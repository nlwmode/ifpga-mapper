module top (ADS_n_pad, \Address[0]_pad , \Address[10]_pad , \Address[11]_pad , \Address[12]_pad , \Address[13]_pad , \Address[14]_pad , \Address[15]_pad , \Address[16]_pad , \Address[17]_pad , \Address[18]_pad , \Address[19]_pad , \Address[1]_pad , \Address[20]_pad , \Address[21]_pad , \Address[22]_pad , \Address[23]_pad , \Address[24]_pad , \Address[25]_pad , \Address[26]_pad , \Address[27]_pad , \Address[28]_pad , \Address[29]_pad , \Address[2]_pad , \Address[3]_pad , \Address[4]_pad , \Address[5]_pad , \Address[6]_pad , \Address[7]_pad , \Address[8]_pad , \Address[9]_pad , \BE_n[0]_pad , \BE_n[1]_pad , \BE_n[2]_pad , \BE_n[3]_pad , \BS16_n_pad , \ByteEnable_reg[0]/NET0131 , \ByteEnable_reg[1]/NET0131 , \ByteEnable_reg[2]/NET0131 , \ByteEnable_reg[3]/NET0131 , \CodeFetch_reg/NET0131 , D_C_n_pad, \DataWidth_reg[0]/NET0131 , \DataWidth_reg[1]/NET0131 , \Datai[0]_pad , \Datai[10]_pad , \Datai[11]_pad , \Datai[12]_pad , \Datai[13]_pad , \Datai[14]_pad , \Datai[15]_pad , \Datai[16]_pad , \Datai[17]_pad , \Datai[18]_pad , \Datai[19]_pad , \Datai[1]_pad , \Datai[20]_pad , \Datai[21]_pad , \Datai[22]_pad , \Datai[23]_pad , \Datai[24]_pad , \Datai[25]_pad , \Datai[26]_pad , \Datai[27]_pad , \Datai[28]_pad , \Datai[29]_pad , \Datai[2]_pad , \Datai[30]_pad , \Datai[31]_pad , \Datai[3]_pad , \Datai[4]_pad , \Datai[5]_pad , \Datai[6]_pad , \Datai[7]_pad , \Datai[8]_pad , \Datai[9]_pad , \Datao[0]_pad , \Datao[10]_pad , \Datao[11]_pad , \Datao[12]_pad , \Datao[13]_pad , \Datao[14]_pad , \Datao[15]_pad , \Datao[16]_pad , \Datao[17]_pad , \Datao[18]_pad , \Datao[19]_pad , \Datao[1]_pad , \Datao[20]_pad , \Datao[21]_pad , \Datao[22]_pad , \Datao[23]_pad , \Datao[24]_pad , \Datao[25]_pad , \Datao[26]_pad , \Datao[27]_pad , \Datao[28]_pad , \Datao[29]_pad , \Datao[2]_pad , \Datao[30]_pad , \Datao[3]_pad , \Datao[4]_pad , \Datao[5]_pad , \Datao[6]_pad , \Datao[7]_pad , \Datao[8]_pad , \Datao[9]_pad , \EAX_reg[0]/NET0131 , \EAX_reg[10]/NET0131 , \EAX_reg[11]/NET0131 , \EAX_reg[12]/NET0131 , \EAX_reg[13]/NET0131 , \EAX_reg[14]/NET0131 , \EAX_reg[15]/NET0131 , \EAX_reg[16]/NET0131 , \EAX_reg[17]/NET0131 , \EAX_reg[18]/NET0131 , \EAX_reg[19]/NET0131 , \EAX_reg[1]/NET0131 , \EAX_reg[20]/NET0131 , \EAX_reg[21]/NET0131 , \EAX_reg[22]/NET0131 , \EAX_reg[23]/NET0131 , \EAX_reg[24]/NET0131 , \EAX_reg[25]/NET0131 , \EAX_reg[26]/NET0131 , \EAX_reg[27]/NET0131 , \EAX_reg[28]/NET0131 , \EAX_reg[29]/NET0131 , \EAX_reg[2]/NET0131 , \EAX_reg[30]/NET0131 , \EAX_reg[31]/NET0131 , \EAX_reg[3]/NET0131 , \EAX_reg[4]/NET0131 , \EAX_reg[5]/NET0131 , \EAX_reg[6]/NET0131 , \EAX_reg[7]/NET0131 , \EAX_reg[8]/NET0131 , \EAX_reg[9]/NET0131 , \EBX_reg[0]/NET0131 , \EBX_reg[10]/NET0131 , \EBX_reg[11]/NET0131 , \EBX_reg[12]/NET0131 , \EBX_reg[13]/NET0131 , \EBX_reg[14]/NET0131 , \EBX_reg[15]/NET0131 , \EBX_reg[16]/NET0131 , \EBX_reg[17]/NET0131 , \EBX_reg[18]/NET0131 , \EBX_reg[19]/NET0131 , \EBX_reg[1]/NET0131 , \EBX_reg[20]/NET0131 , \EBX_reg[21]/NET0131 , \EBX_reg[22]/NET0131 , \EBX_reg[23]/NET0131 , \EBX_reg[24]/NET0131 , \EBX_reg[25]/NET0131 , \EBX_reg[26]/NET0131 , \EBX_reg[27]/NET0131 , \EBX_reg[28]/NET0131 , \EBX_reg[29]/NET0131 , \EBX_reg[2]/NET0131 , \EBX_reg[30]/NET0131 , \EBX_reg[31]/NET0131 , \EBX_reg[3]/NET0131 , \EBX_reg[4]/NET0131 , \EBX_reg[5]/NET0131 , \EBX_reg[6]/NET0131 , \EBX_reg[7]/NET0131 , \EBX_reg[8]/NET0131 , \EBX_reg[9]/NET0131 , \Flush_reg/NET0131 , HOLD_pad, \InstAddrPointer_reg[0]/NET0131 , \InstAddrPointer_reg[10]/NET0131 , \InstAddrPointer_reg[11]/NET0131 , \InstAddrPointer_reg[12]/NET0131 , \InstAddrPointer_reg[13]/NET0131 , \InstAddrPointer_reg[14]/NET0131 , \InstAddrPointer_reg[15]/NET0131 , \InstAddrPointer_reg[16]/NET0131 , \InstAddrPointer_reg[17]/NET0131 , \InstAddrPointer_reg[18]/NET0131 , \InstAddrPointer_reg[19]/NET0131 , \InstAddrPointer_reg[1]/NET0131 , \InstAddrPointer_reg[20]/NET0131 , \InstAddrPointer_reg[21]/NET0131 , \InstAddrPointer_reg[22]/NET0131 , \InstAddrPointer_reg[23]/NET0131 , \InstAddrPointer_reg[24]/NET0131 , \InstAddrPointer_reg[25]/NET0131 , \InstAddrPointer_reg[26]/NET0131 , \InstAddrPointer_reg[27]/NET0131 , \InstAddrPointer_reg[28]/NET0131 , \InstAddrPointer_reg[29]/NET0131 , \InstAddrPointer_reg[2]/NET0131 , \InstAddrPointer_reg[30]/NET0131 , \InstAddrPointer_reg[31]/NET0131 , \InstAddrPointer_reg[3]/NET0131 , \InstAddrPointer_reg[4]/NET0131 , \InstAddrPointer_reg[5]/NET0131 , \InstAddrPointer_reg[6]/NET0131 , \InstAddrPointer_reg[7]/NET0131 , \InstAddrPointer_reg[8]/NET0131 , \InstAddrPointer_reg[9]/NET0131 , \InstQueueRd_Addr_reg[0]/NET0131 , \InstQueueRd_Addr_reg[1]/NET0131 , \InstQueueRd_Addr_reg[2]/NET0131 , \InstQueueRd_Addr_reg[3]/NET0131 , \InstQueueWr_Addr_reg[0]/NET0131 , \InstQueueWr_Addr_reg[1]/NET0131 , \InstQueueWr_Addr_reg[2]/NET0131 , \InstQueueWr_Addr_reg[3]/NET0131 , \InstQueue_reg[0][0]/NET0131 , \InstQueue_reg[0][1]/NET0131 , \InstQueue_reg[0][2]/NET0131 , \InstQueue_reg[0][3]/NET0131 , \InstQueue_reg[0][4]/NET0131 , \InstQueue_reg[0][5]/NET0131 , \InstQueue_reg[0][6]/NET0131 , \InstQueue_reg[0][7]/NET0131 , \InstQueue_reg[10][0]/NET0131 , \InstQueue_reg[10][1]/NET0131 , \InstQueue_reg[10][2]/NET0131 , \InstQueue_reg[10][3]/NET0131 , \InstQueue_reg[10][4]/NET0131 , \InstQueue_reg[10][5]/NET0131 , \InstQueue_reg[10][6]/NET0131 , \InstQueue_reg[10][7]/NET0131 , \InstQueue_reg[11][0]/NET0131 , \InstQueue_reg[11][1]/NET0131 , \InstQueue_reg[11][2]/NET0131 , \InstQueue_reg[11][3]/NET0131 , \InstQueue_reg[11][4]/NET0131 , \InstQueue_reg[11][5]/NET0131 , \InstQueue_reg[11][6]/NET0131 , \InstQueue_reg[11][7]/NET0131 , \InstQueue_reg[12][0]/NET0131 , \InstQueue_reg[12][1]/NET0131 , \InstQueue_reg[12][2]/NET0131 , \InstQueue_reg[12][3]/NET0131 , \InstQueue_reg[12][4]/NET0131 , \InstQueue_reg[12][5]/NET0131 , \InstQueue_reg[12][6]/NET0131 , \InstQueue_reg[12][7]/NET0131 , \InstQueue_reg[13][0]/NET0131 , \InstQueue_reg[13][1]/NET0131 , \InstQueue_reg[13][2]/NET0131 , \InstQueue_reg[13][3]/NET0131 , \InstQueue_reg[13][4]/NET0131 , \InstQueue_reg[13][5]/NET0131 , \InstQueue_reg[13][6]/NET0131 , \InstQueue_reg[13][7]/NET0131 , \InstQueue_reg[14][0]/NET0131 , \InstQueue_reg[14][1]/NET0131 , \InstQueue_reg[14][2]/NET0131 , \InstQueue_reg[14][3]/NET0131 , \InstQueue_reg[14][4]/NET0131 , \InstQueue_reg[14][5]/NET0131 , \InstQueue_reg[14][6]/NET0131 , \InstQueue_reg[14][7]/NET0131 , \InstQueue_reg[15][0]/NET0131 , \InstQueue_reg[15][1]/NET0131 , \InstQueue_reg[15][2]/NET0131 , \InstQueue_reg[15][3]/NET0131 , \InstQueue_reg[15][4]/NET0131 , \InstQueue_reg[15][5]/NET0131 , \InstQueue_reg[15][6]/NET0131 , \InstQueue_reg[15][7]/NET0131 , \InstQueue_reg[1][0]/NET0131 , \InstQueue_reg[1][1]/NET0131 , \InstQueue_reg[1][2]/NET0131 , \InstQueue_reg[1][3]/NET0131 , \InstQueue_reg[1][4]/NET0131 , \InstQueue_reg[1][5]/NET0131 , \InstQueue_reg[1][6]/NET0131 , \InstQueue_reg[1][7]/NET0131 , \InstQueue_reg[2][0]/NET0131 , \InstQueue_reg[2][1]/NET0131 , \InstQueue_reg[2][2]/NET0131 , \InstQueue_reg[2][3]/NET0131 , \InstQueue_reg[2][4]/NET0131 , \InstQueue_reg[2][5]/NET0131 , \InstQueue_reg[2][6]/NET0131 , \InstQueue_reg[2][7]/NET0131 , \InstQueue_reg[3][0]/NET0131 , \InstQueue_reg[3][1]/NET0131 , \InstQueue_reg[3][2]/NET0131 , \InstQueue_reg[3][3]/NET0131 , \InstQueue_reg[3][4]/NET0131 , \InstQueue_reg[3][5]/NET0131 , \InstQueue_reg[3][6]/NET0131 , \InstQueue_reg[3][7]/NET0131 , \InstQueue_reg[4][0]/NET0131 , \InstQueue_reg[4][1]/NET0131 , \InstQueue_reg[4][2]/NET0131 , \InstQueue_reg[4][3]/NET0131 , \InstQueue_reg[4][4]/NET0131 , \InstQueue_reg[4][5]/NET0131 , \InstQueue_reg[4][6]/NET0131 , \InstQueue_reg[4][7]/NET0131 , \InstQueue_reg[5][0]/NET0131 , \InstQueue_reg[5][1]/NET0131 , \InstQueue_reg[5][2]/NET0131 , \InstQueue_reg[5][3]/NET0131 , \InstQueue_reg[5][4]/NET0131 , \InstQueue_reg[5][5]/NET0131 , \InstQueue_reg[5][6]/NET0131 , \InstQueue_reg[5][7]/NET0131 , \InstQueue_reg[6][0]/NET0131 , \InstQueue_reg[6][1]/NET0131 , \InstQueue_reg[6][2]/NET0131 , \InstQueue_reg[6][3]/NET0131 , \InstQueue_reg[6][4]/NET0131 , \InstQueue_reg[6][5]/NET0131 , \InstQueue_reg[6][6]/NET0131 , \InstQueue_reg[6][7]/NET0131 , \InstQueue_reg[7][0]/NET0131 , \InstQueue_reg[7][1]/NET0131 , \InstQueue_reg[7][2]/NET0131 , \InstQueue_reg[7][3]/NET0131 , \InstQueue_reg[7][4]/NET0131 , \InstQueue_reg[7][5]/NET0131 , \InstQueue_reg[7][6]/NET0131 , \InstQueue_reg[7][7]/NET0131 , \InstQueue_reg[8][0]/NET0131 , \InstQueue_reg[8][1]/NET0131 , \InstQueue_reg[8][2]/NET0131 , \InstQueue_reg[8][3]/NET0131 , \InstQueue_reg[8][4]/NET0131 , \InstQueue_reg[8][5]/NET0131 , \InstQueue_reg[8][6]/NET0131 , \InstQueue_reg[8][7]/NET0131 , \InstQueue_reg[9][0]/NET0131 , \InstQueue_reg[9][1]/NET0131 , \InstQueue_reg[9][2]/NET0131 , \InstQueue_reg[9][3]/NET0131 , \InstQueue_reg[9][4]/NET0131 , \InstQueue_reg[9][5]/NET0131 , \InstQueue_reg[9][6]/NET0131 , \InstQueue_reg[9][7]/NET0131 , M_IO_n_pad, \MemoryFetch_reg/NET0131 , \More_reg/NET0131 , NA_n_pad, \PhyAddrPointer_reg[0]/NET0131 , \PhyAddrPointer_reg[10]/NET0131 , \PhyAddrPointer_reg[11]/NET0131 , \PhyAddrPointer_reg[12]/NET0131 , \PhyAddrPointer_reg[13]/NET0131 , \PhyAddrPointer_reg[14]/NET0131 , \PhyAddrPointer_reg[15]/NET0131 , \PhyAddrPointer_reg[16]/NET0131 , \PhyAddrPointer_reg[17]/NET0131 , \PhyAddrPointer_reg[18]/NET0131 , \PhyAddrPointer_reg[19]/NET0131 , \PhyAddrPointer_reg[1]/NET0131 , \PhyAddrPointer_reg[20]/NET0131 , \PhyAddrPointer_reg[21]/NET0131 , \PhyAddrPointer_reg[22]/NET0131 , \PhyAddrPointer_reg[23]/NET0131 , \PhyAddrPointer_reg[24]/NET0131 , \PhyAddrPointer_reg[25]/NET0131 , \PhyAddrPointer_reg[26]/NET0131 , \PhyAddrPointer_reg[27]/NET0131 , \PhyAddrPointer_reg[28]/NET0131 , \PhyAddrPointer_reg[29]/NET0131 , \PhyAddrPointer_reg[2]/NET0131 , \PhyAddrPointer_reg[30]/NET0131 , \PhyAddrPointer_reg[31]/NET0131 , \PhyAddrPointer_reg[3]/NET0131 , \PhyAddrPointer_reg[4]/NET0131 , \PhyAddrPointer_reg[5]/NET0131 , \PhyAddrPointer_reg[6]/NET0131 , \PhyAddrPointer_reg[7]/NET0131 , \PhyAddrPointer_reg[8]/NET0131 , \PhyAddrPointer_reg[9]/NET0131 , READY_n_pad, \ReadRequest_reg/NET0131 , \RequestPending_reg/NET0131 , \State2_reg[0]/NET0131 , \State2_reg[1]/NET0131 , \State2_reg[2]/NET0131 , \State2_reg[3]/NET0131 , \State_reg[0]/NET0131 , \State_reg[1]/NET0131 , \State_reg[2]/NET0131 , W_R_n_pad, \lWord_reg[0]/NET0131 , \lWord_reg[10]/NET0131 , \lWord_reg[11]/NET0131 , \lWord_reg[12]/NET0131 , \lWord_reg[13]/NET0131 , \lWord_reg[14]/NET0131 , \lWord_reg[15]/NET0131 , \lWord_reg[1]/NET0131 , \lWord_reg[2]/NET0131 , \lWord_reg[3]/NET0131 , \lWord_reg[4]/NET0131 , \lWord_reg[5]/NET0131 , \lWord_reg[6]/NET0131 , \lWord_reg[7]/NET0131 , \lWord_reg[8]/NET0131 , \lWord_reg[9]/NET0131 , \rEIP_reg[0]/NET0131 , \rEIP_reg[10]/NET0131 , \rEIP_reg[11]/NET0131 , \rEIP_reg[12]/NET0131 , \rEIP_reg[13]/NET0131 , \rEIP_reg[14]/NET0131 , \rEIP_reg[15]/NET0131 , \rEIP_reg[16]/NET0131 , \rEIP_reg[17]/NET0131 , \rEIP_reg[18]/NET0131 , \rEIP_reg[19]/NET0131 , \rEIP_reg[1]/NET0131 , \rEIP_reg[20]/NET0131 , \rEIP_reg[21]/NET0131 , \rEIP_reg[22]/NET0131 , \rEIP_reg[23]/NET0131 , \rEIP_reg[24]/NET0131 , \rEIP_reg[25]/NET0131 , \rEIP_reg[26]/NET0131 , \rEIP_reg[27]/NET0131 , \rEIP_reg[28]/NET0131 , \rEIP_reg[29]/NET0131 , \rEIP_reg[2]/NET0131 , \rEIP_reg[30]/NET0131 , \rEIP_reg[31]/NET0131 , \rEIP_reg[3]/NET0131 , \rEIP_reg[4]/NET0131 , \rEIP_reg[5]/NET0131 , \rEIP_reg[6]/NET0131 , \rEIP_reg[7]/NET0131 , \rEIP_reg[8]/NET0131 , \rEIP_reg[9]/NET0131 , \uWord_reg[0]/NET0131 , \uWord_reg[10]/NET0131 , \uWord_reg[11]/NET0131 , \uWord_reg[12]/NET0131 , \uWord_reg[13]/NET0131 , \uWord_reg[14]/NET0131 , \uWord_reg[1]/NET0131 , \uWord_reg[2]/NET0131 , \uWord_reg[3]/NET0131 , \uWord_reg[4]/NET0131 , \uWord_reg[5]/NET0131 , \uWord_reg[6]/NET0131 , \uWord_reg[7]/NET0131 , \uWord_reg[8]/NET0131 , \uWord_reg[9]/NET0131 , \_al_n0 , \_al_n1 , \g47406/_2_ , \g47407/_2_ , \g47411/_0_ , \g47413/_0_ , \g47424/_0_ , \g47434/_0_ , \g47437/_0_ , \g47447/_2_ , \g47448/_0_ , \g47451/_0_ , \g47452/_0_ , \g47453/_0_ , \g47465/_2_ , \g47466/_0_ , \g47467/_0_ , \g47471/_0_ , \g47485/_0_ , \g47486/_0_ , \g47487/_2_ , \g47488/_0_ , \g47489/_2_ , \g47491/_0_ , \g47494/_0_ , \g47510/_0_ , \g47511/_0_ , \g47512/_0_ , \g47515/_0_ , \g47516/_0_ , \g47517/_2_ , \g47524/_0_ , \g47525/_0_ , \g47550/_0_ , \g47551/_2_ , \g47552/_0_ , \g47554/_0_ , \g47555/_0_ , \g47556/_0_ , \g47558/_0_ , \g47563/_0_ , \g47564/_0_ , \g47565/_0_ , \g47584/_0_ , \g47592/_0_ , \g47597/_0_ , \g47598/_0_ , \g47601/_0_ , \g47602/_0_ , \g47603/_0_ , \g47604/_0_ , \g47606/_0_ , \g47630/_0_ , \g47636/_0_ , \g47641/_0_ , \g47642/_0_ , \g47643/_0_ , \g47644/_0_ , \g47645/_0_ , \g47646/_0_ , \g47648/_0_ , \g47679/_0_ , \g47680/_0_ , \g47681/_0_ , \g47683/_0_ , \g47687/_0_ , \g47690/_0_ , \g47746/_0_ , \g47747/_0_ , \g47754/_0_ , \g47756/_0_ , \g47804/_0_ , \g47805/_0_ , \g47806/_0_ , \g47807/_0_ , \g47809/_0_ , \g47810/_0_ , \g47812/_0_ , \g47813/_0_ , \g47814/_0_ , \g47815/_0_ , \g47816/_0_ , \g47817/_0_ , \g47818/_0_ , \g47819/_0_ , \g47820/_0_ , \g47821/_0_ , \g47836/_0_ , \g47848/_0_ , \g47851/_0_ , \g47852/_0_ , \g47943/_0_ , \g47944/_0_ , \g47945/_0_ , \g47946/_0_ , \g47947/_0_ , \g47949/_0_ , \g47950/_0_ , \g47952/_0_ , \g47953/_0_ , \g47954/_0_ , \g47955/_0_ , \g47956/_0_ , \g47957/_0_ , \g47958/_0_ , \g47959/_0_ , \g47960/_0_ , \g47999/_0_ , \g48/_0_ , \g48005/_0_ , \g48006/_0_ , \g48007/_0_ , \g48008/_0_ , \g48009/_0_ , \g48010/_0_ , \g48011/_0_ , \g48012/_0_ , \g48013/_0_ , \g48014/_0_ , \g48015/_0_ , \g48057/_0_ , \g48058/_0_ , \g48059/_0_ , \g48060/_0_ , \g48061/_0_ , \g48062/_0_ , \g48063/_0_ , \g48064/_0_ , \g48066/_0_ , \g48067/_0_ , \g48068/_0_ , \g48069/_0_ , \g48070/_0_ , \g48071/_0_ , \g48073/_0_ , \g48074/_0_ , \g48075/_0_ , \g48076/_0_ , \g48077/_0_ , \g48078/_0_ , \g48079/_0_ , \g48080/_0_ , \g48081/_0_ , \g48082/_0_ , \g48084/_0_ , \g48085/_0_ , \g48086/_0_ , \g48087/_0_ , \g48089/_0_ , \g48090/_0_ , \g48091/_0_ , \g48093/_0_ , \g48094/_0_ , \g48119/_0_ , \g48120/_0_ , \g48121/_0_ , \g48122/_0_ , \g48123/_0_ , \g48124/_0_ , \g48125/_0_ , \g48126/_0_ , \g48127/_0_ , \g48128/_0_ , \g48129/_0_ , \g48130/_0_ , \g48131/_0_ , \g48132/_0_ , \g48133/_0_ , \g48134/_0_ , \g48135/_0_ , \g48136/_0_ , \g48137/_0_ , \g48138/_0_ , \g48140/_0_ , \g48144/_0_ , \g48145/_0_ , \g48146/_0_ , \g48147/_0_ , \g48148/_0_ , \g48150/_0_ , \g48151/_0_ , \g48152/_0_ , \g48153/_0_ , \g48154/_0_ , \g48176/_0_ , \g48189/_0_ , \g48192/_0_ , \g48193/_0_ , \g48194/_0_ , \g48195/_0_ , \g48196/_0_ , \g48197/_0_ , \g48198/_0_ , \g48199/_0_ , \g48200/_0_ , \g48263/_0_ , \g48265/_0_ , \g48273/_0_ , \g48313/_0_ , \g48318/_0_ , \g48319/_0_ , \g48321/_0_ , \g48323/_0_ , \g48324/_0_ , \g48325/_0_ , \g48326/_0_ , \g48327/_0_ , \g48328/_0_ , \g48329/_0_ , \g48330/_0_ , \g48331/_0_ , \g48332/_0_ , \g48333/_0_ , \g48472/_0_ , \g48519/_0_ , \g48520/_0_ , \g48521/_0_ , \g48522/_0_ , \g48523/_0_ , \g48524/_0_ , \g48525/_0_ , \g48527/_0_ , \g48529/_0_ , \g48530/_0_ , \g48531/_0_ , \g48532/_0_ , \g48533/_0_ , \g48534/_0_ , \g48535/_0_ , \g48536/_0_ , \g48537/_0_ , \g48538/_0_ , \g48539/_0_ , \g48540/_0_ , \g48541/_0_ , \g48542/_0_ , \g48543/_0_ , \g48545/_0_ , \g48546/_0_ , \g48547/_0_ , \g48639/_0_ , \g48642/_0_ , \g48645/_0_ , \g48648/_0_ , \g48652/_0_ , \g48655/_0_ , \g48658/_0_ , \g48661/_0_ , \g48664/_0_ , \g48667/_0_ , \g48670/_0_ , \g48673/_0_ , \g48678/_0_ , \g48681/_0_ , \g48684/_0_ , \g48688/_0_ , \g48793/_0_ , \g48812/_0_ , \g48813/_0_ , \g48814/_0_ , \g48824/_0_ , \g48825/_0_ , \g48826/_0_ , \g48827/_0_ , \g48828/_0_ , \g48829/_0_ , \g48830/_0_ , \g48831/_0_ , \g48833/_0_ , \g48834/_0_ , \g48835/_0_ , \g48836/_0_ , \g48837/_0_ , \g48838/_0_ , \g48839/_0_ , \g48840/_0_ , \g48841/_0_ , \g48842/_0_ , \g48843/_0_ , \g48844/_0_ , \g48845/_0_ , \g48846/_0_ , \g48847/_0_ , \g48848/_0_ , \g48908/_0_ , \g48909/_0_ , \g48910/_0_ , \g48912/_0_ , \g48913/_0_ , \g48915/_0_ , \g48917/_0_ , \g48932/_0_ , \g48933/_0_ , \g48935/_0_ , \g48937/_0_ , \g48938/_0_ , \g48939/_0_ , \g48940/_0_ , \g48942/_0_ , \g48945/_0_ , \g48971/_0_ , \g49007/_0_ , \g49047/_0_ , \g49048/_0_ , \g49050/_0_ , \g49182/_0_ , \g49280/_0_ , \g49332/_0_ , \g49335/_0_ , \g49336/_0_ , \g49337/_0_ , \g49338/_0_ , \g49339/_0_ , \g49340/_0_ , \g49341/_0_ , \g49342/_0_ , \g49343/_0_ , \g49344/_0_ , \g49345/_0_ , \g49346/_0_ , \g49347/_0_ , \g49348/_0_ , \g49349/_0_ , \g49356/_0_ , \g49375/_0_ , \g49396/_0_ , \g49397/_0_ , \g49400/_0_ , \g49404/_0_ , \g49406/_0_ , \g49414/_0_ , \g49422/_0_ , \g49426/_0_ , \g49430/_0_ , \g49434/_0_ , \g49437/_0_ , \g49440/_0_ , \g49441/_0_ , \g49444/_0_ , \g49448/_0_ , \g49451/_0_ , \g49455/_0_ , \g49456/_0_ , \g49460/_0_ , \g49466/_0_ , \g49563/_0_ , \g49592/_0_ , \g49915/_0_ , \g49941/_0_ , \g50023/_0_ , \g50026/_0_ , \g50029/_0_ , \g50031/_0_ , \g50033/_0_ , \g50035/_0_ , \g50037/_0_ , \g50040/_0_ , \g50050/_0_ , \g50056/_0_ , \g50059/_0_ , \g50065/_0_ , \g50067/_0_ , \g50150/_0_ , \g50283/_0_ , \g50284/_0_ , \g50501/_0_ , \g50594/_0_ , \g50807/_0_ , \g50866/_0_ , \g50875/_0_ , \g51449/_0_ , \g51510/_0_ , \g51534/_0_ , \g52310/_0_ , \g53066/_0_ , \g53087/_0_ , \g53151/_0_ , \g53608/_0_ , \g53634/_0_ , \g54053/_0_ , \g54091/_0_ , \g54103/_0_ , \g54268/_0_ , \g54277/_0_ , \g54287/_0_ , \g54294/_0_ , \g54449/_0_ , \g54453/_0_ , \g54484/_0_ , \g54528/_0_ , \g54582/_0_ , \g55448/_0_ , \g55693/_1_ , \g55874/_0_ , \g56203/_0_ , \g56303/_0_ , \g56329/_0_ , \g56336/_0_ , \g56345/_0_ , \g56367/_0_ , \g56411/_0_ , \g56529/_0_ , \g56858/_0_ , \g60443/_1_ , \g63395/_0_ , \g63442/_0_ , \g63595/_0_ , \g63996/_0_ , \g64048/_0_ , \g64071/_0_ , \g64085/_0_ , \g64096/_0_ , \g64119/_0_ , \g64216/_0_ , \g64513/_0_ , \g64566/_0_ , \g64694/_0_ , \g64913/_0_ );
	input ADS_n_pad ;
	input \Address[0]_pad  ;
	input \Address[10]_pad  ;
	input \Address[11]_pad  ;
	input \Address[12]_pad  ;
	input \Address[13]_pad  ;
	input \Address[14]_pad  ;
	input \Address[15]_pad  ;
	input \Address[16]_pad  ;
	input \Address[17]_pad  ;
	input \Address[18]_pad  ;
	input \Address[19]_pad  ;
	input \Address[1]_pad  ;
	input \Address[20]_pad  ;
	input \Address[21]_pad  ;
	input \Address[22]_pad  ;
	input \Address[23]_pad  ;
	input \Address[24]_pad  ;
	input \Address[25]_pad  ;
	input \Address[26]_pad  ;
	input \Address[27]_pad  ;
	input \Address[28]_pad  ;
	input \Address[29]_pad  ;
	input \Address[2]_pad  ;
	input \Address[3]_pad  ;
	input \Address[4]_pad  ;
	input \Address[5]_pad  ;
	input \Address[6]_pad  ;
	input \Address[7]_pad  ;
	input \Address[8]_pad  ;
	input \Address[9]_pad  ;
	input \BE_n[0]_pad  ;
	input \BE_n[1]_pad  ;
	input \BE_n[2]_pad  ;
	input \BE_n[3]_pad  ;
	input \BS16_n_pad  ;
	input \ByteEnable_reg[0]/NET0131  ;
	input \ByteEnable_reg[1]/NET0131  ;
	input \ByteEnable_reg[2]/NET0131  ;
	input \ByteEnable_reg[3]/NET0131  ;
	input \CodeFetch_reg/NET0131  ;
	input D_C_n_pad ;
	input \DataWidth_reg[0]/NET0131  ;
	input \DataWidth_reg[1]/NET0131  ;
	input \Datai[0]_pad  ;
	input \Datai[10]_pad  ;
	input \Datai[11]_pad  ;
	input \Datai[12]_pad  ;
	input \Datai[13]_pad  ;
	input \Datai[14]_pad  ;
	input \Datai[15]_pad  ;
	input \Datai[16]_pad  ;
	input \Datai[17]_pad  ;
	input \Datai[18]_pad  ;
	input \Datai[19]_pad  ;
	input \Datai[1]_pad  ;
	input \Datai[20]_pad  ;
	input \Datai[21]_pad  ;
	input \Datai[22]_pad  ;
	input \Datai[23]_pad  ;
	input \Datai[24]_pad  ;
	input \Datai[25]_pad  ;
	input \Datai[26]_pad  ;
	input \Datai[27]_pad  ;
	input \Datai[28]_pad  ;
	input \Datai[29]_pad  ;
	input \Datai[2]_pad  ;
	input \Datai[30]_pad  ;
	input \Datai[31]_pad  ;
	input \Datai[3]_pad  ;
	input \Datai[4]_pad  ;
	input \Datai[5]_pad  ;
	input \Datai[6]_pad  ;
	input \Datai[7]_pad  ;
	input \Datai[8]_pad  ;
	input \Datai[9]_pad  ;
	input \Datao[0]_pad  ;
	input \Datao[10]_pad  ;
	input \Datao[11]_pad  ;
	input \Datao[12]_pad  ;
	input \Datao[13]_pad  ;
	input \Datao[14]_pad  ;
	input \Datao[15]_pad  ;
	input \Datao[16]_pad  ;
	input \Datao[17]_pad  ;
	input \Datao[18]_pad  ;
	input \Datao[19]_pad  ;
	input \Datao[1]_pad  ;
	input \Datao[20]_pad  ;
	input \Datao[21]_pad  ;
	input \Datao[22]_pad  ;
	input \Datao[23]_pad  ;
	input \Datao[24]_pad  ;
	input \Datao[25]_pad  ;
	input \Datao[26]_pad  ;
	input \Datao[27]_pad  ;
	input \Datao[28]_pad  ;
	input \Datao[29]_pad  ;
	input \Datao[2]_pad  ;
	input \Datao[30]_pad  ;
	input \Datao[3]_pad  ;
	input \Datao[4]_pad  ;
	input \Datao[5]_pad  ;
	input \Datao[6]_pad  ;
	input \Datao[7]_pad  ;
	input \Datao[8]_pad  ;
	input \Datao[9]_pad  ;
	input \EAX_reg[0]/NET0131  ;
	input \EAX_reg[10]/NET0131  ;
	input \EAX_reg[11]/NET0131  ;
	input \EAX_reg[12]/NET0131  ;
	input \EAX_reg[13]/NET0131  ;
	input \EAX_reg[14]/NET0131  ;
	input \EAX_reg[15]/NET0131  ;
	input \EAX_reg[16]/NET0131  ;
	input \EAX_reg[17]/NET0131  ;
	input \EAX_reg[18]/NET0131  ;
	input \EAX_reg[19]/NET0131  ;
	input \EAX_reg[1]/NET0131  ;
	input \EAX_reg[20]/NET0131  ;
	input \EAX_reg[21]/NET0131  ;
	input \EAX_reg[22]/NET0131  ;
	input \EAX_reg[23]/NET0131  ;
	input \EAX_reg[24]/NET0131  ;
	input \EAX_reg[25]/NET0131  ;
	input \EAX_reg[26]/NET0131  ;
	input \EAX_reg[27]/NET0131  ;
	input \EAX_reg[28]/NET0131  ;
	input \EAX_reg[29]/NET0131  ;
	input \EAX_reg[2]/NET0131  ;
	input \EAX_reg[30]/NET0131  ;
	input \EAX_reg[31]/NET0131  ;
	input \EAX_reg[3]/NET0131  ;
	input \EAX_reg[4]/NET0131  ;
	input \EAX_reg[5]/NET0131  ;
	input \EAX_reg[6]/NET0131  ;
	input \EAX_reg[7]/NET0131  ;
	input \EAX_reg[8]/NET0131  ;
	input \EAX_reg[9]/NET0131  ;
	input \EBX_reg[0]/NET0131  ;
	input \EBX_reg[10]/NET0131  ;
	input \EBX_reg[11]/NET0131  ;
	input \EBX_reg[12]/NET0131  ;
	input \EBX_reg[13]/NET0131  ;
	input \EBX_reg[14]/NET0131  ;
	input \EBX_reg[15]/NET0131  ;
	input \EBX_reg[16]/NET0131  ;
	input \EBX_reg[17]/NET0131  ;
	input \EBX_reg[18]/NET0131  ;
	input \EBX_reg[19]/NET0131  ;
	input \EBX_reg[1]/NET0131  ;
	input \EBX_reg[20]/NET0131  ;
	input \EBX_reg[21]/NET0131  ;
	input \EBX_reg[22]/NET0131  ;
	input \EBX_reg[23]/NET0131  ;
	input \EBX_reg[24]/NET0131  ;
	input \EBX_reg[25]/NET0131  ;
	input \EBX_reg[26]/NET0131  ;
	input \EBX_reg[27]/NET0131  ;
	input \EBX_reg[28]/NET0131  ;
	input \EBX_reg[29]/NET0131  ;
	input \EBX_reg[2]/NET0131  ;
	input \EBX_reg[30]/NET0131  ;
	input \EBX_reg[31]/NET0131  ;
	input \EBX_reg[3]/NET0131  ;
	input \EBX_reg[4]/NET0131  ;
	input \EBX_reg[5]/NET0131  ;
	input \EBX_reg[6]/NET0131  ;
	input \EBX_reg[7]/NET0131  ;
	input \EBX_reg[8]/NET0131  ;
	input \EBX_reg[9]/NET0131  ;
	input \Flush_reg/NET0131  ;
	input HOLD_pad ;
	input \InstAddrPointer_reg[0]/NET0131  ;
	input \InstAddrPointer_reg[10]/NET0131  ;
	input \InstAddrPointer_reg[11]/NET0131  ;
	input \InstAddrPointer_reg[12]/NET0131  ;
	input \InstAddrPointer_reg[13]/NET0131  ;
	input \InstAddrPointer_reg[14]/NET0131  ;
	input \InstAddrPointer_reg[15]/NET0131  ;
	input \InstAddrPointer_reg[16]/NET0131  ;
	input \InstAddrPointer_reg[17]/NET0131  ;
	input \InstAddrPointer_reg[18]/NET0131  ;
	input \InstAddrPointer_reg[19]/NET0131  ;
	input \InstAddrPointer_reg[1]/NET0131  ;
	input \InstAddrPointer_reg[20]/NET0131  ;
	input \InstAddrPointer_reg[21]/NET0131  ;
	input \InstAddrPointer_reg[22]/NET0131  ;
	input \InstAddrPointer_reg[23]/NET0131  ;
	input \InstAddrPointer_reg[24]/NET0131  ;
	input \InstAddrPointer_reg[25]/NET0131  ;
	input \InstAddrPointer_reg[26]/NET0131  ;
	input \InstAddrPointer_reg[27]/NET0131  ;
	input \InstAddrPointer_reg[28]/NET0131  ;
	input \InstAddrPointer_reg[29]/NET0131  ;
	input \InstAddrPointer_reg[2]/NET0131  ;
	input \InstAddrPointer_reg[30]/NET0131  ;
	input \InstAddrPointer_reg[31]/NET0131  ;
	input \InstAddrPointer_reg[3]/NET0131  ;
	input \InstAddrPointer_reg[4]/NET0131  ;
	input \InstAddrPointer_reg[5]/NET0131  ;
	input \InstAddrPointer_reg[6]/NET0131  ;
	input \InstAddrPointer_reg[7]/NET0131  ;
	input \InstAddrPointer_reg[8]/NET0131  ;
	input \InstAddrPointer_reg[9]/NET0131  ;
	input \InstQueueRd_Addr_reg[0]/NET0131  ;
	input \InstQueueRd_Addr_reg[1]/NET0131  ;
	input \InstQueueRd_Addr_reg[2]/NET0131  ;
	input \InstQueueRd_Addr_reg[3]/NET0131  ;
	input \InstQueueWr_Addr_reg[0]/NET0131  ;
	input \InstQueueWr_Addr_reg[1]/NET0131  ;
	input \InstQueueWr_Addr_reg[2]/NET0131  ;
	input \InstQueueWr_Addr_reg[3]/NET0131  ;
	input \InstQueue_reg[0][0]/NET0131  ;
	input \InstQueue_reg[0][1]/NET0131  ;
	input \InstQueue_reg[0][2]/NET0131  ;
	input \InstQueue_reg[0][3]/NET0131  ;
	input \InstQueue_reg[0][4]/NET0131  ;
	input \InstQueue_reg[0][5]/NET0131  ;
	input \InstQueue_reg[0][6]/NET0131  ;
	input \InstQueue_reg[0][7]/NET0131  ;
	input \InstQueue_reg[10][0]/NET0131  ;
	input \InstQueue_reg[10][1]/NET0131  ;
	input \InstQueue_reg[10][2]/NET0131  ;
	input \InstQueue_reg[10][3]/NET0131  ;
	input \InstQueue_reg[10][4]/NET0131  ;
	input \InstQueue_reg[10][5]/NET0131  ;
	input \InstQueue_reg[10][6]/NET0131  ;
	input \InstQueue_reg[10][7]/NET0131  ;
	input \InstQueue_reg[11][0]/NET0131  ;
	input \InstQueue_reg[11][1]/NET0131  ;
	input \InstQueue_reg[11][2]/NET0131  ;
	input \InstQueue_reg[11][3]/NET0131  ;
	input \InstQueue_reg[11][4]/NET0131  ;
	input \InstQueue_reg[11][5]/NET0131  ;
	input \InstQueue_reg[11][6]/NET0131  ;
	input \InstQueue_reg[11][7]/NET0131  ;
	input \InstQueue_reg[12][0]/NET0131  ;
	input \InstQueue_reg[12][1]/NET0131  ;
	input \InstQueue_reg[12][2]/NET0131  ;
	input \InstQueue_reg[12][3]/NET0131  ;
	input \InstQueue_reg[12][4]/NET0131  ;
	input \InstQueue_reg[12][5]/NET0131  ;
	input \InstQueue_reg[12][6]/NET0131  ;
	input \InstQueue_reg[12][7]/NET0131  ;
	input \InstQueue_reg[13][0]/NET0131  ;
	input \InstQueue_reg[13][1]/NET0131  ;
	input \InstQueue_reg[13][2]/NET0131  ;
	input \InstQueue_reg[13][3]/NET0131  ;
	input \InstQueue_reg[13][4]/NET0131  ;
	input \InstQueue_reg[13][5]/NET0131  ;
	input \InstQueue_reg[13][6]/NET0131  ;
	input \InstQueue_reg[13][7]/NET0131  ;
	input \InstQueue_reg[14][0]/NET0131  ;
	input \InstQueue_reg[14][1]/NET0131  ;
	input \InstQueue_reg[14][2]/NET0131  ;
	input \InstQueue_reg[14][3]/NET0131  ;
	input \InstQueue_reg[14][4]/NET0131  ;
	input \InstQueue_reg[14][5]/NET0131  ;
	input \InstQueue_reg[14][6]/NET0131  ;
	input \InstQueue_reg[14][7]/NET0131  ;
	input \InstQueue_reg[15][0]/NET0131  ;
	input \InstQueue_reg[15][1]/NET0131  ;
	input \InstQueue_reg[15][2]/NET0131  ;
	input \InstQueue_reg[15][3]/NET0131  ;
	input \InstQueue_reg[15][4]/NET0131  ;
	input \InstQueue_reg[15][5]/NET0131  ;
	input \InstQueue_reg[15][6]/NET0131  ;
	input \InstQueue_reg[15][7]/NET0131  ;
	input \InstQueue_reg[1][0]/NET0131  ;
	input \InstQueue_reg[1][1]/NET0131  ;
	input \InstQueue_reg[1][2]/NET0131  ;
	input \InstQueue_reg[1][3]/NET0131  ;
	input \InstQueue_reg[1][4]/NET0131  ;
	input \InstQueue_reg[1][5]/NET0131  ;
	input \InstQueue_reg[1][6]/NET0131  ;
	input \InstQueue_reg[1][7]/NET0131  ;
	input \InstQueue_reg[2][0]/NET0131  ;
	input \InstQueue_reg[2][1]/NET0131  ;
	input \InstQueue_reg[2][2]/NET0131  ;
	input \InstQueue_reg[2][3]/NET0131  ;
	input \InstQueue_reg[2][4]/NET0131  ;
	input \InstQueue_reg[2][5]/NET0131  ;
	input \InstQueue_reg[2][6]/NET0131  ;
	input \InstQueue_reg[2][7]/NET0131  ;
	input \InstQueue_reg[3][0]/NET0131  ;
	input \InstQueue_reg[3][1]/NET0131  ;
	input \InstQueue_reg[3][2]/NET0131  ;
	input \InstQueue_reg[3][3]/NET0131  ;
	input \InstQueue_reg[3][4]/NET0131  ;
	input \InstQueue_reg[3][5]/NET0131  ;
	input \InstQueue_reg[3][6]/NET0131  ;
	input \InstQueue_reg[3][7]/NET0131  ;
	input \InstQueue_reg[4][0]/NET0131  ;
	input \InstQueue_reg[4][1]/NET0131  ;
	input \InstQueue_reg[4][2]/NET0131  ;
	input \InstQueue_reg[4][3]/NET0131  ;
	input \InstQueue_reg[4][4]/NET0131  ;
	input \InstQueue_reg[4][5]/NET0131  ;
	input \InstQueue_reg[4][6]/NET0131  ;
	input \InstQueue_reg[4][7]/NET0131  ;
	input \InstQueue_reg[5][0]/NET0131  ;
	input \InstQueue_reg[5][1]/NET0131  ;
	input \InstQueue_reg[5][2]/NET0131  ;
	input \InstQueue_reg[5][3]/NET0131  ;
	input \InstQueue_reg[5][4]/NET0131  ;
	input \InstQueue_reg[5][5]/NET0131  ;
	input \InstQueue_reg[5][6]/NET0131  ;
	input \InstQueue_reg[5][7]/NET0131  ;
	input \InstQueue_reg[6][0]/NET0131  ;
	input \InstQueue_reg[6][1]/NET0131  ;
	input \InstQueue_reg[6][2]/NET0131  ;
	input \InstQueue_reg[6][3]/NET0131  ;
	input \InstQueue_reg[6][4]/NET0131  ;
	input \InstQueue_reg[6][5]/NET0131  ;
	input \InstQueue_reg[6][6]/NET0131  ;
	input \InstQueue_reg[6][7]/NET0131  ;
	input \InstQueue_reg[7][0]/NET0131  ;
	input \InstQueue_reg[7][1]/NET0131  ;
	input \InstQueue_reg[7][2]/NET0131  ;
	input \InstQueue_reg[7][3]/NET0131  ;
	input \InstQueue_reg[7][4]/NET0131  ;
	input \InstQueue_reg[7][5]/NET0131  ;
	input \InstQueue_reg[7][6]/NET0131  ;
	input \InstQueue_reg[7][7]/NET0131  ;
	input \InstQueue_reg[8][0]/NET0131  ;
	input \InstQueue_reg[8][1]/NET0131  ;
	input \InstQueue_reg[8][2]/NET0131  ;
	input \InstQueue_reg[8][3]/NET0131  ;
	input \InstQueue_reg[8][4]/NET0131  ;
	input \InstQueue_reg[8][5]/NET0131  ;
	input \InstQueue_reg[8][6]/NET0131  ;
	input \InstQueue_reg[8][7]/NET0131  ;
	input \InstQueue_reg[9][0]/NET0131  ;
	input \InstQueue_reg[9][1]/NET0131  ;
	input \InstQueue_reg[9][2]/NET0131  ;
	input \InstQueue_reg[9][3]/NET0131  ;
	input \InstQueue_reg[9][4]/NET0131  ;
	input \InstQueue_reg[9][5]/NET0131  ;
	input \InstQueue_reg[9][6]/NET0131  ;
	input \InstQueue_reg[9][7]/NET0131  ;
	input M_IO_n_pad ;
	input \MemoryFetch_reg/NET0131  ;
	input \More_reg/NET0131  ;
	input NA_n_pad ;
	input \PhyAddrPointer_reg[0]/NET0131  ;
	input \PhyAddrPointer_reg[10]/NET0131  ;
	input \PhyAddrPointer_reg[11]/NET0131  ;
	input \PhyAddrPointer_reg[12]/NET0131  ;
	input \PhyAddrPointer_reg[13]/NET0131  ;
	input \PhyAddrPointer_reg[14]/NET0131  ;
	input \PhyAddrPointer_reg[15]/NET0131  ;
	input \PhyAddrPointer_reg[16]/NET0131  ;
	input \PhyAddrPointer_reg[17]/NET0131  ;
	input \PhyAddrPointer_reg[18]/NET0131  ;
	input \PhyAddrPointer_reg[19]/NET0131  ;
	input \PhyAddrPointer_reg[1]/NET0131  ;
	input \PhyAddrPointer_reg[20]/NET0131  ;
	input \PhyAddrPointer_reg[21]/NET0131  ;
	input \PhyAddrPointer_reg[22]/NET0131  ;
	input \PhyAddrPointer_reg[23]/NET0131  ;
	input \PhyAddrPointer_reg[24]/NET0131  ;
	input \PhyAddrPointer_reg[25]/NET0131  ;
	input \PhyAddrPointer_reg[26]/NET0131  ;
	input \PhyAddrPointer_reg[27]/NET0131  ;
	input \PhyAddrPointer_reg[28]/NET0131  ;
	input \PhyAddrPointer_reg[29]/NET0131  ;
	input \PhyAddrPointer_reg[2]/NET0131  ;
	input \PhyAddrPointer_reg[30]/NET0131  ;
	input \PhyAddrPointer_reg[31]/NET0131  ;
	input \PhyAddrPointer_reg[3]/NET0131  ;
	input \PhyAddrPointer_reg[4]/NET0131  ;
	input \PhyAddrPointer_reg[5]/NET0131  ;
	input \PhyAddrPointer_reg[6]/NET0131  ;
	input \PhyAddrPointer_reg[7]/NET0131  ;
	input \PhyAddrPointer_reg[8]/NET0131  ;
	input \PhyAddrPointer_reg[9]/NET0131  ;
	input READY_n_pad ;
	input \ReadRequest_reg/NET0131  ;
	input \RequestPending_reg/NET0131  ;
	input \State2_reg[0]/NET0131  ;
	input \State2_reg[1]/NET0131  ;
	input \State2_reg[2]/NET0131  ;
	input \State2_reg[3]/NET0131  ;
	input \State_reg[0]/NET0131  ;
	input \State_reg[1]/NET0131  ;
	input \State_reg[2]/NET0131  ;
	input W_R_n_pad ;
	input \lWord_reg[0]/NET0131  ;
	input \lWord_reg[10]/NET0131  ;
	input \lWord_reg[11]/NET0131  ;
	input \lWord_reg[12]/NET0131  ;
	input \lWord_reg[13]/NET0131  ;
	input \lWord_reg[14]/NET0131  ;
	input \lWord_reg[15]/NET0131  ;
	input \lWord_reg[1]/NET0131  ;
	input \lWord_reg[2]/NET0131  ;
	input \lWord_reg[3]/NET0131  ;
	input \lWord_reg[4]/NET0131  ;
	input \lWord_reg[5]/NET0131  ;
	input \lWord_reg[6]/NET0131  ;
	input \lWord_reg[7]/NET0131  ;
	input \lWord_reg[8]/NET0131  ;
	input \lWord_reg[9]/NET0131  ;
	input \rEIP_reg[0]/NET0131  ;
	input \rEIP_reg[10]/NET0131  ;
	input \rEIP_reg[11]/NET0131  ;
	input \rEIP_reg[12]/NET0131  ;
	input \rEIP_reg[13]/NET0131  ;
	input \rEIP_reg[14]/NET0131  ;
	input \rEIP_reg[15]/NET0131  ;
	input \rEIP_reg[16]/NET0131  ;
	input \rEIP_reg[17]/NET0131  ;
	input \rEIP_reg[18]/NET0131  ;
	input \rEIP_reg[19]/NET0131  ;
	input \rEIP_reg[1]/NET0131  ;
	input \rEIP_reg[20]/NET0131  ;
	input \rEIP_reg[21]/NET0131  ;
	input \rEIP_reg[22]/NET0131  ;
	input \rEIP_reg[23]/NET0131  ;
	input \rEIP_reg[24]/NET0131  ;
	input \rEIP_reg[25]/NET0131  ;
	input \rEIP_reg[26]/NET0131  ;
	input \rEIP_reg[27]/NET0131  ;
	input \rEIP_reg[28]/NET0131  ;
	input \rEIP_reg[29]/NET0131  ;
	input \rEIP_reg[2]/NET0131  ;
	input \rEIP_reg[30]/NET0131  ;
	input \rEIP_reg[31]/NET0131  ;
	input \rEIP_reg[3]/NET0131  ;
	input \rEIP_reg[4]/NET0131  ;
	input \rEIP_reg[5]/NET0131  ;
	input \rEIP_reg[6]/NET0131  ;
	input \rEIP_reg[7]/NET0131  ;
	input \rEIP_reg[8]/NET0131  ;
	input \rEIP_reg[9]/NET0131  ;
	input \uWord_reg[0]/NET0131  ;
	input \uWord_reg[10]/NET0131  ;
	input \uWord_reg[11]/NET0131  ;
	input \uWord_reg[12]/NET0131  ;
	input \uWord_reg[13]/NET0131  ;
	input \uWord_reg[14]/NET0131  ;
	input \uWord_reg[1]/NET0131  ;
	input \uWord_reg[2]/NET0131  ;
	input \uWord_reg[3]/NET0131  ;
	input \uWord_reg[4]/NET0131  ;
	input \uWord_reg[5]/NET0131  ;
	input \uWord_reg[6]/NET0131  ;
	input \uWord_reg[7]/NET0131  ;
	input \uWord_reg[8]/NET0131  ;
	input \uWord_reg[9]/NET0131  ;
	output \_al_n0  ;
	output \_al_n1  ;
	output \g47406/_2_  ;
	output \g47407/_2_  ;
	output \g47411/_0_  ;
	output \g47413/_0_  ;
	output \g47424/_0_  ;
	output \g47434/_0_  ;
	output \g47437/_0_  ;
	output \g47447/_2_  ;
	output \g47448/_0_  ;
	output \g47451/_0_  ;
	output \g47452/_0_  ;
	output \g47453/_0_  ;
	output \g47465/_2_  ;
	output \g47466/_0_  ;
	output \g47467/_0_  ;
	output \g47471/_0_  ;
	output \g47485/_0_  ;
	output \g47486/_0_  ;
	output \g47487/_2_  ;
	output \g47488/_0_  ;
	output \g47489/_2_  ;
	output \g47491/_0_  ;
	output \g47494/_0_  ;
	output \g47510/_0_  ;
	output \g47511/_0_  ;
	output \g47512/_0_  ;
	output \g47515/_0_  ;
	output \g47516/_0_  ;
	output \g47517/_2_  ;
	output \g47524/_0_  ;
	output \g47525/_0_  ;
	output \g47550/_0_  ;
	output \g47551/_2_  ;
	output \g47552/_0_  ;
	output \g47554/_0_  ;
	output \g47555/_0_  ;
	output \g47556/_0_  ;
	output \g47558/_0_  ;
	output \g47563/_0_  ;
	output \g47564/_0_  ;
	output \g47565/_0_  ;
	output \g47584/_0_  ;
	output \g47592/_0_  ;
	output \g47597/_0_  ;
	output \g47598/_0_  ;
	output \g47601/_0_  ;
	output \g47602/_0_  ;
	output \g47603/_0_  ;
	output \g47604/_0_  ;
	output \g47606/_0_  ;
	output \g47630/_0_  ;
	output \g47636/_0_  ;
	output \g47641/_0_  ;
	output \g47642/_0_  ;
	output \g47643/_0_  ;
	output \g47644/_0_  ;
	output \g47645/_0_  ;
	output \g47646/_0_  ;
	output \g47648/_0_  ;
	output \g47679/_0_  ;
	output \g47680/_0_  ;
	output \g47681/_0_  ;
	output \g47683/_0_  ;
	output \g47687/_0_  ;
	output \g47690/_0_  ;
	output \g47746/_0_  ;
	output \g47747/_0_  ;
	output \g47754/_0_  ;
	output \g47756/_0_  ;
	output \g47804/_0_  ;
	output \g47805/_0_  ;
	output \g47806/_0_  ;
	output \g47807/_0_  ;
	output \g47809/_0_  ;
	output \g47810/_0_  ;
	output \g47812/_0_  ;
	output \g47813/_0_  ;
	output \g47814/_0_  ;
	output \g47815/_0_  ;
	output \g47816/_0_  ;
	output \g47817/_0_  ;
	output \g47818/_0_  ;
	output \g47819/_0_  ;
	output \g47820/_0_  ;
	output \g47821/_0_  ;
	output \g47836/_0_  ;
	output \g47848/_0_  ;
	output \g47851/_0_  ;
	output \g47852/_0_  ;
	output \g47943/_0_  ;
	output \g47944/_0_  ;
	output \g47945/_0_  ;
	output \g47946/_0_  ;
	output \g47947/_0_  ;
	output \g47949/_0_  ;
	output \g47950/_0_  ;
	output \g47952/_0_  ;
	output \g47953/_0_  ;
	output \g47954/_0_  ;
	output \g47955/_0_  ;
	output \g47956/_0_  ;
	output \g47957/_0_  ;
	output \g47958/_0_  ;
	output \g47959/_0_  ;
	output \g47960/_0_  ;
	output \g47999/_0_  ;
	output \g48/_0_  ;
	output \g48005/_0_  ;
	output \g48006/_0_  ;
	output \g48007/_0_  ;
	output \g48008/_0_  ;
	output \g48009/_0_  ;
	output \g48010/_0_  ;
	output \g48011/_0_  ;
	output \g48012/_0_  ;
	output \g48013/_0_  ;
	output \g48014/_0_  ;
	output \g48015/_0_  ;
	output \g48057/_0_  ;
	output \g48058/_0_  ;
	output \g48059/_0_  ;
	output \g48060/_0_  ;
	output \g48061/_0_  ;
	output \g48062/_0_  ;
	output \g48063/_0_  ;
	output \g48064/_0_  ;
	output \g48066/_0_  ;
	output \g48067/_0_  ;
	output \g48068/_0_  ;
	output \g48069/_0_  ;
	output \g48070/_0_  ;
	output \g48071/_0_  ;
	output \g48073/_0_  ;
	output \g48074/_0_  ;
	output \g48075/_0_  ;
	output \g48076/_0_  ;
	output \g48077/_0_  ;
	output \g48078/_0_  ;
	output \g48079/_0_  ;
	output \g48080/_0_  ;
	output \g48081/_0_  ;
	output \g48082/_0_  ;
	output \g48084/_0_  ;
	output \g48085/_0_  ;
	output \g48086/_0_  ;
	output \g48087/_0_  ;
	output \g48089/_0_  ;
	output \g48090/_0_  ;
	output \g48091/_0_  ;
	output \g48093/_0_  ;
	output \g48094/_0_  ;
	output \g48119/_0_  ;
	output \g48120/_0_  ;
	output \g48121/_0_  ;
	output \g48122/_0_  ;
	output \g48123/_0_  ;
	output \g48124/_0_  ;
	output \g48125/_0_  ;
	output \g48126/_0_  ;
	output \g48127/_0_  ;
	output \g48128/_0_  ;
	output \g48129/_0_  ;
	output \g48130/_0_  ;
	output \g48131/_0_  ;
	output \g48132/_0_  ;
	output \g48133/_0_  ;
	output \g48134/_0_  ;
	output \g48135/_0_  ;
	output \g48136/_0_  ;
	output \g48137/_0_  ;
	output \g48138/_0_  ;
	output \g48140/_0_  ;
	output \g48144/_0_  ;
	output \g48145/_0_  ;
	output \g48146/_0_  ;
	output \g48147/_0_  ;
	output \g48148/_0_  ;
	output \g48150/_0_  ;
	output \g48151/_0_  ;
	output \g48152/_0_  ;
	output \g48153/_0_  ;
	output \g48154/_0_  ;
	output \g48176/_0_  ;
	output \g48189/_0_  ;
	output \g48192/_0_  ;
	output \g48193/_0_  ;
	output \g48194/_0_  ;
	output \g48195/_0_  ;
	output \g48196/_0_  ;
	output \g48197/_0_  ;
	output \g48198/_0_  ;
	output \g48199/_0_  ;
	output \g48200/_0_  ;
	output \g48263/_0_  ;
	output \g48265/_0_  ;
	output \g48273/_0_  ;
	output \g48313/_0_  ;
	output \g48318/_0_  ;
	output \g48319/_0_  ;
	output \g48321/_0_  ;
	output \g48323/_0_  ;
	output \g48324/_0_  ;
	output \g48325/_0_  ;
	output \g48326/_0_  ;
	output \g48327/_0_  ;
	output \g48328/_0_  ;
	output \g48329/_0_  ;
	output \g48330/_0_  ;
	output \g48331/_0_  ;
	output \g48332/_0_  ;
	output \g48333/_0_  ;
	output \g48472/_0_  ;
	output \g48519/_0_  ;
	output \g48520/_0_  ;
	output \g48521/_0_  ;
	output \g48522/_0_  ;
	output \g48523/_0_  ;
	output \g48524/_0_  ;
	output \g48525/_0_  ;
	output \g48527/_0_  ;
	output \g48529/_0_  ;
	output \g48530/_0_  ;
	output \g48531/_0_  ;
	output \g48532/_0_  ;
	output \g48533/_0_  ;
	output \g48534/_0_  ;
	output \g48535/_0_  ;
	output \g48536/_0_  ;
	output \g48537/_0_  ;
	output \g48538/_0_  ;
	output \g48539/_0_  ;
	output \g48540/_0_  ;
	output \g48541/_0_  ;
	output \g48542/_0_  ;
	output \g48543/_0_  ;
	output \g48545/_0_  ;
	output \g48546/_0_  ;
	output \g48547/_0_  ;
	output \g48639/_0_  ;
	output \g48642/_0_  ;
	output \g48645/_0_  ;
	output \g48648/_0_  ;
	output \g48652/_0_  ;
	output \g48655/_0_  ;
	output \g48658/_0_  ;
	output \g48661/_0_  ;
	output \g48664/_0_  ;
	output \g48667/_0_  ;
	output \g48670/_0_  ;
	output \g48673/_0_  ;
	output \g48678/_0_  ;
	output \g48681/_0_  ;
	output \g48684/_0_  ;
	output \g48688/_0_  ;
	output \g48793/_0_  ;
	output \g48812/_0_  ;
	output \g48813/_0_  ;
	output \g48814/_0_  ;
	output \g48824/_0_  ;
	output \g48825/_0_  ;
	output \g48826/_0_  ;
	output \g48827/_0_  ;
	output \g48828/_0_  ;
	output \g48829/_0_  ;
	output \g48830/_0_  ;
	output \g48831/_0_  ;
	output \g48833/_0_  ;
	output \g48834/_0_  ;
	output \g48835/_0_  ;
	output \g48836/_0_  ;
	output \g48837/_0_  ;
	output \g48838/_0_  ;
	output \g48839/_0_  ;
	output \g48840/_0_  ;
	output \g48841/_0_  ;
	output \g48842/_0_  ;
	output \g48843/_0_  ;
	output \g48844/_0_  ;
	output \g48845/_0_  ;
	output \g48846/_0_  ;
	output \g48847/_0_  ;
	output \g48848/_0_  ;
	output \g48908/_0_  ;
	output \g48909/_0_  ;
	output \g48910/_0_  ;
	output \g48912/_0_  ;
	output \g48913/_0_  ;
	output \g48915/_0_  ;
	output \g48917/_0_  ;
	output \g48932/_0_  ;
	output \g48933/_0_  ;
	output \g48935/_0_  ;
	output \g48937/_0_  ;
	output \g48938/_0_  ;
	output \g48939/_0_  ;
	output \g48940/_0_  ;
	output \g48942/_0_  ;
	output \g48945/_0_  ;
	output \g48971/_0_  ;
	output \g49007/_0_  ;
	output \g49047/_0_  ;
	output \g49048/_0_  ;
	output \g49050/_0_  ;
	output \g49182/_0_  ;
	output \g49280/_0_  ;
	output \g49332/_0_  ;
	output \g49335/_0_  ;
	output \g49336/_0_  ;
	output \g49337/_0_  ;
	output \g49338/_0_  ;
	output \g49339/_0_  ;
	output \g49340/_0_  ;
	output \g49341/_0_  ;
	output \g49342/_0_  ;
	output \g49343/_0_  ;
	output \g49344/_0_  ;
	output \g49345/_0_  ;
	output \g49346/_0_  ;
	output \g49347/_0_  ;
	output \g49348/_0_  ;
	output \g49349/_0_  ;
	output \g49356/_0_  ;
	output \g49375/_0_  ;
	output \g49396/_0_  ;
	output \g49397/_0_  ;
	output \g49400/_0_  ;
	output \g49404/_0_  ;
	output \g49406/_0_  ;
	output \g49414/_0_  ;
	output \g49422/_0_  ;
	output \g49426/_0_  ;
	output \g49430/_0_  ;
	output \g49434/_0_  ;
	output \g49437/_0_  ;
	output \g49440/_0_  ;
	output \g49441/_0_  ;
	output \g49444/_0_  ;
	output \g49448/_0_  ;
	output \g49451/_0_  ;
	output \g49455/_0_  ;
	output \g49456/_0_  ;
	output \g49460/_0_  ;
	output \g49466/_0_  ;
	output \g49563/_0_  ;
	output \g49592/_0_  ;
	output \g49915/_0_  ;
	output \g49941/_0_  ;
	output \g50023/_0_  ;
	output \g50026/_0_  ;
	output \g50029/_0_  ;
	output \g50031/_0_  ;
	output \g50033/_0_  ;
	output \g50035/_0_  ;
	output \g50037/_0_  ;
	output \g50040/_0_  ;
	output \g50050/_0_  ;
	output \g50056/_0_  ;
	output \g50059/_0_  ;
	output \g50065/_0_  ;
	output \g50067/_0_  ;
	output \g50150/_0_  ;
	output \g50283/_0_  ;
	output \g50284/_0_  ;
	output \g50501/_0_  ;
	output \g50594/_0_  ;
	output \g50807/_0_  ;
	output \g50866/_0_  ;
	output \g50875/_0_  ;
	output \g51449/_0_  ;
	output \g51510/_0_  ;
	output \g51534/_0_  ;
	output \g52310/_0_  ;
	output \g53066/_0_  ;
	output \g53087/_0_  ;
	output \g53151/_0_  ;
	output \g53608/_0_  ;
	output \g53634/_0_  ;
	output \g54053/_0_  ;
	output \g54091/_0_  ;
	output \g54103/_0_  ;
	output \g54268/_0_  ;
	output \g54277/_0_  ;
	output \g54287/_0_  ;
	output \g54294/_0_  ;
	output \g54449/_0_  ;
	output \g54453/_0_  ;
	output \g54484/_0_  ;
	output \g54528/_0_  ;
	output \g54582/_0_  ;
	output \g55448/_0_  ;
	output \g55693/_1_  ;
	output \g55874/_0_  ;
	output \g56203/_0_  ;
	output \g56303/_0_  ;
	output \g56329/_0_  ;
	output \g56336/_0_  ;
	output \g56345/_0_  ;
	output \g56367/_0_  ;
	output \g56411/_0_  ;
	output \g56529/_0_  ;
	output \g56858/_0_  ;
	output \g60443/_1_  ;
	output \g63395/_0_  ;
	output \g63442/_0_  ;
	output \g63595/_0_  ;
	output \g63996/_0_  ;
	output \g64048/_0_  ;
	output \g64071/_0_  ;
	output \g64085/_0_  ;
	output \g64096/_0_  ;
	output \g64119/_0_  ;
	output \g64216/_0_  ;
	output \g64513/_0_  ;
	output \g64566/_0_  ;
	output \g64694/_0_  ;
	output \g64913/_0_  ;
	wire _w5492_ ;
	wire _w5491_ ;
	wire _w5490_ ;
	wire _w5489_ ;
	wire _w5488_ ;
	wire _w5487_ ;
	wire _w5486_ ;
	wire _w5485_ ;
	wire _w5484_ ;
	wire _w5483_ ;
	wire _w5482_ ;
	wire _w5481_ ;
	wire _w5480_ ;
	wire _w5479_ ;
	wire _w5478_ ;
	wire _w5477_ ;
	wire _w5476_ ;
	wire _w5475_ ;
	wire _w5474_ ;
	wire _w5473_ ;
	wire _w5472_ ;
	wire _w5471_ ;
	wire _w5470_ ;
	wire _w5469_ ;
	wire _w5468_ ;
	wire _w5467_ ;
	wire _w5466_ ;
	wire _w5465_ ;
	wire _w5464_ ;
	wire _w5463_ ;
	wire _w5462_ ;
	wire _w5461_ ;
	wire _w5460_ ;
	wire _w5459_ ;
	wire _w5458_ ;
	wire _w5457_ ;
	wire _w5456_ ;
	wire _w5455_ ;
	wire _w5454_ ;
	wire _w5453_ ;
	wire _w5452_ ;
	wire _w5451_ ;
	wire _w5450_ ;
	wire _w5449_ ;
	wire _w5448_ ;
	wire _w5447_ ;
	wire _w5446_ ;
	wire _w5445_ ;
	wire _w5444_ ;
	wire _w5443_ ;
	wire _w5442_ ;
	wire _w5441_ ;
	wire _w5440_ ;
	wire _w5439_ ;
	wire _w5438_ ;
	wire _w5437_ ;
	wire _w5436_ ;
	wire _w5435_ ;
	wire _w5434_ ;
	wire _w5433_ ;
	wire _w5432_ ;
	wire _w5431_ ;
	wire _w5430_ ;
	wire _w5429_ ;
	wire _w5428_ ;
	wire _w5427_ ;
	wire _w5426_ ;
	wire _w5425_ ;
	wire _w5424_ ;
	wire _w5423_ ;
	wire _w5422_ ;
	wire _w5421_ ;
	wire _w5420_ ;
	wire _w5419_ ;
	wire _w5418_ ;
	wire _w5417_ ;
	wire _w5416_ ;
	wire _w5415_ ;
	wire _w5414_ ;
	wire _w5413_ ;
	wire _w5412_ ;
	wire _w5411_ ;
	wire _w5410_ ;
	wire _w5409_ ;
	wire _w5408_ ;
	wire _w5407_ ;
	wire _w5406_ ;
	wire _w5405_ ;
	wire _w5404_ ;
	wire _w5403_ ;
	wire _w5402_ ;
	wire _w5401_ ;
	wire _w5400_ ;
	wire _w5399_ ;
	wire _w5398_ ;
	wire _w5397_ ;
	wire _w5396_ ;
	wire _w5395_ ;
	wire _w5394_ ;
	wire _w5393_ ;
	wire _w5392_ ;
	wire _w5391_ ;
	wire _w5390_ ;
	wire _w5389_ ;
	wire _w5388_ ;
	wire _w5387_ ;
	wire _w5386_ ;
	wire _w5385_ ;
	wire _w5384_ ;
	wire _w5383_ ;
	wire _w5382_ ;
	wire _w5381_ ;
	wire _w5380_ ;
	wire _w5379_ ;
	wire _w5378_ ;
	wire _w5377_ ;
	wire _w5376_ ;
	wire _w5375_ ;
	wire _w5374_ ;
	wire _w5373_ ;
	wire _w5372_ ;
	wire _w5371_ ;
	wire _w5370_ ;
	wire _w5369_ ;
	wire _w5368_ ;
	wire _w5367_ ;
	wire _w5366_ ;
	wire _w5365_ ;
	wire _w5364_ ;
	wire _w5363_ ;
	wire _w5362_ ;
	wire _w5361_ ;
	wire _w5360_ ;
	wire _w5359_ ;
	wire _w5358_ ;
	wire _w5357_ ;
	wire _w5356_ ;
	wire _w5355_ ;
	wire _w5354_ ;
	wire _w5353_ ;
	wire _w5352_ ;
	wire _w5351_ ;
	wire _w5350_ ;
	wire _w5349_ ;
	wire _w5348_ ;
	wire _w5347_ ;
	wire _w5346_ ;
	wire _w5345_ ;
	wire _w5344_ ;
	wire _w5343_ ;
	wire _w5342_ ;
	wire _w5341_ ;
	wire _w5340_ ;
	wire _w5339_ ;
	wire _w5338_ ;
	wire _w5337_ ;
	wire _w5336_ ;
	wire _w5335_ ;
	wire _w5334_ ;
	wire _w5333_ ;
	wire _w5332_ ;
	wire _w5331_ ;
	wire _w5330_ ;
	wire _w5329_ ;
	wire _w5328_ ;
	wire _w5327_ ;
	wire _w5326_ ;
	wire _w5325_ ;
	wire _w5324_ ;
	wire _w5323_ ;
	wire _w5322_ ;
	wire _w5321_ ;
	wire _w5320_ ;
	wire _w5319_ ;
	wire _w5318_ ;
	wire _w5317_ ;
	wire _w5316_ ;
	wire _w5315_ ;
	wire _w5314_ ;
	wire _w5313_ ;
	wire _w5312_ ;
	wire _w5311_ ;
	wire _w5310_ ;
	wire _w5309_ ;
	wire _w5308_ ;
	wire _w5307_ ;
	wire _w5306_ ;
	wire _w5305_ ;
	wire _w5304_ ;
	wire _w5303_ ;
	wire _w5302_ ;
	wire _w5301_ ;
	wire _w5300_ ;
	wire _w5299_ ;
	wire _w5298_ ;
	wire _w5297_ ;
	wire _w5296_ ;
	wire _w5295_ ;
	wire _w5294_ ;
	wire _w5293_ ;
	wire _w5292_ ;
	wire _w5291_ ;
	wire _w5290_ ;
	wire _w5289_ ;
	wire _w5288_ ;
	wire _w5287_ ;
	wire _w5286_ ;
	wire _w5285_ ;
	wire _w5284_ ;
	wire _w5283_ ;
	wire _w5282_ ;
	wire _w5281_ ;
	wire _w5280_ ;
	wire _w5279_ ;
	wire _w5278_ ;
	wire _w5277_ ;
	wire _w5276_ ;
	wire _w5275_ ;
	wire _w5274_ ;
	wire _w5273_ ;
	wire _w5272_ ;
	wire _w5271_ ;
	wire _w5270_ ;
	wire _w5269_ ;
	wire _w5268_ ;
	wire _w5267_ ;
	wire _w5266_ ;
	wire _w5265_ ;
	wire _w5264_ ;
	wire _w5263_ ;
	wire _w5262_ ;
	wire _w5261_ ;
	wire _w5260_ ;
	wire _w5259_ ;
	wire _w5258_ ;
	wire _w5257_ ;
	wire _w5256_ ;
	wire _w5255_ ;
	wire _w5254_ ;
	wire _w5253_ ;
	wire _w5252_ ;
	wire _w5251_ ;
	wire _w5250_ ;
	wire _w5249_ ;
	wire _w5248_ ;
	wire _w5247_ ;
	wire _w5246_ ;
	wire _w5245_ ;
	wire _w5244_ ;
	wire _w5243_ ;
	wire _w5242_ ;
	wire _w5241_ ;
	wire _w5240_ ;
	wire _w5239_ ;
	wire _w5238_ ;
	wire _w5237_ ;
	wire _w5236_ ;
	wire _w5235_ ;
	wire _w5234_ ;
	wire _w5233_ ;
	wire _w5232_ ;
	wire _w5231_ ;
	wire _w5230_ ;
	wire _w5229_ ;
	wire _w5228_ ;
	wire _w5227_ ;
	wire _w5226_ ;
	wire _w5225_ ;
	wire _w5224_ ;
	wire _w5223_ ;
	wire _w5222_ ;
	wire _w5221_ ;
	wire _w5220_ ;
	wire _w5219_ ;
	wire _w5218_ ;
	wire _w5217_ ;
	wire _w5216_ ;
	wire _w5215_ ;
	wire _w5214_ ;
	wire _w5213_ ;
	wire _w5212_ ;
	wire _w5211_ ;
	wire _w5210_ ;
	wire _w5209_ ;
	wire _w5208_ ;
	wire _w5207_ ;
	wire _w5206_ ;
	wire _w5205_ ;
	wire _w5204_ ;
	wire _w5203_ ;
	wire _w5202_ ;
	wire _w5201_ ;
	wire _w5200_ ;
	wire _w5199_ ;
	wire _w5198_ ;
	wire _w5197_ ;
	wire _w5196_ ;
	wire _w5195_ ;
	wire _w5194_ ;
	wire _w5193_ ;
	wire _w5192_ ;
	wire _w5191_ ;
	wire _w5190_ ;
	wire _w5189_ ;
	wire _w5188_ ;
	wire _w5187_ ;
	wire _w5186_ ;
	wire _w5185_ ;
	wire _w5184_ ;
	wire _w5183_ ;
	wire _w5182_ ;
	wire _w5181_ ;
	wire _w5180_ ;
	wire _w5179_ ;
	wire _w5178_ ;
	wire _w5177_ ;
	wire _w5176_ ;
	wire _w5175_ ;
	wire _w5174_ ;
	wire _w5173_ ;
	wire _w5172_ ;
	wire _w5171_ ;
	wire _w5170_ ;
	wire _w5169_ ;
	wire _w5168_ ;
	wire _w5167_ ;
	wire _w5166_ ;
	wire _w5165_ ;
	wire _w5164_ ;
	wire _w5163_ ;
	wire _w5162_ ;
	wire _w5161_ ;
	wire _w5160_ ;
	wire _w5159_ ;
	wire _w5158_ ;
	wire _w5157_ ;
	wire _w5156_ ;
	wire _w5155_ ;
	wire _w5154_ ;
	wire _w5153_ ;
	wire _w5152_ ;
	wire _w5151_ ;
	wire _w5150_ ;
	wire _w5149_ ;
	wire _w5148_ ;
	wire _w5147_ ;
	wire _w5146_ ;
	wire _w5145_ ;
	wire _w5144_ ;
	wire _w5143_ ;
	wire _w5142_ ;
	wire _w5141_ ;
	wire _w5140_ ;
	wire _w5139_ ;
	wire _w5138_ ;
	wire _w5137_ ;
	wire _w5136_ ;
	wire _w5135_ ;
	wire _w5134_ ;
	wire _w5133_ ;
	wire _w5132_ ;
	wire _w5131_ ;
	wire _w5130_ ;
	wire _w5129_ ;
	wire _w5128_ ;
	wire _w5127_ ;
	wire _w5126_ ;
	wire _w5125_ ;
	wire _w5124_ ;
	wire _w5123_ ;
	wire _w5122_ ;
	wire _w5121_ ;
	wire _w5120_ ;
	wire _w5119_ ;
	wire _w5118_ ;
	wire _w5117_ ;
	wire _w5116_ ;
	wire _w5115_ ;
	wire _w5114_ ;
	wire _w5113_ ;
	wire _w5112_ ;
	wire _w5111_ ;
	wire _w5110_ ;
	wire _w5109_ ;
	wire _w5108_ ;
	wire _w5107_ ;
	wire _w5106_ ;
	wire _w5105_ ;
	wire _w5104_ ;
	wire _w5103_ ;
	wire _w5102_ ;
	wire _w5101_ ;
	wire _w5100_ ;
	wire _w5099_ ;
	wire _w5098_ ;
	wire _w5097_ ;
	wire _w5096_ ;
	wire _w5095_ ;
	wire _w5094_ ;
	wire _w5093_ ;
	wire _w5092_ ;
	wire _w5091_ ;
	wire _w5090_ ;
	wire _w5089_ ;
	wire _w5088_ ;
	wire _w5087_ ;
	wire _w5086_ ;
	wire _w5085_ ;
	wire _w5084_ ;
	wire _w5083_ ;
	wire _w5082_ ;
	wire _w5081_ ;
	wire _w5080_ ;
	wire _w5079_ ;
	wire _w5078_ ;
	wire _w5077_ ;
	wire _w5076_ ;
	wire _w5075_ ;
	wire _w5074_ ;
	wire _w5073_ ;
	wire _w5072_ ;
	wire _w5071_ ;
	wire _w5070_ ;
	wire _w5069_ ;
	wire _w5068_ ;
	wire _w5067_ ;
	wire _w5066_ ;
	wire _w5065_ ;
	wire _w5064_ ;
	wire _w5063_ ;
	wire _w5062_ ;
	wire _w5061_ ;
	wire _w5060_ ;
	wire _w5059_ ;
	wire _w5058_ ;
	wire _w5057_ ;
	wire _w5056_ ;
	wire _w5055_ ;
	wire _w5054_ ;
	wire _w5053_ ;
	wire _w5052_ ;
	wire _w5051_ ;
	wire _w5050_ ;
	wire _w5049_ ;
	wire _w5048_ ;
	wire _w5047_ ;
	wire _w5046_ ;
	wire _w5045_ ;
	wire _w5044_ ;
	wire _w5043_ ;
	wire _w5042_ ;
	wire _w5041_ ;
	wire _w5040_ ;
	wire _w5039_ ;
	wire _w5038_ ;
	wire _w5037_ ;
	wire _w5036_ ;
	wire _w5035_ ;
	wire _w5034_ ;
	wire _w5033_ ;
	wire _w5032_ ;
	wire _w5031_ ;
	wire _w5030_ ;
	wire _w5029_ ;
	wire _w5028_ ;
	wire _w5027_ ;
	wire _w5026_ ;
	wire _w5025_ ;
	wire _w5024_ ;
	wire _w5023_ ;
	wire _w5022_ ;
	wire _w5021_ ;
	wire _w5020_ ;
	wire _w5019_ ;
	wire _w5018_ ;
	wire _w5017_ ;
	wire _w5016_ ;
	wire _w5015_ ;
	wire _w5014_ ;
	wire _w5013_ ;
	wire _w5012_ ;
	wire _w5011_ ;
	wire _w5010_ ;
	wire _w5009_ ;
	wire _w5008_ ;
	wire _w5007_ ;
	wire _w5006_ ;
	wire _w5005_ ;
	wire _w5004_ ;
	wire _w5003_ ;
	wire _w5002_ ;
	wire _w5001_ ;
	wire _w5000_ ;
	wire _w4999_ ;
	wire _w4998_ ;
	wire _w4997_ ;
	wire _w4996_ ;
	wire _w4995_ ;
	wire _w4994_ ;
	wire _w4993_ ;
	wire _w4992_ ;
	wire _w4991_ ;
	wire _w4990_ ;
	wire _w4989_ ;
	wire _w4988_ ;
	wire _w4987_ ;
	wire _w4986_ ;
	wire _w4985_ ;
	wire _w4984_ ;
	wire _w4983_ ;
	wire _w4982_ ;
	wire _w4981_ ;
	wire _w4980_ ;
	wire _w4979_ ;
	wire _w4978_ ;
	wire _w4977_ ;
	wire _w4976_ ;
	wire _w4975_ ;
	wire _w4974_ ;
	wire _w4973_ ;
	wire _w4972_ ;
	wire _w4971_ ;
	wire _w4970_ ;
	wire _w4969_ ;
	wire _w4968_ ;
	wire _w4967_ ;
	wire _w4966_ ;
	wire _w4965_ ;
	wire _w4964_ ;
	wire _w4963_ ;
	wire _w4962_ ;
	wire _w4961_ ;
	wire _w4960_ ;
	wire _w4959_ ;
	wire _w4958_ ;
	wire _w4957_ ;
	wire _w4956_ ;
	wire _w4955_ ;
	wire _w4954_ ;
	wire _w4953_ ;
	wire _w4952_ ;
	wire _w4951_ ;
	wire _w4950_ ;
	wire _w4949_ ;
	wire _w4948_ ;
	wire _w4947_ ;
	wire _w4946_ ;
	wire _w4945_ ;
	wire _w4944_ ;
	wire _w4943_ ;
	wire _w4942_ ;
	wire _w4941_ ;
	wire _w4940_ ;
	wire _w4939_ ;
	wire _w4938_ ;
	wire _w4937_ ;
	wire _w4936_ ;
	wire _w4935_ ;
	wire _w4934_ ;
	wire _w4933_ ;
	wire _w4932_ ;
	wire _w4931_ ;
	wire _w4930_ ;
	wire _w4929_ ;
	wire _w4928_ ;
	wire _w4927_ ;
	wire _w4926_ ;
	wire _w4925_ ;
	wire _w4924_ ;
	wire _w4923_ ;
	wire _w4922_ ;
	wire _w4921_ ;
	wire _w4920_ ;
	wire _w4919_ ;
	wire _w4918_ ;
	wire _w4917_ ;
	wire _w4916_ ;
	wire _w4915_ ;
	wire _w4914_ ;
	wire _w4913_ ;
	wire _w4912_ ;
	wire _w4911_ ;
	wire _w4910_ ;
	wire _w4909_ ;
	wire _w4908_ ;
	wire _w4907_ ;
	wire _w4906_ ;
	wire _w4905_ ;
	wire _w4904_ ;
	wire _w4903_ ;
	wire _w4902_ ;
	wire _w4901_ ;
	wire _w4900_ ;
	wire _w4899_ ;
	wire _w4898_ ;
	wire _w4897_ ;
	wire _w4896_ ;
	wire _w4895_ ;
	wire _w4894_ ;
	wire _w4893_ ;
	wire _w4892_ ;
	wire _w4891_ ;
	wire _w4890_ ;
	wire _w4889_ ;
	wire _w4888_ ;
	wire _w4887_ ;
	wire _w4886_ ;
	wire _w4885_ ;
	wire _w4884_ ;
	wire _w4883_ ;
	wire _w4882_ ;
	wire _w4881_ ;
	wire _w4880_ ;
	wire _w4879_ ;
	wire _w4878_ ;
	wire _w4877_ ;
	wire _w4876_ ;
	wire _w4875_ ;
	wire _w4874_ ;
	wire _w4873_ ;
	wire _w4872_ ;
	wire _w4871_ ;
	wire _w4870_ ;
	wire _w4869_ ;
	wire _w4868_ ;
	wire _w4867_ ;
	wire _w4866_ ;
	wire _w4865_ ;
	wire _w4864_ ;
	wire _w4863_ ;
	wire _w4862_ ;
	wire _w4861_ ;
	wire _w4860_ ;
	wire _w4859_ ;
	wire _w4858_ ;
	wire _w4857_ ;
	wire _w4856_ ;
	wire _w4855_ ;
	wire _w4854_ ;
	wire _w4853_ ;
	wire _w4852_ ;
	wire _w4851_ ;
	wire _w4850_ ;
	wire _w4849_ ;
	wire _w4848_ ;
	wire _w4847_ ;
	wire _w4846_ ;
	wire _w4845_ ;
	wire _w4844_ ;
	wire _w4843_ ;
	wire _w4842_ ;
	wire _w4841_ ;
	wire _w4840_ ;
	wire _w4839_ ;
	wire _w4838_ ;
	wire _w4837_ ;
	wire _w4836_ ;
	wire _w4835_ ;
	wire _w4834_ ;
	wire _w4833_ ;
	wire _w4832_ ;
	wire _w4831_ ;
	wire _w4830_ ;
	wire _w4829_ ;
	wire _w4828_ ;
	wire _w4827_ ;
	wire _w4826_ ;
	wire _w4825_ ;
	wire _w4824_ ;
	wire _w4823_ ;
	wire _w4822_ ;
	wire _w4821_ ;
	wire _w4820_ ;
	wire _w4819_ ;
	wire _w4818_ ;
	wire _w4817_ ;
	wire _w4816_ ;
	wire _w4815_ ;
	wire _w4814_ ;
	wire _w4813_ ;
	wire _w4812_ ;
	wire _w4811_ ;
	wire _w4810_ ;
	wire _w4809_ ;
	wire _w4808_ ;
	wire _w4807_ ;
	wire _w4806_ ;
	wire _w4805_ ;
	wire _w4804_ ;
	wire _w4803_ ;
	wire _w4802_ ;
	wire _w4801_ ;
	wire _w4800_ ;
	wire _w4799_ ;
	wire _w4798_ ;
	wire _w4797_ ;
	wire _w4796_ ;
	wire _w4795_ ;
	wire _w4794_ ;
	wire _w4793_ ;
	wire _w4792_ ;
	wire _w4791_ ;
	wire _w4790_ ;
	wire _w4789_ ;
	wire _w4788_ ;
	wire _w4787_ ;
	wire _w4786_ ;
	wire _w4785_ ;
	wire _w4784_ ;
	wire _w4783_ ;
	wire _w4782_ ;
	wire _w4781_ ;
	wire _w4780_ ;
	wire _w4779_ ;
	wire _w4778_ ;
	wire _w4777_ ;
	wire _w4776_ ;
	wire _w4775_ ;
	wire _w4774_ ;
	wire _w4773_ ;
	wire _w4772_ ;
	wire _w4771_ ;
	wire _w4770_ ;
	wire _w4769_ ;
	wire _w4768_ ;
	wire _w4767_ ;
	wire _w4766_ ;
	wire _w4765_ ;
	wire _w4764_ ;
	wire _w4763_ ;
	wire _w4762_ ;
	wire _w4761_ ;
	wire _w4760_ ;
	wire _w4759_ ;
	wire _w4758_ ;
	wire _w4757_ ;
	wire _w4756_ ;
	wire _w4755_ ;
	wire _w4754_ ;
	wire _w4753_ ;
	wire _w4752_ ;
	wire _w4751_ ;
	wire _w4750_ ;
	wire _w4749_ ;
	wire _w4748_ ;
	wire _w4747_ ;
	wire _w4746_ ;
	wire _w4745_ ;
	wire _w4744_ ;
	wire _w4743_ ;
	wire _w4742_ ;
	wire _w4741_ ;
	wire _w4740_ ;
	wire _w4739_ ;
	wire _w4738_ ;
	wire _w4737_ ;
	wire _w4736_ ;
	wire _w4735_ ;
	wire _w4734_ ;
	wire _w4733_ ;
	wire _w4732_ ;
	wire _w4731_ ;
	wire _w4730_ ;
	wire _w4729_ ;
	wire _w4728_ ;
	wire _w4727_ ;
	wire _w4726_ ;
	wire _w4725_ ;
	wire _w4724_ ;
	wire _w4723_ ;
	wire _w4722_ ;
	wire _w4721_ ;
	wire _w4720_ ;
	wire _w4719_ ;
	wire _w4718_ ;
	wire _w4717_ ;
	wire _w4716_ ;
	wire _w4715_ ;
	wire _w4714_ ;
	wire _w4713_ ;
	wire _w4712_ ;
	wire _w4711_ ;
	wire _w4710_ ;
	wire _w4709_ ;
	wire _w4708_ ;
	wire _w4707_ ;
	wire _w4706_ ;
	wire _w4705_ ;
	wire _w4704_ ;
	wire _w4703_ ;
	wire _w4702_ ;
	wire _w4701_ ;
	wire _w4700_ ;
	wire _w4699_ ;
	wire _w4698_ ;
	wire _w4697_ ;
	wire _w4696_ ;
	wire _w4695_ ;
	wire _w4694_ ;
	wire _w4693_ ;
	wire _w4692_ ;
	wire _w4691_ ;
	wire _w4690_ ;
	wire _w4689_ ;
	wire _w4688_ ;
	wire _w4687_ ;
	wire _w4686_ ;
	wire _w4685_ ;
	wire _w4684_ ;
	wire _w4683_ ;
	wire _w4682_ ;
	wire _w4681_ ;
	wire _w4680_ ;
	wire _w4679_ ;
	wire _w4678_ ;
	wire _w4677_ ;
	wire _w4676_ ;
	wire _w4675_ ;
	wire _w4674_ ;
	wire _w4673_ ;
	wire _w4672_ ;
	wire _w4671_ ;
	wire _w4670_ ;
	wire _w4669_ ;
	wire _w4668_ ;
	wire _w4667_ ;
	wire _w4666_ ;
	wire _w4665_ ;
	wire _w4664_ ;
	wire _w4663_ ;
	wire _w4662_ ;
	wire _w4661_ ;
	wire _w4660_ ;
	wire _w4659_ ;
	wire _w4658_ ;
	wire _w4657_ ;
	wire _w4656_ ;
	wire _w4655_ ;
	wire _w4654_ ;
	wire _w4653_ ;
	wire _w4652_ ;
	wire _w4651_ ;
	wire _w4650_ ;
	wire _w4649_ ;
	wire _w4648_ ;
	wire _w4647_ ;
	wire _w4646_ ;
	wire _w4645_ ;
	wire _w4644_ ;
	wire _w4643_ ;
	wire _w4642_ ;
	wire _w4641_ ;
	wire _w4640_ ;
	wire _w4639_ ;
	wire _w4638_ ;
	wire _w4637_ ;
	wire _w4636_ ;
	wire _w4635_ ;
	wire _w4634_ ;
	wire _w4633_ ;
	wire _w4632_ ;
	wire _w4631_ ;
	wire _w4630_ ;
	wire _w4629_ ;
	wire _w4628_ ;
	wire _w4627_ ;
	wire _w4626_ ;
	wire _w4625_ ;
	wire _w4624_ ;
	wire _w4623_ ;
	wire _w4622_ ;
	wire _w4621_ ;
	wire _w4620_ ;
	wire _w4619_ ;
	wire _w4618_ ;
	wire _w4617_ ;
	wire _w4616_ ;
	wire _w4615_ ;
	wire _w4614_ ;
	wire _w4613_ ;
	wire _w4612_ ;
	wire _w4611_ ;
	wire _w4610_ ;
	wire _w4609_ ;
	wire _w4608_ ;
	wire _w4607_ ;
	wire _w4606_ ;
	wire _w4605_ ;
	wire _w4604_ ;
	wire _w4603_ ;
	wire _w4602_ ;
	wire _w4601_ ;
	wire _w4600_ ;
	wire _w4599_ ;
	wire _w4598_ ;
	wire _w4597_ ;
	wire _w4596_ ;
	wire _w4595_ ;
	wire _w4594_ ;
	wire _w4593_ ;
	wire _w4592_ ;
	wire _w4591_ ;
	wire _w4590_ ;
	wire _w4589_ ;
	wire _w4588_ ;
	wire _w4587_ ;
	wire _w4586_ ;
	wire _w4585_ ;
	wire _w4584_ ;
	wire _w4583_ ;
	wire _w4582_ ;
	wire _w4581_ ;
	wire _w4580_ ;
	wire _w4579_ ;
	wire _w4578_ ;
	wire _w4577_ ;
	wire _w4576_ ;
	wire _w4575_ ;
	wire _w4574_ ;
	wire _w4573_ ;
	wire _w4572_ ;
	wire _w4571_ ;
	wire _w4570_ ;
	wire _w4569_ ;
	wire _w4568_ ;
	wire _w4567_ ;
	wire _w4566_ ;
	wire _w4565_ ;
	wire _w4564_ ;
	wire _w4563_ ;
	wire _w4562_ ;
	wire _w4561_ ;
	wire _w4560_ ;
	wire _w4559_ ;
	wire _w4558_ ;
	wire _w4557_ ;
	wire _w4556_ ;
	wire _w4555_ ;
	wire _w4554_ ;
	wire _w4553_ ;
	wire _w4552_ ;
	wire _w4551_ ;
	wire _w4550_ ;
	wire _w4549_ ;
	wire _w4548_ ;
	wire _w4547_ ;
	wire _w4546_ ;
	wire _w4545_ ;
	wire _w4544_ ;
	wire _w4543_ ;
	wire _w4542_ ;
	wire _w4541_ ;
	wire _w4540_ ;
	wire _w4539_ ;
	wire _w4538_ ;
	wire _w4537_ ;
	wire _w4536_ ;
	wire _w4535_ ;
	wire _w4534_ ;
	wire _w4533_ ;
	wire _w4532_ ;
	wire _w4531_ ;
	wire _w4530_ ;
	wire _w4529_ ;
	wire _w4528_ ;
	wire _w4527_ ;
	wire _w4526_ ;
	wire _w4525_ ;
	wire _w4524_ ;
	wire _w4523_ ;
	wire _w4522_ ;
	wire _w4521_ ;
	wire _w4520_ ;
	wire _w4519_ ;
	wire _w4518_ ;
	wire _w4517_ ;
	wire _w4516_ ;
	wire _w4515_ ;
	wire _w4514_ ;
	wire _w4513_ ;
	wire _w4512_ ;
	wire _w4511_ ;
	wire _w4510_ ;
	wire _w4509_ ;
	wire _w4508_ ;
	wire _w4507_ ;
	wire _w4506_ ;
	wire _w4505_ ;
	wire _w4504_ ;
	wire _w4503_ ;
	wire _w4502_ ;
	wire _w4501_ ;
	wire _w4500_ ;
	wire _w4499_ ;
	wire _w4498_ ;
	wire _w4497_ ;
	wire _w4496_ ;
	wire _w4495_ ;
	wire _w4494_ ;
	wire _w4493_ ;
	wire _w4492_ ;
	wire _w4491_ ;
	wire _w4490_ ;
	wire _w4489_ ;
	wire _w4488_ ;
	wire _w4487_ ;
	wire _w4486_ ;
	wire _w4485_ ;
	wire _w4484_ ;
	wire _w4483_ ;
	wire _w4482_ ;
	wire _w4481_ ;
	wire _w4480_ ;
	wire _w4479_ ;
	wire _w4478_ ;
	wire _w4477_ ;
	wire _w4476_ ;
	wire _w4475_ ;
	wire _w4474_ ;
	wire _w4473_ ;
	wire _w4472_ ;
	wire _w4471_ ;
	wire _w4470_ ;
	wire _w4469_ ;
	wire _w4468_ ;
	wire _w4467_ ;
	wire _w4466_ ;
	wire _w4465_ ;
	wire _w4464_ ;
	wire _w4463_ ;
	wire _w4462_ ;
	wire _w4461_ ;
	wire _w4460_ ;
	wire _w4459_ ;
	wire _w4458_ ;
	wire _w4457_ ;
	wire _w4456_ ;
	wire _w4455_ ;
	wire _w4454_ ;
	wire _w4453_ ;
	wire _w4452_ ;
	wire _w4451_ ;
	wire _w4450_ ;
	wire _w4449_ ;
	wire _w4448_ ;
	wire _w4447_ ;
	wire _w4446_ ;
	wire _w4445_ ;
	wire _w4444_ ;
	wire _w4443_ ;
	wire _w4442_ ;
	wire _w4441_ ;
	wire _w4440_ ;
	wire _w4439_ ;
	wire _w4438_ ;
	wire _w4437_ ;
	wire _w4436_ ;
	wire _w4435_ ;
	wire _w4434_ ;
	wire _w4433_ ;
	wire _w4432_ ;
	wire _w4431_ ;
	wire _w4430_ ;
	wire _w4429_ ;
	wire _w4428_ ;
	wire _w4427_ ;
	wire _w4426_ ;
	wire _w4425_ ;
	wire _w4424_ ;
	wire _w4423_ ;
	wire _w4422_ ;
	wire _w4421_ ;
	wire _w4420_ ;
	wire _w4419_ ;
	wire _w4418_ ;
	wire _w4417_ ;
	wire _w4416_ ;
	wire _w4415_ ;
	wire _w4414_ ;
	wire _w4413_ ;
	wire _w4412_ ;
	wire _w4411_ ;
	wire _w4410_ ;
	wire _w4409_ ;
	wire _w4408_ ;
	wire _w4407_ ;
	wire _w4406_ ;
	wire _w4405_ ;
	wire _w4404_ ;
	wire _w4403_ ;
	wire _w4402_ ;
	wire _w4401_ ;
	wire _w4400_ ;
	wire _w4399_ ;
	wire _w4398_ ;
	wire _w4397_ ;
	wire _w4396_ ;
	wire _w4395_ ;
	wire _w4394_ ;
	wire _w4393_ ;
	wire _w4392_ ;
	wire _w4391_ ;
	wire _w4390_ ;
	wire _w4389_ ;
	wire _w4388_ ;
	wire _w4387_ ;
	wire _w4386_ ;
	wire _w4385_ ;
	wire _w4384_ ;
	wire _w4383_ ;
	wire _w4382_ ;
	wire _w4381_ ;
	wire _w4380_ ;
	wire _w4379_ ;
	wire _w4378_ ;
	wire _w4377_ ;
	wire _w4376_ ;
	wire _w4375_ ;
	wire _w4374_ ;
	wire _w4373_ ;
	wire _w4372_ ;
	wire _w4371_ ;
	wire _w4370_ ;
	wire _w4369_ ;
	wire _w4368_ ;
	wire _w4367_ ;
	wire _w4366_ ;
	wire _w4365_ ;
	wire _w4364_ ;
	wire _w4363_ ;
	wire _w4362_ ;
	wire _w4361_ ;
	wire _w4360_ ;
	wire _w4359_ ;
	wire _w4358_ ;
	wire _w4357_ ;
	wire _w4356_ ;
	wire _w4355_ ;
	wire _w4354_ ;
	wire _w4353_ ;
	wire _w4352_ ;
	wire _w4351_ ;
	wire _w4350_ ;
	wire _w4349_ ;
	wire _w4348_ ;
	wire _w4347_ ;
	wire _w4346_ ;
	wire _w4345_ ;
	wire _w4344_ ;
	wire _w4343_ ;
	wire _w4342_ ;
	wire _w4341_ ;
	wire _w4340_ ;
	wire _w4339_ ;
	wire _w4338_ ;
	wire _w4337_ ;
	wire _w4336_ ;
	wire _w4335_ ;
	wire _w4334_ ;
	wire _w4333_ ;
	wire _w4332_ ;
	wire _w4331_ ;
	wire _w4330_ ;
	wire _w4329_ ;
	wire _w4328_ ;
	wire _w4327_ ;
	wire _w4326_ ;
	wire _w4325_ ;
	wire _w4324_ ;
	wire _w4323_ ;
	wire _w4322_ ;
	wire _w4321_ ;
	wire _w4320_ ;
	wire _w4319_ ;
	wire _w4318_ ;
	wire _w4317_ ;
	wire _w4316_ ;
	wire _w4315_ ;
	wire _w4314_ ;
	wire _w4313_ ;
	wire _w4312_ ;
	wire _w4311_ ;
	wire _w4310_ ;
	wire _w4309_ ;
	wire _w4308_ ;
	wire _w4307_ ;
	wire _w4306_ ;
	wire _w4305_ ;
	wire _w4304_ ;
	wire _w4303_ ;
	wire _w4302_ ;
	wire _w4301_ ;
	wire _w4300_ ;
	wire _w4299_ ;
	wire _w4298_ ;
	wire _w4297_ ;
	wire _w4296_ ;
	wire _w4295_ ;
	wire _w4294_ ;
	wire _w4293_ ;
	wire _w4292_ ;
	wire _w4291_ ;
	wire _w4290_ ;
	wire _w4289_ ;
	wire _w4288_ ;
	wire _w4287_ ;
	wire _w4286_ ;
	wire _w4285_ ;
	wire _w4284_ ;
	wire _w4283_ ;
	wire _w4282_ ;
	wire _w4281_ ;
	wire _w4280_ ;
	wire _w4279_ ;
	wire _w4278_ ;
	wire _w4277_ ;
	wire _w4276_ ;
	wire _w4275_ ;
	wire _w4274_ ;
	wire _w4273_ ;
	wire _w4272_ ;
	wire _w4271_ ;
	wire _w4270_ ;
	wire _w4269_ ;
	wire _w4268_ ;
	wire _w4267_ ;
	wire _w4266_ ;
	wire _w4265_ ;
	wire _w4264_ ;
	wire _w4263_ ;
	wire _w4262_ ;
	wire _w4261_ ;
	wire _w4260_ ;
	wire _w4259_ ;
	wire _w4258_ ;
	wire _w4257_ ;
	wire _w4256_ ;
	wire _w4255_ ;
	wire _w4254_ ;
	wire _w4253_ ;
	wire _w4252_ ;
	wire _w4251_ ;
	wire _w4250_ ;
	wire _w4249_ ;
	wire _w4248_ ;
	wire _w4247_ ;
	wire _w4246_ ;
	wire _w4245_ ;
	wire _w4244_ ;
	wire _w4243_ ;
	wire _w4242_ ;
	wire _w4241_ ;
	wire _w4240_ ;
	wire _w4239_ ;
	wire _w4238_ ;
	wire _w4237_ ;
	wire _w4236_ ;
	wire _w4235_ ;
	wire _w4234_ ;
	wire _w4233_ ;
	wire _w4232_ ;
	wire _w4231_ ;
	wire _w4230_ ;
	wire _w4229_ ;
	wire _w4228_ ;
	wire _w4227_ ;
	wire _w4226_ ;
	wire _w4225_ ;
	wire _w4224_ ;
	wire _w4223_ ;
	wire _w4222_ ;
	wire _w4221_ ;
	wire _w4220_ ;
	wire _w4219_ ;
	wire _w4218_ ;
	wire _w4217_ ;
	wire _w4216_ ;
	wire _w4215_ ;
	wire _w4214_ ;
	wire _w4213_ ;
	wire _w4212_ ;
	wire _w4211_ ;
	wire _w4210_ ;
	wire _w4209_ ;
	wire _w4208_ ;
	wire _w4207_ ;
	wire _w4206_ ;
	wire _w4205_ ;
	wire _w4204_ ;
	wire _w4203_ ;
	wire _w4202_ ;
	wire _w4201_ ;
	wire _w4200_ ;
	wire _w4199_ ;
	wire _w4198_ ;
	wire _w4197_ ;
	wire _w4196_ ;
	wire _w4195_ ;
	wire _w4194_ ;
	wire _w4193_ ;
	wire _w4192_ ;
	wire _w4191_ ;
	wire _w4190_ ;
	wire _w4189_ ;
	wire _w4188_ ;
	wire _w4187_ ;
	wire _w4186_ ;
	wire _w4185_ ;
	wire _w4184_ ;
	wire _w4183_ ;
	wire _w4182_ ;
	wire _w4181_ ;
	wire _w4180_ ;
	wire _w4179_ ;
	wire _w4178_ ;
	wire _w4177_ ;
	wire _w4176_ ;
	wire _w4175_ ;
	wire _w4174_ ;
	wire _w4173_ ;
	wire _w4172_ ;
	wire _w4171_ ;
	wire _w4170_ ;
	wire _w4169_ ;
	wire _w4168_ ;
	wire _w4167_ ;
	wire _w4166_ ;
	wire _w4165_ ;
	wire _w4164_ ;
	wire _w4163_ ;
	wire _w4162_ ;
	wire _w4161_ ;
	wire _w4160_ ;
	wire _w4159_ ;
	wire _w4158_ ;
	wire _w4157_ ;
	wire _w4156_ ;
	wire _w4155_ ;
	wire _w4154_ ;
	wire _w4153_ ;
	wire _w4152_ ;
	wire _w4151_ ;
	wire _w4150_ ;
	wire _w4149_ ;
	wire _w4148_ ;
	wire _w4147_ ;
	wire _w4146_ ;
	wire _w4145_ ;
	wire _w4144_ ;
	wire _w4143_ ;
	wire _w4142_ ;
	wire _w4141_ ;
	wire _w4140_ ;
	wire _w4139_ ;
	wire _w4138_ ;
	wire _w4137_ ;
	wire _w4136_ ;
	wire _w4135_ ;
	wire _w4134_ ;
	wire _w4133_ ;
	wire _w4132_ ;
	wire _w4131_ ;
	wire _w4130_ ;
	wire _w4129_ ;
	wire _w4128_ ;
	wire _w4127_ ;
	wire _w4126_ ;
	wire _w4125_ ;
	wire _w4124_ ;
	wire _w4123_ ;
	wire _w4122_ ;
	wire _w4121_ ;
	wire _w4120_ ;
	wire _w4119_ ;
	wire _w4118_ ;
	wire _w4117_ ;
	wire _w4116_ ;
	wire _w4115_ ;
	wire _w4114_ ;
	wire _w4113_ ;
	wire _w4112_ ;
	wire _w4111_ ;
	wire _w4110_ ;
	wire _w4109_ ;
	wire _w4108_ ;
	wire _w4107_ ;
	wire _w4106_ ;
	wire _w4105_ ;
	wire _w4104_ ;
	wire _w4103_ ;
	wire _w4102_ ;
	wire _w4101_ ;
	wire _w4100_ ;
	wire _w4099_ ;
	wire _w4098_ ;
	wire _w4097_ ;
	wire _w4096_ ;
	wire _w4095_ ;
	wire _w4094_ ;
	wire _w4093_ ;
	wire _w4092_ ;
	wire _w4091_ ;
	wire _w4090_ ;
	wire _w4089_ ;
	wire _w4088_ ;
	wire _w4087_ ;
	wire _w4086_ ;
	wire _w4085_ ;
	wire _w4084_ ;
	wire _w4083_ ;
	wire _w4082_ ;
	wire _w4081_ ;
	wire _w4080_ ;
	wire _w4079_ ;
	wire _w4078_ ;
	wire _w4077_ ;
	wire _w4076_ ;
	wire _w4075_ ;
	wire _w4074_ ;
	wire _w4073_ ;
	wire _w4072_ ;
	wire _w4071_ ;
	wire _w4070_ ;
	wire _w4069_ ;
	wire _w4068_ ;
	wire _w4067_ ;
	wire _w4066_ ;
	wire _w4065_ ;
	wire _w4064_ ;
	wire _w4063_ ;
	wire _w4062_ ;
	wire _w4061_ ;
	wire _w4060_ ;
	wire _w4059_ ;
	wire _w4058_ ;
	wire _w4057_ ;
	wire _w4056_ ;
	wire _w4055_ ;
	wire _w4054_ ;
	wire _w4053_ ;
	wire _w4052_ ;
	wire _w4051_ ;
	wire _w4050_ ;
	wire _w4049_ ;
	wire _w4048_ ;
	wire _w4047_ ;
	wire _w4046_ ;
	wire _w4045_ ;
	wire _w4044_ ;
	wire _w4043_ ;
	wire _w4042_ ;
	wire _w4041_ ;
	wire _w4040_ ;
	wire _w4039_ ;
	wire _w4038_ ;
	wire _w4037_ ;
	wire _w4036_ ;
	wire _w4035_ ;
	wire _w4034_ ;
	wire _w4033_ ;
	wire _w4032_ ;
	wire _w4031_ ;
	wire _w4030_ ;
	wire _w4029_ ;
	wire _w4028_ ;
	wire _w4027_ ;
	wire _w4026_ ;
	wire _w4025_ ;
	wire _w4024_ ;
	wire _w4023_ ;
	wire _w4022_ ;
	wire _w4021_ ;
	wire _w4020_ ;
	wire _w4019_ ;
	wire _w4018_ ;
	wire _w4017_ ;
	wire _w4016_ ;
	wire _w4015_ ;
	wire _w4014_ ;
	wire _w4013_ ;
	wire _w4012_ ;
	wire _w4011_ ;
	wire _w4010_ ;
	wire _w4009_ ;
	wire _w4008_ ;
	wire _w4007_ ;
	wire _w4006_ ;
	wire _w4005_ ;
	wire _w4004_ ;
	wire _w4003_ ;
	wire _w4002_ ;
	wire _w4001_ ;
	wire _w4000_ ;
	wire _w3999_ ;
	wire _w3998_ ;
	wire _w3997_ ;
	wire _w3996_ ;
	wire _w3995_ ;
	wire _w3994_ ;
	wire _w3993_ ;
	wire _w3992_ ;
	wire _w3991_ ;
	wire _w3990_ ;
	wire _w3989_ ;
	wire _w3988_ ;
	wire _w3987_ ;
	wire _w3986_ ;
	wire _w3985_ ;
	wire _w3984_ ;
	wire _w3983_ ;
	wire _w3982_ ;
	wire _w3981_ ;
	wire _w3980_ ;
	wire _w3979_ ;
	wire _w3978_ ;
	wire _w3977_ ;
	wire _w3976_ ;
	wire _w3975_ ;
	wire _w3974_ ;
	wire _w3973_ ;
	wire _w3972_ ;
	wire _w3971_ ;
	wire _w3970_ ;
	wire _w3969_ ;
	wire _w3968_ ;
	wire _w3967_ ;
	wire _w3966_ ;
	wire _w3965_ ;
	wire _w3964_ ;
	wire _w3963_ ;
	wire _w3962_ ;
	wire _w3961_ ;
	wire _w3960_ ;
	wire _w3959_ ;
	wire _w3958_ ;
	wire _w3957_ ;
	wire _w3956_ ;
	wire _w3955_ ;
	wire _w3954_ ;
	wire _w3953_ ;
	wire _w3952_ ;
	wire _w3951_ ;
	wire _w3950_ ;
	wire _w3949_ ;
	wire _w3948_ ;
	wire _w3947_ ;
	wire _w3946_ ;
	wire _w3945_ ;
	wire _w3944_ ;
	wire _w3943_ ;
	wire _w3942_ ;
	wire _w3941_ ;
	wire _w3940_ ;
	wire _w3939_ ;
	wire _w3938_ ;
	wire _w3937_ ;
	wire _w3936_ ;
	wire _w3935_ ;
	wire _w3934_ ;
	wire _w3933_ ;
	wire _w3932_ ;
	wire _w3931_ ;
	wire _w3930_ ;
	wire _w3929_ ;
	wire _w3928_ ;
	wire _w3927_ ;
	wire _w3926_ ;
	wire _w3925_ ;
	wire _w3924_ ;
	wire _w3923_ ;
	wire _w3922_ ;
	wire _w3921_ ;
	wire _w3920_ ;
	wire _w3919_ ;
	wire _w3918_ ;
	wire _w3917_ ;
	wire _w3916_ ;
	wire _w3915_ ;
	wire _w3914_ ;
	wire _w3913_ ;
	wire _w3912_ ;
	wire _w3911_ ;
	wire _w3910_ ;
	wire _w3909_ ;
	wire _w3908_ ;
	wire _w3907_ ;
	wire _w3906_ ;
	wire _w3905_ ;
	wire _w3904_ ;
	wire _w3903_ ;
	wire _w3902_ ;
	wire _w3901_ ;
	wire _w3900_ ;
	wire _w3899_ ;
	wire _w3898_ ;
	wire _w3897_ ;
	wire _w3896_ ;
	wire _w3895_ ;
	wire _w3894_ ;
	wire _w3893_ ;
	wire _w3892_ ;
	wire _w3891_ ;
	wire _w3890_ ;
	wire _w3889_ ;
	wire _w3888_ ;
	wire _w3887_ ;
	wire _w3886_ ;
	wire _w3885_ ;
	wire _w3884_ ;
	wire _w3883_ ;
	wire _w3882_ ;
	wire _w3881_ ;
	wire _w3880_ ;
	wire _w3879_ ;
	wire _w3878_ ;
	wire _w3877_ ;
	wire _w3876_ ;
	wire _w3875_ ;
	wire _w3874_ ;
	wire _w3873_ ;
	wire _w3872_ ;
	wire _w3871_ ;
	wire _w3870_ ;
	wire _w3869_ ;
	wire _w3868_ ;
	wire _w3867_ ;
	wire _w3866_ ;
	wire _w3865_ ;
	wire _w3864_ ;
	wire _w3863_ ;
	wire _w3862_ ;
	wire _w3861_ ;
	wire _w3860_ ;
	wire _w3859_ ;
	wire _w3858_ ;
	wire _w3857_ ;
	wire _w3856_ ;
	wire _w3855_ ;
	wire _w3854_ ;
	wire _w3853_ ;
	wire _w3852_ ;
	wire _w3851_ ;
	wire _w3850_ ;
	wire _w3849_ ;
	wire _w3848_ ;
	wire _w3847_ ;
	wire _w3846_ ;
	wire _w3845_ ;
	wire _w3844_ ;
	wire _w3843_ ;
	wire _w3842_ ;
	wire _w3841_ ;
	wire _w3840_ ;
	wire _w3839_ ;
	wire _w3838_ ;
	wire _w3837_ ;
	wire _w3836_ ;
	wire _w3835_ ;
	wire _w3834_ ;
	wire _w3833_ ;
	wire _w3832_ ;
	wire _w3831_ ;
	wire _w3830_ ;
	wire _w3829_ ;
	wire _w3828_ ;
	wire _w3827_ ;
	wire _w3826_ ;
	wire _w3825_ ;
	wire _w3824_ ;
	wire _w3823_ ;
	wire _w3822_ ;
	wire _w3821_ ;
	wire _w3820_ ;
	wire _w3819_ ;
	wire _w3818_ ;
	wire _w3817_ ;
	wire _w3816_ ;
	wire _w3815_ ;
	wire _w3814_ ;
	wire _w3813_ ;
	wire _w3812_ ;
	wire _w3811_ ;
	wire _w3810_ ;
	wire _w3809_ ;
	wire _w3808_ ;
	wire _w3807_ ;
	wire _w3806_ ;
	wire _w3805_ ;
	wire _w3804_ ;
	wire _w3803_ ;
	wire _w3802_ ;
	wire _w3801_ ;
	wire _w3800_ ;
	wire _w3799_ ;
	wire _w3798_ ;
	wire _w3797_ ;
	wire _w3796_ ;
	wire _w3795_ ;
	wire _w3794_ ;
	wire _w3793_ ;
	wire _w3792_ ;
	wire _w3791_ ;
	wire _w3790_ ;
	wire _w3789_ ;
	wire _w3788_ ;
	wire _w3787_ ;
	wire _w3786_ ;
	wire _w3785_ ;
	wire _w3784_ ;
	wire _w3783_ ;
	wire _w3782_ ;
	wire _w3781_ ;
	wire _w3780_ ;
	wire _w3779_ ;
	wire _w3778_ ;
	wire _w3777_ ;
	wire _w3776_ ;
	wire _w3775_ ;
	wire _w3774_ ;
	wire _w3773_ ;
	wire _w3772_ ;
	wire _w3771_ ;
	wire _w3770_ ;
	wire _w3769_ ;
	wire _w3768_ ;
	wire _w3767_ ;
	wire _w3766_ ;
	wire _w3765_ ;
	wire _w3764_ ;
	wire _w3763_ ;
	wire _w3762_ ;
	wire _w3761_ ;
	wire _w3760_ ;
	wire _w3759_ ;
	wire _w3758_ ;
	wire _w3757_ ;
	wire _w3756_ ;
	wire _w3755_ ;
	wire _w3754_ ;
	wire _w3753_ ;
	wire _w3752_ ;
	wire _w3751_ ;
	wire _w3750_ ;
	wire _w3749_ ;
	wire _w3748_ ;
	wire _w3747_ ;
	wire _w3746_ ;
	wire _w3745_ ;
	wire _w3744_ ;
	wire _w3743_ ;
	wire _w3742_ ;
	wire _w3741_ ;
	wire _w3740_ ;
	wire _w3739_ ;
	wire _w3738_ ;
	wire _w3737_ ;
	wire _w3736_ ;
	wire _w3735_ ;
	wire _w3734_ ;
	wire _w3733_ ;
	wire _w3732_ ;
	wire _w3731_ ;
	wire _w3730_ ;
	wire _w3729_ ;
	wire _w3728_ ;
	wire _w3727_ ;
	wire _w3726_ ;
	wire _w3725_ ;
	wire _w3724_ ;
	wire _w3723_ ;
	wire _w3722_ ;
	wire _w3721_ ;
	wire _w3720_ ;
	wire _w3719_ ;
	wire _w3718_ ;
	wire _w3717_ ;
	wire _w3716_ ;
	wire _w3715_ ;
	wire _w3714_ ;
	wire _w3713_ ;
	wire _w3712_ ;
	wire _w3711_ ;
	wire _w3710_ ;
	wire _w3709_ ;
	wire _w3708_ ;
	wire _w3707_ ;
	wire _w3706_ ;
	wire _w3705_ ;
	wire _w3704_ ;
	wire _w3703_ ;
	wire _w3702_ ;
	wire _w3701_ ;
	wire _w3700_ ;
	wire _w3699_ ;
	wire _w3698_ ;
	wire _w3697_ ;
	wire _w3696_ ;
	wire _w3695_ ;
	wire _w3694_ ;
	wire _w3693_ ;
	wire _w3692_ ;
	wire _w3691_ ;
	wire _w3690_ ;
	wire _w3689_ ;
	wire _w3688_ ;
	wire _w3687_ ;
	wire _w3686_ ;
	wire _w3685_ ;
	wire _w3684_ ;
	wire _w3683_ ;
	wire _w3682_ ;
	wire _w3681_ ;
	wire _w3680_ ;
	wire _w3679_ ;
	wire _w3678_ ;
	wire _w3677_ ;
	wire _w3676_ ;
	wire _w3675_ ;
	wire _w3674_ ;
	wire _w3673_ ;
	wire _w3672_ ;
	wire _w3671_ ;
	wire _w3670_ ;
	wire _w3669_ ;
	wire _w3668_ ;
	wire _w3667_ ;
	wire _w3666_ ;
	wire _w3665_ ;
	wire _w3664_ ;
	wire _w3663_ ;
	wire _w3662_ ;
	wire _w3661_ ;
	wire _w3660_ ;
	wire _w3659_ ;
	wire _w3658_ ;
	wire _w3657_ ;
	wire _w3656_ ;
	wire _w3655_ ;
	wire _w3654_ ;
	wire _w3653_ ;
	wire _w3652_ ;
	wire _w3651_ ;
	wire _w3650_ ;
	wire _w3649_ ;
	wire _w3648_ ;
	wire _w3647_ ;
	wire _w3646_ ;
	wire _w3645_ ;
	wire _w3644_ ;
	wire _w3643_ ;
	wire _w3642_ ;
	wire _w3641_ ;
	wire _w3640_ ;
	wire _w3639_ ;
	wire _w3638_ ;
	wire _w3637_ ;
	wire _w3636_ ;
	wire _w3635_ ;
	wire _w3634_ ;
	wire _w3633_ ;
	wire _w3632_ ;
	wire _w3631_ ;
	wire _w3630_ ;
	wire _w3629_ ;
	wire _w3628_ ;
	wire _w3627_ ;
	wire _w3626_ ;
	wire _w3625_ ;
	wire _w3624_ ;
	wire _w3623_ ;
	wire _w3622_ ;
	wire _w3621_ ;
	wire _w3620_ ;
	wire _w3619_ ;
	wire _w3618_ ;
	wire _w3617_ ;
	wire _w3616_ ;
	wire _w3615_ ;
	wire _w3614_ ;
	wire _w3613_ ;
	wire _w3612_ ;
	wire _w3611_ ;
	wire _w3610_ ;
	wire _w3609_ ;
	wire _w3608_ ;
	wire _w3607_ ;
	wire _w3606_ ;
	wire _w3605_ ;
	wire _w3604_ ;
	wire _w3603_ ;
	wire _w3602_ ;
	wire _w3601_ ;
	wire _w3600_ ;
	wire _w3599_ ;
	wire _w3598_ ;
	wire _w3597_ ;
	wire _w3596_ ;
	wire _w3595_ ;
	wire _w3594_ ;
	wire _w3593_ ;
	wire _w3592_ ;
	wire _w3591_ ;
	wire _w3590_ ;
	wire _w3589_ ;
	wire _w3588_ ;
	wire _w3587_ ;
	wire _w3586_ ;
	wire _w3585_ ;
	wire _w3584_ ;
	wire _w3583_ ;
	wire _w3582_ ;
	wire _w3581_ ;
	wire _w3580_ ;
	wire _w3579_ ;
	wire _w3578_ ;
	wire _w3577_ ;
	wire _w3576_ ;
	wire _w3575_ ;
	wire _w3574_ ;
	wire _w3573_ ;
	wire _w3572_ ;
	wire _w3571_ ;
	wire _w3570_ ;
	wire _w3569_ ;
	wire _w3568_ ;
	wire _w3567_ ;
	wire _w3566_ ;
	wire _w3565_ ;
	wire _w3564_ ;
	wire _w3563_ ;
	wire _w3562_ ;
	wire _w3561_ ;
	wire _w3560_ ;
	wire _w3559_ ;
	wire _w3558_ ;
	wire _w3557_ ;
	wire _w3556_ ;
	wire _w3555_ ;
	wire _w3554_ ;
	wire _w3553_ ;
	wire _w3552_ ;
	wire _w3551_ ;
	wire _w3550_ ;
	wire _w3549_ ;
	wire _w3548_ ;
	wire _w3547_ ;
	wire _w3546_ ;
	wire _w3545_ ;
	wire _w3544_ ;
	wire _w3543_ ;
	wire _w3542_ ;
	wire _w3541_ ;
	wire _w3540_ ;
	wire _w3539_ ;
	wire _w3538_ ;
	wire _w3537_ ;
	wire _w3536_ ;
	wire _w3535_ ;
	wire _w3534_ ;
	wire _w3533_ ;
	wire _w3532_ ;
	wire _w3531_ ;
	wire _w3530_ ;
	wire _w3529_ ;
	wire _w3528_ ;
	wire _w3527_ ;
	wire _w3526_ ;
	wire _w3525_ ;
	wire _w3524_ ;
	wire _w3523_ ;
	wire _w3522_ ;
	wire _w3521_ ;
	wire _w3520_ ;
	wire _w3519_ ;
	wire _w3518_ ;
	wire _w3517_ ;
	wire _w3516_ ;
	wire _w3515_ ;
	wire _w3514_ ;
	wire _w3513_ ;
	wire _w3512_ ;
	wire _w3511_ ;
	wire _w3510_ ;
	wire _w3509_ ;
	wire _w3508_ ;
	wire _w3507_ ;
	wire _w3506_ ;
	wire _w3505_ ;
	wire _w3504_ ;
	wire _w3503_ ;
	wire _w3502_ ;
	wire _w3501_ ;
	wire _w3500_ ;
	wire _w3499_ ;
	wire _w3498_ ;
	wire _w3497_ ;
	wire _w3496_ ;
	wire _w3495_ ;
	wire _w3494_ ;
	wire _w3493_ ;
	wire _w3492_ ;
	wire _w3491_ ;
	wire _w3490_ ;
	wire _w3489_ ;
	wire _w3488_ ;
	wire _w3487_ ;
	wire _w3486_ ;
	wire _w3485_ ;
	wire _w3484_ ;
	wire _w3483_ ;
	wire _w3482_ ;
	wire _w3481_ ;
	wire _w3480_ ;
	wire _w3479_ ;
	wire _w3478_ ;
	wire _w3477_ ;
	wire _w3476_ ;
	wire _w3475_ ;
	wire _w3474_ ;
	wire _w3473_ ;
	wire _w3472_ ;
	wire _w3471_ ;
	wire _w3470_ ;
	wire _w3469_ ;
	wire _w3468_ ;
	wire _w3467_ ;
	wire _w3466_ ;
	wire _w3465_ ;
	wire _w3464_ ;
	wire _w3463_ ;
	wire _w3462_ ;
	wire _w3461_ ;
	wire _w3460_ ;
	wire _w3459_ ;
	wire _w3458_ ;
	wire _w3457_ ;
	wire _w3456_ ;
	wire _w3455_ ;
	wire _w3454_ ;
	wire _w3453_ ;
	wire _w3452_ ;
	wire _w3451_ ;
	wire _w3450_ ;
	wire _w3449_ ;
	wire _w3448_ ;
	wire _w3447_ ;
	wire _w3446_ ;
	wire _w3445_ ;
	wire _w3444_ ;
	wire _w3443_ ;
	wire _w3442_ ;
	wire _w3441_ ;
	wire _w3440_ ;
	wire _w3439_ ;
	wire _w3438_ ;
	wire _w3437_ ;
	wire _w3436_ ;
	wire _w3435_ ;
	wire _w3434_ ;
	wire _w3433_ ;
	wire _w3432_ ;
	wire _w3431_ ;
	wire _w3430_ ;
	wire _w3429_ ;
	wire _w3428_ ;
	wire _w3427_ ;
	wire _w3426_ ;
	wire _w3425_ ;
	wire _w3424_ ;
	wire _w3423_ ;
	wire _w3422_ ;
	wire _w3421_ ;
	wire _w3420_ ;
	wire _w3419_ ;
	wire _w3418_ ;
	wire _w3417_ ;
	wire _w3416_ ;
	wire _w3415_ ;
	wire _w3414_ ;
	wire _w3413_ ;
	wire _w3412_ ;
	wire _w3411_ ;
	wire _w3410_ ;
	wire _w3409_ ;
	wire _w3408_ ;
	wire _w3407_ ;
	wire _w3406_ ;
	wire _w3405_ ;
	wire _w3404_ ;
	wire _w3403_ ;
	wire _w3402_ ;
	wire _w3401_ ;
	wire _w3400_ ;
	wire _w3399_ ;
	wire _w3398_ ;
	wire _w3397_ ;
	wire _w3396_ ;
	wire _w3395_ ;
	wire _w3394_ ;
	wire _w3393_ ;
	wire _w3392_ ;
	wire _w3391_ ;
	wire _w3390_ ;
	wire _w3389_ ;
	wire _w3388_ ;
	wire _w3387_ ;
	wire _w3386_ ;
	wire _w3385_ ;
	wire _w3384_ ;
	wire _w3383_ ;
	wire _w3382_ ;
	wire _w3381_ ;
	wire _w3380_ ;
	wire _w3379_ ;
	wire _w3378_ ;
	wire _w3377_ ;
	wire _w3376_ ;
	wire _w3375_ ;
	wire _w3374_ ;
	wire _w3373_ ;
	wire _w3372_ ;
	wire _w3371_ ;
	wire _w3370_ ;
	wire _w3369_ ;
	wire _w3368_ ;
	wire _w3367_ ;
	wire _w3366_ ;
	wire _w3365_ ;
	wire _w3364_ ;
	wire _w3363_ ;
	wire _w3362_ ;
	wire _w3361_ ;
	wire _w3360_ ;
	wire _w3359_ ;
	wire _w3358_ ;
	wire _w3357_ ;
	wire _w3356_ ;
	wire _w3355_ ;
	wire _w3354_ ;
	wire _w3353_ ;
	wire _w3352_ ;
	wire _w3351_ ;
	wire _w3350_ ;
	wire _w3349_ ;
	wire _w3348_ ;
	wire _w3347_ ;
	wire _w3346_ ;
	wire _w3345_ ;
	wire _w3344_ ;
	wire _w3343_ ;
	wire _w3342_ ;
	wire _w3341_ ;
	wire _w3340_ ;
	wire _w3339_ ;
	wire _w3338_ ;
	wire _w3337_ ;
	wire _w3336_ ;
	wire _w3335_ ;
	wire _w3334_ ;
	wire _w3333_ ;
	wire _w3332_ ;
	wire _w3331_ ;
	wire _w3330_ ;
	wire _w3329_ ;
	wire _w3328_ ;
	wire _w3327_ ;
	wire _w3326_ ;
	wire _w3325_ ;
	wire _w3324_ ;
	wire _w3323_ ;
	wire _w3322_ ;
	wire _w3321_ ;
	wire _w3320_ ;
	wire _w3319_ ;
	wire _w3318_ ;
	wire _w3317_ ;
	wire _w3316_ ;
	wire _w3315_ ;
	wire _w3314_ ;
	wire _w3313_ ;
	wire _w3312_ ;
	wire _w3311_ ;
	wire _w3310_ ;
	wire _w3309_ ;
	wire _w3308_ ;
	wire _w3307_ ;
	wire _w3306_ ;
	wire _w3305_ ;
	wire _w3304_ ;
	wire _w3303_ ;
	wire _w3302_ ;
	wire _w3301_ ;
	wire _w3300_ ;
	wire _w3299_ ;
	wire _w3298_ ;
	wire _w3297_ ;
	wire _w3296_ ;
	wire _w3295_ ;
	wire _w3294_ ;
	wire _w3293_ ;
	wire _w3292_ ;
	wire _w3291_ ;
	wire _w3290_ ;
	wire _w3289_ ;
	wire _w3288_ ;
	wire _w3287_ ;
	wire _w3286_ ;
	wire _w3285_ ;
	wire _w3284_ ;
	wire _w3283_ ;
	wire _w3282_ ;
	wire _w3281_ ;
	wire _w3280_ ;
	wire _w3279_ ;
	wire _w3278_ ;
	wire _w3277_ ;
	wire _w3276_ ;
	wire _w3275_ ;
	wire _w3274_ ;
	wire _w3273_ ;
	wire _w3272_ ;
	wire _w3271_ ;
	wire _w3270_ ;
	wire _w3269_ ;
	wire _w3268_ ;
	wire _w3267_ ;
	wire _w3266_ ;
	wire _w3265_ ;
	wire _w3264_ ;
	wire _w3263_ ;
	wire _w3262_ ;
	wire _w3261_ ;
	wire _w3260_ ;
	wire _w3259_ ;
	wire _w3258_ ;
	wire _w3257_ ;
	wire _w3256_ ;
	wire _w3255_ ;
	wire _w3254_ ;
	wire _w3253_ ;
	wire _w3252_ ;
	wire _w3251_ ;
	wire _w3250_ ;
	wire _w3249_ ;
	wire _w3248_ ;
	wire _w3247_ ;
	wire _w3246_ ;
	wire _w3245_ ;
	wire _w3244_ ;
	wire _w3243_ ;
	wire _w3242_ ;
	wire _w3241_ ;
	wire _w3240_ ;
	wire _w3239_ ;
	wire _w3238_ ;
	wire _w3237_ ;
	wire _w3236_ ;
	wire _w3235_ ;
	wire _w3234_ ;
	wire _w3233_ ;
	wire _w3232_ ;
	wire _w3231_ ;
	wire _w3230_ ;
	wire _w3229_ ;
	wire _w3228_ ;
	wire _w3227_ ;
	wire _w3226_ ;
	wire _w3225_ ;
	wire _w3224_ ;
	wire _w3223_ ;
	wire _w3222_ ;
	wire _w3221_ ;
	wire _w3220_ ;
	wire _w3219_ ;
	wire _w3218_ ;
	wire _w3217_ ;
	wire _w3216_ ;
	wire _w3215_ ;
	wire _w3214_ ;
	wire _w3213_ ;
	wire _w3212_ ;
	wire _w3211_ ;
	wire _w3210_ ;
	wire _w3209_ ;
	wire _w3208_ ;
	wire _w3207_ ;
	wire _w3206_ ;
	wire _w3205_ ;
	wire _w3204_ ;
	wire _w3203_ ;
	wire _w3202_ ;
	wire _w3201_ ;
	wire _w3200_ ;
	wire _w3199_ ;
	wire _w3198_ ;
	wire _w3197_ ;
	wire _w3196_ ;
	wire _w3195_ ;
	wire _w3194_ ;
	wire _w3193_ ;
	wire _w3192_ ;
	wire _w3191_ ;
	wire _w3190_ ;
	wire _w3189_ ;
	wire _w3188_ ;
	wire _w3187_ ;
	wire _w3186_ ;
	wire _w3185_ ;
	wire _w3184_ ;
	wire _w3183_ ;
	wire _w3182_ ;
	wire _w3181_ ;
	wire _w3180_ ;
	wire _w3179_ ;
	wire _w3178_ ;
	wire _w3177_ ;
	wire _w3176_ ;
	wire _w3175_ ;
	wire _w3174_ ;
	wire _w3173_ ;
	wire _w3172_ ;
	wire _w3171_ ;
	wire _w3170_ ;
	wire _w3169_ ;
	wire _w3168_ ;
	wire _w3167_ ;
	wire _w3166_ ;
	wire _w3165_ ;
	wire _w3164_ ;
	wire _w3163_ ;
	wire _w3162_ ;
	wire _w3161_ ;
	wire _w3160_ ;
	wire _w3159_ ;
	wire _w3158_ ;
	wire _w3157_ ;
	wire _w3156_ ;
	wire _w3155_ ;
	wire _w3154_ ;
	wire _w3153_ ;
	wire _w3152_ ;
	wire _w3151_ ;
	wire _w3150_ ;
	wire _w3149_ ;
	wire _w3148_ ;
	wire _w3147_ ;
	wire _w3146_ ;
	wire _w3145_ ;
	wire _w3144_ ;
	wire _w3143_ ;
	wire _w3142_ ;
	wire _w3141_ ;
	wire _w3140_ ;
	wire _w3139_ ;
	wire _w3138_ ;
	wire _w3137_ ;
	wire _w3136_ ;
	wire _w3135_ ;
	wire _w3134_ ;
	wire _w3133_ ;
	wire _w3132_ ;
	wire _w3131_ ;
	wire _w3130_ ;
	wire _w3129_ ;
	wire _w3128_ ;
	wire _w3127_ ;
	wire _w3126_ ;
	wire _w3125_ ;
	wire _w3124_ ;
	wire _w3123_ ;
	wire _w3122_ ;
	wire _w3121_ ;
	wire _w3120_ ;
	wire _w3119_ ;
	wire _w3118_ ;
	wire _w3117_ ;
	wire _w3116_ ;
	wire _w3115_ ;
	wire _w3114_ ;
	wire _w3113_ ;
	wire _w3112_ ;
	wire _w3111_ ;
	wire _w3110_ ;
	wire _w3109_ ;
	wire _w3108_ ;
	wire _w3107_ ;
	wire _w3106_ ;
	wire _w3105_ ;
	wire _w3104_ ;
	wire _w3103_ ;
	wire _w3102_ ;
	wire _w3101_ ;
	wire _w3100_ ;
	wire _w3099_ ;
	wire _w3098_ ;
	wire _w3097_ ;
	wire _w3096_ ;
	wire _w3095_ ;
	wire _w3094_ ;
	wire _w3093_ ;
	wire _w3092_ ;
	wire _w3091_ ;
	wire _w3090_ ;
	wire _w3089_ ;
	wire _w3088_ ;
	wire _w3087_ ;
	wire _w3086_ ;
	wire _w3085_ ;
	wire _w3084_ ;
	wire _w3083_ ;
	wire _w3082_ ;
	wire _w3081_ ;
	wire _w3080_ ;
	wire _w3079_ ;
	wire _w3078_ ;
	wire _w3077_ ;
	wire _w3076_ ;
	wire _w3075_ ;
	wire _w3074_ ;
	wire _w3073_ ;
	wire _w3072_ ;
	wire _w3071_ ;
	wire _w3070_ ;
	wire _w3069_ ;
	wire _w3068_ ;
	wire _w3067_ ;
	wire _w3066_ ;
	wire _w3065_ ;
	wire _w3064_ ;
	wire _w3063_ ;
	wire _w3062_ ;
	wire _w3061_ ;
	wire _w3060_ ;
	wire _w3059_ ;
	wire _w3058_ ;
	wire _w3057_ ;
	wire _w3056_ ;
	wire _w3055_ ;
	wire _w3054_ ;
	wire _w3053_ ;
	wire _w3052_ ;
	wire _w3051_ ;
	wire _w3050_ ;
	wire _w3049_ ;
	wire _w3048_ ;
	wire _w3047_ ;
	wire _w3046_ ;
	wire _w3045_ ;
	wire _w3044_ ;
	wire _w3043_ ;
	wire _w3042_ ;
	wire _w3041_ ;
	wire _w3040_ ;
	wire _w3039_ ;
	wire _w3038_ ;
	wire _w3037_ ;
	wire _w3036_ ;
	wire _w3035_ ;
	wire _w3034_ ;
	wire _w3033_ ;
	wire _w3032_ ;
	wire _w3031_ ;
	wire _w3030_ ;
	wire _w3029_ ;
	wire _w3028_ ;
	wire _w3027_ ;
	wire _w3026_ ;
	wire _w3025_ ;
	wire _w3024_ ;
	wire _w3023_ ;
	wire _w3022_ ;
	wire _w3021_ ;
	wire _w3020_ ;
	wire _w3019_ ;
	wire _w3018_ ;
	wire _w3017_ ;
	wire _w3016_ ;
	wire _w3015_ ;
	wire _w3014_ ;
	wire _w3013_ ;
	wire _w3012_ ;
	wire _w3011_ ;
	wire _w3010_ ;
	wire _w3009_ ;
	wire _w3008_ ;
	wire _w3007_ ;
	wire _w3006_ ;
	wire _w3005_ ;
	wire _w3004_ ;
	wire _w3003_ ;
	wire _w3002_ ;
	wire _w3001_ ;
	wire _w3000_ ;
	wire _w2999_ ;
	wire _w2998_ ;
	wire _w2997_ ;
	wire _w2996_ ;
	wire _w2995_ ;
	wire _w2994_ ;
	wire _w2993_ ;
	wire _w2992_ ;
	wire _w2991_ ;
	wire _w2990_ ;
	wire _w2989_ ;
	wire _w2988_ ;
	wire _w2987_ ;
	wire _w2986_ ;
	wire _w2985_ ;
	wire _w2984_ ;
	wire _w2983_ ;
	wire _w2982_ ;
	wire _w2981_ ;
	wire _w2980_ ;
	wire _w2979_ ;
	wire _w2978_ ;
	wire _w2977_ ;
	wire _w2976_ ;
	wire _w2975_ ;
	wire _w2974_ ;
	wire _w2973_ ;
	wire _w2972_ ;
	wire _w2971_ ;
	wire _w2970_ ;
	wire _w2969_ ;
	wire _w2968_ ;
	wire _w2967_ ;
	wire _w2966_ ;
	wire _w2965_ ;
	wire _w2964_ ;
	wire _w2963_ ;
	wire _w2962_ ;
	wire _w2961_ ;
	wire _w2960_ ;
	wire _w2959_ ;
	wire _w2958_ ;
	wire _w2957_ ;
	wire _w2956_ ;
	wire _w2955_ ;
	wire _w2954_ ;
	wire _w2953_ ;
	wire _w2952_ ;
	wire _w2951_ ;
	wire _w2950_ ;
	wire _w2949_ ;
	wire _w2948_ ;
	wire _w2947_ ;
	wire _w2946_ ;
	wire _w2945_ ;
	wire _w2944_ ;
	wire _w2943_ ;
	wire _w2942_ ;
	wire _w2941_ ;
	wire _w2940_ ;
	wire _w2939_ ;
	wire _w2938_ ;
	wire _w2937_ ;
	wire _w2936_ ;
	wire _w2935_ ;
	wire _w2934_ ;
	wire _w2933_ ;
	wire _w2932_ ;
	wire _w2931_ ;
	wire _w2930_ ;
	wire _w2929_ ;
	wire _w2928_ ;
	wire _w2927_ ;
	wire _w2926_ ;
	wire _w2925_ ;
	wire _w2924_ ;
	wire _w2923_ ;
	wire _w2922_ ;
	wire _w2921_ ;
	wire _w2920_ ;
	wire _w2919_ ;
	wire _w2918_ ;
	wire _w2917_ ;
	wire _w2916_ ;
	wire _w2915_ ;
	wire _w2914_ ;
	wire _w2913_ ;
	wire _w2912_ ;
	wire _w2911_ ;
	wire _w2910_ ;
	wire _w2909_ ;
	wire _w2908_ ;
	wire _w2907_ ;
	wire _w2906_ ;
	wire _w2905_ ;
	wire _w2904_ ;
	wire _w2903_ ;
	wire _w2902_ ;
	wire _w2901_ ;
	wire _w2900_ ;
	wire _w2899_ ;
	wire _w2898_ ;
	wire _w2897_ ;
	wire _w2896_ ;
	wire _w2895_ ;
	wire _w2894_ ;
	wire _w2893_ ;
	wire _w2892_ ;
	wire _w2891_ ;
	wire _w2890_ ;
	wire _w2889_ ;
	wire _w2888_ ;
	wire _w2887_ ;
	wire _w2886_ ;
	wire _w2885_ ;
	wire _w2884_ ;
	wire _w2883_ ;
	wire _w2882_ ;
	wire _w2881_ ;
	wire _w2880_ ;
	wire _w2879_ ;
	wire _w2878_ ;
	wire _w2877_ ;
	wire _w2876_ ;
	wire _w2875_ ;
	wire _w2874_ ;
	wire _w2873_ ;
	wire _w2872_ ;
	wire _w2871_ ;
	wire _w2870_ ;
	wire _w2869_ ;
	wire _w2868_ ;
	wire _w2867_ ;
	wire _w2866_ ;
	wire _w2865_ ;
	wire _w2864_ ;
	wire _w2863_ ;
	wire _w2862_ ;
	wire _w2861_ ;
	wire _w2860_ ;
	wire _w2859_ ;
	wire _w2858_ ;
	wire _w2857_ ;
	wire _w2856_ ;
	wire _w2855_ ;
	wire _w2854_ ;
	wire _w2853_ ;
	wire _w2852_ ;
	wire _w2851_ ;
	wire _w2850_ ;
	wire _w2849_ ;
	wire _w2848_ ;
	wire _w2847_ ;
	wire _w2846_ ;
	wire _w2845_ ;
	wire _w2844_ ;
	wire _w2843_ ;
	wire _w2842_ ;
	wire _w2841_ ;
	wire _w2840_ ;
	wire _w2839_ ;
	wire _w2838_ ;
	wire _w2837_ ;
	wire _w2836_ ;
	wire _w2835_ ;
	wire _w2834_ ;
	wire _w2833_ ;
	wire _w2832_ ;
	wire _w2831_ ;
	wire _w2830_ ;
	wire _w2829_ ;
	wire _w2828_ ;
	wire _w2827_ ;
	wire _w2826_ ;
	wire _w2825_ ;
	wire _w2824_ ;
	wire _w2823_ ;
	wire _w2822_ ;
	wire _w2821_ ;
	wire _w2820_ ;
	wire _w2819_ ;
	wire _w2818_ ;
	wire _w2817_ ;
	wire _w2816_ ;
	wire _w2815_ ;
	wire _w2814_ ;
	wire _w2813_ ;
	wire _w2812_ ;
	wire _w2811_ ;
	wire _w2810_ ;
	wire _w1561_ ;
	wire _w1560_ ;
	wire _w1559_ ;
	wire _w1558_ ;
	wire _w1557_ ;
	wire _w1556_ ;
	wire _w1555_ ;
	wire _w1554_ ;
	wire _w1553_ ;
	wire _w1552_ ;
	wire _w1551_ ;
	wire _w1550_ ;
	wire _w1549_ ;
	wire _w1548_ ;
	wire _w1547_ ;
	wire _w1546_ ;
	wire _w1545_ ;
	wire _w1544_ ;
	wire _w1543_ ;
	wire _w1542_ ;
	wire _w1541_ ;
	wire _w1540_ ;
	wire _w1539_ ;
	wire _w1538_ ;
	wire _w1537_ ;
	wire _w1536_ ;
	wire _w1535_ ;
	wire _w1534_ ;
	wire _w1533_ ;
	wire _w1532_ ;
	wire _w1531_ ;
	wire _w1530_ ;
	wire _w1529_ ;
	wire _w1528_ ;
	wire _w1527_ ;
	wire _w1526_ ;
	wire _w1525_ ;
	wire _w1524_ ;
	wire _w1523_ ;
	wire _w1522_ ;
	wire _w1521_ ;
	wire _w1520_ ;
	wire _w1519_ ;
	wire _w1518_ ;
	wire _w1517_ ;
	wire _w1516_ ;
	wire _w1515_ ;
	wire _w1514_ ;
	wire _w1513_ ;
	wire _w1512_ ;
	wire _w1511_ ;
	wire _w1510_ ;
	wire _w1509_ ;
	wire _w1508_ ;
	wire _w1507_ ;
	wire _w1506_ ;
	wire _w1505_ ;
	wire _w1504_ ;
	wire _w1503_ ;
	wire _w1502_ ;
	wire _w1501_ ;
	wire _w1500_ ;
	wire _w1499_ ;
	wire _w1498_ ;
	wire _w1497_ ;
	wire _w1496_ ;
	wire _w1495_ ;
	wire _w1494_ ;
	wire _w1493_ ;
	wire _w1492_ ;
	wire _w1491_ ;
	wire _w1490_ ;
	wire _w1489_ ;
	wire _w1488_ ;
	wire _w1487_ ;
	wire _w1486_ ;
	wire _w1485_ ;
	wire _w1484_ ;
	wire _w1483_ ;
	wire _w1482_ ;
	wire _w1481_ ;
	wire _w1480_ ;
	wire _w1479_ ;
	wire _w1478_ ;
	wire _w1477_ ;
	wire _w1476_ ;
	wire _w1475_ ;
	wire _w1474_ ;
	wire _w1473_ ;
	wire _w1472_ ;
	wire _w1471_ ;
	wire _w1470_ ;
	wire _w1469_ ;
	wire _w1468_ ;
	wire _w1467_ ;
	wire _w1466_ ;
	wire _w1465_ ;
	wire _w1464_ ;
	wire _w1463_ ;
	wire _w1462_ ;
	wire _w1461_ ;
	wire _w1460_ ;
	wire _w1459_ ;
	wire _w1458_ ;
	wire _w1457_ ;
	wire _w1456_ ;
	wire _w1455_ ;
	wire _w1454_ ;
	wire _w1453_ ;
	wire _w1452_ ;
	wire _w1451_ ;
	wire _w1450_ ;
	wire _w1449_ ;
	wire _w1448_ ;
	wire _w1447_ ;
	wire _w1446_ ;
	wire _w1445_ ;
	wire _w1444_ ;
	wire _w1443_ ;
	wire _w1442_ ;
	wire _w1441_ ;
	wire _w1440_ ;
	wire _w1439_ ;
	wire _w1438_ ;
	wire _w1437_ ;
	wire _w1436_ ;
	wire _w1435_ ;
	wire _w1434_ ;
	wire _w1433_ ;
	wire _w1432_ ;
	wire _w1431_ ;
	wire _w1430_ ;
	wire _w1429_ ;
	wire _w1428_ ;
	wire _w1427_ ;
	wire _w1426_ ;
	wire _w1425_ ;
	wire _w1424_ ;
	wire _w1423_ ;
	wire _w1422_ ;
	wire _w1421_ ;
	wire _w1420_ ;
	wire _w1419_ ;
	wire _w1418_ ;
	wire _w1417_ ;
	wire _w1416_ ;
	wire _w1415_ ;
	wire _w1414_ ;
	wire _w1413_ ;
	wire _w1412_ ;
	wire _w1411_ ;
	wire _w1410_ ;
	wire _w1409_ ;
	wire _w1408_ ;
	wire _w1407_ ;
	wire _w1406_ ;
	wire _w1405_ ;
	wire _w1404_ ;
	wire _w1403_ ;
	wire _w1402_ ;
	wire _w1401_ ;
	wire _w1400_ ;
	wire _w1399_ ;
	wire _w1398_ ;
	wire _w1397_ ;
	wire _w1396_ ;
	wire _w1395_ ;
	wire _w1394_ ;
	wire _w1393_ ;
	wire _w1392_ ;
	wire _w1391_ ;
	wire _w1390_ ;
	wire _w1389_ ;
	wire _w1388_ ;
	wire _w1387_ ;
	wire _w1386_ ;
	wire _w1385_ ;
	wire _w1384_ ;
	wire _w1383_ ;
	wire _w1382_ ;
	wire _w1381_ ;
	wire _w1380_ ;
	wire _w1379_ ;
	wire _w1378_ ;
	wire _w1377_ ;
	wire _w1376_ ;
	wire _w1375_ ;
	wire _w1374_ ;
	wire _w1373_ ;
	wire _w1372_ ;
	wire _w1371_ ;
	wire _w1370_ ;
	wire _w1369_ ;
	wire _w1368_ ;
	wire _w1367_ ;
	wire _w1366_ ;
	wire _w1365_ ;
	wire _w1364_ ;
	wire _w1363_ ;
	wire _w1362_ ;
	wire _w1361_ ;
	wire _w1360_ ;
	wire _w1359_ ;
	wire _w1358_ ;
	wire _w1357_ ;
	wire _w1356_ ;
	wire _w1355_ ;
	wire _w1354_ ;
	wire _w1353_ ;
	wire _w1352_ ;
	wire _w1351_ ;
	wire _w1350_ ;
	wire _w1349_ ;
	wire _w1348_ ;
	wire _w1347_ ;
	wire _w1346_ ;
	wire _w1345_ ;
	wire _w1344_ ;
	wire _w1343_ ;
	wire _w1342_ ;
	wire _w1341_ ;
	wire _w1340_ ;
	wire _w1339_ ;
	wire _w1338_ ;
	wire _w1337_ ;
	wire _w1336_ ;
	wire _w1335_ ;
	wire _w1334_ ;
	wire _w1333_ ;
	wire _w1332_ ;
	wire _w1331_ ;
	wire _w1330_ ;
	wire _w1329_ ;
	wire _w1328_ ;
	wire _w1327_ ;
	wire _w1326_ ;
	wire _w1325_ ;
	wire _w1324_ ;
	wire _w1323_ ;
	wire _w1322_ ;
	wire _w1321_ ;
	wire _w1320_ ;
	wire _w1319_ ;
	wire _w1318_ ;
	wire _w1317_ ;
	wire _w1316_ ;
	wire _w1315_ ;
	wire _w1314_ ;
	wire _w1313_ ;
	wire _w1312_ ;
	wire _w1311_ ;
	wire _w1310_ ;
	wire _w1309_ ;
	wire _w1308_ ;
	wire _w1307_ ;
	wire _w1306_ ;
	wire _w1305_ ;
	wire _w1304_ ;
	wire _w1303_ ;
	wire _w1302_ ;
	wire _w1301_ ;
	wire _w1300_ ;
	wire _w1299_ ;
	wire _w1298_ ;
	wire _w1297_ ;
	wire _w1296_ ;
	wire _w1295_ ;
	wire _w1294_ ;
	wire _w1293_ ;
	wire _w1292_ ;
	wire _w1291_ ;
	wire _w1290_ ;
	wire _w1289_ ;
	wire _w1288_ ;
	wire _w1287_ ;
	wire _w1286_ ;
	wire _w1285_ ;
	wire _w1284_ ;
	wire _w1283_ ;
	wire _w1282_ ;
	wire _w1281_ ;
	wire _w1280_ ;
	wire _w1279_ ;
	wire _w1278_ ;
	wire _w1277_ ;
	wire _w1276_ ;
	wire _w1275_ ;
	wire _w1274_ ;
	wire _w1273_ ;
	wire _w1272_ ;
	wire _w1271_ ;
	wire _w1270_ ;
	wire _w1269_ ;
	wire _w1268_ ;
	wire _w1267_ ;
	wire _w1266_ ;
	wire _w1265_ ;
	wire _w1264_ ;
	wire _w1263_ ;
	wire _w1262_ ;
	wire _w1261_ ;
	wire _w1260_ ;
	wire _w1259_ ;
	wire _w1258_ ;
	wire _w1257_ ;
	wire _w1256_ ;
	wire _w1255_ ;
	wire _w1254_ ;
	wire _w1253_ ;
	wire _w1252_ ;
	wire _w1251_ ;
	wire _w1250_ ;
	wire _w1249_ ;
	wire _w1248_ ;
	wire _w1247_ ;
	wire _w1246_ ;
	wire _w1245_ ;
	wire _w1244_ ;
	wire _w1243_ ;
	wire _w1242_ ;
	wire _w1241_ ;
	wire _w1240_ ;
	wire _w1239_ ;
	wire _w1238_ ;
	wire _w1237_ ;
	wire _w1236_ ;
	wire _w1235_ ;
	wire _w1234_ ;
	wire _w1233_ ;
	wire _w1232_ ;
	wire _w1231_ ;
	wire _w1230_ ;
	wire _w1229_ ;
	wire _w1228_ ;
	wire _w1227_ ;
	wire _w1226_ ;
	wire _w1225_ ;
	wire _w1224_ ;
	wire _w1223_ ;
	wire _w1222_ ;
	wire _w1221_ ;
	wire _w1220_ ;
	wire _w1219_ ;
	wire _w1218_ ;
	wire _w1217_ ;
	wire _w1216_ ;
	wire _w1215_ ;
	wire _w1214_ ;
	wire _w1213_ ;
	wire _w1212_ ;
	wire _w1211_ ;
	wire _w1210_ ;
	wire _w1209_ ;
	wire _w1208_ ;
	wire _w1207_ ;
	wire _w1206_ ;
	wire _w1205_ ;
	wire _w1204_ ;
	wire _w1203_ ;
	wire _w1202_ ;
	wire _w1201_ ;
	wire _w1200_ ;
	wire _w1199_ ;
	wire _w1198_ ;
	wire _w1197_ ;
	wire _w1196_ ;
	wire _w1195_ ;
	wire _w1194_ ;
	wire _w1193_ ;
	wire _w1192_ ;
	wire _w1191_ ;
	wire _w1190_ ;
	wire _w1189_ ;
	wire _w1188_ ;
	wire _w1187_ ;
	wire _w1186_ ;
	wire _w1185_ ;
	wire _w1184_ ;
	wire _w1183_ ;
	wire _w1182_ ;
	wire _w1181_ ;
	wire _w1180_ ;
	wire _w1179_ ;
	wire _w1178_ ;
	wire _w1177_ ;
	wire _w1176_ ;
	wire _w1175_ ;
	wire _w1174_ ;
	wire _w1173_ ;
	wire _w1172_ ;
	wire _w1171_ ;
	wire _w1170_ ;
	wire _w1169_ ;
	wire _w1168_ ;
	wire _w1167_ ;
	wire _w1166_ ;
	wire _w1165_ ;
	wire _w1164_ ;
	wire _w1163_ ;
	wire _w1162_ ;
	wire _w1161_ ;
	wire _w1160_ ;
	wire _w1159_ ;
	wire _w1158_ ;
	wire _w1157_ ;
	wire _w1156_ ;
	wire _w1155_ ;
	wire _w1154_ ;
	wire _w1153_ ;
	wire _w1152_ ;
	wire _w1151_ ;
	wire _w1150_ ;
	wire _w1149_ ;
	wire _w1148_ ;
	wire _w1147_ ;
	wire _w1146_ ;
	wire _w1145_ ;
	wire _w1144_ ;
	wire _w1143_ ;
	wire _w1142_ ;
	wire _w1141_ ;
	wire _w1140_ ;
	wire _w1139_ ;
	wire _w1138_ ;
	wire _w1137_ ;
	wire _w1136_ ;
	wire _w1135_ ;
	wire _w1134_ ;
	wire _w1133_ ;
	wire _w1132_ ;
	wire _w1131_ ;
	wire _w1130_ ;
	wire _w1129_ ;
	wire _w1128_ ;
	wire _w1127_ ;
	wire _w1126_ ;
	wire _w1125_ ;
	wire _w1124_ ;
	wire _w1123_ ;
	wire _w1122_ ;
	wire _w1121_ ;
	wire _w1120_ ;
	wire _w1119_ ;
	wire _w1118_ ;
	wire _w1117_ ;
	wire _w1116_ ;
	wire _w1115_ ;
	wire _w1114_ ;
	wire _w1113_ ;
	wire _w1112_ ;
	wire _w1111_ ;
	wire _w1110_ ;
	wire _w1109_ ;
	wire _w1108_ ;
	wire _w1107_ ;
	wire _w1106_ ;
	wire _w1105_ ;
	wire _w1104_ ;
	wire _w1103_ ;
	wire _w1102_ ;
	wire _w1101_ ;
	wire _w1100_ ;
	wire _w1099_ ;
	wire _w1098_ ;
	wire _w1097_ ;
	wire _w1096_ ;
	wire _w1095_ ;
	wire _w1094_ ;
	wire _w1093_ ;
	wire _w1092_ ;
	wire _w1091_ ;
	wire _w1090_ ;
	wire _w1089_ ;
	wire _w1088_ ;
	wire _w1087_ ;
	wire _w1086_ ;
	wire _w1085_ ;
	wire _w1084_ ;
	wire _w1083_ ;
	wire _w1082_ ;
	wire _w1081_ ;
	wire _w1080_ ;
	wire _w1079_ ;
	wire _w1078_ ;
	wire _w1077_ ;
	wire _w1076_ ;
	wire _w1075_ ;
	wire _w1074_ ;
	wire _w1073_ ;
	wire _w1072_ ;
	wire _w1071_ ;
	wire _w1070_ ;
	wire _w1069_ ;
	wire _w1068_ ;
	wire _w1067_ ;
	wire _w1066_ ;
	wire _w1065_ ;
	wire _w1064_ ;
	wire _w1063_ ;
	wire _w1062_ ;
	wire _w1061_ ;
	wire _w1060_ ;
	wire _w1059_ ;
	wire _w1058_ ;
	wire _w1057_ ;
	wire _w1056_ ;
	wire _w1055_ ;
	wire _w1054_ ;
	wire _w1053_ ;
	wire _w1052_ ;
	wire _w1051_ ;
	wire _w1050_ ;
	wire _w1049_ ;
	wire _w1048_ ;
	wire _w1047_ ;
	wire _w1046_ ;
	wire _w1045_ ;
	wire _w1044_ ;
	wire _w1043_ ;
	wire _w1042_ ;
	wire _w1041_ ;
	wire _w1040_ ;
	wire _w1039_ ;
	wire _w1038_ ;
	wire _w1037_ ;
	wire _w1036_ ;
	wire _w1035_ ;
	wire _w1034_ ;
	wire _w1033_ ;
	wire _w1032_ ;
	wire _w1031_ ;
	wire _w1030_ ;
	wire _w1029_ ;
	wire _w1028_ ;
	wire _w1027_ ;
	wire _w1026_ ;
	wire _w1025_ ;
	wire _w1024_ ;
	wire _w1023_ ;
	wire _w1022_ ;
	wire _w1021_ ;
	wire _w1020_ ;
	wire _w1019_ ;
	wire _w1018_ ;
	wire _w1017_ ;
	wire _w1016_ ;
	wire _w1015_ ;
	wire _w1014_ ;
	wire _w1013_ ;
	wire _w1012_ ;
	wire _w1011_ ;
	wire _w1010_ ;
	wire _w1009_ ;
	wire _w1008_ ;
	wire _w1007_ ;
	wire _w1006_ ;
	wire _w1005_ ;
	wire _w1004_ ;
	wire _w1003_ ;
	wire _w1002_ ;
	wire _w1001_ ;
	wire _w1000_ ;
	wire _w999_ ;
	wire _w998_ ;
	wire _w997_ ;
	wire _w996_ ;
	wire _w995_ ;
	wire _w994_ ;
	wire _w709_ ;
	wire _w708_ ;
	wire _w707_ ;
	wire _w706_ ;
	wire _w705_ ;
	wire _w704_ ;
	wire _w703_ ;
	wire _w702_ ;
	wire _w701_ ;
	wire _w700_ ;
	wire _w699_ ;
	wire _w698_ ;
	wire _w697_ ;
	wire _w696_ ;
	wire _w695_ ;
	wire _w694_ ;
	wire _w693_ ;
	wire _w692_ ;
	wire _w691_ ;
	wire _w690_ ;
	wire _w689_ ;
	wire _w688_ ;
	wire _w687_ ;
	wire _w686_ ;
	wire _w685_ ;
	wire _w684_ ;
	wire _w683_ ;
	wire _w682_ ;
	wire _w681_ ;
	wire _w680_ ;
	wire _w679_ ;
	wire _w678_ ;
	wire _w677_ ;
	wire _w676_ ;
	wire _w675_ ;
	wire _w674_ ;
	wire _w673_ ;
	wire _w672_ ;
	wire _w671_ ;
	wire _w670_ ;
	wire _w669_ ;
	wire _w668_ ;
	wire _w667_ ;
	wire _w666_ ;
	wire _w665_ ;
	wire _w664_ ;
	wire _w663_ ;
	wire _w662_ ;
	wire _w661_ ;
	wire _w660_ ;
	wire _w659_ ;
	wire _w658_ ;
	wire _w657_ ;
	wire _w656_ ;
	wire _w655_ ;
	wire _w654_ ;
	wire _w653_ ;
	wire _w652_ ;
	wire _w651_ ;
	wire _w650_ ;
	wire _w649_ ;
	wire _w648_ ;
	wire _w647_ ;
	wire _w646_ ;
	wire _w645_ ;
	wire _w644_ ;
	wire _w643_ ;
	wire _w642_ ;
	wire _w641_ ;
	wire _w640_ ;
	wire _w639_ ;
	wire _w638_ ;
	wire _w637_ ;
	wire _w636_ ;
	wire _w635_ ;
	wire _w634_ ;
	wire _w633_ ;
	wire _w632_ ;
	wire _w631_ ;
	wire _w630_ ;
	wire _w629_ ;
	wire _w628_ ;
	wire _w627_ ;
	wire _w626_ ;
	wire _w625_ ;
	wire _w624_ ;
	wire _w623_ ;
	wire _w622_ ;
	wire _w621_ ;
	wire _w620_ ;
	wire _w619_ ;
	wire _w618_ ;
	wire _w617_ ;
	wire _w616_ ;
	wire _w615_ ;
	wire _w614_ ;
	wire _w613_ ;
	wire _w612_ ;
	wire _w611_ ;
	wire _w610_ ;
	wire _w609_ ;
	wire _w608_ ;
	wire _w607_ ;
	wire _w606_ ;
	wire _w605_ ;
	wire _w604_ ;
	wire _w603_ ;
	wire _w602_ ;
	wire _w601_ ;
	wire _w600_ ;
	wire _w599_ ;
	wire _w598_ ;
	wire _w597_ ;
	wire _w596_ ;
	wire _w595_ ;
	wire _w594_ ;
	wire _w593_ ;
	wire _w592_ ;
	wire _w591_ ;
	wire _w590_ ;
	wire _w589_ ;
	wire _w588_ ;
	wire _w587_ ;
	wire _w586_ ;
	wire _w585_ ;
	wire _w584_ ;
	wire _w583_ ;
	wire _w582_ ;
	wire _w581_ ;
	wire _w580_ ;
	wire _w511_ ;
	wire _w510_ ;
	wire _w509_ ;
	wire _w508_ ;
	wire _w507_ ;
	wire _w506_ ;
	wire _w505_ ;
	wire _w504_ ;
	wire _w503_ ;
	wire _w502_ ;
	wire _w501_ ;
	wire _w500_ ;
	wire _w499_ ;
	wire _w498_ ;
	wire _w497_ ;
	wire _w496_ ;
	wire _w495_ ;
	wire _w494_ ;
	wire _w493_ ;
	wire _w492_ ;
	wire _w491_ ;
	wire _w490_ ;
	wire _w489_ ;
	wire _w488_ ;
	wire _w487_ ;
	wire _w486_ ;
	wire _w485_ ;
	wire _w484_ ;
	wire _w483_ ;
	wire _w482_ ;
	wire _w465_ ;
	wire _w464_ ;
	wire _w463_ ;
	wire _w462_ ;
	wire _w461_ ;
	wire _w460_ ;
	wire _w459_ ;
	wire _w458_ ;
	wire _w457_ ;
	wire _w456_ ;
	wire _w455_ ;
	wire _w454_ ;
	wire _w453_ ;
	wire _w466_ ;
	wire _w467_ ;
	wire _w468_ ;
	wire _w469_ ;
	wire _w470_ ;
	wire _w471_ ;
	wire _w472_ ;
	wire _w473_ ;
	wire _w474_ ;
	wire _w475_ ;
	wire _w476_ ;
	wire _w477_ ;
	wire _w478_ ;
	wire _w479_ ;
	wire _w480_ ;
	wire _w481_ ;
	wire _w512_ ;
	wire _w513_ ;
	wire _w514_ ;
	wire _w515_ ;
	wire _w516_ ;
	wire _w517_ ;
	wire _w518_ ;
	wire _w519_ ;
	wire _w520_ ;
	wire _w521_ ;
	wire _w522_ ;
	wire _w523_ ;
	wire _w524_ ;
	wire _w525_ ;
	wire _w526_ ;
	wire _w527_ ;
	wire _w528_ ;
	wire _w529_ ;
	wire _w530_ ;
	wire _w531_ ;
	wire _w532_ ;
	wire _w533_ ;
	wire _w534_ ;
	wire _w535_ ;
	wire _w536_ ;
	wire _w537_ ;
	wire _w538_ ;
	wire _w539_ ;
	wire _w540_ ;
	wire _w541_ ;
	wire _w542_ ;
	wire _w543_ ;
	wire _w544_ ;
	wire _w545_ ;
	wire _w546_ ;
	wire _w547_ ;
	wire _w548_ ;
	wire _w549_ ;
	wire _w550_ ;
	wire _w551_ ;
	wire _w552_ ;
	wire _w553_ ;
	wire _w554_ ;
	wire _w555_ ;
	wire _w556_ ;
	wire _w557_ ;
	wire _w558_ ;
	wire _w559_ ;
	wire _w560_ ;
	wire _w561_ ;
	wire _w562_ ;
	wire _w563_ ;
	wire _w564_ ;
	wire _w565_ ;
	wire _w566_ ;
	wire _w567_ ;
	wire _w568_ ;
	wire _w569_ ;
	wire _w570_ ;
	wire _w571_ ;
	wire _w572_ ;
	wire _w573_ ;
	wire _w574_ ;
	wire _w575_ ;
	wire _w576_ ;
	wire _w577_ ;
	wire _w578_ ;
	wire _w579_ ;
	wire _w710_ ;
	wire _w711_ ;
	wire _w712_ ;
	wire _w713_ ;
	wire _w714_ ;
	wire _w715_ ;
	wire _w716_ ;
	wire _w717_ ;
	wire _w718_ ;
	wire _w719_ ;
	wire _w720_ ;
	wire _w721_ ;
	wire _w722_ ;
	wire _w723_ ;
	wire _w724_ ;
	wire _w725_ ;
	wire _w726_ ;
	wire _w727_ ;
	wire _w728_ ;
	wire _w729_ ;
	wire _w730_ ;
	wire _w731_ ;
	wire _w732_ ;
	wire _w733_ ;
	wire _w734_ ;
	wire _w735_ ;
	wire _w736_ ;
	wire _w737_ ;
	wire _w738_ ;
	wire _w739_ ;
	wire _w740_ ;
	wire _w741_ ;
	wire _w742_ ;
	wire _w743_ ;
	wire _w744_ ;
	wire _w745_ ;
	wire _w746_ ;
	wire _w747_ ;
	wire _w748_ ;
	wire _w749_ ;
	wire _w750_ ;
	wire _w751_ ;
	wire _w752_ ;
	wire _w753_ ;
	wire _w754_ ;
	wire _w755_ ;
	wire _w756_ ;
	wire _w757_ ;
	wire _w758_ ;
	wire _w759_ ;
	wire _w760_ ;
	wire _w761_ ;
	wire _w762_ ;
	wire _w763_ ;
	wire _w764_ ;
	wire _w765_ ;
	wire _w766_ ;
	wire _w767_ ;
	wire _w768_ ;
	wire _w769_ ;
	wire _w770_ ;
	wire _w771_ ;
	wire _w772_ ;
	wire _w773_ ;
	wire _w774_ ;
	wire _w775_ ;
	wire _w776_ ;
	wire _w777_ ;
	wire _w778_ ;
	wire _w779_ ;
	wire _w780_ ;
	wire _w781_ ;
	wire _w782_ ;
	wire _w783_ ;
	wire _w784_ ;
	wire _w785_ ;
	wire _w786_ ;
	wire _w787_ ;
	wire _w788_ ;
	wire _w789_ ;
	wire _w790_ ;
	wire _w791_ ;
	wire _w792_ ;
	wire _w793_ ;
	wire _w794_ ;
	wire _w795_ ;
	wire _w796_ ;
	wire _w797_ ;
	wire _w798_ ;
	wire _w799_ ;
	wire _w800_ ;
	wire _w801_ ;
	wire _w802_ ;
	wire _w803_ ;
	wire _w804_ ;
	wire _w805_ ;
	wire _w806_ ;
	wire _w807_ ;
	wire _w808_ ;
	wire _w809_ ;
	wire _w810_ ;
	wire _w811_ ;
	wire _w812_ ;
	wire _w813_ ;
	wire _w814_ ;
	wire _w815_ ;
	wire _w816_ ;
	wire _w817_ ;
	wire _w818_ ;
	wire _w819_ ;
	wire _w820_ ;
	wire _w821_ ;
	wire _w822_ ;
	wire _w823_ ;
	wire _w824_ ;
	wire _w825_ ;
	wire _w826_ ;
	wire _w827_ ;
	wire _w828_ ;
	wire _w829_ ;
	wire _w830_ ;
	wire _w831_ ;
	wire _w832_ ;
	wire _w833_ ;
	wire _w834_ ;
	wire _w835_ ;
	wire _w836_ ;
	wire _w837_ ;
	wire _w838_ ;
	wire _w839_ ;
	wire _w840_ ;
	wire _w841_ ;
	wire _w842_ ;
	wire _w843_ ;
	wire _w844_ ;
	wire _w845_ ;
	wire _w846_ ;
	wire _w847_ ;
	wire _w848_ ;
	wire _w849_ ;
	wire _w850_ ;
	wire _w851_ ;
	wire _w852_ ;
	wire _w853_ ;
	wire _w854_ ;
	wire _w855_ ;
	wire _w856_ ;
	wire _w857_ ;
	wire _w858_ ;
	wire _w859_ ;
	wire _w860_ ;
	wire _w861_ ;
	wire _w862_ ;
	wire _w863_ ;
	wire _w864_ ;
	wire _w865_ ;
	wire _w866_ ;
	wire _w867_ ;
	wire _w868_ ;
	wire _w869_ ;
	wire _w870_ ;
	wire _w871_ ;
	wire _w872_ ;
	wire _w873_ ;
	wire _w874_ ;
	wire _w875_ ;
	wire _w876_ ;
	wire _w877_ ;
	wire _w878_ ;
	wire _w879_ ;
	wire _w880_ ;
	wire _w881_ ;
	wire _w882_ ;
	wire _w883_ ;
	wire _w884_ ;
	wire _w885_ ;
	wire _w886_ ;
	wire _w887_ ;
	wire _w888_ ;
	wire _w889_ ;
	wire _w890_ ;
	wire _w891_ ;
	wire _w892_ ;
	wire _w893_ ;
	wire _w894_ ;
	wire _w895_ ;
	wire _w896_ ;
	wire _w897_ ;
	wire _w898_ ;
	wire _w899_ ;
	wire _w900_ ;
	wire _w901_ ;
	wire _w902_ ;
	wire _w903_ ;
	wire _w904_ ;
	wire _w905_ ;
	wire _w906_ ;
	wire _w907_ ;
	wire _w908_ ;
	wire _w909_ ;
	wire _w910_ ;
	wire _w911_ ;
	wire _w912_ ;
	wire _w913_ ;
	wire _w914_ ;
	wire _w915_ ;
	wire _w916_ ;
	wire _w917_ ;
	wire _w918_ ;
	wire _w919_ ;
	wire _w920_ ;
	wire _w921_ ;
	wire _w922_ ;
	wire _w923_ ;
	wire _w924_ ;
	wire _w925_ ;
	wire _w926_ ;
	wire _w927_ ;
	wire _w928_ ;
	wire _w929_ ;
	wire _w930_ ;
	wire _w931_ ;
	wire _w932_ ;
	wire _w933_ ;
	wire _w934_ ;
	wire _w935_ ;
	wire _w936_ ;
	wire _w937_ ;
	wire _w938_ ;
	wire _w939_ ;
	wire _w940_ ;
	wire _w941_ ;
	wire _w942_ ;
	wire _w943_ ;
	wire _w944_ ;
	wire _w945_ ;
	wire _w946_ ;
	wire _w947_ ;
	wire _w948_ ;
	wire _w949_ ;
	wire _w950_ ;
	wire _w951_ ;
	wire _w952_ ;
	wire _w953_ ;
	wire _w954_ ;
	wire _w955_ ;
	wire _w956_ ;
	wire _w957_ ;
	wire _w958_ ;
	wire _w959_ ;
	wire _w960_ ;
	wire _w961_ ;
	wire _w962_ ;
	wire _w963_ ;
	wire _w964_ ;
	wire _w965_ ;
	wire _w966_ ;
	wire _w967_ ;
	wire _w968_ ;
	wire _w969_ ;
	wire _w970_ ;
	wire _w971_ ;
	wire _w972_ ;
	wire _w973_ ;
	wire _w974_ ;
	wire _w975_ ;
	wire _w976_ ;
	wire _w977_ ;
	wire _w978_ ;
	wire _w979_ ;
	wire _w980_ ;
	wire _w981_ ;
	wire _w982_ ;
	wire _w983_ ;
	wire _w984_ ;
	wire _w985_ ;
	wire _w986_ ;
	wire _w987_ ;
	wire _w988_ ;
	wire _w989_ ;
	wire _w990_ ;
	wire _w991_ ;
	wire _w992_ ;
	wire _w993_ ;
	wire _w1562_ ;
	wire _w1563_ ;
	wire _w1564_ ;
	wire _w1565_ ;
	wire _w1566_ ;
	wire _w1567_ ;
	wire _w1568_ ;
	wire _w1569_ ;
	wire _w1570_ ;
	wire _w1571_ ;
	wire _w1572_ ;
	wire _w1573_ ;
	wire _w1574_ ;
	wire _w1575_ ;
	wire _w1576_ ;
	wire _w1577_ ;
	wire _w1578_ ;
	wire _w1579_ ;
	wire _w1580_ ;
	wire _w1581_ ;
	wire _w1582_ ;
	wire _w1583_ ;
	wire _w1584_ ;
	wire _w1585_ ;
	wire _w1586_ ;
	wire _w1587_ ;
	wire _w1588_ ;
	wire _w1589_ ;
	wire _w1590_ ;
	wire _w1591_ ;
	wire _w1592_ ;
	wire _w1593_ ;
	wire _w1594_ ;
	wire _w1595_ ;
	wire _w1596_ ;
	wire _w1597_ ;
	wire _w1598_ ;
	wire _w1599_ ;
	wire _w1600_ ;
	wire _w1601_ ;
	wire _w1602_ ;
	wire _w1603_ ;
	wire _w1604_ ;
	wire _w1605_ ;
	wire _w1606_ ;
	wire _w1607_ ;
	wire _w1608_ ;
	wire _w1609_ ;
	wire _w1610_ ;
	wire _w1611_ ;
	wire _w1612_ ;
	wire _w1613_ ;
	wire _w1614_ ;
	wire _w1615_ ;
	wire _w1616_ ;
	wire _w1617_ ;
	wire _w1618_ ;
	wire _w1619_ ;
	wire _w1620_ ;
	wire _w1621_ ;
	wire _w1622_ ;
	wire _w1623_ ;
	wire _w1624_ ;
	wire _w1625_ ;
	wire _w1626_ ;
	wire _w1627_ ;
	wire _w1628_ ;
	wire _w1629_ ;
	wire _w1630_ ;
	wire _w1631_ ;
	wire _w1632_ ;
	wire _w1633_ ;
	wire _w1634_ ;
	wire _w1635_ ;
	wire _w1636_ ;
	wire _w1637_ ;
	wire _w1638_ ;
	wire _w1639_ ;
	wire _w1640_ ;
	wire _w1641_ ;
	wire _w1642_ ;
	wire _w1643_ ;
	wire _w1644_ ;
	wire _w1645_ ;
	wire _w1646_ ;
	wire _w1647_ ;
	wire _w1648_ ;
	wire _w1649_ ;
	wire _w1650_ ;
	wire _w1651_ ;
	wire _w1652_ ;
	wire _w1653_ ;
	wire _w1654_ ;
	wire _w1655_ ;
	wire _w1656_ ;
	wire _w1657_ ;
	wire _w1658_ ;
	wire _w1659_ ;
	wire _w1660_ ;
	wire _w1661_ ;
	wire _w1662_ ;
	wire _w1663_ ;
	wire _w1664_ ;
	wire _w1665_ ;
	wire _w1666_ ;
	wire _w1667_ ;
	wire _w1668_ ;
	wire _w1669_ ;
	wire _w1670_ ;
	wire _w1671_ ;
	wire _w1672_ ;
	wire _w1673_ ;
	wire _w1674_ ;
	wire _w1675_ ;
	wire _w1676_ ;
	wire _w1677_ ;
	wire _w1678_ ;
	wire _w1679_ ;
	wire _w1680_ ;
	wire _w1681_ ;
	wire _w1682_ ;
	wire _w1683_ ;
	wire _w1684_ ;
	wire _w1685_ ;
	wire _w1686_ ;
	wire _w1687_ ;
	wire _w1688_ ;
	wire _w1689_ ;
	wire _w1690_ ;
	wire _w1691_ ;
	wire _w1692_ ;
	wire _w1693_ ;
	wire _w1694_ ;
	wire _w1695_ ;
	wire _w1696_ ;
	wire _w1697_ ;
	wire _w1698_ ;
	wire _w1699_ ;
	wire _w1700_ ;
	wire _w1701_ ;
	wire _w1702_ ;
	wire _w1703_ ;
	wire _w1704_ ;
	wire _w1705_ ;
	wire _w1706_ ;
	wire _w1707_ ;
	wire _w1708_ ;
	wire _w1709_ ;
	wire _w1710_ ;
	wire _w1711_ ;
	wire _w1712_ ;
	wire _w1713_ ;
	wire _w1714_ ;
	wire _w1715_ ;
	wire _w1716_ ;
	wire _w1717_ ;
	wire _w1718_ ;
	wire _w1719_ ;
	wire _w1720_ ;
	wire _w1721_ ;
	wire _w1722_ ;
	wire _w1723_ ;
	wire _w1724_ ;
	wire _w1725_ ;
	wire _w1726_ ;
	wire _w1727_ ;
	wire _w1728_ ;
	wire _w1729_ ;
	wire _w1730_ ;
	wire _w1731_ ;
	wire _w1732_ ;
	wire _w1733_ ;
	wire _w1734_ ;
	wire _w1735_ ;
	wire _w1736_ ;
	wire _w1737_ ;
	wire _w1738_ ;
	wire _w1739_ ;
	wire _w1740_ ;
	wire _w1741_ ;
	wire _w1742_ ;
	wire _w1743_ ;
	wire _w1744_ ;
	wire _w1745_ ;
	wire _w1746_ ;
	wire _w1747_ ;
	wire _w1748_ ;
	wire _w1749_ ;
	wire _w1750_ ;
	wire _w1751_ ;
	wire _w1752_ ;
	wire _w1753_ ;
	wire _w1754_ ;
	wire _w1755_ ;
	wire _w1756_ ;
	wire _w1757_ ;
	wire _w1758_ ;
	wire _w1759_ ;
	wire _w1760_ ;
	wire _w1761_ ;
	wire _w1762_ ;
	wire _w1763_ ;
	wire _w1764_ ;
	wire _w1765_ ;
	wire _w1766_ ;
	wire _w1767_ ;
	wire _w1768_ ;
	wire _w1769_ ;
	wire _w1770_ ;
	wire _w1771_ ;
	wire _w1772_ ;
	wire _w1773_ ;
	wire _w1774_ ;
	wire _w1775_ ;
	wire _w1776_ ;
	wire _w1777_ ;
	wire _w1778_ ;
	wire _w1779_ ;
	wire _w1780_ ;
	wire _w1781_ ;
	wire _w1782_ ;
	wire _w1783_ ;
	wire _w1784_ ;
	wire _w1785_ ;
	wire _w1786_ ;
	wire _w1787_ ;
	wire _w1788_ ;
	wire _w1789_ ;
	wire _w1790_ ;
	wire _w1791_ ;
	wire _w1792_ ;
	wire _w1793_ ;
	wire _w1794_ ;
	wire _w1795_ ;
	wire _w1796_ ;
	wire _w1797_ ;
	wire _w1798_ ;
	wire _w1799_ ;
	wire _w1800_ ;
	wire _w1801_ ;
	wire _w1802_ ;
	wire _w1803_ ;
	wire _w1804_ ;
	wire _w1805_ ;
	wire _w1806_ ;
	wire _w1807_ ;
	wire _w1808_ ;
	wire _w1809_ ;
	wire _w1810_ ;
	wire _w1811_ ;
	wire _w1812_ ;
	wire _w1813_ ;
	wire _w1814_ ;
	wire _w1815_ ;
	wire _w1816_ ;
	wire _w1817_ ;
	wire _w1818_ ;
	wire _w1819_ ;
	wire _w1820_ ;
	wire _w1821_ ;
	wire _w1822_ ;
	wire _w1823_ ;
	wire _w1824_ ;
	wire _w1825_ ;
	wire _w1826_ ;
	wire _w1827_ ;
	wire _w1828_ ;
	wire _w1829_ ;
	wire _w1830_ ;
	wire _w1831_ ;
	wire _w1832_ ;
	wire _w1833_ ;
	wire _w1834_ ;
	wire _w1835_ ;
	wire _w1836_ ;
	wire _w1837_ ;
	wire _w1838_ ;
	wire _w1839_ ;
	wire _w1840_ ;
	wire _w1841_ ;
	wire _w1842_ ;
	wire _w1843_ ;
	wire _w1844_ ;
	wire _w1845_ ;
	wire _w1846_ ;
	wire _w1847_ ;
	wire _w1848_ ;
	wire _w1849_ ;
	wire _w1850_ ;
	wire _w1851_ ;
	wire _w1852_ ;
	wire _w1853_ ;
	wire _w1854_ ;
	wire _w1855_ ;
	wire _w1856_ ;
	wire _w1857_ ;
	wire _w1858_ ;
	wire _w1859_ ;
	wire _w1860_ ;
	wire _w1861_ ;
	wire _w1862_ ;
	wire _w1863_ ;
	wire _w1864_ ;
	wire _w1865_ ;
	wire _w1866_ ;
	wire _w1867_ ;
	wire _w1868_ ;
	wire _w1869_ ;
	wire _w1870_ ;
	wire _w1871_ ;
	wire _w1872_ ;
	wire _w1873_ ;
	wire _w1874_ ;
	wire _w1875_ ;
	wire _w1876_ ;
	wire _w1877_ ;
	wire _w1878_ ;
	wire _w1879_ ;
	wire _w1880_ ;
	wire _w1881_ ;
	wire _w1882_ ;
	wire _w1883_ ;
	wire _w1884_ ;
	wire _w1885_ ;
	wire _w1886_ ;
	wire _w1887_ ;
	wire _w1888_ ;
	wire _w1889_ ;
	wire _w1890_ ;
	wire _w1891_ ;
	wire _w1892_ ;
	wire _w1893_ ;
	wire _w1894_ ;
	wire _w1895_ ;
	wire _w1896_ ;
	wire _w1897_ ;
	wire _w1898_ ;
	wire _w1899_ ;
	wire _w1900_ ;
	wire _w1901_ ;
	wire _w1902_ ;
	wire _w1903_ ;
	wire _w1904_ ;
	wire _w1905_ ;
	wire _w1906_ ;
	wire _w1907_ ;
	wire _w1908_ ;
	wire _w1909_ ;
	wire _w1910_ ;
	wire _w1911_ ;
	wire _w1912_ ;
	wire _w1913_ ;
	wire _w1914_ ;
	wire _w1915_ ;
	wire _w1916_ ;
	wire _w1917_ ;
	wire _w1918_ ;
	wire _w1919_ ;
	wire _w1920_ ;
	wire _w1921_ ;
	wire _w1922_ ;
	wire _w1923_ ;
	wire _w1924_ ;
	wire _w1925_ ;
	wire _w1926_ ;
	wire _w1927_ ;
	wire _w1928_ ;
	wire _w1929_ ;
	wire _w1930_ ;
	wire _w1931_ ;
	wire _w1932_ ;
	wire _w1933_ ;
	wire _w1934_ ;
	wire _w1935_ ;
	wire _w1936_ ;
	wire _w1937_ ;
	wire _w1938_ ;
	wire _w1939_ ;
	wire _w1940_ ;
	wire _w1941_ ;
	wire _w1942_ ;
	wire _w1943_ ;
	wire _w1944_ ;
	wire _w1945_ ;
	wire _w1946_ ;
	wire _w1947_ ;
	wire _w1948_ ;
	wire _w1949_ ;
	wire _w1950_ ;
	wire _w1951_ ;
	wire _w1952_ ;
	wire _w1953_ ;
	wire _w1954_ ;
	wire _w1955_ ;
	wire _w1956_ ;
	wire _w1957_ ;
	wire _w1958_ ;
	wire _w1959_ ;
	wire _w1960_ ;
	wire _w1961_ ;
	wire _w1962_ ;
	wire _w1963_ ;
	wire _w1964_ ;
	wire _w1965_ ;
	wire _w1966_ ;
	wire _w1967_ ;
	wire _w1968_ ;
	wire _w1969_ ;
	wire _w1970_ ;
	wire _w1971_ ;
	wire _w1972_ ;
	wire _w1973_ ;
	wire _w1974_ ;
	wire _w1975_ ;
	wire _w1976_ ;
	wire _w1977_ ;
	wire _w1978_ ;
	wire _w1979_ ;
	wire _w1980_ ;
	wire _w1981_ ;
	wire _w1982_ ;
	wire _w1983_ ;
	wire _w1984_ ;
	wire _w1985_ ;
	wire _w1986_ ;
	wire _w1987_ ;
	wire _w1988_ ;
	wire _w1989_ ;
	wire _w1990_ ;
	wire _w1991_ ;
	wire _w1992_ ;
	wire _w1993_ ;
	wire _w1994_ ;
	wire _w1995_ ;
	wire _w1996_ ;
	wire _w1997_ ;
	wire _w1998_ ;
	wire _w1999_ ;
	wire _w2000_ ;
	wire _w2001_ ;
	wire _w2002_ ;
	wire _w2003_ ;
	wire _w2004_ ;
	wire _w2005_ ;
	wire _w2006_ ;
	wire _w2007_ ;
	wire _w2008_ ;
	wire _w2009_ ;
	wire _w2010_ ;
	wire _w2011_ ;
	wire _w2012_ ;
	wire _w2013_ ;
	wire _w2014_ ;
	wire _w2015_ ;
	wire _w2016_ ;
	wire _w2017_ ;
	wire _w2018_ ;
	wire _w2019_ ;
	wire _w2020_ ;
	wire _w2021_ ;
	wire _w2022_ ;
	wire _w2023_ ;
	wire _w2024_ ;
	wire _w2025_ ;
	wire _w2026_ ;
	wire _w2027_ ;
	wire _w2028_ ;
	wire _w2029_ ;
	wire _w2030_ ;
	wire _w2031_ ;
	wire _w2032_ ;
	wire _w2033_ ;
	wire _w2034_ ;
	wire _w2035_ ;
	wire _w2036_ ;
	wire _w2037_ ;
	wire _w2038_ ;
	wire _w2039_ ;
	wire _w2040_ ;
	wire _w2041_ ;
	wire _w2042_ ;
	wire _w2043_ ;
	wire _w2044_ ;
	wire _w2045_ ;
	wire _w2046_ ;
	wire _w2047_ ;
	wire _w2048_ ;
	wire _w2049_ ;
	wire _w2050_ ;
	wire _w2051_ ;
	wire _w2052_ ;
	wire _w2053_ ;
	wire _w2054_ ;
	wire _w2055_ ;
	wire _w2056_ ;
	wire _w2057_ ;
	wire _w2058_ ;
	wire _w2059_ ;
	wire _w2060_ ;
	wire _w2061_ ;
	wire _w2062_ ;
	wire _w2063_ ;
	wire _w2064_ ;
	wire _w2065_ ;
	wire _w2066_ ;
	wire _w2067_ ;
	wire _w2068_ ;
	wire _w2069_ ;
	wire _w2070_ ;
	wire _w2071_ ;
	wire _w2072_ ;
	wire _w2073_ ;
	wire _w2074_ ;
	wire _w2075_ ;
	wire _w2076_ ;
	wire _w2077_ ;
	wire _w2078_ ;
	wire _w2079_ ;
	wire _w2080_ ;
	wire _w2081_ ;
	wire _w2082_ ;
	wire _w2083_ ;
	wire _w2084_ ;
	wire _w2085_ ;
	wire _w2086_ ;
	wire _w2087_ ;
	wire _w2088_ ;
	wire _w2089_ ;
	wire _w2090_ ;
	wire _w2091_ ;
	wire _w2092_ ;
	wire _w2093_ ;
	wire _w2094_ ;
	wire _w2095_ ;
	wire _w2096_ ;
	wire _w2097_ ;
	wire _w2098_ ;
	wire _w2099_ ;
	wire _w2100_ ;
	wire _w2101_ ;
	wire _w2102_ ;
	wire _w2103_ ;
	wire _w2104_ ;
	wire _w2105_ ;
	wire _w2106_ ;
	wire _w2107_ ;
	wire _w2108_ ;
	wire _w2109_ ;
	wire _w2110_ ;
	wire _w2111_ ;
	wire _w2112_ ;
	wire _w2113_ ;
	wire _w2114_ ;
	wire _w2115_ ;
	wire _w2116_ ;
	wire _w2117_ ;
	wire _w2118_ ;
	wire _w2119_ ;
	wire _w2120_ ;
	wire _w2121_ ;
	wire _w2122_ ;
	wire _w2123_ ;
	wire _w2124_ ;
	wire _w2125_ ;
	wire _w2126_ ;
	wire _w2127_ ;
	wire _w2128_ ;
	wire _w2129_ ;
	wire _w2130_ ;
	wire _w2131_ ;
	wire _w2132_ ;
	wire _w2133_ ;
	wire _w2134_ ;
	wire _w2135_ ;
	wire _w2136_ ;
	wire _w2137_ ;
	wire _w2138_ ;
	wire _w2139_ ;
	wire _w2140_ ;
	wire _w2141_ ;
	wire _w2142_ ;
	wire _w2143_ ;
	wire _w2144_ ;
	wire _w2145_ ;
	wire _w2146_ ;
	wire _w2147_ ;
	wire _w2148_ ;
	wire _w2149_ ;
	wire _w2150_ ;
	wire _w2151_ ;
	wire _w2152_ ;
	wire _w2153_ ;
	wire _w2154_ ;
	wire _w2155_ ;
	wire _w2156_ ;
	wire _w2157_ ;
	wire _w2158_ ;
	wire _w2159_ ;
	wire _w2160_ ;
	wire _w2161_ ;
	wire _w2162_ ;
	wire _w2163_ ;
	wire _w2164_ ;
	wire _w2165_ ;
	wire _w2166_ ;
	wire _w2167_ ;
	wire _w2168_ ;
	wire _w2169_ ;
	wire _w2170_ ;
	wire _w2171_ ;
	wire _w2172_ ;
	wire _w2173_ ;
	wire _w2174_ ;
	wire _w2175_ ;
	wire _w2176_ ;
	wire _w2177_ ;
	wire _w2178_ ;
	wire _w2179_ ;
	wire _w2180_ ;
	wire _w2181_ ;
	wire _w2182_ ;
	wire _w2183_ ;
	wire _w2184_ ;
	wire _w2185_ ;
	wire _w2186_ ;
	wire _w2187_ ;
	wire _w2188_ ;
	wire _w2189_ ;
	wire _w2190_ ;
	wire _w2191_ ;
	wire _w2192_ ;
	wire _w2193_ ;
	wire _w2194_ ;
	wire _w2195_ ;
	wire _w2196_ ;
	wire _w2197_ ;
	wire _w2198_ ;
	wire _w2199_ ;
	wire _w2200_ ;
	wire _w2201_ ;
	wire _w2202_ ;
	wire _w2203_ ;
	wire _w2204_ ;
	wire _w2205_ ;
	wire _w2206_ ;
	wire _w2207_ ;
	wire _w2208_ ;
	wire _w2209_ ;
	wire _w2210_ ;
	wire _w2211_ ;
	wire _w2212_ ;
	wire _w2213_ ;
	wire _w2214_ ;
	wire _w2215_ ;
	wire _w2216_ ;
	wire _w2217_ ;
	wire _w2218_ ;
	wire _w2219_ ;
	wire _w2220_ ;
	wire _w2221_ ;
	wire _w2222_ ;
	wire _w2223_ ;
	wire _w2224_ ;
	wire _w2225_ ;
	wire _w2226_ ;
	wire _w2227_ ;
	wire _w2228_ ;
	wire _w2229_ ;
	wire _w2230_ ;
	wire _w2231_ ;
	wire _w2232_ ;
	wire _w2233_ ;
	wire _w2234_ ;
	wire _w2235_ ;
	wire _w2236_ ;
	wire _w2237_ ;
	wire _w2238_ ;
	wire _w2239_ ;
	wire _w2240_ ;
	wire _w2241_ ;
	wire _w2242_ ;
	wire _w2243_ ;
	wire _w2244_ ;
	wire _w2245_ ;
	wire _w2246_ ;
	wire _w2247_ ;
	wire _w2248_ ;
	wire _w2249_ ;
	wire _w2250_ ;
	wire _w2251_ ;
	wire _w2252_ ;
	wire _w2253_ ;
	wire _w2254_ ;
	wire _w2255_ ;
	wire _w2256_ ;
	wire _w2257_ ;
	wire _w2258_ ;
	wire _w2259_ ;
	wire _w2260_ ;
	wire _w2261_ ;
	wire _w2262_ ;
	wire _w2263_ ;
	wire _w2264_ ;
	wire _w2265_ ;
	wire _w2266_ ;
	wire _w2267_ ;
	wire _w2268_ ;
	wire _w2269_ ;
	wire _w2270_ ;
	wire _w2271_ ;
	wire _w2272_ ;
	wire _w2273_ ;
	wire _w2274_ ;
	wire _w2275_ ;
	wire _w2276_ ;
	wire _w2277_ ;
	wire _w2278_ ;
	wire _w2279_ ;
	wire _w2280_ ;
	wire _w2281_ ;
	wire _w2282_ ;
	wire _w2283_ ;
	wire _w2284_ ;
	wire _w2285_ ;
	wire _w2286_ ;
	wire _w2287_ ;
	wire _w2288_ ;
	wire _w2289_ ;
	wire _w2290_ ;
	wire _w2291_ ;
	wire _w2292_ ;
	wire _w2293_ ;
	wire _w2294_ ;
	wire _w2295_ ;
	wire _w2296_ ;
	wire _w2297_ ;
	wire _w2298_ ;
	wire _w2299_ ;
	wire _w2300_ ;
	wire _w2301_ ;
	wire _w2302_ ;
	wire _w2303_ ;
	wire _w2304_ ;
	wire _w2305_ ;
	wire _w2306_ ;
	wire _w2307_ ;
	wire _w2308_ ;
	wire _w2309_ ;
	wire _w2310_ ;
	wire _w2311_ ;
	wire _w2312_ ;
	wire _w2313_ ;
	wire _w2314_ ;
	wire _w2315_ ;
	wire _w2316_ ;
	wire _w2317_ ;
	wire _w2318_ ;
	wire _w2319_ ;
	wire _w2320_ ;
	wire _w2321_ ;
	wire _w2322_ ;
	wire _w2323_ ;
	wire _w2324_ ;
	wire _w2325_ ;
	wire _w2326_ ;
	wire _w2327_ ;
	wire _w2328_ ;
	wire _w2329_ ;
	wire _w2330_ ;
	wire _w2331_ ;
	wire _w2332_ ;
	wire _w2333_ ;
	wire _w2334_ ;
	wire _w2335_ ;
	wire _w2336_ ;
	wire _w2337_ ;
	wire _w2338_ ;
	wire _w2339_ ;
	wire _w2340_ ;
	wire _w2341_ ;
	wire _w2342_ ;
	wire _w2343_ ;
	wire _w2344_ ;
	wire _w2345_ ;
	wire _w2346_ ;
	wire _w2347_ ;
	wire _w2348_ ;
	wire _w2349_ ;
	wire _w2350_ ;
	wire _w2351_ ;
	wire _w2352_ ;
	wire _w2353_ ;
	wire _w2354_ ;
	wire _w2355_ ;
	wire _w2356_ ;
	wire _w2357_ ;
	wire _w2358_ ;
	wire _w2359_ ;
	wire _w2360_ ;
	wire _w2361_ ;
	wire _w2362_ ;
	wire _w2363_ ;
	wire _w2364_ ;
	wire _w2365_ ;
	wire _w2366_ ;
	wire _w2367_ ;
	wire _w2368_ ;
	wire _w2369_ ;
	wire _w2370_ ;
	wire _w2371_ ;
	wire _w2372_ ;
	wire _w2373_ ;
	wire _w2374_ ;
	wire _w2375_ ;
	wire _w2376_ ;
	wire _w2377_ ;
	wire _w2378_ ;
	wire _w2379_ ;
	wire _w2380_ ;
	wire _w2381_ ;
	wire _w2382_ ;
	wire _w2383_ ;
	wire _w2384_ ;
	wire _w2385_ ;
	wire _w2386_ ;
	wire _w2387_ ;
	wire _w2388_ ;
	wire _w2389_ ;
	wire _w2390_ ;
	wire _w2391_ ;
	wire _w2392_ ;
	wire _w2393_ ;
	wire _w2394_ ;
	wire _w2395_ ;
	wire _w2396_ ;
	wire _w2397_ ;
	wire _w2398_ ;
	wire _w2399_ ;
	wire _w2400_ ;
	wire _w2401_ ;
	wire _w2402_ ;
	wire _w2403_ ;
	wire _w2404_ ;
	wire _w2405_ ;
	wire _w2406_ ;
	wire _w2407_ ;
	wire _w2408_ ;
	wire _w2409_ ;
	wire _w2410_ ;
	wire _w2411_ ;
	wire _w2412_ ;
	wire _w2413_ ;
	wire _w2414_ ;
	wire _w2415_ ;
	wire _w2416_ ;
	wire _w2417_ ;
	wire _w2418_ ;
	wire _w2419_ ;
	wire _w2420_ ;
	wire _w2421_ ;
	wire _w2422_ ;
	wire _w2423_ ;
	wire _w2424_ ;
	wire _w2425_ ;
	wire _w2426_ ;
	wire _w2427_ ;
	wire _w2428_ ;
	wire _w2429_ ;
	wire _w2430_ ;
	wire _w2431_ ;
	wire _w2432_ ;
	wire _w2433_ ;
	wire _w2434_ ;
	wire _w2435_ ;
	wire _w2436_ ;
	wire _w2437_ ;
	wire _w2438_ ;
	wire _w2439_ ;
	wire _w2440_ ;
	wire _w2441_ ;
	wire _w2442_ ;
	wire _w2443_ ;
	wire _w2444_ ;
	wire _w2445_ ;
	wire _w2446_ ;
	wire _w2447_ ;
	wire _w2448_ ;
	wire _w2449_ ;
	wire _w2450_ ;
	wire _w2451_ ;
	wire _w2452_ ;
	wire _w2453_ ;
	wire _w2454_ ;
	wire _w2455_ ;
	wire _w2456_ ;
	wire _w2457_ ;
	wire _w2458_ ;
	wire _w2459_ ;
	wire _w2460_ ;
	wire _w2461_ ;
	wire _w2462_ ;
	wire _w2463_ ;
	wire _w2464_ ;
	wire _w2465_ ;
	wire _w2466_ ;
	wire _w2467_ ;
	wire _w2468_ ;
	wire _w2469_ ;
	wire _w2470_ ;
	wire _w2471_ ;
	wire _w2472_ ;
	wire _w2473_ ;
	wire _w2474_ ;
	wire _w2475_ ;
	wire _w2476_ ;
	wire _w2477_ ;
	wire _w2478_ ;
	wire _w2479_ ;
	wire _w2480_ ;
	wire _w2481_ ;
	wire _w2482_ ;
	wire _w2483_ ;
	wire _w2484_ ;
	wire _w2485_ ;
	wire _w2486_ ;
	wire _w2487_ ;
	wire _w2488_ ;
	wire _w2489_ ;
	wire _w2490_ ;
	wire _w2491_ ;
	wire _w2492_ ;
	wire _w2493_ ;
	wire _w2494_ ;
	wire _w2495_ ;
	wire _w2496_ ;
	wire _w2497_ ;
	wire _w2498_ ;
	wire _w2499_ ;
	wire _w2500_ ;
	wire _w2501_ ;
	wire _w2502_ ;
	wire _w2503_ ;
	wire _w2504_ ;
	wire _w2505_ ;
	wire _w2506_ ;
	wire _w2507_ ;
	wire _w2508_ ;
	wire _w2509_ ;
	wire _w2510_ ;
	wire _w2511_ ;
	wire _w2512_ ;
	wire _w2513_ ;
	wire _w2514_ ;
	wire _w2515_ ;
	wire _w2516_ ;
	wire _w2517_ ;
	wire _w2518_ ;
	wire _w2519_ ;
	wire _w2520_ ;
	wire _w2521_ ;
	wire _w2522_ ;
	wire _w2523_ ;
	wire _w2524_ ;
	wire _w2525_ ;
	wire _w2526_ ;
	wire _w2527_ ;
	wire _w2528_ ;
	wire _w2529_ ;
	wire _w2530_ ;
	wire _w2531_ ;
	wire _w2532_ ;
	wire _w2533_ ;
	wire _w2534_ ;
	wire _w2535_ ;
	wire _w2536_ ;
	wire _w2537_ ;
	wire _w2538_ ;
	wire _w2539_ ;
	wire _w2540_ ;
	wire _w2541_ ;
	wire _w2542_ ;
	wire _w2543_ ;
	wire _w2544_ ;
	wire _w2545_ ;
	wire _w2546_ ;
	wire _w2547_ ;
	wire _w2548_ ;
	wire _w2549_ ;
	wire _w2550_ ;
	wire _w2551_ ;
	wire _w2552_ ;
	wire _w2553_ ;
	wire _w2554_ ;
	wire _w2555_ ;
	wire _w2556_ ;
	wire _w2557_ ;
	wire _w2558_ ;
	wire _w2559_ ;
	wire _w2560_ ;
	wire _w2561_ ;
	wire _w2562_ ;
	wire _w2563_ ;
	wire _w2564_ ;
	wire _w2565_ ;
	wire _w2566_ ;
	wire _w2567_ ;
	wire _w2568_ ;
	wire _w2569_ ;
	wire _w2570_ ;
	wire _w2571_ ;
	wire _w2572_ ;
	wire _w2573_ ;
	wire _w2574_ ;
	wire _w2575_ ;
	wire _w2576_ ;
	wire _w2577_ ;
	wire _w2578_ ;
	wire _w2579_ ;
	wire _w2580_ ;
	wire _w2581_ ;
	wire _w2582_ ;
	wire _w2583_ ;
	wire _w2584_ ;
	wire _w2585_ ;
	wire _w2586_ ;
	wire _w2587_ ;
	wire _w2588_ ;
	wire _w2589_ ;
	wire _w2590_ ;
	wire _w2591_ ;
	wire _w2592_ ;
	wire _w2593_ ;
	wire _w2594_ ;
	wire _w2595_ ;
	wire _w2596_ ;
	wire _w2597_ ;
	wire _w2598_ ;
	wire _w2599_ ;
	wire _w2600_ ;
	wire _w2601_ ;
	wire _w2602_ ;
	wire _w2603_ ;
	wire _w2604_ ;
	wire _w2605_ ;
	wire _w2606_ ;
	wire _w2607_ ;
	wire _w2608_ ;
	wire _w2609_ ;
	wire _w2610_ ;
	wire _w2611_ ;
	wire _w2612_ ;
	wire _w2613_ ;
	wire _w2614_ ;
	wire _w2615_ ;
	wire _w2616_ ;
	wire _w2617_ ;
	wire _w2618_ ;
	wire _w2619_ ;
	wire _w2620_ ;
	wire _w2621_ ;
	wire _w2622_ ;
	wire _w2623_ ;
	wire _w2624_ ;
	wire _w2625_ ;
	wire _w2626_ ;
	wire _w2627_ ;
	wire _w2628_ ;
	wire _w2629_ ;
	wire _w2630_ ;
	wire _w2631_ ;
	wire _w2632_ ;
	wire _w2633_ ;
	wire _w2634_ ;
	wire _w2635_ ;
	wire _w2636_ ;
	wire _w2637_ ;
	wire _w2638_ ;
	wire _w2639_ ;
	wire _w2640_ ;
	wire _w2641_ ;
	wire _w2642_ ;
	wire _w2643_ ;
	wire _w2644_ ;
	wire _w2645_ ;
	wire _w2646_ ;
	wire _w2647_ ;
	wire _w2648_ ;
	wire _w2649_ ;
	wire _w2650_ ;
	wire _w2651_ ;
	wire _w2652_ ;
	wire _w2653_ ;
	wire _w2654_ ;
	wire _w2655_ ;
	wire _w2656_ ;
	wire _w2657_ ;
	wire _w2658_ ;
	wire _w2659_ ;
	wire _w2660_ ;
	wire _w2661_ ;
	wire _w2662_ ;
	wire _w2663_ ;
	wire _w2664_ ;
	wire _w2665_ ;
	wire _w2666_ ;
	wire _w2667_ ;
	wire _w2668_ ;
	wire _w2669_ ;
	wire _w2670_ ;
	wire _w2671_ ;
	wire _w2672_ ;
	wire _w2673_ ;
	wire _w2674_ ;
	wire _w2675_ ;
	wire _w2676_ ;
	wire _w2677_ ;
	wire _w2678_ ;
	wire _w2679_ ;
	wire _w2680_ ;
	wire _w2681_ ;
	wire _w2682_ ;
	wire _w2683_ ;
	wire _w2684_ ;
	wire _w2685_ ;
	wire _w2686_ ;
	wire _w2687_ ;
	wire _w2688_ ;
	wire _w2689_ ;
	wire _w2690_ ;
	wire _w2691_ ;
	wire _w2692_ ;
	wire _w2693_ ;
	wire _w2694_ ;
	wire _w2695_ ;
	wire _w2696_ ;
	wire _w2697_ ;
	wire _w2698_ ;
	wire _w2699_ ;
	wire _w2700_ ;
	wire _w2701_ ;
	wire _w2702_ ;
	wire _w2703_ ;
	wire _w2704_ ;
	wire _w2705_ ;
	wire _w2706_ ;
	wire _w2707_ ;
	wire _w2708_ ;
	wire _w2709_ ;
	wire _w2710_ ;
	wire _w2711_ ;
	wire _w2712_ ;
	wire _w2713_ ;
	wire _w2714_ ;
	wire _w2715_ ;
	wire _w2716_ ;
	wire _w2717_ ;
	wire _w2718_ ;
	wire _w2719_ ;
	wire _w2720_ ;
	wire _w2721_ ;
	wire _w2722_ ;
	wire _w2723_ ;
	wire _w2724_ ;
	wire _w2725_ ;
	wire _w2726_ ;
	wire _w2727_ ;
	wire _w2728_ ;
	wire _w2729_ ;
	wire _w2730_ ;
	wire _w2731_ ;
	wire _w2732_ ;
	wire _w2733_ ;
	wire _w2734_ ;
	wire _w2735_ ;
	wire _w2736_ ;
	wire _w2737_ ;
	wire _w2738_ ;
	wire _w2739_ ;
	wire _w2740_ ;
	wire _w2741_ ;
	wire _w2742_ ;
	wire _w2743_ ;
	wire _w2744_ ;
	wire _w2745_ ;
	wire _w2746_ ;
	wire _w2747_ ;
	wire _w2748_ ;
	wire _w2749_ ;
	wire _w2750_ ;
	wire _w2751_ ;
	wire _w2752_ ;
	wire _w2753_ ;
	wire _w2754_ ;
	wire _w2755_ ;
	wire _w2756_ ;
	wire _w2757_ ;
	wire _w2758_ ;
	wire _w2759_ ;
	wire _w2760_ ;
	wire _w2761_ ;
	wire _w2762_ ;
	wire _w2763_ ;
	wire _w2764_ ;
	wire _w2765_ ;
	wire _w2766_ ;
	wire _w2767_ ;
	wire _w2768_ ;
	wire _w2769_ ;
	wire _w2770_ ;
	wire _w2771_ ;
	wire _w2772_ ;
	wire _w2773_ ;
	wire _w2774_ ;
	wire _w2775_ ;
	wire _w2776_ ;
	wire _w2777_ ;
	wire _w2778_ ;
	wire _w2779_ ;
	wire _w2780_ ;
	wire _w2781_ ;
	wire _w2782_ ;
	wire _w2783_ ;
	wire _w2784_ ;
	wire _w2785_ ;
	wire _w2786_ ;
	wire _w2787_ ;
	wire _w2788_ ;
	wire _w2789_ ;
	wire _w2790_ ;
	wire _w2791_ ;
	wire _w2792_ ;
	wire _w2793_ ;
	wire _w2794_ ;
	wire _w2795_ ;
	wire _w2796_ ;
	wire _w2797_ ;
	wire _w2798_ ;
	wire _w2799_ ;
	wire _w2800_ ;
	wire _w2801_ ;
	wire _w2802_ ;
	wire _w2803_ ;
	wire _w2804_ ;
	wire _w2805_ ;
	wire _w2806_ ;
	wire _w2807_ ;
	wire _w2808_ ;
	wire _w2809_ ;
	LUT4 #(
		.INIT('h0040)
	) name0 (
		\InstQueueRd_Addr_reg[0]/NET0131 ,
		\InstQueueRd_Addr_reg[1]/NET0131 ,
		\InstQueueRd_Addr_reg[2]/NET0131 ,
		\InstQueueRd_Addr_reg[3]/NET0131 ,
		_w453_
	);
	LUT2 #(
		.INIT('h8)
	) name1 (
		\InstQueueRd_Addr_reg[0]/NET0131 ,
		\InstQueueRd_Addr_reg[1]/NET0131 ,
		_w454_
	);
	LUT4 #(
		.INIT('h8000)
	) name2 (
		\InstQueueRd_Addr_reg[0]/NET0131 ,
		\InstQueueRd_Addr_reg[1]/NET0131 ,
		\InstQueueRd_Addr_reg[2]/NET0131 ,
		\InstQueueRd_Addr_reg[3]/NET0131 ,
		_w455_
	);
	LUT4 #(
		.INIT('h153f)
	) name3 (
		\InstQueue_reg[15][2]/NET0131 ,
		\InstQueue_reg[6][2]/NET0131 ,
		_w453_,
		_w455_,
		_w456_
	);
	LUT4 #(
		.INIT('h0020)
	) name4 (
		\InstQueueRd_Addr_reg[0]/NET0131 ,
		\InstQueueRd_Addr_reg[1]/NET0131 ,
		\InstQueueRd_Addr_reg[2]/NET0131 ,
		\InstQueueRd_Addr_reg[3]/NET0131 ,
		_w457_
	);
	LUT4 #(
		.INIT('h0800)
	) name5 (
		\InstQueueRd_Addr_reg[0]/NET0131 ,
		\InstQueueRd_Addr_reg[1]/NET0131 ,
		\InstQueueRd_Addr_reg[2]/NET0131 ,
		\InstQueueRd_Addr_reg[3]/NET0131 ,
		_w458_
	);
	LUT4 #(
		.INIT('h153f)
	) name6 (
		\InstQueue_reg[11][2]/NET0131 ,
		\InstQueue_reg[5][2]/NET0131 ,
		_w457_,
		_w458_,
		_w459_
	);
	LUT4 #(
		.INIT('h0008)
	) name7 (
		\InstQueueRd_Addr_reg[0]/NET0131 ,
		\InstQueueRd_Addr_reg[1]/NET0131 ,
		\InstQueueRd_Addr_reg[2]/NET0131 ,
		\InstQueueRd_Addr_reg[3]/NET0131 ,
		_w460_
	);
	LUT4 #(
		.INIT('h2000)
	) name8 (
		\InstQueueRd_Addr_reg[0]/NET0131 ,
		\InstQueueRd_Addr_reg[1]/NET0131 ,
		\InstQueueRd_Addr_reg[2]/NET0131 ,
		\InstQueueRd_Addr_reg[3]/NET0131 ,
		_w461_
	);
	LUT4 #(
		.INIT('h135f)
	) name9 (
		\InstQueue_reg[13][2]/NET0131 ,
		\InstQueue_reg[3][2]/NET0131 ,
		_w461_,
		_w460_,
		_w462_
	);
	LUT4 #(
		.INIT('h0100)
	) name10 (
		\InstQueueRd_Addr_reg[0]/NET0131 ,
		\InstQueueRd_Addr_reg[1]/NET0131 ,
		\InstQueueRd_Addr_reg[2]/NET0131 ,
		\InstQueueRd_Addr_reg[3]/NET0131 ,
		_w463_
	);
	LUT4 #(
		.INIT('h0001)
	) name11 (
		\InstQueueRd_Addr_reg[0]/NET0131 ,
		\InstQueueRd_Addr_reg[1]/NET0131 ,
		\InstQueueRd_Addr_reg[2]/NET0131 ,
		\InstQueueRd_Addr_reg[3]/NET0131 ,
		_w464_
	);
	LUT4 #(
		.INIT('h135f)
	) name12 (
		\InstQueue_reg[0][2]/NET0131 ,
		\InstQueue_reg[8][2]/NET0131 ,
		_w464_,
		_w463_,
		_w465_
	);
	LUT4 #(
		.INIT('h8000)
	) name13 (
		_w462_,
		_w465_,
		_w456_,
		_w459_,
		_w466_
	);
	LUT4 #(
		.INIT('h0200)
	) name14 (
		\InstQueueRd_Addr_reg[0]/NET0131 ,
		\InstQueueRd_Addr_reg[1]/NET0131 ,
		\InstQueueRd_Addr_reg[2]/NET0131 ,
		\InstQueueRd_Addr_reg[3]/NET0131 ,
		_w467_
	);
	LUT4 #(
		.INIT('h0010)
	) name15 (
		\InstQueueRd_Addr_reg[0]/NET0131 ,
		\InstQueueRd_Addr_reg[1]/NET0131 ,
		\InstQueueRd_Addr_reg[2]/NET0131 ,
		\InstQueueRd_Addr_reg[3]/NET0131 ,
		_w468_
	);
	LUT4 #(
		.INIT('h135f)
	) name16 (
		\InstQueue_reg[4][2]/NET0131 ,
		\InstQueue_reg[9][2]/NET0131 ,
		_w468_,
		_w467_,
		_w469_
	);
	LUT4 #(
		.INIT('h0080)
	) name17 (
		\InstQueueRd_Addr_reg[0]/NET0131 ,
		\InstQueueRd_Addr_reg[1]/NET0131 ,
		\InstQueueRd_Addr_reg[2]/NET0131 ,
		\InstQueueRd_Addr_reg[3]/NET0131 ,
		_w470_
	);
	LUT4 #(
		.INIT('h0400)
	) name18 (
		\InstQueueRd_Addr_reg[0]/NET0131 ,
		\InstQueueRd_Addr_reg[1]/NET0131 ,
		\InstQueueRd_Addr_reg[2]/NET0131 ,
		\InstQueueRd_Addr_reg[3]/NET0131 ,
		_w471_
	);
	LUT4 #(
		.INIT('h153f)
	) name19 (
		\InstQueue_reg[10][2]/NET0131 ,
		\InstQueue_reg[7][2]/NET0131 ,
		_w470_,
		_w471_,
		_w472_
	);
	LUT4 #(
		.INIT('h0002)
	) name20 (
		\InstQueueRd_Addr_reg[0]/NET0131 ,
		\InstQueueRd_Addr_reg[1]/NET0131 ,
		\InstQueueRd_Addr_reg[2]/NET0131 ,
		\InstQueueRd_Addr_reg[3]/NET0131 ,
		_w473_
	);
	LUT4 #(
		.INIT('h0004)
	) name21 (
		\InstQueueRd_Addr_reg[0]/NET0131 ,
		\InstQueueRd_Addr_reg[1]/NET0131 ,
		\InstQueueRd_Addr_reg[2]/NET0131 ,
		\InstQueueRd_Addr_reg[3]/NET0131 ,
		_w474_
	);
	LUT4 #(
		.INIT('h153f)
	) name22 (
		\InstQueue_reg[1][2]/NET0131 ,
		\InstQueue_reg[2][2]/NET0131 ,
		_w474_,
		_w473_,
		_w475_
	);
	LUT4 #(
		.INIT('h4000)
	) name23 (
		\InstQueueRd_Addr_reg[0]/NET0131 ,
		\InstQueueRd_Addr_reg[1]/NET0131 ,
		\InstQueueRd_Addr_reg[2]/NET0131 ,
		\InstQueueRd_Addr_reg[3]/NET0131 ,
		_w476_
	);
	LUT4 #(
		.INIT('h1000)
	) name24 (
		\InstQueueRd_Addr_reg[0]/NET0131 ,
		\InstQueueRd_Addr_reg[1]/NET0131 ,
		\InstQueueRd_Addr_reg[2]/NET0131 ,
		\InstQueueRd_Addr_reg[3]/NET0131 ,
		_w477_
	);
	LUT4 #(
		.INIT('h135f)
	) name25 (
		\InstQueue_reg[12][2]/NET0131 ,
		\InstQueue_reg[14][2]/NET0131 ,
		_w477_,
		_w476_,
		_w478_
	);
	LUT4 #(
		.INIT('h8000)
	) name26 (
		_w475_,
		_w478_,
		_w469_,
		_w472_,
		_w479_
	);
	LUT2 #(
		.INIT('h8)
	) name27 (
		_w466_,
		_w479_,
		_w480_
	);
	LUT2 #(
		.INIT('h8)
	) name28 (
		\InstQueueRd_Addr_reg[1]/NET0131 ,
		\InstQueueRd_Addr_reg[2]/NET0131 ,
		_w481_
	);
	LUT3 #(
		.INIT('h80)
	) name29 (
		\InstQueueRd_Addr_reg[1]/NET0131 ,
		\InstQueueRd_Addr_reg[2]/NET0131 ,
		\InstQueueRd_Addr_reg[3]/NET0131 ,
		_w482_
	);
	LUT2 #(
		.INIT('h8)
	) name30 (
		\InstQueueRd_Addr_reg[0]/NET0131 ,
		\InstQueue_reg[15][1]/NET0131 ,
		_w483_
	);
	LUT4 #(
		.INIT('h0777)
	) name31 (
		\InstQueue_reg[7][1]/NET0131 ,
		_w470_,
		_w482_,
		_w483_,
		_w484_
	);
	LUT4 #(
		.INIT('h135f)
	) name32 (
		\InstQueue_reg[3][1]/NET0131 ,
		\InstQueue_reg[9][1]/NET0131 ,
		_w460_,
		_w467_,
		_w485_
	);
	LUT4 #(
		.INIT('h135f)
	) name33 (
		\InstQueue_reg[4][1]/NET0131 ,
		\InstQueue_reg[6][1]/NET0131 ,
		_w468_,
		_w453_,
		_w486_
	);
	LUT4 #(
		.INIT('h135f)
	) name34 (
		\InstQueue_reg[0][1]/NET0131 ,
		\InstQueue_reg[8][1]/NET0131 ,
		_w464_,
		_w463_,
		_w487_
	);
	LUT4 #(
		.INIT('h8000)
	) name35 (
		_w486_,
		_w487_,
		_w484_,
		_w485_,
		_w488_
	);
	LUT4 #(
		.INIT('h153f)
	) name36 (
		\InstQueue_reg[12][1]/NET0131 ,
		\InstQueue_reg[2][1]/NET0131 ,
		_w474_,
		_w477_,
		_w489_
	);
	LUT4 #(
		.INIT('h153f)
	) name37 (
		\InstQueue_reg[11][1]/NET0131 ,
		\InstQueue_reg[14][1]/NET0131 ,
		_w476_,
		_w458_,
		_w490_
	);
	LUT4 #(
		.INIT('h135f)
	) name38 (
		\InstQueue_reg[10][1]/NET0131 ,
		\InstQueue_reg[13][1]/NET0131 ,
		_w471_,
		_w461_,
		_w491_
	);
	LUT4 #(
		.INIT('h135f)
	) name39 (
		\InstQueue_reg[1][1]/NET0131 ,
		\InstQueue_reg[5][1]/NET0131 ,
		_w473_,
		_w457_,
		_w492_
	);
	LUT4 #(
		.INIT('h8000)
	) name40 (
		_w491_,
		_w492_,
		_w489_,
		_w490_,
		_w493_
	);
	LUT2 #(
		.INIT('h8)
	) name41 (
		_w488_,
		_w493_,
		_w494_
	);
	LUT4 #(
		.INIT('h8000)
	) name42 (
		_w466_,
		_w479_,
		_w488_,
		_w493_,
		_w495_
	);
	LUT4 #(
		.INIT('h135f)
	) name43 (
		\InstQueue_reg[12][0]/NET0131 ,
		\InstQueue_reg[14][0]/NET0131 ,
		_w477_,
		_w476_,
		_w496_
	);
	LUT4 #(
		.INIT('h153f)
	) name44 (
		\InstQueue_reg[0][0]/NET0131 ,
		\InstQueue_reg[4][0]/NET0131 ,
		_w468_,
		_w464_,
		_w497_
	);
	LUT4 #(
		.INIT('h153f)
	) name45 (
		\InstQueue_reg[2][0]/NET0131 ,
		\InstQueue_reg[7][0]/NET0131 ,
		_w470_,
		_w474_,
		_w498_
	);
	LUT4 #(
		.INIT('h135f)
	) name46 (
		\InstQueue_reg[10][0]/NET0131 ,
		\InstQueue_reg[13][0]/NET0131 ,
		_w471_,
		_w461_,
		_w499_
	);
	LUT4 #(
		.INIT('h8000)
	) name47 (
		_w498_,
		_w499_,
		_w496_,
		_w497_,
		_w500_
	);
	LUT4 #(
		.INIT('h153f)
	) name48 (
		\InstQueue_reg[1][0]/NET0131 ,
		\InstQueue_reg[8][0]/NET0131 ,
		_w463_,
		_w473_,
		_w501_
	);
	LUT4 #(
		.INIT('h153f)
	) name49 (
		\InstQueue_reg[11][0]/NET0131 ,
		\InstQueue_reg[5][0]/NET0131 ,
		_w457_,
		_w458_,
		_w502_
	);
	LUT2 #(
		.INIT('h8)
	) name50 (
		\InstQueueRd_Addr_reg[0]/NET0131 ,
		\InstQueue_reg[15][0]/NET0131 ,
		_w503_
	);
	LUT4 #(
		.INIT('h0777)
	) name51 (
		\InstQueue_reg[3][0]/NET0131 ,
		_w460_,
		_w482_,
		_w503_,
		_w504_
	);
	LUT4 #(
		.INIT('h135f)
	) name52 (
		\InstQueue_reg[6][0]/NET0131 ,
		\InstQueue_reg[9][0]/NET0131 ,
		_w453_,
		_w467_,
		_w505_
	);
	LUT4 #(
		.INIT('h8000)
	) name53 (
		_w504_,
		_w505_,
		_w501_,
		_w502_,
		_w506_
	);
	LUT4 #(
		.INIT('h153f)
	) name54 (
		\InstQueue_reg[1][3]/NET0131 ,
		\InstQueue_reg[4][3]/NET0131 ,
		_w468_,
		_w473_,
		_w507_
	);
	LUT4 #(
		.INIT('h135f)
	) name55 (
		\InstQueue_reg[10][3]/NET0131 ,
		\InstQueue_reg[13][3]/NET0131 ,
		_w471_,
		_w461_,
		_w508_
	);
	LUT4 #(
		.INIT('h135f)
	) name56 (
		\InstQueue_reg[3][3]/NET0131 ,
		\InstQueue_reg[8][3]/NET0131 ,
		_w460_,
		_w463_,
		_w509_
	);
	LUT4 #(
		.INIT('h135f)
	) name57 (
		\InstQueue_reg[12][3]/NET0131 ,
		\InstQueue_reg[5][3]/NET0131 ,
		_w477_,
		_w457_,
		_w510_
	);
	LUT4 #(
		.INIT('h8000)
	) name58 (
		_w509_,
		_w510_,
		_w507_,
		_w508_,
		_w511_
	);
	LUT4 #(
		.INIT('h153f)
	) name59 (
		\InstQueue_reg[15][3]/NET0131 ,
		\InstQueue_reg[2][3]/NET0131 ,
		_w474_,
		_w455_,
		_w512_
	);
	LUT4 #(
		.INIT('h135f)
	) name60 (
		\InstQueue_reg[0][3]/NET0131 ,
		\InstQueue_reg[6][3]/NET0131 ,
		_w464_,
		_w453_,
		_w513_
	);
	LUT4 #(
		.INIT('h135f)
	) name61 (
		\InstQueue_reg[14][3]/NET0131 ,
		\InstQueue_reg[9][3]/NET0131 ,
		_w476_,
		_w467_,
		_w514_
	);
	LUT4 #(
		.INIT('h153f)
	) name62 (
		\InstQueue_reg[11][3]/NET0131 ,
		\InstQueue_reg[7][3]/NET0131 ,
		_w470_,
		_w458_,
		_w515_
	);
	LUT4 #(
		.INIT('h8000)
	) name63 (
		_w514_,
		_w515_,
		_w512_,
		_w513_,
		_w516_
	);
	LUT4 #(
		.INIT('h8000)
	) name64 (
		_w500_,
		_w506_,
		_w511_,
		_w516_,
		_w517_
	);
	LUT2 #(
		.INIT('h8)
	) name65 (
		_w495_,
		_w517_,
		_w518_
	);
	LUT4 #(
		.INIT('h135f)
	) name66 (
		\InstQueue_reg[13][6]/NET0131 ,
		\InstQueue_reg[1][6]/NET0131 ,
		_w461_,
		_w473_,
		_w519_
	);
	LUT4 #(
		.INIT('h135f)
	) name67 (
		\InstQueue_reg[0][6]/NET0131 ,
		\InstQueue_reg[9][6]/NET0131 ,
		_w464_,
		_w467_,
		_w520_
	);
	LUT4 #(
		.INIT('h135f)
	) name68 (
		\InstQueue_reg[3][6]/NET0131 ,
		\InstQueue_reg[8][6]/NET0131 ,
		_w460_,
		_w463_,
		_w521_
	);
	LUT4 #(
		.INIT('h153f)
	) name69 (
		\InstQueue_reg[15][6]/NET0131 ,
		\InstQueue_reg[5][6]/NET0131 ,
		_w457_,
		_w455_,
		_w522_
	);
	LUT4 #(
		.INIT('h8000)
	) name70 (
		_w521_,
		_w522_,
		_w519_,
		_w520_,
		_w523_
	);
	LUT4 #(
		.INIT('h153f)
	) name71 (
		\InstQueue_reg[2][6]/NET0131 ,
		\InstQueue_reg[7][6]/NET0131 ,
		_w470_,
		_w474_,
		_w524_
	);
	LUT4 #(
		.INIT('h135f)
	) name72 (
		\InstQueue_reg[10][6]/NET0131 ,
		\InstQueue_reg[12][6]/NET0131 ,
		_w471_,
		_w477_,
		_w525_
	);
	LUT4 #(
		.INIT('h135f)
	) name73 (
		\InstQueue_reg[14][6]/NET0131 ,
		\InstQueue_reg[6][6]/NET0131 ,
		_w476_,
		_w453_,
		_w526_
	);
	LUT4 #(
		.INIT('h153f)
	) name74 (
		\InstQueue_reg[11][6]/NET0131 ,
		\InstQueue_reg[4][6]/NET0131 ,
		_w468_,
		_w458_,
		_w527_
	);
	LUT4 #(
		.INIT('h8000)
	) name75 (
		_w526_,
		_w527_,
		_w524_,
		_w525_,
		_w528_
	);
	LUT2 #(
		.INIT('h8)
	) name76 (
		_w523_,
		_w528_,
		_w529_
	);
	LUT4 #(
		.INIT('h135f)
	) name77 (
		\InstQueue_reg[0][5]/NET0131 ,
		\InstQueue_reg[1][5]/NET0131 ,
		_w464_,
		_w473_,
		_w530_
	);
	LUT4 #(
		.INIT('h135f)
	) name78 (
		\InstQueue_reg[4][5]/NET0131 ,
		\InstQueue_reg[6][5]/NET0131 ,
		_w468_,
		_w453_,
		_w531_
	);
	LUT4 #(
		.INIT('h153f)
	) name79 (
		\InstQueue_reg[11][5]/NET0131 ,
		\InstQueue_reg[3][5]/NET0131 ,
		_w460_,
		_w458_,
		_w532_
	);
	LUT4 #(
		.INIT('h153f)
	) name80 (
		\InstQueue_reg[15][5]/NET0131 ,
		\InstQueue_reg[5][5]/NET0131 ,
		_w457_,
		_w455_,
		_w533_
	);
	LUT4 #(
		.INIT('h8000)
	) name81 (
		_w532_,
		_w533_,
		_w530_,
		_w531_,
		_w534_
	);
	LUT4 #(
		.INIT('h153f)
	) name82 (
		\InstQueue_reg[13][5]/NET0131 ,
		\InstQueue_reg[2][5]/NET0131 ,
		_w474_,
		_w461_,
		_w535_
	);
	LUT4 #(
		.INIT('h135f)
	) name83 (
		\InstQueue_reg[10][5]/NET0131 ,
		\InstQueue_reg[12][5]/NET0131 ,
		_w471_,
		_w477_,
		_w536_
	);
	LUT4 #(
		.INIT('h135f)
	) name84 (
		\InstQueue_reg[14][5]/NET0131 ,
		\InstQueue_reg[9][5]/NET0131 ,
		_w476_,
		_w467_,
		_w537_
	);
	LUT4 #(
		.INIT('h135f)
	) name85 (
		\InstQueue_reg[7][5]/NET0131 ,
		\InstQueue_reg[8][5]/NET0131 ,
		_w470_,
		_w463_,
		_w538_
	);
	LUT4 #(
		.INIT('h8000)
	) name86 (
		_w537_,
		_w538_,
		_w535_,
		_w536_,
		_w539_
	);
	LUT2 #(
		.INIT('h8)
	) name87 (
		_w534_,
		_w539_,
		_w540_
	);
	LUT2 #(
		.INIT('h8)
	) name88 (
		\InstQueueRd_Addr_reg[0]/NET0131 ,
		\InstQueue_reg[15][7]/NET0131 ,
		_w541_
	);
	LUT4 #(
		.INIT('h0777)
	) name89 (
		\InstQueue_reg[4][7]/NET0131 ,
		_w468_,
		_w482_,
		_w541_,
		_w542_
	);
	LUT4 #(
		.INIT('h153f)
	) name90 (
		\InstQueue_reg[0][7]/NET0131 ,
		\InstQueue_reg[14][7]/NET0131 ,
		_w476_,
		_w464_,
		_w543_
	);
	LUT4 #(
		.INIT('h153f)
	) name91 (
		\InstQueue_reg[12][7]/NET0131 ,
		\InstQueue_reg[13][7]/NET0131 ,
		_w461_,
		_w477_,
		_w544_
	);
	LUT4 #(
		.INIT('h153f)
	) name92 (
		\InstQueue_reg[11][7]/NET0131 ,
		\InstQueue_reg[5][7]/NET0131 ,
		_w457_,
		_w458_,
		_w545_
	);
	LUT4 #(
		.INIT('h8000)
	) name93 (
		_w544_,
		_w545_,
		_w542_,
		_w543_,
		_w546_
	);
	LUT4 #(
		.INIT('h153f)
	) name94 (
		\InstQueue_reg[1][7]/NET0131 ,
		\InstQueue_reg[6][7]/NET0131 ,
		_w453_,
		_w473_,
		_w547_
	);
	LUT4 #(
		.INIT('h153f)
	) name95 (
		\InstQueue_reg[8][7]/NET0131 ,
		\InstQueue_reg[9][7]/NET0131 ,
		_w467_,
		_w463_,
		_w548_
	);
	LUT4 #(
		.INIT('h153f)
	) name96 (
		\InstQueue_reg[3][7]/NET0131 ,
		\InstQueue_reg[7][7]/NET0131 ,
		_w470_,
		_w460_,
		_w549_
	);
	LUT4 #(
		.INIT('h153f)
	) name97 (
		\InstQueue_reg[10][7]/NET0131 ,
		\InstQueue_reg[2][7]/NET0131 ,
		_w474_,
		_w471_,
		_w550_
	);
	LUT4 #(
		.INIT('h8000)
	) name98 (
		_w549_,
		_w550_,
		_w547_,
		_w548_,
		_w551_
	);
	LUT2 #(
		.INIT('h8)
	) name99 (
		_w546_,
		_w551_,
		_w552_
	);
	LUT4 #(
		.INIT('h0888)
	) name100 (
		_w534_,
		_w539_,
		_w546_,
		_w551_,
		_w553_
	);
	LUT4 #(
		.INIT('h4000)
	) name101 (
		_w529_,
		_w495_,
		_w517_,
		_w553_,
		_w554_
	);
	LUT2 #(
		.INIT('h4)
	) name102 (
		\InstQueueRd_Addr_reg[3]/NET0131 ,
		\InstQueueWr_Addr_reg[3]/NET0131 ,
		_w555_
	);
	LUT4 #(
		.INIT('h08ce)
	) name103 (
		\InstQueueRd_Addr_reg[0]/NET0131 ,
		\InstQueueRd_Addr_reg[1]/NET0131 ,
		\InstQueueWr_Addr_reg[0]/NET0131 ,
		\InstQueueWr_Addr_reg[1]/NET0131 ,
		_w556_
	);
	LUT3 #(
		.INIT('hb2)
	) name104 (
		\InstQueueRd_Addr_reg[2]/NET0131 ,
		\InstQueueWr_Addr_reg[2]/NET0131 ,
		_w556_,
		_w557_
	);
	LUT4 #(
		.INIT('h40d0)
	) name105 (
		\InstQueueRd_Addr_reg[2]/NET0131 ,
		\InstQueueWr_Addr_reg[2]/NET0131 ,
		_w555_,
		_w556_,
		_w558_
	);
	LUT2 #(
		.INIT('h2)
	) name106 (
		\InstQueueRd_Addr_reg[3]/NET0131 ,
		\InstQueueWr_Addr_reg[3]/NET0131 ,
		_w559_
	);
	LUT4 #(
		.INIT('h004d)
	) name107 (
		\InstQueueRd_Addr_reg[2]/NET0131 ,
		\InstQueueWr_Addr_reg[2]/NET0131 ,
		_w556_,
		_w559_,
		_w560_
	);
	LUT2 #(
		.INIT('h9)
	) name108 (
		\InstQueueRd_Addr_reg[2]/NET0131 ,
		\InstQueueWr_Addr_reg[2]/NET0131 ,
		_w561_
	);
	LUT2 #(
		.INIT('h9)
	) name109 (
		_w556_,
		_w561_,
		_w562_
	);
	LUT4 #(
		.INIT('hb2fb)
	) name110 (
		\InstQueueRd_Addr_reg[3]/NET0131 ,
		\InstQueueWr_Addr_reg[3]/NET0131 ,
		_w557_,
		_w562_,
		_w563_
	);
	LUT4 #(
		.INIT('h39c6)
	) name111 (
		\InstQueueRd_Addr_reg[0]/NET0131 ,
		\InstQueueRd_Addr_reg[1]/NET0131 ,
		\InstQueueWr_Addr_reg[0]/NET0131 ,
		\InstQueueWr_Addr_reg[1]/NET0131 ,
		_w564_
	);
	LUT3 #(
		.INIT('he0)
	) name112 (
		_w555_,
		_w560_,
		_w564_,
		_w565_
	);
	LUT2 #(
		.INIT('h2)
	) name113 (
		_w563_,
		_w565_,
		_w566_
	);
	LUT4 #(
		.INIT('h0777)
	) name114 (
		_w500_,
		_w506_,
		_w511_,
		_w516_,
		_w567_
	);
	LUT4 #(
		.INIT('h0888)
	) name115 (
		_w466_,
		_w479_,
		_w488_,
		_w493_,
		_w568_
	);
	LUT2 #(
		.INIT('h8)
	) name116 (
		_w567_,
		_w568_,
		_w569_
	);
	LUT4 #(
		.INIT('h153f)
	) name117 (
		\InstQueue_reg[0][4]/NET0131 ,
		\InstQueue_reg[2][4]/NET0131 ,
		_w474_,
		_w464_,
		_w570_
	);
	LUT4 #(
		.INIT('h135f)
	) name118 (
		\InstQueue_reg[12][4]/NET0131 ,
		\InstQueue_reg[4][4]/NET0131 ,
		_w477_,
		_w468_,
		_w571_
	);
	LUT4 #(
		.INIT('h135f)
	) name119 (
		\InstQueue_reg[10][4]/NET0131 ,
		\InstQueue_reg[14][4]/NET0131 ,
		_w471_,
		_w476_,
		_w572_
	);
	LUT4 #(
		.INIT('h153f)
	) name120 (
		\InstQueue_reg[11][4]/NET0131 ,
		\InstQueue_reg[5][4]/NET0131 ,
		_w457_,
		_w458_,
		_w573_
	);
	LUT4 #(
		.INIT('h8000)
	) name121 (
		_w572_,
		_w573_,
		_w570_,
		_w571_,
		_w574_
	);
	LUT4 #(
		.INIT('h153f)
	) name122 (
		\InstQueue_reg[1][4]/NET0131 ,
		\InstQueue_reg[7][4]/NET0131 ,
		_w470_,
		_w473_,
		_w575_
	);
	LUT4 #(
		.INIT('h153f)
	) name123 (
		\InstQueue_reg[15][4]/NET0131 ,
		\InstQueue_reg[9][4]/NET0131 ,
		_w467_,
		_w455_,
		_w576_
	);
	LUT4 #(
		.INIT('h135f)
	) name124 (
		\InstQueue_reg[3][4]/NET0131 ,
		\InstQueue_reg[6][4]/NET0131 ,
		_w460_,
		_w453_,
		_w577_
	);
	LUT4 #(
		.INIT('h135f)
	) name125 (
		\InstQueue_reg[13][4]/NET0131 ,
		\InstQueue_reg[8][4]/NET0131 ,
		_w461_,
		_w463_,
		_w578_
	);
	LUT4 #(
		.INIT('h8000)
	) name126 (
		_w577_,
		_w578_,
		_w575_,
		_w576_,
		_w579_
	);
	LUT2 #(
		.INIT('h8)
	) name127 (
		_w574_,
		_w579_,
		_w580_
	);
	LUT4 #(
		.INIT('h8000)
	) name128 (
		_w574_,
		_w579_,
		_w523_,
		_w528_,
		_w581_
	);
	LUT4 #(
		.INIT('h8000)
	) name129 (
		_w567_,
		_w568_,
		_w581_,
		_w553_,
		_w582_
	);
	LUT4 #(
		.INIT('h0888)
	) name130 (
		_w574_,
		_w579_,
		_w523_,
		_w528_,
		_w583_
	);
	LUT4 #(
		.INIT('h0777)
	) name131 (
		_w534_,
		_w539_,
		_w546_,
		_w551_,
		_w584_
	);
	LUT2 #(
		.INIT('h8)
	) name132 (
		_w583_,
		_w584_,
		_w585_
	);
	LUT4 #(
		.INIT('h4000)
	) name133 (
		_w480_,
		_w583_,
		_w584_,
		_w517_,
		_w586_
	);
	LUT3 #(
		.INIT('h07)
	) name134 (
		_w494_,
		_w586_,
		_w582_,
		_w587_
	);
	LUT4 #(
		.INIT('h00f8)
	) name135 (
		_w494_,
		_w586_,
		_w582_,
		_w566_,
		_w588_
	);
	LUT4 #(
		.INIT('h8000)
	) name136 (
		_w567_,
		_w495_,
		_w581_,
		_w553_,
		_w589_
	);
	LUT3 #(
		.INIT('h10)
	) name137 (
		_w480_,
		_w494_,
		_w517_,
		_w590_
	);
	LUT3 #(
		.INIT('h13)
	) name138 (
		_w585_,
		_w589_,
		_w590_,
		_w591_
	);
	LUT3 #(
		.INIT('h04)
	) name139 (
		\State_reg[0]/NET0131 ,
		\State_reg[1]/NET0131 ,
		\State_reg[2]/NET0131 ,
		_w592_
	);
	LUT3 #(
		.INIT('h10)
	) name140 (
		\State_reg[0]/NET0131 ,
		\State_reg[1]/NET0131 ,
		\State_reg[2]/NET0131 ,
		_w593_
	);
	LUT3 #(
		.INIT('heb)
	) name141 (
		\State_reg[0]/NET0131 ,
		\State_reg[1]/NET0131 ,
		\State_reg[2]/NET0131 ,
		_w594_
	);
	LUT3 #(
		.INIT('h31)
	) name142 (
		_w563_,
		_w594_,
		_w565_,
		_w595_
	);
	LUT4 #(
		.INIT('hec00)
	) name143 (
		_w585_,
		_w589_,
		_w590_,
		_w595_,
		_w596_
	);
	LUT4 #(
		.INIT('h2223)
	) name144 (
		READY_n_pad,
		_w554_,
		_w588_,
		_w596_,
		_w597_
	);
	LUT3 #(
		.INIT('h54)
	) name145 (
		_w481_,
		_w588_,
		_w596_,
		_w598_
	);
	LUT3 #(
		.INIT('h78)
	) name146 (
		\InstQueueRd_Addr_reg[1]/NET0131 ,
		\InstQueueRd_Addr_reg[2]/NET0131 ,
		\InstQueueRd_Addr_reg[3]/NET0131 ,
		_w599_
	);
	LUT3 #(
		.INIT('hd0)
	) name147 (
		_w597_,
		_w598_,
		_w599_,
		_w600_
	);
	LUT4 #(
		.INIT('h0777)
	) name148 (
		_w574_,
		_w579_,
		_w546_,
		_w551_,
		_w601_
	);
	LUT3 #(
		.INIT('h40)
	) name149 (
		_w540_,
		_w529_,
		_w601_,
		_w602_
	);
	LUT4 #(
		.INIT('h0888)
	) name150 (
		_w500_,
		_w506_,
		_w511_,
		_w516_,
		_w603_
	);
	LUT2 #(
		.INIT('h8)
	) name151 (
		_w603_,
		_w495_,
		_w604_
	);
	LUT2 #(
		.INIT('h8)
	) name152 (
		_w602_,
		_w604_,
		_w605_
	);
	LUT3 #(
		.INIT('h37)
	) name153 (
		_w569_,
		_w602_,
		_w604_,
		_w606_
	);
	LUT4 #(
		.INIT('h8000)
	) name154 (
		_w567_,
		_w495_,
		_w583_,
		_w584_,
		_w607_
	);
	LUT4 #(
		.INIT('h8000)
	) name155 (
		_w567_,
		_w568_,
		_w583_,
		_w584_,
		_w608_
	);
	LUT2 #(
		.INIT('h1)
	) name156 (
		_w607_,
		_w608_,
		_w609_
	);
	LUT2 #(
		.INIT('h8)
	) name157 (
		_w606_,
		_w609_,
		_w610_
	);
	LUT3 #(
		.INIT('ha8)
	) name158 (
		READY_n_pad,
		_w588_,
		_w596_,
		_w611_
	);
	LUT4 #(
		.INIT('hf800)
	) name159 (
		_w494_,
		_w586_,
		_w582_,
		_w566_,
		_w612_
	);
	LUT3 #(
		.INIT('h31)
	) name160 (
		_w591_,
		_w595_,
		_w612_,
		_w613_
	);
	LUT4 #(
		.INIT('haaa2)
	) name161 (
		\InstQueueRd_Addr_reg[3]/NET0131 ,
		_w610_,
		_w611_,
		_w613_,
		_w614_
	);
	LUT4 #(
		.INIT('h0001)
	) name162 (
		_w586_,
		_w582_,
		_w589_,
		_w554_,
		_w615_
	);
	LUT3 #(
		.INIT('h80)
	) name163 (
		_w606_,
		_w609_,
		_w615_,
		_w616_
	);
	LUT3 #(
		.INIT('h80)
	) name164 (
		_w540_,
		_w552_,
		_w583_,
		_w617_
	);
	LUT4 #(
		.INIT('hfc7f)
	) name165 (
		_w540_,
		_w580_,
		_w552_,
		_w529_,
		_w618_
	);
	LUT2 #(
		.INIT('h2)
	) name166 (
		_w518_,
		_w618_,
		_w619_
	);
	LUT4 #(
		.INIT('h7000)
	) name167 (
		_w500_,
		_w506_,
		_w511_,
		_w516_,
		_w620_
	);
	LUT2 #(
		.INIT('h8)
	) name168 (
		_w568_,
		_w620_,
		_w621_
	);
	LUT2 #(
		.INIT('h8)
	) name169 (
		_w617_,
		_w621_,
		_w622_
	);
	LUT4 #(
		.INIT('h8000)
	) name170 (
		_w488_,
		_w493_,
		_w534_,
		_w539_,
		_w623_
	);
	LUT4 #(
		.INIT('h0888)
	) name171 (
		_w511_,
		_w516_,
		_w466_,
		_w479_,
		_w624_
	);
	LUT4 #(
		.INIT('h8000)
	) name172 (
		_w552_,
		_w581_,
		_w624_,
		_w623_,
		_w625_
	);
	LUT3 #(
		.INIT('h07)
	) name173 (
		_w617_,
		_w621_,
		_w625_,
		_w626_
	);
	LUT4 #(
		.INIT('h8000)
	) name174 (
		_w568_,
		_w603_,
		_w583_,
		_w584_,
		_w627_
	);
	LUT3 #(
		.INIT('h40)
	) name175 (
		_w540_,
		_w552_,
		_w583_,
		_w628_
	);
	LUT3 #(
		.INIT('h15)
	) name176 (
		_w627_,
		_w590_,
		_w628_,
		_w629_
	);
	LUT3 #(
		.INIT('h40)
	) name177 (
		_w619_,
		_w626_,
		_w629_,
		_w630_
	);
	LUT4 #(
		.INIT('h807f)
	) name178 (
		\InstQueueRd_Addr_reg[0]/NET0131 ,
		\InstQueueRd_Addr_reg[1]/NET0131 ,
		\InstQueueRd_Addr_reg[2]/NET0131 ,
		\InstQueueRd_Addr_reg[3]/NET0131 ,
		_w631_
	);
	LUT4 #(
		.INIT('h8421)
	) name179 (
		\InstQueueRd_Addr_reg[0]/NET0131 ,
		\InstQueueRd_Addr_reg[1]/NET0131 ,
		\InstQueueWr_Addr_reg[0]/NET0131 ,
		\InstQueueWr_Addr_reg[1]/NET0131 ,
		_w632_
	);
	LUT2 #(
		.INIT('h4)
	) name180 (
		_w558_,
		_w632_,
		_w633_
	);
	LUT2 #(
		.INIT('h1)
	) name181 (
		_w563_,
		_w633_,
		_w634_
	);
	LUT4 #(
		.INIT('hc800)
	) name182 (
		_w569_,
		_w602_,
		_w604_,
		_w634_,
		_w635_
	);
	LUT3 #(
		.INIT('h07)
	) name183 (
		\InstQueueRd_Addr_reg[0]/NET0131 ,
		\InstQueueRd_Addr_reg[1]/NET0131 ,
		\InstQueueRd_Addr_reg[2]/NET0131 ,
		_w636_
	);
	LUT2 #(
		.INIT('h2)
	) name184 (
		_w635_,
		_w636_,
		_w637_
	);
	LUT4 #(
		.INIT('h00f4)
	) name185 (
		_w616_,
		_w630_,
		_w631_,
		_w637_,
		_w638_
	);
	LUT3 #(
		.INIT('h10)
	) name186 (
		_w614_,
		_w600_,
		_w638_,
		_w639_
	);
	LUT4 #(
		.INIT('h0200)
	) name187 (
		\InstQueueWr_Addr_reg[3]/NET0131 ,
		_w614_,
		_w600_,
		_w638_,
		_w640_
	);
	LUT4 #(
		.INIT('h0100)
	) name188 (
		\InstQueueRd_Addr_reg[0]/NET0131 ,
		_w635_,
		_w616_,
		_w630_,
		_w641_
	);
	LUT4 #(
		.INIT('h00c8)
	) name189 (
		_w569_,
		_w602_,
		_w604_,
		_w634_,
		_w642_
	);
	LUT4 #(
		.INIT('h0080)
	) name190 (
		\InstQueueRd_Addr_reg[0]/NET0131 ,
		_w609_,
		_w615_,
		_w642_,
		_w643_
	);
	LUT3 #(
		.INIT('ha8)
	) name191 (
		\InstQueueWr_Addr_reg[0]/NET0131 ,
		_w641_,
		_w643_,
		_w644_
	);
	LUT4 #(
		.INIT('h0110)
	) name192 (
		READY_n_pad,
		\State_reg[0]/NET0131 ,
		\State_reg[1]/NET0131 ,
		\State_reg[2]/NET0131 ,
		_w645_
	);
	LUT4 #(
		.INIT('h00ec)
	) name193 (
		_w585_,
		_w589_,
		_w590_,
		_w566_,
		_w646_
	);
	LUT3 #(
		.INIT('h15)
	) name194 (
		_w554_,
		_w645_,
		_w646_,
		_w647_
	);
	LUT2 #(
		.INIT('h4)
	) name195 (
		READY_n_pad,
		_w588_,
		_w648_
	);
	LUT3 #(
		.INIT('h51)
	) name196 (
		\InstQueueRd_Addr_reg[1]/NET0131 ,
		_w647_,
		_w648_,
		_w649_
	);
	LUT2 #(
		.INIT('h9)
	) name197 (
		\InstQueueRd_Addr_reg[0]/NET0131 ,
		\InstQueueRd_Addr_reg[1]/NET0131 ,
		_w650_
	);
	LUT4 #(
		.INIT('h00ef)
	) name198 (
		_w635_,
		_w616_,
		_w630_,
		_w650_,
		_w651_
	);
	LUT3 #(
		.INIT('h51)
	) name199 (
		READY_n_pad,
		_w563_,
		_w565_,
		_w652_
	);
	LUT4 #(
		.INIT('h00f8)
	) name200 (
		_w494_,
		_w586_,
		_w582_,
		_w652_,
		_w653_
	);
	LUT3 #(
		.INIT('hc4)
	) name201 (
		_w563_,
		_w645_,
		_w565_,
		_w654_
	);
	LUT4 #(
		.INIT('h00ec)
	) name202 (
		_w585_,
		_w589_,
		_w590_,
		_w654_,
		_w655_
	);
	LUT4 #(
		.INIT('h0002)
	) name203 (
		_w609_,
		_w642_,
		_w653_,
		_w655_,
		_w656_
	);
	LUT2 #(
		.INIT('h2)
	) name204 (
		\InstQueueRd_Addr_reg[1]/NET0131 ,
		_w656_,
		_w657_
	);
	LUT3 #(
		.INIT('h01)
	) name205 (
		_w651_,
		_w649_,
		_w657_,
		_w658_
	);
	LUT2 #(
		.INIT('h6)
	) name206 (
		\InstQueueRd_Addr_reg[1]/NET0131 ,
		\InstQueueRd_Addr_reg[2]/NET0131 ,
		_w659_
	);
	LUT2 #(
		.INIT('h4)
	) name207 (
		_w597_,
		_w659_,
		_w660_
	);
	LUT3 #(
		.INIT('h78)
	) name208 (
		\InstQueueRd_Addr_reg[0]/NET0131 ,
		\InstQueueRd_Addr_reg[1]/NET0131 ,
		\InstQueueRd_Addr_reg[2]/NET0131 ,
		_w661_
	);
	LUT3 #(
		.INIT('hb0)
	) name209 (
		_w616_,
		_w630_,
		_w661_,
		_w662_
	);
	LUT2 #(
		.INIT('h2)
	) name210 (
		_w635_,
		_w661_,
		_w663_
	);
	LUT3 #(
		.INIT('h0d)
	) name211 (
		\InstQueueRd_Addr_reg[2]/NET0131 ,
		_w656_,
		_w663_,
		_w664_
	);
	LUT4 #(
		.INIT('h0200)
	) name212 (
		\InstQueueWr_Addr_reg[2]/NET0131 ,
		_w660_,
		_w662_,
		_w664_,
		_w665_
	);
	LUT4 #(
		.INIT('h0017)
	) name213 (
		\InstQueueWr_Addr_reg[1]/NET0131 ,
		_w644_,
		_w658_,
		_w665_,
		_w666_
	);
	LUT4 #(
		.INIT('h5455)
	) name214 (
		\InstQueueWr_Addr_reg[2]/NET0131 ,
		_w660_,
		_w662_,
		_w664_,
		_w667_
	);
	LUT4 #(
		.INIT('h0200)
	) name215 (
		\InstQueueWr_Addr_reg[3]/NET0131 ,
		_w660_,
		_w662_,
		_w664_,
		_w668_
	);
	LUT2 #(
		.INIT('h8)
	) name216 (
		READY_n_pad,
		_w588_,
		_w669_
	);
	LUT4 #(
		.INIT('h151f)
	) name217 (
		READY_n_pad,
		_w594_,
		_w646_,
		_w588_,
		_w670_
	);
	LUT2 #(
		.INIT('h8)
	) name218 (
		_w634_,
		_w607_,
		_w671_
	);
	LUT4 #(
		.INIT('h238c)
	) name219 (
		\InstQueueRd_Addr_reg[0]/NET0131 ,
		\InstQueueRd_Addr_reg[1]/NET0131 ,
		\InstQueueWr_Addr_reg[0]/NET0131 ,
		\InstQueueWr_Addr_reg[1]/NET0131 ,
		_w672_
	);
	LUT4 #(
		.INIT('h00e0)
	) name220 (
		_w555_,
		_w560_,
		_w564_,
		_w672_,
		_w673_
	);
	LUT2 #(
		.INIT('h2)
	) name221 (
		_w563_,
		_w673_,
		_w674_
	);
	LUT4 #(
		.INIT('h7707)
	) name222 (
		_w634_,
		_w607_,
		_w608_,
		_w674_,
		_w675_
	);
	LUT3 #(
		.INIT('hd0)
	) name223 (
		\Flush_reg/NET0131 ,
		_w670_,
		_w675_,
		_w676_
	);
	LUT3 #(
		.INIT('h51)
	) name224 (
		\More_reg/NET0131 ,
		_w563_,
		_w565_,
		_w677_
	);
	LUT3 #(
		.INIT('h0e)
	) name225 (
		_w653_,
		_w655_,
		_w677_,
		_w678_
	);
	LUT2 #(
		.INIT('h8)
	) name226 (
		_w608_,
		_w674_,
		_w679_
	);
	LUT2 #(
		.INIT('h4)
	) name227 (
		_w634_,
		_w607_,
		_w680_
	);
	LUT2 #(
		.INIT('h1)
	) name228 (
		_w642_,
		_w680_,
		_w681_
	);
	LUT3 #(
		.INIT('h01)
	) name229 (
		_w642_,
		_w679_,
		_w680_,
		_w682_
	);
	LUT2 #(
		.INIT('h4)
	) name230 (
		_w678_,
		_w682_,
		_w683_
	);
	LUT2 #(
		.INIT('h8)
	) name231 (
		_w676_,
		_w683_,
		_w684_
	);
	LUT3 #(
		.INIT('he0)
	) name232 (
		_w639_,
		_w668_,
		_w684_,
		_w685_
	);
	LUT4 #(
		.INIT('hab00)
	) name233 (
		_w640_,
		_w666_,
		_w667_,
		_w685_,
		_w686_
	);
	LUT2 #(
		.INIT('h2)
	) name234 (
		_w589_,
		_w566_,
		_w687_
	);
	LUT2 #(
		.INIT('h4)
	) name235 (
		\DataWidth_reg[1]/NET0131 ,
		_w645_,
		_w688_
	);
	LUT3 #(
		.INIT('h20)
	) name236 (
		_w589_,
		_w566_,
		_w688_,
		_w689_
	);
	LUT4 #(
		.INIT('h0020)
	) name237 (
		\State2_reg[0]/NET0131 ,
		\State2_reg[1]/NET0131 ,
		\State2_reg[2]/NET0131 ,
		\State2_reg[3]/NET0131 ,
		_w690_
	);
	LUT2 #(
		.INIT('h1)
	) name238 (
		\State2_reg[0]/NET0131 ,
		\State2_reg[3]/NET0131 ,
		_w691_
	);
	LUT3 #(
		.INIT('hf9)
	) name239 (
		\State2_reg[0]/NET0131 ,
		\State2_reg[2]/NET0131 ,
		\State2_reg[3]/NET0131 ,
		_w692_
	);
	LUT2 #(
		.INIT('h8)
	) name240 (
		READY_n_pad,
		\State2_reg[1]/NET0131 ,
		_w693_
	);
	LUT2 #(
		.INIT('h4)
	) name241 (
		_w692_,
		_w693_,
		_w694_
	);
	LUT4 #(
		.INIT('h0004)
	) name242 (
		\State2_reg[0]/NET0131 ,
		\State2_reg[1]/NET0131 ,
		\State2_reg[2]/NET0131 ,
		\State2_reg[3]/NET0131 ,
		_w695_
	);
	LUT4 #(
		.INIT('h0002)
	) name243 (
		\State2_reg[0]/NET0131 ,
		\State2_reg[1]/NET0131 ,
		\State2_reg[2]/NET0131 ,
		\State2_reg[3]/NET0131 ,
		_w696_
	);
	LUT4 #(
		.INIT('h8caf)
	) name244 (
		\DataWidth_reg[1]/NET0131 ,
		READY_n_pad,
		_w695_,
		_w696_,
		_w697_
	);
	LUT2 #(
		.INIT('h4)
	) name245 (
		_w694_,
		_w697_,
		_w698_
	);
	LUT4 #(
		.INIT('hd0ff)
	) name246 (
		_w686_,
		_w689_,
		_w690_,
		_w698_,
		_w699_
	);
	LUT4 #(
		.INIT('h0080)
	) name247 (
		\State2_reg[0]/NET0131 ,
		\State2_reg[1]/NET0131 ,
		\State2_reg[2]/NET0131 ,
		\State2_reg[3]/NET0131 ,
		_w700_
	);
	LUT2 #(
		.INIT('h4)
	) name248 (
		\Flush_reg/NET0131 ,
		\InstQueueRd_Addr_reg[2]/NET0131 ,
		_w701_
	);
	LUT3 #(
		.INIT('he0)
	) name249 (
		\InstQueueRd_Addr_reg[0]/NET0131 ,
		\InstQueueRd_Addr_reg[1]/NET0131 ,
		\InstQueueRd_Addr_reg[3]/NET0131 ,
		_w702_
	);
	LUT3 #(
		.INIT('h2a)
	) name250 (
		_w700_,
		_w701_,
		_w702_,
		_w703_
	);
	LUT4 #(
		.INIT('h0008)
	) name251 (
		READY_n_pad,
		\State2_reg[0]/NET0131 ,
		\State2_reg[2]/NET0131 ,
		\State2_reg[3]/NET0131 ,
		_w704_
	);
	LUT3 #(
		.INIT('h80)
	) name252 (
		READY_n_pad,
		\State2_reg[1]/NET0131 ,
		\State2_reg[2]/NET0131 ,
		_w705_
	);
	LUT4 #(
		.INIT('h0200)
	) name253 (
		\State2_reg[0]/NET0131 ,
		\State2_reg[1]/NET0131 ,
		\State2_reg[2]/NET0131 ,
		\State2_reg[3]/NET0131 ,
		_w706_
	);
	LUT4 #(
		.INIT('h000d)
	) name254 (
		_w691_,
		_w705_,
		_w706_,
		_w704_,
		_w707_
	);
	LUT2 #(
		.INIT('h4)
	) name255 (
		_w703_,
		_w707_,
		_w708_
	);
	LUT4 #(
		.INIT('h70ff)
	) name256 (
		_w686_,
		_w689_,
		_w690_,
		_w708_,
		_w709_
	);
	LUT4 #(
		.INIT('h0100)
	) name257 (
		\State2_reg[0]/NET0131 ,
		\State2_reg[1]/NET0131 ,
		\State2_reg[2]/NET0131 ,
		\State2_reg[3]/NET0131 ,
		_w710_
	);
	LUT4 #(
		.INIT('h0180)
	) name258 (
		\State2_reg[0]/NET0131 ,
		\State2_reg[1]/NET0131 ,
		\State2_reg[2]/NET0131 ,
		\State2_reg[3]/NET0131 ,
		_w711_
	);
	LUT4 #(
		.INIT('h0008)
	) name259 (
		\State2_reg[0]/NET0131 ,
		\State2_reg[1]/NET0131 ,
		\State2_reg[2]/NET0131 ,
		\State2_reg[3]/NET0131 ,
		_w712_
	);
	LUT2 #(
		.INIT('h4)
	) name260 (
		READY_n_pad,
		_w712_,
		_w713_
	);
	LUT2 #(
		.INIT('h8)
	) name261 (
		\DataWidth_reg[1]/NET0131 ,
		_w695_,
		_w714_
	);
	LUT4 #(
		.INIT('hff8f)
	) name262 (
		\State2_reg[0]/NET0131 ,
		\State2_reg[1]/NET0131 ,
		\State2_reg[2]/NET0131 ,
		\State2_reg[3]/NET0131 ,
		_w715_
	);
	LUT3 #(
		.INIT('h70)
	) name263 (
		\DataWidth_reg[1]/NET0131 ,
		_w695_,
		_w715_,
		_w716_
	);
	LUT2 #(
		.INIT('hb)
	) name264 (
		_w713_,
		_w716_,
		_w717_
	);
	LUT2 #(
		.INIT('h8)
	) name265 (
		\InstAddrPointer_reg[17]/NET0131 ,
		\InstAddrPointer_reg[18]/NET0131 ,
		_w718_
	);
	LUT3 #(
		.INIT('h80)
	) name266 (
		\InstAddrPointer_reg[17]/NET0131 ,
		\InstAddrPointer_reg[18]/NET0131 ,
		\InstAddrPointer_reg[19]/NET0131 ,
		_w719_
	);
	LUT2 #(
		.INIT('h8)
	) name267 (
		\InstAddrPointer_reg[6]/NET0131 ,
		\InstAddrPointer_reg[7]/NET0131 ,
		_w720_
	);
	LUT3 #(
		.INIT('h80)
	) name268 (
		\InstAddrPointer_reg[1]/NET0131 ,
		\InstAddrPointer_reg[2]/NET0131 ,
		\InstAddrPointer_reg[3]/NET0131 ,
		_w721_
	);
	LUT4 #(
		.INIT('h8000)
	) name269 (
		\InstAddrPointer_reg[1]/NET0131 ,
		\InstAddrPointer_reg[2]/NET0131 ,
		\InstAddrPointer_reg[3]/NET0131 ,
		\InstAddrPointer_reg[4]/NET0131 ,
		_w722_
	);
	LUT3 #(
		.INIT('h80)
	) name270 (
		\InstAddrPointer_reg[5]/NET0131 ,
		_w722_,
		_w720_,
		_w723_
	);
	LUT2 #(
		.INIT('h8)
	) name271 (
		\InstAddrPointer_reg[8]/NET0131 ,
		\InstAddrPointer_reg[9]/NET0131 ,
		_w724_
	);
	LUT3 #(
		.INIT('h80)
	) name272 (
		\InstAddrPointer_reg[10]/NET0131 ,
		\InstAddrPointer_reg[8]/NET0131 ,
		\InstAddrPointer_reg[9]/NET0131 ,
		_w725_
	);
	LUT4 #(
		.INIT('h8000)
	) name273 (
		\InstAddrPointer_reg[5]/NET0131 ,
		_w722_,
		_w720_,
		_w725_,
		_w726_
	);
	LUT2 #(
		.INIT('h8)
	) name274 (
		\InstAddrPointer_reg[11]/NET0131 ,
		\InstAddrPointer_reg[12]/NET0131 ,
		_w727_
	);
	LUT3 #(
		.INIT('h80)
	) name275 (
		\InstAddrPointer_reg[11]/NET0131 ,
		\InstAddrPointer_reg[12]/NET0131 ,
		\InstAddrPointer_reg[13]/NET0131 ,
		_w728_
	);
	LUT2 #(
		.INIT('h8)
	) name276 (
		_w726_,
		_w728_,
		_w729_
	);
	LUT2 #(
		.INIT('h8)
	) name277 (
		\InstAddrPointer_reg[14]/NET0131 ,
		\InstAddrPointer_reg[15]/NET0131 ,
		_w730_
	);
	LUT3 #(
		.INIT('h80)
	) name278 (
		\InstAddrPointer_reg[14]/NET0131 ,
		\InstAddrPointer_reg[15]/NET0131 ,
		\InstAddrPointer_reg[16]/NET0131 ,
		_w731_
	);
	LUT3 #(
		.INIT('h80)
	) name279 (
		_w726_,
		_w728_,
		_w731_,
		_w732_
	);
	LUT4 #(
		.INIT('h8000)
	) name280 (
		_w726_,
		_w728_,
		_w719_,
		_w731_,
		_w733_
	);
	LUT2 #(
		.INIT('h8)
	) name281 (
		\InstAddrPointer_reg[21]/NET0131 ,
		\InstAddrPointer_reg[22]/NET0131 ,
		_w734_
	);
	LUT3 #(
		.INIT('h80)
	) name282 (
		\InstAddrPointer_reg[21]/NET0131 ,
		\InstAddrPointer_reg[22]/NET0131 ,
		\InstAddrPointer_reg[23]/NET0131 ,
		_w735_
	);
	LUT4 #(
		.INIT('h8000)
	) name283 (
		\InstAddrPointer_reg[20]/NET0131 ,
		\InstAddrPointer_reg[21]/NET0131 ,
		\InstAddrPointer_reg[22]/NET0131 ,
		\InstAddrPointer_reg[23]/NET0131 ,
		_w736_
	);
	LUT3 #(
		.INIT('h80)
	) name284 (
		\InstAddrPointer_reg[24]/NET0131 ,
		_w733_,
		_w736_,
		_w737_
	);
	LUT4 #(
		.INIT('h8000)
	) name285 (
		\InstAddrPointer_reg[24]/NET0131 ,
		\InstAddrPointer_reg[25]/NET0131 ,
		_w733_,
		_w736_,
		_w738_
	);
	LUT2 #(
		.INIT('h8)
	) name286 (
		\InstAddrPointer_reg[26]/NET0131 ,
		\InstAddrPointer_reg[27]/NET0131 ,
		_w739_
	);
	LUT3 #(
		.INIT('h80)
	) name287 (
		\InstAddrPointer_reg[26]/NET0131 ,
		\InstAddrPointer_reg[27]/NET0131 ,
		\InstAddrPointer_reg[28]/NET0131 ,
		_w740_
	);
	LUT2 #(
		.INIT('h8)
	) name288 (
		_w738_,
		_w740_,
		_w741_
	);
	LUT3 #(
		.INIT('h80)
	) name289 (
		\InstAddrPointer_reg[29]/NET0131 ,
		_w738_,
		_w740_,
		_w742_
	);
	LUT4 #(
		.INIT('h8000)
	) name290 (
		\InstAddrPointer_reg[29]/NET0131 ,
		\InstAddrPointer_reg[30]/NET0131 ,
		_w738_,
		_w740_,
		_w743_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name291 (
		\InstAddrPointer_reg[29]/NET0131 ,
		\InstAddrPointer_reg[30]/NET0131 ,
		_w738_,
		_w740_,
		_w744_
	);
	LUT4 #(
		.INIT('h153f)
	) name292 (
		\InstQueue_reg[12][4]/NET0131 ,
		\InstQueue_reg[3][4]/NET0131 ,
		_w474_,
		_w458_,
		_w745_
	);
	LUT4 #(
		.INIT('h135f)
	) name293 (
		\InstQueue_reg[8][4]/NET0131 ,
		\InstQueue_reg[9][4]/NET0131 ,
		_w470_,
		_w463_,
		_w746_
	);
	LUT4 #(
		.INIT('h153f)
	) name294 (
		\InstQueue_reg[2][4]/NET0131 ,
		\InstQueue_reg[4][4]/NET0131 ,
		_w460_,
		_w473_,
		_w747_
	);
	LUT4 #(
		.INIT('h153f)
	) name295 (
		\InstQueue_reg[10][4]/NET0131 ,
		\InstQueue_reg[7][4]/NET0131 ,
		_w453_,
		_w467_,
		_w748_
	);
	LUT4 #(
		.INIT('h8000)
	) name296 (
		_w747_,
		_w748_,
		_w745_,
		_w746_,
		_w749_
	);
	LUT4 #(
		.INIT('h4000)
	) name297 (
		\InstQueueRd_Addr_reg[0]/NET0131 ,
		\InstQueueRd_Addr_reg[1]/NET0131 ,
		\InstQueueRd_Addr_reg[2]/NET0131 ,
		\InstQueue_reg[15][4]/NET0131 ,
		_w750_
	);
	LUT2 #(
		.INIT('h4)
	) name298 (
		_w631_,
		_w750_,
		_w751_
	);
	LUT4 #(
		.INIT('h135f)
	) name299 (
		\InstQueue_reg[11][4]/NET0131 ,
		\InstQueue_reg[5][4]/NET0131 ,
		_w471_,
		_w468_,
		_w752_
	);
	LUT4 #(
		.INIT('h135f)
	) name300 (
		\InstQueue_reg[14][4]/NET0131 ,
		\InstQueue_reg[6][4]/NET0131 ,
		_w461_,
		_w457_,
		_w753_
	);
	LUT3 #(
		.INIT('h40)
	) name301 (
		_w751_,
		_w752_,
		_w753_,
		_w754_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name302 (
		\InstQueueRd_Addr_reg[0]/NET0131 ,
		\InstQueueRd_Addr_reg[1]/NET0131 ,
		\InstQueue_reg[0][4]/NET0131 ,
		\InstQueue_reg[1][4]/NET0131 ,
		_w755_
	);
	LUT3 #(
		.INIT('h02)
	) name303 (
		_w631_,
		_w661_,
		_w755_,
		_w756_
	);
	LUT4 #(
		.INIT('h7800)
	) name304 (
		\InstQueueRd_Addr_reg[0]/NET0131 ,
		\InstQueueRd_Addr_reg[1]/NET0131 ,
		\InstQueueRd_Addr_reg[2]/NET0131 ,
		\InstQueueRd_Addr_reg[3]/NET0131 ,
		_w757_
	);
	LUT3 #(
		.INIT('h10)
	) name305 (
		\InstQueueRd_Addr_reg[0]/NET0131 ,
		\InstQueueRd_Addr_reg[1]/NET0131 ,
		\InstQueue_reg[13][4]/NET0131 ,
		_w758_
	);
	LUT2 #(
		.INIT('h8)
	) name306 (
		_w757_,
		_w758_,
		_w759_
	);
	LUT2 #(
		.INIT('h1)
	) name307 (
		_w756_,
		_w759_,
		_w760_
	);
	LUT3 #(
		.INIT('h80)
	) name308 (
		_w749_,
		_w754_,
		_w760_,
		_w761_
	);
	LUT4 #(
		.INIT('h7f80)
	) name309 (
		\InstAddrPointer_reg[1]/NET0131 ,
		\InstAddrPointer_reg[2]/NET0131 ,
		\InstAddrPointer_reg[3]/NET0131 ,
		\InstAddrPointer_reg[4]/NET0131 ,
		_w762_
	);
	LUT4 #(
		.INIT('h0080)
	) name310 (
		_w749_,
		_w754_,
		_w760_,
		_w762_,
		_w763_
	);
	LUT4 #(
		.INIT('h153f)
	) name311 (
		\InstQueue_reg[13][2]/NET0131 ,
		\InstQueue_reg[8][2]/NET0131 ,
		_w470_,
		_w477_,
		_w764_
	);
	LUT4 #(
		.INIT('h153f)
	) name312 (
		\InstQueue_reg[0][2]/NET0131 ,
		\InstQueue_reg[14][2]/NET0131 ,
		_w461_,
		_w455_,
		_w765_
	);
	LUT4 #(
		.INIT('h135f)
	) name313 (
		\InstQueue_reg[5][2]/NET0131 ,
		\InstQueue_reg[6][2]/NET0131 ,
		_w468_,
		_w457_,
		_w766_
	);
	LUT4 #(
		.INIT('h153f)
	) name314 (
		\InstQueue_reg[12][2]/NET0131 ,
		\InstQueue_reg[9][2]/NET0131 ,
		_w463_,
		_w458_,
		_w767_
	);
	LUT4 #(
		.INIT('h8000)
	) name315 (
		_w766_,
		_w767_,
		_w764_,
		_w765_,
		_w768_
	);
	LUT4 #(
		.INIT('h4000)
	) name316 (
		\InstQueueRd_Addr_reg[0]/NET0131 ,
		\InstQueueRd_Addr_reg[1]/NET0131 ,
		\InstQueueRd_Addr_reg[2]/NET0131 ,
		\InstQueue_reg[7][2]/NET0131 ,
		_w769_
	);
	LUT2 #(
		.INIT('h8)
	) name317 (
		_w631_,
		_w769_,
		_w770_
	);
	LUT2 #(
		.INIT('h8)
	) name318 (
		\InstQueue_reg[2][2]/NET0131 ,
		_w473_,
		_w771_
	);
	LUT4 #(
		.INIT('h153f)
	) name319 (
		\InstQueue_reg[10][2]/NET0131 ,
		\InstQueue_reg[3][2]/NET0131 ,
		_w474_,
		_w467_,
		_w772_
	);
	LUT4 #(
		.INIT('h135f)
	) name320 (
		\InstQueue_reg[1][2]/NET0131 ,
		\InstQueue_reg[4][2]/NET0131 ,
		_w464_,
		_w460_,
		_w773_
	);
	LUT4 #(
		.INIT('h135f)
	) name321 (
		\InstQueue_reg[11][2]/NET0131 ,
		\InstQueue_reg[15][2]/NET0131 ,
		_w471_,
		_w476_,
		_w774_
	);
	LUT4 #(
		.INIT('h4000)
	) name322 (
		_w771_,
		_w773_,
		_w774_,
		_w772_,
		_w775_
	);
	LUT3 #(
		.INIT('h40)
	) name323 (
		_w770_,
		_w768_,
		_w775_,
		_w776_
	);
	LUT2 #(
		.INIT('h6)
	) name324 (
		\InstAddrPointer_reg[1]/NET0131 ,
		\InstAddrPointer_reg[2]/NET0131 ,
		_w777_
	);
	LUT4 #(
		.INIT('h0040)
	) name325 (
		_w770_,
		_w768_,
		_w775_,
		_w777_,
		_w778_
	);
	LUT4 #(
		.INIT('h153f)
	) name326 (
		\InstQueue_reg[14][3]/NET0131 ,
		\InstQueue_reg[8][3]/NET0131 ,
		_w470_,
		_w461_,
		_w779_
	);
	LUT4 #(
		.INIT('h153f)
	) name327 (
		\InstQueue_reg[12][3]/NET0131 ,
		\InstQueue_reg[9][3]/NET0131 ,
		_w463_,
		_w458_,
		_w780_
	);
	LUT4 #(
		.INIT('h153f)
	) name328 (
		\InstQueue_reg[1][3]/NET0131 ,
		\InstQueue_reg[3][3]/NET0131 ,
		_w474_,
		_w464_,
		_w781_
	);
	LUT4 #(
		.INIT('h135f)
	) name329 (
		\InstQueue_reg[13][3]/NET0131 ,
		\InstQueue_reg[6][3]/NET0131 ,
		_w477_,
		_w457_,
		_w782_
	);
	LUT4 #(
		.INIT('h8000)
	) name330 (
		_w781_,
		_w782_,
		_w779_,
		_w780_,
		_w783_
	);
	LUT4 #(
		.INIT('h4000)
	) name331 (
		\InstQueueRd_Addr_reg[0]/NET0131 ,
		\InstQueueRd_Addr_reg[1]/NET0131 ,
		\InstQueueRd_Addr_reg[2]/NET0131 ,
		\InstQueue_reg[7][3]/NET0131 ,
		_w784_
	);
	LUT2 #(
		.INIT('h8)
	) name332 (
		_w631_,
		_w784_,
		_w785_
	);
	LUT2 #(
		.INIT('h8)
	) name333 (
		\InstQueue_reg[0][3]/NET0131 ,
		_w455_,
		_w786_
	);
	LUT4 #(
		.INIT('h135f)
	) name334 (
		\InstQueue_reg[11][3]/NET0131 ,
		\InstQueue_reg[15][3]/NET0131 ,
		_w471_,
		_w476_,
		_w787_
	);
	LUT4 #(
		.INIT('h153f)
	) name335 (
		\InstQueue_reg[2][3]/NET0131 ,
		\InstQueue_reg[4][3]/NET0131 ,
		_w460_,
		_w473_,
		_w788_
	);
	LUT4 #(
		.INIT('h153f)
	) name336 (
		\InstQueue_reg[10][3]/NET0131 ,
		\InstQueue_reg[5][3]/NET0131 ,
		_w468_,
		_w467_,
		_w789_
	);
	LUT4 #(
		.INIT('h4000)
	) name337 (
		_w786_,
		_w788_,
		_w789_,
		_w787_,
		_w790_
	);
	LUT3 #(
		.INIT('h40)
	) name338 (
		_w785_,
		_w783_,
		_w790_,
		_w791_
	);
	LUT3 #(
		.INIT('h78)
	) name339 (
		\InstAddrPointer_reg[1]/NET0131 ,
		\InstAddrPointer_reg[2]/NET0131 ,
		\InstAddrPointer_reg[3]/NET0131 ,
		_w792_
	);
	LUT4 #(
		.INIT('h0040)
	) name340 (
		_w785_,
		_w783_,
		_w790_,
		_w792_,
		_w793_
	);
	LUT2 #(
		.INIT('h1)
	) name341 (
		_w778_,
		_w793_,
		_w794_
	);
	LUT4 #(
		.INIT('hbf00)
	) name342 (
		_w770_,
		_w768_,
		_w775_,
		_w777_,
		_w795_
	);
	LUT4 #(
		.INIT('h135f)
	) name343 (
		\InstQueue_reg[13][1]/NET0131 ,
		\InstQueue_reg[6][1]/NET0131 ,
		_w477_,
		_w457_,
		_w796_
	);
	LUT4 #(
		.INIT('h153f)
	) name344 (
		\InstQueue_reg[0][1]/NET0131 ,
		\InstQueue_reg[11][1]/NET0131 ,
		_w471_,
		_w455_,
		_w797_
	);
	LUT4 #(
		.INIT('h153f)
	) name345 (
		\InstQueue_reg[12][1]/NET0131 ,
		\InstQueue_reg[9][1]/NET0131 ,
		_w463_,
		_w458_,
		_w798_
	);
	LUT4 #(
		.INIT('h135f)
	) name346 (
		\InstQueue_reg[1][1]/NET0131 ,
		\InstQueue_reg[4][1]/NET0131 ,
		_w464_,
		_w460_,
		_w799_
	);
	LUT4 #(
		.INIT('h8000)
	) name347 (
		_w798_,
		_w799_,
		_w796_,
		_w797_,
		_w800_
	);
	LUT4 #(
		.INIT('h153f)
	) name348 (
		\InstQueue_reg[3][1]/NET0131 ,
		\InstQueue_reg[8][1]/NET0131 ,
		_w470_,
		_w474_,
		_w801_
	);
	LUT4 #(
		.INIT('h135f)
	) name349 (
		\InstQueue_reg[14][1]/NET0131 ,
		\InstQueue_reg[5][1]/NET0131 ,
		_w461_,
		_w468_,
		_w802_
	);
	LUT4 #(
		.INIT('h135f)
	) name350 (
		\InstQueue_reg[15][1]/NET0131 ,
		\InstQueue_reg[2][1]/NET0131 ,
		_w476_,
		_w473_,
		_w803_
	);
	LUT4 #(
		.INIT('h153f)
	) name351 (
		\InstQueue_reg[10][1]/NET0131 ,
		\InstQueue_reg[7][1]/NET0131 ,
		_w453_,
		_w467_,
		_w804_
	);
	LUT4 #(
		.INIT('h8000)
	) name352 (
		_w803_,
		_w804_,
		_w801_,
		_w802_,
		_w805_
	);
	LUT2 #(
		.INIT('h8)
	) name353 (
		_w800_,
		_w805_,
		_w806_
	);
	LUT3 #(
		.INIT('h15)
	) name354 (
		\InstAddrPointer_reg[1]/NET0131 ,
		_w800_,
		_w805_,
		_w807_
	);
	LUT4 #(
		.INIT('h135f)
	) name355 (
		\InstQueue_reg[11][0]/NET0131 ,
		\InstQueue_reg[1][0]/NET0131 ,
		_w471_,
		_w464_,
		_w808_
	);
	LUT4 #(
		.INIT('h153f)
	) name356 (
		\InstQueue_reg[0][0]/NET0131 ,
		\InstQueue_reg[6][0]/NET0131 ,
		_w457_,
		_w455_,
		_w809_
	);
	LUT4 #(
		.INIT('h153f)
	) name357 (
		\InstQueue_reg[12][0]/NET0131 ,
		\InstQueue_reg[9][0]/NET0131 ,
		_w463_,
		_w458_,
		_w810_
	);
	LUT4 #(
		.INIT('h135f)
	) name358 (
		\InstQueue_reg[14][0]/NET0131 ,
		\InstQueue_reg[4][0]/NET0131 ,
		_w461_,
		_w460_,
		_w811_
	);
	LUT4 #(
		.INIT('h8000)
	) name359 (
		_w810_,
		_w811_,
		_w808_,
		_w809_,
		_w812_
	);
	LUT4 #(
		.INIT('h153f)
	) name360 (
		\InstQueue_reg[3][0]/NET0131 ,
		\InstQueue_reg[8][0]/NET0131 ,
		_w470_,
		_w474_,
		_w813_
	);
	LUT4 #(
		.INIT('h135f)
	) name361 (
		\InstQueue_reg[13][0]/NET0131 ,
		\InstQueue_reg[5][0]/NET0131 ,
		_w477_,
		_w468_,
		_w814_
	);
	LUT4 #(
		.INIT('h135f)
	) name362 (
		\InstQueue_reg[15][0]/NET0131 ,
		\InstQueue_reg[2][0]/NET0131 ,
		_w476_,
		_w473_,
		_w815_
	);
	LUT4 #(
		.INIT('h153f)
	) name363 (
		\InstQueue_reg[10][0]/NET0131 ,
		\InstQueue_reg[7][0]/NET0131 ,
		_w453_,
		_w467_,
		_w816_
	);
	LUT4 #(
		.INIT('h8000)
	) name364 (
		_w815_,
		_w816_,
		_w813_,
		_w814_,
		_w817_
	);
	LUT2 #(
		.INIT('h8)
	) name365 (
		_w812_,
		_w817_,
		_w818_
	);
	LUT3 #(
		.INIT('h2a)
	) name366 (
		\InstAddrPointer_reg[0]/NET0131 ,
		_w812_,
		_w817_,
		_w819_
	);
	LUT3 #(
		.INIT('h8e)
	) name367 (
		\InstAddrPointer_reg[1]/NET0131 ,
		_w806_,
		_w819_,
		_w820_
	);
	LUT4 #(
		.INIT('h080e)
	) name368 (
		\InstAddrPointer_reg[1]/NET0131 ,
		_w806_,
		_w795_,
		_w819_,
		_w821_
	);
	LUT4 #(
		.INIT('h7f00)
	) name369 (
		_w749_,
		_w754_,
		_w760_,
		_w762_,
		_w822_
	);
	LUT4 #(
		.INIT('hbf00)
	) name370 (
		_w785_,
		_w783_,
		_w790_,
		_w792_,
		_w823_
	);
	LUT2 #(
		.INIT('h1)
	) name371 (
		_w822_,
		_w823_,
		_w824_
	);
	LUT4 #(
		.INIT('h0455)
	) name372 (
		_w763_,
		_w794_,
		_w821_,
		_w824_,
		_w825_
	);
	LUT4 #(
		.INIT('h153f)
	) name373 (
		\InstQueue_reg[1][7]/NET0131 ,
		\InstQueue_reg[8][7]/NET0131 ,
		_w470_,
		_w464_,
		_w826_
	);
	LUT4 #(
		.INIT('h135f)
	) name374 (
		\InstQueue_reg[14][7]/NET0131 ,
		\InstQueue_reg[7][7]/NET0131 ,
		_w461_,
		_w453_,
		_w827_
	);
	LUT4 #(
		.INIT('h153f)
	) name375 (
		\InstQueue_reg[10][7]/NET0131 ,
		\InstQueue_reg[4][7]/NET0131 ,
		_w460_,
		_w467_,
		_w828_
	);
	LUT4 #(
		.INIT('h153f)
	) name376 (
		\InstQueue_reg[12][7]/NET0131 ,
		\InstQueue_reg[3][7]/NET0131 ,
		_w474_,
		_w458_,
		_w829_
	);
	LUT4 #(
		.INIT('h8000)
	) name377 (
		_w828_,
		_w829_,
		_w826_,
		_w827_,
		_w830_
	);
	LUT4 #(
		.INIT('h153f)
	) name378 (
		\InstQueue_reg[0][7]/NET0131 ,
		\InstQueue_reg[11][7]/NET0131 ,
		_w471_,
		_w455_,
		_w831_
	);
	LUT4 #(
		.INIT('h135f)
	) name379 (
		\InstQueue_reg[15][7]/NET0131 ,
		\InstQueue_reg[6][7]/NET0131 ,
		_w476_,
		_w457_,
		_w832_
	);
	LUT4 #(
		.INIT('h153f)
	) name380 (
		\InstQueue_reg[2][7]/NET0131 ,
		\InstQueue_reg[5][7]/NET0131 ,
		_w468_,
		_w473_,
		_w833_
	);
	LUT4 #(
		.INIT('h135f)
	) name381 (
		\InstQueue_reg[13][7]/NET0131 ,
		\InstQueue_reg[9][7]/NET0131 ,
		_w477_,
		_w463_,
		_w834_
	);
	LUT4 #(
		.INIT('h8000)
	) name382 (
		_w833_,
		_w834_,
		_w831_,
		_w832_,
		_w835_
	);
	LUT2 #(
		.INIT('h8)
	) name383 (
		_w830_,
		_w835_,
		_w836_
	);
	LUT4 #(
		.INIT('h78f0)
	) name384 (
		\InstAddrPointer_reg[5]/NET0131 ,
		\InstAddrPointer_reg[6]/NET0131 ,
		\InstAddrPointer_reg[7]/NET0131 ,
		_w722_,
		_w837_
	);
	LUT3 #(
		.INIT('h08)
	) name385 (
		_w830_,
		_w835_,
		_w837_,
		_w838_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name386 (
		\InstAddrPointer_reg[5]/NET0131 ,
		\InstAddrPointer_reg[8]/NET0131 ,
		_w722_,
		_w720_,
		_w839_
	);
	LUT4 #(
		.INIT('hf700)
	) name387 (
		_w830_,
		_w835_,
		_w837_,
		_w839_,
		_w840_
	);
	LUT4 #(
		.INIT('h153f)
	) name388 (
		\InstQueue_reg[0][6]/NET0131 ,
		\InstQueue_reg[14][6]/NET0131 ,
		_w461_,
		_w455_,
		_w841_
	);
	LUT4 #(
		.INIT('h135f)
	) name389 (
		\InstQueue_reg[8][6]/NET0131 ,
		\InstQueue_reg[9][6]/NET0131 ,
		_w470_,
		_w463_,
		_w842_
	);
	LUT4 #(
		.INIT('h135f)
	) name390 (
		\InstQueue_reg[15][6]/NET0131 ,
		\InstQueue_reg[6][6]/NET0131 ,
		_w476_,
		_w457_,
		_w843_
	);
	LUT3 #(
		.INIT('h80)
	) name391 (
		_w841_,
		_w842_,
		_w843_,
		_w844_
	);
	LUT4 #(
		.INIT('h153f)
	) name392 (
		\InstQueue_reg[10][6]/NET0131 ,
		\InstQueue_reg[11][6]/NET0131 ,
		_w471_,
		_w467_,
		_w845_
	);
	LUT4 #(
		.INIT('h153f)
	) name393 (
		\InstQueue_reg[12][6]/NET0131 ,
		\InstQueue_reg[2][6]/NET0131 ,
		_w473_,
		_w458_,
		_w846_
	);
	LUT4 #(
		.INIT('h153f)
	) name394 (
		\InstQueue_reg[1][6]/NET0131 ,
		\InstQueue_reg[3][6]/NET0131 ,
		_w474_,
		_w464_,
		_w847_
	);
	LUT4 #(
		.INIT('h153f)
	) name395 (
		\InstQueue_reg[4][6]/NET0131 ,
		\InstQueue_reg[5][6]/NET0131 ,
		_w468_,
		_w460_,
		_w848_
	);
	LUT4 #(
		.INIT('h8000)
	) name396 (
		_w847_,
		_w848_,
		_w845_,
		_w846_,
		_w849_
	);
	LUT4 #(
		.INIT('h4000)
	) name397 (
		\InstQueueRd_Addr_reg[0]/NET0131 ,
		\InstQueueRd_Addr_reg[1]/NET0131 ,
		\InstQueueRd_Addr_reg[2]/NET0131 ,
		\InstQueue_reg[7][6]/NET0131 ,
		_w850_
	);
	LUT3 #(
		.INIT('h10)
	) name398 (
		\InstQueueRd_Addr_reg[0]/NET0131 ,
		\InstQueueRd_Addr_reg[1]/NET0131 ,
		\InstQueue_reg[13][6]/NET0131 ,
		_w851_
	);
	LUT4 #(
		.INIT('h0777)
	) name399 (
		_w631_,
		_w850_,
		_w757_,
		_w851_,
		_w852_
	);
	LUT3 #(
		.INIT('h80)
	) name400 (
		_w844_,
		_w849_,
		_w852_,
		_w853_
	);
	LUT3 #(
		.INIT('h6c)
	) name401 (
		\InstAddrPointer_reg[5]/NET0131 ,
		\InstAddrPointer_reg[6]/NET0131 ,
		_w722_,
		_w854_
	);
	LUT4 #(
		.INIT('h0080)
	) name402 (
		_w844_,
		_w849_,
		_w852_,
		_w854_,
		_w855_
	);
	LUT4 #(
		.INIT('h153f)
	) name403 (
		\InstQueue_reg[0][5]/NET0131 ,
		\InstQueue_reg[8][5]/NET0131 ,
		_w470_,
		_w455_,
		_w856_
	);
	LUT4 #(
		.INIT('h153f)
	) name404 (
		\InstQueue_reg[10][5]/NET0131 ,
		\InstQueue_reg[4][5]/NET0131 ,
		_w460_,
		_w467_,
		_w857_
	);
	LUT4 #(
		.INIT('h153f)
	) name405 (
		\InstQueue_reg[12][5]/NET0131 ,
		\InstQueue_reg[7][5]/NET0131 ,
		_w453_,
		_w458_,
		_w858_
	);
	LUT4 #(
		.INIT('h153f)
	) name406 (
		\InstQueue_reg[6][5]/NET0131 ,
		\InstQueue_reg[9][5]/NET0131 ,
		_w463_,
		_w457_,
		_w859_
	);
	LUT4 #(
		.INIT('h8000)
	) name407 (
		_w858_,
		_w859_,
		_w856_,
		_w857_,
		_w860_
	);
	LUT4 #(
		.INIT('h135f)
	) name408 (
		\InstQueue_reg[11][5]/NET0131 ,
		\InstQueue_reg[1][5]/NET0131 ,
		_w471_,
		_w464_,
		_w861_
	);
	LUT4 #(
		.INIT('h135f)
	) name409 (
		\InstQueue_reg[3][5]/NET0131 ,
		\InstQueue_reg[5][5]/NET0131 ,
		_w474_,
		_w468_,
		_w862_
	);
	LUT4 #(
		.INIT('h135f)
	) name410 (
		\InstQueue_reg[14][5]/NET0131 ,
		\InstQueue_reg[2][5]/NET0131 ,
		_w461_,
		_w473_,
		_w863_
	);
	LUT4 #(
		.INIT('h135f)
	) name411 (
		\InstQueue_reg[13][5]/NET0131 ,
		\InstQueue_reg[15][5]/NET0131 ,
		_w477_,
		_w476_,
		_w864_
	);
	LUT4 #(
		.INIT('h8000)
	) name412 (
		_w863_,
		_w864_,
		_w861_,
		_w862_,
		_w865_
	);
	LUT2 #(
		.INIT('h8)
	) name413 (
		_w860_,
		_w865_,
		_w866_
	);
	LUT2 #(
		.INIT('h6)
	) name414 (
		\InstAddrPointer_reg[5]/NET0131 ,
		_w722_,
		_w867_
	);
	LUT3 #(
		.INIT('h08)
	) name415 (
		_w860_,
		_w865_,
		_w867_,
		_w868_
	);
	LUT2 #(
		.INIT('h1)
	) name416 (
		_w855_,
		_w868_,
		_w869_
	);
	LUT3 #(
		.INIT('h02)
	) name417 (
		_w840_,
		_w855_,
		_w868_,
		_w870_
	);
	LUT3 #(
		.INIT('h70)
	) name418 (
		_w830_,
		_w835_,
		_w837_,
		_w871_
	);
	LUT4 #(
		.INIT('h7f00)
	) name419 (
		_w844_,
		_w849_,
		_w852_,
		_w854_,
		_w872_
	);
	LUT3 #(
		.INIT('h70)
	) name420 (
		_w860_,
		_w865_,
		_w867_,
		_w873_
	);
	LUT3 #(
		.INIT('h23)
	) name421 (
		_w855_,
		_w872_,
		_w873_,
		_w874_
	);
	LUT4 #(
		.INIT('h020b)
	) name422 (
		_w853_,
		_w854_,
		_w871_,
		_w873_,
		_w875_
	);
	LUT2 #(
		.INIT('h2)
	) name423 (
		_w840_,
		_w875_,
		_w876_
	);
	LUT2 #(
		.INIT('h8)
	) name424 (
		\InstAddrPointer_reg[20]/NET0131 ,
		_w733_,
		_w877_
	);
	LUT2 #(
		.INIT('h6)
	) name425 (
		\InstAddrPointer_reg[20]/NET0131 ,
		_w733_,
		_w878_
	);
	LUT4 #(
		.INIT('h8000)
	) name426 (
		\InstAddrPointer_reg[17]/NET0131 ,
		_w726_,
		_w728_,
		_w731_,
		_w879_
	);
	LUT2 #(
		.INIT('h6)
	) name427 (
		\InstAddrPointer_reg[18]/NET0131 ,
		_w879_,
		_w880_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name428 (
		\InstAddrPointer_reg[14]/NET0131 ,
		\InstAddrPointer_reg[15]/NET0131 ,
		_w726_,
		_w728_,
		_w881_
	);
	LUT3 #(
		.INIT('h80)
	) name429 (
		\InstAddrPointer_reg[16]/NET0131 ,
		\InstAddrPointer_reg[17]/NET0131 ,
		_w881_,
		_w882_
	);
	LUT2 #(
		.INIT('h8)
	) name430 (
		_w880_,
		_w882_,
		_w883_
	);
	LUT4 #(
		.INIT('h78f0)
	) name431 (
		\InstAddrPointer_reg[17]/NET0131 ,
		\InstAddrPointer_reg[18]/NET0131 ,
		\InstAddrPointer_reg[19]/NET0131 ,
		_w732_,
		_w884_
	);
	LUT2 #(
		.INIT('h8)
	) name432 (
		\InstAddrPointer_reg[10]/NET0131 ,
		\InstAddrPointer_reg[11]/NET0131 ,
		_w885_
	);
	LUT3 #(
		.INIT('h6c)
	) name433 (
		\InstAddrPointer_reg[11]/NET0131 ,
		\InstAddrPointer_reg[12]/NET0131 ,
		_w726_,
		_w886_
	);
	LUT2 #(
		.INIT('h8)
	) name434 (
		\InstAddrPointer_reg[13]/NET0131 ,
		\InstAddrPointer_reg[14]/NET0131 ,
		_w887_
	);
	LUT4 #(
		.INIT('h6c00)
	) name435 (
		\InstAddrPointer_reg[11]/NET0131 ,
		\InstAddrPointer_reg[12]/NET0131 ,
		_w726_,
		_w887_,
		_w888_
	);
	LUT4 #(
		.INIT('h8000)
	) name436 (
		\InstAddrPointer_reg[5]/NET0131 ,
		_w722_,
		_w720_,
		_w724_,
		_w889_
	);
	LUT3 #(
		.INIT('h6c)
	) name437 (
		\InstAddrPointer_reg[8]/NET0131 ,
		\InstAddrPointer_reg[9]/NET0131 ,
		_w723_,
		_w890_
	);
	LUT3 #(
		.INIT('h80)
	) name438 (
		_w885_,
		_w888_,
		_w890_,
		_w891_
	);
	LUT4 #(
		.INIT('h8000)
	) name439 (
		_w884_,
		_w880_,
		_w882_,
		_w891_,
		_w892_
	);
	LUT2 #(
		.INIT('h8)
	) name440 (
		_w878_,
		_w892_,
		_w893_
	);
	LUT4 #(
		.INIT('hf800)
	) name441 (
		_w825_,
		_w870_,
		_w876_,
		_w893_,
		_w894_
	);
	LUT3 #(
		.INIT('h6c)
	) name442 (
		\InstAddrPointer_reg[20]/NET0131 ,
		\InstAddrPointer_reg[21]/NET0131 ,
		_w733_,
		_w895_
	);
	LUT4 #(
		.INIT('h60c0)
	) name443 (
		\InstAddrPointer_reg[20]/NET0131 ,
		\InstAddrPointer_reg[21]/NET0131 ,
		\InstAddrPointer_reg[22]/NET0131 ,
		_w733_,
		_w896_
	);
	LUT2 #(
		.INIT('h8)
	) name444 (
		\InstAddrPointer_reg[23]/NET0131 ,
		\InstAddrPointer_reg[24]/NET0131 ,
		_w897_
	);
	LUT3 #(
		.INIT('h80)
	) name445 (
		\InstAddrPointer_reg[23]/NET0131 ,
		\InstAddrPointer_reg[24]/NET0131 ,
		\InstAddrPointer_reg[25]/NET0131 ,
		_w898_
	);
	LUT4 #(
		.INIT('h8000)
	) name446 (
		\InstAddrPointer_reg[23]/NET0131 ,
		\InstAddrPointer_reg[24]/NET0131 ,
		\InstAddrPointer_reg[25]/NET0131 ,
		\InstAddrPointer_reg[26]/NET0131 ,
		_w899_
	);
	LUT4 #(
		.INIT('h8000)
	) name447 (
		\InstAddrPointer_reg[20]/NET0131 ,
		_w733_,
		_w734_,
		_w899_,
		_w900_
	);
	LUT4 #(
		.INIT('h7f4c)
	) name448 (
		\InstAddrPointer_reg[26]/NET0131 ,
		\InstAddrPointer_reg[27]/NET0131 ,
		_w738_,
		_w900_,
		_w901_
	);
	LUT3 #(
		.INIT('h6a)
	) name449 (
		\InstAddrPointer_reg[24]/NET0131 ,
		_w733_,
		_w736_,
		_w902_
	);
	LUT4 #(
		.INIT('h4888)
	) name450 (
		\InstAddrPointer_reg[24]/NET0131 ,
		\InstAddrPointer_reg[25]/NET0131 ,
		_w733_,
		_w736_,
		_w903_
	);
	LUT2 #(
		.INIT('h8)
	) name451 (
		\InstAddrPointer_reg[26]/NET0131 ,
		_w903_,
		_w904_
	);
	LUT2 #(
		.INIT('h8)
	) name452 (
		_w901_,
		_w904_,
		_w905_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name453 (
		\InstAddrPointer_reg[20]/NET0131 ,
		\InstAddrPointer_reg[23]/NET0131 ,
		_w733_,
		_w734_,
		_w906_
	);
	LUT2 #(
		.INIT('h8)
	) name454 (
		\InstAddrPointer_reg[28]/NET0131 ,
		_w906_,
		_w907_
	);
	LUT3 #(
		.INIT('h80)
	) name455 (
		_w901_,
		_w904_,
		_w907_,
		_w908_
	);
	LUT3 #(
		.INIT('h6a)
	) name456 (
		\InstAddrPointer_reg[29]/NET0131 ,
		_w738_,
		_w740_,
		_w909_
	);
	LUT4 #(
		.INIT('h8000)
	) name457 (
		_w901_,
		_w904_,
		_w907_,
		_w909_,
		_w910_
	);
	LUT4 #(
		.INIT('h007f)
	) name458 (
		_w894_,
		_w896_,
		_w910_,
		_w744_,
		_w911_
	);
	LUT2 #(
		.INIT('h8)
	) name459 (
		\InstAddrPointer_reg[30]/NET0131 ,
		_w910_,
		_w912_
	);
	LUT3 #(
		.INIT('h80)
	) name460 (
		_w894_,
		_w896_,
		_w912_,
		_w913_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name461 (
		_w836_,
		_w894_,
		_w896_,
		_w912_,
		_w914_
	);
	LUT2 #(
		.INIT('h4)
	) name462 (
		_w911_,
		_w914_,
		_w915_
	);
	LUT3 #(
		.INIT('h80)
	) name463 (
		\InstAddrPointer_reg[0]/NET0131 ,
		\InstAddrPointer_reg[5]/NET0131 ,
		_w722_,
		_w916_
	);
	LUT4 #(
		.INIT('h8000)
	) name464 (
		\InstAddrPointer_reg[0]/NET0131 ,
		\InstAddrPointer_reg[5]/NET0131 ,
		_w722_,
		_w720_,
		_w917_
	);
	LUT3 #(
		.INIT('h6c)
	) name465 (
		\InstAddrPointer_reg[6]/NET0131 ,
		\InstAddrPointer_reg[7]/NET0131 ,
		_w916_,
		_w918_
	);
	LUT3 #(
		.INIT('h40)
	) name466 (
		_w918_,
		_w830_,
		_w835_,
		_w919_
	);
	LUT4 #(
		.INIT('h78f0)
	) name467 (
		\InstAddrPointer_reg[0]/NET0131 ,
		\InstAddrPointer_reg[5]/NET0131 ,
		\InstAddrPointer_reg[6]/NET0131 ,
		_w722_,
		_w920_
	);
	LUT4 #(
		.INIT('h0080)
	) name468 (
		_w844_,
		_w849_,
		_w852_,
		_w920_,
		_w921_
	);
	LUT2 #(
		.INIT('h1)
	) name469 (
		_w919_,
		_w921_,
		_w922_
	);
	LUT4 #(
		.INIT('h7f00)
	) name470 (
		_w844_,
		_w849_,
		_w852_,
		_w920_,
		_w923_
	);
	LUT2 #(
		.INIT('h8)
	) name471 (
		\InstAddrPointer_reg[0]/NET0131 ,
		\InstAddrPointer_reg[1]/NET0131 ,
		_w924_
	);
	LUT4 #(
		.INIT('h8000)
	) name472 (
		\InstAddrPointer_reg[0]/NET0131 ,
		\InstAddrPointer_reg[1]/NET0131 ,
		\InstAddrPointer_reg[2]/NET0131 ,
		\InstAddrPointer_reg[3]/NET0131 ,
		_w925_
	);
	LUT4 #(
		.INIT('h7f80)
	) name473 (
		\InstAddrPointer_reg[0]/NET0131 ,
		\InstAddrPointer_reg[1]/NET0131 ,
		\InstAddrPointer_reg[2]/NET0131 ,
		\InstAddrPointer_reg[3]/NET0131 ,
		_w926_
	);
	LUT4 #(
		.INIT('h0040)
	) name474 (
		_w785_,
		_w783_,
		_w790_,
		_w926_,
		_w927_
	);
	LUT3 #(
		.INIT('h07)
	) name475 (
		\InstAddrPointer_reg[0]/NET0131 ,
		\InstAddrPointer_reg[1]/NET0131 ,
		\InstAddrPointer_reg[2]/NET0131 ,
		_w928_
	);
	LUT3 #(
		.INIT('h78)
	) name476 (
		\InstAddrPointer_reg[0]/NET0131 ,
		\InstAddrPointer_reg[1]/NET0131 ,
		\InstAddrPointer_reg[2]/NET0131 ,
		_w929_
	);
	LUT4 #(
		.INIT('h0040)
	) name477 (
		_w770_,
		_w768_,
		_w775_,
		_w929_,
		_w930_
	);
	LUT2 #(
		.INIT('h1)
	) name478 (
		_w927_,
		_w930_,
		_w931_
	);
	LUT2 #(
		.INIT('h6)
	) name479 (
		\InstAddrPointer_reg[0]/NET0131 ,
		\InstAddrPointer_reg[1]/NET0131 ,
		_w932_
	);
	LUT3 #(
		.INIT('h08)
	) name480 (
		_w800_,
		_w805_,
		_w932_,
		_w933_
	);
	LUT3 #(
		.INIT('h80)
	) name481 (
		\InstAddrPointer_reg[0]/NET0131 ,
		_w812_,
		_w817_,
		_w934_
	);
	LUT3 #(
		.INIT('h45)
	) name482 (
		_w933_,
		_w807_,
		_w934_,
		_w935_
	);
	LUT4 #(
		.INIT('hbf00)
	) name483 (
		_w785_,
		_w783_,
		_w790_,
		_w926_,
		_w936_
	);
	LUT4 #(
		.INIT('hbf00)
	) name484 (
		_w770_,
		_w768_,
		_w775_,
		_w929_,
		_w937_
	);
	LUT3 #(
		.INIT('h23)
	) name485 (
		_w927_,
		_w936_,
		_w937_,
		_w938_
	);
	LUT3 #(
		.INIT('h6c)
	) name486 (
		\InstAddrPointer_reg[0]/NET0131 ,
		\InstAddrPointer_reg[5]/NET0131 ,
		_w722_,
		_w939_
	);
	LUT3 #(
		.INIT('h40)
	) name487 (
		_w939_,
		_w860_,
		_w865_,
		_w940_
	);
	LUT4 #(
		.INIT('h7f4c)
	) name488 (
		\InstAddrPointer_reg[0]/NET0131 ,
		\InstAddrPointer_reg[4]/NET0131 ,
		_w721_,
		_w925_,
		_w941_
	);
	LUT4 #(
		.INIT('h0080)
	) name489 (
		_w749_,
		_w754_,
		_w760_,
		_w941_,
		_w942_
	);
	LUT2 #(
		.INIT('h1)
	) name490 (
		_w940_,
		_w942_,
		_w943_
	);
	LUT4 #(
		.INIT('h8f00)
	) name491 (
		_w931_,
		_w935_,
		_w938_,
		_w943_,
		_w944_
	);
	LUT3 #(
		.INIT('h2a)
	) name492 (
		_w939_,
		_w860_,
		_w865_,
		_w945_
	);
	LUT4 #(
		.INIT('h7f00)
	) name493 (
		_w749_,
		_w754_,
		_w760_,
		_w941_,
		_w946_
	);
	LUT3 #(
		.INIT('h23)
	) name494 (
		_w940_,
		_w945_,
		_w946_,
		_w947_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name495 (
		_w922_,
		_w923_,
		_w944_,
		_w947_,
		_w948_
	);
	LUT3 #(
		.INIT('h80)
	) name496 (
		\InstAddrPointer_reg[0]/NET0131 ,
		_w726_,
		_w727_,
		_w949_
	);
	LUT4 #(
		.INIT('h8000)
	) name497 (
		\InstAddrPointer_reg[10]/NET0131 ,
		\InstAddrPointer_reg[11]/NET0131 ,
		_w917_,
		_w724_,
		_w950_
	);
	LUT3 #(
		.INIT('h32)
	) name498 (
		\InstAddrPointer_reg[12]/NET0131 ,
		_w949_,
		_w950_,
		_w951_
	);
	LUT3 #(
		.INIT('h6c)
	) name499 (
		\InstAddrPointer_reg[8]/NET0131 ,
		\InstAddrPointer_reg[9]/NET0131 ,
		_w917_,
		_w952_
	);
	LUT3 #(
		.INIT('h6a)
	) name500 (
		\InstAddrPointer_reg[10]/NET0131 ,
		_w917_,
		_w724_,
		_w953_
	);
	LUT4 #(
		.INIT('h8105)
	) name501 (
		\InstAddrPointer_reg[10]/NET0131 ,
		\InstAddrPointer_reg[8]/NET0131 ,
		\InstAddrPointer_reg[9]/NET0131 ,
		_w917_,
		_w954_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name502 (
		\InstAddrPointer_reg[10]/NET0131 ,
		\InstAddrPointer_reg[11]/NET0131 ,
		_w917_,
		_w724_,
		_w955_
	);
	LUT2 #(
		.INIT('h2)
	) name503 (
		_w954_,
		_w955_,
		_w956_
	);
	LUT2 #(
		.INIT('h4)
	) name504 (
		_w951_,
		_w956_,
		_w957_
	);
	LUT2 #(
		.INIT('h6)
	) name505 (
		\InstAddrPointer_reg[8]/NET0131 ,
		_w917_,
		_w958_
	);
	LUT4 #(
		.INIT('h00d5)
	) name506 (
		_w918_,
		_w830_,
		_w835_,
		_w958_,
		_w959_
	);
	LUT3 #(
		.INIT('h80)
	) name507 (
		\InstAddrPointer_reg[0]/NET0131 ,
		_w726_,
		_w728_,
		_w960_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name508 (
		\InstAddrPointer_reg[0]/NET0131 ,
		\InstAddrPointer_reg[14]/NET0131 ,
		_w726_,
		_w728_,
		_w961_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name509 (
		\InstAddrPointer_reg[0]/NET0131 ,
		\InstAddrPointer_reg[13]/NET0131 ,
		_w726_,
		_w727_,
		_w962_
	);
	LUT2 #(
		.INIT('h1)
	) name510 (
		_w961_,
		_w962_,
		_w963_
	);
	LUT4 #(
		.INIT('h0800)
	) name511 (
		_w959_,
		_w963_,
		_w951_,
		_w956_,
		_w964_
	);
	LUT3 #(
		.INIT('h80)
	) name512 (
		\InstAddrPointer_reg[0]/NET0131 ,
		\InstAddrPointer_reg[20]/NET0131 ,
		_w733_,
		_w965_
	);
	LUT4 #(
		.INIT('h78f0)
	) name513 (
		\InstAddrPointer_reg[0]/NET0131 ,
		\InstAddrPointer_reg[20]/NET0131 ,
		\InstAddrPointer_reg[21]/NET0131 ,
		_w733_,
		_w966_
	);
	LUT2 #(
		.INIT('h8)
	) name514 (
		\InstAddrPointer_reg[0]/NET0131 ,
		_w733_,
		_w967_
	);
	LUT3 #(
		.INIT('h6c)
	) name515 (
		\InstAddrPointer_reg[0]/NET0131 ,
		\InstAddrPointer_reg[20]/NET0131 ,
		_w733_,
		_w968_
	);
	LUT4 #(
		.INIT('h8103)
	) name516 (
		\InstAddrPointer_reg[0]/NET0131 ,
		\InstAddrPointer_reg[20]/NET0131 ,
		\InstAddrPointer_reg[21]/NET0131 ,
		_w733_,
		_w969_
	);
	LUT3 #(
		.INIT('h6c)
	) name517 (
		\InstAddrPointer_reg[14]/NET0131 ,
		\InstAddrPointer_reg[15]/NET0131 ,
		_w960_,
		_w970_
	);
	LUT3 #(
		.INIT('h6a)
	) name518 (
		\InstAddrPointer_reg[16]/NET0131 ,
		_w960_,
		_w730_,
		_w971_
	);
	LUT4 #(
		.INIT('h8103)
	) name519 (
		\InstAddrPointer_reg[14]/NET0131 ,
		\InstAddrPointer_reg[15]/NET0131 ,
		\InstAddrPointer_reg[16]/NET0131 ,
		_w960_,
		_w972_
	);
	LUT4 #(
		.INIT('h070f)
	) name520 (
		\InstAddrPointer_reg[0]/NET0131 ,
		\InstAddrPointer_reg[18]/NET0131 ,
		\InstAddrPointer_reg[19]/NET0131 ,
		_w879_,
		_w973_
	);
	LUT2 #(
		.INIT('h1)
	) name521 (
		_w967_,
		_w973_,
		_w974_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name522 (
		\InstAddrPointer_reg[0]/NET0131 ,
		\InstAddrPointer_reg[17]/NET0131 ,
		_w729_,
		_w731_,
		_w975_
	);
	LUT3 #(
		.INIT('h6c)
	) name523 (
		\InstAddrPointer_reg[0]/NET0131 ,
		\InstAddrPointer_reg[18]/NET0131 ,
		_w879_,
		_w976_
	);
	LUT4 #(
		.INIT('h000e)
	) name524 (
		_w967_,
		_w973_,
		_w975_,
		_w976_,
		_w977_
	);
	LUT2 #(
		.INIT('h8)
	) name525 (
		_w972_,
		_w977_,
		_w978_
	);
	LUT3 #(
		.INIT('h80)
	) name526 (
		_w969_,
		_w972_,
		_w977_,
		_w979_
	);
	LUT3 #(
		.INIT('h40)
	) name527 (
		_w948_,
		_w964_,
		_w979_,
		_w980_
	);
	LUT4 #(
		.INIT('h8000)
	) name528 (
		\InstAddrPointer_reg[0]/NET0131 ,
		\InstAddrPointer_reg[20]/NET0131 ,
		_w733_,
		_w734_,
		_w981_
	);
	LUT3 #(
		.INIT('h80)
	) name529 (
		\InstAddrPointer_reg[0]/NET0131 ,
		_w733_,
		_w736_,
		_w982_
	);
	LUT3 #(
		.INIT('h0e)
	) name530 (
		\InstAddrPointer_reg[23]/NET0131 ,
		_w981_,
		_w982_,
		_w983_
	);
	LUT4 #(
		.INIT('h1333)
	) name531 (
		\InstAddrPointer_reg[0]/NET0131 ,
		\InstAddrPointer_reg[24]/NET0131 ,
		_w733_,
		_w736_,
		_w984_
	);
	LUT3 #(
		.INIT('h13)
	) name532 (
		_w981_,
		_w984_,
		_w897_,
		_w985_
	);
	LUT4 #(
		.INIT('h8001)
	) name533 (
		\InstAddrPointer_reg[23]/NET0131 ,
		\InstAddrPointer_reg[24]/NET0131 ,
		_w981_,
		_w982_,
		_w986_
	);
	LUT3 #(
		.INIT('h6c)
	) name534 (
		\InstAddrPointer_reg[21]/NET0131 ,
		\InstAddrPointer_reg[22]/NET0131 ,
		_w965_,
		_w987_
	);
	LUT2 #(
		.INIT('h2)
	) name535 (
		_w986_,
		_w987_,
		_w988_
	);
	LUT3 #(
		.INIT('h6a)
	) name536 (
		\InstAddrPointer_reg[25]/NET0131 ,
		_w981_,
		_w897_,
		_w989_
	);
	LUT3 #(
		.INIT('h02)
	) name537 (
		_w986_,
		_w987_,
		_w989_,
		_w990_
	);
	LUT4 #(
		.INIT('h4000)
	) name538 (
		_w948_,
		_w964_,
		_w979_,
		_w990_,
		_w991_
	);
	LUT3 #(
		.INIT('h15)
	) name539 (
		\InstAddrPointer_reg[27]/NET0131 ,
		_w981_,
		_w899_,
		_w992_
	);
	LUT3 #(
		.INIT('h80)
	) name540 (
		_w981_,
		_w898_,
		_w739_,
		_w993_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name541 (
		\InstAddrPointer_reg[26]/NET0131 ,
		\InstAddrPointer_reg[27]/NET0131 ,
		_w981_,
		_w898_,
		_w994_
	);
	LUT4 #(
		.INIT('h8000)
	) name542 (
		\InstAddrPointer_reg[28]/NET0131 ,
		_w981_,
		_w898_,
		_w739_,
		_w995_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name543 (
		\InstAddrPointer_reg[28]/NET0131 ,
		_w981_,
		_w898_,
		_w739_,
		_w996_
	);
	LUT2 #(
		.INIT('h6)
	) name544 (
		\InstAddrPointer_reg[29]/NET0131 ,
		_w995_,
		_w997_
	);
	LUT4 #(
		.INIT('h8810)
	) name545 (
		\InstAddrPointer_reg[28]/NET0131 ,
		\InstAddrPointer_reg[29]/NET0131 ,
		_w992_,
		_w993_,
		_w998_
	);
	LUT3 #(
		.INIT('h6a)
	) name546 (
		\InstAddrPointer_reg[26]/NET0131 ,
		_w981_,
		_w898_,
		_w999_
	);
	LUT2 #(
		.INIT('h2)
	) name547 (
		_w998_,
		_w999_,
		_w1000_
	);
	LUT3 #(
		.INIT('h6c)
	) name548 (
		\InstAddrPointer_reg[29]/NET0131 ,
		\InstAddrPointer_reg[30]/NET0131 ,
		_w995_,
		_w1001_
	);
	LUT4 #(
		.INIT('heabf)
	) name549 (
		_w836_,
		_w991_,
		_w1000_,
		_w1001_,
		_w1002_
	);
	LUT4 #(
		.INIT('h4744)
	) name550 (
		\InstAddrPointer_reg[30]/NET0131 ,
		_w674_,
		_w915_,
		_w1002_,
		_w1003_
	);
	LUT4 #(
		.INIT('hf800)
	) name551 (
		\InstAddrPointer_reg[0]/NET0131 ,
		\InstAddrPointer_reg[1]/NET0131 ,
		\InstAddrPointer_reg[2]/NET0131 ,
		\InstAddrPointer_reg[3]/NET0131 ,
		_w1004_
	);
	LUT4 #(
		.INIT('h8000)
	) name552 (
		\InstAddrPointer_reg[4]/NET0131 ,
		\InstAddrPointer_reg[5]/NET0131 ,
		\InstAddrPointer_reg[6]/NET0131 ,
		_w1004_,
		_w1005_
	);
	LUT3 #(
		.INIT('h80)
	) name553 (
		\InstAddrPointer_reg[7]/NET0131 ,
		_w725_,
		_w1005_,
		_w1006_
	);
	LUT4 #(
		.INIT('h8000)
	) name554 (
		\InstAddrPointer_reg[7]/NET0131 ,
		_w725_,
		_w728_,
		_w1005_,
		_w1007_
	);
	LUT3 #(
		.INIT('h80)
	) name555 (
		_w719_,
		_w731_,
		_w1007_,
		_w1008_
	);
	LUT4 #(
		.INIT('h8000)
	) name556 (
		\InstAddrPointer_reg[20]/NET0131 ,
		_w719_,
		_w731_,
		_w1007_,
		_w1009_
	);
	LUT4 #(
		.INIT('h8000)
	) name557 (
		\InstAddrPointer_reg[24]/NET0131 ,
		\InstAddrPointer_reg[25]/NET0131 ,
		_w735_,
		_w1009_,
		_w1010_
	);
	LUT3 #(
		.INIT('h80)
	) name558 (
		_w734_,
		_w899_,
		_w1009_,
		_w1011_
	);
	LUT3 #(
		.INIT('h0e)
	) name559 (
		\InstAddrPointer_reg[26]/NET0131 ,
		_w1010_,
		_w1011_,
		_w1012_
	);
	LUT2 #(
		.INIT('h6)
	) name560 (
		\InstAddrPointer_reg[7]/NET0131 ,
		_w1005_,
		_w1013_
	);
	LUT3 #(
		.INIT('h08)
	) name561 (
		_w830_,
		_w835_,
		_w1013_,
		_w1014_
	);
	LUT3 #(
		.INIT('h6c)
	) name562 (
		\InstAddrPointer_reg[7]/NET0131 ,
		\InstAddrPointer_reg[8]/NET0131 ,
		_w1005_,
		_w1015_
	);
	LUT4 #(
		.INIT('hf700)
	) name563 (
		_w830_,
		_w835_,
		_w1013_,
		_w1015_,
		_w1016_
	);
	LUT4 #(
		.INIT('h78f0)
	) name564 (
		\InstAddrPointer_reg[4]/NET0131 ,
		\InstAddrPointer_reg[5]/NET0131 ,
		\InstAddrPointer_reg[6]/NET0131 ,
		_w1004_,
		_w1017_
	);
	LUT4 #(
		.INIT('h0080)
	) name565 (
		_w844_,
		_w849_,
		_w852_,
		_w1017_,
		_w1018_
	);
	LUT3 #(
		.INIT('h6c)
	) name566 (
		\InstAddrPointer_reg[4]/NET0131 ,
		\InstAddrPointer_reg[5]/NET0131 ,
		_w1004_,
		_w1019_
	);
	LUT3 #(
		.INIT('h08)
	) name567 (
		_w860_,
		_w865_,
		_w1019_,
		_w1020_
	);
	LUT2 #(
		.INIT('h1)
	) name568 (
		_w1018_,
		_w1020_,
		_w1021_
	);
	LUT2 #(
		.INIT('h6)
	) name569 (
		\InstAddrPointer_reg[4]/NET0131 ,
		_w1004_,
		_w1022_
	);
	LUT4 #(
		.INIT('h0080)
	) name570 (
		_w749_,
		_w754_,
		_w760_,
		_w1022_,
		_w1023_
	);
	LUT4 #(
		.INIT('h07f8)
	) name571 (
		\InstAddrPointer_reg[0]/NET0131 ,
		\InstAddrPointer_reg[1]/NET0131 ,
		\InstAddrPointer_reg[2]/NET0131 ,
		\InstAddrPointer_reg[3]/NET0131 ,
		_w1024_
	);
	LUT4 #(
		.INIT('h0040)
	) name572 (
		_w785_,
		_w783_,
		_w790_,
		_w1024_,
		_w1025_
	);
	LUT2 #(
		.INIT('h1)
	) name573 (
		_w1023_,
		_w1025_,
		_w1026_
	);
	LUT4 #(
		.INIT('hbf00)
	) name574 (
		_w785_,
		_w783_,
		_w790_,
		_w1024_,
		_w1027_
	);
	LUT4 #(
		.INIT('h4000)
	) name575 (
		_w770_,
		_w768_,
		_w775_,
		_w929_,
		_w1028_
	);
	LUT4 #(
		.INIT('h00bf)
	) name576 (
		_w770_,
		_w768_,
		_w775_,
		_w929_,
		_w1029_
	);
	LUT3 #(
		.INIT('h15)
	) name577 (
		\InstAddrPointer_reg[0]/NET0131 ,
		_w812_,
		_w817_,
		_w1030_
	);
	LUT4 #(
		.INIT('h020b)
	) name578 (
		_w806_,
		_w932_,
		_w1029_,
		_w1030_,
		_w1031_
	);
	LUT4 #(
		.INIT('h888a)
	) name579 (
		_w1026_,
		_w1027_,
		_w1028_,
		_w1031_,
		_w1032_
	);
	LUT4 #(
		.INIT('h7f00)
	) name580 (
		_w749_,
		_w754_,
		_w760_,
		_w1022_,
		_w1033_
	);
	LUT3 #(
		.INIT('h70)
	) name581 (
		_w860_,
		_w865_,
		_w1019_,
		_w1034_
	);
	LUT2 #(
		.INIT('h1)
	) name582 (
		_w1033_,
		_w1034_,
		_w1035_
	);
	LUT4 #(
		.INIT('h7f00)
	) name583 (
		_w844_,
		_w849_,
		_w852_,
		_w1017_,
		_w1036_
	);
	LUT3 #(
		.INIT('h70)
	) name584 (
		_w830_,
		_w835_,
		_w1013_,
		_w1037_
	);
	LUT2 #(
		.INIT('h1)
	) name585 (
		_w1036_,
		_w1037_,
		_w1038_
	);
	LUT4 #(
		.INIT('h7500)
	) name586 (
		_w1021_,
		_w1032_,
		_w1035_,
		_w1038_,
		_w1039_
	);
	LUT3 #(
		.INIT('h6a)
	) name587 (
		\InstAddrPointer_reg[17]/NET0131 ,
		_w731_,
		_w1007_,
		_w1040_
	);
	LUT4 #(
		.INIT('h8000)
	) name588 (
		\InstAddrPointer_reg[7]/NET0131 ,
		\InstAddrPointer_reg[8]/NET0131 ,
		\InstAddrPointer_reg[9]/NET0131 ,
		_w1005_,
		_w1041_
	);
	LUT3 #(
		.INIT('h6a)
	) name589 (
		\InstAddrPointer_reg[12]/NET0131 ,
		_w885_,
		_w1041_,
		_w1042_
	);
	LUT4 #(
		.INIT('h4888)
	) name590 (
		\InstAddrPointer_reg[12]/NET0131 ,
		\InstAddrPointer_reg[13]/NET0131 ,
		_w885_,
		_w1041_,
		_w1043_
	);
	LUT4 #(
		.INIT('h78f0)
	) name591 (
		\InstAddrPointer_reg[7]/NET0131 ,
		\InstAddrPointer_reg[8]/NET0131 ,
		\InstAddrPointer_reg[9]/NET0131 ,
		_w1005_,
		_w1044_
	);
	LUT2 #(
		.INIT('h8)
	) name592 (
		\InstAddrPointer_reg[10]/NET0131 ,
		_w1044_,
		_w1045_
	);
	LUT3 #(
		.INIT('h80)
	) name593 (
		\InstAddrPointer_reg[10]/NET0131 ,
		\InstAddrPointer_reg[14]/NET0131 ,
		_w1044_,
		_w1046_
	);
	LUT4 #(
		.INIT('ha8a0)
	) name594 (
		\InstAddrPointer_reg[11]/NET0131 ,
		\InstAddrPointer_reg[14]/NET0131 ,
		\InstAddrPointer_reg[15]/NET0131 ,
		_w1007_,
		_w1047_
	);
	LUT3 #(
		.INIT('h80)
	) name595 (
		_w1043_,
		_w1046_,
		_w1047_,
		_w1048_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name596 (
		\InstAddrPointer_reg[16]/NET0131 ,
		\InstAddrPointer_reg[7]/NET0131 ,
		_w725_,
		_w1005_,
		_w1049_
	);
	LUT4 #(
		.INIT('h8000)
	) name597 (
		_w1043_,
		_w1046_,
		_w1047_,
		_w1049_,
		_w1050_
	);
	LUT2 #(
		.INIT('h8)
	) name598 (
		_w1040_,
		_w1050_,
		_w1051_
	);
	LUT3 #(
		.INIT('h20)
	) name599 (
		_w1016_,
		_w1039_,
		_w1051_,
		_w1052_
	);
	LUT4 #(
		.INIT('h8000)
	) name600 (
		\InstAddrPointer_reg[17]/NET0131 ,
		\InstAddrPointer_reg[18]/NET0131 ,
		_w731_,
		_w1007_,
		_w1053_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name601 (
		\InstAddrPointer_reg[17]/NET0131 ,
		\InstAddrPointer_reg[18]/NET0131 ,
		_w731_,
		_w1007_,
		_w1054_
	);
	LUT4 #(
		.INIT('h2000)
	) name602 (
		_w1016_,
		_w1039_,
		_w1051_,
		_w1054_,
		_w1055_
	);
	LUT2 #(
		.INIT('h6)
	) name603 (
		\InstAddrPointer_reg[21]/NET0131 ,
		_w1009_,
		_w1056_
	);
	LUT3 #(
		.INIT('h48)
	) name604 (
		\InstAddrPointer_reg[21]/NET0131 ,
		\InstAddrPointer_reg[22]/NET0131 ,
		_w1009_,
		_w1057_
	);
	LUT4 #(
		.INIT('h4080)
	) name605 (
		\InstAddrPointer_reg[21]/NET0131 ,
		\InstAddrPointer_reg[22]/NET0131 ,
		\InstAddrPointer_reg[23]/NET0131 ,
		_w1009_,
		_w1058_
	);
	LUT3 #(
		.INIT('h6a)
	) name606 (
		\InstAddrPointer_reg[24]/NET0131 ,
		_w735_,
		_w1009_,
		_w1059_
	);
	LUT2 #(
		.INIT('h8)
	) name607 (
		_w1058_,
		_w1059_,
		_w1060_
	);
	LUT3 #(
		.INIT('h32)
	) name608 (
		\InstAddrPointer_reg[19]/NET0131 ,
		_w1008_,
		_w1053_,
		_w1061_
	);
	LUT4 #(
		.INIT('h0c08)
	) name609 (
		\InstAddrPointer_reg[19]/NET0131 ,
		\InstAddrPointer_reg[20]/NET0131 ,
		_w1008_,
		_w1053_,
		_w1062_
	);
	LUT4 #(
		.INIT('h8000)
	) name610 (
		\InstAddrPointer_reg[25]/NET0131 ,
		_w1058_,
		_w1059_,
		_w1062_,
		_w1063_
	);
	LUT3 #(
		.INIT('h80)
	) name611 (
		_w1012_,
		_w1055_,
		_w1063_,
		_w1064_
	);
	LUT4 #(
		.INIT('h8000)
	) name612 (
		\InstAddrPointer_reg[27]/NET0131 ,
		_w734_,
		_w899_,
		_w1009_,
		_w1065_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name613 (
		\InstAddrPointer_reg[27]/NET0131 ,
		_w734_,
		_w899_,
		_w1009_,
		_w1066_
	);
	LUT3 #(
		.INIT('h80)
	) name614 (
		\InstAddrPointer_reg[28]/NET0131 ,
		\InstAddrPointer_reg[29]/NET0131 ,
		_w1066_,
		_w1067_
	);
	LUT4 #(
		.INIT('h8000)
	) name615 (
		\InstAddrPointer_reg[29]/NET0131 ,
		\InstAddrPointer_reg[30]/NET0131 ,
		_w740_,
		_w1010_,
		_w1068_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name616 (
		\InstAddrPointer_reg[29]/NET0131 ,
		\InstAddrPointer_reg[30]/NET0131 ,
		_w740_,
		_w1010_,
		_w1069_
	);
	LUT4 #(
		.INIT('h2a80)
	) name617 (
		_w671_,
		_w1064_,
		_w1067_,
		_w1069_,
		_w1070_
	);
	LUT2 #(
		.INIT('h8)
	) name618 (
		_w635_,
		_w1069_,
		_w1071_
	);
	LUT3 #(
		.INIT('hb0)
	) name619 (
		_w616_,
		_w630_,
		_w1001_,
		_w1072_
	);
	LUT4 #(
		.INIT('hec00)
	) name620 (
		_w585_,
		_w589_,
		_w590_,
		_w594_,
		_w1073_
	);
	LUT3 #(
		.INIT('h01)
	) name621 (
		_w642_,
		_w680_,
		_w1073_,
		_w1074_
	);
	LUT4 #(
		.INIT('h00fe)
	) name622 (
		_w586_,
		_w582_,
		_w589_,
		_w652_,
		_w1075_
	);
	LUT4 #(
		.INIT('h0001)
	) name623 (
		_w642_,
		_w680_,
		_w1073_,
		_w1075_,
		_w1076_
	);
	LUT4 #(
		.INIT('hed45)
	) name624 (
		\InstAddrPointer_reg[30]/NET0131 ,
		_w597_,
		_w742_,
		_w1076_,
		_w1077_
	);
	LUT3 #(
		.INIT('h10)
	) name625 (
		_w1072_,
		_w1071_,
		_w1077_,
		_w1078_
	);
	LUT4 #(
		.INIT('h0d00)
	) name626 (
		_w608_,
		_w1003_,
		_w1070_,
		_w1078_,
		_w1079_
	);
	LUT4 #(
		.INIT('h0001)
	) name627 (
		\State2_reg[0]/NET0131 ,
		\State2_reg[1]/NET0131 ,
		\State2_reg[2]/NET0131 ,
		\State2_reg[3]/NET0131 ,
		_w1080_
	);
	LUT4 #(
		.INIT('h03de)
	) name628 (
		\State2_reg[0]/NET0131 ,
		\State2_reg[1]/NET0131 ,
		\State2_reg[2]/NET0131 ,
		\State2_reg[3]/NET0131 ,
		_w1081_
	);
	LUT4 #(
		.INIT('h153f)
	) name629 (
		\InstAddrPointer_reg[30]/NET0131 ,
		\rEIP_reg[30]/NET0131 ,
		_w1080_,
		_w1081_,
		_w1082_
	);
	LUT3 #(
		.INIT('h2f)
	) name630 (
		_w690_,
		_w1079_,
		_w1082_,
		_w1083_
	);
	LUT3 #(
		.INIT('h08)
	) name631 (
		\InstAddrPointer_reg[29]/NET0131 ,
		_w563_,
		_w673_,
		_w1084_
	);
	LUT4 #(
		.INIT('h00ba)
	) name632 (
		_w933_,
		_w807_,
		_w934_,
		_w937_,
		_w1085_
	);
	LUT3 #(
		.INIT('h01)
	) name633 (
		_w942_,
		_w927_,
		_w930_,
		_w1086_
	);
	LUT3 #(
		.INIT('h0b)
	) name634 (
		_w942_,
		_w936_,
		_w946_,
		_w1087_
	);
	LUT3 #(
		.INIT('h01)
	) name635 (
		_w919_,
		_w921_,
		_w940_,
		_w1088_
	);
	LUT4 #(
		.INIT('h4f00)
	) name636 (
		_w1085_,
		_w1086_,
		_w1087_,
		_w1088_,
		_w1089_
	);
	LUT3 #(
		.INIT('h23)
	) name637 (
		_w921_,
		_w923_,
		_w945_,
		_w1090_
	);
	LUT4 #(
		.INIT('h5110)
	) name638 (
		_w919_,
		_w853_,
		_w920_,
		_w945_,
		_w1091_
	);
	LUT2 #(
		.INIT('h2)
	) name639 (
		_w959_,
		_w1091_,
		_w1092_
	);
	LUT2 #(
		.INIT('h8)
	) name640 (
		_w963_,
		_w972_,
		_w1093_
	);
	LUT3 #(
		.INIT('h20)
	) name641 (
		_w963_,
		_w968_,
		_w972_,
		_w1094_
	);
	LUT2 #(
		.INIT('h8)
	) name642 (
		_w977_,
		_w1094_,
		_w1095_
	);
	LUT4 #(
		.INIT('h2000)
	) name643 (
		_w957_,
		_w1089_,
		_w1092_,
		_w1095_,
		_w1096_
	);
	LUT4 #(
		.INIT('h8111)
	) name644 (
		\InstAddrPointer_reg[25]/NET0131 ,
		\InstAddrPointer_reg[26]/NET0131 ,
		_w981_,
		_w897_,
		_w1097_
	);
	LUT3 #(
		.INIT('h10)
	) name645 (
		_w994_,
		_w996_,
		_w1097_,
		_w1098_
	);
	LUT4 #(
		.INIT('h4000)
	) name646 (
		_w966_,
		_w988_,
		_w1096_,
		_w1098_,
		_w1099_
	);
	LUT3 #(
		.INIT('h41)
	) name647 (
		_w836_,
		_w997_,
		_w1099_,
		_w1100_
	);
	LUT3 #(
		.INIT('h80)
	) name648 (
		_w894_,
		_w896_,
		_w908_,
		_w1101_
	);
	LUT4 #(
		.INIT('h1551)
	) name649 (
		_w674_,
		_w836_,
		_w909_,
		_w1101_,
		_w1102_
	);
	LUT4 #(
		.INIT('h8a88)
	) name650 (
		_w608_,
		_w1084_,
		_w1100_,
		_w1102_,
		_w1103_
	);
	LUT3 #(
		.INIT('h6a)
	) name651 (
		\InstAddrPointer_reg[29]/NET0131 ,
		_w740_,
		_w1010_,
		_w1104_
	);
	LUT3 #(
		.INIT('h0b)
	) name652 (
		_w1023_,
		_w1027_,
		_w1033_,
		_w1105_
	);
	LUT4 #(
		.INIT('hfd00)
	) name653 (
		_w1026_,
		_w1028_,
		_w1031_,
		_w1105_,
		_w1106_
	);
	LUT3 #(
		.INIT('h0b)
	) name654 (
		_w1018_,
		_w1034_,
		_w1036_,
		_w1107_
	);
	LUT3 #(
		.INIT('hd0)
	) name655 (
		_w1021_,
		_w1106_,
		_w1107_,
		_w1108_
	);
	LUT4 #(
		.INIT('h3100)
	) name656 (
		_w1021_,
		_w1037_,
		_w1106_,
		_w1107_,
		_w1109_
	);
	LUT3 #(
		.INIT('h08)
	) name657 (
		_w1016_,
		_w1050_,
		_w1109_,
		_w1110_
	);
	LUT4 #(
		.INIT('h4888)
	) name658 (
		\InstAddrPointer_reg[17]/NET0131 ,
		\InstAddrPointer_reg[18]/NET0131 ,
		_w731_,
		_w1007_,
		_w1111_
	);
	LUT2 #(
		.INIT('h8)
	) name659 (
		_w1062_,
		_w1111_,
		_w1112_
	);
	LUT4 #(
		.INIT('h0800)
	) name660 (
		_w1016_,
		_w1050_,
		_w1109_,
		_w1112_,
		_w1113_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name661 (
		\InstAddrPointer_reg[24]/NET0131 ,
		\InstAddrPointer_reg[25]/NET0131 ,
		_w735_,
		_w1009_,
		_w1114_
	);
	LUT4 #(
		.INIT('h8000)
	) name662 (
		\InstAddrPointer_reg[26]/NET0131 ,
		\InstAddrPointer_reg[28]/NET0131 ,
		_w1066_,
		_w1114_,
		_w1115_
	);
	LUT3 #(
		.INIT('h80)
	) name663 (
		_w1060_,
		_w1113_,
		_w1115_,
		_w1116_
	);
	LUT3 #(
		.INIT('h54)
	) name664 (
		\InstAddrPointer_reg[29]/NET0131 ,
		_w563_,
		_w633_,
		_w1117_
	);
	LUT4 #(
		.INIT('h00c8)
	) name665 (
		_w569_,
		_w602_,
		_w604_,
		_w1117_,
		_w1118_
	);
	LUT2 #(
		.INIT('h8)
	) name666 (
		_w1104_,
		_w1118_,
		_w1119_
	);
	LUT4 #(
		.INIT('hfe00)
	) name667 (
		_w586_,
		_w582_,
		_w589_,
		_w566_,
		_w1120_
	);
	LUT4 #(
		.INIT('h0057)
	) name668 (
		READY_n_pad,
		_w588_,
		_w596_,
		_w1120_,
		_w1121_
	);
	LUT3 #(
		.INIT('h2a)
	) name669 (
		\InstAddrPointer_reg[29]/NET0131 ,
		_w1074_,
		_w1121_,
		_w1122_
	);
	LUT3 #(
		.INIT('hb0)
	) name670 (
		_w616_,
		_w630_,
		_w997_,
		_w1123_
	);
	LUT3 #(
		.INIT('h0e)
	) name671 (
		_w588_,
		_w596_,
		_w741_,
		_w1124_
	);
	LUT3 #(
		.INIT('hc4)
	) name672 (
		_w597_,
		_w909_,
		_w1124_,
		_w1125_
	);
	LUT4 #(
		.INIT('h0001)
	) name673 (
		_w1123_,
		_w1125_,
		_w1122_,
		_w1119_,
		_w1126_
	);
	LUT4 #(
		.INIT('hd700)
	) name674 (
		_w671_,
		_w1104_,
		_w1116_,
		_w1126_,
		_w1127_
	);
	LUT4 #(
		.INIT('h153f)
	) name675 (
		\InstAddrPointer_reg[29]/NET0131 ,
		\rEIP_reg[29]/NET0131 ,
		_w1080_,
		_w1081_,
		_w1128_
	);
	LUT4 #(
		.INIT('h8aff)
	) name676 (
		_w690_,
		_w1103_,
		_w1127_,
		_w1128_,
		_w1129_
	);
	LUT3 #(
		.INIT('h08)
	) name677 (
		\InstAddrPointer_reg[27]/NET0131 ,
		_w563_,
		_w673_,
		_w1130_
	);
	LUT2 #(
		.INIT('h6)
	) name678 (
		\InstAddrPointer_reg[11]/NET0131 ,
		_w726_,
		_w1131_
	);
	LUT4 #(
		.INIT('h4800)
	) name679 (
		\InstAddrPointer_reg[11]/NET0131 ,
		\InstAddrPointer_reg[12]/NET0131 ,
		_w726_,
		_w887_,
		_w1132_
	);
	LUT3 #(
		.INIT('h32)
	) name680 (
		\InstAddrPointer_reg[10]/NET0131 ,
		_w726_,
		_w889_,
		_w1133_
	);
	LUT2 #(
		.INIT('h8)
	) name681 (
		\InstAddrPointer_reg[9]/NET0131 ,
		_w839_,
		_w1134_
	);
	LUT4 #(
		.INIT('h2080)
	) name682 (
		\InstAddrPointer_reg[10]/NET0131 ,
		\InstAddrPointer_reg[8]/NET0131 ,
		\InstAddrPointer_reg[9]/NET0131 ,
		_w723_,
		_w1135_
	);
	LUT4 #(
		.INIT('hf700)
	) name683 (
		_w830_,
		_w835_,
		_w837_,
		_w1135_,
		_w1136_
	);
	LUT4 #(
		.INIT('h8f00)
	) name684 (
		_w825_,
		_w869_,
		_w875_,
		_w1136_,
		_w1137_
	);
	LUT3 #(
		.INIT('h0e)
	) name685 (
		\InstAddrPointer_reg[26]/NET0131 ,
		_w738_,
		_w900_,
		_w1138_
	);
	LUT3 #(
		.INIT('h80)
	) name686 (
		_w736_,
		_w884_,
		_w903_,
		_w1139_
	);
	LUT2 #(
		.INIT('h8)
	) name687 (
		_w1138_,
		_w1139_,
		_w1140_
	);
	LUT4 #(
		.INIT('h8000)
	) name688 (
		_w883_,
		_w1132_,
		_w1137_,
		_w1140_,
		_w1141_
	);
	LUT3 #(
		.INIT('h82)
	) name689 (
		_w836_,
		_w901_,
		_w1141_,
		_w1142_
	);
	LUT4 #(
		.INIT('h9300)
	) name690 (
		\InstAddrPointer_reg[21]/NET0131 ,
		\InstAddrPointer_reg[22]/NET0131 ,
		_w965_,
		_w969_,
		_w1143_
	);
	LUT2 #(
		.INIT('h1)
	) name691 (
		_w921_,
		_w940_,
		_w1144_
	);
	LUT3 #(
		.INIT('h40)
	) name692 (
		_w1085_,
		_w1086_,
		_w1144_,
		_w1145_
	);
	LUT3 #(
		.INIT('h8a)
	) name693 (
		_w1090_,
		_w1087_,
		_w1144_,
		_w1146_
	);
	LUT4 #(
		.INIT('h8c88)
	) name694 (
		_w919_,
		_w964_,
		_w1145_,
		_w1146_,
		_w1147_
	);
	LUT2 #(
		.INIT('h8)
	) name695 (
		_w986_,
		_w1097_,
		_w1148_
	);
	LUT4 #(
		.INIT('h8000)
	) name696 (
		_w978_,
		_w1143_,
		_w1147_,
		_w1148_,
		_w1149_
	);
	LUT4 #(
		.INIT('h4554)
	) name697 (
		_w674_,
		_w836_,
		_w994_,
		_w1149_,
		_w1150_
	);
	LUT4 #(
		.INIT('h8a88)
	) name698 (
		_w608_,
		_w1130_,
		_w1142_,
		_w1150_,
		_w1151_
	);
	LUT4 #(
		.INIT('h1555)
	) name699 (
		\InstAddrPointer_reg[11]/NET0131 ,
		\InstAddrPointer_reg[7]/NET0131 ,
		_w725_,
		_w1005_,
		_w1152_
	);
	LUT3 #(
		.INIT('h07)
	) name700 (
		_w885_,
		_w1041_,
		_w1152_,
		_w1153_
	);
	LUT3 #(
		.INIT('h80)
	) name701 (
		_w1043_,
		_w1046_,
		_w1153_,
		_w1154_
	);
	LUT3 #(
		.INIT('h6c)
	) name702 (
		\InstAddrPointer_reg[14]/NET0131 ,
		\InstAddrPointer_reg[15]/NET0131 ,
		_w1007_,
		_w1155_
	);
	LUT3 #(
		.INIT('h6a)
	) name703 (
		\InstAddrPointer_reg[16]/NET0131 ,
		_w730_,
		_w1007_,
		_w1156_
	);
	LUT4 #(
		.INIT('h4888)
	) name704 (
		\InstAddrPointer_reg[16]/NET0131 ,
		_w718_,
		_w730_,
		_w1007_,
		_w1157_
	);
	LUT2 #(
		.INIT('h8)
	) name705 (
		_w1155_,
		_w1157_,
		_w1158_
	);
	LUT4 #(
		.INIT('h2000)
	) name706 (
		_w1016_,
		_w1109_,
		_w1154_,
		_w1158_,
		_w1159_
	);
	LUT2 #(
		.INIT('h8)
	) name707 (
		_w1057_,
		_w1062_,
		_w1160_
	);
	LUT3 #(
		.INIT('h6a)
	) name708 (
		\InstAddrPointer_reg[23]/NET0131 ,
		_w734_,
		_w1009_,
		_w1161_
	);
	LUT4 #(
		.INIT('h4888)
	) name709 (
		\InstAddrPointer_reg[23]/NET0131 ,
		\InstAddrPointer_reg[24]/NET0131 ,
		_w734_,
		_w1009_,
		_w1162_
	);
	LUT3 #(
		.INIT('h80)
	) name710 (
		\InstAddrPointer_reg[26]/NET0131 ,
		_w1114_,
		_w1162_,
		_w1163_
	);
	LUT3 #(
		.INIT('h80)
	) name711 (
		_w1159_,
		_w1160_,
		_w1163_,
		_w1164_
	);
	LUT4 #(
		.INIT('h0001)
	) name712 (
		_w642_,
		_w611_,
		_w613_,
		_w680_,
		_w1165_
	);
	LUT2 #(
		.INIT('h4)
	) name713 (
		_w597_,
		_w901_,
		_w1166_
	);
	LUT2 #(
		.INIT('h8)
	) name714 (
		_w635_,
		_w1066_,
		_w1167_
	);
	LUT4 #(
		.INIT('h004f)
	) name715 (
		_w616_,
		_w630_,
		_w994_,
		_w1167_,
		_w1168_
	);
	LUT4 #(
		.INIT('h0d00)
	) name716 (
		\InstAddrPointer_reg[27]/NET0131 ,
		_w1165_,
		_w1166_,
		_w1168_,
		_w1169_
	);
	LUT4 #(
		.INIT('hd700)
	) name717 (
		_w671_,
		_w1066_,
		_w1164_,
		_w1169_,
		_w1170_
	);
	LUT4 #(
		.INIT('h153f)
	) name718 (
		\InstAddrPointer_reg[27]/NET0131 ,
		\rEIP_reg[27]/NET0131 ,
		_w1080_,
		_w1081_,
		_w1171_
	);
	LUT4 #(
		.INIT('h8aff)
	) name719 (
		_w690_,
		_w1151_,
		_w1170_,
		_w1171_,
		_w1172_
	);
	LUT3 #(
		.INIT('h08)
	) name720 (
		\PhyAddrPointer_reg[31]/NET0131 ,
		_w563_,
		_w673_,
		_w1173_
	);
	LUT2 #(
		.INIT('h2)
	) name721 (
		_w998_,
		_w1001_,
		_w1174_
	);
	LUT4 #(
		.INIT('h78f0)
	) name722 (
		\InstAddrPointer_reg[29]/NET0131 ,
		\InstAddrPointer_reg[30]/NET0131 ,
		\InstAddrPointer_reg[31]/NET0131 ,
		_w995_,
		_w1175_
	);
	LUT4 #(
		.INIT('h4015)
	) name723 (
		_w836_,
		_w1149_,
		_w1174_,
		_w1175_,
		_w1176_
	);
	LUT2 #(
		.INIT('h6)
	) name724 (
		\InstAddrPointer_reg[31]/NET0131 ,
		_w743_,
		_w1177_
	);
	LUT4 #(
		.INIT('h1551)
	) name725 (
		_w674_,
		_w836_,
		_w913_,
		_w1177_,
		_w1178_
	);
	LUT4 #(
		.INIT('h8a88)
	) name726 (
		_w608_,
		_w1173_,
		_w1176_,
		_w1178_,
		_w1179_
	);
	LUT4 #(
		.INIT('h202a)
	) name727 (
		\PhyAddrPointer_reg[31]/NET0131 ,
		_w634_,
		_w607_,
		_w608_,
		_w1180_
	);
	LUT3 #(
		.INIT('h80)
	) name728 (
		_w1067_,
		_w1069_,
		_w1163_,
		_w1181_
	);
	LUT3 #(
		.INIT('h80)
	) name729 (
		_w1159_,
		_w1160_,
		_w1181_,
		_w1182_
	);
	LUT2 #(
		.INIT('h6)
	) name730 (
		\InstAddrPointer_reg[31]/NET0131 ,
		_w1068_,
		_w1183_
	);
	LUT4 #(
		.INIT('h8000)
	) name731 (
		_w1159_,
		_w1160_,
		_w1181_,
		_w1183_,
		_w1184_
	);
	LUT4 #(
		.INIT('h007f)
	) name732 (
		_w1159_,
		_w1160_,
		_w1181_,
		_w1183_,
		_w1185_
	);
	LUT3 #(
		.INIT('h02)
	) name733 (
		_w671_,
		_w1185_,
		_w1184_,
		_w1186_
	);
	LUT4 #(
		.INIT('h3113)
	) name734 (
		_w671_,
		_w1180_,
		_w1182_,
		_w1183_,
		_w1187_
	);
	LUT2 #(
		.INIT('h8)
	) name735 (
		\PhyAddrPointer_reg[22]/NET0131 ,
		\PhyAddrPointer_reg[23]/NET0131 ,
		_w1188_
	);
	LUT3 #(
		.INIT('h80)
	) name736 (
		\PhyAddrPointer_reg[22]/NET0131 ,
		\PhyAddrPointer_reg[23]/NET0131 ,
		\PhyAddrPointer_reg[24]/NET0131 ,
		_w1189_
	);
	LUT3 #(
		.INIT('h80)
	) name737 (
		\PhyAddrPointer_reg[2]/NET0131 ,
		\PhyAddrPointer_reg[3]/NET0131 ,
		\PhyAddrPointer_reg[4]/NET0131 ,
		_w1190_
	);
	LUT4 #(
		.INIT('h8000)
	) name738 (
		\PhyAddrPointer_reg[2]/NET0131 ,
		\PhyAddrPointer_reg[3]/NET0131 ,
		\PhyAddrPointer_reg[4]/NET0131 ,
		\PhyAddrPointer_reg[5]/NET0131 ,
		_w1191_
	);
	LUT2 #(
		.INIT('h8)
	) name739 (
		\PhyAddrPointer_reg[6]/NET0131 ,
		_w1191_,
		_w1192_
	);
	LUT3 #(
		.INIT('h80)
	) name740 (
		\PhyAddrPointer_reg[6]/NET0131 ,
		\PhyAddrPointer_reg[7]/NET0131 ,
		_w1191_,
		_w1193_
	);
	LUT4 #(
		.INIT('h8000)
	) name741 (
		\PhyAddrPointer_reg[6]/NET0131 ,
		\PhyAddrPointer_reg[7]/NET0131 ,
		\PhyAddrPointer_reg[8]/NET0131 ,
		_w1191_,
		_w1194_
	);
	LUT3 #(
		.INIT('h80)
	) name742 (
		\PhyAddrPointer_reg[10]/NET0131 ,
		\PhyAddrPointer_reg[9]/NET0131 ,
		_w1194_,
		_w1195_
	);
	LUT2 #(
		.INIT('h8)
	) name743 (
		\PhyAddrPointer_reg[11]/NET0131 ,
		\PhyAddrPointer_reg[12]/NET0131 ,
		_w1196_
	);
	LUT3 #(
		.INIT('h80)
	) name744 (
		\PhyAddrPointer_reg[11]/NET0131 ,
		\PhyAddrPointer_reg[12]/NET0131 ,
		\PhyAddrPointer_reg[13]/NET0131 ,
		_w1197_
	);
	LUT4 #(
		.INIT('h8000)
	) name745 (
		\PhyAddrPointer_reg[10]/NET0131 ,
		\PhyAddrPointer_reg[9]/NET0131 ,
		_w1194_,
		_w1197_,
		_w1198_
	);
	LUT2 #(
		.INIT('h8)
	) name746 (
		\PhyAddrPointer_reg[15]/NET0131 ,
		\PhyAddrPointer_reg[16]/NET0131 ,
		_w1199_
	);
	LUT3 #(
		.INIT('h80)
	) name747 (
		\PhyAddrPointer_reg[15]/NET0131 ,
		\PhyAddrPointer_reg[16]/NET0131 ,
		\PhyAddrPointer_reg[17]/NET0131 ,
		_w1200_
	);
	LUT3 #(
		.INIT('h80)
	) name748 (
		\PhyAddrPointer_reg[14]/NET0131 ,
		_w1198_,
		_w1200_,
		_w1201_
	);
	LUT2 #(
		.INIT('h8)
	) name749 (
		\PhyAddrPointer_reg[18]/NET0131 ,
		\PhyAddrPointer_reg[19]/NET0131 ,
		_w1202_
	);
	LUT4 #(
		.INIT('h8000)
	) name750 (
		\PhyAddrPointer_reg[18]/NET0131 ,
		\PhyAddrPointer_reg[19]/NET0131 ,
		\PhyAddrPointer_reg[20]/NET0131 ,
		\PhyAddrPointer_reg[21]/NET0131 ,
		_w1203_
	);
	LUT4 #(
		.INIT('h8000)
	) name751 (
		\PhyAddrPointer_reg[14]/NET0131 ,
		_w1198_,
		_w1200_,
		_w1203_,
		_w1204_
	);
	LUT3 #(
		.INIT('h80)
	) name752 (
		\PhyAddrPointer_reg[25]/NET0131 ,
		_w1189_,
		_w1204_,
		_w1205_
	);
	LUT4 #(
		.INIT('h8000)
	) name753 (
		\PhyAddrPointer_reg[25]/NET0131 ,
		\PhyAddrPointer_reg[26]/NET0131 ,
		_w1189_,
		_w1204_,
		_w1206_
	);
	LUT3 #(
		.INIT('h80)
	) name754 (
		\PhyAddrPointer_reg[27]/NET0131 ,
		\PhyAddrPointer_reg[28]/NET0131 ,
		_w1206_,
		_w1207_
	);
	LUT4 #(
		.INIT('h8000)
	) name755 (
		\PhyAddrPointer_reg[27]/NET0131 ,
		\PhyAddrPointer_reg[28]/NET0131 ,
		\PhyAddrPointer_reg[29]/NET0131 ,
		_w1206_,
		_w1208_
	);
	LUT2 #(
		.INIT('h1)
	) name756 (
		\DataWidth_reg[1]/NET0131 ,
		\PhyAddrPointer_reg[1]/NET0131 ,
		_w1209_
	);
	LUT3 #(
		.INIT('h08)
	) name757 (
		\PhyAddrPointer_reg[30]/NET0131 ,
		_w1208_,
		_w1209_,
		_w1210_
	);
	LUT3 #(
		.INIT('h48)
	) name758 (
		\PhyAddrPointer_reg[31]/NET0131 ,
		_w695_,
		_w1210_,
		_w1211_
	);
	LUT4 #(
		.INIT('h0010)
	) name759 (
		\State2_reg[0]/NET0131 ,
		\State2_reg[1]/NET0131 ,
		\State2_reg[2]/NET0131 ,
		\State2_reg[3]/NET0131 ,
		_w1212_
	);
	LUT4 #(
		.INIT('h8000)
	) name760 (
		\PhyAddrPointer_reg[1]/NET0131 ,
		\PhyAddrPointer_reg[27]/NET0131 ,
		\PhyAddrPointer_reg[28]/NET0131 ,
		_w1206_,
		_w1213_
	);
	LUT4 #(
		.INIT('h870f)
	) name761 (
		\PhyAddrPointer_reg[29]/NET0131 ,
		\PhyAddrPointer_reg[30]/NET0131 ,
		\PhyAddrPointer_reg[31]/NET0131 ,
		_w1213_,
		_w1214_
	);
	LUT4 #(
		.INIT('hfc35)
	) name762 (
		\State2_reg[0]/NET0131 ,
		\State2_reg[1]/NET0131 ,
		\State2_reg[2]/NET0131 ,
		\State2_reg[3]/NET0131 ,
		_w1215_
	);
	LUT4 #(
		.INIT('h3f15)
	) name763 (
		\PhyAddrPointer_reg[31]/NET0131 ,
		\rEIP_reg[31]/NET0131 ,
		_w1080_,
		_w1215_,
		_w1216_
	);
	LUT3 #(
		.INIT('hd0)
	) name764 (
		_w1212_,
		_w1214_,
		_w1216_,
		_w1217_
	);
	LUT2 #(
		.INIT('h4)
	) name765 (
		_w1211_,
		_w1217_,
		_w1218_
	);
	LUT4 #(
		.INIT('h8aff)
	) name766 (
		_w690_,
		_w1179_,
		_w1187_,
		_w1218_,
		_w1219_
	);
	LUT3 #(
		.INIT('h08)
	) name767 (
		\InstAddrPointer_reg[15]/NET0131 ,
		_w563_,
		_w673_,
		_w1220_
	);
	LUT4 #(
		.INIT('h8222)
	) name768 (
		_w836_,
		_w881_,
		_w1132_,
		_w1137_,
		_w1221_
	);
	LUT4 #(
		.INIT('h4554)
	) name769 (
		_w674_,
		_w836_,
		_w970_,
		_w1147_,
		_w1222_
	);
	LUT4 #(
		.INIT('h8a88)
	) name770 (
		_w608_,
		_w1220_,
		_w1221_,
		_w1222_,
		_w1223_
	);
	LUT4 #(
		.INIT('h00df)
	) name771 (
		_w1016_,
		_w1109_,
		_w1154_,
		_w1155_,
		_w1224_
	);
	LUT4 #(
		.INIT('haa2a)
	) name772 (
		_w671_,
		_w1016_,
		_w1048_,
		_w1109_,
		_w1225_
	);
	LUT2 #(
		.INIT('h4)
	) name773 (
		_w1224_,
		_w1225_,
		_w1226_
	);
	LUT2 #(
		.INIT('h4)
	) name774 (
		_w597_,
		_w881_,
		_w1227_
	);
	LUT2 #(
		.INIT('h8)
	) name775 (
		_w635_,
		_w1155_,
		_w1228_
	);
	LUT4 #(
		.INIT('h004f)
	) name776 (
		_w616_,
		_w630_,
		_w970_,
		_w1228_,
		_w1229_
	);
	LUT4 #(
		.INIT('h0d00)
	) name777 (
		\InstAddrPointer_reg[15]/NET0131 ,
		_w1165_,
		_w1227_,
		_w1229_,
		_w1230_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name778 (
		_w690_,
		_w1223_,
		_w1226_,
		_w1230_,
		_w1231_
	);
	LUT4 #(
		.INIT('h153f)
	) name779 (
		\InstAddrPointer_reg[15]/NET0131 ,
		\rEIP_reg[15]/NET0131 ,
		_w1080_,
		_w1081_,
		_w1232_
	);
	LUT2 #(
		.INIT('hb)
	) name780 (
		_w1231_,
		_w1232_,
		_w1233_
	);
	LUT3 #(
		.INIT('h08)
	) name781 (
		\InstAddrPointer_reg[22]/NET0131 ,
		_w563_,
		_w673_,
		_w1234_
	);
	LUT4 #(
		.INIT('h78f0)
	) name782 (
		\InstAddrPointer_reg[20]/NET0131 ,
		\InstAddrPointer_reg[21]/NET0131 ,
		\InstAddrPointer_reg[22]/NET0131 ,
		_w733_,
		_w1235_
	);
	LUT4 #(
		.INIT('h366c)
	) name783 (
		\InstAddrPointer_reg[21]/NET0131 ,
		\InstAddrPointer_reg[22]/NET0131 ,
		_w877_,
		_w894_,
		_w1236_
	);
	LUT2 #(
		.INIT('h2)
	) name784 (
		_w836_,
		_w1236_,
		_w1237_
	);
	LUT4 #(
		.INIT('h4554)
	) name785 (
		_w674_,
		_w836_,
		_w980_,
		_w987_,
		_w1238_
	);
	LUT4 #(
		.INIT('h8a88)
	) name786 (
		_w608_,
		_w1234_,
		_w1237_,
		_w1238_,
		_w1239_
	);
	LUT3 #(
		.INIT('h6c)
	) name787 (
		\InstAddrPointer_reg[21]/NET0131 ,
		\InstAddrPointer_reg[22]/NET0131 ,
		_w1009_,
		_w1240_
	);
	LUT4 #(
		.INIT('h007f)
	) name788 (
		_w1055_,
		_w1056_,
		_w1062_,
		_w1240_,
		_w1241_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name789 (
		_w671_,
		_w1055_,
		_w1057_,
		_w1062_,
		_w1242_
	);
	LUT3 #(
		.INIT('hb8)
	) name790 (
		\InstAddrPointer_reg[22]/NET0131 ,
		READY_n_pad,
		_w1235_,
		_w1243_
	);
	LUT3 #(
		.INIT('h80)
	) name791 (
		_w494_,
		_w586_,
		_w1243_,
		_w1244_
	);
	LUT4 #(
		.INIT('haa8a)
	) name792 (
		\InstAddrPointer_reg[22]/NET0131 ,
		_w613_,
		_w681_,
		_w1244_,
		_w1245_
	);
	LUT2 #(
		.INIT('h8)
	) name793 (
		_w554_,
		_w1235_,
		_w1246_
	);
	LUT4 #(
		.INIT('h010f)
	) name794 (
		_w588_,
		_w596_,
		_w1246_,
		_w1243_,
		_w1247_
	);
	LUT2 #(
		.INIT('h8)
	) name795 (
		_w635_,
		_w1240_,
		_w1248_
	);
	LUT4 #(
		.INIT('h004f)
	) name796 (
		_w616_,
		_w630_,
		_w987_,
		_w1248_,
		_w1249_
	);
	LUT3 #(
		.INIT('h40)
	) name797 (
		_w1245_,
		_w1247_,
		_w1249_,
		_w1250_
	);
	LUT3 #(
		.INIT('hb0)
	) name798 (
		_w1241_,
		_w1242_,
		_w1250_,
		_w1251_
	);
	LUT4 #(
		.INIT('h153f)
	) name799 (
		\InstAddrPointer_reg[22]/NET0131 ,
		\rEIP_reg[22]/NET0131 ,
		_w1080_,
		_w1081_,
		_w1252_
	);
	LUT4 #(
		.INIT('h8aff)
	) name800 (
		_w690_,
		_w1239_,
		_w1251_,
		_w1252_,
		_w1253_
	);
	LUT3 #(
		.INIT('h20)
	) name801 (
		_w1016_,
		_w1039_,
		_w1048_,
		_w1254_
	);
	LUT4 #(
		.INIT('h2000)
	) name802 (
		_w1016_,
		_w1039_,
		_w1048_,
		_w1156_,
		_w1255_
	);
	LUT3 #(
		.INIT('h80)
	) name803 (
		_w1058_,
		_w1112_,
		_w1255_,
		_w1256_
	);
	LUT4 #(
		.INIT('h8000)
	) name804 (
		_w1058_,
		_w1059_,
		_w1112_,
		_w1255_,
		_w1257_
	);
	LUT4 #(
		.INIT('h1333)
	) name805 (
		_w1058_,
		_w1059_,
		_w1112_,
		_w1255_,
		_w1258_
	);
	LUT3 #(
		.INIT('h02)
	) name806 (
		_w671_,
		_w1258_,
		_w1257_,
		_w1259_
	);
	LUT3 #(
		.INIT('h08)
	) name807 (
		\InstAddrPointer_reg[24]/NET0131 ,
		_w563_,
		_w673_,
		_w1260_
	);
	LUT4 #(
		.INIT('h0400)
	) name808 (
		_w971_,
		_w977_,
		_w983_,
		_w1143_,
		_w1261_
	);
	LUT4 #(
		.INIT('h0400)
	) name809 (
		_w948_,
		_w964_,
		_w970_,
		_w1261_,
		_w1262_
	);
	LUT3 #(
		.INIT('h41)
	) name810 (
		_w836_,
		_w985_,
		_w1262_,
		_w1263_
	);
	LUT3 #(
		.INIT('h0b)
	) name811 (
		_w793_,
		_w795_,
		_w823_,
		_w1264_
	);
	LUT2 #(
		.INIT('h1)
	) name812 (
		_w763_,
		_w868_,
		_w1265_
	);
	LUT4 #(
		.INIT('h2f00)
	) name813 (
		_w794_,
		_w820_,
		_w1264_,
		_w1265_,
		_w1266_
	);
	LUT3 #(
		.INIT('h0d)
	) name814 (
		_w822_,
		_w868_,
		_w873_,
		_w1267_
	);
	LUT2 #(
		.INIT('h1)
	) name815 (
		_w838_,
		_w855_,
		_w1268_
	);
	LUT3 #(
		.INIT('h23)
	) name816 (
		_w838_,
		_w871_,
		_w872_,
		_w1269_
	);
	LUT4 #(
		.INIT('h4f00)
	) name817 (
		_w1266_,
		_w1267_,
		_w1268_,
		_w1269_,
		_w1270_
	);
	LUT2 #(
		.INIT('h8)
	) name818 (
		_w839_,
		_w892_,
		_w1271_
	);
	LUT2 #(
		.INIT('h4)
	) name819 (
		_w1270_,
		_w1271_,
		_w1272_
	);
	LUT3 #(
		.INIT('h60)
	) name820 (
		\InstAddrPointer_reg[20]/NET0131 ,
		_w733_,
		_w735_,
		_w1273_
	);
	LUT3 #(
		.INIT('h40)
	) name821 (
		_w1270_,
		_w1271_,
		_w1273_,
		_w1274_
	);
	LUT4 #(
		.INIT('h1551)
	) name822 (
		_w674_,
		_w836_,
		_w902_,
		_w1274_,
		_w1275_
	);
	LUT4 #(
		.INIT('h8a88)
	) name823 (
		_w608_,
		_w1260_,
		_w1263_,
		_w1275_,
		_w1276_
	);
	LUT2 #(
		.INIT('h4)
	) name824 (
		_w597_,
		_w902_,
		_w1277_
	);
	LUT2 #(
		.INIT('h8)
	) name825 (
		_w635_,
		_w1059_,
		_w1278_
	);
	LUT4 #(
		.INIT('h004f)
	) name826 (
		_w616_,
		_w630_,
		_w985_,
		_w1278_,
		_w1279_
	);
	LUT4 #(
		.INIT('h0d00)
	) name827 (
		\InstAddrPointer_reg[24]/NET0131 ,
		_w1165_,
		_w1277_,
		_w1279_,
		_w1280_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name828 (
		_w690_,
		_w1276_,
		_w1259_,
		_w1280_,
		_w1281_
	);
	LUT4 #(
		.INIT('h153f)
	) name829 (
		\InstAddrPointer_reg[24]/NET0131 ,
		\rEIP_reg[24]/NET0131 ,
		_w1080_,
		_w1081_,
		_w1282_
	);
	LUT2 #(
		.INIT('hb)
	) name830 (
		_w1281_,
		_w1282_,
		_w1283_
	);
	LUT3 #(
		.INIT('h08)
	) name831 (
		\InstAddrPointer_reg[26]/NET0131 ,
		_w563_,
		_w673_,
		_w1284_
	);
	LUT3 #(
		.INIT('h08)
	) name832 (
		_w1132_,
		_w1135_,
		_w1270_,
		_w1285_
	);
	LUT4 #(
		.INIT('h0080)
	) name833 (
		_w883_,
		_w1132_,
		_w1135_,
		_w1270_,
		_w1286_
	);
	LUT4 #(
		.INIT('h8222)
	) name834 (
		_w836_,
		_w1138_,
		_w1139_,
		_w1286_,
		_w1287_
	);
	LUT4 #(
		.INIT('h4554)
	) name835 (
		_w674_,
		_w836_,
		_w991_,
		_w999_,
		_w1288_
	);
	LUT4 #(
		.INIT('h8a88)
	) name836 (
		_w608_,
		_w1284_,
		_w1287_,
		_w1288_,
		_w1289_
	);
	LUT4 #(
		.INIT('h2888)
	) name837 (
		_w671_,
		_w1012_,
		_w1055_,
		_w1063_,
		_w1290_
	);
	LUT2 #(
		.INIT('h8)
	) name838 (
		_w635_,
		_w1012_,
		_w1291_
	);
	LUT3 #(
		.INIT('hd0)
	) name839 (
		_w647_,
		_w648_,
		_w1138_,
		_w1292_
	);
	LUT3 #(
		.INIT('hb0)
	) name840 (
		_w616_,
		_w630_,
		_w999_,
		_w1293_
	);
	LUT4 #(
		.INIT('hec00)
	) name841 (
		_w585_,
		_w589_,
		_w590_,
		_w1138_,
		_w1294_
	);
	LUT4 #(
		.INIT('h0001)
	) name842 (
		_w642_,
		_w653_,
		_w655_,
		_w680_,
		_w1295_
	);
	LUT3 #(
		.INIT('h8a)
	) name843 (
		\InstAddrPointer_reg[26]/NET0131 ,
		_w1294_,
		_w1295_,
		_w1296_
	);
	LUT4 #(
		.INIT('h0001)
	) name844 (
		_w1293_,
		_w1296_,
		_w1292_,
		_w1291_,
		_w1297_
	);
	LUT2 #(
		.INIT('h4)
	) name845 (
		_w1290_,
		_w1297_,
		_w1298_
	);
	LUT4 #(
		.INIT('h153f)
	) name846 (
		\InstAddrPointer_reg[26]/NET0131 ,
		\rEIP_reg[26]/NET0131 ,
		_w1080_,
		_w1081_,
		_w1299_
	);
	LUT4 #(
		.INIT('h8aff)
	) name847 (
		_w690_,
		_w1289_,
		_w1298_,
		_w1299_,
		_w1300_
	);
	LUT4 #(
		.INIT('h4744)
	) name848 (
		\PhyAddrPointer_reg[30]/NET0131 ,
		_w674_,
		_w915_,
		_w1002_,
		_w1301_
	);
	LUT4 #(
		.INIT('h202a)
	) name849 (
		\PhyAddrPointer_reg[30]/NET0131 ,
		_w634_,
		_w607_,
		_w608_,
		_w1302_
	);
	LUT4 #(
		.INIT('h0031)
	) name850 (
		_w608_,
		_w1070_,
		_w1301_,
		_w1302_,
		_w1303_
	);
	LUT3 #(
		.INIT('h6c)
	) name851 (
		\PhyAddrPointer_reg[29]/NET0131 ,
		\PhyAddrPointer_reg[30]/NET0131 ,
		_w1213_,
		_w1304_
	);
	LUT4 #(
		.INIT('hffeb)
	) name852 (
		\State2_reg[0]/NET0131 ,
		\State2_reg[1]/NET0131 ,
		\State2_reg[2]/NET0131 ,
		\State2_reg[3]/NET0131 ,
		_w1305_
	);
	LUT3 #(
		.INIT('h0d)
	) name853 (
		\DataWidth_reg[1]/NET0131 ,
		_w1212_,
		_w1305_,
		_w1306_
	);
	LUT4 #(
		.INIT('h6c00)
	) name854 (
		\PhyAddrPointer_reg[29]/NET0131 ,
		\PhyAddrPointer_reg[30]/NET0131 ,
		_w1213_,
		_w1306_,
		_w1307_
	);
	LUT4 #(
		.INIT('h3f15)
	) name855 (
		\PhyAddrPointer_reg[30]/NET0131 ,
		\rEIP_reg[30]/NET0131 ,
		_w1080_,
		_w1215_,
		_w1308_
	);
	LUT4 #(
		.INIT('hb700)
	) name856 (
		\PhyAddrPointer_reg[30]/NET0131 ,
		_w714_,
		_w1208_,
		_w1308_,
		_w1309_
	);
	LUT2 #(
		.INIT('h4)
	) name857 (
		_w1307_,
		_w1309_,
		_w1310_
	);
	LUT3 #(
		.INIT('h2f)
	) name858 (
		_w690_,
		_w1303_,
		_w1310_,
		_w1311_
	);
	LUT3 #(
		.INIT('h08)
	) name859 (
		\InstAddrPointer_reg[11]/NET0131 ,
		_w563_,
		_w673_,
		_w1312_
	);
	LUT3 #(
		.INIT('h82)
	) name860 (
		_w836_,
		_w1131_,
		_w1137_,
		_w1313_
	);
	LUT2 #(
		.INIT('h8)
	) name861 (
		_w959_,
		_w954_,
		_w1314_
	);
	LUT3 #(
		.INIT('h10)
	) name862 (
		_w948_,
		_w955_,
		_w1314_,
		_w1315_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name863 (
		_w955_,
		_w1145_,
		_w1146_,
		_w1314_,
		_w1316_
	);
	LUT2 #(
		.INIT('h1)
	) name864 (
		_w836_,
		_w1316_,
		_w1317_
	);
	LUT4 #(
		.INIT('h0045)
	) name865 (
		_w674_,
		_w1315_,
		_w1317_,
		_w1313_,
		_w1318_
	);
	LUT3 #(
		.INIT('ha8)
	) name866 (
		_w608_,
		_w1312_,
		_w1318_,
		_w1319_
	);
	LUT4 #(
		.INIT('h00f7)
	) name867 (
		_w1016_,
		_w1045_,
		_w1109_,
		_w1153_,
		_w1320_
	);
	LUT4 #(
		.INIT('h0080)
	) name868 (
		\InstAddrPointer_reg[11]/NET0131 ,
		_w1016_,
		_w1045_,
		_w1109_,
		_w1321_
	);
	LUT3 #(
		.INIT('h02)
	) name869 (
		_w671_,
		_w1321_,
		_w1320_,
		_w1322_
	);
	LUT3 #(
		.INIT('h0e)
	) name870 (
		_w588_,
		_w596_,
		_w726_,
		_w1323_
	);
	LUT3 #(
		.INIT('ha2)
	) name871 (
		\InstAddrPointer_reg[11]/NET0131 ,
		_w1165_,
		_w1323_,
		_w1324_
	);
	LUT2 #(
		.INIT('h4)
	) name872 (
		_w597_,
		_w1131_,
		_w1325_
	);
	LUT2 #(
		.INIT('h8)
	) name873 (
		_w635_,
		_w1153_,
		_w1326_
	);
	LUT4 #(
		.INIT('h004f)
	) name874 (
		_w616_,
		_w630_,
		_w955_,
		_w1326_,
		_w1327_
	);
	LUT2 #(
		.INIT('h4)
	) name875 (
		_w1325_,
		_w1327_,
		_w1328_
	);
	LUT3 #(
		.INIT('h10)
	) name876 (
		_w1324_,
		_w1322_,
		_w1328_,
		_w1329_
	);
	LUT4 #(
		.INIT('h153f)
	) name877 (
		\InstAddrPointer_reg[11]/NET0131 ,
		\rEIP_reg[11]/NET0131 ,
		_w1080_,
		_w1081_,
		_w1330_
	);
	LUT4 #(
		.INIT('h8aff)
	) name878 (
		_w690_,
		_w1319_,
		_w1329_,
		_w1330_,
		_w1331_
	);
	LUT3 #(
		.INIT('h08)
	) name879 (
		\InstAddrPointer_reg[14]/NET0131 ,
		_w563_,
		_w673_,
		_w1332_
	);
	LUT3 #(
		.INIT('h6a)
	) name880 (
		\InstAddrPointer_reg[14]/NET0131 ,
		_w726_,
		_w728_,
		_w1333_
	);
	LUT4 #(
		.INIT('h0080)
	) name881 (
		\InstAddrPointer_reg[12]/NET0131 ,
		_w1131_,
		_w1135_,
		_w1270_,
		_w1334_
	);
	LUT4 #(
		.INIT('h3230)
	) name882 (
		\InstAddrPointer_reg[13]/NET0131 ,
		_w1285_,
		_w1333_,
		_w1334_,
		_w1335_
	);
	LUT4 #(
		.INIT('h0100)
	) name883 (
		_w948_,
		_w951_,
		_w955_,
		_w1314_,
		_w1336_
	);
	LUT3 #(
		.INIT('h45)
	) name884 (
		_w836_,
		_w948_,
		_w964_,
		_w1337_
	);
	LUT4 #(
		.INIT('h7500)
	) name885 (
		_w961_,
		_w962_,
		_w1336_,
		_w1337_,
		_w1338_
	);
	LUT4 #(
		.INIT('h0051)
	) name886 (
		_w674_,
		_w836_,
		_w1335_,
		_w1338_,
		_w1339_
	);
	LUT2 #(
		.INIT('h6)
	) name887 (
		\InstAddrPointer_reg[14]/NET0131 ,
		_w1007_,
		_w1340_
	);
	LUT4 #(
		.INIT('h0800)
	) name888 (
		\InstAddrPointer_reg[10]/NET0131 ,
		_w1016_,
		_w1039_,
		_w1044_,
		_w1341_
	);
	LUT2 #(
		.INIT('h8)
	) name889 (
		_w1043_,
		_w1153_,
		_w1342_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name890 (
		_w671_,
		_w1016_,
		_w1039_,
		_w1154_,
		_w1343_
	);
	LUT4 #(
		.INIT('hea00)
	) name891 (
		_w1340_,
		_w1341_,
		_w1342_,
		_w1343_,
		_w1344_
	);
	LUT4 #(
		.INIT('haaa8)
	) name892 (
		\InstAddrPointer_reg[14]/NET0131 ,
		_w611_,
		_w613_,
		_w680_,
		_w1345_
	);
	LUT2 #(
		.INIT('h4)
	) name893 (
		_w597_,
		_w1333_,
		_w1346_
	);
	LUT4 #(
		.INIT('h0201)
	) name894 (
		\InstAddrPointer_reg[14]/NET0131 ,
		_w563_,
		_w633_,
		_w1007_,
		_w1347_
	);
	LUT3 #(
		.INIT('h54)
	) name895 (
		\InstAddrPointer_reg[14]/NET0131 ,
		_w563_,
		_w633_,
		_w1348_
	);
	LUT4 #(
		.INIT('h00c8)
	) name896 (
		_w569_,
		_w602_,
		_w604_,
		_w1348_,
		_w1349_
	);
	LUT2 #(
		.INIT('h4)
	) name897 (
		_w1347_,
		_w1349_,
		_w1350_
	);
	LUT4 #(
		.INIT('h004f)
	) name898 (
		_w616_,
		_w630_,
		_w961_,
		_w1350_,
		_w1351_
	);
	LUT3 #(
		.INIT('h10)
	) name899 (
		_w1346_,
		_w1345_,
		_w1351_,
		_w1352_
	);
	LUT2 #(
		.INIT('h4)
	) name900 (
		_w1344_,
		_w1352_,
		_w1353_
	);
	LUT4 #(
		.INIT('h5700)
	) name901 (
		_w608_,
		_w1332_,
		_w1339_,
		_w1353_,
		_w1354_
	);
	LUT4 #(
		.INIT('h153f)
	) name902 (
		\InstAddrPointer_reg[14]/NET0131 ,
		\rEIP_reg[14]/NET0131 ,
		_w1080_,
		_w1081_,
		_w1355_
	);
	LUT3 #(
		.INIT('h2f)
	) name903 (
		_w690_,
		_w1354_,
		_w1355_,
		_w1356_
	);
	LUT3 #(
		.INIT('h08)
	) name904 (
		\InstAddrPointer_reg[25]/NET0131 ,
		_w563_,
		_w673_,
		_w1357_
	);
	LUT4 #(
		.INIT('h0400)
	) name905 (
		_w966_,
		_w988_,
		_w989_,
		_w1096_,
		_w1358_
	);
	LUT4 #(
		.INIT('hb0f0)
	) name906 (
		_w966_,
		_w988_,
		_w989_,
		_w1096_,
		_w1359_
	);
	LUT3 #(
		.INIT('h01)
	) name907 (
		_w836_,
		_w1359_,
		_w1358_,
		_w1360_
	);
	LUT2 #(
		.INIT('h8)
	) name908 (
		\InstAddrPointer_reg[24]/NET0131 ,
		_w906_,
		_w1361_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name909 (
		\InstAddrPointer_reg[24]/NET0131 ,
		\InstAddrPointer_reg[25]/NET0131 ,
		_w733_,
		_w736_,
		_w1362_
	);
	LUT4 #(
		.INIT('h7f00)
	) name910 (
		_w894_,
		_w896_,
		_w1361_,
		_w1362_,
		_w1363_
	);
	LUT4 #(
		.INIT('h4000)
	) name911 (
		\InstAddrPointer_reg[25]/NET0131 ,
		_w894_,
		_w896_,
		_w1361_,
		_w1364_
	);
	LUT4 #(
		.INIT('h5551)
	) name912 (
		_w674_,
		_w836_,
		_w1364_,
		_w1363_,
		_w1365_
	);
	LUT4 #(
		.INIT('h8a88)
	) name913 (
		_w608_,
		_w1357_,
		_w1360_,
		_w1365_,
		_w1366_
	);
	LUT4 #(
		.INIT('h2a80)
	) name914 (
		_w671_,
		_w1060_,
		_w1113_,
		_w1114_,
		_w1367_
	);
	LUT3 #(
		.INIT('ha2)
	) name915 (
		READY_n_pad,
		_w591_,
		_w588_,
		_w1368_
	);
	LUT4 #(
		.INIT('h00ec)
	) name916 (
		_w585_,
		_w589_,
		_w590_,
		_w737_,
		_w1369_
	);
	LUT4 #(
		.INIT('h0004)
	) name917 (
		_w613_,
		_w681_,
		_w1368_,
		_w1369_,
		_w1370_
	);
	LUT2 #(
		.INIT('h4)
	) name918 (
		_w597_,
		_w1362_,
		_w1371_
	);
	LUT2 #(
		.INIT('h8)
	) name919 (
		_w635_,
		_w1114_,
		_w1372_
	);
	LUT4 #(
		.INIT('h004f)
	) name920 (
		_w616_,
		_w630_,
		_w989_,
		_w1372_,
		_w1373_
	);
	LUT4 #(
		.INIT('h0d00)
	) name921 (
		\InstAddrPointer_reg[25]/NET0131 ,
		_w1370_,
		_w1371_,
		_w1373_,
		_w1374_
	);
	LUT2 #(
		.INIT('h4)
	) name922 (
		_w1367_,
		_w1374_,
		_w1375_
	);
	LUT4 #(
		.INIT('h153f)
	) name923 (
		\InstAddrPointer_reg[25]/NET0131 ,
		\rEIP_reg[25]/NET0131 ,
		_w1080_,
		_w1081_,
		_w1376_
	);
	LUT4 #(
		.INIT('h8aff)
	) name924 (
		_w690_,
		_w1366_,
		_w1375_,
		_w1376_,
		_w1377_
	);
	LUT3 #(
		.INIT('h08)
	) name925 (
		\PhyAddrPointer_reg[15]/NET0131 ,
		_w563_,
		_w673_,
		_w1378_
	);
	LUT4 #(
		.INIT('haa20)
	) name926 (
		_w608_,
		_w1221_,
		_w1222_,
		_w1378_,
		_w1379_
	);
	LUT4 #(
		.INIT('h202a)
	) name927 (
		\PhyAddrPointer_reg[15]/NET0131 ,
		_w634_,
		_w607_,
		_w608_,
		_w1380_
	);
	LUT3 #(
		.INIT('h0b)
	) name928 (
		_w1224_,
		_w1225_,
		_w1380_,
		_w1381_
	);
	LUT4 #(
		.INIT('h3313)
	) name929 (
		\PhyAddrPointer_reg[14]/NET0131 ,
		\PhyAddrPointer_reg[15]/NET0131 ,
		_w1198_,
		_w1209_,
		_w1382_
	);
	LUT3 #(
		.INIT('h80)
	) name930 (
		\PhyAddrPointer_reg[14]/NET0131 ,
		\PhyAddrPointer_reg[15]/NET0131 ,
		_w1198_,
		_w1383_
	);
	LUT4 #(
		.INIT('h0080)
	) name931 (
		\PhyAddrPointer_reg[14]/NET0131 ,
		\PhyAddrPointer_reg[15]/NET0131 ,
		_w1198_,
		_w1209_,
		_w1384_
	);
	LUT3 #(
		.INIT('h02)
	) name932 (
		_w695_,
		_w1384_,
		_w1382_,
		_w1385_
	);
	LUT4 #(
		.INIT('h8000)
	) name933 (
		\PhyAddrPointer_reg[1]/NET0131 ,
		\PhyAddrPointer_reg[6]/NET0131 ,
		\PhyAddrPointer_reg[7]/NET0131 ,
		_w1191_,
		_w1386_
	);
	LUT4 #(
		.INIT('h8000)
	) name934 (
		\PhyAddrPointer_reg[10]/NET0131 ,
		\PhyAddrPointer_reg[8]/NET0131 ,
		\PhyAddrPointer_reg[9]/NET0131 ,
		_w1386_,
		_w1387_
	);
	LUT2 #(
		.INIT('h8)
	) name935 (
		_w1197_,
		_w1387_,
		_w1388_
	);
	LUT3 #(
		.INIT('h80)
	) name936 (
		\PhyAddrPointer_reg[14]/NET0131 ,
		_w1197_,
		_w1387_,
		_w1389_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name937 (
		\PhyAddrPointer_reg[14]/NET0131 ,
		\PhyAddrPointer_reg[15]/NET0131 ,
		_w1197_,
		_w1387_,
		_w1390_
	);
	LUT4 #(
		.INIT('h3f15)
	) name938 (
		\PhyAddrPointer_reg[15]/NET0131 ,
		\rEIP_reg[15]/NET0131 ,
		_w1080_,
		_w1215_,
		_w1391_
	);
	LUT3 #(
		.INIT('h70)
	) name939 (
		_w1212_,
		_w1390_,
		_w1391_,
		_w1392_
	);
	LUT2 #(
		.INIT('h4)
	) name940 (
		_w1385_,
		_w1392_,
		_w1393_
	);
	LUT4 #(
		.INIT('h8aff)
	) name941 (
		_w690_,
		_w1379_,
		_w1381_,
		_w1393_,
		_w1394_
	);
	LUT3 #(
		.INIT('h08)
	) name942 (
		\PhyAddrPointer_reg[23]/NET0131 ,
		_w563_,
		_w673_,
		_w1395_
	);
	LUT3 #(
		.INIT('h07)
	) name943 (
		_w894_,
		_w896_,
		_w906_,
		_w1396_
	);
	LUT3 #(
		.INIT('ha8)
	) name944 (
		_w836_,
		_w1274_,
		_w1396_,
		_w1397_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name945 (
		_w978_,
		_w983_,
		_w1143_,
		_w1147_,
		_w1398_
	);
	LUT3 #(
		.INIT('h54)
	) name946 (
		_w674_,
		_w836_,
		_w1398_,
		_w1399_
	);
	LUT4 #(
		.INIT('h8a88)
	) name947 (
		_w608_,
		_w1395_,
		_w1397_,
		_w1399_,
		_w1400_
	);
	LUT4 #(
		.INIT('h202a)
	) name948 (
		\PhyAddrPointer_reg[23]/NET0131 ,
		_w634_,
		_w607_,
		_w608_,
		_w1401_
	);
	LUT3 #(
		.INIT('h07)
	) name949 (
		_w1159_,
		_w1160_,
		_w1161_,
		_w1402_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name950 (
		_w671_,
		_w1058_,
		_w1112_,
		_w1255_,
		_w1403_
	);
	LUT3 #(
		.INIT('h45)
	) name951 (
		_w1401_,
		_w1402_,
		_w1403_,
		_w1404_
	);
	LUT4 #(
		.INIT('h8000)
	) name952 (
		\PhyAddrPointer_reg[14]/NET0131 ,
		\PhyAddrPointer_reg[1]/NET0131 ,
		_w1198_,
		_w1200_,
		_w1405_
	);
	LUT2 #(
		.INIT('h8)
	) name953 (
		_w1203_,
		_w1405_,
		_w1406_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name954 (
		\PhyAddrPointer_reg[22]/NET0131 ,
		\PhyAddrPointer_reg[23]/NET0131 ,
		_w1203_,
		_w1405_,
		_w1407_
	);
	LUT4 #(
		.INIT('h60c0)
	) name955 (
		\PhyAddrPointer_reg[22]/NET0131 ,
		\PhyAddrPointer_reg[23]/NET0131 ,
		_w714_,
		_w1204_,
		_w1408_
	);
	LUT4 #(
		.INIT('h3f15)
	) name956 (
		\PhyAddrPointer_reg[23]/NET0131 ,
		\rEIP_reg[23]/NET0131 ,
		_w1080_,
		_w1215_,
		_w1409_
	);
	LUT4 #(
		.INIT('h1300)
	) name957 (
		_w1306_,
		_w1408_,
		_w1407_,
		_w1409_,
		_w1410_
	);
	LUT4 #(
		.INIT('h8aff)
	) name958 (
		_w690_,
		_w1400_,
		_w1404_,
		_w1410_,
		_w1411_
	);
	LUT3 #(
		.INIT('h08)
	) name959 (
		\PhyAddrPointer_reg[27]/NET0131 ,
		_w563_,
		_w673_,
		_w1412_
	);
	LUT4 #(
		.INIT('haa20)
	) name960 (
		_w608_,
		_w1142_,
		_w1150_,
		_w1412_,
		_w1413_
	);
	LUT4 #(
		.INIT('h202a)
	) name961 (
		\PhyAddrPointer_reg[27]/NET0131 ,
		_w634_,
		_w607_,
		_w608_,
		_w1414_
	);
	LUT4 #(
		.INIT('h00d7)
	) name962 (
		_w671_,
		_w1066_,
		_w1164_,
		_w1414_,
		_w1415_
	);
	LUT3 #(
		.INIT('h6c)
	) name963 (
		\PhyAddrPointer_reg[1]/NET0131 ,
		\PhyAddrPointer_reg[27]/NET0131 ,
		_w1206_,
		_w1416_
	);
	LUT4 #(
		.INIT('h4105)
	) name964 (
		\DataWidth_reg[1]/NET0131 ,
		\PhyAddrPointer_reg[1]/NET0131 ,
		\PhyAddrPointer_reg[27]/NET0131 ,
		_w1206_,
		_w1417_
	);
	LUT4 #(
		.INIT('h70d0)
	) name965 (
		\DataWidth_reg[1]/NET0131 ,
		\PhyAddrPointer_reg[27]/NET0131 ,
		_w695_,
		_w1206_,
		_w1418_
	);
	LUT4 #(
		.INIT('h60c0)
	) name966 (
		\PhyAddrPointer_reg[1]/NET0131 ,
		\PhyAddrPointer_reg[27]/NET0131 ,
		_w1212_,
		_w1206_,
		_w1419_
	);
	LUT4 #(
		.INIT('h3f15)
	) name967 (
		\PhyAddrPointer_reg[27]/NET0131 ,
		\rEIP_reg[27]/NET0131 ,
		_w1080_,
		_w1215_,
		_w1420_
	);
	LUT4 #(
		.INIT('h4500)
	) name968 (
		_w1419_,
		_w1417_,
		_w1418_,
		_w1420_,
		_w1421_
	);
	LUT4 #(
		.INIT('h8aff)
	) name969 (
		_w690_,
		_w1413_,
		_w1415_,
		_w1421_,
		_w1422_
	);
	LUT3 #(
		.INIT('h08)
	) name970 (
		\PhyAddrPointer_reg[28]/NET0131 ,
		_w563_,
		_w673_,
		_w1423_
	);
	LUT3 #(
		.INIT('h10)
	) name971 (
		_w985_,
		_w994_,
		_w1097_,
		_w1424_
	);
	LUT4 #(
		.INIT('h4111)
	) name972 (
		_w836_,
		_w996_,
		_w1262_,
		_w1424_,
		_w1425_
	);
	LUT4 #(
		.INIT('h2000)
	) name973 (
		_w905_,
		_w1270_,
		_w1271_,
		_w1273_,
		_w1426_
	);
	LUT3 #(
		.INIT('h6a)
	) name974 (
		\InstAddrPointer_reg[28]/NET0131 ,
		_w739_,
		_w738_,
		_w1427_
	);
	LUT4 #(
		.INIT('h1551)
	) name975 (
		_w674_,
		_w836_,
		_w1426_,
		_w1427_,
		_w1428_
	);
	LUT4 #(
		.INIT('h8a88)
	) name976 (
		_w608_,
		_w1423_,
		_w1425_,
		_w1428_,
		_w1429_
	);
	LUT4 #(
		.INIT('h202a)
	) name977 (
		\PhyAddrPointer_reg[28]/NET0131 ,
		_w634_,
		_w607_,
		_w608_,
		_w1430_
	);
	LUT4 #(
		.INIT('h7f2a)
	) name978 (
		\InstAddrPointer_reg[28]/NET0131 ,
		_w739_,
		_w1010_,
		_w1065_,
		_w1431_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name979 (
		\InstAddrPointer_reg[20]/NET0131 ,
		_w719_,
		_w731_,
		_w1007_,
		_w1432_
	);
	LUT3 #(
		.INIT('h80)
	) name980 (
		\InstAddrPointer_reg[25]/NET0131 ,
		\InstAddrPointer_reg[26]/NET0131 ,
		\InstAddrPointer_reg[27]/NET0131 ,
		_w1433_
	);
	LUT2 #(
		.INIT('h8)
	) name981 (
		_w1432_,
		_w1433_,
		_w1434_
	);
	LUT3 #(
		.INIT('h80)
	) name982 (
		_w1058_,
		_w1059_,
		_w1434_,
		_w1435_
	);
	LUT3 #(
		.INIT('h80)
	) name983 (
		_w719_,
		_w1255_,
		_w1435_,
		_w1436_
	);
	LUT4 #(
		.INIT('h3113)
	) name984 (
		_w671_,
		_w1430_,
		_w1431_,
		_w1436_,
		_w1437_
	);
	LUT4 #(
		.INIT('h78f0)
	) name985 (
		\PhyAddrPointer_reg[1]/NET0131 ,
		\PhyAddrPointer_reg[27]/NET0131 ,
		\PhyAddrPointer_reg[28]/NET0131 ,
		_w1206_,
		_w1438_
	);
	LUT4 #(
		.INIT('h60c0)
	) name986 (
		\PhyAddrPointer_reg[27]/NET0131 ,
		\PhyAddrPointer_reg[28]/NET0131 ,
		_w714_,
		_w1206_,
		_w1439_
	);
	LUT4 #(
		.INIT('h3f15)
	) name987 (
		\PhyAddrPointer_reg[28]/NET0131 ,
		\rEIP_reg[28]/NET0131 ,
		_w1080_,
		_w1215_,
		_w1440_
	);
	LUT4 #(
		.INIT('h1300)
	) name988 (
		_w1306_,
		_w1439_,
		_w1438_,
		_w1440_,
		_w1441_
	);
	LUT4 #(
		.INIT('h8aff)
	) name989 (
		_w690_,
		_w1429_,
		_w1437_,
		_w1441_,
		_w1442_
	);
	LUT3 #(
		.INIT('h08)
	) name990 (
		\PhyAddrPointer_reg[29]/NET0131 ,
		_w563_,
		_w673_,
		_w1443_
	);
	LUT4 #(
		.INIT('haa20)
	) name991 (
		_w608_,
		_w1100_,
		_w1102_,
		_w1443_,
		_w1444_
	);
	LUT4 #(
		.INIT('h202a)
	) name992 (
		\PhyAddrPointer_reg[29]/NET0131 ,
		_w634_,
		_w607_,
		_w608_,
		_w1445_
	);
	LUT4 #(
		.INIT('h00d7)
	) name993 (
		_w671_,
		_w1104_,
		_w1116_,
		_w1445_,
		_w1446_
	);
	LUT2 #(
		.INIT('h6)
	) name994 (
		\PhyAddrPointer_reg[29]/NET0131 ,
		_w1213_,
		_w1447_
	);
	LUT3 #(
		.INIT('h48)
	) name995 (
		\PhyAddrPointer_reg[29]/NET0131 ,
		_w1212_,
		_w1213_,
		_w1448_
	);
	LUT4 #(
		.INIT('h8848)
	) name996 (
		\PhyAddrPointer_reg[29]/NET0131 ,
		_w695_,
		_w1207_,
		_w1209_,
		_w1449_
	);
	LUT4 #(
		.INIT('h3f15)
	) name997 (
		\PhyAddrPointer_reg[29]/NET0131 ,
		\rEIP_reg[29]/NET0131 ,
		_w1080_,
		_w1215_,
		_w1450_
	);
	LUT3 #(
		.INIT('h10)
	) name998 (
		_w1449_,
		_w1448_,
		_w1450_,
		_w1451_
	);
	LUT4 #(
		.INIT('h8aff)
	) name999 (
		_w690_,
		_w1444_,
		_w1446_,
		_w1451_,
		_w1452_
	);
	LUT3 #(
		.INIT('h08)
	) name1000 (
		\InstAddrPointer_reg[8]/NET0131 ,
		_w563_,
		_w673_,
		_w1453_
	);
	LUT4 #(
		.INIT('h0132)
	) name1001 (
		_w918_,
		_w836_,
		_w948_,
		_w958_,
		_w1454_
	);
	LUT4 #(
		.INIT('h5115)
	) name1002 (
		_w674_,
		_w836_,
		_w839_,
		_w1270_,
		_w1455_
	);
	LUT4 #(
		.INIT('h8a88)
	) name1003 (
		_w608_,
		_w1453_,
		_w1454_,
		_w1455_,
		_w1456_
	);
	LUT4 #(
		.INIT('ha082)
	) name1004 (
		_w671_,
		_w1014_,
		_w1015_,
		_w1039_,
		_w1457_
	);
	LUT2 #(
		.INIT('h4)
	) name1005 (
		_w597_,
		_w839_,
		_w1458_
	);
	LUT2 #(
		.INIT('h8)
	) name1006 (
		_w635_,
		_w1015_,
		_w1459_
	);
	LUT4 #(
		.INIT('h004f)
	) name1007 (
		_w616_,
		_w630_,
		_w958_,
		_w1459_,
		_w1460_
	);
	LUT4 #(
		.INIT('h0d00)
	) name1008 (
		\InstAddrPointer_reg[8]/NET0131 ,
		_w1165_,
		_w1458_,
		_w1460_,
		_w1461_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name1009 (
		_w690_,
		_w1456_,
		_w1457_,
		_w1461_,
		_w1462_
	);
	LUT4 #(
		.INIT('h153f)
	) name1010 (
		\InstAddrPointer_reg[8]/NET0131 ,
		\rEIP_reg[8]/NET0131 ,
		_w1080_,
		_w1081_,
		_w1463_
	);
	LUT2 #(
		.INIT('hb)
	) name1011 (
		_w1462_,
		_w1463_,
		_w1464_
	);
	LUT3 #(
		.INIT('h08)
	) name1012 (
		\InstAddrPointer_reg[13]/NET0131 ,
		_w563_,
		_w673_,
		_w1465_
	);
	LUT3 #(
		.INIT('h6a)
	) name1013 (
		\InstAddrPointer_reg[13]/NET0131 ,
		_w726_,
		_w727_,
		_w1466_
	);
	LUT4 #(
		.INIT('hf800)
	) name1014 (
		_w825_,
		_w870_,
		_w876_,
		_w890_,
		_w1467_
	);
	LUT4 #(
		.INIT('h6a00)
	) name1015 (
		\InstAddrPointer_reg[10]/NET0131 ,
		_w723_,
		_w724_,
		_w727_,
		_w1468_
	);
	LUT4 #(
		.INIT('h8222)
	) name1016 (
		_w836_,
		_w1466_,
		_w1467_,
		_w1468_,
		_w1469_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name1017 (
		_w962_,
		_w957_,
		_w1089_,
		_w1092_,
		_w1470_
	);
	LUT2 #(
		.INIT('h1)
	) name1018 (
		_w836_,
		_w1470_,
		_w1471_
	);
	LUT4 #(
		.INIT('h1055)
	) name1019 (
		_w674_,
		_w962_,
		_w1336_,
		_w1471_,
		_w1472_
	);
	LUT4 #(
		.INIT('h8a88)
	) name1020 (
		_w608_,
		_w1465_,
		_w1469_,
		_w1472_,
		_w1473_
	);
	LUT4 #(
		.INIT('h1333)
	) name1021 (
		\InstAddrPointer_reg[12]/NET0131 ,
		\InstAddrPointer_reg[13]/NET0131 ,
		_w885_,
		_w1041_,
		_w1474_
	);
	LUT2 #(
		.INIT('h1)
	) name1022 (
		_w1007_,
		_w1474_,
		_w1475_
	);
	LUT3 #(
		.INIT('h07)
	) name1023 (
		\InstAddrPointer_reg[12]/NET0131 ,
		_w1321_,
		_w1475_,
		_w1476_
	);
	LUT4 #(
		.INIT('h70f0)
	) name1024 (
		\InstAddrPointer_reg[12]/NET0131 ,
		\InstAddrPointer_reg[13]/NET0131 ,
		_w671_,
		_w1321_,
		_w1477_
	);
	LUT4 #(
		.INIT('ha8a0)
	) name1025 (
		\InstAddrPointer_reg[13]/NET0131 ,
		_w585_,
		_w589_,
		_w590_,
		_w1478_
	);
	LUT3 #(
		.INIT('hc4)
	) name1026 (
		_w597_,
		_w1466_,
		_w1478_,
		_w1479_
	);
	LUT4 #(
		.INIT('haa8a)
	) name1027 (
		\InstAddrPointer_reg[13]/NET0131 ,
		_w613_,
		_w681_,
		_w1368_,
		_w1480_
	);
	LUT2 #(
		.INIT('h8)
	) name1028 (
		_w635_,
		_w1475_,
		_w1481_
	);
	LUT4 #(
		.INIT('h004f)
	) name1029 (
		_w616_,
		_w630_,
		_w962_,
		_w1481_,
		_w1482_
	);
	LUT3 #(
		.INIT('h10)
	) name1030 (
		_w1480_,
		_w1479_,
		_w1482_,
		_w1483_
	);
	LUT3 #(
		.INIT('hb0)
	) name1031 (
		_w1476_,
		_w1477_,
		_w1483_,
		_w1484_
	);
	LUT4 #(
		.INIT('h153f)
	) name1032 (
		\InstAddrPointer_reg[13]/NET0131 ,
		\rEIP_reg[13]/NET0131 ,
		_w1080_,
		_w1081_,
		_w1485_
	);
	LUT4 #(
		.INIT('h8aff)
	) name1033 (
		_w690_,
		_w1473_,
		_w1484_,
		_w1485_,
		_w1486_
	);
	LUT3 #(
		.INIT('h08)
	) name1034 (
		\PhyAddrPointer_reg[11]/NET0131 ,
		_w563_,
		_w673_,
		_w1487_
	);
	LUT4 #(
		.INIT('h202a)
	) name1035 (
		\PhyAddrPointer_reg[11]/NET0131 ,
		_w634_,
		_w607_,
		_w608_,
		_w1488_
	);
	LUT4 #(
		.INIT('h00fd)
	) name1036 (
		_w671_,
		_w1321_,
		_w1320_,
		_w1488_,
		_w1489_
	);
	LUT4 #(
		.INIT('h5700)
	) name1037 (
		_w608_,
		_w1318_,
		_w1487_,
		_w1489_,
		_w1490_
	);
	LUT4 #(
		.INIT('h8000)
	) name1038 (
		\PhyAddrPointer_reg[10]/NET0131 ,
		\PhyAddrPointer_reg[11]/NET0131 ,
		\PhyAddrPointer_reg[9]/NET0131 ,
		_w1194_,
		_w1491_
	);
	LUT4 #(
		.INIT('h7f2a)
	) name1039 (
		\PhyAddrPointer_reg[11]/NET0131 ,
		\PhyAddrPointer_reg[1]/NET0131 ,
		_w1195_,
		_w1387_,
		_w1492_
	);
	LUT4 #(
		.INIT('h3f15)
	) name1040 (
		\PhyAddrPointer_reg[11]/NET0131 ,
		\rEIP_reg[11]/NET0131 ,
		_w1080_,
		_w1215_,
		_w1493_
	);
	LUT4 #(
		.INIT('hb700)
	) name1041 (
		\PhyAddrPointer_reg[11]/NET0131 ,
		_w714_,
		_w1195_,
		_w1493_,
		_w1494_
	);
	LUT3 #(
		.INIT('h70)
	) name1042 (
		_w1306_,
		_w1492_,
		_w1494_,
		_w1495_
	);
	LUT3 #(
		.INIT('h2f)
	) name1043 (
		_w690_,
		_w1490_,
		_w1495_,
		_w1496_
	);
	LUT3 #(
		.INIT('h08)
	) name1044 (
		\PhyAddrPointer_reg[14]/NET0131 ,
		_w563_,
		_w673_,
		_w1497_
	);
	LUT4 #(
		.INIT('h202a)
	) name1045 (
		\PhyAddrPointer_reg[14]/NET0131 ,
		_w634_,
		_w607_,
		_w608_,
		_w1498_
	);
	LUT2 #(
		.INIT('h1)
	) name1046 (
		_w1344_,
		_w1498_,
		_w1499_
	);
	LUT4 #(
		.INIT('h5700)
	) name1047 (
		_w608_,
		_w1339_,
		_w1497_,
		_w1499_,
		_w1500_
	);
	LUT3 #(
		.INIT('h6a)
	) name1048 (
		\PhyAddrPointer_reg[14]/NET0131 ,
		_w1197_,
		_w1387_,
		_w1501_
	);
	LUT4 #(
		.INIT('h4111)
	) name1049 (
		\DataWidth_reg[1]/NET0131 ,
		\PhyAddrPointer_reg[14]/NET0131 ,
		_w1197_,
		_w1387_,
		_w1502_
	);
	LUT4 #(
		.INIT('h70d0)
	) name1050 (
		\DataWidth_reg[1]/NET0131 ,
		\PhyAddrPointer_reg[14]/NET0131 ,
		_w695_,
		_w1198_,
		_w1503_
	);
	LUT4 #(
		.INIT('h4888)
	) name1051 (
		\PhyAddrPointer_reg[14]/NET0131 ,
		_w1212_,
		_w1197_,
		_w1387_,
		_w1504_
	);
	LUT4 #(
		.INIT('h3f15)
	) name1052 (
		\PhyAddrPointer_reg[14]/NET0131 ,
		\rEIP_reg[14]/NET0131 ,
		_w1080_,
		_w1215_,
		_w1505_
	);
	LUT4 #(
		.INIT('h4500)
	) name1053 (
		_w1504_,
		_w1502_,
		_w1503_,
		_w1505_,
		_w1506_
	);
	LUT3 #(
		.INIT('h2f)
	) name1054 (
		_w690_,
		_w1500_,
		_w1506_,
		_w1507_
	);
	LUT3 #(
		.INIT('h08)
	) name1055 (
		\PhyAddrPointer_reg[19]/NET0131 ,
		_w563_,
		_w673_,
		_w1508_
	);
	LUT4 #(
		.INIT('h1555)
	) name1056 (
		_w884_,
		_w883_,
		_w1132_,
		_w1137_,
		_w1509_
	);
	LUT3 #(
		.INIT('ha8)
	) name1057 (
		_w836_,
		_w1272_,
		_w1509_,
		_w1510_
	);
	LUT3 #(
		.INIT('h02)
	) name1058 (
		_w972_,
		_w975_,
		_w976_,
		_w1511_
	);
	LUT3 #(
		.INIT('h2a)
	) name1059 (
		_w974_,
		_w1147_,
		_w1511_,
		_w1512_
	);
	LUT3 #(
		.INIT('h15)
	) name1060 (
		_w836_,
		_w978_,
		_w1147_,
		_w1513_
	);
	LUT3 #(
		.INIT('h45)
	) name1061 (
		_w674_,
		_w1512_,
		_w1513_,
		_w1514_
	);
	LUT4 #(
		.INIT('h8a88)
	) name1062 (
		_w608_,
		_w1508_,
		_w1510_,
		_w1514_,
		_w1515_
	);
	LUT4 #(
		.INIT('h202a)
	) name1063 (
		\PhyAddrPointer_reg[19]/NET0131 ,
		_w634_,
		_w607_,
		_w608_,
		_w1516_
	);
	LUT3 #(
		.INIT('h28)
	) name1064 (
		_w671_,
		_w1061_,
		_w1159_,
		_w1517_
	);
	LUT4 #(
		.INIT('h00d7)
	) name1065 (
		_w671_,
		_w1061_,
		_w1159_,
		_w1516_,
		_w1518_
	);
	LUT4 #(
		.INIT('h8000)
	) name1066 (
		\PhyAddrPointer_reg[14]/NET0131 ,
		\PhyAddrPointer_reg[18]/NET0131 ,
		_w1198_,
		_w1200_,
		_w1519_
	);
	LUT4 #(
		.INIT('h8000)
	) name1067 (
		\PhyAddrPointer_reg[14]/NET0131 ,
		_w1198_,
		_w1200_,
		_w1202_,
		_w1520_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name1068 (
		\PhyAddrPointer_reg[18]/NET0131 ,
		\PhyAddrPointer_reg[19]/NET0131 ,
		\PhyAddrPointer_reg[1]/NET0131 ,
		_w1201_,
		_w1521_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name1069 (
		\PhyAddrPointer_reg[19]/NET0131 ,
		_w714_,
		_w1215_,
		_w1519_,
		_w1522_
	);
	LUT3 #(
		.INIT('h20)
	) name1070 (
		\DataWidth_reg[1]/NET0131 ,
		\PhyAddrPointer_reg[19]/NET0131 ,
		_w695_,
		_w1523_
	);
	LUT2 #(
		.INIT('h8)
	) name1071 (
		\rEIP_reg[19]/NET0131 ,
		_w1080_,
		_w1524_
	);
	LUT3 #(
		.INIT('h07)
	) name1072 (
		_w1519_,
		_w1523_,
		_w1524_,
		_w1525_
	);
	LUT4 #(
		.INIT('h1300)
	) name1073 (
		_w1306_,
		_w1522_,
		_w1521_,
		_w1525_,
		_w1526_
	);
	LUT4 #(
		.INIT('h8aff)
	) name1074 (
		_w690_,
		_w1515_,
		_w1518_,
		_w1526_,
		_w1527_
	);
	LUT3 #(
		.INIT('h08)
	) name1075 (
		\PhyAddrPointer_reg[22]/NET0131 ,
		_w563_,
		_w673_,
		_w1528_
	);
	LUT4 #(
		.INIT('haa20)
	) name1076 (
		_w608_,
		_w1237_,
		_w1238_,
		_w1528_,
		_w1529_
	);
	LUT4 #(
		.INIT('h202a)
	) name1077 (
		\PhyAddrPointer_reg[22]/NET0131 ,
		_w634_,
		_w607_,
		_w608_,
		_w1530_
	);
	LUT3 #(
		.INIT('h0b)
	) name1078 (
		_w1241_,
		_w1242_,
		_w1530_,
		_w1531_
	);
	LUT3 #(
		.INIT('h6a)
	) name1079 (
		\PhyAddrPointer_reg[22]/NET0131 ,
		_w1203_,
		_w1405_,
		_w1532_
	);
	LUT4 #(
		.INIT('h4111)
	) name1080 (
		\DataWidth_reg[1]/NET0131 ,
		\PhyAddrPointer_reg[22]/NET0131 ,
		_w1203_,
		_w1405_,
		_w1533_
	);
	LUT4 #(
		.INIT('h70d0)
	) name1081 (
		\DataWidth_reg[1]/NET0131 ,
		\PhyAddrPointer_reg[22]/NET0131 ,
		_w695_,
		_w1204_,
		_w1534_
	);
	LUT4 #(
		.INIT('h4888)
	) name1082 (
		\PhyAddrPointer_reg[22]/NET0131 ,
		_w1212_,
		_w1203_,
		_w1405_,
		_w1535_
	);
	LUT4 #(
		.INIT('h3f15)
	) name1083 (
		\PhyAddrPointer_reg[22]/NET0131 ,
		\rEIP_reg[22]/NET0131 ,
		_w1080_,
		_w1215_,
		_w1536_
	);
	LUT4 #(
		.INIT('h4500)
	) name1084 (
		_w1535_,
		_w1533_,
		_w1534_,
		_w1536_,
		_w1537_
	);
	LUT4 #(
		.INIT('h8aff)
	) name1085 (
		_w690_,
		_w1529_,
		_w1531_,
		_w1537_,
		_w1538_
	);
	LUT3 #(
		.INIT('h08)
	) name1086 (
		\PhyAddrPointer_reg[24]/NET0131 ,
		_w563_,
		_w673_,
		_w1539_
	);
	LUT4 #(
		.INIT('haa20)
	) name1087 (
		_w608_,
		_w1263_,
		_w1275_,
		_w1539_,
		_w1540_
	);
	LUT4 #(
		.INIT('h202a)
	) name1088 (
		\PhyAddrPointer_reg[24]/NET0131 ,
		_w634_,
		_w607_,
		_w608_,
		_w1541_
	);
	LUT4 #(
		.INIT('h00d7)
	) name1089 (
		_w671_,
		_w1059_,
		_w1256_,
		_w1541_,
		_w1542_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name1090 (
		\PhyAddrPointer_reg[24]/NET0131 ,
		_w1188_,
		_w1203_,
		_w1405_,
		_w1543_
	);
	LUT2 #(
		.INIT('h8)
	) name1091 (
		_w1306_,
		_w1543_,
		_w1544_
	);
	LUT4 #(
		.INIT('h070f)
	) name1092 (
		\PhyAddrPointer_reg[22]/NET0131 ,
		\PhyAddrPointer_reg[23]/NET0131 ,
		\PhyAddrPointer_reg[24]/NET0131 ,
		_w1204_,
		_w1545_
	);
	LUT3 #(
		.INIT('h2a)
	) name1093 (
		_w714_,
		_w1189_,
		_w1204_,
		_w1546_
	);
	LUT4 #(
		.INIT('h3f15)
	) name1094 (
		\PhyAddrPointer_reg[24]/NET0131 ,
		\rEIP_reg[24]/NET0131 ,
		_w1080_,
		_w1215_,
		_w1547_
	);
	LUT3 #(
		.INIT('hb0)
	) name1095 (
		_w1545_,
		_w1546_,
		_w1547_,
		_w1548_
	);
	LUT2 #(
		.INIT('h4)
	) name1096 (
		_w1544_,
		_w1548_,
		_w1549_
	);
	LUT4 #(
		.INIT('h8aff)
	) name1097 (
		_w690_,
		_w1540_,
		_w1542_,
		_w1549_,
		_w1550_
	);
	LUT3 #(
		.INIT('h08)
	) name1098 (
		\PhyAddrPointer_reg[26]/NET0131 ,
		_w563_,
		_w673_,
		_w1551_
	);
	LUT4 #(
		.INIT('haa20)
	) name1099 (
		_w608_,
		_w1287_,
		_w1288_,
		_w1551_,
		_w1552_
	);
	LUT4 #(
		.INIT('h202a)
	) name1100 (
		\PhyAddrPointer_reg[26]/NET0131 ,
		_w634_,
		_w607_,
		_w608_,
		_w1553_
	);
	LUT2 #(
		.INIT('h1)
	) name1101 (
		_w1290_,
		_w1553_,
		_w1554_
	);
	LUT4 #(
		.INIT('h8000)
	) name1102 (
		\PhyAddrPointer_reg[1]/NET0131 ,
		\PhyAddrPointer_reg[25]/NET0131 ,
		_w1189_,
		_w1204_,
		_w1555_
	);
	LUT3 #(
		.INIT('h6c)
	) name1103 (
		\PhyAddrPointer_reg[1]/NET0131 ,
		\PhyAddrPointer_reg[26]/NET0131 ,
		_w1205_,
		_w1556_
	);
	LUT4 #(
		.INIT('h6c00)
	) name1104 (
		\PhyAddrPointer_reg[1]/NET0131 ,
		\PhyAddrPointer_reg[26]/NET0131 ,
		_w1205_,
		_w1306_,
		_w1557_
	);
	LUT4 #(
		.INIT('h3f15)
	) name1105 (
		\PhyAddrPointer_reg[26]/NET0131 ,
		\rEIP_reg[26]/NET0131 ,
		_w1080_,
		_w1215_,
		_w1558_
	);
	LUT4 #(
		.INIT('hb700)
	) name1106 (
		\PhyAddrPointer_reg[26]/NET0131 ,
		_w714_,
		_w1205_,
		_w1558_,
		_w1559_
	);
	LUT2 #(
		.INIT('h4)
	) name1107 (
		_w1557_,
		_w1559_,
		_w1560_
	);
	LUT4 #(
		.INIT('h8aff)
	) name1108 (
		_w690_,
		_w1552_,
		_w1554_,
		_w1560_,
		_w1561_
	);
	LUT3 #(
		.INIT('h87)
	) name1109 (
		_w830_,
		_w835_,
		_w837_,
		_w1562_
	);
	LUT4 #(
		.INIT('h8f70)
	) name1110 (
		_w825_,
		_w869_,
		_w874_,
		_w1562_,
		_w1563_
	);
	LUT4 #(
		.INIT('h808c)
	) name1111 (
		\InstAddrPointer_reg[7]/NET0131 ,
		_w608_,
		_w674_,
		_w1563_,
		_w1564_
	);
	LUT3 #(
		.INIT('h87)
	) name1112 (
		_w830_,
		_w835_,
		_w1013_,
		_w1565_
	);
	LUT4 #(
		.INIT('h2f00)
	) name1113 (
		_w1021_,
		_w1106_,
		_w1107_,
		_w1565_,
		_w1566_
	);
	LUT4 #(
		.INIT('h00d0)
	) name1114 (
		_w1021_,
		_w1106_,
		_w1107_,
		_w1565_,
		_w1567_
	);
	LUT3 #(
		.INIT('h02)
	) name1115 (
		_w671_,
		_w1567_,
		_w1566_,
		_w1568_
	);
	LUT3 #(
		.INIT('h80)
	) name1116 (
		READY_n_pad,
		_w494_,
		_w586_,
		_w1569_
	);
	LUT4 #(
		.INIT('haa8a)
	) name1117 (
		\InstAddrPointer_reg[7]/NET0131 ,
		_w613_,
		_w681_,
		_w1569_,
		_w1570_
	);
	LUT3 #(
		.INIT('hb0)
	) name1118 (
		_w616_,
		_w630_,
		_w918_,
		_w1571_
	);
	LUT4 #(
		.INIT('h00ec)
	) name1119 (
		_w585_,
		_w589_,
		_w590_,
		_w594_,
		_w1572_
	);
	LUT3 #(
		.INIT('hb8)
	) name1120 (
		\InstAddrPointer_reg[7]/NET0131 ,
		READY_n_pad,
		_w837_,
		_w1573_
	);
	LUT3 #(
		.INIT('hd0)
	) name1121 (
		_w563_,
		_w565_,
		_w1573_,
		_w1574_
	);
	LUT3 #(
		.INIT('he0)
	) name1122 (
		_w582_,
		_w1572_,
		_w1574_,
		_w1575_
	);
	LUT4 #(
		.INIT('h070f)
	) name1123 (
		_w494_,
		_w586_,
		_w554_,
		_w652_,
		_w1576_
	);
	LUT4 #(
		.INIT('h5f13)
	) name1124 (
		_w635_,
		_w837_,
		_w1013_,
		_w1576_,
		_w1577_
	);
	LUT2 #(
		.INIT('h4)
	) name1125 (
		_w1575_,
		_w1577_,
		_w1578_
	);
	LUT4 #(
		.INIT('h0100)
	) name1126 (
		_w1570_,
		_w1568_,
		_w1571_,
		_w1578_,
		_w1579_
	);
	LUT4 #(
		.INIT('h153f)
	) name1127 (
		\InstAddrPointer_reg[7]/NET0131 ,
		\rEIP_reg[7]/NET0131 ,
		_w1080_,
		_w1081_,
		_w1580_
	);
	LUT4 #(
		.INIT('h8aff)
	) name1128 (
		_w690_,
		_w1564_,
		_w1579_,
		_w1580_,
		_w1581_
	);
	LUT3 #(
		.INIT('h08)
	) name1129 (
		\InstAddrPointer_reg[9]/NET0131 ,
		_w563_,
		_w673_,
		_w1582_
	);
	LUT4 #(
		.INIT('h07f8)
	) name1130 (
		_w825_,
		_w870_,
		_w876_,
		_w890_,
		_w1583_
	);
	LUT4 #(
		.INIT('h1411)
	) name1131 (
		_w836_,
		_w952_,
		_w1089_,
		_w1092_,
		_w1584_
	);
	LUT4 #(
		.INIT('h0501)
	) name1132 (
		_w674_,
		_w836_,
		_w1584_,
		_w1583_,
		_w1585_
	);
	LUT3 #(
		.INIT('ha8)
	) name1133 (
		_w608_,
		_w1582_,
		_w1585_,
		_w1586_
	);
	LUT4 #(
		.INIT('ha028)
	) name1134 (
		_w671_,
		_w1016_,
		_w1044_,
		_w1109_,
		_w1587_
	);
	LUT2 #(
		.INIT('h4)
	) name1135 (
		_w597_,
		_w890_,
		_w1588_
	);
	LUT3 #(
		.INIT('hb0)
	) name1136 (
		_w616_,
		_w630_,
		_w952_,
		_w1589_
	);
	LUT2 #(
		.INIT('h8)
	) name1137 (
		_w635_,
		_w1044_,
		_w1590_
	);
	LUT3 #(
		.INIT('h0d)
	) name1138 (
		\InstAddrPointer_reg[9]/NET0131 ,
		_w1295_,
		_w1590_,
		_w1591_
	);
	LUT4 #(
		.INIT('h0100)
	) name1139 (
		_w1588_,
		_w1589_,
		_w1587_,
		_w1591_,
		_w1592_
	);
	LUT4 #(
		.INIT('h153f)
	) name1140 (
		\InstAddrPointer_reg[9]/NET0131 ,
		\rEIP_reg[9]/NET0131 ,
		_w1080_,
		_w1081_,
		_w1593_
	);
	LUT4 #(
		.INIT('h8aff)
	) name1141 (
		_w690_,
		_w1586_,
		_w1592_,
		_w1593_,
		_w1594_
	);
	LUT3 #(
		.INIT('h08)
	) name1142 (
		\PhyAddrPointer_reg[13]/NET0131 ,
		_w563_,
		_w673_,
		_w1595_
	);
	LUT4 #(
		.INIT('haa20)
	) name1143 (
		_w608_,
		_w1469_,
		_w1472_,
		_w1595_,
		_w1596_
	);
	LUT4 #(
		.INIT('h202a)
	) name1144 (
		\PhyAddrPointer_reg[13]/NET0131 ,
		_w634_,
		_w607_,
		_w608_,
		_w1597_
	);
	LUT3 #(
		.INIT('h0b)
	) name1145 (
		_w1476_,
		_w1477_,
		_w1597_,
		_w1598_
	);
	LUT4 #(
		.INIT('h1333)
	) name1146 (
		\PhyAddrPointer_reg[12]/NET0131 ,
		\PhyAddrPointer_reg[13]/NET0131 ,
		\PhyAddrPointer_reg[1]/NET0131 ,
		_w1491_,
		_w1599_
	);
	LUT2 #(
		.INIT('h1)
	) name1147 (
		_w1388_,
		_w1599_,
		_w1600_
	);
	LUT3 #(
		.INIT('h02)
	) name1148 (
		_w1306_,
		_w1388_,
		_w1599_,
		_w1601_
	);
	LUT4 #(
		.INIT('h8000)
	) name1149 (
		\PhyAddrPointer_reg[10]/NET0131 ,
		\PhyAddrPointer_reg[9]/NET0131 ,
		_w1194_,
		_w1196_,
		_w1602_
	);
	LUT4 #(
		.INIT('h4888)
	) name1150 (
		\PhyAddrPointer_reg[13]/NET0131 ,
		_w714_,
		_w1195_,
		_w1196_,
		_w1603_
	);
	LUT4 #(
		.INIT('h3f15)
	) name1151 (
		\PhyAddrPointer_reg[13]/NET0131 ,
		\rEIP_reg[13]/NET0131 ,
		_w1080_,
		_w1215_,
		_w1604_
	);
	LUT2 #(
		.INIT('h4)
	) name1152 (
		_w1603_,
		_w1604_,
		_w1605_
	);
	LUT2 #(
		.INIT('h4)
	) name1153 (
		_w1601_,
		_w1605_,
		_w1606_
	);
	LUT4 #(
		.INIT('h8aff)
	) name1154 (
		_w690_,
		_w1596_,
		_w1598_,
		_w1606_,
		_w1607_
	);
	LUT3 #(
		.INIT('h08)
	) name1155 (
		\PhyAddrPointer_reg[16]/NET0131 ,
		_w563_,
		_w673_,
		_w1608_
	);
	LUT4 #(
		.INIT('h0080)
	) name1156 (
		_w881_,
		_w1132_,
		_w1135_,
		_w1270_,
		_w1609_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name1157 (
		\InstAddrPointer_reg[16]/NET0131 ,
		_w726_,
		_w728_,
		_w730_,
		_w1610_
	);
	LUT4 #(
		.INIT('h808c)
	) name1158 (
		\InstAddrPointer_reg[16]/NET0131 ,
		_w836_,
		_w1609_,
		_w1610_,
		_w1611_
	);
	LUT4 #(
		.INIT('hfb00)
	) name1159 (
		_w948_,
		_w964_,
		_w970_,
		_w971_,
		_w1612_
	);
	LUT4 #(
		.INIT('h4555)
	) name1160 (
		_w836_,
		_w948_,
		_w964_,
		_w972_,
		_w1613_
	);
	LUT3 #(
		.INIT('h45)
	) name1161 (
		_w674_,
		_w1612_,
		_w1613_,
		_w1614_
	);
	LUT4 #(
		.INIT('h8a88)
	) name1162 (
		_w608_,
		_w1608_,
		_w1611_,
		_w1614_,
		_w1615_
	);
	LUT4 #(
		.INIT('h202a)
	) name1163 (
		\PhyAddrPointer_reg[16]/NET0131 ,
		_w634_,
		_w607_,
		_w608_,
		_w1616_
	);
	LUT4 #(
		.INIT('h00df)
	) name1164 (
		_w1016_,
		_w1039_,
		_w1048_,
		_w1156_,
		_w1617_
	);
	LUT3 #(
		.INIT('h02)
	) name1165 (
		_w671_,
		_w1255_,
		_w1617_,
		_w1618_
	);
	LUT4 #(
		.INIT('h00d7)
	) name1166 (
		_w671_,
		_w1156_,
		_w1254_,
		_w1616_,
		_w1619_
	);
	LUT4 #(
		.INIT('h8000)
	) name1167 (
		\PhyAddrPointer_reg[14]/NET0131 ,
		_w1197_,
		_w1199_,
		_w1387_,
		_w1620_
	);
	LUT3 #(
		.INIT('h6c)
	) name1168 (
		\PhyAddrPointer_reg[15]/NET0131 ,
		\PhyAddrPointer_reg[16]/NET0131 ,
		_w1389_,
		_w1621_
	);
	LUT4 #(
		.INIT('h60c0)
	) name1169 (
		\PhyAddrPointer_reg[15]/NET0131 ,
		\PhyAddrPointer_reg[16]/NET0131 ,
		_w1306_,
		_w1389_,
		_w1622_
	);
	LUT4 #(
		.INIT('h8000)
	) name1170 (
		\PhyAddrPointer_reg[14]/NET0131 ,
		\PhyAddrPointer_reg[15]/NET0131 ,
		\PhyAddrPointer_reg[16]/NET0131 ,
		_w1198_,
		_w1623_
	);
	LUT4 #(
		.INIT('h3f15)
	) name1171 (
		\PhyAddrPointer_reg[16]/NET0131 ,
		\rEIP_reg[16]/NET0131 ,
		_w1080_,
		_w1215_,
		_w1624_
	);
	LUT4 #(
		.INIT('hb700)
	) name1172 (
		\PhyAddrPointer_reg[16]/NET0131 ,
		_w714_,
		_w1383_,
		_w1624_,
		_w1625_
	);
	LUT2 #(
		.INIT('h4)
	) name1173 (
		_w1622_,
		_w1625_,
		_w1626_
	);
	LUT4 #(
		.INIT('h8aff)
	) name1174 (
		_w690_,
		_w1615_,
		_w1619_,
		_w1626_,
		_w1627_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name1175 (
		\InstAddrPointer_reg[17]/NET0131 ,
		_w726_,
		_w728_,
		_w731_,
		_w1628_
	);
	LUT4 #(
		.INIT('h8000)
	) name1176 (
		\InstAddrPointer_reg[16]/NET0131 ,
		_w885_,
		_w888_,
		_w881_,
		_w1629_
	);
	LUT4 #(
		.INIT('h820a)
	) name1177 (
		_w836_,
		_w1467_,
		_w1628_,
		_w1629_,
		_w1630_
	);
	LUT4 #(
		.INIT('h2000)
	) name1178 (
		_w957_,
		_w1089_,
		_w1092_,
		_w1093_,
		_w1631_
	);
	LUT4 #(
		.INIT('h4554)
	) name1179 (
		_w674_,
		_w836_,
		_w975_,
		_w1631_,
		_w1632_
	);
	LUT3 #(
		.INIT('h20)
	) name1180 (
		_w608_,
		_w1630_,
		_w1632_,
		_w1633_
	);
	LUT4 #(
		.INIT('h08b8)
	) name1181 (
		_w634_,
		_w607_,
		_w608_,
		_w674_,
		_w1634_
	);
	LUT2 #(
		.INIT('h2)
	) name1182 (
		\PhyAddrPointer_reg[17]/NET0131 ,
		_w1634_,
		_w1635_
	);
	LUT4 #(
		.INIT('h0080)
	) name1183 (
		_w1016_,
		_w1040_,
		_w1050_,
		_w1109_,
		_w1636_
	);
	LUT4 #(
		.INIT('h3313)
	) name1184 (
		_w1016_,
		_w1040_,
		_w1050_,
		_w1109_,
		_w1637_
	);
	LUT3 #(
		.INIT('h02)
	) name1185 (
		_w671_,
		_w1637_,
		_w1636_,
		_w1638_
	);
	LUT4 #(
		.INIT('h00d7)
	) name1186 (
		_w671_,
		_w1040_,
		_w1110_,
		_w1635_,
		_w1639_
	);
	LUT3 #(
		.INIT('h32)
	) name1187 (
		\PhyAddrPointer_reg[17]/NET0131 ,
		_w1405_,
		_w1620_,
		_w1640_
	);
	LUT4 #(
		.INIT('h0c08)
	) name1188 (
		\PhyAddrPointer_reg[17]/NET0131 ,
		_w1306_,
		_w1405_,
		_w1620_,
		_w1641_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name1189 (
		\PhyAddrPointer_reg[14]/NET0131 ,
		_w714_,
		_w1198_,
		_w1200_,
		_w1642_
	);
	LUT4 #(
		.INIT('h3f15)
	) name1190 (
		\PhyAddrPointer_reg[17]/NET0131 ,
		\rEIP_reg[17]/NET0131 ,
		_w1080_,
		_w1215_,
		_w1643_
	);
	LUT4 #(
		.INIT('h1f00)
	) name1191 (
		\PhyAddrPointer_reg[17]/NET0131 ,
		_w1623_,
		_w1642_,
		_w1643_,
		_w1644_
	);
	LUT2 #(
		.INIT('h4)
	) name1192 (
		_w1641_,
		_w1644_,
		_w1645_
	);
	LUT4 #(
		.INIT('h8aff)
	) name1193 (
		_w690_,
		_w1633_,
		_w1639_,
		_w1645_,
		_w1646_
	);
	LUT3 #(
		.INIT('h08)
	) name1194 (
		\PhyAddrPointer_reg[18]/NET0131 ,
		_w563_,
		_w673_,
		_w1647_
	);
	LUT4 #(
		.INIT('h8222)
	) name1195 (
		_w836_,
		_w880_,
		_w882_,
		_w1285_,
		_w1648_
	);
	LUT3 #(
		.INIT('h8c)
	) name1196 (
		_w975_,
		_w976_,
		_w1631_,
		_w1649_
	);
	LUT3 #(
		.INIT('h15)
	) name1197 (
		_w836_,
		_w1147_,
		_w1511_,
		_w1650_
	);
	LUT3 #(
		.INIT('h45)
	) name1198 (
		_w674_,
		_w1649_,
		_w1650_,
		_w1651_
	);
	LUT4 #(
		.INIT('h8a88)
	) name1199 (
		_w608_,
		_w1647_,
		_w1648_,
		_w1651_,
		_w1652_
	);
	LUT4 #(
		.INIT('h202a)
	) name1200 (
		\PhyAddrPointer_reg[18]/NET0131 ,
		_w634_,
		_w607_,
		_w608_,
		_w1653_
	);
	LUT4 #(
		.INIT('h00df)
	) name1201 (
		_w1016_,
		_w1039_,
		_w1051_,
		_w1054_,
		_w1654_
	);
	LUT3 #(
		.INIT('h02)
	) name1202 (
		_w671_,
		_w1055_,
		_w1654_,
		_w1655_
	);
	LUT4 #(
		.INIT('h00d7)
	) name1203 (
		_w671_,
		_w1052_,
		_w1054_,
		_w1653_,
		_w1656_
	);
	LUT3 #(
		.INIT('h6a)
	) name1204 (
		\PhyAddrPointer_reg[18]/NET0131 ,
		\PhyAddrPointer_reg[1]/NET0131 ,
		_w1201_,
		_w1657_
	);
	LUT4 #(
		.INIT('h6a00)
	) name1205 (
		\PhyAddrPointer_reg[18]/NET0131 ,
		\PhyAddrPointer_reg[1]/NET0131 ,
		_w1201_,
		_w1306_,
		_w1658_
	);
	LUT4 #(
		.INIT('h3f15)
	) name1206 (
		\PhyAddrPointer_reg[18]/NET0131 ,
		\rEIP_reg[18]/NET0131 ,
		_w1080_,
		_w1215_,
		_w1659_
	);
	LUT4 #(
		.INIT('hb700)
	) name1207 (
		\PhyAddrPointer_reg[18]/NET0131 ,
		_w714_,
		_w1201_,
		_w1659_,
		_w1660_
	);
	LUT2 #(
		.INIT('h4)
	) name1208 (
		_w1658_,
		_w1660_,
		_w1661_
	);
	LUT4 #(
		.INIT('h8aff)
	) name1209 (
		_w690_,
		_w1652_,
		_w1656_,
		_w1661_,
		_w1662_
	);
	LUT3 #(
		.INIT('h08)
	) name1210 (
		\PhyAddrPointer_reg[21]/NET0131 ,
		_w563_,
		_w673_,
		_w1663_
	);
	LUT3 #(
		.INIT('h82)
	) name1211 (
		_w836_,
		_w894_,
		_w895_,
		_w1664_
	);
	LUT4 #(
		.INIT('h4554)
	) name1212 (
		_w674_,
		_w836_,
		_w966_,
		_w1096_,
		_w1665_
	);
	LUT4 #(
		.INIT('h8a88)
	) name1213 (
		_w608_,
		_w1663_,
		_w1664_,
		_w1665_,
		_w1666_
	);
	LUT4 #(
		.INIT('h202a)
	) name1214 (
		\PhyAddrPointer_reg[21]/NET0131 ,
		_w634_,
		_w607_,
		_w608_,
		_w1667_
	);
	LUT3 #(
		.INIT('h28)
	) name1215 (
		_w671_,
		_w1056_,
		_w1113_,
		_w1668_
	);
	LUT4 #(
		.INIT('h00d7)
	) name1216 (
		_w671_,
		_w1056_,
		_w1113_,
		_w1667_,
		_w1669_
	);
	LUT4 #(
		.INIT('h070f)
	) name1217 (
		\PhyAddrPointer_reg[1]/NET0131 ,
		\PhyAddrPointer_reg[20]/NET0131 ,
		\PhyAddrPointer_reg[21]/NET0131 ,
		_w1520_,
		_w1670_
	);
	LUT2 #(
		.INIT('h1)
	) name1218 (
		_w1406_,
		_w1670_,
		_w1671_
	);
	LUT3 #(
		.INIT('h02)
	) name1219 (
		_w1212_,
		_w1406_,
		_w1670_,
		_w1672_
	);
	LUT4 #(
		.INIT('h3133)
	) name1220 (
		\PhyAddrPointer_reg[20]/NET0131 ,
		\PhyAddrPointer_reg[21]/NET0131 ,
		_w1209_,
		_w1520_,
		_w1673_
	);
	LUT3 #(
		.INIT('ha2)
	) name1221 (
		_w695_,
		_w1204_,
		_w1209_,
		_w1674_
	);
	LUT4 #(
		.INIT('h3f15)
	) name1222 (
		\PhyAddrPointer_reg[21]/NET0131 ,
		\rEIP_reg[21]/NET0131 ,
		_w1080_,
		_w1215_,
		_w1675_
	);
	LUT3 #(
		.INIT('hb0)
	) name1223 (
		_w1673_,
		_w1674_,
		_w1675_,
		_w1676_
	);
	LUT2 #(
		.INIT('h4)
	) name1224 (
		_w1672_,
		_w1676_,
		_w1677_
	);
	LUT4 #(
		.INIT('h8aff)
	) name1225 (
		_w690_,
		_w1666_,
		_w1669_,
		_w1677_,
		_w1678_
	);
	LUT3 #(
		.INIT('h08)
	) name1226 (
		\PhyAddrPointer_reg[25]/NET0131 ,
		_w563_,
		_w673_,
		_w1679_
	);
	LUT4 #(
		.INIT('haa20)
	) name1227 (
		_w608_,
		_w1360_,
		_w1365_,
		_w1679_,
		_w1680_
	);
	LUT4 #(
		.INIT('h202a)
	) name1228 (
		\PhyAddrPointer_reg[25]/NET0131 ,
		_w634_,
		_w607_,
		_w608_,
		_w1681_
	);
	LUT2 #(
		.INIT('h1)
	) name1229 (
		_w1367_,
		_w1681_,
		_w1682_
	);
	LUT4 #(
		.INIT('h1555)
	) name1230 (
		\PhyAddrPointer_reg[25]/NET0131 ,
		_w1189_,
		_w1203_,
		_w1405_,
		_w1683_
	);
	LUT2 #(
		.INIT('h1)
	) name1231 (
		_w1555_,
		_w1683_,
		_w1684_
	);
	LUT3 #(
		.INIT('h54)
	) name1232 (
		\DataWidth_reg[1]/NET0131 ,
		_w1555_,
		_w1683_,
		_w1685_
	);
	LUT4 #(
		.INIT('h8222)
	) name1233 (
		\DataWidth_reg[1]/NET0131 ,
		\PhyAddrPointer_reg[25]/NET0131 ,
		_w1189_,
		_w1204_,
		_w1686_
	);
	LUT2 #(
		.INIT('h2)
	) name1234 (
		_w695_,
		_w1686_,
		_w1687_
	);
	LUT4 #(
		.INIT('h3f15)
	) name1235 (
		\PhyAddrPointer_reg[25]/NET0131 ,
		\rEIP_reg[25]/NET0131 ,
		_w1080_,
		_w1215_,
		_w1688_
	);
	LUT4 #(
		.INIT('hfd00)
	) name1236 (
		_w1212_,
		_w1555_,
		_w1683_,
		_w1688_,
		_w1689_
	);
	LUT3 #(
		.INIT('hb0)
	) name1237 (
		_w1685_,
		_w1687_,
		_w1689_,
		_w1690_
	);
	LUT4 #(
		.INIT('h8aff)
	) name1238 (
		_w690_,
		_w1680_,
		_w1682_,
		_w1690_,
		_w1691_
	);
	LUT3 #(
		.INIT('h08)
	) name1239 (
		\PhyAddrPointer_reg[8]/NET0131 ,
		_w563_,
		_w673_,
		_w1692_
	);
	LUT4 #(
		.INIT('haa20)
	) name1240 (
		_w608_,
		_w1454_,
		_w1455_,
		_w1692_,
		_w1693_
	);
	LUT4 #(
		.INIT('h202a)
	) name1241 (
		\PhyAddrPointer_reg[8]/NET0131 ,
		_w634_,
		_w607_,
		_w608_,
		_w1694_
	);
	LUT2 #(
		.INIT('h1)
	) name1242 (
		_w1457_,
		_w1694_,
		_w1695_
	);
	LUT2 #(
		.INIT('h6)
	) name1243 (
		\PhyAddrPointer_reg[8]/NET0131 ,
		_w1386_,
		_w1696_
	);
	LUT3 #(
		.INIT('h48)
	) name1244 (
		\PhyAddrPointer_reg[8]/NET0131 ,
		_w1306_,
		_w1386_,
		_w1697_
	);
	LUT4 #(
		.INIT('h3f15)
	) name1245 (
		\PhyAddrPointer_reg[8]/NET0131 ,
		\rEIP_reg[8]/NET0131 ,
		_w1080_,
		_w1215_,
		_w1698_
	);
	LUT4 #(
		.INIT('hb700)
	) name1246 (
		\PhyAddrPointer_reg[8]/NET0131 ,
		_w714_,
		_w1193_,
		_w1698_,
		_w1699_
	);
	LUT2 #(
		.INIT('h4)
	) name1247 (
		_w1697_,
		_w1699_,
		_w1700_
	);
	LUT4 #(
		.INIT('h8aff)
	) name1248 (
		_w690_,
		_w1693_,
		_w1695_,
		_w1700_,
		_w1701_
	);
	LUT2 #(
		.INIT('h1)
	) name1249 (
		READY_n_pad,
		_w762_,
		_w1702_
	);
	LUT3 #(
		.INIT('h0e)
	) name1250 (
		_w588_,
		_w596_,
		_w1702_,
		_w1703_
	);
	LUT3 #(
		.INIT('h01)
	) name1251 (
		_w655_,
		_w612_,
		_w680_,
		_w1704_
	);
	LUT4 #(
		.INIT('h00ec)
	) name1252 (
		_w585_,
		_w589_,
		_w590_,
		_w721_,
		_w1705_
	);
	LUT4 #(
		.INIT('h0001)
	) name1253 (
		_w655_,
		_w612_,
		_w680_,
		_w1705_,
		_w1706_
	);
	LUT3 #(
		.INIT('h8a)
	) name1254 (
		\InstAddrPointer_reg[4]/NET0131 ,
		_w1703_,
		_w1706_,
		_w1707_
	);
	LUT2 #(
		.INIT('h4)
	) name1255 (
		_w597_,
		_w762_,
		_w1708_
	);
	LUT4 #(
		.INIT('ha9aa)
	) name1256 (
		\InstAddrPointer_reg[4]/NET0131 ,
		_w563_,
		_w633_,
		_w1004_,
		_w1709_
	);
	LUT4 #(
		.INIT('hc800)
	) name1257 (
		_w569_,
		_w602_,
		_w604_,
		_w1709_,
		_w1710_
	);
	LUT4 #(
		.INIT('h004f)
	) name1258 (
		_w616_,
		_w630_,
		_w941_,
		_w1710_,
		_w1711_
	);
	LUT4 #(
		.INIT('h807f)
	) name1259 (
		_w749_,
		_w754_,
		_w760_,
		_w762_,
		_w1712_
	);
	LUT4 #(
		.INIT('h2fd0)
	) name1260 (
		_w794_,
		_w820_,
		_w1264_,
		_w1712_,
		_w1713_
	);
	LUT4 #(
		.INIT('h808c)
	) name1261 (
		\InstAddrPointer_reg[4]/NET0131 ,
		_w608_,
		_w674_,
		_w1713_,
		_w1714_
	);
	LUT4 #(
		.INIT('h807f)
	) name1262 (
		_w749_,
		_w754_,
		_w760_,
		_w1022_,
		_w1715_
	);
	LUT4 #(
		.INIT('h4445)
	) name1263 (
		_w1025_,
		_w1027_,
		_w1028_,
		_w1031_,
		_w1716_
	);
	LUT3 #(
		.INIT('h28)
	) name1264 (
		_w671_,
		_w1715_,
		_w1716_,
		_w1717_
	);
	LUT2 #(
		.INIT('h1)
	) name1265 (
		_w1714_,
		_w1717_,
		_w1718_
	);
	LUT4 #(
		.INIT('h1000)
	) name1266 (
		_w1708_,
		_w1707_,
		_w1711_,
		_w1718_,
		_w1719_
	);
	LUT2 #(
		.INIT('h8)
	) name1267 (
		\rEIP_reg[4]/NET0131 ,
		_w1080_,
		_w1720_
	);
	LUT4 #(
		.INIT('h153f)
	) name1268 (
		\InstAddrPointer_reg[4]/NET0131 ,
		\rEIP_reg[4]/NET0131 ,
		_w1080_,
		_w1081_,
		_w1721_
	);
	LUT3 #(
		.INIT('h2f)
	) name1269 (
		_w690_,
		_w1719_,
		_w1721_,
		_w1722_
	);
	LUT4 #(
		.INIT('h807f)
	) name1270 (
		_w844_,
		_w849_,
		_w852_,
		_w854_,
		_w1723_
	);
	LUT4 #(
		.INIT('h8a20)
	) name1271 (
		_w836_,
		_w1266_,
		_w1267_,
		_w1723_,
		_w1724_
	);
	LUT4 #(
		.INIT('h807f)
	) name1272 (
		_w844_,
		_w849_,
		_w852_,
		_w920_,
		_w1725_
	);
	LUT4 #(
		.INIT('h4510)
	) name1273 (
		_w836_,
		_w944_,
		_w947_,
		_w1725_,
		_w1726_
	);
	LUT4 #(
		.INIT('h7774)
	) name1274 (
		\InstAddrPointer_reg[6]/NET0131 ,
		_w674_,
		_w1726_,
		_w1724_,
		_w1727_
	);
	LUT2 #(
		.INIT('h2)
	) name1275 (
		_w608_,
		_w1727_,
		_w1728_
	);
	LUT4 #(
		.INIT('h008a)
	) name1276 (
		_w1021_,
		_w1032_,
		_w1035_,
		_w1036_,
		_w1729_
	);
	LUT4 #(
		.INIT('h807f)
	) name1277 (
		_w844_,
		_w849_,
		_w852_,
		_w1017_,
		_w1730_
	);
	LUT4 #(
		.INIT('h00ba)
	) name1278 (
		_w1020_,
		_w1032_,
		_w1035_,
		_w1730_,
		_w1731_
	);
	LUT3 #(
		.INIT('h02)
	) name1279 (
		_w671_,
		_w1731_,
		_w1729_,
		_w1732_
	);
	LUT2 #(
		.INIT('h4)
	) name1280 (
		_w597_,
		_w854_,
		_w1733_
	);
	LUT2 #(
		.INIT('h8)
	) name1281 (
		_w635_,
		_w1017_,
		_w1734_
	);
	LUT4 #(
		.INIT('h004f)
	) name1282 (
		_w616_,
		_w630_,
		_w920_,
		_w1734_,
		_w1735_
	);
	LUT4 #(
		.INIT('h0d00)
	) name1283 (
		\InstAddrPointer_reg[6]/NET0131 ,
		_w1165_,
		_w1733_,
		_w1735_,
		_w1736_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name1284 (
		_w690_,
		_w1728_,
		_w1732_,
		_w1736_,
		_w1737_
	);
	LUT4 #(
		.INIT('h153f)
	) name1285 (
		\InstAddrPointer_reg[6]/NET0131 ,
		\rEIP_reg[6]/NET0131 ,
		_w1080_,
		_w1081_,
		_w1738_
	);
	LUT2 #(
		.INIT('hb)
	) name1286 (
		_w1737_,
		_w1738_,
		_w1739_
	);
	LUT3 #(
		.INIT('h80)
	) name1287 (
		_w602_,
		_w604_,
		_w634_,
		_w1740_
	);
	LUT2 #(
		.INIT('h8)
	) name1288 (
		_w518_,
		_w617_,
		_w1741_
	);
	LUT4 #(
		.INIT('h0a0e)
	) name1289 (
		_w605_,
		_w587_,
		_w1740_,
		_w1741_,
		_w1742_
	);
	LUT4 #(
		.INIT('h8000)
	) name1290 (
		\EAX_reg[0]/NET0131 ,
		\EAX_reg[1]/NET0131 ,
		\EAX_reg[2]/NET0131 ,
		\EAX_reg[3]/NET0131 ,
		_w1743_
	);
	LUT4 #(
		.INIT('h8000)
	) name1291 (
		\EAX_reg[4]/NET0131 ,
		\EAX_reg[5]/NET0131 ,
		\EAX_reg[6]/NET0131 ,
		_w1743_,
		_w1744_
	);
	LUT4 #(
		.INIT('h8000)
	) name1292 (
		\EAX_reg[7]/NET0131 ,
		\EAX_reg[8]/NET0131 ,
		\EAX_reg[9]/NET0131 ,
		_w1744_,
		_w1745_
	);
	LUT2 #(
		.INIT('h8)
	) name1293 (
		\EAX_reg[10]/NET0131 ,
		_w1745_,
		_w1746_
	);
	LUT3 #(
		.INIT('h80)
	) name1294 (
		\EAX_reg[10]/NET0131 ,
		\EAX_reg[11]/NET0131 ,
		_w1745_,
		_w1747_
	);
	LUT4 #(
		.INIT('h8000)
	) name1295 (
		\EAX_reg[10]/NET0131 ,
		\EAX_reg[11]/NET0131 ,
		\EAX_reg[12]/NET0131 ,
		_w1745_,
		_w1748_
	);
	LUT2 #(
		.INIT('h8)
	) name1296 (
		\EAX_reg[13]/NET0131 ,
		_w1748_,
		_w1749_
	);
	LUT3 #(
		.INIT('h80)
	) name1297 (
		\EAX_reg[13]/NET0131 ,
		\EAX_reg[14]/NET0131 ,
		_w1748_,
		_w1750_
	);
	LUT4 #(
		.INIT('h8000)
	) name1298 (
		\EAX_reg[13]/NET0131 ,
		\EAX_reg[14]/NET0131 ,
		\EAX_reg[15]/NET0131 ,
		_w1748_,
		_w1751_
	);
	LUT2 #(
		.INIT('h8)
	) name1299 (
		\EAX_reg[16]/NET0131 ,
		_w1751_,
		_w1752_
	);
	LUT3 #(
		.INIT('h80)
	) name1300 (
		\EAX_reg[16]/NET0131 ,
		\EAX_reg[17]/NET0131 ,
		_w1751_,
		_w1753_
	);
	LUT4 #(
		.INIT('h8000)
	) name1301 (
		\EAX_reg[16]/NET0131 ,
		\EAX_reg[17]/NET0131 ,
		\EAX_reg[18]/NET0131 ,
		_w1751_,
		_w1754_
	);
	LUT2 #(
		.INIT('h8)
	) name1302 (
		\EAX_reg[20]/NET0131 ,
		\EAX_reg[21]/NET0131 ,
		_w1755_
	);
	LUT3 #(
		.INIT('h80)
	) name1303 (
		\EAX_reg[19]/NET0131 ,
		\EAX_reg[20]/NET0131 ,
		\EAX_reg[21]/NET0131 ,
		_w1756_
	);
	LUT4 #(
		.INIT('h8000)
	) name1304 (
		\EAX_reg[19]/NET0131 ,
		\EAX_reg[20]/NET0131 ,
		\EAX_reg[21]/NET0131 ,
		\EAX_reg[22]/NET0131 ,
		_w1757_
	);
	LUT2 #(
		.INIT('h8)
	) name1305 (
		\EAX_reg[23]/NET0131 ,
		\EAX_reg[24]/NET0131 ,
		_w1758_
	);
	LUT3 #(
		.INIT('h80)
	) name1306 (
		_w1754_,
		_w1757_,
		_w1758_,
		_w1759_
	);
	LUT4 #(
		.INIT('h8000)
	) name1307 (
		\EAX_reg[25]/NET0131 ,
		_w1754_,
		_w1757_,
		_w1758_,
		_w1760_
	);
	LUT4 #(
		.INIT('h0b03)
	) name1308 (
		\EAX_reg[26]/NET0131 ,
		_w1741_,
		_w1742_,
		_w1760_,
		_w1761_
	);
	LUT3 #(
		.INIT('h40)
	) name1309 (
		\EAX_reg[27]/NET0131 ,
		_w518_,
		_w617_,
		_w1762_
	);
	LUT4 #(
		.INIT('h88a8)
	) name1310 (
		\EAX_reg[27]/NET0131 ,
		READY_n_pad,
		_w563_,
		_w565_,
		_w1763_
	);
	LUT4 #(
		.INIT('h2202)
	) name1311 (
		\Datai[27]_pad ,
		READY_n_pad,
		_w563_,
		_w565_,
		_w1764_
	);
	LUT2 #(
		.INIT('h1)
	) name1312 (
		_w1763_,
		_w1764_,
		_w1765_
	);
	LUT3 #(
		.INIT('h08)
	) name1313 (
		_w494_,
		_w586_,
		_w1765_,
		_w1766_
	);
	LUT4 #(
		.INIT('h135f)
	) name1314 (
		\InstQueue_reg[13][7]/NET0131 ,
		\InstQueue_reg[4][7]/NET0131 ,
		_w471_,
		_w473_,
		_w1767_
	);
	LUT4 #(
		.INIT('h153f)
	) name1315 (
		\InstQueue_reg[11][7]/NET0131 ,
		\InstQueue_reg[7][7]/NET0131 ,
		_w468_,
		_w463_,
		_w1768_
	);
	LUT4 #(
		.INIT('h135f)
	) name1316 (
		\InstQueue_reg[1][7]/NET0131 ,
		\InstQueue_reg[9][7]/NET0131 ,
		_w476_,
		_w453_,
		_w1769_
	);
	LUT4 #(
		.INIT('h153f)
	) name1317 (
		\InstQueue_reg[2][7]/NET0131 ,
		\InstQueue_reg[6][7]/NET0131 ,
		_w460_,
		_w455_,
		_w1770_
	);
	LUT4 #(
		.INIT('h8000)
	) name1318 (
		_w1769_,
		_w1770_,
		_w1767_,
		_w1768_,
		_w1771_
	);
	LUT4 #(
		.INIT('h135f)
	) name1319 (
		\InstQueue_reg[5][7]/NET0131 ,
		\InstQueue_reg[8][7]/NET0131 ,
		_w474_,
		_w457_,
		_w1772_
	);
	LUT4 #(
		.INIT('h153f)
	) name1320 (
		\InstQueue_reg[12][7]/NET0131 ,
		\InstQueue_reg[15][7]/NET0131 ,
		_w477_,
		_w467_,
		_w1773_
	);
	LUT4 #(
		.INIT('h135f)
	) name1321 (
		\InstQueue_reg[0][7]/NET0131 ,
		\InstQueue_reg[3][7]/NET0131 ,
		_w461_,
		_w464_,
		_w1774_
	);
	LUT4 #(
		.INIT('h135f)
	) name1322 (
		\InstQueue_reg[10][7]/NET0131 ,
		\InstQueue_reg[14][7]/NET0131 ,
		_w470_,
		_w458_,
		_w1775_
	);
	LUT4 #(
		.INIT('h8000)
	) name1323 (
		_w1774_,
		_w1775_,
		_w1772_,
		_w1773_,
		_w1776_
	);
	LUT4 #(
		.INIT('h153f)
	) name1324 (
		\InstQueue_reg[14][0]/NET0131 ,
		\InstQueue_reg[6][0]/NET0131 ,
		_w474_,
		_w471_,
		_w1777_
	);
	LUT4 #(
		.INIT('h135f)
	) name1325 (
		\InstQueue_reg[11][0]/NET0131 ,
		\InstQueue_reg[3][0]/NET0131 ,
		_w470_,
		_w455_,
		_w1778_
	);
	LUT4 #(
		.INIT('h153f)
	) name1326 (
		\InstQueue_reg[10][0]/NET0131 ,
		\InstQueue_reg[7][0]/NET0131 ,
		_w460_,
		_w453_,
		_w1779_
	);
	LUT4 #(
		.INIT('h135f)
	) name1327 (
		\InstQueue_reg[1][0]/NET0131 ,
		\InstQueue_reg[2][0]/NET0131 ,
		_w461_,
		_w476_,
		_w1780_
	);
	LUT4 #(
		.INIT('h8000)
	) name1328 (
		_w1779_,
		_w1780_,
		_w1777_,
		_w1778_,
		_w1781_
	);
	LUT4 #(
		.INIT('h135f)
	) name1329 (
		\InstQueue_reg[0][0]/NET0131 ,
		\InstQueue_reg[5][0]/NET0131 ,
		_w477_,
		_w473_,
		_w1782_
	);
	LUT4 #(
		.INIT('h135f)
	) name1330 (
		\InstQueue_reg[13][0]/NET0131 ,
		\InstQueue_reg[9][0]/NET0131 ,
		_w467_,
		_w457_,
		_w1783_
	);
	LUT4 #(
		.INIT('h153f)
	) name1331 (
		\InstQueue_reg[4][0]/NET0131 ,
		\InstQueue_reg[8][0]/NET0131 ,
		_w468_,
		_w464_,
		_w1784_
	);
	LUT4 #(
		.INIT('h135f)
	) name1332 (
		\InstQueue_reg[12][0]/NET0131 ,
		\InstQueue_reg[15][0]/NET0131 ,
		_w463_,
		_w458_,
		_w1785_
	);
	LUT4 #(
		.INIT('h8000)
	) name1333 (
		_w1784_,
		_w1785_,
		_w1782_,
		_w1783_,
		_w1786_
	);
	LUT4 #(
		.INIT('h0777)
	) name1334 (
		_w1771_,
		_w1776_,
		_w1781_,
		_w1786_,
		_w1787_
	);
	LUT4 #(
		.INIT('h153f)
	) name1335 (
		\InstQueue_reg[14][1]/NET0131 ,
		\InstQueue_reg[6][1]/NET0131 ,
		_w474_,
		_w471_,
		_w1788_
	);
	LUT4 #(
		.INIT('h135f)
	) name1336 (
		\InstQueue_reg[11][1]/NET0131 ,
		\InstQueue_reg[3][1]/NET0131 ,
		_w470_,
		_w455_,
		_w1789_
	);
	LUT4 #(
		.INIT('h153f)
	) name1337 (
		\InstQueue_reg[10][1]/NET0131 ,
		\InstQueue_reg[7][1]/NET0131 ,
		_w460_,
		_w453_,
		_w1790_
	);
	LUT4 #(
		.INIT('h135f)
	) name1338 (
		\InstQueue_reg[1][1]/NET0131 ,
		\InstQueue_reg[2][1]/NET0131 ,
		_w461_,
		_w476_,
		_w1791_
	);
	LUT4 #(
		.INIT('h8000)
	) name1339 (
		_w1790_,
		_w1791_,
		_w1788_,
		_w1789_,
		_w1792_
	);
	LUT4 #(
		.INIT('h135f)
	) name1340 (
		\InstQueue_reg[0][1]/NET0131 ,
		\InstQueue_reg[5][1]/NET0131 ,
		_w477_,
		_w473_,
		_w1793_
	);
	LUT4 #(
		.INIT('h135f)
	) name1341 (
		\InstQueue_reg[13][1]/NET0131 ,
		\InstQueue_reg[9][1]/NET0131 ,
		_w467_,
		_w457_,
		_w1794_
	);
	LUT4 #(
		.INIT('h153f)
	) name1342 (
		\InstQueue_reg[4][1]/NET0131 ,
		\InstQueue_reg[8][1]/NET0131 ,
		_w468_,
		_w464_,
		_w1795_
	);
	LUT4 #(
		.INIT('h135f)
	) name1343 (
		\InstQueue_reg[12][1]/NET0131 ,
		\InstQueue_reg[15][1]/NET0131 ,
		_w463_,
		_w458_,
		_w1796_
	);
	LUT4 #(
		.INIT('h8000)
	) name1344 (
		_w1795_,
		_w1796_,
		_w1793_,
		_w1794_,
		_w1797_
	);
	LUT2 #(
		.INIT('h8)
	) name1345 (
		_w1792_,
		_w1797_,
		_w1798_
	);
	LUT4 #(
		.INIT('h135f)
	) name1346 (
		\InstQueue_reg[14][2]/NET0131 ,
		\InstQueue_reg[5][2]/NET0131 ,
		_w471_,
		_w473_,
		_w1799_
	);
	LUT4 #(
		.INIT('h135f)
	) name1347 (
		\InstQueue_reg[0][2]/NET0131 ,
		\InstQueue_reg[2][2]/NET0131 ,
		_w477_,
		_w476_,
		_w1800_
	);
	LUT4 #(
		.INIT('h135f)
	) name1348 (
		\InstQueue_reg[10][2]/NET0131 ,
		\InstQueue_reg[13][2]/NET0131 ,
		_w453_,
		_w467_,
		_w1801_
	);
	LUT4 #(
		.INIT('h135f)
	) name1349 (
		\InstQueue_reg[7][2]/NET0131 ,
		\InstQueue_reg[9][2]/NET0131 ,
		_w460_,
		_w457_,
		_w1802_
	);
	LUT4 #(
		.INIT('h8000)
	) name1350 (
		_w1801_,
		_w1802_,
		_w1799_,
		_w1800_,
		_w1803_
	);
	LUT4 #(
		.INIT('h135f)
	) name1351 (
		\InstQueue_reg[6][2]/NET0131 ,
		\InstQueue_reg[8][2]/NET0131 ,
		_w474_,
		_w468_,
		_w1804_
	);
	LUT4 #(
		.INIT('h153f)
	) name1352 (
		\InstQueue_reg[3][2]/NET0131 ,
		\InstQueue_reg[4][2]/NET0131 ,
		_w464_,
		_w455_,
		_w1805_
	);
	LUT4 #(
		.INIT('h153f)
	) name1353 (
		\InstQueue_reg[12][2]/NET0131 ,
		\InstQueue_reg[1][2]/NET0131 ,
		_w461_,
		_w463_,
		_w1806_
	);
	LUT4 #(
		.INIT('h135f)
	) name1354 (
		\InstQueue_reg[11][2]/NET0131 ,
		\InstQueue_reg[15][2]/NET0131 ,
		_w470_,
		_w458_,
		_w1807_
	);
	LUT4 #(
		.INIT('h8000)
	) name1355 (
		_w1806_,
		_w1807_,
		_w1804_,
		_w1805_,
		_w1808_
	);
	LUT2 #(
		.INIT('h8)
	) name1356 (
		_w1803_,
		_w1808_,
		_w1809_
	);
	LUT4 #(
		.INIT('h153f)
	) name1357 (
		\InstQueue_reg[14][3]/NET0131 ,
		\InstQueue_reg[6][3]/NET0131 ,
		_w474_,
		_w471_,
		_w1810_
	);
	LUT4 #(
		.INIT('h135f)
	) name1358 (
		\InstQueue_reg[11][3]/NET0131 ,
		\InstQueue_reg[3][3]/NET0131 ,
		_w470_,
		_w455_,
		_w1811_
	);
	LUT4 #(
		.INIT('h153f)
	) name1359 (
		\InstQueue_reg[10][3]/NET0131 ,
		\InstQueue_reg[7][3]/NET0131 ,
		_w460_,
		_w453_,
		_w1812_
	);
	LUT4 #(
		.INIT('h135f)
	) name1360 (
		\InstQueue_reg[1][3]/NET0131 ,
		\InstQueue_reg[2][3]/NET0131 ,
		_w461_,
		_w476_,
		_w1813_
	);
	LUT4 #(
		.INIT('h8000)
	) name1361 (
		_w1812_,
		_w1813_,
		_w1810_,
		_w1811_,
		_w1814_
	);
	LUT4 #(
		.INIT('h135f)
	) name1362 (
		\InstQueue_reg[0][3]/NET0131 ,
		\InstQueue_reg[5][3]/NET0131 ,
		_w477_,
		_w473_,
		_w1815_
	);
	LUT4 #(
		.INIT('h135f)
	) name1363 (
		\InstQueue_reg[13][3]/NET0131 ,
		\InstQueue_reg[9][3]/NET0131 ,
		_w467_,
		_w457_,
		_w1816_
	);
	LUT4 #(
		.INIT('h153f)
	) name1364 (
		\InstQueue_reg[4][3]/NET0131 ,
		\InstQueue_reg[8][3]/NET0131 ,
		_w468_,
		_w464_,
		_w1817_
	);
	LUT4 #(
		.INIT('h135f)
	) name1365 (
		\InstQueue_reg[12][3]/NET0131 ,
		\InstQueue_reg[15][3]/NET0131 ,
		_w463_,
		_w458_,
		_w1818_
	);
	LUT4 #(
		.INIT('h8000)
	) name1366 (
		_w1817_,
		_w1818_,
		_w1815_,
		_w1816_,
		_w1819_
	);
	LUT2 #(
		.INIT('h8)
	) name1367 (
		_w1814_,
		_w1819_,
		_w1820_
	);
	LUT4 #(
		.INIT('h0002)
	) name1368 (
		_w1787_,
		_w1798_,
		_w1809_,
		_w1820_,
		_w1821_
	);
	LUT4 #(
		.INIT('h135f)
	) name1369 (
		\InstQueue_reg[14][4]/NET0131 ,
		\InstQueue_reg[5][4]/NET0131 ,
		_w471_,
		_w473_,
		_w1822_
	);
	LUT4 #(
		.INIT('h135f)
	) name1370 (
		\InstQueue_reg[0][4]/NET0131 ,
		\InstQueue_reg[2][4]/NET0131 ,
		_w477_,
		_w476_,
		_w1823_
	);
	LUT4 #(
		.INIT('h135f)
	) name1371 (
		\InstQueue_reg[10][4]/NET0131 ,
		\InstQueue_reg[13][4]/NET0131 ,
		_w453_,
		_w467_,
		_w1824_
	);
	LUT4 #(
		.INIT('h135f)
	) name1372 (
		\InstQueue_reg[7][4]/NET0131 ,
		\InstQueue_reg[9][4]/NET0131 ,
		_w460_,
		_w457_,
		_w1825_
	);
	LUT4 #(
		.INIT('h8000)
	) name1373 (
		_w1824_,
		_w1825_,
		_w1822_,
		_w1823_,
		_w1826_
	);
	LUT4 #(
		.INIT('h135f)
	) name1374 (
		\InstQueue_reg[6][4]/NET0131 ,
		\InstQueue_reg[8][4]/NET0131 ,
		_w474_,
		_w468_,
		_w1827_
	);
	LUT4 #(
		.INIT('h153f)
	) name1375 (
		\InstQueue_reg[3][4]/NET0131 ,
		\InstQueue_reg[4][4]/NET0131 ,
		_w464_,
		_w455_,
		_w1828_
	);
	LUT4 #(
		.INIT('h153f)
	) name1376 (
		\InstQueue_reg[12][4]/NET0131 ,
		\InstQueue_reg[1][4]/NET0131 ,
		_w461_,
		_w463_,
		_w1829_
	);
	LUT4 #(
		.INIT('h135f)
	) name1377 (
		\InstQueue_reg[11][4]/NET0131 ,
		\InstQueue_reg[15][4]/NET0131 ,
		_w470_,
		_w458_,
		_w1830_
	);
	LUT4 #(
		.INIT('h8000)
	) name1378 (
		_w1829_,
		_w1830_,
		_w1827_,
		_w1828_,
		_w1831_
	);
	LUT2 #(
		.INIT('h8)
	) name1379 (
		_w1826_,
		_w1831_,
		_w1832_
	);
	LUT2 #(
		.INIT('h9)
	) name1380 (
		_w1821_,
		_w1832_,
		_w1833_
	);
	LUT4 #(
		.INIT('h2202)
	) name1381 (
		\Datai[11]_pad ,
		READY_n_pad,
		_w563_,
		_w565_,
		_w1834_
	);
	LUT2 #(
		.INIT('h1)
	) name1382 (
		_w1763_,
		_w1834_,
		_w1835_
	);
	LUT2 #(
		.INIT('h2)
	) name1383 (
		_w582_,
		_w1835_,
		_w1836_
	);
	LUT4 #(
		.INIT('h0007)
	) name1384 (
		_w1740_,
		_w1833_,
		_w1836_,
		_w1766_,
		_w1837_
	);
	LUT4 #(
		.INIT('h7f00)
	) name1385 (
		\EAX_reg[26]/NET0131 ,
		_w1760_,
		_w1762_,
		_w1837_,
		_w1838_
	);
	LUT4 #(
		.INIT('h08cc)
	) name1386 (
		\EAX_reg[27]/NET0131 ,
		_w690_,
		_w1761_,
		_w1838_,
		_w1839_
	);
	LUT4 #(
		.INIT('hfc7f)
	) name1387 (
		\State2_reg[0]/NET0131 ,
		\State2_reg[1]/NET0131 ,
		\State2_reg[2]/NET0131 ,
		\State2_reg[3]/NET0131 ,
		_w1840_
	);
	LUT4 #(
		.INIT('hfc20)
	) name1388 (
		\State2_reg[0]/NET0131 ,
		\State2_reg[1]/NET0131 ,
		\State2_reg[2]/NET0131 ,
		\State2_reg[3]/NET0131 ,
		_w1841_
	);
	LUT2 #(
		.INIT('h2)
	) name1389 (
		\EAX_reg[27]/NET0131 ,
		_w1841_,
		_w1842_
	);
	LUT2 #(
		.INIT('he)
	) name1390 (
		_w1839_,
		_w1842_,
		_w1843_
	);
	LUT4 #(
		.INIT('h025f)
	) name1391 (
		\State2_reg[0]/NET0131 ,
		\State2_reg[1]/NET0131 ,
		\State2_reg[2]/NET0131 ,
		\State2_reg[3]/NET0131 ,
		_w1844_
	);
	LUT2 #(
		.INIT('h8)
	) name1392 (
		\InstQueueRd_Addr_reg[0]/NET0131 ,
		_w1844_,
		_w1845_
	);
	LUT3 #(
		.INIT('h72)
	) name1393 (
		\Flush_reg/NET0131 ,
		\InstAddrPointer_reg[0]/NET0131 ,
		\InstQueueRd_Addr_reg[0]/NET0131 ,
		_w1846_
	);
	LUT4 #(
		.INIT('h23af)
	) name1394 (
		\InstQueueRd_Addr_reg[0]/NET0131 ,
		_w700_,
		_w710_,
		_w1846_,
		_w1847_
	);
	LUT2 #(
		.INIT('h4)
	) name1395 (
		_w1845_,
		_w1847_,
		_w1848_
	);
	LUT4 #(
		.INIT('h10ff)
	) name1396 (
		_w641_,
		_w643_,
		_w690_,
		_w1848_,
		_w1849_
	);
	LUT4 #(
		.INIT('h2282)
	) name1397 (
		_w836_,
		_w1133_,
		_w1134_,
		_w1270_,
		_w1850_
	);
	LUT4 #(
		.INIT('hc8cc)
	) name1398 (
		_w952_,
		_w953_,
		_w1089_,
		_w1092_,
		_w1851_
	);
	LUT4 #(
		.INIT('h0045)
	) name1399 (
		_w836_,
		_w948_,
		_w1314_,
		_w1851_,
		_w1852_
	);
	LUT4 #(
		.INIT('h7774)
	) name1400 (
		\PhyAddrPointer_reg[10]/NET0131 ,
		_w674_,
		_w1852_,
		_w1850_,
		_w1853_
	);
	LUT4 #(
		.INIT('h202a)
	) name1401 (
		\PhyAddrPointer_reg[10]/NET0131 ,
		_w634_,
		_w607_,
		_w608_,
		_w1854_
	);
	LUT3 #(
		.INIT('h32)
	) name1402 (
		\InstAddrPointer_reg[10]/NET0131 ,
		_w1006_,
		_w1041_,
		_w1855_
	);
	LUT4 #(
		.INIT('h00df)
	) name1403 (
		_w1016_,
		_w1039_,
		_w1044_,
		_w1855_,
		_w1856_
	);
	LUT3 #(
		.INIT('h02)
	) name1404 (
		_w671_,
		_w1341_,
		_w1856_,
		_w1857_
	);
	LUT4 #(
		.INIT('h0f0d)
	) name1405 (
		_w671_,
		_w1341_,
		_w1854_,
		_w1856_,
		_w1858_
	);
	LUT4 #(
		.INIT('h08cc)
	) name1406 (
		_w608_,
		_w690_,
		_w1853_,
		_w1858_,
		_w1859_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name1407 (
		\PhyAddrPointer_reg[10]/NET0131 ,
		\PhyAddrPointer_reg[8]/NET0131 ,
		\PhyAddrPointer_reg[9]/NET0131 ,
		_w1386_,
		_w1860_
	);
	LUT4 #(
		.INIT('h60a0)
	) name1408 (
		\PhyAddrPointer_reg[10]/NET0131 ,
		\PhyAddrPointer_reg[9]/NET0131 ,
		_w714_,
		_w1194_,
		_w1861_
	);
	LUT4 #(
		.INIT('h3f15)
	) name1409 (
		\PhyAddrPointer_reg[10]/NET0131 ,
		\rEIP_reg[10]/NET0131 ,
		_w1080_,
		_w1215_,
		_w1862_
	);
	LUT4 #(
		.INIT('h1300)
	) name1410 (
		_w1306_,
		_w1861_,
		_w1860_,
		_w1862_,
		_w1863_
	);
	LUT2 #(
		.INIT('hb)
	) name1411 (
		_w1859_,
		_w1863_,
		_w1864_
	);
	LUT4 #(
		.INIT('h808c)
	) name1412 (
		\PhyAddrPointer_reg[7]/NET0131 ,
		_w608_,
		_w674_,
		_w1563_,
		_w1865_
	);
	LUT4 #(
		.INIT('h202a)
	) name1413 (
		\PhyAddrPointer_reg[7]/NET0131 ,
		_w634_,
		_w607_,
		_w608_,
		_w1866_
	);
	LUT4 #(
		.INIT('h007d)
	) name1414 (
		_w671_,
		_w1108_,
		_w1565_,
		_w1866_,
		_w1867_
	);
	LUT4 #(
		.INIT('h78f0)
	) name1415 (
		\PhyAddrPointer_reg[1]/NET0131 ,
		\PhyAddrPointer_reg[6]/NET0131 ,
		\PhyAddrPointer_reg[7]/NET0131 ,
		_w1191_,
		_w1868_
	);
	LUT2 #(
		.INIT('h8)
	) name1416 (
		_w1306_,
		_w1868_,
		_w1869_
	);
	LUT4 #(
		.INIT('h3f15)
	) name1417 (
		\PhyAddrPointer_reg[7]/NET0131 ,
		\rEIP_reg[7]/NET0131 ,
		_w1080_,
		_w1215_,
		_w1870_
	);
	LUT4 #(
		.INIT('hb700)
	) name1418 (
		\PhyAddrPointer_reg[7]/NET0131 ,
		_w714_,
		_w1192_,
		_w1870_,
		_w1871_
	);
	LUT2 #(
		.INIT('h4)
	) name1419 (
		_w1869_,
		_w1871_,
		_w1872_
	);
	LUT4 #(
		.INIT('h8aff)
	) name1420 (
		_w690_,
		_w1865_,
		_w1867_,
		_w1872_,
		_w1873_
	);
	LUT3 #(
		.INIT('h08)
	) name1421 (
		\PhyAddrPointer_reg[9]/NET0131 ,
		_w563_,
		_w673_,
		_w1874_
	);
	LUT3 #(
		.INIT('ha8)
	) name1422 (
		_w608_,
		_w1585_,
		_w1874_,
		_w1875_
	);
	LUT4 #(
		.INIT('h202a)
	) name1423 (
		\PhyAddrPointer_reg[9]/NET0131 ,
		_w634_,
		_w607_,
		_w608_,
		_w1876_
	);
	LUT2 #(
		.INIT('h1)
	) name1424 (
		_w1587_,
		_w1876_,
		_w1877_
	);
	LUT3 #(
		.INIT('h6c)
	) name1425 (
		\PhyAddrPointer_reg[8]/NET0131 ,
		\PhyAddrPointer_reg[9]/NET0131 ,
		_w1386_,
		_w1878_
	);
	LUT4 #(
		.INIT('h60c0)
	) name1426 (
		\PhyAddrPointer_reg[8]/NET0131 ,
		\PhyAddrPointer_reg[9]/NET0131 ,
		_w1306_,
		_w1386_,
		_w1879_
	);
	LUT4 #(
		.INIT('h3f15)
	) name1427 (
		\PhyAddrPointer_reg[9]/NET0131 ,
		\rEIP_reg[9]/NET0131 ,
		_w1080_,
		_w1215_,
		_w1880_
	);
	LUT4 #(
		.INIT('hb700)
	) name1428 (
		\PhyAddrPointer_reg[9]/NET0131 ,
		_w714_,
		_w1194_,
		_w1880_,
		_w1881_
	);
	LUT2 #(
		.INIT('h4)
	) name1429 (
		_w1879_,
		_w1881_,
		_w1882_
	);
	LUT4 #(
		.INIT('h8aff)
	) name1430 (
		_w690_,
		_w1875_,
		_w1877_,
		_w1882_,
		_w1883_
	);
	LUT3 #(
		.INIT('h08)
	) name1431 (
		\InstAddrPointer_reg[3]/NET0131 ,
		_w563_,
		_w673_,
		_w1884_
	);
	LUT4 #(
		.INIT('h40bf)
	) name1432 (
		_w785_,
		_w783_,
		_w790_,
		_w792_,
		_w1885_
	);
	LUT4 #(
		.INIT('h5401)
	) name1433 (
		_w674_,
		_w778_,
		_w821_,
		_w1885_,
		_w1886_
	);
	LUT3 #(
		.INIT('ha8)
	) name1434 (
		_w608_,
		_w1884_,
		_w1886_,
		_w1887_
	);
	LUT4 #(
		.INIT('haaa8)
	) name1435 (
		\InstAddrPointer_reg[3]/NET0131 ,
		_w655_,
		_w612_,
		_w680_,
		_w1888_
	);
	LUT4 #(
		.INIT('h40bf)
	) name1436 (
		_w785_,
		_w783_,
		_w790_,
		_w1024_,
		_w1889_
	);
	LUT3 #(
		.INIT('h0e)
	) name1437 (
		_w1028_,
		_w1031_,
		_w1889_,
		_w1890_
	);
	LUT3 #(
		.INIT('h10)
	) name1438 (
		_w1028_,
		_w1031_,
		_w1889_,
		_w1891_
	);
	LUT3 #(
		.INIT('h02)
	) name1439 (
		_w671_,
		_w1891_,
		_w1890_,
		_w1892_
	);
	LUT4 #(
		.INIT('hf078)
	) name1440 (
		\InstAddrPointer_reg[1]/NET0131 ,
		\InstAddrPointer_reg[2]/NET0131 ,
		\InstAddrPointer_reg[3]/NET0131 ,
		READY_n_pad,
		_w1893_
	);
	LUT4 #(
		.INIT('haaa9)
	) name1441 (
		\InstAddrPointer_reg[3]/NET0131 ,
		_w563_,
		_w633_,
		_w928_,
		_w1894_
	);
	LUT4 #(
		.INIT('hc800)
	) name1442 (
		_w569_,
		_w602_,
		_w604_,
		_w1894_,
		_w1895_
	);
	LUT3 #(
		.INIT('h07)
	) name1443 (
		_w588_,
		_w1893_,
		_w1895_,
		_w1896_
	);
	LUT3 #(
		.INIT('h10)
	) name1444 (
		_w1888_,
		_w1892_,
		_w1896_,
		_w1897_
	);
	LUT4 #(
		.INIT('hea00)
	) name1445 (
		_w554_,
		_w645_,
		_w646_,
		_w792_,
		_w1898_
	);
	LUT4 #(
		.INIT('h004f)
	) name1446 (
		_w616_,
		_w630_,
		_w926_,
		_w1898_,
		_w1899_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name1447 (
		_w690_,
		_w1887_,
		_w1897_,
		_w1899_,
		_w1900_
	);
	LUT4 #(
		.INIT('h153f)
	) name1448 (
		\InstAddrPointer_reg[3]/NET0131 ,
		\rEIP_reg[3]/NET0131 ,
		_w1080_,
		_w1081_,
		_w1901_
	);
	LUT2 #(
		.INIT('hb)
	) name1449 (
		_w1900_,
		_w1901_,
		_w1902_
	);
	LUT3 #(
		.INIT('h87)
	) name1450 (
		_w860_,
		_w865_,
		_w867_,
		_w1903_
	);
	LUT4 #(
		.INIT('h7447)
	) name1451 (
		\InstAddrPointer_reg[5]/NET0131 ,
		_w674_,
		_w825_,
		_w1903_,
		_w1904_
	);
	LUT2 #(
		.INIT('h2)
	) name1452 (
		_w608_,
		_w1904_,
		_w1905_
	);
	LUT2 #(
		.INIT('h2)
	) name1453 (
		\InstAddrPointer_reg[5]/NET0131 ,
		_w1295_,
		_w1906_
	);
	LUT2 #(
		.INIT('h8)
	) name1454 (
		_w635_,
		_w1019_,
		_w1907_
	);
	LUT4 #(
		.INIT('h004f)
	) name1455 (
		_w616_,
		_w630_,
		_w939_,
		_w1907_,
		_w1908_
	);
	LUT3 #(
		.INIT('h87)
	) name1456 (
		_w860_,
		_w865_,
		_w1019_,
		_w1909_
	);
	LUT3 #(
		.INIT('h82)
	) name1457 (
		_w671_,
		_w1106_,
		_w1909_,
		_w1910_
	);
	LUT3 #(
		.INIT('h0b)
	) name1458 (
		_w597_,
		_w867_,
		_w1910_,
		_w1911_
	);
	LUT4 #(
		.INIT('h1000)
	) name1459 (
		_w1906_,
		_w1905_,
		_w1908_,
		_w1911_,
		_w1912_
	);
	LUT2 #(
		.INIT('h8)
	) name1460 (
		\rEIP_reg[5]/NET0131 ,
		_w1080_,
		_w1913_
	);
	LUT4 #(
		.INIT('h153f)
	) name1461 (
		\InstAddrPointer_reg[5]/NET0131 ,
		\rEIP_reg[5]/NET0131 ,
		_w1080_,
		_w1081_,
		_w1914_
	);
	LUT3 #(
		.INIT('h2f)
	) name1462 (
		_w690_,
		_w1912_,
		_w1914_,
		_w1915_
	);
	LUT2 #(
		.INIT('h2)
	) name1463 (
		\EAX_reg[30]/NET0131 ,
		_w1841_,
		_w1916_
	);
	LUT2 #(
		.INIT('h8)
	) name1464 (
		\EAX_reg[26]/NET0131 ,
		\EAX_reg[27]/NET0131 ,
		_w1917_
	);
	LUT2 #(
		.INIT('h8)
	) name1465 (
		\EAX_reg[28]/NET0131 ,
		\EAX_reg[29]/NET0131 ,
		_w1918_
	);
	LUT4 #(
		.INIT('h1555)
	) name1466 (
		\EAX_reg[30]/NET0131 ,
		_w1760_,
		_w1917_,
		_w1918_,
		_w1919_
	);
	LUT3 #(
		.INIT('h80)
	) name1467 (
		\EAX_reg[28]/NET0131 ,
		\EAX_reg[29]/NET0131 ,
		\EAX_reg[30]/NET0131 ,
		_w1920_
	);
	LUT3 #(
		.INIT('h80)
	) name1468 (
		_w1760_,
		_w1917_,
		_w1920_,
		_w1921_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name1469 (
		_w1741_,
		_w1760_,
		_w1917_,
		_w1920_,
		_w1922_
	);
	LUT3 #(
		.INIT('ha8)
	) name1470 (
		\EAX_reg[30]/NET0131 ,
		_w653_,
		_w1742_,
		_w1923_
	);
	LUT4 #(
		.INIT('h153f)
	) name1471 (
		\InstQueue_reg[5][5]/NET0131 ,
		\InstQueue_reg[8][5]/NET0131 ,
		_w468_,
		_w473_,
		_w1924_
	);
	LUT4 #(
		.INIT('h135f)
	) name1472 (
		\InstQueue_reg[0][5]/NET0131 ,
		\InstQueue_reg[15][5]/NET0131 ,
		_w477_,
		_w458_,
		_w1925_
	);
	LUT4 #(
		.INIT('h153f)
	) name1473 (
		\InstQueue_reg[13][5]/NET0131 ,
		\InstQueue_reg[2][5]/NET0131 ,
		_w476_,
		_w467_,
		_w1926_
	);
	LUT4 #(
		.INIT('h135f)
	) name1474 (
		\InstQueue_reg[1][5]/NET0131 ,
		\InstQueue_reg[7][5]/NET0131 ,
		_w461_,
		_w460_,
		_w1927_
	);
	LUT4 #(
		.INIT('h8000)
	) name1475 (
		_w1926_,
		_w1927_,
		_w1924_,
		_w1925_,
		_w1928_
	);
	LUT4 #(
		.INIT('h153f)
	) name1476 (
		\InstQueue_reg[14][5]/NET0131 ,
		\InstQueue_reg[6][5]/NET0131 ,
		_w474_,
		_w471_,
		_w1929_
	);
	LUT4 #(
		.INIT('h135f)
	) name1477 (
		\InstQueue_reg[10][5]/NET0131 ,
		\InstQueue_reg[3][5]/NET0131 ,
		_w453_,
		_w455_,
		_w1930_
	);
	LUT4 #(
		.INIT('h135f)
	) name1478 (
		\InstQueue_reg[4][5]/NET0131 ,
		\InstQueue_reg[9][5]/NET0131 ,
		_w464_,
		_w457_,
		_w1931_
	);
	LUT4 #(
		.INIT('h135f)
	) name1479 (
		\InstQueue_reg[11][5]/NET0131 ,
		\InstQueue_reg[12][5]/NET0131 ,
		_w470_,
		_w463_,
		_w1932_
	);
	LUT4 #(
		.INIT('h8000)
	) name1480 (
		_w1931_,
		_w1932_,
		_w1929_,
		_w1930_,
		_w1933_
	);
	LUT2 #(
		.INIT('h8)
	) name1481 (
		_w1928_,
		_w1933_,
		_w1934_
	);
	LUT4 #(
		.INIT('h153f)
	) name1482 (
		\InstQueue_reg[5][6]/NET0131 ,
		\InstQueue_reg[8][6]/NET0131 ,
		_w468_,
		_w473_,
		_w1935_
	);
	LUT4 #(
		.INIT('h135f)
	) name1483 (
		\InstQueue_reg[0][6]/NET0131 ,
		\InstQueue_reg[15][6]/NET0131 ,
		_w477_,
		_w458_,
		_w1936_
	);
	LUT4 #(
		.INIT('h153f)
	) name1484 (
		\InstQueue_reg[13][6]/NET0131 ,
		\InstQueue_reg[2][6]/NET0131 ,
		_w476_,
		_w467_,
		_w1937_
	);
	LUT4 #(
		.INIT('h135f)
	) name1485 (
		\InstQueue_reg[1][6]/NET0131 ,
		\InstQueue_reg[7][6]/NET0131 ,
		_w461_,
		_w460_,
		_w1938_
	);
	LUT4 #(
		.INIT('h8000)
	) name1486 (
		_w1937_,
		_w1938_,
		_w1935_,
		_w1936_,
		_w1939_
	);
	LUT4 #(
		.INIT('h153f)
	) name1487 (
		\InstQueue_reg[14][6]/NET0131 ,
		\InstQueue_reg[6][6]/NET0131 ,
		_w474_,
		_w471_,
		_w1940_
	);
	LUT4 #(
		.INIT('h135f)
	) name1488 (
		\InstQueue_reg[10][6]/NET0131 ,
		\InstQueue_reg[3][6]/NET0131 ,
		_w453_,
		_w455_,
		_w1941_
	);
	LUT4 #(
		.INIT('h135f)
	) name1489 (
		\InstQueue_reg[4][6]/NET0131 ,
		\InstQueue_reg[9][6]/NET0131 ,
		_w464_,
		_w457_,
		_w1942_
	);
	LUT4 #(
		.INIT('h135f)
	) name1490 (
		\InstQueue_reg[11][6]/NET0131 ,
		\InstQueue_reg[12][6]/NET0131 ,
		_w470_,
		_w463_,
		_w1943_
	);
	LUT4 #(
		.INIT('h8000)
	) name1491 (
		_w1942_,
		_w1943_,
		_w1940_,
		_w1941_,
		_w1944_
	);
	LUT2 #(
		.INIT('h8)
	) name1492 (
		_w1939_,
		_w1944_,
		_w1945_
	);
	LUT4 #(
		.INIT('h0002)
	) name1493 (
		_w1821_,
		_w1832_,
		_w1934_,
		_w1945_,
		_w1946_
	);
	LUT4 #(
		.INIT('h135f)
	) name1494 (
		\InstQueue_reg[14][7]/NET0131 ,
		\InstQueue_reg[5][7]/NET0131 ,
		_w471_,
		_w473_,
		_w1947_
	);
	LUT4 #(
		.INIT('h135f)
	) name1495 (
		\InstQueue_reg[0][7]/NET0131 ,
		\InstQueue_reg[2][7]/NET0131 ,
		_w477_,
		_w476_,
		_w1948_
	);
	LUT4 #(
		.INIT('h135f)
	) name1496 (
		\InstQueue_reg[10][7]/NET0131 ,
		\InstQueue_reg[13][7]/NET0131 ,
		_w453_,
		_w467_,
		_w1949_
	);
	LUT4 #(
		.INIT('h135f)
	) name1497 (
		\InstQueue_reg[7][7]/NET0131 ,
		\InstQueue_reg[9][7]/NET0131 ,
		_w460_,
		_w457_,
		_w1950_
	);
	LUT4 #(
		.INIT('h8000)
	) name1498 (
		_w1949_,
		_w1950_,
		_w1947_,
		_w1948_,
		_w1951_
	);
	LUT4 #(
		.INIT('h135f)
	) name1499 (
		\InstQueue_reg[6][7]/NET0131 ,
		\InstQueue_reg[8][7]/NET0131 ,
		_w474_,
		_w468_,
		_w1952_
	);
	LUT4 #(
		.INIT('h153f)
	) name1500 (
		\InstQueue_reg[3][7]/NET0131 ,
		\InstQueue_reg[4][7]/NET0131 ,
		_w464_,
		_w455_,
		_w1953_
	);
	LUT4 #(
		.INIT('h153f)
	) name1501 (
		\InstQueue_reg[12][7]/NET0131 ,
		\InstQueue_reg[1][7]/NET0131 ,
		_w461_,
		_w463_,
		_w1954_
	);
	LUT4 #(
		.INIT('h135f)
	) name1502 (
		\InstQueue_reg[11][7]/NET0131 ,
		\InstQueue_reg[15][7]/NET0131 ,
		_w470_,
		_w458_,
		_w1955_
	);
	LUT4 #(
		.INIT('h8000)
	) name1503 (
		_w1954_,
		_w1955_,
		_w1952_,
		_w1953_,
		_w1956_
	);
	LUT2 #(
		.INIT('h8)
	) name1504 (
		_w1951_,
		_w1956_,
		_w1957_
	);
	LUT3 #(
		.INIT('h82)
	) name1505 (
		_w1740_,
		_w1946_,
		_w1957_,
		_w1958_
	);
	LUT2 #(
		.INIT('h8)
	) name1506 (
		\Datai[14]_pad ,
		_w582_,
		_w1959_
	);
	LUT3 #(
		.INIT('h80)
	) name1507 (
		\Datai[30]_pad ,
		_w494_,
		_w586_,
		_w1960_
	);
	LUT3 #(
		.INIT('ha8)
	) name1508 (
		_w652_,
		_w1959_,
		_w1960_,
		_w1961_
	);
	LUT2 #(
		.INIT('h1)
	) name1509 (
		_w1958_,
		_w1961_,
		_w1962_
	);
	LUT4 #(
		.INIT('h4500)
	) name1510 (
		_w1923_,
		_w1919_,
		_w1922_,
		_w1962_,
		_w1963_
	);
	LUT3 #(
		.INIT('hce)
	) name1511 (
		_w690_,
		_w1916_,
		_w1963_,
		_w1964_
	);
	LUT4 #(
		.INIT('h8000)
	) name1512 (
		\Datai[31]_pad ,
		_w494_,
		_w586_,
		_w652_,
		_w1965_
	);
	LUT4 #(
		.INIT('h00f7)
	) name1513 (
		_w1740_,
		_w1946_,
		_w1957_,
		_w1965_,
		_w1966_
	);
	LUT4 #(
		.INIT('h5700)
	) name1514 (
		\EAX_reg[31]/NET0131 ,
		_w653_,
		_w1742_,
		_w1966_,
		_w1967_
	);
	LUT4 #(
		.INIT('hb700)
	) name1515 (
		\EAX_reg[31]/NET0131 ,
		_w1741_,
		_w1921_,
		_w1967_,
		_w1968_
	);
	LUT2 #(
		.INIT('h2)
	) name1516 (
		\EAX_reg[31]/NET0131 ,
		_w1841_,
		_w1969_
	);
	LUT3 #(
		.INIT('hf2)
	) name1517 (
		_w690_,
		_w1968_,
		_w1969_,
		_w1970_
	);
	LUT4 #(
		.INIT('h8000)
	) name1518 (
		\EBX_reg[0]/NET0131 ,
		\EBX_reg[1]/NET0131 ,
		\EBX_reg[2]/NET0131 ,
		\EBX_reg[3]/NET0131 ,
		_w1971_
	);
	LUT4 #(
		.INIT('h8000)
	) name1519 (
		\EBX_reg[4]/NET0131 ,
		\EBX_reg[5]/NET0131 ,
		\EBX_reg[6]/NET0131 ,
		_w1971_,
		_w1972_
	);
	LUT4 #(
		.INIT('h8000)
	) name1520 (
		\EBX_reg[7]/NET0131 ,
		\EBX_reg[8]/NET0131 ,
		\EBX_reg[9]/NET0131 ,
		_w1972_,
		_w1973_
	);
	LUT2 #(
		.INIT('h8)
	) name1521 (
		\EBX_reg[10]/NET0131 ,
		_w1973_,
		_w1974_
	);
	LUT3 #(
		.INIT('h80)
	) name1522 (
		\EBX_reg[10]/NET0131 ,
		\EBX_reg[11]/NET0131 ,
		_w1973_,
		_w1975_
	);
	LUT4 #(
		.INIT('h8000)
	) name1523 (
		\EBX_reg[10]/NET0131 ,
		\EBX_reg[11]/NET0131 ,
		\EBX_reg[12]/NET0131 ,
		_w1973_,
		_w1976_
	);
	LUT2 #(
		.INIT('h8)
	) name1524 (
		\EBX_reg[13]/NET0131 ,
		_w1976_,
		_w1977_
	);
	LUT3 #(
		.INIT('h80)
	) name1525 (
		\EBX_reg[13]/NET0131 ,
		\EBX_reg[14]/NET0131 ,
		_w1976_,
		_w1978_
	);
	LUT4 #(
		.INIT('h8000)
	) name1526 (
		\EBX_reg[13]/NET0131 ,
		\EBX_reg[14]/NET0131 ,
		\EBX_reg[15]/NET0131 ,
		_w1976_,
		_w1979_
	);
	LUT2 #(
		.INIT('h8)
	) name1527 (
		\EBX_reg[16]/NET0131 ,
		_w1979_,
		_w1980_
	);
	LUT3 #(
		.INIT('h80)
	) name1528 (
		\EBX_reg[16]/NET0131 ,
		\EBX_reg[17]/NET0131 ,
		_w1979_,
		_w1981_
	);
	LUT4 #(
		.INIT('h8000)
	) name1529 (
		\EBX_reg[16]/NET0131 ,
		\EBX_reg[17]/NET0131 ,
		\EBX_reg[18]/NET0131 ,
		_w1979_,
		_w1982_
	);
	LUT4 #(
		.INIT('h8000)
	) name1530 (
		\EBX_reg[20]/NET0131 ,
		\EBX_reg[21]/NET0131 ,
		\EBX_reg[22]/NET0131 ,
		\EBX_reg[23]/NET0131 ,
		_w1983_
	);
	LUT3 #(
		.INIT('h80)
	) name1531 (
		\EBX_reg[19]/NET0131 ,
		_w1982_,
		_w1983_,
		_w1984_
	);
	LUT2 #(
		.INIT('h8)
	) name1532 (
		\EBX_reg[24]/NET0131 ,
		\EBX_reg[25]/NET0131 ,
		_w1985_
	);
	LUT4 #(
		.INIT('h8000)
	) name1533 (
		\EBX_reg[19]/NET0131 ,
		_w1982_,
		_w1983_,
		_w1985_,
		_w1986_
	);
	LUT2 #(
		.INIT('h8)
	) name1534 (
		\EBX_reg[26]/NET0131 ,
		\EBX_reg[27]/NET0131 ,
		_w1987_
	);
	LUT3 #(
		.INIT('h80)
	) name1535 (
		\EBX_reg[28]/NET0131 ,
		\EBX_reg[29]/NET0131 ,
		\EBX_reg[30]/NET0131 ,
		_w1988_
	);
	LUT3 #(
		.INIT('h80)
	) name1536 (
		_w1986_,
		_w1987_,
		_w1988_,
		_w1989_
	);
	LUT3 #(
		.INIT('h80)
	) name1537 (
		_w569_,
		_w602_,
		_w634_,
		_w1990_
	);
	LUT4 #(
		.INIT('h7000)
	) name1538 (
		_w569_,
		_w602_,
		_w617_,
		_w621_,
		_w1991_
	);
	LUT2 #(
		.INIT('h1)
	) name1539 (
		_w1990_,
		_w1991_,
		_w1992_
	);
	LUT3 #(
		.INIT('h02)
	) name1540 (
		\EBX_reg[31]/NET0131 ,
		_w1990_,
		_w1991_,
		_w1993_
	);
	LUT3 #(
		.INIT('h20)
	) name1541 (
		_w1946_,
		_w1957_,
		_w1990_,
		_w1994_
	);
	LUT2 #(
		.INIT('h1)
	) name1542 (
		_w1993_,
		_w1994_,
		_w1995_
	);
	LUT4 #(
		.INIT('hb700)
	) name1543 (
		\EBX_reg[31]/NET0131 ,
		_w622_,
		_w1989_,
		_w1995_,
		_w1996_
	);
	LUT2 #(
		.INIT('h2)
	) name1544 (
		\EBX_reg[31]/NET0131 ,
		_w1841_,
		_w1997_
	);
	LUT3 #(
		.INIT('hf2)
	) name1545 (
		_w690_,
		_w1996_,
		_w1997_,
		_w1998_
	);
	LUT4 #(
		.INIT('hef00)
	) name1546 (
		_w660_,
		_w662_,
		_w664_,
		_w690_,
		_w1999_
	);
	LUT4 #(
		.INIT('h0880)
	) name1547 (
		\Flush_reg/NET0131 ,
		\InstAddrPointer_reg[0]/NET0131 ,
		\InstAddrPointer_reg[1]/NET0131 ,
		\InstAddrPointer_reg[31]/NET0131 ,
		_w2000_
	);
	LUT3 #(
		.INIT('ha8)
	) name1548 (
		_w700_,
		_w701_,
		_w2000_,
		_w2001_
	);
	LUT4 #(
		.INIT('h159f)
	) name1549 (
		\InstQueueRd_Addr_reg[2]/NET0131 ,
		_w454_,
		_w710_,
		_w1844_,
		_w2002_
	);
	LUT2 #(
		.INIT('h4)
	) name1550 (
		_w2001_,
		_w2002_,
		_w2003_
	);
	LUT2 #(
		.INIT('hb)
	) name1551 (
		_w1999_,
		_w2003_,
		_w2004_
	);
	LUT4 #(
		.INIT('h808c)
	) name1552 (
		\PhyAddrPointer_reg[4]/NET0131 ,
		_w608_,
		_w674_,
		_w1713_,
		_w2005_
	);
	LUT4 #(
		.INIT('h202a)
	) name1553 (
		\PhyAddrPointer_reg[4]/NET0131 ,
		_w634_,
		_w607_,
		_w608_,
		_w2006_
	);
	LUT4 #(
		.INIT('h00d7)
	) name1554 (
		_w671_,
		_w1715_,
		_w1716_,
		_w2006_,
		_w2007_
	);
	LUT3 #(
		.INIT('h80)
	) name1555 (
		\PhyAddrPointer_reg[1]/NET0131 ,
		\PhyAddrPointer_reg[2]/NET0131 ,
		\PhyAddrPointer_reg[3]/NET0131 ,
		_w2008_
	);
	LUT4 #(
		.INIT('h8000)
	) name1556 (
		\PhyAddrPointer_reg[1]/NET0131 ,
		\PhyAddrPointer_reg[2]/NET0131 ,
		\PhyAddrPointer_reg[3]/NET0131 ,
		\PhyAddrPointer_reg[4]/NET0131 ,
		_w2009_
	);
	LUT4 #(
		.INIT('h7f80)
	) name1557 (
		\PhyAddrPointer_reg[1]/NET0131 ,
		\PhyAddrPointer_reg[2]/NET0131 ,
		\PhyAddrPointer_reg[3]/NET0131 ,
		\PhyAddrPointer_reg[4]/NET0131 ,
		_w2010_
	);
	LUT4 #(
		.INIT('hf400)
	) name1558 (
		\DataWidth_reg[1]/NET0131 ,
		_w695_,
		_w1212_,
		_w2010_,
		_w2011_
	);
	LUT2 #(
		.INIT('h2)
	) name1559 (
		\PhyAddrPointer_reg[4]/NET0131 ,
		_w1215_,
		_w2012_
	);
	LUT3 #(
		.INIT('h78)
	) name1560 (
		\PhyAddrPointer_reg[2]/NET0131 ,
		\PhyAddrPointer_reg[3]/NET0131 ,
		\PhyAddrPointer_reg[4]/NET0131 ,
		_w2013_
	);
	LUT3 #(
		.INIT('h80)
	) name1561 (
		\DataWidth_reg[1]/NET0131 ,
		_w695_,
		_w2013_,
		_w2014_
	);
	LUT4 #(
		.INIT('h0001)
	) name1562 (
		_w1720_,
		_w2014_,
		_w2012_,
		_w2011_,
		_w2015_
	);
	LUT4 #(
		.INIT('h8aff)
	) name1563 (
		_w690_,
		_w2005_,
		_w2007_,
		_w2015_,
		_w2016_
	);
	LUT2 #(
		.INIT('h4)
	) name1564 (
		_w597_,
		_w777_,
		_w2017_
	);
	LUT3 #(
		.INIT('h8a)
	) name1565 (
		\InstAddrPointer_reg[2]/NET0131 ,
		_w669_,
		_w1704_,
		_w2018_
	);
	LUT4 #(
		.INIT('h40bf)
	) name1566 (
		_w770_,
		_w768_,
		_w775_,
		_w777_,
		_w2019_
	);
	LUT4 #(
		.INIT('h718e)
	) name1567 (
		\InstAddrPointer_reg[1]/NET0131 ,
		_w806_,
		_w819_,
		_w2019_,
		_w2020_
	);
	LUT4 #(
		.INIT('h808c)
	) name1568 (
		\InstAddrPointer_reg[2]/NET0131 ,
		_w608_,
		_w674_,
		_w2020_,
		_w2021_
	);
	LUT4 #(
		.INIT('haaa9)
	) name1569 (
		\InstAddrPointer_reg[2]/NET0131 ,
		_w563_,
		_w633_,
		_w924_,
		_w2022_
	);
	LUT4 #(
		.INIT('hc800)
	) name1570 (
		_w569_,
		_w602_,
		_w604_,
		_w2022_,
		_w2023_
	);
	LUT4 #(
		.INIT('h40bf)
	) name1571 (
		_w770_,
		_w768_,
		_w775_,
		_w929_,
		_w2024_
	);
	LUT4 #(
		.INIT('h00d4)
	) name1572 (
		_w806_,
		_w932_,
		_w1030_,
		_w2024_,
		_w2025_
	);
	LUT4 #(
		.INIT('h2b00)
	) name1573 (
		_w806_,
		_w932_,
		_w1030_,
		_w2024_,
		_w2026_
	);
	LUT4 #(
		.INIT('h0008)
	) name1574 (
		_w634_,
		_w607_,
		_w2026_,
		_w2025_,
		_w2027_
	);
	LUT3 #(
		.INIT('h01)
	) name1575 (
		_w2023_,
		_w2021_,
		_w2027_,
		_w2028_
	);
	LUT4 #(
		.INIT('h4f00)
	) name1576 (
		_w616_,
		_w630_,
		_w929_,
		_w2028_,
		_w2029_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name1577 (
		_w690_,
		_w2018_,
		_w2017_,
		_w2029_,
		_w2030_
	);
	LUT2 #(
		.INIT('h8)
	) name1578 (
		\rEIP_reg[2]/NET0131 ,
		_w1080_,
		_w2031_
	);
	LUT4 #(
		.INIT('h153f)
	) name1579 (
		\InstAddrPointer_reg[2]/NET0131 ,
		\rEIP_reg[2]/NET0131 ,
		_w1080_,
		_w1081_,
		_w2032_
	);
	LUT2 #(
		.INIT('hb)
	) name1580 (
		_w2030_,
		_w2032_,
		_w2033_
	);
	LUT3 #(
		.INIT('h8a)
	) name1581 (
		\InstAddrPointer_reg[0]/NET0131 ,
		_w634_,
		_w607_,
		_w2034_
	);
	LUT2 #(
		.INIT('h8)
	) name1582 (
		_w615_,
		_w2034_,
		_w2035_
	);
	LUT4 #(
		.INIT('h00ef)
	) name1583 (
		\InstAddrPointer_reg[0]/NET0131 ,
		_w616_,
		_w630_,
		_w2035_,
		_w2036_
	);
	LUT3 #(
		.INIT('ha9)
	) name1584 (
		\InstAddrPointer_reg[0]/NET0131 ,
		_w563_,
		_w633_,
		_w2037_
	);
	LUT4 #(
		.INIT('hc800)
	) name1585 (
		_w569_,
		_w602_,
		_w604_,
		_w2037_,
		_w2038_
	);
	LUT3 #(
		.INIT('h6a)
	) name1586 (
		\InstAddrPointer_reg[0]/NET0131 ,
		_w812_,
		_w817_,
		_w2039_
	);
	LUT2 #(
		.INIT('h1)
	) name1587 (
		_w674_,
		_w2039_,
		_w2040_
	);
	LUT3 #(
		.INIT('h56)
	) name1588 (
		\InstAddrPointer_reg[0]/NET0131 ,
		_w674_,
		_w818_,
		_w2041_
	);
	LUT2 #(
		.INIT('h2)
	) name1589 (
		_w608_,
		_w2041_,
		_w2042_
	);
	LUT3 #(
		.INIT('h80)
	) name1590 (
		_w634_,
		_w607_,
		_w2039_,
		_w2043_
	);
	LUT3 #(
		.INIT('h01)
	) name1591 (
		_w2042_,
		_w2043_,
		_w2038_,
		_w2044_
	);
	LUT2 #(
		.INIT('h8)
	) name1592 (
		\rEIP_reg[0]/NET0131 ,
		_w1080_,
		_w2045_
	);
	LUT4 #(
		.INIT('h153f)
	) name1593 (
		\InstAddrPointer_reg[0]/NET0131 ,
		\rEIP_reg[0]/NET0131 ,
		_w1080_,
		_w1081_,
		_w2046_
	);
	LUT4 #(
		.INIT('h8aff)
	) name1594 (
		_w690_,
		_w2036_,
		_w2044_,
		_w2046_,
		_w2047_
	);
	LUT3 #(
		.INIT('h8a)
	) name1595 (
		\InstAddrPointer_reg[1]/NET0131 ,
		_w679_,
		_w1165_,
		_w2048_
	);
	LUT4 #(
		.INIT('hef00)
	) name1596 (
		_w635_,
		_w616_,
		_w630_,
		_w932_,
		_w2049_
	);
	LUT3 #(
		.INIT('h87)
	) name1597 (
		_w800_,
		_w805_,
		_w932_,
		_w2050_
	);
	LUT3 #(
		.INIT('h6a)
	) name1598 (
		\InstAddrPointer_reg[1]/NET0131 ,
		_w800_,
		_w805_,
		_w2051_
	);
	LUT4 #(
		.INIT('h4051)
	) name1599 (
		_w836_,
		_w934_,
		_w2051_,
		_w2050_,
		_w2052_
	);
	LUT3 #(
		.INIT('h28)
	) name1600 (
		_w836_,
		_w819_,
		_w2051_,
		_w2053_
	);
	LUT4 #(
		.INIT('h2220)
	) name1601 (
		_w608_,
		_w674_,
		_w2052_,
		_w2053_,
		_w2054_
	);
	LUT3 #(
		.INIT('hd8)
	) name1602 (
		_w1030_,
		_w2051_,
		_w2050_,
		_w2055_
	);
	LUT3 #(
		.INIT('h80)
	) name1603 (
		_w634_,
		_w607_,
		_w2055_,
		_w2056_
	);
	LUT2 #(
		.INIT('h1)
	) name1604 (
		_w2054_,
		_w2056_,
		_w2057_
	);
	LUT3 #(
		.INIT('he0)
	) name1605 (
		\InstAddrPointer_reg[1]/NET0131 ,
		_w597_,
		_w2057_,
		_w2058_
	);
	LUT2 #(
		.INIT('h4)
	) name1606 (
		_w2049_,
		_w2058_,
		_w2059_
	);
	LUT2 #(
		.INIT('h8)
	) name1607 (
		\rEIP_reg[1]/NET0131 ,
		_w1080_,
		_w2060_
	);
	LUT4 #(
		.INIT('h153f)
	) name1608 (
		\InstAddrPointer_reg[1]/NET0131 ,
		\rEIP_reg[1]/NET0131 ,
		_w1080_,
		_w1081_,
		_w2061_
	);
	LUT4 #(
		.INIT('h8aff)
	) name1609 (
		_w690_,
		_w2048_,
		_w2059_,
		_w2061_,
		_w2062_
	);
	LUT4 #(
		.INIT('hfe00)
	) name1610 (
		_w651_,
		_w649_,
		_w657_,
		_w690_,
		_w2063_
	);
	LUT2 #(
		.INIT('h4)
	) name1611 (
		\Flush_reg/NET0131 ,
		\InstQueueRd_Addr_reg[1]/NET0131 ,
		_w2064_
	);
	LUT4 #(
		.INIT('h8008)
	) name1612 (
		\Flush_reg/NET0131 ,
		\InstAddrPointer_reg[0]/NET0131 ,
		\InstAddrPointer_reg[1]/NET0131 ,
		\InstAddrPointer_reg[31]/NET0131 ,
		_w2065_
	);
	LUT3 #(
		.INIT('ha8)
	) name1613 (
		_w700_,
		_w2064_,
		_w2065_,
		_w2066_
	);
	LUT4 #(
		.INIT('h139f)
	) name1614 (
		\InstQueueRd_Addr_reg[0]/NET0131 ,
		\InstQueueRd_Addr_reg[1]/NET0131 ,
		_w710_,
		_w1844_,
		_w2067_
	);
	LUT2 #(
		.INIT('h4)
	) name1615 (
		_w2066_,
		_w2067_,
		_w2068_
	);
	LUT2 #(
		.INIT('hb)
	) name1616 (
		_w2063_,
		_w2068_,
		_w2069_
	);
	LUT2 #(
		.INIT('h2)
	) name1617 (
		\EAX_reg[26]/NET0131 ,
		_w1841_,
		_w2070_
	);
	LUT3 #(
		.INIT('h48)
	) name1618 (
		\EAX_reg[26]/NET0131 ,
		_w1741_,
		_w1760_,
		_w2071_
	);
	LUT4 #(
		.INIT('h88a8)
	) name1619 (
		\EAX_reg[26]/NET0131 ,
		READY_n_pad,
		_w563_,
		_w565_,
		_w2072_
	);
	LUT4 #(
		.INIT('h2202)
	) name1620 (
		\Datai[10]_pad ,
		READY_n_pad,
		_w563_,
		_w565_,
		_w2073_
	);
	LUT2 #(
		.INIT('h1)
	) name1621 (
		_w2072_,
		_w2073_,
		_w2074_
	);
	LUT2 #(
		.INIT('h2)
	) name1622 (
		_w582_,
		_w2074_,
		_w2075_
	);
	LUT4 #(
		.INIT('h02fd)
	) name1623 (
		_w1787_,
		_w1798_,
		_w1809_,
		_w1820_,
		_w2076_
	);
	LUT4 #(
		.INIT('h8000)
	) name1624 (
		_w602_,
		_w604_,
		_w634_,
		_w2076_,
		_w2077_
	);
	LUT4 #(
		.INIT('h2202)
	) name1625 (
		\Datai[26]_pad ,
		READY_n_pad,
		_w563_,
		_w565_,
		_w2078_
	);
	LUT2 #(
		.INIT('h1)
	) name1626 (
		_w2072_,
		_w2078_,
		_w2079_
	);
	LUT3 #(
		.INIT('h08)
	) name1627 (
		_w494_,
		_w586_,
		_w2079_,
		_w2080_
	);
	LUT3 #(
		.INIT('h01)
	) name1628 (
		_w2077_,
		_w2080_,
		_w2075_,
		_w2081_
	);
	LUT3 #(
		.INIT('h70)
	) name1629 (
		\EAX_reg[26]/NET0131 ,
		_w1742_,
		_w2081_,
		_w2082_
	);
	LUT4 #(
		.INIT('hecee)
	) name1630 (
		_w690_,
		_w2070_,
		_w2071_,
		_w2082_,
		_w2083_
	);
	LUT4 #(
		.INIT('hfffc)
	) name1631 (
		\State2_reg[0]/NET0131 ,
		\State2_reg[1]/NET0131 ,
		\State2_reg[2]/NET0131 ,
		\State2_reg[3]/NET0131 ,
		_w2084_
	);
	LUT4 #(
		.INIT('hfc23)
	) name1632 (
		\State2_reg[0]/NET0131 ,
		\State2_reg[1]/NET0131 ,
		\State2_reg[2]/NET0131 ,
		\State2_reg[3]/NET0131 ,
		_w2085_
	);
	LUT2 #(
		.INIT('h2)
	) name1633 (
		\uWord_reg[12]/NET0131 ,
		_w1841_,
		_w2086_
	);
	LUT4 #(
		.INIT('h0001)
	) name1634 (
		\EAX_reg[13]/NET0131 ,
		\EAX_reg[14]/NET0131 ,
		\EAX_reg[15]/NET0131 ,
		\EAX_reg[1]/NET0131 ,
		_w2087_
	);
	LUT4 #(
		.INIT('h0001)
	) name1635 (
		\EAX_reg[0]/NET0131 ,
		\EAX_reg[10]/NET0131 ,
		\EAX_reg[11]/NET0131 ,
		\EAX_reg[12]/NET0131 ,
		_w2088_
	);
	LUT4 #(
		.INIT('h0001)
	) name1636 (
		\EAX_reg[6]/NET0131 ,
		\EAX_reg[7]/NET0131 ,
		\EAX_reg[8]/NET0131 ,
		\EAX_reg[9]/NET0131 ,
		_w2089_
	);
	LUT4 #(
		.INIT('h0001)
	) name1637 (
		\EAX_reg[2]/NET0131 ,
		\EAX_reg[3]/NET0131 ,
		\EAX_reg[4]/NET0131 ,
		\EAX_reg[5]/NET0131 ,
		_w2090_
	);
	LUT4 #(
		.INIT('h8000)
	) name1638 (
		_w2089_,
		_w2090_,
		_w2087_,
		_w2088_,
		_w2091_
	);
	LUT4 #(
		.INIT('h0080)
	) name1639 (
		\EAX_reg[16]/NET0131 ,
		\EAX_reg[17]/NET0131 ,
		\EAX_reg[31]/NET0131 ,
		_w2091_,
		_w2092_
	);
	LUT4 #(
		.INIT('h8000)
	) name1640 (
		\EAX_reg[18]/NET0131 ,
		_w1757_,
		_w1758_,
		_w2092_,
		_w2093_
	);
	LUT2 #(
		.INIT('h8)
	) name1641 (
		\EAX_reg[25]/NET0131 ,
		_w2093_,
		_w2094_
	);
	LUT3 #(
		.INIT('h80)
	) name1642 (
		\EAX_reg[25]/NET0131 ,
		_w1917_,
		_w2093_,
		_w2095_
	);
	LUT4 #(
		.INIT('h8000)
	) name1643 (
		\EAX_reg[25]/NET0131 ,
		\EAX_reg[28]/NET0131 ,
		_w1917_,
		_w2093_,
		_w2096_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name1644 (
		\EAX_reg[25]/NET0131 ,
		\EAX_reg[28]/NET0131 ,
		_w1917_,
		_w2093_,
		_w2097_
	);
	LUT3 #(
		.INIT('h20)
	) name1645 (
		_w589_,
		_w566_,
		_w2097_,
		_w2098_
	);
	LUT4 #(
		.INIT('h2202)
	) name1646 (
		\Datai[12]_pad ,
		READY_n_pad,
		_w563_,
		_w565_,
		_w2099_
	);
	LUT2 #(
		.INIT('h8)
	) name1647 (
		_w582_,
		_w2099_,
		_w2100_
	);
	LUT2 #(
		.INIT('h2)
	) name1648 (
		_w582_,
		_w566_,
		_w2101_
	);
	LUT3 #(
		.INIT('hf1)
	) name1649 (
		_w582_,
		_w589_,
		_w566_,
		_w2102_
	);
	LUT4 #(
		.INIT('h0074)
	) name1650 (
		READY_n_pad,
		_w582_,
		_w589_,
		_w566_,
		_w2103_
	);
	LUT4 #(
		.INIT('h0031)
	) name1651 (
		\uWord_reg[12]/NET0131 ,
		_w2100_,
		_w2103_,
		_w2098_,
		_w2104_
	);
	LUT3 #(
		.INIT('hce)
	) name1652 (
		_w690_,
		_w2086_,
		_w2104_,
		_w2105_
	);
	LUT3 #(
		.INIT('h80)
	) name1653 (
		\EBX_reg[28]/NET0131 ,
		_w1986_,
		_w1987_,
		_w2106_
	);
	LUT4 #(
		.INIT('h8000)
	) name1654 (
		\EBX_reg[28]/NET0131 ,
		\EBX_reg[29]/NET0131 ,
		_w1986_,
		_w1987_,
		_w2107_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name1655 (
		_w622_,
		_w1986_,
		_w1987_,
		_w1988_,
		_w2108_
	);
	LUT3 #(
		.INIT('h02)
	) name1656 (
		\EBX_reg[30]/NET0131 ,
		_w1990_,
		_w1991_,
		_w2109_
	);
	LUT3 #(
		.INIT('h90)
	) name1657 (
		_w1946_,
		_w1957_,
		_w1990_,
		_w2110_
	);
	LUT2 #(
		.INIT('h1)
	) name1658 (
		_w2109_,
		_w2110_,
		_w2111_
	);
	LUT4 #(
		.INIT('h1f00)
	) name1659 (
		\EBX_reg[30]/NET0131 ,
		_w2107_,
		_w2108_,
		_w2111_,
		_w2112_
	);
	LUT2 #(
		.INIT('h2)
	) name1660 (
		\EBX_reg[30]/NET0131 ,
		_w1841_,
		_w2113_
	);
	LUT3 #(
		.INIT('hf2)
	) name1661 (
		_w690_,
		_w2112_,
		_w2113_,
		_w2114_
	);
	LUT3 #(
		.INIT('h08)
	) name1662 (
		\PhyAddrPointer_reg[3]/NET0131 ,
		_w563_,
		_w673_,
		_w2115_
	);
	LUT3 #(
		.INIT('ha8)
	) name1663 (
		_w608_,
		_w1886_,
		_w2115_,
		_w2116_
	);
	LUT4 #(
		.INIT('h202a)
	) name1664 (
		\PhyAddrPointer_reg[3]/NET0131 ,
		_w634_,
		_w607_,
		_w608_,
		_w2117_
	);
	LUT4 #(
		.INIT('h00fd)
	) name1665 (
		_w671_,
		_w1891_,
		_w1890_,
		_w2117_,
		_w2118_
	);
	LUT2 #(
		.INIT('h2)
	) name1666 (
		\PhyAddrPointer_reg[3]/NET0131 ,
		_w1215_,
		_w2119_
	);
	LUT4 #(
		.INIT('h001f)
	) name1667 (
		\DataWidth_reg[1]/NET0131 ,
		\PhyAddrPointer_reg[1]/NET0131 ,
		\PhyAddrPointer_reg[2]/NET0131 ,
		\PhyAddrPointer_reg[3]/NET0131 ,
		_w2120_
	);
	LUT4 #(
		.INIT('he000)
	) name1668 (
		\DataWidth_reg[1]/NET0131 ,
		\PhyAddrPointer_reg[1]/NET0131 ,
		\PhyAddrPointer_reg[2]/NET0131 ,
		\PhyAddrPointer_reg[3]/NET0131 ,
		_w2121_
	);
	LUT3 #(
		.INIT('h02)
	) name1669 (
		_w695_,
		_w2121_,
		_w2120_,
		_w2122_
	);
	LUT3 #(
		.INIT('h78)
	) name1670 (
		\PhyAddrPointer_reg[1]/NET0131 ,
		\PhyAddrPointer_reg[2]/NET0131 ,
		\PhyAddrPointer_reg[3]/NET0131 ,
		_w2123_
	);
	LUT4 #(
		.INIT('h0777)
	) name1671 (
		\rEIP_reg[3]/NET0131 ,
		_w1080_,
		_w1212_,
		_w2123_,
		_w2124_
	);
	LUT3 #(
		.INIT('h10)
	) name1672 (
		_w2119_,
		_w2122_,
		_w2124_,
		_w2125_
	);
	LUT4 #(
		.INIT('h8aff)
	) name1673 (
		_w690_,
		_w2116_,
		_w2118_,
		_w2125_,
		_w2126_
	);
	LUT4 #(
		.INIT('h7447)
	) name1674 (
		\PhyAddrPointer_reg[5]/NET0131 ,
		_w674_,
		_w825_,
		_w1903_,
		_w2127_
	);
	LUT4 #(
		.INIT('h202a)
	) name1675 (
		\PhyAddrPointer_reg[5]/NET0131 ,
		_w634_,
		_w607_,
		_w608_,
		_w2128_
	);
	LUT4 #(
		.INIT('h007d)
	) name1676 (
		_w671_,
		_w1106_,
		_w1909_,
		_w2128_,
		_w2129_
	);
	LUT4 #(
		.INIT('h08cc)
	) name1677 (
		_w608_,
		_w690_,
		_w2127_,
		_w2129_,
		_w2130_
	);
	LUT4 #(
		.INIT('h7f4c)
	) name1678 (
		\PhyAddrPointer_reg[1]/NET0131 ,
		\PhyAddrPointer_reg[5]/NET0131 ,
		_w1190_,
		_w2009_,
		_w2131_
	);
	LUT2 #(
		.INIT('h8)
	) name1679 (
		_w1306_,
		_w2131_,
		_w2132_
	);
	LUT2 #(
		.INIT('h2)
	) name1680 (
		\PhyAddrPointer_reg[5]/NET0131 ,
		_w1215_,
		_w2133_
	);
	LUT4 #(
		.INIT('h2080)
	) name1681 (
		\DataWidth_reg[1]/NET0131 ,
		\PhyAddrPointer_reg[5]/NET0131 ,
		_w695_,
		_w1190_,
		_w2134_
	);
	LUT3 #(
		.INIT('h01)
	) name1682 (
		_w1913_,
		_w2134_,
		_w2133_,
		_w2135_
	);
	LUT2 #(
		.INIT('h4)
	) name1683 (
		_w2132_,
		_w2135_,
		_w2136_
	);
	LUT2 #(
		.INIT('hb)
	) name1684 (
		_w2130_,
		_w2136_,
		_w2137_
	);
	LUT4 #(
		.INIT('h7774)
	) name1685 (
		\PhyAddrPointer_reg[6]/NET0131 ,
		_w674_,
		_w1726_,
		_w1724_,
		_w2138_
	);
	LUT4 #(
		.INIT('h202a)
	) name1686 (
		\PhyAddrPointer_reg[6]/NET0131 ,
		_w634_,
		_w607_,
		_w608_,
		_w2139_
	);
	LUT4 #(
		.INIT('h00fd)
	) name1687 (
		_w671_,
		_w1731_,
		_w1729_,
		_w2139_,
		_w2140_
	);
	LUT4 #(
		.INIT('h08cc)
	) name1688 (
		_w608_,
		_w690_,
		_w2138_,
		_w2140_,
		_w2141_
	);
	LUT3 #(
		.INIT('h6c)
	) name1689 (
		\PhyAddrPointer_reg[1]/NET0131 ,
		\PhyAddrPointer_reg[6]/NET0131 ,
		_w1191_,
		_w2142_
	);
	LUT4 #(
		.INIT('h4105)
	) name1690 (
		\DataWidth_reg[1]/NET0131 ,
		\PhyAddrPointer_reg[1]/NET0131 ,
		\PhyAddrPointer_reg[6]/NET0131 ,
		_w1191_,
		_w2143_
	);
	LUT4 #(
		.INIT('h70d0)
	) name1691 (
		\DataWidth_reg[1]/NET0131 ,
		\PhyAddrPointer_reg[6]/NET0131 ,
		_w695_,
		_w1191_,
		_w2144_
	);
	LUT4 #(
		.INIT('h60c0)
	) name1692 (
		\PhyAddrPointer_reg[1]/NET0131 ,
		\PhyAddrPointer_reg[6]/NET0131 ,
		_w1212_,
		_w1191_,
		_w2145_
	);
	LUT4 #(
		.INIT('h3f15)
	) name1693 (
		\PhyAddrPointer_reg[6]/NET0131 ,
		\rEIP_reg[6]/NET0131 ,
		_w1080_,
		_w1215_,
		_w2146_
	);
	LUT4 #(
		.INIT('h4500)
	) name1694 (
		_w2145_,
		_w2143_,
		_w2144_,
		_w2146_,
		_w2147_
	);
	LUT2 #(
		.INIT('hb)
	) name1695 (
		_w2141_,
		_w2147_,
		_w2148_
	);
	LUT4 #(
		.INIT('hef00)
	) name1696 (
		_w614_,
		_w600_,
		_w638_,
		_w690_,
		_w2149_
	);
	LUT2 #(
		.INIT('h4)
	) name1697 (
		\Flush_reg/NET0131 ,
		\InstQueueRd_Addr_reg[3]/NET0131 ,
		_w2150_
	);
	LUT3 #(
		.INIT('ha8)
	) name1698 (
		_w700_,
		_w2000_,
		_w2150_,
		_w2151_
	);
	LUT4 #(
		.INIT('h45cf)
	) name1699 (
		\InstQueueRd_Addr_reg[3]/NET0131 ,
		_w631_,
		_w710_,
		_w1844_,
		_w2152_
	);
	LUT2 #(
		.INIT('h4)
	) name1700 (
		_w2151_,
		_w2152_,
		_w2153_
	);
	LUT2 #(
		.INIT('hb)
	) name1701 (
		_w2149_,
		_w2153_,
		_w2154_
	);
	LUT4 #(
		.INIT('h1333)
	) name1702 (
		\EAX_reg[28]/NET0131 ,
		\EAX_reg[29]/NET0131 ,
		_w1760_,
		_w1917_,
		_w2155_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name1703 (
		_w1741_,
		_w1760_,
		_w1917_,
		_w1918_,
		_w2156_
	);
	LUT3 #(
		.INIT('h08)
	) name1704 (
		_w494_,
		_w586_,
		_w652_,
		_w2157_
	);
	LUT4 #(
		.INIT('h02fd)
	) name1705 (
		_w1821_,
		_w1832_,
		_w1934_,
		_w1945_,
		_w2158_
	);
	LUT4 #(
		.INIT('h8000)
	) name1706 (
		\Datai[29]_pad ,
		_w494_,
		_w586_,
		_w652_,
		_w2159_
	);
	LUT4 #(
		.INIT('h88a8)
	) name1707 (
		\EAX_reg[29]/NET0131 ,
		READY_n_pad,
		_w563_,
		_w565_,
		_w2160_
	);
	LUT4 #(
		.INIT('h2202)
	) name1708 (
		\Datai[13]_pad ,
		READY_n_pad,
		_w563_,
		_w565_,
		_w2161_
	);
	LUT2 #(
		.INIT('h1)
	) name1709 (
		_w2160_,
		_w2161_,
		_w2162_
	);
	LUT2 #(
		.INIT('h2)
	) name1710 (
		_w582_,
		_w2162_,
		_w2163_
	);
	LUT4 #(
		.INIT('h0013)
	) name1711 (
		_w1740_,
		_w2159_,
		_w2158_,
		_w2163_,
		_w2164_
	);
	LUT4 #(
		.INIT('h5700)
	) name1712 (
		\EAX_reg[29]/NET0131 ,
		_w1742_,
		_w2157_,
		_w2164_,
		_w2165_
	);
	LUT4 #(
		.INIT('h20aa)
	) name1713 (
		_w690_,
		_w2155_,
		_w2156_,
		_w2165_,
		_w2166_
	);
	LUT2 #(
		.INIT('h2)
	) name1714 (
		\EAX_reg[29]/NET0131 ,
		_w1841_,
		_w2167_
	);
	LUT2 #(
		.INIT('he)
	) name1715 (
		_w2166_,
		_w2167_,
		_w2168_
	);
	LUT4 #(
		.INIT('h8000)
	) name1716 (
		_w569_,
		_w602_,
		_w634_,
		_w2076_,
		_w2169_
	);
	LUT4 #(
		.INIT('h00fd)
	) name1717 (
		\EBX_reg[26]/NET0131 ,
		_w1990_,
		_w1991_,
		_w2169_,
		_w2170_
	);
	LUT4 #(
		.INIT('hb700)
	) name1718 (
		\EBX_reg[26]/NET0131 ,
		_w622_,
		_w1986_,
		_w2170_,
		_w2171_
	);
	LUT2 #(
		.INIT('h2)
	) name1719 (
		\EBX_reg[26]/NET0131 ,
		_w1841_,
		_w2172_
	);
	LUT3 #(
		.INIT('hf2)
	) name1720 (
		_w690_,
		_w2171_,
		_w2172_,
		_w2173_
	);
	LUT4 #(
		.INIT('h8000)
	) name1721 (
		\EAX_reg[18]/NET0131 ,
		\EAX_reg[23]/NET0131 ,
		_w1757_,
		_w2092_,
		_w2174_
	);
	LUT2 #(
		.INIT('h1)
	) name1722 (
		\EAX_reg[24]/NET0131 ,
		_w2174_,
		_w2175_
	);
	LUT3 #(
		.INIT('h02)
	) name1723 (
		_w589_,
		_w2093_,
		_w2175_,
		_w2176_
	);
	LUT4 #(
		.INIT('h0008)
	) name1724 (
		_w589_,
		_w595_,
		_w2093_,
		_w2175_,
		_w2177_
	);
	LUT4 #(
		.INIT('hf020)
	) name1725 (
		\Datao[24]_pad ,
		_w596_,
		_w690_,
		_w2177_,
		_w2178_
	);
	LUT4 #(
		.INIT('h0040)
	) name1726 (
		\State2_reg[0]/NET0131 ,
		\State2_reg[1]/NET0131 ,
		\State2_reg[2]/NET0131 ,
		\State2_reg[3]/NET0131 ,
		_w2179_
	);
	LUT4 #(
		.INIT('hfc60)
	) name1727 (
		\State2_reg[0]/NET0131 ,
		\State2_reg[1]/NET0131 ,
		\State2_reg[2]/NET0131 ,
		\State2_reg[3]/NET0131 ,
		_w2180_
	);
	LUT4 #(
		.INIT('h3f15)
	) name1728 (
		\Datao[24]_pad ,
		\uWord_reg[8]/NET0131 ,
		_w2179_,
		_w2180_,
		_w2181_
	);
	LUT2 #(
		.INIT('hb)
	) name1729 (
		_w2178_,
		_w2181_,
		_w2182_
	);
	LUT3 #(
		.INIT('h80)
	) name1730 (
		_w585_,
		_w590_,
		_w594_,
		_w2183_
	);
	LUT4 #(
		.INIT('h0a08)
	) name1731 (
		_w589_,
		_w594_,
		_w566_,
		_w2097_,
		_w2184_
	);
	LUT4 #(
		.INIT('haaa2)
	) name1732 (
		\Datao[28]_pad ,
		_w646_,
		_w2183_,
		_w2184_,
		_w2185_
	);
	LUT3 #(
		.INIT('h80)
	) name1733 (
		_w589_,
		_w595_,
		_w2097_,
		_w2186_
	);
	LUT4 #(
		.INIT('h3f15)
	) name1734 (
		\Datao[28]_pad ,
		\uWord_reg[12]/NET0131 ,
		_w2179_,
		_w2180_,
		_w2187_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name1735 (
		_w690_,
		_w2185_,
		_w2186_,
		_w2187_,
		_w2188_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name1736 (
		\uWord_reg[8]/NET0131 ,
		_w690_,
		_w1841_,
		_w2103_,
		_w2189_
	);
	LUT2 #(
		.INIT('h2)
	) name1737 (
		\Datai[8]_pad ,
		READY_n_pad,
		_w2190_
	);
	LUT2 #(
		.INIT('h8)
	) name1738 (
		_w582_,
		_w2190_,
		_w2191_
	);
	LUT3 #(
		.INIT('hd0)
	) name1739 (
		_w563_,
		_w565_,
		_w690_,
		_w2192_
	);
	LUT3 #(
		.INIT('he0)
	) name1740 (
		_w2176_,
		_w2191_,
		_w2192_,
		_w2193_
	);
	LUT2 #(
		.INIT('he)
	) name1741 (
		_w2189_,
		_w2193_,
		_w2194_
	);
	LUT2 #(
		.INIT('h2)
	) name1742 (
		\EBX_reg[29]/NET0131 ,
		_w1841_,
		_w2195_
	);
	LUT4 #(
		.INIT('h31fd)
	) name1743 (
		\EBX_reg[29]/NET0131 ,
		_w1990_,
		_w1991_,
		_w2158_,
		_w2196_
	);
	LUT4 #(
		.INIT('hb700)
	) name1744 (
		\EBX_reg[29]/NET0131 ,
		_w622_,
		_w2106_,
		_w2196_,
		_w2197_
	);
	LUT3 #(
		.INIT('hce)
	) name1745 (
		_w690_,
		_w2195_,
		_w2197_,
		_w2198_
	);
	LUT4 #(
		.INIT('h2000)
	) name1746 (
		\InstQueueWr_Addr_reg[0]/NET0131 ,
		\InstQueueWr_Addr_reg[1]/NET0131 ,
		\InstQueueWr_Addr_reg[2]/NET0131 ,
		\InstQueueWr_Addr_reg[3]/NET0131 ,
		_w2199_
	);
	LUT4 #(
		.INIT('h0001)
	) name1747 (
		\Datai[13]_pad ,
		\Datai[14]_pad ,
		\Datai[15]_pad ,
		\Datai[1]_pad ,
		_w2200_
	);
	LUT4 #(
		.INIT('h0001)
	) name1748 (
		\Datai[0]_pad ,
		\Datai[10]_pad ,
		\Datai[11]_pad ,
		\Datai[12]_pad ,
		_w2201_
	);
	LUT4 #(
		.INIT('h0001)
	) name1749 (
		\Datai[6]_pad ,
		\Datai[7]_pad ,
		\Datai[8]_pad ,
		\Datai[9]_pad ,
		_w2202_
	);
	LUT4 #(
		.INIT('h0001)
	) name1750 (
		\Datai[2]_pad ,
		\Datai[3]_pad ,
		\Datai[4]_pad ,
		\Datai[5]_pad ,
		_w2203_
	);
	LUT4 #(
		.INIT('h8000)
	) name1751 (
		_w2202_,
		_w2203_,
		_w2200_,
		_w2201_,
		_w2204_
	);
	LUT4 #(
		.INIT('h0001)
	) name1752 (
		\Datai[20]_pad ,
		\Datai[21]_pad ,
		\Datai[22]_pad ,
		\Datai[23]_pad ,
		_w2205_
	);
	LUT4 #(
		.INIT('h0001)
	) name1753 (
		\Datai[16]_pad ,
		\Datai[17]_pad ,
		\Datai[18]_pad ,
		\Datai[19]_pad ,
		_w2206_
	);
	LUT2 #(
		.INIT('h8)
	) name1754 (
		_w2205_,
		_w2206_,
		_w2207_
	);
	LUT4 #(
		.INIT('h0888)
	) name1755 (
		\Datai[24]_pad ,
		\Datai[31]_pad ,
		_w2204_,
		_w2207_,
		_w2208_
	);
	LUT4 #(
		.INIT('h8000)
	) name1756 (
		\Datai[25]_pad ,
		\Datai[26]_pad ,
		\Datai[27]_pad ,
		_w2208_,
		_w2209_
	);
	LUT3 #(
		.INIT('h48)
	) name1757 (
		\Datai[28]_pad ,
		_w2199_,
		_w2209_,
		_w2210_
	);
	LUT4 #(
		.INIT('h0080)
	) name1758 (
		\Datai[16]_pad ,
		\Datai[17]_pad ,
		\Datai[31]_pad ,
		_w2204_,
		_w2211_
	);
	LUT4 #(
		.INIT('h8000)
	) name1759 (
		\Datai[18]_pad ,
		\Datai[19]_pad ,
		\Datai[20]_pad ,
		_w2211_,
		_w2212_
	);
	LUT4 #(
		.INIT('h78f0)
	) name1760 (
		\Datai[18]_pad ,
		\Datai[19]_pad ,
		\Datai[20]_pad ,
		_w2211_,
		_w2213_
	);
	LUT2 #(
		.INIT('h4)
	) name1761 (
		\InstQueueWr_Addr_reg[0]/NET0131 ,
		\InstQueueWr_Addr_reg[1]/NET0131 ,
		_w2214_
	);
	LUT4 #(
		.INIT('h4000)
	) name1762 (
		\InstQueueWr_Addr_reg[0]/NET0131 ,
		\InstQueueWr_Addr_reg[1]/NET0131 ,
		\InstQueueWr_Addr_reg[2]/NET0131 ,
		\InstQueueWr_Addr_reg[3]/NET0131 ,
		_w2215_
	);
	LUT2 #(
		.INIT('h8)
	) name1763 (
		_w2213_,
		_w2215_,
		_w2216_
	);
	LUT4 #(
		.INIT('h0001)
	) name1764 (
		\InstQueueWr_Addr_reg[0]/NET0131 ,
		\InstQueueWr_Addr_reg[1]/NET0131 ,
		\InstQueueWr_Addr_reg[2]/NET0131 ,
		\InstQueueWr_Addr_reg[3]/NET0131 ,
		_w2217_
	);
	LUT3 #(
		.INIT('h80)
	) name1765 (
		\InstQueueWr_Addr_reg[0]/NET0131 ,
		\InstQueueWr_Addr_reg[1]/NET0131 ,
		\InstQueueWr_Addr_reg[2]/NET0131 ,
		_w2218_
	);
	LUT4 #(
		.INIT('h8000)
	) name1766 (
		\InstQueueWr_Addr_reg[0]/NET0131 ,
		\InstQueueWr_Addr_reg[1]/NET0131 ,
		\InstQueueWr_Addr_reg[2]/NET0131 ,
		\InstQueueWr_Addr_reg[3]/NET0131 ,
		_w2219_
	);
	LUT4 #(
		.INIT('h7ffe)
	) name1767 (
		\InstQueueWr_Addr_reg[0]/NET0131 ,
		\InstQueueWr_Addr_reg[1]/NET0131 ,
		\InstQueueWr_Addr_reg[2]/NET0131 ,
		\InstQueueWr_Addr_reg[3]/NET0131 ,
		_w2220_
	);
	LUT4 #(
		.INIT('h5553)
	) name1768 (
		\Datai[4]_pad ,
		\InstQueue_reg[0][4]/NET0131 ,
		_w2217_,
		_w2219_,
		_w2221_
	);
	LUT4 #(
		.INIT('h9fff)
	) name1769 (
		\InstQueueWr_Addr_reg[0]/NET0131 ,
		\InstQueueWr_Addr_reg[1]/NET0131 ,
		\InstQueueWr_Addr_reg[2]/NET0131 ,
		\InstQueueWr_Addr_reg[3]/NET0131 ,
		_w2222_
	);
	LUT2 #(
		.INIT('h2)
	) name1770 (
		\DataWidth_reg[1]/NET0131 ,
		_w2222_,
		_w2223_
	);
	LUT2 #(
		.INIT('h1)
	) name1771 (
		_w2221_,
		_w2223_,
		_w2224_
	);
	LUT4 #(
		.INIT('h0057)
	) name1772 (
		\DataWidth_reg[1]/NET0131 ,
		_w2210_,
		_w2216_,
		_w2224_,
		_w2225_
	);
	LUT4 #(
		.INIT('hc055)
	) name1773 (
		\InstQueue_reg[0][4]/NET0131 ,
		_w574_,
		_w579_,
		_w2217_,
		_w2226_
	);
	LUT4 #(
		.INIT('hfd14)
	) name1774 (
		\State2_reg[0]/NET0131 ,
		\State2_reg[1]/NET0131 ,
		\State2_reg[2]/NET0131 ,
		\State2_reg[3]/NET0131 ,
		_w2227_
	);
	LUT2 #(
		.INIT('h2)
	) name1775 (
		\InstQueue_reg[0][4]/NET0131 ,
		_w2227_,
		_w2228_
	);
	LUT3 #(
		.INIT('h0d)
	) name1776 (
		_w1212_,
		_w2221_,
		_w2228_,
		_w2229_
	);
	LUT3 #(
		.INIT('hd0)
	) name1777 (
		_w710_,
		_w2226_,
		_w2229_,
		_w2230_
	);
	LUT3 #(
		.INIT('h2f)
	) name1778 (
		_w695_,
		_w2225_,
		_w2230_,
		_w2231_
	);
	LUT4 #(
		.INIT('h0080)
	) name1779 (
		\InstQueueWr_Addr_reg[0]/NET0131 ,
		\InstQueueWr_Addr_reg[1]/NET0131 ,
		\InstQueueWr_Addr_reg[2]/NET0131 ,
		\InstQueueWr_Addr_reg[3]/NET0131 ,
		_w2232_
	);
	LUT3 #(
		.INIT('h60)
	) name1780 (
		\Datai[28]_pad ,
		_w2209_,
		_w2232_,
		_w2233_
	);
	LUT4 #(
		.INIT('h0100)
	) name1781 (
		\InstQueueWr_Addr_reg[0]/NET0131 ,
		\InstQueueWr_Addr_reg[1]/NET0131 ,
		\InstQueueWr_Addr_reg[2]/NET0131 ,
		\InstQueueWr_Addr_reg[3]/NET0131 ,
		_w2234_
	);
	LUT2 #(
		.INIT('h8)
	) name1782 (
		_w2213_,
		_w2234_,
		_w2235_
	);
	LUT4 #(
		.INIT('h0400)
	) name1783 (
		\InstQueueWr_Addr_reg[0]/NET0131 ,
		\InstQueueWr_Addr_reg[1]/NET0131 ,
		\InstQueueWr_Addr_reg[2]/NET0131 ,
		\InstQueueWr_Addr_reg[3]/NET0131 ,
		_w2236_
	);
	LUT4 #(
		.INIT('h0200)
	) name1784 (
		\InstQueueWr_Addr_reg[0]/NET0131 ,
		\InstQueueWr_Addr_reg[1]/NET0131 ,
		\InstQueueWr_Addr_reg[2]/NET0131 ,
		\InstQueueWr_Addr_reg[3]/NET0131 ,
		_w2237_
	);
	LUT4 #(
		.INIT('hf9ff)
	) name1785 (
		\InstQueueWr_Addr_reg[0]/NET0131 ,
		\InstQueueWr_Addr_reg[1]/NET0131 ,
		\InstQueueWr_Addr_reg[2]/NET0131 ,
		\InstQueueWr_Addr_reg[3]/NET0131 ,
		_w2238_
	);
	LUT4 #(
		.INIT('h5553)
	) name1786 (
		\Datai[4]_pad ,
		\InstQueue_reg[10][4]/NET0131 ,
		_w2236_,
		_w2237_,
		_w2239_
	);
	LUT4 #(
		.INIT('hfe7f)
	) name1787 (
		\InstQueueWr_Addr_reg[0]/NET0131 ,
		\InstQueueWr_Addr_reg[1]/NET0131 ,
		\InstQueueWr_Addr_reg[2]/NET0131 ,
		\InstQueueWr_Addr_reg[3]/NET0131 ,
		_w2240_
	);
	LUT2 #(
		.INIT('h2)
	) name1788 (
		\DataWidth_reg[1]/NET0131 ,
		_w2240_,
		_w2241_
	);
	LUT2 #(
		.INIT('h1)
	) name1789 (
		_w2239_,
		_w2241_,
		_w2242_
	);
	LUT4 #(
		.INIT('h0057)
	) name1790 (
		\DataWidth_reg[1]/NET0131 ,
		_w2233_,
		_w2235_,
		_w2242_,
		_w2243_
	);
	LUT4 #(
		.INIT('hc055)
	) name1791 (
		\InstQueue_reg[10][4]/NET0131 ,
		_w574_,
		_w579_,
		_w2236_,
		_w2244_
	);
	LUT2 #(
		.INIT('h2)
	) name1792 (
		\InstQueue_reg[10][4]/NET0131 ,
		_w2227_,
		_w2245_
	);
	LUT3 #(
		.INIT('h0d)
	) name1793 (
		_w1212_,
		_w2239_,
		_w2245_,
		_w2246_
	);
	LUT3 #(
		.INIT('hd0)
	) name1794 (
		_w710_,
		_w2244_,
		_w2246_,
		_w2247_
	);
	LUT3 #(
		.INIT('h2f)
	) name1795 (
		_w695_,
		_w2243_,
		_w2247_,
		_w2248_
	);
	LUT3 #(
		.INIT('h60)
	) name1796 (
		\Datai[28]_pad ,
		_w2209_,
		_w2234_,
		_w2249_
	);
	LUT2 #(
		.INIT('h8)
	) name1797 (
		_w2213_,
		_w2237_,
		_w2250_
	);
	LUT4 #(
		.INIT('h0800)
	) name1798 (
		\InstQueueWr_Addr_reg[0]/NET0131 ,
		\InstQueueWr_Addr_reg[1]/NET0131 ,
		\InstQueueWr_Addr_reg[2]/NET0131 ,
		\InstQueueWr_Addr_reg[3]/NET0131 ,
		_w2251_
	);
	LUT4 #(
		.INIT('hf3ff)
	) name1799 (
		\InstQueueWr_Addr_reg[0]/NET0131 ,
		\InstQueueWr_Addr_reg[1]/NET0131 ,
		\InstQueueWr_Addr_reg[2]/NET0131 ,
		\InstQueueWr_Addr_reg[3]/NET0131 ,
		_w2252_
	);
	LUT4 #(
		.INIT('h5553)
	) name1800 (
		\Datai[4]_pad ,
		\InstQueue_reg[11][4]/NET0131 ,
		_w2236_,
		_w2251_,
		_w2253_
	);
	LUT4 #(
		.INIT('hfcff)
	) name1801 (
		\InstQueueWr_Addr_reg[0]/NET0131 ,
		\InstQueueWr_Addr_reg[1]/NET0131 ,
		\InstQueueWr_Addr_reg[2]/NET0131 ,
		\InstQueueWr_Addr_reg[3]/NET0131 ,
		_w2254_
	);
	LUT2 #(
		.INIT('h2)
	) name1802 (
		\DataWidth_reg[1]/NET0131 ,
		_w2254_,
		_w2255_
	);
	LUT2 #(
		.INIT('h1)
	) name1803 (
		_w2253_,
		_w2255_,
		_w2256_
	);
	LUT4 #(
		.INIT('h0057)
	) name1804 (
		\DataWidth_reg[1]/NET0131 ,
		_w2249_,
		_w2250_,
		_w2256_,
		_w2257_
	);
	LUT4 #(
		.INIT('hc055)
	) name1805 (
		\InstQueue_reg[11][4]/NET0131 ,
		_w574_,
		_w579_,
		_w2251_,
		_w2258_
	);
	LUT2 #(
		.INIT('h2)
	) name1806 (
		\InstQueue_reg[11][4]/NET0131 ,
		_w2227_,
		_w2259_
	);
	LUT3 #(
		.INIT('h0d)
	) name1807 (
		_w1212_,
		_w2253_,
		_w2259_,
		_w2260_
	);
	LUT3 #(
		.INIT('hd0)
	) name1808 (
		_w710_,
		_w2258_,
		_w2260_,
		_w2261_
	);
	LUT3 #(
		.INIT('h2f)
	) name1809 (
		_w695_,
		_w2257_,
		_w2261_,
		_w2262_
	);
	LUT3 #(
		.INIT('h60)
	) name1810 (
		\Datai[28]_pad ,
		_w2209_,
		_w2237_,
		_w2263_
	);
	LUT2 #(
		.INIT('h8)
	) name1811 (
		_w2213_,
		_w2236_,
		_w2264_
	);
	LUT4 #(
		.INIT('h1000)
	) name1812 (
		\InstQueueWr_Addr_reg[0]/NET0131 ,
		\InstQueueWr_Addr_reg[1]/NET0131 ,
		\InstQueueWr_Addr_reg[2]/NET0131 ,
		\InstQueueWr_Addr_reg[3]/NET0131 ,
		_w2265_
	);
	LUT4 #(
		.INIT('he7ff)
	) name1813 (
		\InstQueueWr_Addr_reg[0]/NET0131 ,
		\InstQueueWr_Addr_reg[1]/NET0131 ,
		\InstQueueWr_Addr_reg[2]/NET0131 ,
		\InstQueueWr_Addr_reg[3]/NET0131 ,
		_w2266_
	);
	LUT4 #(
		.INIT('h5553)
	) name1814 (
		\Datai[4]_pad ,
		\InstQueue_reg[12][4]/NET0131 ,
		_w2251_,
		_w2265_,
		_w2267_
	);
	LUT2 #(
		.INIT('h2)
	) name1815 (
		\DataWidth_reg[1]/NET0131 ,
		_w2238_,
		_w2268_
	);
	LUT2 #(
		.INIT('h1)
	) name1816 (
		_w2267_,
		_w2268_,
		_w2269_
	);
	LUT4 #(
		.INIT('h0057)
	) name1817 (
		\DataWidth_reg[1]/NET0131 ,
		_w2263_,
		_w2264_,
		_w2269_,
		_w2270_
	);
	LUT4 #(
		.INIT('hc055)
	) name1818 (
		\InstQueue_reg[12][4]/NET0131 ,
		_w574_,
		_w579_,
		_w2265_,
		_w2271_
	);
	LUT2 #(
		.INIT('h2)
	) name1819 (
		\InstQueue_reg[12][4]/NET0131 ,
		_w2227_,
		_w2272_
	);
	LUT3 #(
		.INIT('h0d)
	) name1820 (
		_w1212_,
		_w2267_,
		_w2272_,
		_w2273_
	);
	LUT3 #(
		.INIT('hd0)
	) name1821 (
		_w710_,
		_w2271_,
		_w2273_,
		_w2274_
	);
	LUT3 #(
		.INIT('h2f)
	) name1822 (
		_w695_,
		_w2270_,
		_w2274_,
		_w2275_
	);
	LUT3 #(
		.INIT('h60)
	) name1823 (
		\Datai[28]_pad ,
		_w2209_,
		_w2236_,
		_w2276_
	);
	LUT2 #(
		.INIT('h8)
	) name1824 (
		_w2213_,
		_w2251_,
		_w2277_
	);
	LUT4 #(
		.INIT('hcfff)
	) name1825 (
		\InstQueueWr_Addr_reg[0]/NET0131 ,
		\InstQueueWr_Addr_reg[1]/NET0131 ,
		\InstQueueWr_Addr_reg[2]/NET0131 ,
		\InstQueueWr_Addr_reg[3]/NET0131 ,
		_w2278_
	);
	LUT4 #(
		.INIT('h5553)
	) name1826 (
		\Datai[4]_pad ,
		\InstQueue_reg[13][4]/NET0131 ,
		_w2199_,
		_w2265_,
		_w2279_
	);
	LUT2 #(
		.INIT('h2)
	) name1827 (
		\DataWidth_reg[1]/NET0131 ,
		_w2252_,
		_w2280_
	);
	LUT2 #(
		.INIT('h1)
	) name1828 (
		_w2279_,
		_w2280_,
		_w2281_
	);
	LUT4 #(
		.INIT('h0057)
	) name1829 (
		\DataWidth_reg[1]/NET0131 ,
		_w2276_,
		_w2277_,
		_w2281_,
		_w2282_
	);
	LUT4 #(
		.INIT('hc055)
	) name1830 (
		\InstQueue_reg[13][4]/NET0131 ,
		_w574_,
		_w579_,
		_w2199_,
		_w2283_
	);
	LUT2 #(
		.INIT('h2)
	) name1831 (
		\InstQueue_reg[13][4]/NET0131 ,
		_w2227_,
		_w2284_
	);
	LUT3 #(
		.INIT('h0d)
	) name1832 (
		_w1212_,
		_w2279_,
		_w2284_,
		_w2285_
	);
	LUT3 #(
		.INIT('hd0)
	) name1833 (
		_w710_,
		_w2283_,
		_w2285_,
		_w2286_
	);
	LUT3 #(
		.INIT('h2f)
	) name1834 (
		_w695_,
		_w2282_,
		_w2286_,
		_w2287_
	);
	LUT3 #(
		.INIT('h60)
	) name1835 (
		\Datai[28]_pad ,
		_w2209_,
		_w2251_,
		_w2288_
	);
	LUT2 #(
		.INIT('h8)
	) name1836 (
		_w2213_,
		_w2265_,
		_w2289_
	);
	LUT4 #(
		.INIT('h5553)
	) name1837 (
		\Datai[4]_pad ,
		\InstQueue_reg[14][4]/NET0131 ,
		_w2199_,
		_w2215_,
		_w2290_
	);
	LUT2 #(
		.INIT('h2)
	) name1838 (
		\DataWidth_reg[1]/NET0131 ,
		_w2266_,
		_w2291_
	);
	LUT2 #(
		.INIT('h1)
	) name1839 (
		_w2290_,
		_w2291_,
		_w2292_
	);
	LUT4 #(
		.INIT('h0057)
	) name1840 (
		\DataWidth_reg[1]/NET0131 ,
		_w2288_,
		_w2289_,
		_w2292_,
		_w2293_
	);
	LUT4 #(
		.INIT('hc055)
	) name1841 (
		\InstQueue_reg[14][4]/NET0131 ,
		_w574_,
		_w579_,
		_w2215_,
		_w2294_
	);
	LUT2 #(
		.INIT('h2)
	) name1842 (
		\InstQueue_reg[14][4]/NET0131 ,
		_w2227_,
		_w2295_
	);
	LUT3 #(
		.INIT('h0d)
	) name1843 (
		_w1212_,
		_w2290_,
		_w2295_,
		_w2296_
	);
	LUT3 #(
		.INIT('hd0)
	) name1844 (
		_w710_,
		_w2294_,
		_w2296_,
		_w2297_
	);
	LUT3 #(
		.INIT('h2f)
	) name1845 (
		_w695_,
		_w2293_,
		_w2297_,
		_w2298_
	);
	LUT3 #(
		.INIT('h60)
	) name1846 (
		\Datai[28]_pad ,
		_w2209_,
		_w2265_,
		_w2299_
	);
	LUT2 #(
		.INIT('h8)
	) name1847 (
		_w2199_,
		_w2213_,
		_w2300_
	);
	LUT4 #(
		.INIT('h3fff)
	) name1848 (
		\InstQueueWr_Addr_reg[0]/NET0131 ,
		\InstQueueWr_Addr_reg[1]/NET0131 ,
		\InstQueueWr_Addr_reg[2]/NET0131 ,
		\InstQueueWr_Addr_reg[3]/NET0131 ,
		_w2301_
	);
	LUT4 #(
		.INIT('h5553)
	) name1849 (
		\Datai[4]_pad ,
		\InstQueue_reg[15][4]/NET0131 ,
		_w2219_,
		_w2215_,
		_w2302_
	);
	LUT2 #(
		.INIT('h2)
	) name1850 (
		\DataWidth_reg[1]/NET0131 ,
		_w2278_,
		_w2303_
	);
	LUT2 #(
		.INIT('h1)
	) name1851 (
		_w2302_,
		_w2303_,
		_w2304_
	);
	LUT4 #(
		.INIT('h0057)
	) name1852 (
		\DataWidth_reg[1]/NET0131 ,
		_w2299_,
		_w2300_,
		_w2304_,
		_w2305_
	);
	LUT4 #(
		.INIT('hc055)
	) name1853 (
		\InstQueue_reg[15][4]/NET0131 ,
		_w574_,
		_w579_,
		_w2219_,
		_w2306_
	);
	LUT2 #(
		.INIT('h2)
	) name1854 (
		\InstQueue_reg[15][4]/NET0131 ,
		_w2227_,
		_w2307_
	);
	LUT3 #(
		.INIT('h0d)
	) name1855 (
		_w1212_,
		_w2302_,
		_w2307_,
		_w2308_
	);
	LUT3 #(
		.INIT('hd0)
	) name1856 (
		_w710_,
		_w2306_,
		_w2308_,
		_w2309_
	);
	LUT3 #(
		.INIT('h2f)
	) name1857 (
		_w695_,
		_w2305_,
		_w2309_,
		_w2310_
	);
	LUT3 #(
		.INIT('h60)
	) name1858 (
		\Datai[28]_pad ,
		_w2209_,
		_w2215_,
		_w2311_
	);
	LUT2 #(
		.INIT('h8)
	) name1859 (
		_w2219_,
		_w2213_,
		_w2312_
	);
	LUT4 #(
		.INIT('h0002)
	) name1860 (
		\InstQueueWr_Addr_reg[0]/NET0131 ,
		\InstQueueWr_Addr_reg[1]/NET0131 ,
		\InstQueueWr_Addr_reg[2]/NET0131 ,
		\InstQueueWr_Addr_reg[3]/NET0131 ,
		_w2313_
	);
	LUT4 #(
		.INIT('hfffc)
	) name1861 (
		\InstQueueWr_Addr_reg[0]/NET0131 ,
		\InstQueueWr_Addr_reg[1]/NET0131 ,
		\InstQueueWr_Addr_reg[2]/NET0131 ,
		\InstQueueWr_Addr_reg[3]/NET0131 ,
		_w2314_
	);
	LUT4 #(
		.INIT('h5553)
	) name1862 (
		\Datai[4]_pad ,
		\InstQueue_reg[1][4]/NET0131 ,
		_w2217_,
		_w2313_,
		_w2315_
	);
	LUT2 #(
		.INIT('h2)
	) name1863 (
		\DataWidth_reg[1]/NET0131 ,
		_w2301_,
		_w2316_
	);
	LUT2 #(
		.INIT('h1)
	) name1864 (
		_w2315_,
		_w2316_,
		_w2317_
	);
	LUT4 #(
		.INIT('h0057)
	) name1865 (
		\DataWidth_reg[1]/NET0131 ,
		_w2311_,
		_w2312_,
		_w2317_,
		_w2318_
	);
	LUT4 #(
		.INIT('hc055)
	) name1866 (
		\InstQueue_reg[1][4]/NET0131 ,
		_w574_,
		_w579_,
		_w2313_,
		_w2319_
	);
	LUT2 #(
		.INIT('h2)
	) name1867 (
		\InstQueue_reg[1][4]/NET0131 ,
		_w2227_,
		_w2320_
	);
	LUT3 #(
		.INIT('h0d)
	) name1868 (
		_w1212_,
		_w2315_,
		_w2320_,
		_w2321_
	);
	LUT3 #(
		.INIT('hd0)
	) name1869 (
		_w710_,
		_w2319_,
		_w2321_,
		_w2322_
	);
	LUT3 #(
		.INIT('h2f)
	) name1870 (
		_w695_,
		_w2318_,
		_w2322_,
		_w2323_
	);
	LUT2 #(
		.INIT('h8)
	) name1871 (
		_w2217_,
		_w2213_,
		_w2324_
	);
	LUT3 #(
		.INIT('h48)
	) name1872 (
		\Datai[28]_pad ,
		_w2219_,
		_w2209_,
		_w2325_
	);
	LUT4 #(
		.INIT('h0004)
	) name1873 (
		\InstQueueWr_Addr_reg[0]/NET0131 ,
		\InstQueueWr_Addr_reg[1]/NET0131 ,
		\InstQueueWr_Addr_reg[2]/NET0131 ,
		\InstQueueWr_Addr_reg[3]/NET0131 ,
		_w2326_
	);
	LUT4 #(
		.INIT('hfff9)
	) name1874 (
		\InstQueueWr_Addr_reg[0]/NET0131 ,
		\InstQueueWr_Addr_reg[1]/NET0131 ,
		\InstQueueWr_Addr_reg[2]/NET0131 ,
		\InstQueueWr_Addr_reg[3]/NET0131 ,
		_w2327_
	);
	LUT4 #(
		.INIT('h5553)
	) name1875 (
		\Datai[4]_pad ,
		\InstQueue_reg[2][4]/NET0131 ,
		_w2313_,
		_w2326_,
		_w2328_
	);
	LUT2 #(
		.INIT('h2)
	) name1876 (
		\DataWidth_reg[1]/NET0131 ,
		_w2220_,
		_w2329_
	);
	LUT2 #(
		.INIT('h1)
	) name1877 (
		_w2328_,
		_w2329_,
		_w2330_
	);
	LUT4 #(
		.INIT('h0057)
	) name1878 (
		\DataWidth_reg[1]/NET0131 ,
		_w2324_,
		_w2325_,
		_w2330_,
		_w2331_
	);
	LUT4 #(
		.INIT('hc055)
	) name1879 (
		\InstQueue_reg[2][4]/NET0131 ,
		_w574_,
		_w579_,
		_w2326_,
		_w2332_
	);
	LUT2 #(
		.INIT('h2)
	) name1880 (
		\InstQueue_reg[2][4]/NET0131 ,
		_w2227_,
		_w2333_
	);
	LUT3 #(
		.INIT('h0d)
	) name1881 (
		_w1212_,
		_w2328_,
		_w2333_,
		_w2334_
	);
	LUT3 #(
		.INIT('hd0)
	) name1882 (
		_w710_,
		_w2332_,
		_w2334_,
		_w2335_
	);
	LUT3 #(
		.INIT('h2f)
	) name1883 (
		_w695_,
		_w2331_,
		_w2335_,
		_w2336_
	);
	LUT3 #(
		.INIT('h48)
	) name1884 (
		\Datai[28]_pad ,
		_w2217_,
		_w2209_,
		_w2337_
	);
	LUT2 #(
		.INIT('h8)
	) name1885 (
		_w2213_,
		_w2313_,
		_w2338_
	);
	LUT4 #(
		.INIT('h0008)
	) name1886 (
		\InstQueueWr_Addr_reg[0]/NET0131 ,
		\InstQueueWr_Addr_reg[1]/NET0131 ,
		\InstQueueWr_Addr_reg[2]/NET0131 ,
		\InstQueueWr_Addr_reg[3]/NET0131 ,
		_w2339_
	);
	LUT4 #(
		.INIT('hfff3)
	) name1887 (
		\InstQueueWr_Addr_reg[0]/NET0131 ,
		\InstQueueWr_Addr_reg[1]/NET0131 ,
		\InstQueueWr_Addr_reg[2]/NET0131 ,
		\InstQueueWr_Addr_reg[3]/NET0131 ,
		_w2340_
	);
	LUT4 #(
		.INIT('h5553)
	) name1888 (
		\Datai[4]_pad ,
		\InstQueue_reg[3][4]/NET0131 ,
		_w2326_,
		_w2339_,
		_w2341_
	);
	LUT2 #(
		.INIT('h2)
	) name1889 (
		\DataWidth_reg[1]/NET0131 ,
		_w2314_,
		_w2342_
	);
	LUT2 #(
		.INIT('h1)
	) name1890 (
		_w2341_,
		_w2342_,
		_w2343_
	);
	LUT4 #(
		.INIT('h0057)
	) name1891 (
		\DataWidth_reg[1]/NET0131 ,
		_w2337_,
		_w2338_,
		_w2343_,
		_w2344_
	);
	LUT4 #(
		.INIT('hc055)
	) name1892 (
		\InstQueue_reg[3][4]/NET0131 ,
		_w574_,
		_w579_,
		_w2339_,
		_w2345_
	);
	LUT2 #(
		.INIT('h2)
	) name1893 (
		\InstQueue_reg[3][4]/NET0131 ,
		_w2227_,
		_w2346_
	);
	LUT3 #(
		.INIT('h0d)
	) name1894 (
		_w1212_,
		_w2341_,
		_w2346_,
		_w2347_
	);
	LUT3 #(
		.INIT('hd0)
	) name1895 (
		_w710_,
		_w2345_,
		_w2347_,
		_w2348_
	);
	LUT3 #(
		.INIT('h2f)
	) name1896 (
		_w695_,
		_w2344_,
		_w2348_,
		_w2349_
	);
	LUT3 #(
		.INIT('h60)
	) name1897 (
		\Datai[28]_pad ,
		_w2209_,
		_w2313_,
		_w2350_
	);
	LUT2 #(
		.INIT('h8)
	) name1898 (
		_w2213_,
		_w2326_,
		_w2351_
	);
	LUT4 #(
		.INIT('h0010)
	) name1899 (
		\InstQueueWr_Addr_reg[0]/NET0131 ,
		\InstQueueWr_Addr_reg[1]/NET0131 ,
		\InstQueueWr_Addr_reg[2]/NET0131 ,
		\InstQueueWr_Addr_reg[3]/NET0131 ,
		_w2352_
	);
	LUT4 #(
		.INIT('hffe7)
	) name1900 (
		\InstQueueWr_Addr_reg[0]/NET0131 ,
		\InstQueueWr_Addr_reg[1]/NET0131 ,
		\InstQueueWr_Addr_reg[2]/NET0131 ,
		\InstQueueWr_Addr_reg[3]/NET0131 ,
		_w2353_
	);
	LUT4 #(
		.INIT('h5553)
	) name1901 (
		\Datai[4]_pad ,
		\InstQueue_reg[4][4]/NET0131 ,
		_w2339_,
		_w2352_,
		_w2354_
	);
	LUT2 #(
		.INIT('h2)
	) name1902 (
		\DataWidth_reg[1]/NET0131 ,
		_w2327_,
		_w2355_
	);
	LUT2 #(
		.INIT('h1)
	) name1903 (
		_w2354_,
		_w2355_,
		_w2356_
	);
	LUT4 #(
		.INIT('h0057)
	) name1904 (
		\DataWidth_reg[1]/NET0131 ,
		_w2350_,
		_w2351_,
		_w2356_,
		_w2357_
	);
	LUT4 #(
		.INIT('hc055)
	) name1905 (
		\InstQueue_reg[4][4]/NET0131 ,
		_w574_,
		_w579_,
		_w2352_,
		_w2358_
	);
	LUT2 #(
		.INIT('h2)
	) name1906 (
		\InstQueue_reg[4][4]/NET0131 ,
		_w2227_,
		_w2359_
	);
	LUT3 #(
		.INIT('h0d)
	) name1907 (
		_w1212_,
		_w2354_,
		_w2359_,
		_w2360_
	);
	LUT3 #(
		.INIT('hd0)
	) name1908 (
		_w710_,
		_w2358_,
		_w2360_,
		_w2361_
	);
	LUT3 #(
		.INIT('h2f)
	) name1909 (
		_w695_,
		_w2357_,
		_w2361_,
		_w2362_
	);
	LUT3 #(
		.INIT('h60)
	) name1910 (
		\Datai[28]_pad ,
		_w2209_,
		_w2326_,
		_w2363_
	);
	LUT2 #(
		.INIT('h8)
	) name1911 (
		_w2213_,
		_w2339_,
		_w2364_
	);
	LUT4 #(
		.INIT('h0020)
	) name1912 (
		\InstQueueWr_Addr_reg[0]/NET0131 ,
		\InstQueueWr_Addr_reg[1]/NET0131 ,
		\InstQueueWr_Addr_reg[2]/NET0131 ,
		\InstQueueWr_Addr_reg[3]/NET0131 ,
		_w2365_
	);
	LUT4 #(
		.INIT('hffcf)
	) name1913 (
		\InstQueueWr_Addr_reg[0]/NET0131 ,
		\InstQueueWr_Addr_reg[1]/NET0131 ,
		\InstQueueWr_Addr_reg[2]/NET0131 ,
		\InstQueueWr_Addr_reg[3]/NET0131 ,
		_w2366_
	);
	LUT4 #(
		.INIT('h5553)
	) name1914 (
		\Datai[4]_pad ,
		\InstQueue_reg[5][4]/NET0131 ,
		_w2352_,
		_w2365_,
		_w2367_
	);
	LUT2 #(
		.INIT('h2)
	) name1915 (
		\DataWidth_reg[1]/NET0131 ,
		_w2340_,
		_w2368_
	);
	LUT2 #(
		.INIT('h1)
	) name1916 (
		_w2367_,
		_w2368_,
		_w2369_
	);
	LUT4 #(
		.INIT('h0057)
	) name1917 (
		\DataWidth_reg[1]/NET0131 ,
		_w2363_,
		_w2364_,
		_w2369_,
		_w2370_
	);
	LUT4 #(
		.INIT('hc055)
	) name1918 (
		\InstQueue_reg[5][4]/NET0131 ,
		_w574_,
		_w579_,
		_w2365_,
		_w2371_
	);
	LUT2 #(
		.INIT('h2)
	) name1919 (
		\InstQueue_reg[5][4]/NET0131 ,
		_w2227_,
		_w2372_
	);
	LUT3 #(
		.INIT('h0d)
	) name1920 (
		_w1212_,
		_w2367_,
		_w2372_,
		_w2373_
	);
	LUT3 #(
		.INIT('hd0)
	) name1921 (
		_w710_,
		_w2371_,
		_w2373_,
		_w2374_
	);
	LUT3 #(
		.INIT('h2f)
	) name1922 (
		_w695_,
		_w2370_,
		_w2374_,
		_w2375_
	);
	LUT3 #(
		.INIT('h60)
	) name1923 (
		\Datai[28]_pad ,
		_w2209_,
		_w2339_,
		_w2376_
	);
	LUT2 #(
		.INIT('h8)
	) name1924 (
		_w2213_,
		_w2352_,
		_w2377_
	);
	LUT4 #(
		.INIT('h0040)
	) name1925 (
		\InstQueueWr_Addr_reg[0]/NET0131 ,
		\InstQueueWr_Addr_reg[1]/NET0131 ,
		\InstQueueWr_Addr_reg[2]/NET0131 ,
		\InstQueueWr_Addr_reg[3]/NET0131 ,
		_w2378_
	);
	LUT4 #(
		.INIT('hff9f)
	) name1926 (
		\InstQueueWr_Addr_reg[0]/NET0131 ,
		\InstQueueWr_Addr_reg[1]/NET0131 ,
		\InstQueueWr_Addr_reg[2]/NET0131 ,
		\InstQueueWr_Addr_reg[3]/NET0131 ,
		_w2379_
	);
	LUT4 #(
		.INIT('h5553)
	) name1927 (
		\Datai[4]_pad ,
		\InstQueue_reg[6][4]/NET0131 ,
		_w2365_,
		_w2378_,
		_w2380_
	);
	LUT2 #(
		.INIT('h2)
	) name1928 (
		\DataWidth_reg[1]/NET0131 ,
		_w2353_,
		_w2381_
	);
	LUT2 #(
		.INIT('h1)
	) name1929 (
		_w2380_,
		_w2381_,
		_w2382_
	);
	LUT4 #(
		.INIT('h0057)
	) name1930 (
		\DataWidth_reg[1]/NET0131 ,
		_w2376_,
		_w2377_,
		_w2382_,
		_w2383_
	);
	LUT4 #(
		.INIT('hc055)
	) name1931 (
		\InstQueue_reg[6][4]/NET0131 ,
		_w574_,
		_w579_,
		_w2378_,
		_w2384_
	);
	LUT2 #(
		.INIT('h2)
	) name1932 (
		\InstQueue_reg[6][4]/NET0131 ,
		_w2227_,
		_w2385_
	);
	LUT3 #(
		.INIT('h0d)
	) name1933 (
		_w1212_,
		_w2380_,
		_w2385_,
		_w2386_
	);
	LUT3 #(
		.INIT('hd0)
	) name1934 (
		_w710_,
		_w2384_,
		_w2386_,
		_w2387_
	);
	LUT3 #(
		.INIT('h2f)
	) name1935 (
		_w695_,
		_w2383_,
		_w2387_,
		_w2388_
	);
	LUT3 #(
		.INIT('h60)
	) name1936 (
		\Datai[28]_pad ,
		_w2209_,
		_w2352_,
		_w2389_
	);
	LUT2 #(
		.INIT('h8)
	) name1937 (
		_w2213_,
		_w2365_,
		_w2390_
	);
	LUT4 #(
		.INIT('hff3f)
	) name1938 (
		\InstQueueWr_Addr_reg[0]/NET0131 ,
		\InstQueueWr_Addr_reg[1]/NET0131 ,
		\InstQueueWr_Addr_reg[2]/NET0131 ,
		\InstQueueWr_Addr_reg[3]/NET0131 ,
		_w2391_
	);
	LUT4 #(
		.INIT('h5553)
	) name1939 (
		\Datai[4]_pad ,
		\InstQueue_reg[7][4]/NET0131 ,
		_w2232_,
		_w2378_,
		_w2392_
	);
	LUT2 #(
		.INIT('h2)
	) name1940 (
		\DataWidth_reg[1]/NET0131 ,
		_w2366_,
		_w2393_
	);
	LUT2 #(
		.INIT('h1)
	) name1941 (
		_w2392_,
		_w2393_,
		_w2394_
	);
	LUT4 #(
		.INIT('h0057)
	) name1942 (
		\DataWidth_reg[1]/NET0131 ,
		_w2389_,
		_w2390_,
		_w2394_,
		_w2395_
	);
	LUT4 #(
		.INIT('hc055)
	) name1943 (
		\InstQueue_reg[7][4]/NET0131 ,
		_w574_,
		_w579_,
		_w2232_,
		_w2396_
	);
	LUT2 #(
		.INIT('h2)
	) name1944 (
		\InstQueue_reg[7][4]/NET0131 ,
		_w2227_,
		_w2397_
	);
	LUT3 #(
		.INIT('h0d)
	) name1945 (
		_w1212_,
		_w2392_,
		_w2397_,
		_w2398_
	);
	LUT3 #(
		.INIT('hd0)
	) name1946 (
		_w710_,
		_w2396_,
		_w2398_,
		_w2399_
	);
	LUT3 #(
		.INIT('h2f)
	) name1947 (
		_w695_,
		_w2395_,
		_w2399_,
		_w2400_
	);
	LUT3 #(
		.INIT('h60)
	) name1948 (
		\Datai[28]_pad ,
		_w2209_,
		_w2365_,
		_w2401_
	);
	LUT2 #(
		.INIT('h8)
	) name1949 (
		_w2213_,
		_w2378_,
		_w2402_
	);
	LUT4 #(
		.INIT('h5553)
	) name1950 (
		\Datai[4]_pad ,
		\InstQueue_reg[8][4]/NET0131 ,
		_w2232_,
		_w2234_,
		_w2403_
	);
	LUT2 #(
		.INIT('h2)
	) name1951 (
		\DataWidth_reg[1]/NET0131 ,
		_w2379_,
		_w2404_
	);
	LUT2 #(
		.INIT('h1)
	) name1952 (
		_w2403_,
		_w2404_,
		_w2405_
	);
	LUT4 #(
		.INIT('h0057)
	) name1953 (
		\DataWidth_reg[1]/NET0131 ,
		_w2401_,
		_w2402_,
		_w2405_,
		_w2406_
	);
	LUT4 #(
		.INIT('hc055)
	) name1954 (
		\InstQueue_reg[8][4]/NET0131 ,
		_w574_,
		_w579_,
		_w2234_,
		_w2407_
	);
	LUT2 #(
		.INIT('h2)
	) name1955 (
		\InstQueue_reg[8][4]/NET0131 ,
		_w2227_,
		_w2408_
	);
	LUT3 #(
		.INIT('h0d)
	) name1956 (
		_w1212_,
		_w2403_,
		_w2408_,
		_w2409_
	);
	LUT3 #(
		.INIT('hd0)
	) name1957 (
		_w710_,
		_w2407_,
		_w2409_,
		_w2410_
	);
	LUT3 #(
		.INIT('h2f)
	) name1958 (
		_w695_,
		_w2406_,
		_w2410_,
		_w2411_
	);
	LUT3 #(
		.INIT('h60)
	) name1959 (
		\Datai[28]_pad ,
		_w2209_,
		_w2378_,
		_w2412_
	);
	LUT2 #(
		.INIT('h8)
	) name1960 (
		_w2213_,
		_w2232_,
		_w2413_
	);
	LUT4 #(
		.INIT('h5553)
	) name1961 (
		\Datai[4]_pad ,
		\InstQueue_reg[9][4]/NET0131 ,
		_w2237_,
		_w2234_,
		_w2414_
	);
	LUT2 #(
		.INIT('h2)
	) name1962 (
		\DataWidth_reg[1]/NET0131 ,
		_w2391_,
		_w2415_
	);
	LUT2 #(
		.INIT('h1)
	) name1963 (
		_w2414_,
		_w2415_,
		_w2416_
	);
	LUT4 #(
		.INIT('h0057)
	) name1964 (
		\DataWidth_reg[1]/NET0131 ,
		_w2412_,
		_w2413_,
		_w2416_,
		_w2417_
	);
	LUT4 #(
		.INIT('hc055)
	) name1965 (
		\InstQueue_reg[9][4]/NET0131 ,
		_w574_,
		_w579_,
		_w2237_,
		_w2418_
	);
	LUT2 #(
		.INIT('h2)
	) name1966 (
		\InstQueue_reg[9][4]/NET0131 ,
		_w2227_,
		_w2419_
	);
	LUT3 #(
		.INIT('h0d)
	) name1967 (
		_w1212_,
		_w2414_,
		_w2419_,
		_w2420_
	);
	LUT3 #(
		.INIT('hd0)
	) name1968 (
		_w710_,
		_w2418_,
		_w2420_,
		_w2421_
	);
	LUT3 #(
		.INIT('h2f)
	) name1969 (
		_w695_,
		_w2417_,
		_w2421_,
		_w2422_
	);
	LUT3 #(
		.INIT('h02)
	) name1970 (
		_w608_,
		_w674_,
		_w2020_,
		_w2423_
	);
	LUT4 #(
		.INIT('h000d)
	) name1971 (
		\PhyAddrPointer_reg[2]/NET0131 ,
		_w1634_,
		_w2027_,
		_w2423_,
		_w2424_
	);
	LUT2 #(
		.INIT('h2)
	) name1972 (
		\PhyAddrPointer_reg[2]/NET0131 ,
		_w1215_,
		_w2425_
	);
	LUT2 #(
		.INIT('h6)
	) name1973 (
		\PhyAddrPointer_reg[1]/NET0131 ,
		\PhyAddrPointer_reg[2]/NET0131 ,
		_w2426_
	);
	LUT4 #(
		.INIT('hf400)
	) name1974 (
		\DataWidth_reg[1]/NET0131 ,
		_w695_,
		_w1212_,
		_w2426_,
		_w2427_
	);
	LUT3 #(
		.INIT('h20)
	) name1975 (
		\DataWidth_reg[1]/NET0131 ,
		\PhyAddrPointer_reg[2]/NET0131 ,
		_w695_,
		_w2428_
	);
	LUT4 #(
		.INIT('h0001)
	) name1976 (
		_w2031_,
		_w2427_,
		_w2425_,
		_w2428_,
		_w2429_
	);
	LUT3 #(
		.INIT('h2f)
	) name1977 (
		_w690_,
		_w2424_,
		_w2429_,
		_w2430_
	);
	LUT4 #(
		.INIT('h8000)
	) name1978 (
		\EAX_reg[18]/NET0131 ,
		\EAX_reg[19]/NET0131 ,
		\EAX_reg[20]/NET0131 ,
		_w2092_,
		_w2431_
	);
	LUT4 #(
		.INIT('h78f0)
	) name1979 (
		\EAX_reg[18]/NET0131 ,
		\EAX_reg[19]/NET0131 ,
		\EAX_reg[20]/NET0131 ,
		_w2092_,
		_w2432_
	);
	LUT2 #(
		.INIT('h1)
	) name1980 (
		_w594_,
		_w2432_,
		_w2433_
	);
	LUT3 #(
		.INIT('h02)
	) name1981 (
		_w589_,
		_w566_,
		_w2433_,
		_w2434_
	);
	LUT4 #(
		.INIT('haaa2)
	) name1982 (
		\Datao[20]_pad ,
		_w646_,
		_w2183_,
		_w2434_,
		_w2435_
	);
	LUT3 #(
		.INIT('h20)
	) name1983 (
		_w589_,
		_w566_,
		_w2432_,
		_w2436_
	);
	LUT4 #(
		.INIT('h0200)
	) name1984 (
		_w589_,
		_w594_,
		_w566_,
		_w2432_,
		_w2437_
	);
	LUT4 #(
		.INIT('h3f15)
	) name1985 (
		\Datao[20]_pad ,
		\uWord_reg[4]/NET0131 ,
		_w2179_,
		_w2180_,
		_w2438_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name1986 (
		_w690_,
		_w2435_,
		_w2437_,
		_w2438_,
		_w2439_
	);
	LUT2 #(
		.INIT('h2)
	) name1987 (
		\uWord_reg[4]/NET0131 ,
		_w1841_,
		_w2440_
	);
	LUT2 #(
		.INIT('h8)
	) name1988 (
		READY_n_pad,
		\uWord_reg[4]/NET0131 ,
		_w2441_
	);
	LUT4 #(
		.INIT('h2202)
	) name1989 (
		\Datai[4]_pad ,
		READY_n_pad,
		_w563_,
		_w565_,
		_w2442_
	);
	LUT2 #(
		.INIT('h1)
	) name1990 (
		_w2441_,
		_w2442_,
		_w2443_
	);
	LUT2 #(
		.INIT('h2)
	) name1991 (
		_w582_,
		_w2443_,
		_w2444_
	);
	LUT4 #(
		.INIT('haa02)
	) name1992 (
		\uWord_reg[4]/NET0131 ,
		_w582_,
		_w589_,
		_w566_,
		_w2445_
	);
	LUT4 #(
		.INIT('haaa8)
	) name1993 (
		_w690_,
		_w2436_,
		_w2444_,
		_w2445_,
		_w2446_
	);
	LUT2 #(
		.INIT('he)
	) name1994 (
		_w2440_,
		_w2446_,
		_w2447_
	);
	LUT3 #(
		.INIT('h48)
	) name1995 (
		\EAX_reg[25]/NET0131 ,
		_w1741_,
		_w1759_,
		_w2448_
	);
	LUT4 #(
		.INIT('h88a8)
	) name1996 (
		\EAX_reg[25]/NET0131 ,
		READY_n_pad,
		_w563_,
		_w565_,
		_w2449_
	);
	LUT4 #(
		.INIT('h2202)
	) name1997 (
		\Datai[25]_pad ,
		READY_n_pad,
		_w563_,
		_w565_,
		_w2450_
	);
	LUT2 #(
		.INIT('h1)
	) name1998 (
		_w2449_,
		_w2450_,
		_w2451_
	);
	LUT3 #(
		.INIT('h08)
	) name1999 (
		_w494_,
		_w586_,
		_w2451_,
		_w2452_
	);
	LUT3 #(
		.INIT('h2d)
	) name2000 (
		_w1787_,
		_w1798_,
		_w1809_,
		_w2453_
	);
	LUT4 #(
		.INIT('h8000)
	) name2001 (
		_w602_,
		_w604_,
		_w634_,
		_w2453_,
		_w2454_
	);
	LUT4 #(
		.INIT('h2202)
	) name2002 (
		\Datai[9]_pad ,
		READY_n_pad,
		_w563_,
		_w565_,
		_w2455_
	);
	LUT2 #(
		.INIT('h1)
	) name2003 (
		_w2449_,
		_w2455_,
		_w2456_
	);
	LUT2 #(
		.INIT('h2)
	) name2004 (
		_w582_,
		_w2456_,
		_w2457_
	);
	LUT3 #(
		.INIT('h01)
	) name2005 (
		_w2454_,
		_w2457_,
		_w2452_,
		_w2458_
	);
	LUT3 #(
		.INIT('h70)
	) name2006 (
		\EAX_reg[25]/NET0131 ,
		_w1742_,
		_w2458_,
		_w2459_
	);
	LUT2 #(
		.INIT('h2)
	) name2007 (
		\EAX_reg[25]/NET0131 ,
		_w1841_,
		_w2460_
	);
	LUT4 #(
		.INIT('hff8a)
	) name2008 (
		_w690_,
		_w2448_,
		_w2459_,
		_w2460_,
		_w2461_
	);
	LUT4 #(
		.INIT('h8000)
	) name2009 (
		\Datai[28]_pad ,
		\Datai[29]_pad ,
		\Datai[30]_pad ,
		_w2209_,
		_w2462_
	);
	LUT3 #(
		.INIT('h08)
	) name2010 (
		\Datai[31]_pad ,
		_w2199_,
		_w2462_,
		_w2463_
	);
	LUT4 #(
		.INIT('h78f0)
	) name2011 (
		\Datai[21]_pad ,
		\Datai[22]_pad ,
		\Datai[23]_pad ,
		_w2212_,
		_w2464_
	);
	LUT2 #(
		.INIT('h8)
	) name2012 (
		_w2215_,
		_w2464_,
		_w2465_
	);
	LUT4 #(
		.INIT('h5553)
	) name2013 (
		\Datai[7]_pad ,
		\InstQueue_reg[0][7]/NET0131 ,
		_w2217_,
		_w2219_,
		_w2466_
	);
	LUT2 #(
		.INIT('h1)
	) name2014 (
		_w2223_,
		_w2466_,
		_w2467_
	);
	LUT4 #(
		.INIT('h0057)
	) name2015 (
		\DataWidth_reg[1]/NET0131 ,
		_w2463_,
		_w2465_,
		_w2467_,
		_w2468_
	);
	LUT4 #(
		.INIT('hc055)
	) name2016 (
		\InstQueue_reg[0][7]/NET0131 ,
		_w546_,
		_w551_,
		_w2217_,
		_w2469_
	);
	LUT2 #(
		.INIT('h2)
	) name2017 (
		\InstQueue_reg[0][7]/NET0131 ,
		_w2227_,
		_w2470_
	);
	LUT3 #(
		.INIT('h0d)
	) name2018 (
		_w1212_,
		_w2466_,
		_w2470_,
		_w2471_
	);
	LUT3 #(
		.INIT('hd0)
	) name2019 (
		_w710_,
		_w2469_,
		_w2471_,
		_w2472_
	);
	LUT3 #(
		.INIT('h2f)
	) name2020 (
		_w695_,
		_w2468_,
		_w2472_,
		_w2473_
	);
	LUT3 #(
		.INIT('h08)
	) name2021 (
		\Datai[31]_pad ,
		_w2232_,
		_w2462_,
		_w2474_
	);
	LUT2 #(
		.INIT('h8)
	) name2022 (
		_w2234_,
		_w2464_,
		_w2475_
	);
	LUT4 #(
		.INIT('h5553)
	) name2023 (
		\Datai[7]_pad ,
		\InstQueue_reg[10][7]/NET0131 ,
		_w2236_,
		_w2237_,
		_w2476_
	);
	LUT2 #(
		.INIT('h1)
	) name2024 (
		_w2241_,
		_w2476_,
		_w2477_
	);
	LUT4 #(
		.INIT('h0057)
	) name2025 (
		\DataWidth_reg[1]/NET0131 ,
		_w2474_,
		_w2475_,
		_w2477_,
		_w2478_
	);
	LUT4 #(
		.INIT('hc055)
	) name2026 (
		\InstQueue_reg[10][7]/NET0131 ,
		_w546_,
		_w551_,
		_w2236_,
		_w2479_
	);
	LUT2 #(
		.INIT('h2)
	) name2027 (
		\InstQueue_reg[10][7]/NET0131 ,
		_w2227_,
		_w2480_
	);
	LUT3 #(
		.INIT('h0d)
	) name2028 (
		_w1212_,
		_w2476_,
		_w2480_,
		_w2481_
	);
	LUT3 #(
		.INIT('hd0)
	) name2029 (
		_w710_,
		_w2479_,
		_w2481_,
		_w2482_
	);
	LUT3 #(
		.INIT('h2f)
	) name2030 (
		_w695_,
		_w2478_,
		_w2482_,
		_w2483_
	);
	LUT3 #(
		.INIT('h08)
	) name2031 (
		\Datai[31]_pad ,
		_w2234_,
		_w2462_,
		_w2484_
	);
	LUT2 #(
		.INIT('h8)
	) name2032 (
		_w2237_,
		_w2464_,
		_w2485_
	);
	LUT4 #(
		.INIT('h5553)
	) name2033 (
		\Datai[7]_pad ,
		\InstQueue_reg[11][7]/NET0131 ,
		_w2236_,
		_w2251_,
		_w2486_
	);
	LUT2 #(
		.INIT('h1)
	) name2034 (
		_w2255_,
		_w2486_,
		_w2487_
	);
	LUT4 #(
		.INIT('h0057)
	) name2035 (
		\DataWidth_reg[1]/NET0131 ,
		_w2484_,
		_w2485_,
		_w2487_,
		_w2488_
	);
	LUT4 #(
		.INIT('hc055)
	) name2036 (
		\InstQueue_reg[11][7]/NET0131 ,
		_w546_,
		_w551_,
		_w2251_,
		_w2489_
	);
	LUT2 #(
		.INIT('h2)
	) name2037 (
		\InstQueue_reg[11][7]/NET0131 ,
		_w2227_,
		_w2490_
	);
	LUT3 #(
		.INIT('h0d)
	) name2038 (
		_w1212_,
		_w2486_,
		_w2490_,
		_w2491_
	);
	LUT3 #(
		.INIT('hd0)
	) name2039 (
		_w710_,
		_w2489_,
		_w2491_,
		_w2492_
	);
	LUT3 #(
		.INIT('h2f)
	) name2040 (
		_w695_,
		_w2488_,
		_w2492_,
		_w2493_
	);
	LUT3 #(
		.INIT('h08)
	) name2041 (
		\Datai[31]_pad ,
		_w2237_,
		_w2462_,
		_w2494_
	);
	LUT2 #(
		.INIT('h8)
	) name2042 (
		_w2236_,
		_w2464_,
		_w2495_
	);
	LUT4 #(
		.INIT('h5553)
	) name2043 (
		\Datai[7]_pad ,
		\InstQueue_reg[12][7]/NET0131 ,
		_w2251_,
		_w2265_,
		_w2496_
	);
	LUT2 #(
		.INIT('h1)
	) name2044 (
		_w2268_,
		_w2496_,
		_w2497_
	);
	LUT4 #(
		.INIT('h0057)
	) name2045 (
		\DataWidth_reg[1]/NET0131 ,
		_w2494_,
		_w2495_,
		_w2497_,
		_w2498_
	);
	LUT4 #(
		.INIT('hc055)
	) name2046 (
		\InstQueue_reg[12][7]/NET0131 ,
		_w546_,
		_w551_,
		_w2265_,
		_w2499_
	);
	LUT2 #(
		.INIT('h2)
	) name2047 (
		\InstQueue_reg[12][7]/NET0131 ,
		_w2227_,
		_w2500_
	);
	LUT3 #(
		.INIT('h0d)
	) name2048 (
		_w1212_,
		_w2496_,
		_w2500_,
		_w2501_
	);
	LUT3 #(
		.INIT('hd0)
	) name2049 (
		_w710_,
		_w2499_,
		_w2501_,
		_w2502_
	);
	LUT3 #(
		.INIT('h2f)
	) name2050 (
		_w695_,
		_w2498_,
		_w2502_,
		_w2503_
	);
	LUT3 #(
		.INIT('h08)
	) name2051 (
		\Datai[31]_pad ,
		_w2236_,
		_w2462_,
		_w2504_
	);
	LUT2 #(
		.INIT('h8)
	) name2052 (
		_w2251_,
		_w2464_,
		_w2505_
	);
	LUT4 #(
		.INIT('h5553)
	) name2053 (
		\Datai[7]_pad ,
		\InstQueue_reg[13][7]/NET0131 ,
		_w2199_,
		_w2265_,
		_w2506_
	);
	LUT2 #(
		.INIT('h1)
	) name2054 (
		_w2280_,
		_w2506_,
		_w2507_
	);
	LUT4 #(
		.INIT('h0057)
	) name2055 (
		\DataWidth_reg[1]/NET0131 ,
		_w2504_,
		_w2505_,
		_w2507_,
		_w2508_
	);
	LUT4 #(
		.INIT('hc055)
	) name2056 (
		\InstQueue_reg[13][7]/NET0131 ,
		_w546_,
		_w551_,
		_w2199_,
		_w2509_
	);
	LUT2 #(
		.INIT('h2)
	) name2057 (
		\InstQueue_reg[13][7]/NET0131 ,
		_w2227_,
		_w2510_
	);
	LUT3 #(
		.INIT('h0d)
	) name2058 (
		_w1212_,
		_w2506_,
		_w2510_,
		_w2511_
	);
	LUT3 #(
		.INIT('hd0)
	) name2059 (
		_w710_,
		_w2509_,
		_w2511_,
		_w2512_
	);
	LUT3 #(
		.INIT('h2f)
	) name2060 (
		_w695_,
		_w2508_,
		_w2512_,
		_w2513_
	);
	LUT3 #(
		.INIT('h08)
	) name2061 (
		\Datai[31]_pad ,
		_w2251_,
		_w2462_,
		_w2514_
	);
	LUT2 #(
		.INIT('h8)
	) name2062 (
		_w2265_,
		_w2464_,
		_w2515_
	);
	LUT4 #(
		.INIT('h5553)
	) name2063 (
		\Datai[7]_pad ,
		\InstQueue_reg[14][7]/NET0131 ,
		_w2199_,
		_w2215_,
		_w2516_
	);
	LUT2 #(
		.INIT('h1)
	) name2064 (
		_w2291_,
		_w2516_,
		_w2517_
	);
	LUT4 #(
		.INIT('h0057)
	) name2065 (
		\DataWidth_reg[1]/NET0131 ,
		_w2514_,
		_w2515_,
		_w2517_,
		_w2518_
	);
	LUT4 #(
		.INIT('hc055)
	) name2066 (
		\InstQueue_reg[14][7]/NET0131 ,
		_w546_,
		_w551_,
		_w2215_,
		_w2519_
	);
	LUT2 #(
		.INIT('h2)
	) name2067 (
		\InstQueue_reg[14][7]/NET0131 ,
		_w2227_,
		_w2520_
	);
	LUT3 #(
		.INIT('h0d)
	) name2068 (
		_w1212_,
		_w2516_,
		_w2520_,
		_w2521_
	);
	LUT3 #(
		.INIT('hd0)
	) name2069 (
		_w710_,
		_w2519_,
		_w2521_,
		_w2522_
	);
	LUT3 #(
		.INIT('h2f)
	) name2070 (
		_w695_,
		_w2518_,
		_w2522_,
		_w2523_
	);
	LUT3 #(
		.INIT('h08)
	) name2071 (
		\Datai[31]_pad ,
		_w2265_,
		_w2462_,
		_w2524_
	);
	LUT2 #(
		.INIT('h8)
	) name2072 (
		_w2199_,
		_w2464_,
		_w2525_
	);
	LUT4 #(
		.INIT('h5553)
	) name2073 (
		\Datai[7]_pad ,
		\InstQueue_reg[15][7]/NET0131 ,
		_w2219_,
		_w2215_,
		_w2526_
	);
	LUT2 #(
		.INIT('h1)
	) name2074 (
		_w2303_,
		_w2526_,
		_w2527_
	);
	LUT4 #(
		.INIT('h0057)
	) name2075 (
		\DataWidth_reg[1]/NET0131 ,
		_w2524_,
		_w2525_,
		_w2527_,
		_w2528_
	);
	LUT4 #(
		.INIT('hc055)
	) name2076 (
		\InstQueue_reg[15][7]/NET0131 ,
		_w546_,
		_w551_,
		_w2219_,
		_w2529_
	);
	LUT2 #(
		.INIT('h2)
	) name2077 (
		\InstQueue_reg[15][7]/NET0131 ,
		_w2227_,
		_w2530_
	);
	LUT3 #(
		.INIT('h0d)
	) name2078 (
		_w1212_,
		_w2526_,
		_w2530_,
		_w2531_
	);
	LUT3 #(
		.INIT('hd0)
	) name2079 (
		_w710_,
		_w2529_,
		_w2531_,
		_w2532_
	);
	LUT3 #(
		.INIT('h2f)
	) name2080 (
		_w695_,
		_w2528_,
		_w2532_,
		_w2533_
	);
	LUT3 #(
		.INIT('h08)
	) name2081 (
		\Datai[31]_pad ,
		_w2215_,
		_w2462_,
		_w2534_
	);
	LUT2 #(
		.INIT('h8)
	) name2082 (
		_w2219_,
		_w2464_,
		_w2535_
	);
	LUT4 #(
		.INIT('h5553)
	) name2083 (
		\Datai[7]_pad ,
		\InstQueue_reg[1][7]/NET0131 ,
		_w2217_,
		_w2313_,
		_w2536_
	);
	LUT2 #(
		.INIT('h1)
	) name2084 (
		_w2316_,
		_w2536_,
		_w2537_
	);
	LUT4 #(
		.INIT('h0057)
	) name2085 (
		\DataWidth_reg[1]/NET0131 ,
		_w2534_,
		_w2535_,
		_w2537_,
		_w2538_
	);
	LUT4 #(
		.INIT('hc055)
	) name2086 (
		\InstQueue_reg[1][7]/NET0131 ,
		_w546_,
		_w551_,
		_w2313_,
		_w2539_
	);
	LUT2 #(
		.INIT('h2)
	) name2087 (
		\InstQueue_reg[1][7]/NET0131 ,
		_w2227_,
		_w2540_
	);
	LUT3 #(
		.INIT('h0d)
	) name2088 (
		_w1212_,
		_w2536_,
		_w2540_,
		_w2541_
	);
	LUT3 #(
		.INIT('hd0)
	) name2089 (
		_w710_,
		_w2539_,
		_w2541_,
		_w2542_
	);
	LUT3 #(
		.INIT('h2f)
	) name2090 (
		_w695_,
		_w2538_,
		_w2542_,
		_w2543_
	);
	LUT2 #(
		.INIT('h8)
	) name2091 (
		_w2217_,
		_w2464_,
		_w2544_
	);
	LUT3 #(
		.INIT('h08)
	) name2092 (
		\Datai[31]_pad ,
		_w2219_,
		_w2462_,
		_w2545_
	);
	LUT4 #(
		.INIT('h5553)
	) name2093 (
		\Datai[7]_pad ,
		\InstQueue_reg[2][7]/NET0131 ,
		_w2313_,
		_w2326_,
		_w2546_
	);
	LUT2 #(
		.INIT('h1)
	) name2094 (
		_w2329_,
		_w2546_,
		_w2547_
	);
	LUT4 #(
		.INIT('h0057)
	) name2095 (
		\DataWidth_reg[1]/NET0131 ,
		_w2544_,
		_w2545_,
		_w2547_,
		_w2548_
	);
	LUT4 #(
		.INIT('hc055)
	) name2096 (
		\InstQueue_reg[2][7]/NET0131 ,
		_w546_,
		_w551_,
		_w2326_,
		_w2549_
	);
	LUT2 #(
		.INIT('h2)
	) name2097 (
		\InstQueue_reg[2][7]/NET0131 ,
		_w2227_,
		_w2550_
	);
	LUT3 #(
		.INIT('h0d)
	) name2098 (
		_w1212_,
		_w2546_,
		_w2550_,
		_w2551_
	);
	LUT3 #(
		.INIT('hd0)
	) name2099 (
		_w710_,
		_w2549_,
		_w2551_,
		_w2552_
	);
	LUT3 #(
		.INIT('h2f)
	) name2100 (
		_w695_,
		_w2548_,
		_w2552_,
		_w2553_
	);
	LUT3 #(
		.INIT('h08)
	) name2101 (
		\Datai[31]_pad ,
		_w2217_,
		_w2462_,
		_w2554_
	);
	LUT2 #(
		.INIT('h8)
	) name2102 (
		_w2313_,
		_w2464_,
		_w2555_
	);
	LUT4 #(
		.INIT('h5553)
	) name2103 (
		\Datai[7]_pad ,
		\InstQueue_reg[3][7]/NET0131 ,
		_w2326_,
		_w2339_,
		_w2556_
	);
	LUT2 #(
		.INIT('h1)
	) name2104 (
		_w2342_,
		_w2556_,
		_w2557_
	);
	LUT4 #(
		.INIT('h0057)
	) name2105 (
		\DataWidth_reg[1]/NET0131 ,
		_w2554_,
		_w2555_,
		_w2557_,
		_w2558_
	);
	LUT4 #(
		.INIT('hc055)
	) name2106 (
		\InstQueue_reg[3][7]/NET0131 ,
		_w546_,
		_w551_,
		_w2339_,
		_w2559_
	);
	LUT2 #(
		.INIT('h2)
	) name2107 (
		\InstQueue_reg[3][7]/NET0131 ,
		_w2227_,
		_w2560_
	);
	LUT3 #(
		.INIT('h0d)
	) name2108 (
		_w1212_,
		_w2556_,
		_w2560_,
		_w2561_
	);
	LUT3 #(
		.INIT('hd0)
	) name2109 (
		_w710_,
		_w2559_,
		_w2561_,
		_w2562_
	);
	LUT3 #(
		.INIT('h2f)
	) name2110 (
		_w695_,
		_w2558_,
		_w2562_,
		_w2563_
	);
	LUT3 #(
		.INIT('h08)
	) name2111 (
		\Datai[31]_pad ,
		_w2313_,
		_w2462_,
		_w2564_
	);
	LUT2 #(
		.INIT('h8)
	) name2112 (
		_w2326_,
		_w2464_,
		_w2565_
	);
	LUT4 #(
		.INIT('h5553)
	) name2113 (
		\Datai[7]_pad ,
		\InstQueue_reg[4][7]/NET0131 ,
		_w2339_,
		_w2352_,
		_w2566_
	);
	LUT2 #(
		.INIT('h1)
	) name2114 (
		_w2355_,
		_w2566_,
		_w2567_
	);
	LUT4 #(
		.INIT('h0057)
	) name2115 (
		\DataWidth_reg[1]/NET0131 ,
		_w2564_,
		_w2565_,
		_w2567_,
		_w2568_
	);
	LUT4 #(
		.INIT('hc055)
	) name2116 (
		\InstQueue_reg[4][7]/NET0131 ,
		_w546_,
		_w551_,
		_w2352_,
		_w2569_
	);
	LUT2 #(
		.INIT('h2)
	) name2117 (
		\InstQueue_reg[4][7]/NET0131 ,
		_w2227_,
		_w2570_
	);
	LUT3 #(
		.INIT('h0d)
	) name2118 (
		_w1212_,
		_w2566_,
		_w2570_,
		_w2571_
	);
	LUT3 #(
		.INIT('hd0)
	) name2119 (
		_w710_,
		_w2569_,
		_w2571_,
		_w2572_
	);
	LUT3 #(
		.INIT('h2f)
	) name2120 (
		_w695_,
		_w2568_,
		_w2572_,
		_w2573_
	);
	LUT3 #(
		.INIT('h08)
	) name2121 (
		\Datai[31]_pad ,
		_w2326_,
		_w2462_,
		_w2574_
	);
	LUT2 #(
		.INIT('h8)
	) name2122 (
		_w2339_,
		_w2464_,
		_w2575_
	);
	LUT4 #(
		.INIT('h5553)
	) name2123 (
		\Datai[7]_pad ,
		\InstQueue_reg[5][7]/NET0131 ,
		_w2352_,
		_w2365_,
		_w2576_
	);
	LUT2 #(
		.INIT('h1)
	) name2124 (
		_w2368_,
		_w2576_,
		_w2577_
	);
	LUT4 #(
		.INIT('h0057)
	) name2125 (
		\DataWidth_reg[1]/NET0131 ,
		_w2574_,
		_w2575_,
		_w2577_,
		_w2578_
	);
	LUT4 #(
		.INIT('hc055)
	) name2126 (
		\InstQueue_reg[5][7]/NET0131 ,
		_w546_,
		_w551_,
		_w2365_,
		_w2579_
	);
	LUT2 #(
		.INIT('h2)
	) name2127 (
		\InstQueue_reg[5][7]/NET0131 ,
		_w2227_,
		_w2580_
	);
	LUT3 #(
		.INIT('h0d)
	) name2128 (
		_w1212_,
		_w2576_,
		_w2580_,
		_w2581_
	);
	LUT3 #(
		.INIT('hd0)
	) name2129 (
		_w710_,
		_w2579_,
		_w2581_,
		_w2582_
	);
	LUT3 #(
		.INIT('h2f)
	) name2130 (
		_w695_,
		_w2578_,
		_w2582_,
		_w2583_
	);
	LUT3 #(
		.INIT('h08)
	) name2131 (
		\Datai[31]_pad ,
		_w2339_,
		_w2462_,
		_w2584_
	);
	LUT2 #(
		.INIT('h8)
	) name2132 (
		_w2352_,
		_w2464_,
		_w2585_
	);
	LUT4 #(
		.INIT('h5553)
	) name2133 (
		\Datai[7]_pad ,
		\InstQueue_reg[6][7]/NET0131 ,
		_w2365_,
		_w2378_,
		_w2586_
	);
	LUT2 #(
		.INIT('h1)
	) name2134 (
		_w2381_,
		_w2586_,
		_w2587_
	);
	LUT4 #(
		.INIT('h0057)
	) name2135 (
		\DataWidth_reg[1]/NET0131 ,
		_w2584_,
		_w2585_,
		_w2587_,
		_w2588_
	);
	LUT4 #(
		.INIT('hc055)
	) name2136 (
		\InstQueue_reg[6][7]/NET0131 ,
		_w546_,
		_w551_,
		_w2378_,
		_w2589_
	);
	LUT2 #(
		.INIT('h2)
	) name2137 (
		\InstQueue_reg[6][7]/NET0131 ,
		_w2227_,
		_w2590_
	);
	LUT3 #(
		.INIT('h0d)
	) name2138 (
		_w1212_,
		_w2586_,
		_w2590_,
		_w2591_
	);
	LUT3 #(
		.INIT('hd0)
	) name2139 (
		_w710_,
		_w2589_,
		_w2591_,
		_w2592_
	);
	LUT3 #(
		.INIT('h2f)
	) name2140 (
		_w695_,
		_w2588_,
		_w2592_,
		_w2593_
	);
	LUT3 #(
		.INIT('h08)
	) name2141 (
		\Datai[31]_pad ,
		_w2352_,
		_w2462_,
		_w2594_
	);
	LUT2 #(
		.INIT('h8)
	) name2142 (
		_w2365_,
		_w2464_,
		_w2595_
	);
	LUT4 #(
		.INIT('h5553)
	) name2143 (
		\Datai[7]_pad ,
		\InstQueue_reg[7][7]/NET0131 ,
		_w2232_,
		_w2378_,
		_w2596_
	);
	LUT2 #(
		.INIT('h1)
	) name2144 (
		_w2393_,
		_w2596_,
		_w2597_
	);
	LUT4 #(
		.INIT('h0057)
	) name2145 (
		\DataWidth_reg[1]/NET0131 ,
		_w2594_,
		_w2595_,
		_w2597_,
		_w2598_
	);
	LUT4 #(
		.INIT('hc055)
	) name2146 (
		\InstQueue_reg[7][7]/NET0131 ,
		_w546_,
		_w551_,
		_w2232_,
		_w2599_
	);
	LUT2 #(
		.INIT('h2)
	) name2147 (
		\InstQueue_reg[7][7]/NET0131 ,
		_w2227_,
		_w2600_
	);
	LUT3 #(
		.INIT('h0d)
	) name2148 (
		_w1212_,
		_w2596_,
		_w2600_,
		_w2601_
	);
	LUT3 #(
		.INIT('hd0)
	) name2149 (
		_w710_,
		_w2599_,
		_w2601_,
		_w2602_
	);
	LUT3 #(
		.INIT('h2f)
	) name2150 (
		_w695_,
		_w2598_,
		_w2602_,
		_w2603_
	);
	LUT3 #(
		.INIT('h08)
	) name2151 (
		\Datai[31]_pad ,
		_w2365_,
		_w2462_,
		_w2604_
	);
	LUT2 #(
		.INIT('h8)
	) name2152 (
		_w2378_,
		_w2464_,
		_w2605_
	);
	LUT4 #(
		.INIT('h5553)
	) name2153 (
		\Datai[7]_pad ,
		\InstQueue_reg[8][7]/NET0131 ,
		_w2232_,
		_w2234_,
		_w2606_
	);
	LUT2 #(
		.INIT('h1)
	) name2154 (
		_w2404_,
		_w2606_,
		_w2607_
	);
	LUT4 #(
		.INIT('h0057)
	) name2155 (
		\DataWidth_reg[1]/NET0131 ,
		_w2604_,
		_w2605_,
		_w2607_,
		_w2608_
	);
	LUT4 #(
		.INIT('hc055)
	) name2156 (
		\InstQueue_reg[8][7]/NET0131 ,
		_w546_,
		_w551_,
		_w2234_,
		_w2609_
	);
	LUT2 #(
		.INIT('h2)
	) name2157 (
		\InstQueue_reg[8][7]/NET0131 ,
		_w2227_,
		_w2610_
	);
	LUT3 #(
		.INIT('h0d)
	) name2158 (
		_w1212_,
		_w2606_,
		_w2610_,
		_w2611_
	);
	LUT3 #(
		.INIT('hd0)
	) name2159 (
		_w710_,
		_w2609_,
		_w2611_,
		_w2612_
	);
	LUT3 #(
		.INIT('h2f)
	) name2160 (
		_w695_,
		_w2608_,
		_w2612_,
		_w2613_
	);
	LUT3 #(
		.INIT('h08)
	) name2161 (
		\Datai[31]_pad ,
		_w2378_,
		_w2462_,
		_w2614_
	);
	LUT2 #(
		.INIT('h8)
	) name2162 (
		_w2232_,
		_w2464_,
		_w2615_
	);
	LUT4 #(
		.INIT('h5553)
	) name2163 (
		\Datai[7]_pad ,
		\InstQueue_reg[9][7]/NET0131 ,
		_w2237_,
		_w2234_,
		_w2616_
	);
	LUT2 #(
		.INIT('h1)
	) name2164 (
		_w2415_,
		_w2616_,
		_w2617_
	);
	LUT4 #(
		.INIT('h0057)
	) name2165 (
		\DataWidth_reg[1]/NET0131 ,
		_w2614_,
		_w2615_,
		_w2617_,
		_w2618_
	);
	LUT4 #(
		.INIT('hc055)
	) name2166 (
		\InstQueue_reg[9][7]/NET0131 ,
		_w546_,
		_w551_,
		_w2237_,
		_w2619_
	);
	LUT2 #(
		.INIT('h2)
	) name2167 (
		\InstQueue_reg[9][7]/NET0131 ,
		_w2227_,
		_w2620_
	);
	LUT3 #(
		.INIT('h0d)
	) name2168 (
		_w1212_,
		_w2616_,
		_w2620_,
		_w2621_
	);
	LUT3 #(
		.INIT('hd0)
	) name2169 (
		_w710_,
		_w2619_,
		_w2621_,
		_w2622_
	);
	LUT3 #(
		.INIT('h2f)
	) name2170 (
		_w695_,
		_w2618_,
		_w2622_,
		_w2623_
	);
	LUT4 #(
		.INIT('h070f)
	) name2171 (
		\EAX_reg[25]/NET0131 ,
		\EAX_reg[26]/NET0131 ,
		\EAX_reg[27]/NET0131 ,
		_w2093_,
		_w2624_
	);
	LUT4 #(
		.INIT('h0002)
	) name2172 (
		_w589_,
		_w566_,
		_w2095_,
		_w2624_,
		_w2625_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name2173 (
		\Datao[27]_pad ,
		_w594_,
		_w596_,
		_w2625_,
		_w2626_
	);
	LUT4 #(
		.INIT('h3f15)
	) name2174 (
		\Datao[27]_pad ,
		\uWord_reg[11]/NET0131 ,
		_w2179_,
		_w2180_,
		_w2627_
	);
	LUT3 #(
		.INIT('h2f)
	) name2175 (
		_w690_,
		_w2626_,
		_w2627_,
		_w2628_
	);
	LUT2 #(
		.INIT('h2)
	) name2176 (
		\EBX_reg[27]/NET0131 ,
		_w1841_,
		_w2629_
	);
	LUT4 #(
		.INIT('h0b03)
	) name2177 (
		\EBX_reg[26]/NET0131 ,
		_w622_,
		_w1992_,
		_w1986_,
		_w2630_
	);
	LUT2 #(
		.INIT('h8)
	) name2178 (
		_w1833_,
		_w1990_,
		_w2631_
	);
	LUT3 #(
		.INIT('h40)
	) name2179 (
		\EBX_reg[27]/NET0131 ,
		_w617_,
		_w621_,
		_w2632_
	);
	LUT4 #(
		.INIT('h070f)
	) name2180 (
		\EBX_reg[26]/NET0131 ,
		_w1986_,
		_w2631_,
		_w2632_,
		_w2633_
	);
	LUT4 #(
		.INIT('h08cc)
	) name2181 (
		\EBX_reg[27]/NET0131 ,
		_w690_,
		_w2630_,
		_w2633_,
		_w2634_
	);
	LUT2 #(
		.INIT('he)
	) name2182 (
		_w2629_,
		_w2634_,
		_w2635_
	);
	LUT2 #(
		.INIT('h2)
	) name2183 (
		\uWord_reg[11]/NET0131 ,
		_w1841_,
		_w2636_
	);
	LUT2 #(
		.INIT('h8)
	) name2184 (
		READY_n_pad,
		\uWord_reg[11]/NET0131 ,
		_w2637_
	);
	LUT2 #(
		.INIT('h1)
	) name2185 (
		_w1834_,
		_w2637_,
		_w2638_
	);
	LUT2 #(
		.INIT('h2)
	) name2186 (
		_w582_,
		_w2638_,
		_w2639_
	);
	LUT4 #(
		.INIT('haa02)
	) name2187 (
		\uWord_reg[11]/NET0131 ,
		_w582_,
		_w589_,
		_w566_,
		_w2640_
	);
	LUT4 #(
		.INIT('haaa8)
	) name2188 (
		_w690_,
		_w2625_,
		_w2639_,
		_w2640_,
		_w2641_
	);
	LUT2 #(
		.INIT('he)
	) name2189 (
		_w2636_,
		_w2641_,
		_w2642_
	);
	LUT4 #(
		.INIT('h3700)
	) name2190 (
		_w653_,
		_w690_,
		_w1742_,
		_w1841_,
		_w2643_
	);
	LUT4 #(
		.INIT('h2202)
	) name2191 (
		\Datai[7]_pad ,
		READY_n_pad,
		_w563_,
		_w565_,
		_w2644_
	);
	LUT4 #(
		.INIT('hf800)
	) name2192 (
		_w494_,
		_w586_,
		_w582_,
		_w2644_,
		_w2645_
	);
	LUT4 #(
		.INIT('h0080)
	) name2193 (
		_w602_,
		_w604_,
		_w634_,
		_w836_,
		_w2646_
	);
	LUT2 #(
		.INIT('h6)
	) name2194 (
		\EAX_reg[7]/NET0131 ,
		_w1744_,
		_w2647_
	);
	LUT3 #(
		.INIT('h80)
	) name2195 (
		_w518_,
		_w617_,
		_w2647_,
		_w2648_
	);
	LUT4 #(
		.INIT('haaa8)
	) name2196 (
		_w690_,
		_w2646_,
		_w2645_,
		_w2648_,
		_w2649_
	);
	LUT3 #(
		.INIT('hf2)
	) name2197 (
		\EAX_reg[7]/NET0131 ,
		_w2643_,
		_w2649_,
		_w2650_
	);
	LUT4 #(
		.INIT('h153f)
	) name2198 (
		\InstQueue_reg[3][0]/NET0131 ,
		\InstQueue_reg[9][0]/NET0131 ,
		_w470_,
		_w473_,
		_w2651_
	);
	LUT4 #(
		.INIT('h153f)
	) name2199 (
		\InstQueue_reg[10][0]/NET0131 ,
		\InstQueue_reg[15][0]/NET0131 ,
		_w461_,
		_w463_,
		_w2652_
	);
	LUT4 #(
		.INIT('h135f)
	) name2200 (
		\InstQueue_reg[0][0]/NET0131 ,
		\InstQueue_reg[11][0]/NET0131 ,
		_w476_,
		_w467_,
		_w2653_
	);
	LUT4 #(
		.INIT('h153f)
	) name2201 (
		\InstQueue_reg[5][0]/NET0131 ,
		\InstQueue_reg[6][0]/NET0131 ,
		_w468_,
		_w460_,
		_w2654_
	);
	LUT4 #(
		.INIT('h8000)
	) name2202 (
		_w2653_,
		_w2654_,
		_w2651_,
		_w2652_,
		_w2655_
	);
	LUT4 #(
		.INIT('h153f)
	) name2203 (
		\InstQueue_reg[2][0]/NET0131 ,
		\InstQueue_reg[4][0]/NET0131 ,
		_w474_,
		_w464_,
		_w2656_
	);
	LUT4 #(
		.INIT('h153f)
	) name2204 (
		\InstQueue_reg[1][0]/NET0131 ,
		\InstQueue_reg[8][0]/NET0131 ,
		_w453_,
		_w455_,
		_w2657_
	);
	LUT4 #(
		.INIT('h135f)
	) name2205 (
		\InstQueue_reg[14][0]/NET0131 ,
		\InstQueue_reg[7][0]/NET0131 ,
		_w477_,
		_w457_,
		_w2658_
	);
	LUT4 #(
		.INIT('h135f)
	) name2206 (
		\InstQueue_reg[12][0]/NET0131 ,
		\InstQueue_reg[13][0]/NET0131 ,
		_w471_,
		_w458_,
		_w2659_
	);
	LUT4 #(
		.INIT('h8000)
	) name2207 (
		_w2658_,
		_w2659_,
		_w2656_,
		_w2657_,
		_w2660_
	);
	LUT2 #(
		.INIT('h8)
	) name2208 (
		_w2655_,
		_w2660_,
		_w2661_
	);
	LUT4 #(
		.INIT('h0080)
	) name2209 (
		_w602_,
		_w604_,
		_w634_,
		_w2661_,
		_w2662_
	);
	LUT3 #(
		.INIT('h6c)
	) name2210 (
		\EAX_reg[7]/NET0131 ,
		\EAX_reg[8]/NET0131 ,
		_w1744_,
		_w2663_
	);
	LUT3 #(
		.INIT('h80)
	) name2211 (
		_w518_,
		_w617_,
		_w2663_,
		_w2664_
	);
	LUT4 #(
		.INIT('h0007)
	) name2212 (
		_w588_,
		_w2190_,
		_w2662_,
		_w2664_,
		_w2665_
	);
	LUT2 #(
		.INIT('h2)
	) name2213 (
		_w690_,
		_w2665_,
		_w2666_
	);
	LUT3 #(
		.INIT('hf2)
	) name2214 (
		\EAX_reg[8]/NET0131 ,
		_w2643_,
		_w2666_,
		_w2667_
	);
	LUT4 #(
		.INIT('h153f)
	) name2215 (
		\InstQueue_reg[3][1]/NET0131 ,
		\InstQueue_reg[9][1]/NET0131 ,
		_w470_,
		_w473_,
		_w2668_
	);
	LUT4 #(
		.INIT('h153f)
	) name2216 (
		\InstQueue_reg[5][1]/NET0131 ,
		\InstQueue_reg[6][1]/NET0131 ,
		_w468_,
		_w460_,
		_w2669_
	);
	LUT4 #(
		.INIT('h153f)
	) name2217 (
		\InstQueue_reg[11][1]/NET0131 ,
		\InstQueue_reg[8][1]/NET0131 ,
		_w453_,
		_w467_,
		_w2670_
	);
	LUT4 #(
		.INIT('h135f)
	) name2218 (
		\InstQueue_reg[0][1]/NET0131 ,
		\InstQueue_reg[1][1]/NET0131 ,
		_w476_,
		_w455_,
		_w2671_
	);
	LUT4 #(
		.INIT('h8000)
	) name2219 (
		_w2670_,
		_w2671_,
		_w2668_,
		_w2669_,
		_w2672_
	);
	LUT4 #(
		.INIT('h153f)
	) name2220 (
		\InstQueue_reg[12][1]/NET0131 ,
		\InstQueue_reg[4][1]/NET0131 ,
		_w474_,
		_w471_,
		_w2673_
	);
	LUT4 #(
		.INIT('h153f)
	) name2221 (
		\InstQueue_reg[14][1]/NET0131 ,
		\InstQueue_reg[15][1]/NET0131 ,
		_w461_,
		_w477_,
		_w2674_
	);
	LUT4 #(
		.INIT('h135f)
	) name2222 (
		\InstQueue_reg[2][1]/NET0131 ,
		\InstQueue_reg[7][1]/NET0131 ,
		_w464_,
		_w457_,
		_w2675_
	);
	LUT4 #(
		.INIT('h135f)
	) name2223 (
		\InstQueue_reg[10][1]/NET0131 ,
		\InstQueue_reg[13][1]/NET0131 ,
		_w463_,
		_w458_,
		_w2676_
	);
	LUT4 #(
		.INIT('h8000)
	) name2224 (
		_w2675_,
		_w2676_,
		_w2673_,
		_w2674_,
		_w2677_
	);
	LUT2 #(
		.INIT('h8)
	) name2225 (
		_w2672_,
		_w2677_,
		_w2678_
	);
	LUT4 #(
		.INIT('h0080)
	) name2226 (
		_w602_,
		_w604_,
		_w634_,
		_w2678_,
		_w2679_
	);
	LUT4 #(
		.INIT('hf800)
	) name2227 (
		_w494_,
		_w586_,
		_w582_,
		_w2455_,
		_w2680_
	);
	LUT4 #(
		.INIT('h78f0)
	) name2228 (
		\EAX_reg[7]/NET0131 ,
		\EAX_reg[8]/NET0131 ,
		\EAX_reg[9]/NET0131 ,
		_w1744_,
		_w2681_
	);
	LUT3 #(
		.INIT('h80)
	) name2229 (
		_w518_,
		_w617_,
		_w2681_,
		_w2682_
	);
	LUT4 #(
		.INIT('haaa8)
	) name2230 (
		_w690_,
		_w2680_,
		_w2679_,
		_w2682_,
		_w2683_
	);
	LUT3 #(
		.INIT('hf2)
	) name2231 (
		\EAX_reg[9]/NET0131 ,
		_w2643_,
		_w2683_,
		_w2684_
	);
	LUT2 #(
		.INIT('h2)
	) name2232 (
		\EAX_reg[10]/NET0131 ,
		_w1841_,
		_w2685_
	);
	LUT3 #(
		.INIT('h08)
	) name2233 (
		_w518_,
		_w617_,
		_w1746_,
		_w2686_
	);
	LUT4 #(
		.INIT('haaa8)
	) name2234 (
		\EAX_reg[10]/NET0131 ,
		_w653_,
		_w1742_,
		_w2686_,
		_w2687_
	);
	LUT3 #(
		.INIT('h20)
	) name2235 (
		\Datai[10]_pad ,
		READY_n_pad,
		_w588_,
		_w2688_
	);
	LUT4 #(
		.INIT('h4000)
	) name2236 (
		\EAX_reg[10]/NET0131 ,
		_w518_,
		_w617_,
		_w1745_,
		_w2689_
	);
	LUT4 #(
		.INIT('h135f)
	) name2237 (
		\InstQueue_reg[2][2]/NET0131 ,
		\InstQueue_reg[3][2]/NET0131 ,
		_w464_,
		_w473_,
		_w2690_
	);
	LUT4 #(
		.INIT('h153f)
	) name2238 (
		\InstQueue_reg[10][2]/NET0131 ,
		\InstQueue_reg[6][2]/NET0131 ,
		_w468_,
		_w463_,
		_w2691_
	);
	LUT4 #(
		.INIT('h135f)
	) name2239 (
		\InstQueue_reg[0][2]/NET0131 ,
		\InstQueue_reg[8][2]/NET0131 ,
		_w476_,
		_w453_,
		_w2692_
	);
	LUT4 #(
		.INIT('h135f)
	) name2240 (
		\InstQueue_reg[12][2]/NET0131 ,
		\InstQueue_reg[5][2]/NET0131 ,
		_w471_,
		_w460_,
		_w2693_
	);
	LUT4 #(
		.INIT('h8000)
	) name2241 (
		_w2692_,
		_w2693_,
		_w2690_,
		_w2691_,
		_w2694_
	);
	LUT4 #(
		.INIT('h153f)
	) name2242 (
		\InstQueue_reg[14][2]/NET0131 ,
		\InstQueue_reg[4][2]/NET0131 ,
		_w474_,
		_w477_,
		_w2695_
	);
	LUT4 #(
		.INIT('h153f)
	) name2243 (
		\InstQueue_reg[11][2]/NET0131 ,
		\InstQueue_reg[15][2]/NET0131 ,
		_w461_,
		_w467_,
		_w2696_
	);
	LUT4 #(
		.INIT('h153f)
	) name2244 (
		\InstQueue_reg[7][2]/NET0131 ,
		\InstQueue_reg[9][2]/NET0131 ,
		_w470_,
		_w457_,
		_w2697_
	);
	LUT4 #(
		.INIT('h135f)
	) name2245 (
		\InstQueue_reg[13][2]/NET0131 ,
		\InstQueue_reg[1][2]/NET0131 ,
		_w458_,
		_w455_,
		_w2698_
	);
	LUT4 #(
		.INIT('h8000)
	) name2246 (
		_w2697_,
		_w2698_,
		_w2695_,
		_w2696_,
		_w2699_
	);
	LUT2 #(
		.INIT('h8)
	) name2247 (
		_w2694_,
		_w2699_,
		_w2700_
	);
	LUT4 #(
		.INIT('h0080)
	) name2248 (
		_w602_,
		_w604_,
		_w634_,
		_w2700_,
		_w2701_
	);
	LUT2 #(
		.INIT('h1)
	) name2249 (
		_w2689_,
		_w2701_,
		_w2702_
	);
	LUT2 #(
		.INIT('h4)
	) name2250 (
		_w2688_,
		_w2702_,
		_w2703_
	);
	LUT4 #(
		.INIT('hecee)
	) name2251 (
		_w690_,
		_w2685_,
		_w2687_,
		_w2703_,
		_w2704_
	);
	LUT2 #(
		.INIT('h2)
	) name2252 (
		\EAX_reg[11]/NET0131 ,
		_w1841_,
		_w2705_
	);
	LUT4 #(
		.INIT('haaa8)
	) name2253 (
		\EAX_reg[11]/NET0131 ,
		_w653_,
		_w1742_,
		_w2686_,
		_w2706_
	);
	LUT3 #(
		.INIT('h20)
	) name2254 (
		\Datai[11]_pad ,
		READY_n_pad,
		_w588_,
		_w2707_
	);
	LUT4 #(
		.INIT('h135f)
	) name2255 (
		\InstQueue_reg[12][3]/NET0131 ,
		\InstQueue_reg[3][3]/NET0131 ,
		_w471_,
		_w473_,
		_w2708_
	);
	LUT4 #(
		.INIT('h153f)
	) name2256 (
		\InstQueue_reg[10][3]/NET0131 ,
		\InstQueue_reg[6][3]/NET0131 ,
		_w468_,
		_w463_,
		_w2709_
	);
	LUT4 #(
		.INIT('h135f)
	) name2257 (
		\InstQueue_reg[0][3]/NET0131 ,
		\InstQueue_reg[8][3]/NET0131 ,
		_w476_,
		_w453_,
		_w2710_
	);
	LUT4 #(
		.INIT('h135f)
	) name2258 (
		\InstQueue_reg[2][3]/NET0131 ,
		\InstQueue_reg[5][3]/NET0131 ,
		_w464_,
		_w460_,
		_w2711_
	);
	LUT4 #(
		.INIT('h8000)
	) name2259 (
		_w2710_,
		_w2711_,
		_w2708_,
		_w2709_,
		_w2712_
	);
	LUT4 #(
		.INIT('h153f)
	) name2260 (
		\InstQueue_reg[1][3]/NET0131 ,
		\InstQueue_reg[4][3]/NET0131 ,
		_w474_,
		_w455_,
		_w2713_
	);
	LUT4 #(
		.INIT('h153f)
	) name2261 (
		\InstQueue_reg[11][3]/NET0131 ,
		\InstQueue_reg[15][3]/NET0131 ,
		_w461_,
		_w467_,
		_w2714_
	);
	LUT4 #(
		.INIT('h153f)
	) name2262 (
		\InstQueue_reg[7][3]/NET0131 ,
		\InstQueue_reg[9][3]/NET0131 ,
		_w470_,
		_w457_,
		_w2715_
	);
	LUT4 #(
		.INIT('h153f)
	) name2263 (
		\InstQueue_reg[13][3]/NET0131 ,
		\InstQueue_reg[14][3]/NET0131 ,
		_w477_,
		_w458_,
		_w2716_
	);
	LUT4 #(
		.INIT('h8000)
	) name2264 (
		_w2715_,
		_w2716_,
		_w2713_,
		_w2714_,
		_w2717_
	);
	LUT2 #(
		.INIT('h8)
	) name2265 (
		_w2712_,
		_w2717_,
		_w2718_
	);
	LUT4 #(
		.INIT('h0080)
	) name2266 (
		_w602_,
		_w604_,
		_w634_,
		_w2718_,
		_w2719_
	);
	LUT3 #(
		.INIT('h20)
	) name2267 (
		\EAX_reg[10]/NET0131 ,
		\EAX_reg[11]/NET0131 ,
		_w1745_,
		_w2720_
	);
	LUT3 #(
		.INIT('h80)
	) name2268 (
		_w518_,
		_w617_,
		_w2720_,
		_w2721_
	);
	LUT2 #(
		.INIT('h1)
	) name2269 (
		_w2719_,
		_w2721_,
		_w2722_
	);
	LUT2 #(
		.INIT('h4)
	) name2270 (
		_w2707_,
		_w2722_,
		_w2723_
	);
	LUT4 #(
		.INIT('hecee)
	) name2271 (
		_w690_,
		_w2705_,
		_w2706_,
		_w2723_,
		_w2724_
	);
	LUT2 #(
		.INIT('h2)
	) name2272 (
		\EBX_reg[25]/NET0131 ,
		_w1841_,
		_w2725_
	);
	LUT4 #(
		.INIT('h8000)
	) name2273 (
		\EBX_reg[19]/NET0131 ,
		\EBX_reg[24]/NET0131 ,
		_w1982_,
		_w1983_,
		_w2726_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name2274 (
		\EBX_reg[25]/NET0131 ,
		_w622_,
		_w1992_,
		_w2726_,
		_w2727_
	);
	LUT4 #(
		.INIT('h8000)
	) name2275 (
		_w569_,
		_w602_,
		_w634_,
		_w2453_,
		_w2728_
	);
	LUT3 #(
		.INIT('h40)
	) name2276 (
		\EBX_reg[25]/NET0131 ,
		_w617_,
		_w621_,
		_w2729_
	);
	LUT3 #(
		.INIT('h15)
	) name2277 (
		_w2728_,
		_w2726_,
		_w2729_,
		_w2730_
	);
	LUT4 #(
		.INIT('hecee)
	) name2278 (
		_w690_,
		_w2725_,
		_w2727_,
		_w2730_,
		_w2731_
	);
	LUT2 #(
		.INIT('h2)
	) name2279 (
		\EAX_reg[12]/NET0131 ,
		_w1841_,
		_w2732_
	);
	LUT3 #(
		.INIT('h08)
	) name2280 (
		_w518_,
		_w617_,
		_w1747_,
		_w2733_
	);
	LUT4 #(
		.INIT('h88a8)
	) name2281 (
		\EAX_reg[12]/NET0131 ,
		READY_n_pad,
		_w563_,
		_w565_,
		_w2734_
	);
	LUT2 #(
		.INIT('h1)
	) name2282 (
		_w2099_,
		_w2734_,
		_w2735_
	);
	LUT4 #(
		.INIT('h00f8)
	) name2283 (
		_w494_,
		_w586_,
		_w582_,
		_w2735_,
		_w2736_
	);
	LUT4 #(
		.INIT('h4000)
	) name2284 (
		\EAX_reg[12]/NET0131 ,
		_w518_,
		_w617_,
		_w1747_,
		_w2737_
	);
	LUT4 #(
		.INIT('h135f)
	) name2285 (
		\InstQueue_reg[14][4]/NET0131 ,
		\InstQueue_reg[3][4]/NET0131 ,
		_w477_,
		_w473_,
		_w2738_
	);
	LUT4 #(
		.INIT('h135f)
	) name2286 (
		\InstQueue_reg[10][4]/NET0131 ,
		\InstQueue_reg[7][4]/NET0131 ,
		_w463_,
		_w457_,
		_w2739_
	);
	LUT4 #(
		.INIT('h135f)
	) name2287 (
		\InstQueue_reg[0][4]/NET0131 ,
		\InstQueue_reg[8][4]/NET0131 ,
		_w476_,
		_w453_,
		_w2740_
	);
	LUT4 #(
		.INIT('h153f)
	) name2288 (
		\InstQueue_reg[5][4]/NET0131 ,
		\InstQueue_reg[6][4]/NET0131 ,
		_w468_,
		_w460_,
		_w2741_
	);
	LUT4 #(
		.INIT('h8000)
	) name2289 (
		_w2740_,
		_w2741_,
		_w2738_,
		_w2739_,
		_w2742_
	);
	LUT4 #(
		.INIT('h153f)
	) name2290 (
		\InstQueue_reg[12][4]/NET0131 ,
		\InstQueue_reg[4][4]/NET0131 ,
		_w474_,
		_w471_,
		_w2743_
	);
	LUT4 #(
		.INIT('h153f)
	) name2291 (
		\InstQueue_reg[11][4]/NET0131 ,
		\InstQueue_reg[15][4]/NET0131 ,
		_w461_,
		_w467_,
		_w2744_
	);
	LUT4 #(
		.INIT('h153f)
	) name2292 (
		\InstQueue_reg[1][4]/NET0131 ,
		\InstQueue_reg[9][4]/NET0131 ,
		_w470_,
		_w455_,
		_w2745_
	);
	LUT4 #(
		.INIT('h153f)
	) name2293 (
		\InstQueue_reg[13][4]/NET0131 ,
		\InstQueue_reg[2][4]/NET0131 ,
		_w464_,
		_w458_,
		_w2746_
	);
	LUT4 #(
		.INIT('h8000)
	) name2294 (
		_w2745_,
		_w2746_,
		_w2743_,
		_w2744_,
		_w2747_
	);
	LUT2 #(
		.INIT('h8)
	) name2295 (
		_w2742_,
		_w2747_,
		_w2748_
	);
	LUT4 #(
		.INIT('h0080)
	) name2296 (
		_w602_,
		_w604_,
		_w634_,
		_w2748_,
		_w2749_
	);
	LUT3 #(
		.INIT('h01)
	) name2297 (
		_w2737_,
		_w2749_,
		_w2736_,
		_w2750_
	);
	LUT4 #(
		.INIT('h5700)
	) name2298 (
		\EAX_reg[12]/NET0131 ,
		_w1742_,
		_w2733_,
		_w2750_,
		_w2751_
	);
	LUT3 #(
		.INIT('hce)
	) name2299 (
		_w690_,
		_w2732_,
		_w2751_,
		_w2752_
	);
	LUT2 #(
		.INIT('h2)
	) name2300 (
		\EAX_reg[13]/NET0131 ,
		_w1841_,
		_w2753_
	);
	LUT3 #(
		.INIT('h08)
	) name2301 (
		_w518_,
		_w617_,
		_w1748_,
		_w2754_
	);
	LUT4 #(
		.INIT('haaa8)
	) name2302 (
		\EAX_reg[13]/NET0131 ,
		_w653_,
		_w1742_,
		_w2754_,
		_w2755_
	);
	LUT3 #(
		.INIT('h20)
	) name2303 (
		\Datai[13]_pad ,
		READY_n_pad,
		_w588_,
		_w2756_
	);
	LUT4 #(
		.INIT('h153f)
	) name2304 (
		\InstQueue_reg[2][5]/NET0131 ,
		\InstQueue_reg[4][5]/NET0131 ,
		_w474_,
		_w464_,
		_w2757_
	);
	LUT4 #(
		.INIT('h135f)
	) name2305 (
		\InstQueue_reg[6][5]/NET0131 ,
		\InstQueue_reg[8][5]/NET0131 ,
		_w468_,
		_w453_,
		_w2758_
	);
	LUT4 #(
		.INIT('h135f)
	) name2306 (
		\InstQueue_reg[0][5]/NET0131 ,
		\InstQueue_reg[11][5]/NET0131 ,
		_w476_,
		_w467_,
		_w2759_
	);
	LUT4 #(
		.INIT('h135f)
	) name2307 (
		\InstQueue_reg[15][5]/NET0131 ,
		\InstQueue_reg[5][5]/NET0131 ,
		_w461_,
		_w460_,
		_w2760_
	);
	LUT4 #(
		.INIT('h8000)
	) name2308 (
		_w2759_,
		_w2760_,
		_w2757_,
		_w2758_,
		_w2761_
	);
	LUT4 #(
		.INIT('h153f)
	) name2309 (
		\InstQueue_reg[1][5]/NET0131 ,
		\InstQueue_reg[3][5]/NET0131 ,
		_w473_,
		_w455_,
		_w2762_
	);
	LUT4 #(
		.INIT('h153f)
	) name2310 (
		\InstQueue_reg[12][5]/NET0131 ,
		\InstQueue_reg[9][5]/NET0131 ,
		_w470_,
		_w471_,
		_w2763_
	);
	LUT4 #(
		.INIT('h135f)
	) name2311 (
		\InstQueue_reg[14][5]/NET0131 ,
		\InstQueue_reg[7][5]/NET0131 ,
		_w477_,
		_w457_,
		_w2764_
	);
	LUT4 #(
		.INIT('h135f)
	) name2312 (
		\InstQueue_reg[10][5]/NET0131 ,
		\InstQueue_reg[13][5]/NET0131 ,
		_w463_,
		_w458_,
		_w2765_
	);
	LUT4 #(
		.INIT('h8000)
	) name2313 (
		_w2764_,
		_w2765_,
		_w2762_,
		_w2763_,
		_w2766_
	);
	LUT2 #(
		.INIT('h8)
	) name2314 (
		_w2761_,
		_w2766_,
		_w2767_
	);
	LUT4 #(
		.INIT('h0080)
	) name2315 (
		_w602_,
		_w604_,
		_w634_,
		_w2767_,
		_w2768_
	);
	LUT4 #(
		.INIT('h4000)
	) name2316 (
		\EAX_reg[13]/NET0131 ,
		_w518_,
		_w617_,
		_w1748_,
		_w2769_
	);
	LUT2 #(
		.INIT('h1)
	) name2317 (
		_w2768_,
		_w2769_,
		_w2770_
	);
	LUT2 #(
		.INIT('h4)
	) name2318 (
		_w2756_,
		_w2770_,
		_w2771_
	);
	LUT4 #(
		.INIT('hecee)
	) name2319 (
		_w690_,
		_w2753_,
		_w2755_,
		_w2771_,
		_w2772_
	);
	LUT3 #(
		.INIT('ha8)
	) name2320 (
		\EAX_reg[14]/NET0131 ,
		_w653_,
		_w1742_,
		_w2773_
	);
	LUT3 #(
		.INIT('h08)
	) name2321 (
		_w518_,
		_w617_,
		_w1750_,
		_w2774_
	);
	LUT4 #(
		.INIT('h4080)
	) name2322 (
		\EAX_reg[14]/NET0131 ,
		_w518_,
		_w617_,
		_w1749_,
		_w2775_
	);
	LUT4 #(
		.INIT('h135f)
	) name2323 (
		\InstQueue_reg[12][6]/NET0131 ,
		\InstQueue_reg[3][6]/NET0131 ,
		_w471_,
		_w473_,
		_w2776_
	);
	LUT4 #(
		.INIT('h153f)
	) name2324 (
		\InstQueue_reg[10][6]/NET0131 ,
		\InstQueue_reg[6][6]/NET0131 ,
		_w468_,
		_w463_,
		_w2777_
	);
	LUT4 #(
		.INIT('h135f)
	) name2325 (
		\InstQueue_reg[0][6]/NET0131 ,
		\InstQueue_reg[8][6]/NET0131 ,
		_w476_,
		_w453_,
		_w2778_
	);
	LUT4 #(
		.INIT('h135f)
	) name2326 (
		\InstQueue_reg[2][6]/NET0131 ,
		\InstQueue_reg[5][6]/NET0131 ,
		_w464_,
		_w460_,
		_w2779_
	);
	LUT4 #(
		.INIT('h8000)
	) name2327 (
		_w2778_,
		_w2779_,
		_w2776_,
		_w2777_,
		_w2780_
	);
	LUT4 #(
		.INIT('h153f)
	) name2328 (
		\InstQueue_reg[1][6]/NET0131 ,
		\InstQueue_reg[4][6]/NET0131 ,
		_w474_,
		_w455_,
		_w2781_
	);
	LUT4 #(
		.INIT('h153f)
	) name2329 (
		\InstQueue_reg[11][6]/NET0131 ,
		\InstQueue_reg[15][6]/NET0131 ,
		_w461_,
		_w467_,
		_w2782_
	);
	LUT4 #(
		.INIT('h153f)
	) name2330 (
		\InstQueue_reg[7][6]/NET0131 ,
		\InstQueue_reg[9][6]/NET0131 ,
		_w470_,
		_w457_,
		_w2783_
	);
	LUT4 #(
		.INIT('h153f)
	) name2331 (
		\InstQueue_reg[13][6]/NET0131 ,
		\InstQueue_reg[14][6]/NET0131 ,
		_w477_,
		_w458_,
		_w2784_
	);
	LUT4 #(
		.INIT('h8000)
	) name2332 (
		_w2783_,
		_w2784_,
		_w2781_,
		_w2782_,
		_w2785_
	);
	LUT2 #(
		.INIT('h8)
	) name2333 (
		_w2780_,
		_w2785_,
		_w2786_
	);
	LUT4 #(
		.INIT('h0080)
	) name2334 (
		_w602_,
		_w604_,
		_w634_,
		_w2786_,
		_w2787_
	);
	LUT4 #(
		.INIT('h00df)
	) name2335 (
		\Datai[14]_pad ,
		READY_n_pad,
		_w588_,
		_w2787_,
		_w2788_
	);
	LUT2 #(
		.INIT('h4)
	) name2336 (
		_w2775_,
		_w2788_,
		_w2789_
	);
	LUT2 #(
		.INIT('h2)
	) name2337 (
		\EAX_reg[14]/NET0131 ,
		_w1841_,
		_w2790_
	);
	LUT4 #(
		.INIT('hff8a)
	) name2338 (
		_w690_,
		_w2773_,
		_w2789_,
		_w2790_,
		_w2791_
	);
	LUT2 #(
		.INIT('h2)
	) name2339 (
		\EAX_reg[15]/NET0131 ,
		_w1841_,
		_w2792_
	);
	LUT4 #(
		.INIT('haaa8)
	) name2340 (
		\EAX_reg[15]/NET0131 ,
		_w653_,
		_w1742_,
		_w2774_,
		_w2793_
	);
	LUT4 #(
		.INIT('h4000)
	) name2341 (
		\EAX_reg[15]/NET0131 ,
		_w518_,
		_w617_,
		_w1750_,
		_w2794_
	);
	LUT4 #(
		.INIT('h2202)
	) name2342 (
		\Datai[15]_pad ,
		READY_n_pad,
		_w563_,
		_w565_,
		_w2795_
	);
	LUT4 #(
		.INIT('hf800)
	) name2343 (
		_w494_,
		_w586_,
		_w582_,
		_w2795_,
		_w2796_
	);
	LUT4 #(
		.INIT('h135f)
	) name2344 (
		\InstQueue_reg[12][7]/NET0131 ,
		\InstQueue_reg[3][7]/NET0131 ,
		_w471_,
		_w473_,
		_w2797_
	);
	LUT4 #(
		.INIT('h153f)
	) name2345 (
		\InstQueue_reg[10][7]/NET0131 ,
		\InstQueue_reg[6][7]/NET0131 ,
		_w468_,
		_w463_,
		_w2798_
	);
	LUT4 #(
		.INIT('h135f)
	) name2346 (
		\InstQueue_reg[0][7]/NET0131 ,
		\InstQueue_reg[8][7]/NET0131 ,
		_w476_,
		_w453_,
		_w2799_
	);
	LUT4 #(
		.INIT('h135f)
	) name2347 (
		\InstQueue_reg[2][7]/NET0131 ,
		\InstQueue_reg[5][7]/NET0131 ,
		_w464_,
		_w460_,
		_w2800_
	);
	LUT4 #(
		.INIT('h8000)
	) name2348 (
		_w2799_,
		_w2800_,
		_w2797_,
		_w2798_,
		_w2801_
	);
	LUT4 #(
		.INIT('h153f)
	) name2349 (
		\InstQueue_reg[1][7]/NET0131 ,
		\InstQueue_reg[4][7]/NET0131 ,
		_w474_,
		_w455_,
		_w2802_
	);
	LUT4 #(
		.INIT('h153f)
	) name2350 (
		\InstQueue_reg[11][7]/NET0131 ,
		\InstQueue_reg[15][7]/NET0131 ,
		_w461_,
		_w467_,
		_w2803_
	);
	LUT4 #(
		.INIT('h153f)
	) name2351 (
		\InstQueue_reg[7][7]/NET0131 ,
		\InstQueue_reg[9][7]/NET0131 ,
		_w470_,
		_w457_,
		_w2804_
	);
	LUT4 #(
		.INIT('h153f)
	) name2352 (
		\InstQueue_reg[13][7]/NET0131 ,
		\InstQueue_reg[14][7]/NET0131 ,
		_w477_,
		_w458_,
		_w2805_
	);
	LUT4 #(
		.INIT('h8000)
	) name2353 (
		_w2804_,
		_w2805_,
		_w2802_,
		_w2803_,
		_w2806_
	);
	LUT2 #(
		.INIT('h8)
	) name2354 (
		_w2801_,
		_w2806_,
		_w2807_
	);
	LUT4 #(
		.INIT('h0080)
	) name2355 (
		_w602_,
		_w604_,
		_w634_,
		_w2807_,
		_w2808_
	);
	LUT3 #(
		.INIT('h01)
	) name2356 (
		_w2796_,
		_w2808_,
		_w2794_,
		_w2809_
	);
	LUT4 #(
		.INIT('hecee)
	) name2357 (
		_w690_,
		_w2792_,
		_w2793_,
		_w2809_,
		_w2810_
	);
	LUT4 #(
		.INIT('h78f0)
	) name2358 (
		\Datai[25]_pad ,
		\Datai[26]_pad ,
		\Datai[27]_pad ,
		_w2208_,
		_w2811_
	);
	LUT4 #(
		.INIT('h6c00)
	) name2359 (
		\Datai[18]_pad ,
		\Datai[19]_pad ,
		_w2211_,
		_w2215_,
		_w2812_
	);
	LUT4 #(
		.INIT('haa80)
	) name2360 (
		\DataWidth_reg[1]/NET0131 ,
		_w2199_,
		_w2811_,
		_w2812_,
		_w2813_
	);
	LUT4 #(
		.INIT('h5553)
	) name2361 (
		\Datai[3]_pad ,
		\InstQueue_reg[0][3]/NET0131 ,
		_w2217_,
		_w2219_,
		_w2814_
	);
	LUT2 #(
		.INIT('h1)
	) name2362 (
		_w2223_,
		_w2814_,
		_w2815_
	);
	LUT4 #(
		.INIT('hc055)
	) name2363 (
		\InstQueue_reg[0][3]/NET0131 ,
		_w511_,
		_w516_,
		_w2217_,
		_w2816_
	);
	LUT2 #(
		.INIT('h2)
	) name2364 (
		\InstQueue_reg[0][3]/NET0131 ,
		_w2227_,
		_w2817_
	);
	LUT3 #(
		.INIT('h0d)
	) name2365 (
		_w1212_,
		_w2814_,
		_w2817_,
		_w2818_
	);
	LUT3 #(
		.INIT('hd0)
	) name2366 (
		_w710_,
		_w2816_,
		_w2818_,
		_w2819_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name2367 (
		_w695_,
		_w2813_,
		_w2815_,
		_w2819_,
		_w2820_
	);
	LUT4 #(
		.INIT('h78f0)
	) name2368 (
		\Datai[28]_pad ,
		\Datai[29]_pad ,
		\Datai[30]_pad ,
		_w2209_,
		_w2821_
	);
	LUT4 #(
		.INIT('h6c00)
	) name2369 (
		\Datai[21]_pad ,
		\Datai[22]_pad ,
		_w2212_,
		_w2215_,
		_w2822_
	);
	LUT4 #(
		.INIT('haa80)
	) name2370 (
		\DataWidth_reg[1]/NET0131 ,
		_w2199_,
		_w2821_,
		_w2822_,
		_w2823_
	);
	LUT4 #(
		.INIT('h5553)
	) name2371 (
		\Datai[6]_pad ,
		\InstQueue_reg[0][6]/NET0131 ,
		_w2217_,
		_w2219_,
		_w2824_
	);
	LUT2 #(
		.INIT('h1)
	) name2372 (
		_w2223_,
		_w2824_,
		_w2825_
	);
	LUT4 #(
		.INIT('hc055)
	) name2373 (
		\InstQueue_reg[0][6]/NET0131 ,
		_w523_,
		_w528_,
		_w2217_,
		_w2826_
	);
	LUT2 #(
		.INIT('h2)
	) name2374 (
		\InstQueue_reg[0][6]/NET0131 ,
		_w2227_,
		_w2827_
	);
	LUT3 #(
		.INIT('h0d)
	) name2375 (
		_w1212_,
		_w2824_,
		_w2827_,
		_w2828_
	);
	LUT3 #(
		.INIT('hd0)
	) name2376 (
		_w710_,
		_w2826_,
		_w2828_,
		_w2829_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name2377 (
		_w695_,
		_w2823_,
		_w2825_,
		_w2829_,
		_w2830_
	);
	LUT4 #(
		.INIT('h6c00)
	) name2378 (
		\Datai[18]_pad ,
		\Datai[19]_pad ,
		_w2211_,
		_w2234_,
		_w2831_
	);
	LUT4 #(
		.INIT('haa80)
	) name2379 (
		\DataWidth_reg[1]/NET0131 ,
		_w2232_,
		_w2811_,
		_w2831_,
		_w2832_
	);
	LUT4 #(
		.INIT('h5553)
	) name2380 (
		\Datai[3]_pad ,
		\InstQueue_reg[10][3]/NET0131 ,
		_w2236_,
		_w2237_,
		_w2833_
	);
	LUT2 #(
		.INIT('h1)
	) name2381 (
		_w2241_,
		_w2833_,
		_w2834_
	);
	LUT4 #(
		.INIT('hc055)
	) name2382 (
		\InstQueue_reg[10][3]/NET0131 ,
		_w511_,
		_w516_,
		_w2236_,
		_w2835_
	);
	LUT2 #(
		.INIT('h2)
	) name2383 (
		\InstQueue_reg[10][3]/NET0131 ,
		_w2227_,
		_w2836_
	);
	LUT3 #(
		.INIT('h0d)
	) name2384 (
		_w1212_,
		_w2833_,
		_w2836_,
		_w2837_
	);
	LUT3 #(
		.INIT('hd0)
	) name2385 (
		_w710_,
		_w2835_,
		_w2837_,
		_w2838_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name2386 (
		_w695_,
		_w2832_,
		_w2834_,
		_w2838_,
		_w2839_
	);
	LUT4 #(
		.INIT('h6c00)
	) name2387 (
		\Datai[21]_pad ,
		\Datai[22]_pad ,
		_w2212_,
		_w2234_,
		_w2840_
	);
	LUT4 #(
		.INIT('haa80)
	) name2388 (
		\DataWidth_reg[1]/NET0131 ,
		_w2232_,
		_w2821_,
		_w2840_,
		_w2841_
	);
	LUT4 #(
		.INIT('h5553)
	) name2389 (
		\Datai[6]_pad ,
		\InstQueue_reg[10][6]/NET0131 ,
		_w2236_,
		_w2237_,
		_w2842_
	);
	LUT2 #(
		.INIT('h1)
	) name2390 (
		_w2241_,
		_w2842_,
		_w2843_
	);
	LUT4 #(
		.INIT('hc055)
	) name2391 (
		\InstQueue_reg[10][6]/NET0131 ,
		_w523_,
		_w528_,
		_w2236_,
		_w2844_
	);
	LUT2 #(
		.INIT('h2)
	) name2392 (
		\InstQueue_reg[10][6]/NET0131 ,
		_w2227_,
		_w2845_
	);
	LUT3 #(
		.INIT('h0d)
	) name2393 (
		_w1212_,
		_w2842_,
		_w2845_,
		_w2846_
	);
	LUT3 #(
		.INIT('hd0)
	) name2394 (
		_w710_,
		_w2844_,
		_w2846_,
		_w2847_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name2395 (
		_w695_,
		_w2841_,
		_w2843_,
		_w2847_,
		_w2848_
	);
	LUT4 #(
		.INIT('h6c00)
	) name2396 (
		\Datai[18]_pad ,
		\Datai[19]_pad ,
		_w2211_,
		_w2237_,
		_w2849_
	);
	LUT4 #(
		.INIT('haa80)
	) name2397 (
		\DataWidth_reg[1]/NET0131 ,
		_w2234_,
		_w2811_,
		_w2849_,
		_w2850_
	);
	LUT4 #(
		.INIT('h5553)
	) name2398 (
		\Datai[3]_pad ,
		\InstQueue_reg[11][3]/NET0131 ,
		_w2236_,
		_w2251_,
		_w2851_
	);
	LUT2 #(
		.INIT('h1)
	) name2399 (
		_w2255_,
		_w2851_,
		_w2852_
	);
	LUT4 #(
		.INIT('hc055)
	) name2400 (
		\InstQueue_reg[11][3]/NET0131 ,
		_w511_,
		_w516_,
		_w2251_,
		_w2853_
	);
	LUT2 #(
		.INIT('h2)
	) name2401 (
		\InstQueue_reg[11][3]/NET0131 ,
		_w2227_,
		_w2854_
	);
	LUT3 #(
		.INIT('h0d)
	) name2402 (
		_w1212_,
		_w2851_,
		_w2854_,
		_w2855_
	);
	LUT3 #(
		.INIT('hd0)
	) name2403 (
		_w710_,
		_w2853_,
		_w2855_,
		_w2856_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name2404 (
		_w695_,
		_w2850_,
		_w2852_,
		_w2856_,
		_w2857_
	);
	LUT4 #(
		.INIT('h6c00)
	) name2405 (
		\Datai[21]_pad ,
		\Datai[22]_pad ,
		_w2212_,
		_w2237_,
		_w2858_
	);
	LUT4 #(
		.INIT('haa80)
	) name2406 (
		\DataWidth_reg[1]/NET0131 ,
		_w2234_,
		_w2821_,
		_w2858_,
		_w2859_
	);
	LUT4 #(
		.INIT('h5553)
	) name2407 (
		\Datai[6]_pad ,
		\InstQueue_reg[11][6]/NET0131 ,
		_w2236_,
		_w2251_,
		_w2860_
	);
	LUT2 #(
		.INIT('h1)
	) name2408 (
		_w2255_,
		_w2860_,
		_w2861_
	);
	LUT4 #(
		.INIT('hc055)
	) name2409 (
		\InstQueue_reg[11][6]/NET0131 ,
		_w523_,
		_w528_,
		_w2251_,
		_w2862_
	);
	LUT2 #(
		.INIT('h2)
	) name2410 (
		\InstQueue_reg[11][6]/NET0131 ,
		_w2227_,
		_w2863_
	);
	LUT3 #(
		.INIT('h0d)
	) name2411 (
		_w1212_,
		_w2860_,
		_w2863_,
		_w2864_
	);
	LUT3 #(
		.INIT('hd0)
	) name2412 (
		_w710_,
		_w2862_,
		_w2864_,
		_w2865_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name2413 (
		_w695_,
		_w2859_,
		_w2861_,
		_w2865_,
		_w2866_
	);
	LUT4 #(
		.INIT('h6c00)
	) name2414 (
		\Datai[18]_pad ,
		\Datai[19]_pad ,
		_w2211_,
		_w2236_,
		_w2867_
	);
	LUT4 #(
		.INIT('haa80)
	) name2415 (
		\DataWidth_reg[1]/NET0131 ,
		_w2237_,
		_w2811_,
		_w2867_,
		_w2868_
	);
	LUT4 #(
		.INIT('h5553)
	) name2416 (
		\Datai[3]_pad ,
		\InstQueue_reg[12][3]/NET0131 ,
		_w2251_,
		_w2265_,
		_w2869_
	);
	LUT2 #(
		.INIT('h1)
	) name2417 (
		_w2268_,
		_w2869_,
		_w2870_
	);
	LUT4 #(
		.INIT('hc055)
	) name2418 (
		\InstQueue_reg[12][3]/NET0131 ,
		_w511_,
		_w516_,
		_w2265_,
		_w2871_
	);
	LUT2 #(
		.INIT('h2)
	) name2419 (
		\InstQueue_reg[12][3]/NET0131 ,
		_w2227_,
		_w2872_
	);
	LUT3 #(
		.INIT('h0d)
	) name2420 (
		_w1212_,
		_w2869_,
		_w2872_,
		_w2873_
	);
	LUT3 #(
		.INIT('hd0)
	) name2421 (
		_w710_,
		_w2871_,
		_w2873_,
		_w2874_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name2422 (
		_w695_,
		_w2868_,
		_w2870_,
		_w2874_,
		_w2875_
	);
	LUT4 #(
		.INIT('h6c00)
	) name2423 (
		\Datai[21]_pad ,
		\Datai[22]_pad ,
		_w2212_,
		_w2236_,
		_w2876_
	);
	LUT4 #(
		.INIT('haa80)
	) name2424 (
		\DataWidth_reg[1]/NET0131 ,
		_w2237_,
		_w2821_,
		_w2876_,
		_w2877_
	);
	LUT4 #(
		.INIT('h5553)
	) name2425 (
		\Datai[6]_pad ,
		\InstQueue_reg[12][6]/NET0131 ,
		_w2251_,
		_w2265_,
		_w2878_
	);
	LUT2 #(
		.INIT('h1)
	) name2426 (
		_w2268_,
		_w2878_,
		_w2879_
	);
	LUT4 #(
		.INIT('hc055)
	) name2427 (
		\InstQueue_reg[12][6]/NET0131 ,
		_w523_,
		_w528_,
		_w2265_,
		_w2880_
	);
	LUT2 #(
		.INIT('h2)
	) name2428 (
		\InstQueue_reg[12][6]/NET0131 ,
		_w2227_,
		_w2881_
	);
	LUT3 #(
		.INIT('h0d)
	) name2429 (
		_w1212_,
		_w2878_,
		_w2881_,
		_w2882_
	);
	LUT3 #(
		.INIT('hd0)
	) name2430 (
		_w710_,
		_w2880_,
		_w2882_,
		_w2883_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name2431 (
		_w695_,
		_w2877_,
		_w2879_,
		_w2883_,
		_w2884_
	);
	LUT4 #(
		.INIT('h6c00)
	) name2432 (
		\Datai[18]_pad ,
		\Datai[19]_pad ,
		_w2211_,
		_w2251_,
		_w2885_
	);
	LUT4 #(
		.INIT('haa80)
	) name2433 (
		\DataWidth_reg[1]/NET0131 ,
		_w2236_,
		_w2811_,
		_w2885_,
		_w2886_
	);
	LUT4 #(
		.INIT('h5553)
	) name2434 (
		\Datai[3]_pad ,
		\InstQueue_reg[13][3]/NET0131 ,
		_w2199_,
		_w2265_,
		_w2887_
	);
	LUT2 #(
		.INIT('h1)
	) name2435 (
		_w2280_,
		_w2887_,
		_w2888_
	);
	LUT4 #(
		.INIT('hc055)
	) name2436 (
		\InstQueue_reg[13][3]/NET0131 ,
		_w511_,
		_w516_,
		_w2199_,
		_w2889_
	);
	LUT2 #(
		.INIT('h2)
	) name2437 (
		\InstQueue_reg[13][3]/NET0131 ,
		_w2227_,
		_w2890_
	);
	LUT3 #(
		.INIT('h0d)
	) name2438 (
		_w1212_,
		_w2887_,
		_w2890_,
		_w2891_
	);
	LUT3 #(
		.INIT('hd0)
	) name2439 (
		_w710_,
		_w2889_,
		_w2891_,
		_w2892_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name2440 (
		_w695_,
		_w2886_,
		_w2888_,
		_w2892_,
		_w2893_
	);
	LUT4 #(
		.INIT('h6c00)
	) name2441 (
		\Datai[21]_pad ,
		\Datai[22]_pad ,
		_w2212_,
		_w2251_,
		_w2894_
	);
	LUT4 #(
		.INIT('haa80)
	) name2442 (
		\DataWidth_reg[1]/NET0131 ,
		_w2236_,
		_w2821_,
		_w2894_,
		_w2895_
	);
	LUT4 #(
		.INIT('h5553)
	) name2443 (
		\Datai[6]_pad ,
		\InstQueue_reg[13][6]/NET0131 ,
		_w2199_,
		_w2265_,
		_w2896_
	);
	LUT2 #(
		.INIT('h1)
	) name2444 (
		_w2280_,
		_w2896_,
		_w2897_
	);
	LUT4 #(
		.INIT('hc055)
	) name2445 (
		\InstQueue_reg[13][6]/NET0131 ,
		_w523_,
		_w528_,
		_w2199_,
		_w2898_
	);
	LUT2 #(
		.INIT('h2)
	) name2446 (
		\InstQueue_reg[13][6]/NET0131 ,
		_w2227_,
		_w2899_
	);
	LUT3 #(
		.INIT('h0d)
	) name2447 (
		_w1212_,
		_w2896_,
		_w2899_,
		_w2900_
	);
	LUT3 #(
		.INIT('hd0)
	) name2448 (
		_w710_,
		_w2898_,
		_w2900_,
		_w2901_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name2449 (
		_w695_,
		_w2895_,
		_w2897_,
		_w2901_,
		_w2902_
	);
	LUT4 #(
		.INIT('h6c00)
	) name2450 (
		\Datai[18]_pad ,
		\Datai[19]_pad ,
		_w2211_,
		_w2265_,
		_w2903_
	);
	LUT4 #(
		.INIT('haa80)
	) name2451 (
		\DataWidth_reg[1]/NET0131 ,
		_w2251_,
		_w2811_,
		_w2903_,
		_w2904_
	);
	LUT4 #(
		.INIT('h5553)
	) name2452 (
		\Datai[3]_pad ,
		\InstQueue_reg[14][3]/NET0131 ,
		_w2199_,
		_w2215_,
		_w2905_
	);
	LUT2 #(
		.INIT('h1)
	) name2453 (
		_w2291_,
		_w2905_,
		_w2906_
	);
	LUT4 #(
		.INIT('hc055)
	) name2454 (
		\InstQueue_reg[14][3]/NET0131 ,
		_w511_,
		_w516_,
		_w2215_,
		_w2907_
	);
	LUT2 #(
		.INIT('h2)
	) name2455 (
		\InstQueue_reg[14][3]/NET0131 ,
		_w2227_,
		_w2908_
	);
	LUT3 #(
		.INIT('h0d)
	) name2456 (
		_w1212_,
		_w2905_,
		_w2908_,
		_w2909_
	);
	LUT3 #(
		.INIT('hd0)
	) name2457 (
		_w710_,
		_w2907_,
		_w2909_,
		_w2910_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name2458 (
		_w695_,
		_w2904_,
		_w2906_,
		_w2910_,
		_w2911_
	);
	LUT4 #(
		.INIT('h6c00)
	) name2459 (
		\Datai[21]_pad ,
		\Datai[22]_pad ,
		_w2212_,
		_w2265_,
		_w2912_
	);
	LUT4 #(
		.INIT('haa80)
	) name2460 (
		\DataWidth_reg[1]/NET0131 ,
		_w2251_,
		_w2821_,
		_w2912_,
		_w2913_
	);
	LUT4 #(
		.INIT('h5553)
	) name2461 (
		\Datai[6]_pad ,
		\InstQueue_reg[14][6]/NET0131 ,
		_w2199_,
		_w2215_,
		_w2914_
	);
	LUT2 #(
		.INIT('h1)
	) name2462 (
		_w2291_,
		_w2914_,
		_w2915_
	);
	LUT4 #(
		.INIT('hc055)
	) name2463 (
		\InstQueue_reg[14][6]/NET0131 ,
		_w523_,
		_w528_,
		_w2215_,
		_w2916_
	);
	LUT2 #(
		.INIT('h2)
	) name2464 (
		\InstQueue_reg[14][6]/NET0131 ,
		_w2227_,
		_w2917_
	);
	LUT3 #(
		.INIT('h0d)
	) name2465 (
		_w1212_,
		_w2914_,
		_w2917_,
		_w2918_
	);
	LUT3 #(
		.INIT('hd0)
	) name2466 (
		_w710_,
		_w2916_,
		_w2918_,
		_w2919_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name2467 (
		_w695_,
		_w2913_,
		_w2915_,
		_w2919_,
		_w2920_
	);
	LUT4 #(
		.INIT('h60c0)
	) name2468 (
		\Datai[18]_pad ,
		\Datai[19]_pad ,
		_w2199_,
		_w2211_,
		_w2921_
	);
	LUT4 #(
		.INIT('haa80)
	) name2469 (
		\DataWidth_reg[1]/NET0131 ,
		_w2265_,
		_w2811_,
		_w2921_,
		_w2922_
	);
	LUT4 #(
		.INIT('h5553)
	) name2470 (
		\Datai[3]_pad ,
		\InstQueue_reg[15][3]/NET0131 ,
		_w2219_,
		_w2215_,
		_w2923_
	);
	LUT2 #(
		.INIT('h1)
	) name2471 (
		_w2303_,
		_w2923_,
		_w2924_
	);
	LUT4 #(
		.INIT('hc055)
	) name2472 (
		\InstQueue_reg[15][3]/NET0131 ,
		_w511_,
		_w516_,
		_w2219_,
		_w2925_
	);
	LUT2 #(
		.INIT('h2)
	) name2473 (
		\InstQueue_reg[15][3]/NET0131 ,
		_w2227_,
		_w2926_
	);
	LUT3 #(
		.INIT('h0d)
	) name2474 (
		_w1212_,
		_w2923_,
		_w2926_,
		_w2927_
	);
	LUT3 #(
		.INIT('hd0)
	) name2475 (
		_w710_,
		_w2925_,
		_w2927_,
		_w2928_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name2476 (
		_w695_,
		_w2922_,
		_w2924_,
		_w2928_,
		_w2929_
	);
	LUT4 #(
		.INIT('h60c0)
	) name2477 (
		\Datai[21]_pad ,
		\Datai[22]_pad ,
		_w2199_,
		_w2212_,
		_w2930_
	);
	LUT4 #(
		.INIT('haa80)
	) name2478 (
		\DataWidth_reg[1]/NET0131 ,
		_w2265_,
		_w2821_,
		_w2930_,
		_w2931_
	);
	LUT4 #(
		.INIT('h5553)
	) name2479 (
		\Datai[6]_pad ,
		\InstQueue_reg[15][6]/NET0131 ,
		_w2219_,
		_w2215_,
		_w2932_
	);
	LUT2 #(
		.INIT('h1)
	) name2480 (
		_w2303_,
		_w2932_,
		_w2933_
	);
	LUT4 #(
		.INIT('hc055)
	) name2481 (
		\InstQueue_reg[15][6]/NET0131 ,
		_w523_,
		_w528_,
		_w2219_,
		_w2934_
	);
	LUT2 #(
		.INIT('h2)
	) name2482 (
		\InstQueue_reg[15][6]/NET0131 ,
		_w2227_,
		_w2935_
	);
	LUT3 #(
		.INIT('h0d)
	) name2483 (
		_w1212_,
		_w2932_,
		_w2935_,
		_w2936_
	);
	LUT3 #(
		.INIT('hd0)
	) name2484 (
		_w710_,
		_w2934_,
		_w2936_,
		_w2937_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name2485 (
		_w695_,
		_w2931_,
		_w2933_,
		_w2937_,
		_w2938_
	);
	LUT4 #(
		.INIT('h60c0)
	) name2486 (
		\Datai[18]_pad ,
		\Datai[19]_pad ,
		_w2219_,
		_w2211_,
		_w2939_
	);
	LUT4 #(
		.INIT('haa80)
	) name2487 (
		\DataWidth_reg[1]/NET0131 ,
		_w2215_,
		_w2811_,
		_w2939_,
		_w2940_
	);
	LUT4 #(
		.INIT('h5553)
	) name2488 (
		\Datai[3]_pad ,
		\InstQueue_reg[1][3]/NET0131 ,
		_w2217_,
		_w2313_,
		_w2941_
	);
	LUT2 #(
		.INIT('h1)
	) name2489 (
		_w2316_,
		_w2941_,
		_w2942_
	);
	LUT4 #(
		.INIT('hc055)
	) name2490 (
		\InstQueue_reg[1][3]/NET0131 ,
		_w511_,
		_w516_,
		_w2313_,
		_w2943_
	);
	LUT2 #(
		.INIT('h2)
	) name2491 (
		\InstQueue_reg[1][3]/NET0131 ,
		_w2227_,
		_w2944_
	);
	LUT3 #(
		.INIT('h0d)
	) name2492 (
		_w1212_,
		_w2941_,
		_w2944_,
		_w2945_
	);
	LUT3 #(
		.INIT('hd0)
	) name2493 (
		_w710_,
		_w2943_,
		_w2945_,
		_w2946_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name2494 (
		_w695_,
		_w2940_,
		_w2942_,
		_w2946_,
		_w2947_
	);
	LUT4 #(
		.INIT('h60c0)
	) name2495 (
		\Datai[21]_pad ,
		\Datai[22]_pad ,
		_w2219_,
		_w2212_,
		_w2948_
	);
	LUT4 #(
		.INIT('haa80)
	) name2496 (
		\DataWidth_reg[1]/NET0131 ,
		_w2215_,
		_w2821_,
		_w2948_,
		_w2949_
	);
	LUT4 #(
		.INIT('h5553)
	) name2497 (
		\Datai[6]_pad ,
		\InstQueue_reg[1][6]/NET0131 ,
		_w2217_,
		_w2313_,
		_w2950_
	);
	LUT2 #(
		.INIT('h1)
	) name2498 (
		_w2316_,
		_w2950_,
		_w2951_
	);
	LUT4 #(
		.INIT('hc055)
	) name2499 (
		\InstQueue_reg[1][6]/NET0131 ,
		_w523_,
		_w528_,
		_w2313_,
		_w2952_
	);
	LUT2 #(
		.INIT('h2)
	) name2500 (
		\InstQueue_reg[1][6]/NET0131 ,
		_w2227_,
		_w2953_
	);
	LUT3 #(
		.INIT('h0d)
	) name2501 (
		_w1212_,
		_w2950_,
		_w2953_,
		_w2954_
	);
	LUT3 #(
		.INIT('hd0)
	) name2502 (
		_w710_,
		_w2952_,
		_w2954_,
		_w2955_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name2503 (
		_w695_,
		_w2949_,
		_w2951_,
		_w2955_,
		_w2956_
	);
	LUT4 #(
		.INIT('h60c0)
	) name2504 (
		\Datai[18]_pad ,
		\Datai[19]_pad ,
		_w2217_,
		_w2211_,
		_w2957_
	);
	LUT4 #(
		.INIT('haa80)
	) name2505 (
		\DataWidth_reg[1]/NET0131 ,
		_w2219_,
		_w2811_,
		_w2957_,
		_w2958_
	);
	LUT4 #(
		.INIT('h5553)
	) name2506 (
		\Datai[3]_pad ,
		\InstQueue_reg[2][3]/NET0131 ,
		_w2313_,
		_w2326_,
		_w2959_
	);
	LUT2 #(
		.INIT('h1)
	) name2507 (
		_w2329_,
		_w2959_,
		_w2960_
	);
	LUT4 #(
		.INIT('hc055)
	) name2508 (
		\InstQueue_reg[2][3]/NET0131 ,
		_w511_,
		_w516_,
		_w2326_,
		_w2961_
	);
	LUT2 #(
		.INIT('h2)
	) name2509 (
		\InstQueue_reg[2][3]/NET0131 ,
		_w2227_,
		_w2962_
	);
	LUT3 #(
		.INIT('h0d)
	) name2510 (
		_w1212_,
		_w2959_,
		_w2962_,
		_w2963_
	);
	LUT3 #(
		.INIT('hd0)
	) name2511 (
		_w710_,
		_w2961_,
		_w2963_,
		_w2964_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name2512 (
		_w695_,
		_w2958_,
		_w2960_,
		_w2964_,
		_w2965_
	);
	LUT4 #(
		.INIT('h60c0)
	) name2513 (
		\Datai[21]_pad ,
		\Datai[22]_pad ,
		_w2217_,
		_w2212_,
		_w2966_
	);
	LUT4 #(
		.INIT('haa80)
	) name2514 (
		\DataWidth_reg[1]/NET0131 ,
		_w2219_,
		_w2821_,
		_w2966_,
		_w2967_
	);
	LUT4 #(
		.INIT('h5553)
	) name2515 (
		\Datai[6]_pad ,
		\InstQueue_reg[2][6]/NET0131 ,
		_w2313_,
		_w2326_,
		_w2968_
	);
	LUT2 #(
		.INIT('h1)
	) name2516 (
		_w2329_,
		_w2968_,
		_w2969_
	);
	LUT4 #(
		.INIT('hc055)
	) name2517 (
		\InstQueue_reg[2][6]/NET0131 ,
		_w523_,
		_w528_,
		_w2326_,
		_w2970_
	);
	LUT2 #(
		.INIT('h2)
	) name2518 (
		\InstQueue_reg[2][6]/NET0131 ,
		_w2227_,
		_w2971_
	);
	LUT3 #(
		.INIT('h0d)
	) name2519 (
		_w1212_,
		_w2968_,
		_w2971_,
		_w2972_
	);
	LUT3 #(
		.INIT('hd0)
	) name2520 (
		_w710_,
		_w2970_,
		_w2972_,
		_w2973_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name2521 (
		_w695_,
		_w2967_,
		_w2969_,
		_w2973_,
		_w2974_
	);
	LUT4 #(
		.INIT('h6c00)
	) name2522 (
		\Datai[18]_pad ,
		\Datai[19]_pad ,
		_w2211_,
		_w2313_,
		_w2975_
	);
	LUT4 #(
		.INIT('haa80)
	) name2523 (
		\DataWidth_reg[1]/NET0131 ,
		_w2217_,
		_w2811_,
		_w2975_,
		_w2976_
	);
	LUT4 #(
		.INIT('h5553)
	) name2524 (
		\Datai[3]_pad ,
		\InstQueue_reg[3][3]/NET0131 ,
		_w2326_,
		_w2339_,
		_w2977_
	);
	LUT2 #(
		.INIT('h1)
	) name2525 (
		_w2342_,
		_w2977_,
		_w2978_
	);
	LUT4 #(
		.INIT('hc055)
	) name2526 (
		\InstQueue_reg[3][3]/NET0131 ,
		_w511_,
		_w516_,
		_w2339_,
		_w2979_
	);
	LUT2 #(
		.INIT('h2)
	) name2527 (
		\InstQueue_reg[3][3]/NET0131 ,
		_w2227_,
		_w2980_
	);
	LUT3 #(
		.INIT('h0d)
	) name2528 (
		_w1212_,
		_w2977_,
		_w2980_,
		_w2981_
	);
	LUT3 #(
		.INIT('hd0)
	) name2529 (
		_w710_,
		_w2979_,
		_w2981_,
		_w2982_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name2530 (
		_w695_,
		_w2976_,
		_w2978_,
		_w2982_,
		_w2983_
	);
	LUT4 #(
		.INIT('h6c00)
	) name2531 (
		\Datai[21]_pad ,
		\Datai[22]_pad ,
		_w2212_,
		_w2313_,
		_w2984_
	);
	LUT4 #(
		.INIT('haa80)
	) name2532 (
		\DataWidth_reg[1]/NET0131 ,
		_w2217_,
		_w2821_,
		_w2984_,
		_w2985_
	);
	LUT4 #(
		.INIT('h5553)
	) name2533 (
		\Datai[6]_pad ,
		\InstQueue_reg[3][6]/NET0131 ,
		_w2326_,
		_w2339_,
		_w2986_
	);
	LUT2 #(
		.INIT('h1)
	) name2534 (
		_w2342_,
		_w2986_,
		_w2987_
	);
	LUT4 #(
		.INIT('hc055)
	) name2535 (
		\InstQueue_reg[3][6]/NET0131 ,
		_w523_,
		_w528_,
		_w2339_,
		_w2988_
	);
	LUT2 #(
		.INIT('h2)
	) name2536 (
		\InstQueue_reg[3][6]/NET0131 ,
		_w2227_,
		_w2989_
	);
	LUT3 #(
		.INIT('h0d)
	) name2537 (
		_w1212_,
		_w2986_,
		_w2989_,
		_w2990_
	);
	LUT3 #(
		.INIT('hd0)
	) name2538 (
		_w710_,
		_w2988_,
		_w2990_,
		_w2991_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name2539 (
		_w695_,
		_w2985_,
		_w2987_,
		_w2991_,
		_w2992_
	);
	LUT4 #(
		.INIT('h6c00)
	) name2540 (
		\Datai[18]_pad ,
		\Datai[19]_pad ,
		_w2211_,
		_w2326_,
		_w2993_
	);
	LUT4 #(
		.INIT('haa80)
	) name2541 (
		\DataWidth_reg[1]/NET0131 ,
		_w2313_,
		_w2811_,
		_w2993_,
		_w2994_
	);
	LUT4 #(
		.INIT('h5553)
	) name2542 (
		\Datai[3]_pad ,
		\InstQueue_reg[4][3]/NET0131 ,
		_w2339_,
		_w2352_,
		_w2995_
	);
	LUT2 #(
		.INIT('h1)
	) name2543 (
		_w2355_,
		_w2995_,
		_w2996_
	);
	LUT4 #(
		.INIT('hc055)
	) name2544 (
		\InstQueue_reg[4][3]/NET0131 ,
		_w511_,
		_w516_,
		_w2352_,
		_w2997_
	);
	LUT2 #(
		.INIT('h2)
	) name2545 (
		\InstQueue_reg[4][3]/NET0131 ,
		_w2227_,
		_w2998_
	);
	LUT3 #(
		.INIT('h0d)
	) name2546 (
		_w1212_,
		_w2995_,
		_w2998_,
		_w2999_
	);
	LUT3 #(
		.INIT('hd0)
	) name2547 (
		_w710_,
		_w2997_,
		_w2999_,
		_w3000_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name2548 (
		_w695_,
		_w2994_,
		_w2996_,
		_w3000_,
		_w3001_
	);
	LUT4 #(
		.INIT('h6c00)
	) name2549 (
		\Datai[21]_pad ,
		\Datai[22]_pad ,
		_w2212_,
		_w2326_,
		_w3002_
	);
	LUT4 #(
		.INIT('haa80)
	) name2550 (
		\DataWidth_reg[1]/NET0131 ,
		_w2313_,
		_w2821_,
		_w3002_,
		_w3003_
	);
	LUT4 #(
		.INIT('h5553)
	) name2551 (
		\Datai[6]_pad ,
		\InstQueue_reg[4][6]/NET0131 ,
		_w2339_,
		_w2352_,
		_w3004_
	);
	LUT2 #(
		.INIT('h1)
	) name2552 (
		_w2355_,
		_w3004_,
		_w3005_
	);
	LUT4 #(
		.INIT('hc055)
	) name2553 (
		\InstQueue_reg[4][6]/NET0131 ,
		_w523_,
		_w528_,
		_w2352_,
		_w3006_
	);
	LUT2 #(
		.INIT('h2)
	) name2554 (
		\InstQueue_reg[4][6]/NET0131 ,
		_w2227_,
		_w3007_
	);
	LUT3 #(
		.INIT('h0d)
	) name2555 (
		_w1212_,
		_w3004_,
		_w3007_,
		_w3008_
	);
	LUT3 #(
		.INIT('hd0)
	) name2556 (
		_w710_,
		_w3006_,
		_w3008_,
		_w3009_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name2557 (
		_w695_,
		_w3003_,
		_w3005_,
		_w3009_,
		_w3010_
	);
	LUT4 #(
		.INIT('h6c00)
	) name2558 (
		\Datai[18]_pad ,
		\Datai[19]_pad ,
		_w2211_,
		_w2339_,
		_w3011_
	);
	LUT4 #(
		.INIT('haa80)
	) name2559 (
		\DataWidth_reg[1]/NET0131 ,
		_w2326_,
		_w2811_,
		_w3011_,
		_w3012_
	);
	LUT4 #(
		.INIT('h5553)
	) name2560 (
		\Datai[3]_pad ,
		\InstQueue_reg[5][3]/NET0131 ,
		_w2352_,
		_w2365_,
		_w3013_
	);
	LUT2 #(
		.INIT('h1)
	) name2561 (
		_w2368_,
		_w3013_,
		_w3014_
	);
	LUT4 #(
		.INIT('hc055)
	) name2562 (
		\InstQueue_reg[5][3]/NET0131 ,
		_w511_,
		_w516_,
		_w2365_,
		_w3015_
	);
	LUT2 #(
		.INIT('h2)
	) name2563 (
		\InstQueue_reg[5][3]/NET0131 ,
		_w2227_,
		_w3016_
	);
	LUT3 #(
		.INIT('h0d)
	) name2564 (
		_w1212_,
		_w3013_,
		_w3016_,
		_w3017_
	);
	LUT3 #(
		.INIT('hd0)
	) name2565 (
		_w710_,
		_w3015_,
		_w3017_,
		_w3018_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name2566 (
		_w695_,
		_w3012_,
		_w3014_,
		_w3018_,
		_w3019_
	);
	LUT4 #(
		.INIT('h6c00)
	) name2567 (
		\Datai[21]_pad ,
		\Datai[22]_pad ,
		_w2212_,
		_w2339_,
		_w3020_
	);
	LUT4 #(
		.INIT('haa80)
	) name2568 (
		\DataWidth_reg[1]/NET0131 ,
		_w2326_,
		_w2821_,
		_w3020_,
		_w3021_
	);
	LUT4 #(
		.INIT('h5553)
	) name2569 (
		\Datai[6]_pad ,
		\InstQueue_reg[5][6]/NET0131 ,
		_w2352_,
		_w2365_,
		_w3022_
	);
	LUT2 #(
		.INIT('h1)
	) name2570 (
		_w2368_,
		_w3022_,
		_w3023_
	);
	LUT4 #(
		.INIT('hc055)
	) name2571 (
		\InstQueue_reg[5][6]/NET0131 ,
		_w523_,
		_w528_,
		_w2365_,
		_w3024_
	);
	LUT2 #(
		.INIT('h2)
	) name2572 (
		\InstQueue_reg[5][6]/NET0131 ,
		_w2227_,
		_w3025_
	);
	LUT3 #(
		.INIT('h0d)
	) name2573 (
		_w1212_,
		_w3022_,
		_w3025_,
		_w3026_
	);
	LUT3 #(
		.INIT('hd0)
	) name2574 (
		_w710_,
		_w3024_,
		_w3026_,
		_w3027_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name2575 (
		_w695_,
		_w3021_,
		_w3023_,
		_w3027_,
		_w3028_
	);
	LUT4 #(
		.INIT('h6c00)
	) name2576 (
		\Datai[18]_pad ,
		\Datai[19]_pad ,
		_w2211_,
		_w2352_,
		_w3029_
	);
	LUT4 #(
		.INIT('haa80)
	) name2577 (
		\DataWidth_reg[1]/NET0131 ,
		_w2339_,
		_w2811_,
		_w3029_,
		_w3030_
	);
	LUT4 #(
		.INIT('h5553)
	) name2578 (
		\Datai[3]_pad ,
		\InstQueue_reg[6][3]/NET0131 ,
		_w2365_,
		_w2378_,
		_w3031_
	);
	LUT2 #(
		.INIT('h1)
	) name2579 (
		_w2381_,
		_w3031_,
		_w3032_
	);
	LUT4 #(
		.INIT('hc055)
	) name2580 (
		\InstQueue_reg[6][3]/NET0131 ,
		_w511_,
		_w516_,
		_w2378_,
		_w3033_
	);
	LUT2 #(
		.INIT('h2)
	) name2581 (
		\InstQueue_reg[6][3]/NET0131 ,
		_w2227_,
		_w3034_
	);
	LUT3 #(
		.INIT('h0d)
	) name2582 (
		_w1212_,
		_w3031_,
		_w3034_,
		_w3035_
	);
	LUT3 #(
		.INIT('hd0)
	) name2583 (
		_w710_,
		_w3033_,
		_w3035_,
		_w3036_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name2584 (
		_w695_,
		_w3030_,
		_w3032_,
		_w3036_,
		_w3037_
	);
	LUT4 #(
		.INIT('h6c00)
	) name2585 (
		\Datai[21]_pad ,
		\Datai[22]_pad ,
		_w2212_,
		_w2352_,
		_w3038_
	);
	LUT4 #(
		.INIT('haa80)
	) name2586 (
		\DataWidth_reg[1]/NET0131 ,
		_w2339_,
		_w2821_,
		_w3038_,
		_w3039_
	);
	LUT4 #(
		.INIT('h5553)
	) name2587 (
		\Datai[6]_pad ,
		\InstQueue_reg[6][6]/NET0131 ,
		_w2365_,
		_w2378_,
		_w3040_
	);
	LUT2 #(
		.INIT('h1)
	) name2588 (
		_w2381_,
		_w3040_,
		_w3041_
	);
	LUT4 #(
		.INIT('hc055)
	) name2589 (
		\InstQueue_reg[6][6]/NET0131 ,
		_w523_,
		_w528_,
		_w2378_,
		_w3042_
	);
	LUT2 #(
		.INIT('h2)
	) name2590 (
		\InstQueue_reg[6][6]/NET0131 ,
		_w2227_,
		_w3043_
	);
	LUT3 #(
		.INIT('h0d)
	) name2591 (
		_w1212_,
		_w3040_,
		_w3043_,
		_w3044_
	);
	LUT3 #(
		.INIT('hd0)
	) name2592 (
		_w710_,
		_w3042_,
		_w3044_,
		_w3045_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name2593 (
		_w695_,
		_w3039_,
		_w3041_,
		_w3045_,
		_w3046_
	);
	LUT4 #(
		.INIT('h6c00)
	) name2594 (
		\Datai[18]_pad ,
		\Datai[19]_pad ,
		_w2211_,
		_w2365_,
		_w3047_
	);
	LUT4 #(
		.INIT('haa80)
	) name2595 (
		\DataWidth_reg[1]/NET0131 ,
		_w2352_,
		_w2811_,
		_w3047_,
		_w3048_
	);
	LUT4 #(
		.INIT('h5553)
	) name2596 (
		\Datai[3]_pad ,
		\InstQueue_reg[7][3]/NET0131 ,
		_w2232_,
		_w2378_,
		_w3049_
	);
	LUT2 #(
		.INIT('h1)
	) name2597 (
		_w2393_,
		_w3049_,
		_w3050_
	);
	LUT4 #(
		.INIT('hc055)
	) name2598 (
		\InstQueue_reg[7][3]/NET0131 ,
		_w511_,
		_w516_,
		_w2232_,
		_w3051_
	);
	LUT2 #(
		.INIT('h2)
	) name2599 (
		\InstQueue_reg[7][3]/NET0131 ,
		_w2227_,
		_w3052_
	);
	LUT3 #(
		.INIT('h0d)
	) name2600 (
		_w1212_,
		_w3049_,
		_w3052_,
		_w3053_
	);
	LUT3 #(
		.INIT('hd0)
	) name2601 (
		_w710_,
		_w3051_,
		_w3053_,
		_w3054_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name2602 (
		_w695_,
		_w3048_,
		_w3050_,
		_w3054_,
		_w3055_
	);
	LUT4 #(
		.INIT('h6c00)
	) name2603 (
		\Datai[21]_pad ,
		\Datai[22]_pad ,
		_w2212_,
		_w2365_,
		_w3056_
	);
	LUT4 #(
		.INIT('haa80)
	) name2604 (
		\DataWidth_reg[1]/NET0131 ,
		_w2352_,
		_w2821_,
		_w3056_,
		_w3057_
	);
	LUT4 #(
		.INIT('h5553)
	) name2605 (
		\Datai[6]_pad ,
		\InstQueue_reg[7][6]/NET0131 ,
		_w2232_,
		_w2378_,
		_w3058_
	);
	LUT2 #(
		.INIT('h1)
	) name2606 (
		_w2393_,
		_w3058_,
		_w3059_
	);
	LUT4 #(
		.INIT('hc055)
	) name2607 (
		\InstQueue_reg[7][6]/NET0131 ,
		_w523_,
		_w528_,
		_w2232_,
		_w3060_
	);
	LUT2 #(
		.INIT('h2)
	) name2608 (
		\InstQueue_reg[7][6]/NET0131 ,
		_w2227_,
		_w3061_
	);
	LUT3 #(
		.INIT('h0d)
	) name2609 (
		_w1212_,
		_w3058_,
		_w3061_,
		_w3062_
	);
	LUT3 #(
		.INIT('hd0)
	) name2610 (
		_w710_,
		_w3060_,
		_w3062_,
		_w3063_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name2611 (
		_w695_,
		_w3057_,
		_w3059_,
		_w3063_,
		_w3064_
	);
	LUT4 #(
		.INIT('h6c00)
	) name2612 (
		\Datai[18]_pad ,
		\Datai[19]_pad ,
		_w2211_,
		_w2378_,
		_w3065_
	);
	LUT4 #(
		.INIT('haa80)
	) name2613 (
		\DataWidth_reg[1]/NET0131 ,
		_w2365_,
		_w2811_,
		_w3065_,
		_w3066_
	);
	LUT4 #(
		.INIT('h5553)
	) name2614 (
		\Datai[3]_pad ,
		\InstQueue_reg[8][3]/NET0131 ,
		_w2232_,
		_w2234_,
		_w3067_
	);
	LUT2 #(
		.INIT('h1)
	) name2615 (
		_w2404_,
		_w3067_,
		_w3068_
	);
	LUT4 #(
		.INIT('hc055)
	) name2616 (
		\InstQueue_reg[8][3]/NET0131 ,
		_w511_,
		_w516_,
		_w2234_,
		_w3069_
	);
	LUT2 #(
		.INIT('h2)
	) name2617 (
		\InstQueue_reg[8][3]/NET0131 ,
		_w2227_,
		_w3070_
	);
	LUT3 #(
		.INIT('h0d)
	) name2618 (
		_w1212_,
		_w3067_,
		_w3070_,
		_w3071_
	);
	LUT3 #(
		.INIT('hd0)
	) name2619 (
		_w710_,
		_w3069_,
		_w3071_,
		_w3072_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name2620 (
		_w695_,
		_w3066_,
		_w3068_,
		_w3072_,
		_w3073_
	);
	LUT4 #(
		.INIT('h6c00)
	) name2621 (
		\Datai[21]_pad ,
		\Datai[22]_pad ,
		_w2212_,
		_w2378_,
		_w3074_
	);
	LUT4 #(
		.INIT('haa80)
	) name2622 (
		\DataWidth_reg[1]/NET0131 ,
		_w2365_,
		_w2821_,
		_w3074_,
		_w3075_
	);
	LUT4 #(
		.INIT('h5553)
	) name2623 (
		\Datai[6]_pad ,
		\InstQueue_reg[8][6]/NET0131 ,
		_w2232_,
		_w2234_,
		_w3076_
	);
	LUT2 #(
		.INIT('h1)
	) name2624 (
		_w2404_,
		_w3076_,
		_w3077_
	);
	LUT4 #(
		.INIT('hc055)
	) name2625 (
		\InstQueue_reg[8][6]/NET0131 ,
		_w523_,
		_w528_,
		_w2234_,
		_w3078_
	);
	LUT2 #(
		.INIT('h2)
	) name2626 (
		\InstQueue_reg[8][6]/NET0131 ,
		_w2227_,
		_w3079_
	);
	LUT3 #(
		.INIT('h0d)
	) name2627 (
		_w1212_,
		_w3076_,
		_w3079_,
		_w3080_
	);
	LUT3 #(
		.INIT('hd0)
	) name2628 (
		_w710_,
		_w3078_,
		_w3080_,
		_w3081_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name2629 (
		_w695_,
		_w3075_,
		_w3077_,
		_w3081_,
		_w3082_
	);
	LUT4 #(
		.INIT('h6c00)
	) name2630 (
		\Datai[18]_pad ,
		\Datai[19]_pad ,
		_w2211_,
		_w2232_,
		_w3083_
	);
	LUT4 #(
		.INIT('haa80)
	) name2631 (
		\DataWidth_reg[1]/NET0131 ,
		_w2378_,
		_w2811_,
		_w3083_,
		_w3084_
	);
	LUT4 #(
		.INIT('h5553)
	) name2632 (
		\Datai[3]_pad ,
		\InstQueue_reg[9][3]/NET0131 ,
		_w2237_,
		_w2234_,
		_w3085_
	);
	LUT2 #(
		.INIT('h1)
	) name2633 (
		_w2415_,
		_w3085_,
		_w3086_
	);
	LUT4 #(
		.INIT('hc055)
	) name2634 (
		\InstQueue_reg[9][3]/NET0131 ,
		_w511_,
		_w516_,
		_w2237_,
		_w3087_
	);
	LUT2 #(
		.INIT('h2)
	) name2635 (
		\InstQueue_reg[9][3]/NET0131 ,
		_w2227_,
		_w3088_
	);
	LUT3 #(
		.INIT('h0d)
	) name2636 (
		_w1212_,
		_w3085_,
		_w3088_,
		_w3089_
	);
	LUT3 #(
		.INIT('hd0)
	) name2637 (
		_w710_,
		_w3087_,
		_w3089_,
		_w3090_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name2638 (
		_w695_,
		_w3084_,
		_w3086_,
		_w3090_,
		_w3091_
	);
	LUT4 #(
		.INIT('h6c00)
	) name2639 (
		\Datai[21]_pad ,
		\Datai[22]_pad ,
		_w2212_,
		_w2232_,
		_w3092_
	);
	LUT4 #(
		.INIT('haa80)
	) name2640 (
		\DataWidth_reg[1]/NET0131 ,
		_w2378_,
		_w2821_,
		_w3092_,
		_w3093_
	);
	LUT4 #(
		.INIT('h5553)
	) name2641 (
		\Datai[6]_pad ,
		\InstQueue_reg[9][6]/NET0131 ,
		_w2237_,
		_w2234_,
		_w3094_
	);
	LUT2 #(
		.INIT('h1)
	) name2642 (
		_w2415_,
		_w3094_,
		_w3095_
	);
	LUT4 #(
		.INIT('hc055)
	) name2643 (
		\InstQueue_reg[9][6]/NET0131 ,
		_w523_,
		_w528_,
		_w2237_,
		_w3096_
	);
	LUT2 #(
		.INIT('h2)
	) name2644 (
		\InstQueue_reg[9][6]/NET0131 ,
		_w2227_,
		_w3097_
	);
	LUT3 #(
		.INIT('h0d)
	) name2645 (
		_w1212_,
		_w3094_,
		_w3097_,
		_w3098_
	);
	LUT3 #(
		.INIT('hd0)
	) name2646 (
		_w710_,
		_w3096_,
		_w3098_,
		_w3099_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name2647 (
		_w695_,
		_w3093_,
		_w3095_,
		_w3099_,
		_w3100_
	);
	LUT4 #(
		.INIT('hfe25)
	) name2648 (
		\State2_reg[0]/NET0131 ,
		\State2_reg[1]/NET0131 ,
		\State2_reg[2]/NET0131 ,
		\State2_reg[3]/NET0131 ,
		_w3101_
	);
	LUT4 #(
		.INIT('hfc21)
	) name2649 (
		\State2_reg[0]/NET0131 ,
		\State2_reg[1]/NET0131 ,
		\State2_reg[2]/NET0131 ,
		\State2_reg[3]/NET0131 ,
		_w3102_
	);
	LUT4 #(
		.INIT('h08aa)
	) name2650 (
		\PhyAddrPointer_reg[0]/NET0131 ,
		_w690_,
		_w1634_,
		_w3102_,
		_w3103_
	);
	LUT2 #(
		.INIT('h8)
	) name2651 (
		_w608_,
		_w2040_,
		_w3104_
	);
	LUT4 #(
		.INIT('h1113)
	) name2652 (
		_w690_,
		_w2045_,
		_w2043_,
		_w3104_,
		_w3105_
	);
	LUT2 #(
		.INIT('hb)
	) name2653 (
		_w3103_,
		_w3105_,
		_w3106_
	);
	LUT4 #(
		.INIT('h5014)
	) name2654 (
		\DataWidth_reg[1]/NET0131 ,
		\PhyAddrPointer_reg[0]/NET0131 ,
		\PhyAddrPointer_reg[1]/NET0131 ,
		_w1214_,
		_w3107_
	);
	LUT2 #(
		.INIT('h2)
	) name2655 (
		\DataWidth_reg[1]/NET0131 ,
		\rEIP_reg[1]/NET0131 ,
		_w3108_
	);
	LUT2 #(
		.INIT('h2)
	) name2656 (
		_w695_,
		_w3108_,
		_w3109_
	);
	LUT4 #(
		.INIT('h00fe)
	) name2657 (
		_w586_,
		_w582_,
		_w589_,
		_w566_,
		_w3110_
	);
	LUT2 #(
		.INIT('h2)
	) name2658 (
		\rEIP_reg[1]/NET0131 ,
		_w3110_,
		_w3111_
	);
	LUT3 #(
		.INIT('h23)
	) name2659 (
		\DataWidth_reg[1]/NET0131 ,
		\EBX_reg[1]/NET0131 ,
		_w645_,
		_w3112_
	);
	LUT3 #(
		.INIT('h02)
	) name2660 (
		_w589_,
		_w566_,
		_w3112_,
		_w3113_
	);
	LUT2 #(
		.INIT('h6)
	) name2661 (
		\EBX_reg[0]/NET0131 ,
		\EBX_reg[1]/NET0131 ,
		_w3114_
	);
	LUT3 #(
		.INIT('h60)
	) name2662 (
		\EBX_reg[0]/NET0131 ,
		\EBX_reg[1]/NET0131 ,
		\EBX_reg[31]/NET0131 ,
		_w3115_
	);
	LUT2 #(
		.INIT('h1)
	) name2663 (
		\DataWidth_reg[1]/NET0131 ,
		READY_n_pad,
		_w3116_
	);
	LUT4 #(
		.INIT('hf3a2)
	) name2664 (
		\DataWidth_reg[1]/NET0131 ,
		\EBX_reg[1]/NET0131 ,
		\EBX_reg[31]/NET0131 ,
		READY_n_pad,
		_w3117_
	);
	LUT2 #(
		.INIT('h4)
	) name2665 (
		_w3115_,
		_w3117_,
		_w3118_
	);
	LUT3 #(
		.INIT('h02)
	) name2666 (
		_w582_,
		_w566_,
		_w3118_,
		_w3119_
	);
	LUT3 #(
		.INIT('h10)
	) name2667 (
		\DataWidth_reg[1]/NET0131 ,
		READY_n_pad,
		\rEIP_reg[1]/NET0131 ,
		_w3120_
	);
	LUT3 #(
		.INIT('h0e)
	) name2668 (
		_w3113_,
		_w3119_,
		_w3120_,
		_w3121_
	);
	LUT3 #(
		.INIT('h02)
	) name2669 (
		_w586_,
		_w650_,
		_w566_,
		_w3122_
	);
	LUT4 #(
		.INIT('h0008)
	) name2670 (
		_w589_,
		_w594_,
		_w566_,
		_w3112_,
		_w3123_
	);
	LUT2 #(
		.INIT('h1)
	) name2671 (
		_w3122_,
		_w3123_,
		_w3124_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name2672 (
		_w690_,
		_w3121_,
		_w3111_,
		_w3124_,
		_w3125_
	);
	LUT4 #(
		.INIT('h5f13)
	) name2673 (
		\PhyAddrPointer_reg[1]/NET0131 ,
		\rEIP_reg[1]/NET0131 ,
		_w706_,
		_w3101_,
		_w3126_
	);
	LUT4 #(
		.INIT('hbaff)
	) name2674 (
		_w3125_,
		_w3107_,
		_w3109_,
		_w3126_,
		_w3127_
	);
	LUT3 #(
		.INIT('h6c)
	) name2675 (
		\PhyAddrPointer_reg[1]/NET0131 ,
		\PhyAddrPointer_reg[20]/NET0131 ,
		_w1520_,
		_w3128_
	);
	LUT2 #(
		.INIT('h4)
	) name2676 (
		\PhyAddrPointer_reg[0]/NET0131 ,
		_w1386_,
		_w3129_
	);
	LUT2 #(
		.INIT('h8)
	) name2677 (
		_w1198_,
		_w3129_,
		_w3130_
	);
	LUT3 #(
		.INIT('h10)
	) name2678 (
		_w1390_,
		_w1501_,
		_w3130_,
		_w3131_
	);
	LUT2 #(
		.INIT('h4)
	) name2679 (
		_w1621_,
		_w3131_,
		_w3132_
	);
	LUT4 #(
		.INIT('h8111)
	) name2680 (
		\PhyAddrPointer_reg[18]/NET0131 ,
		\PhyAddrPointer_reg[19]/NET0131 ,
		\PhyAddrPointer_reg[1]/NET0131 ,
		_w1201_,
		_w3133_
	);
	LUT4 #(
		.INIT('h1000)
	) name2681 (
		_w1621_,
		_w1640_,
		_w3131_,
		_w3133_,
		_w3134_
	);
	LUT2 #(
		.INIT('h8)
	) name2682 (
		_w2008_,
		_w3134_,
		_w3135_
	);
	LUT4 #(
		.INIT('h0514)
	) name2683 (
		\DataWidth_reg[1]/NET0131 ,
		_w1214_,
		_w3128_,
		_w3135_,
		_w3136_
	);
	LUT2 #(
		.INIT('h2)
	) name2684 (
		\DataWidth_reg[1]/NET0131 ,
		\rEIP_reg[20]/NET0131 ,
		_w3137_
	);
	LUT2 #(
		.INIT('h2)
	) name2685 (
		_w695_,
		_w3137_,
		_w3138_
	);
	LUT4 #(
		.INIT('h0001)
	) name2686 (
		\EBX_reg[0]/NET0131 ,
		\EBX_reg[1]/NET0131 ,
		\EBX_reg[2]/NET0131 ,
		\EBX_reg[3]/NET0131 ,
		_w3139_
	);
	LUT4 #(
		.INIT('h0100)
	) name2687 (
		\EBX_reg[4]/NET0131 ,
		\EBX_reg[5]/NET0131 ,
		\EBX_reg[6]/NET0131 ,
		_w3139_,
		_w3140_
	);
	LUT2 #(
		.INIT('h1)
	) name2688 (
		\EBX_reg[10]/NET0131 ,
		\EBX_reg[9]/NET0131 ,
		_w3141_
	);
	LUT4 #(
		.INIT('h1000)
	) name2689 (
		\EBX_reg[7]/NET0131 ,
		\EBX_reg[8]/NET0131 ,
		_w3140_,
		_w3141_,
		_w3142_
	);
	LUT2 #(
		.INIT('h1)
	) name2690 (
		\EBX_reg[11]/NET0131 ,
		\EBX_reg[12]/NET0131 ,
		_w3143_
	);
	LUT4 #(
		.INIT('h1000)
	) name2691 (
		\EBX_reg[13]/NET0131 ,
		\EBX_reg[14]/NET0131 ,
		_w3142_,
		_w3143_,
		_w3144_
	);
	LUT2 #(
		.INIT('h1)
	) name2692 (
		\EBX_reg[15]/NET0131 ,
		\EBX_reg[16]/NET0131 ,
		_w3145_
	);
	LUT4 #(
		.INIT('h1000)
	) name2693 (
		\EBX_reg[17]/NET0131 ,
		\EBX_reg[18]/NET0131 ,
		_w3144_,
		_w3145_,
		_w3146_
	);
	LUT3 #(
		.INIT('h8c)
	) name2694 (
		\EBX_reg[19]/NET0131 ,
		\EBX_reg[31]/NET0131 ,
		_w3146_,
		_w3147_
	);
	LUT4 #(
		.INIT('h8000)
	) name2695 (
		\rEIP_reg[1]/NET0131 ,
		\rEIP_reg[2]/NET0131 ,
		\rEIP_reg[3]/NET0131 ,
		\rEIP_reg[4]/NET0131 ,
		_w3148_
	);
	LUT4 #(
		.INIT('h8000)
	) name2696 (
		\rEIP_reg[5]/NET0131 ,
		\rEIP_reg[6]/NET0131 ,
		\rEIP_reg[7]/NET0131 ,
		_w3148_,
		_w3149_
	);
	LUT4 #(
		.INIT('h8000)
	) name2697 (
		\rEIP_reg[10]/NET0131 ,
		\rEIP_reg[8]/NET0131 ,
		\rEIP_reg[9]/NET0131 ,
		_w3149_,
		_w3150_
	);
	LUT2 #(
		.INIT('h8)
	) name2698 (
		\rEIP_reg[12]/NET0131 ,
		\rEIP_reg[13]/NET0131 ,
		_w3151_
	);
	LUT3 #(
		.INIT('h80)
	) name2699 (
		\rEIP_reg[12]/NET0131 ,
		\rEIP_reg[13]/NET0131 ,
		\rEIP_reg[14]/NET0131 ,
		_w3152_
	);
	LUT4 #(
		.INIT('h8000)
	) name2700 (
		\rEIP_reg[12]/NET0131 ,
		\rEIP_reg[13]/NET0131 ,
		\rEIP_reg[14]/NET0131 ,
		\rEIP_reg[15]/NET0131 ,
		_w3153_
	);
	LUT3 #(
		.INIT('h80)
	) name2701 (
		\rEIP_reg[11]/NET0131 ,
		_w3150_,
		_w3153_,
		_w3154_
	);
	LUT4 #(
		.INIT('h8000)
	) name2702 (
		\rEIP_reg[11]/NET0131 ,
		\rEIP_reg[16]/NET0131 ,
		_w3150_,
		_w3153_,
		_w3155_
	);
	LUT2 #(
		.INIT('h8)
	) name2703 (
		\rEIP_reg[17]/NET0131 ,
		\rEIP_reg[18]/NET0131 ,
		_w3156_
	);
	LUT2 #(
		.INIT('h8)
	) name2704 (
		\rEIP_reg[19]/NET0131 ,
		\rEIP_reg[20]/NET0131 ,
		_w3157_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name2705 (
		\rEIP_reg[19]/NET0131 ,
		\rEIP_reg[20]/NET0131 ,
		_w3155_,
		_w3156_,
		_w3158_
	);
	LUT4 #(
		.INIT('h2202)
	) name2706 (
		_w582_,
		_w566_,
		_w3116_,
		_w3158_,
		_w3159_
	);
	LUT4 #(
		.INIT('hde00)
	) name2707 (
		\EBX_reg[20]/NET0131 ,
		_w3116_,
		_w3147_,
		_w3159_,
		_w3160_
	);
	LUT3 #(
		.INIT('h04)
	) name2708 (
		_w594_,
		_w3116_,
		_w3158_,
		_w3161_
	);
	LUT3 #(
		.INIT('h23)
	) name2709 (
		\DataWidth_reg[1]/NET0131 ,
		\EBX_reg[20]/NET0131 ,
		_w645_,
		_w3162_
	);
	LUT3 #(
		.INIT('h02)
	) name2710 (
		_w589_,
		_w566_,
		_w3162_,
		_w3163_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name2711 (
		\rEIP_reg[20]/NET0131 ,
		_w3110_,
		_w3161_,
		_w3163_,
		_w3164_
	);
	LUT4 #(
		.INIT('h5f13)
	) name2712 (
		\PhyAddrPointer_reg[20]/NET0131 ,
		\rEIP_reg[20]/NET0131 ,
		_w706_,
		_w3101_,
		_w3165_
	);
	LUT4 #(
		.INIT('h7500)
	) name2713 (
		_w690_,
		_w3160_,
		_w3164_,
		_w3165_,
		_w3166_
	);
	LUT3 #(
		.INIT('h4f)
	) name2714 (
		_w3136_,
		_w3138_,
		_w3166_,
		_w3167_
	);
	LUT2 #(
		.INIT('h4)
	) name2715 (
		_w3128_,
		_w3134_,
		_w3168_
	);
	LUT4 #(
		.INIT('h0514)
	) name2716 (
		\DataWidth_reg[1]/NET0131 ,
		_w1214_,
		_w1671_,
		_w3168_,
		_w3169_
	);
	LUT2 #(
		.INIT('h2)
	) name2717 (
		\DataWidth_reg[1]/NET0131 ,
		\rEIP_reg[21]/NET0131 ,
		_w3170_
	);
	LUT2 #(
		.INIT('h2)
	) name2718 (
		_w695_,
		_w3170_,
		_w3171_
	);
	LUT4 #(
		.INIT('he0f0)
	) name2719 (
		\EBX_reg[19]/NET0131 ,
		\EBX_reg[20]/NET0131 ,
		\EBX_reg[31]/NET0131 ,
		_w3146_,
		_w3172_
	);
	LUT3 #(
		.INIT('h80)
	) name2720 (
		\rEIP_reg[19]/NET0131 ,
		\rEIP_reg[20]/NET0131 ,
		\rEIP_reg[21]/NET0131 ,
		_w3173_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name2721 (
		\rEIP_reg[21]/NET0131 ,
		_w3155_,
		_w3156_,
		_w3157_,
		_w3174_
	);
	LUT4 #(
		.INIT('h2202)
	) name2722 (
		_w582_,
		_w566_,
		_w3116_,
		_w3174_,
		_w3175_
	);
	LUT4 #(
		.INIT('hde00)
	) name2723 (
		\EBX_reg[21]/NET0131 ,
		_w3116_,
		_w3172_,
		_w3175_,
		_w3176_
	);
	LUT3 #(
		.INIT('h04)
	) name2724 (
		_w594_,
		_w3116_,
		_w3174_,
		_w3177_
	);
	LUT3 #(
		.INIT('h23)
	) name2725 (
		\DataWidth_reg[1]/NET0131 ,
		\EBX_reg[21]/NET0131 ,
		_w645_,
		_w3178_
	);
	LUT3 #(
		.INIT('h02)
	) name2726 (
		_w589_,
		_w566_,
		_w3178_,
		_w3179_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name2727 (
		\rEIP_reg[21]/NET0131 ,
		_w3110_,
		_w3177_,
		_w3179_,
		_w3180_
	);
	LUT4 #(
		.INIT('h5f13)
	) name2728 (
		\PhyAddrPointer_reg[21]/NET0131 ,
		\rEIP_reg[21]/NET0131 ,
		_w706_,
		_w3101_,
		_w3181_
	);
	LUT4 #(
		.INIT('h7500)
	) name2729 (
		_w690_,
		_w3176_,
		_w3180_,
		_w3181_,
		_w3182_
	);
	LUT3 #(
		.INIT('h4f)
	) name2730 (
		_w3169_,
		_w3171_,
		_w3182_,
		_w3183_
	);
	LUT3 #(
		.INIT('h0e)
	) name2731 (
		_w1406_,
		_w1670_,
		_w3128_,
		_w3184_
	);
	LUT3 #(
		.INIT('h80)
	) name2732 (
		_w2008_,
		_w3134_,
		_w3184_,
		_w3185_
	);
	LUT4 #(
		.INIT('h0514)
	) name2733 (
		\DataWidth_reg[1]/NET0131 ,
		_w1214_,
		_w1532_,
		_w3185_,
		_w3186_
	);
	LUT2 #(
		.INIT('h2)
	) name2734 (
		\DataWidth_reg[1]/NET0131 ,
		\rEIP_reg[22]/NET0131 ,
		_w3187_
	);
	LUT2 #(
		.INIT('h2)
	) name2735 (
		_w695_,
		_w3187_,
		_w3188_
	);
	LUT2 #(
		.INIT('h4)
	) name2736 (
		_w3186_,
		_w3188_,
		_w3189_
	);
	LUT2 #(
		.INIT('h2)
	) name2737 (
		\rEIP_reg[22]/NET0131 ,
		_w3110_,
		_w3190_
	);
	LUT3 #(
		.INIT('h23)
	) name2738 (
		\DataWidth_reg[1]/NET0131 ,
		\EBX_reg[22]/NET0131 ,
		_w645_,
		_w3191_
	);
	LUT3 #(
		.INIT('h02)
	) name2739 (
		_w589_,
		_w566_,
		_w3191_,
		_w3192_
	);
	LUT4 #(
		.INIT('h0100)
	) name2740 (
		\EBX_reg[19]/NET0131 ,
		\EBX_reg[20]/NET0131 ,
		\EBX_reg[21]/NET0131 ,
		_w3146_,
		_w3193_
	);
	LUT4 #(
		.INIT('h0509)
	) name2741 (
		\EBX_reg[22]/NET0131 ,
		\EBX_reg[31]/NET0131 ,
		_w3116_,
		_w3193_,
		_w3194_
	);
	LUT3 #(
		.INIT('h80)
	) name2742 (
		\rEIP_reg[17]/NET0131 ,
		\rEIP_reg[18]/NET0131 ,
		\rEIP_reg[22]/NET0131 ,
		_w3195_
	);
	LUT2 #(
		.INIT('h8)
	) name2743 (
		_w3173_,
		_w3195_,
		_w3196_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name2744 (
		\rEIP_reg[22]/NET0131 ,
		_w3155_,
		_w3156_,
		_w3173_,
		_w3197_
	);
	LUT4 #(
		.INIT('h0008)
	) name2745 (
		_w589_,
		_w594_,
		_w566_,
		_w3191_,
		_w3198_
	);
	LUT3 #(
		.INIT('h02)
	) name2746 (
		_w3116_,
		_w3197_,
		_w3198_,
		_w3199_
	);
	LUT4 #(
		.INIT('h00ce)
	) name2747 (
		_w2101_,
		_w3192_,
		_w3194_,
		_w3199_,
		_w3200_
	);
	LUT4 #(
		.INIT('h5f13)
	) name2748 (
		\PhyAddrPointer_reg[22]/NET0131 ,
		\rEIP_reg[22]/NET0131 ,
		_w706_,
		_w3101_,
		_w3201_
	);
	LUT4 #(
		.INIT('h5700)
	) name2749 (
		_w690_,
		_w3190_,
		_w3200_,
		_w3201_,
		_w3202_
	);
	LUT2 #(
		.INIT('hb)
	) name2750 (
		_w3189_,
		_w3202_,
		_w3203_
	);
	LUT4 #(
		.INIT('h0098)
	) name2751 (
		\PhyAddrPointer_reg[22]/NET0131 ,
		_w1406_,
		_w1670_,
		_w3128_,
		_w3204_
	);
	LUT3 #(
		.INIT('h80)
	) name2752 (
		_w2008_,
		_w3134_,
		_w3204_,
		_w3205_
	);
	LUT4 #(
		.INIT('h0514)
	) name2753 (
		\DataWidth_reg[1]/NET0131 ,
		_w1214_,
		_w1407_,
		_w3205_,
		_w3206_
	);
	LUT2 #(
		.INIT('h2)
	) name2754 (
		\DataWidth_reg[1]/NET0131 ,
		\rEIP_reg[23]/NET0131 ,
		_w3207_
	);
	LUT2 #(
		.INIT('h2)
	) name2755 (
		_w695_,
		_w3207_,
		_w3208_
	);
	LUT2 #(
		.INIT('h4)
	) name2756 (
		_w3206_,
		_w3208_,
		_w3209_
	);
	LUT3 #(
		.INIT('h8c)
	) name2757 (
		\EBX_reg[22]/NET0131 ,
		\EBX_reg[31]/NET0131 ,
		_w3193_,
		_w3210_
	);
	LUT3 #(
		.INIT('h80)
	) name2758 (
		\rEIP_reg[23]/NET0131 ,
		_w3155_,
		_w3196_,
		_w3211_
	);
	LUT4 #(
		.INIT('h8444)
	) name2759 (
		\rEIP_reg[23]/NET0131 ,
		_w3116_,
		_w3155_,
		_w3196_,
		_w3212_
	);
	LUT3 #(
		.INIT('h02)
	) name2760 (
		_w582_,
		_w566_,
		_w3212_,
		_w3213_
	);
	LUT4 #(
		.INIT('hde00)
	) name2761 (
		\EBX_reg[23]/NET0131 ,
		_w3116_,
		_w3210_,
		_w3213_,
		_w3214_
	);
	LUT4 #(
		.INIT('h8444)
	) name2762 (
		\rEIP_reg[23]/NET0131 ,
		_w688_,
		_w3155_,
		_w3196_,
		_w3215_
	);
	LUT3 #(
		.INIT('h23)
	) name2763 (
		\DataWidth_reg[1]/NET0131 ,
		\EBX_reg[23]/NET0131 ,
		_w645_,
		_w3216_
	);
	LUT4 #(
		.INIT('h0002)
	) name2764 (
		_w589_,
		_w566_,
		_w3216_,
		_w3215_,
		_w3217_
	);
	LUT3 #(
		.INIT('h0d)
	) name2765 (
		\rEIP_reg[23]/NET0131 ,
		_w3110_,
		_w3217_,
		_w3218_
	);
	LUT4 #(
		.INIT('h5f13)
	) name2766 (
		\PhyAddrPointer_reg[23]/NET0131 ,
		\rEIP_reg[23]/NET0131 ,
		_w706_,
		_w3101_,
		_w3219_
	);
	LUT4 #(
		.INIT('h7500)
	) name2767 (
		_w690_,
		_w3214_,
		_w3218_,
		_w3219_,
		_w3220_
	);
	LUT2 #(
		.INIT('hb)
	) name2768 (
		_w3209_,
		_w3220_,
		_w3221_
	);
	LUT4 #(
		.INIT('he0f0)
	) name2769 (
		\EBX_reg[22]/NET0131 ,
		\EBX_reg[23]/NET0131 ,
		\EBX_reg[31]/NET0131 ,
		_w3193_,
		_w3222_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name2770 (
		\rEIP_reg[23]/NET0131 ,
		\rEIP_reg[24]/NET0131 ,
		_w3155_,
		_w3196_,
		_w3223_
	);
	LUT3 #(
		.INIT('h15)
	) name2771 (
		_w566_,
		_w3116_,
		_w3223_,
		_w3224_
	);
	LUT4 #(
		.INIT('hed00)
	) name2772 (
		\EBX_reg[24]/NET0131 ,
		_w3116_,
		_w3222_,
		_w3224_,
		_w3225_
	);
	LUT3 #(
		.INIT('h04)
	) name2773 (
		\rEIP_reg[24]/NET0131 ,
		_w563_,
		_w565_,
		_w3226_
	);
	LUT2 #(
		.INIT('h2)
	) name2774 (
		_w582_,
		_w3226_,
		_w3227_
	);
	LUT2 #(
		.INIT('h2)
	) name2775 (
		_w688_,
		_w3223_,
		_w3228_
	);
	LUT3 #(
		.INIT('h23)
	) name2776 (
		\DataWidth_reg[1]/NET0131 ,
		\EBX_reg[24]/NET0131 ,
		_w645_,
		_w3229_
	);
	LUT3 #(
		.INIT('h02)
	) name2777 (
		_w589_,
		_w566_,
		_w3229_,
		_w3230_
	);
	LUT3 #(
		.INIT('h8a)
	) name2778 (
		\rEIP_reg[24]/NET0131 ,
		_w586_,
		_w582_,
		_w3231_
	);
	LUT4 #(
		.INIT('h8acf)
	) name2779 (
		_w3110_,
		_w3228_,
		_w3230_,
		_w3231_,
		_w3232_
	);
	LUT4 #(
		.INIT('h20aa)
	) name2780 (
		_w690_,
		_w3225_,
		_w3227_,
		_w3232_,
		_w3233_
	);
	LUT4 #(
		.INIT('h4000)
	) name2781 (
		_w1407_,
		_w2008_,
		_w3134_,
		_w3204_,
		_w3234_
	);
	LUT4 #(
		.INIT('h0514)
	) name2782 (
		\DataWidth_reg[1]/NET0131 ,
		_w1214_,
		_w1543_,
		_w3234_,
		_w3235_
	);
	LUT2 #(
		.INIT('h2)
	) name2783 (
		\DataWidth_reg[1]/NET0131 ,
		\rEIP_reg[24]/NET0131 ,
		_w3236_
	);
	LUT2 #(
		.INIT('h2)
	) name2784 (
		_w695_,
		_w3236_,
		_w3237_
	);
	LUT4 #(
		.INIT('h5f13)
	) name2785 (
		\PhyAddrPointer_reg[24]/NET0131 ,
		\rEIP_reg[24]/NET0131 ,
		_w706_,
		_w3101_,
		_w3238_
	);
	LUT3 #(
		.INIT('hb0)
	) name2786 (
		_w3235_,
		_w3237_,
		_w3238_,
		_w3239_
	);
	LUT2 #(
		.INIT('hb)
	) name2787 (
		_w3233_,
		_w3239_,
		_w3240_
	);
	LUT2 #(
		.INIT('h1)
	) name2788 (
		_w1407_,
		_w1543_,
		_w3241_
	);
	LUT3 #(
		.INIT('h80)
	) name2789 (
		_w3134_,
		_w3204_,
		_w3241_,
		_w3242_
	);
	LUT4 #(
		.INIT('h0514)
	) name2790 (
		\DataWidth_reg[1]/NET0131 ,
		_w1214_,
		_w1684_,
		_w3242_,
		_w3243_
	);
	LUT2 #(
		.INIT('h2)
	) name2791 (
		\DataWidth_reg[1]/NET0131 ,
		\rEIP_reg[25]/NET0131 ,
		_w3244_
	);
	LUT2 #(
		.INIT('h2)
	) name2792 (
		_w695_,
		_w3244_,
		_w3245_
	);
	LUT2 #(
		.INIT('h4)
	) name2793 (
		_w3243_,
		_w3245_,
		_w3246_
	);
	LUT2 #(
		.INIT('h1)
	) name2794 (
		\EBX_reg[23]/NET0131 ,
		\EBX_reg[24]/NET0131 ,
		_w3247_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name2795 (
		\EBX_reg[22]/NET0131 ,
		\EBX_reg[31]/NET0131 ,
		_w3193_,
		_w3247_,
		_w3248_
	);
	LUT2 #(
		.INIT('h8)
	) name2796 (
		\rEIP_reg[24]/NET0131 ,
		\rEIP_reg[25]/NET0131 ,
		_w3249_
	);
	LUT4 #(
		.INIT('h8000)
	) name2797 (
		\rEIP_reg[23]/NET0131 ,
		_w3155_,
		_w3196_,
		_w3249_,
		_w3250_
	);
	LUT4 #(
		.INIT('h9030)
	) name2798 (
		\rEIP_reg[24]/NET0131 ,
		\rEIP_reg[25]/NET0131 ,
		_w3116_,
		_w3211_,
		_w3251_
	);
	LUT2 #(
		.INIT('h2)
	) name2799 (
		_w2101_,
		_w3251_,
		_w3252_
	);
	LUT4 #(
		.INIT('hde00)
	) name2800 (
		\EBX_reg[25]/NET0131 ,
		_w3116_,
		_w3248_,
		_w3252_,
		_w3253_
	);
	LUT4 #(
		.INIT('h9030)
	) name2801 (
		\rEIP_reg[24]/NET0131 ,
		\rEIP_reg[25]/NET0131 ,
		_w688_,
		_w3211_,
		_w3254_
	);
	LUT3 #(
		.INIT('h23)
	) name2802 (
		\DataWidth_reg[1]/NET0131 ,
		\EBX_reg[25]/NET0131 ,
		_w645_,
		_w3255_
	);
	LUT3 #(
		.INIT('h02)
	) name2803 (
		_w589_,
		_w566_,
		_w3255_,
		_w3256_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name2804 (
		\rEIP_reg[25]/NET0131 ,
		_w3110_,
		_w3254_,
		_w3256_,
		_w3257_
	);
	LUT4 #(
		.INIT('h5f13)
	) name2805 (
		\PhyAddrPointer_reg[25]/NET0131 ,
		\rEIP_reg[25]/NET0131 ,
		_w706_,
		_w3101_,
		_w3258_
	);
	LUT4 #(
		.INIT('h7500)
	) name2806 (
		_w690_,
		_w3253_,
		_w3257_,
		_w3258_,
		_w3259_
	);
	LUT2 #(
		.INIT('hb)
	) name2807 (
		_w3246_,
		_w3259_,
		_w3260_
	);
	LUT4 #(
		.INIT('h1110)
	) name2808 (
		_w1407_,
		_w1543_,
		_w1555_,
		_w1683_,
		_w3261_
	);
	LUT4 #(
		.INIT('h8000)
	) name2809 (
		_w2008_,
		_w3134_,
		_w3204_,
		_w3261_,
		_w3262_
	);
	LUT4 #(
		.INIT('h0514)
	) name2810 (
		\DataWidth_reg[1]/NET0131 ,
		_w1214_,
		_w1556_,
		_w3262_,
		_w3263_
	);
	LUT2 #(
		.INIT('h2)
	) name2811 (
		\DataWidth_reg[1]/NET0131 ,
		\rEIP_reg[26]/NET0131 ,
		_w3264_
	);
	LUT2 #(
		.INIT('h2)
	) name2812 (
		_w695_,
		_w3264_,
		_w3265_
	);
	LUT2 #(
		.INIT('h4)
	) name2813 (
		_w3263_,
		_w3265_,
		_w3266_
	);
	LUT4 #(
		.INIT('h0001)
	) name2814 (
		\EBX_reg[22]/NET0131 ,
		\EBX_reg[23]/NET0131 ,
		\EBX_reg[24]/NET0131 ,
		\EBX_reg[25]/NET0131 ,
		_w3267_
	);
	LUT3 #(
		.INIT('h2a)
	) name2815 (
		\EBX_reg[31]/NET0131 ,
		_w3193_,
		_w3267_,
		_w3268_
	);
	LUT3 #(
		.INIT('h80)
	) name2816 (
		\rEIP_reg[24]/NET0131 ,
		\rEIP_reg[25]/NET0131 ,
		\rEIP_reg[26]/NET0131 ,
		_w3269_
	);
	LUT4 #(
		.INIT('h8000)
	) name2817 (
		\rEIP_reg[23]/NET0131 ,
		_w3155_,
		_w3196_,
		_w3269_,
		_w3270_
	);
	LUT4 #(
		.INIT('hcc04)
	) name2818 (
		\rEIP_reg[26]/NET0131 ,
		_w3116_,
		_w3250_,
		_w3270_,
		_w3271_
	);
	LUT2 #(
		.INIT('h2)
	) name2819 (
		_w2101_,
		_w3271_,
		_w3272_
	);
	LUT4 #(
		.INIT('hde00)
	) name2820 (
		\EBX_reg[26]/NET0131 ,
		_w3116_,
		_w3268_,
		_w3272_,
		_w3273_
	);
	LUT4 #(
		.INIT('hcc04)
	) name2821 (
		\rEIP_reg[26]/NET0131 ,
		_w688_,
		_w3250_,
		_w3270_,
		_w3274_
	);
	LUT3 #(
		.INIT('h23)
	) name2822 (
		\DataWidth_reg[1]/NET0131 ,
		\EBX_reg[26]/NET0131 ,
		_w645_,
		_w3275_
	);
	LUT3 #(
		.INIT('h02)
	) name2823 (
		_w589_,
		_w566_,
		_w3275_,
		_w3276_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name2824 (
		\rEIP_reg[26]/NET0131 ,
		_w3110_,
		_w3274_,
		_w3276_,
		_w3277_
	);
	LUT4 #(
		.INIT('h5f13)
	) name2825 (
		\PhyAddrPointer_reg[26]/NET0131 ,
		\rEIP_reg[26]/NET0131 ,
		_w706_,
		_w3101_,
		_w3278_
	);
	LUT4 #(
		.INIT('h7500)
	) name2826 (
		_w690_,
		_w3273_,
		_w3277_,
		_w3278_,
		_w3279_
	);
	LUT2 #(
		.INIT('hb)
	) name2827 (
		_w3266_,
		_w3279_,
		_w3280_
	);
	LUT3 #(
		.INIT('h45)
	) name2828 (
		_w1214_,
		_w1556_,
		_w3262_,
		_w3281_
	);
	LUT2 #(
		.INIT('h2)
	) name2829 (
		\DataWidth_reg[1]/NET0131 ,
		\rEIP_reg[27]/NET0131 ,
		_w3282_
	);
	LUT2 #(
		.INIT('h2)
	) name2830 (
		_w695_,
		_w3282_,
		_w3283_
	);
	LUT4 #(
		.INIT('hbe00)
	) name2831 (
		\DataWidth_reg[1]/NET0131 ,
		_w1416_,
		_w3281_,
		_w3283_,
		_w3284_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name2832 (
		\EBX_reg[26]/NET0131 ,
		\EBX_reg[31]/NET0131 ,
		_w3193_,
		_w3267_,
		_w3285_
	);
	LUT3 #(
		.INIT('h84)
	) name2833 (
		\rEIP_reg[27]/NET0131 ,
		_w3116_,
		_w3270_,
		_w3286_
	);
	LUT2 #(
		.INIT('h2)
	) name2834 (
		_w2101_,
		_w3286_,
		_w3287_
	);
	LUT4 #(
		.INIT('hde00)
	) name2835 (
		\EBX_reg[27]/NET0131 ,
		_w3116_,
		_w3285_,
		_w3287_,
		_w3288_
	);
	LUT4 #(
		.INIT('h2010)
	) name2836 (
		\rEIP_reg[27]/NET0131 ,
		_w594_,
		_w3116_,
		_w3270_,
		_w3289_
	);
	LUT3 #(
		.INIT('h23)
	) name2837 (
		\DataWidth_reg[1]/NET0131 ,
		\EBX_reg[27]/NET0131 ,
		_w645_,
		_w3290_
	);
	LUT3 #(
		.INIT('h02)
	) name2838 (
		_w589_,
		_w566_,
		_w3290_,
		_w3291_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name2839 (
		\rEIP_reg[27]/NET0131 ,
		_w3110_,
		_w3289_,
		_w3291_,
		_w3292_
	);
	LUT4 #(
		.INIT('h5f13)
	) name2840 (
		\PhyAddrPointer_reg[27]/NET0131 ,
		\rEIP_reg[27]/NET0131 ,
		_w706_,
		_w3101_,
		_w3293_
	);
	LUT4 #(
		.INIT('h7500)
	) name2841 (
		_w690_,
		_w3288_,
		_w3292_,
		_w3293_,
		_w3294_
	);
	LUT2 #(
		.INIT('hb)
	) name2842 (
		_w3284_,
		_w3294_,
		_w3295_
	);
	LUT4 #(
		.INIT('h1000)
	) name2843 (
		\EBX_reg[26]/NET0131 ,
		\EBX_reg[27]/NET0131 ,
		_w3193_,
		_w3267_,
		_w3296_
	);
	LUT4 #(
		.INIT('h0509)
	) name2844 (
		\EBX_reg[28]/NET0131 ,
		\EBX_reg[31]/NET0131 ,
		_w3116_,
		_w3296_,
		_w3297_
	);
	LUT4 #(
		.INIT('h9030)
	) name2845 (
		\rEIP_reg[27]/NET0131 ,
		\rEIP_reg[28]/NET0131 ,
		_w3116_,
		_w3270_,
		_w3298_
	);
	LUT2 #(
		.INIT('h2)
	) name2846 (
		_w2101_,
		_w3298_,
		_w3299_
	);
	LUT4 #(
		.INIT('h9030)
	) name2847 (
		\rEIP_reg[27]/NET0131 ,
		\rEIP_reg[28]/NET0131 ,
		_w688_,
		_w3270_,
		_w3300_
	);
	LUT3 #(
		.INIT('h23)
	) name2848 (
		\DataWidth_reg[1]/NET0131 ,
		\EBX_reg[28]/NET0131 ,
		_w645_,
		_w3301_
	);
	LUT3 #(
		.INIT('h02)
	) name2849 (
		_w589_,
		_w566_,
		_w3301_,
		_w3302_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name2850 (
		\rEIP_reg[28]/NET0131 ,
		_w3110_,
		_w3300_,
		_w3302_,
		_w3303_
	);
	LUT4 #(
		.INIT('h20aa)
	) name2851 (
		_w690_,
		_w3297_,
		_w3299_,
		_w3303_,
		_w3304_
	);
	LUT4 #(
		.INIT('h5455)
	) name2852 (
		_w1214_,
		_w1416_,
		_w1556_,
		_w3262_,
		_w3305_
	);
	LUT2 #(
		.INIT('h2)
	) name2853 (
		\DataWidth_reg[1]/NET0131 ,
		\rEIP_reg[28]/NET0131 ,
		_w3306_
	);
	LUT2 #(
		.INIT('h2)
	) name2854 (
		_w695_,
		_w3306_,
		_w3307_
	);
	LUT4 #(
		.INIT('hbe00)
	) name2855 (
		\DataWidth_reg[1]/NET0131 ,
		_w1438_,
		_w3305_,
		_w3307_,
		_w3308_
	);
	LUT4 #(
		.INIT('h5f13)
	) name2856 (
		\PhyAddrPointer_reg[28]/NET0131 ,
		\rEIP_reg[28]/NET0131 ,
		_w706_,
		_w3101_,
		_w3309_
	);
	LUT3 #(
		.INIT('hef)
	) name2857 (
		_w3304_,
		_w3308_,
		_w3309_,
		_w3310_
	);
	LUT2 #(
		.INIT('h1)
	) name2858 (
		\EBX_reg[27]/NET0131 ,
		\EBX_reg[28]/NET0131 ,
		_w3311_
	);
	LUT4 #(
		.INIT('h4000)
	) name2859 (
		\EBX_reg[26]/NET0131 ,
		_w3193_,
		_w3267_,
		_w3311_,
		_w3312_
	);
	LUT4 #(
		.INIT('h0509)
	) name2860 (
		\EBX_reg[29]/NET0131 ,
		\EBX_reg[31]/NET0131 ,
		_w3116_,
		_w3312_,
		_w3313_
	);
	LUT4 #(
		.INIT('h8000)
	) name2861 (
		\rEIP_reg[27]/NET0131 ,
		\rEIP_reg[28]/NET0131 ,
		\rEIP_reg[29]/NET0131 ,
		_w3270_,
		_w3314_
	);
	LUT4 #(
		.INIT('h78f0)
	) name2862 (
		\rEIP_reg[27]/NET0131 ,
		\rEIP_reg[28]/NET0131 ,
		\rEIP_reg[29]/NET0131 ,
		_w3270_,
		_w3315_
	);
	LUT3 #(
		.INIT('ha2)
	) name2863 (
		_w2101_,
		_w3116_,
		_w3315_,
		_w3316_
	);
	LUT2 #(
		.INIT('h2)
	) name2864 (
		\rEIP_reg[29]/NET0131 ,
		_w3110_,
		_w3317_
	);
	LUT3 #(
		.INIT('h23)
	) name2865 (
		\DataWidth_reg[1]/NET0131 ,
		\EBX_reg[29]/NET0131 ,
		_w645_,
		_w3318_
	);
	LUT3 #(
		.INIT('h02)
	) name2866 (
		_w589_,
		_w566_,
		_w3318_,
		_w3319_
	);
	LUT3 #(
		.INIT('hd0)
	) name2867 (
		_w688_,
		_w3315_,
		_w3319_,
		_w3320_
	);
	LUT2 #(
		.INIT('h1)
	) name2868 (
		_w3317_,
		_w3320_,
		_w3321_
	);
	LUT4 #(
		.INIT('h20aa)
	) name2869 (
		_w690_,
		_w3313_,
		_w3316_,
		_w3321_,
		_w3322_
	);
	LUT4 #(
		.INIT('h9380)
	) name2870 (
		\PhyAddrPointer_reg[1]/NET0131 ,
		\PhyAddrPointer_reg[26]/NET0131 ,
		_w1205_,
		_w1683_,
		_w3323_
	);
	LUT3 #(
		.INIT('h10)
	) name2871 (
		_w1416_,
		_w1438_,
		_w3323_,
		_w3324_
	);
	LUT3 #(
		.INIT('h15)
	) name2872 (
		_w1214_,
		_w3242_,
		_w3324_,
		_w3325_
	);
	LUT2 #(
		.INIT('h2)
	) name2873 (
		\DataWidth_reg[1]/NET0131 ,
		\rEIP_reg[29]/NET0131 ,
		_w3326_
	);
	LUT2 #(
		.INIT('h2)
	) name2874 (
		_w695_,
		_w3326_,
		_w3327_
	);
	LUT4 #(
		.INIT('hbe00)
	) name2875 (
		\DataWidth_reg[1]/NET0131 ,
		_w1447_,
		_w3325_,
		_w3327_,
		_w3328_
	);
	LUT4 #(
		.INIT('h5f13)
	) name2876 (
		\PhyAddrPointer_reg[29]/NET0131 ,
		\rEIP_reg[29]/NET0131 ,
		_w706_,
		_w3101_,
		_w3329_
	);
	LUT3 #(
		.INIT('hef)
	) name2877 (
		_w3322_,
		_w3328_,
		_w3329_,
		_w3330_
	);
	LUT2 #(
		.INIT('h4)
	) name2878 (
		\PhyAddrPointer_reg[0]/NET0131 ,
		\PhyAddrPointer_reg[1]/NET0131 ,
		_w3331_
	);
	LUT4 #(
		.INIT('h0514)
	) name2879 (
		\DataWidth_reg[1]/NET0131 ,
		_w1214_,
		_w2426_,
		_w3331_,
		_w3332_
	);
	LUT2 #(
		.INIT('h2)
	) name2880 (
		\DataWidth_reg[1]/NET0131 ,
		\rEIP_reg[2]/NET0131 ,
		_w3333_
	);
	LUT2 #(
		.INIT('h2)
	) name2881 (
		_w695_,
		_w3333_,
		_w3334_
	);
	LUT2 #(
		.INIT('h2)
	) name2882 (
		\rEIP_reg[2]/NET0131 ,
		_w3110_,
		_w3335_
	);
	LUT3 #(
		.INIT('h14)
	) name2883 (
		\DataWidth_reg[1]/NET0131 ,
		\rEIP_reg[1]/NET0131 ,
		\rEIP_reg[2]/NET0131 ,
		_w3336_
	);
	LUT4 #(
		.INIT('h0373)
	) name2884 (
		\DataWidth_reg[1]/NET0131 ,
		\EBX_reg[2]/NET0131 ,
		_w645_,
		_w3336_,
		_w3337_
	);
	LUT3 #(
		.INIT('h02)
	) name2885 (
		_w589_,
		_w566_,
		_w3337_,
		_w3338_
	);
	LUT3 #(
		.INIT('h20)
	) name2886 (
		_w586_,
		_w566_,
		_w661_,
		_w3339_
	);
	LUT4 #(
		.INIT('h0110)
	) name2887 (
		\DataWidth_reg[1]/NET0131 ,
		READY_n_pad,
		\rEIP_reg[1]/NET0131 ,
		\rEIP_reg[2]/NET0131 ,
		_w3340_
	);
	LUT3 #(
		.INIT('he0)
	) name2888 (
		\EBX_reg[0]/NET0131 ,
		\EBX_reg[1]/NET0131 ,
		\EBX_reg[31]/NET0131 ,
		_w3341_
	);
	LUT4 #(
		.INIT('h0e0d)
	) name2889 (
		\EBX_reg[2]/NET0131 ,
		_w3116_,
		_w3340_,
		_w3341_,
		_w3342_
	);
	LUT3 #(
		.INIT('h02)
	) name2890 (
		_w582_,
		_w566_,
		_w3342_,
		_w3343_
	);
	LUT3 #(
		.INIT('h01)
	) name2891 (
		_w3339_,
		_w3343_,
		_w3338_,
		_w3344_
	);
	LUT4 #(
		.INIT('h5f13)
	) name2892 (
		\PhyAddrPointer_reg[2]/NET0131 ,
		\rEIP_reg[2]/NET0131 ,
		_w706_,
		_w3101_,
		_w3345_
	);
	LUT4 #(
		.INIT('h7500)
	) name2893 (
		_w690_,
		_w3335_,
		_w3344_,
		_w3345_,
		_w3346_
	);
	LUT3 #(
		.INIT('h4f)
	) name2894 (
		_w3332_,
		_w3334_,
		_w3346_,
		_w3347_
	);
	LUT2 #(
		.INIT('h2)
	) name2895 (
		\rEIP_reg[31]/NET0131 ,
		_w3110_,
		_w3348_
	);
	LUT3 #(
		.INIT('h01)
	) name2896 (
		\EBX_reg[27]/NET0131 ,
		\EBX_reg[28]/NET0131 ,
		\EBX_reg[29]/NET0131 ,
		_w3349_
	);
	LUT4 #(
		.INIT('h4000)
	) name2897 (
		\EBX_reg[26]/NET0131 ,
		_w3193_,
		_w3267_,
		_w3349_,
		_w3350_
	);
	LUT4 #(
		.INIT('h3020)
	) name2898 (
		\DataWidth_reg[1]/NET0131 ,
		\EBX_reg[30]/NET0131 ,
		\EBX_reg[31]/NET0131 ,
		READY_n_pad,
		_w3351_
	);
	LUT4 #(
		.INIT('h60c0)
	) name2899 (
		\rEIP_reg[30]/NET0131 ,
		\rEIP_reg[31]/NET0131 ,
		_w3116_,
		_w3314_,
		_w3352_
	);
	LUT4 #(
		.INIT('haa80)
	) name2900 (
		_w582_,
		_w3350_,
		_w3351_,
		_w3352_,
		_w3353_
	);
	LUT4 #(
		.INIT('h9030)
	) name2901 (
		\rEIP_reg[30]/NET0131 ,
		\rEIP_reg[31]/NET0131 ,
		_w688_,
		_w3314_,
		_w3354_
	);
	LUT3 #(
		.INIT('h23)
	) name2902 (
		\DataWidth_reg[1]/NET0131 ,
		\EBX_reg[31]/NET0131 ,
		_w645_,
		_w3355_
	);
	LUT2 #(
		.INIT('h2)
	) name2903 (
		_w589_,
		_w3355_,
		_w3356_
	);
	LUT2 #(
		.INIT('h4)
	) name2904 (
		_w3354_,
		_w3356_,
		_w3357_
	);
	LUT4 #(
		.INIT('h2223)
	) name2905 (
		_w566_,
		_w3348_,
		_w3353_,
		_w3357_,
		_w3358_
	);
	LUT2 #(
		.INIT('h8)
	) name2906 (
		\DataWidth_reg[1]/NET0131 ,
		\rEIP_reg[31]/NET0131 ,
		_w3359_
	);
	LUT3 #(
		.INIT('h90)
	) name2907 (
		\PhyAddrPointer_reg[29]/NET0131 ,
		_w1213_,
		_w2008_,
		_w3360_
	);
	LUT3 #(
		.INIT('h80)
	) name2908 (
		_w3242_,
		_w3324_,
		_w3360_,
		_w3361_
	);
	LUT4 #(
		.INIT('h4105)
	) name2909 (
		\DataWidth_reg[1]/NET0131 ,
		\PhyAddrPointer_reg[29]/NET0131 ,
		\PhyAddrPointer_reg[30]/NET0131 ,
		_w1213_,
		_w3362_
	);
	LUT2 #(
		.INIT('h4)
	) name2910 (
		_w1214_,
		_w3362_,
		_w3363_
	);
	LUT4 #(
		.INIT('ha888)
	) name2911 (
		_w695_,
		_w3359_,
		_w3361_,
		_w3363_,
		_w3364_
	);
	LUT4 #(
		.INIT('h5f13)
	) name2912 (
		\PhyAddrPointer_reg[31]/NET0131 ,
		\rEIP_reg[31]/NET0131 ,
		_w706_,
		_w3101_,
		_w3365_
	);
	LUT4 #(
		.INIT('hf2ff)
	) name2913 (
		_w690_,
		_w3358_,
		_w3364_,
		_w3365_,
		_w3366_
	);
	LUT3 #(
		.INIT('h40)
	) name2914 (
		\PhyAddrPointer_reg[0]/NET0131 ,
		\PhyAddrPointer_reg[1]/NET0131 ,
		\PhyAddrPointer_reg[2]/NET0131 ,
		_w3367_
	);
	LUT4 #(
		.INIT('h0514)
	) name2915 (
		\DataWidth_reg[1]/NET0131 ,
		_w1214_,
		_w2123_,
		_w3367_,
		_w3368_
	);
	LUT2 #(
		.INIT('h2)
	) name2916 (
		\DataWidth_reg[1]/NET0131 ,
		\rEIP_reg[3]/NET0131 ,
		_w3369_
	);
	LUT2 #(
		.INIT('h2)
	) name2917 (
		_w695_,
		_w3369_,
		_w3370_
	);
	LUT2 #(
		.INIT('h2)
	) name2918 (
		\rEIP_reg[3]/NET0131 ,
		_w3110_,
		_w3371_
	);
	LUT4 #(
		.INIT('hfe00)
	) name2919 (
		\EBX_reg[0]/NET0131 ,
		\EBX_reg[1]/NET0131 ,
		\EBX_reg[2]/NET0131 ,
		\EBX_reg[31]/NET0131 ,
		_w3372_
	);
	LUT3 #(
		.INIT('h12)
	) name2920 (
		\EBX_reg[3]/NET0131 ,
		_w3116_,
		_w3372_,
		_w3373_
	);
	LUT4 #(
		.INIT('h1540)
	) name2921 (
		\DataWidth_reg[1]/NET0131 ,
		\rEIP_reg[1]/NET0131 ,
		\rEIP_reg[2]/NET0131 ,
		\rEIP_reg[3]/NET0131 ,
		_w3374_
	);
	LUT2 #(
		.INIT('h4)
	) name2922 (
		READY_n_pad,
		_w3374_,
		_w3375_
	);
	LUT2 #(
		.INIT('h1)
	) name2923 (
		_w3373_,
		_w3375_,
		_w3376_
	);
	LUT3 #(
		.INIT('h02)
	) name2924 (
		_w582_,
		_w566_,
		_w3376_,
		_w3377_
	);
	LUT3 #(
		.INIT('h02)
	) name2925 (
		_w586_,
		_w566_,
		_w631_,
		_w3378_
	);
	LUT4 #(
		.INIT('h0373)
	) name2926 (
		\DataWidth_reg[1]/NET0131 ,
		\EBX_reg[3]/NET0131 ,
		_w645_,
		_w3374_,
		_w3379_
	);
	LUT3 #(
		.INIT('h02)
	) name2927 (
		_w589_,
		_w566_,
		_w3379_,
		_w3380_
	);
	LUT3 #(
		.INIT('h01)
	) name2928 (
		_w3378_,
		_w3380_,
		_w3377_,
		_w3381_
	);
	LUT4 #(
		.INIT('h5f13)
	) name2929 (
		\PhyAddrPointer_reg[3]/NET0131 ,
		\rEIP_reg[3]/NET0131 ,
		_w706_,
		_w3101_,
		_w3382_
	);
	LUT4 #(
		.INIT('h7500)
	) name2930 (
		_w690_,
		_w3371_,
		_w3381_,
		_w3382_,
		_w3383_
	);
	LUT3 #(
		.INIT('h4f)
	) name2931 (
		_w3368_,
		_w3370_,
		_w3383_,
		_w3384_
	);
	LUT4 #(
		.INIT('h4000)
	) name2932 (
		\PhyAddrPointer_reg[0]/NET0131 ,
		\PhyAddrPointer_reg[1]/NET0131 ,
		\PhyAddrPointer_reg[2]/NET0131 ,
		\PhyAddrPointer_reg[3]/NET0131 ,
		_w3385_
	);
	LUT4 #(
		.INIT('h0514)
	) name2933 (
		\DataWidth_reg[1]/NET0131 ,
		_w1214_,
		_w2010_,
		_w3385_,
		_w3386_
	);
	LUT2 #(
		.INIT('h2)
	) name2934 (
		\DataWidth_reg[1]/NET0131 ,
		\rEIP_reg[4]/NET0131 ,
		_w3387_
	);
	LUT2 #(
		.INIT('h2)
	) name2935 (
		_w695_,
		_w3387_,
		_w3388_
	);
	LUT4 #(
		.INIT('h0309)
	) name2936 (
		\EBX_reg[31]/NET0131 ,
		\EBX_reg[4]/NET0131 ,
		_w3116_,
		_w3139_,
		_w3389_
	);
	LUT4 #(
		.INIT('h7f80)
	) name2937 (
		\rEIP_reg[1]/NET0131 ,
		\rEIP_reg[2]/NET0131 ,
		\rEIP_reg[3]/NET0131 ,
		\rEIP_reg[4]/NET0131 ,
		_w3390_
	);
	LUT2 #(
		.INIT('h2)
	) name2938 (
		_w3116_,
		_w3390_,
		_w3391_
	);
	LUT2 #(
		.INIT('h1)
	) name2939 (
		_w3389_,
		_w3391_,
		_w3392_
	);
	LUT3 #(
		.INIT('h20)
	) name2940 (
		_w582_,
		_w566_,
		_w3392_,
		_w3393_
	);
	LUT4 #(
		.INIT('hdc8c)
	) name2941 (
		\DataWidth_reg[1]/NET0131 ,
		\EBX_reg[4]/NET0131 ,
		_w645_,
		_w3390_,
		_w3394_
	);
	LUT3 #(
		.INIT('h20)
	) name2942 (
		_w589_,
		_w566_,
		_w3394_,
		_w3395_
	);
	LUT4 #(
		.INIT('h000d)
	) name2943 (
		\rEIP_reg[4]/NET0131 ,
		_w3110_,
		_w3393_,
		_w3395_,
		_w3396_
	);
	LUT2 #(
		.INIT('h2)
	) name2944 (
		\rEIP_reg[4]/NET0131 ,
		_w3101_,
		_w3397_
	);
	LUT3 #(
		.INIT('h07)
	) name2945 (
		\PhyAddrPointer_reg[4]/NET0131 ,
		_w706_,
		_w1080_,
		_w3398_
	);
	LUT2 #(
		.INIT('h4)
	) name2946 (
		_w3397_,
		_w3398_,
		_w3399_
	);
	LUT3 #(
		.INIT('hd0)
	) name2947 (
		_w690_,
		_w3396_,
		_w3399_,
		_w3400_
	);
	LUT3 #(
		.INIT('h4f)
	) name2948 (
		_w3386_,
		_w3388_,
		_w3400_,
		_w3401_
	);
	LUT3 #(
		.INIT('hec)
	) name2949 (
		_w1190_,
		_w1214_,
		_w3331_,
		_w3402_
	);
	LUT2 #(
		.INIT('h2)
	) name2950 (
		\DataWidth_reg[1]/NET0131 ,
		\rEIP_reg[5]/NET0131 ,
		_w3403_
	);
	LUT2 #(
		.INIT('h2)
	) name2951 (
		_w695_,
		_w3403_,
		_w3404_
	);
	LUT4 #(
		.INIT('heb00)
	) name2952 (
		\DataWidth_reg[1]/NET0131 ,
		_w2131_,
		_w3402_,
		_w3404_,
		_w3405_
	);
	LUT3 #(
		.INIT('h8a)
	) name2953 (
		\EBX_reg[31]/NET0131 ,
		\EBX_reg[4]/NET0131 ,
		_w3139_,
		_w3406_
	);
	LUT4 #(
		.INIT('h0110)
	) name2954 (
		\DataWidth_reg[1]/NET0131 ,
		READY_n_pad,
		\rEIP_reg[5]/NET0131 ,
		_w3148_,
		_w3407_
	);
	LUT4 #(
		.INIT('h00ed)
	) name2955 (
		\EBX_reg[5]/NET0131 ,
		_w3116_,
		_w3406_,
		_w3407_,
		_w3408_
	);
	LUT3 #(
		.INIT('h02)
	) name2956 (
		_w582_,
		_w566_,
		_w3408_,
		_w3409_
	);
	LUT3 #(
		.INIT('h8c)
	) name2957 (
		\DataWidth_reg[1]/NET0131 ,
		\EBX_reg[5]/NET0131 ,
		_w645_,
		_w3410_
	);
	LUT4 #(
		.INIT('h1040)
	) name2958 (
		\DataWidth_reg[1]/NET0131 ,
		\rEIP_reg[5]/NET0131 ,
		_w645_,
		_w3148_,
		_w3411_
	);
	LUT2 #(
		.INIT('h1)
	) name2959 (
		_w3410_,
		_w3411_,
		_w3412_
	);
	LUT3 #(
		.INIT('h02)
	) name2960 (
		_w589_,
		_w566_,
		_w3412_,
		_w3413_
	);
	LUT4 #(
		.INIT('h000d)
	) name2961 (
		\rEIP_reg[5]/NET0131 ,
		_w3110_,
		_w3409_,
		_w3413_,
		_w3414_
	);
	LUT2 #(
		.INIT('h2)
	) name2962 (
		\rEIP_reg[5]/NET0131 ,
		_w3101_,
		_w3415_
	);
	LUT3 #(
		.INIT('h07)
	) name2963 (
		\PhyAddrPointer_reg[5]/NET0131 ,
		_w706_,
		_w1080_,
		_w3416_
	);
	LUT2 #(
		.INIT('h4)
	) name2964 (
		_w3415_,
		_w3416_,
		_w3417_
	);
	LUT3 #(
		.INIT('hd0)
	) name2965 (
		_w690_,
		_w3414_,
		_w3417_,
		_w3418_
	);
	LUT2 #(
		.INIT('hb)
	) name2966 (
		_w3405_,
		_w3418_,
		_w3419_
	);
	LUT3 #(
		.INIT('h40)
	) name2967 (
		\PhyAddrPointer_reg[0]/NET0131 ,
		\PhyAddrPointer_reg[1]/NET0131 ,
		_w1191_,
		_w3420_
	);
	LUT4 #(
		.INIT('h0514)
	) name2968 (
		\DataWidth_reg[1]/NET0131 ,
		_w1214_,
		_w2142_,
		_w3420_,
		_w3421_
	);
	LUT2 #(
		.INIT('h2)
	) name2969 (
		\DataWidth_reg[1]/NET0131 ,
		\rEIP_reg[6]/NET0131 ,
		_w3422_
	);
	LUT2 #(
		.INIT('h2)
	) name2970 (
		_w695_,
		_w3422_,
		_w3423_
	);
	LUT3 #(
		.INIT('h6c)
	) name2971 (
		\rEIP_reg[5]/NET0131 ,
		\rEIP_reg[6]/NET0131 ,
		_w3148_,
		_w3424_
	);
	LUT3 #(
		.INIT('he2)
	) name2972 (
		\EBX_reg[6]/NET0131 ,
		_w688_,
		_w3424_,
		_w3425_
	);
	LUT3 #(
		.INIT('h20)
	) name2973 (
		_w589_,
		_w566_,
		_w3425_,
		_w3426_
	);
	LUT4 #(
		.INIT('h9030)
	) name2974 (
		\rEIP_reg[5]/NET0131 ,
		\rEIP_reg[6]/NET0131 ,
		_w3116_,
		_w3148_,
		_w3427_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name2975 (
		\EBX_reg[31]/NET0131 ,
		\EBX_reg[4]/NET0131 ,
		\EBX_reg[5]/NET0131 ,
		_w3139_,
		_w3428_
	);
	LUT4 #(
		.INIT('h0d0e)
	) name2976 (
		\EBX_reg[6]/NET0131 ,
		_w3116_,
		_w3427_,
		_w3428_,
		_w3429_
	);
	LUT3 #(
		.INIT('h20)
	) name2977 (
		_w582_,
		_w566_,
		_w3429_,
		_w3430_
	);
	LUT4 #(
		.INIT('h000d)
	) name2978 (
		\rEIP_reg[6]/NET0131 ,
		_w3110_,
		_w3426_,
		_w3430_,
		_w3431_
	);
	LUT2 #(
		.INIT('h2)
	) name2979 (
		\rEIP_reg[6]/NET0131 ,
		_w3101_,
		_w3432_
	);
	LUT3 #(
		.INIT('h07)
	) name2980 (
		\PhyAddrPointer_reg[6]/NET0131 ,
		_w706_,
		_w1080_,
		_w3433_
	);
	LUT2 #(
		.INIT('h4)
	) name2981 (
		_w3432_,
		_w3433_,
		_w3434_
	);
	LUT3 #(
		.INIT('hd0)
	) name2982 (
		_w690_,
		_w3431_,
		_w3434_,
		_w3435_
	);
	LUT3 #(
		.INIT('h4f)
	) name2983 (
		_w3421_,
		_w3423_,
		_w3435_,
		_w3436_
	);
	LUT3 #(
		.INIT('hec)
	) name2984 (
		_w1192_,
		_w1214_,
		_w3331_,
		_w3437_
	);
	LUT2 #(
		.INIT('h2)
	) name2985 (
		\DataWidth_reg[1]/NET0131 ,
		\rEIP_reg[7]/NET0131 ,
		_w3438_
	);
	LUT2 #(
		.INIT('h2)
	) name2986 (
		_w695_,
		_w3438_,
		_w3439_
	);
	LUT4 #(
		.INIT('heb00)
	) name2987 (
		\DataWidth_reg[1]/NET0131 ,
		_w1868_,
		_w3437_,
		_w3439_,
		_w3440_
	);
	LUT2 #(
		.INIT('h2)
	) name2988 (
		\rEIP_reg[7]/NET0131 ,
		_w3110_,
		_w3441_
	);
	LUT4 #(
		.INIT('h78f0)
	) name2989 (
		\rEIP_reg[5]/NET0131 ,
		\rEIP_reg[6]/NET0131 ,
		\rEIP_reg[7]/NET0131 ,
		_w3148_,
		_w3442_
	);
	LUT3 #(
		.INIT('he2)
	) name2990 (
		\EBX_reg[7]/NET0131 ,
		_w688_,
		_w3442_,
		_w3443_
	);
	LUT2 #(
		.INIT('h8)
	) name2991 (
		_w589_,
		_w3443_,
		_w3444_
	);
	LUT4 #(
		.INIT('h0309)
	) name2992 (
		\EBX_reg[31]/NET0131 ,
		\EBX_reg[7]/NET0131 ,
		_w3116_,
		_w3140_,
		_w3445_
	);
	LUT2 #(
		.INIT('h2)
	) name2993 (
		_w3116_,
		_w3442_,
		_w3446_
	);
	LUT3 #(
		.INIT('h02)
	) name2994 (
		_w582_,
		_w3446_,
		_w3445_,
		_w3447_
	);
	LUT3 #(
		.INIT('h54)
	) name2995 (
		_w566_,
		_w3444_,
		_w3447_,
		_w3448_
	);
	LUT2 #(
		.INIT('h2)
	) name2996 (
		\rEIP_reg[7]/NET0131 ,
		_w3101_,
		_w3449_
	);
	LUT3 #(
		.INIT('h07)
	) name2997 (
		\PhyAddrPointer_reg[7]/NET0131 ,
		_w706_,
		_w1080_,
		_w3450_
	);
	LUT2 #(
		.INIT('h4)
	) name2998 (
		_w3449_,
		_w3450_,
		_w3451_
	);
	LUT4 #(
		.INIT('h5700)
	) name2999 (
		_w690_,
		_w3441_,
		_w3448_,
		_w3451_,
		_w3452_
	);
	LUT2 #(
		.INIT('hb)
	) name3000 (
		_w3440_,
		_w3452_,
		_w3453_
	);
	LUT4 #(
		.INIT('h0514)
	) name3001 (
		\DataWidth_reg[1]/NET0131 ,
		_w1214_,
		_w1696_,
		_w3129_,
		_w3454_
	);
	LUT2 #(
		.INIT('h2)
	) name3002 (
		\DataWidth_reg[1]/NET0131 ,
		\rEIP_reg[8]/NET0131 ,
		_w3455_
	);
	LUT2 #(
		.INIT('h2)
	) name3003 (
		_w695_,
		_w3455_,
		_w3456_
	);
	LUT4 #(
		.INIT('h3aca)
	) name3004 (
		\EBX_reg[8]/NET0131 ,
		\rEIP_reg[8]/NET0131 ,
		_w688_,
		_w3149_,
		_w3457_
	);
	LUT3 #(
		.INIT('h20)
	) name3005 (
		_w589_,
		_w566_,
		_w3457_,
		_w3458_
	);
	LUT3 #(
		.INIT('h8a)
	) name3006 (
		\EBX_reg[31]/NET0131 ,
		\EBX_reg[7]/NET0131 ,
		_w3140_,
		_w3459_
	);
	LUT3 #(
		.INIT('h21)
	) name3007 (
		\EBX_reg[8]/NET0131 ,
		_w3116_,
		_w3459_,
		_w3460_
	);
	LUT3 #(
		.INIT('h84)
	) name3008 (
		\rEIP_reg[8]/NET0131 ,
		_w3116_,
		_w3149_,
		_w3461_
	);
	LUT4 #(
		.INIT('h0002)
	) name3009 (
		_w582_,
		_w566_,
		_w3461_,
		_w3460_,
		_w3462_
	);
	LUT4 #(
		.INIT('h000d)
	) name3010 (
		\rEIP_reg[8]/NET0131 ,
		_w3110_,
		_w3458_,
		_w3462_,
		_w3463_
	);
	LUT2 #(
		.INIT('h2)
	) name3011 (
		\rEIP_reg[8]/NET0131 ,
		_w3101_,
		_w3464_
	);
	LUT3 #(
		.INIT('h07)
	) name3012 (
		\PhyAddrPointer_reg[8]/NET0131 ,
		_w706_,
		_w1080_,
		_w3465_
	);
	LUT2 #(
		.INIT('h4)
	) name3013 (
		_w3464_,
		_w3465_,
		_w3466_
	);
	LUT3 #(
		.INIT('hd0)
	) name3014 (
		_w690_,
		_w3463_,
		_w3466_,
		_w3467_
	);
	LUT3 #(
		.INIT('h4f)
	) name3015 (
		_w3454_,
		_w3456_,
		_w3467_,
		_w3468_
	);
	LUT3 #(
		.INIT('h40)
	) name3016 (
		\PhyAddrPointer_reg[0]/NET0131 ,
		\PhyAddrPointer_reg[8]/NET0131 ,
		_w1386_,
		_w3469_
	);
	LUT4 #(
		.INIT('h0514)
	) name3017 (
		\DataWidth_reg[1]/NET0131 ,
		_w1214_,
		_w1878_,
		_w3469_,
		_w3470_
	);
	LUT2 #(
		.INIT('h2)
	) name3018 (
		\DataWidth_reg[1]/NET0131 ,
		\rEIP_reg[9]/NET0131 ,
		_w3471_
	);
	LUT2 #(
		.INIT('h2)
	) name3019 (
		_w695_,
		_w3471_,
		_w3472_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name3020 (
		\EBX_reg[31]/NET0131 ,
		\EBX_reg[7]/NET0131 ,
		\EBX_reg[8]/NET0131 ,
		_w3140_,
		_w3473_
	);
	LUT3 #(
		.INIT('h12)
	) name3021 (
		\EBX_reg[9]/NET0131 ,
		_w3116_,
		_w3473_,
		_w3474_
	);
	LUT4 #(
		.INIT('h1450)
	) name3022 (
		\DataWidth_reg[1]/NET0131 ,
		\rEIP_reg[8]/NET0131 ,
		\rEIP_reg[9]/NET0131 ,
		_w3149_,
		_w3475_
	);
	LUT2 #(
		.INIT('h4)
	) name3023 (
		READY_n_pad,
		_w3475_,
		_w3476_
	);
	LUT2 #(
		.INIT('h1)
	) name3024 (
		_w3474_,
		_w3476_,
		_w3477_
	);
	LUT3 #(
		.INIT('h02)
	) name3025 (
		_w582_,
		_w566_,
		_w3477_,
		_w3478_
	);
	LUT3 #(
		.INIT('h8c)
	) name3026 (
		\DataWidth_reg[1]/NET0131 ,
		\EBX_reg[9]/NET0131 ,
		_w645_,
		_w3479_
	);
	LUT3 #(
		.INIT('h07)
	) name3027 (
		_w645_,
		_w3475_,
		_w3479_,
		_w3480_
	);
	LUT3 #(
		.INIT('h02)
	) name3028 (
		_w589_,
		_w566_,
		_w3480_,
		_w3481_
	);
	LUT4 #(
		.INIT('h000d)
	) name3029 (
		\rEIP_reg[9]/NET0131 ,
		_w3110_,
		_w3478_,
		_w3481_,
		_w3482_
	);
	LUT2 #(
		.INIT('h2)
	) name3030 (
		\rEIP_reg[9]/NET0131 ,
		_w3101_,
		_w3483_
	);
	LUT3 #(
		.INIT('h07)
	) name3031 (
		\PhyAddrPointer_reg[9]/NET0131 ,
		_w706_,
		_w1080_,
		_w3484_
	);
	LUT2 #(
		.INIT('h4)
	) name3032 (
		_w3483_,
		_w3484_,
		_w3485_
	);
	LUT3 #(
		.INIT('hd0)
	) name3033 (
		_w690_,
		_w3482_,
		_w3485_,
		_w3486_
	);
	LUT3 #(
		.INIT('h4f)
	) name3034 (
		_w3470_,
		_w3472_,
		_w3486_,
		_w3487_
	);
	LUT4 #(
		.INIT('h000d)
	) name3035 (
		\PhyAddrPointer_reg[1]/NET0131 ,
		_w1634_,
		_w2054_,
		_w2056_,
		_w3488_
	);
	LUT4 #(
		.INIT('h80cc)
	) name3036 (
		\DataWidth_reg[1]/NET0131 ,
		\PhyAddrPointer_reg[1]/NET0131 ,
		_w695_,
		_w1215_,
		_w3489_
	);
	LUT4 #(
		.INIT('h3310)
	) name3037 (
		\DataWidth_reg[1]/NET0131 ,
		\PhyAddrPointer_reg[1]/NET0131 ,
		_w695_,
		_w1212_,
		_w3490_
	);
	LUT3 #(
		.INIT('h01)
	) name3038 (
		_w2060_,
		_w3490_,
		_w3489_,
		_w3491_
	);
	LUT3 #(
		.INIT('h2f)
	) name3039 (
		_w690_,
		_w3488_,
		_w3491_,
		_w3492_
	);
	LUT4 #(
		.INIT('h4000)
	) name3040 (
		\PhyAddrPointer_reg[0]/NET0131 ,
		\PhyAddrPointer_reg[8]/NET0131 ,
		\PhyAddrPointer_reg[9]/NET0131 ,
		_w1386_,
		_w3493_
	);
	LUT4 #(
		.INIT('h0514)
	) name3041 (
		\DataWidth_reg[1]/NET0131 ,
		_w1214_,
		_w1860_,
		_w3493_,
		_w3494_
	);
	LUT2 #(
		.INIT('h2)
	) name3042 (
		\DataWidth_reg[1]/NET0131 ,
		\rEIP_reg[10]/NET0131 ,
		_w3495_
	);
	LUT2 #(
		.INIT('h2)
	) name3043 (
		_w695_,
		_w3495_,
		_w3496_
	);
	LUT4 #(
		.INIT('h0100)
	) name3044 (
		\EBX_reg[7]/NET0131 ,
		\EBX_reg[8]/NET0131 ,
		\EBX_reg[9]/NET0131 ,
		_w3140_,
		_w3497_
	);
	LUT4 #(
		.INIT('h0509)
	) name3045 (
		\EBX_reg[10]/NET0131 ,
		\EBX_reg[31]/NET0131 ,
		_w3116_,
		_w3497_,
		_w3498_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name3046 (
		\rEIP_reg[10]/NET0131 ,
		\rEIP_reg[8]/NET0131 ,
		\rEIP_reg[9]/NET0131 ,
		_w3149_,
		_w3499_
	);
	LUT2 #(
		.INIT('h2)
	) name3047 (
		_w3116_,
		_w3499_,
		_w3500_
	);
	LUT4 #(
		.INIT('h0002)
	) name3048 (
		_w582_,
		_w566_,
		_w3500_,
		_w3498_,
		_w3501_
	);
	LUT2 #(
		.INIT('h2)
	) name3049 (
		_w688_,
		_w3499_,
		_w3502_
	);
	LUT3 #(
		.INIT('h23)
	) name3050 (
		\DataWidth_reg[1]/NET0131 ,
		\EBX_reg[10]/NET0131 ,
		_w645_,
		_w3503_
	);
	LUT4 #(
		.INIT('h0002)
	) name3051 (
		_w589_,
		_w566_,
		_w3503_,
		_w3502_,
		_w3504_
	);
	LUT4 #(
		.INIT('h000d)
	) name3052 (
		\rEIP_reg[10]/NET0131 ,
		_w3110_,
		_w3504_,
		_w3501_,
		_w3505_
	);
	LUT2 #(
		.INIT('h2)
	) name3053 (
		\rEIP_reg[10]/NET0131 ,
		_w3101_,
		_w3506_
	);
	LUT3 #(
		.INIT('h07)
	) name3054 (
		\PhyAddrPointer_reg[10]/NET0131 ,
		_w706_,
		_w1080_,
		_w3507_
	);
	LUT2 #(
		.INIT('h4)
	) name3055 (
		_w3506_,
		_w3507_,
		_w3508_
	);
	LUT3 #(
		.INIT('hd0)
	) name3056 (
		_w690_,
		_w3505_,
		_w3508_,
		_w3509_
	);
	LUT3 #(
		.INIT('h4f)
	) name3057 (
		_w3494_,
		_w3496_,
		_w3509_,
		_w3510_
	);
	LUT3 #(
		.INIT('h40)
	) name3058 (
		\PhyAddrPointer_reg[0]/NET0131 ,
		_w1386_,
		_w2008_,
		_w3511_
	);
	LUT2 #(
		.INIT('h8)
	) name3059 (
		_w1195_,
		_w3511_,
		_w3512_
	);
	LUT4 #(
		.INIT('h0514)
	) name3060 (
		\DataWidth_reg[1]/NET0131 ,
		_w1214_,
		_w1492_,
		_w3512_,
		_w3513_
	);
	LUT2 #(
		.INIT('h2)
	) name3061 (
		\DataWidth_reg[1]/NET0131 ,
		\rEIP_reg[11]/NET0131 ,
		_w3514_
	);
	LUT2 #(
		.INIT('h2)
	) name3062 (
		_w695_,
		_w3514_,
		_w3515_
	);
	LUT4 #(
		.INIT('h0509)
	) name3063 (
		\EBX_reg[11]/NET0131 ,
		\EBX_reg[31]/NET0131 ,
		_w3116_,
		_w3142_,
		_w3516_
	);
	LUT3 #(
		.INIT('h84)
	) name3064 (
		\rEIP_reg[11]/NET0131 ,
		_w3116_,
		_w3150_,
		_w3517_
	);
	LUT4 #(
		.INIT('h0002)
	) name3065 (
		_w582_,
		_w566_,
		_w3517_,
		_w3516_,
		_w3518_
	);
	LUT3 #(
		.INIT('h84)
	) name3066 (
		\rEIP_reg[11]/NET0131 ,
		_w688_,
		_w3150_,
		_w3519_
	);
	LUT3 #(
		.INIT('h23)
	) name3067 (
		\DataWidth_reg[1]/NET0131 ,
		\EBX_reg[11]/NET0131 ,
		_w645_,
		_w3520_
	);
	LUT4 #(
		.INIT('h0002)
	) name3068 (
		_w589_,
		_w566_,
		_w3520_,
		_w3519_,
		_w3521_
	);
	LUT4 #(
		.INIT('h000d)
	) name3069 (
		\rEIP_reg[11]/NET0131 ,
		_w3110_,
		_w3521_,
		_w3518_,
		_w3522_
	);
	LUT2 #(
		.INIT('h2)
	) name3070 (
		\rEIP_reg[11]/NET0131 ,
		_w3101_,
		_w3523_
	);
	LUT3 #(
		.INIT('h07)
	) name3071 (
		\PhyAddrPointer_reg[11]/NET0131 ,
		_w706_,
		_w1080_,
		_w3524_
	);
	LUT2 #(
		.INIT('h4)
	) name3072 (
		_w3523_,
		_w3524_,
		_w3525_
	);
	LUT3 #(
		.INIT('hd0)
	) name3073 (
		_w690_,
		_w3522_,
		_w3525_,
		_w3526_
	);
	LUT3 #(
		.INIT('h4f)
	) name3074 (
		_w3513_,
		_w3515_,
		_w3526_,
		_w3527_
	);
	LUT3 #(
		.INIT('h6a)
	) name3075 (
		\PhyAddrPointer_reg[12]/NET0131 ,
		\PhyAddrPointer_reg[1]/NET0131 ,
		_w1491_,
		_w3528_
	);
	LUT2 #(
		.INIT('h8)
	) name3076 (
		_w1491_,
		_w3511_,
		_w3529_
	);
	LUT4 #(
		.INIT('h0514)
	) name3077 (
		\DataWidth_reg[1]/NET0131 ,
		_w1214_,
		_w3528_,
		_w3529_,
		_w3530_
	);
	LUT2 #(
		.INIT('h2)
	) name3078 (
		\DataWidth_reg[1]/NET0131 ,
		\rEIP_reg[12]/NET0131 ,
		_w3531_
	);
	LUT2 #(
		.INIT('h2)
	) name3079 (
		_w695_,
		_w3531_,
		_w3532_
	);
	LUT2 #(
		.INIT('h2)
	) name3080 (
		\rEIP_reg[12]/NET0131 ,
		_w3110_,
		_w3533_
	);
	LUT4 #(
		.INIT('h9030)
	) name3081 (
		\rEIP_reg[11]/NET0131 ,
		\rEIP_reg[12]/NET0131 ,
		_w688_,
		_w3150_,
		_w3534_
	);
	LUT3 #(
		.INIT('h23)
	) name3082 (
		\DataWidth_reg[1]/NET0131 ,
		\EBX_reg[12]/NET0131 ,
		_w645_,
		_w3535_
	);
	LUT3 #(
		.INIT('h02)
	) name3083 (
		_w589_,
		_w3535_,
		_w3534_,
		_w3536_
	);
	LUT3 #(
		.INIT('h8c)
	) name3084 (
		\EBX_reg[11]/NET0131 ,
		\EBX_reg[31]/NET0131 ,
		_w3142_,
		_w3537_
	);
	LUT3 #(
		.INIT('h21)
	) name3085 (
		\EBX_reg[12]/NET0131 ,
		_w3116_,
		_w3537_,
		_w3538_
	);
	LUT4 #(
		.INIT('h9030)
	) name3086 (
		\rEIP_reg[11]/NET0131 ,
		\rEIP_reg[12]/NET0131 ,
		_w3116_,
		_w3150_,
		_w3539_
	);
	LUT3 #(
		.INIT('h02)
	) name3087 (
		_w582_,
		_w3539_,
		_w3538_,
		_w3540_
	);
	LUT3 #(
		.INIT('h54)
	) name3088 (
		_w566_,
		_w3536_,
		_w3540_,
		_w3541_
	);
	LUT2 #(
		.INIT('h2)
	) name3089 (
		\rEIP_reg[12]/NET0131 ,
		_w3101_,
		_w3542_
	);
	LUT3 #(
		.INIT('h07)
	) name3090 (
		\PhyAddrPointer_reg[12]/NET0131 ,
		_w706_,
		_w1080_,
		_w3543_
	);
	LUT2 #(
		.INIT('h4)
	) name3091 (
		_w3542_,
		_w3543_,
		_w3544_
	);
	LUT4 #(
		.INIT('h5700)
	) name3092 (
		_w690_,
		_w3533_,
		_w3541_,
		_w3544_,
		_w3545_
	);
	LUT3 #(
		.INIT('h4f)
	) name3093 (
		_w3530_,
		_w3532_,
		_w3545_,
		_w3546_
	);
	LUT3 #(
		.INIT('hea)
	) name3094 (
		_w1214_,
		_w1602_,
		_w3129_,
		_w3547_
	);
	LUT2 #(
		.INIT('h2)
	) name3095 (
		\DataWidth_reg[1]/NET0131 ,
		\rEIP_reg[13]/NET0131 ,
		_w3548_
	);
	LUT2 #(
		.INIT('h2)
	) name3096 (
		_w695_,
		_w3548_,
		_w3549_
	);
	LUT4 #(
		.INIT('heb00)
	) name3097 (
		\DataWidth_reg[1]/NET0131 ,
		_w1600_,
		_w3547_,
		_w3549_,
		_w3550_
	);
	LUT2 #(
		.INIT('h2)
	) name3098 (
		\rEIP_reg[13]/NET0131 ,
		_w3110_,
		_w3551_
	);
	LUT4 #(
		.INIT('h78f0)
	) name3099 (
		\rEIP_reg[11]/NET0131 ,
		\rEIP_reg[12]/NET0131 ,
		\rEIP_reg[13]/NET0131 ,
		_w3150_,
		_w3552_
	);
	LUT2 #(
		.INIT('h2)
	) name3100 (
		_w688_,
		_w3552_,
		_w3553_
	);
	LUT3 #(
		.INIT('h23)
	) name3101 (
		\DataWidth_reg[1]/NET0131 ,
		\EBX_reg[13]/NET0131 ,
		_w645_,
		_w3554_
	);
	LUT3 #(
		.INIT('h02)
	) name3102 (
		_w589_,
		_w3554_,
		_w3553_,
		_w3555_
	);
	LUT3 #(
		.INIT('h2a)
	) name3103 (
		\EBX_reg[31]/NET0131 ,
		_w3142_,
		_w3143_,
		_w3556_
	);
	LUT3 #(
		.INIT('h21)
	) name3104 (
		\EBX_reg[13]/NET0131 ,
		_w3116_,
		_w3556_,
		_w3557_
	);
	LUT2 #(
		.INIT('h2)
	) name3105 (
		_w3116_,
		_w3552_,
		_w3558_
	);
	LUT3 #(
		.INIT('h02)
	) name3106 (
		_w582_,
		_w3558_,
		_w3557_,
		_w3559_
	);
	LUT3 #(
		.INIT('h54)
	) name3107 (
		_w566_,
		_w3555_,
		_w3559_,
		_w3560_
	);
	LUT2 #(
		.INIT('h2)
	) name3108 (
		\rEIP_reg[13]/NET0131 ,
		_w3101_,
		_w3561_
	);
	LUT3 #(
		.INIT('h07)
	) name3109 (
		\PhyAddrPointer_reg[13]/NET0131 ,
		_w706_,
		_w1080_,
		_w3562_
	);
	LUT2 #(
		.INIT('h4)
	) name3110 (
		_w3561_,
		_w3562_,
		_w3563_
	);
	LUT4 #(
		.INIT('h5700)
	) name3111 (
		_w690_,
		_w3551_,
		_w3560_,
		_w3563_,
		_w3564_
	);
	LUT2 #(
		.INIT('hb)
	) name3112 (
		_w3550_,
		_w3564_,
		_w3565_
	);
	LUT2 #(
		.INIT('h8)
	) name3113 (
		_w1198_,
		_w3511_,
		_w3566_
	);
	LUT4 #(
		.INIT('h0514)
	) name3114 (
		\DataWidth_reg[1]/NET0131 ,
		_w1214_,
		_w1501_,
		_w3566_,
		_w3567_
	);
	LUT2 #(
		.INIT('h2)
	) name3115 (
		\DataWidth_reg[1]/NET0131 ,
		\rEIP_reg[14]/NET0131 ,
		_w3568_
	);
	LUT2 #(
		.INIT('h2)
	) name3116 (
		_w695_,
		_w3568_,
		_w3569_
	);
	LUT2 #(
		.INIT('h2)
	) name3117 (
		\rEIP_reg[14]/NET0131 ,
		_w3110_,
		_w3570_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name3118 (
		\rEIP_reg[11]/NET0131 ,
		\rEIP_reg[14]/NET0131 ,
		_w3150_,
		_w3151_,
		_w3571_
	);
	LUT2 #(
		.INIT('h2)
	) name3119 (
		_w688_,
		_w3571_,
		_w3572_
	);
	LUT3 #(
		.INIT('h23)
	) name3120 (
		\DataWidth_reg[1]/NET0131 ,
		\EBX_reg[14]/NET0131 ,
		_w645_,
		_w3573_
	);
	LUT3 #(
		.INIT('h02)
	) name3121 (
		_w589_,
		_w3573_,
		_w3572_,
		_w3574_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name3122 (
		\EBX_reg[13]/NET0131 ,
		\EBX_reg[31]/NET0131 ,
		_w3142_,
		_w3143_,
		_w3575_
	);
	LUT3 #(
		.INIT('h21)
	) name3123 (
		\EBX_reg[14]/NET0131 ,
		_w3116_,
		_w3575_,
		_w3576_
	);
	LUT2 #(
		.INIT('h2)
	) name3124 (
		_w3116_,
		_w3571_,
		_w3577_
	);
	LUT3 #(
		.INIT('h02)
	) name3125 (
		_w582_,
		_w3577_,
		_w3576_,
		_w3578_
	);
	LUT3 #(
		.INIT('h54)
	) name3126 (
		_w566_,
		_w3574_,
		_w3578_,
		_w3579_
	);
	LUT2 #(
		.INIT('h2)
	) name3127 (
		\rEIP_reg[14]/NET0131 ,
		_w3101_,
		_w3580_
	);
	LUT3 #(
		.INIT('h07)
	) name3128 (
		\PhyAddrPointer_reg[14]/NET0131 ,
		_w706_,
		_w1080_,
		_w3581_
	);
	LUT2 #(
		.INIT('h4)
	) name3129 (
		_w3580_,
		_w3581_,
		_w3582_
	);
	LUT4 #(
		.INIT('h5700)
	) name3130 (
		_w690_,
		_w3570_,
		_w3579_,
		_w3582_,
		_w3583_
	);
	LUT3 #(
		.INIT('h4f)
	) name3131 (
		_w3567_,
		_w3569_,
		_w3583_,
		_w3584_
	);
	LUT2 #(
		.INIT('h4)
	) name3132 (
		_w1501_,
		_w3566_,
		_w3585_
	);
	LUT4 #(
		.INIT('h0514)
	) name3133 (
		\DataWidth_reg[1]/NET0131 ,
		_w1214_,
		_w1390_,
		_w3585_,
		_w3586_
	);
	LUT2 #(
		.INIT('h2)
	) name3134 (
		\DataWidth_reg[1]/NET0131 ,
		\rEIP_reg[15]/NET0131 ,
		_w3587_
	);
	LUT2 #(
		.INIT('h2)
	) name3135 (
		_w695_,
		_w3587_,
		_w3588_
	);
	LUT2 #(
		.INIT('h2)
	) name3136 (
		\rEIP_reg[15]/NET0131 ,
		_w3110_,
		_w3589_
	);
	LUT3 #(
		.INIT('h23)
	) name3137 (
		\DataWidth_reg[1]/NET0131 ,
		\EBX_reg[15]/NET0131 ,
		_w645_,
		_w3590_
	);
	LUT4 #(
		.INIT('h0509)
	) name3138 (
		\EBX_reg[15]/NET0131 ,
		\EBX_reg[31]/NET0131 ,
		_w3116_,
		_w3144_,
		_w3591_
	);
	LUT4 #(
		.INIT('hf351)
	) name3139 (
		_w582_,
		_w589_,
		_w3590_,
		_w3591_,
		_w3592_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name3140 (
		\rEIP_reg[11]/NET0131 ,
		\rEIP_reg[15]/NET0131 ,
		_w3150_,
		_w3152_,
		_w3593_
	);
	LUT4 #(
		.INIT('hf070)
	) name3141 (
		_w589_,
		_w594_,
		_w3116_,
		_w3590_,
		_w3594_
	);
	LUT4 #(
		.INIT('h1011)
	) name3142 (
		_w566_,
		_w3592_,
		_w3593_,
		_w3594_,
		_w3595_
	);
	LUT2 #(
		.INIT('h2)
	) name3143 (
		\rEIP_reg[15]/NET0131 ,
		_w3101_,
		_w3596_
	);
	LUT3 #(
		.INIT('h07)
	) name3144 (
		\PhyAddrPointer_reg[15]/NET0131 ,
		_w706_,
		_w1080_,
		_w3597_
	);
	LUT2 #(
		.INIT('h4)
	) name3145 (
		_w3596_,
		_w3597_,
		_w3598_
	);
	LUT4 #(
		.INIT('h5700)
	) name3146 (
		_w690_,
		_w3589_,
		_w3595_,
		_w3598_,
		_w3599_
	);
	LUT3 #(
		.INIT('h4f)
	) name3147 (
		_w3586_,
		_w3588_,
		_w3599_,
		_w3600_
	);
	LUT3 #(
		.INIT('hba)
	) name3148 (
		_w1214_,
		_w1390_,
		_w3585_,
		_w3601_
	);
	LUT2 #(
		.INIT('h2)
	) name3149 (
		\DataWidth_reg[1]/NET0131 ,
		\rEIP_reg[16]/NET0131 ,
		_w3602_
	);
	LUT2 #(
		.INIT('h2)
	) name3150 (
		_w695_,
		_w3602_,
		_w3603_
	);
	LUT4 #(
		.INIT('heb00)
	) name3151 (
		\DataWidth_reg[1]/NET0131 ,
		_w1621_,
		_w3601_,
		_w3603_,
		_w3604_
	);
	LUT2 #(
		.INIT('h2)
	) name3152 (
		\rEIP_reg[16]/NET0131 ,
		_w3110_,
		_w3605_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name3153 (
		\rEIP_reg[11]/NET0131 ,
		\rEIP_reg[16]/NET0131 ,
		_w3150_,
		_w3153_,
		_w3606_
	);
	LUT2 #(
		.INIT('h2)
	) name3154 (
		_w688_,
		_w3606_,
		_w3607_
	);
	LUT3 #(
		.INIT('h23)
	) name3155 (
		\DataWidth_reg[1]/NET0131 ,
		\EBX_reg[16]/NET0131 ,
		_w645_,
		_w3608_
	);
	LUT3 #(
		.INIT('h02)
	) name3156 (
		_w589_,
		_w3608_,
		_w3607_,
		_w3609_
	);
	LUT3 #(
		.INIT('h8c)
	) name3157 (
		\EBX_reg[15]/NET0131 ,
		\EBX_reg[31]/NET0131 ,
		_w3144_,
		_w3610_
	);
	LUT3 #(
		.INIT('h21)
	) name3158 (
		\EBX_reg[16]/NET0131 ,
		_w3116_,
		_w3610_,
		_w3611_
	);
	LUT2 #(
		.INIT('h2)
	) name3159 (
		_w3116_,
		_w3606_,
		_w3612_
	);
	LUT2 #(
		.INIT('h2)
	) name3160 (
		_w582_,
		_w3612_,
		_w3613_
	);
	LUT4 #(
		.INIT('h4544)
	) name3161 (
		_w566_,
		_w3609_,
		_w3611_,
		_w3613_,
		_w3614_
	);
	LUT2 #(
		.INIT('h2)
	) name3162 (
		\rEIP_reg[16]/NET0131 ,
		_w3101_,
		_w3615_
	);
	LUT3 #(
		.INIT('h07)
	) name3163 (
		\PhyAddrPointer_reg[16]/NET0131 ,
		_w706_,
		_w1080_,
		_w3616_
	);
	LUT2 #(
		.INIT('h4)
	) name3164 (
		_w3615_,
		_w3616_,
		_w3617_
	);
	LUT4 #(
		.INIT('h5700)
	) name3165 (
		_w690_,
		_w3605_,
		_w3614_,
		_w3617_,
		_w3618_
	);
	LUT2 #(
		.INIT('hb)
	) name3166 (
		_w3604_,
		_w3618_,
		_w3619_
	);
	LUT4 #(
		.INIT('h0514)
	) name3167 (
		\DataWidth_reg[1]/NET0131 ,
		_w1214_,
		_w1640_,
		_w3132_,
		_w3620_
	);
	LUT2 #(
		.INIT('h2)
	) name3168 (
		\DataWidth_reg[1]/NET0131 ,
		\rEIP_reg[17]/NET0131 ,
		_w3621_
	);
	LUT2 #(
		.INIT('h2)
	) name3169 (
		_w695_,
		_w3621_,
		_w3622_
	);
	LUT3 #(
		.INIT('h2a)
	) name3170 (
		\EBX_reg[31]/NET0131 ,
		_w3144_,
		_w3145_,
		_w3623_
	);
	LUT3 #(
		.INIT('hd0)
	) name3171 (
		_w589_,
		_w594_,
		_w3623_,
		_w3624_
	);
	LUT4 #(
		.INIT('h88a8)
	) name3172 (
		\EBX_reg[17]/NET0131 ,
		_w582_,
		_w589_,
		_w594_,
		_w3625_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name3173 (
		\EBX_reg[17]/NET0131 ,
		_w582_,
		_w3116_,
		_w3623_,
		_w3626_
	);
	LUT3 #(
		.INIT('hb0)
	) name3174 (
		_w3624_,
		_w3625_,
		_w3626_,
		_w3627_
	);
	LUT2 #(
		.INIT('h1)
	) name3175 (
		\rEIP_reg[17]/NET0131 ,
		_w3155_,
		_w3628_
	);
	LUT2 #(
		.INIT('h8)
	) name3176 (
		\rEIP_reg[17]/NET0131 ,
		_w3155_,
		_w3629_
	);
	LUT4 #(
		.INIT('h00ae)
	) name3177 (
		_w582_,
		_w589_,
		_w594_,
		_w3629_,
		_w3630_
	);
	LUT4 #(
		.INIT('h1511)
	) name3178 (
		_w566_,
		_w3116_,
		_w3628_,
		_w3630_,
		_w3631_
	);
	LUT4 #(
		.INIT('ha88a)
	) name3179 (
		\EBX_reg[17]/NET0131 ,
		\State_reg[0]/NET0131 ,
		\State_reg[1]/NET0131 ,
		\State_reg[2]/NET0131 ,
		_w3632_
	);
	LUT3 #(
		.INIT('h20)
	) name3180 (
		_w589_,
		_w566_,
		_w3632_,
		_w3633_
	);
	LUT3 #(
		.INIT('h0d)
	) name3181 (
		\rEIP_reg[17]/NET0131 ,
		_w3110_,
		_w3633_,
		_w3634_
	);
	LUT4 #(
		.INIT('h20aa)
	) name3182 (
		_w690_,
		_w3627_,
		_w3631_,
		_w3634_,
		_w3635_
	);
	LUT2 #(
		.INIT('h2)
	) name3183 (
		\rEIP_reg[17]/NET0131 ,
		_w3101_,
		_w3636_
	);
	LUT3 #(
		.INIT('h07)
	) name3184 (
		\PhyAddrPointer_reg[17]/NET0131 ,
		_w706_,
		_w1080_,
		_w3637_
	);
	LUT2 #(
		.INIT('h4)
	) name3185 (
		_w3636_,
		_w3637_,
		_w3638_
	);
	LUT4 #(
		.INIT('hf4ff)
	) name3186 (
		_w3620_,
		_w3622_,
		_w3635_,
		_w3638_,
		_w3639_
	);
	LUT4 #(
		.INIT('h1000)
	) name3187 (
		_w1621_,
		_w1640_,
		_w2008_,
		_w3131_,
		_w3640_
	);
	LUT4 #(
		.INIT('h0514)
	) name3188 (
		\DataWidth_reg[1]/NET0131 ,
		_w1214_,
		_w1657_,
		_w3640_,
		_w3641_
	);
	LUT2 #(
		.INIT('h2)
	) name3189 (
		\DataWidth_reg[1]/NET0131 ,
		\rEIP_reg[18]/NET0131 ,
		_w3642_
	);
	LUT2 #(
		.INIT('h2)
	) name3190 (
		_w695_,
		_w3642_,
		_w3643_
	);
	LUT2 #(
		.INIT('h2)
	) name3191 (
		\rEIP_reg[18]/NET0131 ,
		_w3110_,
		_w3644_
	);
	LUT3 #(
		.INIT('h23)
	) name3192 (
		\DataWidth_reg[1]/NET0131 ,
		\EBX_reg[18]/NET0131 ,
		_w645_,
		_w3645_
	);
	LUT2 #(
		.INIT('h2)
	) name3193 (
		_w589_,
		_w3645_,
		_w3646_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name3194 (
		\EBX_reg[17]/NET0131 ,
		\EBX_reg[31]/NET0131 ,
		_w3144_,
		_w3145_,
		_w3647_
	);
	LUT4 #(
		.INIT('hc4c8)
	) name3195 (
		\EBX_reg[18]/NET0131 ,
		_w582_,
		_w3116_,
		_w3647_,
		_w3648_
	);
	LUT2 #(
		.INIT('h1)
	) name3196 (
		_w3646_,
		_w3648_,
		_w3649_
	);
	LUT3 #(
		.INIT('h6c)
	) name3197 (
		\rEIP_reg[17]/NET0131 ,
		\rEIP_reg[18]/NET0131 ,
		_w3155_,
		_w3650_
	);
	LUT4 #(
		.INIT('hf070)
	) name3198 (
		_w589_,
		_w594_,
		_w3116_,
		_w3645_,
		_w3651_
	);
	LUT3 #(
		.INIT('h45)
	) name3199 (
		_w566_,
		_w3650_,
		_w3651_,
		_w3652_
	);
	LUT4 #(
		.INIT('h8a88)
	) name3200 (
		_w690_,
		_w3644_,
		_w3649_,
		_w3652_,
		_w3653_
	);
	LUT2 #(
		.INIT('h2)
	) name3201 (
		\rEIP_reg[18]/NET0131 ,
		_w3101_,
		_w3654_
	);
	LUT3 #(
		.INIT('h07)
	) name3202 (
		\PhyAddrPointer_reg[18]/NET0131 ,
		_w706_,
		_w1080_,
		_w3655_
	);
	LUT2 #(
		.INIT('h4)
	) name3203 (
		_w3654_,
		_w3655_,
		_w3656_
	);
	LUT4 #(
		.INIT('hf4ff)
	) name3204 (
		_w3641_,
		_w3643_,
		_w3653_,
		_w3656_,
		_w3657_
	);
	LUT3 #(
		.INIT('hba)
	) name3205 (
		_w1214_,
		_w1657_,
		_w3640_,
		_w3658_
	);
	LUT2 #(
		.INIT('h2)
	) name3206 (
		\DataWidth_reg[1]/NET0131 ,
		\rEIP_reg[19]/NET0131 ,
		_w3659_
	);
	LUT2 #(
		.INIT('h2)
	) name3207 (
		_w695_,
		_w3659_,
		_w3660_
	);
	LUT4 #(
		.INIT('heb00)
	) name3208 (
		\DataWidth_reg[1]/NET0131 ,
		_w1521_,
		_w3658_,
		_w3660_,
		_w3661_
	);
	LUT4 #(
		.INIT('h0509)
	) name3209 (
		\EBX_reg[19]/NET0131 ,
		\EBX_reg[31]/NET0131 ,
		_w3116_,
		_w3146_,
		_w3662_
	);
	LUT4 #(
		.INIT('h8444)
	) name3210 (
		\rEIP_reg[19]/NET0131 ,
		_w3116_,
		_w3155_,
		_w3156_,
		_w3663_
	);
	LUT3 #(
		.INIT('h02)
	) name3211 (
		_w582_,
		_w566_,
		_w3663_,
		_w3664_
	);
	LUT2 #(
		.INIT('h4)
	) name3212 (
		_w3662_,
		_w3664_,
		_w3665_
	);
	LUT2 #(
		.INIT('h4)
	) name3213 (
		_w594_,
		_w3663_,
		_w3666_
	);
	LUT3 #(
		.INIT('h23)
	) name3214 (
		\DataWidth_reg[1]/NET0131 ,
		\EBX_reg[19]/NET0131 ,
		_w645_,
		_w3667_
	);
	LUT3 #(
		.INIT('h02)
	) name3215 (
		_w589_,
		_w566_,
		_w3667_,
		_w3668_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name3216 (
		\rEIP_reg[19]/NET0131 ,
		_w3110_,
		_w3666_,
		_w3668_,
		_w3669_
	);
	LUT2 #(
		.INIT('h2)
	) name3217 (
		\rEIP_reg[19]/NET0131 ,
		_w3101_,
		_w3670_
	);
	LUT3 #(
		.INIT('h07)
	) name3218 (
		\PhyAddrPointer_reg[19]/NET0131 ,
		_w706_,
		_w1080_,
		_w3671_
	);
	LUT2 #(
		.INIT('h4)
	) name3219 (
		_w3670_,
		_w3671_,
		_w3672_
	);
	LUT4 #(
		.INIT('h7500)
	) name3220 (
		_w690_,
		_w3665_,
		_w3669_,
		_w3672_,
		_w3673_
	);
	LUT2 #(
		.INIT('hb)
	) name3221 (
		_w3661_,
		_w3673_,
		_w3674_
	);
	LUT3 #(
		.INIT('h04)
	) name3222 (
		\RequestPending_reg/NET0131 ,
		_w563_,
		_w565_,
		_w3675_
	);
	LUT3 #(
		.INIT('h0e)
	) name3223 (
		_w653_,
		_w655_,
		_w3675_,
		_w3676_
	);
	LUT4 #(
		.INIT('h0002)
	) name3224 (
		\RequestPending_reg/NET0131 ,
		_w586_,
		_w582_,
		_w589_,
		_w3677_
	);
	LUT3 #(
		.INIT('h04)
	) name3225 (
		\DataWidth_reg[1]/NET0131 ,
		_w589_,
		_w566_,
		_w3678_
	);
	LUT2 #(
		.INIT('h1)
	) name3226 (
		_w3677_,
		_w3678_,
		_w3679_
	);
	LUT4 #(
		.INIT('hfff4)
	) name3227 (
		\State2_reg[0]/NET0131 ,
		\State2_reg[1]/NET0131 ,
		\State2_reg[2]/NET0131 ,
		\State2_reg[3]/NET0131 ,
		_w3680_
	);
	LUT4 #(
		.INIT('h80aa)
	) name3228 (
		\RequestPending_reg/NET0131 ,
		_w691_,
		_w705_,
		_w1840_,
		_w3681_
	);
	LUT2 #(
		.INIT('h2)
	) name3229 (
		_w3680_,
		_w3681_,
		_w3682_
	);
	LUT4 #(
		.INIT('h8aff)
	) name3230 (
		_w690_,
		_w3676_,
		_w3679_,
		_w3682_,
		_w3683_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name3231 (
		\EAX_reg[18]/NET0131 ,
		\EAX_reg[23]/NET0131 ,
		_w1757_,
		_w2092_,
		_w3684_
	);
	LUT2 #(
		.INIT('h1)
	) name3232 (
		_w594_,
		_w3684_,
		_w3685_
	);
	LUT3 #(
		.INIT('h02)
	) name3233 (
		_w589_,
		_w566_,
		_w3685_,
		_w3686_
	);
	LUT4 #(
		.INIT('haaa2)
	) name3234 (
		\Datao[23]_pad ,
		_w646_,
		_w2183_,
		_w3686_,
		_w3687_
	);
	LUT3 #(
		.INIT('h20)
	) name3235 (
		_w589_,
		_w566_,
		_w3684_,
		_w3688_
	);
	LUT4 #(
		.INIT('h0200)
	) name3236 (
		_w589_,
		_w594_,
		_w566_,
		_w3684_,
		_w3689_
	);
	LUT4 #(
		.INIT('h3f15)
	) name3237 (
		\Datao[23]_pad ,
		\uWord_reg[7]/NET0131 ,
		_w2179_,
		_w2180_,
		_w3690_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name3238 (
		_w690_,
		_w3687_,
		_w3689_,
		_w3690_,
		_w3691_
	);
	LUT3 #(
		.INIT('h6c)
	) name3239 (
		\EAX_reg[18]/NET0131 ,
		\EAX_reg[19]/NET0131 ,
		_w2092_,
		_w3692_
	);
	LUT4 #(
		.INIT('h0903)
	) name3240 (
		\EAX_reg[18]/NET0131 ,
		\EAX_reg[19]/NET0131 ,
		_w594_,
		_w2092_,
		_w3693_
	);
	LUT3 #(
		.INIT('h02)
	) name3241 (
		_w589_,
		_w566_,
		_w3693_,
		_w3694_
	);
	LUT4 #(
		.INIT('haaa2)
	) name3242 (
		\Datao[19]_pad ,
		_w646_,
		_w2183_,
		_w3694_,
		_w3695_
	);
	LUT3 #(
		.INIT('h20)
	) name3243 (
		_w589_,
		_w566_,
		_w3692_,
		_w3696_
	);
	LUT4 #(
		.INIT('h0200)
	) name3244 (
		_w589_,
		_w594_,
		_w566_,
		_w3692_,
		_w3697_
	);
	LUT4 #(
		.INIT('h3f15)
	) name3245 (
		\Datao[19]_pad ,
		\uWord_reg[3]/NET0131 ,
		_w2179_,
		_w2180_,
		_w3698_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name3246 (
		_w690_,
		_w3695_,
		_w3697_,
		_w3698_,
		_w3699_
	);
	LUT4 #(
		.INIT('h2202)
	) name3247 (
		\Datai[2]_pad ,
		READY_n_pad,
		_w563_,
		_w565_,
		_w3700_
	);
	LUT4 #(
		.INIT('hf800)
	) name3248 (
		_w494_,
		_w586_,
		_w582_,
		_w3700_,
		_w3701_
	);
	LUT4 #(
		.INIT('h0080)
	) name3249 (
		_w602_,
		_w604_,
		_w634_,
		_w776_,
		_w3702_
	);
	LUT3 #(
		.INIT('h78)
	) name3250 (
		\EAX_reg[0]/NET0131 ,
		\EAX_reg[1]/NET0131 ,
		\EAX_reg[2]/NET0131 ,
		_w3703_
	);
	LUT3 #(
		.INIT('h80)
	) name3251 (
		_w518_,
		_w617_,
		_w3703_,
		_w3704_
	);
	LUT4 #(
		.INIT('haaa8)
	) name3252 (
		_w690_,
		_w3702_,
		_w3701_,
		_w3704_,
		_w3705_
	);
	LUT3 #(
		.INIT('hf2)
	) name3253 (
		\EAX_reg[2]/NET0131 ,
		_w2643_,
		_w3705_,
		_w3706_
	);
	LUT2 #(
		.INIT('h2)
	) name3254 (
		\uWord_reg[3]/NET0131 ,
		_w1841_,
		_w3707_
	);
	LUT4 #(
		.INIT('h2202)
	) name3255 (
		\Datai[3]_pad ,
		READY_n_pad,
		_w563_,
		_w565_,
		_w3708_
	);
	LUT2 #(
		.INIT('h8)
	) name3256 (
		READY_n_pad,
		\uWord_reg[3]/NET0131 ,
		_w3709_
	);
	LUT2 #(
		.INIT('h1)
	) name3257 (
		_w3708_,
		_w3709_,
		_w3710_
	);
	LUT2 #(
		.INIT('h2)
	) name3258 (
		_w582_,
		_w3710_,
		_w3711_
	);
	LUT4 #(
		.INIT('haa02)
	) name3259 (
		\uWord_reg[3]/NET0131 ,
		_w582_,
		_w589_,
		_w566_,
		_w3712_
	);
	LUT4 #(
		.INIT('haaa8)
	) name3260 (
		_w690_,
		_w3696_,
		_w3711_,
		_w3712_,
		_w3713_
	);
	LUT2 #(
		.INIT('he)
	) name3261 (
		_w3707_,
		_w3713_,
		_w3714_
	);
	LUT2 #(
		.INIT('h2)
	) name3262 (
		\uWord_reg[7]/NET0131 ,
		_w1841_,
		_w3715_
	);
	LUT2 #(
		.INIT('h8)
	) name3263 (
		READY_n_pad,
		\uWord_reg[7]/NET0131 ,
		_w3716_
	);
	LUT2 #(
		.INIT('h1)
	) name3264 (
		_w2644_,
		_w3716_,
		_w3717_
	);
	LUT2 #(
		.INIT('h2)
	) name3265 (
		_w582_,
		_w3717_,
		_w3718_
	);
	LUT4 #(
		.INIT('haa02)
	) name3266 (
		\uWord_reg[7]/NET0131 ,
		_w582_,
		_w589_,
		_w566_,
		_w3719_
	);
	LUT4 #(
		.INIT('haaa8)
	) name3267 (
		_w690_,
		_w3688_,
		_w3718_,
		_w3719_,
		_w3720_
	);
	LUT2 #(
		.INIT('he)
	) name3268 (
		_w3715_,
		_w3720_,
		_w3721_
	);
	LUT4 #(
		.INIT('hf800)
	) name3269 (
		_w494_,
		_w586_,
		_w582_,
		_w3708_,
		_w3722_
	);
	LUT4 #(
		.INIT('h0080)
	) name3270 (
		_w602_,
		_w604_,
		_w634_,
		_w791_,
		_w3723_
	);
	LUT4 #(
		.INIT('h7f80)
	) name3271 (
		\EAX_reg[0]/NET0131 ,
		\EAX_reg[1]/NET0131 ,
		\EAX_reg[2]/NET0131 ,
		\EAX_reg[3]/NET0131 ,
		_w3724_
	);
	LUT3 #(
		.INIT('h80)
	) name3272 (
		_w518_,
		_w617_,
		_w3724_,
		_w3725_
	);
	LUT4 #(
		.INIT('haaa8)
	) name3273 (
		_w690_,
		_w3723_,
		_w3722_,
		_w3725_,
		_w3726_
	);
	LUT3 #(
		.INIT('hf2)
	) name3274 (
		\EAX_reg[3]/NET0131 ,
		_w2643_,
		_w3726_,
		_w3727_
	);
	LUT4 #(
		.INIT('hf800)
	) name3275 (
		_w494_,
		_w586_,
		_w582_,
		_w2442_,
		_w3728_
	);
	LUT4 #(
		.INIT('h0080)
	) name3276 (
		_w602_,
		_w604_,
		_w634_,
		_w761_,
		_w3729_
	);
	LUT2 #(
		.INIT('h6)
	) name3277 (
		\EAX_reg[4]/NET0131 ,
		_w1743_,
		_w3730_
	);
	LUT3 #(
		.INIT('h80)
	) name3278 (
		_w518_,
		_w617_,
		_w3730_,
		_w3731_
	);
	LUT4 #(
		.INIT('haaa8)
	) name3279 (
		_w690_,
		_w3729_,
		_w3728_,
		_w3731_,
		_w3732_
	);
	LUT3 #(
		.INIT('hf2)
	) name3280 (
		\EAX_reg[4]/NET0131 ,
		_w2643_,
		_w3732_,
		_w3733_
	);
	LUT4 #(
		.INIT('h2202)
	) name3281 (
		\Datai[5]_pad ,
		READY_n_pad,
		_w563_,
		_w565_,
		_w3734_
	);
	LUT4 #(
		.INIT('hf800)
	) name3282 (
		_w494_,
		_w586_,
		_w582_,
		_w3734_,
		_w3735_
	);
	LUT4 #(
		.INIT('h0080)
	) name3283 (
		_w602_,
		_w604_,
		_w634_,
		_w866_,
		_w3736_
	);
	LUT3 #(
		.INIT('h6c)
	) name3284 (
		\EAX_reg[4]/NET0131 ,
		\EAX_reg[5]/NET0131 ,
		_w1743_,
		_w3737_
	);
	LUT3 #(
		.INIT('h80)
	) name3285 (
		_w518_,
		_w617_,
		_w3737_,
		_w3738_
	);
	LUT4 #(
		.INIT('haaa8)
	) name3286 (
		_w690_,
		_w3736_,
		_w3735_,
		_w3738_,
		_w3739_
	);
	LUT3 #(
		.INIT('hf2)
	) name3287 (
		\EAX_reg[5]/NET0131 ,
		_w2643_,
		_w3739_,
		_w3740_
	);
	LUT3 #(
		.INIT('h20)
	) name3288 (
		\Datai[6]_pad ,
		READY_n_pad,
		_w588_,
		_w3741_
	);
	LUT4 #(
		.INIT('h0080)
	) name3289 (
		_w602_,
		_w604_,
		_w634_,
		_w853_,
		_w3742_
	);
	LUT4 #(
		.INIT('h78f0)
	) name3290 (
		\EAX_reg[4]/NET0131 ,
		\EAX_reg[5]/NET0131 ,
		\EAX_reg[6]/NET0131 ,
		_w1743_,
		_w3743_
	);
	LUT3 #(
		.INIT('h80)
	) name3291 (
		_w518_,
		_w617_,
		_w3743_,
		_w3744_
	);
	LUT2 #(
		.INIT('h1)
	) name3292 (
		_w3742_,
		_w3744_,
		_w3745_
	);
	LUT3 #(
		.INIT('h8a)
	) name3293 (
		_w690_,
		_w3741_,
		_w3745_,
		_w3746_
	);
	LUT3 #(
		.INIT('hf2)
	) name3294 (
		\EAX_reg[6]/NET0131 ,
		_w2643_,
		_w3746_,
		_w3747_
	);
	LUT2 #(
		.INIT('h2)
	) name3295 (
		\EAX_reg[1]/NET0131 ,
		_w1841_,
		_w3748_
	);
	LUT3 #(
		.INIT('h40)
	) name3296 (
		\EAX_reg[0]/NET0131 ,
		_w518_,
		_w617_,
		_w3749_
	);
	LUT4 #(
		.INIT('haaa8)
	) name3297 (
		\EAX_reg[1]/NET0131 ,
		_w653_,
		_w1742_,
		_w3749_,
		_w3750_
	);
	LUT4 #(
		.INIT('h0080)
	) name3298 (
		_w602_,
		_w604_,
		_w634_,
		_w806_,
		_w3751_
	);
	LUT4 #(
		.INIT('h2202)
	) name3299 (
		\Datai[1]_pad ,
		READY_n_pad,
		_w563_,
		_w565_,
		_w3752_
	);
	LUT4 #(
		.INIT('hf800)
	) name3300 (
		_w494_,
		_w586_,
		_w582_,
		_w3752_,
		_w3753_
	);
	LUT2 #(
		.INIT('h2)
	) name3301 (
		\EAX_reg[0]/NET0131 ,
		\EAX_reg[1]/NET0131 ,
		_w3754_
	);
	LUT3 #(
		.INIT('h80)
	) name3302 (
		_w518_,
		_w617_,
		_w3754_,
		_w3755_
	);
	LUT3 #(
		.INIT('h01)
	) name3303 (
		_w3753_,
		_w3751_,
		_w3755_,
		_w3756_
	);
	LUT4 #(
		.INIT('hecee)
	) name3304 (
		_w690_,
		_w3748_,
		_w3750_,
		_w3756_,
		_w3757_
	);
	LUT3 #(
		.INIT('ha2)
	) name3305 (
		\MemoryFetch_reg/NET0131 ,
		_w586_,
		_w566_,
		_w3758_
	);
	LUT3 #(
		.INIT('hc4)
	) name3306 (
		\MemoryFetch_reg/NET0131 ,
		_w2084_,
		_w2085_,
		_w3759_
	);
	LUT4 #(
		.INIT('ha2ff)
	) name3307 (
		_w690_,
		_w2102_,
		_w3758_,
		_w3759_,
		_w3760_
	);
	LUT4 #(
		.INIT('hf200)
	) name3308 (
		\ReadRequest_reg/NET0131 ,
		_w646_,
		_w588_,
		_w690_,
		_w3761_
	);
	LUT3 #(
		.INIT('hc4)
	) name3309 (
		\ReadRequest_reg/NET0131 ,
		_w2084_,
		_w2085_,
		_w3762_
	);
	LUT2 #(
		.INIT('hb)
	) name3310 (
		_w3761_,
		_w3762_,
		_w3763_
	);
	LUT2 #(
		.INIT('h2)
	) name3311 (
		\rEIP_reg[0]/NET0131 ,
		_w3110_,
		_w3764_
	);
	LUT4 #(
		.INIT('hcdc8)
	) name3312 (
		\DataWidth_reg[1]/NET0131 ,
		\EBX_reg[0]/NET0131 ,
		READY_n_pad,
		\rEIP_reg[0]/NET0131 ,
		_w3765_
	);
	LUT4 #(
		.INIT('hae00)
	) name3313 (
		_w582_,
		_w589_,
		_w594_,
		_w3765_,
		_w3766_
	);
	LUT4 #(
		.INIT('ha88a)
	) name3314 (
		\EBX_reg[0]/NET0131 ,
		\State_reg[0]/NET0131 ,
		\State_reg[1]/NET0131 ,
		\State_reg[2]/NET0131 ,
		_w3767_
	);
	LUT4 #(
		.INIT('h0bbb)
	) name3315 (
		\InstQueueRd_Addr_reg[0]/NET0131 ,
		_w586_,
		_w589_,
		_w3767_,
		_w3768_
	);
	LUT3 #(
		.INIT('h45)
	) name3316 (
		_w566_,
		_w3766_,
		_w3768_,
		_w3769_
	);
	LUT4 #(
		.INIT('hcc40)
	) name3317 (
		\DataWidth_reg[1]/NET0131 ,
		\PhyAddrPointer_reg[0]/NET0131 ,
		_w695_,
		_w706_,
		_w3770_
	);
	LUT4 #(
		.INIT('h80cc)
	) name3318 (
		\DataWidth_reg[1]/NET0131 ,
		\rEIP_reg[0]/NET0131 ,
		_w695_,
		_w3101_,
		_w3771_
	);
	LUT2 #(
		.INIT('h1)
	) name3319 (
		_w3770_,
		_w3771_,
		_w3772_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name3320 (
		_w690_,
		_w3764_,
		_w3769_,
		_w3772_,
		_w3773_
	);
	LUT4 #(
		.INIT('h8000)
	) name3321 (
		\EAX_reg[25]/NET0131 ,
		_w1917_,
		_w1918_,
		_w2093_,
		_w3774_
	);
	LUT3 #(
		.INIT('h21)
	) name3322 (
		\EAX_reg[30]/NET0131 ,
		_w594_,
		_w3774_,
		_w3775_
	);
	LUT4 #(
		.INIT('h0a02)
	) name3323 (
		_w646_,
		_w687_,
		_w2183_,
		_w3775_,
		_w3776_
	);
	LUT4 #(
		.INIT('h4080)
	) name3324 (
		\EAX_reg[30]/NET0131 ,
		_w589_,
		_w595_,
		_w3774_,
		_w3777_
	);
	LUT4 #(
		.INIT('hcc08)
	) name3325 (
		\Datao[30]_pad ,
		_w690_,
		_w3776_,
		_w3777_,
		_w3778_
	);
	LUT4 #(
		.INIT('h3f15)
	) name3326 (
		\Datao[30]_pad ,
		\uWord_reg[14]/NET0131 ,
		_w2179_,
		_w2180_,
		_w3779_
	);
	LUT2 #(
		.INIT('hb)
	) name3327 (
		_w3778_,
		_w3779_,
		_w3780_
	);
	LUT2 #(
		.INIT('h2)
	) name3328 (
		\EAX_reg[28]/NET0131 ,
		_w1841_,
		_w3781_
	);
	LUT4 #(
		.INIT('h4888)
	) name3329 (
		\EAX_reg[28]/NET0131 ,
		_w1741_,
		_w1760_,
		_w1917_,
		_w3782_
	);
	LUT3 #(
		.INIT('h2d)
	) name3330 (
		_w1821_,
		_w1832_,
		_w1934_,
		_w3783_
	);
	LUT4 #(
		.INIT('h88a8)
	) name3331 (
		\EAX_reg[28]/NET0131 ,
		READY_n_pad,
		_w563_,
		_w565_,
		_w3784_
	);
	LUT4 #(
		.INIT('h2202)
	) name3332 (
		\Datai[28]_pad ,
		READY_n_pad,
		_w563_,
		_w565_,
		_w3785_
	);
	LUT2 #(
		.INIT('h1)
	) name3333 (
		_w3784_,
		_w3785_,
		_w3786_
	);
	LUT3 #(
		.INIT('h08)
	) name3334 (
		_w494_,
		_w586_,
		_w3786_,
		_w3787_
	);
	LUT2 #(
		.INIT('h1)
	) name3335 (
		_w2099_,
		_w3784_,
		_w3788_
	);
	LUT2 #(
		.INIT('h2)
	) name3336 (
		_w582_,
		_w3788_,
		_w3789_
	);
	LUT4 #(
		.INIT('h0013)
	) name3337 (
		_w1740_,
		_w3787_,
		_w3783_,
		_w3789_,
		_w3790_
	);
	LUT3 #(
		.INIT('h70)
	) name3338 (
		\EAX_reg[28]/NET0131 ,
		_w1742_,
		_w3790_,
		_w3791_
	);
	LUT4 #(
		.INIT('hecee)
	) name3339 (
		_w690_,
		_w3781_,
		_w3782_,
		_w3791_,
		_w3792_
	);
	LUT2 #(
		.INIT('h2)
	) name3340 (
		\uWord_reg[14]/NET0131 ,
		_w1841_,
		_w3793_
	);
	LUT4 #(
		.INIT('h0408)
	) name3341 (
		\EAX_reg[30]/NET0131 ,
		_w589_,
		_w566_,
		_w3774_,
		_w3794_
	);
	LUT3 #(
		.INIT('h80)
	) name3342 (
		\Datai[14]_pad ,
		_w582_,
		_w652_,
		_w3795_
	);
	LUT4 #(
		.INIT('h000d)
	) name3343 (
		\uWord_reg[14]/NET0131 ,
		_w2103_,
		_w3795_,
		_w3794_,
		_w3796_
	);
	LUT3 #(
		.INIT('hce)
	) name3344 (
		_w690_,
		_w3793_,
		_w3796_,
		_w3797_
	);
	LUT3 #(
		.INIT('h20)
	) name3345 (
		\Datai[0]_pad ,
		READY_n_pad,
		_w588_,
		_w3798_
	);
	LUT4 #(
		.INIT('h0080)
	) name3346 (
		_w602_,
		_w604_,
		_w634_,
		_w818_,
		_w3799_
	);
	LUT2 #(
		.INIT('h1)
	) name3347 (
		_w3749_,
		_w3799_,
		_w3800_
	);
	LUT3 #(
		.INIT('h8a)
	) name3348 (
		_w690_,
		_w3798_,
		_w3800_,
		_w3801_
	);
	LUT3 #(
		.INIT('hf2)
	) name3349 (
		\EAX_reg[0]/NET0131 ,
		_w2643_,
		_w3801_,
		_w3802_
	);
	LUT4 #(
		.INIT('h4888)
	) name3350 (
		\EBX_reg[28]/NET0131 ,
		_w622_,
		_w1986_,
		_w1987_,
		_w3803_
	);
	LUT4 #(
		.INIT('h31fd)
	) name3351 (
		\EBX_reg[28]/NET0131 ,
		_w1990_,
		_w1991_,
		_w3783_,
		_w3804_
	);
	LUT2 #(
		.INIT('h2)
	) name3352 (
		\EBX_reg[28]/NET0131 ,
		_w1841_,
		_w3805_
	);
	LUT4 #(
		.INIT('hff8a)
	) name3353 (
		_w690_,
		_w3803_,
		_w3804_,
		_w3805_,
		_w3806_
	);
	LUT4 #(
		.INIT('h4080)
	) name3354 (
		\EAX_reg[16]/NET0131 ,
		_w518_,
		_w617_,
		_w1751_,
		_w3807_
	);
	LUT4 #(
		.INIT('h88a8)
	) name3355 (
		\EAX_reg[16]/NET0131 ,
		READY_n_pad,
		_w563_,
		_w565_,
		_w3808_
	);
	LUT4 #(
		.INIT('h2202)
	) name3356 (
		\Datai[16]_pad ,
		READY_n_pad,
		_w563_,
		_w565_,
		_w3809_
	);
	LUT2 #(
		.INIT('h1)
	) name3357 (
		_w3808_,
		_w3809_,
		_w3810_
	);
	LUT3 #(
		.INIT('h08)
	) name3358 (
		_w494_,
		_w586_,
		_w3810_,
		_w3811_
	);
	LUT4 #(
		.INIT('h135f)
	) name3359 (
		\InstQueue_reg[0][0]/NET0131 ,
		\InstQueue_reg[4][0]/NET0131 ,
		_w461_,
		_w473_,
		_w3812_
	);
	LUT4 #(
		.INIT('h153f)
	) name3360 (
		\InstQueue_reg[14][0]/NET0131 ,
		\InstQueue_reg[8][0]/NET0131 ,
		_w457_,
		_w458_,
		_w3813_
	);
	LUT4 #(
		.INIT('h135f)
	) name3361 (
		\InstQueue_reg[1][0]/NET0131 ,
		\InstQueue_reg[9][0]/NET0131 ,
		_w476_,
		_w453_,
		_w3814_
	);
	LUT4 #(
		.INIT('h153f)
	) name3362 (
		\InstQueue_reg[2][0]/NET0131 ,
		\InstQueue_reg[6][0]/NET0131 ,
		_w460_,
		_w455_,
		_w3815_
	);
	LUT4 #(
		.INIT('h8000)
	) name3363 (
		_w3814_,
		_w3815_,
		_w3812_,
		_w3813_,
		_w3816_
	);
	LUT4 #(
		.INIT('h153f)
	) name3364 (
		\InstQueue_reg[15][0]/NET0131 ,
		\InstQueue_reg[5][0]/NET0131 ,
		_w474_,
		_w477_,
		_w3817_
	);
	LUT4 #(
		.INIT('h153f)
	) name3365 (
		\InstQueue_reg[12][0]/NET0131 ,
		\InstQueue_reg[13][0]/NET0131 ,
		_w471_,
		_w467_,
		_w3818_
	);
	LUT4 #(
		.INIT('h153f)
	) name3366 (
		\InstQueue_reg[3][0]/NET0131 ,
		\InstQueue_reg[7][0]/NET0131 ,
		_w468_,
		_w464_,
		_w3819_
	);
	LUT4 #(
		.INIT('h135f)
	) name3367 (
		\InstQueue_reg[10][0]/NET0131 ,
		\InstQueue_reg[11][0]/NET0131 ,
		_w470_,
		_w463_,
		_w3820_
	);
	LUT4 #(
		.INIT('h8000)
	) name3368 (
		_w3819_,
		_w3820_,
		_w3817_,
		_w3818_,
		_w3821_
	);
	LUT2 #(
		.INIT('h8)
	) name3369 (
		_w3816_,
		_w3821_,
		_w3822_
	);
	LUT4 #(
		.INIT('h0080)
	) name3370 (
		_w602_,
		_w604_,
		_w634_,
		_w3822_,
		_w3823_
	);
	LUT4 #(
		.INIT('h2202)
	) name3371 (
		\Datai[0]_pad ,
		READY_n_pad,
		_w563_,
		_w565_,
		_w3824_
	);
	LUT2 #(
		.INIT('h1)
	) name3372 (
		_w3824_,
		_w3808_,
		_w3825_
	);
	LUT2 #(
		.INIT('h2)
	) name3373 (
		_w582_,
		_w3825_,
		_w3826_
	);
	LUT3 #(
		.INIT('h01)
	) name3374 (
		_w3823_,
		_w3826_,
		_w3811_,
		_w3827_
	);
	LUT4 #(
		.INIT('h0700)
	) name3375 (
		\EAX_reg[16]/NET0131 ,
		_w1742_,
		_w3807_,
		_w3827_,
		_w3828_
	);
	LUT2 #(
		.INIT('h2)
	) name3376 (
		\EAX_reg[16]/NET0131 ,
		_w1841_,
		_w3829_
	);
	LUT3 #(
		.INIT('hf2)
	) name3377 (
		_w690_,
		_w3828_,
		_w3829_,
		_w3830_
	);
	LUT2 #(
		.INIT('h2)
	) name3378 (
		\EAX_reg[17]/NET0131 ,
		_w1841_,
		_w3831_
	);
	LUT3 #(
		.INIT('h48)
	) name3379 (
		\EAX_reg[17]/NET0131 ,
		_w1741_,
		_w1752_,
		_w3832_
	);
	LUT4 #(
		.INIT('h88a8)
	) name3380 (
		\EAX_reg[17]/NET0131 ,
		READY_n_pad,
		_w563_,
		_w565_,
		_w3833_
	);
	LUT4 #(
		.INIT('h2202)
	) name3381 (
		\Datai[17]_pad ,
		READY_n_pad,
		_w563_,
		_w565_,
		_w3834_
	);
	LUT2 #(
		.INIT('h1)
	) name3382 (
		_w3833_,
		_w3834_,
		_w3835_
	);
	LUT3 #(
		.INIT('h08)
	) name3383 (
		_w494_,
		_w586_,
		_w3835_,
		_w3836_
	);
	LUT4 #(
		.INIT('h153f)
	) name3384 (
		\InstQueue_reg[3][1]/NET0131 ,
		\InstQueue_reg[5][1]/NET0131 ,
		_w474_,
		_w464_,
		_w3837_
	);
	LUT4 #(
		.INIT('h135f)
	) name3385 (
		\InstQueue_reg[15][1]/NET0131 ,
		\InstQueue_reg[7][1]/NET0131 ,
		_w477_,
		_w468_,
		_w3838_
	);
	LUT4 #(
		.INIT('h135f)
	) name3386 (
		\InstQueue_reg[1][1]/NET0131 ,
		\InstQueue_reg[9][1]/NET0131 ,
		_w476_,
		_w453_,
		_w3839_
	);
	LUT4 #(
		.INIT('h135f)
	) name3387 (
		\InstQueue_reg[13][1]/NET0131 ,
		\InstQueue_reg[6][1]/NET0131 ,
		_w471_,
		_w460_,
		_w3840_
	);
	LUT4 #(
		.INIT('h8000)
	) name3388 (
		_w3839_,
		_w3840_,
		_w3837_,
		_w3838_,
		_w3841_
	);
	LUT4 #(
		.INIT('h153f)
	) name3389 (
		\InstQueue_reg[2][1]/NET0131 ,
		\InstQueue_reg[4][1]/NET0131 ,
		_w473_,
		_w455_,
		_w3842_
	);
	LUT4 #(
		.INIT('h135f)
	) name3390 (
		\InstQueue_reg[12][1]/NET0131 ,
		\InstQueue_reg[8][1]/NET0131 ,
		_w467_,
		_w457_,
		_w3843_
	);
	LUT4 #(
		.INIT('h153f)
	) name3391 (
		\InstQueue_reg[0][1]/NET0131 ,
		\InstQueue_reg[10][1]/NET0131 ,
		_w470_,
		_w461_,
		_w3844_
	);
	LUT4 #(
		.INIT('h135f)
	) name3392 (
		\InstQueue_reg[11][1]/NET0131 ,
		\InstQueue_reg[14][1]/NET0131 ,
		_w463_,
		_w458_,
		_w3845_
	);
	LUT4 #(
		.INIT('h8000)
	) name3393 (
		_w3844_,
		_w3845_,
		_w3842_,
		_w3843_,
		_w3846_
	);
	LUT2 #(
		.INIT('h8)
	) name3394 (
		_w3841_,
		_w3846_,
		_w3847_
	);
	LUT4 #(
		.INIT('h0080)
	) name3395 (
		_w602_,
		_w604_,
		_w634_,
		_w3847_,
		_w3848_
	);
	LUT2 #(
		.INIT('h1)
	) name3396 (
		_w3752_,
		_w3833_,
		_w3849_
	);
	LUT2 #(
		.INIT('h2)
	) name3397 (
		_w582_,
		_w3849_,
		_w3850_
	);
	LUT3 #(
		.INIT('h01)
	) name3398 (
		_w3848_,
		_w3850_,
		_w3836_,
		_w3851_
	);
	LUT4 #(
		.INIT('h0700)
	) name3399 (
		\EAX_reg[17]/NET0131 ,
		_w1742_,
		_w3832_,
		_w3851_,
		_w3852_
	);
	LUT3 #(
		.INIT('hce)
	) name3400 (
		_w690_,
		_w3831_,
		_w3852_,
		_w3853_
	);
	LUT2 #(
		.INIT('h2)
	) name3401 (
		\EAX_reg[18]/NET0131 ,
		_w1841_,
		_w3854_
	);
	LUT3 #(
		.INIT('h48)
	) name3402 (
		\EAX_reg[18]/NET0131 ,
		_w1741_,
		_w1753_,
		_w3855_
	);
	LUT4 #(
		.INIT('h88a8)
	) name3403 (
		\EAX_reg[18]/NET0131 ,
		READY_n_pad,
		_w563_,
		_w565_,
		_w3856_
	);
	LUT2 #(
		.INIT('h1)
	) name3404 (
		_w3700_,
		_w3856_,
		_w3857_
	);
	LUT2 #(
		.INIT('h2)
	) name3405 (
		_w582_,
		_w3857_,
		_w3858_
	);
	LUT4 #(
		.INIT('h153f)
	) name3406 (
		\InstQueue_reg[0][2]/NET0131 ,
		\InstQueue_reg[5][2]/NET0131 ,
		_w474_,
		_w461_,
		_w3859_
	);
	LUT4 #(
		.INIT('h153f)
	) name3407 (
		\InstQueue_reg[12][2]/NET0131 ,
		\InstQueue_reg[7][2]/NET0131 ,
		_w468_,
		_w467_,
		_w3860_
	);
	LUT4 #(
		.INIT('h135f)
	) name3408 (
		\InstQueue_reg[11][2]/NET0131 ,
		\InstQueue_reg[2][2]/NET0131 ,
		_w463_,
		_w455_,
		_w3861_
	);
	LUT4 #(
		.INIT('h135f)
	) name3409 (
		\InstQueue_reg[1][2]/NET0131 ,
		\InstQueue_reg[8][2]/NET0131 ,
		_w476_,
		_w457_,
		_w3862_
	);
	LUT4 #(
		.INIT('h8000)
	) name3410 (
		_w3861_,
		_w3862_,
		_w3859_,
		_w3860_,
		_w3863_
	);
	LUT4 #(
		.INIT('h135f)
	) name3411 (
		\InstQueue_reg[10][2]/NET0131 ,
		\InstQueue_reg[9][2]/NET0131 ,
		_w470_,
		_w453_,
		_w3864_
	);
	LUT4 #(
		.INIT('h153f)
	) name3412 (
		\InstQueue_reg[14][2]/NET0131 ,
		\InstQueue_reg[15][2]/NET0131 ,
		_w477_,
		_w458_,
		_w3865_
	);
	LUT4 #(
		.INIT('h135f)
	) name3413 (
		\InstQueue_reg[13][2]/NET0131 ,
		\InstQueue_reg[6][2]/NET0131 ,
		_w471_,
		_w460_,
		_w3866_
	);
	LUT4 #(
		.INIT('h135f)
	) name3414 (
		\InstQueue_reg[3][2]/NET0131 ,
		\InstQueue_reg[4][2]/NET0131 ,
		_w464_,
		_w473_,
		_w3867_
	);
	LUT4 #(
		.INIT('h8000)
	) name3415 (
		_w3866_,
		_w3867_,
		_w3864_,
		_w3865_,
		_w3868_
	);
	LUT2 #(
		.INIT('h8)
	) name3416 (
		_w3863_,
		_w3868_,
		_w3869_
	);
	LUT4 #(
		.INIT('h0080)
	) name3417 (
		_w602_,
		_w604_,
		_w634_,
		_w3869_,
		_w3870_
	);
	LUT4 #(
		.INIT('h2202)
	) name3418 (
		\Datai[18]_pad ,
		READY_n_pad,
		_w563_,
		_w565_,
		_w3871_
	);
	LUT2 #(
		.INIT('h1)
	) name3419 (
		_w3856_,
		_w3871_,
		_w3872_
	);
	LUT3 #(
		.INIT('h08)
	) name3420 (
		_w494_,
		_w586_,
		_w3872_,
		_w3873_
	);
	LUT3 #(
		.INIT('h01)
	) name3421 (
		_w3870_,
		_w3873_,
		_w3858_,
		_w3874_
	);
	LUT4 #(
		.INIT('h0700)
	) name3422 (
		\EAX_reg[18]/NET0131 ,
		_w1742_,
		_w3855_,
		_w3874_,
		_w3875_
	);
	LUT3 #(
		.INIT('hce)
	) name3423 (
		_w690_,
		_w3854_,
		_w3875_,
		_w3876_
	);
	LUT3 #(
		.INIT('h48)
	) name3424 (
		\EAX_reg[19]/NET0131 ,
		_w1741_,
		_w1754_,
		_w3877_
	);
	LUT4 #(
		.INIT('h88a8)
	) name3425 (
		\EAX_reg[19]/NET0131 ,
		READY_n_pad,
		_w563_,
		_w565_,
		_w3878_
	);
	LUT2 #(
		.INIT('h1)
	) name3426 (
		_w3708_,
		_w3878_,
		_w3879_
	);
	LUT2 #(
		.INIT('h2)
	) name3427 (
		_w582_,
		_w3879_,
		_w3880_
	);
	LUT4 #(
		.INIT('h135f)
	) name3428 (
		\InstQueue_reg[3][3]/NET0131 ,
		\InstQueue_reg[4][3]/NET0131 ,
		_w464_,
		_w473_,
		_w3881_
	);
	LUT4 #(
		.INIT('h135f)
	) name3429 (
		\InstQueue_reg[13][3]/NET0131 ,
		\InstQueue_reg[14][3]/NET0131 ,
		_w471_,
		_w458_,
		_w3882_
	);
	LUT4 #(
		.INIT('h153f)
	) name3430 (
		\InstQueue_reg[12][3]/NET0131 ,
		\InstQueue_reg[1][3]/NET0131 ,
		_w476_,
		_w467_,
		_w3883_
	);
	LUT4 #(
		.INIT('h135f)
	) name3431 (
		\InstQueue_reg[6][3]/NET0131 ,
		\InstQueue_reg[8][3]/NET0131 ,
		_w460_,
		_w457_,
		_w3884_
	);
	LUT4 #(
		.INIT('h8000)
	) name3432 (
		_w3883_,
		_w3884_,
		_w3881_,
		_w3882_,
		_w3885_
	);
	LUT4 #(
		.INIT('h153f)
	) name3433 (
		\InstQueue_reg[2][3]/NET0131 ,
		\InstQueue_reg[5][3]/NET0131 ,
		_w474_,
		_w455_,
		_w3886_
	);
	LUT4 #(
		.INIT('h135f)
	) name3434 (
		\InstQueue_reg[0][3]/NET0131 ,
		\InstQueue_reg[9][3]/NET0131 ,
		_w461_,
		_w453_,
		_w3887_
	);
	LUT4 #(
		.INIT('h135f)
	) name3435 (
		\InstQueue_reg[15][3]/NET0131 ,
		\InstQueue_reg[7][3]/NET0131 ,
		_w477_,
		_w468_,
		_w3888_
	);
	LUT4 #(
		.INIT('h135f)
	) name3436 (
		\InstQueue_reg[10][3]/NET0131 ,
		\InstQueue_reg[11][3]/NET0131 ,
		_w470_,
		_w463_,
		_w3889_
	);
	LUT4 #(
		.INIT('h8000)
	) name3437 (
		_w3888_,
		_w3889_,
		_w3886_,
		_w3887_,
		_w3890_
	);
	LUT2 #(
		.INIT('h8)
	) name3438 (
		_w3885_,
		_w3890_,
		_w3891_
	);
	LUT4 #(
		.INIT('h0080)
	) name3439 (
		_w602_,
		_w604_,
		_w634_,
		_w3891_,
		_w3892_
	);
	LUT4 #(
		.INIT('h2202)
	) name3440 (
		\Datai[19]_pad ,
		READY_n_pad,
		_w563_,
		_w565_,
		_w3893_
	);
	LUT2 #(
		.INIT('h1)
	) name3441 (
		_w3878_,
		_w3893_,
		_w3894_
	);
	LUT3 #(
		.INIT('h08)
	) name3442 (
		_w494_,
		_w586_,
		_w3894_,
		_w3895_
	);
	LUT3 #(
		.INIT('h01)
	) name3443 (
		_w3892_,
		_w3895_,
		_w3880_,
		_w3896_
	);
	LUT4 #(
		.INIT('h0700)
	) name3444 (
		\EAX_reg[19]/NET0131 ,
		_w1742_,
		_w3877_,
		_w3896_,
		_w3897_
	);
	LUT2 #(
		.INIT('h2)
	) name3445 (
		\EAX_reg[19]/NET0131 ,
		_w1841_,
		_w3898_
	);
	LUT3 #(
		.INIT('hf2)
	) name3446 (
		_w690_,
		_w3897_,
		_w3898_,
		_w3899_
	);
	LUT2 #(
		.INIT('h2)
	) name3447 (
		\More_reg/NET0131 ,
		_w1841_,
		_w3900_
	);
	LUT4 #(
		.INIT('hffb0)
	) name3448 (
		_w678_,
		_w682_,
		_w690_,
		_w3900_,
		_w3901_
	);
	LUT4 #(
		.INIT('h70f0)
	) name3449 (
		\EAX_reg[19]/NET0131 ,
		\EAX_reg[20]/NET0131 ,
		_w1741_,
		_w1754_,
		_w3902_
	);
	LUT4 #(
		.INIT('h60c0)
	) name3450 (
		\EAX_reg[19]/NET0131 ,
		\EAX_reg[20]/NET0131 ,
		_w1741_,
		_w1754_,
		_w3903_
	);
	LUT4 #(
		.INIT('h88a8)
	) name3451 (
		\EAX_reg[20]/NET0131 ,
		READY_n_pad,
		_w563_,
		_w565_,
		_w3904_
	);
	LUT2 #(
		.INIT('h1)
	) name3452 (
		_w2442_,
		_w3904_,
		_w3905_
	);
	LUT2 #(
		.INIT('h2)
	) name3453 (
		_w582_,
		_w3905_,
		_w3906_
	);
	LUT4 #(
		.INIT('h135f)
	) name3454 (
		\InstQueue_reg[5][4]/NET0131 ,
		\InstQueue_reg[7][4]/NET0131 ,
		_w474_,
		_w468_,
		_w3907_
	);
	LUT4 #(
		.INIT('h153f)
	) name3455 (
		\InstQueue_reg[2][4]/NET0131 ,
		\InstQueue_reg[9][4]/NET0131 ,
		_w453_,
		_w455_,
		_w3908_
	);
	LUT4 #(
		.INIT('h135f)
	) name3456 (
		\InstQueue_reg[10][4]/NET0131 ,
		\InstQueue_reg[8][4]/NET0131 ,
		_w470_,
		_w457_,
		_w3909_
	);
	LUT4 #(
		.INIT('h153f)
	) name3457 (
		\InstQueue_reg[12][4]/NET0131 ,
		\InstQueue_reg[6][4]/NET0131 ,
		_w460_,
		_w467_,
		_w3910_
	);
	LUT4 #(
		.INIT('h8000)
	) name3458 (
		_w3909_,
		_w3910_,
		_w3907_,
		_w3908_,
		_w3911_
	);
	LUT4 #(
		.INIT('h135f)
	) name3459 (
		\InstQueue_reg[15][4]/NET0131 ,
		\InstQueue_reg[1][4]/NET0131 ,
		_w477_,
		_w476_,
		_w3912_
	);
	LUT4 #(
		.INIT('h135f)
	) name3460 (
		\InstQueue_reg[0][4]/NET0131 ,
		\InstQueue_reg[11][4]/NET0131 ,
		_w461_,
		_w463_,
		_w3913_
	);
	LUT4 #(
		.INIT('h153f)
	) name3461 (
		\InstQueue_reg[14][4]/NET0131 ,
		\InstQueue_reg[3][4]/NET0131 ,
		_w464_,
		_w458_,
		_w3914_
	);
	LUT4 #(
		.INIT('h135f)
	) name3462 (
		\InstQueue_reg[13][4]/NET0131 ,
		\InstQueue_reg[4][4]/NET0131 ,
		_w471_,
		_w473_,
		_w3915_
	);
	LUT4 #(
		.INIT('h8000)
	) name3463 (
		_w3914_,
		_w3915_,
		_w3912_,
		_w3913_,
		_w3916_
	);
	LUT2 #(
		.INIT('h8)
	) name3464 (
		_w3911_,
		_w3916_,
		_w3917_
	);
	LUT4 #(
		.INIT('h0080)
	) name3465 (
		_w602_,
		_w604_,
		_w634_,
		_w3917_,
		_w3918_
	);
	LUT4 #(
		.INIT('h2202)
	) name3466 (
		\Datai[20]_pad ,
		READY_n_pad,
		_w563_,
		_w565_,
		_w3919_
	);
	LUT2 #(
		.INIT('h1)
	) name3467 (
		_w3904_,
		_w3919_,
		_w3920_
	);
	LUT3 #(
		.INIT('h08)
	) name3468 (
		_w494_,
		_w586_,
		_w3920_,
		_w3921_
	);
	LUT3 #(
		.INIT('h01)
	) name3469 (
		_w3918_,
		_w3921_,
		_w3906_,
		_w3922_
	);
	LUT4 #(
		.INIT('h0700)
	) name3470 (
		\EAX_reg[20]/NET0131 ,
		_w1742_,
		_w3903_,
		_w3922_,
		_w3923_
	);
	LUT2 #(
		.INIT('h2)
	) name3471 (
		\EAX_reg[20]/NET0131 ,
		_w1841_,
		_w3924_
	);
	LUT3 #(
		.INIT('hf2)
	) name3472 (
		_w690_,
		_w3923_,
		_w3924_,
		_w3925_
	);
	LUT2 #(
		.INIT('h2)
	) name3473 (
		\EAX_reg[21]/NET0131 ,
		_w1841_,
		_w3926_
	);
	LUT3 #(
		.INIT('ha8)
	) name3474 (
		\EAX_reg[21]/NET0131 ,
		_w1742_,
		_w3902_,
		_w3927_
	);
	LUT3 #(
		.INIT('h40)
	) name3475 (
		\EAX_reg[21]/NET0131 ,
		_w518_,
		_w617_,
		_w3928_
	);
	LUT4 #(
		.INIT('h8000)
	) name3476 (
		\EAX_reg[19]/NET0131 ,
		\EAX_reg[20]/NET0131 ,
		_w1754_,
		_w3928_,
		_w3929_
	);
	LUT4 #(
		.INIT('h88a8)
	) name3477 (
		\EAX_reg[21]/NET0131 ,
		READY_n_pad,
		_w563_,
		_w565_,
		_w3930_
	);
	LUT4 #(
		.INIT('h2202)
	) name3478 (
		\Datai[21]_pad ,
		READY_n_pad,
		_w563_,
		_w565_,
		_w3931_
	);
	LUT2 #(
		.INIT('h1)
	) name3479 (
		_w3930_,
		_w3931_,
		_w3932_
	);
	LUT3 #(
		.INIT('h08)
	) name3480 (
		_w494_,
		_w586_,
		_w3932_,
		_w3933_
	);
	LUT4 #(
		.INIT('h135f)
	) name3481 (
		\InstQueue_reg[15][5]/NET0131 ,
		\InstQueue_reg[4][5]/NET0131 ,
		_w477_,
		_w473_,
		_w3934_
	);
	LUT4 #(
		.INIT('h135f)
	) name3482 (
		\InstQueue_reg[0][5]/NET0131 ,
		\InstQueue_reg[11][5]/NET0131 ,
		_w461_,
		_w463_,
		_w3935_
	);
	LUT4 #(
		.INIT('h135f)
	) name3483 (
		\InstQueue_reg[1][5]/NET0131 ,
		\InstQueue_reg[9][5]/NET0131 ,
		_w476_,
		_w453_,
		_w3936_
	);
	LUT4 #(
		.INIT('h153f)
	) name3484 (
		\InstQueue_reg[6][5]/NET0131 ,
		\InstQueue_reg[7][5]/NET0131 ,
		_w468_,
		_w460_,
		_w3937_
	);
	LUT4 #(
		.INIT('h8000)
	) name3485 (
		_w3936_,
		_w3937_,
		_w3934_,
		_w3935_,
		_w3938_
	);
	LUT4 #(
		.INIT('h153f)
	) name3486 (
		\InstQueue_reg[3][5]/NET0131 ,
		\InstQueue_reg[5][5]/NET0131 ,
		_w474_,
		_w464_,
		_w3939_
	);
	LUT4 #(
		.INIT('h135f)
	) name3487 (
		\InstQueue_reg[12][5]/NET0131 ,
		\InstQueue_reg[2][5]/NET0131 ,
		_w467_,
		_w455_,
		_w3940_
	);
	LUT4 #(
		.INIT('h135f)
	) name3488 (
		\InstQueue_reg[13][5]/NET0131 ,
		\InstQueue_reg[8][5]/NET0131 ,
		_w471_,
		_w457_,
		_w3941_
	);
	LUT4 #(
		.INIT('h135f)
	) name3489 (
		\InstQueue_reg[10][5]/NET0131 ,
		\InstQueue_reg[14][5]/NET0131 ,
		_w470_,
		_w458_,
		_w3942_
	);
	LUT4 #(
		.INIT('h8000)
	) name3490 (
		_w3941_,
		_w3942_,
		_w3939_,
		_w3940_,
		_w3943_
	);
	LUT2 #(
		.INIT('h8)
	) name3491 (
		_w3938_,
		_w3943_,
		_w3944_
	);
	LUT4 #(
		.INIT('h0080)
	) name3492 (
		_w602_,
		_w604_,
		_w634_,
		_w3944_,
		_w3945_
	);
	LUT2 #(
		.INIT('h1)
	) name3493 (
		_w3734_,
		_w3930_,
		_w3946_
	);
	LUT2 #(
		.INIT('h2)
	) name3494 (
		_w582_,
		_w3946_,
		_w3947_
	);
	LUT3 #(
		.INIT('h01)
	) name3495 (
		_w3945_,
		_w3947_,
		_w3933_,
		_w3948_
	);
	LUT2 #(
		.INIT('h4)
	) name3496 (
		_w3929_,
		_w3948_,
		_w3949_
	);
	LUT4 #(
		.INIT('hecee)
	) name3497 (
		_w690_,
		_w3926_,
		_w3927_,
		_w3949_,
		_w3950_
	);
	LUT2 #(
		.INIT('h2)
	) name3498 (
		\EAX_reg[22]/NET0131 ,
		_w1841_,
		_w3951_
	);
	LUT4 #(
		.INIT('h1333)
	) name3499 (
		\EAX_reg[19]/NET0131 ,
		\EAX_reg[22]/NET0131 ,
		_w1754_,
		_w1755_,
		_w3952_
	);
	LUT3 #(
		.INIT('h2a)
	) name3500 (
		_w1741_,
		_w1754_,
		_w1757_,
		_w3953_
	);
	LUT2 #(
		.INIT('h4)
	) name3501 (
		_w3952_,
		_w3953_,
		_w3954_
	);
	LUT4 #(
		.INIT('h153f)
	) name3502 (
		\InstQueue_reg[3][6]/NET0131 ,
		\InstQueue_reg[5][6]/NET0131 ,
		_w474_,
		_w464_,
		_w3955_
	);
	LUT4 #(
		.INIT('h135f)
	) name3503 (
		\InstQueue_reg[12][6]/NET0131 ,
		\InstQueue_reg[2][6]/NET0131 ,
		_w467_,
		_w455_,
		_w3956_
	);
	LUT4 #(
		.INIT('h135f)
	) name3504 (
		\InstQueue_reg[10][6]/NET0131 ,
		\InstQueue_reg[8][6]/NET0131 ,
		_w470_,
		_w457_,
		_w3957_
	);
	LUT4 #(
		.INIT('h135f)
	) name3505 (
		\InstQueue_reg[6][6]/NET0131 ,
		\InstQueue_reg[9][6]/NET0131 ,
		_w460_,
		_w453_,
		_w3958_
	);
	LUT4 #(
		.INIT('h8000)
	) name3506 (
		_w3957_,
		_w3958_,
		_w3955_,
		_w3956_,
		_w3959_
	);
	LUT4 #(
		.INIT('h135f)
	) name3507 (
		\InstQueue_reg[15][6]/NET0131 ,
		\InstQueue_reg[1][6]/NET0131 ,
		_w477_,
		_w476_,
		_w3960_
	);
	LUT4 #(
		.INIT('h135f)
	) name3508 (
		\InstQueue_reg[0][6]/NET0131 ,
		\InstQueue_reg[11][6]/NET0131 ,
		_w461_,
		_w463_,
		_w3961_
	);
	LUT4 #(
		.INIT('h153f)
	) name3509 (
		\InstQueue_reg[14][6]/NET0131 ,
		\InstQueue_reg[7][6]/NET0131 ,
		_w468_,
		_w458_,
		_w3962_
	);
	LUT4 #(
		.INIT('h135f)
	) name3510 (
		\InstQueue_reg[13][6]/NET0131 ,
		\InstQueue_reg[4][6]/NET0131 ,
		_w471_,
		_w473_,
		_w3963_
	);
	LUT4 #(
		.INIT('h8000)
	) name3511 (
		_w3962_,
		_w3963_,
		_w3960_,
		_w3961_,
		_w3964_
	);
	LUT2 #(
		.INIT('h8)
	) name3512 (
		_w3959_,
		_w3964_,
		_w3965_
	);
	LUT4 #(
		.INIT('h0080)
	) name3513 (
		_w602_,
		_w604_,
		_w634_,
		_w3965_,
		_w3966_
	);
	LUT2 #(
		.INIT('h8)
	) name3514 (
		\Datai[6]_pad ,
		_w582_,
		_w3967_
	);
	LUT3 #(
		.INIT('h80)
	) name3515 (
		\Datai[22]_pad ,
		_w494_,
		_w586_,
		_w3968_
	);
	LUT4 #(
		.INIT('h1113)
	) name3516 (
		_w652_,
		_w3966_,
		_w3967_,
		_w3968_,
		_w3969_
	);
	LUT4 #(
		.INIT('h5700)
	) name3517 (
		\EAX_reg[22]/NET0131 ,
		_w653_,
		_w1742_,
		_w3969_,
		_w3970_
	);
	LUT4 #(
		.INIT('hecee)
	) name3518 (
		_w690_,
		_w3951_,
		_w3954_,
		_w3970_,
		_w3971_
	);
	LUT2 #(
		.INIT('h2)
	) name3519 (
		\EAX_reg[23]/NET0131 ,
		_w1841_,
		_w3972_
	);
	LUT4 #(
		.INIT('h4888)
	) name3520 (
		\EAX_reg[23]/NET0131 ,
		_w1741_,
		_w1754_,
		_w1757_,
		_w3973_
	);
	LUT4 #(
		.INIT('h88a8)
	) name3521 (
		\EAX_reg[23]/NET0131 ,
		READY_n_pad,
		_w563_,
		_w565_,
		_w3974_
	);
	LUT2 #(
		.INIT('h1)
	) name3522 (
		_w2644_,
		_w3974_,
		_w3975_
	);
	LUT2 #(
		.INIT('h2)
	) name3523 (
		_w582_,
		_w3975_,
		_w3976_
	);
	LUT4 #(
		.INIT('h7888)
	) name3524 (
		_w1771_,
		_w1776_,
		_w1781_,
		_w1786_,
		_w3977_
	);
	LUT4 #(
		.INIT('h8000)
	) name3525 (
		_w602_,
		_w604_,
		_w634_,
		_w3977_,
		_w3978_
	);
	LUT4 #(
		.INIT('h2202)
	) name3526 (
		\Datai[23]_pad ,
		READY_n_pad,
		_w563_,
		_w565_,
		_w3979_
	);
	LUT2 #(
		.INIT('h1)
	) name3527 (
		_w3974_,
		_w3979_,
		_w3980_
	);
	LUT3 #(
		.INIT('h08)
	) name3528 (
		_w494_,
		_w586_,
		_w3980_,
		_w3981_
	);
	LUT3 #(
		.INIT('h01)
	) name3529 (
		_w3978_,
		_w3981_,
		_w3976_,
		_w3982_
	);
	LUT4 #(
		.INIT('h0700)
	) name3530 (
		\EAX_reg[23]/NET0131 ,
		_w1742_,
		_w3973_,
		_w3982_,
		_w3983_
	);
	LUT3 #(
		.INIT('hce)
	) name3531 (
		_w690_,
		_w3972_,
		_w3983_,
		_w3984_
	);
	LUT4 #(
		.INIT('h1333)
	) name3532 (
		\EAX_reg[23]/NET0131 ,
		\EAX_reg[24]/NET0131 ,
		_w1754_,
		_w1757_,
		_w3985_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name3533 (
		_w1741_,
		_w1754_,
		_w1757_,
		_w1758_,
		_w3986_
	);
	LUT2 #(
		.INIT('h4)
	) name3534 (
		_w3985_,
		_w3986_,
		_w3987_
	);
	LUT4 #(
		.INIT('h88a8)
	) name3535 (
		\EAX_reg[24]/NET0131 ,
		READY_n_pad,
		_w563_,
		_w565_,
		_w3988_
	);
	LUT4 #(
		.INIT('h2202)
	) name3536 (
		\Datai[8]_pad ,
		READY_n_pad,
		_w563_,
		_w565_,
		_w3989_
	);
	LUT2 #(
		.INIT('h1)
	) name3537 (
		_w3988_,
		_w3989_,
		_w3990_
	);
	LUT2 #(
		.INIT('h2)
	) name3538 (
		_w582_,
		_w3990_,
		_w3991_
	);
	LUT2 #(
		.INIT('h9)
	) name3539 (
		_w1787_,
		_w1798_,
		_w3992_
	);
	LUT4 #(
		.INIT('h8000)
	) name3540 (
		_w602_,
		_w604_,
		_w634_,
		_w3992_,
		_w3993_
	);
	LUT4 #(
		.INIT('h2202)
	) name3541 (
		\Datai[24]_pad ,
		READY_n_pad,
		_w563_,
		_w565_,
		_w3994_
	);
	LUT2 #(
		.INIT('h1)
	) name3542 (
		_w3988_,
		_w3994_,
		_w3995_
	);
	LUT3 #(
		.INIT('h08)
	) name3543 (
		_w494_,
		_w586_,
		_w3995_,
		_w3996_
	);
	LUT3 #(
		.INIT('h01)
	) name3544 (
		_w3993_,
		_w3996_,
		_w3991_,
		_w3997_
	);
	LUT3 #(
		.INIT('h70)
	) name3545 (
		\EAX_reg[24]/NET0131 ,
		_w1742_,
		_w3997_,
		_w3998_
	);
	LUT2 #(
		.INIT('h2)
	) name3546 (
		\EAX_reg[24]/NET0131 ,
		_w1841_,
		_w3999_
	);
	LUT4 #(
		.INIT('hff8a)
	) name3547 (
		_w690_,
		_w3987_,
		_w3998_,
		_w3999_,
		_w4000_
	);
	LUT3 #(
		.INIT('h48)
	) name3548 (
		\EAX_reg[26]/NET0131 ,
		_w589_,
		_w2094_,
		_w4001_
	);
	LUT4 #(
		.INIT('h4080)
	) name3549 (
		\EAX_reg[26]/NET0131 ,
		_w589_,
		_w595_,
		_w2094_,
		_w4002_
	);
	LUT4 #(
		.INIT('hf020)
	) name3550 (
		\Datao[26]_pad ,
		_w596_,
		_w690_,
		_w4002_,
		_w4003_
	);
	LUT4 #(
		.INIT('h3f15)
	) name3551 (
		\Datao[26]_pad ,
		\uWord_reg[10]/NET0131 ,
		_w2179_,
		_w2180_,
		_w4004_
	);
	LUT2 #(
		.INIT('hb)
	) name3552 (
		_w4003_,
		_w4004_,
		_w4005_
	);
	LUT2 #(
		.INIT('h2)
	) name3553 (
		\uWord_reg[0]/NET0131 ,
		_w1841_,
		_w4006_
	);
	LUT2 #(
		.INIT('h8)
	) name3554 (
		READY_n_pad,
		\uWord_reg[0]/NET0131 ,
		_w4007_
	);
	LUT2 #(
		.INIT('h1)
	) name3555 (
		_w3824_,
		_w4007_,
		_w4008_
	);
	LUT2 #(
		.INIT('h2)
	) name3556 (
		_w582_,
		_w4008_,
		_w4009_
	);
	LUT4 #(
		.INIT('haa02)
	) name3557 (
		\uWord_reg[0]/NET0131 ,
		_w582_,
		_w589_,
		_w566_,
		_w4010_
	);
	LUT3 #(
		.INIT('ha6)
	) name3558 (
		\EAX_reg[16]/NET0131 ,
		\EAX_reg[31]/NET0131 ,
		_w2091_,
		_w4011_
	);
	LUT3 #(
		.INIT('h20)
	) name3559 (
		_w589_,
		_w566_,
		_w4011_,
		_w4012_
	);
	LUT4 #(
		.INIT('haaa8)
	) name3560 (
		_w690_,
		_w4010_,
		_w4009_,
		_w4012_,
		_w4013_
	);
	LUT2 #(
		.INIT('he)
	) name3561 (
		_w4006_,
		_w4013_,
		_w4014_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name3562 (
		\uWord_reg[10]/NET0131 ,
		_w690_,
		_w1841_,
		_w2103_,
		_w4015_
	);
	LUT2 #(
		.INIT('h2)
	) name3563 (
		\Datai[10]_pad ,
		READY_n_pad,
		_w4016_
	);
	LUT2 #(
		.INIT('h8)
	) name3564 (
		_w582_,
		_w4016_,
		_w4017_
	);
	LUT3 #(
		.INIT('ha8)
	) name3565 (
		_w2192_,
		_w4001_,
		_w4017_,
		_w4018_
	);
	LUT2 #(
		.INIT('he)
	) name3566 (
		_w4015_,
		_w4018_,
		_w4019_
	);
	LUT2 #(
		.INIT('h2)
	) name3567 (
		\uWord_reg[13]/NET0131 ,
		_w1841_,
		_w4020_
	);
	LUT2 #(
		.INIT('h1)
	) name3568 (
		\EAX_reg[29]/NET0131 ,
		_w2096_,
		_w4021_
	);
	LUT3 #(
		.INIT('h02)
	) name3569 (
		_w589_,
		_w566_,
		_w3774_,
		_w4022_
	);
	LUT2 #(
		.INIT('h8)
	) name3570 (
		READY_n_pad,
		\uWord_reg[13]/NET0131 ,
		_w4023_
	);
	LUT2 #(
		.INIT('h1)
	) name3571 (
		_w2161_,
		_w4023_,
		_w4024_
	);
	LUT2 #(
		.INIT('h2)
	) name3572 (
		_w582_,
		_w4024_,
		_w4025_
	);
	LUT4 #(
		.INIT('haa02)
	) name3573 (
		\uWord_reg[13]/NET0131 ,
		_w582_,
		_w589_,
		_w566_,
		_w4026_
	);
	LUT4 #(
		.INIT('h1011)
	) name3574 (
		_w4025_,
		_w4026_,
		_w4021_,
		_w4022_,
		_w4027_
	);
	LUT3 #(
		.INIT('hce)
	) name3575 (
		_w690_,
		_w4020_,
		_w4027_,
		_w4028_
	);
	LUT2 #(
		.INIT('h2)
	) name3576 (
		\uWord_reg[1]/NET0131 ,
		_w1841_,
		_w4029_
	);
	LUT2 #(
		.INIT('h8)
	) name3577 (
		READY_n_pad,
		\uWord_reg[1]/NET0131 ,
		_w4030_
	);
	LUT2 #(
		.INIT('h1)
	) name3578 (
		_w3752_,
		_w4030_,
		_w4031_
	);
	LUT2 #(
		.INIT('h2)
	) name3579 (
		_w582_,
		_w4031_,
		_w4032_
	);
	LUT4 #(
		.INIT('haa02)
	) name3580 (
		\uWord_reg[1]/NET0131 ,
		_w582_,
		_w589_,
		_w566_,
		_w4033_
	);
	LUT4 #(
		.INIT('hcc6c)
	) name3581 (
		\EAX_reg[16]/NET0131 ,
		\EAX_reg[17]/NET0131 ,
		\EAX_reg[31]/NET0131 ,
		_w2091_,
		_w4034_
	);
	LUT3 #(
		.INIT('h20)
	) name3582 (
		_w589_,
		_w566_,
		_w4034_,
		_w4035_
	);
	LUT4 #(
		.INIT('haaa8)
	) name3583 (
		_w690_,
		_w4032_,
		_w4033_,
		_w4035_,
		_w4036_
	);
	LUT2 #(
		.INIT('he)
	) name3584 (
		_w4029_,
		_w4036_,
		_w4037_
	);
	LUT2 #(
		.INIT('h2)
	) name3585 (
		\uWord_reg[2]/NET0131 ,
		_w1841_,
		_w4038_
	);
	LUT2 #(
		.INIT('h8)
	) name3586 (
		READY_n_pad,
		\uWord_reg[2]/NET0131 ,
		_w4039_
	);
	LUT2 #(
		.INIT('h1)
	) name3587 (
		_w3700_,
		_w4039_,
		_w4040_
	);
	LUT2 #(
		.INIT('h2)
	) name3588 (
		_w582_,
		_w4040_,
		_w4041_
	);
	LUT4 #(
		.INIT('haa02)
	) name3589 (
		\uWord_reg[2]/NET0131 ,
		_w582_,
		_w589_,
		_w566_,
		_w4042_
	);
	LUT2 #(
		.INIT('h6)
	) name3590 (
		\EAX_reg[18]/NET0131 ,
		_w2092_,
		_w4043_
	);
	LUT3 #(
		.INIT('h20)
	) name3591 (
		_w589_,
		_w566_,
		_w4043_,
		_w4044_
	);
	LUT4 #(
		.INIT('haaa8)
	) name3592 (
		_w690_,
		_w4041_,
		_w4042_,
		_w4044_,
		_w4045_
	);
	LUT2 #(
		.INIT('he)
	) name3593 (
		_w4038_,
		_w4045_,
		_w4046_
	);
	LUT2 #(
		.INIT('h2)
	) name3594 (
		\uWord_reg[5]/NET0131 ,
		_w1841_,
		_w4047_
	);
	LUT2 #(
		.INIT('h8)
	) name3595 (
		READY_n_pad,
		\uWord_reg[5]/NET0131 ,
		_w4048_
	);
	LUT2 #(
		.INIT('h1)
	) name3596 (
		_w3734_,
		_w4048_,
		_w4049_
	);
	LUT2 #(
		.INIT('h2)
	) name3597 (
		_w582_,
		_w4049_,
		_w4050_
	);
	LUT4 #(
		.INIT('haa02)
	) name3598 (
		\uWord_reg[5]/NET0131 ,
		_w582_,
		_w589_,
		_w566_,
		_w4051_
	);
	LUT2 #(
		.INIT('h1)
	) name3599 (
		\EAX_reg[21]/NET0131 ,
		_w2431_,
		_w4052_
	);
	LUT3 #(
		.INIT('h80)
	) name3600 (
		\EAX_reg[18]/NET0131 ,
		_w1756_,
		_w2092_,
		_w4053_
	);
	LUT4 #(
		.INIT('h0002)
	) name3601 (
		_w589_,
		_w566_,
		_w4053_,
		_w4052_,
		_w4054_
	);
	LUT4 #(
		.INIT('haaa8)
	) name3602 (
		_w690_,
		_w4050_,
		_w4051_,
		_w4054_,
		_w4055_
	);
	LUT2 #(
		.INIT('he)
	) name3603 (
		_w4047_,
		_w4055_,
		_w4056_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name3604 (
		\uWord_reg[6]/NET0131 ,
		_w690_,
		_w1841_,
		_w2103_,
		_w4057_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name3605 (
		\EAX_reg[18]/NET0131 ,
		\EAX_reg[22]/NET0131 ,
		_w1756_,
		_w2092_,
		_w4058_
	);
	LUT2 #(
		.INIT('h8)
	) name3606 (
		_w589_,
		_w4058_,
		_w4059_
	);
	LUT3 #(
		.INIT('h20)
	) name3607 (
		\Datai[6]_pad ,
		READY_n_pad,
		_w582_,
		_w4060_
	);
	LUT3 #(
		.INIT('ha8)
	) name3608 (
		_w2192_,
		_w4059_,
		_w4060_,
		_w4061_
	);
	LUT2 #(
		.INIT('he)
	) name3609 (
		_w4057_,
		_w4061_,
		_w4062_
	);
	LUT2 #(
		.INIT('h2)
	) name3610 (
		\uWord_reg[9]/NET0131 ,
		_w1841_,
		_w4063_
	);
	LUT2 #(
		.INIT('h6)
	) name3611 (
		\EAX_reg[25]/NET0131 ,
		_w2093_,
		_w4064_
	);
	LUT3 #(
		.INIT('h20)
	) name3612 (
		_w589_,
		_w566_,
		_w4064_,
		_w4065_
	);
	LUT2 #(
		.INIT('h8)
	) name3613 (
		_w582_,
		_w2455_,
		_w4066_
	);
	LUT4 #(
		.INIT('h000d)
	) name3614 (
		\uWord_reg[9]/NET0131 ,
		_w2103_,
		_w4065_,
		_w4066_,
		_w4067_
	);
	LUT3 #(
		.INIT('hce)
	) name3615 (
		_w690_,
		_w4063_,
		_w4067_,
		_w4068_
	);
	LUT3 #(
		.INIT('h02)
	) name3616 (
		\EBX_reg[10]/NET0131 ,
		_w1990_,
		_w1991_,
		_w4069_
	);
	LUT4 #(
		.INIT('h0080)
	) name3617 (
		_w569_,
		_w602_,
		_w634_,
		_w2700_,
		_w4070_
	);
	LUT2 #(
		.INIT('h6)
	) name3618 (
		\EBX_reg[10]/NET0131 ,
		_w1973_,
		_w4071_
	);
	LUT3 #(
		.INIT('h80)
	) name3619 (
		_w617_,
		_w621_,
		_w4071_,
		_w4072_
	);
	LUT2 #(
		.INIT('h1)
	) name3620 (
		_w4070_,
		_w4072_,
		_w4073_
	);
	LUT2 #(
		.INIT('h2)
	) name3621 (
		\EBX_reg[10]/NET0131 ,
		_w1841_,
		_w4074_
	);
	LUT4 #(
		.INIT('hff8a)
	) name3622 (
		_w690_,
		_w4069_,
		_w4073_,
		_w4074_,
		_w4075_
	);
	LUT3 #(
		.INIT('h02)
	) name3623 (
		\EBX_reg[11]/NET0131 ,
		_w1990_,
		_w1991_,
		_w4076_
	);
	LUT4 #(
		.INIT('h0080)
	) name3624 (
		_w569_,
		_w602_,
		_w634_,
		_w2718_,
		_w4077_
	);
	LUT4 #(
		.INIT('h4080)
	) name3625 (
		\EBX_reg[11]/NET0131 ,
		_w617_,
		_w621_,
		_w1974_,
		_w4078_
	);
	LUT2 #(
		.INIT('h1)
	) name3626 (
		_w4077_,
		_w4078_,
		_w4079_
	);
	LUT2 #(
		.INIT('h2)
	) name3627 (
		\EBX_reg[11]/NET0131 ,
		_w1841_,
		_w4080_
	);
	LUT4 #(
		.INIT('hff8a)
	) name3628 (
		_w690_,
		_w4076_,
		_w4079_,
		_w4080_,
		_w4081_
	);
	LUT4 #(
		.INIT('h4080)
	) name3629 (
		\EBX_reg[12]/NET0131 ,
		_w617_,
		_w621_,
		_w1975_,
		_w4082_
	);
	LUT4 #(
		.INIT('h0080)
	) name3630 (
		_w569_,
		_w602_,
		_w634_,
		_w2748_,
		_w4083_
	);
	LUT4 #(
		.INIT('h00fd)
	) name3631 (
		\EBX_reg[12]/NET0131 ,
		_w1990_,
		_w1991_,
		_w4083_,
		_w4084_
	);
	LUT2 #(
		.INIT('h2)
	) name3632 (
		\EBX_reg[12]/NET0131 ,
		_w1841_,
		_w4085_
	);
	LUT4 #(
		.INIT('hff8a)
	) name3633 (
		_w690_,
		_w4082_,
		_w4084_,
		_w4085_,
		_w4086_
	);
	LUT4 #(
		.INIT('h4080)
	) name3634 (
		\EBX_reg[14]/NET0131 ,
		_w617_,
		_w621_,
		_w1977_,
		_w4087_
	);
	LUT4 #(
		.INIT('h0080)
	) name3635 (
		_w569_,
		_w602_,
		_w634_,
		_w2786_,
		_w4088_
	);
	LUT4 #(
		.INIT('h00fd)
	) name3636 (
		\EBX_reg[14]/NET0131 ,
		_w1990_,
		_w1991_,
		_w4088_,
		_w4089_
	);
	LUT2 #(
		.INIT('h2)
	) name3637 (
		\EBX_reg[14]/NET0131 ,
		_w1841_,
		_w4090_
	);
	LUT4 #(
		.INIT('hff8a)
	) name3638 (
		_w690_,
		_w4087_,
		_w4089_,
		_w4090_,
		_w4091_
	);
	LUT4 #(
		.INIT('h4080)
	) name3639 (
		\EBX_reg[13]/NET0131 ,
		_w617_,
		_w621_,
		_w1976_,
		_w4092_
	);
	LUT4 #(
		.INIT('h0080)
	) name3640 (
		_w569_,
		_w602_,
		_w634_,
		_w2767_,
		_w4093_
	);
	LUT4 #(
		.INIT('h00fd)
	) name3641 (
		\EBX_reg[13]/NET0131 ,
		_w1990_,
		_w1991_,
		_w4093_,
		_w4094_
	);
	LUT2 #(
		.INIT('h2)
	) name3642 (
		\EBX_reg[13]/NET0131 ,
		_w1841_,
		_w4095_
	);
	LUT4 #(
		.INIT('hff8a)
	) name3643 (
		_w690_,
		_w4092_,
		_w4094_,
		_w4095_,
		_w4096_
	);
	LUT4 #(
		.INIT('h4080)
	) name3644 (
		\EBX_reg[15]/NET0131 ,
		_w617_,
		_w621_,
		_w1978_,
		_w4097_
	);
	LUT4 #(
		.INIT('h0080)
	) name3645 (
		_w569_,
		_w602_,
		_w634_,
		_w2807_,
		_w4098_
	);
	LUT4 #(
		.INIT('h00fd)
	) name3646 (
		\EBX_reg[15]/NET0131 ,
		_w1990_,
		_w1991_,
		_w4098_,
		_w4099_
	);
	LUT2 #(
		.INIT('h2)
	) name3647 (
		\EBX_reg[15]/NET0131 ,
		_w1841_,
		_w4100_
	);
	LUT4 #(
		.INIT('hff8a)
	) name3648 (
		_w690_,
		_w4097_,
		_w4099_,
		_w4100_,
		_w4101_
	);
	LUT4 #(
		.INIT('h4080)
	) name3649 (
		\EBX_reg[16]/NET0131 ,
		_w617_,
		_w621_,
		_w1979_,
		_w4102_
	);
	LUT4 #(
		.INIT('h0080)
	) name3650 (
		_w569_,
		_w602_,
		_w634_,
		_w3822_,
		_w4103_
	);
	LUT4 #(
		.INIT('h00fd)
	) name3651 (
		\EBX_reg[16]/NET0131 ,
		_w1990_,
		_w1991_,
		_w4103_,
		_w4104_
	);
	LUT2 #(
		.INIT('h2)
	) name3652 (
		\EBX_reg[16]/NET0131 ,
		_w1841_,
		_w4105_
	);
	LUT4 #(
		.INIT('hff8a)
	) name3653 (
		_w690_,
		_w4102_,
		_w4104_,
		_w4105_,
		_w4106_
	);
	LUT3 #(
		.INIT('h48)
	) name3654 (
		\EBX_reg[17]/NET0131 ,
		_w622_,
		_w1980_,
		_w4107_
	);
	LUT4 #(
		.INIT('h0080)
	) name3655 (
		_w569_,
		_w602_,
		_w634_,
		_w3847_,
		_w4108_
	);
	LUT4 #(
		.INIT('h00fd)
	) name3656 (
		\EBX_reg[17]/NET0131 ,
		_w1990_,
		_w1991_,
		_w4108_,
		_w4109_
	);
	LUT2 #(
		.INIT('h2)
	) name3657 (
		\EBX_reg[17]/NET0131 ,
		_w1841_,
		_w4110_
	);
	LUT4 #(
		.INIT('hff8a)
	) name3658 (
		_w690_,
		_w4107_,
		_w4109_,
		_w4110_,
		_w4111_
	);
	LUT3 #(
		.INIT('h48)
	) name3659 (
		\EBX_reg[18]/NET0131 ,
		_w622_,
		_w1981_,
		_w4112_
	);
	LUT4 #(
		.INIT('h0080)
	) name3660 (
		_w569_,
		_w602_,
		_w634_,
		_w3869_,
		_w4113_
	);
	LUT4 #(
		.INIT('h00fd)
	) name3661 (
		\EBX_reg[18]/NET0131 ,
		_w1990_,
		_w1991_,
		_w4113_,
		_w4114_
	);
	LUT2 #(
		.INIT('h2)
	) name3662 (
		\EBX_reg[18]/NET0131 ,
		_w1841_,
		_w4115_
	);
	LUT4 #(
		.INIT('hff8a)
	) name3663 (
		_w690_,
		_w4112_,
		_w4114_,
		_w4115_,
		_w4116_
	);
	LUT3 #(
		.INIT('h48)
	) name3664 (
		\EBX_reg[19]/NET0131 ,
		_w622_,
		_w1982_,
		_w4117_
	);
	LUT4 #(
		.INIT('h0080)
	) name3665 (
		_w569_,
		_w602_,
		_w634_,
		_w3891_,
		_w4118_
	);
	LUT4 #(
		.INIT('h00fd)
	) name3666 (
		\EBX_reg[19]/NET0131 ,
		_w1990_,
		_w1991_,
		_w4118_,
		_w4119_
	);
	LUT2 #(
		.INIT('h2)
	) name3667 (
		\EBX_reg[19]/NET0131 ,
		_w1841_,
		_w4120_
	);
	LUT4 #(
		.INIT('hff8a)
	) name3668 (
		_w690_,
		_w4117_,
		_w4119_,
		_w4120_,
		_w4121_
	);
	LUT3 #(
		.INIT('h80)
	) name3669 (
		\EBX_reg[19]/NET0131 ,
		\EBX_reg[20]/NET0131 ,
		_w1982_,
		_w4122_
	);
	LUT4 #(
		.INIT('h60c0)
	) name3670 (
		\EBX_reg[19]/NET0131 ,
		\EBX_reg[20]/NET0131 ,
		_w622_,
		_w1982_,
		_w4123_
	);
	LUT4 #(
		.INIT('h0080)
	) name3671 (
		_w569_,
		_w602_,
		_w634_,
		_w3917_,
		_w4124_
	);
	LUT4 #(
		.INIT('h00fd)
	) name3672 (
		\EBX_reg[20]/NET0131 ,
		_w1990_,
		_w1991_,
		_w4124_,
		_w4125_
	);
	LUT2 #(
		.INIT('h2)
	) name3673 (
		\EBX_reg[20]/NET0131 ,
		_w1841_,
		_w4126_
	);
	LUT4 #(
		.INIT('hff8a)
	) name3674 (
		_w690_,
		_w4123_,
		_w4125_,
		_w4126_,
		_w4127_
	);
	LUT4 #(
		.INIT('h8000)
	) name3675 (
		\EBX_reg[19]/NET0131 ,
		\EBX_reg[20]/NET0131 ,
		\EBX_reg[21]/NET0131 ,
		_w1982_,
		_w4128_
	);
	LUT4 #(
		.INIT('h0080)
	) name3676 (
		_w569_,
		_w602_,
		_w634_,
		_w3944_,
		_w4129_
	);
	LUT4 #(
		.INIT('h00fd)
	) name3677 (
		\EBX_reg[21]/NET0131 ,
		_w1990_,
		_w1991_,
		_w4129_,
		_w4130_
	);
	LUT4 #(
		.INIT('hb700)
	) name3678 (
		\EBX_reg[21]/NET0131 ,
		_w622_,
		_w4122_,
		_w4130_,
		_w4131_
	);
	LUT2 #(
		.INIT('h2)
	) name3679 (
		\EBX_reg[21]/NET0131 ,
		_w1841_,
		_w4132_
	);
	LUT3 #(
		.INIT('hf2)
	) name3680 (
		_w690_,
		_w4131_,
		_w4132_,
		_w4133_
	);
	LUT4 #(
		.INIT('h0080)
	) name3681 (
		_w569_,
		_w602_,
		_w634_,
		_w3965_,
		_w4134_
	);
	LUT4 #(
		.INIT('h00fd)
	) name3682 (
		\EBX_reg[22]/NET0131 ,
		_w1990_,
		_w1991_,
		_w4134_,
		_w4135_
	);
	LUT4 #(
		.INIT('hb700)
	) name3683 (
		\EBX_reg[22]/NET0131 ,
		_w622_,
		_w4128_,
		_w4135_,
		_w4136_
	);
	LUT2 #(
		.INIT('h2)
	) name3684 (
		\EBX_reg[22]/NET0131 ,
		_w1841_,
		_w4137_
	);
	LUT3 #(
		.INIT('hf2)
	) name3685 (
		_w690_,
		_w4136_,
		_w4137_,
		_w4138_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name3686 (
		\EBX_reg[19]/NET0131 ,
		_w622_,
		_w1982_,
		_w1983_,
		_w4139_
	);
	LUT4 #(
		.INIT('hec00)
	) name3687 (
		\EBX_reg[22]/NET0131 ,
		\EBX_reg[23]/NET0131 ,
		_w4128_,
		_w4139_,
		_w4140_
	);
	LUT4 #(
		.INIT('h8000)
	) name3688 (
		_w569_,
		_w602_,
		_w634_,
		_w3977_,
		_w4141_
	);
	LUT4 #(
		.INIT('h00fd)
	) name3689 (
		\EBX_reg[23]/NET0131 ,
		_w1990_,
		_w1991_,
		_w4141_,
		_w4142_
	);
	LUT2 #(
		.INIT('h2)
	) name3690 (
		\EBX_reg[23]/NET0131 ,
		_w1841_,
		_w4143_
	);
	LUT4 #(
		.INIT('hff8a)
	) name3691 (
		_w690_,
		_w4140_,
		_w4142_,
		_w4143_,
		_w4144_
	);
	LUT4 #(
		.INIT('h8000)
	) name3692 (
		_w569_,
		_w602_,
		_w634_,
		_w3992_,
		_w4145_
	);
	LUT4 #(
		.INIT('h00fd)
	) name3693 (
		\EBX_reg[24]/NET0131 ,
		_w1990_,
		_w1991_,
		_w4145_,
		_w4146_
	);
	LUT4 #(
		.INIT('hb700)
	) name3694 (
		\EBX_reg[24]/NET0131 ,
		_w622_,
		_w1984_,
		_w4146_,
		_w4147_
	);
	LUT2 #(
		.INIT('h2)
	) name3695 (
		\EBX_reg[24]/NET0131 ,
		_w1841_,
		_w4148_
	);
	LUT3 #(
		.INIT('hf2)
	) name3696 (
		_w690_,
		_w4147_,
		_w4148_,
		_w4149_
	);
	LUT3 #(
		.INIT('h02)
	) name3697 (
		\EBX_reg[8]/NET0131 ,
		_w1990_,
		_w1991_,
		_w4150_
	);
	LUT4 #(
		.INIT('h0080)
	) name3698 (
		_w569_,
		_w602_,
		_w634_,
		_w2661_,
		_w4151_
	);
	LUT3 #(
		.INIT('h6c)
	) name3699 (
		\EBX_reg[7]/NET0131 ,
		\EBX_reg[8]/NET0131 ,
		_w1972_,
		_w4152_
	);
	LUT3 #(
		.INIT('h80)
	) name3700 (
		_w617_,
		_w621_,
		_w4152_,
		_w4153_
	);
	LUT2 #(
		.INIT('h1)
	) name3701 (
		_w4151_,
		_w4153_,
		_w4154_
	);
	LUT2 #(
		.INIT('h2)
	) name3702 (
		\EBX_reg[8]/NET0131 ,
		_w1841_,
		_w4155_
	);
	LUT4 #(
		.INIT('hff8a)
	) name3703 (
		_w690_,
		_w4150_,
		_w4154_,
		_w4155_,
		_w4156_
	);
	LUT3 #(
		.INIT('h02)
	) name3704 (
		\EBX_reg[9]/NET0131 ,
		_w1990_,
		_w1991_,
		_w4157_
	);
	LUT4 #(
		.INIT('h0080)
	) name3705 (
		_w569_,
		_w602_,
		_w634_,
		_w2678_,
		_w4158_
	);
	LUT4 #(
		.INIT('h78f0)
	) name3706 (
		\EBX_reg[7]/NET0131 ,
		\EBX_reg[8]/NET0131 ,
		\EBX_reg[9]/NET0131 ,
		_w1972_,
		_w4159_
	);
	LUT3 #(
		.INIT('h80)
	) name3707 (
		_w617_,
		_w621_,
		_w4159_,
		_w4160_
	);
	LUT2 #(
		.INIT('h1)
	) name3708 (
		_w4158_,
		_w4160_,
		_w4161_
	);
	LUT2 #(
		.INIT('h2)
	) name3709 (
		\EBX_reg[9]/NET0131 ,
		_w1841_,
		_w4162_
	);
	LUT4 #(
		.INIT('hff8a)
	) name3710 (
		_w690_,
		_w4157_,
		_w4161_,
		_w4162_,
		_w4163_
	);
	LUT4 #(
		.INIT('h2f00)
	) name3711 (
		\Flush_reg/NET0131 ,
		_w670_,
		_w675_,
		_w690_,
		_w4164_
	);
	LUT2 #(
		.INIT('h2)
	) name3712 (
		\Flush_reg/NET0131 ,
		_w1841_,
		_w4165_
	);
	LUT2 #(
		.INIT('he)
	) name3713 (
		_w4164_,
		_w4165_,
		_w4166_
	);
	LUT4 #(
		.INIT('h60c0)
	) name3714 (
		\Datai[25]_pad ,
		\Datai[26]_pad ,
		_w2199_,
		_w2208_,
		_w4167_
	);
	LUT3 #(
		.INIT('h60)
	) name3715 (
		\Datai[18]_pad ,
		_w2211_,
		_w2215_,
		_w4168_
	);
	LUT4 #(
		.INIT('h5553)
	) name3716 (
		\Datai[2]_pad ,
		\InstQueue_reg[0][2]/NET0131 ,
		_w2217_,
		_w2219_,
		_w4169_
	);
	LUT2 #(
		.INIT('h1)
	) name3717 (
		_w2223_,
		_w4169_,
		_w4170_
	);
	LUT4 #(
		.INIT('h0057)
	) name3718 (
		\DataWidth_reg[1]/NET0131 ,
		_w4167_,
		_w4168_,
		_w4170_,
		_w4171_
	);
	LUT4 #(
		.INIT('hc055)
	) name3719 (
		\InstQueue_reg[0][2]/NET0131 ,
		_w466_,
		_w479_,
		_w2217_,
		_w4172_
	);
	LUT2 #(
		.INIT('h2)
	) name3720 (
		\InstQueue_reg[0][2]/NET0131 ,
		_w2227_,
		_w4173_
	);
	LUT3 #(
		.INIT('h0d)
	) name3721 (
		_w1212_,
		_w4169_,
		_w4173_,
		_w4174_
	);
	LUT3 #(
		.INIT('hd0)
	) name3722 (
		_w710_,
		_w4172_,
		_w4174_,
		_w4175_
	);
	LUT3 #(
		.INIT('h2f)
	) name3723 (
		_w695_,
		_w4171_,
		_w4175_,
		_w4176_
	);
	LUT4 #(
		.INIT('h6c00)
	) name3724 (
		\Datai[25]_pad ,
		\Datai[26]_pad ,
		_w2208_,
		_w2232_,
		_w4177_
	);
	LUT3 #(
		.INIT('h60)
	) name3725 (
		\Datai[18]_pad ,
		_w2211_,
		_w2234_,
		_w4178_
	);
	LUT4 #(
		.INIT('h5553)
	) name3726 (
		\Datai[2]_pad ,
		\InstQueue_reg[10][2]/NET0131 ,
		_w2236_,
		_w2237_,
		_w4179_
	);
	LUT2 #(
		.INIT('h1)
	) name3727 (
		_w2241_,
		_w4179_,
		_w4180_
	);
	LUT4 #(
		.INIT('h0057)
	) name3728 (
		\DataWidth_reg[1]/NET0131 ,
		_w4177_,
		_w4178_,
		_w4180_,
		_w4181_
	);
	LUT4 #(
		.INIT('hc055)
	) name3729 (
		\InstQueue_reg[10][2]/NET0131 ,
		_w466_,
		_w479_,
		_w2236_,
		_w4182_
	);
	LUT2 #(
		.INIT('h2)
	) name3730 (
		\InstQueue_reg[10][2]/NET0131 ,
		_w2227_,
		_w4183_
	);
	LUT3 #(
		.INIT('h0d)
	) name3731 (
		_w1212_,
		_w4179_,
		_w4183_,
		_w4184_
	);
	LUT3 #(
		.INIT('hd0)
	) name3732 (
		_w710_,
		_w4182_,
		_w4184_,
		_w4185_
	);
	LUT3 #(
		.INIT('h2f)
	) name3733 (
		_w695_,
		_w4181_,
		_w4185_,
		_w4186_
	);
	LUT4 #(
		.INIT('h6c00)
	) name3734 (
		\Datai[25]_pad ,
		\Datai[26]_pad ,
		_w2208_,
		_w2234_,
		_w4187_
	);
	LUT3 #(
		.INIT('h60)
	) name3735 (
		\Datai[18]_pad ,
		_w2211_,
		_w2237_,
		_w4188_
	);
	LUT4 #(
		.INIT('h5553)
	) name3736 (
		\Datai[2]_pad ,
		\InstQueue_reg[11][2]/NET0131 ,
		_w2236_,
		_w2251_,
		_w4189_
	);
	LUT2 #(
		.INIT('h1)
	) name3737 (
		_w2255_,
		_w4189_,
		_w4190_
	);
	LUT4 #(
		.INIT('h0057)
	) name3738 (
		\DataWidth_reg[1]/NET0131 ,
		_w4187_,
		_w4188_,
		_w4190_,
		_w4191_
	);
	LUT4 #(
		.INIT('hc055)
	) name3739 (
		\InstQueue_reg[11][2]/NET0131 ,
		_w466_,
		_w479_,
		_w2251_,
		_w4192_
	);
	LUT2 #(
		.INIT('h2)
	) name3740 (
		\InstQueue_reg[11][2]/NET0131 ,
		_w2227_,
		_w4193_
	);
	LUT3 #(
		.INIT('h0d)
	) name3741 (
		_w1212_,
		_w4189_,
		_w4193_,
		_w4194_
	);
	LUT3 #(
		.INIT('hd0)
	) name3742 (
		_w710_,
		_w4192_,
		_w4194_,
		_w4195_
	);
	LUT3 #(
		.INIT('h2f)
	) name3743 (
		_w695_,
		_w4191_,
		_w4195_,
		_w4196_
	);
	LUT4 #(
		.INIT('h6c00)
	) name3744 (
		\Datai[25]_pad ,
		\Datai[26]_pad ,
		_w2208_,
		_w2237_,
		_w4197_
	);
	LUT3 #(
		.INIT('h60)
	) name3745 (
		\Datai[18]_pad ,
		_w2211_,
		_w2236_,
		_w4198_
	);
	LUT4 #(
		.INIT('h5553)
	) name3746 (
		\Datai[2]_pad ,
		\InstQueue_reg[12][2]/NET0131 ,
		_w2251_,
		_w2265_,
		_w4199_
	);
	LUT2 #(
		.INIT('h1)
	) name3747 (
		_w2268_,
		_w4199_,
		_w4200_
	);
	LUT4 #(
		.INIT('h0057)
	) name3748 (
		\DataWidth_reg[1]/NET0131 ,
		_w4197_,
		_w4198_,
		_w4200_,
		_w4201_
	);
	LUT4 #(
		.INIT('hc055)
	) name3749 (
		\InstQueue_reg[12][2]/NET0131 ,
		_w466_,
		_w479_,
		_w2265_,
		_w4202_
	);
	LUT2 #(
		.INIT('h2)
	) name3750 (
		\InstQueue_reg[12][2]/NET0131 ,
		_w2227_,
		_w4203_
	);
	LUT3 #(
		.INIT('h0d)
	) name3751 (
		_w1212_,
		_w4199_,
		_w4203_,
		_w4204_
	);
	LUT3 #(
		.INIT('hd0)
	) name3752 (
		_w710_,
		_w4202_,
		_w4204_,
		_w4205_
	);
	LUT3 #(
		.INIT('h2f)
	) name3753 (
		_w695_,
		_w4201_,
		_w4205_,
		_w4206_
	);
	LUT4 #(
		.INIT('h6c00)
	) name3754 (
		\Datai[25]_pad ,
		\Datai[26]_pad ,
		_w2208_,
		_w2236_,
		_w4207_
	);
	LUT3 #(
		.INIT('h60)
	) name3755 (
		\Datai[18]_pad ,
		_w2211_,
		_w2251_,
		_w4208_
	);
	LUT4 #(
		.INIT('h5553)
	) name3756 (
		\Datai[2]_pad ,
		\InstQueue_reg[13][2]/NET0131 ,
		_w2199_,
		_w2265_,
		_w4209_
	);
	LUT2 #(
		.INIT('h1)
	) name3757 (
		_w2280_,
		_w4209_,
		_w4210_
	);
	LUT4 #(
		.INIT('h0057)
	) name3758 (
		\DataWidth_reg[1]/NET0131 ,
		_w4207_,
		_w4208_,
		_w4210_,
		_w4211_
	);
	LUT4 #(
		.INIT('hc055)
	) name3759 (
		\InstQueue_reg[13][2]/NET0131 ,
		_w466_,
		_w479_,
		_w2199_,
		_w4212_
	);
	LUT2 #(
		.INIT('h2)
	) name3760 (
		\InstQueue_reg[13][2]/NET0131 ,
		_w2227_,
		_w4213_
	);
	LUT3 #(
		.INIT('h0d)
	) name3761 (
		_w1212_,
		_w4209_,
		_w4213_,
		_w4214_
	);
	LUT3 #(
		.INIT('hd0)
	) name3762 (
		_w710_,
		_w4212_,
		_w4214_,
		_w4215_
	);
	LUT3 #(
		.INIT('h2f)
	) name3763 (
		_w695_,
		_w4211_,
		_w4215_,
		_w4216_
	);
	LUT4 #(
		.INIT('h6c00)
	) name3764 (
		\Datai[25]_pad ,
		\Datai[26]_pad ,
		_w2208_,
		_w2251_,
		_w4217_
	);
	LUT3 #(
		.INIT('h60)
	) name3765 (
		\Datai[18]_pad ,
		_w2211_,
		_w2265_,
		_w4218_
	);
	LUT4 #(
		.INIT('h5553)
	) name3766 (
		\Datai[2]_pad ,
		\InstQueue_reg[14][2]/NET0131 ,
		_w2199_,
		_w2215_,
		_w4219_
	);
	LUT2 #(
		.INIT('h1)
	) name3767 (
		_w2291_,
		_w4219_,
		_w4220_
	);
	LUT4 #(
		.INIT('h0057)
	) name3768 (
		\DataWidth_reg[1]/NET0131 ,
		_w4217_,
		_w4218_,
		_w4220_,
		_w4221_
	);
	LUT4 #(
		.INIT('hc055)
	) name3769 (
		\InstQueue_reg[14][2]/NET0131 ,
		_w466_,
		_w479_,
		_w2215_,
		_w4222_
	);
	LUT2 #(
		.INIT('h2)
	) name3770 (
		\InstQueue_reg[14][2]/NET0131 ,
		_w2227_,
		_w4223_
	);
	LUT3 #(
		.INIT('h0d)
	) name3771 (
		_w1212_,
		_w4219_,
		_w4223_,
		_w4224_
	);
	LUT3 #(
		.INIT('hd0)
	) name3772 (
		_w710_,
		_w4222_,
		_w4224_,
		_w4225_
	);
	LUT3 #(
		.INIT('h2f)
	) name3773 (
		_w695_,
		_w4221_,
		_w4225_,
		_w4226_
	);
	LUT4 #(
		.INIT('h6c00)
	) name3774 (
		\Datai[25]_pad ,
		\Datai[26]_pad ,
		_w2208_,
		_w2265_,
		_w4227_
	);
	LUT3 #(
		.INIT('h48)
	) name3775 (
		\Datai[18]_pad ,
		_w2199_,
		_w2211_,
		_w4228_
	);
	LUT4 #(
		.INIT('h5553)
	) name3776 (
		\Datai[2]_pad ,
		\InstQueue_reg[15][2]/NET0131 ,
		_w2219_,
		_w2215_,
		_w4229_
	);
	LUT2 #(
		.INIT('h1)
	) name3777 (
		_w2303_,
		_w4229_,
		_w4230_
	);
	LUT4 #(
		.INIT('h0057)
	) name3778 (
		\DataWidth_reg[1]/NET0131 ,
		_w4227_,
		_w4228_,
		_w4230_,
		_w4231_
	);
	LUT4 #(
		.INIT('hc055)
	) name3779 (
		\InstQueue_reg[15][2]/NET0131 ,
		_w466_,
		_w479_,
		_w2219_,
		_w4232_
	);
	LUT2 #(
		.INIT('h2)
	) name3780 (
		\InstQueue_reg[15][2]/NET0131 ,
		_w2227_,
		_w4233_
	);
	LUT3 #(
		.INIT('h0d)
	) name3781 (
		_w1212_,
		_w4229_,
		_w4233_,
		_w4234_
	);
	LUT3 #(
		.INIT('hd0)
	) name3782 (
		_w710_,
		_w4232_,
		_w4234_,
		_w4235_
	);
	LUT3 #(
		.INIT('h2f)
	) name3783 (
		_w695_,
		_w4231_,
		_w4235_,
		_w4236_
	);
	LUT4 #(
		.INIT('h6c00)
	) name3784 (
		\Datai[25]_pad ,
		\Datai[26]_pad ,
		_w2208_,
		_w2215_,
		_w4237_
	);
	LUT3 #(
		.INIT('h48)
	) name3785 (
		\Datai[18]_pad ,
		_w2219_,
		_w2211_,
		_w4238_
	);
	LUT4 #(
		.INIT('h5553)
	) name3786 (
		\Datai[2]_pad ,
		\InstQueue_reg[1][2]/NET0131 ,
		_w2217_,
		_w2313_,
		_w4239_
	);
	LUT2 #(
		.INIT('h1)
	) name3787 (
		_w2316_,
		_w4239_,
		_w4240_
	);
	LUT4 #(
		.INIT('h0057)
	) name3788 (
		\DataWidth_reg[1]/NET0131 ,
		_w4237_,
		_w4238_,
		_w4240_,
		_w4241_
	);
	LUT4 #(
		.INIT('hc055)
	) name3789 (
		\InstQueue_reg[1][2]/NET0131 ,
		_w466_,
		_w479_,
		_w2313_,
		_w4242_
	);
	LUT2 #(
		.INIT('h2)
	) name3790 (
		\InstQueue_reg[1][2]/NET0131 ,
		_w2227_,
		_w4243_
	);
	LUT3 #(
		.INIT('h0d)
	) name3791 (
		_w1212_,
		_w4239_,
		_w4243_,
		_w4244_
	);
	LUT3 #(
		.INIT('hd0)
	) name3792 (
		_w710_,
		_w4242_,
		_w4244_,
		_w4245_
	);
	LUT3 #(
		.INIT('h2f)
	) name3793 (
		_w695_,
		_w4241_,
		_w4245_,
		_w4246_
	);
	LUT3 #(
		.INIT('h48)
	) name3794 (
		\Datai[18]_pad ,
		_w2217_,
		_w2211_,
		_w4247_
	);
	LUT4 #(
		.INIT('h60c0)
	) name3795 (
		\Datai[25]_pad ,
		\Datai[26]_pad ,
		_w2219_,
		_w2208_,
		_w4248_
	);
	LUT4 #(
		.INIT('h5553)
	) name3796 (
		\Datai[2]_pad ,
		\InstQueue_reg[2][2]/NET0131 ,
		_w2313_,
		_w2326_,
		_w4249_
	);
	LUT2 #(
		.INIT('h1)
	) name3797 (
		_w2329_,
		_w4249_,
		_w4250_
	);
	LUT4 #(
		.INIT('h0057)
	) name3798 (
		\DataWidth_reg[1]/NET0131 ,
		_w4247_,
		_w4248_,
		_w4250_,
		_w4251_
	);
	LUT4 #(
		.INIT('hc055)
	) name3799 (
		\InstQueue_reg[2][2]/NET0131 ,
		_w466_,
		_w479_,
		_w2326_,
		_w4252_
	);
	LUT2 #(
		.INIT('h2)
	) name3800 (
		\InstQueue_reg[2][2]/NET0131 ,
		_w2227_,
		_w4253_
	);
	LUT3 #(
		.INIT('h0d)
	) name3801 (
		_w1212_,
		_w4249_,
		_w4253_,
		_w4254_
	);
	LUT3 #(
		.INIT('hd0)
	) name3802 (
		_w710_,
		_w4252_,
		_w4254_,
		_w4255_
	);
	LUT3 #(
		.INIT('h2f)
	) name3803 (
		_w695_,
		_w4251_,
		_w4255_,
		_w4256_
	);
	LUT4 #(
		.INIT('h60c0)
	) name3804 (
		\Datai[25]_pad ,
		\Datai[26]_pad ,
		_w2217_,
		_w2208_,
		_w4257_
	);
	LUT3 #(
		.INIT('h60)
	) name3805 (
		\Datai[18]_pad ,
		_w2211_,
		_w2313_,
		_w4258_
	);
	LUT4 #(
		.INIT('h5553)
	) name3806 (
		\Datai[2]_pad ,
		\InstQueue_reg[3][2]/NET0131 ,
		_w2326_,
		_w2339_,
		_w4259_
	);
	LUT2 #(
		.INIT('h1)
	) name3807 (
		_w2342_,
		_w4259_,
		_w4260_
	);
	LUT4 #(
		.INIT('h0057)
	) name3808 (
		\DataWidth_reg[1]/NET0131 ,
		_w4257_,
		_w4258_,
		_w4260_,
		_w4261_
	);
	LUT4 #(
		.INIT('hc055)
	) name3809 (
		\InstQueue_reg[3][2]/NET0131 ,
		_w466_,
		_w479_,
		_w2339_,
		_w4262_
	);
	LUT2 #(
		.INIT('h2)
	) name3810 (
		\InstQueue_reg[3][2]/NET0131 ,
		_w2227_,
		_w4263_
	);
	LUT3 #(
		.INIT('h0d)
	) name3811 (
		_w1212_,
		_w4259_,
		_w4263_,
		_w4264_
	);
	LUT3 #(
		.INIT('hd0)
	) name3812 (
		_w710_,
		_w4262_,
		_w4264_,
		_w4265_
	);
	LUT3 #(
		.INIT('h2f)
	) name3813 (
		_w695_,
		_w4261_,
		_w4265_,
		_w4266_
	);
	LUT4 #(
		.INIT('h6c00)
	) name3814 (
		\Datai[25]_pad ,
		\Datai[26]_pad ,
		_w2208_,
		_w2313_,
		_w4267_
	);
	LUT3 #(
		.INIT('h60)
	) name3815 (
		\Datai[18]_pad ,
		_w2211_,
		_w2326_,
		_w4268_
	);
	LUT4 #(
		.INIT('h5553)
	) name3816 (
		\Datai[2]_pad ,
		\InstQueue_reg[4][2]/NET0131 ,
		_w2339_,
		_w2352_,
		_w4269_
	);
	LUT2 #(
		.INIT('h1)
	) name3817 (
		_w2355_,
		_w4269_,
		_w4270_
	);
	LUT4 #(
		.INIT('h0057)
	) name3818 (
		\DataWidth_reg[1]/NET0131 ,
		_w4267_,
		_w4268_,
		_w4270_,
		_w4271_
	);
	LUT4 #(
		.INIT('hc055)
	) name3819 (
		\InstQueue_reg[4][2]/NET0131 ,
		_w466_,
		_w479_,
		_w2352_,
		_w4272_
	);
	LUT2 #(
		.INIT('h2)
	) name3820 (
		\InstQueue_reg[4][2]/NET0131 ,
		_w2227_,
		_w4273_
	);
	LUT3 #(
		.INIT('h0d)
	) name3821 (
		_w1212_,
		_w4269_,
		_w4273_,
		_w4274_
	);
	LUT3 #(
		.INIT('hd0)
	) name3822 (
		_w710_,
		_w4272_,
		_w4274_,
		_w4275_
	);
	LUT3 #(
		.INIT('h2f)
	) name3823 (
		_w695_,
		_w4271_,
		_w4275_,
		_w4276_
	);
	LUT4 #(
		.INIT('h6c00)
	) name3824 (
		\Datai[25]_pad ,
		\Datai[26]_pad ,
		_w2208_,
		_w2326_,
		_w4277_
	);
	LUT3 #(
		.INIT('h60)
	) name3825 (
		\Datai[18]_pad ,
		_w2211_,
		_w2339_,
		_w4278_
	);
	LUT4 #(
		.INIT('h5553)
	) name3826 (
		\Datai[2]_pad ,
		\InstQueue_reg[5][2]/NET0131 ,
		_w2352_,
		_w2365_,
		_w4279_
	);
	LUT2 #(
		.INIT('h1)
	) name3827 (
		_w2368_,
		_w4279_,
		_w4280_
	);
	LUT4 #(
		.INIT('h0057)
	) name3828 (
		\DataWidth_reg[1]/NET0131 ,
		_w4277_,
		_w4278_,
		_w4280_,
		_w4281_
	);
	LUT4 #(
		.INIT('hc055)
	) name3829 (
		\InstQueue_reg[5][2]/NET0131 ,
		_w466_,
		_w479_,
		_w2365_,
		_w4282_
	);
	LUT2 #(
		.INIT('h2)
	) name3830 (
		\InstQueue_reg[5][2]/NET0131 ,
		_w2227_,
		_w4283_
	);
	LUT3 #(
		.INIT('h0d)
	) name3831 (
		_w1212_,
		_w4279_,
		_w4283_,
		_w4284_
	);
	LUT3 #(
		.INIT('hd0)
	) name3832 (
		_w710_,
		_w4282_,
		_w4284_,
		_w4285_
	);
	LUT3 #(
		.INIT('h2f)
	) name3833 (
		_w695_,
		_w4281_,
		_w4285_,
		_w4286_
	);
	LUT4 #(
		.INIT('h6c00)
	) name3834 (
		\Datai[25]_pad ,
		\Datai[26]_pad ,
		_w2208_,
		_w2339_,
		_w4287_
	);
	LUT3 #(
		.INIT('h60)
	) name3835 (
		\Datai[18]_pad ,
		_w2211_,
		_w2352_,
		_w4288_
	);
	LUT4 #(
		.INIT('h5553)
	) name3836 (
		\Datai[2]_pad ,
		\InstQueue_reg[6][2]/NET0131 ,
		_w2365_,
		_w2378_,
		_w4289_
	);
	LUT2 #(
		.INIT('h1)
	) name3837 (
		_w2381_,
		_w4289_,
		_w4290_
	);
	LUT4 #(
		.INIT('h0057)
	) name3838 (
		\DataWidth_reg[1]/NET0131 ,
		_w4287_,
		_w4288_,
		_w4290_,
		_w4291_
	);
	LUT4 #(
		.INIT('hc055)
	) name3839 (
		\InstQueue_reg[6][2]/NET0131 ,
		_w466_,
		_w479_,
		_w2378_,
		_w4292_
	);
	LUT2 #(
		.INIT('h2)
	) name3840 (
		\InstQueue_reg[6][2]/NET0131 ,
		_w2227_,
		_w4293_
	);
	LUT3 #(
		.INIT('h0d)
	) name3841 (
		_w1212_,
		_w4289_,
		_w4293_,
		_w4294_
	);
	LUT3 #(
		.INIT('hd0)
	) name3842 (
		_w710_,
		_w4292_,
		_w4294_,
		_w4295_
	);
	LUT3 #(
		.INIT('h2f)
	) name3843 (
		_w695_,
		_w4291_,
		_w4295_,
		_w4296_
	);
	LUT4 #(
		.INIT('h6c00)
	) name3844 (
		\Datai[25]_pad ,
		\Datai[26]_pad ,
		_w2208_,
		_w2352_,
		_w4297_
	);
	LUT3 #(
		.INIT('h60)
	) name3845 (
		\Datai[18]_pad ,
		_w2211_,
		_w2365_,
		_w4298_
	);
	LUT4 #(
		.INIT('h5553)
	) name3846 (
		\Datai[2]_pad ,
		\InstQueue_reg[7][2]/NET0131 ,
		_w2232_,
		_w2378_,
		_w4299_
	);
	LUT2 #(
		.INIT('h1)
	) name3847 (
		_w2393_,
		_w4299_,
		_w4300_
	);
	LUT4 #(
		.INIT('h0057)
	) name3848 (
		\DataWidth_reg[1]/NET0131 ,
		_w4297_,
		_w4298_,
		_w4300_,
		_w4301_
	);
	LUT4 #(
		.INIT('hc055)
	) name3849 (
		\InstQueue_reg[7][2]/NET0131 ,
		_w466_,
		_w479_,
		_w2232_,
		_w4302_
	);
	LUT2 #(
		.INIT('h2)
	) name3850 (
		\InstQueue_reg[7][2]/NET0131 ,
		_w2227_,
		_w4303_
	);
	LUT3 #(
		.INIT('h0d)
	) name3851 (
		_w1212_,
		_w4299_,
		_w4303_,
		_w4304_
	);
	LUT3 #(
		.INIT('hd0)
	) name3852 (
		_w710_,
		_w4302_,
		_w4304_,
		_w4305_
	);
	LUT3 #(
		.INIT('h2f)
	) name3853 (
		_w695_,
		_w4301_,
		_w4305_,
		_w4306_
	);
	LUT4 #(
		.INIT('h6c00)
	) name3854 (
		\Datai[25]_pad ,
		\Datai[26]_pad ,
		_w2208_,
		_w2365_,
		_w4307_
	);
	LUT3 #(
		.INIT('h60)
	) name3855 (
		\Datai[18]_pad ,
		_w2211_,
		_w2378_,
		_w4308_
	);
	LUT4 #(
		.INIT('h5553)
	) name3856 (
		\Datai[2]_pad ,
		\InstQueue_reg[8][2]/NET0131 ,
		_w2232_,
		_w2234_,
		_w4309_
	);
	LUT2 #(
		.INIT('h1)
	) name3857 (
		_w2404_,
		_w4309_,
		_w4310_
	);
	LUT4 #(
		.INIT('h0057)
	) name3858 (
		\DataWidth_reg[1]/NET0131 ,
		_w4307_,
		_w4308_,
		_w4310_,
		_w4311_
	);
	LUT4 #(
		.INIT('hc055)
	) name3859 (
		\InstQueue_reg[8][2]/NET0131 ,
		_w466_,
		_w479_,
		_w2234_,
		_w4312_
	);
	LUT2 #(
		.INIT('h2)
	) name3860 (
		\InstQueue_reg[8][2]/NET0131 ,
		_w2227_,
		_w4313_
	);
	LUT3 #(
		.INIT('h0d)
	) name3861 (
		_w1212_,
		_w4309_,
		_w4313_,
		_w4314_
	);
	LUT3 #(
		.INIT('hd0)
	) name3862 (
		_w710_,
		_w4312_,
		_w4314_,
		_w4315_
	);
	LUT3 #(
		.INIT('h2f)
	) name3863 (
		_w695_,
		_w4311_,
		_w4315_,
		_w4316_
	);
	LUT4 #(
		.INIT('h6c00)
	) name3864 (
		\Datai[25]_pad ,
		\Datai[26]_pad ,
		_w2208_,
		_w2378_,
		_w4317_
	);
	LUT3 #(
		.INIT('h60)
	) name3865 (
		\Datai[18]_pad ,
		_w2211_,
		_w2232_,
		_w4318_
	);
	LUT4 #(
		.INIT('h5553)
	) name3866 (
		\Datai[2]_pad ,
		\InstQueue_reg[9][2]/NET0131 ,
		_w2237_,
		_w2234_,
		_w4319_
	);
	LUT2 #(
		.INIT('h1)
	) name3867 (
		_w2415_,
		_w4319_,
		_w4320_
	);
	LUT4 #(
		.INIT('h0057)
	) name3868 (
		\DataWidth_reg[1]/NET0131 ,
		_w4317_,
		_w4318_,
		_w4320_,
		_w4321_
	);
	LUT4 #(
		.INIT('hc055)
	) name3869 (
		\InstQueue_reg[9][2]/NET0131 ,
		_w466_,
		_w479_,
		_w2237_,
		_w4322_
	);
	LUT2 #(
		.INIT('h2)
	) name3870 (
		\InstQueue_reg[9][2]/NET0131 ,
		_w2227_,
		_w4323_
	);
	LUT3 #(
		.INIT('h0d)
	) name3871 (
		_w1212_,
		_w4319_,
		_w4323_,
		_w4324_
	);
	LUT3 #(
		.INIT('hd0)
	) name3872 (
		_w710_,
		_w4322_,
		_w4324_,
		_w4325_
	);
	LUT3 #(
		.INIT('h2f)
	) name3873 (
		_w695_,
		_w4321_,
		_w4325_,
		_w4326_
	);
	LUT3 #(
		.INIT('h10)
	) name3874 (
		_w594_,
		_w4021_,
		_w4022_,
		_w4327_
	);
	LUT2 #(
		.INIT('h2)
	) name3875 (
		\Datao[29]_pad ,
		_w596_,
		_w4328_
	);
	LUT4 #(
		.INIT('h3f15)
	) name3876 (
		\Datao[29]_pad ,
		\uWord_reg[13]/NET0131 ,
		_w2179_,
		_w2180_,
		_w4329_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name3877 (
		_w690_,
		_w4327_,
		_w4328_,
		_w4329_,
		_w4330_
	);
	LUT2 #(
		.INIT('h8)
	) name3878 (
		\CodeFetch_reg/NET0131 ,
		_w690_,
		_w4331_
	);
	LUT3 #(
		.INIT('h31)
	) name3879 (
		\CodeFetch_reg/NET0131 ,
		_w696_,
		_w1841_,
		_w4332_
	);
	LUT3 #(
		.INIT('h4f)
	) name3880 (
		_w3110_,
		_w4331_,
		_w4332_,
		_w4333_
	);
	LUT4 #(
		.INIT('h0200)
	) name3881 (
		_w589_,
		_w594_,
		_w566_,
		_w4043_,
		_w4334_
	);
	LUT4 #(
		.INIT('hf020)
	) name3882 (
		\Datao[18]_pad ,
		_w596_,
		_w690_,
		_w4334_,
		_w4335_
	);
	LUT4 #(
		.INIT('h3f15)
	) name3883 (
		\Datao[18]_pad ,
		\uWord_reg[2]/NET0131 ,
		_w2179_,
		_w2180_,
		_w4336_
	);
	LUT2 #(
		.INIT('hb)
	) name3884 (
		_w4335_,
		_w4336_,
		_w4337_
	);
	LUT2 #(
		.INIT('h1)
	) name3885 (
		_w594_,
		_w4058_,
		_w4338_
	);
	LUT3 #(
		.INIT('h02)
	) name3886 (
		_w589_,
		_w566_,
		_w4338_,
		_w4339_
	);
	LUT4 #(
		.INIT('haaa2)
	) name3887 (
		\Datao[22]_pad ,
		_w646_,
		_w2183_,
		_w4339_,
		_w4340_
	);
	LUT3 #(
		.INIT('h80)
	) name3888 (
		_w589_,
		_w595_,
		_w4058_,
		_w4341_
	);
	LUT4 #(
		.INIT('h3f15)
	) name3889 (
		\Datao[22]_pad ,
		\uWord_reg[6]/NET0131 ,
		_w2179_,
		_w2180_,
		_w4342_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name3890 (
		_w690_,
		_w4340_,
		_w4341_,
		_w4342_,
		_w4343_
	);
	LUT4 #(
		.INIT('hccc4)
	) name3891 (
		_w690_,
		_w1841_,
		_w1990_,
		_w1991_,
		_w4344_
	);
	LUT4 #(
		.INIT('h8000)
	) name3892 (
		\InstQueue_reg[0][0]/NET0131 ,
		_w569_,
		_w602_,
		_w634_,
		_w4345_
	);
	LUT3 #(
		.INIT('h40)
	) name3893 (
		\EBX_reg[0]/NET0131 ,
		_w617_,
		_w621_,
		_w4346_
	);
	LUT3 #(
		.INIT('ha8)
	) name3894 (
		_w690_,
		_w4345_,
		_w4346_,
		_w4347_
	);
	LUT3 #(
		.INIT('hf2)
	) name3895 (
		\EBX_reg[0]/NET0131 ,
		_w4344_,
		_w4347_,
		_w4348_
	);
	LUT3 #(
		.INIT('h01)
	) name3896 (
		\InstQueue_reg[0][1]/NET0131 ,
		_w563_,
		_w633_,
		_w4349_
	);
	LUT3 #(
		.INIT('h54)
	) name3897 (
		\EBX_reg[1]/NET0131 ,
		_w563_,
		_w633_,
		_w4350_
	);
	LUT4 #(
		.INIT('h0008)
	) name3898 (
		_w569_,
		_w602_,
		_w4350_,
		_w4349_,
		_w4351_
	);
	LUT3 #(
		.INIT('h2a)
	) name3899 (
		\EBX_reg[1]/NET0131 ,
		_w569_,
		_w602_,
		_w4352_
	);
	LUT4 #(
		.INIT('h0027)
	) name3900 (
		_w622_,
		_w3114_,
		_w4352_,
		_w4351_,
		_w4353_
	);
	LUT2 #(
		.INIT('h2)
	) name3901 (
		\EBX_reg[1]/NET0131 ,
		_w1841_,
		_w4354_
	);
	LUT3 #(
		.INIT('hf2)
	) name3902 (
		_w690_,
		_w4353_,
		_w4354_,
		_w4355_
	);
	LUT3 #(
		.INIT('h02)
	) name3903 (
		\EBX_reg[2]/NET0131 ,
		_w1990_,
		_w1991_,
		_w4356_
	);
	LUT4 #(
		.INIT('h8000)
	) name3904 (
		\InstQueue_reg[0][2]/NET0131 ,
		_w569_,
		_w602_,
		_w634_,
		_w4357_
	);
	LUT3 #(
		.INIT('h78)
	) name3905 (
		\EBX_reg[0]/NET0131 ,
		\EBX_reg[1]/NET0131 ,
		\EBX_reg[2]/NET0131 ,
		_w4358_
	);
	LUT3 #(
		.INIT('h80)
	) name3906 (
		_w617_,
		_w621_,
		_w4358_,
		_w4359_
	);
	LUT2 #(
		.INIT('h1)
	) name3907 (
		_w4357_,
		_w4359_,
		_w4360_
	);
	LUT2 #(
		.INIT('h2)
	) name3908 (
		\EBX_reg[2]/NET0131 ,
		_w1841_,
		_w4361_
	);
	LUT4 #(
		.INIT('hff8a)
	) name3909 (
		_w690_,
		_w4356_,
		_w4360_,
		_w4361_,
		_w4362_
	);
	LUT3 #(
		.INIT('h02)
	) name3910 (
		\EBX_reg[3]/NET0131 ,
		_w1990_,
		_w1991_,
		_w4363_
	);
	LUT4 #(
		.INIT('h8000)
	) name3911 (
		\InstQueue_reg[0][3]/NET0131 ,
		_w569_,
		_w602_,
		_w634_,
		_w4364_
	);
	LUT4 #(
		.INIT('h7f80)
	) name3912 (
		\EBX_reg[0]/NET0131 ,
		\EBX_reg[1]/NET0131 ,
		\EBX_reg[2]/NET0131 ,
		\EBX_reg[3]/NET0131 ,
		_w4365_
	);
	LUT3 #(
		.INIT('h80)
	) name3913 (
		_w617_,
		_w621_,
		_w4365_,
		_w4366_
	);
	LUT2 #(
		.INIT('h1)
	) name3914 (
		_w4364_,
		_w4366_,
		_w4367_
	);
	LUT2 #(
		.INIT('h2)
	) name3915 (
		\EBX_reg[3]/NET0131 ,
		_w1841_,
		_w4368_
	);
	LUT4 #(
		.INIT('hff8a)
	) name3916 (
		_w690_,
		_w4363_,
		_w4367_,
		_w4368_,
		_w4369_
	);
	LUT3 #(
		.INIT('h02)
	) name3917 (
		\EBX_reg[4]/NET0131 ,
		_w1990_,
		_w1991_,
		_w4370_
	);
	LUT4 #(
		.INIT('h8000)
	) name3918 (
		\InstQueue_reg[0][4]/NET0131 ,
		_w569_,
		_w602_,
		_w634_,
		_w4371_
	);
	LUT2 #(
		.INIT('h6)
	) name3919 (
		\EBX_reg[4]/NET0131 ,
		_w1971_,
		_w4372_
	);
	LUT3 #(
		.INIT('h80)
	) name3920 (
		_w617_,
		_w621_,
		_w4372_,
		_w4373_
	);
	LUT2 #(
		.INIT('h1)
	) name3921 (
		_w4371_,
		_w4373_,
		_w4374_
	);
	LUT2 #(
		.INIT('h2)
	) name3922 (
		\EBX_reg[4]/NET0131 ,
		_w1841_,
		_w4375_
	);
	LUT4 #(
		.INIT('hff8a)
	) name3923 (
		_w690_,
		_w4370_,
		_w4374_,
		_w4375_,
		_w4376_
	);
	LUT3 #(
		.INIT('h02)
	) name3924 (
		\EBX_reg[5]/NET0131 ,
		_w1990_,
		_w1991_,
		_w4377_
	);
	LUT4 #(
		.INIT('h8000)
	) name3925 (
		\InstQueue_reg[0][5]/NET0131 ,
		_w569_,
		_w602_,
		_w634_,
		_w4378_
	);
	LUT3 #(
		.INIT('h6c)
	) name3926 (
		\EBX_reg[4]/NET0131 ,
		\EBX_reg[5]/NET0131 ,
		_w1971_,
		_w4379_
	);
	LUT3 #(
		.INIT('h80)
	) name3927 (
		_w617_,
		_w621_,
		_w4379_,
		_w4380_
	);
	LUT2 #(
		.INIT('h1)
	) name3928 (
		_w4378_,
		_w4380_,
		_w4381_
	);
	LUT2 #(
		.INIT('h2)
	) name3929 (
		\EBX_reg[5]/NET0131 ,
		_w1841_,
		_w4382_
	);
	LUT4 #(
		.INIT('hff8a)
	) name3930 (
		_w690_,
		_w4377_,
		_w4381_,
		_w4382_,
		_w4383_
	);
	LUT3 #(
		.INIT('h02)
	) name3931 (
		\EBX_reg[6]/NET0131 ,
		_w1990_,
		_w1991_,
		_w4384_
	);
	LUT4 #(
		.INIT('h8000)
	) name3932 (
		\InstQueue_reg[0][6]/NET0131 ,
		_w569_,
		_w602_,
		_w634_,
		_w4385_
	);
	LUT4 #(
		.INIT('h78f0)
	) name3933 (
		\EBX_reg[4]/NET0131 ,
		\EBX_reg[5]/NET0131 ,
		\EBX_reg[6]/NET0131 ,
		_w1971_,
		_w4386_
	);
	LUT3 #(
		.INIT('h80)
	) name3934 (
		_w617_,
		_w621_,
		_w4386_,
		_w4387_
	);
	LUT2 #(
		.INIT('h1)
	) name3935 (
		_w4385_,
		_w4387_,
		_w4388_
	);
	LUT2 #(
		.INIT('h2)
	) name3936 (
		\EBX_reg[6]/NET0131 ,
		_w1841_,
		_w4389_
	);
	LUT4 #(
		.INIT('hff8a)
	) name3937 (
		_w690_,
		_w4384_,
		_w4388_,
		_w4389_,
		_w4390_
	);
	LUT3 #(
		.INIT('h02)
	) name3938 (
		\EBX_reg[7]/NET0131 ,
		_w1990_,
		_w1991_,
		_w4391_
	);
	LUT4 #(
		.INIT('h8000)
	) name3939 (
		\InstQueue_reg[0][7]/NET0131 ,
		_w569_,
		_w602_,
		_w634_,
		_w4392_
	);
	LUT2 #(
		.INIT('h6)
	) name3940 (
		\EBX_reg[7]/NET0131 ,
		_w1972_,
		_w4393_
	);
	LUT3 #(
		.INIT('h80)
	) name3941 (
		_w617_,
		_w621_,
		_w4393_,
		_w4394_
	);
	LUT2 #(
		.INIT('h1)
	) name3942 (
		_w4392_,
		_w4394_,
		_w4395_
	);
	LUT2 #(
		.INIT('h2)
	) name3943 (
		\EBX_reg[7]/NET0131 ,
		_w1841_,
		_w4396_
	);
	LUT4 #(
		.INIT('hff8a)
	) name3944 (
		_w690_,
		_w4391_,
		_w4395_,
		_w4396_,
		_w4397_
	);
	LUT2 #(
		.INIT('h8)
	) name3945 (
		READY_n_pad,
		\lWord_reg[0]/NET0131 ,
		_w4398_
	);
	LUT2 #(
		.INIT('h1)
	) name3946 (
		_w3824_,
		_w4398_,
		_w4399_
	);
	LUT2 #(
		.INIT('h2)
	) name3947 (
		_w582_,
		_w4399_,
		_w4400_
	);
	LUT4 #(
		.INIT('haa02)
	) name3948 (
		\lWord_reg[0]/NET0131 ,
		_w582_,
		_w589_,
		_w566_,
		_w4401_
	);
	LUT3 #(
		.INIT('h08)
	) name3949 (
		\EAX_reg[0]/NET0131 ,
		_w589_,
		_w566_,
		_w4402_
	);
	LUT4 #(
		.INIT('haaa8)
	) name3950 (
		_w690_,
		_w4401_,
		_w4400_,
		_w4402_,
		_w4403_
	);
	LUT2 #(
		.INIT('h2)
	) name3951 (
		\lWord_reg[0]/NET0131 ,
		_w1841_,
		_w4404_
	);
	LUT2 #(
		.INIT('he)
	) name3952 (
		_w4403_,
		_w4404_,
		_w4405_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name3953 (
		\lWord_reg[10]/NET0131 ,
		_w690_,
		_w1841_,
		_w2103_,
		_w4406_
	);
	LUT3 #(
		.INIT('h08)
	) name3954 (
		\EAX_reg[10]/NET0131 ,
		_w589_,
		_w566_,
		_w4407_
	);
	LUT3 #(
		.INIT('h20)
	) name3955 (
		_w582_,
		_w566_,
		_w4016_,
		_w4408_
	);
	LUT3 #(
		.INIT('ha8)
	) name3956 (
		_w690_,
		_w4407_,
		_w4408_,
		_w4409_
	);
	LUT2 #(
		.INIT('he)
	) name3957 (
		_w4406_,
		_w4409_,
		_w4410_
	);
	LUT2 #(
		.INIT('h8)
	) name3958 (
		READY_n_pad,
		\lWord_reg[11]/NET0131 ,
		_w4411_
	);
	LUT2 #(
		.INIT('h1)
	) name3959 (
		_w1834_,
		_w4411_,
		_w4412_
	);
	LUT2 #(
		.INIT('h2)
	) name3960 (
		_w582_,
		_w4412_,
		_w4413_
	);
	LUT4 #(
		.INIT('haa02)
	) name3961 (
		\lWord_reg[11]/NET0131 ,
		_w582_,
		_w589_,
		_w566_,
		_w4414_
	);
	LUT3 #(
		.INIT('h08)
	) name3962 (
		\EAX_reg[11]/NET0131 ,
		_w589_,
		_w566_,
		_w4415_
	);
	LUT4 #(
		.INIT('haaa8)
	) name3963 (
		_w690_,
		_w4414_,
		_w4413_,
		_w4415_,
		_w4416_
	);
	LUT2 #(
		.INIT('h2)
	) name3964 (
		\lWord_reg[11]/NET0131 ,
		_w1841_,
		_w4417_
	);
	LUT2 #(
		.INIT('he)
	) name3965 (
		_w4416_,
		_w4417_,
		_w4418_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name3966 (
		\lWord_reg[12]/NET0131 ,
		_w690_,
		_w1841_,
		_w2103_,
		_w4419_
	);
	LUT3 #(
		.INIT('h08)
	) name3967 (
		\EAX_reg[12]/NET0131 ,
		_w589_,
		_w566_,
		_w4420_
	);
	LUT3 #(
		.INIT('ha8)
	) name3968 (
		_w690_,
		_w2100_,
		_w4420_,
		_w4421_
	);
	LUT2 #(
		.INIT('he)
	) name3969 (
		_w4419_,
		_w4421_,
		_w4422_
	);
	LUT2 #(
		.INIT('h8)
	) name3970 (
		READY_n_pad,
		\lWord_reg[13]/NET0131 ,
		_w4423_
	);
	LUT2 #(
		.INIT('h1)
	) name3971 (
		_w2161_,
		_w4423_,
		_w4424_
	);
	LUT2 #(
		.INIT('h2)
	) name3972 (
		_w582_,
		_w4424_,
		_w4425_
	);
	LUT4 #(
		.INIT('haa02)
	) name3973 (
		\lWord_reg[13]/NET0131 ,
		_w582_,
		_w589_,
		_w566_,
		_w4426_
	);
	LUT3 #(
		.INIT('h08)
	) name3974 (
		\EAX_reg[13]/NET0131 ,
		_w589_,
		_w566_,
		_w4427_
	);
	LUT4 #(
		.INIT('haaa8)
	) name3975 (
		_w690_,
		_w4426_,
		_w4425_,
		_w4427_,
		_w4428_
	);
	LUT2 #(
		.INIT('h2)
	) name3976 (
		\lWord_reg[13]/NET0131 ,
		_w1841_,
		_w4429_
	);
	LUT2 #(
		.INIT('he)
	) name3977 (
		_w4428_,
		_w4429_,
		_w4430_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name3978 (
		\lWord_reg[14]/NET0131 ,
		_w690_,
		_w1841_,
		_w2103_,
		_w4431_
	);
	LUT3 #(
		.INIT('h08)
	) name3979 (
		\EAX_reg[14]/NET0131 ,
		_w589_,
		_w566_,
		_w4432_
	);
	LUT3 #(
		.INIT('ha8)
	) name3980 (
		_w690_,
		_w3795_,
		_w4432_,
		_w4433_
	);
	LUT2 #(
		.INIT('he)
	) name3981 (
		_w4431_,
		_w4433_,
		_w4434_
	);
	LUT2 #(
		.INIT('h8)
	) name3982 (
		READY_n_pad,
		\lWord_reg[15]/NET0131 ,
		_w4435_
	);
	LUT2 #(
		.INIT('h1)
	) name3983 (
		_w2795_,
		_w4435_,
		_w4436_
	);
	LUT2 #(
		.INIT('h2)
	) name3984 (
		_w582_,
		_w4436_,
		_w4437_
	);
	LUT4 #(
		.INIT('haa02)
	) name3985 (
		\lWord_reg[15]/NET0131 ,
		_w582_,
		_w589_,
		_w566_,
		_w4438_
	);
	LUT3 #(
		.INIT('h08)
	) name3986 (
		\EAX_reg[15]/NET0131 ,
		_w589_,
		_w566_,
		_w4439_
	);
	LUT4 #(
		.INIT('haaa8)
	) name3987 (
		_w690_,
		_w4438_,
		_w4437_,
		_w4439_,
		_w4440_
	);
	LUT2 #(
		.INIT('h2)
	) name3988 (
		\lWord_reg[15]/NET0131 ,
		_w1841_,
		_w4441_
	);
	LUT2 #(
		.INIT('he)
	) name3989 (
		_w4440_,
		_w4441_,
		_w4442_
	);
	LUT2 #(
		.INIT('h8)
	) name3990 (
		READY_n_pad,
		\lWord_reg[1]/NET0131 ,
		_w4443_
	);
	LUT2 #(
		.INIT('h1)
	) name3991 (
		_w3752_,
		_w4443_,
		_w4444_
	);
	LUT2 #(
		.INIT('h2)
	) name3992 (
		_w582_,
		_w4444_,
		_w4445_
	);
	LUT4 #(
		.INIT('haa02)
	) name3993 (
		\lWord_reg[1]/NET0131 ,
		_w582_,
		_w589_,
		_w566_,
		_w4446_
	);
	LUT3 #(
		.INIT('h08)
	) name3994 (
		\EAX_reg[1]/NET0131 ,
		_w589_,
		_w566_,
		_w4447_
	);
	LUT4 #(
		.INIT('haaa8)
	) name3995 (
		_w690_,
		_w4446_,
		_w4445_,
		_w4447_,
		_w4448_
	);
	LUT2 #(
		.INIT('h2)
	) name3996 (
		\lWord_reg[1]/NET0131 ,
		_w1841_,
		_w4449_
	);
	LUT2 #(
		.INIT('he)
	) name3997 (
		_w4448_,
		_w4449_,
		_w4450_
	);
	LUT2 #(
		.INIT('h8)
	) name3998 (
		READY_n_pad,
		\lWord_reg[2]/NET0131 ,
		_w4451_
	);
	LUT2 #(
		.INIT('h1)
	) name3999 (
		_w3700_,
		_w4451_,
		_w4452_
	);
	LUT2 #(
		.INIT('h2)
	) name4000 (
		_w582_,
		_w4452_,
		_w4453_
	);
	LUT4 #(
		.INIT('haa02)
	) name4001 (
		\lWord_reg[2]/NET0131 ,
		_w582_,
		_w589_,
		_w566_,
		_w4454_
	);
	LUT3 #(
		.INIT('h08)
	) name4002 (
		\EAX_reg[2]/NET0131 ,
		_w589_,
		_w566_,
		_w4455_
	);
	LUT4 #(
		.INIT('haaa8)
	) name4003 (
		_w690_,
		_w4454_,
		_w4453_,
		_w4455_,
		_w4456_
	);
	LUT2 #(
		.INIT('h2)
	) name4004 (
		\lWord_reg[2]/NET0131 ,
		_w1841_,
		_w4457_
	);
	LUT2 #(
		.INIT('he)
	) name4005 (
		_w4456_,
		_w4457_,
		_w4458_
	);
	LUT2 #(
		.INIT('h8)
	) name4006 (
		READY_n_pad,
		\lWord_reg[3]/NET0131 ,
		_w4459_
	);
	LUT2 #(
		.INIT('h1)
	) name4007 (
		_w3708_,
		_w4459_,
		_w4460_
	);
	LUT2 #(
		.INIT('h2)
	) name4008 (
		_w582_,
		_w4460_,
		_w4461_
	);
	LUT4 #(
		.INIT('haa02)
	) name4009 (
		\lWord_reg[3]/NET0131 ,
		_w582_,
		_w589_,
		_w566_,
		_w4462_
	);
	LUT3 #(
		.INIT('h08)
	) name4010 (
		\EAX_reg[3]/NET0131 ,
		_w589_,
		_w566_,
		_w4463_
	);
	LUT4 #(
		.INIT('haaa8)
	) name4011 (
		_w690_,
		_w4462_,
		_w4461_,
		_w4463_,
		_w4464_
	);
	LUT2 #(
		.INIT('h2)
	) name4012 (
		\lWord_reg[3]/NET0131 ,
		_w1841_,
		_w4465_
	);
	LUT2 #(
		.INIT('he)
	) name4013 (
		_w4464_,
		_w4465_,
		_w4466_
	);
	LUT2 #(
		.INIT('h8)
	) name4014 (
		READY_n_pad,
		\lWord_reg[4]/NET0131 ,
		_w4467_
	);
	LUT2 #(
		.INIT('h1)
	) name4015 (
		_w2442_,
		_w4467_,
		_w4468_
	);
	LUT2 #(
		.INIT('h2)
	) name4016 (
		_w582_,
		_w4468_,
		_w4469_
	);
	LUT4 #(
		.INIT('haa02)
	) name4017 (
		\lWord_reg[4]/NET0131 ,
		_w582_,
		_w589_,
		_w566_,
		_w4470_
	);
	LUT3 #(
		.INIT('h08)
	) name4018 (
		\EAX_reg[4]/NET0131 ,
		_w589_,
		_w566_,
		_w4471_
	);
	LUT4 #(
		.INIT('haaa8)
	) name4019 (
		_w690_,
		_w4470_,
		_w4469_,
		_w4471_,
		_w4472_
	);
	LUT2 #(
		.INIT('h2)
	) name4020 (
		\lWord_reg[4]/NET0131 ,
		_w1841_,
		_w4473_
	);
	LUT2 #(
		.INIT('he)
	) name4021 (
		_w4472_,
		_w4473_,
		_w4474_
	);
	LUT2 #(
		.INIT('h8)
	) name4022 (
		READY_n_pad,
		\lWord_reg[5]/NET0131 ,
		_w4475_
	);
	LUT2 #(
		.INIT('h1)
	) name4023 (
		_w3734_,
		_w4475_,
		_w4476_
	);
	LUT2 #(
		.INIT('h2)
	) name4024 (
		_w582_,
		_w4476_,
		_w4477_
	);
	LUT4 #(
		.INIT('haa02)
	) name4025 (
		\lWord_reg[5]/NET0131 ,
		_w582_,
		_w589_,
		_w566_,
		_w4478_
	);
	LUT3 #(
		.INIT('h08)
	) name4026 (
		\EAX_reg[5]/NET0131 ,
		_w589_,
		_w566_,
		_w4479_
	);
	LUT4 #(
		.INIT('haaa8)
	) name4027 (
		_w690_,
		_w4478_,
		_w4477_,
		_w4479_,
		_w4480_
	);
	LUT2 #(
		.INIT('h2)
	) name4028 (
		\lWord_reg[5]/NET0131 ,
		_w1841_,
		_w4481_
	);
	LUT2 #(
		.INIT('he)
	) name4029 (
		_w4480_,
		_w4481_,
		_w4482_
	);
	LUT4 #(
		.INIT('h2202)
	) name4030 (
		\Datai[6]_pad ,
		READY_n_pad,
		_w563_,
		_w565_,
		_w4483_
	);
	LUT2 #(
		.INIT('h8)
	) name4031 (
		READY_n_pad,
		\lWord_reg[6]/NET0131 ,
		_w4484_
	);
	LUT2 #(
		.INIT('h1)
	) name4032 (
		_w4483_,
		_w4484_,
		_w4485_
	);
	LUT2 #(
		.INIT('h2)
	) name4033 (
		_w582_,
		_w4485_,
		_w4486_
	);
	LUT4 #(
		.INIT('haa02)
	) name4034 (
		\lWord_reg[6]/NET0131 ,
		_w582_,
		_w589_,
		_w566_,
		_w4487_
	);
	LUT3 #(
		.INIT('h08)
	) name4035 (
		\EAX_reg[6]/NET0131 ,
		_w589_,
		_w566_,
		_w4488_
	);
	LUT4 #(
		.INIT('haaa8)
	) name4036 (
		_w690_,
		_w4487_,
		_w4486_,
		_w4488_,
		_w4489_
	);
	LUT2 #(
		.INIT('h2)
	) name4037 (
		\lWord_reg[6]/NET0131 ,
		_w1841_,
		_w4490_
	);
	LUT2 #(
		.INIT('he)
	) name4038 (
		_w4489_,
		_w4490_,
		_w4491_
	);
	LUT2 #(
		.INIT('h8)
	) name4039 (
		READY_n_pad,
		\lWord_reg[7]/NET0131 ,
		_w4492_
	);
	LUT2 #(
		.INIT('h1)
	) name4040 (
		_w2644_,
		_w4492_,
		_w4493_
	);
	LUT2 #(
		.INIT('h2)
	) name4041 (
		_w582_,
		_w4493_,
		_w4494_
	);
	LUT4 #(
		.INIT('haa02)
	) name4042 (
		\lWord_reg[7]/NET0131 ,
		_w582_,
		_w589_,
		_w566_,
		_w4495_
	);
	LUT3 #(
		.INIT('h08)
	) name4043 (
		\EAX_reg[7]/NET0131 ,
		_w589_,
		_w566_,
		_w4496_
	);
	LUT4 #(
		.INIT('haaa8)
	) name4044 (
		_w690_,
		_w4495_,
		_w4494_,
		_w4496_,
		_w4497_
	);
	LUT2 #(
		.INIT('h2)
	) name4045 (
		\lWord_reg[7]/NET0131 ,
		_w1841_,
		_w4498_
	);
	LUT2 #(
		.INIT('he)
	) name4046 (
		_w4497_,
		_w4498_,
		_w4499_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name4047 (
		\lWord_reg[8]/NET0131 ,
		_w690_,
		_w1841_,
		_w2103_,
		_w4500_
	);
	LUT3 #(
		.INIT('h08)
	) name4048 (
		\EAX_reg[8]/NET0131 ,
		_w589_,
		_w566_,
		_w4501_
	);
	LUT3 #(
		.INIT('h20)
	) name4049 (
		_w582_,
		_w566_,
		_w2190_,
		_w4502_
	);
	LUT3 #(
		.INIT('ha8)
	) name4050 (
		_w690_,
		_w4501_,
		_w4502_,
		_w4503_
	);
	LUT2 #(
		.INIT('he)
	) name4051 (
		_w4500_,
		_w4503_,
		_w4504_
	);
	LUT2 #(
		.INIT('h8)
	) name4052 (
		READY_n_pad,
		\lWord_reg[9]/NET0131 ,
		_w4505_
	);
	LUT2 #(
		.INIT('h1)
	) name4053 (
		_w2455_,
		_w4505_,
		_w4506_
	);
	LUT2 #(
		.INIT('h2)
	) name4054 (
		_w582_,
		_w4506_,
		_w4507_
	);
	LUT4 #(
		.INIT('haa02)
	) name4055 (
		\lWord_reg[9]/NET0131 ,
		_w582_,
		_w589_,
		_w566_,
		_w4508_
	);
	LUT3 #(
		.INIT('h08)
	) name4056 (
		\EAX_reg[9]/NET0131 ,
		_w589_,
		_w566_,
		_w4509_
	);
	LUT4 #(
		.INIT('haaa8)
	) name4057 (
		_w690_,
		_w4508_,
		_w4507_,
		_w4509_,
		_w4510_
	);
	LUT2 #(
		.INIT('h2)
	) name4058 (
		\lWord_reg[9]/NET0131 ,
		_w1841_,
		_w4511_
	);
	LUT2 #(
		.INIT('he)
	) name4059 (
		_w4510_,
		_w4511_,
		_w4512_
	);
	LUT4 #(
		.INIT('h60c0)
	) name4060 (
		\Datai[28]_pad ,
		\Datai[29]_pad ,
		_w2199_,
		_w2209_,
		_w4513_
	);
	LUT3 #(
		.INIT('h60)
	) name4061 (
		\Datai[21]_pad ,
		_w2212_,
		_w2215_,
		_w4514_
	);
	LUT4 #(
		.INIT('h5553)
	) name4062 (
		\Datai[5]_pad ,
		\InstQueue_reg[0][5]/NET0131 ,
		_w2217_,
		_w2219_,
		_w4515_
	);
	LUT2 #(
		.INIT('h1)
	) name4063 (
		_w2223_,
		_w4515_,
		_w4516_
	);
	LUT4 #(
		.INIT('h0057)
	) name4064 (
		\DataWidth_reg[1]/NET0131 ,
		_w4513_,
		_w4514_,
		_w4516_,
		_w4517_
	);
	LUT4 #(
		.INIT('hc055)
	) name4065 (
		\InstQueue_reg[0][5]/NET0131 ,
		_w534_,
		_w539_,
		_w2217_,
		_w4518_
	);
	LUT2 #(
		.INIT('h2)
	) name4066 (
		\InstQueue_reg[0][5]/NET0131 ,
		_w2227_,
		_w4519_
	);
	LUT3 #(
		.INIT('h0d)
	) name4067 (
		_w1212_,
		_w4515_,
		_w4519_,
		_w4520_
	);
	LUT3 #(
		.INIT('hd0)
	) name4068 (
		_w710_,
		_w4518_,
		_w4520_,
		_w4521_
	);
	LUT3 #(
		.INIT('h2f)
	) name4069 (
		_w695_,
		_w4517_,
		_w4521_,
		_w4522_
	);
	LUT4 #(
		.INIT('h6c00)
	) name4070 (
		\Datai[28]_pad ,
		\Datai[29]_pad ,
		_w2209_,
		_w2232_,
		_w4523_
	);
	LUT3 #(
		.INIT('h60)
	) name4071 (
		\Datai[21]_pad ,
		_w2212_,
		_w2234_,
		_w4524_
	);
	LUT4 #(
		.INIT('h5553)
	) name4072 (
		\Datai[5]_pad ,
		\InstQueue_reg[10][5]/NET0131 ,
		_w2236_,
		_w2237_,
		_w4525_
	);
	LUT2 #(
		.INIT('h1)
	) name4073 (
		_w2241_,
		_w4525_,
		_w4526_
	);
	LUT4 #(
		.INIT('h0057)
	) name4074 (
		\DataWidth_reg[1]/NET0131 ,
		_w4523_,
		_w4524_,
		_w4526_,
		_w4527_
	);
	LUT4 #(
		.INIT('hc055)
	) name4075 (
		\InstQueue_reg[10][5]/NET0131 ,
		_w534_,
		_w539_,
		_w2236_,
		_w4528_
	);
	LUT2 #(
		.INIT('h2)
	) name4076 (
		\InstQueue_reg[10][5]/NET0131 ,
		_w2227_,
		_w4529_
	);
	LUT3 #(
		.INIT('h0d)
	) name4077 (
		_w1212_,
		_w4525_,
		_w4529_,
		_w4530_
	);
	LUT3 #(
		.INIT('hd0)
	) name4078 (
		_w710_,
		_w4528_,
		_w4530_,
		_w4531_
	);
	LUT3 #(
		.INIT('h2f)
	) name4079 (
		_w695_,
		_w4527_,
		_w4531_,
		_w4532_
	);
	LUT4 #(
		.INIT('h6c00)
	) name4080 (
		\Datai[28]_pad ,
		\Datai[29]_pad ,
		_w2209_,
		_w2234_,
		_w4533_
	);
	LUT3 #(
		.INIT('h60)
	) name4081 (
		\Datai[21]_pad ,
		_w2212_,
		_w2237_,
		_w4534_
	);
	LUT4 #(
		.INIT('h5553)
	) name4082 (
		\Datai[5]_pad ,
		\InstQueue_reg[11][5]/NET0131 ,
		_w2236_,
		_w2251_,
		_w4535_
	);
	LUT2 #(
		.INIT('h1)
	) name4083 (
		_w2255_,
		_w4535_,
		_w4536_
	);
	LUT4 #(
		.INIT('h0057)
	) name4084 (
		\DataWidth_reg[1]/NET0131 ,
		_w4533_,
		_w4534_,
		_w4536_,
		_w4537_
	);
	LUT4 #(
		.INIT('hc055)
	) name4085 (
		\InstQueue_reg[11][5]/NET0131 ,
		_w534_,
		_w539_,
		_w2251_,
		_w4538_
	);
	LUT2 #(
		.INIT('h2)
	) name4086 (
		\InstQueue_reg[11][5]/NET0131 ,
		_w2227_,
		_w4539_
	);
	LUT3 #(
		.INIT('h0d)
	) name4087 (
		_w1212_,
		_w4535_,
		_w4539_,
		_w4540_
	);
	LUT3 #(
		.INIT('hd0)
	) name4088 (
		_w710_,
		_w4538_,
		_w4540_,
		_w4541_
	);
	LUT3 #(
		.INIT('h2f)
	) name4089 (
		_w695_,
		_w4537_,
		_w4541_,
		_w4542_
	);
	LUT4 #(
		.INIT('h6c00)
	) name4090 (
		\Datai[28]_pad ,
		\Datai[29]_pad ,
		_w2209_,
		_w2237_,
		_w4543_
	);
	LUT3 #(
		.INIT('h60)
	) name4091 (
		\Datai[21]_pad ,
		_w2212_,
		_w2236_,
		_w4544_
	);
	LUT4 #(
		.INIT('h5553)
	) name4092 (
		\Datai[5]_pad ,
		\InstQueue_reg[12][5]/NET0131 ,
		_w2251_,
		_w2265_,
		_w4545_
	);
	LUT2 #(
		.INIT('h1)
	) name4093 (
		_w2268_,
		_w4545_,
		_w4546_
	);
	LUT4 #(
		.INIT('h0057)
	) name4094 (
		\DataWidth_reg[1]/NET0131 ,
		_w4543_,
		_w4544_,
		_w4546_,
		_w4547_
	);
	LUT4 #(
		.INIT('hc055)
	) name4095 (
		\InstQueue_reg[12][5]/NET0131 ,
		_w534_,
		_w539_,
		_w2265_,
		_w4548_
	);
	LUT2 #(
		.INIT('h2)
	) name4096 (
		\InstQueue_reg[12][5]/NET0131 ,
		_w2227_,
		_w4549_
	);
	LUT3 #(
		.INIT('h0d)
	) name4097 (
		_w1212_,
		_w4545_,
		_w4549_,
		_w4550_
	);
	LUT3 #(
		.INIT('hd0)
	) name4098 (
		_w710_,
		_w4548_,
		_w4550_,
		_w4551_
	);
	LUT3 #(
		.INIT('h2f)
	) name4099 (
		_w695_,
		_w4547_,
		_w4551_,
		_w4552_
	);
	LUT4 #(
		.INIT('h6c00)
	) name4100 (
		\Datai[28]_pad ,
		\Datai[29]_pad ,
		_w2209_,
		_w2236_,
		_w4553_
	);
	LUT3 #(
		.INIT('h60)
	) name4101 (
		\Datai[21]_pad ,
		_w2212_,
		_w2251_,
		_w4554_
	);
	LUT4 #(
		.INIT('h5553)
	) name4102 (
		\Datai[5]_pad ,
		\InstQueue_reg[13][5]/NET0131 ,
		_w2199_,
		_w2265_,
		_w4555_
	);
	LUT2 #(
		.INIT('h1)
	) name4103 (
		_w2280_,
		_w4555_,
		_w4556_
	);
	LUT4 #(
		.INIT('h0057)
	) name4104 (
		\DataWidth_reg[1]/NET0131 ,
		_w4553_,
		_w4554_,
		_w4556_,
		_w4557_
	);
	LUT4 #(
		.INIT('hc055)
	) name4105 (
		\InstQueue_reg[13][5]/NET0131 ,
		_w534_,
		_w539_,
		_w2199_,
		_w4558_
	);
	LUT2 #(
		.INIT('h2)
	) name4106 (
		\InstQueue_reg[13][5]/NET0131 ,
		_w2227_,
		_w4559_
	);
	LUT3 #(
		.INIT('h0d)
	) name4107 (
		_w1212_,
		_w4555_,
		_w4559_,
		_w4560_
	);
	LUT3 #(
		.INIT('hd0)
	) name4108 (
		_w710_,
		_w4558_,
		_w4560_,
		_w4561_
	);
	LUT3 #(
		.INIT('h2f)
	) name4109 (
		_w695_,
		_w4557_,
		_w4561_,
		_w4562_
	);
	LUT4 #(
		.INIT('h6c00)
	) name4110 (
		\Datai[28]_pad ,
		\Datai[29]_pad ,
		_w2209_,
		_w2251_,
		_w4563_
	);
	LUT3 #(
		.INIT('h60)
	) name4111 (
		\Datai[21]_pad ,
		_w2212_,
		_w2265_,
		_w4564_
	);
	LUT4 #(
		.INIT('h5553)
	) name4112 (
		\Datai[5]_pad ,
		\InstQueue_reg[14][5]/NET0131 ,
		_w2199_,
		_w2215_,
		_w4565_
	);
	LUT2 #(
		.INIT('h1)
	) name4113 (
		_w2291_,
		_w4565_,
		_w4566_
	);
	LUT4 #(
		.INIT('h0057)
	) name4114 (
		\DataWidth_reg[1]/NET0131 ,
		_w4563_,
		_w4564_,
		_w4566_,
		_w4567_
	);
	LUT4 #(
		.INIT('hc055)
	) name4115 (
		\InstQueue_reg[14][5]/NET0131 ,
		_w534_,
		_w539_,
		_w2215_,
		_w4568_
	);
	LUT2 #(
		.INIT('h2)
	) name4116 (
		\InstQueue_reg[14][5]/NET0131 ,
		_w2227_,
		_w4569_
	);
	LUT3 #(
		.INIT('h0d)
	) name4117 (
		_w1212_,
		_w4565_,
		_w4569_,
		_w4570_
	);
	LUT3 #(
		.INIT('hd0)
	) name4118 (
		_w710_,
		_w4568_,
		_w4570_,
		_w4571_
	);
	LUT3 #(
		.INIT('h2f)
	) name4119 (
		_w695_,
		_w4567_,
		_w4571_,
		_w4572_
	);
	LUT4 #(
		.INIT('h6c00)
	) name4120 (
		\Datai[28]_pad ,
		\Datai[29]_pad ,
		_w2209_,
		_w2265_,
		_w4573_
	);
	LUT3 #(
		.INIT('h48)
	) name4121 (
		\Datai[21]_pad ,
		_w2199_,
		_w2212_,
		_w4574_
	);
	LUT4 #(
		.INIT('h5553)
	) name4122 (
		\Datai[5]_pad ,
		\InstQueue_reg[15][5]/NET0131 ,
		_w2219_,
		_w2215_,
		_w4575_
	);
	LUT2 #(
		.INIT('h1)
	) name4123 (
		_w2303_,
		_w4575_,
		_w4576_
	);
	LUT4 #(
		.INIT('h0057)
	) name4124 (
		\DataWidth_reg[1]/NET0131 ,
		_w4573_,
		_w4574_,
		_w4576_,
		_w4577_
	);
	LUT4 #(
		.INIT('hc055)
	) name4125 (
		\InstQueue_reg[15][5]/NET0131 ,
		_w534_,
		_w539_,
		_w2219_,
		_w4578_
	);
	LUT2 #(
		.INIT('h2)
	) name4126 (
		\InstQueue_reg[15][5]/NET0131 ,
		_w2227_,
		_w4579_
	);
	LUT3 #(
		.INIT('h0d)
	) name4127 (
		_w1212_,
		_w4575_,
		_w4579_,
		_w4580_
	);
	LUT3 #(
		.INIT('hd0)
	) name4128 (
		_w710_,
		_w4578_,
		_w4580_,
		_w4581_
	);
	LUT3 #(
		.INIT('h2f)
	) name4129 (
		_w695_,
		_w4577_,
		_w4581_,
		_w4582_
	);
	LUT4 #(
		.INIT('h6c00)
	) name4130 (
		\Datai[28]_pad ,
		\Datai[29]_pad ,
		_w2209_,
		_w2215_,
		_w4583_
	);
	LUT3 #(
		.INIT('h48)
	) name4131 (
		\Datai[21]_pad ,
		_w2219_,
		_w2212_,
		_w4584_
	);
	LUT4 #(
		.INIT('h5553)
	) name4132 (
		\Datai[5]_pad ,
		\InstQueue_reg[1][5]/NET0131 ,
		_w2217_,
		_w2313_,
		_w4585_
	);
	LUT2 #(
		.INIT('h1)
	) name4133 (
		_w2316_,
		_w4585_,
		_w4586_
	);
	LUT4 #(
		.INIT('h0057)
	) name4134 (
		\DataWidth_reg[1]/NET0131 ,
		_w4583_,
		_w4584_,
		_w4586_,
		_w4587_
	);
	LUT4 #(
		.INIT('hc055)
	) name4135 (
		\InstQueue_reg[1][5]/NET0131 ,
		_w534_,
		_w539_,
		_w2313_,
		_w4588_
	);
	LUT2 #(
		.INIT('h2)
	) name4136 (
		\InstQueue_reg[1][5]/NET0131 ,
		_w2227_,
		_w4589_
	);
	LUT3 #(
		.INIT('h0d)
	) name4137 (
		_w1212_,
		_w4585_,
		_w4589_,
		_w4590_
	);
	LUT3 #(
		.INIT('hd0)
	) name4138 (
		_w710_,
		_w4588_,
		_w4590_,
		_w4591_
	);
	LUT3 #(
		.INIT('h2f)
	) name4139 (
		_w695_,
		_w4587_,
		_w4591_,
		_w4592_
	);
	LUT3 #(
		.INIT('h48)
	) name4140 (
		\Datai[21]_pad ,
		_w2217_,
		_w2212_,
		_w4593_
	);
	LUT4 #(
		.INIT('h60c0)
	) name4141 (
		\Datai[28]_pad ,
		\Datai[29]_pad ,
		_w2219_,
		_w2209_,
		_w4594_
	);
	LUT4 #(
		.INIT('h5553)
	) name4142 (
		\Datai[5]_pad ,
		\InstQueue_reg[2][5]/NET0131 ,
		_w2313_,
		_w2326_,
		_w4595_
	);
	LUT2 #(
		.INIT('h1)
	) name4143 (
		_w2329_,
		_w4595_,
		_w4596_
	);
	LUT4 #(
		.INIT('h0057)
	) name4144 (
		\DataWidth_reg[1]/NET0131 ,
		_w4593_,
		_w4594_,
		_w4596_,
		_w4597_
	);
	LUT4 #(
		.INIT('hc055)
	) name4145 (
		\InstQueue_reg[2][5]/NET0131 ,
		_w534_,
		_w539_,
		_w2326_,
		_w4598_
	);
	LUT2 #(
		.INIT('h2)
	) name4146 (
		\InstQueue_reg[2][5]/NET0131 ,
		_w2227_,
		_w4599_
	);
	LUT3 #(
		.INIT('h0d)
	) name4147 (
		_w1212_,
		_w4595_,
		_w4599_,
		_w4600_
	);
	LUT3 #(
		.INIT('hd0)
	) name4148 (
		_w710_,
		_w4598_,
		_w4600_,
		_w4601_
	);
	LUT3 #(
		.INIT('h2f)
	) name4149 (
		_w695_,
		_w4597_,
		_w4601_,
		_w4602_
	);
	LUT4 #(
		.INIT('h60c0)
	) name4150 (
		\Datai[28]_pad ,
		\Datai[29]_pad ,
		_w2217_,
		_w2209_,
		_w4603_
	);
	LUT3 #(
		.INIT('h60)
	) name4151 (
		\Datai[21]_pad ,
		_w2212_,
		_w2313_,
		_w4604_
	);
	LUT4 #(
		.INIT('h5553)
	) name4152 (
		\Datai[5]_pad ,
		\InstQueue_reg[3][5]/NET0131 ,
		_w2326_,
		_w2339_,
		_w4605_
	);
	LUT2 #(
		.INIT('h1)
	) name4153 (
		_w2342_,
		_w4605_,
		_w4606_
	);
	LUT4 #(
		.INIT('h0057)
	) name4154 (
		\DataWidth_reg[1]/NET0131 ,
		_w4603_,
		_w4604_,
		_w4606_,
		_w4607_
	);
	LUT4 #(
		.INIT('hc055)
	) name4155 (
		\InstQueue_reg[3][5]/NET0131 ,
		_w534_,
		_w539_,
		_w2339_,
		_w4608_
	);
	LUT2 #(
		.INIT('h2)
	) name4156 (
		\InstQueue_reg[3][5]/NET0131 ,
		_w2227_,
		_w4609_
	);
	LUT3 #(
		.INIT('h0d)
	) name4157 (
		_w1212_,
		_w4605_,
		_w4609_,
		_w4610_
	);
	LUT3 #(
		.INIT('hd0)
	) name4158 (
		_w710_,
		_w4608_,
		_w4610_,
		_w4611_
	);
	LUT3 #(
		.INIT('h2f)
	) name4159 (
		_w695_,
		_w4607_,
		_w4611_,
		_w4612_
	);
	LUT4 #(
		.INIT('h6c00)
	) name4160 (
		\Datai[28]_pad ,
		\Datai[29]_pad ,
		_w2209_,
		_w2313_,
		_w4613_
	);
	LUT3 #(
		.INIT('h60)
	) name4161 (
		\Datai[21]_pad ,
		_w2212_,
		_w2326_,
		_w4614_
	);
	LUT4 #(
		.INIT('h5553)
	) name4162 (
		\Datai[5]_pad ,
		\InstQueue_reg[4][5]/NET0131 ,
		_w2339_,
		_w2352_,
		_w4615_
	);
	LUT2 #(
		.INIT('h1)
	) name4163 (
		_w2355_,
		_w4615_,
		_w4616_
	);
	LUT4 #(
		.INIT('h0057)
	) name4164 (
		\DataWidth_reg[1]/NET0131 ,
		_w4613_,
		_w4614_,
		_w4616_,
		_w4617_
	);
	LUT4 #(
		.INIT('hc055)
	) name4165 (
		\InstQueue_reg[4][5]/NET0131 ,
		_w534_,
		_w539_,
		_w2352_,
		_w4618_
	);
	LUT2 #(
		.INIT('h2)
	) name4166 (
		\InstQueue_reg[4][5]/NET0131 ,
		_w2227_,
		_w4619_
	);
	LUT3 #(
		.INIT('h0d)
	) name4167 (
		_w1212_,
		_w4615_,
		_w4619_,
		_w4620_
	);
	LUT3 #(
		.INIT('hd0)
	) name4168 (
		_w710_,
		_w4618_,
		_w4620_,
		_w4621_
	);
	LUT3 #(
		.INIT('h2f)
	) name4169 (
		_w695_,
		_w4617_,
		_w4621_,
		_w4622_
	);
	LUT4 #(
		.INIT('h6c00)
	) name4170 (
		\Datai[28]_pad ,
		\Datai[29]_pad ,
		_w2209_,
		_w2326_,
		_w4623_
	);
	LUT3 #(
		.INIT('h60)
	) name4171 (
		\Datai[21]_pad ,
		_w2212_,
		_w2339_,
		_w4624_
	);
	LUT4 #(
		.INIT('h5553)
	) name4172 (
		\Datai[5]_pad ,
		\InstQueue_reg[5][5]/NET0131 ,
		_w2352_,
		_w2365_,
		_w4625_
	);
	LUT2 #(
		.INIT('h1)
	) name4173 (
		_w2368_,
		_w4625_,
		_w4626_
	);
	LUT4 #(
		.INIT('h0057)
	) name4174 (
		\DataWidth_reg[1]/NET0131 ,
		_w4623_,
		_w4624_,
		_w4626_,
		_w4627_
	);
	LUT4 #(
		.INIT('hc055)
	) name4175 (
		\InstQueue_reg[5][5]/NET0131 ,
		_w534_,
		_w539_,
		_w2365_,
		_w4628_
	);
	LUT2 #(
		.INIT('h2)
	) name4176 (
		\InstQueue_reg[5][5]/NET0131 ,
		_w2227_,
		_w4629_
	);
	LUT3 #(
		.INIT('h0d)
	) name4177 (
		_w1212_,
		_w4625_,
		_w4629_,
		_w4630_
	);
	LUT3 #(
		.INIT('hd0)
	) name4178 (
		_w710_,
		_w4628_,
		_w4630_,
		_w4631_
	);
	LUT3 #(
		.INIT('h2f)
	) name4179 (
		_w695_,
		_w4627_,
		_w4631_,
		_w4632_
	);
	LUT4 #(
		.INIT('h6c00)
	) name4180 (
		\Datai[28]_pad ,
		\Datai[29]_pad ,
		_w2209_,
		_w2339_,
		_w4633_
	);
	LUT3 #(
		.INIT('h60)
	) name4181 (
		\Datai[21]_pad ,
		_w2212_,
		_w2352_,
		_w4634_
	);
	LUT4 #(
		.INIT('h5553)
	) name4182 (
		\Datai[5]_pad ,
		\InstQueue_reg[6][5]/NET0131 ,
		_w2365_,
		_w2378_,
		_w4635_
	);
	LUT2 #(
		.INIT('h1)
	) name4183 (
		_w2381_,
		_w4635_,
		_w4636_
	);
	LUT4 #(
		.INIT('h0057)
	) name4184 (
		\DataWidth_reg[1]/NET0131 ,
		_w4633_,
		_w4634_,
		_w4636_,
		_w4637_
	);
	LUT4 #(
		.INIT('hc055)
	) name4185 (
		\InstQueue_reg[6][5]/NET0131 ,
		_w534_,
		_w539_,
		_w2378_,
		_w4638_
	);
	LUT2 #(
		.INIT('h2)
	) name4186 (
		\InstQueue_reg[6][5]/NET0131 ,
		_w2227_,
		_w4639_
	);
	LUT3 #(
		.INIT('h0d)
	) name4187 (
		_w1212_,
		_w4635_,
		_w4639_,
		_w4640_
	);
	LUT3 #(
		.INIT('hd0)
	) name4188 (
		_w710_,
		_w4638_,
		_w4640_,
		_w4641_
	);
	LUT3 #(
		.INIT('h2f)
	) name4189 (
		_w695_,
		_w4637_,
		_w4641_,
		_w4642_
	);
	LUT4 #(
		.INIT('h6c00)
	) name4190 (
		\Datai[28]_pad ,
		\Datai[29]_pad ,
		_w2209_,
		_w2352_,
		_w4643_
	);
	LUT3 #(
		.INIT('h60)
	) name4191 (
		\Datai[21]_pad ,
		_w2212_,
		_w2365_,
		_w4644_
	);
	LUT4 #(
		.INIT('h5553)
	) name4192 (
		\Datai[5]_pad ,
		\InstQueue_reg[7][5]/NET0131 ,
		_w2232_,
		_w2378_,
		_w4645_
	);
	LUT2 #(
		.INIT('h1)
	) name4193 (
		_w2393_,
		_w4645_,
		_w4646_
	);
	LUT4 #(
		.INIT('h0057)
	) name4194 (
		\DataWidth_reg[1]/NET0131 ,
		_w4643_,
		_w4644_,
		_w4646_,
		_w4647_
	);
	LUT4 #(
		.INIT('hc055)
	) name4195 (
		\InstQueue_reg[7][5]/NET0131 ,
		_w534_,
		_w539_,
		_w2232_,
		_w4648_
	);
	LUT2 #(
		.INIT('h2)
	) name4196 (
		\InstQueue_reg[7][5]/NET0131 ,
		_w2227_,
		_w4649_
	);
	LUT3 #(
		.INIT('h0d)
	) name4197 (
		_w1212_,
		_w4645_,
		_w4649_,
		_w4650_
	);
	LUT3 #(
		.INIT('hd0)
	) name4198 (
		_w710_,
		_w4648_,
		_w4650_,
		_w4651_
	);
	LUT3 #(
		.INIT('h2f)
	) name4199 (
		_w695_,
		_w4647_,
		_w4651_,
		_w4652_
	);
	LUT4 #(
		.INIT('h6c00)
	) name4200 (
		\Datai[28]_pad ,
		\Datai[29]_pad ,
		_w2209_,
		_w2365_,
		_w4653_
	);
	LUT3 #(
		.INIT('h60)
	) name4201 (
		\Datai[21]_pad ,
		_w2212_,
		_w2378_,
		_w4654_
	);
	LUT4 #(
		.INIT('h5553)
	) name4202 (
		\Datai[5]_pad ,
		\InstQueue_reg[8][5]/NET0131 ,
		_w2232_,
		_w2234_,
		_w4655_
	);
	LUT2 #(
		.INIT('h1)
	) name4203 (
		_w2404_,
		_w4655_,
		_w4656_
	);
	LUT4 #(
		.INIT('h0057)
	) name4204 (
		\DataWidth_reg[1]/NET0131 ,
		_w4653_,
		_w4654_,
		_w4656_,
		_w4657_
	);
	LUT4 #(
		.INIT('hc055)
	) name4205 (
		\InstQueue_reg[8][5]/NET0131 ,
		_w534_,
		_w539_,
		_w2234_,
		_w4658_
	);
	LUT2 #(
		.INIT('h2)
	) name4206 (
		\InstQueue_reg[8][5]/NET0131 ,
		_w2227_,
		_w4659_
	);
	LUT3 #(
		.INIT('h0d)
	) name4207 (
		_w1212_,
		_w4655_,
		_w4659_,
		_w4660_
	);
	LUT3 #(
		.INIT('hd0)
	) name4208 (
		_w710_,
		_w4658_,
		_w4660_,
		_w4661_
	);
	LUT3 #(
		.INIT('h2f)
	) name4209 (
		_w695_,
		_w4657_,
		_w4661_,
		_w4662_
	);
	LUT4 #(
		.INIT('h6c00)
	) name4210 (
		\Datai[28]_pad ,
		\Datai[29]_pad ,
		_w2209_,
		_w2378_,
		_w4663_
	);
	LUT3 #(
		.INIT('h60)
	) name4211 (
		\Datai[21]_pad ,
		_w2212_,
		_w2232_,
		_w4664_
	);
	LUT4 #(
		.INIT('h5553)
	) name4212 (
		\Datai[5]_pad ,
		\InstQueue_reg[9][5]/NET0131 ,
		_w2237_,
		_w2234_,
		_w4665_
	);
	LUT2 #(
		.INIT('h1)
	) name4213 (
		_w2415_,
		_w4665_,
		_w4666_
	);
	LUT4 #(
		.INIT('h0057)
	) name4214 (
		\DataWidth_reg[1]/NET0131 ,
		_w4663_,
		_w4664_,
		_w4666_,
		_w4667_
	);
	LUT4 #(
		.INIT('hc055)
	) name4215 (
		\InstQueue_reg[9][5]/NET0131 ,
		_w534_,
		_w539_,
		_w2237_,
		_w4668_
	);
	LUT2 #(
		.INIT('h2)
	) name4216 (
		\InstQueue_reg[9][5]/NET0131 ,
		_w2227_,
		_w4669_
	);
	LUT3 #(
		.INIT('h0d)
	) name4217 (
		_w1212_,
		_w4665_,
		_w4669_,
		_w4670_
	);
	LUT3 #(
		.INIT('hd0)
	) name4218 (
		_w710_,
		_w4668_,
		_w4670_,
		_w4671_
	);
	LUT3 #(
		.INIT('h2f)
	) name4219 (
		_w695_,
		_w4667_,
		_w4671_,
		_w4672_
	);
	LUT2 #(
		.INIT('he)
	) name4220 (
		\rEIP_reg[0]/NET0131 ,
		\rEIP_reg[1]/NET0131 ,
		_w4673_
	);
	LUT3 #(
		.INIT('he0)
	) name4221 (
		\rEIP_reg[0]/NET0131 ,
		\rEIP_reg[1]/NET0131 ,
		\rEIP_reg[31]/NET0131 ,
		_w4674_
	);
	LUT4 #(
		.INIT('he000)
	) name4222 (
		\rEIP_reg[0]/NET0131 ,
		\rEIP_reg[1]/NET0131 ,
		\rEIP_reg[2]/NET0131 ,
		\rEIP_reg[31]/NET0131 ,
		_w4675_
	);
	LUT3 #(
		.INIT('h80)
	) name4223 (
		\rEIP_reg[3]/NET0131 ,
		\rEIP_reg[4]/NET0131 ,
		_w4675_,
		_w4676_
	);
	LUT4 #(
		.INIT('h8000)
	) name4224 (
		\rEIP_reg[3]/NET0131 ,
		\rEIP_reg[4]/NET0131 ,
		\rEIP_reg[5]/NET0131 ,
		_w4675_,
		_w4677_
	);
	LUT3 #(
		.INIT('h80)
	) name4225 (
		\rEIP_reg[6]/NET0131 ,
		\rEIP_reg[7]/NET0131 ,
		_w4677_,
		_w4678_
	);
	LUT4 #(
		.INIT('h8000)
	) name4226 (
		\rEIP_reg[6]/NET0131 ,
		\rEIP_reg[7]/NET0131 ,
		\rEIP_reg[8]/NET0131 ,
		_w4677_,
		_w4679_
	);
	LUT3 #(
		.INIT('h80)
	) name4227 (
		\rEIP_reg[10]/NET0131 ,
		\rEIP_reg[9]/NET0131 ,
		_w4679_,
		_w4680_
	);
	LUT4 #(
		.INIT('h8000)
	) name4228 (
		\rEIP_reg[10]/NET0131 ,
		\rEIP_reg[11]/NET0131 ,
		\rEIP_reg[9]/NET0131 ,
		_w4679_,
		_w4681_
	);
	LUT3 #(
		.INIT('h80)
	) name4229 (
		\rEIP_reg[14]/NET0131 ,
		_w3151_,
		_w4681_,
		_w4682_
	);
	LUT4 #(
		.INIT('h8000)
	) name4230 (
		\rEIP_reg[14]/NET0131 ,
		\rEIP_reg[15]/NET0131 ,
		_w3151_,
		_w4681_,
		_w4683_
	);
	LUT3 #(
		.INIT('h80)
	) name4231 (
		\rEIP_reg[16]/NET0131 ,
		_w3196_,
		_w4683_,
		_w4684_
	);
	LUT4 #(
		.INIT('h8000)
	) name4232 (
		\rEIP_reg[16]/NET0131 ,
		\rEIP_reg[23]/NET0131 ,
		_w3196_,
		_w4683_,
		_w4685_
	);
	LUT3 #(
		.INIT('h80)
	) name4233 (
		\rEIP_reg[26]/NET0131 ,
		_w3249_,
		_w4685_,
		_w4686_
	);
	LUT4 #(
		.INIT('h8000)
	) name4234 (
		\rEIP_reg[26]/NET0131 ,
		\rEIP_reg[27]/NET0131 ,
		_w3249_,
		_w4685_,
		_w4687_
	);
	LUT3 #(
		.INIT('h80)
	) name4235 (
		\rEIP_reg[28]/NET0131 ,
		\rEIP_reg[29]/NET0131 ,
		_w4687_,
		_w4688_
	);
	LUT4 #(
		.INIT('h8000)
	) name4236 (
		\rEIP_reg[28]/NET0131 ,
		\rEIP_reg[29]/NET0131 ,
		\rEIP_reg[30]/NET0131 ,
		_w4687_,
		_w4689_
	);
	LUT3 #(
		.INIT('h8a)
	) name4237 (
		\Address[28]_pad ,
		\State_reg[0]/NET0131 ,
		\State_reg[1]/NET0131 ,
		_w4690_
	);
	LUT2 #(
		.INIT('h8)
	) name4238 (
		\rEIP_reg[0]/NET0131 ,
		\rEIP_reg[31]/NET0131 ,
		_w4691_
	);
	LUT4 #(
		.INIT('h8000)
	) name4239 (
		\rEIP_reg[23]/NET0131 ,
		_w3155_,
		_w3196_,
		_w4691_,
		_w4692_
	);
	LUT3 #(
		.INIT('h80)
	) name4240 (
		\rEIP_reg[27]/NET0131 ,
		_w3269_,
		_w4692_,
		_w4693_
	);
	LUT4 #(
		.INIT('h8000)
	) name4241 (
		\rEIP_reg[27]/NET0131 ,
		\rEIP_reg[28]/NET0131 ,
		_w3269_,
		_w4692_,
		_w4694_
	);
	LUT3 #(
		.INIT('h40)
	) name4242 (
		\State_reg[0]/NET0131 ,
		\State_reg[1]/NET0131 ,
		\State_reg[2]/NET0131 ,
		_w4695_
	);
	LUT4 #(
		.INIT('h2313)
	) name4243 (
		\rEIP_reg[29]/NET0131 ,
		_w4690_,
		_w4695_,
		_w4694_,
		_w4696_
	);
	LUT4 #(
		.INIT('h48ff)
	) name4244 (
		\rEIP_reg[30]/NET0131 ,
		_w592_,
		_w4688_,
		_w4696_,
		_w4697_
	);
	LUT3 #(
		.INIT('h21)
	) name4245 (
		\EAX_reg[25]/NET0131 ,
		_w594_,
		_w2093_,
		_w4698_
	);
	LUT3 #(
		.INIT('h02)
	) name4246 (
		_w589_,
		_w566_,
		_w4698_,
		_w4699_
	);
	LUT4 #(
		.INIT('haaa2)
	) name4247 (
		\Datao[25]_pad ,
		_w646_,
		_w2183_,
		_w4699_,
		_w4700_
	);
	LUT4 #(
		.INIT('h0200)
	) name4248 (
		_w589_,
		_w594_,
		_w566_,
		_w4064_,
		_w4701_
	);
	LUT4 #(
		.INIT('h3f15)
	) name4249 (
		\Datao[25]_pad ,
		\uWord_reg[9]/NET0131 ,
		_w2179_,
		_w2180_,
		_w4702_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name4250 (
		_w690_,
		_w4700_,
		_w4701_,
		_w4702_,
		_w4703_
	);
	LUT4 #(
		.INIT('h20aa)
	) name4251 (
		\Datao[17]_pad ,
		_w596_,
		_w690_,
		_w2180_,
		_w4704_
	);
	LUT2 #(
		.INIT('h8)
	) name4252 (
		\uWord_reg[1]/NET0131 ,
		_w2179_,
		_w4705_
	);
	LUT2 #(
		.INIT('h4)
	) name4253 (
		_w594_,
		_w690_,
		_w4706_
	);
	LUT4 #(
		.INIT('h2000)
	) name4254 (
		_w589_,
		_w566_,
		_w4034_,
		_w4706_,
		_w4707_
	);
	LUT2 #(
		.INIT('h1)
	) name4255 (
		_w4705_,
		_w4707_,
		_w4708_
	);
	LUT2 #(
		.INIT('hb)
	) name4256 (
		_w4704_,
		_w4708_,
		_w4709_
	);
	LUT4 #(
		.INIT('h0509)
	) name4257 (
		\EAX_reg[16]/NET0131 ,
		\EAX_reg[31]/NET0131 ,
		_w594_,
		_w2091_,
		_w4710_
	);
	LUT3 #(
		.INIT('h02)
	) name4258 (
		_w589_,
		_w566_,
		_w4710_,
		_w4711_
	);
	LUT4 #(
		.INIT('haaa2)
	) name4259 (
		\Datao[16]_pad ,
		_w646_,
		_w2183_,
		_w4711_,
		_w4712_
	);
	LUT4 #(
		.INIT('h0200)
	) name4260 (
		_w589_,
		_w594_,
		_w566_,
		_w4011_,
		_w4713_
	);
	LUT4 #(
		.INIT('h3f15)
	) name4261 (
		\Datao[16]_pad ,
		\uWord_reg[0]/NET0131 ,
		_w2179_,
		_w2180_,
		_w4714_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name4262 (
		_w690_,
		_w4712_,
		_w4713_,
		_w4714_,
		_w4715_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name4263 (
		\Datao[21]_pad ,
		_w594_,
		_w596_,
		_w4054_,
		_w4716_
	);
	LUT4 #(
		.INIT('h3f15)
	) name4264 (
		\Datao[21]_pad ,
		\uWord_reg[5]/NET0131 ,
		_w2179_,
		_w2180_,
		_w4717_
	);
	LUT3 #(
		.INIT('h2f)
	) name4265 (
		_w690_,
		_w4716_,
		_w4717_,
		_w4718_
	);
	LUT4 #(
		.INIT('h1050)
	) name4266 (
		\Flush_reg/NET0131 ,
		\InstQueueRd_Addr_reg[2]/NET0131 ,
		_w700_,
		_w702_,
		_w4719_
	);
	LUT4 #(
		.INIT('hfd9f)
	) name4267 (
		\State2_reg[0]/NET0131 ,
		\State2_reg[1]/NET0131 ,
		\State2_reg[2]/NET0131 ,
		\State2_reg[3]/NET0131 ,
		_w4720_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name4268 (
		\InstQueueWr_Addr_reg[2]/NET0131 ,
		_w3680_,
		_w4719_,
		_w4720_,
		_w4721_
	);
	LUT4 #(
		.INIT('hcc08)
	) name4269 (
		\DataWidth_reg[1]/NET0131 ,
		\InstQueueWr_Addr_reg[2]/NET0131 ,
		_w1212_,
		_w2214_,
		_w4722_
	);
	LUT3 #(
		.INIT('h54)
	) name4270 (
		_w710_,
		_w1305_,
		_w4722_,
		_w4723_
	);
	LUT2 #(
		.INIT('h4)
	) name4271 (
		_w1305_,
		_w2214_,
		_w4724_
	);
	LUT3 #(
		.INIT('h07)
	) name4272 (
		\InstQueueWr_Addr_reg[0]/NET0131 ,
		\InstQueueWr_Addr_reg[1]/NET0131 ,
		\InstQueueWr_Addr_reg[2]/NET0131 ,
		_w4725_
	);
	LUT3 #(
		.INIT('h70)
	) name4273 (
		\DataWidth_reg[1]/NET0131 ,
		_w695_,
		_w4725_,
		_w4726_
	);
	LUT3 #(
		.INIT('h45)
	) name4274 (
		_w2218_,
		_w4724_,
		_w4726_,
		_w4727_
	);
	LUT3 #(
		.INIT('hba)
	) name4275 (
		_w4721_,
		_w4723_,
		_w4727_,
		_w4728_
	);
	LUT4 #(
		.INIT('h070f)
	) name4276 (
		\rEIP_reg[16]/NET0131 ,
		\rEIP_reg[17]/NET0131 ,
		\rEIP_reg[18]/NET0131 ,
		_w4683_,
		_w4729_
	);
	LUT3 #(
		.INIT('h80)
	) name4277 (
		\rEIP_reg[16]/NET0131 ,
		_w3156_,
		_w4683_,
		_w4730_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name4278 (
		\rEIP_reg[16]/NET0131 ,
		_w592_,
		_w3156_,
		_w4683_,
		_w4731_
	);
	LUT3 #(
		.INIT('h8a)
	) name4279 (
		\Address[16]_pad ,
		\State_reg[0]/NET0131 ,
		\State_reg[1]/NET0131 ,
		_w4732_
	);
	LUT4 #(
		.INIT('h60a0)
	) name4280 (
		\rEIP_reg[17]/NET0131 ,
		_w3155_,
		_w4695_,
		_w4691_,
		_w4733_
	);
	LUT2 #(
		.INIT('h1)
	) name4281 (
		_w4732_,
		_w4733_,
		_w4734_
	);
	LUT3 #(
		.INIT('h4f)
	) name4282 (
		_w4729_,
		_w4731_,
		_w4734_,
		_w4735_
	);
	LUT4 #(
		.INIT('hca00)
	) name4283 (
		\Datao[2]_pad ,
		\EAX_reg[2]/NET0131 ,
		_w596_,
		_w690_,
		_w4736_
	);
	LUT4 #(
		.INIT('h3f15)
	) name4284 (
		\Datao[2]_pad ,
		\lWord_reg[2]/NET0131 ,
		_w2179_,
		_w2180_,
		_w4737_
	);
	LUT2 #(
		.INIT('hb)
	) name4285 (
		_w4736_,
		_w4737_,
		_w4738_
	);
	LUT4 #(
		.INIT('hca00)
	) name4286 (
		\Datao[4]_pad ,
		\EAX_reg[4]/NET0131 ,
		_w596_,
		_w690_,
		_w4739_
	);
	LUT4 #(
		.INIT('h3f15)
	) name4287 (
		\Datao[4]_pad ,
		\lWord_reg[4]/NET0131 ,
		_w2179_,
		_w2180_,
		_w4740_
	);
	LUT2 #(
		.INIT('hb)
	) name4288 (
		_w4739_,
		_w4740_,
		_w4741_
	);
	LUT4 #(
		.INIT('hca00)
	) name4289 (
		\Datao[3]_pad ,
		\EAX_reg[3]/NET0131 ,
		_w596_,
		_w690_,
		_w4742_
	);
	LUT4 #(
		.INIT('h3f15)
	) name4290 (
		\Datao[3]_pad ,
		\lWord_reg[3]/NET0131 ,
		_w2179_,
		_w2180_,
		_w4743_
	);
	LUT2 #(
		.INIT('hb)
	) name4291 (
		_w4742_,
		_w4743_,
		_w4744_
	);
	LUT4 #(
		.INIT('hca00)
	) name4292 (
		\Datao[5]_pad ,
		\EAX_reg[5]/NET0131 ,
		_w596_,
		_w690_,
		_w4745_
	);
	LUT4 #(
		.INIT('h3f15)
	) name4293 (
		\Datao[5]_pad ,
		\lWord_reg[5]/NET0131 ,
		_w2179_,
		_w2180_,
		_w4746_
	);
	LUT2 #(
		.INIT('hb)
	) name4294 (
		_w4745_,
		_w4746_,
		_w4747_
	);
	LUT4 #(
		.INIT('hca00)
	) name4295 (
		\Datao[6]_pad ,
		\EAX_reg[6]/NET0131 ,
		_w596_,
		_w690_,
		_w4748_
	);
	LUT4 #(
		.INIT('h3f15)
	) name4296 (
		\Datao[6]_pad ,
		\lWord_reg[6]/NET0131 ,
		_w2179_,
		_w2180_,
		_w4749_
	);
	LUT2 #(
		.INIT('hb)
	) name4297 (
		_w4748_,
		_w4749_,
		_w4750_
	);
	LUT4 #(
		.INIT('hca00)
	) name4298 (
		\Datao[7]_pad ,
		\EAX_reg[7]/NET0131 ,
		_w596_,
		_w690_,
		_w4751_
	);
	LUT4 #(
		.INIT('h3f15)
	) name4299 (
		\Datao[7]_pad ,
		\lWord_reg[7]/NET0131 ,
		_w2179_,
		_w2180_,
		_w4752_
	);
	LUT2 #(
		.INIT('hb)
	) name4300 (
		_w4751_,
		_w4752_,
		_w4753_
	);
	LUT4 #(
		.INIT('hca00)
	) name4301 (
		\Datao[8]_pad ,
		\EAX_reg[8]/NET0131 ,
		_w596_,
		_w690_,
		_w4754_
	);
	LUT4 #(
		.INIT('h3f15)
	) name4302 (
		\Datao[8]_pad ,
		\lWord_reg[8]/NET0131 ,
		_w2179_,
		_w2180_,
		_w4755_
	);
	LUT2 #(
		.INIT('hb)
	) name4303 (
		_w4754_,
		_w4755_,
		_w4756_
	);
	LUT4 #(
		.INIT('hca00)
	) name4304 (
		\Datao[9]_pad ,
		\EAX_reg[9]/NET0131 ,
		_w596_,
		_w690_,
		_w4757_
	);
	LUT4 #(
		.INIT('h3f15)
	) name4305 (
		\Datao[9]_pad ,
		\lWord_reg[9]/NET0131 ,
		_w2179_,
		_w2180_,
		_w4758_
	);
	LUT2 #(
		.INIT('hb)
	) name4306 (
		_w4757_,
		_w4758_,
		_w4759_
	);
	LUT4 #(
		.INIT('hca00)
	) name4307 (
		\Datao[0]_pad ,
		\EAX_reg[0]/NET0131 ,
		_w596_,
		_w690_,
		_w4760_
	);
	LUT4 #(
		.INIT('h3f15)
	) name4308 (
		\Datao[0]_pad ,
		\lWord_reg[0]/NET0131 ,
		_w2179_,
		_w2180_,
		_w4761_
	);
	LUT2 #(
		.INIT('hb)
	) name4309 (
		_w4760_,
		_w4761_,
		_w4762_
	);
	LUT4 #(
		.INIT('hca00)
	) name4310 (
		\Datao[10]_pad ,
		\EAX_reg[10]/NET0131 ,
		_w596_,
		_w690_,
		_w4763_
	);
	LUT4 #(
		.INIT('h3f15)
	) name4311 (
		\Datao[10]_pad ,
		\lWord_reg[10]/NET0131 ,
		_w2179_,
		_w2180_,
		_w4764_
	);
	LUT2 #(
		.INIT('hb)
	) name4312 (
		_w4763_,
		_w4764_,
		_w4765_
	);
	LUT4 #(
		.INIT('hca00)
	) name4313 (
		\Datao[12]_pad ,
		\EAX_reg[12]/NET0131 ,
		_w596_,
		_w690_,
		_w4766_
	);
	LUT4 #(
		.INIT('h3f15)
	) name4314 (
		\Datao[12]_pad ,
		\lWord_reg[12]/NET0131 ,
		_w2179_,
		_w2180_,
		_w4767_
	);
	LUT2 #(
		.INIT('hb)
	) name4315 (
		_w4766_,
		_w4767_,
		_w4768_
	);
	LUT4 #(
		.INIT('hca00)
	) name4316 (
		\Datao[11]_pad ,
		\EAX_reg[11]/NET0131 ,
		_w596_,
		_w690_,
		_w4769_
	);
	LUT4 #(
		.INIT('h3f15)
	) name4317 (
		\Datao[11]_pad ,
		\lWord_reg[11]/NET0131 ,
		_w2179_,
		_w2180_,
		_w4770_
	);
	LUT2 #(
		.INIT('hb)
	) name4318 (
		_w4769_,
		_w4770_,
		_w4771_
	);
	LUT4 #(
		.INIT('hca00)
	) name4319 (
		\Datao[13]_pad ,
		\EAX_reg[13]/NET0131 ,
		_w596_,
		_w690_,
		_w4772_
	);
	LUT4 #(
		.INIT('h3f15)
	) name4320 (
		\Datao[13]_pad ,
		\lWord_reg[13]/NET0131 ,
		_w2179_,
		_w2180_,
		_w4773_
	);
	LUT2 #(
		.INIT('hb)
	) name4321 (
		_w4772_,
		_w4773_,
		_w4774_
	);
	LUT4 #(
		.INIT('hca00)
	) name4322 (
		\Datao[14]_pad ,
		\EAX_reg[14]/NET0131 ,
		_w596_,
		_w690_,
		_w4775_
	);
	LUT4 #(
		.INIT('h3f15)
	) name4323 (
		\Datao[14]_pad ,
		\lWord_reg[14]/NET0131 ,
		_w2179_,
		_w2180_,
		_w4776_
	);
	LUT2 #(
		.INIT('hb)
	) name4324 (
		_w4775_,
		_w4776_,
		_w4777_
	);
	LUT4 #(
		.INIT('hca00)
	) name4325 (
		\Datao[15]_pad ,
		\EAX_reg[15]/NET0131 ,
		_w596_,
		_w690_,
		_w4778_
	);
	LUT4 #(
		.INIT('h3f15)
	) name4326 (
		\Datao[15]_pad ,
		\lWord_reg[15]/NET0131 ,
		_w2179_,
		_w2180_,
		_w4779_
	);
	LUT2 #(
		.INIT('hb)
	) name4327 (
		_w4778_,
		_w4779_,
		_w4780_
	);
	LUT4 #(
		.INIT('hca00)
	) name4328 (
		\Datao[1]_pad ,
		\EAX_reg[1]/NET0131 ,
		_w596_,
		_w690_,
		_w4781_
	);
	LUT4 #(
		.INIT('h3f15)
	) name4329 (
		\Datao[1]_pad ,
		\lWord_reg[1]/NET0131 ,
		_w2179_,
		_w2180_,
		_w4782_
	);
	LUT2 #(
		.INIT('hb)
	) name4330 (
		_w4781_,
		_w4782_,
		_w4783_
	);
	LUT4 #(
		.INIT('h807f)
	) name4331 (
		\InstQueueWr_Addr_reg[0]/NET0131 ,
		\InstQueueWr_Addr_reg[1]/NET0131 ,
		\InstQueueWr_Addr_reg[2]/NET0131 ,
		\InstQueueWr_Addr_reg[3]/NET0131 ,
		_w4784_
	);
	LUT4 #(
		.INIT('hc03f)
	) name4332 (
		\InstQueueWr_Addr_reg[0]/NET0131 ,
		\InstQueueWr_Addr_reg[1]/NET0131 ,
		\InstQueueWr_Addr_reg[2]/NET0131 ,
		\InstQueueWr_Addr_reg[3]/NET0131 ,
		_w4785_
	);
	LUT4 #(
		.INIT('he00f)
	) name4333 (
		\InstQueueWr_Addr_reg[0]/NET0131 ,
		\InstQueueWr_Addr_reg[1]/NET0131 ,
		\InstQueueWr_Addr_reg[2]/NET0131 ,
		\InstQueueWr_Addr_reg[3]/NET0131 ,
		_w4786_
	);
	LUT4 #(
		.INIT('h0008)
	) name4334 (
		\DataWidth_reg[1]/NET0131 ,
		_w695_,
		_w2265_,
		_w4786_,
		_w4787_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name4335 (
		\InstQueueWr_Addr_reg[3]/NET0131 ,
		_w3680_,
		_w4719_,
		_w4720_,
		_w4788_
	);
	LUT2 #(
		.INIT('h2)
	) name4336 (
		_w710_,
		_w4784_,
		_w4789_
	);
	LUT4 #(
		.INIT('h00f4)
	) name4337 (
		\DataWidth_reg[1]/NET0131 ,
		_w695_,
		_w1212_,
		_w4785_,
		_w4790_
	);
	LUT2 #(
		.INIT('h1)
	) name4338 (
		_w4789_,
		_w4790_,
		_w4791_
	);
	LUT3 #(
		.INIT('hef)
	) name4339 (
		_w4787_,
		_w4788_,
		_w4791_,
		_w4792_
	);
	LUT3 #(
		.INIT('h8a)
	) name4340 (
		\InstQueueWr_Addr_reg[1]/NET0131 ,
		_w4719_,
		_w4720_,
		_w4793_
	);
	LUT2 #(
		.INIT('h4)
	) name4341 (
		\InstQueueWr_Addr_reg[0]/NET0131 ,
		_w710_,
		_w4794_
	);
	LUT4 #(
		.INIT('h4c00)
	) name4342 (
		\DataWidth_reg[1]/NET0131 ,
		\InstQueueWr_Addr_reg[1]/NET0131 ,
		_w695_,
		_w3680_,
		_w4795_
	);
	LUT3 #(
		.INIT('h13)
	) name4343 (
		\InstQueueWr_Addr_reg[0]/NET0131 ,
		\InstQueueWr_Addr_reg[1]/NET0131 ,
		_w710_,
		_w4796_
	);
	LUT4 #(
		.INIT('h8acf)
	) name4344 (
		_w1306_,
		_w4794_,
		_w4795_,
		_w4796_,
		_w4797_
	);
	LUT2 #(
		.INIT('he)
	) name4345 (
		_w4793_,
		_w4797_,
		_w4798_
	);
	LUT4 #(
		.INIT('hfd80)
	) name4346 (
		\State2_reg[0]/NET0131 ,
		\State2_reg[1]/NET0131 ,
		\State2_reg[2]/NET0131 ,
		\State2_reg[3]/NET0131 ,
		_w4799_
	);
	LUT2 #(
		.INIT('h2)
	) name4347 (
		\InstQueueWr_Addr_reg[0]/NET0131 ,
		_w4799_,
		_w4800_
	);
	LUT2 #(
		.INIT('h1)
	) name4348 (
		\Flush_reg/NET0131 ,
		\InstQueueWr_Addr_reg[0]/NET0131 ,
		_w4801_
	);
	LUT4 #(
		.INIT('h002a)
	) name4349 (
		_w700_,
		_w701_,
		_w702_,
		_w4801_,
		_w4802_
	);
	LUT3 #(
		.INIT('hfe)
	) name4350 (
		_w4794_,
		_w4802_,
		_w4800_,
		_w4803_
	);
	LUT3 #(
		.INIT('h48)
	) name4351 (
		\Datai[25]_pad ,
		_w2199_,
		_w2208_,
		_w4804_
	);
	LUT4 #(
		.INIT('hcc6c)
	) name4352 (
		\Datai[16]_pad ,
		\Datai[17]_pad ,
		\Datai[31]_pad ,
		_w2204_,
		_w4805_
	);
	LUT2 #(
		.INIT('h8)
	) name4353 (
		_w2215_,
		_w4805_,
		_w4806_
	);
	LUT4 #(
		.INIT('h5553)
	) name4354 (
		\Datai[1]_pad ,
		\InstQueue_reg[0][1]/NET0131 ,
		_w2217_,
		_w2219_,
		_w4807_
	);
	LUT2 #(
		.INIT('h1)
	) name4355 (
		_w2223_,
		_w4807_,
		_w4808_
	);
	LUT4 #(
		.INIT('h0057)
	) name4356 (
		\DataWidth_reg[1]/NET0131 ,
		_w4804_,
		_w4806_,
		_w4808_,
		_w4809_
	);
	LUT4 #(
		.INIT('hc055)
	) name4357 (
		\InstQueue_reg[0][1]/NET0131 ,
		_w488_,
		_w493_,
		_w2217_,
		_w4810_
	);
	LUT2 #(
		.INIT('h2)
	) name4358 (
		\InstQueue_reg[0][1]/NET0131 ,
		_w2227_,
		_w4811_
	);
	LUT3 #(
		.INIT('h0d)
	) name4359 (
		_w1212_,
		_w4807_,
		_w4811_,
		_w4812_
	);
	LUT3 #(
		.INIT('hd0)
	) name4360 (
		_w710_,
		_w4810_,
		_w4812_,
		_w4813_
	);
	LUT3 #(
		.INIT('h2f)
	) name4361 (
		_w695_,
		_w4809_,
		_w4813_,
		_w4814_
	);
	LUT3 #(
		.INIT('h60)
	) name4362 (
		\Datai[25]_pad ,
		_w2208_,
		_w2232_,
		_w4815_
	);
	LUT2 #(
		.INIT('h8)
	) name4363 (
		_w2234_,
		_w4805_,
		_w4816_
	);
	LUT4 #(
		.INIT('h5553)
	) name4364 (
		\Datai[1]_pad ,
		\InstQueue_reg[10][1]/NET0131 ,
		_w2236_,
		_w2237_,
		_w4817_
	);
	LUT2 #(
		.INIT('h1)
	) name4365 (
		_w2241_,
		_w4817_,
		_w4818_
	);
	LUT4 #(
		.INIT('h0057)
	) name4366 (
		\DataWidth_reg[1]/NET0131 ,
		_w4815_,
		_w4816_,
		_w4818_,
		_w4819_
	);
	LUT4 #(
		.INIT('hc055)
	) name4367 (
		\InstQueue_reg[10][1]/NET0131 ,
		_w488_,
		_w493_,
		_w2236_,
		_w4820_
	);
	LUT2 #(
		.INIT('h2)
	) name4368 (
		\InstQueue_reg[10][1]/NET0131 ,
		_w2227_,
		_w4821_
	);
	LUT3 #(
		.INIT('h0d)
	) name4369 (
		_w1212_,
		_w4817_,
		_w4821_,
		_w4822_
	);
	LUT3 #(
		.INIT('hd0)
	) name4370 (
		_w710_,
		_w4820_,
		_w4822_,
		_w4823_
	);
	LUT3 #(
		.INIT('h2f)
	) name4371 (
		_w695_,
		_w4819_,
		_w4823_,
		_w4824_
	);
	LUT4 #(
		.INIT('ha666)
	) name4372 (
		\Datai[24]_pad ,
		\Datai[31]_pad ,
		_w2204_,
		_w2207_,
		_w4825_
	);
	LUT4 #(
		.INIT('ha600)
	) name4373 (
		\Datai[16]_pad ,
		\Datai[31]_pad ,
		_w2204_,
		_w2237_,
		_w4826_
	);
	LUT4 #(
		.INIT('haa80)
	) name4374 (
		\DataWidth_reg[1]/NET0131 ,
		_w2234_,
		_w4825_,
		_w4826_,
		_w4827_
	);
	LUT4 #(
		.INIT('h5553)
	) name4375 (
		\Datai[0]_pad ,
		\InstQueue_reg[11][0]/NET0131 ,
		_w2236_,
		_w2251_,
		_w4828_
	);
	LUT2 #(
		.INIT('h1)
	) name4376 (
		_w2255_,
		_w4828_,
		_w4829_
	);
	LUT3 #(
		.INIT('ha8)
	) name4377 (
		_w695_,
		_w4827_,
		_w4829_,
		_w4830_
	);
	LUT4 #(
		.INIT('hc055)
	) name4378 (
		\InstQueue_reg[11][0]/NET0131 ,
		_w500_,
		_w506_,
		_w2251_,
		_w4831_
	);
	LUT2 #(
		.INIT('h2)
	) name4379 (
		\InstQueue_reg[11][0]/NET0131 ,
		_w2227_,
		_w4832_
	);
	LUT3 #(
		.INIT('h0d)
	) name4380 (
		_w1212_,
		_w4828_,
		_w4832_,
		_w4833_
	);
	LUT3 #(
		.INIT('hd0)
	) name4381 (
		_w710_,
		_w4831_,
		_w4833_,
		_w4834_
	);
	LUT2 #(
		.INIT('hb)
	) name4382 (
		_w4830_,
		_w4834_,
		_w4835_
	);
	LUT3 #(
		.INIT('h60)
	) name4383 (
		\Datai[25]_pad ,
		_w2208_,
		_w2234_,
		_w4836_
	);
	LUT2 #(
		.INIT('h8)
	) name4384 (
		_w2237_,
		_w4805_,
		_w4837_
	);
	LUT4 #(
		.INIT('h5553)
	) name4385 (
		\Datai[1]_pad ,
		\InstQueue_reg[11][1]/NET0131 ,
		_w2236_,
		_w2251_,
		_w4838_
	);
	LUT2 #(
		.INIT('h1)
	) name4386 (
		_w2255_,
		_w4838_,
		_w4839_
	);
	LUT4 #(
		.INIT('h0057)
	) name4387 (
		\DataWidth_reg[1]/NET0131 ,
		_w4836_,
		_w4837_,
		_w4839_,
		_w4840_
	);
	LUT4 #(
		.INIT('hc055)
	) name4388 (
		\InstQueue_reg[11][1]/NET0131 ,
		_w488_,
		_w493_,
		_w2251_,
		_w4841_
	);
	LUT2 #(
		.INIT('h2)
	) name4389 (
		\InstQueue_reg[11][1]/NET0131 ,
		_w2227_,
		_w4842_
	);
	LUT3 #(
		.INIT('h0d)
	) name4390 (
		_w1212_,
		_w4838_,
		_w4842_,
		_w4843_
	);
	LUT3 #(
		.INIT('hd0)
	) name4391 (
		_w710_,
		_w4841_,
		_w4843_,
		_w4844_
	);
	LUT3 #(
		.INIT('h2f)
	) name4392 (
		_w695_,
		_w4840_,
		_w4844_,
		_w4845_
	);
	LUT3 #(
		.INIT('h60)
	) name4393 (
		\Datai[25]_pad ,
		_w2208_,
		_w2237_,
		_w4846_
	);
	LUT2 #(
		.INIT('h8)
	) name4394 (
		_w2236_,
		_w4805_,
		_w4847_
	);
	LUT4 #(
		.INIT('h5553)
	) name4395 (
		\Datai[1]_pad ,
		\InstQueue_reg[12][1]/NET0131 ,
		_w2251_,
		_w2265_,
		_w4848_
	);
	LUT2 #(
		.INIT('h1)
	) name4396 (
		_w2268_,
		_w4848_,
		_w4849_
	);
	LUT4 #(
		.INIT('h0057)
	) name4397 (
		\DataWidth_reg[1]/NET0131 ,
		_w4846_,
		_w4847_,
		_w4849_,
		_w4850_
	);
	LUT4 #(
		.INIT('hc055)
	) name4398 (
		\InstQueue_reg[12][1]/NET0131 ,
		_w488_,
		_w493_,
		_w2265_,
		_w4851_
	);
	LUT2 #(
		.INIT('h2)
	) name4399 (
		\InstQueue_reg[12][1]/NET0131 ,
		_w2227_,
		_w4852_
	);
	LUT3 #(
		.INIT('h0d)
	) name4400 (
		_w1212_,
		_w4848_,
		_w4852_,
		_w4853_
	);
	LUT3 #(
		.INIT('hd0)
	) name4401 (
		_w710_,
		_w4851_,
		_w4853_,
		_w4854_
	);
	LUT3 #(
		.INIT('h2f)
	) name4402 (
		_w695_,
		_w4850_,
		_w4854_,
		_w4855_
	);
	LUT3 #(
		.INIT('h60)
	) name4403 (
		\Datai[25]_pad ,
		_w2208_,
		_w2236_,
		_w4856_
	);
	LUT2 #(
		.INIT('h8)
	) name4404 (
		_w2251_,
		_w4805_,
		_w4857_
	);
	LUT4 #(
		.INIT('h5553)
	) name4405 (
		\Datai[1]_pad ,
		\InstQueue_reg[13][1]/NET0131 ,
		_w2199_,
		_w2265_,
		_w4858_
	);
	LUT2 #(
		.INIT('h1)
	) name4406 (
		_w2280_,
		_w4858_,
		_w4859_
	);
	LUT4 #(
		.INIT('h0057)
	) name4407 (
		\DataWidth_reg[1]/NET0131 ,
		_w4856_,
		_w4857_,
		_w4859_,
		_w4860_
	);
	LUT4 #(
		.INIT('hc055)
	) name4408 (
		\InstQueue_reg[13][1]/NET0131 ,
		_w488_,
		_w493_,
		_w2199_,
		_w4861_
	);
	LUT2 #(
		.INIT('h2)
	) name4409 (
		\InstQueue_reg[13][1]/NET0131 ,
		_w2227_,
		_w4862_
	);
	LUT3 #(
		.INIT('h0d)
	) name4410 (
		_w1212_,
		_w4858_,
		_w4862_,
		_w4863_
	);
	LUT3 #(
		.INIT('hd0)
	) name4411 (
		_w710_,
		_w4861_,
		_w4863_,
		_w4864_
	);
	LUT3 #(
		.INIT('h2f)
	) name4412 (
		_w695_,
		_w4860_,
		_w4864_,
		_w4865_
	);
	LUT3 #(
		.INIT('h60)
	) name4413 (
		\Datai[25]_pad ,
		_w2208_,
		_w2251_,
		_w4866_
	);
	LUT2 #(
		.INIT('h8)
	) name4414 (
		_w2265_,
		_w4805_,
		_w4867_
	);
	LUT4 #(
		.INIT('h5553)
	) name4415 (
		\Datai[1]_pad ,
		\InstQueue_reg[14][1]/NET0131 ,
		_w2199_,
		_w2215_,
		_w4868_
	);
	LUT2 #(
		.INIT('h1)
	) name4416 (
		_w2291_,
		_w4868_,
		_w4869_
	);
	LUT4 #(
		.INIT('h0057)
	) name4417 (
		\DataWidth_reg[1]/NET0131 ,
		_w4866_,
		_w4867_,
		_w4869_,
		_w4870_
	);
	LUT4 #(
		.INIT('hc055)
	) name4418 (
		\InstQueue_reg[14][1]/NET0131 ,
		_w488_,
		_w493_,
		_w2215_,
		_w4871_
	);
	LUT2 #(
		.INIT('h2)
	) name4419 (
		\InstQueue_reg[14][1]/NET0131 ,
		_w2227_,
		_w4872_
	);
	LUT3 #(
		.INIT('h0d)
	) name4420 (
		_w1212_,
		_w4868_,
		_w4872_,
		_w4873_
	);
	LUT3 #(
		.INIT('hd0)
	) name4421 (
		_w710_,
		_w4871_,
		_w4873_,
		_w4874_
	);
	LUT3 #(
		.INIT('h2f)
	) name4422 (
		_w695_,
		_w4870_,
		_w4874_,
		_w4875_
	);
	LUT3 #(
		.INIT('h60)
	) name4423 (
		\Datai[25]_pad ,
		_w2208_,
		_w2265_,
		_w4876_
	);
	LUT2 #(
		.INIT('h8)
	) name4424 (
		_w2199_,
		_w4805_,
		_w4877_
	);
	LUT4 #(
		.INIT('h5553)
	) name4425 (
		\Datai[1]_pad ,
		\InstQueue_reg[15][1]/NET0131 ,
		_w2219_,
		_w2215_,
		_w4878_
	);
	LUT2 #(
		.INIT('h1)
	) name4426 (
		_w2303_,
		_w4878_,
		_w4879_
	);
	LUT4 #(
		.INIT('h0057)
	) name4427 (
		\DataWidth_reg[1]/NET0131 ,
		_w4876_,
		_w4877_,
		_w4879_,
		_w4880_
	);
	LUT4 #(
		.INIT('hc055)
	) name4428 (
		\InstQueue_reg[15][1]/NET0131 ,
		_w488_,
		_w493_,
		_w2219_,
		_w4881_
	);
	LUT2 #(
		.INIT('h2)
	) name4429 (
		\InstQueue_reg[15][1]/NET0131 ,
		_w2227_,
		_w4882_
	);
	LUT3 #(
		.INIT('h0d)
	) name4430 (
		_w1212_,
		_w4878_,
		_w4882_,
		_w4883_
	);
	LUT3 #(
		.INIT('hd0)
	) name4431 (
		_w710_,
		_w4881_,
		_w4883_,
		_w4884_
	);
	LUT3 #(
		.INIT('h2f)
	) name4432 (
		_w695_,
		_w4880_,
		_w4884_,
		_w4885_
	);
	LUT3 #(
		.INIT('h60)
	) name4433 (
		\Datai[25]_pad ,
		_w2208_,
		_w2215_,
		_w4886_
	);
	LUT2 #(
		.INIT('h8)
	) name4434 (
		_w2219_,
		_w4805_,
		_w4887_
	);
	LUT4 #(
		.INIT('h5553)
	) name4435 (
		\Datai[1]_pad ,
		\InstQueue_reg[1][1]/NET0131 ,
		_w2217_,
		_w2313_,
		_w4888_
	);
	LUT2 #(
		.INIT('h1)
	) name4436 (
		_w2316_,
		_w4888_,
		_w4889_
	);
	LUT4 #(
		.INIT('h0057)
	) name4437 (
		\DataWidth_reg[1]/NET0131 ,
		_w4886_,
		_w4887_,
		_w4889_,
		_w4890_
	);
	LUT4 #(
		.INIT('hc055)
	) name4438 (
		\InstQueue_reg[1][1]/NET0131 ,
		_w488_,
		_w493_,
		_w2313_,
		_w4891_
	);
	LUT2 #(
		.INIT('h2)
	) name4439 (
		\InstQueue_reg[1][1]/NET0131 ,
		_w2227_,
		_w4892_
	);
	LUT3 #(
		.INIT('h0d)
	) name4440 (
		_w1212_,
		_w4888_,
		_w4892_,
		_w4893_
	);
	LUT3 #(
		.INIT('hd0)
	) name4441 (
		_w710_,
		_w4891_,
		_w4893_,
		_w4894_
	);
	LUT3 #(
		.INIT('h2f)
	) name4442 (
		_w695_,
		_w4890_,
		_w4894_,
		_w4895_
	);
	LUT2 #(
		.INIT('h8)
	) name4443 (
		_w2217_,
		_w4805_,
		_w4896_
	);
	LUT3 #(
		.INIT('h48)
	) name4444 (
		\Datai[25]_pad ,
		_w2219_,
		_w2208_,
		_w4897_
	);
	LUT4 #(
		.INIT('h5553)
	) name4445 (
		\Datai[1]_pad ,
		\InstQueue_reg[2][1]/NET0131 ,
		_w2313_,
		_w2326_,
		_w4898_
	);
	LUT2 #(
		.INIT('h1)
	) name4446 (
		_w2329_,
		_w4898_,
		_w4899_
	);
	LUT4 #(
		.INIT('h0057)
	) name4447 (
		\DataWidth_reg[1]/NET0131 ,
		_w4896_,
		_w4897_,
		_w4899_,
		_w4900_
	);
	LUT4 #(
		.INIT('hc055)
	) name4448 (
		\InstQueue_reg[2][1]/NET0131 ,
		_w488_,
		_w493_,
		_w2326_,
		_w4901_
	);
	LUT2 #(
		.INIT('h2)
	) name4449 (
		\InstQueue_reg[2][1]/NET0131 ,
		_w2227_,
		_w4902_
	);
	LUT3 #(
		.INIT('h0d)
	) name4450 (
		_w1212_,
		_w4898_,
		_w4902_,
		_w4903_
	);
	LUT3 #(
		.INIT('hd0)
	) name4451 (
		_w710_,
		_w4901_,
		_w4903_,
		_w4904_
	);
	LUT3 #(
		.INIT('h2f)
	) name4452 (
		_w695_,
		_w4900_,
		_w4904_,
		_w4905_
	);
	LUT4 #(
		.INIT('ha600)
	) name4453 (
		\Datai[16]_pad ,
		\Datai[31]_pad ,
		_w2204_,
		_w2313_,
		_w4906_
	);
	LUT4 #(
		.INIT('haa80)
	) name4454 (
		\DataWidth_reg[1]/NET0131 ,
		_w2217_,
		_w4825_,
		_w4906_,
		_w4907_
	);
	LUT4 #(
		.INIT('h5553)
	) name4455 (
		\Datai[0]_pad ,
		\InstQueue_reg[3][0]/NET0131 ,
		_w2326_,
		_w2339_,
		_w4908_
	);
	LUT2 #(
		.INIT('h1)
	) name4456 (
		_w2342_,
		_w4908_,
		_w4909_
	);
	LUT3 #(
		.INIT('ha8)
	) name4457 (
		_w695_,
		_w4907_,
		_w4909_,
		_w4910_
	);
	LUT4 #(
		.INIT('hc055)
	) name4458 (
		\InstQueue_reg[3][0]/NET0131 ,
		_w500_,
		_w506_,
		_w2339_,
		_w4911_
	);
	LUT2 #(
		.INIT('h2)
	) name4459 (
		\InstQueue_reg[3][0]/NET0131 ,
		_w2227_,
		_w4912_
	);
	LUT3 #(
		.INIT('h0d)
	) name4460 (
		_w1212_,
		_w4908_,
		_w4912_,
		_w4913_
	);
	LUT3 #(
		.INIT('hd0)
	) name4461 (
		_w710_,
		_w4911_,
		_w4913_,
		_w4914_
	);
	LUT2 #(
		.INIT('hb)
	) name4462 (
		_w4910_,
		_w4914_,
		_w4915_
	);
	LUT3 #(
		.INIT('h48)
	) name4463 (
		\Datai[25]_pad ,
		_w2217_,
		_w2208_,
		_w4916_
	);
	LUT2 #(
		.INIT('h8)
	) name4464 (
		_w2313_,
		_w4805_,
		_w4917_
	);
	LUT4 #(
		.INIT('h5553)
	) name4465 (
		\Datai[1]_pad ,
		\InstQueue_reg[3][1]/NET0131 ,
		_w2326_,
		_w2339_,
		_w4918_
	);
	LUT2 #(
		.INIT('h1)
	) name4466 (
		_w2342_,
		_w4918_,
		_w4919_
	);
	LUT4 #(
		.INIT('h0057)
	) name4467 (
		\DataWidth_reg[1]/NET0131 ,
		_w4916_,
		_w4917_,
		_w4919_,
		_w4920_
	);
	LUT4 #(
		.INIT('hc055)
	) name4468 (
		\InstQueue_reg[3][1]/NET0131 ,
		_w488_,
		_w493_,
		_w2339_,
		_w4921_
	);
	LUT2 #(
		.INIT('h2)
	) name4469 (
		\InstQueue_reg[3][1]/NET0131 ,
		_w2227_,
		_w4922_
	);
	LUT3 #(
		.INIT('h0d)
	) name4470 (
		_w1212_,
		_w4918_,
		_w4922_,
		_w4923_
	);
	LUT3 #(
		.INIT('hd0)
	) name4471 (
		_w710_,
		_w4921_,
		_w4923_,
		_w4924_
	);
	LUT3 #(
		.INIT('h2f)
	) name4472 (
		_w695_,
		_w4920_,
		_w4924_,
		_w4925_
	);
	LUT3 #(
		.INIT('h60)
	) name4473 (
		\Datai[25]_pad ,
		_w2208_,
		_w2313_,
		_w4926_
	);
	LUT2 #(
		.INIT('h8)
	) name4474 (
		_w2326_,
		_w4805_,
		_w4927_
	);
	LUT4 #(
		.INIT('h5553)
	) name4475 (
		\Datai[1]_pad ,
		\InstQueue_reg[4][1]/NET0131 ,
		_w2339_,
		_w2352_,
		_w4928_
	);
	LUT2 #(
		.INIT('h1)
	) name4476 (
		_w2355_,
		_w4928_,
		_w4929_
	);
	LUT4 #(
		.INIT('h0057)
	) name4477 (
		\DataWidth_reg[1]/NET0131 ,
		_w4926_,
		_w4927_,
		_w4929_,
		_w4930_
	);
	LUT4 #(
		.INIT('hc055)
	) name4478 (
		\InstQueue_reg[4][1]/NET0131 ,
		_w488_,
		_w493_,
		_w2352_,
		_w4931_
	);
	LUT2 #(
		.INIT('h2)
	) name4479 (
		\InstQueue_reg[4][1]/NET0131 ,
		_w2227_,
		_w4932_
	);
	LUT3 #(
		.INIT('h0d)
	) name4480 (
		_w1212_,
		_w4928_,
		_w4932_,
		_w4933_
	);
	LUT3 #(
		.INIT('hd0)
	) name4481 (
		_w710_,
		_w4931_,
		_w4933_,
		_w4934_
	);
	LUT3 #(
		.INIT('h2f)
	) name4482 (
		_w695_,
		_w4930_,
		_w4934_,
		_w4935_
	);
	LUT3 #(
		.INIT('h60)
	) name4483 (
		\Datai[25]_pad ,
		_w2208_,
		_w2326_,
		_w4936_
	);
	LUT2 #(
		.INIT('h8)
	) name4484 (
		_w2339_,
		_w4805_,
		_w4937_
	);
	LUT4 #(
		.INIT('h5553)
	) name4485 (
		\Datai[1]_pad ,
		\InstQueue_reg[5][1]/NET0131 ,
		_w2352_,
		_w2365_,
		_w4938_
	);
	LUT2 #(
		.INIT('h1)
	) name4486 (
		_w2368_,
		_w4938_,
		_w4939_
	);
	LUT4 #(
		.INIT('h0057)
	) name4487 (
		\DataWidth_reg[1]/NET0131 ,
		_w4936_,
		_w4937_,
		_w4939_,
		_w4940_
	);
	LUT4 #(
		.INIT('hc055)
	) name4488 (
		\InstQueue_reg[5][1]/NET0131 ,
		_w488_,
		_w493_,
		_w2365_,
		_w4941_
	);
	LUT2 #(
		.INIT('h2)
	) name4489 (
		\InstQueue_reg[5][1]/NET0131 ,
		_w2227_,
		_w4942_
	);
	LUT3 #(
		.INIT('h0d)
	) name4490 (
		_w1212_,
		_w4938_,
		_w4942_,
		_w4943_
	);
	LUT3 #(
		.INIT('hd0)
	) name4491 (
		_w710_,
		_w4941_,
		_w4943_,
		_w4944_
	);
	LUT3 #(
		.INIT('h2f)
	) name4492 (
		_w695_,
		_w4940_,
		_w4944_,
		_w4945_
	);
	LUT3 #(
		.INIT('h60)
	) name4493 (
		\Datai[25]_pad ,
		_w2208_,
		_w2339_,
		_w4946_
	);
	LUT2 #(
		.INIT('h8)
	) name4494 (
		_w2352_,
		_w4805_,
		_w4947_
	);
	LUT4 #(
		.INIT('h5553)
	) name4495 (
		\Datai[1]_pad ,
		\InstQueue_reg[6][1]/NET0131 ,
		_w2365_,
		_w2378_,
		_w4948_
	);
	LUT2 #(
		.INIT('h1)
	) name4496 (
		_w2381_,
		_w4948_,
		_w4949_
	);
	LUT4 #(
		.INIT('h0057)
	) name4497 (
		\DataWidth_reg[1]/NET0131 ,
		_w4946_,
		_w4947_,
		_w4949_,
		_w4950_
	);
	LUT4 #(
		.INIT('hc055)
	) name4498 (
		\InstQueue_reg[6][1]/NET0131 ,
		_w488_,
		_w493_,
		_w2378_,
		_w4951_
	);
	LUT2 #(
		.INIT('h2)
	) name4499 (
		\InstQueue_reg[6][1]/NET0131 ,
		_w2227_,
		_w4952_
	);
	LUT3 #(
		.INIT('h0d)
	) name4500 (
		_w1212_,
		_w4948_,
		_w4952_,
		_w4953_
	);
	LUT3 #(
		.INIT('hd0)
	) name4501 (
		_w710_,
		_w4951_,
		_w4953_,
		_w4954_
	);
	LUT3 #(
		.INIT('h2f)
	) name4502 (
		_w695_,
		_w4950_,
		_w4954_,
		_w4955_
	);
	LUT4 #(
		.INIT('ha600)
	) name4503 (
		\Datai[16]_pad ,
		\Datai[31]_pad ,
		_w2204_,
		_w2365_,
		_w4956_
	);
	LUT4 #(
		.INIT('haa80)
	) name4504 (
		\DataWidth_reg[1]/NET0131 ,
		_w2352_,
		_w4825_,
		_w4956_,
		_w4957_
	);
	LUT4 #(
		.INIT('h5553)
	) name4505 (
		\Datai[0]_pad ,
		\InstQueue_reg[7][0]/NET0131 ,
		_w2232_,
		_w2378_,
		_w4958_
	);
	LUT2 #(
		.INIT('h1)
	) name4506 (
		_w2393_,
		_w4958_,
		_w4959_
	);
	LUT3 #(
		.INIT('ha8)
	) name4507 (
		_w695_,
		_w4957_,
		_w4959_,
		_w4960_
	);
	LUT4 #(
		.INIT('hc055)
	) name4508 (
		\InstQueue_reg[7][0]/NET0131 ,
		_w500_,
		_w506_,
		_w2232_,
		_w4961_
	);
	LUT2 #(
		.INIT('h2)
	) name4509 (
		\InstQueue_reg[7][0]/NET0131 ,
		_w2227_,
		_w4962_
	);
	LUT3 #(
		.INIT('h0d)
	) name4510 (
		_w1212_,
		_w4958_,
		_w4962_,
		_w4963_
	);
	LUT3 #(
		.INIT('hd0)
	) name4511 (
		_w710_,
		_w4961_,
		_w4963_,
		_w4964_
	);
	LUT2 #(
		.INIT('hb)
	) name4512 (
		_w4960_,
		_w4964_,
		_w4965_
	);
	LUT3 #(
		.INIT('h60)
	) name4513 (
		\Datai[25]_pad ,
		_w2208_,
		_w2352_,
		_w4966_
	);
	LUT2 #(
		.INIT('h8)
	) name4514 (
		_w2365_,
		_w4805_,
		_w4967_
	);
	LUT4 #(
		.INIT('h5553)
	) name4515 (
		\Datai[1]_pad ,
		\InstQueue_reg[7][1]/NET0131 ,
		_w2232_,
		_w2378_,
		_w4968_
	);
	LUT2 #(
		.INIT('h1)
	) name4516 (
		_w2393_,
		_w4968_,
		_w4969_
	);
	LUT4 #(
		.INIT('h0057)
	) name4517 (
		\DataWidth_reg[1]/NET0131 ,
		_w4966_,
		_w4967_,
		_w4969_,
		_w4970_
	);
	LUT4 #(
		.INIT('hc055)
	) name4518 (
		\InstQueue_reg[7][1]/NET0131 ,
		_w488_,
		_w493_,
		_w2232_,
		_w4971_
	);
	LUT2 #(
		.INIT('h2)
	) name4519 (
		\InstQueue_reg[7][1]/NET0131 ,
		_w2227_,
		_w4972_
	);
	LUT3 #(
		.INIT('h0d)
	) name4520 (
		_w1212_,
		_w4968_,
		_w4972_,
		_w4973_
	);
	LUT3 #(
		.INIT('hd0)
	) name4521 (
		_w710_,
		_w4971_,
		_w4973_,
		_w4974_
	);
	LUT3 #(
		.INIT('h2f)
	) name4522 (
		_w695_,
		_w4970_,
		_w4974_,
		_w4975_
	);
	LUT3 #(
		.INIT('h60)
	) name4523 (
		\Datai[25]_pad ,
		_w2208_,
		_w2365_,
		_w4976_
	);
	LUT2 #(
		.INIT('h8)
	) name4524 (
		_w2378_,
		_w4805_,
		_w4977_
	);
	LUT4 #(
		.INIT('h5553)
	) name4525 (
		\Datai[1]_pad ,
		\InstQueue_reg[8][1]/NET0131 ,
		_w2232_,
		_w2234_,
		_w4978_
	);
	LUT2 #(
		.INIT('h1)
	) name4526 (
		_w2404_,
		_w4978_,
		_w4979_
	);
	LUT4 #(
		.INIT('h0057)
	) name4527 (
		\DataWidth_reg[1]/NET0131 ,
		_w4976_,
		_w4977_,
		_w4979_,
		_w4980_
	);
	LUT4 #(
		.INIT('hc055)
	) name4528 (
		\InstQueue_reg[8][1]/NET0131 ,
		_w488_,
		_w493_,
		_w2234_,
		_w4981_
	);
	LUT2 #(
		.INIT('h2)
	) name4529 (
		\InstQueue_reg[8][1]/NET0131 ,
		_w2227_,
		_w4982_
	);
	LUT3 #(
		.INIT('h0d)
	) name4530 (
		_w1212_,
		_w4978_,
		_w4982_,
		_w4983_
	);
	LUT3 #(
		.INIT('hd0)
	) name4531 (
		_w710_,
		_w4981_,
		_w4983_,
		_w4984_
	);
	LUT3 #(
		.INIT('h2f)
	) name4532 (
		_w695_,
		_w4980_,
		_w4984_,
		_w4985_
	);
	LUT3 #(
		.INIT('h60)
	) name4533 (
		\Datai[25]_pad ,
		_w2208_,
		_w2378_,
		_w4986_
	);
	LUT2 #(
		.INIT('h8)
	) name4534 (
		_w2232_,
		_w4805_,
		_w4987_
	);
	LUT4 #(
		.INIT('h5553)
	) name4535 (
		\Datai[1]_pad ,
		\InstQueue_reg[9][1]/NET0131 ,
		_w2237_,
		_w2234_,
		_w4988_
	);
	LUT2 #(
		.INIT('h1)
	) name4536 (
		_w2415_,
		_w4988_,
		_w4989_
	);
	LUT4 #(
		.INIT('h0057)
	) name4537 (
		\DataWidth_reg[1]/NET0131 ,
		_w4986_,
		_w4987_,
		_w4989_,
		_w4990_
	);
	LUT4 #(
		.INIT('hc055)
	) name4538 (
		\InstQueue_reg[9][1]/NET0131 ,
		_w488_,
		_w493_,
		_w2237_,
		_w4991_
	);
	LUT2 #(
		.INIT('h2)
	) name4539 (
		\InstQueue_reg[9][1]/NET0131 ,
		_w2227_,
		_w4992_
	);
	LUT3 #(
		.INIT('h0d)
	) name4540 (
		_w1212_,
		_w4988_,
		_w4992_,
		_w4993_
	);
	LUT3 #(
		.INIT('hd0)
	) name4541 (
		_w710_,
		_w4991_,
		_w4993_,
		_w4994_
	);
	LUT3 #(
		.INIT('h2f)
	) name4542 (
		_w695_,
		_w4990_,
		_w4994_,
		_w4995_
	);
	LUT4 #(
		.INIT('h4888)
	) name4543 (
		\rEIP_reg[26]/NET0131 ,
		_w592_,
		_w3249_,
		_w4685_,
		_w4996_
	);
	LUT3 #(
		.INIT('h8a)
	) name4544 (
		\Address[24]_pad ,
		\State_reg[0]/NET0131 ,
		\State_reg[1]/NET0131 ,
		_w4997_
	);
	LUT3 #(
		.INIT('h13)
	) name4545 (
		\rEIP_reg[24]/NET0131 ,
		\rEIP_reg[25]/NET0131 ,
		_w4692_,
		_w4998_
	);
	LUT3 #(
		.INIT('h4c)
	) name4546 (
		_w3250_,
		_w4695_,
		_w4691_,
		_w4999_
	);
	LUT3 #(
		.INIT('h45)
	) name4547 (
		_w4997_,
		_w4998_,
		_w4999_,
		_w5000_
	);
	LUT2 #(
		.INIT('hb)
	) name4548 (
		_w4996_,
		_w5000_,
		_w5001_
	);
	LUT4 #(
		.INIT('h4888)
	) name4549 (
		\rEIP_reg[14]/NET0131 ,
		_w592_,
		_w3151_,
		_w4681_,
		_w5002_
	);
	LUT3 #(
		.INIT('h8a)
	) name4550 (
		\Address[12]_pad ,
		\State_reg[0]/NET0131 ,
		\State_reg[1]/NET0131 ,
		_w5003_
	);
	LUT3 #(
		.INIT('h13)
	) name4551 (
		\rEIP_reg[0]/NET0131 ,
		\rEIP_reg[13]/NET0131 ,
		\rEIP_reg[31]/NET0131 ,
		_w5004_
	);
	LUT2 #(
		.INIT('h2)
	) name4552 (
		_w4695_,
		_w5004_,
		_w5005_
	);
	LUT4 #(
		.INIT('h040f)
	) name4553 (
		_w3552_,
		_w4691_,
		_w5003_,
		_w5005_,
		_w5006_
	);
	LUT2 #(
		.INIT('hb)
	) name4554 (
		_w5002_,
		_w5006_,
		_w5007_
	);
	LUT4 #(
		.INIT('h8000)
	) name4555 (
		\rEIP_reg[16]/NET0131 ,
		_w3156_,
		_w3157_,
		_w4683_,
		_w5008_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name4556 (
		\rEIP_reg[16]/NET0131 ,
		_w592_,
		_w3196_,
		_w4683_,
		_w5009_
	);
	LUT4 #(
		.INIT('hec00)
	) name4557 (
		\rEIP_reg[21]/NET0131 ,
		\rEIP_reg[22]/NET0131 ,
		_w5008_,
		_w5009_,
		_w5010_
	);
	LUT3 #(
		.INIT('h8a)
	) name4558 (
		\Address[20]_pad ,
		\State_reg[0]/NET0131 ,
		\State_reg[1]/NET0131 ,
		_w5011_
	);
	LUT4 #(
		.INIT('h8000)
	) name4559 (
		_w3155_,
		_w3156_,
		_w3157_,
		_w4691_,
		_w5012_
	);
	LUT4 #(
		.INIT('h0b07)
	) name4560 (
		\rEIP_reg[21]/NET0131 ,
		_w4695_,
		_w5011_,
		_w5012_,
		_w5013_
	);
	LUT2 #(
		.INIT('hb)
	) name4561 (
		_w5010_,
		_w5013_,
		_w5014_
	);
	LUT4 #(
		.INIT('h60a0)
	) name4562 (
		\rEIP_reg[10]/NET0131 ,
		\rEIP_reg[9]/NET0131 ,
		_w592_,
		_w4679_,
		_w5015_
	);
	LUT3 #(
		.INIT('h8a)
	) name4563 (
		\Address[8]_pad ,
		\State_reg[0]/NET0131 ,
		\State_reg[1]/NET0131 ,
		_w5016_
	);
	LUT4 #(
		.INIT('h9300)
	) name4564 (
		\rEIP_reg[8]/NET0131 ,
		\rEIP_reg[9]/NET0131 ,
		_w3149_,
		_w4691_,
		_w5017_
	);
	LUT3 #(
		.INIT('h07)
	) name4565 (
		\rEIP_reg[0]/NET0131 ,
		\rEIP_reg[31]/NET0131 ,
		\rEIP_reg[9]/NET0131 ,
		_w5018_
	);
	LUT2 #(
		.INIT('h2)
	) name4566 (
		_w4695_,
		_w5018_,
		_w5019_
	);
	LUT3 #(
		.INIT('h45)
	) name4567 (
		_w5016_,
		_w5017_,
		_w5019_,
		_w5020_
	);
	LUT2 #(
		.INIT('hb)
	) name4568 (
		_w5015_,
		_w5020_,
		_w5021_
	);
	LUT4 #(
		.INIT('ha600)
	) name4569 (
		\Datai[16]_pad ,
		\Datai[31]_pad ,
		_w2204_,
		_w2215_,
		_w5022_
	);
	LUT4 #(
		.INIT('haa80)
	) name4570 (
		\DataWidth_reg[1]/NET0131 ,
		_w2199_,
		_w4825_,
		_w5022_,
		_w5023_
	);
	LUT4 #(
		.INIT('h5553)
	) name4571 (
		\Datai[0]_pad ,
		\InstQueue_reg[0][0]/NET0131 ,
		_w2217_,
		_w2219_,
		_w5024_
	);
	LUT2 #(
		.INIT('h1)
	) name4572 (
		_w2223_,
		_w5024_,
		_w5025_
	);
	LUT3 #(
		.INIT('ha8)
	) name4573 (
		_w695_,
		_w5023_,
		_w5025_,
		_w5026_
	);
	LUT4 #(
		.INIT('hc055)
	) name4574 (
		\InstQueue_reg[0][0]/NET0131 ,
		_w500_,
		_w506_,
		_w2217_,
		_w5027_
	);
	LUT2 #(
		.INIT('h2)
	) name4575 (
		\InstQueue_reg[0][0]/NET0131 ,
		_w2227_,
		_w5028_
	);
	LUT3 #(
		.INIT('h0d)
	) name4576 (
		_w1212_,
		_w5024_,
		_w5028_,
		_w5029_
	);
	LUT3 #(
		.INIT('hd0)
	) name4577 (
		_w710_,
		_w5027_,
		_w5029_,
		_w5030_
	);
	LUT2 #(
		.INIT('hb)
	) name4578 (
		_w5026_,
		_w5030_,
		_w5031_
	);
	LUT4 #(
		.INIT('ha600)
	) name4579 (
		\Datai[16]_pad ,
		\Datai[31]_pad ,
		_w2204_,
		_w2234_,
		_w5032_
	);
	LUT4 #(
		.INIT('haa80)
	) name4580 (
		\DataWidth_reg[1]/NET0131 ,
		_w2232_,
		_w4825_,
		_w5032_,
		_w5033_
	);
	LUT4 #(
		.INIT('h5553)
	) name4581 (
		\Datai[0]_pad ,
		\InstQueue_reg[10][0]/NET0131 ,
		_w2236_,
		_w2237_,
		_w5034_
	);
	LUT2 #(
		.INIT('h1)
	) name4582 (
		_w2241_,
		_w5034_,
		_w5035_
	);
	LUT3 #(
		.INIT('ha8)
	) name4583 (
		_w695_,
		_w5033_,
		_w5035_,
		_w5036_
	);
	LUT4 #(
		.INIT('hc055)
	) name4584 (
		\InstQueue_reg[10][0]/NET0131 ,
		_w500_,
		_w506_,
		_w2236_,
		_w5037_
	);
	LUT2 #(
		.INIT('h2)
	) name4585 (
		\InstQueue_reg[10][0]/NET0131 ,
		_w2227_,
		_w5038_
	);
	LUT3 #(
		.INIT('h0d)
	) name4586 (
		_w1212_,
		_w5034_,
		_w5038_,
		_w5039_
	);
	LUT3 #(
		.INIT('hd0)
	) name4587 (
		_w710_,
		_w5037_,
		_w5039_,
		_w5040_
	);
	LUT2 #(
		.INIT('hb)
	) name4588 (
		_w5036_,
		_w5040_,
		_w5041_
	);
	LUT4 #(
		.INIT('ha600)
	) name4589 (
		\Datai[16]_pad ,
		\Datai[31]_pad ,
		_w2204_,
		_w2236_,
		_w5042_
	);
	LUT4 #(
		.INIT('haa80)
	) name4590 (
		\DataWidth_reg[1]/NET0131 ,
		_w2237_,
		_w4825_,
		_w5042_,
		_w5043_
	);
	LUT4 #(
		.INIT('h5553)
	) name4591 (
		\Datai[0]_pad ,
		\InstQueue_reg[12][0]/NET0131 ,
		_w2251_,
		_w2265_,
		_w5044_
	);
	LUT2 #(
		.INIT('h1)
	) name4592 (
		_w2268_,
		_w5044_,
		_w5045_
	);
	LUT3 #(
		.INIT('ha8)
	) name4593 (
		_w695_,
		_w5043_,
		_w5045_,
		_w5046_
	);
	LUT4 #(
		.INIT('hc055)
	) name4594 (
		\InstQueue_reg[12][0]/NET0131 ,
		_w500_,
		_w506_,
		_w2265_,
		_w5047_
	);
	LUT2 #(
		.INIT('h2)
	) name4595 (
		\InstQueue_reg[12][0]/NET0131 ,
		_w2227_,
		_w5048_
	);
	LUT3 #(
		.INIT('h0d)
	) name4596 (
		_w1212_,
		_w5044_,
		_w5048_,
		_w5049_
	);
	LUT3 #(
		.INIT('hd0)
	) name4597 (
		_w710_,
		_w5047_,
		_w5049_,
		_w5050_
	);
	LUT2 #(
		.INIT('hb)
	) name4598 (
		_w5046_,
		_w5050_,
		_w5051_
	);
	LUT4 #(
		.INIT('ha600)
	) name4599 (
		\Datai[16]_pad ,
		\Datai[31]_pad ,
		_w2204_,
		_w2251_,
		_w5052_
	);
	LUT4 #(
		.INIT('haa80)
	) name4600 (
		\DataWidth_reg[1]/NET0131 ,
		_w2236_,
		_w4825_,
		_w5052_,
		_w5053_
	);
	LUT4 #(
		.INIT('h5553)
	) name4601 (
		\Datai[0]_pad ,
		\InstQueue_reg[13][0]/NET0131 ,
		_w2199_,
		_w2265_,
		_w5054_
	);
	LUT2 #(
		.INIT('h1)
	) name4602 (
		_w2280_,
		_w5054_,
		_w5055_
	);
	LUT3 #(
		.INIT('ha8)
	) name4603 (
		_w695_,
		_w5053_,
		_w5055_,
		_w5056_
	);
	LUT4 #(
		.INIT('hc055)
	) name4604 (
		\InstQueue_reg[13][0]/NET0131 ,
		_w500_,
		_w506_,
		_w2199_,
		_w5057_
	);
	LUT2 #(
		.INIT('h2)
	) name4605 (
		\InstQueue_reg[13][0]/NET0131 ,
		_w2227_,
		_w5058_
	);
	LUT3 #(
		.INIT('h0d)
	) name4606 (
		_w1212_,
		_w5054_,
		_w5058_,
		_w5059_
	);
	LUT3 #(
		.INIT('hd0)
	) name4607 (
		_w710_,
		_w5057_,
		_w5059_,
		_w5060_
	);
	LUT2 #(
		.INIT('hb)
	) name4608 (
		_w5056_,
		_w5060_,
		_w5061_
	);
	LUT4 #(
		.INIT('ha600)
	) name4609 (
		\Datai[16]_pad ,
		\Datai[31]_pad ,
		_w2204_,
		_w2265_,
		_w5062_
	);
	LUT4 #(
		.INIT('haa80)
	) name4610 (
		\DataWidth_reg[1]/NET0131 ,
		_w2251_,
		_w4825_,
		_w5062_,
		_w5063_
	);
	LUT4 #(
		.INIT('h5553)
	) name4611 (
		\Datai[0]_pad ,
		\InstQueue_reg[14][0]/NET0131 ,
		_w2199_,
		_w2215_,
		_w5064_
	);
	LUT2 #(
		.INIT('h1)
	) name4612 (
		_w2291_,
		_w5064_,
		_w5065_
	);
	LUT3 #(
		.INIT('ha8)
	) name4613 (
		_w695_,
		_w5063_,
		_w5065_,
		_w5066_
	);
	LUT4 #(
		.INIT('hc055)
	) name4614 (
		\InstQueue_reg[14][0]/NET0131 ,
		_w500_,
		_w506_,
		_w2215_,
		_w5067_
	);
	LUT2 #(
		.INIT('h2)
	) name4615 (
		\InstQueue_reg[14][0]/NET0131 ,
		_w2227_,
		_w5068_
	);
	LUT3 #(
		.INIT('h0d)
	) name4616 (
		_w1212_,
		_w5064_,
		_w5068_,
		_w5069_
	);
	LUT3 #(
		.INIT('hd0)
	) name4617 (
		_w710_,
		_w5067_,
		_w5069_,
		_w5070_
	);
	LUT2 #(
		.INIT('hb)
	) name4618 (
		_w5066_,
		_w5070_,
		_w5071_
	);
	LUT4 #(
		.INIT('ha060)
	) name4619 (
		\Datai[16]_pad ,
		\Datai[31]_pad ,
		_w2199_,
		_w2204_,
		_w5072_
	);
	LUT4 #(
		.INIT('haa80)
	) name4620 (
		\DataWidth_reg[1]/NET0131 ,
		_w2265_,
		_w4825_,
		_w5072_,
		_w5073_
	);
	LUT4 #(
		.INIT('h5553)
	) name4621 (
		\Datai[0]_pad ,
		\InstQueue_reg[15][0]/NET0131 ,
		_w2219_,
		_w2215_,
		_w5074_
	);
	LUT2 #(
		.INIT('h1)
	) name4622 (
		_w2303_,
		_w5074_,
		_w5075_
	);
	LUT3 #(
		.INIT('ha8)
	) name4623 (
		_w695_,
		_w5073_,
		_w5075_,
		_w5076_
	);
	LUT4 #(
		.INIT('hc055)
	) name4624 (
		\InstQueue_reg[15][0]/NET0131 ,
		_w500_,
		_w506_,
		_w2219_,
		_w5077_
	);
	LUT2 #(
		.INIT('h2)
	) name4625 (
		\InstQueue_reg[15][0]/NET0131 ,
		_w2227_,
		_w5078_
	);
	LUT3 #(
		.INIT('h0d)
	) name4626 (
		_w1212_,
		_w5074_,
		_w5078_,
		_w5079_
	);
	LUT3 #(
		.INIT('hd0)
	) name4627 (
		_w710_,
		_w5077_,
		_w5079_,
		_w5080_
	);
	LUT2 #(
		.INIT('hb)
	) name4628 (
		_w5076_,
		_w5080_,
		_w5081_
	);
	LUT4 #(
		.INIT('ha060)
	) name4629 (
		\Datai[16]_pad ,
		\Datai[31]_pad ,
		_w2219_,
		_w2204_,
		_w5082_
	);
	LUT4 #(
		.INIT('haa80)
	) name4630 (
		\DataWidth_reg[1]/NET0131 ,
		_w2215_,
		_w4825_,
		_w5082_,
		_w5083_
	);
	LUT4 #(
		.INIT('h5553)
	) name4631 (
		\Datai[0]_pad ,
		\InstQueue_reg[1][0]/NET0131 ,
		_w2217_,
		_w2313_,
		_w5084_
	);
	LUT2 #(
		.INIT('h1)
	) name4632 (
		_w2316_,
		_w5084_,
		_w5085_
	);
	LUT3 #(
		.INIT('ha8)
	) name4633 (
		_w695_,
		_w5083_,
		_w5085_,
		_w5086_
	);
	LUT4 #(
		.INIT('hc055)
	) name4634 (
		\InstQueue_reg[1][0]/NET0131 ,
		_w500_,
		_w506_,
		_w2313_,
		_w5087_
	);
	LUT2 #(
		.INIT('h2)
	) name4635 (
		\InstQueue_reg[1][0]/NET0131 ,
		_w2227_,
		_w5088_
	);
	LUT3 #(
		.INIT('h0d)
	) name4636 (
		_w1212_,
		_w5084_,
		_w5088_,
		_w5089_
	);
	LUT3 #(
		.INIT('hd0)
	) name4637 (
		_w710_,
		_w5087_,
		_w5089_,
		_w5090_
	);
	LUT2 #(
		.INIT('hb)
	) name4638 (
		_w5086_,
		_w5090_,
		_w5091_
	);
	LUT4 #(
		.INIT('ha060)
	) name4639 (
		\Datai[16]_pad ,
		\Datai[31]_pad ,
		_w2217_,
		_w2204_,
		_w5092_
	);
	LUT4 #(
		.INIT('haa80)
	) name4640 (
		\DataWidth_reg[1]/NET0131 ,
		_w2219_,
		_w4825_,
		_w5092_,
		_w5093_
	);
	LUT4 #(
		.INIT('h5553)
	) name4641 (
		\Datai[0]_pad ,
		\InstQueue_reg[2][0]/NET0131 ,
		_w2313_,
		_w2326_,
		_w5094_
	);
	LUT2 #(
		.INIT('h1)
	) name4642 (
		_w2329_,
		_w5094_,
		_w5095_
	);
	LUT3 #(
		.INIT('ha8)
	) name4643 (
		_w695_,
		_w5093_,
		_w5095_,
		_w5096_
	);
	LUT4 #(
		.INIT('hc055)
	) name4644 (
		\InstQueue_reg[2][0]/NET0131 ,
		_w500_,
		_w506_,
		_w2326_,
		_w5097_
	);
	LUT2 #(
		.INIT('h2)
	) name4645 (
		\InstQueue_reg[2][0]/NET0131 ,
		_w2227_,
		_w5098_
	);
	LUT3 #(
		.INIT('h0d)
	) name4646 (
		_w1212_,
		_w5094_,
		_w5098_,
		_w5099_
	);
	LUT3 #(
		.INIT('hd0)
	) name4647 (
		_w710_,
		_w5097_,
		_w5099_,
		_w5100_
	);
	LUT2 #(
		.INIT('hb)
	) name4648 (
		_w5096_,
		_w5100_,
		_w5101_
	);
	LUT4 #(
		.INIT('ha600)
	) name4649 (
		\Datai[16]_pad ,
		\Datai[31]_pad ,
		_w2204_,
		_w2326_,
		_w5102_
	);
	LUT4 #(
		.INIT('haa80)
	) name4650 (
		\DataWidth_reg[1]/NET0131 ,
		_w2313_,
		_w4825_,
		_w5102_,
		_w5103_
	);
	LUT4 #(
		.INIT('h5553)
	) name4651 (
		\Datai[0]_pad ,
		\InstQueue_reg[4][0]/NET0131 ,
		_w2339_,
		_w2352_,
		_w5104_
	);
	LUT2 #(
		.INIT('h1)
	) name4652 (
		_w2355_,
		_w5104_,
		_w5105_
	);
	LUT3 #(
		.INIT('ha8)
	) name4653 (
		_w695_,
		_w5103_,
		_w5105_,
		_w5106_
	);
	LUT4 #(
		.INIT('hc055)
	) name4654 (
		\InstQueue_reg[4][0]/NET0131 ,
		_w500_,
		_w506_,
		_w2352_,
		_w5107_
	);
	LUT2 #(
		.INIT('h2)
	) name4655 (
		\InstQueue_reg[4][0]/NET0131 ,
		_w2227_,
		_w5108_
	);
	LUT3 #(
		.INIT('h0d)
	) name4656 (
		_w1212_,
		_w5104_,
		_w5108_,
		_w5109_
	);
	LUT3 #(
		.INIT('hd0)
	) name4657 (
		_w710_,
		_w5107_,
		_w5109_,
		_w5110_
	);
	LUT2 #(
		.INIT('hb)
	) name4658 (
		_w5106_,
		_w5110_,
		_w5111_
	);
	LUT4 #(
		.INIT('ha600)
	) name4659 (
		\Datai[16]_pad ,
		\Datai[31]_pad ,
		_w2204_,
		_w2339_,
		_w5112_
	);
	LUT4 #(
		.INIT('haa80)
	) name4660 (
		\DataWidth_reg[1]/NET0131 ,
		_w2326_,
		_w4825_,
		_w5112_,
		_w5113_
	);
	LUT4 #(
		.INIT('h5553)
	) name4661 (
		\Datai[0]_pad ,
		\InstQueue_reg[5][0]/NET0131 ,
		_w2352_,
		_w2365_,
		_w5114_
	);
	LUT2 #(
		.INIT('h1)
	) name4662 (
		_w2368_,
		_w5114_,
		_w5115_
	);
	LUT3 #(
		.INIT('ha8)
	) name4663 (
		_w695_,
		_w5113_,
		_w5115_,
		_w5116_
	);
	LUT4 #(
		.INIT('hc055)
	) name4664 (
		\InstQueue_reg[5][0]/NET0131 ,
		_w500_,
		_w506_,
		_w2365_,
		_w5117_
	);
	LUT2 #(
		.INIT('h2)
	) name4665 (
		\InstQueue_reg[5][0]/NET0131 ,
		_w2227_,
		_w5118_
	);
	LUT3 #(
		.INIT('h0d)
	) name4666 (
		_w1212_,
		_w5114_,
		_w5118_,
		_w5119_
	);
	LUT3 #(
		.INIT('hd0)
	) name4667 (
		_w710_,
		_w5117_,
		_w5119_,
		_w5120_
	);
	LUT2 #(
		.INIT('hb)
	) name4668 (
		_w5116_,
		_w5120_,
		_w5121_
	);
	LUT4 #(
		.INIT('ha600)
	) name4669 (
		\Datai[16]_pad ,
		\Datai[31]_pad ,
		_w2204_,
		_w2352_,
		_w5122_
	);
	LUT4 #(
		.INIT('haa80)
	) name4670 (
		\DataWidth_reg[1]/NET0131 ,
		_w2339_,
		_w4825_,
		_w5122_,
		_w5123_
	);
	LUT4 #(
		.INIT('h5553)
	) name4671 (
		\Datai[0]_pad ,
		\InstQueue_reg[6][0]/NET0131 ,
		_w2365_,
		_w2378_,
		_w5124_
	);
	LUT2 #(
		.INIT('h1)
	) name4672 (
		_w2381_,
		_w5124_,
		_w5125_
	);
	LUT3 #(
		.INIT('ha8)
	) name4673 (
		_w695_,
		_w5123_,
		_w5125_,
		_w5126_
	);
	LUT4 #(
		.INIT('hc055)
	) name4674 (
		\InstQueue_reg[6][0]/NET0131 ,
		_w500_,
		_w506_,
		_w2378_,
		_w5127_
	);
	LUT2 #(
		.INIT('h2)
	) name4675 (
		\InstQueue_reg[6][0]/NET0131 ,
		_w2227_,
		_w5128_
	);
	LUT3 #(
		.INIT('h0d)
	) name4676 (
		_w1212_,
		_w5124_,
		_w5128_,
		_w5129_
	);
	LUT3 #(
		.INIT('hd0)
	) name4677 (
		_w710_,
		_w5127_,
		_w5129_,
		_w5130_
	);
	LUT2 #(
		.INIT('hb)
	) name4678 (
		_w5126_,
		_w5130_,
		_w5131_
	);
	LUT4 #(
		.INIT('ha600)
	) name4679 (
		\Datai[16]_pad ,
		\Datai[31]_pad ,
		_w2204_,
		_w2378_,
		_w5132_
	);
	LUT4 #(
		.INIT('haa80)
	) name4680 (
		\DataWidth_reg[1]/NET0131 ,
		_w2365_,
		_w4825_,
		_w5132_,
		_w5133_
	);
	LUT4 #(
		.INIT('h5553)
	) name4681 (
		\Datai[0]_pad ,
		\InstQueue_reg[8][0]/NET0131 ,
		_w2232_,
		_w2234_,
		_w5134_
	);
	LUT2 #(
		.INIT('h1)
	) name4682 (
		_w2404_,
		_w5134_,
		_w5135_
	);
	LUT3 #(
		.INIT('ha8)
	) name4683 (
		_w695_,
		_w5133_,
		_w5135_,
		_w5136_
	);
	LUT4 #(
		.INIT('hc055)
	) name4684 (
		\InstQueue_reg[8][0]/NET0131 ,
		_w500_,
		_w506_,
		_w2234_,
		_w5137_
	);
	LUT2 #(
		.INIT('h2)
	) name4685 (
		\InstQueue_reg[8][0]/NET0131 ,
		_w2227_,
		_w5138_
	);
	LUT3 #(
		.INIT('h0d)
	) name4686 (
		_w1212_,
		_w5134_,
		_w5138_,
		_w5139_
	);
	LUT3 #(
		.INIT('hd0)
	) name4687 (
		_w710_,
		_w5137_,
		_w5139_,
		_w5140_
	);
	LUT2 #(
		.INIT('hb)
	) name4688 (
		_w5136_,
		_w5140_,
		_w5141_
	);
	LUT4 #(
		.INIT('ha600)
	) name4689 (
		\Datai[16]_pad ,
		\Datai[31]_pad ,
		_w2204_,
		_w2232_,
		_w5142_
	);
	LUT4 #(
		.INIT('haa80)
	) name4690 (
		\DataWidth_reg[1]/NET0131 ,
		_w2378_,
		_w4825_,
		_w5142_,
		_w5143_
	);
	LUT4 #(
		.INIT('h5553)
	) name4691 (
		\Datai[0]_pad ,
		\InstQueue_reg[9][0]/NET0131 ,
		_w2237_,
		_w2234_,
		_w5144_
	);
	LUT2 #(
		.INIT('h1)
	) name4692 (
		_w2415_,
		_w5144_,
		_w5145_
	);
	LUT3 #(
		.INIT('ha8)
	) name4693 (
		_w695_,
		_w5143_,
		_w5145_,
		_w5146_
	);
	LUT4 #(
		.INIT('hc055)
	) name4694 (
		\InstQueue_reg[9][0]/NET0131 ,
		_w500_,
		_w506_,
		_w2237_,
		_w5147_
	);
	LUT2 #(
		.INIT('h2)
	) name4695 (
		\InstQueue_reg[9][0]/NET0131 ,
		_w2227_,
		_w5148_
	);
	LUT3 #(
		.INIT('h0d)
	) name4696 (
		_w1212_,
		_w5144_,
		_w5148_,
		_w5149_
	);
	LUT3 #(
		.INIT('hd0)
	) name4697 (
		_w710_,
		_w5147_,
		_w5149_,
		_w5150_
	);
	LUT2 #(
		.INIT('hb)
	) name4698 (
		_w5146_,
		_w5150_,
		_w5151_
	);
	LUT3 #(
		.INIT('h48)
	) name4699 (
		\rEIP_reg[6]/NET0131 ,
		_w592_,
		_w4677_,
		_w5152_
	);
	LUT3 #(
		.INIT('h8a)
	) name4700 (
		\Address[4]_pad ,
		\State_reg[0]/NET0131 ,
		\State_reg[1]/NET0131 ,
		_w5153_
	);
	LUT4 #(
		.INIT('h60a0)
	) name4701 (
		\rEIP_reg[5]/NET0131 ,
		_w3148_,
		_w4695_,
		_w4691_,
		_w5154_
	);
	LUT2 #(
		.INIT('h1)
	) name4702 (
		_w5153_,
		_w5154_,
		_w5155_
	);
	LUT2 #(
		.INIT('hb)
	) name4703 (
		_w5152_,
		_w5155_,
		_w5156_
	);
	LUT4 #(
		.INIT('h60c0)
	) name4704 (
		\rEIP_reg[28]/NET0131 ,
		\rEIP_reg[29]/NET0131 ,
		_w592_,
		_w4687_,
		_w5157_
	);
	LUT3 #(
		.INIT('h8a)
	) name4705 (
		\Address[27]_pad ,
		\State_reg[0]/NET0131 ,
		\State_reg[1]/NET0131 ,
		_w5158_
	);
	LUT4 #(
		.INIT('h00b7)
	) name4706 (
		\rEIP_reg[28]/NET0131 ,
		_w4695_,
		_w4693_,
		_w5158_,
		_w5159_
	);
	LUT2 #(
		.INIT('hb)
	) name4707 (
		_w5157_,
		_w5159_,
		_w5160_
	);
	LUT4 #(
		.INIT('h60c0)
	) name4708 (
		\rEIP_reg[16]/NET0131 ,
		\rEIP_reg[17]/NET0131 ,
		_w592_,
		_w4683_,
		_w5161_
	);
	LUT3 #(
		.INIT('h8a)
	) name4709 (
		\Address[15]_pad ,
		\State_reg[0]/NET0131 ,
		\State_reg[1]/NET0131 ,
		_w5162_
	);
	LUT4 #(
		.INIT('h8000)
	) name4710 (
		\rEIP_reg[11]/NET0131 ,
		_w3150_,
		_w3153_,
		_w4691_,
		_w5163_
	);
	LUT4 #(
		.INIT('h60a0)
	) name4711 (
		\rEIP_reg[16]/NET0131 ,
		_w3154_,
		_w4695_,
		_w4691_,
		_w5164_
	);
	LUT2 #(
		.INIT('h1)
	) name4712 (
		_w5162_,
		_w5164_,
		_w5165_
	);
	LUT2 #(
		.INIT('hb)
	) name4713 (
		_w5161_,
		_w5165_,
		_w5166_
	);
	LUT4 #(
		.INIT('h60c0)
	) name4714 (
		\rEIP_reg[24]/NET0131 ,
		\rEIP_reg[25]/NET0131 ,
		_w592_,
		_w4685_,
		_w5167_
	);
	LUT3 #(
		.INIT('h8a)
	) name4715 (
		\Address[23]_pad ,
		\State_reg[0]/NET0131 ,
		\State_reg[1]/NET0131 ,
		_w5168_
	);
	LUT4 #(
		.INIT('h00b7)
	) name4716 (
		\rEIP_reg[24]/NET0131 ,
		_w4695_,
		_w4692_,
		_w5168_,
		_w5169_
	);
	LUT2 #(
		.INIT('hb)
	) name4717 (
		_w5167_,
		_w5169_,
		_w5170_
	);
	LUT4 #(
		.INIT('h60c0)
	) name4718 (
		\rEIP_reg[12]/NET0131 ,
		\rEIP_reg[13]/NET0131 ,
		_w592_,
		_w4681_,
		_w5171_
	);
	LUT3 #(
		.INIT('h8a)
	) name4719 (
		\Address[11]_pad ,
		\State_reg[0]/NET0131 ,
		\State_reg[1]/NET0131 ,
		_w5172_
	);
	LUT4 #(
		.INIT('h9300)
	) name4720 (
		\rEIP_reg[11]/NET0131 ,
		\rEIP_reg[12]/NET0131 ,
		_w3150_,
		_w4691_,
		_w5173_
	);
	LUT3 #(
		.INIT('h13)
	) name4721 (
		\rEIP_reg[0]/NET0131 ,
		\rEIP_reg[12]/NET0131 ,
		\rEIP_reg[31]/NET0131 ,
		_w5174_
	);
	LUT2 #(
		.INIT('h2)
	) name4722 (
		_w4695_,
		_w5174_,
		_w5175_
	);
	LUT3 #(
		.INIT('h45)
	) name4723 (
		_w5172_,
		_w5173_,
		_w5175_,
		_w5176_
	);
	LUT2 #(
		.INIT('hb)
	) name4724 (
		_w5171_,
		_w5176_,
		_w5177_
	);
	LUT3 #(
		.INIT('h48)
	) name4725 (
		\rEIP_reg[5]/NET0131 ,
		_w592_,
		_w4676_,
		_w5178_
	);
	LUT3 #(
		.INIT('h8a)
	) name4726 (
		\Address[3]_pad ,
		\State_reg[0]/NET0131 ,
		\State_reg[1]/NET0131 ,
		_w5179_
	);
	LUT3 #(
		.INIT('h80)
	) name4727 (
		\rEIP_reg[0]/NET0131 ,
		\rEIP_reg[1]/NET0131 ,
		\rEIP_reg[31]/NET0131 ,
		_w5180_
	);
	LUT4 #(
		.INIT('h8000)
	) name4728 (
		\rEIP_reg[0]/NET0131 ,
		\rEIP_reg[1]/NET0131 ,
		\rEIP_reg[2]/NET0131 ,
		\rEIP_reg[31]/NET0131 ,
		_w5181_
	);
	LUT4 #(
		.INIT('h60c0)
	) name4729 (
		\rEIP_reg[3]/NET0131 ,
		\rEIP_reg[4]/NET0131 ,
		_w4695_,
		_w5181_,
		_w5182_
	);
	LUT2 #(
		.INIT('h1)
	) name4730 (
		_w5179_,
		_w5182_,
		_w5183_
	);
	LUT2 #(
		.INIT('hb)
	) name4731 (
		_w5178_,
		_w5183_,
		_w5184_
	);
	LUT3 #(
		.INIT('h48)
	) name4732 (
		\rEIP_reg[21]/NET0131 ,
		_w592_,
		_w5008_,
		_w5185_
	);
	LUT3 #(
		.INIT('h8a)
	) name4733 (
		\Address[19]_pad ,
		\State_reg[0]/NET0131 ,
		\State_reg[1]/NET0131 ,
		_w5186_
	);
	LUT4 #(
		.INIT('h8000)
	) name4734 (
		\rEIP_reg[19]/NET0131 ,
		_w3155_,
		_w3156_,
		_w4691_,
		_w5187_
	);
	LUT4 #(
		.INIT('h0c08)
	) name4735 (
		\rEIP_reg[20]/NET0131 ,
		_w4695_,
		_w5012_,
		_w5187_,
		_w5188_
	);
	LUT2 #(
		.INIT('h1)
	) name4736 (
		_w5186_,
		_w5188_,
		_w5189_
	);
	LUT2 #(
		.INIT('hb)
	) name4737 (
		_w5185_,
		_w5189_,
		_w5190_
	);
	LUT3 #(
		.INIT('h48)
	) name4738 (
		\rEIP_reg[9]/NET0131 ,
		_w592_,
		_w4679_,
		_w5191_
	);
	LUT3 #(
		.INIT('h8a)
	) name4739 (
		\Address[7]_pad ,
		\State_reg[0]/NET0131 ,
		\State_reg[1]/NET0131 ,
		_w5192_
	);
	LUT3 #(
		.INIT('h07)
	) name4740 (
		\rEIP_reg[0]/NET0131 ,
		\rEIP_reg[31]/NET0131 ,
		\rEIP_reg[8]/NET0131 ,
		_w5193_
	);
	LUT2 #(
		.INIT('h2)
	) name4741 (
		_w4695_,
		_w5193_,
		_w5194_
	);
	LUT4 #(
		.INIT('h6f00)
	) name4742 (
		\rEIP_reg[8]/NET0131 ,
		_w3149_,
		_w4691_,
		_w5194_,
		_w5195_
	);
	LUT2 #(
		.INIT('h1)
	) name4743 (
		_w5192_,
		_w5195_,
		_w5196_
	);
	LUT2 #(
		.INIT('hb)
	) name4744 (
		_w5191_,
		_w5196_,
		_w5197_
	);
	LUT3 #(
		.INIT('h48)
	) name4745 (
		\rEIP_reg[16]/NET0131 ,
		_w592_,
		_w4683_,
		_w5198_
	);
	LUT3 #(
		.INIT('h8a)
	) name4746 (
		\Address[14]_pad ,
		\State_reg[0]/NET0131 ,
		\State_reg[1]/NET0131 ,
		_w5199_
	);
	LUT4 #(
		.INIT('h8000)
	) name4747 (
		\rEIP_reg[11]/NET0131 ,
		_w3150_,
		_w3152_,
		_w4691_,
		_w5200_
	);
	LUT4 #(
		.INIT('h0c08)
	) name4748 (
		\rEIP_reg[15]/NET0131 ,
		_w4695_,
		_w5163_,
		_w5200_,
		_w5201_
	);
	LUT2 #(
		.INIT('h1)
	) name4749 (
		_w5199_,
		_w5201_,
		_w5202_
	);
	LUT2 #(
		.INIT('hb)
	) name4750 (
		_w5198_,
		_w5202_,
		_w5203_
	);
	LUT3 #(
		.INIT('h8a)
	) name4751 (
		\Address[26]_pad ,
		\State_reg[0]/NET0131 ,
		\State_reg[1]/NET0131 ,
		_w5204_
	);
	LUT4 #(
		.INIT('h60a0)
	) name4752 (
		\rEIP_reg[27]/NET0131 ,
		_w3269_,
		_w4695_,
		_w4692_,
		_w5205_
	);
	LUT2 #(
		.INIT('h1)
	) name4753 (
		_w5204_,
		_w5205_,
		_w5206_
	);
	LUT4 #(
		.INIT('h48ff)
	) name4754 (
		\rEIP_reg[28]/NET0131 ,
		_w592_,
		_w4687_,
		_w5206_,
		_w5207_
	);
	LUT3 #(
		.INIT('h8a)
	) name4755 (
		\Address[22]_pad ,
		\State_reg[0]/NET0131 ,
		\State_reg[1]/NET0131 ,
		_w5208_
	);
	LUT4 #(
		.INIT('h1555)
	) name4756 (
		\rEIP_reg[23]/NET0131 ,
		_w3155_,
		_w3196_,
		_w4691_,
		_w5209_
	);
	LUT4 #(
		.INIT('h0f0d)
	) name4757 (
		_w4695_,
		_w4692_,
		_w5208_,
		_w5209_,
		_w5210_
	);
	LUT4 #(
		.INIT('h48ff)
	) name4758 (
		\rEIP_reg[24]/NET0131 ,
		_w592_,
		_w4685_,
		_w5210_,
		_w5211_
	);
	LUT3 #(
		.INIT('h48)
	) name4759 (
		\rEIP_reg[12]/NET0131 ,
		_w592_,
		_w4681_,
		_w5212_
	);
	LUT3 #(
		.INIT('h8a)
	) name4760 (
		\Address[10]_pad ,
		\State_reg[0]/NET0131 ,
		\State_reg[1]/NET0131 ,
		_w5213_
	);
	LUT4 #(
		.INIT('h60a0)
	) name4761 (
		\rEIP_reg[11]/NET0131 ,
		_w3150_,
		_w4695_,
		_w4691_,
		_w5214_
	);
	LUT2 #(
		.INIT('h1)
	) name4762 (
		_w5213_,
		_w5214_,
		_w5215_
	);
	LUT2 #(
		.INIT('hb)
	) name4763 (
		_w5212_,
		_w5215_,
		_w5216_
	);
	LUT4 #(
		.INIT('h60c0)
	) name4764 (
		\rEIP_reg[3]/NET0131 ,
		\rEIP_reg[4]/NET0131 ,
		_w592_,
		_w4675_,
		_w5217_
	);
	LUT3 #(
		.INIT('h8a)
	) name4765 (
		\Address[2]_pad ,
		\State_reg[0]/NET0131 ,
		\State_reg[1]/NET0131 ,
		_w5218_
	);
	LUT4 #(
		.INIT('h00b7)
	) name4766 (
		\rEIP_reg[3]/NET0131 ,
		_w4695_,
		_w5181_,
		_w5218_,
		_w5219_
	);
	LUT2 #(
		.INIT('hb)
	) name4767 (
		_w5217_,
		_w5219_,
		_w5220_
	);
	LUT4 #(
		.INIT('h60c0)
	) name4768 (
		\rEIP_reg[19]/NET0131 ,
		\rEIP_reg[20]/NET0131 ,
		_w592_,
		_w4730_,
		_w5221_
	);
	LUT3 #(
		.INIT('h8a)
	) name4769 (
		\Address[18]_pad ,
		\State_reg[0]/NET0131 ,
		\State_reg[1]/NET0131 ,
		_w5222_
	);
	LUT4 #(
		.INIT('h1555)
	) name4770 (
		\rEIP_reg[19]/NET0131 ,
		_w3155_,
		_w3156_,
		_w4691_,
		_w5223_
	);
	LUT4 #(
		.INIT('h0f0d)
	) name4771 (
		_w4695_,
		_w5187_,
		_w5222_,
		_w5223_,
		_w5224_
	);
	LUT2 #(
		.INIT('hb)
	) name4772 (
		_w5221_,
		_w5224_,
		_w5225_
	);
	LUT3 #(
		.INIT('h8a)
	) name4773 (
		\Address[6]_pad ,
		\State_reg[0]/NET0131 ,
		\State_reg[1]/NET0131 ,
		_w5226_
	);
	LUT3 #(
		.INIT('h07)
	) name4774 (
		\rEIP_reg[0]/NET0131 ,
		\rEIP_reg[31]/NET0131 ,
		\rEIP_reg[7]/NET0131 ,
		_w5227_
	);
	LUT2 #(
		.INIT('h2)
	) name4775 (
		_w4695_,
		_w5227_,
		_w5228_
	);
	LUT4 #(
		.INIT('h040f)
	) name4776 (
		_w3442_,
		_w4691_,
		_w5226_,
		_w5228_,
		_w5229_
	);
	LUT4 #(
		.INIT('h48ff)
	) name4777 (
		\rEIP_reg[8]/NET0131 ,
		_w592_,
		_w4678_,
		_w5229_,
		_w5230_
	);
	LUT3 #(
		.INIT('h8a)
	) name4778 (
		\Address[25]_pad ,
		\State_reg[0]/NET0131 ,
		\State_reg[1]/NET0131 ,
		_w5231_
	);
	LUT3 #(
		.INIT('h15)
	) name4779 (
		\rEIP_reg[26]/NET0131 ,
		_w3250_,
		_w4691_,
		_w5232_
	);
	LUT3 #(
		.INIT('h4c)
	) name4780 (
		_w3269_,
		_w4695_,
		_w4692_,
		_w5233_
	);
	LUT3 #(
		.INIT('h45)
	) name4781 (
		_w5231_,
		_w5232_,
		_w5233_,
		_w5234_
	);
	LUT4 #(
		.INIT('h48ff)
	) name4782 (
		\rEIP_reg[27]/NET0131 ,
		_w592_,
		_w4686_,
		_w5234_,
		_w5235_
	);
	LUT3 #(
		.INIT('h8a)
	) name4783 (
		\Address[29]_pad ,
		\State_reg[0]/NET0131 ,
		\State_reg[1]/NET0131 ,
		_w5236_
	);
	LUT3 #(
		.INIT('h13)
	) name4784 (
		\rEIP_reg[0]/NET0131 ,
		\rEIP_reg[30]/NET0131 ,
		\rEIP_reg[31]/NET0131 ,
		_w5237_
	);
	LUT2 #(
		.INIT('h2)
	) name4785 (
		_w4695_,
		_w5237_,
		_w5238_
	);
	LUT4 #(
		.INIT('h6f00)
	) name4786 (
		\rEIP_reg[30]/NET0131 ,
		_w3314_,
		_w4691_,
		_w5238_,
		_w5239_
	);
	LUT2 #(
		.INIT('h1)
	) name4787 (
		_w5236_,
		_w5239_,
		_w5240_
	);
	LUT4 #(
		.INIT('h48ff)
	) name4788 (
		\rEIP_reg[31]/NET0131 ,
		_w592_,
		_w4689_,
		_w5240_,
		_w5241_
	);
	LUT3 #(
		.INIT('h8a)
	) name4789 (
		\Address[13]_pad ,
		\State_reg[0]/NET0131 ,
		\State_reg[1]/NET0131 ,
		_w5242_
	);
	LUT3 #(
		.INIT('h13)
	) name4790 (
		\rEIP_reg[0]/NET0131 ,
		\rEIP_reg[14]/NET0131 ,
		\rEIP_reg[31]/NET0131 ,
		_w5243_
	);
	LUT2 #(
		.INIT('h2)
	) name4791 (
		_w4695_,
		_w5243_,
		_w5244_
	);
	LUT4 #(
		.INIT('h040f)
	) name4792 (
		_w3571_,
		_w4691_,
		_w5242_,
		_w5244_,
		_w5245_
	);
	LUT4 #(
		.INIT('h48ff)
	) name4793 (
		\rEIP_reg[15]/NET0131 ,
		_w592_,
		_w4682_,
		_w5245_,
		_w5246_
	);
	LUT3 #(
		.INIT('h8a)
	) name4794 (
		\Address[9]_pad ,
		\State_reg[0]/NET0131 ,
		\State_reg[1]/NET0131 ,
		_w5247_
	);
	LUT3 #(
		.INIT('h13)
	) name4795 (
		\rEIP_reg[0]/NET0131 ,
		\rEIP_reg[10]/NET0131 ,
		\rEIP_reg[31]/NET0131 ,
		_w5248_
	);
	LUT2 #(
		.INIT('h2)
	) name4796 (
		_w4695_,
		_w5248_,
		_w5249_
	);
	LUT4 #(
		.INIT('h040f)
	) name4797 (
		_w3499_,
		_w4691_,
		_w5247_,
		_w5249_,
		_w5250_
	);
	LUT4 #(
		.INIT('h48ff)
	) name4798 (
		\rEIP_reg[11]/NET0131 ,
		_w592_,
		_w4680_,
		_w5250_,
		_w5251_
	);
	LUT3 #(
		.INIT('h13)
	) name4799 (
		\rEIP_reg[0]/NET0131 ,
		\rEIP_reg[22]/NET0131 ,
		\rEIP_reg[31]/NET0131 ,
		_w5252_
	);
	LUT2 #(
		.INIT('h2)
	) name4800 (
		_w4695_,
		_w5252_,
		_w5253_
	);
	LUT3 #(
		.INIT('h8a)
	) name4801 (
		\Address[21]_pad ,
		\State_reg[0]/NET0131 ,
		\State_reg[1]/NET0131 ,
		_w5254_
	);
	LUT4 #(
		.INIT('h004f)
	) name4802 (
		_w3197_,
		_w4691_,
		_w5253_,
		_w5254_,
		_w5255_
	);
	LUT4 #(
		.INIT('h48ff)
	) name4803 (
		\rEIP_reg[23]/NET0131 ,
		_w592_,
		_w4684_,
		_w5255_,
		_w5256_
	);
	LUT2 #(
		.INIT('h7)
	) name4804 (
		\DataWidth_reg[0]/NET0131 ,
		\DataWidth_reg[1]/NET0131 ,
		_w5257_
	);
	LUT3 #(
		.INIT('h80)
	) name4805 (
		\ByteEnable_reg[2]/NET0131 ,
		\DataWidth_reg[0]/NET0131 ,
		\DataWidth_reg[1]/NET0131 ,
		_w5258_
	);
	LUT4 #(
		.INIT('h7013)
	) name4806 (
		\DataWidth_reg[0]/NET0131 ,
		\DataWidth_reg[1]/NET0131 ,
		\rEIP_reg[0]/NET0131 ,
		\rEIP_reg[1]/NET0131 ,
		_w5259_
	);
	LUT2 #(
		.INIT('he)
	) name4807 (
		_w5258_,
		_w5259_,
		_w5260_
	);
	LUT4 #(
		.INIT('h3310)
	) name4808 (
		HOLD_pad,
		READY_n_pad,
		\State_reg[0]/NET0131 ,
		\State_reg[2]/NET0131 ,
		_w5261_
	);
	LUT4 #(
		.INIT('h40c0)
	) name4809 (
		HOLD_pad,
		\RequestPending_reg/NET0131 ,
		\State_reg[0]/NET0131 ,
		\State_reg[2]/NET0131 ,
		_w5262_
	);
	LUT4 #(
		.INIT('hfcfe)
	) name4810 (
		\State_reg[1]/NET0131 ,
		_w593_,
		_w5262_,
		_w5261_,
		_w5263_
	);
	LUT3 #(
		.INIT('h01)
	) name4811 (
		\DataWidth_reg[0]/NET0131 ,
		\DataWidth_reg[1]/NET0131 ,
		\rEIP_reg[0]/NET0131 ,
		_w5264_
	);
	LUT4 #(
		.INIT('h407f)
	) name4812 (
		\ByteEnable_reg[1]/NET0131 ,
		\DataWidth_reg[0]/NET0131 ,
		\DataWidth_reg[1]/NET0131 ,
		\rEIP_reg[1]/NET0131 ,
		_w5265_
	);
	LUT2 #(
		.INIT('hb)
	) name4813 (
		_w5264_,
		_w5265_,
		_w5266_
	);
	LUT4 #(
		.INIT('h0acf)
	) name4814 (
		NA_n_pad,
		READY_n_pad,
		\State_reg[0]/NET0131 ,
		\State_reg[2]/NET0131 ,
		_w5267_
	);
	LUT3 #(
		.INIT('h02)
	) name4815 (
		\State_reg[0]/NET0131 ,
		\State_reg[1]/NET0131 ,
		\State_reg[2]/NET0131 ,
		_w5268_
	);
	LUT4 #(
		.INIT('hcc04)
	) name4816 (
		HOLD_pad,
		\RequestPending_reg/NET0131 ,
		_w5267_,
		_w5268_,
		_w5269_
	);
	LUT2 #(
		.INIT('h1)
	) name4817 (
		_w4695_,
		_w5269_,
		_w5270_
	);
	LUT3 #(
		.INIT('h48)
	) name4818 (
		\rEIP_reg[3]/NET0131 ,
		_w592_,
		_w4675_,
		_w5271_
	);
	LUT3 #(
		.INIT('h8a)
	) name4819 (
		\Address[1]_pad ,
		\State_reg[0]/NET0131 ,
		\State_reg[1]/NET0131 ,
		_w5272_
	);
	LUT4 #(
		.INIT('h00b7)
	) name4820 (
		\rEIP_reg[2]/NET0131 ,
		_w4695_,
		_w5180_,
		_w5272_,
		_w5273_
	);
	LUT2 #(
		.INIT('hb)
	) name4821 (
		_w5271_,
		_w5273_,
		_w5274_
	);
	LUT3 #(
		.INIT('h8a)
	) name4822 (
		\Address[17]_pad ,
		\State_reg[0]/NET0131 ,
		\State_reg[1]/NET0131 ,
		_w5275_
	);
	LUT4 #(
		.INIT('h1333)
	) name4823 (
		\rEIP_reg[17]/NET0131 ,
		\rEIP_reg[18]/NET0131 ,
		_w3155_,
		_w4691_,
		_w5276_
	);
	LUT4 #(
		.INIT('h70f0)
	) name4824 (
		_w3155_,
		_w3156_,
		_w4695_,
		_w4691_,
		_w5277_
	);
	LUT3 #(
		.INIT('h45)
	) name4825 (
		_w5275_,
		_w5276_,
		_w5277_,
		_w5278_
	);
	LUT4 #(
		.INIT('h48ff)
	) name4826 (
		\rEIP_reg[19]/NET0131 ,
		_w592_,
		_w4730_,
		_w5278_,
		_w5279_
	);
	LUT4 #(
		.INIT('h60c0)
	) name4827 (
		\rEIP_reg[6]/NET0131 ,
		\rEIP_reg[7]/NET0131 ,
		_w592_,
		_w4677_,
		_w5280_
	);
	LUT3 #(
		.INIT('h8a)
	) name4828 (
		\Address[5]_pad ,
		\State_reg[0]/NET0131 ,
		\State_reg[1]/NET0131 ,
		_w5281_
	);
	LUT4 #(
		.INIT('h9300)
	) name4829 (
		\rEIP_reg[5]/NET0131 ,
		\rEIP_reg[6]/NET0131 ,
		_w3148_,
		_w4691_,
		_w5282_
	);
	LUT3 #(
		.INIT('h07)
	) name4830 (
		\rEIP_reg[0]/NET0131 ,
		\rEIP_reg[31]/NET0131 ,
		\rEIP_reg[6]/NET0131 ,
		_w5283_
	);
	LUT2 #(
		.INIT('h2)
	) name4831 (
		_w4695_,
		_w5283_,
		_w5284_
	);
	LUT3 #(
		.INIT('h45)
	) name4832 (
		_w5281_,
		_w5282_,
		_w5284_,
		_w5285_
	);
	LUT2 #(
		.INIT('hb)
	) name4833 (
		_w5280_,
		_w5285_,
		_w5286_
	);
	LUT3 #(
		.INIT('h08)
	) name4834 (
		\State_reg[0]/NET0131 ,
		\State_reg[1]/NET0131 ,
		\State_reg[2]/NET0131 ,
		_w5287_
	);
	LUT3 #(
		.INIT('hc8)
	) name4835 (
		HOLD_pad,
		READY_n_pad,
		\RequestPending_reg/NET0131 ,
		_w5288_
	);
	LUT4 #(
		.INIT('h5444)
	) name4836 (
		NA_n_pad,
		_w593_,
		_w5287_,
		_w5288_,
		_w5289_
	);
	LUT3 #(
		.INIT('h0e)
	) name4837 (
		\RequestPending_reg/NET0131 ,
		\State_reg[1]/NET0131 ,
		\State_reg[2]/NET0131 ,
		_w5290_
	);
	LUT2 #(
		.INIT('h8)
	) name4838 (
		HOLD_pad,
		\State_reg[0]/NET0131 ,
		_w5291_
	);
	LUT4 #(
		.INIT('hb000)
	) name4839 (
		READY_n_pad,
		\State_reg[0]/NET0131 ,
		\State_reg[1]/NET0131 ,
		\State_reg[2]/NET0131 ,
		_w5292_
	);
	LUT3 #(
		.INIT('h0b)
	) name4840 (
		_w5290_,
		_w5291_,
		_w5292_,
		_w5293_
	);
	LUT2 #(
		.INIT('hb)
	) name4841 (
		_w5289_,
		_w5293_,
		_w5294_
	);
	LUT3 #(
		.INIT('h80)
	) name4842 (
		\ByteEnable_reg[3]/NET0131 ,
		\DataWidth_reg[0]/NET0131 ,
		\DataWidth_reg[1]/NET0131 ,
		_w5295_
	);
	LUT4 #(
		.INIT('h0133)
	) name4843 (
		\DataWidth_reg[0]/NET0131 ,
		\DataWidth_reg[1]/NET0131 ,
		\rEIP_reg[0]/NET0131 ,
		\rEIP_reg[1]/NET0131 ,
		_w5296_
	);
	LUT2 #(
		.INIT('he)
	) name4844 (
		_w5295_,
		_w5296_,
		_w5297_
	);
	LUT3 #(
		.INIT('h48)
	) name4845 (
		\rEIP_reg[2]/NET0131 ,
		_w592_,
		_w4674_,
		_w5298_
	);
	LUT3 #(
		.INIT('h8a)
	) name4846 (
		\Address[0]_pad ,
		\State_reg[0]/NET0131 ,
		\State_reg[1]/NET0131 ,
		_w5299_
	);
	LUT4 #(
		.INIT('h00b7)
	) name4847 (
		\rEIP_reg[1]/NET0131 ,
		_w4695_,
		_w4691_,
		_w5299_,
		_w5300_
	);
	LUT2 #(
		.INIT('hb)
	) name4848 (
		_w5298_,
		_w5300_,
		_w5301_
	);
	LUT4 #(
		.INIT('h0140)
	) name4849 (
		\BS16_n_pad ,
		\State_reg[0]/NET0131 ,
		\State_reg[1]/NET0131 ,
		\State_reg[2]/NET0131 ,
		_w5302_
	);
	LUT4 #(
		.INIT('h5414)
	) name4850 (
		\DataWidth_reg[1]/NET0131 ,
		\State_reg[0]/NET0131 ,
		\State_reg[1]/NET0131 ,
		\State_reg[2]/NET0131 ,
		_w5303_
	);
	LUT2 #(
		.INIT('h1)
	) name4851 (
		_w5302_,
		_w5303_,
		_w5304_
	);
	LUT4 #(
		.INIT('hacaa)
	) name4852 (
		\BE_n[2]_pad ,
		\ByteEnable_reg[2]/NET0131 ,
		\State_reg[0]/NET0131 ,
		\State_reg[1]/NET0131 ,
		_w5305_
	);
	LUT4 #(
		.INIT('h8bcb)
	) name4853 (
		ADS_n_pad,
		\State_reg[0]/NET0131 ,
		\State_reg[1]/NET0131 ,
		\State_reg[2]/NET0131 ,
		_w5306_
	);
	LUT4 #(
		.INIT('hacaa)
	) name4854 (
		\BE_n[0]_pad ,
		\ByteEnable_reg[0]/NET0131 ,
		\State_reg[0]/NET0131 ,
		\State_reg[1]/NET0131 ,
		_w5307_
	);
	LUT4 #(
		.INIT('hacaa)
	) name4855 (
		\BE_n[1]_pad ,
		\ByteEnable_reg[1]/NET0131 ,
		\State_reg[0]/NET0131 ,
		\State_reg[1]/NET0131 ,
		_w5308_
	);
	LUT4 #(
		.INIT('hacaa)
	) name4856 (
		\BE_n[3]_pad ,
		\ByteEnable_reg[3]/NET0131 ,
		\State_reg[0]/NET0131 ,
		\State_reg[1]/NET0131 ,
		_w5309_
	);
	LUT4 #(
		.INIT('hacaa)
	) name4857 (
		M_IO_n_pad,
		\MemoryFetch_reg/NET0131 ,
		\State_reg[0]/NET0131 ,
		\State_reg[1]/NET0131 ,
		_w5310_
	);
	LUT4 #(
		.INIT('hdf10)
	) name4858 (
		\ReadRequest_reg/NET0131 ,
		\State_reg[0]/NET0131 ,
		\State_reg[1]/NET0131 ,
		W_R_n_pad,
		_w5311_
	);
	LUT4 #(
		.INIT('h4544)
	) name4859 (
		D_C_n_pad,
		\State_reg[0]/NET0131 ,
		\State_reg[1]/NET0131 ,
		\State_reg[2]/NET0131 ,
		_w5312_
	);
	LUT3 #(
		.INIT('h20)
	) name4860 (
		\CodeFetch_reg/NET0131 ,
		\State_reg[0]/NET0131 ,
		\State_reg[1]/NET0131 ,
		_w5313_
	);
	LUT2 #(
		.INIT('h1)
	) name4861 (
		_w5312_,
		_w5313_,
		_w5314_
	);
	LUT4 #(
		.INIT('ha828)
	) name4862 (
		\DataWidth_reg[0]/NET0131 ,
		\State_reg[0]/NET0131 ,
		\State_reg[1]/NET0131 ,
		\State_reg[2]/NET0131 ,
		_w5315_
	);
	LUT2 #(
		.INIT('he)
	) name4863 (
		_w5302_,
		_w5315_,
		_w5316_
	);
	LUT3 #(
		.INIT('h08)
	) name4864 (
		\InstAddrPointer_reg[28]/NET0131 ,
		_w563_,
		_w673_,
		_w5317_
	);
	LUT4 #(
		.INIT('haa20)
	) name4865 (
		_w608_,
		_w1425_,
		_w1428_,
		_w5317_,
		_w5318_
	);
	LUT3 #(
		.INIT('h54)
	) name4866 (
		\InstAddrPointer_reg[28]/NET0131 ,
		_w563_,
		_w633_,
		_w5319_
	);
	LUT4 #(
		.INIT('h00c8)
	) name4867 (
		_w569_,
		_w602_,
		_w604_,
		_w5319_,
		_w5320_
	);
	LUT2 #(
		.INIT('h8)
	) name4868 (
		_w1431_,
		_w5320_,
		_w5321_
	);
	LUT3 #(
		.INIT('hb0)
	) name4869 (
		_w616_,
		_w630_,
		_w996_,
		_w5322_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name4870 (
		\InstAddrPointer_reg[28]/NET0131 ,
		_w597_,
		_w1076_,
		_w1427_,
		_w5323_
	);
	LUT3 #(
		.INIT('h10)
	) name4871 (
		_w5321_,
		_w5322_,
		_w5323_,
		_w5324_
	);
	LUT4 #(
		.INIT('hd700)
	) name4872 (
		_w671_,
		_w1431_,
		_w1436_,
		_w5324_,
		_w5325_
	);
	LUT4 #(
		.INIT('h153f)
	) name4873 (
		\InstAddrPointer_reg[28]/NET0131 ,
		\rEIP_reg[28]/NET0131 ,
		_w1080_,
		_w1081_,
		_w5326_
	);
	LUT4 #(
		.INIT('h8aff)
	) name4874 (
		_w690_,
		_w5318_,
		_w5325_,
		_w5326_,
		_w5327_
	);
	LUT3 #(
		.INIT('h08)
	) name4875 (
		\PhyAddrPointer_reg[12]/NET0131 ,
		_w563_,
		_w673_,
		_w5328_
	);
	LUT4 #(
		.INIT('h5515)
	) name4876 (
		_w886_,
		_w1131_,
		_w1135_,
		_w1270_,
		_w5329_
	);
	LUT3 #(
		.INIT('ha8)
	) name4877 (
		_w836_,
		_w1334_,
		_w5329_,
		_w5330_
	);
	LUT4 #(
		.INIT('h4554)
	) name4878 (
		_w674_,
		_w836_,
		_w951_,
		_w1315_,
		_w5331_
	);
	LUT4 #(
		.INIT('h8a88)
	) name4879 (
		_w608_,
		_w5328_,
		_w5330_,
		_w5331_,
		_w5332_
	);
	LUT4 #(
		.INIT('h202a)
	) name4880 (
		\PhyAddrPointer_reg[12]/NET0131 ,
		_w634_,
		_w607_,
		_w608_,
		_w5333_
	);
	LUT4 #(
		.INIT('h48c0)
	) name4881 (
		\InstAddrPointer_reg[11]/NET0131 ,
		_w671_,
		_w1042_,
		_w1341_,
		_w5334_
	);
	LUT2 #(
		.INIT('h1)
	) name4882 (
		_w5333_,
		_w5334_,
		_w5335_
	);
	LUT4 #(
		.INIT('h4111)
	) name4883 (
		\DataWidth_reg[1]/NET0131 ,
		\PhyAddrPointer_reg[12]/NET0131 ,
		\PhyAddrPointer_reg[1]/NET0131 ,
		_w1491_,
		_w5336_
	);
	LUT4 #(
		.INIT('h820a)
	) name4884 (
		\DataWidth_reg[1]/NET0131 ,
		\PhyAddrPointer_reg[11]/NET0131 ,
		\PhyAddrPointer_reg[12]/NET0131 ,
		_w1195_,
		_w5337_
	);
	LUT3 #(
		.INIT('h02)
	) name4885 (
		_w695_,
		_w5337_,
		_w5336_,
		_w5338_
	);
	LUT4 #(
		.INIT('h60a0)
	) name4886 (
		\PhyAddrPointer_reg[12]/NET0131 ,
		\PhyAddrPointer_reg[1]/NET0131 ,
		_w1212_,
		_w1491_,
		_w5339_
	);
	LUT4 #(
		.INIT('h3f15)
	) name4887 (
		\PhyAddrPointer_reg[12]/NET0131 ,
		\rEIP_reg[12]/NET0131 ,
		_w1080_,
		_w1215_,
		_w5340_
	);
	LUT2 #(
		.INIT('h4)
	) name4888 (
		_w5339_,
		_w5340_,
		_w5341_
	);
	LUT2 #(
		.INIT('h4)
	) name4889 (
		_w5338_,
		_w5341_,
		_w5342_
	);
	LUT4 #(
		.INIT('h8aff)
	) name4890 (
		_w690_,
		_w5332_,
		_w5335_,
		_w5342_,
		_w5343_
	);
	LUT3 #(
		.INIT('h08)
	) name4891 (
		\InstAddrPointer_reg[17]/NET0131 ,
		_w563_,
		_w673_,
		_w5344_
	);
	LUT4 #(
		.INIT('haa20)
	) name4892 (
		_w608_,
		_w1630_,
		_w1632_,
		_w5344_,
		_w5345_
	);
	LUT2 #(
		.INIT('h4)
	) name4893 (
		_w597_,
		_w1628_,
		_w5346_
	);
	LUT2 #(
		.INIT('h8)
	) name4894 (
		_w635_,
		_w1040_,
		_w5347_
	);
	LUT4 #(
		.INIT('h004f)
	) name4895 (
		_w616_,
		_w630_,
		_w975_,
		_w5347_,
		_w5348_
	);
	LUT4 #(
		.INIT('h0d00)
	) name4896 (
		\InstAddrPointer_reg[17]/NET0131 ,
		_w1165_,
		_w5346_,
		_w5348_,
		_w5349_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name4897 (
		_w690_,
		_w1638_,
		_w5345_,
		_w5349_,
		_w5350_
	);
	LUT4 #(
		.INIT('h153f)
	) name4898 (
		\InstAddrPointer_reg[17]/NET0131 ,
		\rEIP_reg[17]/NET0131 ,
		_w1080_,
		_w1081_,
		_w5351_
	);
	LUT2 #(
		.INIT('hb)
	) name4899 (
		_w5350_,
		_w5351_,
		_w5352_
	);
	LUT3 #(
		.INIT('h08)
	) name4900 (
		\InstAddrPointer_reg[19]/NET0131 ,
		_w563_,
		_w673_,
		_w5353_
	);
	LUT4 #(
		.INIT('haa20)
	) name4901 (
		_w608_,
		_w1510_,
		_w1514_,
		_w5353_,
		_w5354_
	);
	LUT4 #(
		.INIT('hec00)
	) name4902 (
		_w585_,
		_w589_,
		_w590_,
		_w884_,
		_w5355_
	);
	LUT4 #(
		.INIT('h0004)
	) name4903 (
		_w613_,
		_w681_,
		_w1368_,
		_w5355_,
		_w5356_
	);
	LUT2 #(
		.INIT('h4)
	) name4904 (
		_w597_,
		_w884_,
		_w5357_
	);
	LUT2 #(
		.INIT('h8)
	) name4905 (
		_w635_,
		_w1061_,
		_w5358_
	);
	LUT4 #(
		.INIT('h004f)
	) name4906 (
		_w616_,
		_w630_,
		_w974_,
		_w5358_,
		_w5359_
	);
	LUT4 #(
		.INIT('h0d00)
	) name4907 (
		\InstAddrPointer_reg[19]/NET0131 ,
		_w5356_,
		_w5357_,
		_w5359_,
		_w5360_
	);
	LUT2 #(
		.INIT('h4)
	) name4908 (
		_w1517_,
		_w5360_,
		_w5361_
	);
	LUT4 #(
		.INIT('h153f)
	) name4909 (
		\InstAddrPointer_reg[19]/NET0131 ,
		\rEIP_reg[19]/NET0131 ,
		_w1080_,
		_w1081_,
		_w5362_
	);
	LUT4 #(
		.INIT('h8aff)
	) name4910 (
		_w690_,
		_w5354_,
		_w5361_,
		_w5362_,
		_w5363_
	);
	LUT3 #(
		.INIT('h08)
	) name4911 (
		\InstAddrPointer_reg[16]/NET0131 ,
		_w563_,
		_w673_,
		_w5364_
	);
	LUT4 #(
		.INIT('haa20)
	) name4912 (
		_w608_,
		_w1611_,
		_w1614_,
		_w5364_,
		_w5365_
	);
	LUT2 #(
		.INIT('h4)
	) name4913 (
		_w597_,
		_w1610_,
		_w5366_
	);
	LUT2 #(
		.INIT('h2)
	) name4914 (
		\InstAddrPointer_reg[16]/NET0131 ,
		_w1295_,
		_w5367_
	);
	LUT2 #(
		.INIT('h8)
	) name4915 (
		_w635_,
		_w1156_,
		_w5368_
	);
	LUT4 #(
		.INIT('h004f)
	) name4916 (
		_w616_,
		_w630_,
		_w971_,
		_w5368_,
		_w5369_
	);
	LUT3 #(
		.INIT('h10)
	) name4917 (
		_w5366_,
		_w5367_,
		_w5369_,
		_w5370_
	);
	LUT2 #(
		.INIT('h4)
	) name4918 (
		_w1618_,
		_w5370_,
		_w5371_
	);
	LUT4 #(
		.INIT('h153f)
	) name4919 (
		\InstAddrPointer_reg[16]/NET0131 ,
		\rEIP_reg[16]/NET0131 ,
		_w1080_,
		_w1081_,
		_w5372_
	);
	LUT4 #(
		.INIT('h8aff)
	) name4920 (
		_w690_,
		_w5365_,
		_w5371_,
		_w5372_,
		_w5373_
	);
	LUT3 #(
		.INIT('h08)
	) name4921 (
		\InstAddrPointer_reg[20]/NET0131 ,
		_w563_,
		_w673_,
		_w5374_
	);
	LUT4 #(
		.INIT('h4000)
	) name4922 (
		_w948_,
		_w964_,
		_w972_,
		_w977_,
		_w5375_
	);
	LUT3 #(
		.INIT('h41)
	) name4923 (
		_w836_,
		_w968_,
		_w5375_,
		_w5376_
	);
	LUT4 #(
		.INIT('h2322)
	) name4924 (
		_w878_,
		_w894_,
		_w1270_,
		_w1271_,
		_w5377_
	);
	LUT3 #(
		.INIT('h51)
	) name4925 (
		_w674_,
		_w836_,
		_w5377_,
		_w5378_
	);
	LUT4 #(
		.INIT('h8a88)
	) name4926 (
		_w608_,
		_w5374_,
		_w5376_,
		_w5378_,
		_w5379_
	);
	LUT3 #(
		.INIT('h07)
	) name4927 (
		_w719_,
		_w1255_,
		_w1432_,
		_w5380_
	);
	LUT3 #(
		.INIT('h2a)
	) name4928 (
		_w671_,
		_w1112_,
		_w1255_,
		_w5381_
	);
	LUT3 #(
		.INIT('h21)
	) name4929 (
		\InstAddrPointer_reg[20]/NET0131 ,
		READY_n_pad,
		_w733_,
		_w5382_
	);
	LUT3 #(
		.INIT('h08)
	) name4930 (
		_w494_,
		_w586_,
		_w5382_,
		_w5383_
	);
	LUT2 #(
		.INIT('h1)
	) name4931 (
		_w680_,
		_w5383_,
		_w5384_
	);
	LUT3 #(
		.INIT('h8a)
	) name4932 (
		\InstAddrPointer_reg[20]/NET0131 ,
		_w613_,
		_w5384_,
		_w5385_
	);
	LUT3 #(
		.INIT('hb0)
	) name4933 (
		_w616_,
		_w630_,
		_w968_,
		_w5386_
	);
	LUT3 #(
		.INIT('h9a)
	) name4934 (
		\InstAddrPointer_reg[20]/NET0131 ,
		READY_n_pad,
		_w733_,
		_w5387_
	);
	LUT3 #(
		.INIT('he0)
	) name4935 (
		_w588_,
		_w596_,
		_w5387_,
		_w5388_
	);
	LUT2 #(
		.INIT('h8)
	) name4936 (
		_w554_,
		_w878_,
		_w5389_
	);
	LUT2 #(
		.INIT('h2)
	) name4937 (
		_w634_,
		_w1432_,
		_w5390_
	);
	LUT3 #(
		.INIT('h54)
	) name4938 (
		\InstAddrPointer_reg[20]/NET0131 ,
		_w563_,
		_w633_,
		_w5391_
	);
	LUT4 #(
		.INIT('h00c8)
	) name4939 (
		_w569_,
		_w602_,
		_w604_,
		_w5391_,
		_w5392_
	);
	LUT3 #(
		.INIT('h45)
	) name4940 (
		_w5389_,
		_w5390_,
		_w5392_,
		_w5393_
	);
	LUT2 #(
		.INIT('h4)
	) name4941 (
		_w5388_,
		_w5393_,
		_w5394_
	);
	LUT3 #(
		.INIT('h10)
	) name4942 (
		_w5386_,
		_w5385_,
		_w5394_,
		_w5395_
	);
	LUT3 #(
		.INIT('hb0)
	) name4943 (
		_w5380_,
		_w5381_,
		_w5395_,
		_w5396_
	);
	LUT4 #(
		.INIT('h153f)
	) name4944 (
		\InstAddrPointer_reg[20]/NET0131 ,
		\rEIP_reg[20]/NET0131 ,
		_w1080_,
		_w1081_,
		_w5397_
	);
	LUT4 #(
		.INIT('h8aff)
	) name4945 (
		_w690_,
		_w5379_,
		_w5396_,
		_w5397_,
		_w5398_
	);
	LUT3 #(
		.INIT('h08)
	) name4946 (
		\InstAddrPointer_reg[18]/NET0131 ,
		_w563_,
		_w673_,
		_w5399_
	);
	LUT4 #(
		.INIT('haa20)
	) name4947 (
		_w608_,
		_w1648_,
		_w1651_,
		_w5399_,
		_w5400_
	);
	LUT2 #(
		.INIT('h4)
	) name4948 (
		_w597_,
		_w880_,
		_w5401_
	);
	LUT2 #(
		.INIT('h8)
	) name4949 (
		_w635_,
		_w1054_,
		_w5402_
	);
	LUT4 #(
		.INIT('h004f)
	) name4950 (
		_w616_,
		_w630_,
		_w976_,
		_w5402_,
		_w5403_
	);
	LUT4 #(
		.INIT('h0d00)
	) name4951 (
		\InstAddrPointer_reg[18]/NET0131 ,
		_w1165_,
		_w5401_,
		_w5403_,
		_w5404_
	);
	LUT2 #(
		.INIT('h4)
	) name4952 (
		_w1655_,
		_w5404_,
		_w5405_
	);
	LUT4 #(
		.INIT('h153f)
	) name4953 (
		\InstAddrPointer_reg[18]/NET0131 ,
		\rEIP_reg[18]/NET0131 ,
		_w1080_,
		_w1081_,
		_w5406_
	);
	LUT4 #(
		.INIT('h8aff)
	) name4954 (
		_w690_,
		_w5400_,
		_w5405_,
		_w5406_,
		_w5407_
	);
	LUT3 #(
		.INIT('h08)
	) name4955 (
		\InstAddrPointer_reg[31]/NET0131 ,
		_w563_,
		_w673_,
		_w5408_
	);
	LUT4 #(
		.INIT('haa20)
	) name4956 (
		_w608_,
		_w1176_,
		_w1178_,
		_w5408_,
		_w5409_
	);
	LUT3 #(
		.INIT('h48)
	) name4957 (
		\InstAddrPointer_reg[31]/NET0131 ,
		_w635_,
		_w1068_,
		_w5410_
	);
	LUT3 #(
		.INIT('hb0)
	) name4958 (
		_w616_,
		_w630_,
		_w1175_,
		_w5411_
	);
	LUT4 #(
		.INIT('h00ec)
	) name4959 (
		_w585_,
		_w589_,
		_w590_,
		_w743_,
		_w5412_
	);
	LUT4 #(
		.INIT('h0004)
	) name4960 (
		_w613_,
		_w681_,
		_w1368_,
		_w5412_,
		_w5413_
	);
	LUT2 #(
		.INIT('h4)
	) name4961 (
		_w597_,
		_w1177_,
		_w5414_
	);
	LUT4 #(
		.INIT('h0031)
	) name4962 (
		\InstAddrPointer_reg[31]/NET0131 ,
		_w5411_,
		_w5413_,
		_w5414_,
		_w5415_
	);
	LUT2 #(
		.INIT('h4)
	) name4963 (
		_w5410_,
		_w5415_,
		_w5416_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name4964 (
		_w690_,
		_w1186_,
		_w5409_,
		_w5416_,
		_w5417_
	);
	LUT4 #(
		.INIT('h153f)
	) name4965 (
		\InstAddrPointer_reg[31]/NET0131 ,
		\rEIP_reg[31]/NET0131 ,
		_w1080_,
		_w1081_,
		_w5418_
	);
	LUT2 #(
		.INIT('hb)
	) name4966 (
		_w5417_,
		_w5418_,
		_w5419_
	);
	LUT3 #(
		.INIT('h08)
	) name4967 (
		\InstAddrPointer_reg[23]/NET0131 ,
		_w563_,
		_w673_,
		_w5420_
	);
	LUT4 #(
		.INIT('haa20)
	) name4968 (
		_w608_,
		_w1397_,
		_w1399_,
		_w5420_,
		_w5421_
	);
	LUT3 #(
		.INIT('hb8)
	) name4969 (
		\InstAddrPointer_reg[23]/NET0131 ,
		READY_n_pad,
		_w906_,
		_w5422_
	);
	LUT4 #(
		.INIT('hec00)
	) name4970 (
		_w585_,
		_w589_,
		_w590_,
		_w5422_,
		_w5423_
	);
	LUT4 #(
		.INIT('haa8a)
	) name4971 (
		\InstAddrPointer_reg[23]/NET0131 ,
		_w613_,
		_w681_,
		_w5423_,
		_w5424_
	);
	LUT2 #(
		.INIT('h8)
	) name4972 (
		_w554_,
		_w906_,
		_w5425_
	);
	LUT3 #(
		.INIT('h07)
	) name4973 (
		_w635_,
		_w1161_,
		_w5425_,
		_w5426_
	);
	LUT3 #(
		.INIT('he0)
	) name4974 (
		_w588_,
		_w596_,
		_w5422_,
		_w5427_
	);
	LUT4 #(
		.INIT('h004f)
	) name4975 (
		_w616_,
		_w630_,
		_w983_,
		_w5427_,
		_w5428_
	);
	LUT3 #(
		.INIT('h40)
	) name4976 (
		_w5424_,
		_w5426_,
		_w5428_,
		_w5429_
	);
	LUT3 #(
		.INIT('hb0)
	) name4977 (
		_w1402_,
		_w1403_,
		_w5429_,
		_w5430_
	);
	LUT4 #(
		.INIT('h153f)
	) name4978 (
		\InstAddrPointer_reg[23]/NET0131 ,
		\rEIP_reg[23]/NET0131 ,
		_w1080_,
		_w1081_,
		_w5431_
	);
	LUT4 #(
		.INIT('h8aff)
	) name4979 (
		_w690_,
		_w5421_,
		_w5430_,
		_w5431_,
		_w5432_
	);
	LUT3 #(
		.INIT('h08)
	) name4980 (
		\InstAddrPointer_reg[12]/NET0131 ,
		_w563_,
		_w673_,
		_w5433_
	);
	LUT4 #(
		.INIT('haa20)
	) name4981 (
		_w608_,
		_w5330_,
		_w5331_,
		_w5433_,
		_w5434_
	);
	LUT4 #(
		.INIT('hc6cc)
	) name4982 (
		\InstAddrPointer_reg[11]/NET0131 ,
		\InstAddrPointer_reg[12]/NET0131 ,
		READY_n_pad,
		_w726_,
		_w5435_
	);
	LUT4 #(
		.INIT('hec00)
	) name4983 (
		_w585_,
		_w589_,
		_w590_,
		_w5435_,
		_w5436_
	);
	LUT4 #(
		.INIT('haa8a)
	) name4984 (
		\InstAddrPointer_reg[12]/NET0131 ,
		_w613_,
		_w681_,
		_w5436_,
		_w5437_
	);
	LUT3 #(
		.INIT('hb0)
	) name4985 (
		_w616_,
		_w630_,
		_w951_,
		_w5438_
	);
	LUT3 #(
		.INIT('he0)
	) name4986 (
		_w588_,
		_w596_,
		_w5435_,
		_w5439_
	);
	LUT2 #(
		.INIT('h8)
	) name4987 (
		_w554_,
		_w886_,
		_w5440_
	);
	LUT3 #(
		.INIT('h07)
	) name4988 (
		_w635_,
		_w1042_,
		_w5440_,
		_w5441_
	);
	LUT2 #(
		.INIT('h4)
	) name4989 (
		_w5439_,
		_w5441_,
		_w5442_
	);
	LUT3 #(
		.INIT('h10)
	) name4990 (
		_w5438_,
		_w5437_,
		_w5442_,
		_w5443_
	);
	LUT2 #(
		.INIT('h4)
	) name4991 (
		_w5334_,
		_w5443_,
		_w5444_
	);
	LUT4 #(
		.INIT('h153f)
	) name4992 (
		\InstAddrPointer_reg[12]/NET0131 ,
		\rEIP_reg[12]/NET0131 ,
		_w1080_,
		_w1081_,
		_w5445_
	);
	LUT4 #(
		.INIT('h8aff)
	) name4993 (
		_w690_,
		_w5434_,
		_w5444_,
		_w5445_,
		_w5446_
	);
	LUT3 #(
		.INIT('h08)
	) name4994 (
		\PhyAddrPointer_reg[20]/NET0131 ,
		_w563_,
		_w673_,
		_w5447_
	);
	LUT4 #(
		.INIT('haa20)
	) name4995 (
		_w608_,
		_w5376_,
		_w5378_,
		_w5447_,
		_w5448_
	);
	LUT4 #(
		.INIT('h202a)
	) name4996 (
		\PhyAddrPointer_reg[20]/NET0131 ,
		_w634_,
		_w607_,
		_w608_,
		_w5449_
	);
	LUT3 #(
		.INIT('h0b)
	) name4997 (
		_w5380_,
		_w5381_,
		_w5449_,
		_w5450_
	);
	LUT4 #(
		.INIT('h60c0)
	) name4998 (
		\PhyAddrPointer_reg[1]/NET0131 ,
		\PhyAddrPointer_reg[20]/NET0131 ,
		_w1306_,
		_w1520_,
		_w5451_
	);
	LUT4 #(
		.INIT('h3f15)
	) name4999 (
		\PhyAddrPointer_reg[20]/NET0131 ,
		\rEIP_reg[20]/NET0131 ,
		_w1080_,
		_w1215_,
		_w5452_
	);
	LUT4 #(
		.INIT('hb700)
	) name5000 (
		\PhyAddrPointer_reg[20]/NET0131 ,
		_w714_,
		_w1520_,
		_w5452_,
		_w5453_
	);
	LUT2 #(
		.INIT('h4)
	) name5001 (
		_w5451_,
		_w5453_,
		_w5454_
	);
	LUT4 #(
		.INIT('h8aff)
	) name5002 (
		_w690_,
		_w5448_,
		_w5450_,
		_w5454_,
		_w5455_
	);
	LUT4 #(
		.INIT('h7774)
	) name5003 (
		\InstAddrPointer_reg[10]/NET0131 ,
		_w674_,
		_w1852_,
		_w1850_,
		_w5456_
	);
	LUT2 #(
		.INIT('h4)
	) name5004 (
		_w597_,
		_w1133_,
		_w5457_
	);
	LUT2 #(
		.INIT('h2)
	) name5005 (
		\InstAddrPointer_reg[10]/NET0131 ,
		_w1295_,
		_w5458_
	);
	LUT2 #(
		.INIT('h8)
	) name5006 (
		_w635_,
		_w1855_,
		_w5459_
	);
	LUT4 #(
		.INIT('h004f)
	) name5007 (
		_w616_,
		_w630_,
		_w953_,
		_w5459_,
		_w5460_
	);
	LUT3 #(
		.INIT('h10)
	) name5008 (
		_w5457_,
		_w5458_,
		_w5460_,
		_w5461_
	);
	LUT4 #(
		.INIT('h3100)
	) name5009 (
		_w608_,
		_w1857_,
		_w5456_,
		_w5461_,
		_w5462_
	);
	LUT4 #(
		.INIT('h153f)
	) name5010 (
		\InstAddrPointer_reg[10]/NET0131 ,
		\rEIP_reg[10]/NET0131 ,
		_w1080_,
		_w1081_,
		_w5463_
	);
	LUT3 #(
		.INIT('h2f)
	) name5011 (
		_w690_,
		_w5462_,
		_w5463_,
		_w5464_
	);
	LUT4 #(
		.INIT('h1555)
	) name5012 (
		_w1214_,
		_w3242_,
		_w3324_,
		_w3360_,
		_w5465_
	);
	LUT2 #(
		.INIT('h2)
	) name5013 (
		\DataWidth_reg[1]/NET0131 ,
		\rEIP_reg[30]/NET0131 ,
		_w5466_
	);
	LUT2 #(
		.INIT('h2)
	) name5014 (
		_w695_,
		_w5466_,
		_w5467_
	);
	LUT4 #(
		.INIT('hbe00)
	) name5015 (
		\DataWidth_reg[1]/NET0131 ,
		_w1304_,
		_w5465_,
		_w5467_,
		_w5468_
	);
	LUT4 #(
		.INIT('h0509)
	) name5016 (
		\EBX_reg[30]/NET0131 ,
		\EBX_reg[31]/NET0131 ,
		_w3116_,
		_w3350_,
		_w5469_
	);
	LUT4 #(
		.INIT('h4c8c)
	) name5017 (
		\rEIP_reg[30]/NET0131 ,
		_w2101_,
		_w3116_,
		_w3314_,
		_w5470_
	);
	LUT2 #(
		.INIT('h2)
	) name5018 (
		\rEIP_reg[30]/NET0131 ,
		_w3110_,
		_w5471_
	);
	LUT3 #(
		.INIT('h23)
	) name5019 (
		\DataWidth_reg[1]/NET0131 ,
		\EBX_reg[30]/NET0131 ,
		_w645_,
		_w5472_
	);
	LUT3 #(
		.INIT('h02)
	) name5020 (
		_w589_,
		_w566_,
		_w5472_,
		_w5473_
	);
	LUT4 #(
		.INIT('h7b00)
	) name5021 (
		\rEIP_reg[30]/NET0131 ,
		_w688_,
		_w3314_,
		_w5473_,
		_w5474_
	);
	LUT2 #(
		.INIT('h1)
	) name5022 (
		_w5471_,
		_w5474_,
		_w5475_
	);
	LUT4 #(
		.INIT('h20aa)
	) name5023 (
		_w690_,
		_w5469_,
		_w5470_,
		_w5475_,
		_w5476_
	);
	LUT4 #(
		.INIT('h5f13)
	) name5024 (
		\PhyAddrPointer_reg[30]/NET0131 ,
		\rEIP_reg[30]/NET0131 ,
		_w706_,
		_w3101_,
		_w5477_
	);
	LUT3 #(
		.INIT('hef)
	) name5025 (
		_w5476_,
		_w5468_,
		_w5477_,
		_w5478_
	);
	LUT3 #(
		.INIT('h08)
	) name5026 (
		\InstAddrPointer_reg[21]/NET0131 ,
		_w563_,
		_w673_,
		_w5479_
	);
	LUT4 #(
		.INIT('haa20)
	) name5027 (
		_w608_,
		_w1664_,
		_w1665_,
		_w5479_,
		_w5480_
	);
	LUT4 #(
		.INIT('hc6cc)
	) name5028 (
		\InstAddrPointer_reg[20]/NET0131 ,
		\InstAddrPointer_reg[21]/NET0131 ,
		READY_n_pad,
		_w733_,
		_w5481_
	);
	LUT4 #(
		.INIT('hec00)
	) name5029 (
		_w585_,
		_w589_,
		_w590_,
		_w5481_,
		_w5482_
	);
	LUT4 #(
		.INIT('haa8a)
	) name5030 (
		\InstAddrPointer_reg[21]/NET0131 ,
		_w613_,
		_w681_,
		_w5482_,
		_w5483_
	);
	LUT3 #(
		.INIT('hb0)
	) name5031 (
		_w616_,
		_w630_,
		_w966_,
		_w5484_
	);
	LUT2 #(
		.INIT('h8)
	) name5032 (
		_w635_,
		_w1056_,
		_w5485_
	);
	LUT2 #(
		.INIT('h8)
	) name5033 (
		_w554_,
		_w895_,
		_w5486_
	);
	LUT4 #(
		.INIT('h010f)
	) name5034 (
		_w588_,
		_w596_,
		_w5486_,
		_w5481_,
		_w5487_
	);
	LUT2 #(
		.INIT('h4)
	) name5035 (
		_w5485_,
		_w5487_,
		_w5488_
	);
	LUT3 #(
		.INIT('h10)
	) name5036 (
		_w5484_,
		_w5483_,
		_w5488_,
		_w5489_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name5037 (
		_w690_,
		_w1668_,
		_w5480_,
		_w5489_,
		_w5490_
	);
	LUT4 #(
		.INIT('h153f)
	) name5038 (
		\InstAddrPointer_reg[21]/NET0131 ,
		\rEIP_reg[21]/NET0131 ,
		_w1080_,
		_w1081_,
		_w5491_
	);
	LUT2 #(
		.INIT('hb)
	) name5039 (
		_w5490_,
		_w5491_,
		_w5492_
	);
	assign \_al_n0  = 1'b0;
	assign \_al_n1  = 1'b1;
	assign \g47406/_2_  = _w699_ ;
	assign \g47407/_2_  = _w709_ ;
	assign \g47411/_0_  = _w711_ ;
	assign \g47413/_0_  = _w717_ ;
	assign \g47424/_0_  = _w1083_ ;
	assign \g47434/_0_  = _w1129_ ;
	assign \g47437/_0_  = _w1172_ ;
	assign \g47447/_2_  = _w1219_ ;
	assign \g47448/_0_  = _w1233_ ;
	assign \g47451/_0_  = _w1253_ ;
	assign \g47452/_0_  = _w1283_ ;
	assign \g47453/_0_  = _w1300_ ;
	assign \g47465/_2_  = _w1311_ ;
	assign \g47466/_0_  = _w1331_ ;
	assign \g47467/_0_  = _w1356_ ;
	assign \g47471/_0_  = _w1377_ ;
	assign \g47485/_0_  = _w1394_ ;
	assign \g47486/_0_  = _w1411_ ;
	assign \g47487/_2_  = _w1422_ ;
	assign \g47488/_0_  = _w1442_ ;
	assign \g47489/_2_  = _w1452_ ;
	assign \g47491/_0_  = _w1464_ ;
	assign \g47494/_0_  = _w1486_ ;
	assign \g47510/_0_  = _w1496_ ;
	assign \g47511/_0_  = _w1507_ ;
	assign \g47512/_0_  = _w1527_ ;
	assign \g47515/_0_  = _w1538_ ;
	assign \g47516/_0_  = _w1550_ ;
	assign \g47517/_2_  = _w1561_ ;
	assign \g47524/_0_  = _w1581_ ;
	assign \g47525/_0_  = _w1594_ ;
	assign \g47550/_0_  = _w1607_ ;
	assign \g47551/_2_  = _w1627_ ;
	assign \g47552/_0_  = _w1646_ ;
	assign \g47554/_0_  = _w1662_ ;
	assign \g47555/_0_  = _w1678_ ;
	assign \g47556/_0_  = _w1691_ ;
	assign \g47558/_0_  = _w1701_ ;
	assign \g47563/_0_  = _w1722_ ;
	assign \g47564/_0_  = _w1739_ ;
	assign \g47565/_0_  = _w1843_ ;
	assign \g47584/_0_  = _w1849_ ;
	assign \g47592/_0_  = _w1864_ ;
	assign \g47597/_0_  = _w1873_ ;
	assign \g47598/_0_  = _w1883_ ;
	assign \g47601/_0_  = _w1902_ ;
	assign \g47602/_0_  = _w1915_ ;
	assign \g47603/_0_  = _w1964_ ;
	assign \g47604/_0_  = _w1970_ ;
	assign \g47606/_0_  = _w1998_ ;
	assign \g47630/_0_  = _w2004_ ;
	assign \g47636/_0_  = _w2016_ ;
	assign \g47641/_0_  = _w2033_ ;
	assign \g47642/_0_  = _w2047_ ;
	assign \g47643/_0_  = _w2062_ ;
	assign \g47644/_0_  = _w2069_ ;
	assign \g47645/_0_  = _w2083_ ;
	assign \g47646/_0_  = _w2105_ ;
	assign \g47648/_0_  = _w2114_ ;
	assign \g47679/_0_  = _w2126_ ;
	assign \g47680/_0_  = _w2137_ ;
	assign \g47681/_0_  = _w2148_ ;
	assign \g47683/_0_  = _w2154_ ;
	assign \g47687/_0_  = _w2168_ ;
	assign \g47690/_0_  = _w2173_ ;
	assign \g47746/_0_  = _w2182_ ;
	assign \g47747/_0_  = _w2188_ ;
	assign \g47754/_0_  = _w2194_ ;
	assign \g47756/_0_  = _w2198_ ;
	assign \g47804/_0_  = _w2231_ ;
	assign \g47805/_0_  = _w2248_ ;
	assign \g47806/_0_  = _w2262_ ;
	assign \g47807/_0_  = _w2275_ ;
	assign \g47809/_0_  = _w2287_ ;
	assign \g47810/_0_  = _w2298_ ;
	assign \g47812/_0_  = _w2310_ ;
	assign \g47813/_0_  = _w2323_ ;
	assign \g47814/_0_  = _w2336_ ;
	assign \g47815/_0_  = _w2349_ ;
	assign \g47816/_0_  = _w2362_ ;
	assign \g47817/_0_  = _w2375_ ;
	assign \g47818/_0_  = _w2388_ ;
	assign \g47819/_0_  = _w2400_ ;
	assign \g47820/_0_  = _w2411_ ;
	assign \g47821/_0_  = _w2422_ ;
	assign \g47836/_0_  = _w2430_ ;
	assign \g47848/_0_  = _w2439_ ;
	assign \g47851/_0_  = _w2447_ ;
	assign \g47852/_0_  = _w2461_ ;
	assign \g47943/_0_  = _w2473_ ;
	assign \g47944/_0_  = _w2483_ ;
	assign \g47945/_0_  = _w2493_ ;
	assign \g47946/_0_  = _w2503_ ;
	assign \g47947/_0_  = _w2513_ ;
	assign \g47949/_0_  = _w2523_ ;
	assign \g47950/_0_  = _w2533_ ;
	assign \g47952/_0_  = _w2543_ ;
	assign \g47953/_0_  = _w2553_ ;
	assign \g47954/_0_  = _w2563_ ;
	assign \g47955/_0_  = _w2573_ ;
	assign \g47956/_0_  = _w2583_ ;
	assign \g47957/_0_  = _w2593_ ;
	assign \g47958/_0_  = _w2603_ ;
	assign \g47959/_0_  = _w2613_ ;
	assign \g47960/_0_  = _w2623_ ;
	assign \g47999/_0_  = _w2628_ ;
	assign \g48/_0_  = _w2635_ ;
	assign \g48005/_0_  = _w2642_ ;
	assign \g48006/_0_  = _w2650_ ;
	assign \g48007/_0_  = _w2667_ ;
	assign \g48008/_0_  = _w2684_ ;
	assign \g48009/_0_  = _w2704_ ;
	assign \g48010/_0_  = _w2724_ ;
	assign \g48011/_0_  = _w2731_ ;
	assign \g48012/_0_  = _w2752_ ;
	assign \g48013/_0_  = _w2772_ ;
	assign \g48014/_0_  = _w2791_ ;
	assign \g48015/_0_  = _w2810_ ;
	assign \g48057/_0_  = _w2820_ ;
	assign \g48058/_0_  = _w2830_ ;
	assign \g48059/_0_  = _w2839_ ;
	assign \g48060/_0_  = _w2848_ ;
	assign \g48061/_0_  = _w2857_ ;
	assign \g48062/_0_  = _w2866_ ;
	assign \g48063/_0_  = _w2875_ ;
	assign \g48064/_0_  = _w2884_ ;
	assign \g48066/_0_  = _w2893_ ;
	assign \g48067/_0_  = _w2902_ ;
	assign \g48068/_0_  = _w2911_ ;
	assign \g48069/_0_  = _w2920_ ;
	assign \g48070/_0_  = _w2929_ ;
	assign \g48071/_0_  = _w2938_ ;
	assign \g48073/_0_  = _w2947_ ;
	assign \g48074/_0_  = _w2956_ ;
	assign \g48075/_0_  = _w2965_ ;
	assign \g48076/_0_  = _w2974_ ;
	assign \g48077/_0_  = _w2983_ ;
	assign \g48078/_0_  = _w2992_ ;
	assign \g48079/_0_  = _w3001_ ;
	assign \g48080/_0_  = _w3010_ ;
	assign \g48081/_0_  = _w3019_ ;
	assign \g48082/_0_  = _w3028_ ;
	assign \g48084/_0_  = _w3037_ ;
	assign \g48085/_0_  = _w3046_ ;
	assign \g48086/_0_  = _w3055_ ;
	assign \g48087/_0_  = _w3064_ ;
	assign \g48089/_0_  = _w3073_ ;
	assign \g48090/_0_  = _w3082_ ;
	assign \g48091/_0_  = _w3091_ ;
	assign \g48093/_0_  = _w3100_ ;
	assign \g48094/_0_  = _w3106_ ;
	assign \g48119/_0_  = _w3127_ ;
	assign \g48120/_0_  = _w3167_ ;
	assign \g48121/_0_  = _w3183_ ;
	assign \g48122/_0_  = _w3203_ ;
	assign \g48123/_0_  = _w3221_ ;
	assign \g48124/_0_  = _w3240_ ;
	assign \g48125/_0_  = _w3260_ ;
	assign \g48126/_0_  = _w3280_ ;
	assign \g48127/_0_  = _w3295_ ;
	assign \g48128/_0_  = _w3310_ ;
	assign \g48129/_0_  = _w3330_ ;
	assign \g48130/_0_  = _w3347_ ;
	assign \g48131/_0_  = _w3366_ ;
	assign \g48132/_0_  = _w3384_ ;
	assign \g48133/_0_  = _w3401_ ;
	assign \g48134/_0_  = _w3419_ ;
	assign \g48135/_0_  = _w3436_ ;
	assign \g48136/_0_  = _w3453_ ;
	assign \g48137/_0_  = _w3468_ ;
	assign \g48138/_0_  = _w3487_ ;
	assign \g48140/_0_  = _w3492_ ;
	assign \g48144/_0_  = _w3510_ ;
	assign \g48145/_0_  = _w3527_ ;
	assign \g48146/_0_  = _w3546_ ;
	assign \g48147/_0_  = _w3565_ ;
	assign \g48148/_0_  = _w3584_ ;
	assign \g48150/_0_  = _w3600_ ;
	assign \g48151/_0_  = _w3619_ ;
	assign \g48152/_0_  = _w3639_ ;
	assign \g48153/_0_  = _w3657_ ;
	assign \g48154/_0_  = _w3674_ ;
	assign \g48176/_0_  = _w3683_ ;
	assign \g48189/_0_  = _w3691_ ;
	assign \g48192/_0_  = _w3699_ ;
	assign \g48193/_0_  = _w3706_ ;
	assign \g48194/_0_  = _w3714_ ;
	assign \g48195/_0_  = _w3721_ ;
	assign \g48196/_0_  = _w3727_ ;
	assign \g48197/_0_  = _w3733_ ;
	assign \g48198/_0_  = _w3740_ ;
	assign \g48199/_0_  = _w3747_ ;
	assign \g48200/_0_  = _w3757_ ;
	assign \g48263/_0_  = _w3760_ ;
	assign \g48265/_0_  = _w3763_ ;
	assign \g48273/_0_  = _w3773_ ;
	assign \g48313/_0_  = _w3780_ ;
	assign \g48318/_0_  = _w3792_ ;
	assign \g48319/_0_  = _w3797_ ;
	assign \g48321/_0_  = _w3802_ ;
	assign \g48323/_0_  = _w3806_ ;
	assign \g48324/_0_  = _w3830_ ;
	assign \g48325/_0_  = _w3853_ ;
	assign \g48326/_0_  = _w3876_ ;
	assign \g48327/_0_  = _w3899_ ;
	assign \g48328/_0_  = _w3901_ ;
	assign \g48329/_0_  = _w3925_ ;
	assign \g48330/_0_  = _w3950_ ;
	assign \g48331/_0_  = _w3971_ ;
	assign \g48332/_0_  = _w3984_ ;
	assign \g48333/_0_  = _w4000_ ;
	assign \g48472/_0_  = _w4005_ ;
	assign \g48519/_0_  = _w4014_ ;
	assign \g48520/_0_  = _w4019_ ;
	assign \g48521/_0_  = _w4028_ ;
	assign \g48522/_0_  = _w4037_ ;
	assign \g48523/_0_  = _w4046_ ;
	assign \g48524/_0_  = _w4056_ ;
	assign \g48525/_0_  = _w4062_ ;
	assign \g48527/_0_  = _w4068_ ;
	assign \g48529/_0_  = _w4075_ ;
	assign \g48530/_0_  = _w4081_ ;
	assign \g48531/_0_  = _w4086_ ;
	assign \g48532/_0_  = _w4091_ ;
	assign \g48533/_0_  = _w4096_ ;
	assign \g48534/_0_  = _w4101_ ;
	assign \g48535/_0_  = _w4106_ ;
	assign \g48536/_0_  = _w4111_ ;
	assign \g48537/_0_  = _w4116_ ;
	assign \g48538/_0_  = _w4121_ ;
	assign \g48539/_0_  = _w4127_ ;
	assign \g48540/_0_  = _w4133_ ;
	assign \g48541/_0_  = _w4138_ ;
	assign \g48542/_0_  = _w4144_ ;
	assign \g48543/_0_  = _w4149_ ;
	assign \g48545/_0_  = _w4156_ ;
	assign \g48546/_0_  = _w4163_ ;
	assign \g48547/_0_  = _w4166_ ;
	assign \g48639/_0_  = _w4176_ ;
	assign \g48642/_0_  = _w4186_ ;
	assign \g48645/_0_  = _w4196_ ;
	assign \g48648/_0_  = _w4206_ ;
	assign \g48652/_0_  = _w4216_ ;
	assign \g48655/_0_  = _w4226_ ;
	assign \g48658/_0_  = _w4236_ ;
	assign \g48661/_0_  = _w4246_ ;
	assign \g48664/_0_  = _w4256_ ;
	assign \g48667/_0_  = _w4266_ ;
	assign \g48670/_0_  = _w4276_ ;
	assign \g48673/_0_  = _w4286_ ;
	assign \g48678/_0_  = _w4296_ ;
	assign \g48681/_0_  = _w4306_ ;
	assign \g48684/_0_  = _w4316_ ;
	assign \g48688/_0_  = _w4326_ ;
	assign \g48793/_0_  = _w4330_ ;
	assign \g48812/_0_  = _w4333_ ;
	assign \g48813/_0_  = _w4337_ ;
	assign \g48814/_0_  = _w4343_ ;
	assign \g48824/_0_  = _w4348_ ;
	assign \g48825/_0_  = _w4355_ ;
	assign \g48826/_0_  = _w4362_ ;
	assign \g48827/_0_  = _w4369_ ;
	assign \g48828/_0_  = _w4376_ ;
	assign \g48829/_0_  = _w4383_ ;
	assign \g48830/_0_  = _w4390_ ;
	assign \g48831/_0_  = _w4397_ ;
	assign \g48833/_0_  = _w4405_ ;
	assign \g48834/_0_  = _w4410_ ;
	assign \g48835/_0_  = _w4418_ ;
	assign \g48836/_0_  = _w4422_ ;
	assign \g48837/_0_  = _w4430_ ;
	assign \g48838/_0_  = _w4434_ ;
	assign \g48839/_0_  = _w4442_ ;
	assign \g48840/_0_  = _w4450_ ;
	assign \g48841/_0_  = _w4458_ ;
	assign \g48842/_0_  = _w4466_ ;
	assign \g48843/_0_  = _w4474_ ;
	assign \g48844/_0_  = _w4482_ ;
	assign \g48845/_0_  = _w4491_ ;
	assign \g48846/_0_  = _w4499_ ;
	assign \g48847/_0_  = _w4504_ ;
	assign \g48848/_0_  = _w4512_ ;
	assign \g48908/_0_  = _w4522_ ;
	assign \g48909/_0_  = _w4532_ ;
	assign \g48910/_0_  = _w4542_ ;
	assign \g48912/_0_  = _w4552_ ;
	assign \g48913/_0_  = _w4562_ ;
	assign \g48915/_0_  = _w4572_ ;
	assign \g48917/_0_  = _w4582_ ;
	assign \g48932/_0_  = _w4592_ ;
	assign \g48933/_0_  = _w4602_ ;
	assign \g48935/_0_  = _w4612_ ;
	assign \g48937/_0_  = _w4622_ ;
	assign \g48938/_0_  = _w4632_ ;
	assign \g48939/_0_  = _w4642_ ;
	assign \g48940/_0_  = _w4652_ ;
	assign \g48942/_0_  = _w4662_ ;
	assign \g48945/_0_  = _w4672_ ;
	assign \g48971/_0_  = _w4697_ ;
	assign \g49007/_0_  = _w4703_ ;
	assign \g49047/_0_  = _w4709_ ;
	assign \g49048/_0_  = _w4715_ ;
	assign \g49050/_0_  = _w4718_ ;
	assign \g49182/_0_  = _w4728_ ;
	assign \g49280/_0_  = _w4735_ ;
	assign \g49332/_0_  = _w4738_ ;
	assign \g49335/_0_  = _w4741_ ;
	assign \g49336/_0_  = _w4744_ ;
	assign \g49337/_0_  = _w4747_ ;
	assign \g49338/_0_  = _w4750_ ;
	assign \g49339/_0_  = _w4753_ ;
	assign \g49340/_0_  = _w4756_ ;
	assign \g49341/_0_  = _w4759_ ;
	assign \g49342/_0_  = _w4762_ ;
	assign \g49343/_0_  = _w4765_ ;
	assign \g49344/_0_  = _w4768_ ;
	assign \g49345/_0_  = _w4771_ ;
	assign \g49346/_0_  = _w4774_ ;
	assign \g49347/_0_  = _w4777_ ;
	assign \g49348/_0_  = _w4780_ ;
	assign \g49349/_0_  = _w4783_ ;
	assign \g49356/_0_  = _w4792_ ;
	assign \g49375/_0_  = _w4798_ ;
	assign \g49396/_0_  = _w4803_ ;
	assign \g49397/_0_  = _w4814_ ;
	assign \g49400/_0_  = _w4824_ ;
	assign \g49404/_0_  = _w4835_ ;
	assign \g49406/_0_  = _w4845_ ;
	assign \g49414/_0_  = _w4855_ ;
	assign \g49422/_0_  = _w4865_ ;
	assign \g49426/_0_  = _w4875_ ;
	assign \g49430/_0_  = _w4885_ ;
	assign \g49434/_0_  = _w4895_ ;
	assign \g49437/_0_  = _w4905_ ;
	assign \g49440/_0_  = _w4915_ ;
	assign \g49441/_0_  = _w4925_ ;
	assign \g49444/_0_  = _w4935_ ;
	assign \g49448/_0_  = _w4945_ ;
	assign \g49451/_0_  = _w4955_ ;
	assign \g49455/_0_  = _w4965_ ;
	assign \g49456/_0_  = _w4975_ ;
	assign \g49460/_0_  = _w4985_ ;
	assign \g49466/_0_  = _w4995_ ;
	assign \g49563/_0_  = _w5001_ ;
	assign \g49592/_0_  = _w5007_ ;
	assign \g49915/_0_  = _w5014_ ;
	assign \g49941/_0_  = _w5021_ ;
	assign \g50023/_0_  = _w5031_ ;
	assign \g50026/_0_  = _w5041_ ;
	assign \g50029/_0_  = _w5051_ ;
	assign \g50031/_0_  = _w5061_ ;
	assign \g50033/_0_  = _w5071_ ;
	assign \g50035/_0_  = _w5081_ ;
	assign \g50037/_0_  = _w5091_ ;
	assign \g50040/_0_  = _w5101_ ;
	assign \g50050/_0_  = _w5111_ ;
	assign \g50056/_0_  = _w5121_ ;
	assign \g50059/_0_  = _w5131_ ;
	assign \g50065/_0_  = _w5141_ ;
	assign \g50067/_0_  = _w5151_ ;
	assign \g50150/_0_  = _w5156_ ;
	assign \g50283/_0_  = _w5160_ ;
	assign \g50284/_0_  = _w5166_ ;
	assign \g50501/_0_  = _w5170_ ;
	assign \g50594/_0_  = _w5177_ ;
	assign \g50807/_0_  = _w5184_ ;
	assign \g50866/_0_  = _w5190_ ;
	assign \g50875/_0_  = _w5197_ ;
	assign \g51449/_0_  = _w5203_ ;
	assign \g51510/_0_  = _w5207_ ;
	assign \g51534/_0_  = _w5211_ ;
	assign \g52310/_0_  = _w5216_ ;
	assign \g53066/_0_  = _w5220_ ;
	assign \g53087/_0_  = _w5225_ ;
	assign \g53151/_0_  = _w5230_ ;
	assign \g53608/_0_  = _w5235_ ;
	assign \g53634/_0_  = _w5241_ ;
	assign \g54053/_0_  = _w5246_ ;
	assign \g54091/_0_  = _w5251_ ;
	assign \g54103/_0_  = _w5256_ ;
	assign \g54268/_0_  = _w5260_ ;
	assign \g54277/_0_  = _w5263_ ;
	assign \g54287/_0_  = _w5266_ ;
	assign \g54294/_0_  = _w5270_ ;
	assign \g54449/_0_  = _w5274_ ;
	assign \g54453/_0_  = _w5279_ ;
	assign \g54484/_0_  = _w5286_ ;
	assign \g54528/_0_  = _w5294_ ;
	assign \g54582/_0_  = _w5297_ ;
	assign \g55448/_0_  = _w5301_ ;
	assign \g55693/_1_  = _w5257_ ;
	assign \g55874/_0_  = _w5304_ ;
	assign \g56203/_0_  = _w5305_ ;
	assign \g56303/_0_  = _w5306_ ;
	assign \g56329/_0_  = _w5307_ ;
	assign \g56336/_0_  = _w5308_ ;
	assign \g56345/_0_  = _w5309_ ;
	assign \g56367/_0_  = _w5310_ ;
	assign \g56411/_0_  = _w5311_ ;
	assign \g56529/_0_  = _w5314_ ;
	assign \g56858/_0_  = _w5316_ ;
	assign \g60443/_1_  = _w4673_ ;
	assign \g63395/_0_  = _w5327_ ;
	assign \g63442/_0_  = _w5343_ ;
	assign \g63595/_0_  = _w5352_ ;
	assign \g63996/_0_  = _w5363_ ;
	assign \g64048/_0_  = _w5373_ ;
	assign \g64071/_0_  = _w5398_ ;
	assign \g64085/_0_  = _w5407_ ;
	assign \g64096/_0_  = _w5419_ ;
	assign \g64119/_0_  = _w5432_ ;
	assign \g64216/_0_  = _w5446_ ;
	assign \g64513/_0_  = _w5455_ ;
	assign \g64566/_0_  = _w5464_ ;
	assign \g64694/_0_  = _w5478_ ;
	assign \g64913/_0_  = _w5492_ ;
endmodule;