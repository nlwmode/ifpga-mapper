module top( CLR_pad , \v0_pad  , \v10_reg/NET0131  , \v11_reg/NET0131  , \v12_reg/NET0131  , \v1_pad  , \v2_pad  , \v3_pad  , \v4_pad  , \v5_pad  , \v6_pad  , \v7_reg/NET0131  , \v8_reg/NET0131  , \v9_reg/NET0131  , \_al_n0  , \_al_n1  , \g1759/_1_  , \g1762/_1_  , \g1764/_1_  , \g1765/_0_  , \g1786/_2_  , \g1791/_3_  , \g1808/_3_  , \g1822/_2_  , \g1929/_3_  , \g2713/_1_  , \g2744/_0_  , \v13_D_11_pad  , \v13_D_12_pad  , \v13_D_13_pad  , \v13_D_14_pad  , \v13_D_16_pad  , \v13_D_18_pad  , \v13_D_19_pad  , \v13_D_21_pad  , \v13_D_22_pad  , \v13_D_23_pad  , \v13_D_24_pad  , \v13_D_7_pad  , \v13_D_8_pad  , \v13_D_9_pad  );
  input CLR_pad ;
  input \v0_pad  ;
  input \v10_reg/NET0131  ;
  input \v11_reg/NET0131  ;
  input \v12_reg/NET0131  ;
  input \v1_pad  ;
  input \v2_pad  ;
  input \v3_pad  ;
  input \v4_pad  ;
  input \v5_pad  ;
  input \v6_pad  ;
  input \v7_reg/NET0131  ;
  input \v8_reg/NET0131  ;
  input \v9_reg/NET0131  ;
  output \_al_n0  ;
  output \_al_n1  ;
  output \g1759/_1_  ;
  output \g1762/_1_  ;
  output \g1764/_1_  ;
  output \g1765/_0_  ;
  output \g1786/_2_  ;
  output \g1791/_3_  ;
  output \g1808/_3_  ;
  output \g1822/_2_  ;
  output \g1929/_3_  ;
  output \g2713/_1_  ;
  output \g2744/_0_  ;
  output \v13_D_11_pad  ;
  output \v13_D_12_pad  ;
  output \v13_D_13_pad  ;
  output \v13_D_14_pad  ;
  output \v13_D_16_pad  ;
  output \v13_D_18_pad  ;
  output \v13_D_19_pad  ;
  output \v13_D_21_pad  ;
  output \v13_D_22_pad  ;
  output \v13_D_23_pad  ;
  output \v13_D_24_pad  ;
  output \v13_D_7_pad  ;
  output \v13_D_8_pad  ;
  output \v13_D_9_pad  ;
  wire n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 ;
  assign n15 = ~\v0_pad  & \v10_reg/NET0131  ;
  assign n16 = ~\v12_reg/NET0131  & ~\v9_reg/NET0131  ;
  assign n17 = \v4_pad  & \v5_pad  ;
  assign n18 = n16 & n17 ;
  assign n19 = \v11_reg/NET0131  & \v12_reg/NET0131  ;
  assign n20 = \v8_reg/NET0131  & n19 ;
  assign n21 = ~\v1_pad  & \v6_pad  ;
  assign n22 = \v3_pad  & n21 ;
  assign n23 = n20 & n22 ;
  assign n24 = ~n18 & ~n23 ;
  assign n25 = n15 & ~n24 ;
  assign n39 = \v6_pad  & ~\v8_reg/NET0131  ;
  assign n40 = \v12_reg/NET0131  & ~\v9_reg/NET0131  ;
  assign n41 = ~\v10_reg/NET0131  & n40 ;
  assign n42 = ~\v11_reg/NET0131  & n41 ;
  assign n43 = n39 & n42 ;
  assign n36 = \v10_reg/NET0131  & \v11_reg/NET0131  ;
  assign n37 = ~\v8_reg/NET0131  & n36 ;
  assign n38 = \v9_reg/NET0131  & n37 ;
  assign n44 = \v10_reg/NET0131  & ~\v9_reg/NET0131  ;
  assign n45 = ~\v11_reg/NET0131  & ~\v12_reg/NET0131  ;
  assign n46 = n44 & n45 ;
  assign n55 = ~n38 & ~n46 ;
  assign n56 = ~n43 & n55 ;
  assign n57 = ~n25 & n56 ;
  assign n26 = \v12_reg/NET0131  & \v3_pad  ;
  assign n27 = \v0_pad  & \v11_reg/NET0131  ;
  assign n28 = \v10_reg/NET0131  & \v8_reg/NET0131  ;
  assign n29 = ~n21 & n28 ;
  assign n30 = n27 & n29 ;
  assign n31 = ~\v11_reg/NET0131  & ~\v8_reg/NET0131  ;
  assign n32 = ~\v9_reg/NET0131  & n31 ;
  assign n33 = ~\v10_reg/NET0131  & n32 ;
  assign n34 = ~n30 & ~n33 ;
  assign n35 = n26 & ~n34 ;
  assign n48 = \v11_reg/NET0131  & ~\v12_reg/NET0131  ;
  assign n49 = \v10_reg/NET0131  & ~\v2_pad  ;
  assign n50 = ~n17 & n49 ;
  assign n51 = n48 & ~n50 ;
  assign n52 = \v9_reg/NET0131  & ~n51 ;
  assign n47 = ~\v10_reg/NET0131  & ~\v9_reg/NET0131  ;
  assign n53 = \v8_reg/NET0131  & ~n47 ;
  assign n54 = ~n52 & n53 ;
  assign n58 = ~n35 & ~n54 ;
  assign n59 = n57 & n58 ;
  assign n60 = ~\v7_reg/NET0131  & ~n59 ;
  assign n64 = \v10_reg/NET0131  & \v9_reg/NET0131  ;
  assign n65 = n48 & n64 ;
  assign n66 = \v7_reg/NET0131  & n65 ;
  assign n61 = ~\v2_pad  & \v8_reg/NET0131  ;
  assign n62 = ~\v9_reg/NET0131  & n36 ;
  assign n63 = n61 & n62 ;
  assign n67 = n16 & n28 ;
  assign n82 = ~n63 & ~n67 ;
  assign n83 = ~n66 & n82 ;
  assign n68 = ~\v10_reg/NET0131  & \v7_reg/NET0131  ;
  assign n69 = ~\v11_reg/NET0131  & \v8_reg/NET0131  ;
  assign n70 = ~n16 & n69 ;
  assign n71 = \v11_reg/NET0131  & ~\v8_reg/NET0131  ;
  assign n72 = ~\v12_reg/NET0131  & n71 ;
  assign n73 = ~n70 & ~n72 ;
  assign n74 = n68 & ~n73 ;
  assign n76 = ~\v12_reg/NET0131  & \v9_reg/NET0131  ;
  assign n77 = ~\v7_reg/NET0131  & n76 ;
  assign n75 = ~\v10_reg/NET0131  & ~\v11_reg/NET0131  ;
  assign n78 = \v1_pad  & ~\v2_pad  ;
  assign n79 = n39 & n78 ;
  assign n80 = n75 & n79 ;
  assign n81 = n77 & n80 ;
  assign n84 = ~n74 & ~n81 ;
  assign n85 = n83 & n84 ;
  assign n86 = ~n60 & n85 ;
  assign n87 = CLR_pad & ~n86 ;
  assign n101 = \v10_reg/NET0131  & ~\v12_reg/NET0131  ;
  assign n102 = ~\v11_reg/NET0131  & n101 ;
  assign n103 = \v9_reg/NET0131  & ~n102 ;
  assign n96 = ~n36 & ~n75 ;
  assign n97 = \v12_reg/NET0131  & n96 ;
  assign n98 = \v12_reg/NET0131  & ~\v6_pad  ;
  assign n99 = ~\v3_pad  & n98 ;
  assign n100 = ~\v10_reg/NET0131  & n99 ;
  assign n104 = ~n97 & ~n100 ;
  assign n105 = ~n103 & n104 ;
  assign n88 = ~\v12_reg/NET0131  & n17 ;
  assign n89 = ~\v0_pad  & n36 ;
  assign n90 = ~n75 & ~n89 ;
  assign n91 = n88 & ~n90 ;
  assign n92 = \v10_reg/NET0131  & \v12_reg/NET0131  ;
  assign n93 = ~\v3_pad  & n92 ;
  assign n94 = ~\v9_reg/NET0131  & ~n93 ;
  assign n95 = \v2_pad  & ~n94 ;
  assign n106 = ~n91 & ~n95 ;
  assign n107 = n105 & n106 ;
  assign n108 = ~\v8_reg/NET0131  & ~n107 ;
  assign n109 = ~\v10_reg/NET0131  & ~\v1_pad  ;
  assign n110 = \v2_pad  & n109 ;
  assign n111 = ~\v9_reg/NET0131  & ~n110 ;
  assign n112 = n19 & ~n111 ;
  assign n113 = ~\v12_reg/NET0131  & \v8_reg/NET0131  ;
  assign n114 = n47 & n113 ;
  assign n115 = ~n112 & ~n114 ;
  assign n116 = ~n108 & n115 ;
  assign n117 = ~\v7_reg/NET0131  & ~n116 ;
  assign n122 = \v10_reg/NET0131  & n48 ;
  assign n136 = ~\v8_reg/NET0131  & ~\v9_reg/NET0131  ;
  assign n137 = n122 & ~n136 ;
  assign n133 = ~\v10_reg/NET0131  & \v8_reg/NET0131  ;
  assign n134 = \v11_reg/NET0131  & ~n40 ;
  assign n135 = n133 & ~n134 ;
  assign n138 = ~\v10_reg/NET0131  & ~\v8_reg/NET0131  ;
  assign n139 = n48 & n138 ;
  assign n140 = ~n135 & ~n139 ;
  assign n141 = ~n137 & n140 ;
  assign n142 = \v7_reg/NET0131  & ~n141 ;
  assign n127 = \v12_reg/NET0131  & \v1_pad  ;
  assign n128 = ~\v10_reg/NET0131  & n127 ;
  assign n129 = n17 & n113 ;
  assign n130 = ~n128 & ~n129 ;
  assign n126 = ~\v2_pad  & ~\v7_reg/NET0131  ;
  assign n131 = \v11_reg/NET0131  & n126 ;
  assign n132 = ~n130 & n131 ;
  assign n118 = ~\v10_reg/NET0131  & ~\v12_reg/NET0131  ;
  assign n119 = \v3_pad  & n118 ;
  assign n120 = ~n40 & ~n119 ;
  assign n121 = n69 & ~n120 ;
  assign n123 = \v7_reg/NET0131  & n40 ;
  assign n124 = ~n122 & ~n123 ;
  assign n125 = n61 & ~n124 ;
  assign n143 = ~n121 & ~n125 ;
  assign n144 = ~n132 & n143 ;
  assign n145 = ~n142 & n144 ;
  assign n146 = ~n117 & n145 ;
  assign n147 = CLR_pad & ~n146 ;
  assign n150 = n31 & n76 ;
  assign n151 = n19 & n61 ;
  assign n152 = ~n150 & ~n151 ;
  assign n153 = ~\v1_pad  & ~n152 ;
  assign n148 = ~\v11_reg/NET0131  & \v3_pad  ;
  assign n149 = n113 & n148 ;
  assign n154 = ~\v6_pad  & \v9_reg/NET0131  ;
  assign n155 = n45 & n154 ;
  assign n156 = ~\v8_reg/NET0131  & n155 ;
  assign n157 = ~n149 & ~n156 ;
  assign n158 = ~n153 & n157 ;
  assign n159 = ~\v10_reg/NET0131  & ~n158 ;
  assign n171 = ~\v9_reg/NET0131  & ~n92 ;
  assign n172 = ~\v8_reg/NET0131  & ~n118 ;
  assign n173 = n171 & n172 ;
  assign n174 = n90 & n173 ;
  assign n175 = n18 & n75 ;
  assign n176 = \v8_reg/NET0131  & \v9_reg/NET0131  ;
  assign n177 = \v12_reg/NET0131  & ~n36 ;
  assign n178 = n176 & n177 ;
  assign n184 = ~n175 & ~n178 ;
  assign n179 = ~\v11_reg/NET0131  & n92 ;
  assign n180 = \v9_reg/NET0131  & n179 ;
  assign n181 = \v10_reg/NET0131  & ~\v11_reg/NET0131  ;
  assign n182 = \v2_pad  & n181 ;
  assign n183 = n16 & n182 ;
  assign n185 = ~n180 & ~n183 ;
  assign n186 = n184 & n185 ;
  assign n187 = ~n174 & n186 ;
  assign n160 = ~\v10_reg/NET0131  & n150 ;
  assign n161 = \v11_reg/NET0131  & n133 ;
  assign n162 = ~\v9_reg/NET0131  & ~n127 ;
  assign n163 = n161 & ~n162 ;
  assign n164 = ~n160 & ~n163 ;
  assign n165 = \v2_pad  & ~n164 ;
  assign n166 = ~\v12_reg/NET0131  & ~\v8_reg/NET0131  ;
  assign n167 = n44 & n166 ;
  assign n168 = \v9_reg/NET0131  & n161 ;
  assign n169 = ~n167 & ~n168 ;
  assign n170 = ~n17 & ~n169 ;
  assign n188 = ~n165 & ~n170 ;
  assign n189 = n187 & n188 ;
  assign n190 = ~n159 & n189 ;
  assign n191 = ~\v7_reg/NET0131  & ~n190 ;
  assign n192 = \v7_reg/NET0131  & \v8_reg/NET0131  ;
  assign n193 = ~n75 & n192 ;
  assign n194 = \v2_pad  & n36 ;
  assign n195 = ~\v9_reg/NET0131  & ~n194 ;
  assign n196 = \v12_reg/NET0131  & ~n195 ;
  assign n197 = n193 & ~n196 ;
  assign n203 = ~\v7_reg/NET0131  & ~\v8_reg/NET0131  ;
  assign n204 = n47 & n203 ;
  assign n205 = n99 & n204 ;
  assign n198 = \v11_reg/NET0131  & \v3_pad  ;
  assign n199 = n114 & ~n198 ;
  assign n200 = ~\v12_reg/NET0131  & \v7_reg/NET0131  ;
  assign n201 = \v11_reg/NET0131  & ~n44 ;
  assign n202 = n200 & n201 ;
  assign n206 = ~n199 & ~n202 ;
  assign n207 = ~n205 & n206 ;
  assign n208 = ~n197 & n207 ;
  assign n209 = ~n191 & n208 ;
  assign n210 = CLR_pad & ~n209 ;
  assign n211 = \v2_pad  & n77 ;
  assign n212 = ~n19 & ~n31 ;
  assign n213 = ~n113 & ~n136 ;
  assign n214 = n212 & n213 ;
  assign n215 = ~n211 & ~n214 ;
  assign n216 = ~\v10_reg/NET0131  & ~n215 ;
  assign n227 = ~\v9_reg/NET0131  & n98 ;
  assign n228 = ~n92 & ~n227 ;
  assign n229 = ~\v11_reg/NET0131  & ~n228 ;
  assign n217 = \v9_reg/NET0131  & n109 ;
  assign n218 = ~n62 & ~n217 ;
  assign n219 = n166 & ~n218 ;
  assign n224 = ~\v3_pad  & ~\v9_reg/NET0131  ;
  assign n225 = n48 & ~n224 ;
  assign n226 = n133 & ~n225 ;
  assign n238 = ~\v7_reg/NET0131  & ~n226 ;
  assign n241 = ~n219 & n238 ;
  assign n242 = ~n229 & n241 ;
  assign n220 = ~\v12_reg/NET0131  & n176 ;
  assign n221 = n17 & n220 ;
  assign n222 = ~n67 & ~n221 ;
  assign n223 = ~\v2_pad  & ~n222 ;
  assign n235 = ~\v8_reg/NET0131  & \v9_reg/NET0131  ;
  assign n236 = ~\v6_pad  & n118 ;
  assign n237 = n235 & n236 ;
  assign n230 = \v0_pad  & n21 ;
  assign n231 = n26 & n176 ;
  assign n232 = ~n230 & n231 ;
  assign n233 = \v9_reg/NET0131  & ~n48 ;
  assign n234 = n96 & n233 ;
  assign n239 = ~n232 & ~n234 ;
  assign n240 = ~n237 & n239 ;
  assign n243 = ~n223 & n240 ;
  assign n244 = n242 & n243 ;
  assign n248 = ~\v12_reg/NET0131  & ~n31 ;
  assign n247 = \v11_reg/NET0131  & ~n138 ;
  assign n249 = ~n64 & ~n133 ;
  assign n250 = ~n247 & n249 ;
  assign n251 = n248 & n250 ;
  assign n245 = \v2_pad  & n44 ;
  assign n246 = n20 & n245 ;
  assign n252 = \v7_reg/NET0131  & ~n246 ;
  assign n253 = ~n251 & n252 ;
  assign n254 = ~n244 & ~n253 ;
  assign n255 = ~n216 & ~n254 ;
  assign n256 = CLR_pad & ~n255 ;
  assign n257 = \v12_reg/NET0131  & n44 ;
  assign n258 = ~\v12_reg/NET0131  & ~n47 ;
  assign n259 = ~n126 & n258 ;
  assign n260 = ~n257 & ~n259 ;
  assign n261 = \v11_reg/NET0131  & ~n260 ;
  assign n262 = ~n118 & ~n171 ;
  assign n263 = ~\v11_reg/NET0131  & \v7_reg/NET0131  ;
  assign n264 = ~n262 & n263 ;
  assign n265 = ~n261 & ~n264 ;
  assign n266 = \v8_reg/NET0131  & ~n265 ;
  assign n274 = \v8_reg/NET0131  & ~n182 ;
  assign n273 = ~\v7_reg/NET0131  & ~\v9_reg/NET0131  ;
  assign n275 = ~n27 & ~n181 ;
  assign n276 = n273 & ~n275 ;
  assign n277 = ~n274 & n276 ;
  assign n267 = ~n47 & ~n64 ;
  assign n268 = n71 & ~n267 ;
  assign n269 = \v11_reg/NET0131  & \v9_reg/NET0131  ;
  assign n270 = ~n203 & ~n269 ;
  assign n271 = n17 & ~n235 ;
  assign n272 = ~n270 & n271 ;
  assign n278 = ~n268 & ~n272 ;
  assign n279 = ~n277 & n278 ;
  assign n280 = ~\v12_reg/NET0131  & ~n279 ;
  assign n281 = ~n266 & ~n280 ;
  assign n282 = n175 & n203 ;
  assign n283 = \v12_reg/NET0131  & ~n62 ;
  assign n284 = \v8_reg/NET0131  & ~n283 ;
  assign n285 = ~\v10_reg/NET0131  & n48 ;
  assign n286 = ~n284 & ~n285 ;
  assign n287 = \v7_reg/NET0131  & ~n286 ;
  assign n288 = ~n27 & n273 ;
  assign n289 = ~n269 & ~n288 ;
  assign n290 = \v10_reg/NET0131  & ~n289 ;
  assign n291 = \v11_reg/NET0131  & \v8_reg/NET0131  ;
  assign n292 = ~n47 & n291 ;
  assign n293 = ~n290 & ~n292 ;
  assign n294 = ~\v12_reg/NET0131  & ~n293 ;
  assign n295 = ~n287 & ~n294 ;
  assign n296 = \v2_pad  & ~n295 ;
  assign n297 = ~n282 & ~n296 ;
  assign n298 = ~\v4_pad  & \v5_pad  ;
  assign n299 = ~\v10_reg/NET0131  & ~n298 ;
  assign n300 = ~\v9_reg/NET0131  & ~n299 ;
  assign n301 = ~n247 & ~n300 ;
  assign n302 = ~\v12_reg/NET0131  & ~n301 ;
  assign n303 = \v11_reg/NET0131  & n47 ;
  assign n304 = ~n302 & ~n303 ;
  assign n305 = \v11_reg/NET0131  & ~\v2_pad  ;
  assign n306 = \v9_reg/NET0131  & n305 ;
  assign n307 = n274 & ~n306 ;
  assign n308 = ~n304 & ~n307 ;
  assign n309 = ~\v7_reg/NET0131  & ~n308 ;
  assign n312 = \v7_reg/NET0131  & n47 ;
  assign n313 = ~\v12_reg/NET0131  & ~n312 ;
  assign n310 = \v9_reg/NET0131  & ~n75 ;
  assign n311 = \v8_reg/NET0131  & ~n310 ;
  assign n314 = ~n42 & n311 ;
  assign n315 = ~n313 & n314 ;
  assign n316 = ~n309 & ~n315 ;
  assign n317 = ~n90 & n136 ;
  assign n318 = n176 & n305 ;
  assign n319 = ~n317 & ~n318 ;
  assign n320 = ~\v12_reg/NET0131  & ~\v7_reg/NET0131  ;
  assign n321 = \v4_pad  & ~\v5_pad  ;
  assign n322 = n320 & n321 ;
  assign n323 = ~n319 & n322 ;
  assign n324 = n26 & n269 ;
  assign n325 = ~\v7_reg/NET0131  & n29 ;
  assign n326 = n324 & n325 ;
  assign n342 = ~\v12_reg/NET0131  & \v1_pad  ;
  assign n343 = ~n21 & n36 ;
  assign n344 = ~n342 & ~n343 ;
  assign n345 = \v3_pad  & ~n344 ;
  assign n346 = n31 & n92 ;
  assign n347 = \v9_reg/NET0131  & ~n248 ;
  assign n348 = ~n346 & n347 ;
  assign n349 = ~n345 & n348 ;
  assign n333 = n15 & n136 ;
  assign n334 = n88 & n333 ;
  assign n335 = ~\v8_reg/NET0131  & ~n101 ;
  assign n336 = \v9_reg/NET0131  & n335 ;
  assign n337 = ~n334 & ~n336 ;
  assign n338 = \v11_reg/NET0131  & ~n337 ;
  assign n339 = n76 & n181 ;
  assign n340 = ~n155 & ~n339 ;
  assign n341 = ~\v8_reg/NET0131  & ~n340 ;
  assign n350 = ~n338 & ~n341 ;
  assign n351 = ~n349 & n350 ;
  assign n352 = ~\v7_reg/NET0131  & ~n351 ;
  assign n327 = n17 & n291 ;
  assign n328 = ~n31 & ~n327 ;
  assign n329 = n77 & ~n328 ;
  assign n330 = n40 & n192 ;
  assign n331 = ~n329 & ~n330 ;
  assign n332 = ~\v2_pad  & ~n331 ;
  assign n353 = ~n16 & n192 ;
  assign n354 = ~n62 & n353 ;
  assign n355 = ~n310 & n354 ;
  assign n356 = ~n332 & ~n355 ;
  assign n357 = ~n352 & n356 ;
  assign n358 = CLR_pad & ~n357 ;
  assign n359 = ~\v12_reg/NET0131  & \v2_pad  ;
  assign n360 = ~\v11_reg/NET0131  & ~n359 ;
  assign n361 = \v10_reg/NET0131  & ~n360 ;
  assign n362 = ~\v9_reg/NET0131  & ~n361 ;
  assign n365 = ~n230 & n324 ;
  assign n363 = n17 & ~n19 ;
  assign n364 = ~\v10_reg/NET0131  & ~n363 ;
  assign n366 = ~n155 & ~n364 ;
  assign n367 = ~n365 & n366 ;
  assign n368 = ~n362 & n367 ;
  assign n369 = \v8_reg/NET0131  & ~n368 ;
  assign n370 = ~\v10_reg/NET0131  & \v12_reg/NET0131  ;
  assign n371 = ~n220 & ~n370 ;
  assign n372 = ~\v3_pad  & ~n371 ;
  assign n373 = ~\v10_reg/NET0131  & n18 ;
  assign n374 = ~n372 & ~n373 ;
  assign n375 = ~\v11_reg/NET0131  & ~n374 ;
  assign n380 = ~\v11_reg/NET0131  & \v6_pad  ;
  assign n381 = ~\v9_reg/NET0131  & ~n380 ;
  assign n382 = \v12_reg/NET0131  & n138 ;
  assign n383 = ~n381 & n382 ;
  assign n376 = n37 & n40 ;
  assign n377 = \v10_reg/NET0131  & ~n235 ;
  assign n378 = ~n138 & n359 ;
  assign n379 = ~n377 & n378 ;
  assign n384 = ~n376 & ~n379 ;
  assign n385 = ~n383 & n384 ;
  assign n386 = ~n375 & n385 ;
  assign n387 = ~n369 & n386 ;
  assign n388 = ~\v7_reg/NET0131  & ~n387 ;
  assign n389 = n200 & n269 ;
  assign n390 = \v10_reg/NET0131  & ~n40 ;
  assign n391 = ~n41 & n69 ;
  assign n392 = ~n390 & n391 ;
  assign n393 = ~n389 & ~n392 ;
  assign n394 = ~n388 & n393 ;
  assign n395 = CLR_pad & ~n394 ;
  assign n396 = \v3_pad  & n380 ;
  assign n397 = ~n305 & ~n396 ;
  assign n398 = \v8_reg/NET0131  & ~n397 ;
  assign n399 = n136 & n275 ;
  assign n400 = ~n398 & ~n399 ;
  assign n401 = n17 & ~n69 ;
  assign n402 = ~\v12_reg/NET0131  & ~n401 ;
  assign n403 = ~n400 & n402 ;
  assign n404 = ~\v7_reg/NET0131  & ~n403 ;
  assign n405 = ~n139 & ~n311 ;
  assign n406 = ~n404 & n405 ;
  assign n407 = ~\v10_reg/NET0131  & n17 ;
  assign n408 = ~n27 & ~n407 ;
  assign n409 = ~\v12_reg/NET0131  & ~n408 ;
  assign n410 = ~n179 & ~n409 ;
  assign n411 = ~\v9_reg/NET0131  & ~n410 ;
  assign n412 = ~n65 & ~n411 ;
  assign n413 = ~\v7_reg/NET0131  & ~n412 ;
  assign n414 = ~\v9_reg/NET0131  & n285 ;
  assign n415 = ~n413 & ~n414 ;
  assign n416 = ~\v8_reg/NET0131  & ~n415 ;
  assign n417 = ~n47 & n359 ;
  assign n418 = ~n257 & ~n417 ;
  assign n419 = \v11_reg/NET0131  & ~n418 ;
  assign n420 = ~n200 & ~n419 ;
  assign n421 = \v8_reg/NET0131  & ~n420 ;
  assign n422 = ~n416 & ~n421 ;
  assign n423 = ~n291 & ~n320 ;
  assign n424 = ~\v1_pad  & ~n423 ;
  assign n425 = ~n20 & ~n424 ;
  assign n426 = ~\v9_reg/NET0131  & ~n425 ;
  assign n427 = \v9_reg/NET0131  & n48 ;
  assign n428 = \v1_pad  & n427 ;
  assign n429 = ~n426 & ~n428 ;
  assign n430 = \v10_reg/NET0131  & ~n429 ;
  assign n431 = ~n19 & n47 ;
  assign n432 = ~n339 & ~n431 ;
  assign n433 = \v8_reg/NET0131  & ~n432 ;
  assign n434 = \v7_reg/NET0131  & ~n139 ;
  assign n435 = ~n433 & n434 ;
  assign n436 = \v11_reg/NET0131  & ~n15 ;
  assign n437 = n136 & ~n436 ;
  assign n438 = ~n318 & ~n437 ;
  assign n439 = n17 & ~n438 ;
  assign n440 = \v2_pad  & n292 ;
  assign n441 = ~n439 & ~n440 ;
  assign n442 = ~\v12_reg/NET0131  & ~n441 ;
  assign n443 = ~n45 & ~n172 ;
  assign n444 = ~\v9_reg/NET0131  & n96 ;
  assign n445 = ~n443 & n444 ;
  assign n446 = ~\v7_reg/NET0131  & ~n445 ;
  assign n447 = ~n442 & n446 ;
  assign n448 = ~n435 & ~n447 ;
  assign n449 = ~n430 & ~n448 ;
  assign n452 = ~\v9_reg/NET0131  & ~n436 ;
  assign n453 = ~\v8_reg/NET0131  & ~n452 ;
  assign n456 = ~\v12_reg/NET0131  & ~n17 ;
  assign n455 = \v2_pad  & \v8_reg/NET0131  ;
  assign n454 = ~\v4_pad  & ~\v5_pad  ;
  assign n457 = ~n181 & ~n454 ;
  assign n458 = ~n455 & n457 ;
  assign n459 = n456 & n458 ;
  assign n460 = ~n453 & n459 ;
  assign n461 = ~\v7_reg/NET0131  & ~n460 ;
  assign n450 = ~n200 & n310 ;
  assign n451 = \v8_reg/NET0131  & ~n450 ;
  assign n462 = ~n202 & ~n451 ;
  assign n463 = ~n461 & n462 ;
  assign n464 = n77 & n396 ;
  assign n465 = \v11_reg/NET0131  & \v2_pad  ;
  assign n466 = n123 & n465 ;
  assign n467 = ~n464 & ~n466 ;
  assign n468 = n28 & ~n467 ;
  assign n469 = ~\v2_pad  & \v9_reg/NET0131  ;
  assign n470 = \v8_reg/NET0131  & n469 ;
  assign n471 = ~n333 & ~n470 ;
  assign n472 = \v11_reg/NET0131  & ~n454 ;
  assign n473 = ~n471 & n472 ;
  assign n474 = n32 & n407 ;
  assign n475 = ~n473 & ~n474 ;
  assign n476 = n320 & ~n475 ;
  assign n477 = n28 & n466 ;
  assign n478 = n138 & n227 ;
  assign n479 = \v6_pad  & n101 ;
  assign n480 = n176 & n479 ;
  assign n481 = ~n478 & ~n480 ;
  assign n482 = ~\v7_reg/NET0131  & n148 ;
  assign n483 = ~n481 & n482 ;
  assign n484 = ~n477 & ~n483 ;
  assign n485 = n17 & n32 ;
  assign n486 = \v2_pad  & n176 ;
  assign n487 = ~n485 & ~n486 ;
  assign n488 = ~\v7_reg/NET0131  & n118 ;
  assign n489 = ~n487 & n488 ;
  assign n490 = \v7_reg/NET0131  & n176 ;
  assign n491 = n102 & n490 ;
  assign n492 = n45 & n61 ;
  assign n493 = \v12_reg/NET0131  & n235 ;
  assign n494 = ~n492 & ~n493 ;
  assign n495 = ~\v10_reg/NET0131  & ~\v7_reg/NET0131  ;
  assign n496 = ~n494 & n495 ;
  assign n497 = ~n491 & ~n496 ;
  assign n498 = n370 & n380 ;
  assign n499 = \v0_pad  & n122 ;
  assign n500 = ~n498 & ~n499 ;
  assign n501 = ~\v9_reg/NET0131  & ~n500 ;
  assign n502 = n19 & n64 ;
  assign n503 = ~n501 & ~n502 ;
  assign n504 = n203 & ~n503 ;
  assign n505 = ~\v5_pad  & n45 ;
  assign n506 = ~n19 & ~n505 ;
  assign n507 = ~\v10_reg/NET0131  & ~n506 ;
  assign n508 = ~n179 & ~n507 ;
  assign n509 = n136 & ~n508 ;
  assign n510 = n148 & n480 ;
  assign n511 = ~n509 & ~n510 ;
  assign n512 = ~\v7_reg/NET0131  & ~n511 ;
  assign n514 = ~\v10_reg/NET0131  & n176 ;
  assign n513 = \v10_reg/NET0131  & ~n176 ;
  assign n515 = n200 & ~n513 ;
  assign n516 = ~n514 & n515 ;
  assign n517 = ~\v5_pad  & n76 ;
  assign n518 = ~n123 & ~n517 ;
  assign n519 = n61 & ~n68 ;
  assign n520 = ~n518 & n519 ;
  assign n521 = ~n516 & ~n520 ;
  assign n522 = \v11_reg/NET0131  & ~n521 ;
  assign n523 = n61 & n68 ;
  assign n524 = ~\v5_pad  & n36 ;
  assign n525 = n203 & n524 ;
  assign n526 = ~n523 & ~n525 ;
  assign n527 = ~\v0_pad  & n16 ;
  assign n528 = ~n526 & n527 ;
  assign n529 = ~n522 & ~n528 ;
  assign n530 = ~n512 & n529 ;
  assign n531 = ~n41 & ~n258 ;
  assign n532 = n69 & ~n531 ;
  assign n533 = ~n133 & n427 ;
  assign n534 = ~n532 & ~n533 ;
  assign n535 = \v7_reg/NET0131  & ~n534 ;
  assign n536 = n181 & n359 ;
  assign n537 = ~n19 & ~n101 ;
  assign n538 = ~\v8_reg/NET0131  & ~n36 ;
  assign n539 = ~n537 & n538 ;
  assign n540 = ~n536 & ~n539 ;
  assign n541 = ~\v9_reg/NET0131  & ~n540 ;
  assign n542 = ~n318 & ~n333 ;
  assign n543 = ~\v12_reg/NET0131  & ~n298 ;
  assign n544 = ~n542 & n543 ;
  assign n545 = ~n541 & ~n544 ;
  assign n546 = ~\v7_reg/NET0131  & ~n545 ;
  assign n547 = ~n535 & ~n546 ;
  assign n550 = ~\v0_pad  & ~\v12_reg/NET0131  ;
  assign n551 = \v11_reg/NET0131  & ~n550 ;
  assign n552 = ~\v9_reg/NET0131  & ~n102 ;
  assign n553 = ~n551 & n552 ;
  assign n554 = ~\v8_reg/NET0131  & ~n553 ;
  assign n556 = ~\v2_pad  & n101 ;
  assign n557 = ~\v11_reg/NET0131  & ~n335 ;
  assign n558 = ~n556 & n557 ;
  assign n548 = ~n71 & ~n469 ;
  assign n549 = ~n298 & ~n548 ;
  assign n555 = ~n45 & n47 ;
  assign n559 = ~\v7_reg/NET0131  & ~n233 ;
  assign n560 = ~n555 & n559 ;
  assign n561 = ~n549 & n560 ;
  assign n562 = ~n558 & n561 ;
  assign n563 = ~n554 & n562 ;
  assign n564 = \v9_reg/NET0131  & ~n45 ;
  assign n565 = ~n19 & n28 ;
  assign n566 = ~n564 & n565 ;
  assign n567 = n434 & ~n566 ;
  assign n568 = ~n563 & ~n567 ;
  assign n569 = ~n16 & n133 ;
  assign n570 = ~n269 & n569 ;
  assign n571 = ~n568 & ~n570 ;
  assign n572 = ~n37 & ~n193 ;
  assign n573 = \v9_reg/NET0131  & ~n572 ;
  assign n574 = ~\v9_reg/NET0131  & n61 ;
  assign n575 = \v0_pad  & n71 ;
  assign n576 = ~n574 & ~n575 ;
  assign n577 = \v10_reg/NET0131  & ~\v7_reg/NET0131  ;
  assign n578 = ~n576 & n577 ;
  assign n579 = ~n573 & ~n578 ;
  assign n580 = ~\v12_reg/NET0131  & ~n579 ;
  assign \_al_n0  = 1'b0 ;
  assign \_al_n1  = ~1'b0 ;
  assign \g1759/_1_  = n87 ;
  assign \g1762/_1_  = n147 ;
  assign \g1764/_1_  = n210 ;
  assign \g1765/_0_  = n256 ;
  assign \g1786/_2_  = ~n281 ;
  assign \g1791/_3_  = ~n297 ;
  assign \g1808/_3_  = ~n316 ;
  assign \g1822/_2_  = n323 ;
  assign \g1929/_3_  = n326 ;
  assign \g2713/_1_  = n358 ;
  assign \g2744/_0_  = n395 ;
  assign \v13_D_11_pad  = ~n406 ;
  assign \v13_D_12_pad  = ~n422 ;
  assign \v13_D_13_pad  = ~n449 ;
  assign \v13_D_14_pad  = ~n463 ;
  assign \v13_D_16_pad  = n468 ;
  assign \v13_D_18_pad  = n476 ;
  assign \v13_D_19_pad  = ~n484 ;
  assign \v13_D_21_pad  = n489 ;
  assign \v13_D_22_pad  = ~n497 ;
  assign \v13_D_23_pad  = n504 ;
  assign \v13_D_24_pad  = ~n530 ;
  assign \v13_D_7_pad  = ~n547 ;
  assign \v13_D_8_pad  = ~n571 ;
  assign \v13_D_9_pad  = n580 ;
endmodule
