module top (\1(0)_pad , \100(77)_pad , \101(78)_pad , \102(79)_pad , \103(80)_pad , \104(81)_pad , \105(82)_pad , \106(83)_pad , \107(84)_pad , \108(85)_pad , \11(8)_pad , \111(86)_pad , \112(87)_pad , \113(88)_pad , \114(89)_pad , \115(90)_pad , \116(91)_pad , \117(92)_pad , \118(93)_pad , \119(94)_pad , \120(95)_pad , \123(96)_pad , \124(97)_pad , \125(98)_pad , \126(99)_pad , \127(100)_pad , \128(101)_pad , \129(102)_pad , \130(103)_pad , \131(104)_pad , \132(105)_pad , \1341(200)_pad , \1348(201)_pad , \135(106)_pad , \136(107)_pad , \137(108)_pad , \138(109)_pad , \1384(202)_pad , \139(110)_pad , \14(9)_pad , \140(111)_pad , \141(112)_pad , \142(113)_pad , \15(10)_pad , \16(11)_pad , \19(12)_pad , \1956(203)_pad , \1961(204)_pad , \1966(205)_pad , \1971(206)_pad , \1976(207)_pad , \1981(208)_pad , \1986(209)_pad , \1991(210)_pad , \1996(211)_pad , \2(1)_pad , \20(13)_pad , \2067(213)_pad , \2072(214)_pad , \2078(215)_pad , \2084(216)_pad , \2090(217)_pad , \2096(218)_pad , \21(14)_pad , \2100(219)_pad , \2104(220)_pad , \2105(221)_pad , \2106(222)_pad , \22(15)_pad , \23(16)_pad , \24(17)_pad , \2427(223)_pad , \2430(224)_pad , \2435(225)_pad , \2438(226)_pad , \2443(227)_pad , \2446(228)_pad , \2451(229)_pad , \2454(230)_pad , \2474(231)_pad , \25(18)_pad , \26(19)_pad , \2678(232)_pad , \27(20)_pad , \28(21)_pad , \29(22)_pad , \3(2)_pad , \32(23)_pad , \33(24)_pad , \34(25)_pad , \35(26)_pad , \36(27)_pad , \37(28)_pad , \4(3)_pad , \40(29)_pad , \409(298)_pad , \43(30)_pad , \44(31)_pad , \47(32)_pad , \48(33)_pad , \483(191)_pad , \49(34)_pad , \5(4)_pad , \50(35)_pad , \51(36)_pad , \52(37)_pad , \53(38)_pad , \54(39)_pad , \543(192)_pad , \55(40)_pad , \559(193)_pad , \56(41)_pad , \567(194)_pad , \57(42)_pad , \6(5)_pad , \60(43)_pad , \61(44)_pad , \62(45)_pad , \63(46)_pad , \64(47)_pad , \65(48)_pad , \651(195)_pad , \66(49)_pad , \661(196)_pad , \67(50)_pad , \68(51)_pad , \69(52)_pad , \7(6)_pad , \72(53)_pad , \73(54)_pad , \74(55)_pad , \75(56)_pad , \76(57)_pad , \77(58)_pad , \78(59)_pad , \79(60)_pad , \8(7)_pad , \80(61)_pad , \81(62)_pad , \82(63)_pad , \85(64)_pad , \86(65)_pad , \860(197)_pad , \868(198)_pad , \87(66)_pad , \88(67)_pad , \89(68)_pad , \90(69)_pad , \91(70)_pad , \92(71)_pad , \93(72)_pad , \94(73)_pad , \95(74)_pad , \96(75)_pad , \99(76)_pad , \145(1358)_pad , \148(851)_pad , \150(1277)_pad , \153(671)_pad , \156(1046)_pad , \158(349)_pad , \160(609)_pad , \162(612)_pad , \164(607)_pad , \166(625)_pad , \168(623)_pad , \171(621)_pad , \173(389)_pad , \176(803)_pad , \188(761)_pad , \217(423)_pad , \218(311)_pad , \219(302)_pad , \220(306)_pad , \221(305)_pad , \223(413)_pad , \225(1424)_pad , \227(1179)_pad , \229(1180)_pad , \234(376)_pad , \235(307)_pad , \236(303)_pad , \237(309)_pad , \238(304)_pad , \259(414)_pad , \261(506)_pad , \282(922)_pad , \284(847)_pad , \286(696)_pad , \288(700)_pad , \290(704)_pad , \295(1400)_pad , \297(849)_pad , \299(692)_pad , \301(694)_pad , \303(698)_pad , \305(702)_pad , \325(507)_pad , \329(1414)_pad , \_al_n0 , \u1082_syn_3 , \u1396_syn_3 , \u1414_syn_3 , \u1447_syn_3 , \u538_syn_3 , \u539_syn_3 );
	input \1(0)_pad  ;
	input \100(77)_pad  ;
	input \101(78)_pad  ;
	input \102(79)_pad  ;
	input \103(80)_pad  ;
	input \104(81)_pad  ;
	input \105(82)_pad  ;
	input \106(83)_pad  ;
	input \107(84)_pad  ;
	input \108(85)_pad  ;
	input \11(8)_pad  ;
	input \111(86)_pad  ;
	input \112(87)_pad  ;
	input \113(88)_pad  ;
	input \114(89)_pad  ;
	input \115(90)_pad  ;
	input \116(91)_pad  ;
	input \117(92)_pad  ;
	input \118(93)_pad  ;
	input \119(94)_pad  ;
	input \120(95)_pad  ;
	input \123(96)_pad  ;
	input \124(97)_pad  ;
	input \125(98)_pad  ;
	input \126(99)_pad  ;
	input \127(100)_pad  ;
	input \128(101)_pad  ;
	input \129(102)_pad  ;
	input \130(103)_pad  ;
	input \131(104)_pad  ;
	input \132(105)_pad  ;
	input \1341(200)_pad  ;
	input \1348(201)_pad  ;
	input \135(106)_pad  ;
	input \136(107)_pad  ;
	input \137(108)_pad  ;
	input \138(109)_pad  ;
	input \1384(202)_pad  ;
	input \139(110)_pad  ;
	input \14(9)_pad  ;
	input \140(111)_pad  ;
	input \141(112)_pad  ;
	input \142(113)_pad  ;
	input \15(10)_pad  ;
	input \16(11)_pad  ;
	input \19(12)_pad  ;
	input \1956(203)_pad  ;
	input \1961(204)_pad  ;
	input \1966(205)_pad  ;
	input \1971(206)_pad  ;
	input \1976(207)_pad  ;
	input \1981(208)_pad  ;
	input \1986(209)_pad  ;
	input \1991(210)_pad  ;
	input \1996(211)_pad  ;
	input \2(1)_pad  ;
	input \20(13)_pad  ;
	input \2067(213)_pad  ;
	input \2072(214)_pad  ;
	input \2078(215)_pad  ;
	input \2084(216)_pad  ;
	input \2090(217)_pad  ;
	input \2096(218)_pad  ;
	input \21(14)_pad  ;
	input \2100(219)_pad  ;
	input \2104(220)_pad  ;
	input \2105(221)_pad  ;
	input \2106(222)_pad  ;
	input \22(15)_pad  ;
	input \23(16)_pad  ;
	input \24(17)_pad  ;
	input \2427(223)_pad  ;
	input \2430(224)_pad  ;
	input \2435(225)_pad  ;
	input \2438(226)_pad  ;
	input \2443(227)_pad  ;
	input \2446(228)_pad  ;
	input \2451(229)_pad  ;
	input \2454(230)_pad  ;
	input \2474(231)_pad  ;
	input \25(18)_pad  ;
	input \26(19)_pad  ;
	input \2678(232)_pad  ;
	input \27(20)_pad  ;
	input \28(21)_pad  ;
	input \29(22)_pad  ;
	input \3(2)_pad  ;
	input \32(23)_pad  ;
	input \33(24)_pad  ;
	input \34(25)_pad  ;
	input \35(26)_pad  ;
	input \36(27)_pad  ;
	input \37(28)_pad  ;
	input \4(3)_pad  ;
	input \40(29)_pad  ;
	input \409(298)_pad  ;
	input \43(30)_pad  ;
	input \44(31)_pad  ;
	input \47(32)_pad  ;
	input \48(33)_pad  ;
	input \483(191)_pad  ;
	input \49(34)_pad  ;
	input \5(4)_pad  ;
	input \50(35)_pad  ;
	input \51(36)_pad  ;
	input \52(37)_pad  ;
	input \53(38)_pad  ;
	input \54(39)_pad  ;
	input \543(192)_pad  ;
	input \55(40)_pad  ;
	input \559(193)_pad  ;
	input \56(41)_pad  ;
	input \567(194)_pad  ;
	input \57(42)_pad  ;
	input \6(5)_pad  ;
	input \60(43)_pad  ;
	input \61(44)_pad  ;
	input \62(45)_pad  ;
	input \63(46)_pad  ;
	input \64(47)_pad  ;
	input \65(48)_pad  ;
	input \651(195)_pad  ;
	input \66(49)_pad  ;
	input \661(196)_pad  ;
	input \67(50)_pad  ;
	input \68(51)_pad  ;
	input \69(52)_pad  ;
	input \7(6)_pad  ;
	input \72(53)_pad  ;
	input \73(54)_pad  ;
	input \74(55)_pad  ;
	input \75(56)_pad  ;
	input \76(57)_pad  ;
	input \77(58)_pad  ;
	input \78(59)_pad  ;
	input \79(60)_pad  ;
	input \8(7)_pad  ;
	input \80(61)_pad  ;
	input \81(62)_pad  ;
	input \82(63)_pad  ;
	input \85(64)_pad  ;
	input \86(65)_pad  ;
	input \860(197)_pad  ;
	input \868(198)_pad  ;
	input \87(66)_pad  ;
	input \88(67)_pad  ;
	input \89(68)_pad  ;
	input \90(69)_pad  ;
	input \91(70)_pad  ;
	input \92(71)_pad  ;
	input \93(72)_pad  ;
	input \94(73)_pad  ;
	input \95(74)_pad  ;
	input \96(75)_pad  ;
	input \99(76)_pad  ;
	output \145(1358)_pad  ;
	output \148(851)_pad  ;
	output \150(1277)_pad  ;
	output \153(671)_pad  ;
	output \156(1046)_pad  ;
	output \158(349)_pad  ;
	output \160(609)_pad  ;
	output \162(612)_pad  ;
	output \164(607)_pad  ;
	output \166(625)_pad  ;
	output \168(623)_pad  ;
	output \171(621)_pad  ;
	output \173(389)_pad  ;
	output \176(803)_pad  ;
	output \188(761)_pad  ;
	output \217(423)_pad  ;
	output \218(311)_pad  ;
	output \219(302)_pad  ;
	output \220(306)_pad  ;
	output \221(305)_pad  ;
	output \223(413)_pad  ;
	output \225(1424)_pad  ;
	output \227(1179)_pad  ;
	output \229(1180)_pad  ;
	output \234(376)_pad  ;
	output \235(307)_pad  ;
	output \236(303)_pad  ;
	output \237(309)_pad  ;
	output \238(304)_pad  ;
	output \259(414)_pad  ;
	output \261(506)_pad  ;
	output \282(922)_pad  ;
	output \284(847)_pad  ;
	output \286(696)_pad  ;
	output \288(700)_pad  ;
	output \290(704)_pad  ;
	output \295(1400)_pad  ;
	output \297(849)_pad  ;
	output \299(692)_pad  ;
	output \301(694)_pad  ;
	output \303(698)_pad  ;
	output \305(702)_pad  ;
	output \325(507)_pad  ;
	output \329(1414)_pad  ;
	output \_al_n0  ;
	output \u1082_syn_3  ;
	output \u1396_syn_3  ;
	output \u1414_syn_3  ;
	output \u1447_syn_3  ;
	output \u538_syn_3  ;
	output \u539_syn_3  ;
	wire _w380_ ;
	wire _w379_ ;
	wire _w378_ ;
	wire _w376_ ;
	wire _w375_ ;
	wire _w374_ ;
	wire _w373_ ;
	wire _w372_ ;
	wire _w371_ ;
	wire _w370_ ;
	wire _w369_ ;
	wire _w368_ ;
	wire _w367_ ;
	wire _w366_ ;
	wire _w365_ ;
	wire _w364_ ;
	wire _w363_ ;
	wire _w362_ ;
	wire _w361_ ;
	wire _w359_ ;
	wire _w358_ ;
	wire _w357_ ;
	wire _w356_ ;
	wire _w355_ ;
	wire _w354_ ;
	wire _w353_ ;
	wire _w352_ ;
	wire _w351_ ;
	wire _w350_ ;
	wire _w349_ ;
	wire _w348_ ;
	wire _w347_ ;
	wire _w346_ ;
	wire _w345_ ;
	wire _w344_ ;
	wire _w343_ ;
	wire _w342_ ;
	wire _w341_ ;
	wire _w340_ ;
	wire _w339_ ;
	wire _w338_ ;
	wire _w337_ ;
	wire _w336_ ;
	wire _w335_ ;
	wire _w334_ ;
	wire _w333_ ;
	wire _w332_ ;
	wire _w331_ ;
	wire _w330_ ;
	wire _w329_ ;
	wire _w328_ ;
	wire _w327_ ;
	wire _w326_ ;
	wire _w325_ ;
	wire _w324_ ;
	wire _w323_ ;
	wire _w322_ ;
	wire _w321_ ;
	wire _w320_ ;
	wire _w319_ ;
	wire _w318_ ;
	wire _w317_ ;
	wire _w316_ ;
	wire _w315_ ;
	wire _w314_ ;
	wire _w313_ ;
	wire _w312_ ;
	wire _w311_ ;
	wire _w310_ ;
	wire _w309_ ;
	wire _w308_ ;
	wire _w307_ ;
	wire _w306_ ;
	wire _w305_ ;
	wire _w304_ ;
	wire _w303_ ;
	wire _w302_ ;
	wire _w301_ ;
	wire _w300_ ;
	wire _w299_ ;
	wire _w298_ ;
	wire _w297_ ;
	wire _w296_ ;
	wire _w295_ ;
	wire _w294_ ;
	wire _w293_ ;
	wire _w291_ ;
	wire _w290_ ;
	wire _w289_ ;
	wire _w288_ ;
	wire _w287_ ;
	wire _w286_ ;
	wire _w285_ ;
	wire _w284_ ;
	wire _w215_ ;
	wire _w214_ ;
	wire _w213_ ;
	wire _w211_ ;
	wire _w210_ ;
	wire _w209_ ;
	wire _w208_ ;
	wire _w206_ ;
	wire _w205_ ;
	wire _w204_ ;
	wire _w203_ ;
	wire _w202_ ;
	wire _w200_ ;
	wire _w199_ ;
	wire _w198_ ;
	wire _w197_ ;
	wire _w196_ ;
	wire _w195_ ;
	wire _w194_ ;
	wire _w192_ ;
	wire _w191_ ;
	wire _w190_ ;
	wire _w188_ ;
	wire _w187_ ;
	wire _w186_ ;
	wire _w169_ ;
	wire _w201_ ;
	wire _w278_ ;
	wire _w166_ ;
	wire _w163_ ;
	wire _w193_ ;
	wire _w134_ ;
	wire _w261_ ;
	wire _w207_ ;
	wire _w148_ ;
	wire _w275_ ;
	wire _w177_ ;
	wire _w178_ ;
	wire _w165_ ;
	wire _w212_ ;
	wire _w292_ ;
	wire _w35_ ;
	wire _w180_ ;
	wire _w167_ ;
	wire _w168_ ;
	wire _w360_ ;
	wire _w103_ ;
	wire _w230_ ;
	wire _w189_ ;
	wire _w266_ ;
	wire _w170_ ;
	wire _w171_ ;
	wire _w172_ ;
	wire _w173_ ;
	wire _w174_ ;
	wire _w175_ ;
	wire _w176_ ;
	wire _w377_ ;
	wire _w120_ ;
	wire _w247_ ;
	wire _w179_ ;
	wire _w181_ ;
	wire _w182_ ;
	wire _w183_ ;
	wire _w184_ ;
	wire _w185_ ;
	wire _w216_ ;
	wire _w217_ ;
	wire _w218_ ;
	wire _w219_ ;
	wire _w220_ ;
	wire _w221_ ;
	wire _w222_ ;
	wire _w223_ ;
	wire _w224_ ;
	wire _w225_ ;
	wire _w226_ ;
	wire _w227_ ;
	wire _w228_ ;
	wire _w229_ ;
	wire _w231_ ;
	wire _w232_ ;
	wire _w233_ ;
	wire _w234_ ;
	wire _w235_ ;
	wire _w236_ ;
	wire _w237_ ;
	wire _w238_ ;
	wire _w239_ ;
	wire _w240_ ;
	wire _w241_ ;
	wire _w242_ ;
	wire _w243_ ;
	wire _w244_ ;
	wire _w245_ ;
	wire _w246_ ;
	wire _w248_ ;
	wire _w249_ ;
	wire _w250_ ;
	wire _w251_ ;
	wire _w252_ ;
	wire _w253_ ;
	wire _w254_ ;
	wire _w255_ ;
	wire _w256_ ;
	wire _w257_ ;
	wire _w258_ ;
	wire _w259_ ;
	wire _w260_ ;
	wire _w262_ ;
	wire _w263_ ;
	wire _w264_ ;
	wire _w265_ ;
	wire _w267_ ;
	wire _w268_ ;
	wire _w12_ ;
	wire _w269_ ;
	wire _w270_ ;
	wire _w271_ ;
	wire _w272_ ;
	wire _w273_ ;
	wire _w274_ ;
	wire _w276_ ;
	wire _w277_ ;
	wire _w279_ ;
	wire _w280_ ;
	wire _w24_ ;
	wire _w281_ ;
	wire _w282_ ;
	wire _w283_ ;
	LUT1 #(
		.INIT('h1)
	) name0 (
		\108(85)_pad ,
		_w12_
	);
	LUT1 #(
		.INIT('h1)
	) name1 (
		\120(95)_pad ,
		_w24_
	);
	LUT1 #(
		.INIT('h1)
	) name2 (
		\132(105)_pad ,
		_w35_
	);
	LUT1 #(
		.INIT('h1)
	) name3 (
		\44(31)_pad ,
		_w103_
	);
	LUT1 #(
		.INIT('h1)
	) name4 (
		\57(42)_pad ,
		_w120_
	);
	LUT1 #(
		.INIT('h1)
	) name5 (
		\69(52)_pad ,
		_w134_
	);
	LUT1 #(
		.INIT('h1)
	) name6 (
		\82(63)_pad ,
		_w148_
	);
	LUT1 #(
		.INIT('h1)
	) name7 (
		\96(75)_pad ,
		_w163_
	);
	LUT4 #(
		.INIT('h37f7)
	) name8 (
		\54(39)_pad ,
		\543(192)_pad ,
		\651(195)_pad ,
		\79(60)_pad ,
		_w165_
	);
	LUT4 #(
		.INIT('haebf)
	) name9 (
		\543(192)_pad ,
		\651(195)_pad ,
		\66(49)_pad ,
		\92(71)_pad ,
		_w166_
	);
	LUT2 #(
		.INIT('h8)
	) name10 (
		_w165_,
		_w166_,
		_w167_
	);
	LUT3 #(
		.INIT('h80)
	) name11 (
		\559(193)_pad ,
		_w165_,
		_w166_,
		_w168_
	);
	LUT4 #(
		.INIT('h2000)
	) name12 (
		\559(193)_pad ,
		\860(197)_pad ,
		_w165_,
		_w166_,
		_w169_
	);
	LUT4 #(
		.INIT('h37f7)
	) name13 (
		\43(30)_pad ,
		\543(192)_pad ,
		\651(195)_pad ,
		\68(51)_pad ,
		_w170_
	);
	LUT4 #(
		.INIT('hbabf)
	) name14 (
		\543(192)_pad ,
		\56(41)_pad ,
		\651(195)_pad ,
		\81(62)_pad ,
		_w171_
	);
	LUT2 #(
		.INIT('h8)
	) name15 (
		_w170_,
		_w171_,
		_w172_
	);
	LUT3 #(
		.INIT('h80)
	) name16 (
		\860(197)_pad ,
		_w170_,
		_w171_,
		_w173_
	);
	LUT3 #(
		.INIT('h7f)
	) name17 (
		\860(197)_pad ,
		_w170_,
		_w171_,
		_w174_
	);
	LUT4 #(
		.INIT('h57f7)
	) name18 (
		\543(192)_pad ,
		\55(40)_pad ,
		\651(195)_pad ,
		\80(61)_pad ,
		_w175_
	);
	LUT4 #(
		.INIT('haebf)
	) name19 (
		\543(192)_pad ,
		\651(195)_pad ,
		\67(50)_pad ,
		\93(72)_pad ,
		_w176_
	);
	LUT4 #(
		.INIT('h8777)
	) name20 (
		_w170_,
		_w171_,
		_w175_,
		_w176_,
		_w177_
	);
	LUT3 #(
		.INIT('h1e)
	) name21 (
		_w169_,
		_w173_,
		_w177_,
		_w178_
	);
	LUT4 #(
		.INIT('h2fff)
	) name22 (
		\559(193)_pad ,
		\860(197)_pad ,
		_w165_,
		_w166_,
		_w179_
	);
	LUT4 #(
		.INIT('hb111)
	) name23 (
		\16(11)_pad ,
		\19(12)_pad ,
		_w170_,
		_w171_,
		_w180_
	);
	LUT3 #(
		.INIT('hab)
	) name24 (
		\543(192)_pad ,
		\651(195)_pad ,
		\87(66)_pad ,
		_w181_
	);
	LUT4 #(
		.INIT('h37f7)
	) name25 (
		\49(34)_pad ,
		\543(192)_pad ,
		\651(195)_pad ,
		\74(55)_pad ,
		_w182_
	);
	LUT2 #(
		.INIT('h8)
	) name26 (
		_w181_,
		_w182_,
		_w183_
	);
	LUT2 #(
		.INIT('h7)
	) name27 (
		_w181_,
		_w182_,
		_w184_
	);
	LUT4 #(
		.INIT('h4eee)
	) name28 (
		\16(11)_pad ,
		\23(16)_pad ,
		_w181_,
		_w182_,
		_w185_
	);
	LUT4 #(
		.INIT('ha854)
	) name29 (
		\1341(200)_pad ,
		\1976(207)_pad ,
		_w185_,
		_w180_,
		_w186_
	);
	LUT4 #(
		.INIT('h37f7)
	) name30 (
		\50(35)_pad ,
		\543(192)_pad ,
		\651(195)_pad ,
		\75(56)_pad ,
		_w187_
	);
	LUT4 #(
		.INIT('hbabf)
	) name31 (
		\543(192)_pad ,
		\62(45)_pad ,
		\651(195)_pad ,
		\88(67)_pad ,
		_w188_
	);
	LUT2 #(
		.INIT('h8)
	) name32 (
		_w187_,
		_w188_,
		_w189_
	);
	LUT2 #(
		.INIT('h7)
	) name33 (
		_w187_,
		_w188_,
		_w190_
	);
	LUT4 #(
		.INIT('h4eee)
	) name34 (
		\16(11)_pad ,
		\22(15)_pad ,
		_w187_,
		_w188_,
		_w191_
	);
	LUT4 #(
		.INIT('h37f7)
	) name35 (
		\51(36)_pad ,
		\543(192)_pad ,
		\651(195)_pad ,
		\76(57)_pad ,
		_w192_
	);
	LUT4 #(
		.INIT('hbabf)
	) name36 (
		\543(192)_pad ,
		\63(46)_pad ,
		\651(195)_pad ,
		\89(68)_pad ,
		_w193_
	);
	LUT2 #(
		.INIT('h8)
	) name37 (
		_w192_,
		_w193_,
		_w194_
	);
	LUT2 #(
		.INIT('h7)
	) name38 (
		_w192_,
		_w193_,
		_w195_
	);
	LUT4 #(
		.INIT('hb111)
	) name39 (
		\16(11)_pad ,
		\21(14)_pad ,
		_w192_,
		_w193_,
		_w196_
	);
	LUT4 #(
		.INIT('hf5c4)
	) name40 (
		\1966(205)_pad ,
		\1971(206)_pad ,
		_w196_,
		_w191_,
		_w197_
	);
	LUT4 #(
		.INIT('h37f7)
	) name41 (
		\52(37)_pad ,
		\543(192)_pad ,
		\651(195)_pad ,
		\77(58)_pad ,
		_w198_
	);
	LUT4 #(
		.INIT('hbabf)
	) name42 (
		\543(192)_pad ,
		\64(47)_pad ,
		\651(195)_pad ,
		\90(69)_pad ,
		_w199_
	);
	LUT2 #(
		.INIT('h8)
	) name43 (
		_w198_,
		_w199_,
		_w200_
	);
	LUT2 #(
		.INIT('h7)
	) name44 (
		_w198_,
		_w199_,
		_w201_
	);
	LUT4 #(
		.INIT('hb111)
	) name45 (
		\16(11)_pad ,
		\5(4)_pad ,
		_w198_,
		_w199_,
		_w202_
	);
	LUT2 #(
		.INIT('h9)
	) name46 (
		\1961(204)_pad ,
		_w202_,
		_w203_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name47 (
		\105(82)_pad ,
		\117(92)_pad ,
		\2104(220)_pad ,
		\2105(221)_pad ,
		_w204_
	);
	LUT4 #(
		.INIT('hf5f3)
	) name48 (
		\129(102)_pad ,
		\141(112)_pad ,
		\2104(220)_pad ,
		\2105(221)_pad ,
		_w205_
	);
	LUT2 #(
		.INIT('h8)
	) name49 (
		_w204_,
		_w205_,
		_w206_
	);
	LUT4 #(
		.INIT('h4eee)
	) name50 (
		\29(22)_pad ,
		\32(23)_pad ,
		_w204_,
		_w205_,
		_w207_
	);
	LUT4 #(
		.INIT('h153f)
	) name51 (
		\1971(206)_pad ,
		\1996(211)_pad ,
		_w207_,
		_w191_,
		_w208_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name52 (
		\103(80)_pad ,
		\115(90)_pad ,
		\2104(220)_pad ,
		\2105(221)_pad ,
		_w209_
	);
	LUT4 #(
		.INIT('hf5f3)
	) name53 (
		\127(100)_pad ,
		\139(110)_pad ,
		\2104(220)_pad ,
		\2105(221)_pad ,
		_w210_
	);
	LUT2 #(
		.INIT('h8)
	) name54 (
		_w209_,
		_w210_,
		_w211_
	);
	LUT4 #(
		.INIT('h4eee)
	) name55 (
		\29(22)_pad ,
		\33(24)_pad ,
		_w209_,
		_w210_,
		_w212_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name56 (
		\104(81)_pad ,
		\116(91)_pad ,
		\2104(220)_pad ,
		\2105(221)_pad ,
		_w213_
	);
	LUT4 #(
		.INIT('hf5f3)
	) name57 (
		\128(101)_pad ,
		\140(111)_pad ,
		\2104(220)_pad ,
		\2105(221)_pad ,
		_w214_
	);
	LUT4 #(
		.INIT('h2eee)
	) name58 (
		\26(19)_pad ,
		\29(22)_pad ,
		_w213_,
		_w214_,
		_w215_
	);
	LUT4 #(
		.INIT('h3f2a)
	) name59 (
		\2067(213)_pad ,
		\2072(214)_pad ,
		_w212_,
		_w215_,
		_w216_
	);
	LUT4 #(
		.INIT('h8000)
	) name60 (
		_w208_,
		_w216_,
		_w197_,
		_w203_,
		_w217_
	);
	LUT2 #(
		.INIT('h8)
	) name61 (
		_w186_,
		_w217_,
		_w218_
	);
	LUT4 #(
		.INIT('h37f7)
	) name62 (
		\48(33)_pad ,
		\543(192)_pad ,
		\651(195)_pad ,
		\73(54)_pad ,
		_w219_
	);
	LUT4 #(
		.INIT('hbabf)
	) name63 (
		\543(192)_pad ,
		\61(44)_pad ,
		\651(195)_pad ,
		\86(65)_pad ,
		_w220_
	);
	LUT2 #(
		.INIT('h8)
	) name64 (
		_w219_,
		_w220_,
		_w221_
	);
	LUT2 #(
		.INIT('h7)
	) name65 (
		_w219_,
		_w220_,
		_w222_
	);
	LUT4 #(
		.INIT('hb111)
	) name66 (
		\16(11)_pad ,
		\6(5)_pad ,
		_w219_,
		_w220_,
		_w223_
	);
	LUT2 #(
		.INIT('h6)
	) name67 (
		\1981(208)_pad ,
		_w223_,
		_w224_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name68 (
		\100(77)_pad ,
		\112(87)_pad ,
		\2104(220)_pad ,
		\2105(221)_pad ,
		_w225_
	);
	LUT4 #(
		.INIT('hf5f3)
	) name69 (
		\124(97)_pad ,
		\136(107)_pad ,
		\2104(220)_pad ,
		\2105(221)_pad ,
		_w226_
	);
	LUT2 #(
		.INIT('h8)
	) name70 (
		_w225_,
		_w226_,
		_w227_
	);
	LUT4 #(
		.INIT('hb111)
	) name71 (
		\29(22)_pad ,
		\35(26)_pad ,
		_w225_,
		_w226_,
		_w228_
	);
	LUT2 #(
		.INIT('h6)
	) name72 (
		\2090(217)_pad ,
		_w228_,
		_w229_
	);
	LUT4 #(
		.INIT('h737f)
	) name73 (
		\111(86)_pad ,
		\2104(220)_pad ,
		\2105(221)_pad ,
		\99(76)_pad ,
		_w230_
	);
	LUT4 #(
		.INIT('hf5f3)
	) name74 (
		\123(96)_pad ,
		\135(106)_pad ,
		\2104(220)_pad ,
		\2105(221)_pad ,
		_w231_
	);
	LUT3 #(
		.INIT('ha8)
	) name75 (
		\11(8)_pad ,
		\28(21)_pad ,
		\29(22)_pad ,
		_w232_
	);
	LUT4 #(
		.INIT('h7f00)
	) name76 (
		\29(22)_pad ,
		_w230_,
		_w231_,
		_w232_,
		_w233_
	);
	LUT3 #(
		.INIT('he0)
	) name77 (
		\2072(214)_pad ,
		_w212_,
		_w233_,
		_w234_
	);
	LUT3 #(
		.INIT('h10)
	) name78 (
		_w229_,
		_w224_,
		_w234_,
		_w235_
	);
	LUT4 #(
		.INIT('hb111)
	) name79 (
		\16(11)_pad ,
		\4(3)_pad ,
		_w165_,
		_w166_,
		_w236_
	);
	LUT4 #(
		.INIT('h37f7)
	) name80 (
		\47(32)_pad ,
		\543(192)_pad ,
		\651(195)_pad ,
		\72(53)_pad ,
		_w237_
	);
	LUT4 #(
		.INIT('hbabf)
	) name81 (
		\543(192)_pad ,
		\60(43)_pad ,
		\651(195)_pad ,
		\85(64)_pad ,
		_w238_
	);
	LUT2 #(
		.INIT('h8)
	) name82 (
		_w237_,
		_w238_,
		_w239_
	);
	LUT2 #(
		.INIT('h7)
	) name83 (
		_w237_,
		_w238_,
		_w240_
	);
	LUT4 #(
		.INIT('hb111)
	) name84 (
		\16(11)_pad ,
		\24(17)_pad ,
		_w237_,
		_w238_,
		_w241_
	);
	LUT4 #(
		.INIT('haf23)
	) name85 (
		\1348(201)_pad ,
		\1986(209)_pad ,
		_w236_,
		_w241_,
		_w242_
	);
	LUT4 #(
		.INIT('h737f)
	) name86 (
		\107(84)_pad ,
		\2104(220)_pad ,
		\2105(221)_pad ,
		\95(74)_pad ,
		_w243_
	);
	LUT4 #(
		.INIT('hf5f3)
	) name87 (
		\119(94)_pad ,
		\131(104)_pad ,
		\2104(220)_pad ,
		\2105(221)_pad ,
		_w244_
	);
	LUT2 #(
		.INIT('h8)
	) name88 (
		_w243_,
		_w244_,
		_w245_
	);
	LUT4 #(
		.INIT('hd111)
	) name89 (
		\25(18)_pad ,
		\29(22)_pad ,
		_w243_,
		_w244_,
		_w246_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name90 (
		\101(78)_pad ,
		\113(88)_pad ,
		\2104(220)_pad ,
		\2105(221)_pad ,
		_w247_
	);
	LUT4 #(
		.INIT('hf5f3)
	) name91 (
		\125(98)_pad ,
		\137(108)_pad ,
		\2104(220)_pad ,
		\2105(221)_pad ,
		_w248_
	);
	LUT2 #(
		.INIT('h8)
	) name92 (
		_w247_,
		_w248_,
		_w249_
	);
	LUT4 #(
		.INIT('h4eee)
	) name93 (
		\29(22)_pad ,
		\34(25)_pad ,
		_w247_,
		_w248_,
		_w250_
	);
	LUT4 #(
		.INIT('h31f5)
	) name94 (
		\1991(210)_pad ,
		\2084(216)_pad ,
		_w246_,
		_w250_,
		_w251_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name95 (
		\102(79)_pad ,
		\114(89)_pad ,
		\2104(220)_pad ,
		\2105(221)_pad ,
		_w252_
	);
	LUT4 #(
		.INIT('hf5f3)
	) name96 (
		\126(99)_pad ,
		\138(109)_pad ,
		\2104(220)_pad ,
		\2105(221)_pad ,
		_w253_
	);
	LUT2 #(
		.INIT('h8)
	) name97 (
		_w252_,
		_w253_,
		_w254_
	);
	LUT4 #(
		.INIT('hd111)
	) name98 (
		\27(20)_pad ,
		\29(22)_pad ,
		_w252_,
		_w253_,
		_w255_
	);
	LUT4 #(
		.INIT('h8acf)
	) name99 (
		\1966(205)_pad ,
		\2078(215)_pad ,
		_w255_,
		_w196_,
		_w256_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name100 (
		\1348(201)_pad ,
		\1986(209)_pad ,
		_w236_,
		_w241_,
		_w257_
	);
	LUT4 #(
		.INIT('h8000)
	) name101 (
		_w256_,
		_w257_,
		_w242_,
		_w251_,
		_w258_
	);
	LUT4 #(
		.INIT('haf8c)
	) name102 (
		\1991(210)_pad ,
		\1996(211)_pad ,
		_w246_,
		_w207_,
		_w259_
	);
	LUT4 #(
		.INIT('h51f3)
	) name103 (
		\1976(207)_pad ,
		\2078(215)_pad ,
		_w255_,
		_w185_,
		_w260_
	);
	LUT4 #(
		.INIT('h37f7)
	) name104 (
		\53(38)_pad ,
		\543(192)_pad ,
		\651(195)_pad ,
		\78(59)_pad ,
		_w261_
	);
	LUT4 #(
		.INIT('hbabf)
	) name105 (
		\543(192)_pad ,
		\65(48)_pad ,
		\651(195)_pad ,
		\91(70)_pad ,
		_w262_
	);
	LUT2 #(
		.INIT('h8)
	) name106 (
		_w261_,
		_w262_,
		_w263_
	);
	LUT2 #(
		.INIT('h7)
	) name107 (
		_w261_,
		_w262_,
		_w264_
	);
	LUT4 #(
		.INIT('hb111)
	) name108 (
		\16(11)_pad ,
		\20(13)_pad ,
		_w261_,
		_w262_,
		_w265_
	);
	LUT2 #(
		.INIT('h9)
	) name109 (
		\1956(203)_pad ,
		_w265_,
		_w266_
	);
	LUT4 #(
		.INIT('h54fc)
	) name110 (
		\2067(213)_pad ,
		\2084(216)_pad ,
		_w250_,
		_w215_,
		_w267_
	);
	LUT4 #(
		.INIT('h8000)
	) name111 (
		_w266_,
		_w267_,
		_w259_,
		_w260_,
		_w268_
	);
	LUT3 #(
		.INIT('h80)
	) name112 (
		_w235_,
		_w258_,
		_w268_,
		_w269_
	);
	LUT2 #(
		.INIT('h8)
	) name113 (
		_w218_,
		_w269_,
		_w270_
	);
	LUT2 #(
		.INIT('h7)
	) name114 (
		_w218_,
		_w269_,
		_w271_
	);
	LUT4 #(
		.INIT('hdeee)
	) name115 (
		\2096(218)_pad ,
		\2100(219)_pad ,
		_w230_,
		_w231_,
		_w272_
	);
	LUT4 #(
		.INIT('h7fff)
	) name116 (
		\2072(214)_pad ,
		\2078(215)_pad ,
		\2084(216)_pad ,
		\2090(217)_pad ,
		_w273_
	);
	LUT2 #(
		.INIT('h8)
	) name117 (
		\409(298)_pad ,
		\94(73)_pad ,
		_w274_
	);
	LUT4 #(
		.INIT('h8000)
	) name118 (
		\108(85)_pad ,
		\120(95)_pad ,
		\57(42)_pad ,
		\69(52)_pad ,
		_w275_
	);
	LUT4 #(
		.INIT('h8000)
	) name119 (
		\132(105)_pad ,
		\44(31)_pad ,
		\82(63)_pad ,
		\96(75)_pad ,
		_w276_
	);
	LUT4 #(
		.INIT('hf351)
	) name120 (
		\2106(222)_pad ,
		\567(194)_pad ,
		_w275_,
		_w276_,
		_w277_
	);
	LUT3 #(
		.INIT('h80)
	) name121 (
		\36(27)_pad ,
		\483(191)_pad ,
		\661(196)_pad ,
		_w278_
	);
	LUT2 #(
		.INIT('h7)
	) name122 (
		_w277_,
		_w278_,
		_w279_
	);
	LUT4 #(
		.INIT('h7000)
	) name123 (
		\1(0)_pad ,
		\3(2)_pad ,
		\483(191)_pad ,
		\661(196)_pad ,
		_w280_
	);
	LUT2 #(
		.INIT('h7)
	) name124 (
		_w277_,
		_w280_,
		_w281_
	);
	LUT2 #(
		.INIT('h7)
	) name125 (
		\661(196)_pad ,
		\7(6)_pad ,
		_w282_
	);
	LUT3 #(
		.INIT('h7f)
	) name126 (
		\2106(222)_pad ,
		\661(196)_pad ,
		\7(6)_pad ,
		_w283_
	);
	LUT4 #(
		.INIT('h8777)
	) name127 (
		_w261_,
		_w262_,
		_w187_,
		_w188_,
		_w284_
	);
	LUT4 #(
		.INIT('h6996)
	) name128 (
		_w177_,
		_w221_,
		_w239_,
		_w183_,
		_w285_
	);
	LUT4 #(
		.INIT('h8777)
	) name129 (
		_w165_,
		_w166_,
		_w198_,
		_w199_,
		_w286_
	);
	LUT2 #(
		.INIT('h6)
	) name130 (
		_w194_,
		_w286_,
		_w287_
	);
	LUT4 #(
		.INIT('h4114)
	) name131 (
		\37(28)_pad ,
		_w284_,
		_w285_,
		_w287_,
		_w288_
	);
	LUT4 #(
		.INIT('h8777)
	) name132 (
		_w225_,
		_w226_,
		_w230_,
		_w231_,
		_w289_
	);
	LUT2 #(
		.INIT('h6)
	) name133 (
		_w249_,
		_w289_,
		_w290_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name134 (
		\106(83)_pad ,
		\118(93)_pad ,
		\2104(220)_pad ,
		\2105(221)_pad ,
		_w291_
	);
	LUT4 #(
		.INIT('hf5f3)
	) name135 (
		\130(103)_pad ,
		\142(113)_pad ,
		\2104(220)_pad ,
		\2105(221)_pad ,
		_w292_
	);
	LUT4 #(
		.INIT('h8777)
	) name136 (
		_w252_,
		_w253_,
		_w291_,
		_w292_,
		_w293_
	);
	LUT4 #(
		.INIT('h8777)
	) name137 (
		_w213_,
		_w214_,
		_w204_,
		_w205_,
		_w294_
	);
	LUT4 #(
		.INIT('h9669)
	) name138 (
		_w211_,
		_w245_,
		_w293_,
		_w294_,
		_w295_
	);
	LUT3 #(
		.INIT('h41)
	) name139 (
		\37(28)_pad ,
		_w290_,
		_w295_,
		_w296_
	);
	LUT4 #(
		.INIT('h6996)
	) name140 (
		\1341(200)_pad ,
		\1348(201)_pad ,
		\2435(225)_pad ,
		\2438(226)_pad ,
		_w297_
	);
	LUT2 #(
		.INIT('h6)
	) name141 (
		\2446(228)_pad ,
		\2454(230)_pad ,
		_w298_
	);
	LUT4 #(
		.INIT('h6996)
	) name142 (
		\2427(223)_pad ,
		\2430(224)_pad ,
		\2443(227)_pad ,
		\2451(229)_pad ,
		_w299_
	);
	LUT4 #(
		.INIT('h2882)
	) name143 (
		\14(9)_pad ,
		_w297_,
		_w298_,
		_w299_,
		_w300_
	);
	LUT4 #(
		.INIT('h6996)
	) name144 (
		\1971(206)_pad ,
		\1976(207)_pad ,
		\1981(208)_pad ,
		\2474(231)_pad ,
		_w301_
	);
	LUT4 #(
		.INIT('h9669)
	) name145 (
		\1961(204)_pad ,
		\1966(205)_pad ,
		\1986(209)_pad ,
		\1991(210)_pad ,
		_w302_
	);
	LUT2 #(
		.INIT('h9)
	) name146 (
		\1956(203)_pad ,
		\1996(211)_pad ,
		_w303_
	);
	LUT3 #(
		.INIT('h69)
	) name147 (
		_w301_,
		_w302_,
		_w303_,
		_w304_
	);
	LUT4 #(
		.INIT('h6996)
	) name148 (
		\2072(214)_pad ,
		\2078(215)_pad ,
		\2084(216)_pad ,
		\2096(218)_pad ,
		_w305_
	);
	LUT4 #(
		.INIT('h9669)
	) name149 (
		\2067(213)_pad ,
		\2090(217)_pad ,
		\2100(219)_pad ,
		\2678(232)_pad ,
		_w306_
	);
	LUT2 #(
		.INIT('h6)
	) name150 (
		_w305_,
		_w306_,
		_w307_
	);
	LUT4 #(
		.INIT('h0002)
	) name151 (
		_w277_,
		_w300_,
		_w307_,
		_w304_,
		_w308_
	);
	LUT4 #(
		.INIT('hbe00)
	) name152 (
		\37(28)_pad ,
		_w290_,
		_w295_,
		_w308_,
		_w309_
	);
	LUT2 #(
		.INIT('h4)
	) name153 (
		_w288_,
		_w309_,
		_w310_
	);
	LUT2 #(
		.INIT('hb)
	) name154 (
		_w288_,
		_w309_,
		_w311_
	);
	LUT3 #(
		.INIT('h7f)
	) name155 (
		\567(194)_pad ,
		\661(196)_pad ,
		\7(6)_pad ,
		_w312_
	);
	LUT3 #(
		.INIT('h7f)
	) name156 (
		\15(10)_pad ,
		\2(1)_pad ,
		\661(196)_pad ,
		_w313_
	);
	LUT2 #(
		.INIT('h8)
	) name157 (
		_w275_,
		_w276_,
		_w314_
	);
	LUT2 #(
		.INIT('h7)
	) name158 (
		_w275_,
		_w276_,
		_w315_
	);
	LUT3 #(
		.INIT('h40)
	) name159 (
		\868(198)_pad ,
		_w170_,
		_w171_,
		_w316_
	);
	LUT2 #(
		.INIT('h4)
	) name160 (
		\559(193)_pad ,
		\868(198)_pad ,
		_w317_
	);
	LUT3 #(
		.INIT('h80)
	) name161 (
		_w165_,
		_w166_,
		_w317_,
		_w318_
	);
	LUT2 #(
		.INIT('h1)
	) name162 (
		_w316_,
		_w318_,
		_w319_
	);
	LUT3 #(
		.INIT('h2a)
	) name163 (
		\868(198)_pad ,
		_w198_,
		_w199_,
		_w320_
	);
	LUT3 #(
		.INIT('h15)
	) name164 (
		\868(198)_pad ,
		_w165_,
		_w166_,
		_w321_
	);
	LUT2 #(
		.INIT('he)
	) name165 (
		_w320_,
		_w321_,
		_w322_
	);
	LUT4 #(
		.INIT('h2882)
	) name166 (
		\868(198)_pad ,
		_w168_,
		_w284_,
		_w285_,
		_w323_
	);
	LUT3 #(
		.INIT('h15)
	) name167 (
		\868(198)_pad ,
		_w175_,
		_w176_,
		_w324_
	);
	LUT2 #(
		.INIT('he)
	) name168 (
		_w323_,
		_w324_,
		_w325_
	);
	LUT3 #(
		.INIT('h2a)
	) name169 (
		\868(198)_pad ,
		_w192_,
		_w193_,
		_w326_
	);
	LUT3 #(
		.INIT('h15)
	) name170 (
		\868(198)_pad ,
		_w261_,
		_w262_,
		_w327_
	);
	LUT2 #(
		.INIT('he)
	) name171 (
		_w326_,
		_w327_,
		_w328_
	);
	LUT3 #(
		.INIT('h15)
	) name172 (
		\1384(202)_pad ,
		_w252_,
		_w253_,
		_w329_
	);
	LUT3 #(
		.INIT('h80)
	) name173 (
		\40(29)_pad ,
		_w247_,
		_w248_,
		_w330_
	);
	LUT4 #(
		.INIT('h3555)
	) name174 (
		\1348(201)_pad ,
		\2067(213)_pad ,
		_w329_,
		_w330_,
		_w331_
	);
	LUT3 #(
		.INIT('h2a)
	) name175 (
		\1341(200)_pad ,
		_w329_,
		_w330_,
		_w332_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name176 (
		\1996(211)_pad ,
		_w172_,
		_w329_,
		_w330_,
		_w333_
	);
	LUT4 #(
		.INIT('h0e00)
	) name177 (
		_w167_,
		_w331_,
		_w332_,
		_w333_,
		_w334_
	);
	LUT4 #(
		.INIT('h3555)
	) name178 (
		\1956(203)_pad ,
		\2072(214)_pad ,
		_w329_,
		_w330_,
		_w335_
	);
	LUT4 #(
		.INIT('h153f)
	) name179 (
		_w167_,
		_w263_,
		_w335_,
		_w331_,
		_w336_
	);
	LUT4 #(
		.INIT('h3555)
	) name180 (
		\1961(204)_pad ,
		\2078(215)_pad ,
		_w329_,
		_w330_,
		_w337_
	);
	LUT2 #(
		.INIT('h8)
	) name181 (
		_w200_,
		_w337_,
		_w338_
	);
	LUT4 #(
		.INIT('h32c8)
	) name182 (
		_w263_,
		_w200_,
		_w335_,
		_w337_,
		_w339_
	);
	LUT3 #(
		.INIT('h2a)
	) name183 (
		\1966(205)_pad ,
		_w329_,
		_w330_,
		_w340_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name184 (
		\2084(216)_pad ,
		\8(7)_pad ,
		_w329_,
		_w330_,
		_w341_
	);
	LUT3 #(
		.INIT('h2a)
	) name185 (
		\8(7)_pad ,
		_w192_,
		_w193_,
		_w342_
	);
	LUT3 #(
		.INIT('hb0)
	) name186 (
		_w340_,
		_w341_,
		_w342_,
		_w343_
	);
	LUT3 #(
		.INIT('h20)
	) name187 (
		_w194_,
		_w340_,
		_w341_,
		_w344_
	);
	LUT4 #(
		.INIT('hd3dd)
	) name188 (
		\8(7)_pad ,
		_w194_,
		_w340_,
		_w341_,
		_w345_
	);
	LUT4 #(
		.INIT('hb000)
	) name189 (
		_w334_,
		_w336_,
		_w339_,
		_w345_,
		_w346_
	);
	LUT3 #(
		.INIT('h0b)
	) name190 (
		_w343_,
		_w338_,
		_w344_,
		_w347_
	);
	LUT3 #(
		.INIT('h2a)
	) name191 (
		\1971(206)_pad ,
		_w329_,
		_w330_,
		_w348_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name192 (
		\2090(217)_pad ,
		\8(7)_pad ,
		_w329_,
		_w330_,
		_w349_
	);
	LUT3 #(
		.INIT('h2a)
	) name193 (
		\8(7)_pad ,
		_w187_,
		_w188_,
		_w350_
	);
	LUT3 #(
		.INIT('hb0)
	) name194 (
		_w348_,
		_w349_,
		_w350_,
		_w351_
	);
	LUT3 #(
		.INIT('h20)
	) name195 (
		_w189_,
		_w348_,
		_w349_,
		_w352_
	);
	LUT3 #(
		.INIT('h40)
	) name196 (
		\1976(207)_pad ,
		_w181_,
		_w182_,
		_w353_
	);
	LUT4 #(
		.INIT('h2a00)
	) name197 (
		\8(7)_pad ,
		_w329_,
		_w330_,
		_w353_,
		_w354_
	);
	LUT3 #(
		.INIT('h2a)
	) name198 (
		\1981(208)_pad ,
		_w219_,
		_w220_,
		_w355_
	);
	LUT4 #(
		.INIT('h2a00)
	) name199 (
		\8(7)_pad ,
		_w329_,
		_w330_,
		_w355_,
		_w356_
	);
	LUT3 #(
		.INIT('h2a)
	) name200 (
		\1976(207)_pad ,
		_w181_,
		_w182_,
		_w357_
	);
	LUT4 #(
		.INIT('h2a00)
	) name201 (
		\8(7)_pad ,
		_w329_,
		_w330_,
		_w357_,
		_w358_
	);
	LUT3 #(
		.INIT('h40)
	) name202 (
		\1981(208)_pad ,
		_w219_,
		_w220_,
		_w359_
	);
	LUT4 #(
		.INIT('h2a00)
	) name203 (
		\8(7)_pad ,
		_w329_,
		_w330_,
		_w359_,
		_w360_
	);
	LUT4 #(
		.INIT('h0001)
	) name204 (
		_w354_,
		_w356_,
		_w358_,
		_w360_,
		_w361_
	);
	LUT3 #(
		.INIT('h10)
	) name205 (
		_w352_,
		_w351_,
		_w361_,
		_w362_
	);
	LUT4 #(
		.INIT('h0200)
	) name206 (
		_w189_,
		_w358_,
		_w348_,
		_w349_,
		_w363_
	);
	LUT4 #(
		.INIT('h0c0d)
	) name207 (
		_w354_,
		_w356_,
		_w360_,
		_w363_,
		_w364_
	);
	LUT4 #(
		.INIT('h4f00)
	) name208 (
		_w346_,
		_w347_,
		_w362_,
		_w364_,
		_w365_
	);
	LUT2 #(
		.INIT('h4)
	) name209 (
		_w329_,
		_w330_,
		_w366_
	);
	LUT3 #(
		.INIT('h40)
	) name210 (
		\2067(213)_pad ,
		_w213_,
		_w214_,
		_w367_
	);
	LUT3 #(
		.INIT('h2a)
	) name211 (
		\1991(210)_pad ,
		_w243_,
		_w244_,
		_w368_
	);
	LUT3 #(
		.INIT('h40)
	) name212 (
		\1986(209)_pad ,
		_w237_,
		_w238_,
		_w369_
	);
	LUT4 #(
		.INIT('h0009)
	) name213 (
		\1986(209)_pad ,
		_w239_,
		_w367_,
		_w368_,
		_w370_
	);
	LUT3 #(
		.INIT('h2a)
	) name214 (
		\2067(213)_pad ,
		_w213_,
		_w214_,
		_w371_
	);
	LUT3 #(
		.INIT('h2a)
	) name215 (
		\1996(211)_pad ,
		_w204_,
		_w205_,
		_w372_
	);
	LUT2 #(
		.INIT('h1)
	) name216 (
		_w371_,
		_w372_,
		_w373_
	);
	LUT3 #(
		.INIT('h40)
	) name217 (
		\1991(210)_pad ,
		_w243_,
		_w244_,
		_w374_
	);
	LUT3 #(
		.INIT('h40)
	) name218 (
		\1996(211)_pad ,
		_w204_,
		_w205_,
		_w375_
	);
	LUT4 #(
		.INIT('h0009)
	) name219 (
		\1996(211)_pad ,
		_w206_,
		_w371_,
		_w374_,
		_w376_
	);
	LUT3 #(
		.INIT('h2a)
	) name220 (
		_w366_,
		_w370_,
		_w376_,
		_w377_
	);
	LUT4 #(
		.INIT('h002b)
	) name221 (
		\1991(210)_pad ,
		_w245_,
		_w369_,
		_w375_,
		_w378_
	);
	LUT4 #(
		.INIT('h88a8)
	) name222 (
		_w366_,
		_w367_,
		_w373_,
		_w378_,
		_w379_
	);
	LUT3 #(
		.INIT('hf1)
	) name223 (
		_w365_,
		_w377_,
		_w379_,
		_w380_
	);
	assign \145(1358)_pad  = _w178_ ;
	assign \148(851)_pad  = _w179_ ;
	assign \150(1277)_pad  = _w271_ ;
	assign \153(671)_pad  = _w174_ ;
	assign \156(1046)_pad  = _w272_ ;
	assign \158(349)_pad  = _w273_ ;
	assign \160(609)_pad  = _w249_ ;
	assign \162(612)_pad  = _w227_ ;
	assign \164(607)_pad  = _w254_ ;
	assign \166(625)_pad  = _w189_ ;
	assign \168(623)_pad  = _w194_ ;
	assign \171(621)_pad  = _w200_ ;
	assign \173(389)_pad  = _w274_ ;
	assign \176(803)_pad  = _w279_ ;
	assign \188(761)_pad  = _w281_ ;
	assign \217(423)_pad  = _w283_ ;
	assign \218(311)_pad  = _w103_ ;
	assign \219(302)_pad  = _w35_ ;
	assign \220(306)_pad  = _w148_ ;
	assign \221(305)_pad  = _w163_ ;
	assign \223(413)_pad  = _w282_ ;
	assign \225(1424)_pad  = _w311_ ;
	assign \227(1179)_pad  = _w307_ ;
	assign \229(1180)_pad  = _w304_ ;
	assign \234(376)_pad  = _w312_ ;
	assign \235(307)_pad  = _w134_ ;
	assign \236(303)_pad  = _w24_ ;
	assign \237(309)_pad  = _w120_ ;
	assign \238(304)_pad  = _w12_ ;
	assign \259(414)_pad  = _w313_ ;
	assign \261(506)_pad  = _w315_ ;
	assign \282(922)_pad  = _w319_ ;
	assign \284(847)_pad  = _w322_ ;
	assign \286(696)_pad  = _w195_ ;
	assign \288(700)_pad  = _w184_ ;
	assign \290(704)_pad  = _w240_ ;
	assign \295(1400)_pad  = _w325_ ;
	assign \297(849)_pad  = _w328_ ;
	assign \299(692)_pad  = _w264_ ;
	assign \301(694)_pad  = _w201_ ;
	assign \303(698)_pad  = _w190_ ;
	assign \305(702)_pad  = _w222_ ;
	assign \325(507)_pad  = _w314_ ;
	assign \329(1414)_pad  = _w380_ ;
	assign \_al_n0  = 1'b0;
	assign \u1082_syn_3  = _w277_ ;
	assign \u1396_syn_3  = _w310_ ;
	assign \u1414_syn_3  = _w288_ ;
	assign \u1447_syn_3  = _w296_ ;
	assign \u538_syn_3  = _w270_ ;
	assign \u539_syn_3  = _w300_ ;
endmodule;