module top (\count[0] , \count[1] , \count[2] , \count[3] , \count[4] , \count[5] , \count[6] , \count[7] , \selectp1[0] , \selectp1[1] , \selectp1[2] , \selectp1[3] , \selectp1[4] , \selectp1[5] , \selectp1[6] , \selectp1[7] , \selectp1[8] , \selectp1[9] , \selectp1[10] , \selectp1[11] , \selectp1[12] , \selectp1[13] , \selectp1[14] , \selectp1[15] , \selectp1[16] , \selectp1[17] , \selectp1[18] , \selectp1[19] , \selectp1[20] , \selectp1[21] , \selectp1[22] , \selectp1[23] , \selectp1[24] , \selectp1[25] , \selectp1[26] , \selectp1[27] , \selectp1[28] , \selectp1[29] , \selectp1[30] , \selectp1[31] , \selectp1[32] , \selectp1[33] , \selectp1[34] , \selectp1[35] , \selectp1[36] , \selectp1[37] , \selectp1[38] , \selectp1[39] , \selectp1[40] , \selectp1[41] , \selectp1[42] , \selectp1[43] , \selectp1[44] , \selectp1[45] , \selectp1[46] , \selectp1[47] , \selectp1[48] , \selectp1[49] , \selectp1[50] , \selectp1[51] , \selectp1[52] , \selectp1[53] , \selectp1[54] , \selectp1[55] , \selectp1[56] , \selectp1[57] , \selectp1[58] , \selectp1[59] , \selectp1[60] , \selectp1[61] , \selectp1[62] , \selectp1[63] , \selectp1[64] , \selectp1[65] , \selectp1[66] , \selectp1[67] , \selectp1[68] , \selectp1[69] , \selectp1[70] , \selectp1[71] , \selectp1[72] , \selectp1[73] , \selectp1[74] , \selectp1[75] , \selectp1[76] , \selectp1[77] , \selectp1[78] , \selectp1[79] , \selectp1[80] , \selectp1[81] , \selectp1[82] , \selectp1[83] , \selectp1[84] , \selectp1[85] , \selectp1[86] , \selectp1[87] , \selectp1[88] , \selectp1[89] , \selectp1[90] , \selectp1[91] , \selectp1[92] , \selectp1[93] , \selectp1[94] , \selectp1[95] , \selectp1[96] , \selectp1[97] , \selectp1[98] , \selectp1[99] , \selectp1[100] , \selectp1[101] , \selectp1[102] , \selectp1[103] , \selectp1[104] , \selectp1[105] , \selectp1[106] , \selectp1[107] , \selectp1[108] , \selectp1[109] , \selectp1[110] , \selectp1[111] , \selectp1[112] , \selectp1[113] , \selectp1[114] , \selectp1[115] , \selectp1[116] , \selectp1[117] , \selectp1[118] , \selectp1[119] , \selectp1[120] , \selectp1[121] , \selectp1[122] , \selectp1[123] , \selectp1[124] , \selectp1[125] , \selectp1[126] , \selectp1[127] , \selectp2[0] , \selectp2[1] , \selectp2[2] , \selectp2[3] , \selectp2[4] , \selectp2[5] , \selectp2[6] , \selectp2[7] , \selectp2[8] , \selectp2[9] , \selectp2[10] , \selectp2[11] , \selectp2[12] , \selectp2[13] , \selectp2[14] , \selectp2[15] , \selectp2[16] , \selectp2[17] , \selectp2[18] , \selectp2[19] , \selectp2[20] , \selectp2[21] , \selectp2[22] , \selectp2[23] , \selectp2[24] , \selectp2[25] , \selectp2[26] , \selectp2[27] , \selectp2[28] , \selectp2[29] , \selectp2[30] , \selectp2[31] , \selectp2[32] , \selectp2[33] , \selectp2[34] , \selectp2[35] , \selectp2[36] , \selectp2[37] , \selectp2[38] , \selectp2[39] , \selectp2[40] , \selectp2[41] , \selectp2[42] , \selectp2[43] , \selectp2[44] , \selectp2[45] , \selectp2[46] , \selectp2[47] , \selectp2[48] , \selectp2[49] , \selectp2[50] , \selectp2[51] , \selectp2[52] , \selectp2[53] , \selectp2[54] , \selectp2[55] , \selectp2[56] , \selectp2[57] , \selectp2[58] , \selectp2[59] , \selectp2[60] , \selectp2[61] , \selectp2[62] , \selectp2[63] , \selectp2[64] , \selectp2[65] , \selectp2[66] , \selectp2[67] , \selectp2[68] , \selectp2[69] , \selectp2[70] , \selectp2[71] , \selectp2[72] , \selectp2[73] , \selectp2[74] , \selectp2[75] , \selectp2[76] , \selectp2[77] , \selectp2[78] , \selectp2[79] , \selectp2[80] , \selectp2[81] , \selectp2[82] , \selectp2[83] , \selectp2[84] , \selectp2[85] , \selectp2[86] , \selectp2[87] , \selectp2[88] , \selectp2[89] , \selectp2[90] , \selectp2[91] , \selectp2[92] , \selectp2[93] , \selectp2[94] , \selectp2[95] , \selectp2[96] , \selectp2[97] , \selectp2[98] , \selectp2[99] , \selectp2[100] , \selectp2[101] , \selectp2[102] , \selectp2[103] , \selectp2[104] , \selectp2[105] , \selectp2[106] , \selectp2[107] , \selectp2[108] , \selectp2[109] , \selectp2[110] , \selectp2[111] , \selectp2[112] , \selectp2[113] , \selectp2[114] , \selectp2[115] , \selectp2[116] , \selectp2[117] , \selectp2[118] , \selectp2[119] , \selectp2[120] , \selectp2[121] , \selectp2[122] , \selectp2[123] , \selectp2[124] , \selectp2[125] , \selectp2[126] , \selectp2[127] );
	input \count[0]  ;
	input \count[1]  ;
	input \count[2]  ;
	input \count[3]  ;
	input \count[4]  ;
	input \count[5]  ;
	input \count[6]  ;
	input \count[7]  ;
	output \selectp1[0]  ;
	output \selectp1[1]  ;
	output \selectp1[2]  ;
	output \selectp1[3]  ;
	output \selectp1[4]  ;
	output \selectp1[5]  ;
	output \selectp1[6]  ;
	output \selectp1[7]  ;
	output \selectp1[8]  ;
	output \selectp1[9]  ;
	output \selectp1[10]  ;
	output \selectp1[11]  ;
	output \selectp1[12]  ;
	output \selectp1[13]  ;
	output \selectp1[14]  ;
	output \selectp1[15]  ;
	output \selectp1[16]  ;
	output \selectp1[17]  ;
	output \selectp1[18]  ;
	output \selectp1[19]  ;
	output \selectp1[20]  ;
	output \selectp1[21]  ;
	output \selectp1[22]  ;
	output \selectp1[23]  ;
	output \selectp1[24]  ;
	output \selectp1[25]  ;
	output \selectp1[26]  ;
	output \selectp1[27]  ;
	output \selectp1[28]  ;
	output \selectp1[29]  ;
	output \selectp1[30]  ;
	output \selectp1[31]  ;
	output \selectp1[32]  ;
	output \selectp1[33]  ;
	output \selectp1[34]  ;
	output \selectp1[35]  ;
	output \selectp1[36]  ;
	output \selectp1[37]  ;
	output \selectp1[38]  ;
	output \selectp1[39]  ;
	output \selectp1[40]  ;
	output \selectp1[41]  ;
	output \selectp1[42]  ;
	output \selectp1[43]  ;
	output \selectp1[44]  ;
	output \selectp1[45]  ;
	output \selectp1[46]  ;
	output \selectp1[47]  ;
	output \selectp1[48]  ;
	output \selectp1[49]  ;
	output \selectp1[50]  ;
	output \selectp1[51]  ;
	output \selectp1[52]  ;
	output \selectp1[53]  ;
	output \selectp1[54]  ;
	output \selectp1[55]  ;
	output \selectp1[56]  ;
	output \selectp1[57]  ;
	output \selectp1[58]  ;
	output \selectp1[59]  ;
	output \selectp1[60]  ;
	output \selectp1[61]  ;
	output \selectp1[62]  ;
	output \selectp1[63]  ;
	output \selectp1[64]  ;
	output \selectp1[65]  ;
	output \selectp1[66]  ;
	output \selectp1[67]  ;
	output \selectp1[68]  ;
	output \selectp1[69]  ;
	output \selectp1[70]  ;
	output \selectp1[71]  ;
	output \selectp1[72]  ;
	output \selectp1[73]  ;
	output \selectp1[74]  ;
	output \selectp1[75]  ;
	output \selectp1[76]  ;
	output \selectp1[77]  ;
	output \selectp1[78]  ;
	output \selectp1[79]  ;
	output \selectp1[80]  ;
	output \selectp1[81]  ;
	output \selectp1[82]  ;
	output \selectp1[83]  ;
	output \selectp1[84]  ;
	output \selectp1[85]  ;
	output \selectp1[86]  ;
	output \selectp1[87]  ;
	output \selectp1[88]  ;
	output \selectp1[89]  ;
	output \selectp1[90]  ;
	output \selectp1[91]  ;
	output \selectp1[92]  ;
	output \selectp1[93]  ;
	output \selectp1[94]  ;
	output \selectp1[95]  ;
	output \selectp1[96]  ;
	output \selectp1[97]  ;
	output \selectp1[98]  ;
	output \selectp1[99]  ;
	output \selectp1[100]  ;
	output \selectp1[101]  ;
	output \selectp1[102]  ;
	output \selectp1[103]  ;
	output \selectp1[104]  ;
	output \selectp1[105]  ;
	output \selectp1[106]  ;
	output \selectp1[107]  ;
	output \selectp1[108]  ;
	output \selectp1[109]  ;
	output \selectp1[110]  ;
	output \selectp1[111]  ;
	output \selectp1[112]  ;
	output \selectp1[113]  ;
	output \selectp1[114]  ;
	output \selectp1[115]  ;
	output \selectp1[116]  ;
	output \selectp1[117]  ;
	output \selectp1[118]  ;
	output \selectp1[119]  ;
	output \selectp1[120]  ;
	output \selectp1[121]  ;
	output \selectp1[122]  ;
	output \selectp1[123]  ;
	output \selectp1[124]  ;
	output \selectp1[125]  ;
	output \selectp1[126]  ;
	output \selectp1[127]  ;
	output \selectp2[0]  ;
	output \selectp2[1]  ;
	output \selectp2[2]  ;
	output \selectp2[3]  ;
	output \selectp2[4]  ;
	output \selectp2[5]  ;
	output \selectp2[6]  ;
	output \selectp2[7]  ;
	output \selectp2[8]  ;
	output \selectp2[9]  ;
	output \selectp2[10]  ;
	output \selectp2[11]  ;
	output \selectp2[12]  ;
	output \selectp2[13]  ;
	output \selectp2[14]  ;
	output \selectp2[15]  ;
	output \selectp2[16]  ;
	output \selectp2[17]  ;
	output \selectp2[18]  ;
	output \selectp2[19]  ;
	output \selectp2[20]  ;
	output \selectp2[21]  ;
	output \selectp2[22]  ;
	output \selectp2[23]  ;
	output \selectp2[24]  ;
	output \selectp2[25]  ;
	output \selectp2[26]  ;
	output \selectp2[27]  ;
	output \selectp2[28]  ;
	output \selectp2[29]  ;
	output \selectp2[30]  ;
	output \selectp2[31]  ;
	output \selectp2[32]  ;
	output \selectp2[33]  ;
	output \selectp2[34]  ;
	output \selectp2[35]  ;
	output \selectp2[36]  ;
	output \selectp2[37]  ;
	output \selectp2[38]  ;
	output \selectp2[39]  ;
	output \selectp2[40]  ;
	output \selectp2[41]  ;
	output \selectp2[42]  ;
	output \selectp2[43]  ;
	output \selectp2[44]  ;
	output \selectp2[45]  ;
	output \selectp2[46]  ;
	output \selectp2[47]  ;
	output \selectp2[48]  ;
	output \selectp2[49]  ;
	output \selectp2[50]  ;
	output \selectp2[51]  ;
	output \selectp2[52]  ;
	output \selectp2[53]  ;
	output \selectp2[54]  ;
	output \selectp2[55]  ;
	output \selectp2[56]  ;
	output \selectp2[57]  ;
	output \selectp2[58]  ;
	output \selectp2[59]  ;
	output \selectp2[60]  ;
	output \selectp2[61]  ;
	output \selectp2[62]  ;
	output \selectp2[63]  ;
	output \selectp2[64]  ;
	output \selectp2[65]  ;
	output \selectp2[66]  ;
	output \selectp2[67]  ;
	output \selectp2[68]  ;
	output \selectp2[69]  ;
	output \selectp2[70]  ;
	output \selectp2[71]  ;
	output \selectp2[72]  ;
	output \selectp2[73]  ;
	output \selectp2[74]  ;
	output \selectp2[75]  ;
	output \selectp2[76]  ;
	output \selectp2[77]  ;
	output \selectp2[78]  ;
	output \selectp2[79]  ;
	output \selectp2[80]  ;
	output \selectp2[81]  ;
	output \selectp2[82]  ;
	output \selectp2[83]  ;
	output \selectp2[84]  ;
	output \selectp2[85]  ;
	output \selectp2[86]  ;
	output \selectp2[87]  ;
	output \selectp2[88]  ;
	output \selectp2[89]  ;
	output \selectp2[90]  ;
	output \selectp2[91]  ;
	output \selectp2[92]  ;
	output \selectp2[93]  ;
	output \selectp2[94]  ;
	output \selectp2[95]  ;
	output \selectp2[96]  ;
	output \selectp2[97]  ;
	output \selectp2[98]  ;
	output \selectp2[99]  ;
	output \selectp2[100]  ;
	output \selectp2[101]  ;
	output \selectp2[102]  ;
	output \selectp2[103]  ;
	output \selectp2[104]  ;
	output \selectp2[105]  ;
	output \selectp2[106]  ;
	output \selectp2[107]  ;
	output \selectp2[108]  ;
	output \selectp2[109]  ;
	output \selectp2[110]  ;
	output \selectp2[111]  ;
	output \selectp2[112]  ;
	output \selectp2[113]  ;
	output \selectp2[114]  ;
	output \selectp2[115]  ;
	output \selectp2[116]  ;
	output \selectp2[117]  ;
	output \selectp2[118]  ;
	output \selectp2[119]  ;
	output \selectp2[120]  ;
	output \selectp2[121]  ;
	output \selectp2[122]  ;
	output \selectp2[123]  ;
	output \selectp2[124]  ;
	output \selectp2[125]  ;
	output \selectp2[126]  ;
	output \selectp2[127]  ;
	wire _w312_ ;
	wire _w311_ ;
	wire _w310_ ;
	wire _w309_ ;
	wire _w308_ ;
	wire _w307_ ;
	wire _w306_ ;
	wire _w305_ ;
	wire _w304_ ;
	wire _w303_ ;
	wire _w302_ ;
	wire _w301_ ;
	wire _w300_ ;
	wire _w299_ ;
	wire _w298_ ;
	wire _w297_ ;
	wire _w296_ ;
	wire _w295_ ;
	wire _w294_ ;
	wire _w293_ ;
	wire _w292_ ;
	wire _w291_ ;
	wire _w290_ ;
	wire _w289_ ;
	wire _w288_ ;
	wire _w287_ ;
	wire _w286_ ;
	wire _w285_ ;
	wire _w284_ ;
	wire _w283_ ;
	wire _w282_ ;
	wire _w281_ ;
	wire _w280_ ;
	wire _w279_ ;
	wire _w278_ ;
	wire _w277_ ;
	wire _w276_ ;
	wire _w275_ ;
	wire _w274_ ;
	wire _w273_ ;
	wire _w272_ ;
	wire _w271_ ;
	wire _w270_ ;
	wire _w269_ ;
	wire _w268_ ;
	wire _w267_ ;
	wire _w266_ ;
	wire _w135_ ;
	wire _w134_ ;
	wire _w133_ ;
	wire _w132_ ;
	wire _w131_ ;
	wire _w130_ ;
	wire _w129_ ;
	wire _w128_ ;
	wire _w127_ ;
	wire _w126_ ;
	wire _w125_ ;
	wire _w124_ ;
	wire _w123_ ;
	wire _w122_ ;
	wire _w121_ ;
	wire _w120_ ;
	wire _w119_ ;
	wire _w118_ ;
	wire _w117_ ;
	wire _w116_ ;
	wire _w115_ ;
	wire _w114_ ;
	wire _w113_ ;
	wire _w112_ ;
	wire _w111_ ;
	wire _w110_ ;
	wire _w109_ ;
	wire _w108_ ;
	wire _w107_ ;
	wire _w106_ ;
	wire _w105_ ;
	wire _w104_ ;
	wire _w103_ ;
	wire _w102_ ;
	wire _w101_ ;
	wire _w100_ ;
	wire _w99_ ;
	wire _w98_ ;
	wire _w97_ ;
	wire _w96_ ;
	wire _w95_ ;
	wire _w94_ ;
	wire _w93_ ;
	wire _w92_ ;
	wire _w91_ ;
	wire _w90_ ;
	wire _w89_ ;
	wire _w88_ ;
	wire _w87_ ;
	wire _w86_ ;
	wire _w85_ ;
	wire _w84_ ;
	wire _w83_ ;
	wire _w82_ ;
	wire _w81_ ;
	wire _w80_ ;
	wire _w79_ ;
	wire _w78_ ;
	wire _w77_ ;
	wire _w76_ ;
	wire _w75_ ;
	wire _w74_ ;
	wire _w73_ ;
	wire _w72_ ;
	wire _w71_ ;
	wire _w70_ ;
	wire _w69_ ;
	wire _w68_ ;
	wire _w37_ ;
	wire _w36_ ;
	wire _w35_ ;
	wire _w34_ ;
	wire _w33_ ;
	wire _w32_ ;
	wire _w31_ ;
	wire _w30_ ;
	wire _w29_ ;
	wire _w28_ ;
	wire _w27_ ;
	wire _w26_ ;
	wire _w25_ ;
	wire _w24_ ;
	wire _w23_ ;
	wire _w22_ ;
	wire _w9_ ;
	wire _w10_ ;
	wire _w11_ ;
	wire _w12_ ;
	wire _w13_ ;
	wire _w14_ ;
	wire _w15_ ;
	wire _w16_ ;
	wire _w17_ ;
	wire _w18_ ;
	wire _w19_ ;
	wire _w20_ ;
	wire _w21_ ;
	wire _w38_ ;
	wire _w39_ ;
	wire _w40_ ;
	wire _w41_ ;
	wire _w42_ ;
	wire _w43_ ;
	wire _w44_ ;
	wire _w45_ ;
	wire _w46_ ;
	wire _w47_ ;
	wire _w48_ ;
	wire _w49_ ;
	wire _w50_ ;
	wire _w51_ ;
	wire _w52_ ;
	wire _w53_ ;
	wire _w54_ ;
	wire _w55_ ;
	wire _w56_ ;
	wire _w57_ ;
	wire _w58_ ;
	wire _w59_ ;
	wire _w60_ ;
	wire _w61_ ;
	wire _w62_ ;
	wire _w63_ ;
	wire _w64_ ;
	wire _w65_ ;
	wire _w66_ ;
	wire _w67_ ;
	wire _w136_ ;
	wire _w137_ ;
	wire _w138_ ;
	wire _w139_ ;
	wire _w140_ ;
	wire _w141_ ;
	wire _w142_ ;
	wire _w143_ ;
	wire _w144_ ;
	wire _w145_ ;
	wire _w146_ ;
	wire _w147_ ;
	wire _w148_ ;
	wire _w149_ ;
	wire _w150_ ;
	wire _w151_ ;
	wire _w152_ ;
	wire _w153_ ;
	wire _w154_ ;
	wire _w155_ ;
	wire _w156_ ;
	wire _w157_ ;
	wire _w158_ ;
	wire _w159_ ;
	wire _w160_ ;
	wire _w161_ ;
	wire _w162_ ;
	wire _w163_ ;
	wire _w164_ ;
	wire _w165_ ;
	wire _w166_ ;
	wire _w167_ ;
	wire _w168_ ;
	wire _w169_ ;
	wire _w170_ ;
	wire _w171_ ;
	wire _w172_ ;
	wire _w173_ ;
	wire _w174_ ;
	wire _w175_ ;
	wire _w176_ ;
	wire _w177_ ;
	wire _w178_ ;
	wire _w179_ ;
	wire _w180_ ;
	wire _w181_ ;
	wire _w182_ ;
	wire _w183_ ;
	wire _w184_ ;
	wire _w185_ ;
	wire _w186_ ;
	wire _w187_ ;
	wire _w188_ ;
	wire _w189_ ;
	wire _w190_ ;
	wire _w191_ ;
	wire _w192_ ;
	wire _w193_ ;
	wire _w194_ ;
	wire _w195_ ;
	wire _w196_ ;
	wire _w197_ ;
	wire _w198_ ;
	wire _w199_ ;
	wire _w200_ ;
	wire _w201_ ;
	wire _w202_ ;
	wire _w203_ ;
	wire _w204_ ;
	wire _w205_ ;
	wire _w206_ ;
	wire _w207_ ;
	wire _w208_ ;
	wire _w209_ ;
	wire _w210_ ;
	wire _w211_ ;
	wire _w212_ ;
	wire _w213_ ;
	wire _w214_ ;
	wire _w215_ ;
	wire _w216_ ;
	wire _w217_ ;
	wire _w218_ ;
	wire _w219_ ;
	wire _w220_ ;
	wire _w221_ ;
	wire _w222_ ;
	wire _w223_ ;
	wire _w224_ ;
	wire _w225_ ;
	wire _w226_ ;
	wire _w227_ ;
	wire _w228_ ;
	wire _w229_ ;
	wire _w230_ ;
	wire _w231_ ;
	wire _w232_ ;
	wire _w233_ ;
	wire _w234_ ;
	wire _w235_ ;
	wire _w236_ ;
	wire _w237_ ;
	wire _w238_ ;
	wire _w239_ ;
	wire _w240_ ;
	wire _w241_ ;
	wire _w242_ ;
	wire _w243_ ;
	wire _w244_ ;
	wire _w245_ ;
	wire _w246_ ;
	wire _w247_ ;
	wire _w248_ ;
	wire _w249_ ;
	wire _w250_ ;
	wire _w251_ ;
	wire _w252_ ;
	wire _w253_ ;
	wire _w254_ ;
	wire _w255_ ;
	wire _w256_ ;
	wire _w257_ ;
	wire _w258_ ;
	wire _w259_ ;
	wire _w260_ ;
	wire _w261_ ;
	wire _w262_ ;
	wire _w263_ ;
	wire _w264_ ;
	wire _w265_ ;
	LUT2 #(
		.INIT('h1)
	) name0 (
		\count[4] ,
		\count[5] ,
		_w9_
	);
	LUT2 #(
		.INIT('h4)
	) name1 (
		\count[6] ,
		\count[7] ,
		_w10_
	);
	LUT2 #(
		.INIT('h8)
	) name2 (
		_w9_,
		_w10_,
		_w11_
	);
	LUT2 #(
		.INIT('h1)
	) name3 (
		\count[0] ,
		\count[2] ,
		_w12_
	);
	LUT2 #(
		.INIT('h1)
	) name4 (
		\count[1] ,
		\count[3] ,
		_w13_
	);
	LUT2 #(
		.INIT('h8)
	) name5 (
		_w12_,
		_w13_,
		_w14_
	);
	LUT2 #(
		.INIT('h8)
	) name6 (
		_w11_,
		_w14_,
		_w15_
	);
	LUT2 #(
		.INIT('h2)
	) name7 (
		\count[0] ,
		\count[2] ,
		_w16_
	);
	LUT2 #(
		.INIT('h8)
	) name8 (
		_w13_,
		_w16_,
		_w17_
	);
	LUT2 #(
		.INIT('h8)
	) name9 (
		_w11_,
		_w17_,
		_w18_
	);
	LUT2 #(
		.INIT('h2)
	) name10 (
		\count[1] ,
		\count[3] ,
		_w19_
	);
	LUT2 #(
		.INIT('h8)
	) name11 (
		_w12_,
		_w19_,
		_w20_
	);
	LUT2 #(
		.INIT('h8)
	) name12 (
		_w11_,
		_w20_,
		_w21_
	);
	LUT2 #(
		.INIT('h8)
	) name13 (
		_w16_,
		_w19_,
		_w22_
	);
	LUT2 #(
		.INIT('h8)
	) name14 (
		_w11_,
		_w22_,
		_w23_
	);
	LUT2 #(
		.INIT('h4)
	) name15 (
		\count[0] ,
		\count[2] ,
		_w24_
	);
	LUT2 #(
		.INIT('h8)
	) name16 (
		_w13_,
		_w24_,
		_w25_
	);
	LUT2 #(
		.INIT('h8)
	) name17 (
		_w11_,
		_w25_,
		_w26_
	);
	LUT2 #(
		.INIT('h8)
	) name18 (
		\count[0] ,
		\count[2] ,
		_w27_
	);
	LUT2 #(
		.INIT('h8)
	) name19 (
		_w13_,
		_w27_,
		_w28_
	);
	LUT2 #(
		.INIT('h8)
	) name20 (
		_w11_,
		_w28_,
		_w29_
	);
	LUT2 #(
		.INIT('h8)
	) name21 (
		_w19_,
		_w24_,
		_w30_
	);
	LUT2 #(
		.INIT('h8)
	) name22 (
		_w11_,
		_w30_,
		_w31_
	);
	LUT2 #(
		.INIT('h8)
	) name23 (
		_w19_,
		_w27_,
		_w32_
	);
	LUT2 #(
		.INIT('h8)
	) name24 (
		_w11_,
		_w32_,
		_w33_
	);
	LUT2 #(
		.INIT('h4)
	) name25 (
		\count[1] ,
		\count[3] ,
		_w34_
	);
	LUT2 #(
		.INIT('h8)
	) name26 (
		_w12_,
		_w34_,
		_w35_
	);
	LUT2 #(
		.INIT('h8)
	) name27 (
		_w11_,
		_w35_,
		_w36_
	);
	LUT2 #(
		.INIT('h8)
	) name28 (
		_w16_,
		_w34_,
		_w37_
	);
	LUT2 #(
		.INIT('h8)
	) name29 (
		_w11_,
		_w37_,
		_w38_
	);
	LUT2 #(
		.INIT('h8)
	) name30 (
		\count[1] ,
		\count[3] ,
		_w39_
	);
	LUT2 #(
		.INIT('h8)
	) name31 (
		_w12_,
		_w39_,
		_w40_
	);
	LUT2 #(
		.INIT('h8)
	) name32 (
		_w11_,
		_w40_,
		_w41_
	);
	LUT2 #(
		.INIT('h8)
	) name33 (
		_w16_,
		_w39_,
		_w42_
	);
	LUT2 #(
		.INIT('h8)
	) name34 (
		_w11_,
		_w42_,
		_w43_
	);
	LUT2 #(
		.INIT('h8)
	) name35 (
		_w24_,
		_w34_,
		_w44_
	);
	LUT2 #(
		.INIT('h8)
	) name36 (
		_w11_,
		_w44_,
		_w45_
	);
	LUT2 #(
		.INIT('h8)
	) name37 (
		_w27_,
		_w34_,
		_w46_
	);
	LUT2 #(
		.INIT('h8)
	) name38 (
		_w11_,
		_w46_,
		_w47_
	);
	LUT2 #(
		.INIT('h8)
	) name39 (
		_w24_,
		_w39_,
		_w48_
	);
	LUT2 #(
		.INIT('h8)
	) name40 (
		_w11_,
		_w48_,
		_w49_
	);
	LUT2 #(
		.INIT('h8)
	) name41 (
		_w27_,
		_w39_,
		_w50_
	);
	LUT2 #(
		.INIT('h8)
	) name42 (
		_w11_,
		_w50_,
		_w51_
	);
	LUT2 #(
		.INIT('h2)
	) name43 (
		\count[4] ,
		\count[5] ,
		_w52_
	);
	LUT2 #(
		.INIT('h8)
	) name44 (
		_w10_,
		_w52_,
		_w53_
	);
	LUT2 #(
		.INIT('h8)
	) name45 (
		_w14_,
		_w53_,
		_w54_
	);
	LUT2 #(
		.INIT('h8)
	) name46 (
		_w17_,
		_w53_,
		_w55_
	);
	LUT2 #(
		.INIT('h8)
	) name47 (
		_w20_,
		_w53_,
		_w56_
	);
	LUT2 #(
		.INIT('h8)
	) name48 (
		_w22_,
		_w53_,
		_w57_
	);
	LUT2 #(
		.INIT('h8)
	) name49 (
		_w25_,
		_w53_,
		_w58_
	);
	LUT2 #(
		.INIT('h8)
	) name50 (
		_w28_,
		_w53_,
		_w59_
	);
	LUT2 #(
		.INIT('h8)
	) name51 (
		_w30_,
		_w53_,
		_w60_
	);
	LUT2 #(
		.INIT('h8)
	) name52 (
		_w32_,
		_w53_,
		_w61_
	);
	LUT2 #(
		.INIT('h8)
	) name53 (
		_w35_,
		_w53_,
		_w62_
	);
	LUT2 #(
		.INIT('h8)
	) name54 (
		_w37_,
		_w53_,
		_w63_
	);
	LUT2 #(
		.INIT('h8)
	) name55 (
		_w40_,
		_w53_,
		_w64_
	);
	LUT2 #(
		.INIT('h8)
	) name56 (
		_w42_,
		_w53_,
		_w65_
	);
	LUT2 #(
		.INIT('h8)
	) name57 (
		_w44_,
		_w53_,
		_w66_
	);
	LUT2 #(
		.INIT('h8)
	) name58 (
		_w46_,
		_w53_,
		_w67_
	);
	LUT2 #(
		.INIT('h8)
	) name59 (
		_w48_,
		_w53_,
		_w68_
	);
	LUT2 #(
		.INIT('h8)
	) name60 (
		_w50_,
		_w53_,
		_w69_
	);
	LUT2 #(
		.INIT('h4)
	) name61 (
		\count[4] ,
		\count[5] ,
		_w70_
	);
	LUT2 #(
		.INIT('h8)
	) name62 (
		_w10_,
		_w70_,
		_w71_
	);
	LUT2 #(
		.INIT('h8)
	) name63 (
		_w14_,
		_w71_,
		_w72_
	);
	LUT2 #(
		.INIT('h8)
	) name64 (
		_w17_,
		_w71_,
		_w73_
	);
	LUT2 #(
		.INIT('h8)
	) name65 (
		_w20_,
		_w71_,
		_w74_
	);
	LUT2 #(
		.INIT('h8)
	) name66 (
		_w22_,
		_w71_,
		_w75_
	);
	LUT2 #(
		.INIT('h8)
	) name67 (
		_w25_,
		_w71_,
		_w76_
	);
	LUT2 #(
		.INIT('h8)
	) name68 (
		_w28_,
		_w71_,
		_w77_
	);
	LUT2 #(
		.INIT('h8)
	) name69 (
		_w30_,
		_w71_,
		_w78_
	);
	LUT2 #(
		.INIT('h8)
	) name70 (
		_w32_,
		_w71_,
		_w79_
	);
	LUT2 #(
		.INIT('h8)
	) name71 (
		_w35_,
		_w71_,
		_w80_
	);
	LUT2 #(
		.INIT('h8)
	) name72 (
		_w37_,
		_w71_,
		_w81_
	);
	LUT2 #(
		.INIT('h8)
	) name73 (
		_w40_,
		_w71_,
		_w82_
	);
	LUT2 #(
		.INIT('h8)
	) name74 (
		_w42_,
		_w71_,
		_w83_
	);
	LUT2 #(
		.INIT('h8)
	) name75 (
		_w44_,
		_w71_,
		_w84_
	);
	LUT2 #(
		.INIT('h8)
	) name76 (
		_w46_,
		_w71_,
		_w85_
	);
	LUT2 #(
		.INIT('h8)
	) name77 (
		_w48_,
		_w71_,
		_w86_
	);
	LUT2 #(
		.INIT('h8)
	) name78 (
		_w50_,
		_w71_,
		_w87_
	);
	LUT2 #(
		.INIT('h8)
	) name79 (
		\count[4] ,
		\count[5] ,
		_w88_
	);
	LUT2 #(
		.INIT('h8)
	) name80 (
		_w10_,
		_w88_,
		_w89_
	);
	LUT2 #(
		.INIT('h8)
	) name81 (
		_w14_,
		_w89_,
		_w90_
	);
	LUT2 #(
		.INIT('h8)
	) name82 (
		_w17_,
		_w89_,
		_w91_
	);
	LUT2 #(
		.INIT('h8)
	) name83 (
		_w20_,
		_w89_,
		_w92_
	);
	LUT2 #(
		.INIT('h8)
	) name84 (
		_w22_,
		_w89_,
		_w93_
	);
	LUT2 #(
		.INIT('h8)
	) name85 (
		_w25_,
		_w89_,
		_w94_
	);
	LUT2 #(
		.INIT('h8)
	) name86 (
		_w28_,
		_w89_,
		_w95_
	);
	LUT2 #(
		.INIT('h8)
	) name87 (
		_w30_,
		_w89_,
		_w96_
	);
	LUT2 #(
		.INIT('h8)
	) name88 (
		_w32_,
		_w89_,
		_w97_
	);
	LUT2 #(
		.INIT('h8)
	) name89 (
		_w35_,
		_w89_,
		_w98_
	);
	LUT2 #(
		.INIT('h8)
	) name90 (
		_w37_,
		_w89_,
		_w99_
	);
	LUT2 #(
		.INIT('h8)
	) name91 (
		_w40_,
		_w89_,
		_w100_
	);
	LUT2 #(
		.INIT('h8)
	) name92 (
		_w42_,
		_w89_,
		_w101_
	);
	LUT2 #(
		.INIT('h8)
	) name93 (
		_w44_,
		_w89_,
		_w102_
	);
	LUT2 #(
		.INIT('h8)
	) name94 (
		_w46_,
		_w89_,
		_w103_
	);
	LUT2 #(
		.INIT('h8)
	) name95 (
		_w48_,
		_w89_,
		_w104_
	);
	LUT2 #(
		.INIT('h8)
	) name96 (
		_w50_,
		_w89_,
		_w105_
	);
	LUT2 #(
		.INIT('h8)
	) name97 (
		\count[6] ,
		\count[7] ,
		_w106_
	);
	LUT2 #(
		.INIT('h8)
	) name98 (
		_w9_,
		_w106_,
		_w107_
	);
	LUT2 #(
		.INIT('h8)
	) name99 (
		_w14_,
		_w107_,
		_w108_
	);
	LUT2 #(
		.INIT('h8)
	) name100 (
		_w17_,
		_w107_,
		_w109_
	);
	LUT2 #(
		.INIT('h8)
	) name101 (
		_w20_,
		_w107_,
		_w110_
	);
	LUT2 #(
		.INIT('h8)
	) name102 (
		_w22_,
		_w107_,
		_w111_
	);
	LUT2 #(
		.INIT('h8)
	) name103 (
		_w25_,
		_w107_,
		_w112_
	);
	LUT2 #(
		.INIT('h8)
	) name104 (
		_w28_,
		_w107_,
		_w113_
	);
	LUT2 #(
		.INIT('h8)
	) name105 (
		_w30_,
		_w107_,
		_w114_
	);
	LUT2 #(
		.INIT('h8)
	) name106 (
		_w32_,
		_w107_,
		_w115_
	);
	LUT2 #(
		.INIT('h8)
	) name107 (
		_w35_,
		_w107_,
		_w116_
	);
	LUT2 #(
		.INIT('h8)
	) name108 (
		_w37_,
		_w107_,
		_w117_
	);
	LUT2 #(
		.INIT('h8)
	) name109 (
		_w40_,
		_w107_,
		_w118_
	);
	LUT2 #(
		.INIT('h8)
	) name110 (
		_w42_,
		_w107_,
		_w119_
	);
	LUT2 #(
		.INIT('h8)
	) name111 (
		_w44_,
		_w107_,
		_w120_
	);
	LUT2 #(
		.INIT('h8)
	) name112 (
		_w46_,
		_w107_,
		_w121_
	);
	LUT2 #(
		.INIT('h8)
	) name113 (
		_w48_,
		_w107_,
		_w122_
	);
	LUT2 #(
		.INIT('h8)
	) name114 (
		_w50_,
		_w107_,
		_w123_
	);
	LUT2 #(
		.INIT('h8)
	) name115 (
		_w52_,
		_w106_,
		_w124_
	);
	LUT2 #(
		.INIT('h8)
	) name116 (
		_w14_,
		_w124_,
		_w125_
	);
	LUT2 #(
		.INIT('h8)
	) name117 (
		_w17_,
		_w124_,
		_w126_
	);
	LUT2 #(
		.INIT('h8)
	) name118 (
		_w20_,
		_w124_,
		_w127_
	);
	LUT2 #(
		.INIT('h8)
	) name119 (
		_w22_,
		_w124_,
		_w128_
	);
	LUT2 #(
		.INIT('h8)
	) name120 (
		_w25_,
		_w124_,
		_w129_
	);
	LUT2 #(
		.INIT('h8)
	) name121 (
		_w28_,
		_w124_,
		_w130_
	);
	LUT2 #(
		.INIT('h8)
	) name122 (
		_w30_,
		_w124_,
		_w131_
	);
	LUT2 #(
		.INIT('h8)
	) name123 (
		_w32_,
		_w124_,
		_w132_
	);
	LUT2 #(
		.INIT('h8)
	) name124 (
		_w35_,
		_w124_,
		_w133_
	);
	LUT2 #(
		.INIT('h8)
	) name125 (
		_w37_,
		_w124_,
		_w134_
	);
	LUT2 #(
		.INIT('h8)
	) name126 (
		_w40_,
		_w124_,
		_w135_
	);
	LUT2 #(
		.INIT('h8)
	) name127 (
		_w42_,
		_w124_,
		_w136_
	);
	LUT2 #(
		.INIT('h8)
	) name128 (
		_w44_,
		_w124_,
		_w137_
	);
	LUT2 #(
		.INIT('h8)
	) name129 (
		_w46_,
		_w124_,
		_w138_
	);
	LUT2 #(
		.INIT('h8)
	) name130 (
		_w48_,
		_w124_,
		_w139_
	);
	LUT2 #(
		.INIT('h8)
	) name131 (
		_w50_,
		_w124_,
		_w140_
	);
	LUT2 #(
		.INIT('h8)
	) name132 (
		_w70_,
		_w106_,
		_w141_
	);
	LUT2 #(
		.INIT('h8)
	) name133 (
		_w14_,
		_w141_,
		_w142_
	);
	LUT2 #(
		.INIT('h8)
	) name134 (
		_w17_,
		_w141_,
		_w143_
	);
	LUT2 #(
		.INIT('h8)
	) name135 (
		_w20_,
		_w141_,
		_w144_
	);
	LUT2 #(
		.INIT('h8)
	) name136 (
		_w22_,
		_w141_,
		_w145_
	);
	LUT2 #(
		.INIT('h8)
	) name137 (
		_w25_,
		_w141_,
		_w146_
	);
	LUT2 #(
		.INIT('h8)
	) name138 (
		_w28_,
		_w141_,
		_w147_
	);
	LUT2 #(
		.INIT('h8)
	) name139 (
		_w30_,
		_w141_,
		_w148_
	);
	LUT2 #(
		.INIT('h8)
	) name140 (
		_w32_,
		_w141_,
		_w149_
	);
	LUT2 #(
		.INIT('h8)
	) name141 (
		_w35_,
		_w141_,
		_w150_
	);
	LUT2 #(
		.INIT('h8)
	) name142 (
		_w37_,
		_w141_,
		_w151_
	);
	LUT2 #(
		.INIT('h8)
	) name143 (
		_w40_,
		_w141_,
		_w152_
	);
	LUT2 #(
		.INIT('h8)
	) name144 (
		_w42_,
		_w141_,
		_w153_
	);
	LUT2 #(
		.INIT('h8)
	) name145 (
		_w44_,
		_w141_,
		_w154_
	);
	LUT2 #(
		.INIT('h8)
	) name146 (
		_w46_,
		_w141_,
		_w155_
	);
	LUT2 #(
		.INIT('h8)
	) name147 (
		_w48_,
		_w141_,
		_w156_
	);
	LUT2 #(
		.INIT('h8)
	) name148 (
		_w50_,
		_w141_,
		_w157_
	);
	LUT2 #(
		.INIT('h8)
	) name149 (
		_w88_,
		_w106_,
		_w158_
	);
	LUT2 #(
		.INIT('h8)
	) name150 (
		_w14_,
		_w158_,
		_w159_
	);
	LUT2 #(
		.INIT('h8)
	) name151 (
		_w17_,
		_w158_,
		_w160_
	);
	LUT2 #(
		.INIT('h8)
	) name152 (
		_w20_,
		_w158_,
		_w161_
	);
	LUT2 #(
		.INIT('h8)
	) name153 (
		_w22_,
		_w158_,
		_w162_
	);
	LUT2 #(
		.INIT('h8)
	) name154 (
		_w25_,
		_w158_,
		_w163_
	);
	LUT2 #(
		.INIT('h8)
	) name155 (
		_w28_,
		_w158_,
		_w164_
	);
	LUT2 #(
		.INIT('h8)
	) name156 (
		_w30_,
		_w158_,
		_w165_
	);
	LUT2 #(
		.INIT('h8)
	) name157 (
		_w32_,
		_w158_,
		_w166_
	);
	LUT2 #(
		.INIT('h8)
	) name158 (
		_w35_,
		_w158_,
		_w167_
	);
	LUT2 #(
		.INIT('h8)
	) name159 (
		_w37_,
		_w158_,
		_w168_
	);
	LUT2 #(
		.INIT('h8)
	) name160 (
		_w40_,
		_w158_,
		_w169_
	);
	LUT2 #(
		.INIT('h8)
	) name161 (
		_w42_,
		_w158_,
		_w170_
	);
	LUT2 #(
		.INIT('h8)
	) name162 (
		_w44_,
		_w158_,
		_w171_
	);
	LUT2 #(
		.INIT('h8)
	) name163 (
		_w46_,
		_w158_,
		_w172_
	);
	LUT2 #(
		.INIT('h8)
	) name164 (
		_w48_,
		_w158_,
		_w173_
	);
	LUT2 #(
		.INIT('h8)
	) name165 (
		_w50_,
		_w158_,
		_w174_
	);
	LUT2 #(
		.INIT('h1)
	) name166 (
		\count[6] ,
		\count[7] ,
		_w175_
	);
	LUT2 #(
		.INIT('h8)
	) name167 (
		_w9_,
		_w175_,
		_w176_
	);
	LUT2 #(
		.INIT('h8)
	) name168 (
		_w14_,
		_w176_,
		_w177_
	);
	LUT2 #(
		.INIT('h8)
	) name169 (
		_w17_,
		_w176_,
		_w178_
	);
	LUT2 #(
		.INIT('h8)
	) name170 (
		_w20_,
		_w176_,
		_w179_
	);
	LUT2 #(
		.INIT('h8)
	) name171 (
		_w22_,
		_w176_,
		_w180_
	);
	LUT2 #(
		.INIT('h8)
	) name172 (
		_w25_,
		_w176_,
		_w181_
	);
	LUT2 #(
		.INIT('h8)
	) name173 (
		_w28_,
		_w176_,
		_w182_
	);
	LUT2 #(
		.INIT('h8)
	) name174 (
		_w30_,
		_w176_,
		_w183_
	);
	LUT2 #(
		.INIT('h8)
	) name175 (
		_w32_,
		_w176_,
		_w184_
	);
	LUT2 #(
		.INIT('h8)
	) name176 (
		_w35_,
		_w176_,
		_w185_
	);
	LUT2 #(
		.INIT('h8)
	) name177 (
		_w37_,
		_w176_,
		_w186_
	);
	LUT2 #(
		.INIT('h8)
	) name178 (
		_w40_,
		_w176_,
		_w187_
	);
	LUT2 #(
		.INIT('h8)
	) name179 (
		_w42_,
		_w176_,
		_w188_
	);
	LUT2 #(
		.INIT('h8)
	) name180 (
		_w44_,
		_w176_,
		_w189_
	);
	LUT2 #(
		.INIT('h8)
	) name181 (
		_w46_,
		_w176_,
		_w190_
	);
	LUT2 #(
		.INIT('h8)
	) name182 (
		_w48_,
		_w176_,
		_w191_
	);
	LUT2 #(
		.INIT('h8)
	) name183 (
		_w50_,
		_w176_,
		_w192_
	);
	LUT2 #(
		.INIT('h8)
	) name184 (
		_w52_,
		_w175_,
		_w193_
	);
	LUT2 #(
		.INIT('h8)
	) name185 (
		_w14_,
		_w193_,
		_w194_
	);
	LUT2 #(
		.INIT('h8)
	) name186 (
		_w17_,
		_w193_,
		_w195_
	);
	LUT2 #(
		.INIT('h8)
	) name187 (
		_w20_,
		_w193_,
		_w196_
	);
	LUT2 #(
		.INIT('h8)
	) name188 (
		_w22_,
		_w193_,
		_w197_
	);
	LUT2 #(
		.INIT('h8)
	) name189 (
		_w25_,
		_w193_,
		_w198_
	);
	LUT2 #(
		.INIT('h8)
	) name190 (
		_w28_,
		_w193_,
		_w199_
	);
	LUT2 #(
		.INIT('h8)
	) name191 (
		_w30_,
		_w193_,
		_w200_
	);
	LUT2 #(
		.INIT('h8)
	) name192 (
		_w32_,
		_w193_,
		_w201_
	);
	LUT2 #(
		.INIT('h8)
	) name193 (
		_w35_,
		_w193_,
		_w202_
	);
	LUT2 #(
		.INIT('h8)
	) name194 (
		_w37_,
		_w193_,
		_w203_
	);
	LUT2 #(
		.INIT('h8)
	) name195 (
		_w40_,
		_w193_,
		_w204_
	);
	LUT2 #(
		.INIT('h8)
	) name196 (
		_w42_,
		_w193_,
		_w205_
	);
	LUT2 #(
		.INIT('h8)
	) name197 (
		_w44_,
		_w193_,
		_w206_
	);
	LUT2 #(
		.INIT('h8)
	) name198 (
		_w46_,
		_w193_,
		_w207_
	);
	LUT2 #(
		.INIT('h8)
	) name199 (
		_w48_,
		_w193_,
		_w208_
	);
	LUT2 #(
		.INIT('h8)
	) name200 (
		_w50_,
		_w193_,
		_w209_
	);
	LUT2 #(
		.INIT('h8)
	) name201 (
		_w70_,
		_w175_,
		_w210_
	);
	LUT2 #(
		.INIT('h8)
	) name202 (
		_w14_,
		_w210_,
		_w211_
	);
	LUT2 #(
		.INIT('h8)
	) name203 (
		_w17_,
		_w210_,
		_w212_
	);
	LUT2 #(
		.INIT('h8)
	) name204 (
		_w20_,
		_w210_,
		_w213_
	);
	LUT2 #(
		.INIT('h8)
	) name205 (
		_w22_,
		_w210_,
		_w214_
	);
	LUT2 #(
		.INIT('h8)
	) name206 (
		_w25_,
		_w210_,
		_w215_
	);
	LUT2 #(
		.INIT('h8)
	) name207 (
		_w28_,
		_w210_,
		_w216_
	);
	LUT2 #(
		.INIT('h8)
	) name208 (
		_w30_,
		_w210_,
		_w217_
	);
	LUT2 #(
		.INIT('h8)
	) name209 (
		_w32_,
		_w210_,
		_w218_
	);
	LUT2 #(
		.INIT('h8)
	) name210 (
		_w35_,
		_w210_,
		_w219_
	);
	LUT2 #(
		.INIT('h8)
	) name211 (
		_w37_,
		_w210_,
		_w220_
	);
	LUT2 #(
		.INIT('h8)
	) name212 (
		_w40_,
		_w210_,
		_w221_
	);
	LUT2 #(
		.INIT('h8)
	) name213 (
		_w42_,
		_w210_,
		_w222_
	);
	LUT2 #(
		.INIT('h8)
	) name214 (
		_w44_,
		_w210_,
		_w223_
	);
	LUT2 #(
		.INIT('h8)
	) name215 (
		_w46_,
		_w210_,
		_w224_
	);
	LUT2 #(
		.INIT('h8)
	) name216 (
		_w48_,
		_w210_,
		_w225_
	);
	LUT2 #(
		.INIT('h8)
	) name217 (
		_w50_,
		_w210_,
		_w226_
	);
	LUT2 #(
		.INIT('h8)
	) name218 (
		_w88_,
		_w175_,
		_w227_
	);
	LUT2 #(
		.INIT('h8)
	) name219 (
		_w14_,
		_w227_,
		_w228_
	);
	LUT2 #(
		.INIT('h8)
	) name220 (
		_w17_,
		_w227_,
		_w229_
	);
	LUT2 #(
		.INIT('h8)
	) name221 (
		_w20_,
		_w227_,
		_w230_
	);
	LUT2 #(
		.INIT('h8)
	) name222 (
		_w22_,
		_w227_,
		_w231_
	);
	LUT2 #(
		.INIT('h8)
	) name223 (
		_w25_,
		_w227_,
		_w232_
	);
	LUT2 #(
		.INIT('h8)
	) name224 (
		_w28_,
		_w227_,
		_w233_
	);
	LUT2 #(
		.INIT('h8)
	) name225 (
		_w30_,
		_w227_,
		_w234_
	);
	LUT2 #(
		.INIT('h8)
	) name226 (
		_w32_,
		_w227_,
		_w235_
	);
	LUT2 #(
		.INIT('h8)
	) name227 (
		_w35_,
		_w227_,
		_w236_
	);
	LUT2 #(
		.INIT('h8)
	) name228 (
		_w37_,
		_w227_,
		_w237_
	);
	LUT2 #(
		.INIT('h8)
	) name229 (
		_w40_,
		_w227_,
		_w238_
	);
	LUT2 #(
		.INIT('h8)
	) name230 (
		_w42_,
		_w227_,
		_w239_
	);
	LUT2 #(
		.INIT('h8)
	) name231 (
		_w44_,
		_w227_,
		_w240_
	);
	LUT2 #(
		.INIT('h8)
	) name232 (
		_w46_,
		_w227_,
		_w241_
	);
	LUT2 #(
		.INIT('h8)
	) name233 (
		_w48_,
		_w227_,
		_w242_
	);
	LUT2 #(
		.INIT('h8)
	) name234 (
		_w50_,
		_w227_,
		_w243_
	);
	LUT2 #(
		.INIT('h2)
	) name235 (
		\count[6] ,
		\count[7] ,
		_w244_
	);
	LUT2 #(
		.INIT('h8)
	) name236 (
		_w9_,
		_w244_,
		_w245_
	);
	LUT2 #(
		.INIT('h8)
	) name237 (
		_w14_,
		_w245_,
		_w246_
	);
	LUT2 #(
		.INIT('h8)
	) name238 (
		_w17_,
		_w245_,
		_w247_
	);
	LUT2 #(
		.INIT('h8)
	) name239 (
		_w20_,
		_w245_,
		_w248_
	);
	LUT2 #(
		.INIT('h8)
	) name240 (
		_w22_,
		_w245_,
		_w249_
	);
	LUT2 #(
		.INIT('h8)
	) name241 (
		_w25_,
		_w245_,
		_w250_
	);
	LUT2 #(
		.INIT('h8)
	) name242 (
		_w28_,
		_w245_,
		_w251_
	);
	LUT2 #(
		.INIT('h8)
	) name243 (
		_w30_,
		_w245_,
		_w252_
	);
	LUT2 #(
		.INIT('h8)
	) name244 (
		_w32_,
		_w245_,
		_w253_
	);
	LUT2 #(
		.INIT('h8)
	) name245 (
		_w35_,
		_w245_,
		_w254_
	);
	LUT2 #(
		.INIT('h8)
	) name246 (
		_w37_,
		_w245_,
		_w255_
	);
	LUT2 #(
		.INIT('h8)
	) name247 (
		_w40_,
		_w245_,
		_w256_
	);
	LUT2 #(
		.INIT('h8)
	) name248 (
		_w42_,
		_w245_,
		_w257_
	);
	LUT2 #(
		.INIT('h8)
	) name249 (
		_w44_,
		_w245_,
		_w258_
	);
	LUT2 #(
		.INIT('h8)
	) name250 (
		_w46_,
		_w245_,
		_w259_
	);
	LUT2 #(
		.INIT('h8)
	) name251 (
		_w48_,
		_w245_,
		_w260_
	);
	LUT2 #(
		.INIT('h8)
	) name252 (
		_w50_,
		_w245_,
		_w261_
	);
	LUT2 #(
		.INIT('h8)
	) name253 (
		_w52_,
		_w244_,
		_w262_
	);
	LUT2 #(
		.INIT('h8)
	) name254 (
		_w14_,
		_w262_,
		_w263_
	);
	LUT2 #(
		.INIT('h8)
	) name255 (
		_w17_,
		_w262_,
		_w264_
	);
	LUT2 #(
		.INIT('h8)
	) name256 (
		_w20_,
		_w262_,
		_w265_
	);
	LUT2 #(
		.INIT('h8)
	) name257 (
		_w22_,
		_w262_,
		_w266_
	);
	LUT2 #(
		.INIT('h8)
	) name258 (
		_w25_,
		_w262_,
		_w267_
	);
	LUT2 #(
		.INIT('h8)
	) name259 (
		_w28_,
		_w262_,
		_w268_
	);
	LUT2 #(
		.INIT('h8)
	) name260 (
		_w30_,
		_w262_,
		_w269_
	);
	LUT2 #(
		.INIT('h8)
	) name261 (
		_w32_,
		_w262_,
		_w270_
	);
	LUT2 #(
		.INIT('h8)
	) name262 (
		_w35_,
		_w262_,
		_w271_
	);
	LUT2 #(
		.INIT('h8)
	) name263 (
		_w37_,
		_w262_,
		_w272_
	);
	LUT2 #(
		.INIT('h8)
	) name264 (
		_w40_,
		_w262_,
		_w273_
	);
	LUT2 #(
		.INIT('h8)
	) name265 (
		_w42_,
		_w262_,
		_w274_
	);
	LUT2 #(
		.INIT('h8)
	) name266 (
		_w44_,
		_w262_,
		_w275_
	);
	LUT2 #(
		.INIT('h8)
	) name267 (
		_w46_,
		_w262_,
		_w276_
	);
	LUT2 #(
		.INIT('h8)
	) name268 (
		_w48_,
		_w262_,
		_w277_
	);
	LUT2 #(
		.INIT('h8)
	) name269 (
		_w50_,
		_w262_,
		_w278_
	);
	LUT2 #(
		.INIT('h8)
	) name270 (
		_w70_,
		_w244_,
		_w279_
	);
	LUT2 #(
		.INIT('h8)
	) name271 (
		_w14_,
		_w279_,
		_w280_
	);
	LUT2 #(
		.INIT('h8)
	) name272 (
		_w17_,
		_w279_,
		_w281_
	);
	LUT2 #(
		.INIT('h8)
	) name273 (
		_w20_,
		_w279_,
		_w282_
	);
	LUT2 #(
		.INIT('h8)
	) name274 (
		_w22_,
		_w279_,
		_w283_
	);
	LUT2 #(
		.INIT('h8)
	) name275 (
		_w25_,
		_w279_,
		_w284_
	);
	LUT2 #(
		.INIT('h8)
	) name276 (
		_w28_,
		_w279_,
		_w285_
	);
	LUT2 #(
		.INIT('h8)
	) name277 (
		_w30_,
		_w279_,
		_w286_
	);
	LUT2 #(
		.INIT('h8)
	) name278 (
		_w32_,
		_w279_,
		_w287_
	);
	LUT2 #(
		.INIT('h8)
	) name279 (
		_w35_,
		_w279_,
		_w288_
	);
	LUT2 #(
		.INIT('h8)
	) name280 (
		_w37_,
		_w279_,
		_w289_
	);
	LUT2 #(
		.INIT('h8)
	) name281 (
		_w40_,
		_w279_,
		_w290_
	);
	LUT2 #(
		.INIT('h8)
	) name282 (
		_w42_,
		_w279_,
		_w291_
	);
	LUT2 #(
		.INIT('h8)
	) name283 (
		_w44_,
		_w279_,
		_w292_
	);
	LUT2 #(
		.INIT('h8)
	) name284 (
		_w46_,
		_w279_,
		_w293_
	);
	LUT2 #(
		.INIT('h8)
	) name285 (
		_w48_,
		_w279_,
		_w294_
	);
	LUT2 #(
		.INIT('h8)
	) name286 (
		_w50_,
		_w279_,
		_w295_
	);
	LUT2 #(
		.INIT('h8)
	) name287 (
		_w88_,
		_w244_,
		_w296_
	);
	LUT2 #(
		.INIT('h8)
	) name288 (
		_w14_,
		_w296_,
		_w297_
	);
	LUT2 #(
		.INIT('h8)
	) name289 (
		_w17_,
		_w296_,
		_w298_
	);
	LUT2 #(
		.INIT('h8)
	) name290 (
		_w20_,
		_w296_,
		_w299_
	);
	LUT2 #(
		.INIT('h8)
	) name291 (
		_w22_,
		_w296_,
		_w300_
	);
	LUT2 #(
		.INIT('h8)
	) name292 (
		_w25_,
		_w296_,
		_w301_
	);
	LUT2 #(
		.INIT('h8)
	) name293 (
		_w28_,
		_w296_,
		_w302_
	);
	LUT2 #(
		.INIT('h8)
	) name294 (
		_w30_,
		_w296_,
		_w303_
	);
	LUT2 #(
		.INIT('h8)
	) name295 (
		_w32_,
		_w296_,
		_w304_
	);
	LUT2 #(
		.INIT('h8)
	) name296 (
		_w35_,
		_w296_,
		_w305_
	);
	LUT2 #(
		.INIT('h8)
	) name297 (
		_w37_,
		_w296_,
		_w306_
	);
	LUT2 #(
		.INIT('h8)
	) name298 (
		_w40_,
		_w296_,
		_w307_
	);
	LUT2 #(
		.INIT('h8)
	) name299 (
		_w42_,
		_w296_,
		_w308_
	);
	LUT2 #(
		.INIT('h8)
	) name300 (
		_w44_,
		_w296_,
		_w309_
	);
	LUT2 #(
		.INIT('h8)
	) name301 (
		_w46_,
		_w296_,
		_w310_
	);
	LUT2 #(
		.INIT('h8)
	) name302 (
		_w48_,
		_w296_,
		_w311_
	);
	LUT2 #(
		.INIT('h8)
	) name303 (
		_w50_,
		_w296_,
		_w312_
	);
	assign \selectp1[0]  = _w15_ ;
	assign \selectp1[1]  = _w18_ ;
	assign \selectp1[2]  = _w21_ ;
	assign \selectp1[3]  = _w23_ ;
	assign \selectp1[4]  = _w26_ ;
	assign \selectp1[5]  = _w29_ ;
	assign \selectp1[6]  = _w31_ ;
	assign \selectp1[7]  = _w33_ ;
	assign \selectp1[8]  = _w36_ ;
	assign \selectp1[9]  = _w38_ ;
	assign \selectp1[10]  = _w41_ ;
	assign \selectp1[11]  = _w43_ ;
	assign \selectp1[12]  = _w45_ ;
	assign \selectp1[13]  = _w47_ ;
	assign \selectp1[14]  = _w49_ ;
	assign \selectp1[15]  = _w51_ ;
	assign \selectp1[16]  = _w54_ ;
	assign \selectp1[17]  = _w55_ ;
	assign \selectp1[18]  = _w56_ ;
	assign \selectp1[19]  = _w57_ ;
	assign \selectp1[20]  = _w58_ ;
	assign \selectp1[21]  = _w59_ ;
	assign \selectp1[22]  = _w60_ ;
	assign \selectp1[23]  = _w61_ ;
	assign \selectp1[24]  = _w62_ ;
	assign \selectp1[25]  = _w63_ ;
	assign \selectp1[26]  = _w64_ ;
	assign \selectp1[27]  = _w65_ ;
	assign \selectp1[28]  = _w66_ ;
	assign \selectp1[29]  = _w67_ ;
	assign \selectp1[30]  = _w68_ ;
	assign \selectp1[31]  = _w69_ ;
	assign \selectp1[32]  = _w72_ ;
	assign \selectp1[33]  = _w73_ ;
	assign \selectp1[34]  = _w74_ ;
	assign \selectp1[35]  = _w75_ ;
	assign \selectp1[36]  = _w76_ ;
	assign \selectp1[37]  = _w77_ ;
	assign \selectp1[38]  = _w78_ ;
	assign \selectp1[39]  = _w79_ ;
	assign \selectp1[40]  = _w80_ ;
	assign \selectp1[41]  = _w81_ ;
	assign \selectp1[42]  = _w82_ ;
	assign \selectp1[43]  = _w83_ ;
	assign \selectp1[44]  = _w84_ ;
	assign \selectp1[45]  = _w85_ ;
	assign \selectp1[46]  = _w86_ ;
	assign \selectp1[47]  = _w87_ ;
	assign \selectp1[48]  = _w90_ ;
	assign \selectp1[49]  = _w91_ ;
	assign \selectp1[50]  = _w92_ ;
	assign \selectp1[51]  = _w93_ ;
	assign \selectp1[52]  = _w94_ ;
	assign \selectp1[53]  = _w95_ ;
	assign \selectp1[54]  = _w96_ ;
	assign \selectp1[55]  = _w97_ ;
	assign \selectp1[56]  = _w98_ ;
	assign \selectp1[57]  = _w99_ ;
	assign \selectp1[58]  = _w100_ ;
	assign \selectp1[59]  = _w101_ ;
	assign \selectp1[60]  = _w102_ ;
	assign \selectp1[61]  = _w103_ ;
	assign \selectp1[62]  = _w104_ ;
	assign \selectp1[63]  = _w105_ ;
	assign \selectp1[64]  = _w108_ ;
	assign \selectp1[65]  = _w109_ ;
	assign \selectp1[66]  = _w110_ ;
	assign \selectp1[67]  = _w111_ ;
	assign \selectp1[68]  = _w112_ ;
	assign \selectp1[69]  = _w113_ ;
	assign \selectp1[70]  = _w114_ ;
	assign \selectp1[71]  = _w115_ ;
	assign \selectp1[72]  = _w116_ ;
	assign \selectp1[73]  = _w117_ ;
	assign \selectp1[74]  = _w118_ ;
	assign \selectp1[75]  = _w119_ ;
	assign \selectp1[76]  = _w120_ ;
	assign \selectp1[77]  = _w121_ ;
	assign \selectp1[78]  = _w122_ ;
	assign \selectp1[79]  = _w123_ ;
	assign \selectp1[80]  = _w125_ ;
	assign \selectp1[81]  = _w126_ ;
	assign \selectp1[82]  = _w127_ ;
	assign \selectp1[83]  = _w128_ ;
	assign \selectp1[84]  = _w129_ ;
	assign \selectp1[85]  = _w130_ ;
	assign \selectp1[86]  = _w131_ ;
	assign \selectp1[87]  = _w132_ ;
	assign \selectp1[88]  = _w133_ ;
	assign \selectp1[89]  = _w134_ ;
	assign \selectp1[90]  = _w135_ ;
	assign \selectp1[91]  = _w136_ ;
	assign \selectp1[92]  = _w137_ ;
	assign \selectp1[93]  = _w138_ ;
	assign \selectp1[94]  = _w139_ ;
	assign \selectp1[95]  = _w140_ ;
	assign \selectp1[96]  = _w142_ ;
	assign \selectp1[97]  = _w143_ ;
	assign \selectp1[98]  = _w144_ ;
	assign \selectp1[99]  = _w145_ ;
	assign \selectp1[100]  = _w146_ ;
	assign \selectp1[101]  = _w147_ ;
	assign \selectp1[102]  = _w148_ ;
	assign \selectp1[103]  = _w149_ ;
	assign \selectp1[104]  = _w150_ ;
	assign \selectp1[105]  = _w151_ ;
	assign \selectp1[106]  = _w152_ ;
	assign \selectp1[107]  = _w153_ ;
	assign \selectp1[108]  = _w154_ ;
	assign \selectp1[109]  = _w155_ ;
	assign \selectp1[110]  = _w156_ ;
	assign \selectp1[111]  = _w157_ ;
	assign \selectp1[112]  = _w159_ ;
	assign \selectp1[113]  = _w160_ ;
	assign \selectp1[114]  = _w161_ ;
	assign \selectp1[115]  = _w162_ ;
	assign \selectp1[116]  = _w163_ ;
	assign \selectp1[117]  = _w164_ ;
	assign \selectp1[118]  = _w165_ ;
	assign \selectp1[119]  = _w166_ ;
	assign \selectp1[120]  = _w167_ ;
	assign \selectp1[121]  = _w168_ ;
	assign \selectp1[122]  = _w169_ ;
	assign \selectp1[123]  = _w170_ ;
	assign \selectp1[124]  = _w171_ ;
	assign \selectp1[125]  = _w172_ ;
	assign \selectp1[126]  = _w173_ ;
	assign \selectp1[127]  = _w174_ ;
	assign \selectp2[0]  = _w177_ ;
	assign \selectp2[1]  = _w178_ ;
	assign \selectp2[2]  = _w179_ ;
	assign \selectp2[3]  = _w180_ ;
	assign \selectp2[4]  = _w181_ ;
	assign \selectp2[5]  = _w182_ ;
	assign \selectp2[6]  = _w183_ ;
	assign \selectp2[7]  = _w184_ ;
	assign \selectp2[8]  = _w185_ ;
	assign \selectp2[9]  = _w186_ ;
	assign \selectp2[10]  = _w187_ ;
	assign \selectp2[11]  = _w188_ ;
	assign \selectp2[12]  = _w189_ ;
	assign \selectp2[13]  = _w190_ ;
	assign \selectp2[14]  = _w191_ ;
	assign \selectp2[15]  = _w192_ ;
	assign \selectp2[16]  = _w194_ ;
	assign \selectp2[17]  = _w195_ ;
	assign \selectp2[18]  = _w196_ ;
	assign \selectp2[19]  = _w197_ ;
	assign \selectp2[20]  = _w198_ ;
	assign \selectp2[21]  = _w199_ ;
	assign \selectp2[22]  = _w200_ ;
	assign \selectp2[23]  = _w201_ ;
	assign \selectp2[24]  = _w202_ ;
	assign \selectp2[25]  = _w203_ ;
	assign \selectp2[26]  = _w204_ ;
	assign \selectp2[27]  = _w205_ ;
	assign \selectp2[28]  = _w206_ ;
	assign \selectp2[29]  = _w207_ ;
	assign \selectp2[30]  = _w208_ ;
	assign \selectp2[31]  = _w209_ ;
	assign \selectp2[32]  = _w211_ ;
	assign \selectp2[33]  = _w212_ ;
	assign \selectp2[34]  = _w213_ ;
	assign \selectp2[35]  = _w214_ ;
	assign \selectp2[36]  = _w215_ ;
	assign \selectp2[37]  = _w216_ ;
	assign \selectp2[38]  = _w217_ ;
	assign \selectp2[39]  = _w218_ ;
	assign \selectp2[40]  = _w219_ ;
	assign \selectp2[41]  = _w220_ ;
	assign \selectp2[42]  = _w221_ ;
	assign \selectp2[43]  = _w222_ ;
	assign \selectp2[44]  = _w223_ ;
	assign \selectp2[45]  = _w224_ ;
	assign \selectp2[46]  = _w225_ ;
	assign \selectp2[47]  = _w226_ ;
	assign \selectp2[48]  = _w228_ ;
	assign \selectp2[49]  = _w229_ ;
	assign \selectp2[50]  = _w230_ ;
	assign \selectp2[51]  = _w231_ ;
	assign \selectp2[52]  = _w232_ ;
	assign \selectp2[53]  = _w233_ ;
	assign \selectp2[54]  = _w234_ ;
	assign \selectp2[55]  = _w235_ ;
	assign \selectp2[56]  = _w236_ ;
	assign \selectp2[57]  = _w237_ ;
	assign \selectp2[58]  = _w238_ ;
	assign \selectp2[59]  = _w239_ ;
	assign \selectp2[60]  = _w240_ ;
	assign \selectp2[61]  = _w241_ ;
	assign \selectp2[62]  = _w242_ ;
	assign \selectp2[63]  = _w243_ ;
	assign \selectp2[64]  = _w246_ ;
	assign \selectp2[65]  = _w247_ ;
	assign \selectp2[66]  = _w248_ ;
	assign \selectp2[67]  = _w249_ ;
	assign \selectp2[68]  = _w250_ ;
	assign \selectp2[69]  = _w251_ ;
	assign \selectp2[70]  = _w252_ ;
	assign \selectp2[71]  = _w253_ ;
	assign \selectp2[72]  = _w254_ ;
	assign \selectp2[73]  = _w255_ ;
	assign \selectp2[74]  = _w256_ ;
	assign \selectp2[75]  = _w257_ ;
	assign \selectp2[76]  = _w258_ ;
	assign \selectp2[77]  = _w259_ ;
	assign \selectp2[78]  = _w260_ ;
	assign \selectp2[79]  = _w261_ ;
	assign \selectp2[80]  = _w263_ ;
	assign \selectp2[81]  = _w264_ ;
	assign \selectp2[82]  = _w265_ ;
	assign \selectp2[83]  = _w266_ ;
	assign \selectp2[84]  = _w267_ ;
	assign \selectp2[85]  = _w268_ ;
	assign \selectp2[86]  = _w269_ ;
	assign \selectp2[87]  = _w270_ ;
	assign \selectp2[88]  = _w271_ ;
	assign \selectp2[89]  = _w272_ ;
	assign \selectp2[90]  = _w273_ ;
	assign \selectp2[91]  = _w274_ ;
	assign \selectp2[92]  = _w275_ ;
	assign \selectp2[93]  = _w276_ ;
	assign \selectp2[94]  = _w277_ ;
	assign \selectp2[95]  = _w278_ ;
	assign \selectp2[96]  = _w280_ ;
	assign \selectp2[97]  = _w281_ ;
	assign \selectp2[98]  = _w282_ ;
	assign \selectp2[99]  = _w283_ ;
	assign \selectp2[100]  = _w284_ ;
	assign \selectp2[101]  = _w285_ ;
	assign \selectp2[102]  = _w286_ ;
	assign \selectp2[103]  = _w287_ ;
	assign \selectp2[104]  = _w288_ ;
	assign \selectp2[105]  = _w289_ ;
	assign \selectp2[106]  = _w290_ ;
	assign \selectp2[107]  = _w291_ ;
	assign \selectp2[108]  = _w292_ ;
	assign \selectp2[109]  = _w293_ ;
	assign \selectp2[110]  = _w294_ ;
	assign \selectp2[111]  = _w295_ ;
	assign \selectp2[112]  = _w297_ ;
	assign \selectp2[113]  = _w298_ ;
	assign \selectp2[114]  = _w299_ ;
	assign \selectp2[115]  = _w300_ ;
	assign \selectp2[116]  = _w301_ ;
	assign \selectp2[117]  = _w302_ ;
	assign \selectp2[118]  = _w303_ ;
	assign \selectp2[119]  = _w304_ ;
	assign \selectp2[120]  = _w305_ ;
	assign \selectp2[121]  = _w306_ ;
	assign \selectp2[122]  = _w307_ ;
	assign \selectp2[123]  = _w308_ ;
	assign \selectp2[124]  = _w309_ ;
	assign \selectp2[125]  = _w310_ ;
	assign \selectp2[126]  = _w311_ ;
	assign \selectp2[127]  = _w312_ ;
endmodule;