module top (\a0_pad , \a1_pad , \a2_pad , \a3_pad , \a4_pad , \b0_pad , \b1_pad , \b2_pad , \b3_pad , \b4_pad , \b5_pad , b_pad, \c0_pad , \c1_pad , \c2_pad , \c3_pad , \c4_pad , \c5_pad , c_pad, \d0_pad , \d1_pad , \d2_pad , \d3_pad , \d4_pad , \d5_pad , d_pad, \e0_pad , \e2_pad , \e3_pad , \e4_pad , \e5_pad , e_pad, \f0_pad , \f1_pad , \f2_pad , \f3_pad , \f4_pad , \f5_pad , f_pad, \g0_pad , \g1_pad , \g2_pad , \g3_pad , \g4_pad , g_pad, \h0_pad , \h1_pad , \h2_pad , \h3_pad , \h4_pad , \h5_pad , h_pad, \i0_pad , \i10_pad , \i1_pad , \i2_pad , \i3_pad , \i4_pad , \i5_pad , i_pad, \j0_pad , \j2_pad , \j3_pad , \j4_pad , \j5_pad , j_pad, \k0_pad , \k1_pad , \k2_pad , \k3_pad , \k4_pad , \k5_pad , k_pad, \l0_pad , \l1_pad , \l2_pad , \l3_pad , \l4_pad , \l5_pad , \l6_pad , l_pad, \m0_pad , \m1_pad , \m2_pad , \m3_pad , \m4_pad , \m5_pad , \m6_pad , m_pad, \n0_pad , \n1_pad , \n2_pad , \n3_pad , \n4_pad , \n5_pad , n_pad, \o0_pad , \o1_pad , \o2_pad , \o3_pad , \o4_pad , \o5_pad , o_pad, \p0_pad , \p10_pad , \p1_pad , \p2_pad , \p3_pad , \p4_pad , \p5_pad , p_pad, \q0_pad , \q1_pad , \q2_pad , \q3_pad , \q4_pad , \q5_pad , q_pad, \r0_pad , \r1_pad , \r2_pad , \r3_pad , \r4_pad , \r5_pad , \r6_pad , r_pad, \s0_pad , \s1_pad , \s2_pad , \s3_pad , \s4_pad , s_pad, \t0_pad , \t1_pad , \t2_pad , \t3_pad , \t4_pad , t_pad, \u0_pad , \u1_pad , \u2_pad , \u3_pad , \u4_pad , u_pad, \v0_pad , \v1_pad , \v2_pad , \v3_pad , \v4_pad , v_pad, \w0_pad , \w1_pad , \w2_pad , \w3_pad , \w4_pad , w_pad, \x0_pad , \x1_pad , \x2_pad , \x3_pad , \x4_pad , \y0_pad , \y1_pad , \y2_pad , \y3_pad , \y4_pad , \z0_pad , \z1_pad , \z2_pad , \z3_pad , \z4_pad , z_pad, \a10_pad , \a6_pad , \a7_pad , \a8_pad , \a9_pad , \b10_pad , \b6_pad , \b7_pad , \b8_pad , \b9_pad , \c10_pad , \c53 , \c6_pad , \c7_pad , \c8_pad , \c9_pad , \d10_pad , \d6_pad , \d7_pad , \d8_pad , \d9_pad , \e10_pad , \e6_pad , \e7_pad , \e8_pad , \e9_pad , \f10_pad , \f22 , \f6_pad , \f7_pad , \f8_pad , \f9_pad , \g10_pad , \g6_pad , \g7_pad , \g8_pad , \g9_pad , \h6_pad , \h7_pad , \h8_pad , \h9_pad , \i6_pad , \i7_pad , \i8_pad , \i9_pad , \j10_pad , \j6_pad , \j7_pad , \j8_pad , \j9_pad , \k10_pad , \k53 , \k6_pad , \k7_pad , \k8_pad , \k9_pad , \l10_pad , \l7_pad , \l8_pad , \l9_pad , \m10_pad , \m7_pad , \m8_pad , \m9_pad , \n10_pad , \n6_pad , \n7_pad , \n8_pad , \n9_pad , \o10_pad , \o6_pad , \o7_pad , \o8_pad , \o9_pad , \p6_pad , \p7_pad , \p8_pad , \p9_pad , \q10_pad , \q6_pad , \q7_pad , \q8_pad , \q9_pad , \r10_pad , \r7_pad , \r8_pad , \r9_pad , \s5_pad , \s7_pad , \s8_pad , \s9_pad , \t10_pad , \t5_pad , \t6_pad , \t7_pad , \t8_pad , \t9_pad , \u5_pad , \u7_pad , \u8_pad , \u9_pad , \v10_pad , \v5_pad , \v6_pad , \v7_pad , \v8_pad , \v9_pad , \w10_pad , \w5_pad , \w6_pad , \w7_pad , \w8_pad , \w9_pad , \x10_pad , \x21 , \x5_pad , \x6_pad , \x7_pad , \x8_pad , \x9_pad , \y10_pad , \y5_pad , \y6_pad , \y7_pad , \y8_pad , \y9_pad , \z5_pad , \z6_pad , \z7_pad , \z8_pad , \z9_pad );
	input \a0_pad  ;
	input \a1_pad  ;
	input \a2_pad  ;
	input \a3_pad  ;
	input \a4_pad  ;
	input \b0_pad  ;
	input \b1_pad  ;
	input \b2_pad  ;
	input \b3_pad  ;
	input \b4_pad  ;
	input \b5_pad  ;
	input b_pad ;
	input \c0_pad  ;
	input \c1_pad  ;
	input \c2_pad  ;
	input \c3_pad  ;
	input \c4_pad  ;
	input \c5_pad  ;
	input c_pad ;
	input \d0_pad  ;
	input \d1_pad  ;
	input \d2_pad  ;
	input \d3_pad  ;
	input \d4_pad  ;
	input \d5_pad  ;
	input d_pad ;
	input \e0_pad  ;
	input \e2_pad  ;
	input \e3_pad  ;
	input \e4_pad  ;
	input \e5_pad  ;
	input e_pad ;
	input \f0_pad  ;
	input \f1_pad  ;
	input \f2_pad  ;
	input \f3_pad  ;
	input \f4_pad  ;
	input \f5_pad  ;
	input f_pad ;
	input \g0_pad  ;
	input \g1_pad  ;
	input \g2_pad  ;
	input \g3_pad  ;
	input \g4_pad  ;
	input g_pad ;
	input \h0_pad  ;
	input \h1_pad  ;
	input \h2_pad  ;
	input \h3_pad  ;
	input \h4_pad  ;
	input \h5_pad  ;
	input h_pad ;
	input \i0_pad  ;
	input \i10_pad  ;
	input \i1_pad  ;
	input \i2_pad  ;
	input \i3_pad  ;
	input \i4_pad  ;
	input \i5_pad  ;
	input i_pad ;
	input \j0_pad  ;
	input \j2_pad  ;
	input \j3_pad  ;
	input \j4_pad  ;
	input \j5_pad  ;
	input j_pad ;
	input \k0_pad  ;
	input \k1_pad  ;
	input \k2_pad  ;
	input \k3_pad  ;
	input \k4_pad  ;
	input \k5_pad  ;
	input k_pad ;
	input \l0_pad  ;
	input \l1_pad  ;
	input \l2_pad  ;
	input \l3_pad  ;
	input \l4_pad  ;
	input \l5_pad  ;
	input \l6_pad  ;
	input l_pad ;
	input \m0_pad  ;
	input \m1_pad  ;
	input \m2_pad  ;
	input \m3_pad  ;
	input \m4_pad  ;
	input \m5_pad  ;
	input \m6_pad  ;
	input m_pad ;
	input \n0_pad  ;
	input \n1_pad  ;
	input \n2_pad  ;
	input \n3_pad  ;
	input \n4_pad  ;
	input \n5_pad  ;
	input n_pad ;
	input \o0_pad  ;
	input \o1_pad  ;
	input \o2_pad  ;
	input \o3_pad  ;
	input \o4_pad  ;
	input \o5_pad  ;
	input o_pad ;
	input \p0_pad  ;
	input \p10_pad  ;
	input \p1_pad  ;
	input \p2_pad  ;
	input \p3_pad  ;
	input \p4_pad  ;
	input \p5_pad  ;
	input p_pad ;
	input \q0_pad  ;
	input \q1_pad  ;
	input \q2_pad  ;
	input \q3_pad  ;
	input \q4_pad  ;
	input \q5_pad  ;
	input q_pad ;
	input \r0_pad  ;
	input \r1_pad  ;
	input \r2_pad  ;
	input \r3_pad  ;
	input \r4_pad  ;
	input \r5_pad  ;
	input \r6_pad  ;
	input r_pad ;
	input \s0_pad  ;
	input \s1_pad  ;
	input \s2_pad  ;
	input \s3_pad  ;
	input \s4_pad  ;
	input s_pad ;
	input \t0_pad  ;
	input \t1_pad  ;
	input \t2_pad  ;
	input \t3_pad  ;
	input \t4_pad  ;
	input t_pad ;
	input \u0_pad  ;
	input \u1_pad  ;
	input \u2_pad  ;
	input \u3_pad  ;
	input \u4_pad  ;
	input u_pad ;
	input \v0_pad  ;
	input \v1_pad  ;
	input \v2_pad  ;
	input \v3_pad  ;
	input \v4_pad  ;
	input v_pad ;
	input \w0_pad  ;
	input \w1_pad  ;
	input \w2_pad  ;
	input \w3_pad  ;
	input \w4_pad  ;
	input w_pad ;
	input \x0_pad  ;
	input \x1_pad  ;
	input \x2_pad  ;
	input \x3_pad  ;
	input \x4_pad  ;
	input \y0_pad  ;
	input \y1_pad  ;
	input \y2_pad  ;
	input \y3_pad  ;
	input \y4_pad  ;
	input \z0_pad  ;
	input \z1_pad  ;
	input \z2_pad  ;
	input \z3_pad  ;
	input \z4_pad  ;
	input z_pad ;
	output \a10_pad  ;
	output \a6_pad  ;
	output \a7_pad  ;
	output \a8_pad  ;
	output \a9_pad  ;
	output \b10_pad  ;
	output \b6_pad  ;
	output \b7_pad  ;
	output \b8_pad  ;
	output \b9_pad  ;
	output \c10_pad  ;
	output \c53  ;
	output \c6_pad  ;
	output \c7_pad  ;
	output \c8_pad  ;
	output \c9_pad  ;
	output \d10_pad  ;
	output \d6_pad  ;
	output \d7_pad  ;
	output \d8_pad  ;
	output \d9_pad  ;
	output \e10_pad  ;
	output \e6_pad  ;
	output \e7_pad  ;
	output \e8_pad  ;
	output \e9_pad  ;
	output \f10_pad  ;
	output \f22  ;
	output \f6_pad  ;
	output \f7_pad  ;
	output \f8_pad  ;
	output \f9_pad  ;
	output \g10_pad  ;
	output \g6_pad  ;
	output \g7_pad  ;
	output \g8_pad  ;
	output \g9_pad  ;
	output \h6_pad  ;
	output \h7_pad  ;
	output \h8_pad  ;
	output \h9_pad  ;
	output \i6_pad  ;
	output \i7_pad  ;
	output \i8_pad  ;
	output \i9_pad  ;
	output \j10_pad  ;
	output \j6_pad  ;
	output \j7_pad  ;
	output \j8_pad  ;
	output \j9_pad  ;
	output \k10_pad  ;
	output \k53  ;
	output \k6_pad  ;
	output \k7_pad  ;
	output \k8_pad  ;
	output \k9_pad  ;
	output \l10_pad  ;
	output \l7_pad  ;
	output \l8_pad  ;
	output \l9_pad  ;
	output \m10_pad  ;
	output \m7_pad  ;
	output \m8_pad  ;
	output \m9_pad  ;
	output \n10_pad  ;
	output \n6_pad  ;
	output \n7_pad  ;
	output \n8_pad  ;
	output \n9_pad  ;
	output \o10_pad  ;
	output \o6_pad  ;
	output \o7_pad  ;
	output \o8_pad  ;
	output \o9_pad  ;
	output \p6_pad  ;
	output \p7_pad  ;
	output \p8_pad  ;
	output \p9_pad  ;
	output \q10_pad  ;
	output \q6_pad  ;
	output \q7_pad  ;
	output \q8_pad  ;
	output \q9_pad  ;
	output \r10_pad  ;
	output \r7_pad  ;
	output \r8_pad  ;
	output \r9_pad  ;
	output \s5_pad  ;
	output \s7_pad  ;
	output \s8_pad  ;
	output \s9_pad  ;
	output \t10_pad  ;
	output \t5_pad  ;
	output \t6_pad  ;
	output \t7_pad  ;
	output \t8_pad  ;
	output \t9_pad  ;
	output \u5_pad  ;
	output \u7_pad  ;
	output \u8_pad  ;
	output \u9_pad  ;
	output \v10_pad  ;
	output \v5_pad  ;
	output \v6_pad  ;
	output \v7_pad  ;
	output \v8_pad  ;
	output \v9_pad  ;
	output \w10_pad  ;
	output \w5_pad  ;
	output \w6_pad  ;
	output \w7_pad  ;
	output \w8_pad  ;
	output \w9_pad  ;
	output \x10_pad  ;
	output \x21  ;
	output \x5_pad  ;
	output \x6_pad  ;
	output \x7_pad  ;
	output \x8_pad  ;
	output \x9_pad  ;
	output \y10_pad  ;
	output \y5_pad  ;
	output \y6_pad  ;
	output \y7_pad  ;
	output \y8_pad  ;
	output \y9_pad  ;
	output \z5_pad  ;
	output \z6_pad  ;
	output \z7_pad  ;
	output \z8_pad  ;
	output \z9_pad  ;
	wire _w1431_ ;
	wire _w1430_ ;
	wire _w1429_ ;
	wire _w1428_ ;
	wire _w1427_ ;
	wire _w1426_ ;
	wire _w1425_ ;
	wire _w1424_ ;
	wire _w1423_ ;
	wire _w1422_ ;
	wire _w1421_ ;
	wire _w1420_ ;
	wire _w1419_ ;
	wire _w1418_ ;
	wire _w1417_ ;
	wire _w1416_ ;
	wire _w1415_ ;
	wire _w1414_ ;
	wire _w1413_ ;
	wire _w1412_ ;
	wire _w1411_ ;
	wire _w1410_ ;
	wire _w1409_ ;
	wire _w1408_ ;
	wire _w1407_ ;
	wire _w1406_ ;
	wire _w1405_ ;
	wire _w1404_ ;
	wire _w1403_ ;
	wire _w1402_ ;
	wire _w1401_ ;
	wire _w1400_ ;
	wire _w1399_ ;
	wire _w1398_ ;
	wire _w1397_ ;
	wire _w1396_ ;
	wire _w1395_ ;
	wire _w1394_ ;
	wire _w1393_ ;
	wire _w1392_ ;
	wire _w1391_ ;
	wire _w1390_ ;
	wire _w1389_ ;
	wire _w1388_ ;
	wire _w1387_ ;
	wire _w1386_ ;
	wire _w1385_ ;
	wire _w1384_ ;
	wire _w1383_ ;
	wire _w1382_ ;
	wire _w1381_ ;
	wire _w1380_ ;
	wire _w1379_ ;
	wire _w1378_ ;
	wire _w1377_ ;
	wire _w1376_ ;
	wire _w1375_ ;
	wire _w1374_ ;
	wire _w1373_ ;
	wire _w1372_ ;
	wire _w1371_ ;
	wire _w1370_ ;
	wire _w1369_ ;
	wire _w1368_ ;
	wire _w1367_ ;
	wire _w1366_ ;
	wire _w1365_ ;
	wire _w1364_ ;
	wire _w1363_ ;
	wire _w1362_ ;
	wire _w1361_ ;
	wire _w1360_ ;
	wire _w1359_ ;
	wire _w1358_ ;
	wire _w1357_ ;
	wire _w1356_ ;
	wire _w1355_ ;
	wire _w1354_ ;
	wire _w1353_ ;
	wire _w1352_ ;
	wire _w1351_ ;
	wire _w1350_ ;
	wire _w1349_ ;
	wire _w1348_ ;
	wire _w1347_ ;
	wire _w1346_ ;
	wire _w1345_ ;
	wire _w1344_ ;
	wire _w1343_ ;
	wire _w1342_ ;
	wire _w1341_ ;
	wire _w1340_ ;
	wire _w1339_ ;
	wire _w1338_ ;
	wire _w1337_ ;
	wire _w1336_ ;
	wire _w1335_ ;
	wire _w1334_ ;
	wire _w1333_ ;
	wire _w1332_ ;
	wire _w1331_ ;
	wire _w1330_ ;
	wire _w1329_ ;
	wire _w1328_ ;
	wire _w1327_ ;
	wire _w1326_ ;
	wire _w1325_ ;
	wire _w1324_ ;
	wire _w1323_ ;
	wire _w1322_ ;
	wire _w1321_ ;
	wire _w1320_ ;
	wire _w1319_ ;
	wire _w1318_ ;
	wire _w1317_ ;
	wire _w1316_ ;
	wire _w1315_ ;
	wire _w1314_ ;
	wire _w1313_ ;
	wire _w1312_ ;
	wire _w1311_ ;
	wire _w1310_ ;
	wire _w1309_ ;
	wire _w1308_ ;
	wire _w1307_ ;
	wire _w1306_ ;
	wire _w1305_ ;
	wire _w1304_ ;
	wire _w1303_ ;
	wire _w1302_ ;
	wire _w1301_ ;
	wire _w1300_ ;
	wire _w1299_ ;
	wire _w1298_ ;
	wire _w1297_ ;
	wire _w1296_ ;
	wire _w1295_ ;
	wire _w1294_ ;
	wire _w1293_ ;
	wire _w1292_ ;
	wire _w1291_ ;
	wire _w1290_ ;
	wire _w1289_ ;
	wire _w1288_ ;
	wire _w1287_ ;
	wire _w1286_ ;
	wire _w1285_ ;
	wire _w1284_ ;
	wire _w1283_ ;
	wire _w1282_ ;
	wire _w713_ ;
	wire _w712_ ;
	wire _w711_ ;
	wire _w710_ ;
	wire _w709_ ;
	wire _w708_ ;
	wire _w707_ ;
	wire _w706_ ;
	wire _w705_ ;
	wire _w704_ ;
	wire _w703_ ;
	wire _w702_ ;
	wire _w701_ ;
	wire _w700_ ;
	wire _w699_ ;
	wire _w698_ ;
	wire _w697_ ;
	wire _w696_ ;
	wire _w695_ ;
	wire _w694_ ;
	wire _w693_ ;
	wire _w692_ ;
	wire _w691_ ;
	wire _w690_ ;
	wire _w689_ ;
	wire _w688_ ;
	wire _w687_ ;
	wire _w686_ ;
	wire _w685_ ;
	wire _w684_ ;
	wire _w683_ ;
	wire _w682_ ;
	wire _w681_ ;
	wire _w680_ ;
	wire _w679_ ;
	wire _w678_ ;
	wire _w677_ ;
	wire _w676_ ;
	wire _w675_ ;
	wire _w674_ ;
	wire _w673_ ;
	wire _w672_ ;
	wire _w671_ ;
	wire _w670_ ;
	wire _w669_ ;
	wire _w668_ ;
	wire _w667_ ;
	wire _w666_ ;
	wire _w665_ ;
	wire _w664_ ;
	wire _w663_ ;
	wire _w662_ ;
	wire _w661_ ;
	wire _w660_ ;
	wire _w659_ ;
	wire _w658_ ;
	wire _w657_ ;
	wire _w656_ ;
	wire _w655_ ;
	wire _w654_ ;
	wire _w653_ ;
	wire _w652_ ;
	wire _w651_ ;
	wire _w650_ ;
	wire _w649_ ;
	wire _w648_ ;
	wire _w647_ ;
	wire _w646_ ;
	wire _w645_ ;
	wire _w644_ ;
	wire _w643_ ;
	wire _w642_ ;
	wire _w641_ ;
	wire _w640_ ;
	wire _w639_ ;
	wire _w638_ ;
	wire _w637_ ;
	wire _w636_ ;
	wire _w635_ ;
	wire _w634_ ;
	wire _w633_ ;
	wire _w632_ ;
	wire _w631_ ;
	wire _w630_ ;
	wire _w629_ ;
	wire _w628_ ;
	wire _w627_ ;
	wire _w626_ ;
	wire _w625_ ;
	wire _w624_ ;
	wire _w623_ ;
	wire _w622_ ;
	wire _w621_ ;
	wire _w620_ ;
	wire _w619_ ;
	wire _w618_ ;
	wire _w617_ ;
	wire _w616_ ;
	wire _w615_ ;
	wire _w614_ ;
	wire _w613_ ;
	wire _w612_ ;
	wire _w611_ ;
	wire _w610_ ;
	wire _w609_ ;
	wire _w608_ ;
	wire _w607_ ;
	wire _w606_ ;
	wire _w605_ ;
	wire _w604_ ;
	wire _w603_ ;
	wire _w602_ ;
	wire _w601_ ;
	wire _w600_ ;
	wire _w599_ ;
	wire _w598_ ;
	wire _w597_ ;
	wire _w596_ ;
	wire _w595_ ;
	wire _w594_ ;
	wire _w593_ ;
	wire _w592_ ;
	wire _w591_ ;
	wire _w590_ ;
	wire _w589_ ;
	wire _w588_ ;
	wire _w587_ ;
	wire _w586_ ;
	wire _w585_ ;
	wire _w584_ ;
	wire _w583_ ;
	wire _w582_ ;
	wire _w581_ ;
	wire _w580_ ;
	wire _w579_ ;
	wire _w578_ ;
	wire _w577_ ;
	wire _w576_ ;
	wire _w575_ ;
	wire _w574_ ;
	wire _w573_ ;
	wire _w572_ ;
	wire _w571_ ;
	wire _w570_ ;
	wire _w569_ ;
	wire _w568_ ;
	wire _w567_ ;
	wire _w566_ ;
	wire _w565_ ;
	wire _w564_ ;
	wire _w563_ ;
	wire _w562_ ;
	wire _w561_ ;
	wire _w560_ ;
	wire _w559_ ;
	wire _w558_ ;
	wire _w557_ ;
	wire _w556_ ;
	wire _w555_ ;
	wire _w554_ ;
	wire _w553_ ;
	wire _w552_ ;
	wire _w551_ ;
	wire _w550_ ;
	wire _w549_ ;
	wire _w548_ ;
	wire _w547_ ;
	wire _w546_ ;
	wire _w545_ ;
	wire _w544_ ;
	wire _w543_ ;
	wire _w542_ ;
	wire _w541_ ;
	wire _w540_ ;
	wire _w539_ ;
	wire _w538_ ;
	wire _w537_ ;
	wire _w536_ ;
	wire _w535_ ;
	wire _w534_ ;
	wire _w533_ ;
	wire _w532_ ;
	wire _w531_ ;
	wire _w530_ ;
	wire _w529_ ;
	wire _w528_ ;
	wire _w527_ ;
	wire _w526_ ;
	wire _w525_ ;
	wire _w524_ ;
	wire _w523_ ;
	wire _w522_ ;
	wire _w521_ ;
	wire _w520_ ;
	wire _w519_ ;
	wire _w518_ ;
	wire _w517_ ;
	wire _w516_ ;
	wire _w515_ ;
	wire _w514_ ;
	wire _w513_ ;
	wire _w512_ ;
	wire _w511_ ;
	wire _w510_ ;
	wire _w509_ ;
	wire _w508_ ;
	wire _w507_ ;
	wire _w506_ ;
	wire _w505_ ;
	wire _w504_ ;
	wire _w503_ ;
	wire _w502_ ;
	wire _w501_ ;
	wire _w500_ ;
	wire _w499_ ;
	wire _w498_ ;
	wire _w497_ ;
	wire _w496_ ;
	wire _w495_ ;
	wire _w494_ ;
	wire _w493_ ;
	wire _w492_ ;
	wire _w491_ ;
	wire _w490_ ;
	wire _w489_ ;
	wire _w488_ ;
	wire _w487_ ;
	wire _w486_ ;
	wire _w485_ ;
	wire _w484_ ;
	wire _w483_ ;
	wire _w482_ ;
	wire _w481_ ;
	wire _w480_ ;
	wire _w479_ ;
	wire _w478_ ;
	wire _w477_ ;
	wire _w476_ ;
	wire _w475_ ;
	wire _w474_ ;
	wire _w473_ ;
	wire _w472_ ;
	wire _w471_ ;
	wire _w470_ ;
	wire _w469_ ;
	wire _w468_ ;
	wire _w467_ ;
	wire _w466_ ;
	wire _w465_ ;
	wire _w464_ ;
	wire _w463_ ;
	wire _w462_ ;
	wire _w461_ ;
	wire _w460_ ;
	wire _w459_ ;
	wire _w458_ ;
	wire _w457_ ;
	wire _w456_ ;
	wire _w455_ ;
	wire _w454_ ;
	wire _w453_ ;
	wire _w452_ ;
	wire _w451_ ;
	wire _w450_ ;
	wire _w449_ ;
	wire _w448_ ;
	wire _w447_ ;
	wire _w446_ ;
	wire _w445_ ;
	wire _w444_ ;
	wire _w443_ ;
	wire _w442_ ;
	wire _w441_ ;
	wire _w440_ ;
	wire _w439_ ;
	wire _w438_ ;
	wire _w437_ ;
	wire _w436_ ;
	wire _w435_ ;
	wire _w434_ ;
	wire _w433_ ;
	wire _w432_ ;
	wire _w431_ ;
	wire _w430_ ;
	wire _w299_ ;
	wire _w298_ ;
	wire _w297_ ;
	wire _w296_ ;
	wire _w295_ ;
	wire _w294_ ;
	wire _w293_ ;
	wire _w292_ ;
	wire _w291_ ;
	wire _w290_ ;
	wire _w289_ ;
	wire _w288_ ;
	wire _w287_ ;
	wire _w286_ ;
	wire _w285_ ;
	wire _w284_ ;
	wire _w283_ ;
	wire _w282_ ;
	wire _w281_ ;
	wire _w280_ ;
	wire _w279_ ;
	wire _w278_ ;
	wire _w277_ ;
	wire _w276_ ;
	wire _w275_ ;
	wire _w274_ ;
	wire _w273_ ;
	wire _w272_ ;
	wire _w271_ ;
	wire _w270_ ;
	wire _w269_ ;
	wire _w268_ ;
	wire _w267_ ;
	wire _w266_ ;
	wire _w265_ ;
	wire _w264_ ;
	wire _w263_ ;
	wire _w262_ ;
	wire _w261_ ;
	wire _w260_ ;
	wire _w259_ ;
	wire _w258_ ;
	wire _w257_ ;
	wire _w256_ ;
	wire _w255_ ;
	wire _w254_ ;
	wire _w253_ ;
	wire _w252_ ;
	wire _w251_ ;
	wire _w250_ ;
	wire _w249_ ;
	wire _w248_ ;
	wire _w247_ ;
	wire _w246_ ;
	wire _w245_ ;
	wire _w244_ ;
	wire _w243_ ;
	wire _w242_ ;
	wire _w241_ ;
	wire _w240_ ;
	wire _w239_ ;
	wire _w238_ ;
	wire _w237_ ;
	wire _w236_ ;
	wire _w235_ ;
	wire _w234_ ;
	wire _w233_ ;
	wire _w232_ ;
	wire _w201_ ;
	wire _w200_ ;
	wire _w199_ ;
	wire _w198_ ;
	wire _w197_ ;
	wire _w196_ ;
	wire _w195_ ;
	wire _w194_ ;
	wire _w193_ ;
	wire _w192_ ;
	wire _w191_ ;
	wire _w190_ ;
	wire _w189_ ;
	wire _w188_ ;
	wire _w187_ ;
	wire _w186_ ;
	wire _w173_ ;
	wire _w174_ ;
	wire _w175_ ;
	wire _w176_ ;
	wire _w177_ ;
	wire _w178_ ;
	wire _w179_ ;
	wire _w180_ ;
	wire _w181_ ;
	wire _w182_ ;
	wire _w183_ ;
	wire _w184_ ;
	wire _w185_ ;
	wire _w202_ ;
	wire _w203_ ;
	wire _w204_ ;
	wire _w205_ ;
	wire _w206_ ;
	wire _w207_ ;
	wire _w208_ ;
	wire _w209_ ;
	wire _w210_ ;
	wire _w211_ ;
	wire _w212_ ;
	wire _w213_ ;
	wire _w214_ ;
	wire _w215_ ;
	wire _w216_ ;
	wire _w217_ ;
	wire _w218_ ;
	wire _w219_ ;
	wire _w220_ ;
	wire _w221_ ;
	wire _w222_ ;
	wire _w223_ ;
	wire _w224_ ;
	wire _w225_ ;
	wire _w226_ ;
	wire _w227_ ;
	wire _w228_ ;
	wire _w229_ ;
	wire _w230_ ;
	wire _w231_ ;
	wire _w300_ ;
	wire _w301_ ;
	wire _w302_ ;
	wire _w303_ ;
	wire _w304_ ;
	wire _w305_ ;
	wire _w306_ ;
	wire _w307_ ;
	wire _w308_ ;
	wire _w309_ ;
	wire _w310_ ;
	wire _w311_ ;
	wire _w312_ ;
	wire _w313_ ;
	wire _w314_ ;
	wire _w315_ ;
	wire _w316_ ;
	wire _w317_ ;
	wire _w318_ ;
	wire _w319_ ;
	wire _w320_ ;
	wire _w321_ ;
	wire _w322_ ;
	wire _w323_ ;
	wire _w324_ ;
	wire _w325_ ;
	wire _w326_ ;
	wire _w327_ ;
	wire _w328_ ;
	wire _w329_ ;
	wire _w330_ ;
	wire _w331_ ;
	wire _w332_ ;
	wire _w333_ ;
	wire _w334_ ;
	wire _w335_ ;
	wire _w336_ ;
	wire _w337_ ;
	wire _w338_ ;
	wire _w339_ ;
	wire _w340_ ;
	wire _w341_ ;
	wire _w342_ ;
	wire _w343_ ;
	wire _w344_ ;
	wire _w345_ ;
	wire _w346_ ;
	wire _w347_ ;
	wire _w348_ ;
	wire _w349_ ;
	wire _w350_ ;
	wire _w351_ ;
	wire _w352_ ;
	wire _w353_ ;
	wire _w354_ ;
	wire _w355_ ;
	wire _w356_ ;
	wire _w357_ ;
	wire _w358_ ;
	wire _w359_ ;
	wire _w360_ ;
	wire _w361_ ;
	wire _w362_ ;
	wire _w363_ ;
	wire _w364_ ;
	wire _w365_ ;
	wire _w366_ ;
	wire _w367_ ;
	wire _w368_ ;
	wire _w369_ ;
	wire _w370_ ;
	wire _w371_ ;
	wire _w372_ ;
	wire _w373_ ;
	wire _w374_ ;
	wire _w375_ ;
	wire _w376_ ;
	wire _w377_ ;
	wire _w378_ ;
	wire _w379_ ;
	wire _w380_ ;
	wire _w381_ ;
	wire _w382_ ;
	wire _w383_ ;
	wire _w384_ ;
	wire _w385_ ;
	wire _w386_ ;
	wire _w387_ ;
	wire _w388_ ;
	wire _w389_ ;
	wire _w390_ ;
	wire _w391_ ;
	wire _w392_ ;
	wire _w393_ ;
	wire _w394_ ;
	wire _w395_ ;
	wire _w396_ ;
	wire _w397_ ;
	wire _w398_ ;
	wire _w399_ ;
	wire _w400_ ;
	wire _w401_ ;
	wire _w402_ ;
	wire _w403_ ;
	wire _w404_ ;
	wire _w405_ ;
	wire _w406_ ;
	wire _w407_ ;
	wire _w408_ ;
	wire _w409_ ;
	wire _w410_ ;
	wire _w411_ ;
	wire _w412_ ;
	wire _w413_ ;
	wire _w414_ ;
	wire _w415_ ;
	wire _w416_ ;
	wire _w417_ ;
	wire _w418_ ;
	wire _w419_ ;
	wire _w420_ ;
	wire _w421_ ;
	wire _w422_ ;
	wire _w423_ ;
	wire _w424_ ;
	wire _w425_ ;
	wire _w426_ ;
	wire _w427_ ;
	wire _w428_ ;
	wire _w429_ ;
	wire _w714_ ;
	wire _w715_ ;
	wire _w716_ ;
	wire _w717_ ;
	wire _w718_ ;
	wire _w719_ ;
	wire _w720_ ;
	wire _w721_ ;
	wire _w722_ ;
	wire _w723_ ;
	wire _w724_ ;
	wire _w725_ ;
	wire _w726_ ;
	wire _w727_ ;
	wire _w728_ ;
	wire _w729_ ;
	wire _w730_ ;
	wire _w731_ ;
	wire _w732_ ;
	wire _w733_ ;
	wire _w734_ ;
	wire _w735_ ;
	wire _w736_ ;
	wire _w737_ ;
	wire _w738_ ;
	wire _w739_ ;
	wire _w740_ ;
	wire _w741_ ;
	wire _w742_ ;
	wire _w743_ ;
	wire _w744_ ;
	wire _w745_ ;
	wire _w746_ ;
	wire _w747_ ;
	wire _w748_ ;
	wire _w749_ ;
	wire _w750_ ;
	wire _w751_ ;
	wire _w752_ ;
	wire _w753_ ;
	wire _w754_ ;
	wire _w755_ ;
	wire _w756_ ;
	wire _w757_ ;
	wire _w758_ ;
	wire _w759_ ;
	wire _w760_ ;
	wire _w761_ ;
	wire _w762_ ;
	wire _w763_ ;
	wire _w764_ ;
	wire _w765_ ;
	wire _w766_ ;
	wire _w767_ ;
	wire _w768_ ;
	wire _w769_ ;
	wire _w770_ ;
	wire _w771_ ;
	wire _w772_ ;
	wire _w773_ ;
	wire _w774_ ;
	wire _w775_ ;
	wire _w776_ ;
	wire _w777_ ;
	wire _w778_ ;
	wire _w779_ ;
	wire _w780_ ;
	wire _w781_ ;
	wire _w782_ ;
	wire _w783_ ;
	wire _w784_ ;
	wire _w785_ ;
	wire _w786_ ;
	wire _w787_ ;
	wire _w788_ ;
	wire _w789_ ;
	wire _w790_ ;
	wire _w791_ ;
	wire _w792_ ;
	wire _w793_ ;
	wire _w794_ ;
	wire _w795_ ;
	wire _w796_ ;
	wire _w797_ ;
	wire _w798_ ;
	wire _w799_ ;
	wire _w800_ ;
	wire _w801_ ;
	wire _w802_ ;
	wire _w803_ ;
	wire _w804_ ;
	wire _w805_ ;
	wire _w806_ ;
	wire _w807_ ;
	wire _w808_ ;
	wire _w809_ ;
	wire _w810_ ;
	wire _w811_ ;
	wire _w812_ ;
	wire _w813_ ;
	wire _w814_ ;
	wire _w815_ ;
	wire _w816_ ;
	wire _w817_ ;
	wire _w818_ ;
	wire _w819_ ;
	wire _w820_ ;
	wire _w821_ ;
	wire _w822_ ;
	wire _w823_ ;
	wire _w824_ ;
	wire _w825_ ;
	wire _w826_ ;
	wire _w827_ ;
	wire _w828_ ;
	wire _w829_ ;
	wire _w830_ ;
	wire _w831_ ;
	wire _w832_ ;
	wire _w833_ ;
	wire _w834_ ;
	wire _w835_ ;
	wire _w836_ ;
	wire _w837_ ;
	wire _w838_ ;
	wire _w839_ ;
	wire _w840_ ;
	wire _w841_ ;
	wire _w842_ ;
	wire _w843_ ;
	wire _w844_ ;
	wire _w845_ ;
	wire _w846_ ;
	wire _w847_ ;
	wire _w848_ ;
	wire _w849_ ;
	wire _w850_ ;
	wire _w851_ ;
	wire _w852_ ;
	wire _w853_ ;
	wire _w854_ ;
	wire _w855_ ;
	wire _w856_ ;
	wire _w857_ ;
	wire _w858_ ;
	wire _w859_ ;
	wire _w860_ ;
	wire _w861_ ;
	wire _w862_ ;
	wire _w863_ ;
	wire _w864_ ;
	wire _w865_ ;
	wire _w866_ ;
	wire _w867_ ;
	wire _w868_ ;
	wire _w869_ ;
	wire _w870_ ;
	wire _w871_ ;
	wire _w872_ ;
	wire _w873_ ;
	wire _w874_ ;
	wire _w875_ ;
	wire _w876_ ;
	wire _w877_ ;
	wire _w878_ ;
	wire _w879_ ;
	wire _w880_ ;
	wire _w881_ ;
	wire _w882_ ;
	wire _w883_ ;
	wire _w884_ ;
	wire _w885_ ;
	wire _w886_ ;
	wire _w887_ ;
	wire _w888_ ;
	wire _w889_ ;
	wire _w890_ ;
	wire _w891_ ;
	wire _w892_ ;
	wire _w893_ ;
	wire _w894_ ;
	wire _w895_ ;
	wire _w896_ ;
	wire _w897_ ;
	wire _w898_ ;
	wire _w899_ ;
	wire _w900_ ;
	wire _w901_ ;
	wire _w902_ ;
	wire _w903_ ;
	wire _w904_ ;
	wire _w905_ ;
	wire _w906_ ;
	wire _w907_ ;
	wire _w908_ ;
	wire _w909_ ;
	wire _w910_ ;
	wire _w911_ ;
	wire _w912_ ;
	wire _w913_ ;
	wire _w914_ ;
	wire _w915_ ;
	wire _w916_ ;
	wire _w917_ ;
	wire _w918_ ;
	wire _w919_ ;
	wire _w920_ ;
	wire _w921_ ;
	wire _w922_ ;
	wire _w923_ ;
	wire _w924_ ;
	wire _w925_ ;
	wire _w926_ ;
	wire _w927_ ;
	wire _w928_ ;
	wire _w929_ ;
	wire _w930_ ;
	wire _w931_ ;
	wire _w932_ ;
	wire _w933_ ;
	wire _w934_ ;
	wire _w935_ ;
	wire _w936_ ;
	wire _w937_ ;
	wire _w938_ ;
	wire _w939_ ;
	wire _w940_ ;
	wire _w941_ ;
	wire _w942_ ;
	wire _w943_ ;
	wire _w944_ ;
	wire _w945_ ;
	wire _w946_ ;
	wire _w947_ ;
	wire _w948_ ;
	wire _w949_ ;
	wire _w950_ ;
	wire _w951_ ;
	wire _w952_ ;
	wire _w953_ ;
	wire _w954_ ;
	wire _w955_ ;
	wire _w956_ ;
	wire _w957_ ;
	wire _w958_ ;
	wire _w959_ ;
	wire _w960_ ;
	wire _w961_ ;
	wire _w962_ ;
	wire _w963_ ;
	wire _w964_ ;
	wire _w965_ ;
	wire _w966_ ;
	wire _w967_ ;
	wire _w968_ ;
	wire _w969_ ;
	wire _w970_ ;
	wire _w971_ ;
	wire _w972_ ;
	wire _w973_ ;
	wire _w974_ ;
	wire _w975_ ;
	wire _w976_ ;
	wire _w977_ ;
	wire _w978_ ;
	wire _w979_ ;
	wire _w980_ ;
	wire _w981_ ;
	wire _w982_ ;
	wire _w983_ ;
	wire _w984_ ;
	wire _w985_ ;
	wire _w986_ ;
	wire _w987_ ;
	wire _w988_ ;
	wire _w989_ ;
	wire _w990_ ;
	wire _w991_ ;
	wire _w992_ ;
	wire _w993_ ;
	wire _w994_ ;
	wire _w995_ ;
	wire _w996_ ;
	wire _w997_ ;
	wire _w998_ ;
	wire _w999_ ;
	wire _w1000_ ;
	wire _w1001_ ;
	wire _w1002_ ;
	wire _w1003_ ;
	wire _w1004_ ;
	wire _w1005_ ;
	wire _w1006_ ;
	wire _w1007_ ;
	wire _w1008_ ;
	wire _w1009_ ;
	wire _w1010_ ;
	wire _w1011_ ;
	wire _w1012_ ;
	wire _w1013_ ;
	wire _w1014_ ;
	wire _w1015_ ;
	wire _w1016_ ;
	wire _w1017_ ;
	wire _w1018_ ;
	wire _w1019_ ;
	wire _w1020_ ;
	wire _w1021_ ;
	wire _w1022_ ;
	wire _w1023_ ;
	wire _w1024_ ;
	wire _w1025_ ;
	wire _w1026_ ;
	wire _w1027_ ;
	wire _w1028_ ;
	wire _w1029_ ;
	wire _w1030_ ;
	wire _w1031_ ;
	wire _w1032_ ;
	wire _w1033_ ;
	wire _w1034_ ;
	wire _w1035_ ;
	wire _w1036_ ;
	wire _w1037_ ;
	wire _w1038_ ;
	wire _w1039_ ;
	wire _w1040_ ;
	wire _w1041_ ;
	wire _w1042_ ;
	wire _w1043_ ;
	wire _w1044_ ;
	wire _w1045_ ;
	wire _w1046_ ;
	wire _w1047_ ;
	wire _w1048_ ;
	wire _w1049_ ;
	wire _w1050_ ;
	wire _w1051_ ;
	wire _w1052_ ;
	wire _w1053_ ;
	wire _w1054_ ;
	wire _w1055_ ;
	wire _w1056_ ;
	wire _w1057_ ;
	wire _w1058_ ;
	wire _w1059_ ;
	wire _w1060_ ;
	wire _w1061_ ;
	wire _w1062_ ;
	wire _w1063_ ;
	wire _w1064_ ;
	wire _w1065_ ;
	wire _w1066_ ;
	wire _w1067_ ;
	wire _w1068_ ;
	wire _w1069_ ;
	wire _w1070_ ;
	wire _w1071_ ;
	wire _w1072_ ;
	wire _w1073_ ;
	wire _w1074_ ;
	wire _w1075_ ;
	wire _w1076_ ;
	wire _w1077_ ;
	wire _w1078_ ;
	wire _w1079_ ;
	wire _w1080_ ;
	wire _w1081_ ;
	wire _w1082_ ;
	wire _w1083_ ;
	wire _w1084_ ;
	wire _w1085_ ;
	wire _w1086_ ;
	wire _w1087_ ;
	wire _w1088_ ;
	wire _w1089_ ;
	wire _w1090_ ;
	wire _w1091_ ;
	wire _w1092_ ;
	wire _w1093_ ;
	wire _w1094_ ;
	wire _w1095_ ;
	wire _w1096_ ;
	wire _w1097_ ;
	wire _w1098_ ;
	wire _w1099_ ;
	wire _w1100_ ;
	wire _w1101_ ;
	wire _w1102_ ;
	wire _w1103_ ;
	wire _w1104_ ;
	wire _w1105_ ;
	wire _w1106_ ;
	wire _w1107_ ;
	wire _w1108_ ;
	wire _w1109_ ;
	wire _w1110_ ;
	wire _w1111_ ;
	wire _w1112_ ;
	wire _w1113_ ;
	wire _w1114_ ;
	wire _w1115_ ;
	wire _w1116_ ;
	wire _w1117_ ;
	wire _w1118_ ;
	wire _w1119_ ;
	wire _w1120_ ;
	wire _w1121_ ;
	wire _w1122_ ;
	wire _w1123_ ;
	wire _w1124_ ;
	wire _w1125_ ;
	wire _w1126_ ;
	wire _w1127_ ;
	wire _w1128_ ;
	wire _w1129_ ;
	wire _w1130_ ;
	wire _w1131_ ;
	wire _w1132_ ;
	wire _w1133_ ;
	wire _w1134_ ;
	wire _w1135_ ;
	wire _w1136_ ;
	wire _w1137_ ;
	wire _w1138_ ;
	wire _w1139_ ;
	wire _w1140_ ;
	wire _w1141_ ;
	wire _w1142_ ;
	wire _w1143_ ;
	wire _w1144_ ;
	wire _w1145_ ;
	wire _w1146_ ;
	wire _w1147_ ;
	wire _w1148_ ;
	wire _w1149_ ;
	wire _w1150_ ;
	wire _w1151_ ;
	wire _w1152_ ;
	wire _w1153_ ;
	wire _w1154_ ;
	wire _w1155_ ;
	wire _w1156_ ;
	wire _w1157_ ;
	wire _w1158_ ;
	wire _w1159_ ;
	wire _w1160_ ;
	wire _w1161_ ;
	wire _w1162_ ;
	wire _w1163_ ;
	wire _w1164_ ;
	wire _w1165_ ;
	wire _w1166_ ;
	wire _w1167_ ;
	wire _w1168_ ;
	wire _w1169_ ;
	wire _w1170_ ;
	wire _w1171_ ;
	wire _w1172_ ;
	wire _w1173_ ;
	wire _w1174_ ;
	wire _w1175_ ;
	wire _w1176_ ;
	wire _w1177_ ;
	wire _w1178_ ;
	wire _w1179_ ;
	wire _w1180_ ;
	wire _w1181_ ;
	wire _w1182_ ;
	wire _w1183_ ;
	wire _w1184_ ;
	wire _w1185_ ;
	wire _w1186_ ;
	wire _w1187_ ;
	wire _w1188_ ;
	wire _w1189_ ;
	wire _w1190_ ;
	wire _w1191_ ;
	wire _w1192_ ;
	wire _w1193_ ;
	wire _w1194_ ;
	wire _w1195_ ;
	wire _w1196_ ;
	wire _w1197_ ;
	wire _w1198_ ;
	wire _w1199_ ;
	wire _w1200_ ;
	wire _w1201_ ;
	wire _w1202_ ;
	wire _w1203_ ;
	wire _w1204_ ;
	wire _w1205_ ;
	wire _w1206_ ;
	wire _w1207_ ;
	wire _w1208_ ;
	wire _w1209_ ;
	wire _w1210_ ;
	wire _w1211_ ;
	wire _w1212_ ;
	wire _w1213_ ;
	wire _w1214_ ;
	wire _w1215_ ;
	wire _w1216_ ;
	wire _w1217_ ;
	wire _w1218_ ;
	wire _w1219_ ;
	wire _w1220_ ;
	wire _w1221_ ;
	wire _w1222_ ;
	wire _w1223_ ;
	wire _w1224_ ;
	wire _w1225_ ;
	wire _w1226_ ;
	wire _w1227_ ;
	wire _w1228_ ;
	wire _w1229_ ;
	wire _w1230_ ;
	wire _w1231_ ;
	wire _w1232_ ;
	wire _w1233_ ;
	wire _w1234_ ;
	wire _w1235_ ;
	wire _w1236_ ;
	wire _w1237_ ;
	wire _w1238_ ;
	wire _w1239_ ;
	wire _w1240_ ;
	wire _w1241_ ;
	wire _w1242_ ;
	wire _w1243_ ;
	wire _w1244_ ;
	wire _w1245_ ;
	wire _w1246_ ;
	wire _w1247_ ;
	wire _w1248_ ;
	wire _w1249_ ;
	wire _w1250_ ;
	wire _w1251_ ;
	wire _w1252_ ;
	wire _w1253_ ;
	wire _w1254_ ;
	wire _w1255_ ;
	wire _w1256_ ;
	wire _w1257_ ;
	wire _w1258_ ;
	wire _w1259_ ;
	wire _w1260_ ;
	wire _w1261_ ;
	wire _w1262_ ;
	wire _w1263_ ;
	wire _w1264_ ;
	wire _w1265_ ;
	wire _w1266_ ;
	wire _w1267_ ;
	wire _w1268_ ;
	wire _w1269_ ;
	wire _w1270_ ;
	wire _w1271_ ;
	wire _w1272_ ;
	wire _w1273_ ;
	wire _w1274_ ;
	wire _w1275_ ;
	wire _w1276_ ;
	wire _w1277_ ;
	wire _w1278_ ;
	wire _w1279_ ;
	wire _w1280_ ;
	wire _w1281_ ;
	LUT2 #(
		.INIT('h1)
	) name0 (
		\n5_pad ,
		z_pad,
		_w173_
	);
	LUT2 #(
		.INIT('h8)
	) name1 (
		\l5_pad ,
		\m5_pad ,
		_w174_
	);
	LUT2 #(
		.INIT('h8)
	) name2 (
		_w173_,
		_w174_,
		_w175_
	);
	LUT2 #(
		.INIT('h8)
	) name3 (
		\r5_pad ,
		_w175_,
		_w176_
	);
	LUT2 #(
		.INIT('h8)
	) name4 (
		\r4_pad ,
		_w176_,
		_w177_
	);
	LUT2 #(
		.INIT('h2)
	) name5 (
		\l5_pad ,
		\m5_pad ,
		_w178_
	);
	LUT2 #(
		.INIT('h2)
	) name6 (
		\n5_pad ,
		z_pad,
		_w179_
	);
	LUT2 #(
		.INIT('h8)
	) name7 (
		_w178_,
		_w179_,
		_w180_
	);
	LUT2 #(
		.INIT('h1)
	) name8 (
		z_pad,
		_w180_,
		_w181_
	);
	LUT2 #(
		.INIT('h4)
	) name9 (
		\i5_pad ,
		\o5_pad ,
		_w182_
	);
	LUT2 #(
		.INIT('h8)
	) name10 (
		\p10_pad ,
		_w182_,
		_w183_
	);
	LUT2 #(
		.INIT('h1)
	) name11 (
		\d5_pad ,
		\e5_pad ,
		_w184_
	);
	LUT2 #(
		.INIT('h4)
	) name12 (
		\b5_pad ,
		\i10_pad ,
		_w185_
	);
	LUT2 #(
		.INIT('h8)
	) name13 (
		_w184_,
		_w185_,
		_w186_
	);
	LUT2 #(
		.INIT('h4)
	) name14 (
		_w183_,
		_w186_,
		_w187_
	);
	LUT2 #(
		.INIT('h1)
	) name15 (
		\e5_pad ,
		_w187_,
		_w188_
	);
	LUT2 #(
		.INIT('h4)
	) name16 (
		\c5_pad ,
		_w188_,
		_w189_
	);
	LUT2 #(
		.INIT('h2)
	) name17 (
		_w184_,
		_w185_,
		_w190_
	);
	LUT2 #(
		.INIT('h8)
	) name18 (
		_w183_,
		_w190_,
		_w191_
	);
	LUT2 #(
		.INIT('h1)
	) name19 (
		\d5_pad ,
		_w191_,
		_w192_
	);
	LUT2 #(
		.INIT('h8)
	) name20 (
		_w189_,
		_w192_,
		_w193_
	);
	LUT2 #(
		.INIT('h1)
	) name21 (
		\l5_pad ,
		\m5_pad ,
		_w194_
	);
	LUT2 #(
		.INIT('h4)
	) name22 (
		\n5_pad ,
		_w194_,
		_w195_
	);
	LUT2 #(
		.INIT('h8)
	) name23 (
		_w193_,
		_w195_,
		_w196_
	);
	LUT2 #(
		.INIT('h2)
	) name24 (
		_w181_,
		_w196_,
		_w197_
	);
	LUT2 #(
		.INIT('h4)
	) name25 (
		_w177_,
		_w197_,
		_w198_
	);
	LUT2 #(
		.INIT('h4)
	) name26 (
		_w176_,
		_w193_,
		_w199_
	);
	LUT2 #(
		.INIT('h2)
	) name27 (
		\r4_pad ,
		_w199_,
		_w200_
	);
	LUT2 #(
		.INIT('h8)
	) name28 (
		\s4_pad ,
		_w200_,
		_w201_
	);
	LUT2 #(
		.INIT('h8)
	) name29 (
		\t4_pad ,
		_w201_,
		_w202_
	);
	LUT2 #(
		.INIT('h1)
	) name30 (
		\t4_pad ,
		_w201_,
		_w203_
	);
	LUT2 #(
		.INIT('h2)
	) name31 (
		_w198_,
		_w202_,
		_w204_
	);
	LUT2 #(
		.INIT('h4)
	) name32 (
		_w203_,
		_w204_,
		_w205_
	);
	LUT2 #(
		.INIT('h8)
	) name33 (
		\o0_pad ,
		\r5_pad ,
		_w206_
	);
	LUT2 #(
		.INIT('h8)
	) name34 (
		\r4_pad ,
		\u0_pad ,
		_w207_
	);
	LUT2 #(
		.INIT('h8)
	) name35 (
		\t0_pad ,
		\w4_pad ,
		_w208_
	);
	LUT2 #(
		.INIT('h8)
	) name36 (
		\d4_pad ,
		\s0_pad ,
		_w209_
	);
	LUT2 #(
		.INIT('h8)
	) name37 (
		\m5_pad ,
		\p0_pad ,
		_w210_
	);
	LUT2 #(
		.INIT('h8)
	) name38 (
		\h4_pad ,
		\r0_pad ,
		_w211_
	);
	LUT2 #(
		.INIT('h8)
	) name39 (
		\k0_pad ,
		\q3_pad ,
		_w212_
	);
	LUT2 #(
		.INIT('h8)
	) name40 (
		\l0_pad ,
		\m3_pad ,
		_w213_
	);
	LUT2 #(
		.INIT('h8)
	) name41 (
		\n0_pad ,
		\p5_pad ,
		_w214_
	);
	LUT2 #(
		.INIT('h8)
	) name42 (
		\f3_pad ,
		\m0_pad ,
		_w215_
	);
	LUT2 #(
		.INIT('h8)
	) name43 (
		\m4_pad ,
		\q0_pad ,
		_w216_
	);
	LUT2 #(
		.INIT('h1)
	) name44 (
		_w206_,
		_w207_,
		_w217_
	);
	LUT2 #(
		.INIT('h1)
	) name45 (
		_w208_,
		_w209_,
		_w218_
	);
	LUT2 #(
		.INIT('h1)
	) name46 (
		_w210_,
		_w211_,
		_w219_
	);
	LUT2 #(
		.INIT('h1)
	) name47 (
		_w212_,
		_w213_,
		_w220_
	);
	LUT2 #(
		.INIT('h1)
	) name48 (
		_w214_,
		_w215_,
		_w221_
	);
	LUT2 #(
		.INIT('h4)
	) name49 (
		_w216_,
		_w221_,
		_w222_
	);
	LUT2 #(
		.INIT('h8)
	) name50 (
		_w219_,
		_w220_,
		_w223_
	);
	LUT2 #(
		.INIT('h8)
	) name51 (
		_w217_,
		_w218_,
		_w224_
	);
	LUT2 #(
		.INIT('h8)
	) name52 (
		_w223_,
		_w224_,
		_w225_
	);
	LUT2 #(
		.INIT('h8)
	) name53 (
		_w222_,
		_w225_,
		_w226_
	);
	LUT2 #(
		.INIT('h4)
	) name54 (
		b_pad,
		\l1_pad ,
		_w227_
	);
	LUT2 #(
		.INIT('h4)
	) name55 (
		\m1_pad ,
		_w227_,
		_w228_
	);
	LUT2 #(
		.INIT('h4)
	) name56 (
		\n1_pad ,
		_w228_,
		_w229_
	);
	LUT2 #(
		.INIT('h1)
	) name57 (
		\a1_pad ,
		\b1_pad ,
		_w230_
	);
	LUT2 #(
		.INIT('h4)
	) name58 (
		\c1_pad ,
		_w230_,
		_w231_
	);
	LUT2 #(
		.INIT('h1)
	) name59 (
		\x0_pad ,
		\y0_pad ,
		_w232_
	);
	LUT2 #(
		.INIT('h1)
	) name60 (
		\d1_pad ,
		\w0_pad ,
		_w233_
	);
	LUT2 #(
		.INIT('h4)
	) name61 (
		\z0_pad ,
		_w233_,
		_w234_
	);
	LUT2 #(
		.INIT('h8)
	) name62 (
		_w232_,
		_w234_,
		_w235_
	);
	LUT2 #(
		.INIT('h8)
	) name63 (
		_w231_,
		_w235_,
		_w236_
	);
	LUT2 #(
		.INIT('h1)
	) name64 (
		\l1_pad ,
		\m1_pad ,
		_w237_
	);
	LUT2 #(
		.INIT('h4)
	) name65 (
		\n1_pad ,
		_w237_,
		_w238_
	);
	LUT2 #(
		.INIT('h1)
	) name66 (
		b_pad,
		_w238_,
		_w239_
	);
	LUT2 #(
		.INIT('h2)
	) name67 (
		\v0_pad ,
		_w239_,
		_w240_
	);
	LUT2 #(
		.INIT('h8)
	) name68 (
		_w236_,
		_w240_,
		_w241_
	);
	LUT2 #(
		.INIT('h1)
	) name69 (
		_w229_,
		_w241_,
		_w242_
	);
	LUT2 #(
		.INIT('h1)
	) name70 (
		\x2_pad ,
		_w242_,
		_w243_
	);
	LUT2 #(
		.INIT('h4)
	) name71 (
		\k1_pad ,
		\o1_pad ,
		_w244_
	);
	LUT2 #(
		.INIT('h8)
	) name72 (
		\r6_pad ,
		_w244_,
		_w245_
	);
	LUT2 #(
		.INIT('h1)
	) name73 (
		\h1_pad ,
		\i1_pad ,
		_w246_
	);
	LUT2 #(
		.INIT('h4)
	) name74 (
		\f1_pad ,
		\m6_pad ,
		_w247_
	);
	LUT2 #(
		.INIT('h8)
	) name75 (
		_w246_,
		_w247_,
		_w248_
	);
	LUT2 #(
		.INIT('h4)
	) name76 (
		_w245_,
		_w248_,
		_w249_
	);
	LUT2 #(
		.INIT('h1)
	) name77 (
		\i1_pad ,
		_w249_,
		_w250_
	);
	LUT2 #(
		.INIT('h4)
	) name78 (
		\g1_pad ,
		_w250_,
		_w251_
	);
	LUT2 #(
		.INIT('h4)
	) name79 (
		i_pad,
		_w251_,
		_w252_
	);
	LUT2 #(
		.INIT('h8)
	) name80 (
		\s1_pad ,
		_w252_,
		_w253_
	);
	LUT2 #(
		.INIT('h1)
	) name81 (
		\s1_pad ,
		_w252_,
		_w254_
	);
	LUT2 #(
		.INIT('h1)
	) name82 (
		\v0_pad ,
		_w239_,
		_w255_
	);
	LUT2 #(
		.INIT('h8)
	) name83 (
		\r1_pad ,
		_w231_,
		_w256_
	);
	LUT2 #(
		.INIT('h1)
	) name84 (
		\q1_pad ,
		_w256_,
		_w257_
	);
	LUT2 #(
		.INIT('h1)
	) name85 (
		\z0_pad ,
		_w257_,
		_w258_
	);
	LUT2 #(
		.INIT('h1)
	) name86 (
		\p1_pad ,
		_w258_,
		_w259_
	);
	LUT2 #(
		.INIT('h8)
	) name87 (
		\w0_pad ,
		_w232_,
		_w260_
	);
	LUT2 #(
		.INIT('h8)
	) name88 (
		_w255_,
		_w260_,
		_w261_
	);
	LUT2 #(
		.INIT('h4)
	) name89 (
		_w259_,
		_w261_,
		_w262_
	);
	LUT2 #(
		.INIT('h1)
	) name90 (
		h_pad,
		_w262_,
		_w263_
	);
	LUT2 #(
		.INIT('h1)
	) name91 (
		_w254_,
		_w263_,
		_w264_
	);
	LUT2 #(
		.INIT('h4)
	) name92 (
		_w253_,
		_w264_,
		_w265_
	);
	LUT2 #(
		.INIT('h2)
	) name93 (
		\t1_pad ,
		_w265_,
		_w266_
	);
	LUT2 #(
		.INIT('h4)
	) name94 (
		\t1_pad ,
		_w265_,
		_w267_
	);
	LUT2 #(
		.INIT('h2)
	) name95 (
		_w242_,
		_w266_,
		_w268_
	);
	LUT2 #(
		.INIT('h4)
	) name96 (
		_w267_,
		_w268_,
		_w269_
	);
	LUT2 #(
		.INIT('h1)
	) name97 (
		b_pad,
		_w243_,
		_w270_
	);
	LUT2 #(
		.INIT('h4)
	) name98 (
		_w269_,
		_w270_,
		_w271_
	);
	LUT2 #(
		.INIT('h1)
	) name99 (
		_w239_,
		_w251_,
		_w272_
	);
	LUT2 #(
		.INIT('h1)
	) name100 (
		g_pad,
		_w272_,
		_w273_
	);
	LUT2 #(
		.INIT('h4)
	) name101 (
		b_pad,
		\m1_pad ,
		_w274_
	);
	LUT2 #(
		.INIT('h4)
	) name102 (
		\n1_pad ,
		_w274_,
		_w275_
	);
	LUT2 #(
		.INIT('h4)
	) name103 (
		\l1_pad ,
		_w275_,
		_w276_
	);
	LUT2 #(
		.INIT('h1)
	) name104 (
		b_pad,
		_w276_,
		_w277_
	);
	LUT2 #(
		.INIT('h1)
	) name105 (
		_w273_,
		_w277_,
		_w278_
	);
	LUT2 #(
		.INIT('h8)
	) name106 (
		\l1_pad ,
		_w275_,
		_w279_
	);
	LUT2 #(
		.INIT('h4)
	) name107 (
		j_pad,
		\q1_pad ,
		_w280_
	);
	LUT2 #(
		.INIT('h8)
	) name108 (
		_w279_,
		_w280_,
		_w281_
	);
	LUT2 #(
		.INIT('h8)
	) name109 (
		\q2_pad ,
		\r2_pad ,
		_w282_
	);
	LUT2 #(
		.INIT('h1)
	) name110 (
		_w281_,
		_w282_,
		_w283_
	);
	LUT2 #(
		.INIT('h2)
	) name111 (
		\s2_pad ,
		_w283_,
		_w284_
	);
	LUT2 #(
		.INIT('h4)
	) name112 (
		j_pad,
		\p1_pad ,
		_w285_
	);
	LUT2 #(
		.INIT('h8)
	) name113 (
		_w279_,
		_w285_,
		_w286_
	);
	LUT2 #(
		.INIT('h1)
	) name114 (
		_w284_,
		_w286_,
		_w287_
	);
	LUT2 #(
		.INIT('h4)
	) name115 (
		_w273_,
		_w287_,
		_w288_
	);
	LUT2 #(
		.INIT('h1)
	) name116 (
		\q2_pad ,
		\r2_pad ,
		_w289_
	);
	LUT2 #(
		.INIT('h1)
	) name117 (
		_w281_,
		_w289_,
		_w290_
	);
	LUT2 #(
		.INIT('h1)
	) name118 (
		\s2_pad ,
		_w290_,
		_w291_
	);
	LUT2 #(
		.INIT('h1)
	) name119 (
		_w286_,
		_w291_,
		_w292_
	);
	LUT2 #(
		.INIT('h8)
	) name120 (
		_w273_,
		_w292_,
		_w293_
	);
	LUT2 #(
		.INIT('h2)
	) name121 (
		\r1_pad ,
		\v0_pad ,
		_w294_
	);
	LUT2 #(
		.INIT('h2)
	) name122 (
		_w279_,
		_w294_,
		_w295_
	);
	LUT2 #(
		.INIT('h2)
	) name123 (
		_w246_,
		_w247_,
		_w296_
	);
	LUT2 #(
		.INIT('h8)
	) name124 (
		_w245_,
		_w296_,
		_w297_
	);
	LUT2 #(
		.INIT('h1)
	) name125 (
		\h1_pad ,
		_w297_,
		_w298_
	);
	LUT2 #(
		.INIT('h8)
	) name126 (
		_w251_,
		_w298_,
		_w299_
	);
	LUT2 #(
		.INIT('h8)
	) name127 (
		_w236_,
		_w255_,
		_w300_
	);
	LUT2 #(
		.INIT('h4)
	) name128 (
		_w299_,
		_w300_,
		_w301_
	);
	LUT2 #(
		.INIT('h1)
	) name129 (
		f_pad,
		_w295_,
		_w302_
	);
	LUT2 #(
		.INIT('h4)
	) name130 (
		_w301_,
		_w302_,
		_w303_
	);
	LUT2 #(
		.INIT('h1)
	) name131 (
		_w288_,
		_w293_,
		_w304_
	);
	LUT2 #(
		.INIT('h4)
	) name132 (
		_w303_,
		_w304_,
		_w305_
	);
	LUT2 #(
		.INIT('h1)
	) name133 (
		\t2_pad ,
		_w305_,
		_w306_
	);
	LUT2 #(
		.INIT('h8)
	) name134 (
		\t2_pad ,
		_w305_,
		_w307_
	);
	LUT2 #(
		.INIT('h2)
	) name135 (
		_w277_,
		_w306_,
		_w308_
	);
	LUT2 #(
		.INIT('h4)
	) name136 (
		_w307_,
		_w308_,
		_w309_
	);
	LUT2 #(
		.INIT('h1)
	) name137 (
		_w278_,
		_w309_,
		_w310_
	);
	LUT2 #(
		.INIT('h1)
	) name138 (
		z_pad,
		_w195_,
		_w311_
	);
	LUT2 #(
		.INIT('h1)
	) name139 (
		_w189_,
		_w311_,
		_w312_
	);
	LUT2 #(
		.INIT('h1)
	) name140 (
		\e0_pad ,
		_w312_,
		_w313_
	);
	LUT2 #(
		.INIT('h4)
	) name141 (
		\l5_pad ,
		\m5_pad ,
		_w314_
	);
	LUT2 #(
		.INIT('h8)
	) name142 (
		_w173_,
		_w314_,
		_w315_
	);
	LUT2 #(
		.INIT('h1)
	) name143 (
		z_pad,
		_w315_,
		_w316_
	);
	LUT2 #(
		.INIT('h1)
	) name144 (
		_w313_,
		_w316_,
		_w317_
	);
	LUT2 #(
		.INIT('h1)
	) name145 (
		\f3_pad ,
		\g3_pad ,
		_w318_
	);
	LUT2 #(
		.INIT('h4)
	) name146 (
		\h0_pad ,
		\q5_pad ,
		_w319_
	);
	LUT2 #(
		.INIT('h8)
	) name147 (
		_w175_,
		_w319_,
		_w320_
	);
	LUT2 #(
		.INIT('h1)
	) name148 (
		_w318_,
		_w320_,
		_w321_
	);
	LUT2 #(
		.INIT('h1)
	) name149 (
		\h3_pad ,
		_w321_,
		_w322_
	);
	LUT2 #(
		.INIT('h4)
	) name150 (
		\h0_pad ,
		\p5_pad ,
		_w323_
	);
	LUT2 #(
		.INIT('h8)
	) name151 (
		_w175_,
		_w323_,
		_w324_
	);
	LUT2 #(
		.INIT('h1)
	) name152 (
		_w322_,
		_w324_,
		_w325_
	);
	LUT2 #(
		.INIT('h1)
	) name153 (
		\i3_pad ,
		_w325_,
		_w326_
	);
	LUT2 #(
		.INIT('h1)
	) name154 (
		\h0_pad ,
		_w326_,
		_w327_
	);
	LUT2 #(
		.INIT('h2)
	) name155 (
		\j3_pad ,
		_w327_,
		_w328_
	);
	LUT2 #(
		.INIT('h4)
	) name156 (
		\p3_pad ,
		_w328_,
		_w329_
	);
	LUT2 #(
		.INIT('h1)
	) name157 (
		\h0_pad ,
		_w329_,
		_w330_
	);
	LUT2 #(
		.INIT('h1)
	) name158 (
		\q3_pad ,
		_w330_,
		_w331_
	);
	LUT2 #(
		.INIT('h4)
	) name159 (
		\r3_pad ,
		_w331_,
		_w332_
	);
	LUT2 #(
		.INIT('h2)
	) name160 (
		_w313_,
		_w332_,
		_w333_
	);
	LUT2 #(
		.INIT('h8)
	) name161 (
		\q3_pad ,
		\r3_pad ,
		_w334_
	);
	LUT2 #(
		.INIT('h1)
	) name162 (
		_w313_,
		_w334_,
		_w335_
	);
	LUT2 #(
		.INIT('h4)
	) name163 (
		\j5_pad ,
		\k5_pad ,
		_w336_
	);
	LUT2 #(
		.INIT('h4)
	) name164 (
		\r4_pad ,
		\r5_pad ,
		_w337_
	);
	LUT2 #(
		.INIT('h2)
	) name165 (
		_w336_,
		_w337_,
		_w338_
	);
	LUT2 #(
		.INIT('h1)
	) name166 (
		\t4_pad ,
		\u4_pad ,
		_w339_
	);
	LUT2 #(
		.INIT('h1)
	) name167 (
		\v4_pad ,
		\w4_pad ,
		_w340_
	);
	LUT2 #(
		.INIT('h1)
	) name168 (
		\x4_pad ,
		\y4_pad ,
		_w341_
	);
	LUT2 #(
		.INIT('h8)
	) name169 (
		_w340_,
		_w341_,
		_w342_
	);
	LUT2 #(
		.INIT('h8)
	) name170 (
		_w339_,
		_w342_,
		_w343_
	);
	LUT2 #(
		.INIT('h1)
	) name171 (
		\s4_pad ,
		\z4_pad ,
		_w344_
	);
	LUT2 #(
		.INIT('h4)
	) name172 (
		_w311_,
		_w344_,
		_w345_
	);
	LUT2 #(
		.INIT('h8)
	) name173 (
		_w343_,
		_w345_,
		_w346_
	);
	LUT2 #(
		.INIT('h4)
	) name174 (
		\r4_pad ,
		_w346_,
		_w347_
	);
	LUT2 #(
		.INIT('h4)
	) name175 (
		_w193_,
		_w347_,
		_w348_
	);
	LUT2 #(
		.INIT('h1)
	) name176 (
		\d0_pad ,
		_w338_,
		_w349_
	);
	LUT2 #(
		.INIT('h4)
	) name177 (
		_w348_,
		_w349_,
		_w350_
	);
	LUT2 #(
		.INIT('h8)
	) name178 (
		\f3_pad ,
		\g3_pad ,
		_w351_
	);
	LUT2 #(
		.INIT('h1)
	) name179 (
		_w320_,
		_w351_,
		_w352_
	);
	LUT2 #(
		.INIT('h2)
	) name180 (
		\h3_pad ,
		_w352_,
		_w353_
	);
	LUT2 #(
		.INIT('h1)
	) name181 (
		_w324_,
		_w353_,
		_w354_
	);
	LUT2 #(
		.INIT('h2)
	) name182 (
		\i3_pad ,
		_w354_,
		_w355_
	);
	LUT2 #(
		.INIT('h1)
	) name183 (
		\h0_pad ,
		_w355_,
		_w356_
	);
	LUT2 #(
		.INIT('h2)
	) name184 (
		\k3_pad ,
		_w356_,
		_w357_
	);
	LUT2 #(
		.INIT('h8)
	) name185 (
		\p3_pad ,
		_w357_,
		_w358_
	);
	LUT2 #(
		.INIT('h1)
	) name186 (
		\h0_pad ,
		_w313_,
		_w359_
	);
	LUT2 #(
		.INIT('h4)
	) name187 (
		_w358_,
		_w359_,
		_w360_
	);
	LUT2 #(
		.INIT('h1)
	) name188 (
		_w350_,
		_w360_,
		_w361_
	);
	LUT2 #(
		.INIT('h4)
	) name189 (
		_w335_,
		_w361_,
		_w362_
	);
	LUT2 #(
		.INIT('h4)
	) name190 (
		_w333_,
		_w362_,
		_w363_
	);
	LUT2 #(
		.INIT('h1)
	) name191 (
		\s3_pad ,
		_w313_,
		_w364_
	);
	LUT2 #(
		.INIT('h8)
	) name192 (
		\s3_pad ,
		_w313_,
		_w365_
	);
	LUT2 #(
		.INIT('h1)
	) name193 (
		_w364_,
		_w365_,
		_w366_
	);
	LUT2 #(
		.INIT('h8)
	) name194 (
		_w363_,
		_w366_,
		_w367_
	);
	LUT2 #(
		.INIT('h1)
	) name195 (
		\t3_pad ,
		_w367_,
		_w368_
	);
	LUT2 #(
		.INIT('h8)
	) name196 (
		\t3_pad ,
		_w367_,
		_w369_
	);
	LUT2 #(
		.INIT('h2)
	) name197 (
		_w316_,
		_w368_,
		_w370_
	);
	LUT2 #(
		.INIT('h4)
	) name198 (
		_w369_,
		_w370_,
		_w371_
	);
	LUT2 #(
		.INIT('h1)
	) name199 (
		_w317_,
		_w371_,
		_w372_
	);
	LUT2 #(
		.INIT('h8)
	) name200 (
		\u4_pad ,
		_w202_,
		_w373_
	);
	LUT2 #(
		.INIT('h1)
	) name201 (
		\u4_pad ,
		_w202_,
		_w374_
	);
	LUT2 #(
		.INIT('h2)
	) name202 (
		_w198_,
		_w373_,
		_w375_
	);
	LUT2 #(
		.INIT('h4)
	) name203 (
		_w374_,
		_w375_,
		_w376_
	);
	LUT2 #(
		.INIT('h8)
	) name204 (
		\n5_pad ,
		\p0_pad ,
		_w377_
	);
	LUT2 #(
		.INIT('h8)
	) name205 (
		\l0_pad ,
		\l3_pad ,
		_w378_
	);
	LUT2 #(
		.INIT('h8)
	) name206 (
		\g4_pad ,
		\r0_pad ,
		_w379_
	);
	LUT2 #(
		.INIT('h8)
	) name207 (
		\p3_pad ,
		\s3_pad ,
		_w380_
	);
	LUT2 #(
		.INIT('h8)
	) name208 (
		\t3_pad ,
		_w380_,
		_w381_
	);
	LUT2 #(
		.INIT('h8)
	) name209 (
		_w334_,
		_w381_,
		_w382_
	);
	LUT2 #(
		.INIT('h8)
	) name210 (
		\m0_pad ,
		_w382_,
		_w383_
	);
	LUT2 #(
		.INIT('h2)
	) name211 (
		\n3_pad ,
		\o3_pad ,
		_w384_
	);
	LUT2 #(
		.INIT('h1)
	) name212 (
		\p3_pad ,
		\q3_pad ,
		_w385_
	);
	LUT2 #(
		.INIT('h1)
	) name213 (
		\r3_pad ,
		\s3_pad ,
		_w386_
	);
	LUT2 #(
		.INIT('h4)
	) name214 (
		\t3_pad ,
		_w386_,
		_w387_
	);
	LUT2 #(
		.INIT('h8)
	) name215 (
		_w384_,
		_w385_,
		_w388_
	);
	LUT2 #(
		.INIT('h8)
	) name216 (
		_w387_,
		_w388_,
		_w389_
	);
	LUT2 #(
		.INIT('h8)
	) name217 (
		\k0_pad ,
		_w389_,
		_w390_
	);
	LUT2 #(
		.INIT('h8)
	) name218 (
		\l5_pad ,
		\u0_pad ,
		_w391_
	);
	LUT2 #(
		.INIT('h2)
	) name219 (
		\o0_pad ,
		_w316_,
		_w392_
	);
	LUT2 #(
		.INIT('h8)
	) name220 (
		\s0_pad ,
		_w350_,
		_w393_
	);
	LUT2 #(
		.INIT('h4)
	) name221 (
		\j0_pad ,
		\q5_pad ,
		_w394_
	);
	LUT2 #(
		.INIT('h8)
	) name222 (
		\d4_pad ,
		\e4_pad ,
		_w395_
	);
	LUT2 #(
		.INIT('h8)
	) name223 (
		\f4_pad ,
		_w395_,
		_w396_
	);
	LUT2 #(
		.INIT('h1)
	) name224 (
		_w394_,
		_w396_,
		_w397_
	);
	LUT2 #(
		.INIT('h2)
	) name225 (
		\i4_pad ,
		_w397_,
		_w398_
	);
	LUT2 #(
		.INIT('h1)
	) name226 (
		\j0_pad ,
		\p5_pad ,
		_w399_
	);
	LUT2 #(
		.INIT('h4)
	) name227 (
		_w398_,
		_w399_,
		_w400_
	);
	LUT2 #(
		.INIT('h2)
	) name228 (
		\g4_pad ,
		_w400_,
		_w401_
	);
	LUT2 #(
		.INIT('h8)
	) name229 (
		\p4_pad ,
		_w401_,
		_w402_
	);
	LUT2 #(
		.INIT('h8)
	) name230 (
		\q0_pad ,
		_w402_,
		_w403_
	);
	LUT2 #(
		.INIT('h8)
	) name231 (
		\t0_pad ,
		\v4_pad ,
		_w404_
	);
	LUT2 #(
		.INIT('h8)
	) name232 (
		\n0_pad ,
		\q5_pad ,
		_w405_
	);
	LUT2 #(
		.INIT('h1)
	) name233 (
		_w377_,
		_w378_,
		_w406_
	);
	LUT2 #(
		.INIT('h1)
	) name234 (
		_w379_,
		_w391_,
		_w407_
	);
	LUT2 #(
		.INIT('h1)
	) name235 (
		_w404_,
		_w405_,
		_w408_
	);
	LUT2 #(
		.INIT('h8)
	) name236 (
		_w407_,
		_w408_,
		_w409_
	);
	LUT2 #(
		.INIT('h8)
	) name237 (
		_w406_,
		_w409_,
		_w410_
	);
	LUT2 #(
		.INIT('h4)
	) name238 (
		_w383_,
		_w410_,
		_w411_
	);
	LUT2 #(
		.INIT('h1)
	) name239 (
		_w390_,
		_w392_,
		_w412_
	);
	LUT2 #(
		.INIT('h8)
	) name240 (
		_w411_,
		_w412_,
		_w413_
	);
	LUT2 #(
		.INIT('h4)
	) name241 (
		_w403_,
		_w413_,
		_w414_
	);
	LUT2 #(
		.INIT('h4)
	) name242 (
		_w393_,
		_w414_,
		_w415_
	);
	LUT2 #(
		.INIT('h1)
	) name243 (
		\y2_pad ,
		_w242_,
		_w416_
	);
	LUT2 #(
		.INIT('h1)
	) name244 (
		\s1_pad ,
		\t1_pad ,
		_w417_
	);
	LUT2 #(
		.INIT('h2)
	) name245 (
		\t1_pad ,
		_w252_,
		_w418_
	);
	LUT2 #(
		.INIT('h1)
	) name246 (
		_w417_,
		_w418_,
		_w419_
	);
	LUT2 #(
		.INIT('h2)
	) name247 (
		_w264_,
		_w419_,
		_w420_
	);
	LUT2 #(
		.INIT('h2)
	) name248 (
		\u1_pad ,
		_w420_,
		_w421_
	);
	LUT2 #(
		.INIT('h4)
	) name249 (
		\u1_pad ,
		_w420_,
		_w422_
	);
	LUT2 #(
		.INIT('h2)
	) name250 (
		_w242_,
		_w421_,
		_w423_
	);
	LUT2 #(
		.INIT('h4)
	) name251 (
		_w422_,
		_w423_,
		_w424_
	);
	LUT2 #(
		.INIT('h1)
	) name252 (
		b_pad,
		_w416_,
		_w425_
	);
	LUT2 #(
		.INIT('h4)
	) name253 (
		_w424_,
		_w425_,
		_w426_
	);
	LUT2 #(
		.INIT('h1)
	) name254 (
		\w2_pad ,
		\x2_pad ,
		_w427_
	);
	LUT2 #(
		.INIT('h1)
	) name255 (
		\y2_pad ,
		\z2_pad ,
		_w428_
	);
	LUT2 #(
		.INIT('h8)
	) name256 (
		_w427_,
		_w428_,
		_w429_
	);
	LUT2 #(
		.INIT('h2)
	) name257 (
		_w277_,
		_w429_,
		_w430_
	);
	LUT2 #(
		.INIT('h1)
	) name258 (
		_w278_,
		_w430_,
		_w431_
	);
	LUT2 #(
		.INIT('h8)
	) name259 (
		\r4_pad ,
		_w346_,
		_w432_
	);
	LUT2 #(
		.INIT('h8)
	) name260 (
		_w173_,
		_w178_,
		_w433_
	);
	LUT2 #(
		.INIT('h1)
	) name261 (
		_w432_,
		_w433_,
		_w434_
	);
	LUT2 #(
		.INIT('h1)
	) name262 (
		\l3_pad ,
		_w434_,
		_w435_
	);
	LUT2 #(
		.INIT('h2)
	) name263 (
		\q5_pad ,
		\v4_pad ,
		_w436_
	);
	LUT2 #(
		.INIT('h8)
	) name264 (
		\r5_pad ,
		_w343_,
		_w437_
	);
	LUT2 #(
		.INIT('h1)
	) name265 (
		\p5_pad ,
		_w436_,
		_w438_
	);
	LUT2 #(
		.INIT('h4)
	) name266 (
		_w437_,
		_w438_,
		_w439_
	);
	LUT2 #(
		.INIT('h4)
	) name267 (
		\r4_pad ,
		\s4_pad ,
		_w440_
	);
	LUT2 #(
		.INIT('h8)
	) name268 (
		_w339_,
		_w440_,
		_w441_
	);
	LUT2 #(
		.INIT('h4)
	) name269 (
		_w311_,
		_w441_,
		_w442_
	);
	LUT2 #(
		.INIT('h4)
	) name270 (
		_w439_,
		_w442_,
		_w443_
	);
	LUT2 #(
		.INIT('h1)
	) name271 (
		\f0_pad ,
		_w443_,
		_w444_
	);
	LUT2 #(
		.INIT('h2)
	) name272 (
		\u3_pad ,
		_w444_,
		_w445_
	);
	LUT2 #(
		.INIT('h4)
	) name273 (
		\u3_pad ,
		_w444_,
		_w446_
	);
	LUT2 #(
		.INIT('h1)
	) name274 (
		_w445_,
		_w446_,
		_w447_
	);
	LUT2 #(
		.INIT('h2)
	) name275 (
		_w434_,
		_w447_,
		_w448_
	);
	LUT2 #(
		.INIT('h1)
	) name276 (
		z_pad,
		_w435_,
		_w449_
	);
	LUT2 #(
		.INIT('h4)
	) name277 (
		_w448_,
		_w449_,
		_w450_
	);
	LUT2 #(
		.INIT('h1)
	) name278 (
		\v4_pad ,
		_w373_,
		_w451_
	);
	LUT2 #(
		.INIT('h8)
	) name279 (
		\v4_pad ,
		_w373_,
		_w452_
	);
	LUT2 #(
		.INIT('h2)
	) name280 (
		_w198_,
		_w451_,
		_w453_
	);
	LUT2 #(
		.INIT('h4)
	) name281 (
		_w452_,
		_w453_,
		_w454_
	);
	LUT2 #(
		.INIT('h8)
	) name282 (
		_w179_,
		_w194_,
		_w455_
	);
	LUT2 #(
		.INIT('h8)
	) name283 (
		_w175_,
		_w389_,
		_w456_
	);
	LUT2 #(
		.INIT('h1)
	) name284 (
		_w455_,
		_w456_,
		_w457_
	);
	LUT2 #(
		.INIT('h8)
	) name285 (
		_w175_,
		_w185_,
		_w458_
	);
	LUT2 #(
		.INIT('h8)
	) name286 (
		_w382_,
		_w458_,
		_w459_
	);
	LUT2 #(
		.INIT('h8)
	) name287 (
		_w174_,
		_w179_,
		_w460_
	);
	LUT2 #(
		.INIT('h1)
	) name288 (
		_w433_,
		_w460_,
		_w461_
	);
	LUT2 #(
		.INIT('h4)
	) name289 (
		_w459_,
		_w461_,
		_w462_
	);
	LUT2 #(
		.INIT('h8)
	) name290 (
		_w457_,
		_w462_,
		_w463_
	);
	LUT2 #(
		.INIT('h8)
	) name291 (
		\n1_pad ,
		_w228_,
		_w464_
	);
	LUT2 #(
		.INIT('h1)
	) name292 (
		b_pad,
		_w464_,
		_w465_
	);
	LUT2 #(
		.INIT('h8)
	) name293 (
		_w238_,
		_w299_,
		_w466_
	);
	LUT2 #(
		.INIT('h2)
	) name294 (
		_w465_,
		_w466_,
		_w467_
	);
	LUT2 #(
		.INIT('h8)
	) name295 (
		\r1_pad ,
		_w279_,
		_w468_
	);
	LUT2 #(
		.INIT('h2)
	) name296 (
		_w299_,
		_w468_,
		_w469_
	);
	LUT2 #(
		.INIT('h2)
	) name297 (
		\v0_pad ,
		_w469_,
		_w470_
	);
	LUT2 #(
		.INIT('h4)
	) name298 (
		\v0_pad ,
		_w469_,
		_w471_
	);
	LUT2 #(
		.INIT('h2)
	) name299 (
		_w467_,
		_w470_,
		_w472_
	);
	LUT2 #(
		.INIT('h4)
	) name300 (
		_w471_,
		_w472_,
		_w473_
	);
	LUT2 #(
		.INIT('h2)
	) name301 (
		\z2_pad ,
		_w242_,
		_w474_
	);
	LUT2 #(
		.INIT('h8)
	) name302 (
		\s1_pad ,
		\t1_pad ,
		_w475_
	);
	LUT2 #(
		.INIT('h8)
	) name303 (
		\u1_pad ,
		_w475_,
		_w476_
	);
	LUT2 #(
		.INIT('h1)
	) name304 (
		k_pad,
		_w476_,
		_w477_
	);
	LUT2 #(
		.INIT('h4)
	) name305 (
		_w252_,
		_w477_,
		_w478_
	);
	LUT2 #(
		.INIT('h4)
	) name306 (
		\u1_pad ,
		_w417_,
		_w479_
	);
	LUT2 #(
		.INIT('h1)
	) name307 (
		k_pad,
		_w479_,
		_w480_
	);
	LUT2 #(
		.INIT('h8)
	) name308 (
		_w252_,
		_w480_,
		_w481_
	);
	LUT2 #(
		.INIT('h1)
	) name309 (
		_w478_,
		_w481_,
		_w482_
	);
	LUT2 #(
		.INIT('h4)
	) name310 (
		_w263_,
		_w482_,
		_w483_
	);
	LUT2 #(
		.INIT('h1)
	) name311 (
		\v1_pad ,
		_w483_,
		_w484_
	);
	LUT2 #(
		.INIT('h8)
	) name312 (
		\v1_pad ,
		_w483_,
		_w485_
	);
	LUT2 #(
		.INIT('h2)
	) name313 (
		_w242_,
		_w484_,
		_w486_
	);
	LUT2 #(
		.INIT('h4)
	) name314 (
		_w485_,
		_w486_,
		_w487_
	);
	LUT2 #(
		.INIT('h1)
	) name315 (
		b_pad,
		_w474_,
		_w488_
	);
	LUT2 #(
		.INIT('h4)
	) name316 (
		_w487_,
		_w488_,
		_w489_
	);
	LUT2 #(
		.INIT('h8)
	) name317 (
		\w2_pad ,
		\x2_pad ,
		_w490_
	);
	LUT2 #(
		.INIT('h8)
	) name318 (
		\y2_pad ,
		\z2_pad ,
		_w491_
	);
	LUT2 #(
		.INIT('h8)
	) name319 (
		_w490_,
		_w491_,
		_w492_
	);
	LUT2 #(
		.INIT('h8)
	) name320 (
		_w277_,
		_w492_,
		_w493_
	);
	LUT2 #(
		.INIT('h1)
	) name321 (
		\m3_pad ,
		_w434_,
		_w494_
	);
	LUT2 #(
		.INIT('h4)
	) name322 (
		\g0_pad ,
		_w189_,
		_w495_
	);
	LUT2 #(
		.INIT('h8)
	) name323 (
		\u3_pad ,
		_w495_,
		_w496_
	);
	LUT2 #(
		.INIT('h1)
	) name324 (
		\u3_pad ,
		_w495_,
		_w497_
	);
	LUT2 #(
		.INIT('h1)
	) name325 (
		_w444_,
		_w497_,
		_w498_
	);
	LUT2 #(
		.INIT('h4)
	) name326 (
		_w496_,
		_w498_,
		_w499_
	);
	LUT2 #(
		.INIT('h2)
	) name327 (
		\v3_pad ,
		_w499_,
		_w500_
	);
	LUT2 #(
		.INIT('h4)
	) name328 (
		\v3_pad ,
		_w499_,
		_w501_
	);
	LUT2 #(
		.INIT('h2)
	) name329 (
		_w434_,
		_w500_,
		_w502_
	);
	LUT2 #(
		.INIT('h4)
	) name330 (
		_w501_,
		_w502_,
		_w503_
	);
	LUT2 #(
		.INIT('h1)
	) name331 (
		z_pad,
		_w494_,
		_w504_
	);
	LUT2 #(
		.INIT('h4)
	) name332 (
		_w503_,
		_w504_,
		_w505_
	);
	LUT2 #(
		.INIT('h1)
	) name333 (
		\w4_pad ,
		_w452_,
		_w506_
	);
	LUT2 #(
		.INIT('h8)
	) name334 (
		\w4_pad ,
		_w452_,
		_w507_
	);
	LUT2 #(
		.INIT('h2)
	) name335 (
		_w198_,
		_w506_,
		_w508_
	);
	LUT2 #(
		.INIT('h4)
	) name336 (
		_w507_,
		_w508_,
		_w509_
	);
	LUT2 #(
		.INIT('h8)
	) name337 (
		\v0_pad ,
		_w468_,
		_w510_
	);
	LUT2 #(
		.INIT('h2)
	) name338 (
		_w467_,
		_w510_,
		_w511_
	);
	LUT2 #(
		.INIT('h1)
	) name339 (
		\w0_pad ,
		_w470_,
		_w512_
	);
	LUT2 #(
		.INIT('h8)
	) name340 (
		\w0_pad ,
		_w470_,
		_w513_
	);
	LUT2 #(
		.INIT('h2)
	) name341 (
		_w511_,
		_w512_,
		_w514_
	);
	LUT2 #(
		.INIT('h4)
	) name342 (
		_w513_,
		_w514_,
		_w515_
	);
	LUT2 #(
		.INIT('h2)
	) name343 (
		\a3_pad ,
		_w242_,
		_w516_
	);
	LUT2 #(
		.INIT('h1)
	) name344 (
		\v1_pad ,
		_w480_,
		_w517_
	);
	LUT2 #(
		.INIT('h2)
	) name345 (
		_w252_,
		_w517_,
		_w518_
	);
	LUT2 #(
		.INIT('h2)
	) name346 (
		\v1_pad ,
		_w477_,
		_w519_
	);
	LUT2 #(
		.INIT('h1)
	) name347 (
		_w252_,
		_w519_,
		_w520_
	);
	LUT2 #(
		.INIT('h1)
	) name348 (
		_w518_,
		_w520_,
		_w521_
	);
	LUT2 #(
		.INIT('h4)
	) name349 (
		_w263_,
		_w521_,
		_w522_
	);
	LUT2 #(
		.INIT('h1)
	) name350 (
		\w1_pad ,
		_w522_,
		_w523_
	);
	LUT2 #(
		.INIT('h8)
	) name351 (
		\w1_pad ,
		_w522_,
		_w524_
	);
	LUT2 #(
		.INIT('h2)
	) name352 (
		_w242_,
		_w523_,
		_w525_
	);
	LUT2 #(
		.INIT('h4)
	) name353 (
		_w524_,
		_w525_,
		_w526_
	);
	LUT2 #(
		.INIT('h1)
	) name354 (
		b_pad,
		_w516_,
		_w527_
	);
	LUT2 #(
		.INIT('h4)
	) name355 (
		_w526_,
		_w527_,
		_w528_
	);
	LUT2 #(
		.INIT('h1)
	) name356 (
		\t2_pad ,
		_w292_,
		_w529_
	);
	LUT2 #(
		.INIT('h1)
	) name357 (
		j_pad,
		_w529_,
		_w530_
	);
	LUT2 #(
		.INIT('h2)
	) name358 (
		_w273_,
		_w530_,
		_w531_
	);
	LUT2 #(
		.INIT('h2)
	) name359 (
		\t2_pad ,
		_w287_,
		_w532_
	);
	LUT2 #(
		.INIT('h1)
	) name360 (
		j_pad,
		_w532_,
		_w533_
	);
	LUT2 #(
		.INIT('h1)
	) name361 (
		_w273_,
		_w533_,
		_w534_
	);
	LUT2 #(
		.INIT('h1)
	) name362 (
		_w531_,
		_w534_,
		_w535_
	);
	LUT2 #(
		.INIT('h1)
	) name363 (
		_w303_,
		_w535_,
		_w536_
	);
	LUT2 #(
		.INIT('h8)
	) name364 (
		\w2_pad ,
		_w536_,
		_w537_
	);
	LUT2 #(
		.INIT('h1)
	) name365 (
		\w2_pad ,
		_w536_,
		_w538_
	);
	LUT2 #(
		.INIT('h2)
	) name366 (
		_w277_,
		_w537_,
		_w539_
	);
	LUT2 #(
		.INIT('h4)
	) name367 (
		_w538_,
		_w539_,
		_w540_
	);
	LUT2 #(
		.INIT('h1)
	) name368 (
		\n3_pad ,
		_w434_,
		_w541_
	);
	LUT2 #(
		.INIT('h1)
	) name369 (
		\u3_pad ,
		\v3_pad ,
		_w542_
	);
	LUT2 #(
		.INIT('h2)
	) name370 (
		\v3_pad ,
		_w495_,
		_w543_
	);
	LUT2 #(
		.INIT('h1)
	) name371 (
		_w542_,
		_w543_,
		_w544_
	);
	LUT2 #(
		.INIT('h2)
	) name372 (
		_w498_,
		_w544_,
		_w545_
	);
	LUT2 #(
		.INIT('h2)
	) name373 (
		\w3_pad ,
		_w545_,
		_w546_
	);
	LUT2 #(
		.INIT('h4)
	) name374 (
		\w3_pad ,
		_w545_,
		_w547_
	);
	LUT2 #(
		.INIT('h2)
	) name375 (
		_w434_,
		_w546_,
		_w548_
	);
	LUT2 #(
		.INIT('h4)
	) name376 (
		_w547_,
		_w548_,
		_w549_
	);
	LUT2 #(
		.INIT('h1)
	) name377 (
		z_pad,
		_w541_,
		_w550_
	);
	LUT2 #(
		.INIT('h4)
	) name378 (
		_w549_,
		_w550_,
		_w551_
	);
	LUT2 #(
		.INIT('h8)
	) name379 (
		\w4_pad ,
		\x4_pad ,
		_w552_
	);
	LUT2 #(
		.INIT('h8)
	) name380 (
		_w452_,
		_w552_,
		_w553_
	);
	LUT2 #(
		.INIT('h1)
	) name381 (
		\x4_pad ,
		_w507_,
		_w554_
	);
	LUT2 #(
		.INIT('h2)
	) name382 (
		_w198_,
		_w553_,
		_w555_
	);
	LUT2 #(
		.INIT('h4)
	) name383 (
		_w554_,
		_w555_,
		_w556_
	);
	LUT2 #(
		.INIT('h1)
	) name384 (
		\x0_pad ,
		_w513_,
		_w557_
	);
	LUT2 #(
		.INIT('h8)
	) name385 (
		\x0_pad ,
		_w513_,
		_w558_
	);
	LUT2 #(
		.INIT('h2)
	) name386 (
		_w511_,
		_w557_,
		_w559_
	);
	LUT2 #(
		.INIT('h4)
	) name387 (
		_w558_,
		_w559_,
		_w560_
	);
	LUT2 #(
		.INIT('h2)
	) name388 (
		\b3_pad ,
		_w242_,
		_w561_
	);
	LUT2 #(
		.INIT('h4)
	) name389 (
		\w1_pad ,
		_w517_,
		_w562_
	);
	LUT2 #(
		.INIT('h2)
	) name390 (
		_w252_,
		_w562_,
		_w563_
	);
	LUT2 #(
		.INIT('h8)
	) name391 (
		\w1_pad ,
		_w519_,
		_w564_
	);
	LUT2 #(
		.INIT('h1)
	) name392 (
		_w252_,
		_w564_,
		_w565_
	);
	LUT2 #(
		.INIT('h1)
	) name393 (
		_w563_,
		_w565_,
		_w566_
	);
	LUT2 #(
		.INIT('h4)
	) name394 (
		_w263_,
		_w566_,
		_w567_
	);
	LUT2 #(
		.INIT('h1)
	) name395 (
		\x1_pad ,
		_w567_,
		_w568_
	);
	LUT2 #(
		.INIT('h8)
	) name396 (
		\x1_pad ,
		_w567_,
		_w569_
	);
	LUT2 #(
		.INIT('h2)
	) name397 (
		_w242_,
		_w568_,
		_w570_
	);
	LUT2 #(
		.INIT('h4)
	) name398 (
		_w569_,
		_w570_,
		_w571_
	);
	LUT2 #(
		.INIT('h1)
	) name399 (
		b_pad,
		_w561_,
		_w572_
	);
	LUT2 #(
		.INIT('h4)
	) name400 (
		_w571_,
		_w572_,
		_w573_
	);
	LUT2 #(
		.INIT('h2)
	) name401 (
		\w2_pad ,
		_w534_,
		_w574_
	);
	LUT2 #(
		.INIT('h1)
	) name402 (
		\w2_pad ,
		_w531_,
		_w575_
	);
	LUT2 #(
		.INIT('h1)
	) name403 (
		_w303_,
		_w574_,
		_w576_
	);
	LUT2 #(
		.INIT('h4)
	) name404 (
		_w575_,
		_w576_,
		_w577_
	);
	LUT2 #(
		.INIT('h8)
	) name405 (
		\x2_pad ,
		_w577_,
		_w578_
	);
	LUT2 #(
		.INIT('h1)
	) name406 (
		\x2_pad ,
		_w577_,
		_w579_
	);
	LUT2 #(
		.INIT('h2)
	) name407 (
		_w277_,
		_w578_,
		_w580_
	);
	LUT2 #(
		.INIT('h4)
	) name408 (
		_w579_,
		_w580_,
		_w581_
	);
	LUT2 #(
		.INIT('h2)
	) name409 (
		\o3_pad ,
		_w434_,
		_w582_
	);
	LUT2 #(
		.INIT('h4)
	) name410 (
		\w3_pad ,
		_w542_,
		_w583_
	);
	LUT2 #(
		.INIT('h4)
	) name411 (
		\i0_pad ,
		_w495_,
		_w584_
	);
	LUT2 #(
		.INIT('h4)
	) name412 (
		_w583_,
		_w584_,
		_w585_
	);
	LUT2 #(
		.INIT('h8)
	) name413 (
		\u3_pad ,
		\v3_pad ,
		_w586_
	);
	LUT2 #(
		.INIT('h8)
	) name414 (
		\w3_pad ,
		_w586_,
		_w587_
	);
	LUT2 #(
		.INIT('h1)
	) name415 (
		\i0_pad ,
		_w587_,
		_w588_
	);
	LUT2 #(
		.INIT('h4)
	) name416 (
		_w495_,
		_w588_,
		_w589_
	);
	LUT2 #(
		.INIT('h1)
	) name417 (
		_w444_,
		_w589_,
		_w590_
	);
	LUT2 #(
		.INIT('h4)
	) name418 (
		_w585_,
		_w590_,
		_w591_
	);
	LUT2 #(
		.INIT('h1)
	) name419 (
		\x3_pad ,
		_w591_,
		_w592_
	);
	LUT2 #(
		.INIT('h8)
	) name420 (
		\x3_pad ,
		_w591_,
		_w593_
	);
	LUT2 #(
		.INIT('h2)
	) name421 (
		_w434_,
		_w592_,
		_w594_
	);
	LUT2 #(
		.INIT('h4)
	) name422 (
		_w593_,
		_w594_,
		_w595_
	);
	LUT2 #(
		.INIT('h1)
	) name423 (
		z_pad,
		_w582_,
		_w596_
	);
	LUT2 #(
		.INIT('h4)
	) name424 (
		_w595_,
		_w596_,
		_w597_
	);
	LUT2 #(
		.INIT('h1)
	) name425 (
		\y4_pad ,
		_w553_,
		_w598_
	);
	LUT2 #(
		.INIT('h8)
	) name426 (
		\y4_pad ,
		_w553_,
		_w599_
	);
	LUT2 #(
		.INIT('h2)
	) name427 (
		_w198_,
		_w598_,
		_w600_
	);
	LUT2 #(
		.INIT('h4)
	) name428 (
		_w599_,
		_w600_,
		_w601_
	);
	LUT2 #(
		.INIT('h8)
	) name429 (
		_w247_,
		_w276_,
		_w602_
	);
	LUT2 #(
		.INIT('h8)
	) name430 (
		\c3_pad ,
		\d3_pad ,
		_w603_
	);
	LUT2 #(
		.INIT('h8)
	) name431 (
		\e3_pad ,
		_w603_,
		_w604_
	);
	LUT2 #(
		.INIT('h8)
	) name432 (
		_w247_,
		_w604_,
		_w605_
	);
	LUT2 #(
		.INIT('h2)
	) name433 (
		_w279_,
		_w605_,
		_w606_
	);
	LUT2 #(
		.INIT('h1)
	) name434 (
		_w229_,
		_w602_,
		_w607_
	);
	LUT2 #(
		.INIT('h4)
	) name435 (
		_w606_,
		_w607_,
		_w608_
	);
	LUT2 #(
		.INIT('h1)
	) name436 (
		\y0_pad ,
		_w558_,
		_w609_
	);
	LUT2 #(
		.INIT('h8)
	) name437 (
		\y0_pad ,
		_w558_,
		_w610_
	);
	LUT2 #(
		.INIT('h2)
	) name438 (
		_w511_,
		_w609_,
		_w611_
	);
	LUT2 #(
		.INIT('h4)
	) name439 (
		_w610_,
		_w611_,
		_w612_
	);
	LUT2 #(
		.INIT('h1)
	) name440 (
		\c3_pad ,
		_w242_,
		_w613_
	);
	LUT2 #(
		.INIT('h4)
	) name441 (
		\x1_pad ,
		_w562_,
		_w614_
	);
	LUT2 #(
		.INIT('h1)
	) name442 (
		k_pad,
		_w614_,
		_w615_
	);
	LUT2 #(
		.INIT('h8)
	) name443 (
		_w252_,
		_w615_,
		_w616_
	);
	LUT2 #(
		.INIT('h8)
	) name444 (
		\x1_pad ,
		_w564_,
		_w617_
	);
	LUT2 #(
		.INIT('h1)
	) name445 (
		k_pad,
		_w617_,
		_w618_
	);
	LUT2 #(
		.INIT('h4)
	) name446 (
		_w252_,
		_w618_,
		_w619_
	);
	LUT2 #(
		.INIT('h1)
	) name447 (
		_w263_,
		_w616_,
		_w620_
	);
	LUT2 #(
		.INIT('h4)
	) name448 (
		_w619_,
		_w620_,
		_w621_
	);
	LUT2 #(
		.INIT('h2)
	) name449 (
		\y1_pad ,
		_w621_,
		_w622_
	);
	LUT2 #(
		.INIT('h4)
	) name450 (
		\y1_pad ,
		_w621_,
		_w623_
	);
	LUT2 #(
		.INIT('h2)
	) name451 (
		_w242_,
		_w622_,
		_w624_
	);
	LUT2 #(
		.INIT('h4)
	) name452 (
		_w623_,
		_w624_,
		_w625_
	);
	LUT2 #(
		.INIT('h1)
	) name453 (
		b_pad,
		_w613_,
		_w626_
	);
	LUT2 #(
		.INIT('h4)
	) name454 (
		_w625_,
		_w626_,
		_w627_
	);
	LUT2 #(
		.INIT('h8)
	) name455 (
		_w427_,
		_w531_,
		_w628_
	);
	LUT2 #(
		.INIT('h8)
	) name456 (
		_w490_,
		_w534_,
		_w629_
	);
	LUT2 #(
		.INIT('h1)
	) name457 (
		_w628_,
		_w629_,
		_w630_
	);
	LUT2 #(
		.INIT('h1)
	) name458 (
		_w303_,
		_w630_,
		_w631_
	);
	LUT2 #(
		.INIT('h8)
	) name459 (
		\y2_pad ,
		_w631_,
		_w632_
	);
	LUT2 #(
		.INIT('h1)
	) name460 (
		\y2_pad ,
		_w631_,
		_w633_
	);
	LUT2 #(
		.INIT('h2)
	) name461 (
		_w277_,
		_w632_,
		_w634_
	);
	LUT2 #(
		.INIT('h4)
	) name462 (
		_w633_,
		_w634_,
		_w635_
	);
	LUT2 #(
		.INIT('h2)
	) name463 (
		\p3_pad ,
		_w434_,
		_w636_
	);
	LUT2 #(
		.INIT('h1)
	) name464 (
		\i0_pad ,
		_w583_,
		_w637_
	);
	LUT2 #(
		.INIT('h1)
	) name465 (
		\x3_pad ,
		_w637_,
		_w638_
	);
	LUT2 #(
		.INIT('h2)
	) name466 (
		_w495_,
		_w638_,
		_w639_
	);
	LUT2 #(
		.INIT('h2)
	) name467 (
		\x3_pad ,
		_w588_,
		_w640_
	);
	LUT2 #(
		.INIT('h1)
	) name468 (
		_w495_,
		_w640_,
		_w641_
	);
	LUT2 #(
		.INIT('h1)
	) name469 (
		_w444_,
		_w639_,
		_w642_
	);
	LUT2 #(
		.INIT('h4)
	) name470 (
		_w641_,
		_w642_,
		_w643_
	);
	LUT2 #(
		.INIT('h1)
	) name471 (
		\y3_pad ,
		_w643_,
		_w644_
	);
	LUT2 #(
		.INIT('h8)
	) name472 (
		\y3_pad ,
		_w643_,
		_w645_
	);
	LUT2 #(
		.INIT('h2)
	) name473 (
		_w434_,
		_w644_,
		_w646_
	);
	LUT2 #(
		.INIT('h4)
	) name474 (
		_w645_,
		_w646_,
		_w647_
	);
	LUT2 #(
		.INIT('h1)
	) name475 (
		z_pad,
		_w636_,
		_w648_
	);
	LUT2 #(
		.INIT('h4)
	) name476 (
		_w647_,
		_w648_,
		_w649_
	);
	LUT2 #(
		.INIT('h1)
	) name477 (
		\z4_pad ,
		_w599_,
		_w650_
	);
	LUT2 #(
		.INIT('h8)
	) name478 (
		\z4_pad ,
		_w599_,
		_w651_
	);
	LUT2 #(
		.INIT('h2)
	) name479 (
		_w198_,
		_w650_,
		_w652_
	);
	LUT2 #(
		.INIT('h4)
	) name480 (
		_w651_,
		_w652_,
		_w653_
	);
	LUT2 #(
		.INIT('h8)
	) name481 (
		\y0_pad ,
		\z0_pad ,
		_w654_
	);
	LUT2 #(
		.INIT('h8)
	) name482 (
		_w558_,
		_w654_,
		_w655_
	);
	LUT2 #(
		.INIT('h1)
	) name483 (
		\z0_pad ,
		_w610_,
		_w656_
	);
	LUT2 #(
		.INIT('h2)
	) name484 (
		_w511_,
		_w655_,
		_w657_
	);
	LUT2 #(
		.INIT('h4)
	) name485 (
		_w656_,
		_w657_,
		_w658_
	);
	LUT2 #(
		.INIT('h2)
	) name486 (
		\d3_pad ,
		_w242_,
		_w659_
	);
	LUT2 #(
		.INIT('h2)
	) name487 (
		\y1_pad ,
		_w252_,
		_w660_
	);
	LUT2 #(
		.INIT('h4)
	) name488 (
		_w618_,
		_w660_,
		_w661_
	);
	LUT2 #(
		.INIT('h4)
	) name489 (
		\y1_pad ,
		_w252_,
		_w662_
	);
	LUT2 #(
		.INIT('h4)
	) name490 (
		_w615_,
		_w662_,
		_w663_
	);
	LUT2 #(
		.INIT('h1)
	) name491 (
		_w661_,
		_w663_,
		_w664_
	);
	LUT2 #(
		.INIT('h1)
	) name492 (
		_w263_,
		_w664_,
		_w665_
	);
	LUT2 #(
		.INIT('h1)
	) name493 (
		\z1_pad ,
		_w665_,
		_w666_
	);
	LUT2 #(
		.INIT('h8)
	) name494 (
		\z1_pad ,
		_w665_,
		_w667_
	);
	LUT2 #(
		.INIT('h2)
	) name495 (
		_w242_,
		_w666_,
		_w668_
	);
	LUT2 #(
		.INIT('h4)
	) name496 (
		_w667_,
		_w668_,
		_w669_
	);
	LUT2 #(
		.INIT('h1)
	) name497 (
		b_pad,
		_w659_,
		_w670_
	);
	LUT2 #(
		.INIT('h4)
	) name498 (
		_w669_,
		_w670_,
		_w671_
	);
	LUT2 #(
		.INIT('h1)
	) name499 (
		\y2_pad ,
		_w628_,
		_w672_
	);
	LUT2 #(
		.INIT('h2)
	) name500 (
		\y2_pad ,
		_w629_,
		_w673_
	);
	LUT2 #(
		.INIT('h1)
	) name501 (
		_w303_,
		_w672_,
		_w674_
	);
	LUT2 #(
		.INIT('h4)
	) name502 (
		_w673_,
		_w674_,
		_w675_
	);
	LUT2 #(
		.INIT('h1)
	) name503 (
		\z2_pad ,
		_w675_,
		_w676_
	);
	LUT2 #(
		.INIT('h8)
	) name504 (
		\z2_pad ,
		_w675_,
		_w677_
	);
	LUT2 #(
		.INIT('h2)
	) name505 (
		_w277_,
		_w676_,
		_w678_
	);
	LUT2 #(
		.INIT('h4)
	) name506 (
		_w677_,
		_w678_,
		_w679_
	);
	LUT2 #(
		.INIT('h1)
	) name507 (
		_w278_,
		_w679_,
		_w680_
	);
	LUT2 #(
		.INIT('h2)
	) name508 (
		\q3_pad ,
		_w434_,
		_w681_
	);
	LUT2 #(
		.INIT('h4)
	) name509 (
		\y3_pad ,
		_w638_,
		_w682_
	);
	LUT2 #(
		.INIT('h2)
	) name510 (
		_w495_,
		_w682_,
		_w683_
	);
	LUT2 #(
		.INIT('h8)
	) name511 (
		\y3_pad ,
		_w640_,
		_w684_
	);
	LUT2 #(
		.INIT('h1)
	) name512 (
		_w495_,
		_w684_,
		_w685_
	);
	LUT2 #(
		.INIT('h1)
	) name513 (
		_w444_,
		_w683_,
		_w686_
	);
	LUT2 #(
		.INIT('h4)
	) name514 (
		_w685_,
		_w686_,
		_w687_
	);
	LUT2 #(
		.INIT('h1)
	) name515 (
		\z3_pad ,
		_w687_,
		_w688_
	);
	LUT2 #(
		.INIT('h8)
	) name516 (
		\z3_pad ,
		_w687_,
		_w689_
	);
	LUT2 #(
		.INIT('h2)
	) name517 (
		_w434_,
		_w688_,
		_w690_
	);
	LUT2 #(
		.INIT('h4)
	) name518 (
		_w689_,
		_w690_,
		_w691_
	);
	LUT2 #(
		.INIT('h1)
	) name519 (
		z_pad,
		_w681_,
		_w692_
	);
	LUT2 #(
		.INIT('h4)
	) name520 (
		_w691_,
		_w692_,
		_w693_
	);
	LUT2 #(
		.INIT('h1)
	) name521 (
		\a1_pad ,
		_w655_,
		_w694_
	);
	LUT2 #(
		.INIT('h8)
	) name522 (
		\a1_pad ,
		_w655_,
		_w695_
	);
	LUT2 #(
		.INIT('h2)
	) name523 (
		_w511_,
		_w694_,
		_w696_
	);
	LUT2 #(
		.INIT('h4)
	) name524 (
		_w695_,
		_w696_,
		_w697_
	);
	LUT2 #(
		.INIT('h2)
	) name525 (
		\e3_pad ,
		_w242_,
		_w698_
	);
	LUT2 #(
		.INIT('h1)
	) name526 (
		\z1_pad ,
		_w663_,
		_w699_
	);
	LUT2 #(
		.INIT('h2)
	) name527 (
		\z1_pad ,
		_w661_,
		_w700_
	);
	LUT2 #(
		.INIT('h1)
	) name528 (
		_w263_,
		_w699_,
		_w701_
	);
	LUT2 #(
		.INIT('h4)
	) name529 (
		_w700_,
		_w701_,
		_w702_
	);
	LUT2 #(
		.INIT('h1)
	) name530 (
		\a2_pad ,
		_w702_,
		_w703_
	);
	LUT2 #(
		.INIT('h8)
	) name531 (
		\a2_pad ,
		_w702_,
		_w704_
	);
	LUT2 #(
		.INIT('h2)
	) name532 (
		_w242_,
		_w703_,
		_w705_
	);
	LUT2 #(
		.INIT('h4)
	) name533 (
		_w704_,
		_w705_,
		_w706_
	);
	LUT2 #(
		.INIT('h1)
	) name534 (
		b_pad,
		_w698_,
		_w707_
	);
	LUT2 #(
		.INIT('h4)
	) name535 (
		_w706_,
		_w707_,
		_w708_
	);
	LUT2 #(
		.INIT('h2)
	) name536 (
		\u2_pad ,
		_w530_,
		_w709_
	);
	LUT2 #(
		.INIT('h2)
	) name537 (
		_w273_,
		_w709_,
		_w710_
	);
	LUT2 #(
		.INIT('h2)
	) name538 (
		\v2_pad ,
		_w533_,
		_w711_
	);
	LUT2 #(
		.INIT('h1)
	) name539 (
		_w273_,
		_w711_,
		_w712_
	);
	LUT2 #(
		.INIT('h1)
	) name540 (
		_w303_,
		_w710_,
		_w713_
	);
	LUT2 #(
		.INIT('h4)
	) name541 (
		_w712_,
		_w713_,
		_w714_
	);
	LUT2 #(
		.INIT('h1)
	) name542 (
		\a3_pad ,
		_w714_,
		_w715_
	);
	LUT2 #(
		.INIT('h8)
	) name543 (
		\a3_pad ,
		_w714_,
		_w716_
	);
	LUT2 #(
		.INIT('h2)
	) name544 (
		_w277_,
		_w715_,
		_w717_
	);
	LUT2 #(
		.INIT('h4)
	) name545 (
		_w716_,
		_w717_,
		_w718_
	);
	LUT2 #(
		.INIT('h1)
	) name546 (
		_w278_,
		_w718_,
		_w719_
	);
	LUT2 #(
		.INIT('h1)
	) name547 (
		\r3_pad ,
		_w434_,
		_w720_
	);
	LUT2 #(
		.INIT('h4)
	) name548 (
		\z3_pad ,
		_w682_,
		_w721_
	);
	LUT2 #(
		.INIT('h2)
	) name549 (
		_w584_,
		_w721_,
		_w722_
	);
	LUT2 #(
		.INIT('h8)
	) name550 (
		\z3_pad ,
		_w684_,
		_w723_
	);
	LUT2 #(
		.INIT('h1)
	) name551 (
		\i0_pad ,
		_w495_,
		_w724_
	);
	LUT2 #(
		.INIT('h4)
	) name552 (
		_w723_,
		_w724_,
		_w725_
	);
	LUT2 #(
		.INIT('h1)
	) name553 (
		_w444_,
		_w722_,
		_w726_
	);
	LUT2 #(
		.INIT('h4)
	) name554 (
		_w725_,
		_w726_,
		_w727_
	);
	LUT2 #(
		.INIT('h1)
	) name555 (
		\a4_pad ,
		_w727_,
		_w728_
	);
	LUT2 #(
		.INIT('h8)
	) name556 (
		\a4_pad ,
		_w727_,
		_w729_
	);
	LUT2 #(
		.INIT('h1)
	) name557 (
		_w728_,
		_w729_,
		_w730_
	);
	LUT2 #(
		.INIT('h2)
	) name558 (
		_w434_,
		_w730_,
		_w731_
	);
	LUT2 #(
		.INIT('h1)
	) name559 (
		z_pad,
		_w720_,
		_w732_
	);
	LUT2 #(
		.INIT('h4)
	) name560 (
		_w731_,
		_w732_,
		_w733_
	);
	LUT2 #(
		.INIT('h1)
	) name561 (
		\b1_pad ,
		_w695_,
		_w734_
	);
	LUT2 #(
		.INIT('h8)
	) name562 (
		\b1_pad ,
		_w695_,
		_w735_
	);
	LUT2 #(
		.INIT('h2)
	) name563 (
		_w511_,
		_w734_,
		_w736_
	);
	LUT2 #(
		.INIT('h4)
	) name564 (
		_w735_,
		_w736_,
		_w737_
	);
	LUT2 #(
		.INIT('h2)
	) name565 (
		\b2_pad ,
		b_pad,
		_w738_
	);
	LUT2 #(
		.INIT('h4)
	) name566 (
		\a3_pad ,
		_w709_,
		_w739_
	);
	LUT2 #(
		.INIT('h1)
	) name567 (
		j_pad,
		_w739_,
		_w740_
	);
	LUT2 #(
		.INIT('h8)
	) name568 (
		_w273_,
		_w740_,
		_w741_
	);
	LUT2 #(
		.INIT('h8)
	) name569 (
		\a3_pad ,
		_w711_,
		_w742_
	);
	LUT2 #(
		.INIT('h1)
	) name570 (
		j_pad,
		_w273_,
		_w743_
	);
	LUT2 #(
		.INIT('h4)
	) name571 (
		_w742_,
		_w743_,
		_w744_
	);
	LUT2 #(
		.INIT('h1)
	) name572 (
		_w303_,
		_w744_,
		_w745_
	);
	LUT2 #(
		.INIT('h4)
	) name573 (
		_w741_,
		_w745_,
		_w746_
	);
	LUT2 #(
		.INIT('h1)
	) name574 (
		\b3_pad ,
		_w746_,
		_w747_
	);
	LUT2 #(
		.INIT('h8)
	) name575 (
		\b3_pad ,
		_w746_,
		_w748_
	);
	LUT2 #(
		.INIT('h2)
	) name576 (
		_w277_,
		_w747_,
		_w749_
	);
	LUT2 #(
		.INIT('h4)
	) name577 (
		_w748_,
		_w749_,
		_w750_
	);
	LUT2 #(
		.INIT('h1)
	) name578 (
		_w278_,
		_w750_,
		_w751_
	);
	LUT2 #(
		.INIT('h2)
	) name579 (
		\s3_pad ,
		_w434_,
		_w752_
	);
	LUT2 #(
		.INIT('h1)
	) name580 (
		\a4_pad ,
		_w495_,
		_w753_
	);
	LUT2 #(
		.INIT('h8)
	) name581 (
		\a4_pad ,
		_w495_,
		_w754_
	);
	LUT2 #(
		.INIT('h1)
	) name582 (
		_w753_,
		_w754_,
		_w755_
	);
	LUT2 #(
		.INIT('h8)
	) name583 (
		_w727_,
		_w755_,
		_w756_
	);
	LUT2 #(
		.INIT('h2)
	) name584 (
		\b4_pad ,
		_w756_,
		_w757_
	);
	LUT2 #(
		.INIT('h4)
	) name585 (
		\b4_pad ,
		_w756_,
		_w758_
	);
	LUT2 #(
		.INIT('h1)
	) name586 (
		_w757_,
		_w758_,
		_w759_
	);
	LUT2 #(
		.INIT('h2)
	) name587 (
		_w434_,
		_w759_,
		_w760_
	);
	LUT2 #(
		.INIT('h1)
	) name588 (
		z_pad,
		_w752_,
		_w761_
	);
	LUT2 #(
		.INIT('h4)
	) name589 (
		_w760_,
		_w761_,
		_w762_
	);
	LUT2 #(
		.INIT('h1)
	) name590 (
		\c1_pad ,
		_w735_,
		_w763_
	);
	LUT2 #(
		.INIT('h8)
	) name591 (
		\c1_pad ,
		_w735_,
		_w764_
	);
	LUT2 #(
		.INIT('h2)
	) name592 (
		_w511_,
		_w763_,
		_w765_
	);
	LUT2 #(
		.INIT('h4)
	) name593 (
		_w764_,
		_w765_,
		_w766_
	);
	LUT2 #(
		.INIT('h1)
	) name594 (
		\b2_pad ,
		\c2_pad ,
		_w767_
	);
	LUT2 #(
		.INIT('h8)
	) name595 (
		\b2_pad ,
		\c2_pad ,
		_w768_
	);
	LUT2 #(
		.INIT('h1)
	) name596 (
		_w767_,
		_w768_,
		_w769_
	);
	LUT2 #(
		.INIT('h1)
	) name597 (
		b_pad,
		_w769_,
		_w770_
	);
	LUT2 #(
		.INIT('h1)
	) name598 (
		\b3_pad ,
		_w740_,
		_w771_
	);
	LUT2 #(
		.INIT('h2)
	) name599 (
		_w273_,
		_w771_,
		_w772_
	);
	LUT2 #(
		.INIT('h1)
	) name600 (
		\b3_pad ,
		_w273_,
		_w773_
	);
	LUT2 #(
		.INIT('h2)
	) name601 (
		_w745_,
		_w773_,
		_w774_
	);
	LUT2 #(
		.INIT('h4)
	) name602 (
		_w772_,
		_w774_,
		_w775_
	);
	LUT2 #(
		.INIT('h1)
	) name603 (
		\c3_pad ,
		_w775_,
		_w776_
	);
	LUT2 #(
		.INIT('h8)
	) name604 (
		\c3_pad ,
		_w775_,
		_w777_
	);
	LUT2 #(
		.INIT('h2)
	) name605 (
		_w277_,
		_w776_,
		_w778_
	);
	LUT2 #(
		.INIT('h4)
	) name606 (
		_w777_,
		_w778_,
		_w779_
	);
	LUT2 #(
		.INIT('h2)
	) name607 (
		\t3_pad ,
		_w434_,
		_w780_
	);
	LUT2 #(
		.INIT('h1)
	) name608 (
		\b4_pad ,
		_w495_,
		_w781_
	);
	LUT2 #(
		.INIT('h8)
	) name609 (
		\b4_pad ,
		_w495_,
		_w782_
	);
	LUT2 #(
		.INIT('h1)
	) name610 (
		_w781_,
		_w782_,
		_w783_
	);
	LUT2 #(
		.INIT('h8)
	) name611 (
		_w756_,
		_w783_,
		_w784_
	);
	LUT2 #(
		.INIT('h1)
	) name612 (
		\c4_pad ,
		_w784_,
		_w785_
	);
	LUT2 #(
		.INIT('h8)
	) name613 (
		\c4_pad ,
		_w784_,
		_w786_
	);
	LUT2 #(
		.INIT('h2)
	) name614 (
		_w434_,
		_w785_,
		_w787_
	);
	LUT2 #(
		.INIT('h4)
	) name615 (
		_w786_,
		_w787_,
		_w788_
	);
	LUT2 #(
		.INIT('h1)
	) name616 (
		z_pad,
		_w780_,
		_w789_
	);
	LUT2 #(
		.INIT('h4)
	) name617 (
		_w788_,
		_w789_,
		_w790_
	);
	LUT2 #(
		.INIT('h2)
	) name618 (
		\d5_pad ,
		_w185_,
		_w791_
	);
	LUT2 #(
		.INIT('h8)
	) name619 (
		_w181_,
		_w791_,
		_w792_
	);
	LUT2 #(
		.INIT('h1)
	) name620 (
		_w191_,
		_w792_,
		_w793_
	);
	LUT2 #(
		.INIT('h8)
	) name621 (
		_w185_,
		_w315_,
		_w794_
	);
	LUT2 #(
		.INIT('h2)
	) name622 (
		_w175_,
		_w459_,
		_w795_
	);
	LUT2 #(
		.INIT('h1)
	) name623 (
		_w433_,
		_w794_,
		_w796_
	);
	LUT2 #(
		.INIT('h4)
	) name624 (
		_w795_,
		_w796_,
		_w797_
	);
	LUT2 #(
		.INIT('h1)
	) name625 (
		\d1_pad ,
		_w764_,
		_w798_
	);
	LUT2 #(
		.INIT('h8)
	) name626 (
		\d1_pad ,
		_w764_,
		_w799_
	);
	LUT2 #(
		.INIT('h2)
	) name627 (
		_w511_,
		_w798_,
		_w800_
	);
	LUT2 #(
		.INIT('h4)
	) name628 (
		_w799_,
		_w800_,
		_w801_
	);
	LUT2 #(
		.INIT('h8)
	) name629 (
		\d2_pad ,
		_w768_,
		_w802_
	);
	LUT2 #(
		.INIT('h1)
	) name630 (
		\d2_pad ,
		_w768_,
		_w803_
	);
	LUT2 #(
		.INIT('h1)
	) name631 (
		_w802_,
		_w803_,
		_w804_
	);
	LUT2 #(
		.INIT('h1)
	) name632 (
		b_pad,
		_w804_,
		_w805_
	);
	LUT2 #(
		.INIT('h1)
	) name633 (
		\c3_pad ,
		_w273_,
		_w806_
	);
	LUT2 #(
		.INIT('h8)
	) name634 (
		\c3_pad ,
		_w273_,
		_w807_
	);
	LUT2 #(
		.INIT('h1)
	) name635 (
		_w806_,
		_w807_,
		_w808_
	);
	LUT2 #(
		.INIT('h8)
	) name636 (
		_w775_,
		_w808_,
		_w809_
	);
	LUT2 #(
		.INIT('h1)
	) name637 (
		\d3_pad ,
		_w809_,
		_w810_
	);
	LUT2 #(
		.INIT('h8)
	) name638 (
		\d3_pad ,
		_w809_,
		_w811_
	);
	LUT2 #(
		.INIT('h2)
	) name639 (
		_w277_,
		_w810_,
		_w812_
	);
	LUT2 #(
		.INIT('h4)
	) name640 (
		_w811_,
		_w812_,
		_w813_
	);
	LUT2 #(
		.INIT('h1)
	) name641 (
		_w278_,
		_w813_,
		_w814_
	);
	LUT2 #(
		.INIT('h2)
	) name642 (
		\d4_pad ,
		z_pad,
		_w815_
	);
	LUT2 #(
		.INIT('h2)
	) name643 (
		\e5_pad ,
		_w183_,
		_w816_
	);
	LUT2 #(
		.INIT('h8)
	) name644 (
		_w181_,
		_w816_,
		_w817_
	);
	LUT2 #(
		.INIT('h1)
	) name645 (
		_w187_,
		_w817_,
		_w818_
	);
	LUT2 #(
		.INIT('h4)
	) name646 (
		l_pad,
		\q1_pad ,
		_w819_
	);
	LUT2 #(
		.INIT('h1)
	) name647 (
		_w802_,
		_w819_,
		_w820_
	);
	LUT2 #(
		.INIT('h2)
	) name648 (
		\g2_pad ,
		_w820_,
		_w821_
	);
	LUT2 #(
		.INIT('h1)
	) name649 (
		l_pad,
		\p1_pad ,
		_w822_
	);
	LUT2 #(
		.INIT('h4)
	) name650 (
		_w821_,
		_w822_,
		_w823_
	);
	LUT2 #(
		.INIT('h2)
	) name651 (
		\e2_pad ,
		_w823_,
		_w824_
	);
	LUT2 #(
		.INIT('h8)
	) name652 (
		\n2_pad ,
		_w824_,
		_w825_
	);
	LUT2 #(
		.INIT('h1)
	) name653 (
		_w464_,
		_w825_,
		_w826_
	);
	LUT2 #(
		.INIT('h2)
	) name654 (
		\s1_pad ,
		_w826_,
		_w827_
	);
	LUT2 #(
		.INIT('h4)
	) name655 (
		\e2_pad ,
		_w823_,
		_w828_
	);
	LUT2 #(
		.INIT('h1)
	) name656 (
		_w824_,
		_w828_,
		_w829_
	);
	LUT2 #(
		.INIT('h8)
	) name657 (
		_w826_,
		_w829_,
		_w830_
	);
	LUT2 #(
		.INIT('h1)
	) name658 (
		b_pad,
		_w827_,
		_w831_
	);
	LUT2 #(
		.INIT('h4)
	) name659 (
		_w830_,
		_w831_,
		_w832_
	);
	LUT2 #(
		.INIT('h1)
	) name660 (
		\c3_pad ,
		\d3_pad ,
		_w833_
	);
	LUT2 #(
		.INIT('h8)
	) name661 (
		_w771_,
		_w833_,
		_w834_
	);
	LUT2 #(
		.INIT('h2)
	) name662 (
		_w273_,
		_w834_,
		_w835_
	);
	LUT2 #(
		.INIT('h1)
	) name663 (
		_w273_,
		_w603_,
		_w836_
	);
	LUT2 #(
		.INIT('h2)
	) name664 (
		_w774_,
		_w836_,
		_w837_
	);
	LUT2 #(
		.INIT('h4)
	) name665 (
		_w835_,
		_w837_,
		_w838_
	);
	LUT2 #(
		.INIT('h1)
	) name666 (
		\e3_pad ,
		_w838_,
		_w839_
	);
	LUT2 #(
		.INIT('h8)
	) name667 (
		\e3_pad ,
		_w838_,
		_w840_
	);
	LUT2 #(
		.INIT('h2)
	) name668 (
		_w277_,
		_w839_,
		_w841_
	);
	LUT2 #(
		.INIT('h4)
	) name669 (
		_w840_,
		_w841_,
		_w842_
	);
	LUT2 #(
		.INIT('h1)
	) name670 (
		_w278_,
		_w842_,
		_w843_
	);
	LUT2 #(
		.INIT('h1)
	) name671 (
		\d4_pad ,
		\e4_pad ,
		_w844_
	);
	LUT2 #(
		.INIT('h1)
	) name672 (
		_w395_,
		_w844_,
		_w845_
	);
	LUT2 #(
		.INIT('h1)
	) name673 (
		z_pad,
		_w845_,
		_w846_
	);
	LUT2 #(
		.INIT('h2)
	) name674 (
		\h5_pad ,
		_w402_,
		_w847_
	);
	LUT2 #(
		.INIT('h4)
	) name675 (
		\h5_pad ,
		_w402_,
		_w848_
	);
	LUT2 #(
		.INIT('h1)
	) name676 (
		_w178_,
		_w847_,
		_w849_
	);
	LUT2 #(
		.INIT('h4)
	) name677 (
		_w848_,
		_w849_,
		_w850_
	);
	LUT2 #(
		.INIT('h1)
	) name678 (
		z_pad,
		_w850_,
		_w851_
	);
	LUT2 #(
		.INIT('h4)
	) name679 (
		\h5_pad ,
		_w851_,
		_w852_
	);
	LUT2 #(
		.INIT('h4)
	) name680 (
		\p10_pad ,
		_w852_,
		_w853_
	);
	LUT2 #(
		.INIT('h1)
	) name681 (
		\f5_pad ,
		_w853_,
		_w854_
	);
	LUT2 #(
		.INIT('h8)
	) name682 (
		\f5_pad ,
		_w852_,
		_w855_
	);
	LUT2 #(
		.INIT('h1)
	) name683 (
		_w178_,
		_w855_,
		_w856_
	);
	LUT2 #(
		.INIT('h4)
	) name684 (
		_w854_,
		_w856_,
		_w857_
	);
	LUT2 #(
		.INIT('h1)
	) name685 (
		z_pad,
		_w857_,
		_w858_
	);
	LUT2 #(
		.INIT('h2)
	) name686 (
		\t1_pad ,
		_w826_,
		_w859_
	);
	LUT2 #(
		.INIT('h8)
	) name687 (
		\f2_pad ,
		_w824_,
		_w860_
	);
	LUT2 #(
		.INIT('h1)
	) name688 (
		\f2_pad ,
		_w824_,
		_w861_
	);
	LUT2 #(
		.INIT('h1)
	) name689 (
		_w860_,
		_w861_,
		_w862_
	);
	LUT2 #(
		.INIT('h8)
	) name690 (
		_w826_,
		_w862_,
		_w863_
	);
	LUT2 #(
		.INIT('h1)
	) name691 (
		b_pad,
		_w859_,
		_w864_
	);
	LUT2 #(
		.INIT('h4)
	) name692 (
		_w863_,
		_w864_,
		_w865_
	);
	LUT2 #(
		.INIT('h2)
	) name693 (
		\f3_pad ,
		_w350_,
		_w866_
	);
	LUT2 #(
		.INIT('h4)
	) name694 (
		\f3_pad ,
		_w350_,
		_w867_
	);
	LUT2 #(
		.INIT('h2)
	) name695 (
		_w316_,
		_w866_,
		_w868_
	);
	LUT2 #(
		.INIT('h4)
	) name696 (
		_w867_,
		_w868_,
		_w869_
	);
	LUT2 #(
		.INIT('h1)
	) name697 (
		\f4_pad ,
		_w395_,
		_w870_
	);
	LUT2 #(
		.INIT('h1)
	) name698 (
		_w396_,
		_w870_,
		_w871_
	);
	LUT2 #(
		.INIT('h1)
	) name699 (
		z_pad,
		_w871_,
		_w872_
	);
	LUT2 #(
		.INIT('h2)
	) name700 (
		\p10_pad ,
		_w852_,
		_w873_
	);
	LUT2 #(
		.INIT('h2)
	) name701 (
		_w856_,
		_w873_,
		_w874_
	);
	LUT2 #(
		.INIT('h1)
	) name702 (
		z_pad,
		_w874_,
		_w875_
	);
	LUT2 #(
		.INIT('h4)
	) name703 (
		\g2_pad ,
		_w820_,
		_w876_
	);
	LUT2 #(
		.INIT('h1)
	) name704 (
		_w821_,
		_w876_,
		_w877_
	);
	LUT2 #(
		.INIT('h1)
	) name705 (
		b_pad,
		_w877_,
		_w878_
	);
	LUT2 #(
		.INIT('h1)
	) name706 (
		\f3_pad ,
		_w313_,
		_w879_
	);
	LUT2 #(
		.INIT('h8)
	) name707 (
		\f3_pad ,
		_w313_,
		_w880_
	);
	LUT2 #(
		.INIT('h1)
	) name708 (
		_w350_,
		_w879_,
		_w881_
	);
	LUT2 #(
		.INIT('h4)
	) name709 (
		_w880_,
		_w881_,
		_w882_
	);
	LUT2 #(
		.INIT('h8)
	) name710 (
		\g3_pad ,
		_w882_,
		_w883_
	);
	LUT2 #(
		.INIT('h1)
	) name711 (
		\g3_pad ,
		_w882_,
		_w884_
	);
	LUT2 #(
		.INIT('h2)
	) name712 (
		_w316_,
		_w883_,
		_w885_
	);
	LUT2 #(
		.INIT('h4)
	) name713 (
		_w884_,
		_w885_,
		_w886_
	);
	LUT2 #(
		.INIT('h1)
	) name714 (
		_w180_,
		_w402_,
		_w887_
	);
	LUT2 #(
		.INIT('h2)
	) name715 (
		\u3_pad ,
		_w887_,
		_w888_
	);
	LUT2 #(
		.INIT('h4)
	) name716 (
		\g4_pad ,
		_w400_,
		_w889_
	);
	LUT2 #(
		.INIT('h1)
	) name717 (
		_w401_,
		_w889_,
		_w890_
	);
	LUT2 #(
		.INIT('h8)
	) name718 (
		_w887_,
		_w890_,
		_w891_
	);
	LUT2 #(
		.INIT('h1)
	) name719 (
		z_pad,
		_w888_,
		_w892_
	);
	LUT2 #(
		.INIT('h4)
	) name720 (
		_w891_,
		_w892_,
		_w893_
	);
	LUT2 #(
		.INIT('h2)
	) name721 (
		\h1_pad ,
		_w247_,
		_w894_
	);
	LUT2 #(
		.INIT('h8)
	) name722 (
		_w465_,
		_w894_,
		_w895_
	);
	LUT2 #(
		.INIT('h1)
	) name723 (
		_w297_,
		_w895_,
		_w896_
	);
	LUT2 #(
		.INIT('h1)
	) name724 (
		\h2_pad ,
		_w860_,
		_w897_
	);
	LUT2 #(
		.INIT('h8)
	) name725 (
		\f2_pad ,
		\h2_pad ,
		_w898_
	);
	LUT2 #(
		.INIT('h8)
	) name726 (
		_w824_,
		_w898_,
		_w899_
	);
	LUT2 #(
		.INIT('h2)
	) name727 (
		_w826_,
		_w899_,
		_w900_
	);
	LUT2 #(
		.INIT('h4)
	) name728 (
		_w897_,
		_w900_,
		_w901_
	);
	LUT2 #(
		.INIT('h2)
	) name729 (
		\u1_pad ,
		_w826_,
		_w902_
	);
	LUT2 #(
		.INIT('h1)
	) name730 (
		b_pad,
		_w902_,
		_w903_
	);
	LUT2 #(
		.INIT('h4)
	) name731 (
		_w901_,
		_w903_,
		_w904_
	);
	LUT2 #(
		.INIT('h8)
	) name732 (
		_w313_,
		_w321_,
		_w905_
	);
	LUT2 #(
		.INIT('h4)
	) name733 (
		_w313_,
		_w352_,
		_w906_
	);
	LUT2 #(
		.INIT('h1)
	) name734 (
		_w350_,
		_w905_,
		_w907_
	);
	LUT2 #(
		.INIT('h4)
	) name735 (
		_w906_,
		_w907_,
		_w908_
	);
	LUT2 #(
		.INIT('h8)
	) name736 (
		\h3_pad ,
		_w908_,
		_w909_
	);
	LUT2 #(
		.INIT('h1)
	) name737 (
		\h3_pad ,
		_w908_,
		_w910_
	);
	LUT2 #(
		.INIT('h2)
	) name738 (
		_w316_,
		_w909_,
		_w911_
	);
	LUT2 #(
		.INIT('h4)
	) name739 (
		_w910_,
		_w911_,
		_w912_
	);
	LUT2 #(
		.INIT('h2)
	) name740 (
		\v3_pad ,
		_w887_,
		_w913_
	);
	LUT2 #(
		.INIT('h8)
	) name741 (
		\h4_pad ,
		_w401_,
		_w914_
	);
	LUT2 #(
		.INIT('h1)
	) name742 (
		\h4_pad ,
		_w401_,
		_w915_
	);
	LUT2 #(
		.INIT('h1)
	) name743 (
		_w914_,
		_w915_,
		_w916_
	);
	LUT2 #(
		.INIT('h8)
	) name744 (
		_w887_,
		_w916_,
		_w917_
	);
	LUT2 #(
		.INIT('h1)
	) name745 (
		z_pad,
		_w913_,
		_w918_
	);
	LUT2 #(
		.INIT('h4)
	) name746 (
		_w917_,
		_w918_,
		_w919_
	);
	LUT2 #(
		.INIT('h2)
	) name747 (
		\i1_pad ,
		_w245_,
		_w920_
	);
	LUT2 #(
		.INIT('h8)
	) name748 (
		_w465_,
		_w920_,
		_w921_
	);
	LUT2 #(
		.INIT('h1)
	) name749 (
		_w249_,
		_w921_,
		_w922_
	);
	LUT2 #(
		.INIT('h2)
	) name750 (
		\v1_pad ,
		_w826_,
		_w923_
	);
	LUT2 #(
		.INIT('h8)
	) name751 (
		\i2_pad ,
		_w899_,
		_w924_
	);
	LUT2 #(
		.INIT('h1)
	) name752 (
		\i2_pad ,
		_w899_,
		_w925_
	);
	LUT2 #(
		.INIT('h2)
	) name753 (
		_w826_,
		_w924_,
		_w926_
	);
	LUT2 #(
		.INIT('h4)
	) name754 (
		_w925_,
		_w926_,
		_w927_
	);
	LUT2 #(
		.INIT('h1)
	) name755 (
		b_pad,
		_w923_,
		_w928_
	);
	LUT2 #(
		.INIT('h4)
	) name756 (
		_w927_,
		_w928_,
		_w929_
	);
	LUT2 #(
		.INIT('h8)
	) name757 (
		_w313_,
		_w325_,
		_w930_
	);
	LUT2 #(
		.INIT('h4)
	) name758 (
		_w313_,
		_w354_,
		_w931_
	);
	LUT2 #(
		.INIT('h1)
	) name759 (
		_w350_,
		_w930_,
		_w932_
	);
	LUT2 #(
		.INIT('h4)
	) name760 (
		_w931_,
		_w932_,
		_w933_
	);
	LUT2 #(
		.INIT('h1)
	) name761 (
		\i3_pad ,
		_w933_,
		_w934_
	);
	LUT2 #(
		.INIT('h8)
	) name762 (
		\i3_pad ,
		_w933_,
		_w935_
	);
	LUT2 #(
		.INIT('h2)
	) name763 (
		_w316_,
		_w934_,
		_w936_
	);
	LUT2 #(
		.INIT('h4)
	) name764 (
		_w935_,
		_w936_,
		_w937_
	);
	LUT2 #(
		.INIT('h1)
	) name765 (
		_w317_,
		_w937_,
		_w938_
	);
	LUT2 #(
		.INIT('h4)
	) name766 (
		\i4_pad ,
		_w397_,
		_w939_
	);
	LUT2 #(
		.INIT('h1)
	) name767 (
		_w398_,
		_w939_,
		_w940_
	);
	LUT2 #(
		.INIT('h1)
	) name768 (
		z_pad,
		_w940_,
		_w941_
	);
	LUT2 #(
		.INIT('h1)
	) name769 (
		z_pad,
		_w336_,
		_w942_
	);
	LUT2 #(
		.INIT('h1)
	) name770 (
		\j5_pad ,
		_w175_,
		_w943_
	);
	LUT2 #(
		.INIT('h8)
	) name771 (
		\j5_pad ,
		_w175_,
		_w944_
	);
	LUT2 #(
		.INIT('h2)
	) name772 (
		_w942_,
		_w943_,
		_w945_
	);
	LUT2 #(
		.INIT('h4)
	) name773 (
		_w944_,
		_w945_,
		_w946_
	);
	LUT2 #(
		.INIT('h8)
	) name774 (
		\r6_pad ,
		_w825_,
		_w947_
	);
	LUT2 #(
		.INIT('h1)
	) name775 (
		\r6_pad ,
		_w825_,
		_w948_
	);
	LUT2 #(
		.INIT('h1)
	) name776 (
		b_pad,
		_w947_,
		_w949_
	);
	LUT2 #(
		.INIT('h4)
	) name777 (
		_w948_,
		_w949_,
		_w950_
	);
	LUT2 #(
		.INIT('h1)
	) name778 (
		_w228_,
		_w950_,
		_w951_
	);
	LUT2 #(
		.INIT('h2)
	) name779 (
		\w1_pad ,
		_w826_,
		_w952_
	);
	LUT2 #(
		.INIT('h1)
	) name780 (
		\j2_pad ,
		_w924_,
		_w953_
	);
	LUT2 #(
		.INIT('h8)
	) name781 (
		\i2_pad ,
		\j2_pad ,
		_w954_
	);
	LUT2 #(
		.INIT('h8)
	) name782 (
		_w898_,
		_w954_,
		_w955_
	);
	LUT2 #(
		.INIT('h8)
	) name783 (
		_w824_,
		_w955_,
		_w956_
	);
	LUT2 #(
		.INIT('h2)
	) name784 (
		_w826_,
		_w956_,
		_w957_
	);
	LUT2 #(
		.INIT('h4)
	) name785 (
		_w953_,
		_w957_,
		_w958_
	);
	LUT2 #(
		.INIT('h1)
	) name786 (
		b_pad,
		_w952_,
		_w959_
	);
	LUT2 #(
		.INIT('h4)
	) name787 (
		_w958_,
		_w959_,
		_w960_
	);
	LUT2 #(
		.INIT('h1)
	) name788 (
		\l3_pad ,
		\m3_pad ,
		_w961_
	);
	LUT2 #(
		.INIT('h1)
	) name789 (
		\n3_pad ,
		\o3_pad ,
		_w962_
	);
	LUT2 #(
		.INIT('h8)
	) name790 (
		_w961_,
		_w962_,
		_w963_
	);
	LUT2 #(
		.INIT('h2)
	) name791 (
		_w316_,
		_w963_,
		_w964_
	);
	LUT2 #(
		.INIT('h1)
	) name792 (
		_w317_,
		_w964_,
		_w965_
	);
	LUT2 #(
		.INIT('h1)
	) name793 (
		\j4_pad ,
		_w914_,
		_w966_
	);
	LUT2 #(
		.INIT('h8)
	) name794 (
		\h4_pad ,
		\j4_pad ,
		_w967_
	);
	LUT2 #(
		.INIT('h8)
	) name795 (
		_w401_,
		_w967_,
		_w968_
	);
	LUT2 #(
		.INIT('h2)
	) name796 (
		_w887_,
		_w968_,
		_w969_
	);
	LUT2 #(
		.INIT('h4)
	) name797 (
		_w966_,
		_w969_,
		_w970_
	);
	LUT2 #(
		.INIT('h2)
	) name798 (
		\w3_pad ,
		_w887_,
		_w971_
	);
	LUT2 #(
		.INIT('h1)
	) name799 (
		z_pad,
		_w971_,
		_w972_
	);
	LUT2 #(
		.INIT('h4)
	) name800 (
		_w970_,
		_w972_,
		_w973_
	);
	LUT2 #(
		.INIT('h1)
	) name801 (
		\k5_pad ,
		_w944_,
		_w974_
	);
	LUT2 #(
		.INIT('h8)
	) name802 (
		\k5_pad ,
		_w944_,
		_w975_
	);
	LUT2 #(
		.INIT('h2)
	) name803 (
		_w942_,
		_w974_,
		_w976_
	);
	LUT2 #(
		.INIT('h4)
	) name804 (
		_w975_,
		_w976_,
		_w977_
	);
	LUT2 #(
		.INIT('h2)
	) name805 (
		\x1_pad ,
		_w826_,
		_w978_
	);
	LUT2 #(
		.INIT('h1)
	) name806 (
		l_pad,
		_w956_,
		_w979_
	);
	LUT2 #(
		.INIT('h2)
	) name807 (
		\k2_pad ,
		_w979_,
		_w980_
	);
	LUT2 #(
		.INIT('h4)
	) name808 (
		\k2_pad ,
		_w979_,
		_w981_
	);
	LUT2 #(
		.INIT('h2)
	) name809 (
		_w826_,
		_w980_,
		_w982_
	);
	LUT2 #(
		.INIT('h4)
	) name810 (
		_w981_,
		_w982_,
		_w983_
	);
	LUT2 #(
		.INIT('h1)
	) name811 (
		b_pad,
		_w978_,
		_w984_
	);
	LUT2 #(
		.INIT('h4)
	) name812 (
		_w983_,
		_w984_,
		_w985_
	);
	LUT2 #(
		.INIT('h8)
	) name813 (
		\l3_pad ,
		\m3_pad ,
		_w986_
	);
	LUT2 #(
		.INIT('h8)
	) name814 (
		\n3_pad ,
		\o3_pad ,
		_w987_
	);
	LUT2 #(
		.INIT('h8)
	) name815 (
		_w986_,
		_w987_,
		_w988_
	);
	LUT2 #(
		.INIT('h8)
	) name816 (
		_w316_,
		_w988_,
		_w989_
	);
	LUT2 #(
		.INIT('h2)
	) name817 (
		\x3_pad ,
		_w887_,
		_w990_
	);
	LUT2 #(
		.INIT('h8)
	) name818 (
		\k4_pad ,
		_w968_,
		_w991_
	);
	LUT2 #(
		.INIT('h1)
	) name819 (
		\k4_pad ,
		_w968_,
		_w992_
	);
	LUT2 #(
		.INIT('h2)
	) name820 (
		_w887_,
		_w991_,
		_w993_
	);
	LUT2 #(
		.INIT('h4)
	) name821 (
		_w992_,
		_w993_,
		_w994_
	);
	LUT2 #(
		.INIT('h1)
	) name822 (
		z_pad,
		_w990_,
		_w995_
	);
	LUT2 #(
		.INIT('h4)
	) name823 (
		_w994_,
		_w995_,
		_w996_
	);
	LUT2 #(
		.INIT('h8)
	) name824 (
		\a2_pad ,
		p_pad,
		_w997_
	);
	LUT2 #(
		.INIT('h8)
	) name825 (
		w_pad,
		\y0_pad ,
		_w998_
	);
	LUT2 #(
		.INIT('h8)
	) name826 (
		\d1_pad ,
		v_pad,
		_w999_
	);
	LUT2 #(
		.INIT('h8)
	) name827 (
		\g2_pad ,
		u_pad,
		_w1000_
	);
	LUT2 #(
		.INIT('h8)
	) name828 (
		q_pad,
		\x1_pad ,
		_w1001_
	);
	LUT2 #(
		.INIT('h8)
	) name829 (
		\j2_pad ,
		t_pad,
		_w1002_
	);
	LUT2 #(
		.INIT('h8)
	) name830 (
		\a3_pad ,
		n_pad,
		_w1003_
	);
	LUT2 #(
		.INIT('h8)
	) name831 (
		\e3_pad ,
		m_pad,
		_w1004_
	);
	LUT2 #(
		.INIT('h8)
	) name832 (
		r_pad,
		\u1_pad ,
		_w1005_
	);
	LUT2 #(
		.INIT('h8)
	) name833 (
		o_pad,
		\t2_pad ,
		_w1006_
	);
	LUT2 #(
		.INIT('h8)
	) name834 (
		\o2_pad ,
		s_pad,
		_w1007_
	);
	LUT2 #(
		.INIT('h1)
	) name835 (
		_w997_,
		_w998_,
		_w1008_
	);
	LUT2 #(
		.INIT('h1)
	) name836 (
		_w999_,
		_w1000_,
		_w1009_
	);
	LUT2 #(
		.INIT('h1)
	) name837 (
		_w1001_,
		_w1002_,
		_w1010_
	);
	LUT2 #(
		.INIT('h1)
	) name838 (
		_w1003_,
		_w1004_,
		_w1011_
	);
	LUT2 #(
		.INIT('h1)
	) name839 (
		_w1005_,
		_w1006_,
		_w1012_
	);
	LUT2 #(
		.INIT('h4)
	) name840 (
		_w1007_,
		_w1012_,
		_w1013_
	);
	LUT2 #(
		.INIT('h8)
	) name841 (
		_w1010_,
		_w1011_,
		_w1014_
	);
	LUT2 #(
		.INIT('h8)
	) name842 (
		_w1008_,
		_w1009_,
		_w1015_
	);
	LUT2 #(
		.INIT('h8)
	) name843 (
		_w1014_,
		_w1015_,
		_w1016_
	);
	LUT2 #(
		.INIT('h8)
	) name844 (
		_w1013_,
		_w1016_,
		_w1017_
	);
	LUT2 #(
		.INIT('h2)
	) name845 (
		\y1_pad ,
		_w826_,
		_w1018_
	);
	LUT2 #(
		.INIT('h1)
	) name846 (
		\l2_pad ,
		_w980_,
		_w1019_
	);
	LUT2 #(
		.INIT('h8)
	) name847 (
		\l2_pad ,
		_w980_,
		_w1020_
	);
	LUT2 #(
		.INIT('h2)
	) name848 (
		_w826_,
		_w1019_,
		_w1021_
	);
	LUT2 #(
		.INIT('h4)
	) name849 (
		_w1020_,
		_w1021_,
		_w1022_
	);
	LUT2 #(
		.INIT('h1)
	) name850 (
		b_pad,
		_w1018_,
		_w1023_
	);
	LUT2 #(
		.INIT('h4)
	) name851 (
		_w1022_,
		_w1023_,
		_w1024_
	);
	LUT2 #(
		.INIT('h4)
	) name852 (
		_w313_,
		_w356_,
		_w1025_
	);
	LUT2 #(
		.INIT('h8)
	) name853 (
		_w313_,
		_w327_,
		_w1026_
	);
	LUT2 #(
		.INIT('h1)
	) name854 (
		_w350_,
		_w1025_,
		_w1027_
	);
	LUT2 #(
		.INIT('h4)
	) name855 (
		_w1026_,
		_w1027_,
		_w1028_
	);
	LUT2 #(
		.INIT('h1)
	) name856 (
		\l3_pad ,
		_w1028_,
		_w1029_
	);
	LUT2 #(
		.INIT('h8)
	) name857 (
		\l3_pad ,
		_w1028_,
		_w1030_
	);
	LUT2 #(
		.INIT('h2)
	) name858 (
		_w316_,
		_w1029_,
		_w1031_
	);
	LUT2 #(
		.INIT('h4)
	) name859 (
		_w1030_,
		_w1031_,
		_w1032_
	);
	LUT2 #(
		.INIT('h2)
	) name860 (
		\y3_pad ,
		_w887_,
		_w1033_
	);
	LUT2 #(
		.INIT('h1)
	) name861 (
		\l4_pad ,
		_w991_,
		_w1034_
	);
	LUT2 #(
		.INIT('h8)
	) name862 (
		\k4_pad ,
		\l4_pad ,
		_w1035_
	);
	LUT2 #(
		.INIT('h8)
	) name863 (
		_w967_,
		_w1035_,
		_w1036_
	);
	LUT2 #(
		.INIT('h8)
	) name864 (
		_w401_,
		_w1036_,
		_w1037_
	);
	LUT2 #(
		.INIT('h2)
	) name865 (
		_w887_,
		_w1037_,
		_w1038_
	);
	LUT2 #(
		.INIT('h4)
	) name866 (
		_w1034_,
		_w1038_,
		_w1039_
	);
	LUT2 #(
		.INIT('h1)
	) name867 (
		z_pad,
		_w1033_,
		_w1040_
	);
	LUT2 #(
		.INIT('h4)
	) name868 (
		_w1039_,
		_w1040_,
		_w1041_
	);
	LUT2 #(
		.INIT('h2)
	) name869 (
		\r5_pad ,
		_w599_,
		_w1042_
	);
	LUT2 #(
		.INIT('h2)
	) name870 (
		\z4_pad ,
		_w1042_,
		_w1043_
	);
	LUT2 #(
		.INIT('h1)
	) name871 (
		\a0_pad ,
		_w1043_,
		_w1044_
	);
	LUT2 #(
		.INIT('h2)
	) name872 (
		_w195_,
		_w1044_,
		_w1045_
	);
	LUT2 #(
		.INIT('h8)
	) name873 (
		\m5_pad ,
		\n5_pad ,
		_w1046_
	);
	LUT2 #(
		.INIT('h2)
	) name874 (
		_w175_,
		_w185_,
		_w1047_
	);
	LUT2 #(
		.INIT('h4)
	) name875 (
		_w389_,
		_w1047_,
		_w1048_
	);
	LUT2 #(
		.INIT('h1)
	) name876 (
		_w315_,
		_w1046_,
		_w1049_
	);
	LUT2 #(
		.INIT('h4)
	) name877 (
		_w1048_,
		_w1049_,
		_w1050_
	);
	LUT2 #(
		.INIT('h8)
	) name878 (
		_w457_,
		_w1050_,
		_w1051_
	);
	LUT2 #(
		.INIT('h4)
	) name879 (
		_w1045_,
		_w1051_,
		_w1052_
	);
	LUT2 #(
		.INIT('h1)
	) name880 (
		z_pad,
		_w1052_,
		_w1053_
	);
	LUT2 #(
		.INIT('h8)
	) name881 (
		p_pad,
		\z1_pad ,
		_w1054_
	);
	LUT2 #(
		.INIT('h8)
	) name882 (
		w_pad,
		\x0_pad ,
		_w1055_
	);
	LUT2 #(
		.INIT('h8)
	) name883 (
		\c1_pad ,
		v_pad,
		_w1056_
	);
	LUT2 #(
		.INIT('h8)
	) name884 (
		\d2_pad ,
		u_pad,
		_w1057_
	);
	LUT2 #(
		.INIT('h8)
	) name885 (
		r_pad,
		\t1_pad ,
		_w1058_
	);
	LUT2 #(
		.INIT('h8)
	) name886 (
		\i2_pad ,
		t_pad,
		_w1059_
	);
	LUT2 #(
		.INIT('h8)
	) name887 (
		n_pad,
		\z2_pad ,
		_w1060_
	);
	LUT2 #(
		.INIT('h8)
	) name888 (
		\d3_pad ,
		m_pad,
		_w1061_
	);
	LUT2 #(
		.INIT('h8)
	) name889 (
		q_pad,
		\w1_pad ,
		_w1062_
	);
	LUT2 #(
		.INIT('h8)
	) name890 (
		o_pad,
		\s2_pad ,
		_w1063_
	);
	LUT2 #(
		.INIT('h8)
	) name891 (
		\m2_pad ,
		s_pad,
		_w1064_
	);
	LUT2 #(
		.INIT('h1)
	) name892 (
		_w1054_,
		_w1055_,
		_w1065_
	);
	LUT2 #(
		.INIT('h1)
	) name893 (
		_w1056_,
		_w1057_,
		_w1066_
	);
	LUT2 #(
		.INIT('h1)
	) name894 (
		_w1058_,
		_w1059_,
		_w1067_
	);
	LUT2 #(
		.INIT('h1)
	) name895 (
		_w1060_,
		_w1061_,
		_w1068_
	);
	LUT2 #(
		.INIT('h1)
	) name896 (
		_w1062_,
		_w1063_,
		_w1069_
	);
	LUT2 #(
		.INIT('h4)
	) name897 (
		_w1064_,
		_w1069_,
		_w1070_
	);
	LUT2 #(
		.INIT('h8)
	) name898 (
		_w1067_,
		_w1068_,
		_w1071_
	);
	LUT2 #(
		.INIT('h8)
	) name899 (
		_w1065_,
		_w1066_,
		_w1072_
	);
	LUT2 #(
		.INIT('h8)
	) name900 (
		_w1071_,
		_w1072_,
		_w1073_
	);
	LUT2 #(
		.INIT('h8)
	) name901 (
		_w1070_,
		_w1073_,
		_w1074_
	);
	LUT2 #(
		.INIT('h2)
	) name902 (
		\r1_pad ,
		_w764_,
		_w1075_
	);
	LUT2 #(
		.INIT('h2)
	) name903 (
		\d1_pad ,
		_w1075_,
		_w1076_
	);
	LUT2 #(
		.INIT('h1)
	) name904 (
		c_pad,
		_w1076_,
		_w1077_
	);
	LUT2 #(
		.INIT('h2)
	) name905 (
		_w238_,
		_w1077_,
		_w1078_
	);
	LUT2 #(
		.INIT('h8)
	) name906 (
		\m1_pad ,
		\n1_pad ,
		_w1079_
	);
	LUT2 #(
		.INIT('h1)
	) name907 (
		\a3_pad ,
		\b3_pad ,
		_w1080_
	);
	LUT2 #(
		.INIT('h4)
	) name908 (
		\e3_pad ,
		\y2_pad ,
		_w1081_
	);
	LUT2 #(
		.INIT('h4)
	) name909 (
		\z2_pad ,
		_w1081_,
		_w1082_
	);
	LUT2 #(
		.INIT('h8)
	) name910 (
		_w833_,
		_w1080_,
		_w1083_
	);
	LUT2 #(
		.INIT('h8)
	) name911 (
		_w1082_,
		_w1083_,
		_w1084_
	);
	LUT2 #(
		.INIT('h8)
	) name912 (
		_w279_,
		_w1084_,
		_w1085_
	);
	LUT2 #(
		.INIT('h4)
	) name913 (
		b_pad,
		\n1_pad ,
		_w1086_
	);
	LUT2 #(
		.INIT('h8)
	) name914 (
		_w237_,
		_w1086_,
		_w1087_
	);
	LUT2 #(
		.INIT('h1)
	) name915 (
		_w1085_,
		_w1087_,
		_w1088_
	);
	LUT2 #(
		.INIT('h4)
	) name916 (
		_w247_,
		_w279_,
		_w1089_
	);
	LUT2 #(
		.INIT('h4)
	) name917 (
		_w1084_,
		_w1089_,
		_w1090_
	);
	LUT2 #(
		.INIT('h1)
	) name918 (
		_w276_,
		_w1079_,
		_w1091_
	);
	LUT2 #(
		.INIT('h8)
	) name919 (
		_w1088_,
		_w1091_,
		_w1092_
	);
	LUT2 #(
		.INIT('h4)
	) name920 (
		_w1090_,
		_w1092_,
		_w1093_
	);
	LUT2 #(
		.INIT('h4)
	) name921 (
		_w1078_,
		_w1093_,
		_w1094_
	);
	LUT2 #(
		.INIT('h1)
	) name922 (
		b_pad,
		_w1094_,
		_w1095_
	);
	LUT2 #(
		.INIT('h2)
	) name923 (
		\z1_pad ,
		_w826_,
		_w1096_
	);
	LUT2 #(
		.INIT('h1)
	) name924 (
		\m2_pad ,
		_w1020_,
		_w1097_
	);
	LUT2 #(
		.INIT('h8)
	) name925 (
		\m2_pad ,
		_w1020_,
		_w1098_
	);
	LUT2 #(
		.INIT('h2)
	) name926 (
		_w826_,
		_w1097_,
		_w1099_
	);
	LUT2 #(
		.INIT('h4)
	) name927 (
		_w1098_,
		_w1099_,
		_w1100_
	);
	LUT2 #(
		.INIT('h1)
	) name928 (
		b_pad,
		_w1096_,
		_w1101_
	);
	LUT2 #(
		.INIT('h4)
	) name929 (
		_w1100_,
		_w1101_,
		_w1102_
	);
	LUT2 #(
		.INIT('h1)
	) name930 (
		\l3_pad ,
		_w313_,
		_w1103_
	);
	LUT2 #(
		.INIT('h8)
	) name931 (
		\l3_pad ,
		_w313_,
		_w1104_
	);
	LUT2 #(
		.INIT('h1)
	) name932 (
		_w1103_,
		_w1104_,
		_w1105_
	);
	LUT2 #(
		.INIT('h8)
	) name933 (
		_w1028_,
		_w1105_,
		_w1106_
	);
	LUT2 #(
		.INIT('h1)
	) name934 (
		\m3_pad ,
		_w1106_,
		_w1107_
	);
	LUT2 #(
		.INIT('h8)
	) name935 (
		\m3_pad ,
		_w1106_,
		_w1108_
	);
	LUT2 #(
		.INIT('h2)
	) name936 (
		_w316_,
		_w1107_,
		_w1109_
	);
	LUT2 #(
		.INIT('h4)
	) name937 (
		_w1108_,
		_w1109_,
		_w1110_
	);
	LUT2 #(
		.INIT('h2)
	) name938 (
		\z3_pad ,
		_w887_,
		_w1111_
	);
	LUT2 #(
		.INIT('h1)
	) name939 (
		\j0_pad ,
		_w1037_,
		_w1112_
	);
	LUT2 #(
		.INIT('h2)
	) name940 (
		\m4_pad ,
		_w1112_,
		_w1113_
	);
	LUT2 #(
		.INIT('h4)
	) name941 (
		\m4_pad ,
		_w1112_,
		_w1114_
	);
	LUT2 #(
		.INIT('h2)
	) name942 (
		_w887_,
		_w1113_,
		_w1115_
	);
	LUT2 #(
		.INIT('h4)
	) name943 (
		_w1114_,
		_w1115_,
		_w1116_
	);
	LUT2 #(
		.INIT('h1)
	) name944 (
		z_pad,
		_w1111_,
		_w1117_
	);
	LUT2 #(
		.INIT('h4)
	) name945 (
		_w1116_,
		_w1117_,
		_w1118_
	);
	LUT2 #(
		.INIT('h8)
	) name946 (
		p_pad,
		\y1_pad ,
		_w1119_
	);
	LUT2 #(
		.INIT('h8)
	) name947 (
		\w0_pad ,
		w_pad,
		_w1120_
	);
	LUT2 #(
		.INIT('h8)
	) name948 (
		\b1_pad ,
		v_pad,
		_w1121_
	);
	LUT2 #(
		.INIT('h8)
	) name949 (
		\c2_pad ,
		u_pad,
		_w1122_
	);
	LUT2 #(
		.INIT('h8)
	) name950 (
		r_pad,
		\s1_pad ,
		_w1123_
	);
	LUT2 #(
		.INIT('h8)
	) name951 (
		\h2_pad ,
		t_pad,
		_w1124_
	);
	LUT2 #(
		.INIT('h8)
	) name952 (
		n_pad,
		\y2_pad ,
		_w1125_
	);
	LUT2 #(
		.INIT('h8)
	) name953 (
		\c3_pad ,
		m_pad,
		_w1126_
	);
	LUT2 #(
		.INIT('h8)
	) name954 (
		q_pad,
		\v1_pad ,
		_w1127_
	);
	LUT2 #(
		.INIT('h8)
	) name955 (
		o_pad,
		\r2_pad ,
		_w1128_
	);
	LUT2 #(
		.INIT('h8)
	) name956 (
		\l2_pad ,
		s_pad,
		_w1129_
	);
	LUT2 #(
		.INIT('h1)
	) name957 (
		_w1119_,
		_w1120_,
		_w1130_
	);
	LUT2 #(
		.INIT('h1)
	) name958 (
		_w1121_,
		_w1122_,
		_w1131_
	);
	LUT2 #(
		.INIT('h1)
	) name959 (
		_w1123_,
		_w1124_,
		_w1132_
	);
	LUT2 #(
		.INIT('h1)
	) name960 (
		_w1125_,
		_w1126_,
		_w1133_
	);
	LUT2 #(
		.INIT('h1)
	) name961 (
		_w1127_,
		_w1128_,
		_w1134_
	);
	LUT2 #(
		.INIT('h4)
	) name962 (
		_w1129_,
		_w1134_,
		_w1135_
	);
	LUT2 #(
		.INIT('h8)
	) name963 (
		_w1132_,
		_w1133_,
		_w1136_
	);
	LUT2 #(
		.INIT('h8)
	) name964 (
		_w1130_,
		_w1131_,
		_w1137_
	);
	LUT2 #(
		.INIT('h8)
	) name965 (
		_w1136_,
		_w1137_,
		_w1138_
	);
	LUT2 #(
		.INIT('h8)
	) name966 (
		_w1135_,
		_w1138_,
		_w1139_
	);
	LUT2 #(
		.INIT('h1)
	) name967 (
		b_pad,
		_w826_,
		_w1140_
	);
	LUT2 #(
		.INIT('h8)
	) name968 (
		\k2_pad ,
		\l2_pad ,
		_w1141_
	);
	LUT2 #(
		.INIT('h8)
	) name969 (
		\m2_pad ,
		\o2_pad ,
		_w1142_
	);
	LUT2 #(
		.INIT('h8)
	) name970 (
		_w1141_,
		_w1142_,
		_w1143_
	);
	LUT2 #(
		.INIT('h8)
	) name971 (
		_w955_,
		_w1143_,
		_w1144_
	);
	LUT2 #(
		.INIT('h4)
	) name972 (
		_w1140_,
		_w1144_,
		_w1145_
	);
	LUT2 #(
		.INIT('h1)
	) name973 (
		\m3_pad ,
		_w313_,
		_w1146_
	);
	LUT2 #(
		.INIT('h8)
	) name974 (
		\m3_pad ,
		_w313_,
		_w1147_
	);
	LUT2 #(
		.INIT('h1)
	) name975 (
		_w1146_,
		_w1147_,
		_w1148_
	);
	LUT2 #(
		.INIT('h8)
	) name976 (
		_w1106_,
		_w1148_,
		_w1149_
	);
	LUT2 #(
		.INIT('h1)
	) name977 (
		\n3_pad ,
		_w1149_,
		_w1150_
	);
	LUT2 #(
		.INIT('h8)
	) name978 (
		\n3_pad ,
		_w1149_,
		_w1151_
	);
	LUT2 #(
		.INIT('h2)
	) name979 (
		_w316_,
		_w1150_,
		_w1152_
	);
	LUT2 #(
		.INIT('h4)
	) name980 (
		_w1151_,
		_w1152_,
		_w1153_
	);
	LUT2 #(
		.INIT('h2)
	) name981 (
		\a4_pad ,
		_w887_,
		_w1154_
	);
	LUT2 #(
		.INIT('h1)
	) name982 (
		\n4_pad ,
		_w1113_,
		_w1155_
	);
	LUT2 #(
		.INIT('h8)
	) name983 (
		\n4_pad ,
		_w1113_,
		_w1156_
	);
	LUT2 #(
		.INIT('h2)
	) name984 (
		_w887_,
		_w1155_,
		_w1157_
	);
	LUT2 #(
		.INIT('h4)
	) name985 (
		_w1156_,
		_w1157_,
		_w1158_
	);
	LUT2 #(
		.INIT('h1)
	) name986 (
		z_pad,
		_w1154_,
		_w1159_
	);
	LUT2 #(
		.INIT('h4)
	) name987 (
		_w1158_,
		_w1159_,
		_w1160_
	);
	LUT2 #(
		.INIT('h8)
	) name988 (
		\p1_pad ,
		p_pad,
		_w1161_
	);
	LUT2 #(
		.INIT('h8)
	) name989 (
		\v0_pad ,
		w_pad,
		_w1162_
	);
	LUT2 #(
		.INIT('h8)
	) name990 (
		\a1_pad ,
		v_pad,
		_w1163_
	);
	LUT2 #(
		.INIT('h8)
	) name991 (
		\b2_pad ,
		u_pad,
		_w1164_
	);
	LUT2 #(
		.INIT('h8)
	) name992 (
		q_pad,
		\r1_pad ,
		_w1165_
	);
	LUT2 #(
		.INIT('h8)
	) name993 (
		\f2_pad ,
		t_pad,
		_w1166_
	);
	LUT2 #(
		.INIT('h8)
	) name994 (
		n_pad,
		\x2_pad ,
		_w1167_
	);
	LUT2 #(
		.INIT('h8)
	) name995 (
		\b3_pad ,
		m_pad,
		_w1168_
	);
	LUT2 #(
		.INIT('h8)
	) name996 (
		\m1_pad ,
		r_pad,
		_w1169_
	);
	LUT2 #(
		.INIT('h8)
	) name997 (
		o_pad,
		\q2_pad ,
		_w1170_
	);
	LUT2 #(
		.INIT('h8)
	) name998 (
		\k2_pad ,
		s_pad,
		_w1171_
	);
	LUT2 #(
		.INIT('h1)
	) name999 (
		_w1161_,
		_w1162_,
		_w1172_
	);
	LUT2 #(
		.INIT('h1)
	) name1000 (
		_w1163_,
		_w1164_,
		_w1173_
	);
	LUT2 #(
		.INIT('h1)
	) name1001 (
		_w1165_,
		_w1166_,
		_w1174_
	);
	LUT2 #(
		.INIT('h1)
	) name1002 (
		_w1167_,
		_w1168_,
		_w1175_
	);
	LUT2 #(
		.INIT('h1)
	) name1003 (
		_w1169_,
		_w1170_,
		_w1176_
	);
	LUT2 #(
		.INIT('h4)
	) name1004 (
		_w1171_,
		_w1176_,
		_w1177_
	);
	LUT2 #(
		.INIT('h8)
	) name1005 (
		_w1174_,
		_w1175_,
		_w1178_
	);
	LUT2 #(
		.INIT('h8)
	) name1006 (
		_w1172_,
		_w1173_,
		_w1179_
	);
	LUT2 #(
		.INIT('h8)
	) name1007 (
		_w1178_,
		_w1179_,
		_w1180_
	);
	LUT2 #(
		.INIT('h8)
	) name1008 (
		_w1177_,
		_w1180_,
		_w1181_
	);
	LUT2 #(
		.INIT('h2)
	) name1009 (
		\a2_pad ,
		_w826_,
		_w1182_
	);
	LUT2 #(
		.INIT('h4)
	) name1010 (
		_w979_,
		_w1143_,
		_w1183_
	);
	LUT2 #(
		.INIT('h1)
	) name1011 (
		\o2_pad ,
		_w1098_,
		_w1184_
	);
	LUT2 #(
		.INIT('h2)
	) name1012 (
		_w826_,
		_w1183_,
		_w1185_
	);
	LUT2 #(
		.INIT('h4)
	) name1013 (
		_w1184_,
		_w1185_,
		_w1186_
	);
	LUT2 #(
		.INIT('h1)
	) name1014 (
		b_pad,
		_w1182_,
		_w1187_
	);
	LUT2 #(
		.INIT('h4)
	) name1015 (
		_w1186_,
		_w1187_,
		_w1188_
	);
	LUT2 #(
		.INIT('h1)
	) name1016 (
		\n3_pad ,
		_w313_,
		_w1189_
	);
	LUT2 #(
		.INIT('h8)
	) name1017 (
		\n3_pad ,
		_w313_,
		_w1190_
	);
	LUT2 #(
		.INIT('h1)
	) name1018 (
		_w1189_,
		_w1190_,
		_w1191_
	);
	LUT2 #(
		.INIT('h8)
	) name1019 (
		_w1149_,
		_w1191_,
		_w1192_
	);
	LUT2 #(
		.INIT('h1)
	) name1020 (
		\o3_pad ,
		_w1192_,
		_w1193_
	);
	LUT2 #(
		.INIT('h8)
	) name1021 (
		\o3_pad ,
		_w1192_,
		_w1194_
	);
	LUT2 #(
		.INIT('h2)
	) name1022 (
		_w316_,
		_w1193_,
		_w1195_
	);
	LUT2 #(
		.INIT('h4)
	) name1023 (
		_w1194_,
		_w1195_,
		_w1196_
	);
	LUT2 #(
		.INIT('h1)
	) name1024 (
		_w317_,
		_w1196_,
		_w1197_
	);
	LUT2 #(
		.INIT('h2)
	) name1025 (
		\b4_pad ,
		_w887_,
		_w1198_
	);
	LUT2 #(
		.INIT('h1)
	) name1026 (
		\o4_pad ,
		_w1156_,
		_w1199_
	);
	LUT2 #(
		.INIT('h8)
	) name1027 (
		\o4_pad ,
		_w1156_,
		_w1200_
	);
	LUT2 #(
		.INIT('h2)
	) name1028 (
		_w887_,
		_w1199_,
		_w1201_
	);
	LUT2 #(
		.INIT('h4)
	) name1029 (
		_w1200_,
		_w1201_,
		_w1202_
	);
	LUT2 #(
		.INIT('h1)
	) name1030 (
		z_pad,
		_w1198_,
		_w1203_
	);
	LUT2 #(
		.INIT('h4)
	) name1031 (
		_w1202_,
		_w1203_,
		_w1204_
	);
	LUT2 #(
		.INIT('h1)
	) name1032 (
		\c0_pad ,
		_w460_,
		_w1205_
	);
	LUT2 #(
		.INIT('h2)
	) name1033 (
		\r5_pad ,
		_w1205_,
		_w1206_
	);
	LUT2 #(
		.INIT('h1)
	) name1034 (
		\b0_pad ,
		_w455_,
		_w1207_
	);
	LUT2 #(
		.INIT('h2)
	) name1035 (
		\q5_pad ,
		_w1207_,
		_w1208_
	);
	LUT2 #(
		.INIT('h8)
	) name1036 (
		\p5_pad ,
		\q5_pad ,
		_w1209_
	);
	LUT2 #(
		.INIT('h1)
	) name1037 (
		\p5_pad ,
		\q5_pad ,
		_w1210_
	);
	LUT2 #(
		.INIT('h1)
	) name1038 (
		\r5_pad ,
		_w1210_,
		_w1211_
	);
	LUT2 #(
		.INIT('h8)
	) name1039 (
		\r5_pad ,
		_w1210_,
		_w1212_
	);
	LUT2 #(
		.INIT('h1)
	) name1040 (
		_w1211_,
		_w1212_,
		_w1213_
	);
	LUT2 #(
		.INIT('h1)
	) name1041 (
		z_pad,
		_w1209_,
		_w1214_
	);
	LUT2 #(
		.INIT('h4)
	) name1042 (
		_w1213_,
		_w1214_,
		_w1215_
	);
	LUT2 #(
		.INIT('h8)
	) name1043 (
		\p5_pad ,
		_w1205_,
		_w1216_
	);
	LUT2 #(
		.INIT('h8)
	) name1044 (
		_w1207_,
		_w1216_,
		_w1217_
	);
	LUT2 #(
		.INIT('h1)
	) name1045 (
		_w1206_,
		_w1208_,
		_w1218_
	);
	LUT2 #(
		.INIT('h8)
	) name1046 (
		_w1215_,
		_w1218_,
		_w1219_
	);
	LUT2 #(
		.INIT('h4)
	) name1047 (
		_w1217_,
		_w1219_,
		_w1220_
	);
	LUT2 #(
		.INIT('h8)
	) name1048 (
		p_pad,
		\q1_pad ,
		_w1221_
	);
	LUT2 #(
		.INIT('h8)
	) name1049 (
		\e2_pad ,
		t_pad,
		_w1222_
	);
	LUT2 #(
		.INIT('h8)
	) name1050 (
		\l1_pad ,
		w_pad,
		_w1223_
	);
	LUT2 #(
		.INIT('h8)
	) name1051 (
		v_pad,
		\z0_pad ,
		_w1224_
	);
	LUT2 #(
		.INIT('h8)
	) name1052 (
		n_pad,
		\w2_pad ,
		_w1225_
	);
	LUT2 #(
		.INIT('h2)
	) name1053 (
		q_pad,
		_w277_,
		_w1226_
	);
	LUT2 #(
		.INIT('h8)
	) name1054 (
		\n1_pad ,
		r_pad,
		_w1227_
	);
	LUT2 #(
		.INIT('h8)
	) name1055 (
		u_pad,
		_w303_,
		_w1228_
	);
	LUT2 #(
		.INIT('h8)
	) name1056 (
		s_pad,
		_w825_,
		_w1229_
	);
	LUT2 #(
		.INIT('h8)
	) name1057 (
		m_pad,
		_w1084_,
		_w1230_
	);
	LUT2 #(
		.INIT('h8)
	) name1058 (
		o_pad,
		_w604_,
		_w1231_
	);
	LUT2 #(
		.INIT('h1)
	) name1059 (
		_w1221_,
		_w1222_,
		_w1232_
	);
	LUT2 #(
		.INIT('h1)
	) name1060 (
		_w1223_,
		_w1224_,
		_w1233_
	);
	LUT2 #(
		.INIT('h1)
	) name1061 (
		_w1225_,
		_w1227_,
		_w1234_
	);
	LUT2 #(
		.INIT('h8)
	) name1062 (
		_w1233_,
		_w1234_,
		_w1235_
	);
	LUT2 #(
		.INIT('h8)
	) name1063 (
		_w1232_,
		_w1235_,
		_w1236_
	);
	LUT2 #(
		.INIT('h4)
	) name1064 (
		_w1231_,
		_w1236_,
		_w1237_
	);
	LUT2 #(
		.INIT('h4)
	) name1065 (
		_w1230_,
		_w1237_,
		_w1238_
	);
	LUT2 #(
		.INIT('h4)
	) name1066 (
		_w1226_,
		_w1238_,
		_w1239_
	);
	LUT2 #(
		.INIT('h4)
	) name1067 (
		_w1229_,
		_w1239_,
		_w1240_
	);
	LUT2 #(
		.INIT('h4)
	) name1068 (
		_w1228_,
		_w1240_,
		_w1241_
	);
	LUT2 #(
		.INIT('h8)
	) name1069 (
		_w227_,
		_w1079_,
		_w1242_
	);
	LUT2 #(
		.INIT('h1)
	) name1070 (
		e_pad,
		_w1242_,
		_w1243_
	);
	LUT2 #(
		.INIT('h2)
	) name1071 (
		\r1_pad ,
		_w1243_,
		_w1244_
	);
	LUT2 #(
		.INIT('h1)
	) name1072 (
		d_pad,
		_w1087_,
		_w1245_
	);
	LUT2 #(
		.INIT('h2)
	) name1073 (
		\q1_pad ,
		_w1245_,
		_w1246_
	);
	LUT2 #(
		.INIT('h8)
	) name1074 (
		\p1_pad ,
		\q1_pad ,
		_w1247_
	);
	LUT2 #(
		.INIT('h1)
	) name1075 (
		\p1_pad ,
		\q1_pad ,
		_w1248_
	);
	LUT2 #(
		.INIT('h1)
	) name1076 (
		\r1_pad ,
		_w1248_,
		_w1249_
	);
	LUT2 #(
		.INIT('h8)
	) name1077 (
		\r1_pad ,
		_w1248_,
		_w1250_
	);
	LUT2 #(
		.INIT('h1)
	) name1078 (
		_w1249_,
		_w1250_,
		_w1251_
	);
	LUT2 #(
		.INIT('h1)
	) name1079 (
		b_pad,
		_w1247_,
		_w1252_
	);
	LUT2 #(
		.INIT('h4)
	) name1080 (
		_w1251_,
		_w1252_,
		_w1253_
	);
	LUT2 #(
		.INIT('h8)
	) name1081 (
		\p1_pad ,
		_w1243_,
		_w1254_
	);
	LUT2 #(
		.INIT('h8)
	) name1082 (
		_w1245_,
		_w1254_,
		_w1255_
	);
	LUT2 #(
		.INIT('h1)
	) name1083 (
		_w1244_,
		_w1246_,
		_w1256_
	);
	LUT2 #(
		.INIT('h8)
	) name1084 (
		_w1253_,
		_w1256_,
		_w1257_
	);
	LUT2 #(
		.INIT('h4)
	) name1085 (
		_w1255_,
		_w1257_,
		_w1258_
	);
	LUT2 #(
		.INIT('h2)
	) name1086 (
		\p2_pad ,
		_w947_,
		_w1259_
	);
	LUT2 #(
		.INIT('h4)
	) name1087 (
		\l6_pad ,
		_w947_,
		_w1260_
	);
	LUT2 #(
		.INIT('h1)
	) name1088 (
		_w1259_,
		_w1260_,
		_w1261_
	);
	LUT2 #(
		.INIT('h1)
	) name1089 (
		_w313_,
		_w357_,
		_w1262_
	);
	LUT2 #(
		.INIT('h2)
	) name1090 (
		_w313_,
		_w328_,
		_w1263_
	);
	LUT2 #(
		.INIT('h1)
	) name1091 (
		_w350_,
		_w1262_,
		_w1264_
	);
	LUT2 #(
		.INIT('h4)
	) name1092 (
		_w1263_,
		_w1264_,
		_w1265_
	);
	LUT2 #(
		.INIT('h1)
	) name1093 (
		\p3_pad ,
		_w1265_,
		_w1266_
	);
	LUT2 #(
		.INIT('h8)
	) name1094 (
		\p3_pad ,
		_w1265_,
		_w1267_
	);
	LUT2 #(
		.INIT('h2)
	) name1095 (
		_w316_,
		_w1266_,
		_w1268_
	);
	LUT2 #(
		.INIT('h4)
	) name1096 (
		_w1267_,
		_w1268_,
		_w1269_
	);
	LUT2 #(
		.INIT('h1)
	) name1097 (
		_w317_,
		_w1269_,
		_w1270_
	);
	LUT2 #(
		.INIT('h1)
	) name1098 (
		z_pad,
		_w887_,
		_w1271_
	);
	LUT2 #(
		.INIT('h8)
	) name1099 (
		\m4_pad ,
		\n4_pad ,
		_w1272_
	);
	LUT2 #(
		.INIT('h8)
	) name1100 (
		\o4_pad ,
		\q4_pad ,
		_w1273_
	);
	LUT2 #(
		.INIT('h8)
	) name1101 (
		_w1272_,
		_w1273_,
		_w1274_
	);
	LUT2 #(
		.INIT('h8)
	) name1102 (
		_w1036_,
		_w1274_,
		_w1275_
	);
	LUT2 #(
		.INIT('h4)
	) name1103 (
		_w1271_,
		_w1275_,
		_w1276_
	);
	LUT2 #(
		.INIT('h2)
	) name1104 (
		\r5_pad ,
		_w1207_,
		_w1277_
	);
	LUT2 #(
		.INIT('h2)
	) name1105 (
		\p5_pad ,
		_w1205_,
		_w1278_
	);
	LUT2 #(
		.INIT('h8)
	) name1106 (
		\q5_pad ,
		_w1205_,
		_w1279_
	);
	LUT2 #(
		.INIT('h8)
	) name1107 (
		_w1207_,
		_w1279_,
		_w1280_
	);
	LUT2 #(
		.INIT('h1)
	) name1108 (
		_w1277_,
		_w1278_,
		_w1281_
	);
	LUT2 #(
		.INIT('h4)
	) name1109 (
		_w1280_,
		_w1281_,
		_w1282_
	);
	LUT2 #(
		.INIT('h2)
	) name1110 (
		_w1215_,
		_w1282_,
		_w1283_
	);
	LUT2 #(
		.INIT('h8)
	) name1111 (
		_w279_,
		_w605_,
		_w1284_
	);
	LUT2 #(
		.INIT('h1)
	) name1112 (
		_w229_,
		_w1242_,
		_w1285_
	);
	LUT2 #(
		.INIT('h4)
	) name1113 (
		_w1284_,
		_w1285_,
		_w1286_
	);
	LUT2 #(
		.INIT('h8)
	) name1114 (
		_w1088_,
		_w1286_,
		_w1287_
	);
	LUT2 #(
		.INIT('h8)
	) name1115 (
		\c4_pad ,
		\n0_pad ,
		_w1288_
	);
	LUT2 #(
		.INIT('h8)
	) name1116 (
		\u0_pad ,
		\u4_pad ,
		_w1289_
	);
	LUT2 #(
		.INIT('h8)
	) name1117 (
		\t0_pad ,
		\z4_pad ,
		_w1290_
	);
	LUT2 #(
		.INIT('h8)
	) name1118 (
		\i4_pad ,
		\s0_pad ,
		_w1291_
	);
	LUT2 #(
		.INIT('h8)
	) name1119 (
		\o0_pad ,
		\z3_pad ,
		_w1292_
	);
	LUT2 #(
		.INIT('h8)
	) name1120 (
		\l4_pad ,
		\r0_pad ,
		_w1293_
	);
	LUT2 #(
		.INIT('h8)
	) name1121 (
		\k0_pad ,
		\t3_pad ,
		_w1294_
	);
	LUT2 #(
		.INIT('h8)
	) name1122 (
		\l0_pad ,
		\p3_pad ,
		_w1295_
	);
	LUT2 #(
		.INIT('h8)
	) name1123 (
		\p0_pad ,
		\w3_pad ,
		_w1296_
	);
	LUT2 #(
		.INIT('h8)
	) name1124 (
		\i3_pad ,
		\m0_pad ,
		_w1297_
	);
	LUT2 #(
		.INIT('h8)
	) name1125 (
		\q0_pad ,
		\q4_pad ,
		_w1298_
	);
	LUT2 #(
		.INIT('h1)
	) name1126 (
		_w1288_,
		_w1289_,
		_w1299_
	);
	LUT2 #(
		.INIT('h1)
	) name1127 (
		_w1290_,
		_w1291_,
		_w1300_
	);
	LUT2 #(
		.INIT('h1)
	) name1128 (
		_w1292_,
		_w1293_,
		_w1301_
	);
	LUT2 #(
		.INIT('h1)
	) name1129 (
		_w1294_,
		_w1295_,
		_w1302_
	);
	LUT2 #(
		.INIT('h1)
	) name1130 (
		_w1296_,
		_w1297_,
		_w1303_
	);
	LUT2 #(
		.INIT('h4)
	) name1131 (
		_w1298_,
		_w1303_,
		_w1304_
	);
	LUT2 #(
		.INIT('h8)
	) name1132 (
		_w1301_,
		_w1302_,
		_w1305_
	);
	LUT2 #(
		.INIT('h8)
	) name1133 (
		_w1299_,
		_w1300_,
		_w1306_
	);
	LUT2 #(
		.INIT('h8)
	) name1134 (
		_w1305_,
		_w1306_,
		_w1307_
	);
	LUT2 #(
		.INIT('h8)
	) name1135 (
		_w1304_,
		_w1307_,
		_w1308_
	);
	LUT2 #(
		.INIT('h2)
	) name1136 (
		\r1_pad ,
		_w1245_,
		_w1309_
	);
	LUT2 #(
		.INIT('h2)
	) name1137 (
		\p1_pad ,
		_w1243_,
		_w1310_
	);
	LUT2 #(
		.INIT('h8)
	) name1138 (
		\q1_pad ,
		_w1243_,
		_w1311_
	);
	LUT2 #(
		.INIT('h8)
	) name1139 (
		_w1245_,
		_w1311_,
		_w1312_
	);
	LUT2 #(
		.INIT('h1)
	) name1140 (
		_w1309_,
		_w1310_,
		_w1313_
	);
	LUT2 #(
		.INIT('h4)
	) name1141 (
		_w1312_,
		_w1313_,
		_w1314_
	);
	LUT2 #(
		.INIT('h2)
	) name1142 (
		_w1253_,
		_w1314_,
		_w1315_
	);
	LUT2 #(
		.INIT('h2)
	) name1143 (
		\q2_pad ,
		_w303_,
		_w1316_
	);
	LUT2 #(
		.INIT('h4)
	) name1144 (
		\q2_pad ,
		_w303_,
		_w1317_
	);
	LUT2 #(
		.INIT('h2)
	) name1145 (
		_w277_,
		_w1316_,
		_w1318_
	);
	LUT2 #(
		.INIT('h4)
	) name1146 (
		_w1317_,
		_w1318_,
		_w1319_
	);
	LUT2 #(
		.INIT('h8)
	) name1147 (
		_w313_,
		_w330_,
		_w1320_
	);
	LUT2 #(
		.INIT('h2)
	) name1148 (
		_w361_,
		_w1320_,
		_w1321_
	);
	LUT2 #(
		.INIT('h1)
	) name1149 (
		\q3_pad ,
		_w1321_,
		_w1322_
	);
	LUT2 #(
		.INIT('h8)
	) name1150 (
		\q3_pad ,
		_w1321_,
		_w1323_
	);
	LUT2 #(
		.INIT('h2)
	) name1151 (
		_w316_,
		_w1322_,
		_w1324_
	);
	LUT2 #(
		.INIT('h4)
	) name1152 (
		_w1323_,
		_w1324_,
		_w1325_
	);
	LUT2 #(
		.INIT('h1)
	) name1153 (
		_w317_,
		_w1325_,
		_w1326_
	);
	LUT2 #(
		.INIT('h2)
	) name1154 (
		\c4_pad ,
		_w887_,
		_w1327_
	);
	LUT2 #(
		.INIT('h4)
	) name1155 (
		_w1112_,
		_w1274_,
		_w1328_
	);
	LUT2 #(
		.INIT('h1)
	) name1156 (
		\q4_pad ,
		_w1200_,
		_w1329_
	);
	LUT2 #(
		.INIT('h2)
	) name1157 (
		_w887_,
		_w1328_,
		_w1330_
	);
	LUT2 #(
		.INIT('h4)
	) name1158 (
		_w1329_,
		_w1330_,
		_w1331_
	);
	LUT2 #(
		.INIT('h1)
	) name1159 (
		z_pad,
		_w1327_,
		_w1332_
	);
	LUT2 #(
		.INIT('h4)
	) name1160 (
		_w1331_,
		_w1332_,
		_w1333_
	);
	LUT2 #(
		.INIT('h2)
	) name1161 (
		\p5_pad ,
		_w1207_,
		_w1334_
	);
	LUT2 #(
		.INIT('h2)
	) name1162 (
		\q5_pad ,
		_w1205_,
		_w1335_
	);
	LUT2 #(
		.INIT('h8)
	) name1163 (
		\r5_pad ,
		_w1205_,
		_w1336_
	);
	LUT2 #(
		.INIT('h8)
	) name1164 (
		_w1207_,
		_w1336_,
		_w1337_
	);
	LUT2 #(
		.INIT('h1)
	) name1165 (
		_w1334_,
		_w1335_,
		_w1338_
	);
	LUT2 #(
		.INIT('h4)
	) name1166 (
		_w1337_,
		_w1338_,
		_w1339_
	);
	LUT2 #(
		.INIT('h2)
	) name1167 (
		_w1215_,
		_w1339_,
		_w1340_
	);
	LUT2 #(
		.INIT('h8)
	) name1168 (
		\b4_pad ,
		\n0_pad ,
		_w1341_
	);
	LUT2 #(
		.INIT('h8)
	) name1169 (
		\t4_pad ,
		\u0_pad ,
		_w1342_
	);
	LUT2 #(
		.INIT('h8)
	) name1170 (
		\t0_pad ,
		\y4_pad ,
		_w1343_
	);
	LUT2 #(
		.INIT('h8)
	) name1171 (
		\f4_pad ,
		\s0_pad ,
		_w1344_
	);
	LUT2 #(
		.INIT('h8)
	) name1172 (
		\o0_pad ,
		\y3_pad ,
		_w1345_
	);
	LUT2 #(
		.INIT('h8)
	) name1173 (
		\k4_pad ,
		\r0_pad ,
		_w1346_
	);
	LUT2 #(
		.INIT('h8)
	) name1174 (
		\k0_pad ,
		\s3_pad ,
		_w1347_
	);
	LUT2 #(
		.INIT('h8)
	) name1175 (
		\l0_pad ,
		\o3_pad ,
		_w1348_
	);
	LUT2 #(
		.INIT('h8)
	) name1176 (
		\p0_pad ,
		\v3_pad ,
		_w1349_
	);
	LUT2 #(
		.INIT('h8)
	) name1177 (
		\h3_pad ,
		\m0_pad ,
		_w1350_
	);
	LUT2 #(
		.INIT('h8)
	) name1178 (
		\o4_pad ,
		\q0_pad ,
		_w1351_
	);
	LUT2 #(
		.INIT('h1)
	) name1179 (
		_w1341_,
		_w1342_,
		_w1352_
	);
	LUT2 #(
		.INIT('h1)
	) name1180 (
		_w1343_,
		_w1344_,
		_w1353_
	);
	LUT2 #(
		.INIT('h1)
	) name1181 (
		_w1345_,
		_w1346_,
		_w1354_
	);
	LUT2 #(
		.INIT('h1)
	) name1182 (
		_w1347_,
		_w1348_,
		_w1355_
	);
	LUT2 #(
		.INIT('h1)
	) name1183 (
		_w1349_,
		_w1350_,
		_w1356_
	);
	LUT2 #(
		.INIT('h4)
	) name1184 (
		_w1351_,
		_w1356_,
		_w1357_
	);
	LUT2 #(
		.INIT('h8)
	) name1185 (
		_w1354_,
		_w1355_,
		_w1358_
	);
	LUT2 #(
		.INIT('h8)
	) name1186 (
		_w1352_,
		_w1353_,
		_w1359_
	);
	LUT2 #(
		.INIT('h8)
	) name1187 (
		_w1358_,
		_w1359_,
		_w1360_
	);
	LUT2 #(
		.INIT('h8)
	) name1188 (
		_w1357_,
		_w1360_,
		_w1361_
	);
	LUT2 #(
		.INIT('h2)
	) name1189 (
		\p1_pad ,
		_w1245_,
		_w1362_
	);
	LUT2 #(
		.INIT('h2)
	) name1190 (
		\q1_pad ,
		_w1243_,
		_w1363_
	);
	LUT2 #(
		.INIT('h8)
	) name1191 (
		\r1_pad ,
		_w1243_,
		_w1364_
	);
	LUT2 #(
		.INIT('h8)
	) name1192 (
		_w1245_,
		_w1364_,
		_w1365_
	);
	LUT2 #(
		.INIT('h1)
	) name1193 (
		_w1362_,
		_w1363_,
		_w1366_
	);
	LUT2 #(
		.INIT('h4)
	) name1194 (
		_w1365_,
		_w1366_,
		_w1367_
	);
	LUT2 #(
		.INIT('h2)
	) name1195 (
		_w1253_,
		_w1367_,
		_w1368_
	);
	LUT2 #(
		.INIT('h1)
	) name1196 (
		\q2_pad ,
		_w273_,
		_w1369_
	);
	LUT2 #(
		.INIT('h8)
	) name1197 (
		\q2_pad ,
		_w273_,
		_w1370_
	);
	LUT2 #(
		.INIT('h1)
	) name1198 (
		_w303_,
		_w1369_,
		_w1371_
	);
	LUT2 #(
		.INIT('h4)
	) name1199 (
		_w1370_,
		_w1371_,
		_w1372_
	);
	LUT2 #(
		.INIT('h8)
	) name1200 (
		\r2_pad ,
		_w1372_,
		_w1373_
	);
	LUT2 #(
		.INIT('h1)
	) name1201 (
		\r2_pad ,
		_w1372_,
		_w1374_
	);
	LUT2 #(
		.INIT('h2)
	) name1202 (
		_w277_,
		_w1373_,
		_w1375_
	);
	LUT2 #(
		.INIT('h4)
	) name1203 (
		_w1374_,
		_w1375_,
		_w1376_
	);
	LUT2 #(
		.INIT('h1)
	) name1204 (
		\q3_pad ,
		_w313_,
		_w1377_
	);
	LUT2 #(
		.INIT('h2)
	) name1205 (
		_w313_,
		_w331_,
		_w1378_
	);
	LUT2 #(
		.INIT('h2)
	) name1206 (
		_w361_,
		_w1377_,
		_w1379_
	);
	LUT2 #(
		.INIT('h4)
	) name1207 (
		_w1378_,
		_w1379_,
		_w1380_
	);
	LUT2 #(
		.INIT('h8)
	) name1208 (
		\r3_pad ,
		_w1380_,
		_w1381_
	);
	LUT2 #(
		.INIT('h1)
	) name1209 (
		\r3_pad ,
		_w1380_,
		_w1382_
	);
	LUT2 #(
		.INIT('h2)
	) name1210 (
		_w316_,
		_w1381_,
		_w1383_
	);
	LUT2 #(
		.INIT('h4)
	) name1211 (
		_w1382_,
		_w1383_,
		_w1384_
	);
	LUT2 #(
		.INIT('h4)
	) name1212 (
		\r4_pad ,
		_w199_,
		_w1385_
	);
	LUT2 #(
		.INIT('h2)
	) name1213 (
		_w197_,
		_w200_,
		_w1386_
	);
	LUT2 #(
		.INIT('h4)
	) name1214 (
		_w1385_,
		_w1386_,
		_w1387_
	);
	LUT2 #(
		.INIT('h8)
	) name1215 (
		\a4_pad ,
		\n0_pad ,
		_w1388_
	);
	LUT2 #(
		.INIT('h8)
	) name1216 (
		\s4_pad ,
		\u0_pad ,
		_w1389_
	);
	LUT2 #(
		.INIT('h8)
	) name1217 (
		\t0_pad ,
		\x4_pad ,
		_w1390_
	);
	LUT2 #(
		.INIT('h8)
	) name1218 (
		\e4_pad ,
		\s0_pad ,
		_w1391_
	);
	LUT2 #(
		.INIT('h8)
	) name1219 (
		\o0_pad ,
		\x3_pad ,
		_w1392_
	);
	LUT2 #(
		.INIT('h8)
	) name1220 (
		\j4_pad ,
		\r0_pad ,
		_w1393_
	);
	LUT2 #(
		.INIT('h8)
	) name1221 (
		\k0_pad ,
		\r3_pad ,
		_w1394_
	);
	LUT2 #(
		.INIT('h8)
	) name1222 (
		\l0_pad ,
		\n3_pad ,
		_w1395_
	);
	LUT2 #(
		.INIT('h8)
	) name1223 (
		\p0_pad ,
		\u3_pad ,
		_w1396_
	);
	LUT2 #(
		.INIT('h8)
	) name1224 (
		\g3_pad ,
		\m0_pad ,
		_w1397_
	);
	LUT2 #(
		.INIT('h8)
	) name1225 (
		\n4_pad ,
		\q0_pad ,
		_w1398_
	);
	LUT2 #(
		.INIT('h1)
	) name1226 (
		_w1388_,
		_w1389_,
		_w1399_
	);
	LUT2 #(
		.INIT('h1)
	) name1227 (
		_w1390_,
		_w1391_,
		_w1400_
	);
	LUT2 #(
		.INIT('h1)
	) name1228 (
		_w1392_,
		_w1393_,
		_w1401_
	);
	LUT2 #(
		.INIT('h1)
	) name1229 (
		_w1394_,
		_w1395_,
		_w1402_
	);
	LUT2 #(
		.INIT('h1)
	) name1230 (
		_w1396_,
		_w1397_,
		_w1403_
	);
	LUT2 #(
		.INIT('h4)
	) name1231 (
		_w1398_,
		_w1403_,
		_w1404_
	);
	LUT2 #(
		.INIT('h8)
	) name1232 (
		_w1401_,
		_w1402_,
		_w1405_
	);
	LUT2 #(
		.INIT('h8)
	) name1233 (
		_w1399_,
		_w1400_,
		_w1406_
	);
	LUT2 #(
		.INIT('h8)
	) name1234 (
		_w1405_,
		_w1406_,
		_w1407_
	);
	LUT2 #(
		.INIT('h8)
	) name1235 (
		_w1404_,
		_w1407_,
		_w1408_
	);
	LUT2 #(
		.INIT('h1)
	) name1236 (
		\w2_pad ,
		_w242_,
		_w1409_
	);
	LUT2 #(
		.INIT('h2)
	) name1237 (
		\s1_pad ,
		_w263_,
		_w1410_
	);
	LUT2 #(
		.INIT('h4)
	) name1238 (
		\s1_pad ,
		_w263_,
		_w1411_
	);
	LUT2 #(
		.INIT('h1)
	) name1239 (
		_w1410_,
		_w1411_,
		_w1412_
	);
	LUT2 #(
		.INIT('h2)
	) name1240 (
		_w242_,
		_w1412_,
		_w1413_
	);
	LUT2 #(
		.INIT('h1)
	) name1241 (
		b_pad,
		_w1409_,
		_w1414_
	);
	LUT2 #(
		.INIT('h4)
	) name1242 (
		_w1413_,
		_w1414_,
		_w1415_
	);
	LUT2 #(
		.INIT('h8)
	) name1243 (
		_w273_,
		_w290_,
		_w1416_
	);
	LUT2 #(
		.INIT('h4)
	) name1244 (
		_w273_,
		_w283_,
		_w1417_
	);
	LUT2 #(
		.INIT('h1)
	) name1245 (
		_w303_,
		_w1416_,
		_w1418_
	);
	LUT2 #(
		.INIT('h4)
	) name1246 (
		_w1417_,
		_w1418_,
		_w1419_
	);
	LUT2 #(
		.INIT('h8)
	) name1247 (
		\s2_pad ,
		_w1419_,
		_w1420_
	);
	LUT2 #(
		.INIT('h1)
	) name1248 (
		\s2_pad ,
		_w1419_,
		_w1421_
	);
	LUT2 #(
		.INIT('h2)
	) name1249 (
		_w277_,
		_w1420_,
		_w1422_
	);
	LUT2 #(
		.INIT('h4)
	) name1250 (
		_w1421_,
		_w1422_,
		_w1423_
	);
	LUT2 #(
		.INIT('h8)
	) name1251 (
		\s3_pad ,
		_w363_,
		_w1424_
	);
	LUT2 #(
		.INIT('h1)
	) name1252 (
		\s3_pad ,
		_w363_,
		_w1425_
	);
	LUT2 #(
		.INIT('h2)
	) name1253 (
		_w316_,
		_w1424_,
		_w1426_
	);
	LUT2 #(
		.INIT('h4)
	) name1254 (
		_w1425_,
		_w1426_,
		_w1427_
	);
	LUT2 #(
		.INIT('h1)
	) name1255 (
		_w317_,
		_w1427_,
		_w1428_
	);
	LUT2 #(
		.INIT('h1)
	) name1256 (
		\s4_pad ,
		_w200_,
		_w1429_
	);
	LUT2 #(
		.INIT('h2)
	) name1257 (
		_w198_,
		_w201_,
		_w1430_
	);
	LUT2 #(
		.INIT('h4)
	) name1258 (
		_w1429_,
		_w1430_,
		_w1431_
	);
	assign \a10_pad  = _w205_ ;
	assign \a6_pad  = _w226_ ;
	assign \a7_pad  = _w271_ ;
	assign \a8_pad  = _w310_ ;
	assign \a9_pad  = _w372_ ;
	assign \b10_pad  = _w376_ ;
	assign \b6_pad  = _w415_ ;
	assign \b7_pad  = _w426_ ;
	assign \b8_pad  = _w431_ ;
	assign \b9_pad  = _w450_ ;
	assign \c10_pad  = _w454_ ;
	assign \c53  = _w463_ ;
	assign \c6_pad  = _w473_ ;
	assign \c7_pad  = _w489_ ;
	assign \c8_pad  = _w493_ ;
	assign \c9_pad  = _w505_ ;
	assign \d10_pad  = _w509_ ;
	assign \d6_pad  = _w515_ ;
	assign \d7_pad  = _w528_ ;
	assign \d8_pad  = _w540_ ;
	assign \d9_pad  = _w551_ ;
	assign \e10_pad  = _w556_ ;
	assign \e6_pad  = _w560_ ;
	assign \e7_pad  = _w573_ ;
	assign \e8_pad  = _w581_ ;
	assign \e9_pad  = _w597_ ;
	assign \f10_pad  = _w601_ ;
	assign \f22  = _w608_ ;
	assign \f6_pad  = _w612_ ;
	assign \f7_pad  = _w627_ ;
	assign \f8_pad  = _w635_ ;
	assign \f9_pad  = _w649_ ;
	assign \g10_pad  = _w653_ ;
	assign \g6_pad  = _w658_ ;
	assign \g7_pad  = _w671_ ;
	assign \g8_pad  = _w680_ ;
	assign \g9_pad  = _w693_ ;
	assign \h6_pad  = _w697_ ;
	assign \h7_pad  = _w708_ ;
	assign \h8_pad  = _w719_ ;
	assign \h9_pad  = _w733_ ;
	assign \i6_pad  = _w737_ ;
	assign \i7_pad  = _w738_ ;
	assign \i8_pad  = _w751_ ;
	assign \i9_pad  = _w762_ ;
	assign \j10_pad  = _w188_ ;
	assign \j6_pad  = _w766_ ;
	assign \j7_pad  = _w770_ ;
	assign \j8_pad  = _w779_ ;
	assign \j9_pad  = _w790_ ;
	assign \k10_pad  = _w793_ ;
	assign \k53  = _w797_ ;
	assign \k6_pad  = _w801_ ;
	assign \k7_pad  = _w805_ ;
	assign \k8_pad  = _w814_ ;
	assign \k9_pad  = _w815_ ;
	assign \l10_pad  = _w818_ ;
	assign \l7_pad  = _w832_ ;
	assign \l8_pad  = _w843_ ;
	assign \l9_pad  = _w846_ ;
	assign \m10_pad  = _w858_ ;
	assign \m7_pad  = _w865_ ;
	assign \m8_pad  = _w869_ ;
	assign \m9_pad  = _w872_ ;
	assign \n10_pad  = _w875_ ;
	assign \n6_pad  = _w250_ ;
	assign \n7_pad  = _w878_ ;
	assign \n8_pad  = _w886_ ;
	assign \n9_pad  = _w893_ ;
	assign \o10_pad  = _w851_ ;
	assign \o6_pad  = _w896_ ;
	assign \o7_pad  = _w904_ ;
	assign \o8_pad  = _w912_ ;
	assign \o9_pad  = _w919_ ;
	assign \p6_pad  = _w922_ ;
	assign \p7_pad  = _w929_ ;
	assign \p8_pad  = _w938_ ;
	assign \p9_pad  = _w941_ ;
	assign \q10_pad  = _w946_ ;
	assign \q6_pad  = _w951_ ;
	assign \q7_pad  = _w960_ ;
	assign \q8_pad  = _w965_ ;
	assign \q9_pad  = _w973_ ;
	assign \r10_pad  = _w977_ ;
	assign \r7_pad  = _w985_ ;
	assign \r8_pad  = _w989_ ;
	assign \r9_pad  = _w996_ ;
	assign \s5_pad  = _w1017_ ;
	assign \s7_pad  = _w1024_ ;
	assign \s8_pad  = _w1032_ ;
	assign \s9_pad  = _w1041_ ;
	assign \t10_pad  = _w1053_ ;
	assign \t5_pad  = _w1074_ ;
	assign \t6_pad  = _w1095_ ;
	assign \t7_pad  = _w1102_ ;
	assign \t8_pad  = _w1110_ ;
	assign \t9_pad  = _w1118_ ;
	assign \u5_pad  = _w1139_ ;
	assign \u7_pad  = _w1145_ ;
	assign \u8_pad  = _w1153_ ;
	assign \u9_pad  = _w1160_ ;
	assign \v10_pad  = _w311_ ;
	assign \v5_pad  = _w1181_ ;
	assign \v6_pad  = _w239_ ;
	assign \v7_pad  = _w1188_ ;
	assign \v8_pad  = _w1197_ ;
	assign \v9_pad  = _w1204_ ;
	assign \w10_pad  = _w1220_ ;
	assign \w5_pad  = _w1241_ ;
	assign \w6_pad  = _w1258_ ;
	assign \w7_pad  = _w1261_ ;
	assign \w8_pad  = _w1270_ ;
	assign \w9_pad  = _w1276_ ;
	assign \x10_pad  = _w1283_ ;
	assign \x21  = _w1287_ ;
	assign \x5_pad  = _w1308_ ;
	assign \x6_pad  = _w1315_ ;
	assign \x7_pad  = _w1319_ ;
	assign \x8_pad  = _w1326_ ;
	assign \x9_pad  = _w1333_ ;
	assign \y10_pad  = _w1340_ ;
	assign \y5_pad  = _w1361_ ;
	assign \y6_pad  = _w1368_ ;
	assign \y7_pad  = _w1376_ ;
	assign \y8_pad  = _w1384_ ;
	assign \y9_pad  = _w1387_ ;
	assign \z5_pad  = _w1408_ ;
	assign \z6_pad  = _w1415_ ;
	assign \z7_pad  = _w1423_ ;
	assign \z8_pad  = _w1428_ ;
	assign \z9_pad  = _w1431_ ;
endmodule;