module top( \IC0(32)_pad  , \IC1(33)_pad  , \IC2(34)_pad  , \IC3(35)_pad  , \IC4(36)_pad  , \IC5(37)_pad  , \IC6(38)_pad  , \IC7(39)_pad  , \ID0(0)_pad  , \ID1(1)_pad  , \ID10(10)_pad  , \ID11(11)_pad  , \ID12(12)_pad  , \ID13(13)_pad  , \ID14(14)_pad  , \ID15(15)_pad  , \ID16(16)_pad  , \ID17(17)_pad  , \ID18(18)_pad  , \ID19(19)_pad  , \ID2(2)_pad  , \ID20(20)_pad  , \ID21(21)_pad  , \ID22(22)_pad  , \ID23(23)_pad  , \ID24(24)_pad  , \ID25(25)_pad  , \ID26(26)_pad  , \ID27(27)_pad  , \ID28(28)_pad  , \ID29(29)_pad  , \ID3(3)_pad  , \ID30(30)_pad  , \ID31(31)_pad  , \ID4(4)_pad  , \ID5(5)_pad  , \ID6(6)_pad  , \ID7(7)_pad  , \ID8(8)_pad  , \ID9(9)_pad  , \R(40)_pad  , \OD0(242)_pad  , \OD1(241)_pad  , \OD10(232)_pad  , \OD11(231)_pad  , \OD12(230)_pad  , \OD13(229)_pad  , \OD14(228)_pad  , \OD15(227)_pad  , \OD16(226)_pad  , \OD17(225)_pad  , \OD18(224)_pad  , \OD19(223)_pad  , \OD2(240)_pad  , \OD20(222)_pad  , \OD21(221)_pad  , \OD22(220)_pad  , \OD23(219)_pad  , \OD24(218)_pad  , \OD25(217)_pad  , \OD26(216)_pad  , \OD27(215)_pad  , \OD28(214)_pad  , \OD29(213)_pad  , \OD3(239)_pad  , \OD30(212)_pad  , \OD31(211)_pad  , \OD4(238)_pad  , \OD5(237)_pad  , \OD6(236)_pad  , \OD7(235)_pad  , \OD8(234)_pad  , \OD9(233)_pad  );
  input \IC0(32)_pad  ;
  input \IC1(33)_pad  ;
  input \IC2(34)_pad  ;
  input \IC3(35)_pad  ;
  input \IC4(36)_pad  ;
  input \IC5(37)_pad  ;
  input \IC6(38)_pad  ;
  input \IC7(39)_pad  ;
  input \ID0(0)_pad  ;
  input \ID1(1)_pad  ;
  input \ID10(10)_pad  ;
  input \ID11(11)_pad  ;
  input \ID12(12)_pad  ;
  input \ID13(13)_pad  ;
  input \ID14(14)_pad  ;
  input \ID15(15)_pad  ;
  input \ID16(16)_pad  ;
  input \ID17(17)_pad  ;
  input \ID18(18)_pad  ;
  input \ID19(19)_pad  ;
  input \ID2(2)_pad  ;
  input \ID20(20)_pad  ;
  input \ID21(21)_pad  ;
  input \ID22(22)_pad  ;
  input \ID23(23)_pad  ;
  input \ID24(24)_pad  ;
  input \ID25(25)_pad  ;
  input \ID26(26)_pad  ;
  input \ID27(27)_pad  ;
  input \ID28(28)_pad  ;
  input \ID29(29)_pad  ;
  input \ID3(3)_pad  ;
  input \ID30(30)_pad  ;
  input \ID31(31)_pad  ;
  input \ID4(4)_pad  ;
  input \ID5(5)_pad  ;
  input \ID6(6)_pad  ;
  input \ID7(7)_pad  ;
  input \ID8(8)_pad  ;
  input \ID9(9)_pad  ;
  input \R(40)_pad  ;
  output \OD0(242)_pad  ;
  output \OD1(241)_pad  ;
  output \OD10(232)_pad  ;
  output \OD11(231)_pad  ;
  output \OD12(230)_pad  ;
  output \OD13(229)_pad  ;
  output \OD14(228)_pad  ;
  output \OD15(227)_pad  ;
  output \OD16(226)_pad  ;
  output \OD17(225)_pad  ;
  output \OD18(224)_pad  ;
  output \OD19(223)_pad  ;
  output \OD2(240)_pad  ;
  output \OD20(222)_pad  ;
  output \OD21(221)_pad  ;
  output \OD22(220)_pad  ;
  output \OD23(219)_pad  ;
  output \OD24(218)_pad  ;
  output \OD25(217)_pad  ;
  output \OD26(216)_pad  ;
  output \OD27(215)_pad  ;
  output \OD28(214)_pad  ;
  output \OD29(213)_pad  ;
  output \OD3(239)_pad  ;
  output \OD30(212)_pad  ;
  output \OD31(211)_pad  ;
  output \OD4(238)_pad  ;
  output \OD5(237)_pad  ;
  output \OD6(236)_pad  ;
  output \OD7(235)_pad  ;
  output \OD8(234)_pad  ;
  output \OD9(233)_pad  ;
  wire n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 ;
  assign n42 = ~\ID21(21)_pad  & ~\ID22(22)_pad  ;
  assign n43 = \ID21(21)_pad  & \ID22(22)_pad  ;
  assign n44 = ~n42 & ~n43 ;
  assign n45 = \ID20(20)_pad  & ~\ID23(23)_pad  ;
  assign n46 = ~\ID20(20)_pad  & \ID23(23)_pad  ;
  assign n47 = ~n45 & ~n46 ;
  assign n48 = n44 & n47 ;
  assign n49 = ~n44 & ~n47 ;
  assign n50 = ~n48 & ~n49 ;
  assign n51 = \IC0(32)_pad  & \R(40)_pad  ;
  assign n52 = n50 & n51 ;
  assign n53 = ~n50 & ~n51 ;
  assign n54 = ~n52 & ~n53 ;
  assign n55 = ~\ID17(17)_pad  & ~\ID18(18)_pad  ;
  assign n56 = \ID17(17)_pad  & \ID18(18)_pad  ;
  assign n57 = ~n55 & ~n56 ;
  assign n58 = \ID16(16)_pad  & ~\ID19(19)_pad  ;
  assign n59 = ~\ID16(16)_pad  & \ID19(19)_pad  ;
  assign n60 = ~n58 & ~n59 ;
  assign n61 = n57 & n60 ;
  assign n62 = ~n57 & ~n60 ;
  assign n63 = ~n61 & ~n62 ;
  assign n64 = n54 & n63 ;
  assign n65 = ~n54 & ~n63 ;
  assign n66 = ~n64 & ~n65 ;
  assign n67 = \ID12(12)_pad  & ~\ID8(8)_pad  ;
  assign n68 = ~\ID12(12)_pad  & \ID8(8)_pad  ;
  assign n69 = ~n67 & ~n68 ;
  assign n70 = \ID0(0)_pad  & ~\ID4(4)_pad  ;
  assign n71 = ~\ID0(0)_pad  & \ID4(4)_pad  ;
  assign n72 = ~n70 & ~n71 ;
  assign n73 = n69 & ~n72 ;
  assign n74 = ~n69 & n72 ;
  assign n75 = ~n73 & ~n74 ;
  assign n76 = n66 & n75 ;
  assign n77 = ~n66 & ~n75 ;
  assign n78 = ~n76 & ~n77 ;
  assign n153 = \IC3(35)_pad  & \R(40)_pad  ;
  assign n154 = ~n50 & n153 ;
  assign n155 = n50 & ~n153 ;
  assign n156 = ~n154 & ~n155 ;
  assign n157 = ~\ID11(11)_pad  & ~\ID15(15)_pad  ;
  assign n158 = \ID11(11)_pad  & \ID15(15)_pad  ;
  assign n159 = ~n157 & ~n158 ;
  assign n160 = \ID3(3)_pad  & n159 ;
  assign n161 = ~\ID3(3)_pad  & ~n159 ;
  assign n162 = ~n160 & ~n161 ;
  assign n163 = ~\ID29(29)_pad  & ~\ID30(30)_pad  ;
  assign n164 = \ID29(29)_pad  & \ID30(30)_pad  ;
  assign n165 = ~n163 & ~n164 ;
  assign n166 = \ID28(28)_pad  & ~\ID31(31)_pad  ;
  assign n167 = ~\ID28(28)_pad  & \ID31(31)_pad  ;
  assign n168 = ~n166 & ~n167 ;
  assign n169 = n165 & n168 ;
  assign n170 = ~n165 & ~n168 ;
  assign n171 = ~n169 & ~n170 ;
  assign n172 = \ID7(7)_pad  & ~n171 ;
  assign n173 = ~\ID7(7)_pad  & n171 ;
  assign n174 = ~n172 & ~n173 ;
  assign n175 = n162 & ~n174 ;
  assign n176 = ~n162 & n174 ;
  assign n177 = ~n175 & ~n176 ;
  assign n178 = n156 & n177 ;
  assign n179 = ~n156 & ~n177 ;
  assign n180 = ~n178 & ~n179 ;
  assign n185 = \ID26(26)_pad  & ~\ID27(27)_pad  ;
  assign n186 = ~\ID26(26)_pad  & \ID27(27)_pad  ;
  assign n187 = ~n185 & ~n186 ;
  assign n188 = \ID24(24)_pad  & ~\ID25(25)_pad  ;
  assign n189 = ~\ID24(24)_pad  & \ID25(25)_pad  ;
  assign n190 = ~n188 & ~n189 ;
  assign n191 = n187 & n190 ;
  assign n192 = ~n187 & ~n190 ;
  assign n193 = ~n191 & ~n192 ;
  assign n210 = \IC2(34)_pad  & \R(40)_pad  ;
  assign n211 = n63 & n210 ;
  assign n212 = ~n63 & ~n210 ;
  assign n213 = ~n211 & ~n212 ;
  assign n214 = n193 & n213 ;
  assign n215 = ~n193 & ~n213 ;
  assign n216 = ~n214 & ~n215 ;
  assign n217 = \ID10(10)_pad  & ~\ID14(14)_pad  ;
  assign n218 = ~\ID10(10)_pad  & \ID14(14)_pad  ;
  assign n219 = ~n217 & ~n218 ;
  assign n220 = \ID2(2)_pad  & ~\ID6(6)_pad  ;
  assign n221 = ~\ID2(2)_pad  & \ID6(6)_pad  ;
  assign n222 = ~n220 & ~n221 ;
  assign n223 = n219 & ~n222 ;
  assign n224 = ~n219 & n222 ;
  assign n225 = ~n223 & ~n224 ;
  assign n226 = n216 & n225 ;
  assign n227 = ~n216 & ~n225 ;
  assign n228 = ~n226 & ~n227 ;
  assign n181 = \IC1(33)_pad  & \R(40)_pad  ;
  assign n182 = n171 & n181 ;
  assign n183 = ~n171 & ~n181 ;
  assign n184 = ~n182 & ~n183 ;
  assign n194 = n184 & n193 ;
  assign n195 = ~n184 & ~n193 ;
  assign n196 = ~n194 & ~n195 ;
  assign n197 = \ID13(13)_pad  & ~\ID9(9)_pad  ;
  assign n198 = ~\ID13(13)_pad  & \ID9(9)_pad  ;
  assign n199 = ~n197 & ~n198 ;
  assign n200 = \ID1(1)_pad  & ~\ID5(5)_pad  ;
  assign n201 = ~\ID1(1)_pad  & \ID5(5)_pad  ;
  assign n202 = ~n200 & ~n201 ;
  assign n203 = n199 & ~n202 ;
  assign n204 = ~n199 & n202 ;
  assign n205 = ~n203 & ~n204 ;
  assign n206 = n196 & n205 ;
  assign n207 = ~n196 & ~n205 ;
  assign n208 = ~n206 & ~n207 ;
  assign n232 = ~n78 & ~n208 ;
  assign n233 = ~n228 & n232 ;
  assign n209 = n78 & ~n208 ;
  assign n229 = n209 & n228 ;
  assign n230 = n78 & n208 ;
  assign n231 = ~n228 & n230 ;
  assign n234 = ~n229 & ~n231 ;
  assign n235 = ~n233 & n234 ;
  assign n236 = n180 & ~n235 ;
  assign n237 = ~n180 & ~n228 ;
  assign n238 = n209 & n237 ;
  assign n239 = ~n236 & ~n238 ;
  assign n79 = ~\ID5(5)_pad  & ~\ID6(6)_pad  ;
  assign n80 = \ID5(5)_pad  & \ID6(6)_pad  ;
  assign n81 = ~n79 & ~n80 ;
  assign n82 = \ID4(4)_pad  & ~\ID7(7)_pad  ;
  assign n83 = ~\ID4(4)_pad  & \ID7(7)_pad  ;
  assign n84 = ~n82 & ~n83 ;
  assign n85 = n81 & n84 ;
  assign n86 = ~n81 & ~n84 ;
  assign n87 = ~n85 & ~n86 ;
  assign n88 = \ID12(12)_pad  & ~\ID15(15)_pad  ;
  assign n89 = ~\ID12(12)_pad  & \ID15(15)_pad  ;
  assign n90 = ~n88 & ~n89 ;
  assign n91 = \ID13(13)_pad  & ~\ID14(14)_pad  ;
  assign n92 = ~\ID13(13)_pad  & \ID14(14)_pad  ;
  assign n93 = ~n91 & ~n92 ;
  assign n94 = n90 & n93 ;
  assign n95 = ~n90 & ~n93 ;
  assign n96 = ~n94 & ~n95 ;
  assign n97 = \ID23(23)_pad  & n96 ;
  assign n98 = ~\ID23(23)_pad  & ~n96 ;
  assign n99 = ~n97 & ~n98 ;
  assign n100 = \ID19(19)_pad  & ~\ID31(31)_pad  ;
  assign n101 = ~\ID19(19)_pad  & \ID31(31)_pad  ;
  assign n102 = ~n100 & ~n101 ;
  assign n103 = \IC7(39)_pad  & \R(40)_pad  ;
  assign n104 = \ID27(27)_pad  & ~n103 ;
  assign n105 = ~\ID27(27)_pad  & n103 ;
  assign n106 = ~n104 & ~n105 ;
  assign n107 = n102 & n106 ;
  assign n108 = ~n102 & ~n106 ;
  assign n109 = ~n107 & ~n108 ;
  assign n110 = n99 & ~n109 ;
  assign n111 = ~n99 & n109 ;
  assign n112 = ~n110 & ~n111 ;
  assign n113 = n87 & n112 ;
  assign n114 = ~n87 & ~n112 ;
  assign n115 = ~n113 & ~n114 ;
  assign n116 = \ID2(2)_pad  & ~\ID3(3)_pad  ;
  assign n117 = ~\ID2(2)_pad  & \ID3(3)_pad  ;
  assign n118 = ~n116 & ~n117 ;
  assign n119 = \ID0(0)_pad  & ~\ID1(1)_pad  ;
  assign n120 = ~\ID0(0)_pad  & \ID1(1)_pad  ;
  assign n121 = ~n119 & ~n120 ;
  assign n122 = n118 & n121 ;
  assign n123 = ~n118 & ~n121 ;
  assign n124 = ~n122 & ~n123 ;
  assign n125 = \IC6(38)_pad  & \R(40)_pad  ;
  assign n126 = ~\ID11(11)_pad  & ~\ID8(8)_pad  ;
  assign n127 = \ID11(11)_pad  & \ID8(8)_pad  ;
  assign n128 = ~n126 & ~n127 ;
  assign n129 = \ID10(10)_pad  & ~\ID9(9)_pad  ;
  assign n130 = ~\ID10(10)_pad  & \ID9(9)_pad  ;
  assign n131 = ~n129 & ~n130 ;
  assign n132 = n128 & n131 ;
  assign n133 = ~n128 & ~n131 ;
  assign n134 = ~n132 & ~n133 ;
  assign n135 = n125 & ~n134 ;
  assign n136 = ~n125 & n134 ;
  assign n137 = ~n135 & ~n136 ;
  assign n138 = n124 & n137 ;
  assign n139 = ~n124 & ~n137 ;
  assign n140 = ~n138 & ~n139 ;
  assign n141 = \ID26(26)_pad  & ~\ID30(30)_pad  ;
  assign n142 = ~\ID26(26)_pad  & \ID30(30)_pad  ;
  assign n143 = ~n141 & ~n142 ;
  assign n144 = \ID18(18)_pad  & ~\ID22(22)_pad  ;
  assign n145 = ~\ID18(18)_pad  & \ID22(22)_pad  ;
  assign n146 = ~n144 & ~n145 ;
  assign n147 = n143 & ~n146 ;
  assign n148 = ~n143 & n146 ;
  assign n149 = ~n147 & ~n148 ;
  assign n150 = n140 & n149 ;
  assign n151 = ~n140 & ~n149 ;
  assign n152 = ~n150 & ~n151 ;
  assign n240 = ~n115 & ~n152 ;
  assign n241 = ~n239 & n240 ;
  assign n242 = \IC5(37)_pad  & \R(40)_pad  ;
  assign n243 = n134 & n242 ;
  assign n244 = ~n134 & ~n242 ;
  assign n245 = ~n243 & ~n244 ;
  assign n246 = n96 & n245 ;
  assign n247 = ~n96 & ~n245 ;
  assign n248 = ~n246 & ~n247 ;
  assign n249 = \ID25(25)_pad  & ~\ID29(29)_pad  ;
  assign n250 = ~\ID25(25)_pad  & \ID29(29)_pad  ;
  assign n251 = ~n249 & ~n250 ;
  assign n252 = \ID17(17)_pad  & ~\ID21(21)_pad  ;
  assign n253 = ~\ID17(17)_pad  & \ID21(21)_pad  ;
  assign n254 = ~n252 & ~n253 ;
  assign n255 = n251 & ~n254 ;
  assign n256 = ~n251 & n254 ;
  assign n257 = ~n255 & ~n256 ;
  assign n258 = n248 & n257 ;
  assign n259 = ~n248 & ~n257 ;
  assign n260 = ~n258 & ~n259 ;
  assign n261 = \IC4(36)_pad  & \R(40)_pad  ;
  assign n262 = n87 & n261 ;
  assign n263 = ~n87 & ~n261 ;
  assign n264 = ~n262 & ~n263 ;
  assign n265 = n124 & n264 ;
  assign n266 = ~n124 & ~n264 ;
  assign n267 = ~n265 & ~n266 ;
  assign n268 = \ID24(24)_pad  & ~\ID28(28)_pad  ;
  assign n269 = ~\ID24(24)_pad  & \ID28(28)_pad  ;
  assign n270 = ~n268 & ~n269 ;
  assign n271 = \ID16(16)_pad  & ~\ID20(20)_pad  ;
  assign n272 = ~\ID16(16)_pad  & \ID20(20)_pad  ;
  assign n273 = ~n271 & ~n272 ;
  assign n274 = n270 & ~n273 ;
  assign n275 = ~n270 & n273 ;
  assign n276 = ~n274 & ~n275 ;
  assign n277 = n267 & n276 ;
  assign n278 = ~n267 & ~n276 ;
  assign n279 = ~n277 & ~n278 ;
  assign n280 = ~n260 & n279 ;
  assign n281 = n241 & n280 ;
  assign n282 = ~n78 & n281 ;
  assign n283 = \ID0(0)_pad  & ~n282 ;
  assign n284 = ~\ID0(0)_pad  & n282 ;
  assign n285 = ~n283 & ~n284 ;
  assign n286 = n208 & n281 ;
  assign n287 = \ID1(1)_pad  & ~n286 ;
  assign n288 = ~\ID1(1)_pad  & n286 ;
  assign n289 = ~n287 & ~n288 ;
  assign n290 = n260 & ~n279 ;
  assign n291 = n241 & n290 ;
  assign n292 = n228 & n291 ;
  assign n293 = \ID10(10)_pad  & ~n292 ;
  assign n294 = ~\ID10(10)_pad  & n292 ;
  assign n295 = ~n293 & ~n294 ;
  assign n296 = ~n180 & n291 ;
  assign n297 = \ID11(11)_pad  & ~n296 ;
  assign n298 = ~\ID11(11)_pad  & n296 ;
  assign n299 = ~n297 & ~n298 ;
  assign n300 = n115 & ~n239 ;
  assign n301 = n152 & n290 ;
  assign n302 = n300 & n301 ;
  assign n303 = ~n78 & n302 ;
  assign n304 = \ID12(12)_pad  & ~n303 ;
  assign n305 = ~\ID12(12)_pad  & n303 ;
  assign n306 = ~n304 & ~n305 ;
  assign n307 = n208 & n302 ;
  assign n308 = \ID13(13)_pad  & ~n307 ;
  assign n309 = ~\ID13(13)_pad  & n307 ;
  assign n310 = ~n308 & ~n309 ;
  assign n311 = n228 & n302 ;
  assign n312 = \ID14(14)_pad  & ~n311 ;
  assign n313 = ~\ID14(14)_pad  & n311 ;
  assign n314 = ~n312 & ~n313 ;
  assign n315 = ~n180 & n302 ;
  assign n316 = \ID15(15)_pad  & ~n315 ;
  assign n317 = ~\ID15(15)_pad  & n315 ;
  assign n318 = ~n316 & ~n317 ;
  assign n320 = ~n260 & ~n279 ;
  assign n321 = ~n152 & n320 ;
  assign n319 = n152 & n280 ;
  assign n322 = ~n301 & ~n319 ;
  assign n323 = ~n321 & n322 ;
  assign n324 = ~n115 & ~n323 ;
  assign n325 = n115 & n152 ;
  assign n326 = n320 & n325 ;
  assign n327 = ~n324 & ~n326 ;
  assign n328 = n180 & n228 ;
  assign n329 = ~n327 & n328 ;
  assign n330 = n232 & n329 ;
  assign n331 = n279 & n330 ;
  assign n332 = \ID16(16)_pad  & ~n331 ;
  assign n333 = ~\ID16(16)_pad  & n331 ;
  assign n334 = ~n332 & ~n333 ;
  assign n335 = n260 & n330 ;
  assign n336 = \ID17(17)_pad  & ~n335 ;
  assign n337 = ~\ID17(17)_pad  & n335 ;
  assign n338 = ~n336 & ~n337 ;
  assign n339 = ~n152 & n330 ;
  assign n340 = \ID18(18)_pad  & ~n339 ;
  assign n341 = ~\ID18(18)_pad  & n339 ;
  assign n342 = ~n340 & ~n341 ;
  assign n343 = n115 & n330 ;
  assign n344 = \ID19(19)_pad  & ~n343 ;
  assign n345 = ~\ID19(19)_pad  & n343 ;
  assign n346 = ~n344 & ~n345 ;
  assign n347 = n228 & n281 ;
  assign n348 = \ID2(2)_pad  & ~n347 ;
  assign n349 = ~\ID2(2)_pad  & n347 ;
  assign n350 = ~n348 & ~n349 ;
  assign n351 = ~n180 & ~n327 ;
  assign n352 = n233 & n351 ;
  assign n353 = n279 & n352 ;
  assign n354 = \ID20(20)_pad  & ~n353 ;
  assign n355 = ~\ID20(20)_pad  & n353 ;
  assign n356 = ~n354 & ~n355 ;
  assign n357 = n260 & n352 ;
  assign n358 = \ID21(21)_pad  & ~n357 ;
  assign n359 = ~\ID21(21)_pad  & n357 ;
  assign n360 = ~n358 & ~n359 ;
  assign n361 = ~n152 & n352 ;
  assign n362 = \ID22(22)_pad  & ~n361 ;
  assign n363 = ~\ID22(22)_pad  & n361 ;
  assign n364 = ~n362 & ~n363 ;
  assign n365 = n115 & n352 ;
  assign n366 = \ID23(23)_pad  & ~n365 ;
  assign n367 = ~\ID23(23)_pad  & n365 ;
  assign n368 = ~n366 & ~n367 ;
  assign n369 = n230 & n329 ;
  assign n370 = n279 & n369 ;
  assign n371 = \ID24(24)_pad  & ~n370 ;
  assign n372 = ~\ID24(24)_pad  & n370 ;
  assign n373 = ~n371 & ~n372 ;
  assign n374 = n260 & n369 ;
  assign n375 = \ID25(25)_pad  & ~n374 ;
  assign n376 = ~\ID25(25)_pad  & n374 ;
  assign n377 = ~n375 & ~n376 ;
  assign n378 = ~n152 & n369 ;
  assign n379 = \ID26(26)_pad  & ~n378 ;
  assign n380 = ~\ID26(26)_pad  & n378 ;
  assign n381 = ~n379 & ~n380 ;
  assign n382 = n115 & n369 ;
  assign n383 = \ID27(27)_pad  & ~n382 ;
  assign n384 = ~\ID27(27)_pad  & n382 ;
  assign n385 = ~n383 & ~n384 ;
  assign n386 = n231 & n351 ;
  assign n387 = n279 & n386 ;
  assign n388 = \ID28(28)_pad  & ~n387 ;
  assign n389 = ~\ID28(28)_pad  & n387 ;
  assign n390 = ~n388 & ~n389 ;
  assign n391 = n260 & n386 ;
  assign n392 = \ID29(29)_pad  & ~n391 ;
  assign n393 = ~\ID29(29)_pad  & n391 ;
  assign n394 = ~n392 & ~n393 ;
  assign n395 = ~n180 & n281 ;
  assign n396 = \ID3(3)_pad  & ~n395 ;
  assign n397 = ~\ID3(3)_pad  & n395 ;
  assign n398 = ~n396 & ~n397 ;
  assign n399 = ~n152 & n386 ;
  assign n400 = \ID30(30)_pad  & ~n399 ;
  assign n401 = ~\ID30(30)_pad  & n399 ;
  assign n402 = ~n400 & ~n401 ;
  assign n403 = n115 & n386 ;
  assign n404 = \ID31(31)_pad  & ~n403 ;
  assign n405 = ~\ID31(31)_pad  & n403 ;
  assign n406 = ~n404 & ~n405 ;
  assign n407 = n300 & n319 ;
  assign n408 = ~n78 & n407 ;
  assign n409 = \ID4(4)_pad  & ~n408 ;
  assign n410 = ~\ID4(4)_pad  & n408 ;
  assign n411 = ~n409 & ~n410 ;
  assign n412 = n208 & n407 ;
  assign n413 = \ID5(5)_pad  & ~n412 ;
  assign n414 = ~\ID5(5)_pad  & n412 ;
  assign n415 = ~n413 & ~n414 ;
  assign n416 = n228 & n407 ;
  assign n417 = \ID6(6)_pad  & ~n416 ;
  assign n418 = ~\ID6(6)_pad  & n416 ;
  assign n419 = ~n417 & ~n418 ;
  assign n420 = ~n180 & n407 ;
  assign n421 = \ID7(7)_pad  & ~n420 ;
  assign n422 = ~\ID7(7)_pad  & n420 ;
  assign n423 = ~n421 & ~n422 ;
  assign n424 = ~n78 & n291 ;
  assign n425 = \ID8(8)_pad  & ~n424 ;
  assign n426 = ~\ID8(8)_pad  & n424 ;
  assign n427 = ~n425 & ~n426 ;
  assign n428 = n208 & n291 ;
  assign n429 = \ID9(9)_pad  & ~n428 ;
  assign n430 = ~\ID9(9)_pad  & n428 ;
  assign n431 = ~n429 & ~n430 ;
  assign \OD0(242)_pad  = ~n285 ;
  assign \OD1(241)_pad  = ~n289 ;
  assign \OD10(232)_pad  = ~n295 ;
  assign \OD11(231)_pad  = ~n299 ;
  assign \OD12(230)_pad  = ~n306 ;
  assign \OD13(229)_pad  = ~n310 ;
  assign \OD14(228)_pad  = ~n314 ;
  assign \OD15(227)_pad  = ~n318 ;
  assign \OD16(226)_pad  = ~n334 ;
  assign \OD17(225)_pad  = ~n338 ;
  assign \OD18(224)_pad  = ~n342 ;
  assign \OD19(223)_pad  = ~n346 ;
  assign \OD2(240)_pad  = ~n350 ;
  assign \OD20(222)_pad  = ~n356 ;
  assign \OD21(221)_pad  = ~n360 ;
  assign \OD22(220)_pad  = ~n364 ;
  assign \OD23(219)_pad  = ~n368 ;
  assign \OD24(218)_pad  = ~n373 ;
  assign \OD25(217)_pad  = ~n377 ;
  assign \OD26(216)_pad  = ~n381 ;
  assign \OD27(215)_pad  = ~n385 ;
  assign \OD28(214)_pad  = ~n390 ;
  assign \OD29(213)_pad  = ~n394 ;
  assign \OD3(239)_pad  = ~n398 ;
  assign \OD30(212)_pad  = ~n402 ;
  assign \OD31(211)_pad  = ~n406 ;
  assign \OD4(238)_pad  = ~n411 ;
  assign \OD5(237)_pad  = ~n415 ;
  assign \OD6(236)_pad  = ~n419 ;
  assign \OD7(235)_pad  = ~n423 ;
  assign \OD8(234)_pad  = ~n427 ;
  assign \OD9(233)_pad  = ~n431 ;
endmodule
