module top( a_pad , b_pad , c_pad , d_pad , e_pad , f_pad , g_pad , h_pad , i_pad , j_pad , k_pad , l_pad , m_pad , n_pad );
  input a_pad ;
  input b_pad ;
  input c_pad ;
  input d_pad ;
  input e_pad ;
  input f_pad ;
  input g_pad ;
  input h_pad ;
  input i_pad ;
  input j_pad ;
  input k_pad ;
  output l_pad ;
  output m_pad ;
  output n_pad ;
  wire n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 ;
  assign n12 = ~f_pad & g_pad ;
  assign n13 = ~h_pad & i_pad ;
  assign n14 = ~j_pad & k_pad ;
  assign n15 = ~n13 & ~n14 ;
  assign n16 = h_pad & ~i_pad ;
  assign n17 = f_pad & ~g_pad ;
  assign n18 = ~n16 & ~n17 ;
  assign n19 = ~n15 & n18 ;
  assign n20 = ~n12 & ~n19 ;
  assign n21 = ~d_pad & ~e_pad ;
  assign n22 = d_pad & e_pad ;
  assign n23 = ~n21 & ~n22 ;
  assign n24 = b_pad & ~n23 ;
  assign n25 = ~n20 & n24 ;
  assign n26 = b_pad & ~d_pad ;
  assign n27 = e_pad & n26 ;
  assign n28 = ~a_pad & ~n27 ;
  assign n29 = ~n25 & n28 ;
  assign n31 = j_pad & ~k_pad ;
  assign n32 = n18 & ~n31 ;
  assign n30 = ~n12 & ~n13 ;
  assign n33 = ~n14 & n30 ;
  assign n34 = n24 & n33 ;
  assign n35 = n32 & n34 ;
  assign n38 = ~n17 & ~n30 ;
  assign n39 = n24 & ~n32 ;
  assign n40 = ~n38 & n39 ;
  assign n36 = b_pad & d_pad ;
  assign n37 = ~e_pad & n36 ;
  assign n41 = ~c_pad & ~n37 ;
  assign n42 = ~n40 & n41 ;
  assign l_pad = ~n29 ;
  assign m_pad = n35 ;
  assign n_pad = ~n42 ;
endmodule
