module top (\a0_pad , \a1_pad , \a2_pad , \a3_pad , \a4_pad , \b0_pad , \b1_pad , \b2_pad , \b3_pad , \b4_pad , b_pad, \c0_pad , \c1_pad , \c2_pad , \c3_pad , \c4_pad , c_pad, \d0_pad , \d1_pad , \d2_pad , \d3_pad , \d4_pad , d_pad, \e0_pad , \e1_pad , \e2_pad , \e3_pad , \e4_pad , e_pad, \f0_pad , \f1_pad , \f2_pad , \f3_pad , \f4_pad , f_pad, \g0_pad , \g1_pad , \g2_pad , \g3_pad , \g4_pad , g_pad, \h0_pad , \h1_pad , \h2_pad , \h3_pad , \h4_pad , h_pad, \i0_pad , \i1_pad , \i2_pad , \i3_pad , i_pad, \j0_pad , \j1_pad , \j2_pad , \j3_pad , j_pad, \k0_pad , \k1_pad , \k2_pad , \k3_pad , k_pad, \l0_pad , \l1_pad , \l2_pad , \l3_pad , l_pad, \m0_pad , \m1_pad , \m2_pad , \m3_pad , m_pad, \n0_pad , \n1_pad , \n2_pad , \n3_pad , n_pad, \o0_pad , \o1_pad , \o2_pad , \o3_pad , o_pad, \p1_pad , \p2_pad , \p3_pad , p_pad, \q1_pad , \q2_pad , \q3_pad , q_pad, \r0_pad , \r1_pad , \r2_pad , \r3_pad , r_pad, \s0_pad , \s1_pad , \s2_pad , \s3_pad , s_pad, \t0_pad , \t1_pad , \t2_pad , \t3_pad , t_pad, \u0_pad , \u1_pad , \u2_pad , \u3_pad , u_pad, \v0_pad , \v1_pad , \v2_pad , \v3_pad , v_pad, \w0_pad , \w1_pad , \w2_pad , \w3_pad , w_pad, \x0_pad , \x1_pad , \x2_pad , \x3_pad , x_pad, \y0_pad , \y1_pad , \y2_pad , \y3_pad , y_pad, \z0_pad , \z1_pad , \z2_pad , \z3_pad , z_pad, \a5_pad , \a6_pad , \a7_pad , \a8_pad , \b5_pad , \b6_pad , \b7_pad , \b8_pad , \c5_pad , \c6_pad , \c7_pad , \c8_pad , \d5_pad , \d6_pad , \d7_pad , \e5_pad , \e6_pad , \e7_pad , \f5_pad , \f6_pad , \f7_pad , \g5_pad , \g6_pad , \g7_pad , \h5_pad , \h6_pad , \h7_pad , \i4_pad , \i5_pad , \i6_pad , \i7_pad , \j4_pad , \j5_pad , \j6_pad , \j7_pad , \k4_pad , \k5_pad , \k6_pad , \k7_pad , \l4_pad , \l5_pad , \l6_pad , \l7_pad , \m4_pad , \m5_pad , \m6_pad , \m7_pad , \n4_pad , \n5_pad , \n6_pad , \n7_pad , \o4_pad , \o5_pad , \o6_pad , \o7_pad , \p4_pad , \p5_pad , \p6_pad , \p7_pad , \q4_pad , \q5_pad , \q6_pad , \q7_pad , \r4_pad , \r5_pad , \r6_pad , \r7_pad , \s4_pad , \s5_pad , \s6_pad , \s7_pad , \t4_pad , \t5_pad , \t6_pad , \t7_pad , \u4_pad , \u5_pad , \u6_pad , \u7_pad , \v4_pad , \v5_pad , \v6_pad , \v7_pad , \w4_pad , \w5_pad , \w6_pad , \w7_pad , \x4_pad , \x5_pad , \x6_pad , \x7_pad , \y4_pad , \y5_pad , \y6_pad , \y7_pad , \z4_pad , \z5_pad , \z6_pad , \z7_pad );
	input \a0_pad  ;
	input \a1_pad  ;
	input \a2_pad  ;
	input \a3_pad  ;
	input \a4_pad  ;
	input \b0_pad  ;
	input \b1_pad  ;
	input \b2_pad  ;
	input \b3_pad  ;
	input \b4_pad  ;
	input b_pad ;
	input \c0_pad  ;
	input \c1_pad  ;
	input \c2_pad  ;
	input \c3_pad  ;
	input \c4_pad  ;
	input c_pad ;
	input \d0_pad  ;
	input \d1_pad  ;
	input \d2_pad  ;
	input \d3_pad  ;
	input \d4_pad  ;
	input d_pad ;
	input \e0_pad  ;
	input \e1_pad  ;
	input \e2_pad  ;
	input \e3_pad  ;
	input \e4_pad  ;
	input e_pad ;
	input \f0_pad  ;
	input \f1_pad  ;
	input \f2_pad  ;
	input \f3_pad  ;
	input \f4_pad  ;
	input f_pad ;
	input \g0_pad  ;
	input \g1_pad  ;
	input \g2_pad  ;
	input \g3_pad  ;
	input \g4_pad  ;
	input g_pad ;
	input \h0_pad  ;
	input \h1_pad  ;
	input \h2_pad  ;
	input \h3_pad  ;
	input \h4_pad  ;
	input h_pad ;
	input \i0_pad  ;
	input \i1_pad  ;
	input \i2_pad  ;
	input \i3_pad  ;
	input i_pad ;
	input \j0_pad  ;
	input \j1_pad  ;
	input \j2_pad  ;
	input \j3_pad  ;
	input j_pad ;
	input \k0_pad  ;
	input \k1_pad  ;
	input \k2_pad  ;
	input \k3_pad  ;
	input k_pad ;
	input \l0_pad  ;
	input \l1_pad  ;
	input \l2_pad  ;
	input \l3_pad  ;
	input l_pad ;
	input \m0_pad  ;
	input \m1_pad  ;
	input \m2_pad  ;
	input \m3_pad  ;
	input m_pad ;
	input \n0_pad  ;
	input \n1_pad  ;
	input \n2_pad  ;
	input \n3_pad  ;
	input n_pad ;
	input \o0_pad  ;
	input \o1_pad  ;
	input \o2_pad  ;
	input \o3_pad  ;
	input o_pad ;
	input \p1_pad  ;
	input \p2_pad  ;
	input \p3_pad  ;
	input p_pad ;
	input \q1_pad  ;
	input \q2_pad  ;
	input \q3_pad  ;
	input q_pad ;
	input \r0_pad  ;
	input \r1_pad  ;
	input \r2_pad  ;
	input \r3_pad  ;
	input r_pad ;
	input \s0_pad  ;
	input \s1_pad  ;
	input \s2_pad  ;
	input \s3_pad  ;
	input s_pad ;
	input \t0_pad  ;
	input \t1_pad  ;
	input \t2_pad  ;
	input \t3_pad  ;
	input t_pad ;
	input \u0_pad  ;
	input \u1_pad  ;
	input \u2_pad  ;
	input \u3_pad  ;
	input u_pad ;
	input \v0_pad  ;
	input \v1_pad  ;
	input \v2_pad  ;
	input \v3_pad  ;
	input v_pad ;
	input \w0_pad  ;
	input \w1_pad  ;
	input \w2_pad  ;
	input \w3_pad  ;
	input w_pad ;
	input \x0_pad  ;
	input \x1_pad  ;
	input \x2_pad  ;
	input \x3_pad  ;
	input x_pad ;
	input \y0_pad  ;
	input \y1_pad  ;
	input \y2_pad  ;
	input \y3_pad  ;
	input y_pad ;
	input \z0_pad  ;
	input \z1_pad  ;
	input \z2_pad  ;
	input \z3_pad  ;
	input z_pad ;
	output \a5_pad  ;
	output \a6_pad  ;
	output \a7_pad  ;
	output \a8_pad  ;
	output \b5_pad  ;
	output \b6_pad  ;
	output \b7_pad  ;
	output \b8_pad  ;
	output \c5_pad  ;
	output \c6_pad  ;
	output \c7_pad  ;
	output \c8_pad  ;
	output \d5_pad  ;
	output \d6_pad  ;
	output \d7_pad  ;
	output \e5_pad  ;
	output \e6_pad  ;
	output \e7_pad  ;
	output \f5_pad  ;
	output \f6_pad  ;
	output \f7_pad  ;
	output \g5_pad  ;
	output \g6_pad  ;
	output \g7_pad  ;
	output \h5_pad  ;
	output \h6_pad  ;
	output \h7_pad  ;
	output \i4_pad  ;
	output \i5_pad  ;
	output \i6_pad  ;
	output \i7_pad  ;
	output \j4_pad  ;
	output \j5_pad  ;
	output \j6_pad  ;
	output \j7_pad  ;
	output \k4_pad  ;
	output \k5_pad  ;
	output \k6_pad  ;
	output \k7_pad  ;
	output \l4_pad  ;
	output \l5_pad  ;
	output \l6_pad  ;
	output \l7_pad  ;
	output \m4_pad  ;
	output \m5_pad  ;
	output \m6_pad  ;
	output \m7_pad  ;
	output \n4_pad  ;
	output \n5_pad  ;
	output \n6_pad  ;
	output \n7_pad  ;
	output \o4_pad  ;
	output \o5_pad  ;
	output \o6_pad  ;
	output \o7_pad  ;
	output \p4_pad  ;
	output \p5_pad  ;
	output \p6_pad  ;
	output \p7_pad  ;
	output \q4_pad  ;
	output \q5_pad  ;
	output \q6_pad  ;
	output \q7_pad  ;
	output \r4_pad  ;
	output \r5_pad  ;
	output \r6_pad  ;
	output \r7_pad  ;
	output \s4_pad  ;
	output \s5_pad  ;
	output \s6_pad  ;
	output \s7_pad  ;
	output \t4_pad  ;
	output \t5_pad  ;
	output \t6_pad  ;
	output \t7_pad  ;
	output \u4_pad  ;
	output \u5_pad  ;
	output \u6_pad  ;
	output \u7_pad  ;
	output \v4_pad  ;
	output \v5_pad  ;
	output \v6_pad  ;
	output \v7_pad  ;
	output \w4_pad  ;
	output \w5_pad  ;
	output \w6_pad  ;
	output \w7_pad  ;
	output \x4_pad  ;
	output \x5_pad  ;
	output \x6_pad  ;
	output \x7_pad  ;
	output \y4_pad  ;
	output \y5_pad  ;
	output \y6_pad  ;
	output \y7_pad  ;
	output \z4_pad  ;
	output \z5_pad  ;
	output \z6_pad  ;
	output \z7_pad  ;
	wire _w741_ ;
	wire _w740_ ;
	wire _w739_ ;
	wire _w738_ ;
	wire _w737_ ;
	wire _w736_ ;
	wire _w735_ ;
	wire _w734_ ;
	wire _w733_ ;
	wire _w732_ ;
	wire _w731_ ;
	wire _w730_ ;
	wire _w729_ ;
	wire _w728_ ;
	wire _w727_ ;
	wire _w726_ ;
	wire _w725_ ;
	wire _w724_ ;
	wire _w723_ ;
	wire _w722_ ;
	wire _w721_ ;
	wire _w720_ ;
	wire _w719_ ;
	wire _w718_ ;
	wire _w717_ ;
	wire _w716_ ;
	wire _w715_ ;
	wire _w714_ ;
	wire _w713_ ;
	wire _w712_ ;
	wire _w711_ ;
	wire _w710_ ;
	wire _w709_ ;
	wire _w708_ ;
	wire _w707_ ;
	wire _w706_ ;
	wire _w705_ ;
	wire _w704_ ;
	wire _w703_ ;
	wire _w702_ ;
	wire _w701_ ;
	wire _w700_ ;
	wire _w699_ ;
	wire _w698_ ;
	wire _w697_ ;
	wire _w696_ ;
	wire _w695_ ;
	wire _w694_ ;
	wire _w693_ ;
	wire _w692_ ;
	wire _w691_ ;
	wire _w690_ ;
	wire _w689_ ;
	wire _w688_ ;
	wire _w687_ ;
	wire _w686_ ;
	wire _w685_ ;
	wire _w684_ ;
	wire _w683_ ;
	wire _w682_ ;
	wire _w681_ ;
	wire _w680_ ;
	wire _w679_ ;
	wire _w678_ ;
	wire _w677_ ;
	wire _w392_ ;
	wire _w391_ ;
	wire _w390_ ;
	wire _w389_ ;
	wire _w388_ ;
	wire _w387_ ;
	wire _w386_ ;
	wire _w385_ ;
	wire _w384_ ;
	wire _w383_ ;
	wire _w382_ ;
	wire _w381_ ;
	wire _w380_ ;
	wire _w379_ ;
	wire _w378_ ;
	wire _w377_ ;
	wire _w376_ ;
	wire _w375_ ;
	wire _w374_ ;
	wire _w373_ ;
	wire _w372_ ;
	wire _w371_ ;
	wire _w370_ ;
	wire _w369_ ;
	wire _w368_ ;
	wire _w367_ ;
	wire _w366_ ;
	wire _w365_ ;
	wire _w364_ ;
	wire _w363_ ;
	wire _w362_ ;
	wire _w361_ ;
	wire _w360_ ;
	wire _w359_ ;
	wire _w358_ ;
	wire _w357_ ;
	wire _w356_ ;
	wire _w355_ ;
	wire _w354_ ;
	wire _w353_ ;
	wire _w352_ ;
	wire _w351_ ;
	wire _w350_ ;
	wire _w349_ ;
	wire _w348_ ;
	wire _w347_ ;
	wire _w346_ ;
	wire _w345_ ;
	wire _w344_ ;
	wire _w343_ ;
	wire _w342_ ;
	wire _w341_ ;
	wire _w340_ ;
	wire _w339_ ;
	wire _w338_ ;
	wire _w337_ ;
	wire _w336_ ;
	wire _w335_ ;
	wire _w334_ ;
	wire _w333_ ;
	wire _w332_ ;
	wire _w331_ ;
	wire _w330_ ;
	wire _w329_ ;
	wire _w328_ ;
	wire _w327_ ;
	wire _w326_ ;
	wire _w325_ ;
	wire _w324_ ;
	wire _w323_ ;
	wire _w322_ ;
	wire _w321_ ;
	wire _w320_ ;
	wire _w319_ ;
	wire _w318_ ;
	wire _w317_ ;
	wire _w316_ ;
	wire _w315_ ;
	wire _w314_ ;
	wire _w313_ ;
	wire _w312_ ;
	wire _w311_ ;
	wire _w310_ ;
	wire _w309_ ;
	wire _w308_ ;
	wire _w307_ ;
	wire _w306_ ;
	wire _w305_ ;
	wire _w304_ ;
	wire _w303_ ;
	wire _w302_ ;
	wire _w301_ ;
	wire _w300_ ;
	wire _w299_ ;
	wire _w298_ ;
	wire _w297_ ;
	wire _w296_ ;
	wire _w295_ ;
	wire _w294_ ;
	wire _w293_ ;
	wire _w292_ ;
	wire _w291_ ;
	wire _w290_ ;
	wire _w289_ ;
	wire _w288_ ;
	wire _w287_ ;
	wire _w286_ ;
	wire _w285_ ;
	wire _w284_ ;
	wire _w283_ ;
	wire _w282_ ;
	wire _w281_ ;
	wire _w280_ ;
	wire _w279_ ;
	wire _w278_ ;
	wire _w277_ ;
	wire _w276_ ;
	wire _w275_ ;
	wire _w274_ ;
	wire _w273_ ;
	wire _w272_ ;
	wire _w271_ ;
	wire _w270_ ;
	wire _w269_ ;
	wire _w268_ ;
	wire _w267_ ;
	wire _w266_ ;
	wire _w265_ ;
	wire _w264_ ;
	wire _w263_ ;
	wire _w194_ ;
	wire _w193_ ;
	wire _w192_ ;
	wire _w191_ ;
	wire _w190_ ;
	wire _w189_ ;
	wire _w188_ ;
	wire _w187_ ;
	wire _w186_ ;
	wire _w185_ ;
	wire _w184_ ;
	wire _w183_ ;
	wire _w182_ ;
	wire _w181_ ;
	wire _w180_ ;
	wire _w179_ ;
	wire _w178_ ;
	wire _w177_ ;
	wire _w176_ ;
	wire _w175_ ;
	wire _w174_ ;
	wire _w173_ ;
	wire _w172_ ;
	wire _w171_ ;
	wire _w170_ ;
	wire _w169_ ;
	wire _w168_ ;
	wire _w167_ ;
	wire _w166_ ;
	wire _w165_ ;
	wire _w148_ ;
	wire _w147_ ;
	wire _w146_ ;
	wire _w145_ ;
	wire _w144_ ;
	wire _w143_ ;
	wire _w142_ ;
	wire _w141_ ;
	wire _w140_ ;
	wire _w139_ ;
	wire _w138_ ;
	wire _w137_ ;
	wire _w136_ ;
	wire _w149_ ;
	wire _w150_ ;
	wire _w151_ ;
	wire _w152_ ;
	wire _w153_ ;
	wire _w154_ ;
	wire _w155_ ;
	wire _w156_ ;
	wire _w157_ ;
	wire _w158_ ;
	wire _w159_ ;
	wire _w160_ ;
	wire _w161_ ;
	wire _w162_ ;
	wire _w163_ ;
	wire _w164_ ;
	wire _w195_ ;
	wire _w196_ ;
	wire _w197_ ;
	wire _w198_ ;
	wire _w199_ ;
	wire _w200_ ;
	wire _w201_ ;
	wire _w202_ ;
	wire _w203_ ;
	wire _w204_ ;
	wire _w205_ ;
	wire _w206_ ;
	wire _w207_ ;
	wire _w208_ ;
	wire _w209_ ;
	wire _w210_ ;
	wire _w211_ ;
	wire _w212_ ;
	wire _w213_ ;
	wire _w214_ ;
	wire _w215_ ;
	wire _w216_ ;
	wire _w217_ ;
	wire _w218_ ;
	wire _w219_ ;
	wire _w220_ ;
	wire _w221_ ;
	wire _w222_ ;
	wire _w223_ ;
	wire _w224_ ;
	wire _w225_ ;
	wire _w226_ ;
	wire _w227_ ;
	wire _w228_ ;
	wire _w229_ ;
	wire _w230_ ;
	wire _w231_ ;
	wire _w232_ ;
	wire _w233_ ;
	wire _w234_ ;
	wire _w235_ ;
	wire _w236_ ;
	wire _w237_ ;
	wire _w238_ ;
	wire _w239_ ;
	wire _w240_ ;
	wire _w241_ ;
	wire _w242_ ;
	wire _w243_ ;
	wire _w244_ ;
	wire _w245_ ;
	wire _w246_ ;
	wire _w247_ ;
	wire _w248_ ;
	wire _w249_ ;
	wire _w250_ ;
	wire _w251_ ;
	wire _w252_ ;
	wire _w253_ ;
	wire _w254_ ;
	wire _w255_ ;
	wire _w256_ ;
	wire _w257_ ;
	wire _w258_ ;
	wire _w259_ ;
	wire _w260_ ;
	wire _w261_ ;
	wire _w262_ ;
	wire _w393_ ;
	wire _w394_ ;
	wire _w395_ ;
	wire _w396_ ;
	wire _w397_ ;
	wire _w398_ ;
	wire _w399_ ;
	wire _w400_ ;
	wire _w401_ ;
	wire _w402_ ;
	wire _w403_ ;
	wire _w404_ ;
	wire _w405_ ;
	wire _w406_ ;
	wire _w407_ ;
	wire _w408_ ;
	wire _w409_ ;
	wire _w410_ ;
	wire _w411_ ;
	wire _w412_ ;
	wire _w413_ ;
	wire _w414_ ;
	wire _w415_ ;
	wire _w416_ ;
	wire _w417_ ;
	wire _w418_ ;
	wire _w419_ ;
	wire _w420_ ;
	wire _w421_ ;
	wire _w422_ ;
	wire _w423_ ;
	wire _w424_ ;
	wire _w425_ ;
	wire _w426_ ;
	wire _w427_ ;
	wire _w428_ ;
	wire _w429_ ;
	wire _w430_ ;
	wire _w431_ ;
	wire _w432_ ;
	wire _w433_ ;
	wire _w434_ ;
	wire _w435_ ;
	wire _w436_ ;
	wire _w437_ ;
	wire _w438_ ;
	wire _w439_ ;
	wire _w440_ ;
	wire _w441_ ;
	wire _w442_ ;
	wire _w443_ ;
	wire _w444_ ;
	wire _w445_ ;
	wire _w446_ ;
	wire _w447_ ;
	wire _w448_ ;
	wire _w449_ ;
	wire _w450_ ;
	wire _w451_ ;
	wire _w452_ ;
	wire _w453_ ;
	wire _w454_ ;
	wire _w455_ ;
	wire _w456_ ;
	wire _w457_ ;
	wire _w458_ ;
	wire _w459_ ;
	wire _w460_ ;
	wire _w461_ ;
	wire _w462_ ;
	wire _w463_ ;
	wire _w464_ ;
	wire _w465_ ;
	wire _w466_ ;
	wire _w467_ ;
	wire _w468_ ;
	wire _w469_ ;
	wire _w470_ ;
	wire _w471_ ;
	wire _w472_ ;
	wire _w473_ ;
	wire _w474_ ;
	wire _w475_ ;
	wire _w476_ ;
	wire _w477_ ;
	wire _w478_ ;
	wire _w479_ ;
	wire _w480_ ;
	wire _w481_ ;
	wire _w482_ ;
	wire _w483_ ;
	wire _w484_ ;
	wire _w485_ ;
	wire _w486_ ;
	wire _w487_ ;
	wire _w488_ ;
	wire _w489_ ;
	wire _w490_ ;
	wire _w491_ ;
	wire _w492_ ;
	wire _w493_ ;
	wire _w494_ ;
	wire _w495_ ;
	wire _w496_ ;
	wire _w497_ ;
	wire _w498_ ;
	wire _w499_ ;
	wire _w500_ ;
	wire _w501_ ;
	wire _w502_ ;
	wire _w503_ ;
	wire _w504_ ;
	wire _w505_ ;
	wire _w506_ ;
	wire _w507_ ;
	wire _w508_ ;
	wire _w509_ ;
	wire _w510_ ;
	wire _w511_ ;
	wire _w512_ ;
	wire _w513_ ;
	wire _w514_ ;
	wire _w515_ ;
	wire _w516_ ;
	wire _w517_ ;
	wire _w518_ ;
	wire _w519_ ;
	wire _w520_ ;
	wire _w521_ ;
	wire _w522_ ;
	wire _w523_ ;
	wire _w524_ ;
	wire _w525_ ;
	wire _w526_ ;
	wire _w527_ ;
	wire _w528_ ;
	wire _w529_ ;
	wire _w530_ ;
	wire _w531_ ;
	wire _w532_ ;
	wire _w533_ ;
	wire _w534_ ;
	wire _w535_ ;
	wire _w536_ ;
	wire _w537_ ;
	wire _w538_ ;
	wire _w539_ ;
	wire _w540_ ;
	wire _w541_ ;
	wire _w542_ ;
	wire _w543_ ;
	wire _w544_ ;
	wire _w545_ ;
	wire _w546_ ;
	wire _w547_ ;
	wire _w548_ ;
	wire _w549_ ;
	wire _w550_ ;
	wire _w551_ ;
	wire _w552_ ;
	wire _w553_ ;
	wire _w554_ ;
	wire _w555_ ;
	wire _w556_ ;
	wire _w557_ ;
	wire _w558_ ;
	wire _w559_ ;
	wire _w560_ ;
	wire _w561_ ;
	wire _w562_ ;
	wire _w563_ ;
	wire _w564_ ;
	wire _w565_ ;
	wire _w566_ ;
	wire _w567_ ;
	wire _w568_ ;
	wire _w569_ ;
	wire _w570_ ;
	wire _w571_ ;
	wire _w572_ ;
	wire _w573_ ;
	wire _w574_ ;
	wire _w575_ ;
	wire _w576_ ;
	wire _w577_ ;
	wire _w578_ ;
	wire _w579_ ;
	wire _w580_ ;
	wire _w581_ ;
	wire _w582_ ;
	wire _w583_ ;
	wire _w584_ ;
	wire _w585_ ;
	wire _w586_ ;
	wire _w587_ ;
	wire _w588_ ;
	wire _w589_ ;
	wire _w590_ ;
	wire _w591_ ;
	wire _w592_ ;
	wire _w593_ ;
	wire _w594_ ;
	wire _w595_ ;
	wire _w596_ ;
	wire _w597_ ;
	wire _w598_ ;
	wire _w599_ ;
	wire _w600_ ;
	wire _w601_ ;
	wire _w602_ ;
	wire _w603_ ;
	wire _w604_ ;
	wire _w605_ ;
	wire _w606_ ;
	wire _w607_ ;
	wire _w608_ ;
	wire _w609_ ;
	wire _w610_ ;
	wire _w611_ ;
	wire _w612_ ;
	wire _w613_ ;
	wire _w614_ ;
	wire _w615_ ;
	wire _w616_ ;
	wire _w617_ ;
	wire _w618_ ;
	wire _w619_ ;
	wire _w620_ ;
	wire _w621_ ;
	wire _w622_ ;
	wire _w623_ ;
	wire _w624_ ;
	wire _w625_ ;
	wire _w626_ ;
	wire _w627_ ;
	wire _w628_ ;
	wire _w629_ ;
	wire _w630_ ;
	wire _w631_ ;
	wire _w632_ ;
	wire _w633_ ;
	wire _w634_ ;
	wire _w635_ ;
	wire _w636_ ;
	wire _w637_ ;
	wire _w638_ ;
	wire _w639_ ;
	wire _w640_ ;
	wire _w641_ ;
	wire _w642_ ;
	wire _w643_ ;
	wire _w644_ ;
	wire _w645_ ;
	wire _w646_ ;
	wire _w647_ ;
	wire _w648_ ;
	wire _w649_ ;
	wire _w650_ ;
	wire _w651_ ;
	wire _w652_ ;
	wire _w653_ ;
	wire _w654_ ;
	wire _w655_ ;
	wire _w656_ ;
	wire _w657_ ;
	wire _w658_ ;
	wire _w659_ ;
	wire _w660_ ;
	wire _w661_ ;
	wire _w662_ ;
	wire _w663_ ;
	wire _w664_ ;
	wire _w665_ ;
	wire _w666_ ;
	wire _w667_ ;
	wire _w668_ ;
	wire _w669_ ;
	wire _w670_ ;
	wire _w671_ ;
	wire _w672_ ;
	wire _w673_ ;
	wire _w674_ ;
	wire _w675_ ;
	wire _w676_ ;
	LUT2 #(
		.INIT('h8)
	) name0 (
		i_pad,
		r_pad,
		_w136_
	);
	LUT2 #(
		.INIT('h1)
	) name1 (
		\f1_pad ,
		_w136_,
		_w137_
	);
	LUT2 #(
		.INIT('h4)
	) name2 (
		p_pad,
		_w136_,
		_w138_
	);
	LUT2 #(
		.INIT('h1)
	) name3 (
		\y1_pad ,
		_w137_,
		_w139_
	);
	LUT2 #(
		.INIT('h4)
	) name4 (
		_w138_,
		_w139_,
		_w140_
	);
	LUT2 #(
		.INIT('h8)
	) name5 (
		\a4_pad ,
		\y3_pad ,
		_w141_
	);
	LUT2 #(
		.INIT('h8)
	) name6 (
		\z3_pad ,
		_w141_,
		_w142_
	);
	LUT2 #(
		.INIT('h8)
	) name7 (
		\b4_pad ,
		_w142_,
		_w143_
	);
	LUT2 #(
		.INIT('h8)
	) name8 (
		\c4_pad ,
		_w143_,
		_w144_
	);
	LUT2 #(
		.INIT('h2)
	) name9 (
		\f4_pad ,
		\j0_pad ,
		_w145_
	);
	LUT2 #(
		.INIT('h1)
	) name10 (
		\d4_pad ,
		\h0_pad ,
		_w146_
	);
	LUT2 #(
		.INIT('h8)
	) name11 (
		\d4_pad ,
		\h0_pad ,
		_w147_
	);
	LUT2 #(
		.INIT('h4)
	) name12 (
		\f4_pad ,
		\j0_pad ,
		_w148_
	);
	LUT2 #(
		.INIT('h1)
	) name13 (
		\e4_pad ,
		\i0_pad ,
		_w149_
	);
	LUT2 #(
		.INIT('h8)
	) name14 (
		\e4_pad ,
		\i0_pad ,
		_w150_
	);
	LUT2 #(
		.INIT('h1)
	) name15 (
		_w149_,
		_w150_,
		_w151_
	);
	LUT2 #(
		.INIT('h1)
	) name16 (
		\g4_pad ,
		\k0_pad ,
		_w152_
	);
	LUT2 #(
		.INIT('h8)
	) name17 (
		\g4_pad ,
		\k0_pad ,
		_w153_
	);
	LUT2 #(
		.INIT('h1)
	) name18 (
		_w152_,
		_w153_,
		_w154_
	);
	LUT2 #(
		.INIT('h2)
	) name19 (
		\h4_pad ,
		_w145_,
		_w155_
	);
	LUT2 #(
		.INIT('h1)
	) name20 (
		_w146_,
		_w147_,
		_w156_
	);
	LUT2 #(
		.INIT('h4)
	) name21 (
		_w148_,
		_w156_,
		_w157_
	);
	LUT2 #(
		.INIT('h4)
	) name22 (
		_w151_,
		_w155_,
		_w158_
	);
	LUT2 #(
		.INIT('h4)
	) name23 (
		_w154_,
		_w158_,
		_w159_
	);
	LUT2 #(
		.INIT('h8)
	) name24 (
		_w157_,
		_w159_,
		_w160_
	);
	LUT2 #(
		.INIT('h8)
	) name25 (
		_w144_,
		_w160_,
		_w161_
	);
	LUT2 #(
		.INIT('h8)
	) name26 (
		\d2_pad ,
		\l0_pad ,
		_w162_
	);
	LUT2 #(
		.INIT('h1)
	) name27 (
		\h0_pad ,
		\i0_pad ,
		_w163_
	);
	LUT2 #(
		.INIT('h1)
	) name28 (
		\j0_pad ,
		\k0_pad ,
		_w164_
	);
	LUT2 #(
		.INIT('h8)
	) name29 (
		_w163_,
		_w164_,
		_w165_
	);
	LUT2 #(
		.INIT('h8)
	) name30 (
		_w162_,
		_w165_,
		_w166_
	);
	LUT2 #(
		.INIT('h1)
	) name31 (
		_w161_,
		_w166_,
		_w167_
	);
	LUT2 #(
		.INIT('h4)
	) name32 (
		\a2_pad ,
		_w167_,
		_w168_
	);
	LUT2 #(
		.INIT('h2)
	) name33 (
		\e2_pad ,
		_w168_,
		_w169_
	);
	LUT2 #(
		.INIT('h1)
	) name34 (
		\f2_pad ,
		_w169_,
		_w170_
	);
	LUT2 #(
		.INIT('h8)
	) name35 (
		\f2_pad ,
		_w169_,
		_w171_
	);
	LUT2 #(
		.INIT('h1)
	) name36 (
		\n0_pad ,
		_w170_,
		_w172_
	);
	LUT2 #(
		.INIT('h4)
	) name37 (
		_w171_,
		_w172_,
		_w173_
	);
	LUT2 #(
		.INIT('h8)
	) name38 (
		f_pad,
		h_pad,
		_w174_
	);
	LUT2 #(
		.INIT('h1)
	) name39 (
		\f3_pad ,
		_w174_,
		_w175_
	);
	LUT2 #(
		.INIT('h4)
	) name40 (
		\g3_pad ,
		_w174_,
		_w176_
	);
	LUT2 #(
		.INIT('h1)
	) name41 (
		\y1_pad ,
		_w175_,
		_w177_
	);
	LUT2 #(
		.INIT('h4)
	) name42 (
		_w176_,
		_w177_,
		_w178_
	);
	LUT2 #(
		.INIT('h1)
	) name43 (
		\l0_pad ,
		\n0_pad ,
		_w179_
	);
	LUT2 #(
		.INIT('h4)
	) name44 (
		\d4_pad ,
		_w144_,
		_w180_
	);
	LUT2 #(
		.INIT('h8)
	) name45 (
		\e4_pad ,
		_w180_,
		_w181_
	);
	LUT2 #(
		.INIT('h1)
	) name46 (
		\f4_pad ,
		_w181_,
		_w182_
	);
	LUT2 #(
		.INIT('h8)
	) name47 (
		\f4_pad ,
		_w181_,
		_w183_
	);
	LUT2 #(
		.INIT('h2)
	) name48 (
		_w179_,
		_w182_,
		_w184_
	);
	LUT2 #(
		.INIT('h4)
	) name49 (
		_w183_,
		_w184_,
		_w185_
	);
	LUT2 #(
		.INIT('h1)
	) name50 (
		\g1_pad ,
		_w136_,
		_w186_
	);
	LUT2 #(
		.INIT('h4)
	) name51 (
		q_pad,
		_w136_,
		_w187_
	);
	LUT2 #(
		.INIT('h1)
	) name52 (
		\y1_pad ,
		_w186_,
		_w188_
	);
	LUT2 #(
		.INIT('h4)
	) name53 (
		_w187_,
		_w188_,
		_w189_
	);
	LUT2 #(
		.INIT('h2)
	) name54 (
		\h2_pad ,
		\n0_pad ,
		_w190_
	);
	LUT2 #(
		.INIT('h1)
	) name55 (
		\g3_pad ,
		_w174_,
		_w191_
	);
	LUT2 #(
		.INIT('h4)
	) name56 (
		\h3_pad ,
		_w174_,
		_w192_
	);
	LUT2 #(
		.INIT('h1)
	) name57 (
		\y1_pad ,
		_w191_,
		_w193_
	);
	LUT2 #(
		.INIT('h4)
	) name58 (
		_w192_,
		_w193_,
		_w194_
	);
	LUT2 #(
		.INIT('h1)
	) name59 (
		\g4_pad ,
		_w183_,
		_w195_
	);
	LUT2 #(
		.INIT('h8)
	) name60 (
		\g4_pad ,
		_w183_,
		_w196_
	);
	LUT2 #(
		.INIT('h2)
	) name61 (
		_w179_,
		_w195_,
		_w197_
	);
	LUT2 #(
		.INIT('h4)
	) name62 (
		_w196_,
		_w197_,
		_w198_
	);
	LUT2 #(
		.INIT('h4)
	) name63 (
		\b0_pad ,
		s_pad,
		_w199_
	);
	LUT2 #(
		.INIT('h1)
	) name64 (
		\h1_pad ,
		_w199_,
		_w200_
	);
	LUT2 #(
		.INIT('h4)
	) name65 (
		t_pad,
		_w199_,
		_w201_
	);
	LUT2 #(
		.INIT('h1)
	) name66 (
		\y1_pad ,
		_w200_,
		_w202_
	);
	LUT2 #(
		.INIT('h4)
	) name67 (
		_w201_,
		_w202_,
		_w203_
	);
	LUT2 #(
		.INIT('h2)
	) name68 (
		\l0_pad ,
		\n0_pad ,
		_w204_
	);
	LUT2 #(
		.INIT('h1)
	) name69 (
		\h3_pad ,
		_w174_,
		_w205_
	);
	LUT2 #(
		.INIT('h4)
	) name70 (
		g_pad,
		_w174_,
		_w206_
	);
	LUT2 #(
		.INIT('h1)
	) name71 (
		\y1_pad ,
		_w205_,
		_w207_
	);
	LUT2 #(
		.INIT('h4)
	) name72 (
		_w206_,
		_w207_,
		_w208_
	);
	LUT2 #(
		.INIT('h1)
	) name73 (
		\h4_pad ,
		_w162_,
		_w209_
	);
	LUT2 #(
		.INIT('h8)
	) name74 (
		\g2_pad ,
		\h2_pad ,
		_w210_
	);
	LUT2 #(
		.INIT('h2)
	) name75 (
		b_pad,
		\n0_pad ,
		_w211_
	);
	LUT2 #(
		.INIT('h4)
	) name76 (
		_w210_,
		_w211_,
		_w212_
	);
	LUT2 #(
		.INIT('h4)
	) name77 (
		_w209_,
		_w212_,
		_w213_
	);
	LUT2 #(
		.INIT('h1)
	) name78 (
		\i1_pad ,
		_w199_,
		_w214_
	);
	LUT2 #(
		.INIT('h4)
	) name79 (
		u_pad,
		_w199_,
		_w215_
	);
	LUT2 #(
		.INIT('h1)
	) name80 (
		\y1_pad ,
		_w214_,
		_w216_
	);
	LUT2 #(
		.INIT('h4)
	) name81 (
		_w215_,
		_w216_,
		_w217_
	);
	LUT2 #(
		.INIT('h2)
	) name82 (
		\j2_pad ,
		\p2_pad ,
		_w218_
	);
	LUT2 #(
		.INIT('h2)
	) name83 (
		\o2_pad ,
		_w218_,
		_w219_
	);
	LUT2 #(
		.INIT('h2)
	) name84 (
		\l2_pad ,
		\m2_pad ,
		_w220_
	);
	LUT2 #(
		.INIT('h8)
	) name85 (
		\n2_pad ,
		_w220_,
		_w221_
	);
	LUT2 #(
		.INIT('h1)
	) name86 (
		\o2_pad ,
		\p2_pad ,
		_w222_
	);
	LUT2 #(
		.INIT('h8)
	) name87 (
		\g0_pad ,
		_w222_,
		_w223_
	);
	LUT2 #(
		.INIT('h4)
	) name88 (
		_w219_,
		_w221_,
		_w224_
	);
	LUT2 #(
		.INIT('h4)
	) name89 (
		_w223_,
		_w224_,
		_w225_
	);
	LUT2 #(
		.INIT('h4)
	) name90 (
		\x1_pad ,
		_w225_,
		_w226_
	);
	LUT2 #(
		.INIT('h1)
	) name91 (
		\i2_pad ,
		_w226_,
		_w227_
	);
	LUT2 #(
		.INIT('h1)
	) name92 (
		\y1_pad ,
		_w227_,
		_w228_
	);
	LUT2 #(
		.INIT('h2)
	) name93 (
		d_pad,
		e_pad,
		_w229_
	);
	LUT2 #(
		.INIT('h4)
	) name94 (
		\r0_pad ,
		_w229_,
		_w230_
	);
	LUT2 #(
		.INIT('h1)
	) name95 (
		\j2_pad ,
		\k2_pad ,
		_w231_
	);
	LUT2 #(
		.INIT('h1)
	) name96 (
		\x1_pad ,
		_w231_,
		_w232_
	);
	LUT2 #(
		.INIT('h8)
	) name97 (
		\j3_pad ,
		_w232_,
		_w233_
	);
	LUT2 #(
		.INIT('h1)
	) name98 (
		c_pad,
		d_pad,
		_w234_
	);
	LUT2 #(
		.INIT('h4)
	) name99 (
		e_pad,
		_w234_,
		_w235_
	);
	LUT2 #(
		.INIT('h2)
	) name100 (
		\i3_pad ,
		_w232_,
		_w236_
	);
	LUT2 #(
		.INIT('h4)
	) name101 (
		_w233_,
		_w235_,
		_w237_
	);
	LUT2 #(
		.INIT('h4)
	) name102 (
		_w236_,
		_w237_,
		_w238_
	);
	LUT2 #(
		.INIT('h2)
	) name103 (
		e_pad,
		\h1_pad ,
		_w239_
	);
	LUT2 #(
		.INIT('h2)
	) name104 (
		c_pad,
		d_pad,
		_w240_
	);
	LUT2 #(
		.INIT('h4)
	) name105 (
		e_pad,
		_w240_,
		_w241_
	);
	LUT2 #(
		.INIT('h4)
	) name106 (
		\s2_pad ,
		_w241_,
		_w242_
	);
	LUT2 #(
		.INIT('h1)
	) name107 (
		\y1_pad ,
		_w239_,
		_w243_
	);
	LUT2 #(
		.INIT('h4)
	) name108 (
		_w230_,
		_w243_,
		_w244_
	);
	LUT2 #(
		.INIT('h4)
	) name109 (
		_w242_,
		_w244_,
		_w245_
	);
	LUT2 #(
		.INIT('h4)
	) name110 (
		_w238_,
		_w245_,
		_w246_
	);
	LUT2 #(
		.INIT('h1)
	) name111 (
		\j1_pad ,
		_w199_,
		_w247_
	);
	LUT2 #(
		.INIT('h4)
	) name112 (
		v_pad,
		_w199_,
		_w248_
	);
	LUT2 #(
		.INIT('h1)
	) name113 (
		\y1_pad ,
		_w247_,
		_w249_
	);
	LUT2 #(
		.INIT('h4)
	) name114 (
		_w248_,
		_w249_,
		_w250_
	);
	LUT2 #(
		.INIT('h1)
	) name115 (
		\j2_pad ,
		\o2_pad ,
		_w251_
	);
	LUT2 #(
		.INIT('h1)
	) name116 (
		\e0_pad ,
		\f0_pad ,
		_w252_
	);
	LUT2 #(
		.INIT('h2)
	) name117 (
		\g0_pad ,
		_w252_,
		_w253_
	);
	LUT2 #(
		.INIT('h1)
	) name118 (
		\o2_pad ,
		_w253_,
		_w254_
	);
	LUT2 #(
		.INIT('h1)
	) name119 (
		\p2_pad ,
		\x1_pad ,
		_w255_
	);
	LUT2 #(
		.INIT('h8)
	) name120 (
		_w221_,
		_w255_,
		_w256_
	);
	LUT2 #(
		.INIT('h4)
	) name121 (
		_w254_,
		_w256_,
		_w257_
	);
	LUT2 #(
		.INIT('h4)
	) name122 (
		_w251_,
		_w257_,
		_w258_
	);
	LUT2 #(
		.INIT('h1)
	) name123 (
		\j2_pad ,
		_w257_,
		_w259_
	);
	LUT2 #(
		.INIT('h1)
	) name124 (
		\y1_pad ,
		_w258_,
		_w260_
	);
	LUT2 #(
		.INIT('h4)
	) name125 (
		_w259_,
		_w260_,
		_w261_
	);
	LUT2 #(
		.INIT('h4)
	) name126 (
		\s0_pad ,
		_w229_,
		_w262_
	);
	LUT2 #(
		.INIT('h8)
	) name127 (
		\k3_pad ,
		_w232_,
		_w263_
	);
	LUT2 #(
		.INIT('h2)
	) name128 (
		\j3_pad ,
		_w232_,
		_w264_
	);
	LUT2 #(
		.INIT('h2)
	) name129 (
		_w235_,
		_w263_,
		_w265_
	);
	LUT2 #(
		.INIT('h4)
	) name130 (
		_w264_,
		_w265_,
		_w266_
	);
	LUT2 #(
		.INIT('h2)
	) name131 (
		e_pad,
		\i1_pad ,
		_w267_
	);
	LUT2 #(
		.INIT('h4)
	) name132 (
		\t2_pad ,
		_w241_,
		_w268_
	);
	LUT2 #(
		.INIT('h1)
	) name133 (
		\y1_pad ,
		_w267_,
		_w269_
	);
	LUT2 #(
		.INIT('h4)
	) name134 (
		_w262_,
		_w269_,
		_w270_
	);
	LUT2 #(
		.INIT('h4)
	) name135 (
		_w268_,
		_w270_,
		_w271_
	);
	LUT2 #(
		.INIT('h4)
	) name136 (
		_w266_,
		_w271_,
		_w272_
	);
	LUT2 #(
		.INIT('h1)
	) name137 (
		\k1_pad ,
		_w199_,
		_w273_
	);
	LUT2 #(
		.INIT('h4)
	) name138 (
		w_pad,
		_w199_,
		_w274_
	);
	LUT2 #(
		.INIT('h1)
	) name139 (
		\y1_pad ,
		_w273_,
		_w275_
	);
	LUT2 #(
		.INIT('h4)
	) name140 (
		_w274_,
		_w275_,
		_w276_
	);
	LUT2 #(
		.INIT('h8)
	) name141 (
		\g0_pad ,
		_w252_,
		_w277_
	);
	LUT2 #(
		.INIT('h1)
	) name142 (
		\p2_pad ,
		_w277_,
		_w278_
	);
	LUT2 #(
		.INIT('h1)
	) name143 (
		\o2_pad ,
		\x1_pad ,
		_w279_
	);
	LUT2 #(
		.INIT('h8)
	) name144 (
		_w221_,
		_w279_,
		_w280_
	);
	LUT2 #(
		.INIT('h4)
	) name145 (
		_w278_,
		_w280_,
		_w281_
	);
	LUT2 #(
		.INIT('h1)
	) name146 (
		\k2_pad ,
		_w281_,
		_w282_
	);
	LUT2 #(
		.INIT('h8)
	) name147 (
		\k2_pad ,
		_w281_,
		_w283_
	);
	LUT2 #(
		.INIT('h1)
	) name148 (
		\y1_pad ,
		_w282_,
		_w284_
	);
	LUT2 #(
		.INIT('h4)
	) name149 (
		_w283_,
		_w284_,
		_w285_
	);
	LUT2 #(
		.INIT('h4)
	) name150 (
		\t0_pad ,
		_w229_,
		_w286_
	);
	LUT2 #(
		.INIT('h8)
	) name151 (
		\l3_pad ,
		_w232_,
		_w287_
	);
	LUT2 #(
		.INIT('h2)
	) name152 (
		\k3_pad ,
		_w232_,
		_w288_
	);
	LUT2 #(
		.INIT('h2)
	) name153 (
		_w235_,
		_w287_,
		_w289_
	);
	LUT2 #(
		.INIT('h4)
	) name154 (
		_w288_,
		_w289_,
		_w290_
	);
	LUT2 #(
		.INIT('h2)
	) name155 (
		e_pad,
		\j1_pad ,
		_w291_
	);
	LUT2 #(
		.INIT('h4)
	) name156 (
		\u2_pad ,
		_w241_,
		_w292_
	);
	LUT2 #(
		.INIT('h1)
	) name157 (
		\y1_pad ,
		_w291_,
		_w293_
	);
	LUT2 #(
		.INIT('h4)
	) name158 (
		_w286_,
		_w293_,
		_w294_
	);
	LUT2 #(
		.INIT('h4)
	) name159 (
		_w292_,
		_w294_,
		_w295_
	);
	LUT2 #(
		.INIT('h4)
	) name160 (
		_w290_,
		_w295_,
		_w296_
	);
	LUT2 #(
		.INIT('h1)
	) name161 (
		\l1_pad ,
		_w199_,
		_w297_
	);
	LUT2 #(
		.INIT('h4)
	) name162 (
		x_pad,
		_w199_,
		_w298_
	);
	LUT2 #(
		.INIT('h1)
	) name163 (
		\y1_pad ,
		_w297_,
		_w299_
	);
	LUT2 #(
		.INIT('h4)
	) name164 (
		_w298_,
		_w299_,
		_w300_
	);
	LUT2 #(
		.INIT('h8)
	) name165 (
		\x1_pad ,
		_w235_,
		_w301_
	);
	LUT2 #(
		.INIT('h2)
	) name166 (
		\l2_pad ,
		_w301_,
		_w302_
	);
	LUT2 #(
		.INIT('h4)
	) name167 (
		\l2_pad ,
		_w301_,
		_w303_
	);
	LUT2 #(
		.INIT('h1)
	) name168 (
		\y1_pad ,
		_w302_,
		_w304_
	);
	LUT2 #(
		.INIT('h4)
	) name169 (
		_w303_,
		_w304_,
		_w305_
	);
	LUT2 #(
		.INIT('h4)
	) name170 (
		\u0_pad ,
		_w229_,
		_w306_
	);
	LUT2 #(
		.INIT('h8)
	) name171 (
		\m3_pad ,
		_w232_,
		_w307_
	);
	LUT2 #(
		.INIT('h2)
	) name172 (
		\l3_pad ,
		_w232_,
		_w308_
	);
	LUT2 #(
		.INIT('h2)
	) name173 (
		_w235_,
		_w307_,
		_w309_
	);
	LUT2 #(
		.INIT('h4)
	) name174 (
		_w308_,
		_w309_,
		_w310_
	);
	LUT2 #(
		.INIT('h2)
	) name175 (
		e_pad,
		\k1_pad ,
		_w311_
	);
	LUT2 #(
		.INIT('h4)
	) name176 (
		\v2_pad ,
		_w241_,
		_w312_
	);
	LUT2 #(
		.INIT('h1)
	) name177 (
		\y1_pad ,
		_w311_,
		_w313_
	);
	LUT2 #(
		.INIT('h4)
	) name178 (
		_w306_,
		_w313_,
		_w314_
	);
	LUT2 #(
		.INIT('h4)
	) name179 (
		_w312_,
		_w314_,
		_w315_
	);
	LUT2 #(
		.INIT('h4)
	) name180 (
		_w310_,
		_w315_,
		_w316_
	);
	LUT2 #(
		.INIT('h1)
	) name181 (
		\m1_pad ,
		_w199_,
		_w317_
	);
	LUT2 #(
		.INIT('h4)
	) name182 (
		y_pad,
		_w199_,
		_w318_
	);
	LUT2 #(
		.INIT('h1)
	) name183 (
		\y1_pad ,
		_w317_,
		_w319_
	);
	LUT2 #(
		.INIT('h4)
	) name184 (
		_w318_,
		_w319_,
		_w320_
	);
	LUT2 #(
		.INIT('h1)
	) name185 (
		\m2_pad ,
		_w302_,
		_w321_
	);
	LUT2 #(
		.INIT('h8)
	) name186 (
		\m2_pad ,
		_w302_,
		_w322_
	);
	LUT2 #(
		.INIT('h1)
	) name187 (
		\y1_pad ,
		_w321_,
		_w323_
	);
	LUT2 #(
		.INIT('h4)
	) name188 (
		_w322_,
		_w323_,
		_w324_
	);
	LUT2 #(
		.INIT('h4)
	) name189 (
		\v0_pad ,
		_w229_,
		_w325_
	);
	LUT2 #(
		.INIT('h8)
	) name190 (
		\n3_pad ,
		_w232_,
		_w326_
	);
	LUT2 #(
		.INIT('h2)
	) name191 (
		\m3_pad ,
		_w232_,
		_w327_
	);
	LUT2 #(
		.INIT('h2)
	) name192 (
		_w235_,
		_w326_,
		_w328_
	);
	LUT2 #(
		.INIT('h4)
	) name193 (
		_w327_,
		_w328_,
		_w329_
	);
	LUT2 #(
		.INIT('h2)
	) name194 (
		e_pad,
		\l1_pad ,
		_w330_
	);
	LUT2 #(
		.INIT('h4)
	) name195 (
		\w2_pad ,
		_w241_,
		_w331_
	);
	LUT2 #(
		.INIT('h1)
	) name196 (
		\y1_pad ,
		_w330_,
		_w332_
	);
	LUT2 #(
		.INIT('h4)
	) name197 (
		_w325_,
		_w332_,
		_w333_
	);
	LUT2 #(
		.INIT('h4)
	) name198 (
		_w331_,
		_w333_,
		_w334_
	);
	LUT2 #(
		.INIT('h4)
	) name199 (
		_w329_,
		_w334_,
		_w335_
	);
	LUT2 #(
		.INIT('h4)
	) name200 (
		\a2_pad ,
		\x1_pad ,
		_w336_
	);
	LUT2 #(
		.INIT('h1)
	) name201 (
		\n1_pad ,
		_w199_,
		_w337_
	);
	LUT2 #(
		.INIT('h4)
	) name202 (
		z_pad,
		_w199_,
		_w338_
	);
	LUT2 #(
		.INIT('h1)
	) name203 (
		\y1_pad ,
		_w337_,
		_w339_
	);
	LUT2 #(
		.INIT('h4)
	) name204 (
		_w338_,
		_w339_,
		_w340_
	);
	LUT2 #(
		.INIT('h1)
	) name205 (
		\n2_pad ,
		_w322_,
		_w341_
	);
	LUT2 #(
		.INIT('h8)
	) name206 (
		\n2_pad ,
		_w322_,
		_w342_
	);
	LUT2 #(
		.INIT('h1)
	) name207 (
		\y1_pad ,
		_w341_,
		_w343_
	);
	LUT2 #(
		.INIT('h4)
	) name208 (
		_w342_,
		_w343_,
		_w344_
	);
	LUT2 #(
		.INIT('h4)
	) name209 (
		\w0_pad ,
		_w229_,
		_w345_
	);
	LUT2 #(
		.INIT('h8)
	) name210 (
		\o3_pad ,
		_w232_,
		_w346_
	);
	LUT2 #(
		.INIT('h2)
	) name211 (
		\n3_pad ,
		_w232_,
		_w347_
	);
	LUT2 #(
		.INIT('h2)
	) name212 (
		_w235_,
		_w346_,
		_w348_
	);
	LUT2 #(
		.INIT('h4)
	) name213 (
		_w347_,
		_w348_,
		_w349_
	);
	LUT2 #(
		.INIT('h2)
	) name214 (
		e_pad,
		\m1_pad ,
		_w350_
	);
	LUT2 #(
		.INIT('h4)
	) name215 (
		\x2_pad ,
		_w241_,
		_w351_
	);
	LUT2 #(
		.INIT('h1)
	) name216 (
		\y1_pad ,
		_w350_,
		_w352_
	);
	LUT2 #(
		.INIT('h4)
	) name217 (
		_w345_,
		_w352_,
		_w353_
	);
	LUT2 #(
		.INIT('h4)
	) name218 (
		_w351_,
		_w353_,
		_w354_
	);
	LUT2 #(
		.INIT('h4)
	) name219 (
		_w349_,
		_w354_,
		_w355_
	);
	LUT2 #(
		.INIT('h8)
	) name220 (
		\i2_pad ,
		\r2_pad ,
		_w356_
	);
	LUT2 #(
		.INIT('h2)
	) name221 (
		\q2_pad ,
		\x1_pad ,
		_w357_
	);
	LUT2 #(
		.INIT('h8)
	) name222 (
		_w356_,
		_w357_,
		_w358_
	);
	LUT2 #(
		.INIT('h1)
	) name223 (
		\o0_pad ,
		_w358_,
		_w359_
	);
	LUT2 #(
		.INIT('h2)
	) name224 (
		_w235_,
		_w359_,
		_w360_
	);
	LUT2 #(
		.INIT('h1)
	) name225 (
		\y1_pad ,
		_w360_,
		_w361_
	);
	LUT2 #(
		.INIT('h1)
	) name226 (
		\o1_pad ,
		_w199_,
		_w362_
	);
	LUT2 #(
		.INIT('h4)
	) name227 (
		\a0_pad ,
		_w199_,
		_w363_
	);
	LUT2 #(
		.INIT('h1)
	) name228 (
		\y1_pad ,
		_w362_,
		_w364_
	);
	LUT2 #(
		.INIT('h4)
	) name229 (
		_w363_,
		_w364_,
		_w365_
	);
	LUT2 #(
		.INIT('h1)
	) name230 (
		\o2_pad ,
		_w342_,
		_w366_
	);
	LUT2 #(
		.INIT('h8)
	) name231 (
		\o2_pad ,
		_w342_,
		_w367_
	);
	LUT2 #(
		.INIT('h1)
	) name232 (
		\y1_pad ,
		_w366_,
		_w368_
	);
	LUT2 #(
		.INIT('h4)
	) name233 (
		_w367_,
		_w368_,
		_w369_
	);
	LUT2 #(
		.INIT('h4)
	) name234 (
		\x0_pad ,
		_w229_,
		_w370_
	);
	LUT2 #(
		.INIT('h8)
	) name235 (
		\p3_pad ,
		_w232_,
		_w371_
	);
	LUT2 #(
		.INIT('h2)
	) name236 (
		\o3_pad ,
		_w232_,
		_w372_
	);
	LUT2 #(
		.INIT('h2)
	) name237 (
		_w235_,
		_w371_,
		_w373_
	);
	LUT2 #(
		.INIT('h4)
	) name238 (
		_w372_,
		_w373_,
		_w374_
	);
	LUT2 #(
		.INIT('h2)
	) name239 (
		e_pad,
		\n1_pad ,
		_w375_
	);
	LUT2 #(
		.INIT('h4)
	) name240 (
		\y2_pad ,
		_w241_,
		_w376_
	);
	LUT2 #(
		.INIT('h1)
	) name241 (
		\y1_pad ,
		_w375_,
		_w377_
	);
	LUT2 #(
		.INIT('h4)
	) name242 (
		_w370_,
		_w377_,
		_w378_
	);
	LUT2 #(
		.INIT('h4)
	) name243 (
		_w376_,
		_w378_,
		_w379_
	);
	LUT2 #(
		.INIT('h4)
	) name244 (
		_w374_,
		_w379_,
		_w380_
	);
	LUT2 #(
		.INIT('h1)
	) name245 (
		\q2_pad ,
		\r2_pad ,
		_w381_
	);
	LUT2 #(
		.INIT('h2)
	) name246 (
		\i2_pad ,
		_w381_,
		_w382_
	);
	LUT2 #(
		.INIT('h2)
	) name247 (
		_w231_,
		_w382_,
		_w383_
	);
	LUT2 #(
		.INIT('h1)
	) name248 (
		\x1_pad ,
		_w383_,
		_w384_
	);
	LUT2 #(
		.INIT('h8)
	) name249 (
		\d0_pad ,
		\r2_pad ,
		_w385_
	);
	LUT2 #(
		.INIT('h1)
	) name250 (
		\q2_pad ,
		_w385_,
		_w386_
	);
	LUT2 #(
		.INIT('h2)
	) name251 (
		\i2_pad ,
		_w386_,
		_w387_
	);
	LUT2 #(
		.INIT('h2)
	) name252 (
		\i3_pad ,
		_w356_,
		_w388_
	);
	LUT2 #(
		.INIT('h1)
	) name253 (
		_w387_,
		_w388_,
		_w389_
	);
	LUT2 #(
		.INIT('h2)
	) name254 (
		\r2_pad ,
		\z1_pad ,
		_w390_
	);
	LUT2 #(
		.INIT('h1)
	) name255 (
		\c0_pad ,
		\r2_pad ,
		_w391_
	);
	LUT2 #(
		.INIT('h8)
	) name256 (
		\i2_pad ,
		\q2_pad ,
		_w392_
	);
	LUT2 #(
		.INIT('h4)
	) name257 (
		_w390_,
		_w392_,
		_w393_
	);
	LUT2 #(
		.INIT('h4)
	) name258 (
		_w391_,
		_w393_,
		_w394_
	);
	LUT2 #(
		.INIT('h1)
	) name259 (
		_w389_,
		_w394_,
		_w395_
	);
	LUT2 #(
		.INIT('h2)
	) name260 (
		_w384_,
		_w395_,
		_w396_
	);
	LUT2 #(
		.INIT('h1)
	) name261 (
		\i0_pad ,
		\l2_pad ,
		_w397_
	);
	LUT2 #(
		.INIT('h4)
	) name262 (
		\h0_pad ,
		\l2_pad ,
		_w398_
	);
	LUT2 #(
		.INIT('h2)
	) name263 (
		\n2_pad ,
		_w397_,
		_w399_
	);
	LUT2 #(
		.INIT('h4)
	) name264 (
		_w398_,
		_w399_,
		_w400_
	);
	LUT2 #(
		.INIT('h1)
	) name265 (
		\m2_pad ,
		_w400_,
		_w401_
	);
	LUT2 #(
		.INIT('h1)
	) name266 (
		\k0_pad ,
		\l2_pad ,
		_w402_
	);
	LUT2 #(
		.INIT('h4)
	) name267 (
		\j0_pad ,
		\l2_pad ,
		_w403_
	);
	LUT2 #(
		.INIT('h1)
	) name268 (
		\n2_pad ,
		_w402_,
		_w404_
	);
	LUT2 #(
		.INIT('h4)
	) name269 (
		_w403_,
		_w404_,
		_w405_
	);
	LUT2 #(
		.INIT('h2)
	) name270 (
		\m2_pad ,
		_w405_,
		_w406_
	);
	LUT2 #(
		.INIT('h2)
	) name271 (
		_w222_,
		_w401_,
		_w407_
	);
	LUT2 #(
		.INIT('h4)
	) name272 (
		_w406_,
		_w407_,
		_w408_
	);
	LUT2 #(
		.INIT('h1)
	) name273 (
		_w384_,
		_w408_,
		_w409_
	);
	LUT2 #(
		.INIT('h1)
	) name274 (
		\a2_pad ,
		\y1_pad ,
		_w410_
	);
	LUT2 #(
		.INIT('h4)
	) name275 (
		_w396_,
		_w410_,
		_w411_
	);
	LUT2 #(
		.INIT('h4)
	) name276 (
		_w409_,
		_w411_,
		_w412_
	);
	LUT2 #(
		.INIT('h2)
	) name277 (
		\d0_pad ,
		\f2_pad ,
		_w413_
	);
	LUT2 #(
		.INIT('h8)
	) name278 (
		\e2_pad ,
		\f2_pad ,
		_w414_
	);
	LUT2 #(
		.INIT('h2)
	) name279 (
		\a2_pad ,
		_w414_,
		_w415_
	);
	LUT2 #(
		.INIT('h1)
	) name280 (
		\d0_pad ,
		\e2_pad ,
		_w416_
	);
	LUT2 #(
		.INIT('h2)
	) name281 (
		\m0_pad ,
		\y1_pad ,
		_w417_
	);
	LUT2 #(
		.INIT('h4)
	) name282 (
		_w413_,
		_w417_,
		_w418_
	);
	LUT2 #(
		.INIT('h4)
	) name283 (
		_w416_,
		_w418_,
		_w419_
	);
	LUT2 #(
		.INIT('h8)
	) name284 (
		_w415_,
		_w419_,
		_w420_
	);
	LUT2 #(
		.INIT('h1)
	) name285 (
		_w412_,
		_w420_,
		_w421_
	);
	LUT2 #(
		.INIT('h8)
	) name286 (
		\b0_pad ,
		s_pad,
		_w422_
	);
	LUT2 #(
		.INIT('h1)
	) name287 (
		\p1_pad ,
		_w422_,
		_w423_
	);
	LUT2 #(
		.INIT('h4)
	) name288 (
		t_pad,
		_w422_,
		_w424_
	);
	LUT2 #(
		.INIT('h1)
	) name289 (
		\y1_pad ,
		_w423_,
		_w425_
	);
	LUT2 #(
		.INIT('h4)
	) name290 (
		_w424_,
		_w425_,
		_w426_
	);
	LUT2 #(
		.INIT('h1)
	) name291 (
		\p2_pad ,
		_w367_,
		_w427_
	);
	LUT2 #(
		.INIT('h8)
	) name292 (
		\p2_pad ,
		_w367_,
		_w428_
	);
	LUT2 #(
		.INIT('h1)
	) name293 (
		\y1_pad ,
		_w427_,
		_w429_
	);
	LUT2 #(
		.INIT('h4)
	) name294 (
		_w428_,
		_w429_,
		_w430_
	);
	LUT2 #(
		.INIT('h4)
	) name295 (
		\y0_pad ,
		_w229_,
		_w431_
	);
	LUT2 #(
		.INIT('h8)
	) name296 (
		\q3_pad ,
		_w232_,
		_w432_
	);
	LUT2 #(
		.INIT('h2)
	) name297 (
		\p3_pad ,
		_w232_,
		_w433_
	);
	LUT2 #(
		.INIT('h2)
	) name298 (
		_w235_,
		_w432_,
		_w434_
	);
	LUT2 #(
		.INIT('h4)
	) name299 (
		_w433_,
		_w434_,
		_w435_
	);
	LUT2 #(
		.INIT('h2)
	) name300 (
		e_pad,
		\o1_pad ,
		_w436_
	);
	LUT2 #(
		.INIT('h4)
	) name301 (
		\z2_pad ,
		_w241_,
		_w437_
	);
	LUT2 #(
		.INIT('h1)
	) name302 (
		\y1_pad ,
		_w436_,
		_w438_
	);
	LUT2 #(
		.INIT('h4)
	) name303 (
		_w431_,
		_w438_,
		_w439_
	);
	LUT2 #(
		.INIT('h4)
	) name304 (
		_w437_,
		_w439_,
		_w440_
	);
	LUT2 #(
		.INIT('h4)
	) name305 (
		_w435_,
		_w440_,
		_w441_
	);
	LUT2 #(
		.INIT('h1)
	) name306 (
		\c2_pad ,
		_w210_,
		_w442_
	);
	LUT2 #(
		.INIT('h1)
	) name307 (
		\n0_pad ,
		_w442_,
		_w443_
	);
	LUT2 #(
		.INIT('h1)
	) name308 (
		\q1_pad ,
		_w422_,
		_w444_
	);
	LUT2 #(
		.INIT('h4)
	) name309 (
		u_pad,
		_w422_,
		_w445_
	);
	LUT2 #(
		.INIT('h1)
	) name310 (
		\y1_pad ,
		_w444_,
		_w446_
	);
	LUT2 #(
		.INIT('h4)
	) name311 (
		_w445_,
		_w446_,
		_w447_
	);
	LUT2 #(
		.INIT('h1)
	) name312 (
		\i2_pad ,
		_w225_,
		_w448_
	);
	LUT2 #(
		.INIT('h1)
	) name313 (
		\x1_pad ,
		_w448_,
		_w449_
	);
	LUT2 #(
		.INIT('h8)
	) name314 (
		\q2_pad ,
		_w449_,
		_w450_
	);
	LUT2 #(
		.INIT('h1)
	) name315 (
		\q2_pad ,
		_w449_,
		_w451_
	);
	LUT2 #(
		.INIT('h1)
	) name316 (
		\y1_pad ,
		_w450_,
		_w452_
	);
	LUT2 #(
		.INIT('h4)
	) name317 (
		_w451_,
		_w452_,
		_w453_
	);
	LUT2 #(
		.INIT('h4)
	) name318 (
		\z0_pad ,
		_w229_,
		_w454_
	);
	LUT2 #(
		.INIT('h8)
	) name319 (
		\r3_pad ,
		_w232_,
		_w455_
	);
	LUT2 #(
		.INIT('h2)
	) name320 (
		\q3_pad ,
		_w232_,
		_w456_
	);
	LUT2 #(
		.INIT('h2)
	) name321 (
		_w235_,
		_w455_,
		_w457_
	);
	LUT2 #(
		.INIT('h4)
	) name322 (
		_w456_,
		_w457_,
		_w458_
	);
	LUT2 #(
		.INIT('h2)
	) name323 (
		e_pad,
		\p1_pad ,
		_w459_
	);
	LUT2 #(
		.INIT('h4)
	) name324 (
		\a3_pad ,
		_w241_,
		_w460_
	);
	LUT2 #(
		.INIT('h1)
	) name325 (
		\y1_pad ,
		_w459_,
		_w461_
	);
	LUT2 #(
		.INIT('h4)
	) name326 (
		_w454_,
		_w461_,
		_w462_
	);
	LUT2 #(
		.INIT('h4)
	) name327 (
		_w460_,
		_w462_,
		_w463_
	);
	LUT2 #(
		.INIT('h4)
	) name328 (
		_w458_,
		_w463_,
		_w464_
	);
	LUT2 #(
		.INIT('h2)
	) name329 (
		i_pad,
		r_pad,
		_w465_
	);
	LUT2 #(
		.INIT('h1)
	) name330 (
		\r0_pad ,
		_w465_,
		_w466_
	);
	LUT2 #(
		.INIT('h4)
	) name331 (
		j_pad,
		_w465_,
		_w467_
	);
	LUT2 #(
		.INIT('h1)
	) name332 (
		\y1_pad ,
		_w466_,
		_w468_
	);
	LUT2 #(
		.INIT('h4)
	) name333 (
		_w467_,
		_w468_,
		_w469_
	);
	LUT2 #(
		.INIT('h1)
	) name334 (
		\r1_pad ,
		_w422_,
		_w470_
	);
	LUT2 #(
		.INIT('h4)
	) name335 (
		v_pad,
		_w422_,
		_w471_
	);
	LUT2 #(
		.INIT('h1)
	) name336 (
		\y1_pad ,
		_w470_,
		_w472_
	);
	LUT2 #(
		.INIT('h4)
	) name337 (
		_w471_,
		_w472_,
		_w473_
	);
	LUT2 #(
		.INIT('h1)
	) name338 (
		\r2_pad ,
		_w450_,
		_w474_
	);
	LUT2 #(
		.INIT('h8)
	) name339 (
		\r2_pad ,
		_w450_,
		_w475_
	);
	LUT2 #(
		.INIT('h1)
	) name340 (
		\y1_pad ,
		_w474_,
		_w476_
	);
	LUT2 #(
		.INIT('h4)
	) name341 (
		_w475_,
		_w476_,
		_w477_
	);
	LUT2 #(
		.INIT('h4)
	) name342 (
		\a1_pad ,
		_w229_,
		_w478_
	);
	LUT2 #(
		.INIT('h8)
	) name343 (
		\s3_pad ,
		_w232_,
		_w479_
	);
	LUT2 #(
		.INIT('h2)
	) name344 (
		\r3_pad ,
		_w232_,
		_w480_
	);
	LUT2 #(
		.INIT('h2)
	) name345 (
		_w235_,
		_w479_,
		_w481_
	);
	LUT2 #(
		.INIT('h4)
	) name346 (
		_w480_,
		_w481_,
		_w482_
	);
	LUT2 #(
		.INIT('h2)
	) name347 (
		e_pad,
		\q1_pad ,
		_w483_
	);
	LUT2 #(
		.INIT('h4)
	) name348 (
		\b3_pad ,
		_w241_,
		_w484_
	);
	LUT2 #(
		.INIT('h1)
	) name349 (
		\y1_pad ,
		_w483_,
		_w485_
	);
	LUT2 #(
		.INIT('h4)
	) name350 (
		_w478_,
		_w485_,
		_w486_
	);
	LUT2 #(
		.INIT('h4)
	) name351 (
		_w484_,
		_w486_,
		_w487_
	);
	LUT2 #(
		.INIT('h4)
	) name352 (
		_w482_,
		_w487_,
		_w488_
	);
	LUT2 #(
		.INIT('h1)
	) name353 (
		\s0_pad ,
		_w465_,
		_w489_
	);
	LUT2 #(
		.INIT('h4)
	) name354 (
		k_pad,
		_w465_,
		_w490_
	);
	LUT2 #(
		.INIT('h1)
	) name355 (
		\y1_pad ,
		_w489_,
		_w491_
	);
	LUT2 #(
		.INIT('h4)
	) name356 (
		_w490_,
		_w491_,
		_w492_
	);
	LUT2 #(
		.INIT('h1)
	) name357 (
		\s1_pad ,
		_w422_,
		_w493_
	);
	LUT2 #(
		.INIT('h4)
	) name358 (
		w_pad,
		_w422_,
		_w494_
	);
	LUT2 #(
		.INIT('h1)
	) name359 (
		\y1_pad ,
		_w493_,
		_w495_
	);
	LUT2 #(
		.INIT('h4)
	) name360 (
		_w494_,
		_w495_,
		_w496_
	);
	LUT2 #(
		.INIT('h2)
	) name361 (
		f_pad,
		h_pad,
		_w497_
	);
	LUT2 #(
		.INIT('h1)
	) name362 (
		\s2_pad ,
		_w497_,
		_w498_
	);
	LUT2 #(
		.INIT('h4)
	) name363 (
		\t2_pad ,
		_w497_,
		_w499_
	);
	LUT2 #(
		.INIT('h1)
	) name364 (
		\y1_pad ,
		_w498_,
		_w500_
	);
	LUT2 #(
		.INIT('h4)
	) name365 (
		_w499_,
		_w500_,
		_w501_
	);
	LUT2 #(
		.INIT('h4)
	) name366 (
		\b1_pad ,
		_w229_,
		_w502_
	);
	LUT2 #(
		.INIT('h8)
	) name367 (
		\t3_pad ,
		_w232_,
		_w503_
	);
	LUT2 #(
		.INIT('h2)
	) name368 (
		\s3_pad ,
		_w232_,
		_w504_
	);
	LUT2 #(
		.INIT('h2)
	) name369 (
		_w235_,
		_w503_,
		_w505_
	);
	LUT2 #(
		.INIT('h4)
	) name370 (
		_w504_,
		_w505_,
		_w506_
	);
	LUT2 #(
		.INIT('h2)
	) name371 (
		e_pad,
		\r1_pad ,
		_w507_
	);
	LUT2 #(
		.INIT('h4)
	) name372 (
		\c3_pad ,
		_w241_,
		_w508_
	);
	LUT2 #(
		.INIT('h1)
	) name373 (
		\y1_pad ,
		_w507_,
		_w509_
	);
	LUT2 #(
		.INIT('h4)
	) name374 (
		_w502_,
		_w509_,
		_w510_
	);
	LUT2 #(
		.INIT('h4)
	) name375 (
		_w508_,
		_w510_,
		_w511_
	);
	LUT2 #(
		.INIT('h4)
	) name376 (
		_w506_,
		_w511_,
		_w512_
	);
	LUT2 #(
		.INIT('h1)
	) name377 (
		\t0_pad ,
		_w465_,
		_w513_
	);
	LUT2 #(
		.INIT('h4)
	) name378 (
		l_pad,
		_w465_,
		_w514_
	);
	LUT2 #(
		.INIT('h1)
	) name379 (
		\y1_pad ,
		_w513_,
		_w515_
	);
	LUT2 #(
		.INIT('h4)
	) name380 (
		_w514_,
		_w515_,
		_w516_
	);
	LUT2 #(
		.INIT('h1)
	) name381 (
		\t1_pad ,
		_w422_,
		_w517_
	);
	LUT2 #(
		.INIT('h4)
	) name382 (
		x_pad,
		_w422_,
		_w518_
	);
	LUT2 #(
		.INIT('h1)
	) name383 (
		\y1_pad ,
		_w517_,
		_w519_
	);
	LUT2 #(
		.INIT('h4)
	) name384 (
		_w518_,
		_w519_,
		_w520_
	);
	LUT2 #(
		.INIT('h1)
	) name385 (
		\t2_pad ,
		_w497_,
		_w521_
	);
	LUT2 #(
		.INIT('h4)
	) name386 (
		\u2_pad ,
		_w497_,
		_w522_
	);
	LUT2 #(
		.INIT('h1)
	) name387 (
		\y1_pad ,
		_w521_,
		_w523_
	);
	LUT2 #(
		.INIT('h4)
	) name388 (
		_w522_,
		_w523_,
		_w524_
	);
	LUT2 #(
		.INIT('h4)
	) name389 (
		\c1_pad ,
		_w229_,
		_w525_
	);
	LUT2 #(
		.INIT('h8)
	) name390 (
		\u3_pad ,
		_w232_,
		_w526_
	);
	LUT2 #(
		.INIT('h2)
	) name391 (
		\t3_pad ,
		_w232_,
		_w527_
	);
	LUT2 #(
		.INIT('h2)
	) name392 (
		_w235_,
		_w526_,
		_w528_
	);
	LUT2 #(
		.INIT('h4)
	) name393 (
		_w527_,
		_w528_,
		_w529_
	);
	LUT2 #(
		.INIT('h2)
	) name394 (
		e_pad,
		\s1_pad ,
		_w530_
	);
	LUT2 #(
		.INIT('h4)
	) name395 (
		\d3_pad ,
		_w241_,
		_w531_
	);
	LUT2 #(
		.INIT('h1)
	) name396 (
		\y1_pad ,
		_w530_,
		_w532_
	);
	LUT2 #(
		.INIT('h4)
	) name397 (
		_w525_,
		_w532_,
		_w533_
	);
	LUT2 #(
		.INIT('h4)
	) name398 (
		_w531_,
		_w533_,
		_w534_
	);
	LUT2 #(
		.INIT('h4)
	) name399 (
		_w529_,
		_w534_,
		_w535_
	);
	LUT2 #(
		.INIT('h1)
	) name400 (
		\u0_pad ,
		_w465_,
		_w536_
	);
	LUT2 #(
		.INIT('h4)
	) name401 (
		m_pad,
		_w465_,
		_w537_
	);
	LUT2 #(
		.INIT('h1)
	) name402 (
		\y1_pad ,
		_w536_,
		_w538_
	);
	LUT2 #(
		.INIT('h4)
	) name403 (
		_w537_,
		_w538_,
		_w539_
	);
	LUT2 #(
		.INIT('h1)
	) name404 (
		\u1_pad ,
		_w422_,
		_w540_
	);
	LUT2 #(
		.INIT('h4)
	) name405 (
		y_pad,
		_w422_,
		_w541_
	);
	LUT2 #(
		.INIT('h1)
	) name406 (
		\y1_pad ,
		_w540_,
		_w542_
	);
	LUT2 #(
		.INIT('h4)
	) name407 (
		_w541_,
		_w542_,
		_w543_
	);
	LUT2 #(
		.INIT('h1)
	) name408 (
		\u2_pad ,
		_w497_,
		_w544_
	);
	LUT2 #(
		.INIT('h4)
	) name409 (
		\v2_pad ,
		_w497_,
		_w545_
	);
	LUT2 #(
		.INIT('h1)
	) name410 (
		\y1_pad ,
		_w544_,
		_w546_
	);
	LUT2 #(
		.INIT('h4)
	) name411 (
		_w545_,
		_w546_,
		_w547_
	);
	LUT2 #(
		.INIT('h4)
	) name412 (
		\d1_pad ,
		_w229_,
		_w548_
	);
	LUT2 #(
		.INIT('h8)
	) name413 (
		\v3_pad ,
		_w232_,
		_w549_
	);
	LUT2 #(
		.INIT('h2)
	) name414 (
		\u3_pad ,
		_w232_,
		_w550_
	);
	LUT2 #(
		.INIT('h2)
	) name415 (
		_w235_,
		_w549_,
		_w551_
	);
	LUT2 #(
		.INIT('h4)
	) name416 (
		_w550_,
		_w551_,
		_w552_
	);
	LUT2 #(
		.INIT('h2)
	) name417 (
		e_pad,
		\t1_pad ,
		_w553_
	);
	LUT2 #(
		.INIT('h4)
	) name418 (
		\e3_pad ,
		_w241_,
		_w554_
	);
	LUT2 #(
		.INIT('h1)
	) name419 (
		\y1_pad ,
		_w553_,
		_w555_
	);
	LUT2 #(
		.INIT('h4)
	) name420 (
		_w548_,
		_w555_,
		_w556_
	);
	LUT2 #(
		.INIT('h4)
	) name421 (
		_w554_,
		_w556_,
		_w557_
	);
	LUT2 #(
		.INIT('h4)
	) name422 (
		_w552_,
		_w557_,
		_w558_
	);
	LUT2 #(
		.INIT('h1)
	) name423 (
		\v0_pad ,
		_w465_,
		_w559_
	);
	LUT2 #(
		.INIT('h4)
	) name424 (
		n_pad,
		_w465_,
		_w560_
	);
	LUT2 #(
		.INIT('h1)
	) name425 (
		\y1_pad ,
		_w559_,
		_w561_
	);
	LUT2 #(
		.INIT('h4)
	) name426 (
		_w560_,
		_w561_,
		_w562_
	);
	LUT2 #(
		.INIT('h1)
	) name427 (
		\v1_pad ,
		_w422_,
		_w563_
	);
	LUT2 #(
		.INIT('h4)
	) name428 (
		z_pad,
		_w422_,
		_w564_
	);
	LUT2 #(
		.INIT('h1)
	) name429 (
		\y1_pad ,
		_w563_,
		_w565_
	);
	LUT2 #(
		.INIT('h4)
	) name430 (
		_w564_,
		_w565_,
		_w566_
	);
	LUT2 #(
		.INIT('h1)
	) name431 (
		\v2_pad ,
		_w497_,
		_w567_
	);
	LUT2 #(
		.INIT('h4)
	) name432 (
		\w2_pad ,
		_w497_,
		_w568_
	);
	LUT2 #(
		.INIT('h1)
	) name433 (
		\y1_pad ,
		_w567_,
		_w569_
	);
	LUT2 #(
		.INIT('h4)
	) name434 (
		_w568_,
		_w569_,
		_w570_
	);
	LUT2 #(
		.INIT('h4)
	) name435 (
		\e1_pad ,
		_w229_,
		_w571_
	);
	LUT2 #(
		.INIT('h8)
	) name436 (
		\w3_pad ,
		_w232_,
		_w572_
	);
	LUT2 #(
		.INIT('h2)
	) name437 (
		\v3_pad ,
		_w232_,
		_w573_
	);
	LUT2 #(
		.INIT('h2)
	) name438 (
		_w235_,
		_w572_,
		_w574_
	);
	LUT2 #(
		.INIT('h4)
	) name439 (
		_w573_,
		_w574_,
		_w575_
	);
	LUT2 #(
		.INIT('h2)
	) name440 (
		e_pad,
		\u1_pad ,
		_w576_
	);
	LUT2 #(
		.INIT('h4)
	) name441 (
		\f3_pad ,
		_w241_,
		_w577_
	);
	LUT2 #(
		.INIT('h1)
	) name442 (
		\y1_pad ,
		_w576_,
		_w578_
	);
	LUT2 #(
		.INIT('h4)
	) name443 (
		_w571_,
		_w578_,
		_w579_
	);
	LUT2 #(
		.INIT('h4)
	) name444 (
		_w577_,
		_w579_,
		_w580_
	);
	LUT2 #(
		.INIT('h4)
	) name445 (
		_w575_,
		_w580_,
		_w581_
	);
	LUT2 #(
		.INIT('h1)
	) name446 (
		\w0_pad ,
		_w465_,
		_w582_
	);
	LUT2 #(
		.INIT('h4)
	) name447 (
		o_pad,
		_w465_,
		_w583_
	);
	LUT2 #(
		.INIT('h1)
	) name448 (
		\y1_pad ,
		_w582_,
		_w584_
	);
	LUT2 #(
		.INIT('h4)
	) name449 (
		_w583_,
		_w584_,
		_w585_
	);
	LUT2 #(
		.INIT('h1)
	) name450 (
		\w1_pad ,
		_w422_,
		_w586_
	);
	LUT2 #(
		.INIT('h4)
	) name451 (
		\a0_pad ,
		_w422_,
		_w587_
	);
	LUT2 #(
		.INIT('h1)
	) name452 (
		\y1_pad ,
		_w586_,
		_w588_
	);
	LUT2 #(
		.INIT('h4)
	) name453 (
		_w587_,
		_w588_,
		_w589_
	);
	LUT2 #(
		.INIT('h1)
	) name454 (
		\w2_pad ,
		_w497_,
		_w590_
	);
	LUT2 #(
		.INIT('h4)
	) name455 (
		\x2_pad ,
		_w497_,
		_w591_
	);
	LUT2 #(
		.INIT('h1)
	) name456 (
		\y1_pad ,
		_w590_,
		_w592_
	);
	LUT2 #(
		.INIT('h4)
	) name457 (
		_w591_,
		_w592_,
		_w593_
	);
	LUT2 #(
		.INIT('h4)
	) name458 (
		\f1_pad ,
		_w229_,
		_w594_
	);
	LUT2 #(
		.INIT('h8)
	) name459 (
		\x3_pad ,
		_w232_,
		_w595_
	);
	LUT2 #(
		.INIT('h2)
	) name460 (
		\w3_pad ,
		_w232_,
		_w596_
	);
	LUT2 #(
		.INIT('h2)
	) name461 (
		_w235_,
		_w595_,
		_w597_
	);
	LUT2 #(
		.INIT('h4)
	) name462 (
		_w596_,
		_w597_,
		_w598_
	);
	LUT2 #(
		.INIT('h2)
	) name463 (
		e_pad,
		\v1_pad ,
		_w599_
	);
	LUT2 #(
		.INIT('h4)
	) name464 (
		\g3_pad ,
		_w241_,
		_w600_
	);
	LUT2 #(
		.INIT('h1)
	) name465 (
		\y1_pad ,
		_w599_,
		_w601_
	);
	LUT2 #(
		.INIT('h4)
	) name466 (
		_w594_,
		_w601_,
		_w602_
	);
	LUT2 #(
		.INIT('h4)
	) name467 (
		_w600_,
		_w602_,
		_w603_
	);
	LUT2 #(
		.INIT('h4)
	) name468 (
		_w598_,
		_w603_,
		_w604_
	);
	LUT2 #(
		.INIT('h1)
	) name469 (
		\x0_pad ,
		_w465_,
		_w605_
	);
	LUT2 #(
		.INIT('h4)
	) name470 (
		p_pad,
		_w465_,
		_w606_
	);
	LUT2 #(
		.INIT('h1)
	) name471 (
		\y1_pad ,
		_w605_,
		_w607_
	);
	LUT2 #(
		.INIT('h4)
	) name472 (
		_w606_,
		_w607_,
		_w608_
	);
	LUT2 #(
		.INIT('h1)
	) name473 (
		\y1_pad ,
		_w301_,
		_w609_
	);
	LUT2 #(
		.INIT('h1)
	) name474 (
		\x2_pad ,
		_w497_,
		_w610_
	);
	LUT2 #(
		.INIT('h4)
	) name475 (
		\y2_pad ,
		_w497_,
		_w611_
	);
	LUT2 #(
		.INIT('h1)
	) name476 (
		\y1_pad ,
		_w610_,
		_w612_
	);
	LUT2 #(
		.INIT('h4)
	) name477 (
		_w611_,
		_w612_,
		_w613_
	);
	LUT2 #(
		.INIT('h2)
	) name478 (
		e_pad,
		\w1_pad ,
		_w614_
	);
	LUT2 #(
		.INIT('h2)
	) name479 (
		\x3_pad ,
		_w232_,
		_w615_
	);
	LUT2 #(
		.INIT('h2)
	) name480 (
		_w235_,
		_w615_,
		_w616_
	);
	LUT2 #(
		.INIT('h4)
	) name481 (
		\h3_pad ,
		_w241_,
		_w617_
	);
	LUT2 #(
		.INIT('h4)
	) name482 (
		\g1_pad ,
		_w229_,
		_w618_
	);
	LUT2 #(
		.INIT('h1)
	) name483 (
		\y1_pad ,
		_w614_,
		_w619_
	);
	LUT2 #(
		.INIT('h4)
	) name484 (
		_w618_,
		_w619_,
		_w620_
	);
	LUT2 #(
		.INIT('h4)
	) name485 (
		_w617_,
		_w620_,
		_w621_
	);
	LUT2 #(
		.INIT('h4)
	) name486 (
		_w616_,
		_w621_,
		_w622_
	);
	LUT2 #(
		.INIT('h1)
	) name487 (
		\y0_pad ,
		_w465_,
		_w623_
	);
	LUT2 #(
		.INIT('h4)
	) name488 (
		q_pad,
		_w465_,
		_w624_
	);
	LUT2 #(
		.INIT('h1)
	) name489 (
		\y1_pad ,
		_w623_,
		_w625_
	);
	LUT2 #(
		.INIT('h4)
	) name490 (
		_w624_,
		_w625_,
		_w626_
	);
	LUT2 #(
		.INIT('h1)
	) name491 (
		\n0_pad ,
		_w358_,
		_w627_
	);
	LUT2 #(
		.INIT('h1)
	) name492 (
		\y2_pad ,
		_w497_,
		_w628_
	);
	LUT2 #(
		.INIT('h4)
	) name493 (
		\z2_pad ,
		_w497_,
		_w629_
	);
	LUT2 #(
		.INIT('h1)
	) name494 (
		\y1_pad ,
		_w628_,
		_w630_
	);
	LUT2 #(
		.INIT('h4)
	) name495 (
		_w629_,
		_w630_,
		_w631_
	);
	LUT2 #(
		.INIT('h4)
	) name496 (
		\y3_pad ,
		_w179_,
		_w632_
	);
	LUT2 #(
		.INIT('h1)
	) name497 (
		\z0_pad ,
		_w136_,
		_w633_
	);
	LUT2 #(
		.INIT('h4)
	) name498 (
		j_pad,
		_w136_,
		_w634_
	);
	LUT2 #(
		.INIT('h1)
	) name499 (
		\y1_pad ,
		_w633_,
		_w635_
	);
	LUT2 #(
		.INIT('h4)
	) name500 (
		_w634_,
		_w635_,
		_w636_
	);
	LUT2 #(
		.INIT('h2)
	) name501 (
		_w383_,
		_w408_,
		_w637_
	);
	LUT2 #(
		.INIT('h4)
	) name502 (
		\d0_pad ,
		\r2_pad ,
		_w638_
	);
	LUT2 #(
		.INIT('h8)
	) name503 (
		\c0_pad ,
		\q2_pad ,
		_w639_
	);
	LUT2 #(
		.INIT('h1)
	) name504 (
		_w638_,
		_w639_,
		_w640_
	);
	LUT2 #(
		.INIT('h2)
	) name505 (
		\i2_pad ,
		_w640_,
		_w641_
	);
	LUT2 #(
		.INIT('h1)
	) name506 (
		_w231_,
		_w382_,
		_w642_
	);
	LUT2 #(
		.INIT('h4)
	) name507 (
		\i3_pad ,
		_w642_,
		_w643_
	);
	LUT2 #(
		.INIT('h1)
	) name508 (
		\x1_pad ,
		_w641_,
		_w644_
	);
	LUT2 #(
		.INIT('h4)
	) name509 (
		_w643_,
		_w644_,
		_w645_
	);
	LUT2 #(
		.INIT('h4)
	) name510 (
		_w637_,
		_w645_,
		_w646_
	);
	LUT2 #(
		.INIT('h2)
	) name511 (
		\z1_pad ,
		_w646_,
		_w647_
	);
	LUT2 #(
		.INIT('h1)
	) name512 (
		_w358_,
		_w647_,
		_w648_
	);
	LUT2 #(
		.INIT('h1)
	) name513 (
		\y1_pad ,
		_w648_,
		_w649_
	);
	LUT2 #(
		.INIT('h8)
	) name514 (
		\i3_pad ,
		_w642_,
		_w650_
	);
	LUT2 #(
		.INIT('h8)
	) name515 (
		_w383_,
		_w408_,
		_w651_
	);
	LUT2 #(
		.INIT('h2)
	) name516 (
		\c0_pad ,
		_w385_,
		_w652_
	);
	LUT2 #(
		.INIT('h2)
	) name517 (
		_w387_,
		_w652_,
		_w653_
	);
	LUT2 #(
		.INIT('h1)
	) name518 (
		_w650_,
		_w653_,
		_w654_
	);
	LUT2 #(
		.INIT('h4)
	) name519 (
		_w651_,
		_w654_,
		_w655_
	);
	LUT2 #(
		.INIT('h1)
	) name520 (
		\x1_pad ,
		\y1_pad ,
		_w656_
	);
	LUT2 #(
		.INIT('h4)
	) name521 (
		\z1_pad ,
		_w656_,
		_w657_
	);
	LUT2 #(
		.INIT('h4)
	) name522 (
		_w655_,
		_w657_,
		_w658_
	);
	LUT2 #(
		.INIT('h1)
	) name523 (
		_w649_,
		_w658_,
		_w659_
	);
	LUT2 #(
		.INIT('h1)
	) name524 (
		\z2_pad ,
		_w497_,
		_w660_
	);
	LUT2 #(
		.INIT('h4)
	) name525 (
		g_pad,
		_w497_,
		_w661_
	);
	LUT2 #(
		.INIT('h1)
	) name526 (
		\y1_pad ,
		_w660_,
		_w662_
	);
	LUT2 #(
		.INIT('h4)
	) name527 (
		_w661_,
		_w662_,
		_w663_
	);
	LUT2 #(
		.INIT('h8)
	) name528 (
		\y3_pad ,
		\z3_pad ,
		_w664_
	);
	LUT2 #(
		.INIT('h1)
	) name529 (
		\y3_pad ,
		\z3_pad ,
		_w665_
	);
	LUT2 #(
		.INIT('h2)
	) name530 (
		_w179_,
		_w664_,
		_w666_
	);
	LUT2 #(
		.INIT('h4)
	) name531 (
		_w665_,
		_w666_,
		_w667_
	);
	LUT2 #(
		.INIT('h1)
	) name532 (
		\a1_pad ,
		_w136_,
		_w668_
	);
	LUT2 #(
		.INIT('h4)
	) name533 (
		k_pad,
		_w136_,
		_w669_
	);
	LUT2 #(
		.INIT('h1)
	) name534 (
		\y1_pad ,
		_w668_,
		_w670_
	);
	LUT2 #(
		.INIT('h4)
	) name535 (
		_w669_,
		_w670_,
		_w671_
	);
	LUT2 #(
		.INIT('h2)
	) name536 (
		_w167_,
		_w415_,
		_w672_
	);
	LUT2 #(
		.INIT('h1)
	) name537 (
		\y1_pad ,
		_w672_,
		_w673_
	);
	LUT2 #(
		.INIT('h1)
	) name538 (
		\a3_pad ,
		_w174_,
		_w674_
	);
	LUT2 #(
		.INIT('h4)
	) name539 (
		\b3_pad ,
		_w174_,
		_w675_
	);
	LUT2 #(
		.INIT('h1)
	) name540 (
		\y1_pad ,
		_w674_,
		_w676_
	);
	LUT2 #(
		.INIT('h4)
	) name541 (
		_w675_,
		_w676_,
		_w677_
	);
	LUT2 #(
		.INIT('h1)
	) name542 (
		\a4_pad ,
		_w664_,
		_w678_
	);
	LUT2 #(
		.INIT('h4)
	) name543 (
		_w142_,
		_w179_,
		_w679_
	);
	LUT2 #(
		.INIT('h4)
	) name544 (
		_w678_,
		_w679_,
		_w680_
	);
	LUT2 #(
		.INIT('h1)
	) name545 (
		\b1_pad ,
		_w136_,
		_w681_
	);
	LUT2 #(
		.INIT('h4)
	) name546 (
		l_pad,
		_w136_,
		_w682_
	);
	LUT2 #(
		.INIT('h1)
	) name547 (
		\y1_pad ,
		_w681_,
		_w683_
	);
	LUT2 #(
		.INIT('h4)
	) name548 (
		_w682_,
		_w683_,
		_w684_
	);
	LUT2 #(
		.INIT('h8)
	) name549 (
		\d4_pad ,
		_w144_,
		_w685_
	);
	LUT2 #(
		.INIT('h1)
	) name550 (
		\e4_pad ,
		\f4_pad ,
		_w686_
	);
	LUT2 #(
		.INIT('h4)
	) name551 (
		\g4_pad ,
		_w686_,
		_w687_
	);
	LUT2 #(
		.INIT('h8)
	) name552 (
		_w685_,
		_w687_,
		_w688_
	);
	LUT2 #(
		.INIT('h8)
	) name553 (
		\b2_pad ,
		_w688_,
		_w689_
	);
	LUT2 #(
		.INIT('h1)
	) name554 (
		\b2_pad ,
		_w688_,
		_w690_
	);
	LUT2 #(
		.INIT('h2)
	) name555 (
		_w179_,
		_w689_,
		_w691_
	);
	LUT2 #(
		.INIT('h4)
	) name556 (
		_w690_,
		_w691_,
		_w692_
	);
	LUT2 #(
		.INIT('h1)
	) name557 (
		\b3_pad ,
		_w174_,
		_w693_
	);
	LUT2 #(
		.INIT('h4)
	) name558 (
		\c3_pad ,
		_w174_,
		_w694_
	);
	LUT2 #(
		.INIT('h1)
	) name559 (
		\y1_pad ,
		_w693_,
		_w695_
	);
	LUT2 #(
		.INIT('h4)
	) name560 (
		_w694_,
		_w695_,
		_w696_
	);
	LUT2 #(
		.INIT('h1)
	) name561 (
		\b4_pad ,
		_w142_,
		_w697_
	);
	LUT2 #(
		.INIT('h4)
	) name562 (
		_w143_,
		_w179_,
		_w698_
	);
	LUT2 #(
		.INIT('h4)
	) name563 (
		_w697_,
		_w698_,
		_w699_
	);
	LUT2 #(
		.INIT('h1)
	) name564 (
		\c1_pad ,
		_w136_,
		_w700_
	);
	LUT2 #(
		.INIT('h4)
	) name565 (
		m_pad,
		_w136_,
		_w701_
	);
	LUT2 #(
		.INIT('h1)
	) name566 (
		\y1_pad ,
		_w700_,
		_w702_
	);
	LUT2 #(
		.INIT('h4)
	) name567 (
		_w701_,
		_w702_,
		_w703_
	);
	LUT2 #(
		.INIT('h1)
	) name568 (
		\c2_pad ,
		_w689_,
		_w704_
	);
	LUT2 #(
		.INIT('h8)
	) name569 (
		\c2_pad ,
		_w689_,
		_w705_
	);
	LUT2 #(
		.INIT('h2)
	) name570 (
		_w179_,
		_w704_,
		_w706_
	);
	LUT2 #(
		.INIT('h4)
	) name571 (
		_w705_,
		_w706_,
		_w707_
	);
	LUT2 #(
		.INIT('h1)
	) name572 (
		\c3_pad ,
		_w174_,
		_w708_
	);
	LUT2 #(
		.INIT('h4)
	) name573 (
		\d3_pad ,
		_w174_,
		_w709_
	);
	LUT2 #(
		.INIT('h1)
	) name574 (
		\y1_pad ,
		_w708_,
		_w710_
	);
	LUT2 #(
		.INIT('h4)
	) name575 (
		_w709_,
		_w710_,
		_w711_
	);
	LUT2 #(
		.INIT('h1)
	) name576 (
		\c4_pad ,
		_w143_,
		_w712_
	);
	LUT2 #(
		.INIT('h4)
	) name577 (
		_w144_,
		_w179_,
		_w713_
	);
	LUT2 #(
		.INIT('h4)
	) name578 (
		_w712_,
		_w713_,
		_w714_
	);
	LUT2 #(
		.INIT('h1)
	) name579 (
		\d1_pad ,
		_w136_,
		_w715_
	);
	LUT2 #(
		.INIT('h4)
	) name580 (
		n_pad,
		_w136_,
		_w716_
	);
	LUT2 #(
		.INIT('h1)
	) name581 (
		\y1_pad ,
		_w715_,
		_w717_
	);
	LUT2 #(
		.INIT('h4)
	) name582 (
		_w716_,
		_w717_,
		_w718_
	);
	LUT2 #(
		.INIT('h1)
	) name583 (
		\d2_pad ,
		\l0_pad ,
		_w719_
	);
	LUT2 #(
		.INIT('h2)
	) name584 (
		_w212_,
		_w719_,
		_w720_
	);
	LUT2 #(
		.INIT('h1)
	) name585 (
		\d3_pad ,
		_w174_,
		_w721_
	);
	LUT2 #(
		.INIT('h4)
	) name586 (
		\e3_pad ,
		_w174_,
		_w722_
	);
	LUT2 #(
		.INIT('h1)
	) name587 (
		\y1_pad ,
		_w721_,
		_w723_
	);
	LUT2 #(
		.INIT('h4)
	) name588 (
		_w722_,
		_w723_,
		_w724_
	);
	LUT2 #(
		.INIT('h1)
	) name589 (
		\d4_pad ,
		_w144_,
		_w725_
	);
	LUT2 #(
		.INIT('h2)
	) name590 (
		_w179_,
		_w685_,
		_w726_
	);
	LUT2 #(
		.INIT('h4)
	) name591 (
		_w725_,
		_w726_,
		_w727_
	);
	LUT2 #(
		.INIT('h1)
	) name592 (
		\e1_pad ,
		_w136_,
		_w728_
	);
	LUT2 #(
		.INIT('h4)
	) name593 (
		o_pad,
		_w136_,
		_w729_
	);
	LUT2 #(
		.INIT('h1)
	) name594 (
		\y1_pad ,
		_w728_,
		_w730_
	);
	LUT2 #(
		.INIT('h4)
	) name595 (
		_w729_,
		_w730_,
		_w731_
	);
	LUT2 #(
		.INIT('h4)
	) name596 (
		\e2_pad ,
		_w168_,
		_w732_
	);
	LUT2 #(
		.INIT('h1)
	) name597 (
		\n0_pad ,
		_w169_,
		_w733_
	);
	LUT2 #(
		.INIT('h4)
	) name598 (
		_w732_,
		_w733_,
		_w734_
	);
	LUT2 #(
		.INIT('h1)
	) name599 (
		\e3_pad ,
		_w174_,
		_w735_
	);
	LUT2 #(
		.INIT('h4)
	) name600 (
		\f3_pad ,
		_w174_,
		_w736_
	);
	LUT2 #(
		.INIT('h1)
	) name601 (
		\y1_pad ,
		_w735_,
		_w737_
	);
	LUT2 #(
		.INIT('h4)
	) name602 (
		_w736_,
		_w737_,
		_w738_
	);
	LUT2 #(
		.INIT('h1)
	) name603 (
		\e4_pad ,
		_w180_,
		_w739_
	);
	LUT2 #(
		.INIT('h2)
	) name604 (
		_w179_,
		_w181_,
		_w740_
	);
	LUT2 #(
		.INIT('h4)
	) name605 (
		_w739_,
		_w740_,
		_w741_
	);
	assign \a5_pad  = _w140_ ;
	assign \a6_pad  = _w173_ ;
	assign \a7_pad  = _w178_ ;
	assign \a8_pad  = _w185_ ;
	assign \b5_pad  = _w189_ ;
	assign \b6_pad  = _w190_ ;
	assign \b7_pad  = _w194_ ;
	assign \b8_pad  = _w198_ ;
	assign \c5_pad  = _w203_ ;
	assign \c6_pad  = _w204_ ;
	assign \c7_pad  = _w208_ ;
	assign \c8_pad  = _w213_ ;
	assign \d5_pad  = _w217_ ;
	assign \d6_pad  = _w228_ ;
	assign \d7_pad  = _w246_ ;
	assign \e5_pad  = _w250_ ;
	assign \e6_pad  = _w261_ ;
	assign \e7_pad  = _w272_ ;
	assign \f5_pad  = _w276_ ;
	assign \f6_pad  = _w285_ ;
	assign \f7_pad  = _w296_ ;
	assign \g5_pad  = _w300_ ;
	assign \g6_pad  = _w305_ ;
	assign \g7_pad  = _w316_ ;
	assign \h5_pad  = _w320_ ;
	assign \h6_pad  = _w324_ ;
	assign \h7_pad  = _w335_ ;
	assign \i4_pad  = _w336_ ;
	assign \i5_pad  = _w340_ ;
	assign \i6_pad  = _w344_ ;
	assign \i7_pad  = _w355_ ;
	assign \j4_pad  = _w361_ ;
	assign \j5_pad  = _w365_ ;
	assign \j6_pad  = _w369_ ;
	assign \j7_pad  = _w380_ ;
	assign \k4_pad  = _w421_ ;
	assign \k5_pad  = _w426_ ;
	assign \k6_pad  = _w430_ ;
	assign \k7_pad  = _w441_ ;
	assign \l4_pad  = _w443_ ;
	assign \l5_pad  = _w447_ ;
	assign \l6_pad  = _w453_ ;
	assign \l7_pad  = _w464_ ;
	assign \m4_pad  = _w469_ ;
	assign \m5_pad  = _w473_ ;
	assign \m6_pad  = _w477_ ;
	assign \m7_pad  = _w488_ ;
	assign \n4_pad  = _w492_ ;
	assign \n5_pad  = _w496_ ;
	assign \n6_pad  = _w501_ ;
	assign \n7_pad  = _w512_ ;
	assign \o4_pad  = _w516_ ;
	assign \o5_pad  = _w520_ ;
	assign \o6_pad  = _w524_ ;
	assign \o7_pad  = _w535_ ;
	assign \p4_pad  = _w539_ ;
	assign \p5_pad  = _w543_ ;
	assign \p6_pad  = _w547_ ;
	assign \p7_pad  = _w558_ ;
	assign \q4_pad  = _w562_ ;
	assign \q5_pad  = _w566_ ;
	assign \q6_pad  = _w570_ ;
	assign \q7_pad  = _w581_ ;
	assign \r4_pad  = _w585_ ;
	assign \r5_pad  = _w589_ ;
	assign \r6_pad  = _w593_ ;
	assign \r7_pad  = _w604_ ;
	assign \s4_pad  = _w608_ ;
	assign \s5_pad  = _w609_ ;
	assign \s6_pad  = _w613_ ;
	assign \s7_pad  = _w622_ ;
	assign \t4_pad  = _w626_ ;
	assign \t5_pad  = _w627_ ;
	assign \t6_pad  = _w631_ ;
	assign \t7_pad  = _w632_ ;
	assign \u4_pad  = _w636_ ;
	assign \u5_pad  = _w659_ ;
	assign \u6_pad  = _w663_ ;
	assign \u7_pad  = _w667_ ;
	assign \v4_pad  = _w671_ ;
	assign \v5_pad  = _w673_ ;
	assign \v6_pad  = _w677_ ;
	assign \v7_pad  = _w680_ ;
	assign \w4_pad  = _w684_ ;
	assign \w5_pad  = _w692_ ;
	assign \w6_pad  = _w696_ ;
	assign \w7_pad  = _w699_ ;
	assign \x4_pad  = _w703_ ;
	assign \x5_pad  = _w707_ ;
	assign \x6_pad  = _w711_ ;
	assign \x7_pad  = _w714_ ;
	assign \y4_pad  = _w718_ ;
	assign \y5_pad  = _w720_ ;
	assign \y6_pad  = _w724_ ;
	assign \y7_pad  = _w727_ ;
	assign \z4_pad  = _w731_ ;
	assign \z5_pad  = _w734_ ;
	assign \z6_pad  = _w738_ ;
	assign \z7_pad  = _w741_ ;
endmodule;