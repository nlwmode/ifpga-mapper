module top (\n1035gat_reg/NET0131 , \n1045gat_reg/NET0131 , \n1068gat_reg/NET0131 , \n1072gat_reg/NET0131 , \n1080gat_reg/NET0131 , \n1121gat_reg/NET0131 , \n1135gat_reg/NET0131 , \n1148gat_reg/NET0131 , \n1197gat_reg/NET0131 , \n1226gat_reg/NET0131 , \n1241gat_reg/NET0131 , \n1282gat_reg/NET0131 , \n1294gat_reg/NET0131 , \n1312gat_reg/NET0131 , \n1316gat_reg/NET0131 , \n1332gat_reg/NET0131 , \n1336gat_reg/NET0131 , \n1340gat_reg/NET0131 , \n1363gat_reg/NET0131 , \n1389gat_reg/NET0131 , \n1394gat_reg/NET0131 , \n1433gat_reg/NET0131 , \n1456gat_reg/NET0131 , \n1462gat_reg/NET0131 , \n148gat_reg/NET0131 , \n1496gat_reg/NET0131 , \n1508gat_reg/NET0131 , \n1525gat_reg/NET0131 , \n152gat_reg/NET0131 , \n156gat_reg/NET0131 , \n1588gat_reg/NET0131 , \n1596gat_reg/NET0131 , \n160gat_reg/NET0131 , \n1675gat_reg/NET0131 , \n1678gat_reg/NET0131 , \n1740gat_reg/NET0131 , \n1748gat_reg/NET0131 , \n1763gat_reg/NET0131 , \n1767gat_reg/NET0131 , \n1771gat_reg/NET0131 , \n1775gat_reg/NET0131 , \n1807gat_reg/NET0131 , \n1821gat_reg/NET0131 , \n1829gat_reg/NET0131 , \n1834gat_reg/NET0131 , \n1850gat_reg/NET0131 , \n1871gat_reg/NET0131 , \n1880gat_reg/NET0131 , \n1899gat_reg/NET0131 , \n1975gat_reg/NET0131 , \n2021gat_reg/NET0131 , \n2025gat_reg/NET0131 , \n2029gat_reg/NET0131 , \n2033gat_reg/NET0131 , \n2037gat_reg/NET0131 , \n2040gat_reg/NET0131 , \n2044gat_reg/NET0131 , \n2061gat_reg/NET0131 , \n2084gat_reg/NET0131 , \n2091gat_reg/NET0131 , \n2095gat_reg/NET0131 , \n2099gat_reg/NET0131 , \n2102gat_reg/NET0131 , \n2110gat_reg/NET0131 , \n2117gat_reg/NET0131 , \n2121gat_reg/NET0131 , \n2125gat_reg/NET0131 , \n2135gat_reg/NET0131 , \n2139gat_reg/NET0131 , \n2143gat_reg/NET0131 , \n2155gat_reg/NET0131 , \n2169gat_reg/NET0131 , \n2176gat_reg/NET0131 , \n2179gat_reg/NET0131 , \n2182gat_reg/NET0131 , \n2190gat_reg/NET0131 , \n2203gat_reg/NET0131 , \n2207gat_reg/NET0131 , \n2262gat_reg/NET0131 , \n2266gat_reg/NET0131 , \n2270gat_reg/NET0131 , \n2319gat_reg/NET0131 , \n2339gat_reg/NET0131 , \n2343gat_reg/NET0131 , \n2347gat_reg/NET0131 , \n2390gat_reg/NET0131 , \n2394gat_reg/NET0131 , \n2399gat_reg/NET0131 , \n2403gat_reg/NET0131 , \n2407gat_reg/NET0131 , \n2440gat_reg/NET0131 , \n2446gat_reg/NET0131 , \n2450gat_reg/NET0131 , \n2454gat_reg/NET0131 , \n2458gat_reg/NET0131 , \n2464gat_reg/NET0131 , \n2468gat_reg/NET0131 , \n2472gat_reg/NET0131 , \n2476gat_reg/NET0131 , \n2490gat_reg/NET0131 , \n2495gat_reg/NET0131 , \n2502gat_reg/NET0131 , \n2506gat_reg/NET0131 , \n2510gat_reg/NET0131 , \n2514gat_reg/NET0131 , \n2518gat_reg/NET0131 , \n2526gat_reg/NET0131 , \n2543gat_reg/NET0131 , \n2562gat_reg/NET0131 , \n256gat_reg/NET0131 , \n2588gat_reg/NET0131 , \n2592gat_reg/NET0131 , \n2599gat_reg/NET0131 , \n2622gat_reg/NET0131 , \n2626gat_reg/NET0131 , \n2630gat_reg/NET0131 , \n2634gat_reg/NET0131 , \n2640gat_reg/NET0131 , \n2644gat_reg/NET0131 , \n2658gat_reg/NET0131 , \n271gat_reg/NET0131 , \n3065gat_pad , \n3066gat_pad , \n3067gat_pad , \n3068gat_pad , \n3069gat_pad , \n3070gat_pad , \n3071gat_pad , \n3072gat_pad , \n3073gat_pad , \n3074gat_pad , \n3075gat_pad , \n3076gat_pad , \n3077gat_pad , \n3078gat_pad , \n3079gat_pad , \n3080gat_pad , \n3081gat_pad , \n3082gat_pad , \n3083gat_pad , \n3084gat_pad , \n3085gat_pad , \n3086gat_pad , \n3087gat_pad , \n3088gat_pad , \n3089gat_pad , \n3090gat_pad , \n3091gat_pad , \n3092gat_pad , \n3093gat_pad , \n3094gat_pad , \n3095gat_pad , \n3097gat_pad , \n3098gat_pad , \n3099gat_pad , \n3100gat_pad , \n314gat_reg/NET0131 , \n318gat_reg/NET0131 , \n322gat_reg/NET0131 , \n327gat_reg/NET0131 , \n331gat_reg/NET0131 , \n337gat_reg/NET0131 , \n341gat_reg/NET0131 , \n366gat_reg/NET0131 , \n384gat_reg/NET0131 , \n388gat_reg/NET0131 , \n398gat_reg/NET0131 , \n402gat_reg/NET0131 , \n463gat_reg/NET0131 , \n470gat_reg/NET0131 , \n553gat_reg/NET0131 , \n561gat_reg/NET0131 , \n580gat_reg/NET0131 , \n584gat_reg/NET0131 , \n614gat_reg/NET0131 , \n659gat_reg/NET0131 , \n667gat_reg/NET0131 , \n673gat_reg/NET0131 , \n680gat_reg/NET0131 , \n684gat_reg/NET0131 , \n699gat_reg/NET0131 , \n707gat_reg/NET0131 , \n777gat_reg/NET0131 , \n816gat_reg/NET0131 , \n820gat_reg/NET0131 , \n824gat_reg/NET0131 , \n830gat_reg/NET0131 , \n834gat_reg/NET0131 , \n838gat_reg/NET0131 , \n842gat_reg/NET0131 , \n846gat_reg/NET0131 , \n861gat_reg/NET0131 , \n865gat_reg/NET0131 , \n883gat_reg/NET0131 , \n919gat_reg/NET0131 , \n931gat_reg/NET0131 , \n957gat_reg/NET0131 , \_al_n0 , \g17_dup/_0_ , \g6952/_2_ , \g6953/_2_ , \g6961/_0_ , \g7076/_0_ , \g7077/_0_ , \g7079/_0_ , \g7081/_0_ , \g7082/_0_ , \g7083/_0_ , \g7146/_0_ , \g7147/_0_ , \g7148/_0_ , \g7149/_0_ , \g7150/_0_ , \g7151/_0_ , \g7152/_0_ , \g7153/_0_ , \g7154/_0_ , \g7156/_2_ , \g7161/_2_ , \g7165/_2_ , \g7174/_0_ , \g7180/_00_ , \g7182/_3_ , \g7191/_0_ , \g7204/_0_ , \g7209/_3_ , \g7220/_0_ , \g7229/_0_ , \g7233/_0_ , \g7234/_0_ , \g7235/_0_ , \g7236/_0_ , \g7237/_0_ , \g7238/_0_ , \g7241/_3_ , \g7264/_0_ , \g7265/_0_ , \g7266/_0_ , \g7267/_0_ , \g7268/_0_ , \g7301/_0_ , \g7326/_3_ , \g7350/_2_ , \g7352/_0_ , \g7356/_0_ , \g7359/_0_ , \g7389/_3_ , \g7417/_0_ , \g7418/_0_ , \g7419/_0_ , \g7444/_0_ , \g7445/_0_ , \g7449/_3_ , \g7451/_3_ , \g7454/_0_ , \g7467/_3_ , \g7476/_0_ , \g7480/_0_ , \g7494/_0_ , \g7509/_0_ , \g7514/_0_ , \g7517/_3_ , \g7524/_0_ , \g7558/_0_ , \g7560/_0_ , \g7561/_0_ , \g7563/_0_ , \g7567/_0_ , \g7572/_0_ , \g7579/_0_ , \g7605/_0_ , \g7625/_0_ , \g7627/_0_ , \g7671/_0_ , \g7675/_0_ , \g7689/_0_ , \g7697/_0_ , \g7743/_1_ , \g7764/_1_ , \g7769/_0_ , \g7771/_2_ , \g7779/_0_ , \g7852/_0_ , \g7873/_0_ , \g7884/_3_ , \g7889/_0_ , \g7902/_1_ , \g7992/_3_ , \g7994/_3_ , \g7996/_3_ , \g7998/_3_ , \g8000/_3_ , \g8002/_3_ , \g8004/_3_ , \g8006/_3_ , \g8008/_3_ , \g8150/_0_ , \g8151/_0_ , \g8157/_0_ , \g8163/_0_ , \g8172/_0_ , \g8197/_0_ , \g8211/_0_ , \g8223/_0_ , \g8237/_0_ , \g8251/_0_ , \g8261/_0_ , \g8272/_0_ , \g8287/_0_ , \g8647/_0_ , \g8671/_0_ , \g8672/_0_ , \g8735/_0_ , \g8766/_0_ , \g8811/_0_ , \g8821/_0_ , \g8856/_0_ , \g8858/_3_ , \g8868/_0_ , \g8880/_2_ , \g8886/_0_ , \g8900/_0_ , \g8932/_0_ , \g8991/_3_ , \g9014/_3_ , \g9074/_0_ , \g9091/_0_ , \g9105/_0_ , \g9107/_1_ , \g9111/_0_ , \n1332gat_reg/P0001 , \n1363gat_reg/P0001 , \n1394gat_reg/P0001 , \n1433gat_reg/P0001 , \n1775gat_reg/P0001 , \n2025gat_reg/P0001 , \n2029gat_reg/P0001 , \n2033gat_reg/P0001 , \n2044gat_reg/P0001 , \n2121gat_reg/P0001 , \n2125gat_reg/P0001 , \n2458gat_reg/P0001 , \n2472gat_reg/P0001 , \n2592gat_reg/P0001 , \n3104gat_pad , \n3105gat_pad , \n3106gat_pad , \n3107gat_pad , \n3108gat_pad , \n3109gat_pad , \n3110gat_pad , \n3111gat_pad , \n3112gat_pad , \n3113gat_pad , \n3114gat_pad , \n3116gat_pad , \n3117gat_pad , \n3118gat_pad , \n3119gat_pad , \n3120gat_pad , \n3121gat_pad , \n3122gat_pad , \n3123gat_pad , \n3124gat_pad , \n3125gat_pad , \n3126gat_pad , \n3127gat_pad , \n3128gat_pad , \n3130gat_pad , \n3131gat_pad , \n3132gat_pad , \n3133gat_pad , \n3134gat_pad , \n3135gat_pad , \n3136gat_pad , \n3137gat_pad , \n3138gat_pad , \n3140gat_pad , \n3142gat_pad , \n3143gat_pad , \n3144gat_pad , \n3145gat_pad , \n3146gat_pad , \n3147gat_pad , \n3148gat_pad , \n3149gat_pad , \n3150gat_pad , \n3151gat_pad , \n684gat_reg/P0001 , \n824gat_reg/P0001 , \n883gat_reg/P0001 );
	input \n1035gat_reg/NET0131  ;
	input \n1045gat_reg/NET0131  ;
	input \n1068gat_reg/NET0131  ;
	input \n1072gat_reg/NET0131  ;
	input \n1080gat_reg/NET0131  ;
	input \n1121gat_reg/NET0131  ;
	input \n1135gat_reg/NET0131  ;
	input \n1148gat_reg/NET0131  ;
	input \n1197gat_reg/NET0131  ;
	input \n1226gat_reg/NET0131  ;
	input \n1241gat_reg/NET0131  ;
	input \n1282gat_reg/NET0131  ;
	input \n1294gat_reg/NET0131  ;
	input \n1312gat_reg/NET0131  ;
	input \n1316gat_reg/NET0131  ;
	input \n1332gat_reg/NET0131  ;
	input \n1336gat_reg/NET0131  ;
	input \n1340gat_reg/NET0131  ;
	input \n1363gat_reg/NET0131  ;
	input \n1389gat_reg/NET0131  ;
	input \n1394gat_reg/NET0131  ;
	input \n1433gat_reg/NET0131  ;
	input \n1456gat_reg/NET0131  ;
	input \n1462gat_reg/NET0131  ;
	input \n148gat_reg/NET0131  ;
	input \n1496gat_reg/NET0131  ;
	input \n1508gat_reg/NET0131  ;
	input \n1525gat_reg/NET0131  ;
	input \n152gat_reg/NET0131  ;
	input \n156gat_reg/NET0131  ;
	input \n1588gat_reg/NET0131  ;
	input \n1596gat_reg/NET0131  ;
	input \n160gat_reg/NET0131  ;
	input \n1675gat_reg/NET0131  ;
	input \n1678gat_reg/NET0131  ;
	input \n1740gat_reg/NET0131  ;
	input \n1748gat_reg/NET0131  ;
	input \n1763gat_reg/NET0131  ;
	input \n1767gat_reg/NET0131  ;
	input \n1771gat_reg/NET0131  ;
	input \n1775gat_reg/NET0131  ;
	input \n1807gat_reg/NET0131  ;
	input \n1821gat_reg/NET0131  ;
	input \n1829gat_reg/NET0131  ;
	input \n1834gat_reg/NET0131  ;
	input \n1850gat_reg/NET0131  ;
	input \n1871gat_reg/NET0131  ;
	input \n1880gat_reg/NET0131  ;
	input \n1899gat_reg/NET0131  ;
	input \n1975gat_reg/NET0131  ;
	input \n2021gat_reg/NET0131  ;
	input \n2025gat_reg/NET0131  ;
	input \n2029gat_reg/NET0131  ;
	input \n2033gat_reg/NET0131  ;
	input \n2037gat_reg/NET0131  ;
	input \n2040gat_reg/NET0131  ;
	input \n2044gat_reg/NET0131  ;
	input \n2061gat_reg/NET0131  ;
	input \n2084gat_reg/NET0131  ;
	input \n2091gat_reg/NET0131  ;
	input \n2095gat_reg/NET0131  ;
	input \n2099gat_reg/NET0131  ;
	input \n2102gat_reg/NET0131  ;
	input \n2110gat_reg/NET0131  ;
	input \n2117gat_reg/NET0131  ;
	input \n2121gat_reg/NET0131  ;
	input \n2125gat_reg/NET0131  ;
	input \n2135gat_reg/NET0131  ;
	input \n2139gat_reg/NET0131  ;
	input \n2143gat_reg/NET0131  ;
	input \n2155gat_reg/NET0131  ;
	input \n2169gat_reg/NET0131  ;
	input \n2176gat_reg/NET0131  ;
	input \n2179gat_reg/NET0131  ;
	input \n2182gat_reg/NET0131  ;
	input \n2190gat_reg/NET0131  ;
	input \n2203gat_reg/NET0131  ;
	input \n2207gat_reg/NET0131  ;
	input \n2262gat_reg/NET0131  ;
	input \n2266gat_reg/NET0131  ;
	input \n2270gat_reg/NET0131  ;
	input \n2319gat_reg/NET0131  ;
	input \n2339gat_reg/NET0131  ;
	input \n2343gat_reg/NET0131  ;
	input \n2347gat_reg/NET0131  ;
	input \n2390gat_reg/NET0131  ;
	input \n2394gat_reg/NET0131  ;
	input \n2399gat_reg/NET0131  ;
	input \n2403gat_reg/NET0131  ;
	input \n2407gat_reg/NET0131  ;
	input \n2440gat_reg/NET0131  ;
	input \n2446gat_reg/NET0131  ;
	input \n2450gat_reg/NET0131  ;
	input \n2454gat_reg/NET0131  ;
	input \n2458gat_reg/NET0131  ;
	input \n2464gat_reg/NET0131  ;
	input \n2468gat_reg/NET0131  ;
	input \n2472gat_reg/NET0131  ;
	input \n2476gat_reg/NET0131  ;
	input \n2490gat_reg/NET0131  ;
	input \n2495gat_reg/NET0131  ;
	input \n2502gat_reg/NET0131  ;
	input \n2506gat_reg/NET0131  ;
	input \n2510gat_reg/NET0131  ;
	input \n2514gat_reg/NET0131  ;
	input \n2518gat_reg/NET0131  ;
	input \n2526gat_reg/NET0131  ;
	input \n2543gat_reg/NET0131  ;
	input \n2562gat_reg/NET0131  ;
	input \n256gat_reg/NET0131  ;
	input \n2588gat_reg/NET0131  ;
	input \n2592gat_reg/NET0131  ;
	input \n2599gat_reg/NET0131  ;
	input \n2622gat_reg/NET0131  ;
	input \n2626gat_reg/NET0131  ;
	input \n2630gat_reg/NET0131  ;
	input \n2634gat_reg/NET0131  ;
	input \n2640gat_reg/NET0131  ;
	input \n2644gat_reg/NET0131  ;
	input \n2658gat_reg/NET0131  ;
	input \n271gat_reg/NET0131  ;
	input \n3065gat_pad  ;
	input \n3066gat_pad  ;
	input \n3067gat_pad  ;
	input \n3068gat_pad  ;
	input \n3069gat_pad  ;
	input \n3070gat_pad  ;
	input \n3071gat_pad  ;
	input \n3072gat_pad  ;
	input \n3073gat_pad  ;
	input \n3074gat_pad  ;
	input \n3075gat_pad  ;
	input \n3076gat_pad  ;
	input \n3077gat_pad  ;
	input \n3078gat_pad  ;
	input \n3079gat_pad  ;
	input \n3080gat_pad  ;
	input \n3081gat_pad  ;
	input \n3082gat_pad  ;
	input \n3083gat_pad  ;
	input \n3084gat_pad  ;
	input \n3085gat_pad  ;
	input \n3086gat_pad  ;
	input \n3087gat_pad  ;
	input \n3088gat_pad  ;
	input \n3089gat_pad  ;
	input \n3090gat_pad  ;
	input \n3091gat_pad  ;
	input \n3092gat_pad  ;
	input \n3093gat_pad  ;
	input \n3094gat_pad  ;
	input \n3095gat_pad  ;
	input \n3097gat_pad  ;
	input \n3098gat_pad  ;
	input \n3099gat_pad  ;
	input \n3100gat_pad  ;
	input \n314gat_reg/NET0131  ;
	input \n318gat_reg/NET0131  ;
	input \n322gat_reg/NET0131  ;
	input \n327gat_reg/NET0131  ;
	input \n331gat_reg/NET0131  ;
	input \n337gat_reg/NET0131  ;
	input \n341gat_reg/NET0131  ;
	input \n366gat_reg/NET0131  ;
	input \n384gat_reg/NET0131  ;
	input \n388gat_reg/NET0131  ;
	input \n398gat_reg/NET0131  ;
	input \n402gat_reg/NET0131  ;
	input \n463gat_reg/NET0131  ;
	input \n470gat_reg/NET0131  ;
	input \n553gat_reg/NET0131  ;
	input \n561gat_reg/NET0131  ;
	input \n580gat_reg/NET0131  ;
	input \n584gat_reg/NET0131  ;
	input \n614gat_reg/NET0131  ;
	input \n659gat_reg/NET0131  ;
	input \n667gat_reg/NET0131  ;
	input \n673gat_reg/NET0131  ;
	input \n680gat_reg/NET0131  ;
	input \n684gat_reg/NET0131  ;
	input \n699gat_reg/NET0131  ;
	input \n707gat_reg/NET0131  ;
	input \n777gat_reg/NET0131  ;
	input \n816gat_reg/NET0131  ;
	input \n820gat_reg/NET0131  ;
	input \n824gat_reg/NET0131  ;
	input \n830gat_reg/NET0131  ;
	input \n834gat_reg/NET0131  ;
	input \n838gat_reg/NET0131  ;
	input \n842gat_reg/NET0131  ;
	input \n846gat_reg/NET0131  ;
	input \n861gat_reg/NET0131  ;
	input \n865gat_reg/NET0131  ;
	input \n883gat_reg/NET0131  ;
	input \n919gat_reg/NET0131  ;
	input \n931gat_reg/NET0131  ;
	input \n957gat_reg/NET0131  ;
	output \_al_n0  ;
	output \g17_dup/_0_  ;
	output \g6952/_2_  ;
	output \g6953/_2_  ;
	output \g6961/_0_  ;
	output \g7076/_0_  ;
	output \g7077/_0_  ;
	output \g7079/_0_  ;
	output \g7081/_0_  ;
	output \g7082/_0_  ;
	output \g7083/_0_  ;
	output \g7146/_0_  ;
	output \g7147/_0_  ;
	output \g7148/_0_  ;
	output \g7149/_0_  ;
	output \g7150/_0_  ;
	output \g7151/_0_  ;
	output \g7152/_0_  ;
	output \g7153/_0_  ;
	output \g7154/_0_  ;
	output \g7156/_2_  ;
	output \g7161/_2_  ;
	output \g7165/_2_  ;
	output \g7174/_0_  ;
	output \g7180/_00_  ;
	output \g7182/_3_  ;
	output \g7191/_0_  ;
	output \g7204/_0_  ;
	output \g7209/_3_  ;
	output \g7220/_0_  ;
	output \g7229/_0_  ;
	output \g7233/_0_  ;
	output \g7234/_0_  ;
	output \g7235/_0_  ;
	output \g7236/_0_  ;
	output \g7237/_0_  ;
	output \g7238/_0_  ;
	output \g7241/_3_  ;
	output \g7264/_0_  ;
	output \g7265/_0_  ;
	output \g7266/_0_  ;
	output \g7267/_0_  ;
	output \g7268/_0_  ;
	output \g7301/_0_  ;
	output \g7326/_3_  ;
	output \g7350/_2_  ;
	output \g7352/_0_  ;
	output \g7356/_0_  ;
	output \g7359/_0_  ;
	output \g7389/_3_  ;
	output \g7417/_0_  ;
	output \g7418/_0_  ;
	output \g7419/_0_  ;
	output \g7444/_0_  ;
	output \g7445/_0_  ;
	output \g7449/_3_  ;
	output \g7451/_3_  ;
	output \g7454/_0_  ;
	output \g7467/_3_  ;
	output \g7476/_0_  ;
	output \g7480/_0_  ;
	output \g7494/_0_  ;
	output \g7509/_0_  ;
	output \g7514/_0_  ;
	output \g7517/_3_  ;
	output \g7524/_0_  ;
	output \g7558/_0_  ;
	output \g7560/_0_  ;
	output \g7561/_0_  ;
	output \g7563/_0_  ;
	output \g7567/_0_  ;
	output \g7572/_0_  ;
	output \g7579/_0_  ;
	output \g7605/_0_  ;
	output \g7625/_0_  ;
	output \g7627/_0_  ;
	output \g7671/_0_  ;
	output \g7675/_0_  ;
	output \g7689/_0_  ;
	output \g7697/_0_  ;
	output \g7743/_1_  ;
	output \g7764/_1_  ;
	output \g7769/_0_  ;
	output \g7771/_2_  ;
	output \g7779/_0_  ;
	output \g7852/_0_  ;
	output \g7873/_0_  ;
	output \g7884/_3_  ;
	output \g7889/_0_  ;
	output \g7902/_1_  ;
	output \g7992/_3_  ;
	output \g7994/_3_  ;
	output \g7996/_3_  ;
	output \g7998/_3_  ;
	output \g8000/_3_  ;
	output \g8002/_3_  ;
	output \g8004/_3_  ;
	output \g8006/_3_  ;
	output \g8008/_3_  ;
	output \g8150/_0_  ;
	output \g8151/_0_  ;
	output \g8157/_0_  ;
	output \g8163/_0_  ;
	output \g8172/_0_  ;
	output \g8197/_0_  ;
	output \g8211/_0_  ;
	output \g8223/_0_  ;
	output \g8237/_0_  ;
	output \g8251/_0_  ;
	output \g8261/_0_  ;
	output \g8272/_0_  ;
	output \g8287/_0_  ;
	output \g8647/_0_  ;
	output \g8671/_0_  ;
	output \g8672/_0_  ;
	output \g8735/_0_  ;
	output \g8766/_0_  ;
	output \g8811/_0_  ;
	output \g8821/_0_  ;
	output \g8856/_0_  ;
	output \g8858/_3_  ;
	output \g8868/_0_  ;
	output \g8880/_2_  ;
	output \g8886/_0_  ;
	output \g8900/_0_  ;
	output \g8932/_0_  ;
	output \g8991/_3_  ;
	output \g9014/_3_  ;
	output \g9074/_0_  ;
	output \g9091/_0_  ;
	output \g9105/_0_  ;
	output \g9107/_1_  ;
	output \g9111/_0_  ;
	output \n1332gat_reg/P0001  ;
	output \n1363gat_reg/P0001  ;
	output \n1394gat_reg/P0001  ;
	output \n1433gat_reg/P0001  ;
	output \n1775gat_reg/P0001  ;
	output \n2025gat_reg/P0001  ;
	output \n2029gat_reg/P0001  ;
	output \n2033gat_reg/P0001  ;
	output \n2044gat_reg/P0001  ;
	output \n2121gat_reg/P0001  ;
	output \n2125gat_reg/P0001  ;
	output \n2458gat_reg/P0001  ;
	output \n2472gat_reg/P0001  ;
	output \n2592gat_reg/P0001  ;
	output \n3104gat_pad  ;
	output \n3105gat_pad  ;
	output \n3106gat_pad  ;
	output \n3107gat_pad  ;
	output \n3108gat_pad  ;
	output \n3109gat_pad  ;
	output \n3110gat_pad  ;
	output \n3111gat_pad  ;
	output \n3112gat_pad  ;
	output \n3113gat_pad  ;
	output \n3114gat_pad  ;
	output \n3116gat_pad  ;
	output \n3117gat_pad  ;
	output \n3118gat_pad  ;
	output \n3119gat_pad  ;
	output \n3120gat_pad  ;
	output \n3121gat_pad  ;
	output \n3122gat_pad  ;
	output \n3123gat_pad  ;
	output \n3124gat_pad  ;
	output \n3125gat_pad  ;
	output \n3126gat_pad  ;
	output \n3127gat_pad  ;
	output \n3128gat_pad  ;
	output \n3130gat_pad  ;
	output \n3131gat_pad  ;
	output \n3132gat_pad  ;
	output \n3133gat_pad  ;
	output \n3134gat_pad  ;
	output \n3135gat_pad  ;
	output \n3136gat_pad  ;
	output \n3137gat_pad  ;
	output \n3138gat_pad  ;
	output \n3140gat_pad  ;
	output \n3142gat_pad  ;
	output \n3143gat_pad  ;
	output \n3144gat_pad  ;
	output \n3145gat_pad  ;
	output \n3146gat_pad  ;
	output \n3147gat_pad  ;
	output \n3148gat_pad  ;
	output \n3149gat_pad  ;
	output \n3150gat_pad  ;
	output \n3151gat_pad  ;
	output \n684gat_reg/P0001  ;
	output \n824gat_reg/P0001  ;
	output \n883gat_reg/P0001  ;
	wire _w896_ ;
	wire _w895_ ;
	wire _w894_ ;
	wire _w893_ ;
	wire _w892_ ;
	wire _w891_ ;
	wire _w890_ ;
	wire _w889_ ;
	wire _w888_ ;
	wire _w887_ ;
	wire _w886_ ;
	wire _w885_ ;
	wire _w884_ ;
	wire _w883_ ;
	wire _w882_ ;
	wire _w881_ ;
	wire _w880_ ;
	wire _w879_ ;
	wire _w878_ ;
	wire _w877_ ;
	wire _w876_ ;
	wire _w875_ ;
	wire _w874_ ;
	wire _w873_ ;
	wire _w872_ ;
	wire _w871_ ;
	wire _w870_ ;
	wire _w869_ ;
	wire _w868_ ;
	wire _w867_ ;
	wire _w866_ ;
	wire _w865_ ;
	wire _w864_ ;
	wire _w863_ ;
	wire _w862_ ;
	wire _w861_ ;
	wire _w860_ ;
	wire _w859_ ;
	wire _w858_ ;
	wire _w857_ ;
	wire _w856_ ;
	wire _w855_ ;
	wire _w854_ ;
	wire _w853_ ;
	wire _w852_ ;
	wire _w851_ ;
	wire _w850_ ;
	wire _w849_ ;
	wire _w848_ ;
	wire _w847_ ;
	wire _w846_ ;
	wire _w845_ ;
	wire _w844_ ;
	wire _w843_ ;
	wire _w842_ ;
	wire _w841_ ;
	wire _w840_ ;
	wire _w839_ ;
	wire _w838_ ;
	wire _w837_ ;
	wire _w836_ ;
	wire _w835_ ;
	wire _w834_ ;
	wire _w833_ ;
	wire _w832_ ;
	wire _w831_ ;
	wire _w830_ ;
	wire _w829_ ;
	wire _w828_ ;
	wire _w827_ ;
	wire _w826_ ;
	wire _w825_ ;
	wire _w824_ ;
	wire _w823_ ;
	wire _w822_ ;
	wire _w821_ ;
	wire _w820_ ;
	wire _w819_ ;
	wire _w818_ ;
	wire _w817_ ;
	wire _w816_ ;
	wire _w815_ ;
	wire _w814_ ;
	wire _w813_ ;
	wire _w812_ ;
	wire _w811_ ;
	wire _w810_ ;
	wire _w809_ ;
	wire _w808_ ;
	wire _w807_ ;
	wire _w806_ ;
	wire _w805_ ;
	wire _w804_ ;
	wire _w803_ ;
	wire _w802_ ;
	wire _w801_ ;
	wire _w800_ ;
	wire _w799_ ;
	wire _w798_ ;
	wire _w797_ ;
	wire _w796_ ;
	wire _w795_ ;
	wire _w794_ ;
	wire _w793_ ;
	wire _w792_ ;
	wire _w791_ ;
	wire _w790_ ;
	wire _w789_ ;
	wire _w788_ ;
	wire _w787_ ;
	wire _w786_ ;
	wire _w785_ ;
	wire _w784_ ;
	wire _w783_ ;
	wire _w782_ ;
	wire _w781_ ;
	wire _w780_ ;
	wire _w779_ ;
	wire _w778_ ;
	wire _w777_ ;
	wire _w776_ ;
	wire _w775_ ;
	wire _w774_ ;
	wire _w773_ ;
	wire _w772_ ;
	wire _w771_ ;
	wire _w770_ ;
	wire _w769_ ;
	wire _w768_ ;
	wire _w767_ ;
	wire _w766_ ;
	wire _w765_ ;
	wire _w764_ ;
	wire _w763_ ;
	wire _w762_ ;
	wire _w761_ ;
	wire _w760_ ;
	wire _w759_ ;
	wire _w758_ ;
	wire _w757_ ;
	wire _w756_ ;
	wire _w755_ ;
	wire _w754_ ;
	wire _w753_ ;
	wire _w752_ ;
	wire _w751_ ;
	wire _w750_ ;
	wire _w749_ ;
	wire _w748_ ;
	wire _w747_ ;
	wire _w746_ ;
	wire _w745_ ;
	wire _w744_ ;
	wire _w743_ ;
	wire _w742_ ;
	wire _w741_ ;
	wire _w740_ ;
	wire _w455_ ;
	wire _w454_ ;
	wire _w453_ ;
	wire _w452_ ;
	wire _w451_ ;
	wire _w450_ ;
	wire _w449_ ;
	wire _w448_ ;
	wire _w447_ ;
	wire _w446_ ;
	wire _w445_ ;
	wire _w444_ ;
	wire _w443_ ;
	wire _w442_ ;
	wire _w441_ ;
	wire _w440_ ;
	wire _w439_ ;
	wire _w438_ ;
	wire _w437_ ;
	wire _w436_ ;
	wire _w435_ ;
	wire _w434_ ;
	wire _w433_ ;
	wire _w432_ ;
	wire _w431_ ;
	wire _w430_ ;
	wire _w429_ ;
	wire _w428_ ;
	wire _w427_ ;
	wire _w426_ ;
	wire _w425_ ;
	wire _w424_ ;
	wire _w423_ ;
	wire _w422_ ;
	wire _w421_ ;
	wire _w420_ ;
	wire _w419_ ;
	wire _w418_ ;
	wire _w417_ ;
	wire _w416_ ;
	wire _w415_ ;
	wire _w413_ ;
	wire _w411_ ;
	wire _w409_ ;
	wire _w407_ ;
	wire _w405_ ;
	wire _w404_ ;
	wire _w402_ ;
	wire _w401_ ;
	wire _w400_ ;
	wire _w398_ ;
	wire _w396_ ;
	wire _w395_ ;
	wire _w394_ ;
	wire _w393_ ;
	wire _w392_ ;
	wire _w391_ ;
	wire _w390_ ;
	wire _w388_ ;
	wire _w386_ ;
	wire _w385_ ;
	wire _w383_ ;
	wire _w382_ ;
	wire _w381_ ;
	wire _w379_ ;
	wire _w378_ ;
	wire _w376_ ;
	wire _w375_ ;
	wire _w374_ ;
	wire _w373_ ;
	wire _w372_ ;
	wire _w370_ ;
	wire _w369_ ;
	wire _w367_ ;
	wire _w366_ ;
	wire _w364_ ;
	wire _w362_ ;
	wire _w361_ ;
	wire _w359_ ;
	wire _w358_ ;
	wire _w357_ ;
	wire _w355_ ;
	wire _w353_ ;
	wire _w352_ ;
	wire _w351_ ;
	wire _w350_ ;
	wire _w348_ ;
	wire _w347_ ;
	wire _w346_ ;
	wire _w345_ ;
	wire _w344_ ;
	wire _w343_ ;
	wire _w341_ ;
	wire _w339_ ;
	wire _w338_ ;
	wire _w336_ ;
	wire _w335_ ;
	wire _w334_ ;
	wire _w332_ ;
	wire _w331_ ;
	wire _w330_ ;
	wire _w329_ ;
	wire _w327_ ;
	wire _w326_ ;
	wire _w256_ ;
	wire _w254_ ;
	wire _w384_ ;
	wire _w127_ ;
	wire _w668_ ;
	wire _w252_ ;
	wire _w251_ ;
	wire _w249_ ;
	wire _w247_ ;
	wire _w377_ ;
	wire _w120_ ;
	wire _w661_ ;
	wire _w237_ ;
	wire _w235_ ;
	wire _w365_ ;
	wire _w108_ ;
	wire _w649_ ;
	wire _w231_ ;
	wire _w223_ ;
	wire _w414_ ;
	wire _w157_ ;
	wire _w698_ ;
	wire _w284_ ;
	wire _w412_ ;
	wire _w155_ ;
	wire _w696_ ;
	wire _w282_ ;
	wire _w410_ ;
	wire _w153_ ;
	wire _w694_ ;
	wire _w406_ ;
	wire _w149_ ;
	wire _w690_ ;
	wire _w397_ ;
	wire _w140_ ;
	wire _w681_ ;
	wire _w267_ ;
	wire _w250_ ;
	wire _w380_ ;
	wire _w123_ ;
	wire _w664_ ;
	wire _w389_ ;
	wire _w132_ ;
	wire _w673_ ;
	wire _w259_ ;
	wire _w215_ ;
	wire _w354_ ;
	wire _w97_ ;
	wire _w638_ ;
	wire _w243_ ;
	wire _w320_ ;
	wire _w257_ ;
	wire _w387_ ;
	wire _w130_ ;
	wire _w671_ ;
	wire _w337_ ;
	wire _w80_ ;
	wire _w621_ ;
	wire _w225_ ;
	wire _w305_ ;
	wire _w48_ ;
	wire _w589_ ;
	wire _w302_ ;
	wire _w255_ ;
	wire _w276_ ;
	wire _w19_ ;
	wire _w560_ ;
	wire _w403_ ;
	wire _w146_ ;
	wire _w687_ ;
	wire _w273_ ;
	wire _w363_ ;
	wire _w106_ ;
	wire _w647_ ;
	wire _w233_ ;
	wire _w316_ ;
	wire _w280_ ;
	wire _w23_ ;
	wire _w564_ ;
	wire _w277_ ;
	wire _w310_ ;
	wire _w342_ ;
	wire _w85_ ;
	wire _w626_ ;
	wire _w371_ ;
	wire _w114_ ;
	wire _w655_ ;
	wire _w253_ ;
	wire _w271_ ;
	wire _w333_ ;
	wire _w76_ ;
	wire _w617_ ;
	wire _w399_ ;
	wire _w142_ ;
	wire _w683_ ;
	wire _w269_ ;
	wire _w340_ ;
	wire _w83_ ;
	wire _w624_ ;
	wire _w408_ ;
	wire _w151_ ;
	wire _w692_ ;
	wire _w278_ ;
	wire _w349_ ;
	wire _w92_ ;
	wire _w633_ ;
	wire _w356_ ;
	wire _w99_ ;
	wire _w640_ ;
	wire _w221_ ;
	wire _w360_ ;
	wire _w103_ ;
	wire _w644_ ;
	wire _w229_ ;
	wire _w368_ ;
	wire _w111_ ;
	wire _w652_ ;
	wire _w318_ ;
	wire _w322_ ;
	wire _w248_ ;
	wire _w328_ ;
	wire _w71_ ;
	wire _w612_ ;
	wire _w68_ ;
	wire _w609_ ;
	wire _w325_ ;
	wire _w258_ ;
	wire _w260_ ;
	wire _w261_ ;
	wire _w262_ ;
	wire _w263_ ;
	wire _w264_ ;
	wire _w265_ ;
	wire _w266_ ;
	wire _w268_ ;
	wire _w270_ ;
	wire _w272_ ;
	wire _w17_ ;
	wire _w558_ ;
	wire _w274_ ;
	wire _w275_ ;
	wire _w279_ ;
	wire _w281_ ;
	wire _w26_ ;
	wire _w567_ ;
	wire _w283_ ;
	wire _w28_ ;
	wire _w569_ ;
	wire _w285_ ;
	wire _w286_ ;
	wire _w287_ ;
	wire _w288_ ;
	wire _w289_ ;
	wire _w290_ ;
	wire _w291_ ;
	wire _w292_ ;
	wire _w293_ ;
	wire _w294_ ;
	wire _w295_ ;
	wire _w296_ ;
	wire _w297_ ;
	wire _w298_ ;
	wire _w299_ ;
	wire _w300_ ;
	wire _w301_ ;
	wire _w303_ ;
	wire _w304_ ;
	wire _w306_ ;
	wire _w307_ ;
	wire _w51_ ;
	wire _w592_ ;
	wire _w308_ ;
	wire _w309_ ;
	wire _w311_ ;
	wire _w312_ ;
	wire _w56_ ;
	wire _w597_ ;
	wire _w313_ ;
	wire _w314_ ;
	wire _w315_ ;
	wire _w317_ ;
	wire _w62_ ;
	wire _w603_ ;
	wire _w319_ ;
	wire _w64_ ;
	wire _w605_ ;
	wire _w321_ ;
	wire _w66_ ;
	wire _w607_ ;
	wire _w323_ ;
	wire _w324_ ;
	wire _w456_ ;
	wire _w457_ ;
	wire _w458_ ;
	wire _w459_ ;
	wire _w460_ ;
	wire _w461_ ;
	wire _w462_ ;
	wire _w463_ ;
	wire _w464_ ;
	wire _w465_ ;
	wire _w466_ ;
	wire _w467_ ;
	wire _w468_ ;
	wire _w469_ ;
	wire _w470_ ;
	wire _w471_ ;
	wire _w472_ ;
	wire _w473_ ;
	wire _w474_ ;
	wire _w475_ ;
	wire _w476_ ;
	wire _w477_ ;
	wire _w478_ ;
	wire _w479_ ;
	wire _w480_ ;
	wire _w481_ ;
	wire _w482_ ;
	wire _w483_ ;
	wire _w484_ ;
	wire _w485_ ;
	wire _w486_ ;
	wire _w487_ ;
	wire _w488_ ;
	wire _w489_ ;
	wire _w490_ ;
	wire _w491_ ;
	wire _w492_ ;
	wire _w493_ ;
	wire _w494_ ;
	wire _w495_ ;
	wire _w496_ ;
	wire _w497_ ;
	wire _w498_ ;
	wire _w499_ ;
	wire _w500_ ;
	wire _w501_ ;
	wire _w502_ ;
	wire _w503_ ;
	wire _w504_ ;
	wire _w505_ ;
	wire _w506_ ;
	wire _w507_ ;
	wire _w508_ ;
	wire _w509_ ;
	wire _w510_ ;
	wire _w511_ ;
	wire _w512_ ;
	wire _w513_ ;
	wire _w514_ ;
	wire _w515_ ;
	wire _w516_ ;
	wire _w517_ ;
	wire _w518_ ;
	wire _w519_ ;
	wire _w520_ ;
	wire _w521_ ;
	wire _w522_ ;
	wire _w523_ ;
	wire _w524_ ;
	wire _w525_ ;
	wire _w526_ ;
	wire _w527_ ;
	wire _w528_ ;
	wire _w529_ ;
	wire _w530_ ;
	wire _w531_ ;
	wire _w532_ ;
	wire _w533_ ;
	wire _w534_ ;
	wire _w535_ ;
	wire _w536_ ;
	wire _w537_ ;
	wire _w538_ ;
	wire _w539_ ;
	wire _w540_ ;
	wire _w541_ ;
	wire _w542_ ;
	wire _w543_ ;
	wire _w544_ ;
	wire _w545_ ;
	wire _w546_ ;
	wire _w547_ ;
	wire _w548_ ;
	wire _w549_ ;
	wire _w550_ ;
	wire _w551_ ;
	wire _w552_ ;
	wire _w553_ ;
	wire _w554_ ;
	wire _w555_ ;
	wire _w556_ ;
	wire _w557_ ;
	wire _w559_ ;
	wire _w561_ ;
	wire _w562_ ;
	wire _w563_ ;
	wire _w565_ ;
	wire _w566_ ;
	wire _w568_ ;
	wire _w570_ ;
	wire _w571_ ;
	wire _w572_ ;
	wire _w573_ ;
	wire _w574_ ;
	wire _w575_ ;
	wire _w576_ ;
	wire _w577_ ;
	wire _w578_ ;
	wire _w579_ ;
	wire _w580_ ;
	wire _w581_ ;
	wire _w582_ ;
	wire _w583_ ;
	wire _w584_ ;
	wire _w585_ ;
	wire _w586_ ;
	wire _w587_ ;
	wire _w588_ ;
	wire _w590_ ;
	wire _w591_ ;
	wire _w593_ ;
	wire _w594_ ;
	wire _w595_ ;
	wire _w596_ ;
	wire _w598_ ;
	wire _w599_ ;
	wire _w600_ ;
	wire _w601_ ;
	wire _w602_ ;
	wire _w604_ ;
	wire _w606_ ;
	wire _w608_ ;
	wire _w610_ ;
	wire _w611_ ;
	wire _w613_ ;
	wire _w614_ ;
	wire _w615_ ;
	wire _w616_ ;
	wire _w618_ ;
	wire _w619_ ;
	wire _w620_ ;
	wire _w622_ ;
	wire _w623_ ;
	wire _w625_ ;
	wire _w627_ ;
	wire _w628_ ;
	wire _w629_ ;
	wire _w630_ ;
	wire _w631_ ;
	wire _w632_ ;
	wire _w634_ ;
	wire _w635_ ;
	wire _w636_ ;
	wire _w637_ ;
	wire _w639_ ;
	wire _w641_ ;
	wire _w642_ ;
	wire _w643_ ;
	wire _w645_ ;
	wire _w646_ ;
	wire _w648_ ;
	wire _w650_ ;
	wire _w651_ ;
	wire _w653_ ;
	wire _w654_ ;
	wire _w656_ ;
	wire _w657_ ;
	wire _w658_ ;
	wire _w659_ ;
	wire _w660_ ;
	wire _w662_ ;
	wire _w663_ ;
	wire _w665_ ;
	wire _w666_ ;
	wire _w667_ ;
	wire _w669_ ;
	wire _w670_ ;
	wire _w672_ ;
	wire _w674_ ;
	wire _w675_ ;
	wire _w676_ ;
	wire _w677_ ;
	wire _w678_ ;
	wire _w679_ ;
	wire _w680_ ;
	wire _w682_ ;
	wire _w684_ ;
	wire _w685_ ;
	wire _w686_ ;
	wire _w688_ ;
	wire _w689_ ;
	wire _w691_ ;
	wire _w693_ ;
	wire _w695_ ;
	wire _w697_ ;
	wire _w699_ ;
	wire _w700_ ;
	wire _w701_ ;
	wire _w702_ ;
	wire _w703_ ;
	wire _w704_ ;
	wire _w705_ ;
	wire _w706_ ;
	wire _w707_ ;
	wire _w708_ ;
	wire _w709_ ;
	wire _w710_ ;
	wire _w711_ ;
	wire _w712_ ;
	wire _w713_ ;
	wire _w714_ ;
	wire _w715_ ;
	wire _w716_ ;
	wire _w717_ ;
	wire _w718_ ;
	wire _w719_ ;
	wire _w720_ ;
	wire _w721_ ;
	wire _w722_ ;
	wire _w723_ ;
	wire _w724_ ;
	wire _w725_ ;
	wire _w726_ ;
	wire _w727_ ;
	wire _w728_ ;
	wire _w729_ ;
	wire _w730_ ;
	wire _w731_ ;
	wire _w732_ ;
	wire _w733_ ;
	wire _w734_ ;
	wire _w735_ ;
	wire _w736_ ;
	wire _w737_ ;
	wire _w738_ ;
	wire _w739_ ;
	LUT1 #(
		.INIT('h1)
	) name0 (
		\n1316gat_reg/NET0131 ,
		_w17_
	);
	LUT1 #(
		.INIT('h1)
	) name1 (
		\n1332gat_reg/NET0131 ,
		_w19_
	);
	LUT1 #(
		.INIT('h1)
	) name2 (
		\n1363gat_reg/NET0131 ,
		_w23_
	);
	LUT1 #(
		.INIT('h1)
	) name3 (
		\n1394gat_reg/NET0131 ,
		_w26_
	);
	LUT1 #(
		.INIT('h1)
	) name4 (
		\n1433gat_reg/NET0131 ,
		_w28_
	);
	LUT1 #(
		.INIT('h1)
	) name5 (
		\n1775gat_reg/NET0131 ,
		_w48_
	);
	LUT1 #(
		.INIT('h1)
	) name6 (
		\n1821gat_reg/NET0131 ,
		_w51_
	);
	LUT1 #(
		.INIT('h1)
	) name7 (
		\n1871gat_reg/NET0131 ,
		_w56_
	);
	LUT1 #(
		.INIT('h1)
	) name8 (
		\n2025gat_reg/NET0131 ,
		_w62_
	);
	LUT1 #(
		.INIT('h1)
	) name9 (
		\n2029gat_reg/NET0131 ,
		_w64_
	);
	LUT1 #(
		.INIT('h1)
	) name10 (
		\n2033gat_reg/NET0131 ,
		_w66_
	);
	LUT1 #(
		.INIT('h1)
	) name11 (
		\n2037gat_reg/NET0131 ,
		_w68_
	);
	LUT1 #(
		.INIT('h1)
	) name12 (
		\n2044gat_reg/NET0131 ,
		_w71_
	);
	LUT1 #(
		.INIT('h1)
	) name13 (
		\n2095gat_reg/NET0131 ,
		_w76_
	);
	LUT1 #(
		.INIT('h1)
	) name14 (
		\n2110gat_reg/NET0131 ,
		_w80_
	);
	LUT1 #(
		.INIT('h1)
	) name15 (
		\n2121gat_reg/NET0131 ,
		_w83_
	);
	LUT1 #(
		.INIT('h1)
	) name16 (
		\n2125gat_reg/NET0131 ,
		_w85_
	);
	LUT1 #(
		.INIT('h1)
	) name17 (
		\n2176gat_reg/NET0131 ,
		_w92_
	);
	LUT1 #(
		.INIT('h1)
	) name18 (
		\n2203gat_reg/NET0131 ,
		_w97_
	);
	LUT1 #(
		.INIT('h1)
	) name19 (
		\n2207gat_reg/NET0131 ,
		_w99_
	);
	LUT1 #(
		.INIT('h1)
	) name20 (
		\n2270gat_reg/NET0131 ,
		_w103_
	);
	LUT1 #(
		.INIT('h1)
	) name21 (
		\n2339gat_reg/NET0131 ,
		_w106_
	);
	LUT1 #(
		.INIT('h1)
	) name22 (
		\n2343gat_reg/NET0131 ,
		_w108_
	);
	LUT1 #(
		.INIT('h1)
	) name23 (
		\n2390gat_reg/NET0131 ,
		_w111_
	);
	LUT1 #(
		.INIT('h1)
	) name24 (
		\n2399gat_reg/NET0131 ,
		_w114_
	);
	LUT1 #(
		.INIT('h1)
	) name25 (
		\n2450gat_reg/NET0131 ,
		_w120_
	);
	LUT1 #(
		.INIT('h1)
	) name26 (
		\n2458gat_reg/NET0131 ,
		_w123_
	);
	LUT1 #(
		.INIT('h1)
	) name27 (
		\n2472gat_reg/NET0131 ,
		_w127_
	);
	LUT1 #(
		.INIT('h1)
	) name28 (
		\n2490gat_reg/NET0131 ,
		_w130_
	);
	LUT1 #(
		.INIT('h1)
	) name29 (
		\n2495gat_reg/NET0131 ,
		_w132_
	);
	LUT1 #(
		.INIT('h1)
	) name30 (
		\n2543gat_reg/NET0131 ,
		_w140_
	);
	LUT1 #(
		.INIT('h1)
	) name31 (
		\n2562gat_reg/NET0131 ,
		_w142_
	);
	LUT1 #(
		.INIT('h1)
	) name32 (
		\n2592gat_reg/NET0131 ,
		_w146_
	);
	LUT1 #(
		.INIT('h1)
	) name33 (
		\n2622gat_reg/NET0131 ,
		_w149_
	);
	LUT1 #(
		.INIT('h1)
	) name34 (
		\n2626gat_reg/NET0131 ,
		_w151_
	);
	LUT1 #(
		.INIT('h1)
	) name35 (
		\n2630gat_reg/NET0131 ,
		_w153_
	);
	LUT1 #(
		.INIT('h1)
	) name36 (
		\n2634gat_reg/NET0131 ,
		_w155_
	);
	LUT1 #(
		.INIT('h1)
	) name37 (
		\n2640gat_reg/NET0131 ,
		_w157_
	);
	LUT1 #(
		.INIT('h1)
	) name38 (
		\n614gat_reg/NET0131 ,
		_w215_
	);
	LUT1 #(
		.INIT('h1)
	) name39 (
		\n684gat_reg/NET0131 ,
		_w221_
	);
	LUT1 #(
		.INIT('h1)
	) name40 (
		\n699gat_reg/NET0131 ,
		_w223_
	);
	LUT1 #(
		.INIT('h1)
	) name41 (
		\n707gat_reg/NET0131 ,
		_w225_
	);
	LUT1 #(
		.INIT('h1)
	) name42 (
		\n820gat_reg/NET0131 ,
		_w229_
	);
	LUT1 #(
		.INIT('h1)
	) name43 (
		\n824gat_reg/NET0131 ,
		_w231_
	);
	LUT1 #(
		.INIT('h1)
	) name44 (
		\n830gat_reg/NET0131 ,
		_w233_
	);
	LUT1 #(
		.INIT('h1)
	) name45 (
		\n834gat_reg/NET0131 ,
		_w235_
	);
	LUT1 #(
		.INIT('h1)
	) name46 (
		\n838gat_reg/NET0131 ,
		_w237_
	);
	LUT1 #(
		.INIT('h1)
	) name47 (
		\n883gat_reg/NET0131 ,
		_w243_
	);
	LUT2 #(
		.INIT('h2)
	) name48 (
		\n398gat_reg/NET0131 ,
		\n402gat_reg/NET0131 ,
		_w247_
	);
	LUT2 #(
		.INIT('h4)
	) name49 (
		\n2454gat_reg/NET0131 ,
		\n846gat_reg/NET0131 ,
		_w248_
	);
	LUT4 #(
		.INIT('h0400)
	) name50 (
		\n2454gat_reg/NET0131 ,
		\n398gat_reg/NET0131 ,
		\n402gat_reg/NET0131 ,
		\n846gat_reg/NET0131 ,
		_w249_
	);
	LUT2 #(
		.INIT('h6)
	) name51 (
		\n553gat_reg/NET0131 ,
		\n777gat_reg/NET0131 ,
		_w250_
	);
	LUT3 #(
		.INIT('h69)
	) name52 (
		\n314gat_reg/NET0131 ,
		\n366gat_reg/NET0131 ,
		\n561gat_reg/NET0131 ,
		_w251_
	);
	LUT2 #(
		.INIT('h6)
	) name53 (
		_w250_,
		_w251_,
		_w252_
	);
	LUT4 #(
		.INIT('h135f)
	) name54 (
		\n3087gat_pad ,
		\n3088gat_pad ,
		\n3093gat_pad ,
		\n3095gat_pad ,
		_w253_
	);
	LUT2 #(
		.INIT('h8)
	) name55 (
		\n3087gat_pad ,
		\n3095gat_pad ,
		_w254_
	);
	LUT4 #(
		.INIT('h135f)
	) name56 (
		\n3086gat_pad ,
		\n3087gat_pad ,
		\n3093gat_pad ,
		\n3095gat_pad ,
		_w255_
	);
	LUT4 #(
		.INIT('h135f)
	) name57 (
		\n3085gat_pad ,
		\n3086gat_pad ,
		\n3093gat_pad ,
		\n3095gat_pad ,
		_w256_
	);
	LUT3 #(
		.INIT('h02)
	) name58 (
		_w253_,
		_w255_,
		_w256_,
		_w257_
	);
	LUT3 #(
		.INIT('h69)
	) name59 (
		\n318gat_reg/NET0131 ,
		\n322gat_reg/NET0131 ,
		\n659gat_reg/NET0131 ,
		_w258_
	);
	LUT3 #(
		.INIT('h7b)
	) name60 (
		_w252_,
		_w257_,
		_w258_,
		_w259_
	);
	LUT4 #(
		.INIT('h0afc)
	) name61 (
		\n820gat_reg/NET0131 ,
		\n842gat_reg/NET0131 ,
		_w253_,
		_w255_,
		_w260_
	);
	LUT4 #(
		.INIT('h0100)
	) name62 (
		\n1241gat_reg/NET0131 ,
		_w253_,
		_w255_,
		_w256_,
		_w261_
	);
	LUT4 #(
		.INIT('h0800)
	) name63 (
		\n673gat_reg/NET0131 ,
		_w253_,
		_w255_,
		_w256_,
		_w262_
	);
	LUT4 #(
		.INIT('h000e)
	) name64 (
		_w256_,
		_w260_,
		_w261_,
		_w262_,
		_w263_
	);
	LUT3 #(
		.INIT('h10)
	) name65 (
		\n3083gat_pad ,
		\n3084gat_pad ,
		\n3093gat_pad ,
		_w264_
	);
	LUT2 #(
		.INIT('h1)
	) name66 (
		\n3085gat_pad ,
		\n3086gat_pad ,
		_w265_
	);
	LUT3 #(
		.INIT('h0e)
	) name67 (
		\n3085gat_pad ,
		\n3086gat_pad ,
		\n3088gat_pad ,
		_w266_
	);
	LUT3 #(
		.INIT('h01)
	) name68 (
		\n3083gat_pad ,
		\n3084gat_pad ,
		\n3085gat_pad ,
		_w267_
	);
	LUT4 #(
		.INIT('h8000)
	) name69 (
		\n3086gat_pad ,
		\n3087gat_pad ,
		\n3088gat_pad ,
		\n3095gat_pad ,
		_w268_
	);
	LUT4 #(
		.INIT('h0777)
	) name70 (
		_w264_,
		_w266_,
		_w267_,
		_w268_,
		_w269_
	);
	LUT3 #(
		.INIT('h07)
	) name71 (
		_w259_,
		_w263_,
		_w269_,
		_w270_
	);
	LUT3 #(
		.INIT('he0)
	) name72 (
		\n3086gat_pad ,
		\n3087gat_pad ,
		\n3095gat_pad ,
		_w271_
	);
	LUT2 #(
		.INIT('h8)
	) name73 (
		_w267_,
		_w271_,
		_w272_
	);
	LUT4 #(
		.INIT('h8000)
	) name74 (
		\n3085gat_pad ,
		\n3086gat_pad ,
		\n3087gat_pad ,
		\n3093gat_pad ,
		_w273_
	);
	LUT4 #(
		.INIT('h0008)
	) name75 (
		\n3088gat_pad ,
		_w264_,
		_w265_,
		_w273_,
		_w274_
	);
	LUT2 #(
		.INIT('h1)
	) name76 (
		_w272_,
		_w274_,
		_w275_
	);
	LUT4 #(
		.INIT('h9669)
	) name77 (
		\n1035gat_reg/NET0131 ,
		\n1121gat_reg/NET0131 ,
		\n1226gat_reg/NET0131 ,
		\n1282gat_reg/NET0131 ,
		_w276_
	);
	LUT2 #(
		.INIT('h9)
	) name78 (
		\n1135gat_reg/NET0131 ,
		\n931gat_reg/NET0131 ,
		_w277_
	);
	LUT2 #(
		.INIT('h9)
	) name79 (
		\n1045gat_reg/NET0131 ,
		\n1072gat_reg/NET0131 ,
		_w278_
	);
	LUT4 #(
		.INIT('h0200)
	) name80 (
		_w253_,
		_w255_,
		_w256_,
		_w278_,
		_w279_
	);
	LUT3 #(
		.INIT('h6f)
	) name81 (
		_w276_,
		_w277_,
		_w279_,
		_w280_
	);
	LUT4 #(
		.INIT('h6006)
	) name82 (
		\n1045gat_reg/NET0131 ,
		\n1072gat_reg/NET0131 ,
		\n1135gat_reg/NET0131 ,
		\n931gat_reg/NET0131 ,
		_w281_
	);
	LUT4 #(
		.INIT('h0200)
	) name83 (
		_w253_,
		_w255_,
		_w256_,
		_w281_,
		_w282_
	);
	LUT4 #(
		.INIT('h0660)
	) name84 (
		\n1045gat_reg/NET0131 ,
		\n1072gat_reg/NET0131 ,
		\n1135gat_reg/NET0131 ,
		\n931gat_reg/NET0131 ,
		_w283_
	);
	LUT4 #(
		.INIT('h0200)
	) name85 (
		_w253_,
		_w255_,
		_w256_,
		_w283_,
		_w284_
	);
	LUT3 #(
		.INIT('h1b)
	) name86 (
		_w276_,
		_w282_,
		_w284_,
		_w285_
	);
	LUT4 #(
		.INIT('h0100)
	) name87 (
		\n842gat_reg/NET0131 ,
		_w253_,
		_w255_,
		_w256_,
		_w286_
	);
	LUT4 #(
		.INIT('h0010)
	) name88 (
		\n830gat_reg/NET0131 ,
		_w253_,
		_w255_,
		_w256_,
		_w287_
	);
	LUT2 #(
		.INIT('h1)
	) name89 (
		_w286_,
		_w287_,
		_w288_
	);
	LUT4 #(
		.INIT('h1555)
	) name90 (
		_w275_,
		_w280_,
		_w285_,
		_w288_,
		_w289_
	);
	LUT2 #(
		.INIT('he)
	) name91 (
		_w270_,
		_w289_,
		_w290_
	);
	LUT3 #(
		.INIT('h80)
	) name92 (
		\n2464gat_reg/NET0131 ,
		\n2476gat_reg/NET0131 ,
		\n2518gat_reg/NET0131 ,
		_w291_
	);
	LUT4 #(
		.INIT('h0080)
	) name93 (
		\n2468gat_reg/NET0131 ,
		\n2526gat_reg/NET0131 ,
		\n2599gat_reg/NET0131 ,
		\n3090gat_pad ,
		_w292_
	);
	LUT2 #(
		.INIT('h7)
	) name94 (
		_w291_,
		_w292_,
		_w293_
	);
	LUT4 #(
		.INIT('h96ff)
	) name95 (
		\n318gat_reg/NET0131 ,
		\n322gat_reg/NET0131 ,
		\n659gat_reg/NET0131 ,
		\n667gat_reg/NET0131 ,
		_w294_
	);
	LUT4 #(
		.INIT('h9600)
	) name96 (
		\n318gat_reg/NET0131 ,
		\n322gat_reg/NET0131 ,
		\n659gat_reg/NET0131 ,
		\n667gat_reg/NET0131 ,
		_w295_
	);
	LUT4 #(
		.INIT('h90f6)
	) name97 (
		_w250_,
		_w251_,
		_w294_,
		_w295_,
		_w296_
	);
	LUT4 #(
		.INIT('h0096)
	) name98 (
		\n318gat_reg/NET0131 ,
		\n322gat_reg/NET0131 ,
		\n659gat_reg/NET0131 ,
		\n667gat_reg/NET0131 ,
		_w297_
	);
	LUT4 #(
		.INIT('hff96)
	) name99 (
		\n318gat_reg/NET0131 ,
		\n322gat_reg/NET0131 ,
		\n659gat_reg/NET0131 ,
		\n667gat_reg/NET0131 ,
		_w298_
	);
	LUT4 #(
		.INIT('h6f09)
	) name100 (
		_w250_,
		_w251_,
		_w297_,
		_w298_,
		_w299_
	);
	LUT2 #(
		.INIT('h8)
	) name101 (
		_w296_,
		_w299_,
		_w300_
	);
	LUT4 #(
		.INIT('h135f)
	) name102 (
		\n3069gat_pad ,
		\n3078gat_pad ,
		\n3093gat_pad ,
		\n3095gat_pad ,
		_w301_
	);
	LUT4 #(
		.INIT('heca0)
	) name103 (
		\n3069gat_pad ,
		\n3078gat_pad ,
		\n3093gat_pad ,
		\n3095gat_pad ,
		_w302_
	);
	LUT2 #(
		.INIT('h2)
	) name104 (
		\n2155gat_reg/NET0131 ,
		\n2622gat_reg/NET0131 ,
		_w303_
	);
	LUT4 #(
		.INIT('h0800)
	) name105 (
		\n2490gat_reg/NET0131 ,
		\n2543gat_reg/NET0131 ,
		\n2626gat_reg/NET0131 ,
		\n2630gat_reg/NET0131 ,
		_w304_
	);
	LUT2 #(
		.INIT('h4)
	) name106 (
		\n2543gat_reg/NET0131 ,
		\n2630gat_reg/NET0131 ,
		_w305_
	);
	LUT4 #(
		.INIT('h0100)
	) name107 (
		\n2155gat_reg/NET0131 ,
		\n2490gat_reg/NET0131 ,
		\n2622gat_reg/NET0131 ,
		\n2626gat_reg/NET0131 ,
		_w306_
	);
	LUT4 #(
		.INIT('h0777)
	) name108 (
		_w303_,
		_w304_,
		_w305_,
		_w306_,
		_w307_
	);
	LUT2 #(
		.INIT('h1)
	) name109 (
		\n2203gat_reg/NET0131 ,
		\n2207gat_reg/NET0131 ,
		_w308_
	);
	LUT3 #(
		.INIT('h40)
	) name110 (
		\n2343gat_reg/NET0131 ,
		\n2399gat_reg/NET0131 ,
		\n2562gat_reg/NET0131 ,
		_w309_
	);
	LUT2 #(
		.INIT('h8)
	) name111 (
		_w308_,
		_w309_,
		_w310_
	);
	LUT2 #(
		.INIT('h8)
	) name112 (
		\n398gat_reg/NET0131 ,
		\n402gat_reg/NET0131 ,
		_w311_
	);
	LUT3 #(
		.INIT('h04)
	) name113 (
		\n2454gat_reg/NET0131 ,
		\n846gat_reg/NET0131 ,
		\n919gat_reg/NET0131 ,
		_w312_
	);
	LUT2 #(
		.INIT('h8)
	) name114 (
		_w311_,
		_w312_,
		_w313_
	);
	LUT4 #(
		.INIT('h95ff)
	) name115 (
		\n398gat_reg/NET0131 ,
		\n402gat_reg/NET0131 ,
		\n919gat_reg/NET0131 ,
		_w248_,
		_w314_
	);
	LUT4 #(
		.INIT('h6a00)
	) name116 (
		\n398gat_reg/NET0131 ,
		\n402gat_reg/NET0131 ,
		\n919gat_reg/NET0131 ,
		_w248_,
		_w315_
	);
	LUT3 #(
		.INIT('h15)
	) name117 (
		\n2207gat_reg/NET0131 ,
		\n2343gat_reg/NET0131 ,
		\n2399gat_reg/NET0131 ,
		_w316_
	);
	LUT2 #(
		.INIT('h2)
	) name118 (
		\n2203gat_reg/NET0131 ,
		\n2207gat_reg/NET0131 ,
		_w317_
	);
	LUT3 #(
		.INIT('hcd)
	) name119 (
		\n2203gat_reg/NET0131 ,
		\n2207gat_reg/NET0131 ,
		\n2562gat_reg/NET0131 ,
		_w318_
	);
	LUT2 #(
		.INIT('h4)
	) name120 (
		_w316_,
		_w318_,
		_w319_
	);
	LUT4 #(
		.INIT('h0001)
	) name121 (
		_w307_,
		_w310_,
		_w314_,
		_w319_,
		_w320_
	);
	LUT2 #(
		.INIT('hd)
	) name122 (
		_w301_,
		_w320_,
		_w321_
	);
	LUT4 #(
		.INIT('h135f)
	) name123 (
		\n3070gat_pad ,
		\n3079gat_pad ,
		\n3093gat_pad ,
		\n3095gat_pad ,
		_w322_
	);
	LUT4 #(
		.INIT('heca0)
	) name124 (
		\n3070gat_pad ,
		\n3079gat_pad ,
		\n3093gat_pad ,
		\n3095gat_pad ,
		_w323_
	);
	LUT2 #(
		.INIT('hb)
	) name125 (
		_w320_,
		_w322_,
		_w324_
	);
	LUT4 #(
		.INIT('h135f)
	) name126 (
		\n3072gat_pad ,
		\n3081gat_pad ,
		\n3093gat_pad ,
		\n3095gat_pad ,
		_w325_
	);
	LUT4 #(
		.INIT('heca0)
	) name127 (
		\n3072gat_pad ,
		\n3081gat_pad ,
		\n3093gat_pad ,
		\n3095gat_pad ,
		_w326_
	);
	LUT2 #(
		.INIT('hb)
	) name128 (
		_w320_,
		_w325_,
		_w327_
	);
	LUT4 #(
		.INIT('h135f)
	) name129 (
		\n3071gat_pad ,
		\n3080gat_pad ,
		\n3093gat_pad ,
		\n3095gat_pad ,
		_w328_
	);
	LUT4 #(
		.INIT('heca0)
	) name130 (
		\n3071gat_pad ,
		\n3080gat_pad ,
		\n3093gat_pad ,
		\n3095gat_pad ,
		_w329_
	);
	LUT2 #(
		.INIT('hb)
	) name131 (
		_w320_,
		_w328_,
		_w330_
	);
	LUT4 #(
		.INIT('h135f)
	) name132 (
		\n3065gat_pad ,
		\n3074gat_pad ,
		\n3093gat_pad ,
		\n3095gat_pad ,
		_w331_
	);
	LUT4 #(
		.INIT('heca0)
	) name133 (
		\n3065gat_pad ,
		\n3074gat_pad ,
		\n3093gat_pad ,
		\n3095gat_pad ,
		_w332_
	);
	LUT2 #(
		.INIT('hb)
	) name134 (
		_w320_,
		_w331_,
		_w333_
	);
	LUT4 #(
		.INIT('h135f)
	) name135 (
		\n3073gat_pad ,
		\n3082gat_pad ,
		\n3093gat_pad ,
		\n3095gat_pad ,
		_w334_
	);
	LUT4 #(
		.INIT('heca0)
	) name136 (
		\n3073gat_pad ,
		\n3082gat_pad ,
		\n3093gat_pad ,
		\n3095gat_pad ,
		_w335_
	);
	LUT2 #(
		.INIT('hb)
	) name137 (
		_w320_,
		_w334_,
		_w336_
	);
	LUT4 #(
		.INIT('h0002)
	) name138 (
		\n1871gat_reg/NET0131 ,
		\n3083gat_pad ,
		\n3084gat_pad ,
		\n3085gat_pad ,
		_w337_
	);
	LUT3 #(
		.INIT('h80)
	) name139 (
		\n3087gat_pad ,
		\n3094gat_pad ,
		\n3095gat_pad ,
		_w338_
	);
	LUT3 #(
		.INIT('h20)
	) name140 (
		\n3086gat_pad ,
		\n3088gat_pad ,
		\n3095gat_pad ,
		_w339_
	);
	LUT3 #(
		.INIT('h80)
	) name141 (
		_w337_,
		_w338_,
		_w339_,
		_w340_
	);
	LUT4 #(
		.INIT('h0200)
	) name142 (
		\n1871gat_reg/NET0131 ,
		\n3083gat_pad ,
		\n3084gat_pad ,
		\n3093gat_pad ,
		_w341_
	);
	LUT2 #(
		.INIT('h4)
	) name143 (
		\n3087gat_pad ,
		\n3088gat_pad ,
		_w342_
	);
	LUT2 #(
		.INIT('h1)
	) name144 (
		\n3091gat_pad ,
		\n3092gat_pad ,
		_w343_
	);
	LUT4 #(
		.INIT('h8880)
	) name145 (
		\n3085gat_pad ,
		\n3086gat_pad ,
		\n3091gat_pad ,
		\n3092gat_pad ,
		_w344_
	);
	LUT3 #(
		.INIT('h80)
	) name146 (
		_w341_,
		_w342_,
		_w344_,
		_w345_
	);
	LUT3 #(
		.INIT('ha8)
	) name147 (
		\n3068gat_pad ,
		_w340_,
		_w345_,
		_w346_
	);
	LUT2 #(
		.INIT('he)
	) name148 (
		_w320_,
		_w346_,
		_w347_
	);
	LUT3 #(
		.INIT('ha8)
	) name149 (
		\n3065gat_pad ,
		_w340_,
		_w345_,
		_w348_
	);
	LUT2 #(
		.INIT('he)
	) name150 (
		_w320_,
		_w348_,
		_w349_
	);
	LUT3 #(
		.INIT('ha8)
	) name151 (
		\n3069gat_pad ,
		_w340_,
		_w345_,
		_w350_
	);
	LUT2 #(
		.INIT('he)
	) name152 (
		_w320_,
		_w350_,
		_w351_
	);
	LUT3 #(
		.INIT('ha8)
	) name153 (
		\n3066gat_pad ,
		_w340_,
		_w345_,
		_w352_
	);
	LUT2 #(
		.INIT('he)
	) name154 (
		_w320_,
		_w352_,
		_w353_
	);
	LUT3 #(
		.INIT('ha8)
	) name155 (
		\n3067gat_pad ,
		_w340_,
		_w345_,
		_w354_
	);
	LUT2 #(
		.INIT('he)
	) name156 (
		_w320_,
		_w354_,
		_w355_
	);
	LUT3 #(
		.INIT('ha8)
	) name157 (
		\n3070gat_pad ,
		_w340_,
		_w345_,
		_w356_
	);
	LUT2 #(
		.INIT('he)
	) name158 (
		_w320_,
		_w356_,
		_w357_
	);
	LUT3 #(
		.INIT('ha8)
	) name159 (
		\n3073gat_pad ,
		_w340_,
		_w345_,
		_w358_
	);
	LUT2 #(
		.INIT('he)
	) name160 (
		_w320_,
		_w358_,
		_w359_
	);
	LUT3 #(
		.INIT('ha8)
	) name161 (
		\n3072gat_pad ,
		_w340_,
		_w345_,
		_w360_
	);
	LUT2 #(
		.INIT('he)
	) name162 (
		_w320_,
		_w360_,
		_w361_
	);
	LUT3 #(
		.INIT('ha8)
	) name163 (
		\n3071gat_pad ,
		_w340_,
		_w345_,
		_w362_
	);
	LUT2 #(
		.INIT('he)
	) name164 (
		_w320_,
		_w362_,
		_w363_
	);
	LUT2 #(
		.INIT('h6)
	) name165 (
		\n2403gat_reg/NET0131 ,
		\n402gat_reg/NET0131 ,
		_w364_
	);
	LUT3 #(
		.INIT('h20)
	) name166 (
		\n2347gat_reg/NET0131 ,
		\n2407gat_reg/NET0131 ,
		\n398gat_reg/NET0131 ,
		_w365_
	);
	LUT2 #(
		.INIT('h1)
	) name167 (
		\n2394gat_reg/NET0131 ,
		\n2440gat_reg/NET0131 ,
		_w366_
	);
	LUT2 #(
		.INIT('h1)
	) name168 (
		\n846gat_reg/NET0131 ,
		\n919gat_reg/NET0131 ,
		_w367_
	);
	LUT2 #(
		.INIT('h4)
	) name169 (
		\n846gat_reg/NET0131 ,
		\n919gat_reg/NET0131 ,
		_w368_
	);
	LUT2 #(
		.INIT('h4)
	) name170 (
		\n2394gat_reg/NET0131 ,
		\n2440gat_reg/NET0131 ,
		_w369_
	);
	LUT2 #(
		.INIT('h2)
	) name171 (
		\n2394gat_reg/NET0131 ,
		\n2440gat_reg/NET0131 ,
		_w370_
	);
	LUT4 #(
		.INIT('hfbde)
	) name172 (
		\n2394gat_reg/NET0131 ,
		\n2440gat_reg/NET0131 ,
		\n846gat_reg/NET0131 ,
		\n919gat_reg/NET0131 ,
		_w371_
	);
	LUT3 #(
		.INIT('h04)
	) name173 (
		_w364_,
		_w365_,
		_w371_,
		_w372_
	);
	LUT2 #(
		.INIT('h8)
	) name174 (
		\n846gat_reg/NET0131 ,
		\n919gat_reg/NET0131 ,
		_w373_
	);
	LUT2 #(
		.INIT('h8)
	) name175 (
		\n2394gat_reg/NET0131 ,
		\n2440gat_reg/NET0131 ,
		_w374_
	);
	LUT4 #(
		.INIT('h8000)
	) name176 (
		\n2394gat_reg/NET0131 ,
		\n2440gat_reg/NET0131 ,
		\n846gat_reg/NET0131 ,
		\n919gat_reg/NET0131 ,
		_w375_
	);
	LUT3 #(
		.INIT('h40)
	) name177 (
		_w364_,
		_w365_,
		_w375_,
		_w376_
	);
	LUT3 #(
		.INIT('h04)
	) name178 (
		\n2347gat_reg/NET0131 ,
		\n2403gat_reg/NET0131 ,
		\n2407gat_reg/NET0131 ,
		_w377_
	);
	LUT2 #(
		.INIT('h8)
	) name179 (
		_w374_,
		_w377_,
		_w378_
	);
	LUT3 #(
		.INIT('h01)
	) name180 (
		_w372_,
		_w376_,
		_w378_,
		_w379_
	);
	LUT3 #(
		.INIT('he0)
	) name181 (
		\n1763gat_reg/NET0131 ,
		\n1880gat_reg/NET0131 ,
		\n2102gat_reg/NET0131 ,
		_w380_
	);
	LUT3 #(
		.INIT('h1f)
	) name182 (
		\n1763gat_reg/NET0131 ,
		\n1880gat_reg/NET0131 ,
		\n2102gat_reg/NET0131 ,
		_w381_
	);
	LUT2 #(
		.INIT('h8)
	) name183 (
		\n1850gat_reg/NET0131 ,
		\n2143gat_reg/NET0131 ,
		_w382_
	);
	LUT3 #(
		.INIT('h01)
	) name184 (
		\n1899gat_reg/NET0131 ,
		\n2061gat_reg/NET0131 ,
		\n2139gat_reg/NET0131 ,
		_w383_
	);
	LUT2 #(
		.INIT('h8)
	) name185 (
		_w382_,
		_w383_,
		_w384_
	);
	LUT3 #(
		.INIT('h80)
	) name186 (
		_w380_,
		_w382_,
		_w383_,
		_w385_
	);
	LUT4 #(
		.INIT('h10f0)
	) name187 (
		\n1763gat_reg/NET0131 ,
		\n1880gat_reg/NET0131 ,
		\n2061gat_reg/NET0131 ,
		\n2102gat_reg/NET0131 ,
		_w386_
	);
	LUT2 #(
		.INIT('h4)
	) name188 (
		\n1899gat_reg/NET0131 ,
		\n2139gat_reg/NET0131 ,
		_w387_
	);
	LUT4 #(
		.INIT('h1000)
	) name189 (
		\n1850gat_reg/NET0131 ,
		\n1899gat_reg/NET0131 ,
		\n2139gat_reg/NET0131 ,
		\n2143gat_reg/NET0131 ,
		_w388_
	);
	LUT2 #(
		.INIT('h8)
	) name190 (
		_w386_,
		_w388_,
		_w389_
	);
	LUT3 #(
		.INIT('h80)
	) name191 (
		\n1767gat_reg/NET0131 ,
		\n1834gat_reg/NET0131 ,
		\n1880gat_reg/NET0131 ,
		_w390_
	);
	LUT3 #(
		.INIT('h7f)
	) name192 (
		\n1767gat_reg/NET0131 ,
		\n1834gat_reg/NET0131 ,
		\n1880gat_reg/NET0131 ,
		_w391_
	);
	LUT3 #(
		.INIT('h0e)
	) name193 (
		_w385_,
		_w389_,
		_w390_,
		_w392_
	);
	LUT2 #(
		.INIT('h8)
	) name194 (
		\n1880gat_reg/NET0131 ,
		\n2021gat_reg/NET0131 ,
		_w393_
	);
	LUT3 #(
		.INIT('hb0)
	) name195 (
		\n1312gat_reg/NET0131 ,
		\n1775gat_reg/NET0131 ,
		\n3100gat_pad ,
		_w394_
	);
	LUT3 #(
		.INIT('h80)
	) name196 (
		\n2510gat_reg/NET0131 ,
		\n2588gat_reg/NET0131 ,
		\n2658gat_reg/NET0131 ,
		_w395_
	);
	LUT2 #(
		.INIT('h8)
	) name197 (
		\n2502gat_reg/NET0131 ,
		\n2506gat_reg/NET0131 ,
		_w396_
	);
	LUT4 #(
		.INIT('hb000)
	) name198 (
		\n1312gat_reg/NET0131 ,
		\n1775gat_reg/NET0131 ,
		\n2502gat_reg/NET0131 ,
		\n2506gat_reg/NET0131 ,
		_w397_
	);
	LUT4 #(
		.INIT('h5444)
	) name199 (
		_w393_,
		_w394_,
		_w395_,
		_w397_,
		_w398_
	);
	LUT3 #(
		.INIT('hb0)
	) name200 (
		_w379_,
		_w392_,
		_w398_,
		_w399_
	);
	LUT4 #(
		.INIT('h7000)
	) name201 (
		_w369_,
		_w377_,
		_w386_,
		_w388_,
		_w400_
	);
	LUT3 #(
		.INIT('hb0)
	) name202 (
		_w379_,
		_w392_,
		_w400_,
		_w401_
	);
	LUT2 #(
		.INIT('h6)
	) name203 (
		\n2490gat_reg/NET0131 ,
		\n2634gat_reg/NET0131 ,
		_w402_
	);
	LUT2 #(
		.INIT('h2)
	) name204 (
		\n2622gat_reg/NET0131 ,
		\n2626gat_reg/NET0131 ,
		_w403_
	);
	LUT4 #(
		.INIT('h6996)
	) name205 (
		\n2543gat_reg/NET0131 ,
		\n2622gat_reg/NET0131 ,
		\n2626gat_reg/NET0131 ,
		\n2630gat_reg/NET0131 ,
		_w404_
	);
	LUT2 #(
		.INIT('h6)
	) name206 (
		_w402_,
		_w404_,
		_w405_
	);
	LUT2 #(
		.INIT('h9)
	) name207 (
		_w402_,
		_w404_,
		_w406_
	);
	LUT3 #(
		.INIT('h8c)
	) name208 (
		_w379_,
		_w384_,
		_w392_,
		_w407_
	);
	LUT3 #(
		.INIT('h40)
	) name209 (
		\n1740gat_reg/NET0131 ,
		_w386_,
		_w388_,
		_w408_
	);
	LUT2 #(
		.INIT('h1)
	) name210 (
		\n1496gat_reg/NET0131 ,
		\n2091gat_reg/NET0131 ,
		_w409_
	);
	LUT4 #(
		.INIT('h0080)
	) name211 (
		_w380_,
		_w382_,
		_w383_,
		_w409_,
		_w410_
	);
	LUT3 #(
		.INIT('h20)
	) name212 (
		\n1850gat_reg/NET0131 ,
		\n2061gat_reg/NET0131 ,
		\n2143gat_reg/NET0131 ,
		_w411_
	);
	LUT2 #(
		.INIT('h8)
	) name213 (
		_w387_,
		_w411_,
		_w412_
	);
	LUT4 #(
		.INIT('h8000)
	) name214 (
		_w380_,
		_w387_,
		_w409_,
		_w411_,
		_w413_
	);
	LUT4 #(
		.INIT('h0001)
	) name215 (
		\n1899gat_reg/NET0131 ,
		\n2061gat_reg/NET0131 ,
		\n2139gat_reg/NET0131 ,
		\n2143gat_reg/NET0131 ,
		_w414_
	);
	LUT2 #(
		.INIT('h8)
	) name216 (
		\n1850gat_reg/NET0131 ,
		_w414_,
		_w415_
	);
	LUT4 #(
		.INIT('h02aa)
	) name217 (
		\n1740gat_reg/NET0131 ,
		\n1763gat_reg/NET0131 ,
		\n1880gat_reg/NET0131 ,
		\n2102gat_reg/NET0131 ,
		_w416_
	);
	LUT3 #(
		.INIT('h80)
	) name218 (
		\n1850gat_reg/NET0131 ,
		_w414_,
		_w416_,
		_w417_
	);
	LUT4 #(
		.INIT('h0001)
	) name219 (
		_w408_,
		_w410_,
		_w413_,
		_w417_,
		_w418_
	);
	LUT3 #(
		.INIT('hc8)
	) name220 (
		_w369_,
		_w377_,
		_w380_,
		_w419_
	);
	LUT4 #(
		.INIT('h0001)
	) name221 (
		\n2135gat_reg/NET0131 ,
		\n2179gat_reg/NET0131 ,
		\n2190gat_reg/NET0131 ,
		\n2262gat_reg/NET0131 ,
		_w420_
	);
	LUT2 #(
		.INIT('h2)
	) name222 (
		\n2182gat_reg/NET0131 ,
		_w420_,
		_w421_
	);
	LUT2 #(
		.INIT('h4)
	) name223 (
		_w370_,
		_w380_,
		_w422_
	);
	LUT3 #(
		.INIT('h02)
	) name224 (
		_w419_,
		_w421_,
		_w422_,
		_w423_
	);
	LUT2 #(
		.INIT('h4)
	) name225 (
		_w418_,
		_w423_,
		_w424_
	);
	LUT3 #(
		.INIT('h80)
	) name226 (
		\n2490gat_reg/NET0131 ,
		\n2543gat_reg/NET0131 ,
		\n2630gat_reg/NET0131 ,
		_w425_
	);
	LUT2 #(
		.INIT('h8)
	) name227 (
		_w403_,
		_w425_,
		_w426_
	);
	LUT3 #(
		.INIT('h80)
	) name228 (
		\n2343gat_reg/NET0131 ,
		\n2399gat_reg/NET0131 ,
		\n2562gat_reg/NET0131 ,
		_w427_
	);
	LUT4 #(
		.INIT('h8000)
	) name229 (
		_w317_,
		_w403_,
		_w425_,
		_w427_,
		_w428_
	);
	LUT2 #(
		.INIT('h7)
	) name230 (
		_w395_,
		_w396_,
		_w429_
	);
	LUT3 #(
		.INIT('h15)
	) name231 (
		\n3100gat_pad ,
		_w395_,
		_w396_,
		_w430_
	);
	LUT3 #(
		.INIT('h56)
	) name232 (
		\n2135gat_reg/NET0131 ,
		\n2190gat_reg/NET0131 ,
		\n2262gat_reg/NET0131 ,
		_w431_
	);
	LUT3 #(
		.INIT('h70)
	) name233 (
		\n1880gat_reg/NET0131 ,
		\n2021gat_reg/NET0131 ,
		\n2099gat_reg/NET0131 ,
		_w432_
	);
	LUT2 #(
		.INIT('h8)
	) name234 (
		\n2037gat_reg/NET0131 ,
		\n2095gat_reg/NET0131 ,
		_w433_
	);
	LUT2 #(
		.INIT('h4)
	) name235 (
		_w432_,
		_w433_,
		_w434_
	);
	LUT3 #(
		.INIT('h20)
	) name236 (
		_w431_,
		_w432_,
		_w433_,
		_w435_
	);
	LUT2 #(
		.INIT('h4)
	) name237 (
		_w430_,
		_w435_,
		_w436_
	);
	LUT3 #(
		.INIT('h2d)
	) name238 (
		\n2190gat_reg/NET0131 ,
		\n2262gat_reg/NET0131 ,
		\n2266gat_reg/NET0131 ,
		_w437_
	);
	LUT3 #(
		.INIT('h40)
	) name239 (
		_w432_,
		_w433_,
		_w437_,
		_w438_
	);
	LUT2 #(
		.INIT('hb)
	) name240 (
		_w430_,
		_w438_,
		_w439_
	);
	LUT2 #(
		.INIT('h9)
	) name241 (
		\n684gat_reg/NET0131 ,
		\n816gat_reg/NET0131 ,
		_w440_
	);
	LUT4 #(
		.INIT('h9669)
	) name242 (
		\n680gat_reg/NET0131 ,
		\n699gat_reg/NET0131 ,
		\n824gat_reg/NET0131 ,
		\n883gat_reg/NET0131 ,
		_w441_
	);
	LUT3 #(
		.INIT('h96)
	) name243 (
		\n580gat_reg/NET0131 ,
		\n584gat_reg/NET0131 ,
		\n820gat_reg/NET0131 ,
		_w442_
	);
	LUT3 #(
		.INIT('h96)
	) name244 (
		_w440_,
		_w441_,
		_w442_,
		_w443_
	);
	LUT4 #(
		.INIT('h9669)
	) name245 (
		\n2270gat_reg/NET0131 ,
		\n2339gat_reg/NET0131 ,
		\n2390gat_reg/NET0131 ,
		\n2495gat_reg/NET0131 ,
		_w444_
	);
	LUT2 #(
		.INIT('h8)
	) name246 (
		\n2190gat_reg/NET0131 ,
		\n2262gat_reg/NET0131 ,
		_w445_
	);
	LUT3 #(
		.INIT('h04)
	) name247 (
		_w432_,
		_w433_,
		_w445_,
		_w446_
	);
	LUT2 #(
		.INIT('h4)
	) name248 (
		_w430_,
		_w446_,
		_w447_
	);
	LUT2 #(
		.INIT('h4)
	) name249 (
		_w430_,
		_w434_,
		_w448_
	);
	LUT2 #(
		.INIT('h8)
	) name250 (
		\n1899gat_reg/NET0131 ,
		\n2139gat_reg/NET0131 ,
		_w449_
	);
	LUT3 #(
		.INIT('h04)
	) name251 (
		_w430_,
		_w434_,
		_w449_,
		_w450_
	);
	LUT2 #(
		.INIT('h8)
	) name252 (
		_w418_,
		_w450_,
		_w451_
	);
	LUT4 #(
		.INIT('h01fe)
	) name253 (
		\n1899gat_reg/NET0131 ,
		\n2061gat_reg/NET0131 ,
		\n2139gat_reg/NET0131 ,
		\n2143gat_reg/NET0131 ,
		_w452_
	);
	LUT3 #(
		.INIT('h40)
	) name254 (
		_w430_,
		_w434_,
		_w452_,
		_w453_
	);
	LUT2 #(
		.INIT('h8)
	) name255 (
		_w418_,
		_w453_,
		_w454_
	);
	LUT3 #(
		.INIT('h04)
	) name256 (
		\n1899gat_reg/NET0131 ,
		\n2061gat_reg/NET0131 ,
		\n2139gat_reg/NET0131 ,
		_w455_
	);
	LUT3 #(
		.INIT('hc9)
	) name257 (
		\n1899gat_reg/NET0131 ,
		\n2061gat_reg/NET0131 ,
		\n2139gat_reg/NET0131 ,
		_w456_
	);
	LUT3 #(
		.INIT('h04)
	) name258 (
		_w430_,
		_w434_,
		_w456_,
		_w457_
	);
	LUT2 #(
		.INIT('h8)
	) name259 (
		_w418_,
		_w457_,
		_w458_
	);
	LUT2 #(
		.INIT('h6)
	) name260 (
		\n1850gat_reg/NET0131 ,
		_w414_,
		_w459_
	);
	LUT3 #(
		.INIT('h04)
	) name261 (
		_w430_,
		_w434_,
		_w459_,
		_w460_
	);
	LUT2 #(
		.INIT('h8)
	) name262 (
		_w418_,
		_w460_,
		_w461_
	);
	LUT4 #(
		.INIT('h5150)
	) name263 (
		\n1899gat_reg/NET0131 ,
		\n2061gat_reg/NET0131 ,
		\n2139gat_reg/NET0131 ,
		\n2143gat_reg/NET0131 ,
		_w462_
	);
	LUT2 #(
		.INIT('h6)
	) name264 (
		\n1975gat_reg/NET0131 ,
		_w462_,
		_w463_
	);
	LUT3 #(
		.INIT('h04)
	) name265 (
		_w430_,
		_w434_,
		_w463_,
		_w464_
	);
	LUT2 #(
		.INIT('h7)
	) name266 (
		_w418_,
		_w464_,
		_w465_
	);
	LUT4 #(
		.INIT('h9669)
	) name267 (
		\n398gat_reg/NET0131 ,
		\n402gat_reg/NET0131 ,
		\n846gat_reg/NET0131 ,
		\n919gat_reg/NET0131 ,
		_w466_
	);
	LUT2 #(
		.INIT('h6)
	) name268 (
		\n830gat_reg/NET0131 ,
		\n834gat_reg/NET0131 ,
		_w467_
	);
	LUT2 #(
		.INIT('h9)
	) name269 (
		\n614gat_reg/NET0131 ,
		\n838gat_reg/NET0131 ,
		_w468_
	);
	LUT4 #(
		.INIT('h6996)
	) name270 (
		\n707gat_reg/NET0131 ,
		_w466_,
		_w467_,
		_w468_,
		_w469_
	);
	LUT4 #(
		.INIT('h2040)
	) name271 (
		\n2394gat_reg/NET0131 ,
		\n2440gat_reg/NET0131 ,
		_w377_,
		_w380_,
		_w470_
	);
	LUT3 #(
		.INIT('h04)
	) name272 (
		_w430_,
		_w434_,
		_w470_,
		_w471_
	);
	LUT4 #(
		.INIT('h5554)
	) name273 (
		\n2347gat_reg/NET0131 ,
		\n2394gat_reg/NET0131 ,
		\n2403gat_reg/NET0131 ,
		\n2440gat_reg/NET0131 ,
		_w472_
	);
	LUT4 #(
		.INIT('h0002)
	) name274 (
		\n2347gat_reg/NET0131 ,
		\n2394gat_reg/NET0131 ,
		\n2403gat_reg/NET0131 ,
		\n2440gat_reg/NET0131 ,
		_w473_
	);
	LUT4 #(
		.INIT('haaa9)
	) name275 (
		\n2347gat_reg/NET0131 ,
		\n2394gat_reg/NET0131 ,
		\n2403gat_reg/NET0131 ,
		\n2440gat_reg/NET0131 ,
		_w474_
	);
	LUT4 #(
		.INIT('h0004)
	) name276 (
		_w430_,
		_w434_,
		_w470_,
		_w474_,
		_w475_
	);
	LUT4 #(
		.INIT('h1e0f)
	) name277 (
		\n2347gat_reg/NET0131 ,
		\n2403gat_reg/NET0131 ,
		\n2407gat_reg/NET0131 ,
		_w366_,
		_w476_
	);
	LUT4 #(
		.INIT('h0400)
	) name278 (
		_w430_,
		_w434_,
		_w470_,
		_w476_,
		_w477_
	);
	LUT3 #(
		.INIT('h02)
	) name279 (
		\n2394gat_reg/NET0131 ,
		\n2440gat_reg/NET0131 ,
		\n2644gat_reg/NET0131 ,
		_w478_
	);
	LUT4 #(
		.INIT('h0002)
	) name280 (
		\n2347gat_reg/NET0131 ,
		\n2403gat_reg/NET0131 ,
		\n2440gat_reg/NET0131 ,
		\n2644gat_reg/NET0131 ,
		_w479_
	);
	LUT2 #(
		.INIT('h1)
	) name281 (
		_w478_,
		_w479_,
		_w480_
	);
	LUT3 #(
		.INIT('h02)
	) name282 (
		\n2347gat_reg/NET0131 ,
		\n2403gat_reg/NET0131 ,
		\n2440gat_reg/NET0131 ,
		_w481_
	);
	LUT3 #(
		.INIT('hd0)
	) name283 (
		\n2394gat_reg/NET0131 ,
		\n2440gat_reg/NET0131 ,
		\n2644gat_reg/NET0131 ,
		_w482_
	);
	LUT4 #(
		.INIT('h4044)
	) name284 (
		_w432_,
		_w433_,
		_w481_,
		_w482_,
		_w483_
	);
	LUT4 #(
		.INIT('hefff)
	) name285 (
		_w430_,
		_w470_,
		_w480_,
		_w483_,
		_w484_
	);
	LUT3 #(
		.INIT('h36)
	) name286 (
		\n2394gat_reg/NET0131 ,
		\n2403gat_reg/NET0131 ,
		\n2440gat_reg/NET0131 ,
		_w485_
	);
	LUT3 #(
		.INIT('h40)
	) name287 (
		_w432_,
		_w433_,
		_w485_,
		_w486_
	);
	LUT3 #(
		.INIT('h10)
	) name288 (
		_w430_,
		_w470_,
		_w486_,
		_w487_
	);
	LUT4 #(
		.INIT('ha8c8)
	) name289 (
		\n2394gat_reg/NET0131 ,
		\n2440gat_reg/NET0131 ,
		_w377_,
		_w380_,
		_w488_
	);
	LUT3 #(
		.INIT('h04)
	) name290 (
		_w430_,
		_w434_,
		_w488_,
		_w489_
	);
	LUT3 #(
		.INIT('h10)
	) name291 (
		\n2347gat_reg/NET0131 ,
		\n2403gat_reg/NET0131 ,
		\n2407gat_reg/NET0131 ,
		_w490_
	);
	LUT2 #(
		.INIT('h8)
	) name292 (
		_w369_,
		_w490_,
		_w491_
	);
	LUT3 #(
		.INIT('he0)
	) name293 (
		_w385_,
		_w389_,
		_w491_,
		_w492_
	);
	LUT2 #(
		.INIT('h2)
	) name294 (
		\n1850gat_reg/NET0131 ,
		\n2143gat_reg/NET0131 ,
		_w493_
	);
	LUT3 #(
		.INIT('h40)
	) name295 (
		\n1899gat_reg/NET0131 ,
		\n2061gat_reg/NET0131 ,
		\n2139gat_reg/NET0131 ,
		_w494_
	);
	LUT3 #(
		.INIT('h40)
	) name296 (
		_w380_,
		_w493_,
		_w494_,
		_w495_
	);
	LUT4 #(
		.INIT('h0040)
	) name297 (
		\n2454gat_reg/NET0131 ,
		\n398gat_reg/NET0131 ,
		\n402gat_reg/NET0131 ,
		\n846gat_reg/NET0131 ,
		_w496_
	);
	LUT2 #(
		.INIT('hd)
	) name298 (
		_w314_,
		_w496_,
		_w497_
	);
	LUT3 #(
		.INIT('h01)
	) name299 (
		\n1316gat_reg/NET0131 ,
		\n1775gat_reg/NET0131 ,
		\n2040gat_reg/NET0131 ,
		_w498_
	);
	LUT2 #(
		.INIT('h9)
	) name300 (
		\n1241gat_reg/NET0131 ,
		\n957gat_reg/NET0131 ,
		_w499_
	);
	LUT4 #(
		.INIT('h9669)
	) name301 (
		\n1068gat_reg/NET0131 ,
		\n1294gat_reg/NET0131 ,
		\n673gat_reg/NET0131 ,
		\n861gat_reg/NET0131 ,
		_w500_
	);
	LUT3 #(
		.INIT('h96)
	) name302 (
		\n1080gat_reg/NET0131 ,
		\n1148gat_reg/NET0131 ,
		\n865gat_reg/NET0131 ,
		_w501_
	);
	LUT3 #(
		.INIT('h96)
	) name303 (
		_w499_,
		_w500_,
		_w501_,
		_w502_
	);
	LUT3 #(
		.INIT('h04)
	) name304 (
		\n2454gat_reg/NET0131 ,
		\n398gat_reg/NET0131 ,
		\n402gat_reg/NET0131 ,
		_w503_
	);
	LUT2 #(
		.INIT('h8)
	) name305 (
		_w368_,
		_w503_,
		_w504_
	);
	LUT2 #(
		.INIT('h7)
	) name306 (
		\n2446gat_reg/NET0131 ,
		\n2450gat_reg/NET0131 ,
		_w505_
	);
	LUT3 #(
		.INIT('h07)
	) name307 (
		\n2446gat_reg/NET0131 ,
		\n2450gat_reg/NET0131 ,
		\n3100gat_pad ,
		_w506_
	);
	LUT3 #(
		.INIT('hd0)
	) name308 (
		\n1821gat_reg/NET0131 ,
		\n1829gat_reg/NET0131 ,
		\n2472gat_reg/NET0131 ,
		_w507_
	);
	LUT4 #(
		.INIT('h0800)
	) name309 (
		_w368_,
		_w503_,
		_w506_,
		_w507_,
		_w508_
	);
	LUT2 #(
		.INIT('h1)
	) name310 (
		\n2454gat_reg/NET0131 ,
		\n271gat_reg/NET0131 ,
		_w509_
	);
	LUT3 #(
		.INIT('h40)
	) name311 (
		_w506_,
		_w507_,
		_w509_,
		_w510_
	);
	LUT2 #(
		.INIT('h8)
	) name312 (
		_w367_,
		_w503_,
		_w511_
	);
	LUT4 #(
		.INIT('h0800)
	) name313 (
		_w367_,
		_w503_,
		_w506_,
		_w507_,
		_w512_
	);
	LUT4 #(
		.INIT('h0010)
	) name314 (
		\n2454gat_reg/NET0131 ,
		\n388gat_reg/NET0131 ,
		\n398gat_reg/NET0131 ,
		\n402gat_reg/NET0131 ,
		_w513_
	);
	LUT3 #(
		.INIT('h2a)
	) name315 (
		\n331gat_reg/NET0131 ,
		_w373_,
		_w513_,
		_w514_
	);
	LUT3 #(
		.INIT('h2a)
	) name316 (
		\n3094gat_pad ,
		_w254_,
		_w337_,
		_w515_
	);
	LUT3 #(
		.INIT('h80)
	) name317 (
		\n3086gat_pad ,
		\n3088gat_pad ,
		\n3095gat_pad ,
		_w516_
	);
	LUT4 #(
		.INIT('h2000)
	) name318 (
		\n3094gat_pad ,
		_w254_,
		_w337_,
		_w516_,
		_w517_
	);
	LUT4 #(
		.INIT('h2220)
	) name319 (
		\n3085gat_pad ,
		\n3086gat_pad ,
		\n3091gat_pad ,
		\n3092gat_pad ,
		_w518_
	);
	LUT4 #(
		.INIT('h2000)
	) name320 (
		\n3087gat_pad ,
		\n3088gat_pad ,
		_w341_,
		_w518_,
		_w519_
	);
	LUT4 #(
		.INIT('h1000)
	) name321 (
		\n331gat_reg/NET0131 ,
		\n388gat_reg/NET0131 ,
		\n846gat_reg/NET0131 ,
		\n919gat_reg/NET0131 ,
		_w520_
	);
	LUT2 #(
		.INIT('h8)
	) name322 (
		_w503_,
		_w520_,
		_w521_
	);
	LUT4 #(
		.INIT('h0001)
	) name323 (
		_w514_,
		_w517_,
		_w519_,
		_w521_,
		_w522_
	);
	LUT3 #(
		.INIT('h80)
	) name324 (
		\n3080gat_pad ,
		_w337_,
		_w516_,
		_w523_
	);
	LUT2 #(
		.INIT('h2)
	) name325 (
		\n3071gat_pad ,
		\n3088gat_pad ,
		_w524_
	);
	LUT4 #(
		.INIT('h8000)
	) name326 (
		\n3087gat_pad ,
		_w341_,
		_w518_,
		_w524_,
		_w525_
	);
	LUT3 #(
		.INIT('h07)
	) name327 (
		_w515_,
		_w523_,
		_w525_,
		_w526_
	);
	LUT2 #(
		.INIT('hb)
	) name328 (
		_w522_,
		_w526_,
		_w527_
	);
	LUT2 #(
		.INIT('h8)
	) name329 (
		\n3087gat_pad ,
		\n3088gat_pad ,
		_w528_
	);
	LUT3 #(
		.INIT('h80)
	) name330 (
		_w341_,
		_w518_,
		_w528_,
		_w529_
	);
	LUT4 #(
		.INIT('h8000)
	) name331 (
		\n3065gat_pad ,
		_w341_,
		_w518_,
		_w528_,
		_w530_
	);
	LUT3 #(
		.INIT('h80)
	) name332 (
		\n3065gat_pad ,
		_w337_,
		_w516_,
		_w531_
	);
	LUT3 #(
		.INIT('h13)
	) name333 (
		_w515_,
		_w530_,
		_w531_,
		_w532_
	);
	LUT4 #(
		.INIT('h0010)
	) name334 (
		\n152gat_reg/NET0131 ,
		\n156gat_reg/NET0131 ,
		\n398gat_reg/NET0131 ,
		\n402gat_reg/NET0131 ,
		_w533_
	);
	LUT4 #(
		.INIT('h0010)
	) name335 (
		\n2454gat_reg/NET0131 ,
		\n256gat_reg/NET0131 ,
		\n846gat_reg/NET0131 ,
		\n919gat_reg/NET0131 ,
		_w534_
	);
	LUT3 #(
		.INIT('h6a)
	) name336 (
		\n148gat_reg/NET0131 ,
		_w533_,
		_w534_,
		_w535_
	);
	LUT3 #(
		.INIT('h01)
	) name337 (
		_w517_,
		_w529_,
		_w535_,
		_w536_
	);
	LUT2 #(
		.INIT('hd)
	) name338 (
		_w532_,
		_w536_,
		_w537_
	);
	LUT3 #(
		.INIT('h23)
	) name339 (
		\n152gat_reg/NET0131 ,
		\n156gat_reg/NET0131 ,
		\n256gat_reg/NET0131 ,
		_w538_
	);
	LUT4 #(
		.INIT('haa6a)
	) name340 (
		\n470gat_reg/NET0131 ,
		_w247_,
		_w312_,
		_w538_,
		_w539_
	);
	LUT3 #(
		.INIT('h01)
	) name341 (
		_w517_,
		_w529_,
		_w539_,
		_w540_
	);
	LUT4 #(
		.INIT('h8000)
	) name342 (
		\n3073gat_pad ,
		_w341_,
		_w518_,
		_w528_,
		_w541_
	);
	LUT3 #(
		.INIT('h80)
	) name343 (
		\n3073gat_pad ,
		_w337_,
		_w516_,
		_w542_
	);
	LUT3 #(
		.INIT('h13)
	) name344 (
		_w515_,
		_w541_,
		_w542_,
		_w543_
	);
	LUT2 #(
		.INIT('hb)
	) name345 (
		_w540_,
		_w543_,
		_w544_
	);
	LUT3 #(
		.INIT('h96)
	) name346 (
		\n3084gat_pad ,
		\n3085gat_pad ,
		\n3089gat_pad ,
		_w545_
	);
	LUT2 #(
		.INIT('h6)
	) name347 (
		\n3083gat_pad ,
		\n3088gat_pad ,
		_w546_
	);
	LUT2 #(
		.INIT('h6)
	) name348 (
		\n3086gat_pad ,
		\n3087gat_pad ,
		_w547_
	);
	LUT3 #(
		.INIT('h69)
	) name349 (
		_w545_,
		_w546_,
		_w547_,
		_w548_
	);
	LUT2 #(
		.INIT('h8)
	) name350 (
		_w312_,
		_w533_,
		_w549_
	);
	LUT4 #(
		.INIT('h6555)
	) name351 (
		\n256gat_reg/NET0131 ,
		\n919gat_reg/NET0131 ,
		_w248_,
		_w533_,
		_w550_
	);
	LUT3 #(
		.INIT('h10)
	) name352 (
		_w517_,
		_w529_,
		_w550_,
		_w551_
	);
	LUT4 #(
		.INIT('h8000)
	) name353 (
		\n3066gat_pad ,
		_w341_,
		_w518_,
		_w528_,
		_w552_
	);
	LUT3 #(
		.INIT('h80)
	) name354 (
		\n3066gat_pad ,
		_w337_,
		_w516_,
		_w553_
	);
	LUT3 #(
		.INIT('h13)
	) name355 (
		_w515_,
		_w552_,
		_w553_,
		_w554_
	);
	LUT2 #(
		.INIT('hb)
	) name356 (
		_w551_,
		_w554_,
		_w555_
	);
	LUT4 #(
		.INIT('h0010)
	) name357 (
		\n2454gat_reg/NET0131 ,
		\n327gat_reg/NET0131 ,
		\n398gat_reg/NET0131 ,
		\n402gat_reg/NET0131 ,
		_w556_
	);
	LUT4 #(
		.INIT('h6333)
	) name358 (
		\n2454gat_reg/NET0131 ,
		\n327gat_reg/NET0131 ,
		_w247_,
		_w520_,
		_w557_
	);
	LUT3 #(
		.INIT('h10)
	) name359 (
		_w517_,
		_w519_,
		_w557_,
		_w558_
	);
	LUT3 #(
		.INIT('h80)
	) name360 (
		\n3079gat_pad ,
		_w337_,
		_w516_,
		_w559_
	);
	LUT2 #(
		.INIT('h8)
	) name361 (
		\n3070gat_pad ,
		\n3087gat_pad ,
		_w560_
	);
	LUT4 #(
		.INIT('h4000)
	) name362 (
		\n3088gat_pad ,
		_w341_,
		_w518_,
		_w560_,
		_w561_
	);
	LUT3 #(
		.INIT('h07)
	) name363 (
		_w515_,
		_w559_,
		_w561_,
		_w562_
	);
	LUT2 #(
		.INIT('hb)
	) name364 (
		_w558_,
		_w562_,
		_w563_
	);
	LUT3 #(
		.INIT('h04)
	) name365 (
		\n156gat_reg/NET0131 ,
		\n398gat_reg/NET0131 ,
		\n402gat_reg/NET0131 ,
		_w564_
	);
	LUT3 #(
		.INIT('h2a)
	) name366 (
		\n152gat_reg/NET0131 ,
		_w312_,
		_w564_,
		_w565_
	);
	LUT4 #(
		.INIT('h0001)
	) name367 (
		_w517_,
		_w529_,
		_w549_,
		_w565_,
		_w566_
	);
	LUT4 #(
		.INIT('h8000)
	) name368 (
		\n3067gat_pad ,
		_w341_,
		_w518_,
		_w528_,
		_w567_
	);
	LUT3 #(
		.INIT('h80)
	) name369 (
		\n3067gat_pad ,
		_w337_,
		_w516_,
		_w568_
	);
	LUT3 #(
		.INIT('h13)
	) name370 (
		_w515_,
		_w567_,
		_w568_,
		_w569_
	);
	LUT2 #(
		.INIT('hb)
	) name371 (
		_w566_,
		_w569_,
		_w570_
	);
	LUT3 #(
		.INIT('h40)
	) name372 (
		\n398gat_reg/NET0131 ,
		\n402gat_reg/NET0131 ,
		\n919gat_reg/NET0131 ,
		_w571_
	);
	LUT3 #(
		.INIT('h13)
	) name373 (
		_w248_,
		_w496_,
		_w571_,
		_w572_
	);
	LUT3 #(
		.INIT('h07)
	) name374 (
		_w311_,
		_w312_,
		_w503_,
		_w573_
	);
	LUT2 #(
		.INIT('h7)
	) name375 (
		_w572_,
		_w573_,
		_w574_
	);
	LUT3 #(
		.INIT('h95)
	) name376 (
		\n156gat_reg/NET0131 ,
		_w247_,
		_w312_,
		_w575_
	);
	LUT3 #(
		.INIT('h10)
	) name377 (
		_w517_,
		_w529_,
		_w575_,
		_w576_
	);
	LUT4 #(
		.INIT('h8000)
	) name378 (
		\n3068gat_pad ,
		_w341_,
		_w518_,
		_w528_,
		_w577_
	);
	LUT3 #(
		.INIT('h80)
	) name379 (
		\n3068gat_pad ,
		_w337_,
		_w516_,
		_w578_
	);
	LUT3 #(
		.INIT('h13)
	) name380 (
		_w515_,
		_w577_,
		_w578_,
		_w579_
	);
	LUT2 #(
		.INIT('hb)
	) name381 (
		_w576_,
		_w579_,
		_w580_
	);
	LUT2 #(
		.INIT('h8)
	) name382 (
		\n3067gat_pad ,
		\n3087gat_pad ,
		_w581_
	);
	LUT4 #(
		.INIT('h4000)
	) name383 (
		\n3088gat_pad ,
		_w341_,
		_w518_,
		_w581_,
		_w582_
	);
	LUT3 #(
		.INIT('h80)
	) name384 (
		\n3076gat_pad ,
		_w337_,
		_w516_,
		_w583_
	);
	LUT3 #(
		.INIT('hec)
	) name385 (
		_w515_,
		_w582_,
		_w583_,
		_w584_
	);
	LUT2 #(
		.INIT('h8)
	) name386 (
		\n3068gat_pad ,
		\n3087gat_pad ,
		_w585_
	);
	LUT4 #(
		.INIT('h4000)
	) name387 (
		\n3088gat_pad ,
		_w341_,
		_w518_,
		_w585_,
		_w586_
	);
	LUT3 #(
		.INIT('h80)
	) name388 (
		\n3077gat_pad ,
		_w337_,
		_w516_,
		_w587_
	);
	LUT3 #(
		.INIT('hec)
	) name389 (
		_w515_,
		_w586_,
		_w587_,
		_w588_
	);
	LUT2 #(
		.INIT('h8)
	) name390 (
		\n3065gat_pad ,
		\n3087gat_pad ,
		_w589_
	);
	LUT4 #(
		.INIT('h4000)
	) name391 (
		\n3088gat_pad ,
		_w341_,
		_w518_,
		_w589_,
		_w590_
	);
	LUT3 #(
		.INIT('h80)
	) name392 (
		\n3074gat_pad ,
		_w337_,
		_w516_,
		_w591_
	);
	LUT3 #(
		.INIT('hec)
	) name393 (
		_w515_,
		_w590_,
		_w591_,
		_w592_
	);
	LUT2 #(
		.INIT('h8)
	) name394 (
		\n3066gat_pad ,
		\n3087gat_pad ,
		_w593_
	);
	LUT4 #(
		.INIT('h4000)
	) name395 (
		\n3088gat_pad ,
		_w341_,
		_w518_,
		_w593_,
		_w594_
	);
	LUT3 #(
		.INIT('h80)
	) name396 (
		\n3075gat_pad ,
		_w337_,
		_w516_,
		_w595_
	);
	LUT3 #(
		.INIT('hec)
	) name397 (
		_w515_,
		_w594_,
		_w595_,
		_w596_
	);
	LUT2 #(
		.INIT('h8)
	) name398 (
		\n2203gat_reg/NET0131 ,
		\n2207gat_reg/NET0131 ,
		_w597_
	);
	LUT2 #(
		.INIT('h6)
	) name399 (
		\n2203gat_reg/NET0131 ,
		\n2207gat_reg/NET0131 ,
		_w598_
	);
	LUT4 #(
		.INIT('h9669)
	) name400 (
		\n2343gat_reg/NET0131 ,
		\n2399gat_reg/NET0131 ,
		\n2562gat_reg/NET0131 ,
		\n2640gat_reg/NET0131 ,
		_w599_
	);
	LUT2 #(
		.INIT('h6)
	) name401 (
		_w598_,
		_w599_,
		_w600_
	);
	LUT2 #(
		.INIT('h2)
	) name402 (
		\n2117gat_reg/NET0131 ,
		\n2125gat_reg/NET0131 ,
		_w601_
	);
	LUT2 #(
		.INIT('h4)
	) name403 (
		_w506_,
		_w601_,
		_w602_
	);
	LUT3 #(
		.INIT('h80)
	) name404 (
		_w337_,
		_w338_,
		_w516_,
		_w603_
	);
	LUT2 #(
		.INIT('h2)
	) name405 (
		\n3087gat_pad ,
		\n3088gat_pad ,
		_w604_
	);
	LUT3 #(
		.INIT('h80)
	) name406 (
		_w341_,
		_w344_,
		_w604_,
		_w605_
	);
	LUT2 #(
		.INIT('he)
	) name407 (
		_w603_,
		_w605_,
		_w606_
	);
	LUT2 #(
		.INIT('h2)
	) name408 (
		\n2319gat_reg/NET0131 ,
		\n3099gat_pad ,
		_w607_
	);
	LUT2 #(
		.INIT('hb)
	) name409 (
		_w313_,
		_w572_,
		_w608_
	);
	LUT4 #(
		.INIT('h8000)
	) name410 (
		\n1850gat_reg/NET0131 ,
		_w370_,
		_w414_,
		_w490_,
		_w609_
	);
	LUT3 #(
		.INIT('h80)
	) name411 (
		\n2394gat_reg/NET0131 ,
		\n2403gat_reg/NET0131 ,
		\n2440gat_reg/NET0131 ,
		_w610_
	);
	LUT3 #(
		.INIT('h80)
	) name412 (
		\n1850gat_reg/NET0131 ,
		\n2061gat_reg/NET0131 ,
		\n2143gat_reg/NET0131 ,
		_w611_
	);
	LUT4 #(
		.INIT('h0040)
	) name413 (
		\n1899gat_reg/NET0131 ,
		\n2139gat_reg/NET0131 ,
		\n2347gat_reg/NET0131 ,
		\n2407gat_reg/NET0131 ,
		_w612_
	);
	LUT3 #(
		.INIT('h80)
	) name414 (
		_w610_,
		_w611_,
		_w612_,
		_w613_
	);
	LUT4 #(
		.INIT('h8000)
	) name415 (
		_w370_,
		_w382_,
		_w383_,
		_w490_,
		_w614_
	);
	LUT2 #(
		.INIT('h8)
	) name416 (
		_w411_,
		_w449_,
		_w615_
	);
	LUT4 #(
		.INIT('h8000)
	) name417 (
		_w369_,
		_w411_,
		_w449_,
		_w490_,
		_w616_
	);
	LUT4 #(
		.INIT('h8000)
	) name418 (
		_w369_,
		_w382_,
		_w455_,
		_w490_,
		_w617_
	);
	LUT3 #(
		.INIT('h20)
	) name419 (
		\n1312gat_reg/NET0131 ,
		\n1899gat_reg/NET0131 ,
		\n2139gat_reg/NET0131 ,
		_w618_
	);
	LUT2 #(
		.INIT('h8)
	) name420 (
		_w611_,
		_w618_,
		_w619_
	);
	LUT2 #(
		.INIT('h2)
	) name421 (
		\n1899gat_reg/NET0131 ,
		\n2139gat_reg/NET0131 ,
		_w620_
	);
	LUT2 #(
		.INIT('h8)
	) name422 (
		_w611_,
		_w620_,
		_w621_
	);
	LUT4 #(
		.INIT('h8000)
	) name423 (
		\n398gat_reg/NET0131 ,
		\n402gat_reg/NET0131 ,
		\n846gat_reg/NET0131 ,
		\n919gat_reg/NET0131 ,
		_w622_
	);
	LUT4 #(
		.INIT('h135f)
	) name424 (
		\n3066gat_pad ,
		\n3075gat_pad ,
		\n3093gat_pad ,
		\n3095gat_pad ,
		_w623_
	);
	LUT4 #(
		.INIT('heca0)
	) name425 (
		\n3066gat_pad ,
		\n3075gat_pad ,
		\n3093gat_pad ,
		\n3095gat_pad ,
		_w624_
	);
	LUT4 #(
		.INIT('h135f)
	) name426 (
		\n3068gat_pad ,
		\n3077gat_pad ,
		\n3093gat_pad ,
		\n3095gat_pad ,
		_w625_
	);
	LUT4 #(
		.INIT('heca0)
	) name427 (
		\n3068gat_pad ,
		\n3077gat_pad ,
		\n3093gat_pad ,
		\n3095gat_pad ,
		_w626_
	);
	LUT4 #(
		.INIT('h135f)
	) name428 (
		\n3067gat_pad ,
		\n3076gat_pad ,
		\n3093gat_pad ,
		\n3095gat_pad ,
		_w627_
	);
	LUT4 #(
		.INIT('heca0)
	) name429 (
		\n3067gat_pad ,
		\n3076gat_pad ,
		\n3093gat_pad ,
		\n3095gat_pad ,
		_w628_
	);
	LUT2 #(
		.INIT('h6)
	) name430 (
		\n271gat_reg/NET0131 ,
		\n842gat_reg/NET0131 ,
		_w629_
	);
	LUT2 #(
		.INIT('h9)
	) name431 (
		\n337gat_reg/NET0131 ,
		\n341gat_reg/NET0131 ,
		_w630_
	);
	LUT4 #(
		.INIT('h6996)
	) name432 (
		\n160gat_reg/NET0131 ,
		_w466_,
		_w629_,
		_w630_,
		_w631_
	);
	LUT2 #(
		.INIT('hb)
	) name433 (
		_w320_,
		_w627_,
		_w632_
	);
	LUT2 #(
		.INIT('hb)
	) name434 (
		_w320_,
		_w625_,
		_w633_
	);
	LUT3 #(
		.INIT('h2a)
	) name435 (
		\n384gat_reg/NET0131 ,
		_w520_,
		_w556_,
		_w634_
	);
	LUT2 #(
		.INIT('h1)
	) name436 (
		\n327gat_reg/NET0131 ,
		\n384gat_reg/NET0131 ,
		_w635_
	);
	LUT3 #(
		.INIT('h80)
	) name437 (
		_w503_,
		_w520_,
		_w635_,
		_w636_
	);
	LUT4 #(
		.INIT('h0001)
	) name438 (
		_w517_,
		_w519_,
		_w634_,
		_w636_,
		_w637_
	);
	LUT3 #(
		.INIT('h80)
	) name439 (
		\n3078gat_pad ,
		_w337_,
		_w516_,
		_w638_
	);
	LUT2 #(
		.INIT('h8)
	) name440 (
		\n3069gat_pad ,
		\n3087gat_pad ,
		_w639_
	);
	LUT4 #(
		.INIT('h4000)
	) name441 (
		\n3088gat_pad ,
		_w341_,
		_w518_,
		_w639_,
		_w640_
	);
	LUT3 #(
		.INIT('h07)
	) name442 (
		_w515_,
		_w638_,
		_w640_,
		_w641_
	);
	LUT2 #(
		.INIT('hb)
	) name443 (
		_w637_,
		_w641_,
		_w642_
	);
	LUT2 #(
		.INIT('h8)
	) name444 (
		_w418_,
		_w448_,
		_w643_
	);
	LUT3 #(
		.INIT('h0d)
	) name445 (
		\n327gat_reg/NET0131 ,
		\n331gat_reg/NET0131 ,
		\n388gat_reg/NET0131 ,
		_w644_
	);
	LUT4 #(
		.INIT('haa6a)
	) name446 (
		\n463gat_reg/NET0131 ,
		_w373_,
		_w503_,
		_w644_,
		_w645_
	);
	LUT3 #(
		.INIT('h01)
	) name447 (
		_w517_,
		_w519_,
		_w645_,
		_w646_
	);
	LUT3 #(
		.INIT('h80)
	) name448 (
		\n3082gat_pad ,
		_w337_,
		_w516_,
		_w647_
	);
	LUT2 #(
		.INIT('h8)
	) name449 (
		\n3073gat_pad ,
		\n3087gat_pad ,
		_w648_
	);
	LUT4 #(
		.INIT('h4000)
	) name450 (
		\n3088gat_pad ,
		_w341_,
		_w518_,
		_w648_,
		_w649_
	);
	LUT3 #(
		.INIT('h07)
	) name451 (
		_w515_,
		_w647_,
		_w649_,
		_w650_
	);
	LUT2 #(
		.INIT('hb)
	) name452 (
		_w646_,
		_w650_,
		_w651_
	);
	LUT2 #(
		.INIT('hb)
	) name453 (
		_w320_,
		_w623_,
		_w652_
	);
	LUT4 #(
		.INIT('h6333)
	) name454 (
		\n2454gat_reg/NET0131 ,
		\n388gat_reg/NET0131 ,
		_w247_,
		_w373_,
		_w653_
	);
	LUT3 #(
		.INIT('h10)
	) name455 (
		_w517_,
		_w519_,
		_w653_,
		_w654_
	);
	LUT3 #(
		.INIT('h80)
	) name456 (
		\n3081gat_pad ,
		_w337_,
		_w516_,
		_w655_
	);
	LUT2 #(
		.INIT('h8)
	) name457 (
		\n3072gat_pad ,
		\n3087gat_pad ,
		_w656_
	);
	LUT4 #(
		.INIT('h4000)
	) name458 (
		\n3088gat_pad ,
		_w341_,
		_w518_,
		_w656_,
		_w657_
	);
	LUT3 #(
		.INIT('h07)
	) name459 (
		_w515_,
		_w655_,
		_w657_,
		_w658_
	);
	LUT2 #(
		.INIT('hb)
	) name460 (
		_w654_,
		_w658_,
		_w659_
	);
	LUT3 #(
		.INIT('h0b)
	) name461 (
		_w379_,
		_w392_,
		_w393_,
		_w660_
	);
	LUT3 #(
		.INIT('h20)
	) name462 (
		\n1312gat_reg/NET0131 ,
		\n2169gat_reg/NET0131 ,
		\n3100gat_pad ,
		_w661_
	);
	LUT4 #(
		.INIT('h2000)
	) name463 (
		\n1312gat_reg/NET0131 ,
		\n2169gat_reg/NET0131 ,
		\n2502gat_reg/NET0131 ,
		\n2506gat_reg/NET0131 ,
		_w662_
	);
	LUT3 #(
		.INIT('h13)
	) name464 (
		_w395_,
		_w661_,
		_w662_,
		_w663_
	);
	LUT3 #(
		.INIT('h0b)
	) name465 (
		_w379_,
		_w392_,
		_w663_,
		_w664_
	);
	LUT4 #(
		.INIT('h6996)
	) name466 (
		\n1197gat_reg/NET0131 ,
		_w276_,
		_w277_,
		_w278_,
		_w665_
	);
	LUT4 #(
		.INIT('h9669)
	) name467 (
		\n1197gat_reg/NET0131 ,
		_w276_,
		_w277_,
		_w278_,
		_w666_
	);
	LUT4 #(
		.INIT('h0400)
	) name468 (
		\n3085gat_pad ,
		\n3086gat_pad ,
		\n3087gat_pad ,
		\n3088gat_pad ,
		_w667_
	);
	LUT3 #(
		.INIT('h20)
	) name469 (
		_w341_,
		_w343_,
		_w667_,
		_w668_
	);
	LUT3 #(
		.INIT('h15)
	) name470 (
		\n3086gat_pad ,
		\n3088gat_pad ,
		\n3095gat_pad ,
		_w669_
	);
	LUT3 #(
		.INIT('h80)
	) name471 (
		_w337_,
		_w338_,
		_w669_,
		_w670_
	);
	LUT3 #(
		.INIT('hfd)
	) name472 (
		_w459_,
		_w668_,
		_w670_,
		_w671_
	);
	LUT4 #(
		.INIT('h2000)
	) name473 (
		\n3094gat_pad ,
		_w254_,
		_w337_,
		_w339_,
		_w672_
	);
	LUT4 #(
		.INIT('h070f)
	) name474 (
		_w341_,
		_w342_,
		_w452_,
		_w518_,
		_w673_
	);
	LUT2 #(
		.INIT('hb)
	) name475 (
		_w672_,
		_w673_,
		_w674_
	);
	LUT3 #(
		.INIT('h70)
	) name476 (
		\n1771gat_reg/NET0131 ,
		\n1775gat_reg/NET0131 ,
		\n1871gat_reg/NET0131 ,
		_w675_
	);
	LUT2 #(
		.INIT('hd)
	) name477 (
		\n1035gat_reg/NET0131 ,
		_w476_,
		_w676_
	);
	LUT3 #(
		.INIT('hfd)
	) name478 (
		\n1072gat_reg/NET0131 ,
		_w472_,
		_w473_,
		_w677_
	);
	LUT4 #(
		.INIT('h5f7d)
	) name479 (
		\n1121gat_reg/NET0131 ,
		\n2394gat_reg/NET0131 ,
		\n2403gat_reg/NET0131 ,
		\n2440gat_reg/NET0131 ,
		_w678_
	);
	LUT3 #(
		.INIT('h7f)
	) name480 (
		\n2394gat_reg/NET0131 ,
		\n2440gat_reg/NET0131 ,
		\n931gat_reg/NET0131 ,
		_w679_
	);
	LUT4 #(
		.INIT('h777d)
	) name481 (
		\n1135gat_reg/NET0131 ,
		\n2135gat_reg/NET0131 ,
		\n2190gat_reg/NET0131 ,
		\n2262gat_reg/NET0131 ,
		_w680_
	);
	LUT3 #(
		.INIT('h7f)
	) name482 (
		\n1282gat_reg/NET0131 ,
		\n2190gat_reg/NET0131 ,
		\n2262gat_reg/NET0131 ,
		_w681_
	);
	LUT3 #(
		.INIT('h96)
	) name483 (
		_w276_,
		_w277_,
		_w278_,
		_w682_
	);
	LUT4 #(
		.INIT('h0004)
	) name484 (
		\n659gat_reg/NET0131 ,
		_w253_,
		_w255_,
		_w256_,
		_w683_
	);
	LUT4 #(
		.INIT('h0100)
	) name485 (
		\n1068gat_reg/NET0131 ,
		_w253_,
		_w255_,
		_w256_,
		_w684_
	);
	LUT4 #(
		.INIT('h0010)
	) name486 (
		\n680gat_reg/NET0131 ,
		_w253_,
		_w255_,
		_w256_,
		_w685_
	);
	LUT4 #(
		.INIT('h0001)
	) name487 (
		\n271gat_reg/NET0131 ,
		_w253_,
		_w255_,
		_w256_,
		_w686_
	);
	LUT4 #(
		.INIT('h0001)
	) name488 (
		_w683_,
		_w684_,
		_w685_,
		_w686_,
		_w687_
	);
	LUT3 #(
		.INIT('h3b)
	) name489 (
		_w272_,
		_w548_,
		_w687_,
		_w688_
	);
	LUT4 #(
		.INIT('h0010)
	) name490 (
		\n580gat_reg/NET0131 ,
		_w253_,
		_w255_,
		_w256_,
		_w689_
	);
	LUT4 #(
		.INIT('h0001)
	) name491 (
		\n337gat_reg/NET0131 ,
		_w253_,
		_w255_,
		_w256_,
		_w690_
	);
	LUT4 #(
		.INIT('h0100)
	) name492 (
		\n861gat_reg/NET0131 ,
		_w253_,
		_w255_,
		_w256_,
		_w691_
	);
	LUT4 #(
		.INIT('h0004)
	) name493 (
		\n777gat_reg/NET0131 ,
		_w253_,
		_w255_,
		_w256_,
		_w692_
	);
	LUT4 #(
		.INIT('h0001)
	) name494 (
		_w689_,
		_w690_,
		_w691_,
		_w692_,
		_w693_
	);
	LUT3 #(
		.INIT('h3b)
	) name495 (
		_w272_,
		_w631_,
		_w693_,
		_w694_
	);
	LUT4 #(
		.INIT('h0010)
	) name496 (
		\n816gat_reg/NET0131 ,
		_w253_,
		_w255_,
		_w256_,
		_w695_
	);
	LUT4 #(
		.INIT('h0001)
	) name497 (
		\n160gat_reg/NET0131 ,
		_w253_,
		_w255_,
		_w256_,
		_w696_
	);
	LUT4 #(
		.INIT('h0100)
	) name498 (
		\n957gat_reg/NET0131 ,
		_w253_,
		_w255_,
		_w256_,
		_w697_
	);
	LUT4 #(
		.INIT('h0004)
	) name499 (
		\n553gat_reg/NET0131 ,
		_w253_,
		_w255_,
		_w256_,
		_w698_
	);
	LUT4 #(
		.INIT('h0001)
	) name500 (
		_w695_,
		_w696_,
		_w697_,
		_w698_,
		_w699_
	);
	LUT3 #(
		.INIT('h3b)
	) name501 (
		_w272_,
		_w502_,
		_w699_,
		_w700_
	);
	LUT4 #(
		.INIT('h0004)
	) name502 (
		\n322gat_reg/NET0131 ,
		_w253_,
		_w255_,
		_w256_,
		_w701_
	);
	LUT4 #(
		.INIT('h0100)
	) name503 (
		\n865gat_reg/NET0131 ,
		_w253_,
		_w255_,
		_w256_,
		_w702_
	);
	LUT4 #(
		.INIT('h0010)
	) name504 (
		\n584gat_reg/NET0131 ,
		_w253_,
		_w255_,
		_w256_,
		_w703_
	);
	LUT4 #(
		.INIT('h0001)
	) name505 (
		\n341gat_reg/NET0131 ,
		_w253_,
		_w255_,
		_w256_,
		_w704_
	);
	LUT4 #(
		.INIT('h0001)
	) name506 (
		_w701_,
		_w702_,
		_w703_,
		_w704_,
		_w705_
	);
	LUT3 #(
		.INIT('h3b)
	) name507 (
		_w272_,
		_w631_,
		_w705_,
		_w706_
	);
	LUT4 #(
		.INIT('h0004)
	) name508 (
		\n314gat_reg/NET0131 ,
		_w253_,
		_w255_,
		_w256_,
		_w707_
	);
	LUT4 #(
		.INIT('h0100)
	) name509 (
		\n1148gat_reg/NET0131 ,
		_w253_,
		_w255_,
		_w256_,
		_w708_
	);
	LUT4 #(
		.INIT('h0001)
	) name510 (
		\n398gat_reg/NET0131 ,
		_w253_,
		_w255_,
		_w256_,
		_w709_
	);
	LUT4 #(
		.INIT('h0010)
	) name511 (
		\n699gat_reg/NET0131 ,
		_w253_,
		_w255_,
		_w256_,
		_w710_
	);
	LUT4 #(
		.INIT('h0001)
	) name512 (
		_w707_,
		_w708_,
		_w709_,
		_w710_,
		_w711_
	);
	LUT3 #(
		.INIT('h3b)
	) name513 (
		_w272_,
		_w443_,
		_w711_,
		_w712_
	);
	LUT4 #(
		.INIT('h0004)
	) name514 (
		\n318gat_reg/NET0131 ,
		_w253_,
		_w255_,
		_w256_,
		_w713_
	);
	LUT4 #(
		.INIT('h0100)
	) name515 (
		\n1080gat_reg/NET0131 ,
		_w253_,
		_w255_,
		_w256_,
		_w714_
	);
	LUT4 #(
		.INIT('h0001)
	) name516 (
		\n402gat_reg/NET0131 ,
		_w253_,
		_w255_,
		_w256_,
		_w715_
	);
	LUT4 #(
		.INIT('h0010)
	) name517 (
		\n684gat_reg/NET0131 ,
		_w253_,
		_w255_,
		_w256_,
		_w716_
	);
	LUT4 #(
		.INIT('h0001)
	) name518 (
		_w713_,
		_w714_,
		_w715_,
		_w716_,
		_w717_
	);
	LUT3 #(
		.INIT('h3b)
	) name519 (
		_w272_,
		_w469_,
		_w717_,
		_w718_
	);
	LUT4 #(
		.INIT('h0004)
	) name520 (
		\n561gat_reg/NET0131 ,
		_w253_,
		_w255_,
		_w256_,
		_w719_
	);
	LUT4 #(
		.INIT('h0100)
	) name521 (
		\n1294gat_reg/NET0131 ,
		_w253_,
		_w255_,
		_w256_,
		_w720_
	);
	LUT4 #(
		.INIT('h0010)
	) name522 (
		\n824gat_reg/NET0131 ,
		_w253_,
		_w255_,
		_w256_,
		_w721_
	);
	LUT4 #(
		.INIT('h0001)
	) name523 (
		\n846gat_reg/NET0131 ,
		_w253_,
		_w255_,
		_w256_,
		_w722_
	);
	LUT4 #(
		.INIT('h0001)
	) name524 (
		_w719_,
		_w720_,
		_w721_,
		_w722_,
		_w723_
	);
	LUT3 #(
		.INIT('h3b)
	) name525 (
		_w272_,
		_w300_,
		_w723_,
		_w724_
	);
	LUT3 #(
		.INIT('h0e)
	) name526 (
		\n919gat_reg/NET0131 ,
		_w253_,
		_w256_,
		_w725_
	);
	LUT3 #(
		.INIT('h13)
	) name527 (
		\n673gat_reg/NET0131 ,
		_w255_,
		_w256_,
		_w726_
	);
	LUT4 #(
		.INIT('h0004)
	) name528 (
		\n366gat_reg/NET0131 ,
		_w253_,
		_w255_,
		_w256_,
		_w727_
	);
	LUT4 #(
		.INIT('h0010)
	) name529 (
		\n883gat_reg/NET0131 ,
		_w253_,
		_w255_,
		_w256_,
		_w728_
	);
	LUT4 #(
		.INIT('h000b)
	) name530 (
		_w725_,
		_w726_,
		_w727_,
		_w728_,
		_w729_
	);
	LUT3 #(
		.INIT('hce)
	) name531 (
		_w272_,
		_w665_,
		_w729_,
		_w730_
	);
	LUT3 #(
		.INIT('h70)
	) name532 (
		_w267_,
		_w271_,
		_w444_,
		_w731_
	);
	LUT4 #(
		.INIT('h007f)
	) name533 (
		_w259_,
		_w263_,
		_w444_,
		_w731_,
		_w732_
	);
	LUT4 #(
		.INIT('h0100)
	) name534 (
		\n271gat_reg/NET0131 ,
		_w253_,
		_w255_,
		_w256_,
		_w733_
	);
	LUT4 #(
		.INIT('h0004)
	) name535 (
		\n1035gat_reg/NET0131 ,
		_w253_,
		_w255_,
		_w256_,
		_w734_
	);
	LUT4 #(
		.INIT('h0010)
	) name536 (
		\n834gat_reg/NET0131 ,
		_w253_,
		_w255_,
		_w256_,
		_w735_
	);
	LUT3 #(
		.INIT('h01)
	) name537 (
		_w733_,
		_w734_,
		_w735_,
		_w736_
	);
	LUT4 #(
		.INIT('h0537)
	) name538 (
		_w269_,
		_w275_,
		_w687_,
		_w736_,
		_w737_
	);
	LUT4 #(
		.INIT('h0004)
	) name539 (
		\n1072gat_reg/NET0131 ,
		_w253_,
		_w255_,
		_w256_,
		_w738_
	);
	LUT4 #(
		.INIT('h0100)
	) name540 (
		\n337gat_reg/NET0131 ,
		_w253_,
		_w255_,
		_w256_,
		_w739_
	);
	LUT4 #(
		.INIT('h0010)
	) name541 (
		\n838gat_reg/NET0131 ,
		_w253_,
		_w255_,
		_w256_,
		_w740_
	);
	LUT3 #(
		.INIT('h01)
	) name542 (
		_w738_,
		_w739_,
		_w740_,
		_w741_
	);
	LUT4 #(
		.INIT('h0537)
	) name543 (
		_w269_,
		_w275_,
		_w693_,
		_w741_,
		_w742_
	);
	LUT4 #(
		.INIT('h0004)
	) name544 (
		\n1121gat_reg/NET0131 ,
		_w253_,
		_w255_,
		_w256_,
		_w743_
	);
	LUT4 #(
		.INIT('h0100)
	) name545 (
		\n160gat_reg/NET0131 ,
		_w253_,
		_w255_,
		_w256_,
		_w744_
	);
	LUT4 #(
		.INIT('h0010)
	) name546 (
		\n707gat_reg/NET0131 ,
		_w253_,
		_w255_,
		_w256_,
		_w745_
	);
	LUT3 #(
		.INIT('h01)
	) name547 (
		_w743_,
		_w744_,
		_w745_,
		_w746_
	);
	LUT4 #(
		.INIT('h0537)
	) name548 (
		_w269_,
		_w275_,
		_w699_,
		_w746_,
		_w747_
	);
	LUT4 #(
		.INIT('h0004)
	) name549 (
		\n931gat_reg/NET0131 ,
		_w253_,
		_w255_,
		_w256_,
		_w748_
	);
	LUT4 #(
		.INIT('h0100)
	) name550 (
		\n341gat_reg/NET0131 ,
		_w253_,
		_w255_,
		_w256_,
		_w749_
	);
	LUT4 #(
		.INIT('h0010)
	) name551 (
		\n614gat_reg/NET0131 ,
		_w253_,
		_w255_,
		_w256_,
		_w750_
	);
	LUT3 #(
		.INIT('h01)
	) name552 (
		_w748_,
		_w749_,
		_w750_,
		_w751_
	);
	LUT4 #(
		.INIT('h0537)
	) name553 (
		_w269_,
		_w275_,
		_w705_,
		_w751_,
		_w752_
	);
	LUT4 #(
		.INIT('h0004)
	) name554 (
		\n1045gat_reg/NET0131 ,
		_w253_,
		_w255_,
		_w256_,
		_w753_
	);
	LUT4 #(
		.INIT('hfeef)
	) name555 (
		\n398gat_reg/NET0131 ,
		_w253_,
		_w255_,
		_w256_,
		_w754_
	);
	LUT4 #(
		.INIT('he0ee)
	) name556 (
		_w272_,
		_w274_,
		_w753_,
		_w754_,
		_w755_
	);
	LUT3 #(
		.INIT('hf1)
	) name557 (
		_w269_,
		_w711_,
		_w755_,
		_w756_
	);
	LUT4 #(
		.INIT('h0004)
	) name558 (
		\n1135gat_reg/NET0131 ,
		_w253_,
		_w255_,
		_w256_,
		_w757_
	);
	LUT4 #(
		.INIT('hfeef)
	) name559 (
		\n402gat_reg/NET0131 ,
		_w253_,
		_w255_,
		_w256_,
		_w758_
	);
	LUT4 #(
		.INIT('he0ee)
	) name560 (
		_w272_,
		_w274_,
		_w757_,
		_w758_,
		_w759_
	);
	LUT3 #(
		.INIT('hf1)
	) name561 (
		_w269_,
		_w717_,
		_w759_,
		_w760_
	);
	LUT4 #(
		.INIT('h0004)
	) name562 (
		\n1282gat_reg/NET0131 ,
		_w253_,
		_w255_,
		_w256_,
		_w761_
	);
	LUT4 #(
		.INIT('hfeef)
	) name563 (
		\n846gat_reg/NET0131 ,
		_w253_,
		_w255_,
		_w256_,
		_w762_
	);
	LUT4 #(
		.INIT('he0ee)
	) name564 (
		_w272_,
		_w274_,
		_w761_,
		_w762_,
		_w763_
	);
	LUT3 #(
		.INIT('hf1)
	) name565 (
		_w269_,
		_w723_,
		_w763_,
		_w764_
	);
	LUT4 #(
		.INIT('h0004)
	) name566 (
		\n1226gat_reg/NET0131 ,
		_w253_,
		_w255_,
		_w256_,
		_w765_
	);
	LUT4 #(
		.INIT('hfeef)
	) name567 (
		\n919gat_reg/NET0131 ,
		_w253_,
		_w255_,
		_w256_,
		_w766_
	);
	LUT4 #(
		.INIT('he0ee)
	) name568 (
		_w272_,
		_w274_,
		_w765_,
		_w766_,
		_w767_
	);
	LUT3 #(
		.INIT('hf1)
	) name569 (
		_w269_,
		_w729_,
		_w767_,
		_w768_
	);
	LUT3 #(
		.INIT('h08)
	) name570 (
		\n2343gat_reg/NET0131 ,
		\n2399gat_reg/NET0131 ,
		\n2562gat_reg/NET0131 ,
		_w769_
	);
	LUT3 #(
		.INIT('h80)
	) name571 (
		_w249_,
		_w308_,
		_w769_,
		_w770_
	);
	LUT2 #(
		.INIT('h8)
	) name572 (
		_w426_,
		_w770_,
		_w771_
	);
	LUT4 #(
		.INIT('h0155)
	) name573 (
		\n1462gat_reg/NET0131 ,
		\n1763gat_reg/NET0131 ,
		\n1880gat_reg/NET0131 ,
		\n2102gat_reg/NET0131 ,
		_w772_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name574 (
		\n1394gat_reg/NET0131 ,
		\n1767gat_reg/NET0131 ,
		\n1834gat_reg/NET0131 ,
		\n1880gat_reg/NET0131 ,
		_w773_
	);
	LUT3 #(
		.INIT('h40)
	) name575 (
		\n1508gat_reg/NET0131 ,
		_w772_,
		_w773_,
		_w774_
	);
	LUT4 #(
		.INIT('h0155)
	) name576 (
		\n1340gat_reg/NET0131 ,
		\n1763gat_reg/NET0131 ,
		\n1880gat_reg/NET0131 ,
		\n2102gat_reg/NET0131 ,
		_w775_
	);
	LUT4 #(
		.INIT('h1500)
	) name577 (
		\n1508gat_reg/NET0131 ,
		_w308_,
		_w309_,
		_w775_,
		_w776_
	);
	LUT4 #(
		.INIT('h020f)
	) name578 (
		_w314_,
		_w496_,
		_w774_,
		_w776_,
		_w777_
	);
	LUT4 #(
		.INIT('hc0d0)
	) name579 (
		\n1394gat_reg/NET0131 ,
		\n1596gat_reg/NET0131 ,
		_w380_,
		_w496_,
		_w778_
	);
	LUT2 #(
		.INIT('h2)
	) name580 (
		\n1462gat_reg/NET0131 ,
		\n1678gat_reg/NET0131 ,
		_w779_
	);
	LUT4 #(
		.INIT('h5400)
	) name581 (
		\n1678gat_reg/NET0131 ,
		\n1763gat_reg/NET0131 ,
		\n1880gat_reg/NET0131 ,
		\n2102gat_reg/NET0131 ,
		_w780_
	);
	LUT2 #(
		.INIT('h1)
	) name582 (
		_w779_,
		_w780_,
		_w781_
	);
	LUT2 #(
		.INIT('h1)
	) name583 (
		_w778_,
		_w781_,
		_w782_
	);
	LUT4 #(
		.INIT('h5400)
	) name584 (
		\n1394gat_reg/NET0131 ,
		\n1763gat_reg/NET0131 ,
		\n1880gat_reg/NET0131 ,
		\n2102gat_reg/NET0131 ,
		_w783_
	);
	LUT2 #(
		.INIT('h4)
	) name585 (
		\n1525gat_reg/NET0131 ,
		_w783_,
		_w784_
	);
	LUT4 #(
		.INIT('h8000)
	) name586 (
		\n1829gat_reg/NET0131 ,
		\n1880gat_reg/NET0131 ,
		\n2021gat_reg/NET0131 ,
		\n3097gat_pad ,
		_w785_
	);
	LUT3 #(
		.INIT('h04)
	) name587 (
		\n1775gat_reg/NET0131 ,
		\n1871gat_reg/NET0131 ,
		\n3098gat_pad ,
		_w786_
	);
	LUT3 #(
		.INIT('hd0)
	) name588 (
		\n1821gat_reg/NET0131 ,
		_w785_,
		_w786_,
		_w787_
	);
	LUT4 #(
		.INIT('h5400)
	) name589 (
		\n1588gat_reg/NET0131 ,
		\n1763gat_reg/NET0131 ,
		\n1880gat_reg/NET0131 ,
		\n2102gat_reg/NET0131 ,
		_w788_
	);
	LUT2 #(
		.INIT('h8)
	) name590 (
		\n1596gat_reg/NET0131 ,
		_w788_,
		_w789_
	);
	LUT4 #(
		.INIT('h000b)
	) name591 (
		_w314_,
		_w784_,
		_w787_,
		_w789_,
		_w790_
	);
	LUT3 #(
		.INIT('hdf)
	) name592 (
		_w777_,
		_w782_,
		_w790_,
		_w791_
	);
	LUT3 #(
		.INIT('h51)
	) name593 (
		\n1748gat_reg/NET0131 ,
		_w390_,
		_w496_,
		_w792_
	);
	LUT2 #(
		.INIT('h2)
	) name594 (
		\n1336gat_reg/NET0131 ,
		\n1748gat_reg/NET0131 ,
		_w793_
	);
	LUT4 #(
		.INIT('hc4c0)
	) name595 (
		_w314_,
		_w380_,
		_w792_,
		_w793_,
		_w794_
	);
	LUT2 #(
		.INIT('h4)
	) name596 (
		\n1675gat_reg/NET0131 ,
		_w783_,
		_w795_
	);
	LUT3 #(
		.INIT('h8c)
	) name597 (
		_w314_,
		_w380_,
		_w795_,
		_w796_
	);
	LUT4 #(
		.INIT('h1555)
	) name598 (
		\n1456gat_reg/NET0131 ,
		\n1767gat_reg/NET0131 ,
		\n1834gat_reg/NET0131 ,
		\n1880gat_reg/NET0131 ,
		_w797_
	);
	LUT2 #(
		.INIT('h1)
	) name599 (
		\n1340gat_reg/NET0131 ,
		\n1456gat_reg/NET0131 ,
		_w798_
	);
	LUT2 #(
		.INIT('h1)
	) name600 (
		_w797_,
		_w798_,
		_w799_
	);
	LUT2 #(
		.INIT('h1)
	) name601 (
		_w496_,
		_w797_,
		_w800_
	);
	LUT3 #(
		.INIT('h13)
	) name602 (
		_w314_,
		_w799_,
		_w800_,
		_w801_
	);
	LUT2 #(
		.INIT('h2)
	) name603 (
		\n1340gat_reg/NET0131 ,
		\n1807gat_reg/NET0131 ,
		_w802_
	);
	LUT3 #(
		.INIT('h0b)
	) name604 (
		_w314_,
		_w795_,
		_w802_,
		_w803_
	);
	LUT4 #(
		.INIT('hbabb)
	) name605 (
		_w794_,
		_w796_,
		_w801_,
		_w803_,
		_w804_
	);
	LUT4 #(
		.INIT('ha800)
	) name606 (
		\n1678gat_reg/NET0131 ,
		\n1763gat_reg/NET0131 ,
		\n1880gat_reg/NET0131 ,
		\n2102gat_reg/NET0131 ,
		_w805_
	);
	LUT4 #(
		.INIT('h02aa)
	) name607 (
		\n1508gat_reg/NET0131 ,
		\n1763gat_reg/NET0131 ,
		\n1880gat_reg/NET0131 ,
		\n2102gat_reg/NET0131 ,
		_w806_
	);
	LUT4 #(
		.INIT('h1555)
	) name608 (
		\n1394gat_reg/NET0131 ,
		\n1767gat_reg/NET0131 ,
		\n1834gat_reg/NET0131 ,
		\n1880gat_reg/NET0131 ,
		_w807_
	);
	LUT3 #(
		.INIT('h02)
	) name609 (
		\n1871gat_reg/NET0131 ,
		\n2592gat_reg/NET0131 ,
		\n673gat_reg/NET0131 ,
		_w808_
	);
	LUT4 #(
		.INIT('h5551)
	) name610 (
		\n1389gat_reg/NET0131 ,
		\n1871gat_reg/NET0131 ,
		\n2592gat_reg/NET0131 ,
		\n673gat_reg/NET0131 ,
		_w809_
	);
	LUT4 #(
		.INIT('hef00)
	) name611 (
		_w805_,
		_w806_,
		_w807_,
		_w809_,
		_w810_
	);
	LUT4 #(
		.INIT('hec00)
	) name612 (
		_w248_,
		_w496_,
		_w571_,
		_w769_,
		_w811_
	);
	LUT4 #(
		.INIT('hd050)
	) name613 (
		\n2084gat_reg/NET0131 ,
		_w248_,
		_w427_,
		_w571_,
		_w812_
	);
	LUT2 #(
		.INIT('h1)
	) name614 (
		_w811_,
		_w812_,
		_w813_
	);
	LUT4 #(
		.INIT('h1000)
	) name615 (
		\n1068gat_reg/NET0131 ,
		\n2343gat_reg/NET0131 ,
		\n2399gat_reg/NET0131 ,
		\n2562gat_reg/NET0131 ,
		_w814_
	);
	LUT4 #(
		.INIT('h0002)
	) name616 (
		\n2343gat_reg/NET0131 ,
		\n2399gat_reg/NET0131 ,
		\n2562gat_reg/NET0131 ,
		\n865gat_reg/NET0131 ,
		_w815_
	);
	LUT4 #(
		.INIT('h0020)
	) name617 (
		\n2343gat_reg/NET0131 ,
		\n2399gat_reg/NET0131 ,
		\n2562gat_reg/NET0131 ,
		\n957gat_reg/NET0131 ,
		_w816_
	);
	LUT4 #(
		.INIT('h0004)
	) name618 (
		\n2343gat_reg/NET0131 ,
		\n2399gat_reg/NET0131 ,
		\n2562gat_reg/NET0131 ,
		\n861gat_reg/NET0131 ,
		_w817_
	);
	LUT4 #(
		.INIT('h0001)
	) name619 (
		_w814_,
		_w815_,
		_w816_,
		_w817_,
		_w818_
	);
	LUT4 #(
		.INIT('h0020)
	) name620 (
		\n2343gat_reg/NET0131 ,
		\n2399gat_reg/NET0131 ,
		\n2562gat_reg/NET0131 ,
		\n816gat_reg/NET0131 ,
		_w819_
	);
	LUT4 #(
		.INIT('h0040)
	) name621 (
		\n2343gat_reg/NET0131 ,
		\n2399gat_reg/NET0131 ,
		\n2562gat_reg/NET0131 ,
		\n680gat_reg/NET0131 ,
		_w820_
	);
	LUT4 #(
		.INIT('h0004)
	) name622 (
		\n2343gat_reg/NET0131 ,
		\n2399gat_reg/NET0131 ,
		\n2562gat_reg/NET0131 ,
		\n580gat_reg/NET0131 ,
		_w821_
	);
	LUT4 #(
		.INIT('h0002)
	) name623 (
		\n2343gat_reg/NET0131 ,
		\n2399gat_reg/NET0131 ,
		\n2562gat_reg/NET0131 ,
		\n584gat_reg/NET0131 ,
		_w822_
	);
	LUT4 #(
		.INIT('h0001)
	) name624 (
		_w819_,
		_w820_,
		_w821_,
		_w822_,
		_w823_
	);
	LUT3 #(
		.INIT('he4)
	) name625 (
		_w390_,
		_w818_,
		_w823_,
		_w824_
	);
	LUT4 #(
		.INIT('h8000)
	) name626 (
		\n1767gat_reg/NET0131 ,
		\n1834gat_reg/NET0131 ,
		\n1880gat_reg/NET0131 ,
		\n699gat_reg/NET0131 ,
		_w825_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name627 (
		\n1148gat_reg/NET0131 ,
		\n1767gat_reg/NET0131 ,
		\n1834gat_reg/NET0131 ,
		\n1880gat_reg/NET0131 ,
		_w826_
	);
	LUT2 #(
		.INIT('h1)
	) name628 (
		\n2343gat_reg/NET0131 ,
		\n2399gat_reg/NET0131 ,
		_w827_
	);
	LUT3 #(
		.INIT('h80)
	) name629 (
		\n2203gat_reg/NET0131 ,
		\n2207gat_reg/NET0131 ,
		\n2562gat_reg/NET0131 ,
		_w828_
	);
	LUT4 #(
		.INIT('h1000)
	) name630 (
		_w825_,
		_w826_,
		_w827_,
		_w828_,
		_w829_
	);
	LUT4 #(
		.INIT('h8000)
	) name631 (
		\n1767gat_reg/NET0131 ,
		\n1834gat_reg/NET0131 ,
		\n1880gat_reg/NET0131 ,
		\n684gat_reg/NET0131 ,
		_w830_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name632 (
		\n1080gat_reg/NET0131 ,
		\n1767gat_reg/NET0131 ,
		\n1834gat_reg/NET0131 ,
		\n1880gat_reg/NET0131 ,
		_w831_
	);
	LUT3 #(
		.INIT('h08)
	) name633 (
		\n2203gat_reg/NET0131 ,
		\n2207gat_reg/NET0131 ,
		\n2562gat_reg/NET0131 ,
		_w832_
	);
	LUT4 #(
		.INIT('h0200)
	) name634 (
		_w827_,
		_w830_,
		_w831_,
		_w832_,
		_w833_
	);
	LUT2 #(
		.INIT('h1)
	) name635 (
		_w829_,
		_w833_,
		_w834_
	);
	LUT4 #(
		.INIT('hd500)
	) name636 (
		_w597_,
		_w813_,
		_w824_,
		_w834_,
		_w835_
	);
	LUT4 #(
		.INIT('h00ef)
	) name637 (
		_w805_,
		_w806_,
		_w807_,
		_w808_,
		_w836_
	);
	LUT4 #(
		.INIT('h0400)
	) name638 (
		\n160gat_reg/NET0131 ,
		\n2343gat_reg/NET0131 ,
		\n2399gat_reg/NET0131 ,
		\n2562gat_reg/NET0131 ,
		_w837_
	);
	LUT4 #(
		.INIT('h0040)
	) name639 (
		\n2343gat_reg/NET0131 ,
		\n2399gat_reg/NET0131 ,
		\n2562gat_reg/NET0131 ,
		\n271gat_reg/NET0131 ,
		_w838_
	);
	LUT2 #(
		.INIT('h1)
	) name640 (
		_w837_,
		_w838_,
		_w839_
	);
	LUT4 #(
		.INIT('h0004)
	) name641 (
		\n2343gat_reg/NET0131 ,
		\n2399gat_reg/NET0131 ,
		\n2562gat_reg/NET0131 ,
		\n337gat_reg/NET0131 ,
		_w840_
	);
	LUT4 #(
		.INIT('h0002)
	) name642 (
		\n2343gat_reg/NET0131 ,
		\n2399gat_reg/NET0131 ,
		\n2562gat_reg/NET0131 ,
		\n341gat_reg/NET0131 ,
		_w841_
	);
	LUT3 #(
		.INIT('h01)
	) name643 (
		_w390_,
		_w840_,
		_w841_,
		_w842_
	);
	LUT4 #(
		.INIT('h0002)
	) name644 (
		\n2343gat_reg/NET0131 ,
		\n2399gat_reg/NET0131 ,
		\n2562gat_reg/NET0131 ,
		\n614gat_reg/NET0131 ,
		_w843_
	);
	LUT2 #(
		.INIT('h2)
	) name645 (
		_w390_,
		_w843_,
		_w844_
	);
	LUT4 #(
		.INIT('h0020)
	) name646 (
		\n2343gat_reg/NET0131 ,
		\n2399gat_reg/NET0131 ,
		\n2562gat_reg/NET0131 ,
		\n707gat_reg/NET0131 ,
		_w845_
	);
	LUT4 #(
		.INIT('h0004)
	) name647 (
		\n2343gat_reg/NET0131 ,
		\n2399gat_reg/NET0131 ,
		\n2562gat_reg/NET0131 ,
		\n838gat_reg/NET0131 ,
		_w846_
	);
	LUT4 #(
		.INIT('h0040)
	) name648 (
		\n2343gat_reg/NET0131 ,
		\n2399gat_reg/NET0131 ,
		\n2562gat_reg/NET0131 ,
		\n834gat_reg/NET0131 ,
		_w847_
	);
	LUT3 #(
		.INIT('h01)
	) name649 (
		_w845_,
		_w846_,
		_w847_,
		_w848_
	);
	LUT4 #(
		.INIT('h0777)
	) name650 (
		_w839_,
		_w842_,
		_w844_,
		_w848_,
		_w849_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name651 (
		\n1294gat_reg/NET0131 ,
		\n1767gat_reg/NET0131 ,
		\n1834gat_reg/NET0131 ,
		\n1880gat_reg/NET0131 ,
		_w850_
	);
	LUT4 #(
		.INIT('h8000)
	) name652 (
		\n1767gat_reg/NET0131 ,
		\n1834gat_reg/NET0131 ,
		\n1880gat_reg/NET0131 ,
		\n824gat_reg/NET0131 ,
		_w851_
	);
	LUT3 #(
		.INIT('h02)
	) name653 (
		_w427_,
		_w850_,
		_w851_,
		_w852_
	);
	LUT4 #(
		.INIT('h7f00)
	) name654 (
		\n1767gat_reg/NET0131 ,
		\n1834gat_reg/NET0131 ,
		\n1880gat_reg/NET0131 ,
		\n673gat_reg/NET0131 ,
		_w853_
	);
	LUT4 #(
		.INIT('h8000)
	) name655 (
		\n1767gat_reg/NET0131 ,
		\n1834gat_reg/NET0131 ,
		\n1880gat_reg/NET0131 ,
		\n883gat_reg/NET0131 ,
		_w854_
	);
	LUT3 #(
		.INIT('h02)
	) name656 (
		_w769_,
		_w853_,
		_w854_,
		_w855_
	);
	LUT2 #(
		.INIT('h1)
	) name657 (
		_w852_,
		_w855_,
		_w856_
	);
	LUT2 #(
		.INIT('h4)
	) name658 (
		\n2203gat_reg/NET0131 ,
		\n2207gat_reg/NET0131 ,
		_w857_
	);
	LUT4 #(
		.INIT('h20aa)
	) name659 (
		_w836_,
		_w849_,
		_w856_,
		_w857_,
		_w858_
	);
	LUT4 #(
		.INIT('h0096)
	) name660 (
		\n318gat_reg/NET0131 ,
		\n322gat_reg/NET0131 ,
		\n659gat_reg/NET0131 ,
		\n919gat_reg/NET0131 ,
		_w859_
	);
	LUT4 #(
		.INIT('hff96)
	) name661 (
		\n318gat_reg/NET0131 ,
		\n322gat_reg/NET0131 ,
		\n659gat_reg/NET0131 ,
		\n919gat_reg/NET0131 ,
		_w860_
	);
	LUT4 #(
		.INIT('h6f09)
	) name662 (
		_w250_,
		_w251_,
		_w859_,
		_w860_,
		_w861_
	);
	LUT2 #(
		.INIT('h8)
	) name663 (
		_w308_,
		_w427_,
		_w862_
	);
	LUT4 #(
		.INIT('h9600)
	) name664 (
		\n318gat_reg/NET0131 ,
		\n322gat_reg/NET0131 ,
		\n659gat_reg/NET0131 ,
		\n919gat_reg/NET0131 ,
		_w863_
	);
	LUT3 #(
		.INIT('h60)
	) name665 (
		_w250_,
		_w251_,
		_w863_,
		_w864_
	);
	LUT4 #(
		.INIT('h96ff)
	) name666 (
		\n318gat_reg/NET0131 ,
		\n322gat_reg/NET0131 ,
		\n659gat_reg/NET0131 ,
		\n919gat_reg/NET0131 ,
		_w865_
	);
	LUT4 #(
		.INIT('h0f9f)
	) name667 (
		_w250_,
		_w251_,
		_w496_,
		_w865_,
		_w866_
	);
	LUT4 #(
		.INIT('h0008)
	) name668 (
		_w861_,
		_w862_,
		_w864_,
		_w866_,
		_w867_
	);
	LUT4 #(
		.INIT('h0010)
	) name669 (
		\n2343gat_reg/NET0131 ,
		\n2399gat_reg/NET0131 ,
		\n2562gat_reg/NET0131 ,
		\n561gat_reg/NET0131 ,
		_w868_
	);
	LUT4 #(
		.INIT('h0080)
	) name670 (
		\n2343gat_reg/NET0131 ,
		\n2399gat_reg/NET0131 ,
		\n2562gat_reg/NET0131 ,
		\n659gat_reg/NET0131 ,
		_w869_
	);
	LUT4 #(
		.INIT('h0002)
	) name671 (
		\n2343gat_reg/NET0131 ,
		\n2399gat_reg/NET0131 ,
		\n2562gat_reg/NET0131 ,
		\n318gat_reg/NET0131 ,
		_w870_
	);
	LUT4 #(
		.INIT('h0008)
	) name672 (
		\n2343gat_reg/NET0131 ,
		\n2399gat_reg/NET0131 ,
		\n2562gat_reg/NET0131 ,
		\n777gat_reg/NET0131 ,
		_w871_
	);
	LUT4 #(
		.INIT('h0001)
	) name673 (
		_w868_,
		_w869_,
		_w870_,
		_w871_,
		_w872_
	);
	LUT4 #(
		.INIT('h0004)
	) name674 (
		\n2343gat_reg/NET0131 ,
		\n2399gat_reg/NET0131 ,
		\n2562gat_reg/NET0131 ,
		\n322gat_reg/NET0131 ,
		_w873_
	);
	LUT4 #(
		.INIT('h0020)
	) name675 (
		\n2343gat_reg/NET0131 ,
		\n2399gat_reg/NET0131 ,
		\n2562gat_reg/NET0131 ,
		\n314gat_reg/NET0131 ,
		_w874_
	);
	LUT4 #(
		.INIT('h0040)
	) name676 (
		\n2343gat_reg/NET0131 ,
		\n2399gat_reg/NET0131 ,
		\n2562gat_reg/NET0131 ,
		\n553gat_reg/NET0131 ,
		_w875_
	);
	LUT4 #(
		.INIT('h0001)
	) name677 (
		\n2343gat_reg/NET0131 ,
		\n2399gat_reg/NET0131 ,
		\n2562gat_reg/NET0131 ,
		\n366gat_reg/NET0131 ,
		_w876_
	);
	LUT4 #(
		.INIT('h0001)
	) name678 (
		_w873_,
		_w874_,
		_w875_,
		_w876_,
		_w877_
	);
	LUT2 #(
		.INIT('h8)
	) name679 (
		_w317_,
		_w496_,
		_w878_
	);
	LUT4 #(
		.INIT('h4055)
	) name680 (
		_w405_,
		_w872_,
		_w877_,
		_w878_,
		_w879_
	);
	LUT2 #(
		.INIT('h4)
	) name681 (
		_w867_,
		_w879_,
		_w880_
	);
	LUT4 #(
		.INIT('h15ff)
	) name682 (
		_w810_,
		_w835_,
		_w858_,
		_w880_,
		_w881_
	);
	LUT4 #(
		.INIT('h80aa)
	) name683 (
		_w600_,
		_w872_,
		_w877_,
		_w878_,
		_w882_
	);
	LUT2 #(
		.INIT('h4)
	) name684 (
		_w867_,
		_w882_,
		_w883_
	);
	LUT4 #(
		.INIT('h15ff)
	) name685 (
		_w810_,
		_w835_,
		_w858_,
		_w883_,
		_w884_
	);
	LUT3 #(
		.INIT('h80)
	) name686 (
		\n1771gat_reg/NET0131 ,
		\n1775gat_reg/NET0131 ,
		\n2514gat_reg/NET0131 ,
		_w885_
	);
	LUT2 #(
		.INIT('h1)
	) name687 (
		_w496_,
		_w885_,
		_w886_
	);
	LUT2 #(
		.INIT('h8)
	) name688 (
		_w314_,
		_w886_,
		_w887_
	);
	LUT4 #(
		.INIT('h8000)
	) name689 (
		\n1771gat_reg/NET0131 ,
		\n1775gat_reg/NET0131 ,
		\n1871gat_reg/NET0131 ,
		\n2514gat_reg/NET0131 ,
		_w888_
	);
	LUT3 #(
		.INIT('h80)
	) name690 (
		\n2033gat_reg/NET0131 ,
		\n2169gat_reg/NET0131 ,
		\n2176gat_reg/NET0131 ,
		_w889_
	);
	LUT3 #(
		.INIT('h80)
	) name691 (
		\n2037gat_reg/NET0131 ,
		\n2095gat_reg/NET0131 ,
		\n2110gat_reg/NET0131 ,
		_w890_
	);
	LUT3 #(
		.INIT('h40)
	) name692 (
		_w888_,
		_w889_,
		_w890_,
		_w891_
	);
	LUT2 #(
		.INIT('h1)
	) name693 (
		\n2454gat_reg/NET0131 ,
		\n337gat_reg/NET0131 ,
		_w892_
	);
	LUT2 #(
		.INIT('hd)
	) name694 (
		_w456_,
		_w892_,
		_w893_
	);
	LUT3 #(
		.INIT('h80)
	) name695 (
		_w254_,
		_w337_,
		_w669_,
		_w894_
	);
	LUT3 #(
		.INIT('h4c)
	) name696 (
		_w341_,
		_w449_,
		_w667_,
		_w895_
	);
	LUT2 #(
		.INIT('hb)
	) name697 (
		_w894_,
		_w895_,
		_w896_
	);
	assign \_al_n0  = 1'b0;
	assign \g17_dup/_0_  = _w249_ ;
	assign \g6952/_2_  = _w290_ ;
	assign \g6953/_2_  = _w293_ ;
	assign \g6961/_0_  = _w300_ ;
	assign \g7076/_0_  = _w321_ ;
	assign \g7077/_0_  = _w324_ ;
	assign \g7079/_0_  = _w327_ ;
	assign \g7081/_0_  = _w330_ ;
	assign \g7082/_0_  = _w333_ ;
	assign \g7083/_0_  = _w336_ ;
	assign \g7146/_0_  = _w347_ ;
	assign \g7147/_0_  = _w349_ ;
	assign \g7148/_0_  = _w351_ ;
	assign \g7149/_0_  = _w353_ ;
	assign \g7150/_0_  = _w355_ ;
	assign \g7151/_0_  = _w357_ ;
	assign \g7152/_0_  = _w359_ ;
	assign \g7153/_0_  = _w361_ ;
	assign \g7154/_0_  = _w363_ ;
	assign \g7156/_2_  = _w399_ ;
	assign \g7161/_2_  = _w401_ ;
	assign \g7165/_2_  = _w406_ ;
	assign \g7174/_0_  = _w407_ ;
	assign \g7180/_00_  = _w424_ ;
	assign \g7182/_3_  = _w428_ ;
	assign \g7191/_0_  = _w436_ ;
	assign \g7204/_0_  = _w439_ ;
	assign \g7209/_3_  = _w443_ ;
	assign \g7220/_0_  = _w140_ ;
	assign \g7229/_0_  = _w444_ ;
	assign \g7233/_0_  = _w447_ ;
	assign \g7234/_0_  = _w451_ ;
	assign \g7235/_0_  = _w454_ ;
	assign \g7236/_0_  = _w458_ ;
	assign \g7237/_0_  = _w461_ ;
	assign \g7238/_0_  = _w465_ ;
	assign \g7241/_3_  = _w469_ ;
	assign \g7264/_0_  = _w475_ ;
	assign \g7265/_0_  = _w477_ ;
	assign \g7266/_0_  = _w484_ ;
	assign \g7267/_0_  = _w487_ ;
	assign \g7268/_0_  = _w489_ ;
	assign \g7301/_0_  = _w492_ ;
	assign \g7326/_3_  = _w495_ ;
	assign \g7350/_2_  = _w497_ ;
	assign \g7352/_0_  = _w237_ ;
	assign \g7356/_0_  = _w498_ ;
	assign \g7359/_0_  = _w429_ ;
	assign \g7389/_3_  = _w502_ ;
	assign \g7417/_0_  = _w508_ ;
	assign \g7418/_0_  = _w510_ ;
	assign \g7419/_0_  = _w512_ ;
	assign \g7444/_0_  = _w527_ ;
	assign \g7445/_0_  = _w537_ ;
	assign \g7449/_3_  = _w544_ ;
	assign \g7451/_3_  = _w548_ ;
	assign \g7454/_0_  = _w225_ ;
	assign \g7467/_3_  = _w555_ ;
	assign \g7476/_0_  = _w215_ ;
	assign \g7480/_0_  = _w563_ ;
	assign \g7494/_0_  = _w570_ ;
	assign \g7509/_0_  = _w92_ ;
	assign \g7514/_0_  = _w574_ ;
	assign \g7517/_3_  = _w580_ ;
	assign \g7524/_0_  = _w76_ ;
	assign \g7558/_0_  = _w584_ ;
	assign \g7560/_0_  = _w588_ ;
	assign \g7561/_0_  = _w592_ ;
	assign \g7563/_0_  = _w596_ ;
	assign \g7567/_0_  = _w600_ ;
	assign \g7572/_0_  = _w51_ ;
	assign \g7579/_0_  = _w602_ ;
	assign \g7605/_0_  = _w606_ ;
	assign \g7625/_0_  = _w607_ ;
	assign \g7627/_0_  = _w608_ ;
	assign \g7671/_0_  = _w609_ ;
	assign \g7675/_0_  = _w613_ ;
	assign \g7689/_0_  = _w614_ ;
	assign \g7697/_0_  = _w616_ ;
	assign \g7743/_1_  = _w504_ ;
	assign \g7764/_1_  = _w511_ ;
	assign \g7769/_0_  = _w617_ ;
	assign \g7771/_2_  = _w615_ ;
	assign \g7779/_0_  = _w619_ ;
	assign \g7852/_0_  = _w621_ ;
	assign \g7873/_0_  = _w622_ ;
	assign \g7884/_3_  = _w412_ ;
	assign \g7889/_0_  = _w80_ ;
	assign \g7902/_1_  = _w509_ ;
	assign \g7992/_3_  = _w624_ ;
	assign \g7994/_3_  = _w323_ ;
	assign \g7996/_3_  = _w329_ ;
	assign \g7998/_3_  = _w626_ ;
	assign \g8000/_3_  = _w628_ ;
	assign \g8002/_3_  = _w302_ ;
	assign \g8004/_3_  = _w335_ ;
	assign \g8006/_3_  = _w332_ ;
	assign \g8008/_3_  = _w326_ ;
	assign \g8150/_0_  = _w151_ ;
	assign \g8151/_0_  = _w132_ ;
	assign \g8157/_0_  = _w68_ ;
	assign \g8163/_0_  = _w233_ ;
	assign \g8172/_0_  = _w130_ ;
	assign \g8197/_0_  = _w235_ ;
	assign \g8211/_0_  = _w142_ ;
	assign \g8223/_0_  = _w155_ ;
	assign \g8237/_0_  = _w97_ ;
	assign \g8251/_0_  = _w157_ ;
	assign \g8261/_0_  = _w229_ ;
	assign \g8272/_0_  = _w17_ ;
	assign \g8287/_0_  = _w223_ ;
	assign \g8647/_0_  = _w99_ ;
	assign \g8671/_0_  = _w108_ ;
	assign \g8672/_0_  = _w114_ ;
	assign \g8735/_0_  = _w631_ ;
	assign \g8766/_0_  = _w632_ ;
	assign \g8811/_0_  = _w633_ ;
	assign \g8821/_0_  = _w642_ ;
	assign \g8856/_0_  = _w471_ ;
	assign \g8858/_3_  = _w448_ ;
	assign \g8868/_0_  = _w381_ ;
	assign \g8880/_2_  = _w643_ ;
	assign \g8886/_0_  = _w651_ ;
	assign \g8900/_0_  = _w652_ ;
	assign \g8932/_0_  = _w659_ ;
	assign \g8991/_3_  = _w660_ ;
	assign \g9014/_3_  = _w664_ ;
	assign \g9074/_0_  = _w415_ ;
	assign \g9091/_0_  = _w149_ ;
	assign \g9105/_0_  = _w153_ ;
	assign \g9107/_1_  = _w315_ ;
	assign \g9111/_0_  = _w666_ ;
	assign \n1332gat_reg/P0001  = _w19_ ;
	assign \n1363gat_reg/P0001  = _w23_ ;
	assign \n1394gat_reg/P0001  = _w26_ ;
	assign \n1433gat_reg/P0001  = _w28_ ;
	assign \n1775gat_reg/P0001  = _w48_ ;
	assign \n2025gat_reg/P0001  = _w62_ ;
	assign \n2029gat_reg/P0001  = _w64_ ;
	assign \n2033gat_reg/P0001  = _w66_ ;
	assign \n2044gat_reg/P0001  = _w71_ ;
	assign \n2121gat_reg/P0001  = _w83_ ;
	assign \n2125gat_reg/P0001  = _w85_ ;
	assign \n2458gat_reg/P0001  = _w123_ ;
	assign \n2472gat_reg/P0001  = _w127_ ;
	assign \n2592gat_reg/P0001  = _w146_ ;
	assign \n3104gat_pad  = _w671_ ;
	assign \n3105gat_pad  = _w674_ ;
	assign \n3106gat_pad  = _w56_ ;
	assign \n3107gat_pad  = _w675_ ;
	assign \n3108gat_pad  = _w676_ ;
	assign \n3109gat_pad  = _w677_ ;
	assign \n3110gat_pad  = _w678_ ;
	assign \n3111gat_pad  = _w679_ ;
	assign \n3112gat_pad  = 1'b1;
	assign \n3113gat_pad  = _w680_ ;
	assign \n3114gat_pad  = _w681_ ;
	assign \n3116gat_pad  = _w682_ ;
	assign \n3117gat_pad  = _w688_ ;
	assign \n3118gat_pad  = _w694_ ;
	assign \n3119gat_pad  = _w700_ ;
	assign \n3120gat_pad  = _w706_ ;
	assign \n3121gat_pad  = _w712_ ;
	assign \n3122gat_pad  = _w718_ ;
	assign \n3123gat_pad  = _w724_ ;
	assign \n3124gat_pad  = _w730_ ;
	assign \n3125gat_pad  = _w732_ ;
	assign \n3126gat_pad  = _w106_ ;
	assign \n3127gat_pad  = _w103_ ;
	assign \n3128gat_pad  = _w111_ ;
	assign \n3130gat_pad  = _w737_ ;
	assign \n3131gat_pad  = _w742_ ;
	assign \n3132gat_pad  = _w747_ ;
	assign \n3133gat_pad  = _w752_ ;
	assign \n3134gat_pad  = _w756_ ;
	assign \n3135gat_pad  = _w760_ ;
	assign \n3136gat_pad  = _w764_ ;
	assign \n3137gat_pad  = _w768_ ;
	assign \n3138gat_pad  = _w771_ ;
	assign \n3140gat_pad  = _w791_ ;
	assign \n3142gat_pad  = _w804_ ;
	assign \n3143gat_pad  = _w881_ ;
	assign \n3144gat_pad  = _w884_ ;
	assign \n3145gat_pad  = _w887_ ;
	assign \n3146gat_pad  = _w891_ ;
	assign \n3147gat_pad  = _w505_ ;
	assign \n3148gat_pad  = _w120_ ;
	assign \n3149gat_pad  = _w391_ ;
	assign \n3150gat_pad  = _w893_ ;
	assign \n3151gat_pad  = _w896_ ;
	assign \n684gat_reg/P0001  = _w221_ ;
	assign \n824gat_reg/P0001  = _w231_ ;
	assign \n883gat_reg/P0001  = _w243_ ;
endmodule;