module top (ADS_n_pad, \Address[0]_pad , \Address[10]_pad , \Address[11]_pad , \Address[12]_pad , \Address[13]_pad , \Address[14]_pad , \Address[15]_pad , \Address[16]_pad , \Address[17]_pad , \Address[18]_pad , \Address[19]_pad , \Address[1]_pad , \Address[20]_pad , \Address[21]_pad , \Address[22]_pad , \Address[23]_pad , \Address[24]_pad , \Address[25]_pad , \Address[26]_pad , \Address[27]_pad , \Address[28]_pad , \Address[29]_pad , \Address[2]_pad , \Address[3]_pad , \Address[4]_pad , \Address[5]_pad , \Address[6]_pad , \Address[7]_pad , \Address[8]_pad , \Address[9]_pad , \BE_n[0]_pad , \BE_n[1]_pad , \BE_n[2]_pad , \BE_n[3]_pad , \BS16_n_pad , \ByteEnable_reg[0]/NET0131 , \ByteEnable_reg[1]/NET0131 , \ByteEnable_reg[2]/NET0131 , \ByteEnable_reg[3]/NET0131 , \CodeFetch_reg/NET0131 , D_C_n_pad, \DataWidth_reg[0]/NET0131 , \DataWidth_reg[1]/NET0131 , \Datai[0]_pad , \Datai[10]_pad , \Datai[11]_pad , \Datai[12]_pad , \Datai[13]_pad , \Datai[14]_pad , \Datai[15]_pad , \Datai[16]_pad , \Datai[17]_pad , \Datai[18]_pad , \Datai[19]_pad , \Datai[1]_pad , \Datai[20]_pad , \Datai[21]_pad , \Datai[22]_pad , \Datai[23]_pad , \Datai[24]_pad , \Datai[25]_pad , \Datai[26]_pad , \Datai[27]_pad , \Datai[28]_pad , \Datai[29]_pad , \Datai[2]_pad , \Datai[30]_pad , \Datai[31]_pad , \Datai[3]_pad , \Datai[4]_pad , \Datai[5]_pad , \Datai[6]_pad , \Datai[7]_pad , \Datai[8]_pad , \Datai[9]_pad , \Datao[0]_pad , \Datao[10]_pad , \Datao[11]_pad , \Datao[12]_pad , \Datao[13]_pad , \Datao[14]_pad , \Datao[15]_pad , \Datao[16]_pad , \Datao[17]_pad , \Datao[18]_pad , \Datao[19]_pad , \Datao[1]_pad , \Datao[20]_pad , \Datao[21]_pad , \Datao[23]_pad , \Datao[24]_pad , \Datao[25]_pad , \Datao[26]_pad , \Datao[27]_pad , \Datao[28]_pad , \Datao[29]_pad , \Datao[2]_pad , \Datao[30]_pad , \Datao[3]_pad , \Datao[4]_pad , \Datao[5]_pad , \Datao[6]_pad , \Datao[7]_pad , \Datao[8]_pad , \Datao[9]_pad , \Datao_reg[22]/NET0131 , \EAX_reg[0]/NET0131 , \EAX_reg[10]/NET0131 , \EAX_reg[11]/NET0131 , \EAX_reg[12]/NET0131 , \EAX_reg[13]/NET0131 , \EAX_reg[14]/NET0131 , \EAX_reg[15]/NET0131 , \EAX_reg[16]/NET0131 , \EAX_reg[17]/NET0131 , \EAX_reg[18]/NET0131 , \EAX_reg[19]/NET0131 , \EAX_reg[1]/NET0131 , \EAX_reg[20]/NET0131 , \EAX_reg[21]/NET0131 , \EAX_reg[22]/NET0131 , \EAX_reg[23]/NET0131 , \EAX_reg[24]/NET0131 , \EAX_reg[25]/NET0131 , \EAX_reg[26]/NET0131 , \EAX_reg[27]/NET0131 , \EAX_reg[28]/NET0131 , \EAX_reg[29]/NET0131 , \EAX_reg[2]/NET0131 , \EAX_reg[30]/NET0131 , \EAX_reg[31]/NET0131 , \EAX_reg[3]/NET0131 , \EAX_reg[4]/NET0131 , \EAX_reg[5]/NET0131 , \EAX_reg[6]/NET0131 , \EAX_reg[7]/NET0131 , \EAX_reg[8]/NET0131 , \EAX_reg[9]/NET0131 , \EBX_reg[0]/NET0131 , \EBX_reg[10]/NET0131 , \EBX_reg[11]/NET0131 , \EBX_reg[12]/NET0131 , \EBX_reg[13]/NET0131 , \EBX_reg[14]/NET0131 , \EBX_reg[15]/NET0131 , \EBX_reg[16]/NET0131 , \EBX_reg[17]/NET0131 , \EBX_reg[18]/NET0131 , \EBX_reg[19]/NET0131 , \EBX_reg[1]/NET0131 , \EBX_reg[20]/NET0131 , \EBX_reg[21]/NET0131 , \EBX_reg[22]/NET0131 , \EBX_reg[23]/NET0131 , \EBX_reg[24]/NET0131 , \EBX_reg[25]/NET0131 , \EBX_reg[26]/NET0131 , \EBX_reg[27]/NET0131 , \EBX_reg[28]/NET0131 , \EBX_reg[29]/NET0131 , \EBX_reg[2]/NET0131 , \EBX_reg[30]/NET0131 , \EBX_reg[31]/NET0131 , \EBX_reg[3]/NET0131 , \EBX_reg[4]/NET0131 , \EBX_reg[5]/NET0131 , \EBX_reg[6]/NET0131 , \EBX_reg[7]/NET0131 , \EBX_reg[8]/NET0131 , \EBX_reg[9]/NET0131 , \Flush_reg/NET0131 , HOLD_pad, \InstAddrPointer_reg[0]/NET0131 , \InstAddrPointer_reg[10]/NET0131 , \InstAddrPointer_reg[11]/NET0131 , \InstAddrPointer_reg[12]/NET0131 , \InstAddrPointer_reg[13]/NET0131 , \InstAddrPointer_reg[14]/NET0131 , \InstAddrPointer_reg[15]/NET0131 , \InstAddrPointer_reg[16]/NET0131 , \InstAddrPointer_reg[17]/NET0131 , \InstAddrPointer_reg[18]/NET0131 , \InstAddrPointer_reg[19]/NET0131 , \InstAddrPointer_reg[1]/NET0131 , \InstAddrPointer_reg[20]/NET0131 , \InstAddrPointer_reg[21]/NET0131 , \InstAddrPointer_reg[22]/NET0131 , \InstAddrPointer_reg[23]/NET0131 , \InstAddrPointer_reg[24]/NET0131 , \InstAddrPointer_reg[25]/NET0131 , \InstAddrPointer_reg[26]/NET0131 , \InstAddrPointer_reg[27]/NET0131 , \InstAddrPointer_reg[28]/NET0131 , \InstAddrPointer_reg[29]/NET0131 , \InstAddrPointer_reg[2]/NET0131 , \InstAddrPointer_reg[30]/NET0131 , \InstAddrPointer_reg[31]/NET0131 , \InstAddrPointer_reg[3]/NET0131 , \InstAddrPointer_reg[4]/NET0131 , \InstAddrPointer_reg[5]/NET0131 , \InstAddrPointer_reg[6]/NET0131 , \InstAddrPointer_reg[7]/NET0131 , \InstAddrPointer_reg[8]/NET0131 , \InstAddrPointer_reg[9]/NET0131 , \InstQueueRd_Addr_reg[0]/NET0131 , \InstQueueRd_Addr_reg[1]/NET0131 , \InstQueueRd_Addr_reg[2]/NET0131 , \InstQueueRd_Addr_reg[3]/NET0131 , \InstQueueWr_Addr_reg[0]/NET0131 , \InstQueueWr_Addr_reg[1]/NET0131 , \InstQueueWr_Addr_reg[2]/NET0131 , \InstQueueWr_Addr_reg[3]/NET0131 , \InstQueue_reg[0][0]/NET0131 , \InstQueue_reg[0][1]/NET0131 , \InstQueue_reg[0][2]/NET0131 , \InstQueue_reg[0][3]/NET0131 , \InstQueue_reg[0][4]/NET0131 , \InstQueue_reg[0][5]/NET0131 , \InstQueue_reg[0][6]/NET0131 , \InstQueue_reg[0][7]/NET0131 , \InstQueue_reg[10][0]/NET0131 , \InstQueue_reg[10][1]/NET0131 , \InstQueue_reg[10][2]/NET0131 , \InstQueue_reg[10][3]/NET0131 , \InstQueue_reg[10][4]/NET0131 , \InstQueue_reg[10][5]/NET0131 , \InstQueue_reg[10][6]/NET0131 , \InstQueue_reg[10][7]/NET0131 , \InstQueue_reg[11][0]/NET0131 , \InstQueue_reg[11][1]/NET0131 , \InstQueue_reg[11][2]/NET0131 , \InstQueue_reg[11][3]/NET0131 , \InstQueue_reg[11][4]/NET0131 , \InstQueue_reg[11][5]/NET0131 , \InstQueue_reg[11][6]/NET0131 , \InstQueue_reg[11][7]/NET0131 , \InstQueue_reg[12][0]/NET0131 , \InstQueue_reg[12][1]/NET0131 , \InstQueue_reg[12][2]/NET0131 , \InstQueue_reg[12][3]/NET0131 , \InstQueue_reg[12][4]/NET0131 , \InstQueue_reg[12][5]/NET0131 , \InstQueue_reg[12][6]/NET0131 , \InstQueue_reg[12][7]/NET0131 , \InstQueue_reg[13][0]/NET0131 , \InstQueue_reg[13][1]/NET0131 , \InstQueue_reg[13][2]/NET0131 , \InstQueue_reg[13][3]/NET0131 , \InstQueue_reg[13][4]/NET0131 , \InstQueue_reg[13][5]/NET0131 , \InstQueue_reg[13][6]/NET0131 , \InstQueue_reg[13][7]/NET0131 , \InstQueue_reg[14][0]/NET0131 , \InstQueue_reg[14][1]/NET0131 , \InstQueue_reg[14][2]/NET0131 , \InstQueue_reg[14][3]/NET0131 , \InstQueue_reg[14][4]/NET0131 , \InstQueue_reg[14][5]/NET0131 , \InstQueue_reg[14][6]/NET0131 , \InstQueue_reg[14][7]/NET0131 , \InstQueue_reg[15][0]/NET0131 , \InstQueue_reg[15][1]/NET0131 , \InstQueue_reg[15][2]/NET0131 , \InstQueue_reg[15][3]/NET0131 , \InstQueue_reg[15][4]/NET0131 , \InstQueue_reg[15][5]/NET0131 , \InstQueue_reg[15][6]/NET0131 , \InstQueue_reg[15][7]/NET0131 , \InstQueue_reg[1][0]/NET0131 , \InstQueue_reg[1][1]/NET0131 , \InstQueue_reg[1][2]/NET0131 , \InstQueue_reg[1][3]/NET0131 , \InstQueue_reg[1][4]/NET0131 , \InstQueue_reg[1][5]/NET0131 , \InstQueue_reg[1][6]/NET0131 , \InstQueue_reg[1][7]/NET0131 , \InstQueue_reg[2][0]/NET0131 , \InstQueue_reg[2][1]/NET0131 , \InstQueue_reg[2][2]/NET0131 , \InstQueue_reg[2][3]/NET0131 , \InstQueue_reg[2][4]/NET0131 , \InstQueue_reg[2][5]/NET0131 , \InstQueue_reg[2][6]/NET0131 , \InstQueue_reg[2][7]/NET0131 , \InstQueue_reg[3][0]/NET0131 , \InstQueue_reg[3][1]/NET0131 , \InstQueue_reg[3][2]/NET0131 , \InstQueue_reg[3][3]/NET0131 , \InstQueue_reg[3][4]/NET0131 , \InstQueue_reg[3][5]/NET0131 , \InstQueue_reg[3][6]/NET0131 , \InstQueue_reg[3][7]/NET0131 , \InstQueue_reg[4][0]/NET0131 , \InstQueue_reg[4][1]/NET0131 , \InstQueue_reg[4][2]/NET0131 , \InstQueue_reg[4][3]/NET0131 , \InstQueue_reg[4][4]/NET0131 , \InstQueue_reg[4][5]/NET0131 , \InstQueue_reg[4][6]/NET0131 , \InstQueue_reg[4][7]/NET0131 , \InstQueue_reg[5][0]/NET0131 , \InstQueue_reg[5][1]/NET0131 , \InstQueue_reg[5][2]/NET0131 , \InstQueue_reg[5][3]/NET0131 , \InstQueue_reg[5][4]/NET0131 , \InstQueue_reg[5][5]/NET0131 , \InstQueue_reg[5][6]/NET0131 , \InstQueue_reg[5][7]/NET0131 , \InstQueue_reg[6][0]/NET0131 , \InstQueue_reg[6][1]/NET0131 , \InstQueue_reg[6][2]/NET0131 , \InstQueue_reg[6][3]/NET0131 , \InstQueue_reg[6][4]/NET0131 , \InstQueue_reg[6][5]/NET0131 , \InstQueue_reg[6][6]/NET0131 , \InstQueue_reg[6][7]/NET0131 , \InstQueue_reg[7][0]/NET0131 , \InstQueue_reg[7][1]/NET0131 , \InstQueue_reg[7][2]/NET0131 , \InstQueue_reg[7][3]/NET0131 , \InstQueue_reg[7][4]/NET0131 , \InstQueue_reg[7][5]/NET0131 , \InstQueue_reg[7][6]/NET0131 , \InstQueue_reg[7][7]/NET0131 , \InstQueue_reg[8][0]/NET0131 , \InstQueue_reg[8][1]/NET0131 , \InstQueue_reg[8][2]/NET0131 , \InstQueue_reg[8][3]/NET0131 , \InstQueue_reg[8][4]/NET0131 , \InstQueue_reg[8][5]/NET0131 , \InstQueue_reg[8][6]/NET0131 , \InstQueue_reg[8][7]/NET0131 , \InstQueue_reg[9][0]/NET0131 , \InstQueue_reg[9][1]/NET0131 , \InstQueue_reg[9][2]/NET0131 , \InstQueue_reg[9][3]/NET0131 , \InstQueue_reg[9][4]/NET0131 , \InstQueue_reg[9][5]/NET0131 , \InstQueue_reg[9][6]/NET0131 , \InstQueue_reg[9][7]/NET0131 , M_IO_n_pad, \MemoryFetch_reg/NET0131 , \More_reg/NET0131 , NA_n_pad, \PhyAddrPointer_reg[0]/NET0131 , \PhyAddrPointer_reg[10]/NET0131 , \PhyAddrPointer_reg[11]/NET0131 , \PhyAddrPointer_reg[12]/NET0131 , \PhyAddrPointer_reg[13]/NET0131 , \PhyAddrPointer_reg[14]/NET0131 , \PhyAddrPointer_reg[15]/NET0131 , \PhyAddrPointer_reg[16]/NET0131 , \PhyAddrPointer_reg[17]/NET0131 , \PhyAddrPointer_reg[18]/NET0131 , \PhyAddrPointer_reg[19]/NET0131 , \PhyAddrPointer_reg[1]/NET0131 , \PhyAddrPointer_reg[20]/NET0131 , \PhyAddrPointer_reg[21]/NET0131 , \PhyAddrPointer_reg[22]/NET0131 , \PhyAddrPointer_reg[23]/NET0131 , \PhyAddrPointer_reg[24]/NET0131 , \PhyAddrPointer_reg[25]/NET0131 , \PhyAddrPointer_reg[26]/NET0131 , \PhyAddrPointer_reg[27]/NET0131 , \PhyAddrPointer_reg[28]/NET0131 , \PhyAddrPointer_reg[29]/NET0131 , \PhyAddrPointer_reg[2]/NET0131 , \PhyAddrPointer_reg[30]/NET0131 , \PhyAddrPointer_reg[31]/NET0131 , \PhyAddrPointer_reg[3]/NET0131 , \PhyAddrPointer_reg[4]/NET0131 , \PhyAddrPointer_reg[5]/NET0131 , \PhyAddrPointer_reg[6]/NET0131 , \PhyAddrPointer_reg[7]/NET0131 , \PhyAddrPointer_reg[8]/NET0131 , \PhyAddrPointer_reg[9]/NET0131 , READY_n_pad, \ReadRequest_reg/NET0131 , \RequestPending_reg/NET0131 , \State2_reg[0]/NET0131 , \State2_reg[1]/NET0131 , \State2_reg[2]/NET0131 , \State2_reg[3]/NET0131 , \State_reg[0]/NET0131 , \State_reg[1]/NET0131 , \State_reg[2]/NET0131 , W_R_n_pad, \lWord_reg[0]/NET0131 , \lWord_reg[10]/NET0131 , \lWord_reg[11]/NET0131 , \lWord_reg[12]/NET0131 , \lWord_reg[13]/NET0131 , \lWord_reg[14]/NET0131 , \lWord_reg[15]/NET0131 , \lWord_reg[1]/NET0131 , \lWord_reg[2]/NET0131 , \lWord_reg[3]/NET0131 , \lWord_reg[4]/NET0131 , \lWord_reg[5]/NET0131 , \lWord_reg[6]/NET0131 , \lWord_reg[7]/NET0131 , \lWord_reg[8]/NET0131 , \lWord_reg[9]/NET0131 , \rEIP_reg[0]/NET0131 , \rEIP_reg[10]/NET0131 , \rEIP_reg[11]/NET0131 , \rEIP_reg[12]/NET0131 , \rEIP_reg[13]/NET0131 , \rEIP_reg[14]/NET0131 , \rEIP_reg[15]/NET0131 , \rEIP_reg[16]/NET0131 , \rEIP_reg[17]/NET0131 , \rEIP_reg[18]/NET0131 , \rEIP_reg[19]/NET0131 , \rEIP_reg[1]/NET0131 , \rEIP_reg[20]/NET0131 , \rEIP_reg[21]/NET0131 , \rEIP_reg[22]/NET0131 , \rEIP_reg[23]/NET0131 , \rEIP_reg[24]/NET0131 , \rEIP_reg[25]/NET0131 , \rEIP_reg[26]/NET0131 , \rEIP_reg[27]/NET0131 , \rEIP_reg[28]/NET0131 , \rEIP_reg[29]/NET0131 , \rEIP_reg[2]/NET0131 , \rEIP_reg[30]/NET0131 , \rEIP_reg[31]/NET0131 , \rEIP_reg[3]/NET0131 , \rEIP_reg[4]/NET0131 , \rEIP_reg[5]/NET0131 , \rEIP_reg[6]/NET0131 , \rEIP_reg[7]/NET0131 , \rEIP_reg[8]/NET0131 , \rEIP_reg[9]/NET0131 , \uWord_reg[0]/NET0131 , \uWord_reg[10]/NET0131 , \uWord_reg[11]/NET0131 , \uWord_reg[12]/NET0131 , \uWord_reg[13]/NET0131 , \uWord_reg[14]/NET0131 , \uWord_reg[1]/NET0131 , \uWord_reg[2]/NET0131 , \uWord_reg[3]/NET0131 , \uWord_reg[4]/NET0131 , \uWord_reg[5]/NET0131 , \uWord_reg[6]/NET0131 , \uWord_reg[7]/NET0131 , \uWord_reg[8]/NET0131 , \uWord_reg[9]/NET0131 , \_al_n0 , \_al_n1 , \g47521/_2_ , \g47523/_0_ , \g47526/_0_ , \g47529/_0_ , \g47533/_0_ , \g47540/_0_ , \g47551/_0_ , \g47552/_0_ , \g47553/_0_ , \g47563/_2_ , \g47566/_0_ , \g47567/_0_ , \g47568/_0_ , \g47569/_0_ , \g47583/_2_ , \g47584/_0_ , \g47585/_0_ , \g47589/_0_ , \g47602/_0_ , \g47603/_0_ , \g47604/_2_ , \g47605/_0_ , \g47606/_2_ , \g47609/_0_ , \g47611/_0_ , \g47631/_0_ , \g47632/_0_ , \g47633/_0_ , \g47635/_0_ , \g47636/_0_ , \g47637/_0_ , \g47638/_2_ , \g47643/_0_ , \g47665/_2_ , \g47666/_0_ , \g47667/_0_ , \g47670/_0_ , \g47672/_0_ , \g47677/_0_ , \g47678/_0_ , \g47706/_0_ , \g47711/_0_ , \g47717/_0_ , \g47718/_0_ , \g47721/_0_ , \g47722/_0_ , \g47751/_0_ , \g47755/_0_ , \g47756/_0_ , \g47757/_0_ , \g47759/_0_ , \g47789/_0_ , \g47793/_0_ , \g47797/_0_ , \g47798/_0_ , \g47799/_0_ , \g47802/_0_ , \g47804/_0_ , \g47807/_0_ , \g47809/_0_ , \g47862/_0_ , \g47863/_0_ , \g47864/_0_ , \g47869/_0_ , \g47870/_0_ , \g47924/_0_ , \g47925/_0_ , \g47926/_0_ , \g47927/_0_ , \g47928/_0_ , \g47930/_0_ , \g47932/_0_ , \g47933/_0_ , \g47934/_0_ , \g47935/_0_ , \g47936/_0_ , \g47937/_0_ , \g47938/_0_ , \g47939/_0_ , \g47940/_0_ , \g47941/_0_ , \g47957/_0_ , \g47970/_0_ , \g47973/_0_ , \g47975/_0_ , \g48058/_0_ , \g48059/_0_ , \g48060/_0_ , \g48061/_0_ , \g48062/_0_ , \g48064/_0_ , \g48065/_0_ , \g48066/_0_ , \g48067/_0_ , \g48068/_0_ , \g48069/_0_ , \g48070/_0_ , \g48071/_0_ , \g48072/_0_ , \g48073/_0_ , \g48074/_0_ , \g48087/_0_ , \g48110/_0_ , \g48117/_0_ , \g48118/_0_ , \g48119/_0_ , \g48120/_0_ , \g48121/_0_ , \g48122/_0_ , \g48124/_0_ , \g48125/_0_ , \g48126/_0_ , \g48127/_0_ , \g48128/_0_ , \g48129/_0_ , \g48130/_0_ , \g48131/_0_ , \g48132/_0_ , \g48133/_0_ , \g48134/_0_ , \g48168/_0_ , \g48169/_0_ , \g48170/_0_ , \g48171/_0_ , \g48172/_0_ , \g48173/_0_ , \g48174/_0_ , \g48175/_0_ , \g48177/_0_ , \g48178/_0_ , \g48179/_0_ , \g48180/_0_ , \g48181/_0_ , \g48182/_0_ , \g48183/_0_ , \g48184/_0_ , \g48185/_0_ , \g48186/_0_ , \g48187/_0_ , \g48188/_0_ , \g48189/_0_ , \g48192/_0_ , \g48193/_0_ , \g48194/_0_ , \g48195/_0_ , \g48196/_0_ , \g48197/_0_ , \g48198/_0_ , \g48199/_0_ , \g48200/_0_ , \g48201/_0_ , \g48202/_0_ , \g48203/_0_ , \g48213/_0_ , \g48214/_0_ , \g48215/_0_ , \g48216/_0_ , \g48217/_0_ , \g48218/_0_ , \g48219/_0_ , \g48220/_0_ , \g48221/_0_ , \g48222/_0_ , \g48223/_0_ , \g48224/_0_ , \g48225/_0_ , \g48226/_0_ , \g48227/_0_ , \g48228/_0_ , \g48229/_0_ , \g48230/_0_ , \g48231/_0_ , \g48232/_0_ , \g48234/_0_ , \g48236/_0_ , \g48237/_0_ , \g48238/_0_ , \g48239/_0_ , \g48240/_0_ , \g48241/_0_ , \g48243/_0_ , \g48244/_0_ , \g48245/_0_ , \g48246/_0_ , \g48263/_0_ , \g48270/_0_ , \g48273/_0_ , \g48276/_0_ , \g48277/_0_ , \g48370/_0_ , \g48377/_0_ , \g48391/_0_ , \g48423/_0_ , \g48428/_0_ , \g48429/_0_ , \g48431/_0_ , \g48433/_0_ , \g48434/_0_ , \g48435/_0_ , \g48436/_0_ , \g48437/_0_ , \g48438/_0_ , \g48439/_0_ , \g48440/_0_ , \g48441/_0_ , \g48442/_0_ , \g48443/_0_ , \g48610/_0_ , \g48634/_0_ , \g48635/_0_ , \g48636/_0_ , \g48637/_0_ , \g48638/_0_ , \g48639/_0_ , \g48640/_0_ , \g48642/_0_ , \g48643/_0_ , \g48644/_0_ , \g48645/_0_ , \g48646/_0_ , \g48647/_0_ , \g48648/_0_ , \g48649/_0_ , \g48650/_0_ , \g48651/_0_ , \g48652/_0_ , \g48653/_0_ , \g48654/_0_ , \g48655/_0_ , \g48656/_0_ , \g48657/_0_ , \g48658/_0_ , \g48659/_0_ , \g48660/_0_ , \g48662/_0_ , \g48663/_0_ , \g48664/_0_ , \g48665/_0_ , \g48666/_0_ , \g48667/_0_ , \g48668/_0_ , \g48669/_0_ , \g48750/_0_ , \g48753/_0_ , \g48756/_0_ , \g48759/_0_ , \g48763/_0_ , \g48766/_0_ , \g48769/_0_ , \g48772/_0_ , \g48775/_0_ , \g48778/_0_ , \g48781/_0_ , \g48785/_0_ , \g48789/_0_ , \g48792/_0_ , \g48796/_0_ , \g48799/_0_ , \g48937/_0_ , \g48958/_0_ , \g48959/_0_ , \g48964/_0_ , \g48965/_0_ , \g48966/_0_ , \g48967/_0_ , \g48968/_0_ , \g48969/_0_ , \g48970/_0_ , \g48971/_0_ , \g48972/_0_ , \g48973/_0_ , \g48974/_0_ , \g48975/_0_ , \g48976/_0_ , \g48977/_0_ , \g48978/_0_ , \g48979/_0_ , \g49/_0_ , \g49069/_0_ , \g49070/_0_ , \g49071/_0_ , \g49073/_0_ , \g49074/_0_ , \g49076/_0_ , \g49078/_0_ , \g49081/_0_ , \g49083/_0_ , \g49085/_0_ , \g49087/_0_ , \g49088/_0_ , \g49090/_0_ , \g49092/_0_ , \g49095/_0_ , \g49098/_0_ , \g49125/_0_ , \g49162/_0_ , \g49202/_0_ , \g49203/_0_ , \g49206/_0_ , \g49340/_0_ , \g49457/_0_ , \g49512/_0_ , \g49513/_0_ , \g49514/_0_ , \g49515/_0_ , \g49516/_0_ , \g49517/_0_ , \g49518/_0_ , \g49519/_0_ , \g49520/_0_ , \g49521/_0_ , \g49522/_0_ , \g49523/_0_ , \g49524/_0_ , \g49525/_0_ , \g49526/_0_ , \g49527/_0_ , \g49534/_0_ , \g49551/_0_ , \g49573/_0_ , \g49574/_0_ , \g49578/_0_ , \g49582/_0_ , \g49584/_0_ , \g49592/_0_ , \g49600/_0_ , \g49604/_0_ , \g49608/_0_ , \g49612/_0_ , \g49616/_0_ , \g49619/_0_ , \g49620/_0_ , \g49623/_0_ , \g49627/_0_ , \g49630/_0_ , \g49634/_0_ , \g49635/_0_ , \g49639/_0_ , \g49645/_0_ , \g49744/_0_ , \g49766/_0_ , \g50098/_0_ , \g50124/_0_ , \g50195/_0_ , \g50198/_0_ , \g50201/_0_ , \g50203/_0_ , \g50205/_0_ , \g50207/_0_ , \g50209/_0_ , \g50213/_0_ , \g50222/_0_ , \g50228/_0_ , \g50231/_0_ , \g50237/_0_ , \g50240/_0_ , \g50335/_0_ , \g50477/_0_ , \g50478/_0_ , \g50671/_0_ , \g50757/_0_ , \g50938/_0_ , \g50998/_0_ , \g51008/_0_ , \g51579/_0_ , \g51637/_0_ , \g51662/_0_ , \g52424/_0_ , \g53184/_0_ , \g53206/_0_ , \g53270/_0_ , \g53730/_0_ , \g53754/_0_ , \g54176/_0_ , \g54214/_0_ , \g54229/_0_ , \g54392/_0_ , \g54400/_0_ , \g54415/_0_ , \g54421/_0_ , \g54604/_0_ , \g54607/_0_ , \g54638/_0_ , \g54694/_0_ , \g54759/_0_ , \g55607/_0_ , \g55863/_1_ , \g56073/_0_ , \g56292/_0_ , \g56320/_0_ , \g56527/_0_ , \g56531/_0_ , \g56533/_0_ , \g56562/_0_ , \g56615/_0_ , \g56720/_0_ , \g57044/_0_ , \g60635/_1_ , \g62873/_0_ , \g62886/_0_ , \g63001/_0_ , \g63101/_0_ , \g63129/_0_ , \g63198/_0_ , \g63449/_0_ , \g63471/_0_ , \g63493/_0_ , \g63626/_0_ , \g63688/_0_ , \g63800/_0_ , \g63934/_0_ , \g63954/_0_ , \g64060/_0_ , \g64375/_0_ , \g65/_0_ , \g67/_0_ );
	input ADS_n_pad ;
	input \Address[0]_pad  ;
	input \Address[10]_pad  ;
	input \Address[11]_pad  ;
	input \Address[12]_pad  ;
	input \Address[13]_pad  ;
	input \Address[14]_pad  ;
	input \Address[15]_pad  ;
	input \Address[16]_pad  ;
	input \Address[17]_pad  ;
	input \Address[18]_pad  ;
	input \Address[19]_pad  ;
	input \Address[1]_pad  ;
	input \Address[20]_pad  ;
	input \Address[21]_pad  ;
	input \Address[22]_pad  ;
	input \Address[23]_pad  ;
	input \Address[24]_pad  ;
	input \Address[25]_pad  ;
	input \Address[26]_pad  ;
	input \Address[27]_pad  ;
	input \Address[28]_pad  ;
	input \Address[29]_pad  ;
	input \Address[2]_pad  ;
	input \Address[3]_pad  ;
	input \Address[4]_pad  ;
	input \Address[5]_pad  ;
	input \Address[6]_pad  ;
	input \Address[7]_pad  ;
	input \Address[8]_pad  ;
	input \Address[9]_pad  ;
	input \BE_n[0]_pad  ;
	input \BE_n[1]_pad  ;
	input \BE_n[2]_pad  ;
	input \BE_n[3]_pad  ;
	input \BS16_n_pad  ;
	input \ByteEnable_reg[0]/NET0131  ;
	input \ByteEnable_reg[1]/NET0131  ;
	input \ByteEnable_reg[2]/NET0131  ;
	input \ByteEnable_reg[3]/NET0131  ;
	input \CodeFetch_reg/NET0131  ;
	input D_C_n_pad ;
	input \DataWidth_reg[0]/NET0131  ;
	input \DataWidth_reg[1]/NET0131  ;
	input \Datai[0]_pad  ;
	input \Datai[10]_pad  ;
	input \Datai[11]_pad  ;
	input \Datai[12]_pad  ;
	input \Datai[13]_pad  ;
	input \Datai[14]_pad  ;
	input \Datai[15]_pad  ;
	input \Datai[16]_pad  ;
	input \Datai[17]_pad  ;
	input \Datai[18]_pad  ;
	input \Datai[19]_pad  ;
	input \Datai[1]_pad  ;
	input \Datai[20]_pad  ;
	input \Datai[21]_pad  ;
	input \Datai[22]_pad  ;
	input \Datai[23]_pad  ;
	input \Datai[24]_pad  ;
	input \Datai[25]_pad  ;
	input \Datai[26]_pad  ;
	input \Datai[27]_pad  ;
	input \Datai[28]_pad  ;
	input \Datai[29]_pad  ;
	input \Datai[2]_pad  ;
	input \Datai[30]_pad  ;
	input \Datai[31]_pad  ;
	input \Datai[3]_pad  ;
	input \Datai[4]_pad  ;
	input \Datai[5]_pad  ;
	input \Datai[6]_pad  ;
	input \Datai[7]_pad  ;
	input \Datai[8]_pad  ;
	input \Datai[9]_pad  ;
	input \Datao[0]_pad  ;
	input \Datao[10]_pad  ;
	input \Datao[11]_pad  ;
	input \Datao[12]_pad  ;
	input \Datao[13]_pad  ;
	input \Datao[14]_pad  ;
	input \Datao[15]_pad  ;
	input \Datao[16]_pad  ;
	input \Datao[17]_pad  ;
	input \Datao[18]_pad  ;
	input \Datao[19]_pad  ;
	input \Datao[1]_pad  ;
	input \Datao[20]_pad  ;
	input \Datao[21]_pad  ;
	input \Datao[23]_pad  ;
	input \Datao[24]_pad  ;
	input \Datao[25]_pad  ;
	input \Datao[26]_pad  ;
	input \Datao[27]_pad  ;
	input \Datao[28]_pad  ;
	input \Datao[29]_pad  ;
	input \Datao[2]_pad  ;
	input \Datao[30]_pad  ;
	input \Datao[3]_pad  ;
	input \Datao[4]_pad  ;
	input \Datao[5]_pad  ;
	input \Datao[6]_pad  ;
	input \Datao[7]_pad  ;
	input \Datao[8]_pad  ;
	input \Datao[9]_pad  ;
	input \Datao_reg[22]/NET0131  ;
	input \EAX_reg[0]/NET0131  ;
	input \EAX_reg[10]/NET0131  ;
	input \EAX_reg[11]/NET0131  ;
	input \EAX_reg[12]/NET0131  ;
	input \EAX_reg[13]/NET0131  ;
	input \EAX_reg[14]/NET0131  ;
	input \EAX_reg[15]/NET0131  ;
	input \EAX_reg[16]/NET0131  ;
	input \EAX_reg[17]/NET0131  ;
	input \EAX_reg[18]/NET0131  ;
	input \EAX_reg[19]/NET0131  ;
	input \EAX_reg[1]/NET0131  ;
	input \EAX_reg[20]/NET0131  ;
	input \EAX_reg[21]/NET0131  ;
	input \EAX_reg[22]/NET0131  ;
	input \EAX_reg[23]/NET0131  ;
	input \EAX_reg[24]/NET0131  ;
	input \EAX_reg[25]/NET0131  ;
	input \EAX_reg[26]/NET0131  ;
	input \EAX_reg[27]/NET0131  ;
	input \EAX_reg[28]/NET0131  ;
	input \EAX_reg[29]/NET0131  ;
	input \EAX_reg[2]/NET0131  ;
	input \EAX_reg[30]/NET0131  ;
	input \EAX_reg[31]/NET0131  ;
	input \EAX_reg[3]/NET0131  ;
	input \EAX_reg[4]/NET0131  ;
	input \EAX_reg[5]/NET0131  ;
	input \EAX_reg[6]/NET0131  ;
	input \EAX_reg[7]/NET0131  ;
	input \EAX_reg[8]/NET0131  ;
	input \EAX_reg[9]/NET0131  ;
	input \EBX_reg[0]/NET0131  ;
	input \EBX_reg[10]/NET0131  ;
	input \EBX_reg[11]/NET0131  ;
	input \EBX_reg[12]/NET0131  ;
	input \EBX_reg[13]/NET0131  ;
	input \EBX_reg[14]/NET0131  ;
	input \EBX_reg[15]/NET0131  ;
	input \EBX_reg[16]/NET0131  ;
	input \EBX_reg[17]/NET0131  ;
	input \EBX_reg[18]/NET0131  ;
	input \EBX_reg[19]/NET0131  ;
	input \EBX_reg[1]/NET0131  ;
	input \EBX_reg[20]/NET0131  ;
	input \EBX_reg[21]/NET0131  ;
	input \EBX_reg[22]/NET0131  ;
	input \EBX_reg[23]/NET0131  ;
	input \EBX_reg[24]/NET0131  ;
	input \EBX_reg[25]/NET0131  ;
	input \EBX_reg[26]/NET0131  ;
	input \EBX_reg[27]/NET0131  ;
	input \EBX_reg[28]/NET0131  ;
	input \EBX_reg[29]/NET0131  ;
	input \EBX_reg[2]/NET0131  ;
	input \EBX_reg[30]/NET0131  ;
	input \EBX_reg[31]/NET0131  ;
	input \EBX_reg[3]/NET0131  ;
	input \EBX_reg[4]/NET0131  ;
	input \EBX_reg[5]/NET0131  ;
	input \EBX_reg[6]/NET0131  ;
	input \EBX_reg[7]/NET0131  ;
	input \EBX_reg[8]/NET0131  ;
	input \EBX_reg[9]/NET0131  ;
	input \Flush_reg/NET0131  ;
	input HOLD_pad ;
	input \InstAddrPointer_reg[0]/NET0131  ;
	input \InstAddrPointer_reg[10]/NET0131  ;
	input \InstAddrPointer_reg[11]/NET0131  ;
	input \InstAddrPointer_reg[12]/NET0131  ;
	input \InstAddrPointer_reg[13]/NET0131  ;
	input \InstAddrPointer_reg[14]/NET0131  ;
	input \InstAddrPointer_reg[15]/NET0131  ;
	input \InstAddrPointer_reg[16]/NET0131  ;
	input \InstAddrPointer_reg[17]/NET0131  ;
	input \InstAddrPointer_reg[18]/NET0131  ;
	input \InstAddrPointer_reg[19]/NET0131  ;
	input \InstAddrPointer_reg[1]/NET0131  ;
	input \InstAddrPointer_reg[20]/NET0131  ;
	input \InstAddrPointer_reg[21]/NET0131  ;
	input \InstAddrPointer_reg[22]/NET0131  ;
	input \InstAddrPointer_reg[23]/NET0131  ;
	input \InstAddrPointer_reg[24]/NET0131  ;
	input \InstAddrPointer_reg[25]/NET0131  ;
	input \InstAddrPointer_reg[26]/NET0131  ;
	input \InstAddrPointer_reg[27]/NET0131  ;
	input \InstAddrPointer_reg[28]/NET0131  ;
	input \InstAddrPointer_reg[29]/NET0131  ;
	input \InstAddrPointer_reg[2]/NET0131  ;
	input \InstAddrPointer_reg[30]/NET0131  ;
	input \InstAddrPointer_reg[31]/NET0131  ;
	input \InstAddrPointer_reg[3]/NET0131  ;
	input \InstAddrPointer_reg[4]/NET0131  ;
	input \InstAddrPointer_reg[5]/NET0131  ;
	input \InstAddrPointer_reg[6]/NET0131  ;
	input \InstAddrPointer_reg[7]/NET0131  ;
	input \InstAddrPointer_reg[8]/NET0131  ;
	input \InstAddrPointer_reg[9]/NET0131  ;
	input \InstQueueRd_Addr_reg[0]/NET0131  ;
	input \InstQueueRd_Addr_reg[1]/NET0131  ;
	input \InstQueueRd_Addr_reg[2]/NET0131  ;
	input \InstQueueRd_Addr_reg[3]/NET0131  ;
	input \InstQueueWr_Addr_reg[0]/NET0131  ;
	input \InstQueueWr_Addr_reg[1]/NET0131  ;
	input \InstQueueWr_Addr_reg[2]/NET0131  ;
	input \InstQueueWr_Addr_reg[3]/NET0131  ;
	input \InstQueue_reg[0][0]/NET0131  ;
	input \InstQueue_reg[0][1]/NET0131  ;
	input \InstQueue_reg[0][2]/NET0131  ;
	input \InstQueue_reg[0][3]/NET0131  ;
	input \InstQueue_reg[0][4]/NET0131  ;
	input \InstQueue_reg[0][5]/NET0131  ;
	input \InstQueue_reg[0][6]/NET0131  ;
	input \InstQueue_reg[0][7]/NET0131  ;
	input \InstQueue_reg[10][0]/NET0131  ;
	input \InstQueue_reg[10][1]/NET0131  ;
	input \InstQueue_reg[10][2]/NET0131  ;
	input \InstQueue_reg[10][3]/NET0131  ;
	input \InstQueue_reg[10][4]/NET0131  ;
	input \InstQueue_reg[10][5]/NET0131  ;
	input \InstQueue_reg[10][6]/NET0131  ;
	input \InstQueue_reg[10][7]/NET0131  ;
	input \InstQueue_reg[11][0]/NET0131  ;
	input \InstQueue_reg[11][1]/NET0131  ;
	input \InstQueue_reg[11][2]/NET0131  ;
	input \InstQueue_reg[11][3]/NET0131  ;
	input \InstQueue_reg[11][4]/NET0131  ;
	input \InstQueue_reg[11][5]/NET0131  ;
	input \InstQueue_reg[11][6]/NET0131  ;
	input \InstQueue_reg[11][7]/NET0131  ;
	input \InstQueue_reg[12][0]/NET0131  ;
	input \InstQueue_reg[12][1]/NET0131  ;
	input \InstQueue_reg[12][2]/NET0131  ;
	input \InstQueue_reg[12][3]/NET0131  ;
	input \InstQueue_reg[12][4]/NET0131  ;
	input \InstQueue_reg[12][5]/NET0131  ;
	input \InstQueue_reg[12][6]/NET0131  ;
	input \InstQueue_reg[12][7]/NET0131  ;
	input \InstQueue_reg[13][0]/NET0131  ;
	input \InstQueue_reg[13][1]/NET0131  ;
	input \InstQueue_reg[13][2]/NET0131  ;
	input \InstQueue_reg[13][3]/NET0131  ;
	input \InstQueue_reg[13][4]/NET0131  ;
	input \InstQueue_reg[13][5]/NET0131  ;
	input \InstQueue_reg[13][6]/NET0131  ;
	input \InstQueue_reg[13][7]/NET0131  ;
	input \InstQueue_reg[14][0]/NET0131  ;
	input \InstQueue_reg[14][1]/NET0131  ;
	input \InstQueue_reg[14][2]/NET0131  ;
	input \InstQueue_reg[14][3]/NET0131  ;
	input \InstQueue_reg[14][4]/NET0131  ;
	input \InstQueue_reg[14][5]/NET0131  ;
	input \InstQueue_reg[14][6]/NET0131  ;
	input \InstQueue_reg[14][7]/NET0131  ;
	input \InstQueue_reg[15][0]/NET0131  ;
	input \InstQueue_reg[15][1]/NET0131  ;
	input \InstQueue_reg[15][2]/NET0131  ;
	input \InstQueue_reg[15][3]/NET0131  ;
	input \InstQueue_reg[15][4]/NET0131  ;
	input \InstQueue_reg[15][5]/NET0131  ;
	input \InstQueue_reg[15][6]/NET0131  ;
	input \InstQueue_reg[15][7]/NET0131  ;
	input \InstQueue_reg[1][0]/NET0131  ;
	input \InstQueue_reg[1][1]/NET0131  ;
	input \InstQueue_reg[1][2]/NET0131  ;
	input \InstQueue_reg[1][3]/NET0131  ;
	input \InstQueue_reg[1][4]/NET0131  ;
	input \InstQueue_reg[1][5]/NET0131  ;
	input \InstQueue_reg[1][6]/NET0131  ;
	input \InstQueue_reg[1][7]/NET0131  ;
	input \InstQueue_reg[2][0]/NET0131  ;
	input \InstQueue_reg[2][1]/NET0131  ;
	input \InstQueue_reg[2][2]/NET0131  ;
	input \InstQueue_reg[2][3]/NET0131  ;
	input \InstQueue_reg[2][4]/NET0131  ;
	input \InstQueue_reg[2][5]/NET0131  ;
	input \InstQueue_reg[2][6]/NET0131  ;
	input \InstQueue_reg[2][7]/NET0131  ;
	input \InstQueue_reg[3][0]/NET0131  ;
	input \InstQueue_reg[3][1]/NET0131  ;
	input \InstQueue_reg[3][2]/NET0131  ;
	input \InstQueue_reg[3][3]/NET0131  ;
	input \InstQueue_reg[3][4]/NET0131  ;
	input \InstQueue_reg[3][5]/NET0131  ;
	input \InstQueue_reg[3][6]/NET0131  ;
	input \InstQueue_reg[3][7]/NET0131  ;
	input \InstQueue_reg[4][0]/NET0131  ;
	input \InstQueue_reg[4][1]/NET0131  ;
	input \InstQueue_reg[4][2]/NET0131  ;
	input \InstQueue_reg[4][3]/NET0131  ;
	input \InstQueue_reg[4][4]/NET0131  ;
	input \InstQueue_reg[4][5]/NET0131  ;
	input \InstQueue_reg[4][6]/NET0131  ;
	input \InstQueue_reg[4][7]/NET0131  ;
	input \InstQueue_reg[5][0]/NET0131  ;
	input \InstQueue_reg[5][1]/NET0131  ;
	input \InstQueue_reg[5][2]/NET0131  ;
	input \InstQueue_reg[5][3]/NET0131  ;
	input \InstQueue_reg[5][4]/NET0131  ;
	input \InstQueue_reg[5][5]/NET0131  ;
	input \InstQueue_reg[5][6]/NET0131  ;
	input \InstQueue_reg[5][7]/NET0131  ;
	input \InstQueue_reg[6][0]/NET0131  ;
	input \InstQueue_reg[6][1]/NET0131  ;
	input \InstQueue_reg[6][2]/NET0131  ;
	input \InstQueue_reg[6][3]/NET0131  ;
	input \InstQueue_reg[6][4]/NET0131  ;
	input \InstQueue_reg[6][5]/NET0131  ;
	input \InstQueue_reg[6][6]/NET0131  ;
	input \InstQueue_reg[6][7]/NET0131  ;
	input \InstQueue_reg[7][0]/NET0131  ;
	input \InstQueue_reg[7][1]/NET0131  ;
	input \InstQueue_reg[7][2]/NET0131  ;
	input \InstQueue_reg[7][3]/NET0131  ;
	input \InstQueue_reg[7][4]/NET0131  ;
	input \InstQueue_reg[7][5]/NET0131  ;
	input \InstQueue_reg[7][6]/NET0131  ;
	input \InstQueue_reg[7][7]/NET0131  ;
	input \InstQueue_reg[8][0]/NET0131  ;
	input \InstQueue_reg[8][1]/NET0131  ;
	input \InstQueue_reg[8][2]/NET0131  ;
	input \InstQueue_reg[8][3]/NET0131  ;
	input \InstQueue_reg[8][4]/NET0131  ;
	input \InstQueue_reg[8][5]/NET0131  ;
	input \InstQueue_reg[8][6]/NET0131  ;
	input \InstQueue_reg[8][7]/NET0131  ;
	input \InstQueue_reg[9][0]/NET0131  ;
	input \InstQueue_reg[9][1]/NET0131  ;
	input \InstQueue_reg[9][2]/NET0131  ;
	input \InstQueue_reg[9][3]/NET0131  ;
	input \InstQueue_reg[9][4]/NET0131  ;
	input \InstQueue_reg[9][5]/NET0131  ;
	input \InstQueue_reg[9][6]/NET0131  ;
	input \InstQueue_reg[9][7]/NET0131  ;
	input M_IO_n_pad ;
	input \MemoryFetch_reg/NET0131  ;
	input \More_reg/NET0131  ;
	input NA_n_pad ;
	input \PhyAddrPointer_reg[0]/NET0131  ;
	input \PhyAddrPointer_reg[10]/NET0131  ;
	input \PhyAddrPointer_reg[11]/NET0131  ;
	input \PhyAddrPointer_reg[12]/NET0131  ;
	input \PhyAddrPointer_reg[13]/NET0131  ;
	input \PhyAddrPointer_reg[14]/NET0131  ;
	input \PhyAddrPointer_reg[15]/NET0131  ;
	input \PhyAddrPointer_reg[16]/NET0131  ;
	input \PhyAddrPointer_reg[17]/NET0131  ;
	input \PhyAddrPointer_reg[18]/NET0131  ;
	input \PhyAddrPointer_reg[19]/NET0131  ;
	input \PhyAddrPointer_reg[1]/NET0131  ;
	input \PhyAddrPointer_reg[20]/NET0131  ;
	input \PhyAddrPointer_reg[21]/NET0131  ;
	input \PhyAddrPointer_reg[22]/NET0131  ;
	input \PhyAddrPointer_reg[23]/NET0131  ;
	input \PhyAddrPointer_reg[24]/NET0131  ;
	input \PhyAddrPointer_reg[25]/NET0131  ;
	input \PhyAddrPointer_reg[26]/NET0131  ;
	input \PhyAddrPointer_reg[27]/NET0131  ;
	input \PhyAddrPointer_reg[28]/NET0131  ;
	input \PhyAddrPointer_reg[29]/NET0131  ;
	input \PhyAddrPointer_reg[2]/NET0131  ;
	input \PhyAddrPointer_reg[30]/NET0131  ;
	input \PhyAddrPointer_reg[31]/NET0131  ;
	input \PhyAddrPointer_reg[3]/NET0131  ;
	input \PhyAddrPointer_reg[4]/NET0131  ;
	input \PhyAddrPointer_reg[5]/NET0131  ;
	input \PhyAddrPointer_reg[6]/NET0131  ;
	input \PhyAddrPointer_reg[7]/NET0131  ;
	input \PhyAddrPointer_reg[8]/NET0131  ;
	input \PhyAddrPointer_reg[9]/NET0131  ;
	input READY_n_pad ;
	input \ReadRequest_reg/NET0131  ;
	input \RequestPending_reg/NET0131  ;
	input \State2_reg[0]/NET0131  ;
	input \State2_reg[1]/NET0131  ;
	input \State2_reg[2]/NET0131  ;
	input \State2_reg[3]/NET0131  ;
	input \State_reg[0]/NET0131  ;
	input \State_reg[1]/NET0131  ;
	input \State_reg[2]/NET0131  ;
	input W_R_n_pad ;
	input \lWord_reg[0]/NET0131  ;
	input \lWord_reg[10]/NET0131  ;
	input \lWord_reg[11]/NET0131  ;
	input \lWord_reg[12]/NET0131  ;
	input \lWord_reg[13]/NET0131  ;
	input \lWord_reg[14]/NET0131  ;
	input \lWord_reg[15]/NET0131  ;
	input \lWord_reg[1]/NET0131  ;
	input \lWord_reg[2]/NET0131  ;
	input \lWord_reg[3]/NET0131  ;
	input \lWord_reg[4]/NET0131  ;
	input \lWord_reg[5]/NET0131  ;
	input \lWord_reg[6]/NET0131  ;
	input \lWord_reg[7]/NET0131  ;
	input \lWord_reg[8]/NET0131  ;
	input \lWord_reg[9]/NET0131  ;
	input \rEIP_reg[0]/NET0131  ;
	input \rEIP_reg[10]/NET0131  ;
	input \rEIP_reg[11]/NET0131  ;
	input \rEIP_reg[12]/NET0131  ;
	input \rEIP_reg[13]/NET0131  ;
	input \rEIP_reg[14]/NET0131  ;
	input \rEIP_reg[15]/NET0131  ;
	input \rEIP_reg[16]/NET0131  ;
	input \rEIP_reg[17]/NET0131  ;
	input \rEIP_reg[18]/NET0131  ;
	input \rEIP_reg[19]/NET0131  ;
	input \rEIP_reg[1]/NET0131  ;
	input \rEIP_reg[20]/NET0131  ;
	input \rEIP_reg[21]/NET0131  ;
	input \rEIP_reg[22]/NET0131  ;
	input \rEIP_reg[23]/NET0131  ;
	input \rEIP_reg[24]/NET0131  ;
	input \rEIP_reg[25]/NET0131  ;
	input \rEIP_reg[26]/NET0131  ;
	input \rEIP_reg[27]/NET0131  ;
	input \rEIP_reg[28]/NET0131  ;
	input \rEIP_reg[29]/NET0131  ;
	input \rEIP_reg[2]/NET0131  ;
	input \rEIP_reg[30]/NET0131  ;
	input \rEIP_reg[31]/NET0131  ;
	input \rEIP_reg[3]/NET0131  ;
	input \rEIP_reg[4]/NET0131  ;
	input \rEIP_reg[5]/NET0131  ;
	input \rEIP_reg[6]/NET0131  ;
	input \rEIP_reg[7]/NET0131  ;
	input \rEIP_reg[8]/NET0131  ;
	input \rEIP_reg[9]/NET0131  ;
	input \uWord_reg[0]/NET0131  ;
	input \uWord_reg[10]/NET0131  ;
	input \uWord_reg[11]/NET0131  ;
	input \uWord_reg[12]/NET0131  ;
	input \uWord_reg[13]/NET0131  ;
	input \uWord_reg[14]/NET0131  ;
	input \uWord_reg[1]/NET0131  ;
	input \uWord_reg[2]/NET0131  ;
	input \uWord_reg[3]/NET0131  ;
	input \uWord_reg[4]/NET0131  ;
	input \uWord_reg[5]/NET0131  ;
	input \uWord_reg[6]/NET0131  ;
	input \uWord_reg[7]/NET0131  ;
	input \uWord_reg[8]/NET0131  ;
	input \uWord_reg[9]/NET0131  ;
	output \_al_n0  ;
	output \_al_n1  ;
	output \g47521/_2_  ;
	output \g47523/_0_  ;
	output \g47526/_0_  ;
	output \g47529/_0_  ;
	output \g47533/_0_  ;
	output \g47540/_0_  ;
	output \g47551/_0_  ;
	output \g47552/_0_  ;
	output \g47553/_0_  ;
	output \g47563/_2_  ;
	output \g47566/_0_  ;
	output \g47567/_0_  ;
	output \g47568/_0_  ;
	output \g47569/_0_  ;
	output \g47583/_2_  ;
	output \g47584/_0_  ;
	output \g47585/_0_  ;
	output \g47589/_0_  ;
	output \g47602/_0_  ;
	output \g47603/_0_  ;
	output \g47604/_2_  ;
	output \g47605/_0_  ;
	output \g47606/_2_  ;
	output \g47609/_0_  ;
	output \g47611/_0_  ;
	output \g47631/_0_  ;
	output \g47632/_0_  ;
	output \g47633/_0_  ;
	output \g47635/_0_  ;
	output \g47636/_0_  ;
	output \g47637/_0_  ;
	output \g47638/_2_  ;
	output \g47643/_0_  ;
	output \g47665/_2_  ;
	output \g47666/_0_  ;
	output \g47667/_0_  ;
	output \g47670/_0_  ;
	output \g47672/_0_  ;
	output \g47677/_0_  ;
	output \g47678/_0_  ;
	output \g47706/_0_  ;
	output \g47711/_0_  ;
	output \g47717/_0_  ;
	output \g47718/_0_  ;
	output \g47721/_0_  ;
	output \g47722/_0_  ;
	output \g47751/_0_  ;
	output \g47755/_0_  ;
	output \g47756/_0_  ;
	output \g47757/_0_  ;
	output \g47759/_0_  ;
	output \g47789/_0_  ;
	output \g47793/_0_  ;
	output \g47797/_0_  ;
	output \g47798/_0_  ;
	output \g47799/_0_  ;
	output \g47802/_0_  ;
	output \g47804/_0_  ;
	output \g47807/_0_  ;
	output \g47809/_0_  ;
	output \g47862/_0_  ;
	output \g47863/_0_  ;
	output \g47864/_0_  ;
	output \g47869/_0_  ;
	output \g47870/_0_  ;
	output \g47924/_0_  ;
	output \g47925/_0_  ;
	output \g47926/_0_  ;
	output \g47927/_0_  ;
	output \g47928/_0_  ;
	output \g47930/_0_  ;
	output \g47932/_0_  ;
	output \g47933/_0_  ;
	output \g47934/_0_  ;
	output \g47935/_0_  ;
	output \g47936/_0_  ;
	output \g47937/_0_  ;
	output \g47938/_0_  ;
	output \g47939/_0_  ;
	output \g47940/_0_  ;
	output \g47941/_0_  ;
	output \g47957/_0_  ;
	output \g47970/_0_  ;
	output \g47973/_0_  ;
	output \g47975/_0_  ;
	output \g48058/_0_  ;
	output \g48059/_0_  ;
	output \g48060/_0_  ;
	output \g48061/_0_  ;
	output \g48062/_0_  ;
	output \g48064/_0_  ;
	output \g48065/_0_  ;
	output \g48066/_0_  ;
	output \g48067/_0_  ;
	output \g48068/_0_  ;
	output \g48069/_0_  ;
	output \g48070/_0_  ;
	output \g48071/_0_  ;
	output \g48072/_0_  ;
	output \g48073/_0_  ;
	output \g48074/_0_  ;
	output \g48087/_0_  ;
	output \g48110/_0_  ;
	output \g48117/_0_  ;
	output \g48118/_0_  ;
	output \g48119/_0_  ;
	output \g48120/_0_  ;
	output \g48121/_0_  ;
	output \g48122/_0_  ;
	output \g48124/_0_  ;
	output \g48125/_0_  ;
	output \g48126/_0_  ;
	output \g48127/_0_  ;
	output \g48128/_0_  ;
	output \g48129/_0_  ;
	output \g48130/_0_  ;
	output \g48131/_0_  ;
	output \g48132/_0_  ;
	output \g48133/_0_  ;
	output \g48134/_0_  ;
	output \g48168/_0_  ;
	output \g48169/_0_  ;
	output \g48170/_0_  ;
	output \g48171/_0_  ;
	output \g48172/_0_  ;
	output \g48173/_0_  ;
	output \g48174/_0_  ;
	output \g48175/_0_  ;
	output \g48177/_0_  ;
	output \g48178/_0_  ;
	output \g48179/_0_  ;
	output \g48180/_0_  ;
	output \g48181/_0_  ;
	output \g48182/_0_  ;
	output \g48183/_0_  ;
	output \g48184/_0_  ;
	output \g48185/_0_  ;
	output \g48186/_0_  ;
	output \g48187/_0_  ;
	output \g48188/_0_  ;
	output \g48189/_0_  ;
	output \g48192/_0_  ;
	output \g48193/_0_  ;
	output \g48194/_0_  ;
	output \g48195/_0_  ;
	output \g48196/_0_  ;
	output \g48197/_0_  ;
	output \g48198/_0_  ;
	output \g48199/_0_  ;
	output \g48200/_0_  ;
	output \g48201/_0_  ;
	output \g48202/_0_  ;
	output \g48203/_0_  ;
	output \g48213/_0_  ;
	output \g48214/_0_  ;
	output \g48215/_0_  ;
	output \g48216/_0_  ;
	output \g48217/_0_  ;
	output \g48218/_0_  ;
	output \g48219/_0_  ;
	output \g48220/_0_  ;
	output \g48221/_0_  ;
	output \g48222/_0_  ;
	output \g48223/_0_  ;
	output \g48224/_0_  ;
	output \g48225/_0_  ;
	output \g48226/_0_  ;
	output \g48227/_0_  ;
	output \g48228/_0_  ;
	output \g48229/_0_  ;
	output \g48230/_0_  ;
	output \g48231/_0_  ;
	output \g48232/_0_  ;
	output \g48234/_0_  ;
	output \g48236/_0_  ;
	output \g48237/_0_  ;
	output \g48238/_0_  ;
	output \g48239/_0_  ;
	output \g48240/_0_  ;
	output \g48241/_0_  ;
	output \g48243/_0_  ;
	output \g48244/_0_  ;
	output \g48245/_0_  ;
	output \g48246/_0_  ;
	output \g48263/_0_  ;
	output \g48270/_0_  ;
	output \g48273/_0_  ;
	output \g48276/_0_  ;
	output \g48277/_0_  ;
	output \g48370/_0_  ;
	output \g48377/_0_  ;
	output \g48391/_0_  ;
	output \g48423/_0_  ;
	output \g48428/_0_  ;
	output \g48429/_0_  ;
	output \g48431/_0_  ;
	output \g48433/_0_  ;
	output \g48434/_0_  ;
	output \g48435/_0_  ;
	output \g48436/_0_  ;
	output \g48437/_0_  ;
	output \g48438/_0_  ;
	output \g48439/_0_  ;
	output \g48440/_0_  ;
	output \g48441/_0_  ;
	output \g48442/_0_  ;
	output \g48443/_0_  ;
	output \g48610/_0_  ;
	output \g48634/_0_  ;
	output \g48635/_0_  ;
	output \g48636/_0_  ;
	output \g48637/_0_  ;
	output \g48638/_0_  ;
	output \g48639/_0_  ;
	output \g48640/_0_  ;
	output \g48642/_0_  ;
	output \g48643/_0_  ;
	output \g48644/_0_  ;
	output \g48645/_0_  ;
	output \g48646/_0_  ;
	output \g48647/_0_  ;
	output \g48648/_0_  ;
	output \g48649/_0_  ;
	output \g48650/_0_  ;
	output \g48651/_0_  ;
	output \g48652/_0_  ;
	output \g48653/_0_  ;
	output \g48654/_0_  ;
	output \g48655/_0_  ;
	output \g48656/_0_  ;
	output \g48657/_0_  ;
	output \g48658/_0_  ;
	output \g48659/_0_  ;
	output \g48660/_0_  ;
	output \g48662/_0_  ;
	output \g48663/_0_  ;
	output \g48664/_0_  ;
	output \g48665/_0_  ;
	output \g48666/_0_  ;
	output \g48667/_0_  ;
	output \g48668/_0_  ;
	output \g48669/_0_  ;
	output \g48750/_0_  ;
	output \g48753/_0_  ;
	output \g48756/_0_  ;
	output \g48759/_0_  ;
	output \g48763/_0_  ;
	output \g48766/_0_  ;
	output \g48769/_0_  ;
	output \g48772/_0_  ;
	output \g48775/_0_  ;
	output \g48778/_0_  ;
	output \g48781/_0_  ;
	output \g48785/_0_  ;
	output \g48789/_0_  ;
	output \g48792/_0_  ;
	output \g48796/_0_  ;
	output \g48799/_0_  ;
	output \g48937/_0_  ;
	output \g48958/_0_  ;
	output \g48959/_0_  ;
	output \g48964/_0_  ;
	output \g48965/_0_  ;
	output \g48966/_0_  ;
	output \g48967/_0_  ;
	output \g48968/_0_  ;
	output \g48969/_0_  ;
	output \g48970/_0_  ;
	output \g48971/_0_  ;
	output \g48972/_0_  ;
	output \g48973/_0_  ;
	output \g48974/_0_  ;
	output \g48975/_0_  ;
	output \g48976/_0_  ;
	output \g48977/_0_  ;
	output \g48978/_0_  ;
	output \g48979/_0_  ;
	output \g49/_0_  ;
	output \g49069/_0_  ;
	output \g49070/_0_  ;
	output \g49071/_0_  ;
	output \g49073/_0_  ;
	output \g49074/_0_  ;
	output \g49076/_0_  ;
	output \g49078/_0_  ;
	output \g49081/_0_  ;
	output \g49083/_0_  ;
	output \g49085/_0_  ;
	output \g49087/_0_  ;
	output \g49088/_0_  ;
	output \g49090/_0_  ;
	output \g49092/_0_  ;
	output \g49095/_0_  ;
	output \g49098/_0_  ;
	output \g49125/_0_  ;
	output \g49162/_0_  ;
	output \g49202/_0_  ;
	output \g49203/_0_  ;
	output \g49206/_0_  ;
	output \g49340/_0_  ;
	output \g49457/_0_  ;
	output \g49512/_0_  ;
	output \g49513/_0_  ;
	output \g49514/_0_  ;
	output \g49515/_0_  ;
	output \g49516/_0_  ;
	output \g49517/_0_  ;
	output \g49518/_0_  ;
	output \g49519/_0_  ;
	output \g49520/_0_  ;
	output \g49521/_0_  ;
	output \g49522/_0_  ;
	output \g49523/_0_  ;
	output \g49524/_0_  ;
	output \g49525/_0_  ;
	output \g49526/_0_  ;
	output \g49527/_0_  ;
	output \g49534/_0_  ;
	output \g49551/_0_  ;
	output \g49573/_0_  ;
	output \g49574/_0_  ;
	output \g49578/_0_  ;
	output \g49582/_0_  ;
	output \g49584/_0_  ;
	output \g49592/_0_  ;
	output \g49600/_0_  ;
	output \g49604/_0_  ;
	output \g49608/_0_  ;
	output \g49612/_0_  ;
	output \g49616/_0_  ;
	output \g49619/_0_  ;
	output \g49620/_0_  ;
	output \g49623/_0_  ;
	output \g49627/_0_  ;
	output \g49630/_0_  ;
	output \g49634/_0_  ;
	output \g49635/_0_  ;
	output \g49639/_0_  ;
	output \g49645/_0_  ;
	output \g49744/_0_  ;
	output \g49766/_0_  ;
	output \g50098/_0_  ;
	output \g50124/_0_  ;
	output \g50195/_0_  ;
	output \g50198/_0_  ;
	output \g50201/_0_  ;
	output \g50203/_0_  ;
	output \g50205/_0_  ;
	output \g50207/_0_  ;
	output \g50209/_0_  ;
	output \g50213/_0_  ;
	output \g50222/_0_  ;
	output \g50228/_0_  ;
	output \g50231/_0_  ;
	output \g50237/_0_  ;
	output \g50240/_0_  ;
	output \g50335/_0_  ;
	output \g50477/_0_  ;
	output \g50478/_0_  ;
	output \g50671/_0_  ;
	output \g50757/_0_  ;
	output \g50938/_0_  ;
	output \g50998/_0_  ;
	output \g51008/_0_  ;
	output \g51579/_0_  ;
	output \g51637/_0_  ;
	output \g51662/_0_  ;
	output \g52424/_0_  ;
	output \g53184/_0_  ;
	output \g53206/_0_  ;
	output \g53270/_0_  ;
	output \g53730/_0_  ;
	output \g53754/_0_  ;
	output \g54176/_0_  ;
	output \g54214/_0_  ;
	output \g54229/_0_  ;
	output \g54392/_0_  ;
	output \g54400/_0_  ;
	output \g54415/_0_  ;
	output \g54421/_0_  ;
	output \g54604/_0_  ;
	output \g54607/_0_  ;
	output \g54638/_0_  ;
	output \g54694/_0_  ;
	output \g54759/_0_  ;
	output \g55607/_0_  ;
	output \g55863/_1_  ;
	output \g56073/_0_  ;
	output \g56292/_0_  ;
	output \g56320/_0_  ;
	output \g56527/_0_  ;
	output \g56531/_0_  ;
	output \g56533/_0_  ;
	output \g56562/_0_  ;
	output \g56615/_0_  ;
	output \g56720/_0_  ;
	output \g57044/_0_  ;
	output \g60635/_1_  ;
	output \g62873/_0_  ;
	output \g62886/_0_  ;
	output \g63001/_0_  ;
	output \g63101/_0_  ;
	output \g63129/_0_  ;
	output \g63198/_0_  ;
	output \g63449/_0_  ;
	output \g63471/_0_  ;
	output \g63493/_0_  ;
	output \g63626/_0_  ;
	output \g63688/_0_  ;
	output \g63800/_0_  ;
	output \g63934/_0_  ;
	output \g63954/_0_  ;
	output \g64060/_0_  ;
	output \g64375/_0_  ;
	output \g65/_0_  ;
	output \g67/_0_  ;
	wire _w5394_ ;
	wire _w5393_ ;
	wire _w5392_ ;
	wire _w5391_ ;
	wire _w5390_ ;
	wire _w5389_ ;
	wire _w5388_ ;
	wire _w5387_ ;
	wire _w5386_ ;
	wire _w5385_ ;
	wire _w5384_ ;
	wire _w5383_ ;
	wire _w5382_ ;
	wire _w5381_ ;
	wire _w5380_ ;
	wire _w5379_ ;
	wire _w5378_ ;
	wire _w5377_ ;
	wire _w5376_ ;
	wire _w5375_ ;
	wire _w5374_ ;
	wire _w5373_ ;
	wire _w5372_ ;
	wire _w5371_ ;
	wire _w5370_ ;
	wire _w5369_ ;
	wire _w5368_ ;
	wire _w5367_ ;
	wire _w5366_ ;
	wire _w5365_ ;
	wire _w5364_ ;
	wire _w5363_ ;
	wire _w5362_ ;
	wire _w5361_ ;
	wire _w5360_ ;
	wire _w5359_ ;
	wire _w5358_ ;
	wire _w5357_ ;
	wire _w5356_ ;
	wire _w5355_ ;
	wire _w5354_ ;
	wire _w5353_ ;
	wire _w5352_ ;
	wire _w5351_ ;
	wire _w5350_ ;
	wire _w5349_ ;
	wire _w5348_ ;
	wire _w5347_ ;
	wire _w5346_ ;
	wire _w5345_ ;
	wire _w5344_ ;
	wire _w5343_ ;
	wire _w5342_ ;
	wire _w5341_ ;
	wire _w5340_ ;
	wire _w5339_ ;
	wire _w5338_ ;
	wire _w5337_ ;
	wire _w5336_ ;
	wire _w5335_ ;
	wire _w5334_ ;
	wire _w5333_ ;
	wire _w5332_ ;
	wire _w5331_ ;
	wire _w5330_ ;
	wire _w5329_ ;
	wire _w5328_ ;
	wire _w5327_ ;
	wire _w5326_ ;
	wire _w5325_ ;
	wire _w5324_ ;
	wire _w5323_ ;
	wire _w5322_ ;
	wire _w5321_ ;
	wire _w5320_ ;
	wire _w5319_ ;
	wire _w5318_ ;
	wire _w5317_ ;
	wire _w5316_ ;
	wire _w5315_ ;
	wire _w5314_ ;
	wire _w5313_ ;
	wire _w5312_ ;
	wire _w5311_ ;
	wire _w5310_ ;
	wire _w5309_ ;
	wire _w5308_ ;
	wire _w5307_ ;
	wire _w5306_ ;
	wire _w5305_ ;
	wire _w5304_ ;
	wire _w5303_ ;
	wire _w5302_ ;
	wire _w5301_ ;
	wire _w5300_ ;
	wire _w5299_ ;
	wire _w5298_ ;
	wire _w5297_ ;
	wire _w5296_ ;
	wire _w5295_ ;
	wire _w5294_ ;
	wire _w5293_ ;
	wire _w5292_ ;
	wire _w5291_ ;
	wire _w5290_ ;
	wire _w5289_ ;
	wire _w5288_ ;
	wire _w5287_ ;
	wire _w5286_ ;
	wire _w5285_ ;
	wire _w5284_ ;
	wire _w5283_ ;
	wire _w5282_ ;
	wire _w5281_ ;
	wire _w5280_ ;
	wire _w5279_ ;
	wire _w5278_ ;
	wire _w5277_ ;
	wire _w5276_ ;
	wire _w5275_ ;
	wire _w5274_ ;
	wire _w5273_ ;
	wire _w5272_ ;
	wire _w5271_ ;
	wire _w5270_ ;
	wire _w5269_ ;
	wire _w5268_ ;
	wire _w5267_ ;
	wire _w5266_ ;
	wire _w5265_ ;
	wire _w5264_ ;
	wire _w5263_ ;
	wire _w5262_ ;
	wire _w5261_ ;
	wire _w5260_ ;
	wire _w5259_ ;
	wire _w5258_ ;
	wire _w5257_ ;
	wire _w5256_ ;
	wire _w5255_ ;
	wire _w5254_ ;
	wire _w5253_ ;
	wire _w5252_ ;
	wire _w5251_ ;
	wire _w5250_ ;
	wire _w5249_ ;
	wire _w5248_ ;
	wire _w5247_ ;
	wire _w5246_ ;
	wire _w5245_ ;
	wire _w5244_ ;
	wire _w5243_ ;
	wire _w5242_ ;
	wire _w5241_ ;
	wire _w5240_ ;
	wire _w5239_ ;
	wire _w5238_ ;
	wire _w5237_ ;
	wire _w5236_ ;
	wire _w5235_ ;
	wire _w5234_ ;
	wire _w5233_ ;
	wire _w5232_ ;
	wire _w5231_ ;
	wire _w5230_ ;
	wire _w5229_ ;
	wire _w5228_ ;
	wire _w5227_ ;
	wire _w5226_ ;
	wire _w5225_ ;
	wire _w5224_ ;
	wire _w5223_ ;
	wire _w5222_ ;
	wire _w5221_ ;
	wire _w5220_ ;
	wire _w5219_ ;
	wire _w5218_ ;
	wire _w5217_ ;
	wire _w5216_ ;
	wire _w5215_ ;
	wire _w5214_ ;
	wire _w5213_ ;
	wire _w5212_ ;
	wire _w5211_ ;
	wire _w5210_ ;
	wire _w5209_ ;
	wire _w5208_ ;
	wire _w5207_ ;
	wire _w5206_ ;
	wire _w5205_ ;
	wire _w5204_ ;
	wire _w5203_ ;
	wire _w5202_ ;
	wire _w5201_ ;
	wire _w5200_ ;
	wire _w5199_ ;
	wire _w5198_ ;
	wire _w5197_ ;
	wire _w5196_ ;
	wire _w5195_ ;
	wire _w5194_ ;
	wire _w5193_ ;
	wire _w5192_ ;
	wire _w5191_ ;
	wire _w5190_ ;
	wire _w5189_ ;
	wire _w5188_ ;
	wire _w5187_ ;
	wire _w5186_ ;
	wire _w5185_ ;
	wire _w5184_ ;
	wire _w5183_ ;
	wire _w5182_ ;
	wire _w5181_ ;
	wire _w5180_ ;
	wire _w5179_ ;
	wire _w5178_ ;
	wire _w5177_ ;
	wire _w5176_ ;
	wire _w5175_ ;
	wire _w5174_ ;
	wire _w5173_ ;
	wire _w5172_ ;
	wire _w5171_ ;
	wire _w5170_ ;
	wire _w5169_ ;
	wire _w5168_ ;
	wire _w5167_ ;
	wire _w5166_ ;
	wire _w5165_ ;
	wire _w5164_ ;
	wire _w5163_ ;
	wire _w5162_ ;
	wire _w5161_ ;
	wire _w5160_ ;
	wire _w5159_ ;
	wire _w5158_ ;
	wire _w5157_ ;
	wire _w5156_ ;
	wire _w5155_ ;
	wire _w5154_ ;
	wire _w5153_ ;
	wire _w5152_ ;
	wire _w5151_ ;
	wire _w5150_ ;
	wire _w5149_ ;
	wire _w5148_ ;
	wire _w5147_ ;
	wire _w5146_ ;
	wire _w5145_ ;
	wire _w5144_ ;
	wire _w5143_ ;
	wire _w5142_ ;
	wire _w5141_ ;
	wire _w5140_ ;
	wire _w5139_ ;
	wire _w5138_ ;
	wire _w5137_ ;
	wire _w5136_ ;
	wire _w5135_ ;
	wire _w5134_ ;
	wire _w5133_ ;
	wire _w5132_ ;
	wire _w5131_ ;
	wire _w5130_ ;
	wire _w5129_ ;
	wire _w5128_ ;
	wire _w5127_ ;
	wire _w5126_ ;
	wire _w5125_ ;
	wire _w5124_ ;
	wire _w5123_ ;
	wire _w5122_ ;
	wire _w5121_ ;
	wire _w5120_ ;
	wire _w5119_ ;
	wire _w5118_ ;
	wire _w5117_ ;
	wire _w5116_ ;
	wire _w5115_ ;
	wire _w5114_ ;
	wire _w5113_ ;
	wire _w5112_ ;
	wire _w5111_ ;
	wire _w5110_ ;
	wire _w5109_ ;
	wire _w5108_ ;
	wire _w5107_ ;
	wire _w5106_ ;
	wire _w5105_ ;
	wire _w5104_ ;
	wire _w5103_ ;
	wire _w5102_ ;
	wire _w5101_ ;
	wire _w5100_ ;
	wire _w5099_ ;
	wire _w5098_ ;
	wire _w5097_ ;
	wire _w5096_ ;
	wire _w5095_ ;
	wire _w5094_ ;
	wire _w5093_ ;
	wire _w5092_ ;
	wire _w5091_ ;
	wire _w5090_ ;
	wire _w5089_ ;
	wire _w5088_ ;
	wire _w5087_ ;
	wire _w5086_ ;
	wire _w5085_ ;
	wire _w5084_ ;
	wire _w5083_ ;
	wire _w5082_ ;
	wire _w5081_ ;
	wire _w5080_ ;
	wire _w5079_ ;
	wire _w5078_ ;
	wire _w5077_ ;
	wire _w5076_ ;
	wire _w5075_ ;
	wire _w5074_ ;
	wire _w5073_ ;
	wire _w5072_ ;
	wire _w5071_ ;
	wire _w5070_ ;
	wire _w5069_ ;
	wire _w5068_ ;
	wire _w5067_ ;
	wire _w5066_ ;
	wire _w5065_ ;
	wire _w5064_ ;
	wire _w5063_ ;
	wire _w5062_ ;
	wire _w5061_ ;
	wire _w5060_ ;
	wire _w5059_ ;
	wire _w5058_ ;
	wire _w5057_ ;
	wire _w5056_ ;
	wire _w5055_ ;
	wire _w5054_ ;
	wire _w5053_ ;
	wire _w5052_ ;
	wire _w5051_ ;
	wire _w5050_ ;
	wire _w5049_ ;
	wire _w5048_ ;
	wire _w5047_ ;
	wire _w5046_ ;
	wire _w5045_ ;
	wire _w5044_ ;
	wire _w5043_ ;
	wire _w5042_ ;
	wire _w5041_ ;
	wire _w5040_ ;
	wire _w5039_ ;
	wire _w5038_ ;
	wire _w5037_ ;
	wire _w5036_ ;
	wire _w5035_ ;
	wire _w5034_ ;
	wire _w5033_ ;
	wire _w5032_ ;
	wire _w5031_ ;
	wire _w5030_ ;
	wire _w5029_ ;
	wire _w5028_ ;
	wire _w5027_ ;
	wire _w5026_ ;
	wire _w5025_ ;
	wire _w5024_ ;
	wire _w5023_ ;
	wire _w5022_ ;
	wire _w5021_ ;
	wire _w5020_ ;
	wire _w5019_ ;
	wire _w5018_ ;
	wire _w5017_ ;
	wire _w5016_ ;
	wire _w5015_ ;
	wire _w5014_ ;
	wire _w5013_ ;
	wire _w5012_ ;
	wire _w5011_ ;
	wire _w5010_ ;
	wire _w5009_ ;
	wire _w5008_ ;
	wire _w5007_ ;
	wire _w5006_ ;
	wire _w5005_ ;
	wire _w5004_ ;
	wire _w5003_ ;
	wire _w5002_ ;
	wire _w5001_ ;
	wire _w5000_ ;
	wire _w4999_ ;
	wire _w4998_ ;
	wire _w4997_ ;
	wire _w4996_ ;
	wire _w4995_ ;
	wire _w4994_ ;
	wire _w4993_ ;
	wire _w4992_ ;
	wire _w4991_ ;
	wire _w4990_ ;
	wire _w4989_ ;
	wire _w4988_ ;
	wire _w4987_ ;
	wire _w4986_ ;
	wire _w4985_ ;
	wire _w4984_ ;
	wire _w4983_ ;
	wire _w4982_ ;
	wire _w4981_ ;
	wire _w4980_ ;
	wire _w4979_ ;
	wire _w4978_ ;
	wire _w4977_ ;
	wire _w4976_ ;
	wire _w4975_ ;
	wire _w4974_ ;
	wire _w4973_ ;
	wire _w4972_ ;
	wire _w4971_ ;
	wire _w4970_ ;
	wire _w4969_ ;
	wire _w4968_ ;
	wire _w4967_ ;
	wire _w4966_ ;
	wire _w4965_ ;
	wire _w4964_ ;
	wire _w4963_ ;
	wire _w4962_ ;
	wire _w4961_ ;
	wire _w4960_ ;
	wire _w4959_ ;
	wire _w4958_ ;
	wire _w4957_ ;
	wire _w4956_ ;
	wire _w4955_ ;
	wire _w4954_ ;
	wire _w4953_ ;
	wire _w4952_ ;
	wire _w4951_ ;
	wire _w4950_ ;
	wire _w4949_ ;
	wire _w4948_ ;
	wire _w4947_ ;
	wire _w4946_ ;
	wire _w4945_ ;
	wire _w4944_ ;
	wire _w4943_ ;
	wire _w4942_ ;
	wire _w4941_ ;
	wire _w4940_ ;
	wire _w4939_ ;
	wire _w4938_ ;
	wire _w4937_ ;
	wire _w4936_ ;
	wire _w4935_ ;
	wire _w4934_ ;
	wire _w4933_ ;
	wire _w4932_ ;
	wire _w4931_ ;
	wire _w4930_ ;
	wire _w4929_ ;
	wire _w4928_ ;
	wire _w4927_ ;
	wire _w4926_ ;
	wire _w4925_ ;
	wire _w4924_ ;
	wire _w4923_ ;
	wire _w4922_ ;
	wire _w4921_ ;
	wire _w4920_ ;
	wire _w4919_ ;
	wire _w4918_ ;
	wire _w4917_ ;
	wire _w4916_ ;
	wire _w4915_ ;
	wire _w4914_ ;
	wire _w4913_ ;
	wire _w4912_ ;
	wire _w4911_ ;
	wire _w4910_ ;
	wire _w4909_ ;
	wire _w4908_ ;
	wire _w4907_ ;
	wire _w4906_ ;
	wire _w4905_ ;
	wire _w4904_ ;
	wire _w4903_ ;
	wire _w4902_ ;
	wire _w4901_ ;
	wire _w4900_ ;
	wire _w4899_ ;
	wire _w4898_ ;
	wire _w4897_ ;
	wire _w4896_ ;
	wire _w4895_ ;
	wire _w4894_ ;
	wire _w4893_ ;
	wire _w4892_ ;
	wire _w4891_ ;
	wire _w4890_ ;
	wire _w4889_ ;
	wire _w4888_ ;
	wire _w4887_ ;
	wire _w4886_ ;
	wire _w4885_ ;
	wire _w4884_ ;
	wire _w4883_ ;
	wire _w4882_ ;
	wire _w4881_ ;
	wire _w4880_ ;
	wire _w4879_ ;
	wire _w4878_ ;
	wire _w4877_ ;
	wire _w4876_ ;
	wire _w4875_ ;
	wire _w4874_ ;
	wire _w4873_ ;
	wire _w4872_ ;
	wire _w4871_ ;
	wire _w4870_ ;
	wire _w4869_ ;
	wire _w4868_ ;
	wire _w4867_ ;
	wire _w4866_ ;
	wire _w4865_ ;
	wire _w4864_ ;
	wire _w4863_ ;
	wire _w4862_ ;
	wire _w4861_ ;
	wire _w4860_ ;
	wire _w4859_ ;
	wire _w4858_ ;
	wire _w4857_ ;
	wire _w4856_ ;
	wire _w4855_ ;
	wire _w4854_ ;
	wire _w4853_ ;
	wire _w4852_ ;
	wire _w4851_ ;
	wire _w4850_ ;
	wire _w4849_ ;
	wire _w4848_ ;
	wire _w4847_ ;
	wire _w4846_ ;
	wire _w4845_ ;
	wire _w4844_ ;
	wire _w4843_ ;
	wire _w4842_ ;
	wire _w4841_ ;
	wire _w4840_ ;
	wire _w4839_ ;
	wire _w4838_ ;
	wire _w4837_ ;
	wire _w4836_ ;
	wire _w4835_ ;
	wire _w4834_ ;
	wire _w4833_ ;
	wire _w4832_ ;
	wire _w4831_ ;
	wire _w4830_ ;
	wire _w4829_ ;
	wire _w4828_ ;
	wire _w4827_ ;
	wire _w4826_ ;
	wire _w4825_ ;
	wire _w4824_ ;
	wire _w4823_ ;
	wire _w4822_ ;
	wire _w4821_ ;
	wire _w4820_ ;
	wire _w4819_ ;
	wire _w4818_ ;
	wire _w4817_ ;
	wire _w4816_ ;
	wire _w4815_ ;
	wire _w4814_ ;
	wire _w4813_ ;
	wire _w4812_ ;
	wire _w4811_ ;
	wire _w4810_ ;
	wire _w4809_ ;
	wire _w4808_ ;
	wire _w4807_ ;
	wire _w4806_ ;
	wire _w4805_ ;
	wire _w4804_ ;
	wire _w4803_ ;
	wire _w4802_ ;
	wire _w4801_ ;
	wire _w4800_ ;
	wire _w4799_ ;
	wire _w4798_ ;
	wire _w4797_ ;
	wire _w4796_ ;
	wire _w4795_ ;
	wire _w4794_ ;
	wire _w4793_ ;
	wire _w4792_ ;
	wire _w4791_ ;
	wire _w4790_ ;
	wire _w4789_ ;
	wire _w4788_ ;
	wire _w4787_ ;
	wire _w4786_ ;
	wire _w4785_ ;
	wire _w4784_ ;
	wire _w4783_ ;
	wire _w4782_ ;
	wire _w4781_ ;
	wire _w4780_ ;
	wire _w4779_ ;
	wire _w4778_ ;
	wire _w4777_ ;
	wire _w4776_ ;
	wire _w4775_ ;
	wire _w4774_ ;
	wire _w4773_ ;
	wire _w4772_ ;
	wire _w4771_ ;
	wire _w4770_ ;
	wire _w4769_ ;
	wire _w4768_ ;
	wire _w4767_ ;
	wire _w4766_ ;
	wire _w4765_ ;
	wire _w4764_ ;
	wire _w4763_ ;
	wire _w4762_ ;
	wire _w4761_ ;
	wire _w4760_ ;
	wire _w4759_ ;
	wire _w4758_ ;
	wire _w4757_ ;
	wire _w4756_ ;
	wire _w4755_ ;
	wire _w4754_ ;
	wire _w4753_ ;
	wire _w4752_ ;
	wire _w4751_ ;
	wire _w4750_ ;
	wire _w4749_ ;
	wire _w4748_ ;
	wire _w4747_ ;
	wire _w4746_ ;
	wire _w4745_ ;
	wire _w4744_ ;
	wire _w4743_ ;
	wire _w4742_ ;
	wire _w4741_ ;
	wire _w4740_ ;
	wire _w4739_ ;
	wire _w4738_ ;
	wire _w4737_ ;
	wire _w4736_ ;
	wire _w4735_ ;
	wire _w4734_ ;
	wire _w4733_ ;
	wire _w4732_ ;
	wire _w4731_ ;
	wire _w4730_ ;
	wire _w4729_ ;
	wire _w4728_ ;
	wire _w4727_ ;
	wire _w4726_ ;
	wire _w4725_ ;
	wire _w4724_ ;
	wire _w4723_ ;
	wire _w4722_ ;
	wire _w4721_ ;
	wire _w4720_ ;
	wire _w4719_ ;
	wire _w4718_ ;
	wire _w4717_ ;
	wire _w4716_ ;
	wire _w4715_ ;
	wire _w4714_ ;
	wire _w4713_ ;
	wire _w4712_ ;
	wire _w4711_ ;
	wire _w4710_ ;
	wire _w4709_ ;
	wire _w4708_ ;
	wire _w4707_ ;
	wire _w4706_ ;
	wire _w4705_ ;
	wire _w4704_ ;
	wire _w4703_ ;
	wire _w4702_ ;
	wire _w4701_ ;
	wire _w4700_ ;
	wire _w4699_ ;
	wire _w4698_ ;
	wire _w4697_ ;
	wire _w4696_ ;
	wire _w4695_ ;
	wire _w4694_ ;
	wire _w4693_ ;
	wire _w4692_ ;
	wire _w4691_ ;
	wire _w4690_ ;
	wire _w4689_ ;
	wire _w4688_ ;
	wire _w4687_ ;
	wire _w4686_ ;
	wire _w4685_ ;
	wire _w4684_ ;
	wire _w4683_ ;
	wire _w4682_ ;
	wire _w4681_ ;
	wire _w4680_ ;
	wire _w4679_ ;
	wire _w4678_ ;
	wire _w4677_ ;
	wire _w4676_ ;
	wire _w4675_ ;
	wire _w4674_ ;
	wire _w4673_ ;
	wire _w4672_ ;
	wire _w4671_ ;
	wire _w4670_ ;
	wire _w4669_ ;
	wire _w4668_ ;
	wire _w4667_ ;
	wire _w4666_ ;
	wire _w4665_ ;
	wire _w4664_ ;
	wire _w4663_ ;
	wire _w4662_ ;
	wire _w4661_ ;
	wire _w4660_ ;
	wire _w4659_ ;
	wire _w4658_ ;
	wire _w4657_ ;
	wire _w4656_ ;
	wire _w4655_ ;
	wire _w4654_ ;
	wire _w4653_ ;
	wire _w4652_ ;
	wire _w4651_ ;
	wire _w4650_ ;
	wire _w4649_ ;
	wire _w4648_ ;
	wire _w4647_ ;
	wire _w4646_ ;
	wire _w4645_ ;
	wire _w4644_ ;
	wire _w4643_ ;
	wire _w4642_ ;
	wire _w4641_ ;
	wire _w4640_ ;
	wire _w4639_ ;
	wire _w4638_ ;
	wire _w4637_ ;
	wire _w4636_ ;
	wire _w4635_ ;
	wire _w4634_ ;
	wire _w4633_ ;
	wire _w4632_ ;
	wire _w4631_ ;
	wire _w4630_ ;
	wire _w4629_ ;
	wire _w4628_ ;
	wire _w4627_ ;
	wire _w4626_ ;
	wire _w4625_ ;
	wire _w4624_ ;
	wire _w4623_ ;
	wire _w4622_ ;
	wire _w4621_ ;
	wire _w4620_ ;
	wire _w4619_ ;
	wire _w4618_ ;
	wire _w4617_ ;
	wire _w4616_ ;
	wire _w4615_ ;
	wire _w4614_ ;
	wire _w4613_ ;
	wire _w4612_ ;
	wire _w4611_ ;
	wire _w4610_ ;
	wire _w4609_ ;
	wire _w4608_ ;
	wire _w4607_ ;
	wire _w4606_ ;
	wire _w4605_ ;
	wire _w4604_ ;
	wire _w4603_ ;
	wire _w4602_ ;
	wire _w4601_ ;
	wire _w4600_ ;
	wire _w4599_ ;
	wire _w4598_ ;
	wire _w4597_ ;
	wire _w4596_ ;
	wire _w4595_ ;
	wire _w4594_ ;
	wire _w4593_ ;
	wire _w4592_ ;
	wire _w4591_ ;
	wire _w4590_ ;
	wire _w4589_ ;
	wire _w4588_ ;
	wire _w4587_ ;
	wire _w4586_ ;
	wire _w4585_ ;
	wire _w4584_ ;
	wire _w4583_ ;
	wire _w4582_ ;
	wire _w4581_ ;
	wire _w4580_ ;
	wire _w4579_ ;
	wire _w4578_ ;
	wire _w4577_ ;
	wire _w4576_ ;
	wire _w4575_ ;
	wire _w4574_ ;
	wire _w4573_ ;
	wire _w4572_ ;
	wire _w4571_ ;
	wire _w4570_ ;
	wire _w4569_ ;
	wire _w4568_ ;
	wire _w4567_ ;
	wire _w4566_ ;
	wire _w4565_ ;
	wire _w4564_ ;
	wire _w4563_ ;
	wire _w4562_ ;
	wire _w4561_ ;
	wire _w4560_ ;
	wire _w4559_ ;
	wire _w4558_ ;
	wire _w4557_ ;
	wire _w4556_ ;
	wire _w4555_ ;
	wire _w4554_ ;
	wire _w4553_ ;
	wire _w4552_ ;
	wire _w4551_ ;
	wire _w4550_ ;
	wire _w4549_ ;
	wire _w4548_ ;
	wire _w4547_ ;
	wire _w4546_ ;
	wire _w4545_ ;
	wire _w4544_ ;
	wire _w4543_ ;
	wire _w4542_ ;
	wire _w4541_ ;
	wire _w4540_ ;
	wire _w4539_ ;
	wire _w4538_ ;
	wire _w4537_ ;
	wire _w4536_ ;
	wire _w4535_ ;
	wire _w4534_ ;
	wire _w4533_ ;
	wire _w4532_ ;
	wire _w4531_ ;
	wire _w4530_ ;
	wire _w4529_ ;
	wire _w4528_ ;
	wire _w4527_ ;
	wire _w4526_ ;
	wire _w4525_ ;
	wire _w4524_ ;
	wire _w4523_ ;
	wire _w4522_ ;
	wire _w4521_ ;
	wire _w4520_ ;
	wire _w4519_ ;
	wire _w4518_ ;
	wire _w4517_ ;
	wire _w4516_ ;
	wire _w4515_ ;
	wire _w4514_ ;
	wire _w4513_ ;
	wire _w4512_ ;
	wire _w4511_ ;
	wire _w4510_ ;
	wire _w4509_ ;
	wire _w4508_ ;
	wire _w4507_ ;
	wire _w4506_ ;
	wire _w4505_ ;
	wire _w4504_ ;
	wire _w4503_ ;
	wire _w4502_ ;
	wire _w4501_ ;
	wire _w4500_ ;
	wire _w4499_ ;
	wire _w4498_ ;
	wire _w4497_ ;
	wire _w4496_ ;
	wire _w4495_ ;
	wire _w4494_ ;
	wire _w4493_ ;
	wire _w4492_ ;
	wire _w4491_ ;
	wire _w4490_ ;
	wire _w4489_ ;
	wire _w4488_ ;
	wire _w4487_ ;
	wire _w4486_ ;
	wire _w4485_ ;
	wire _w4484_ ;
	wire _w4483_ ;
	wire _w4482_ ;
	wire _w4481_ ;
	wire _w4480_ ;
	wire _w4479_ ;
	wire _w4478_ ;
	wire _w4477_ ;
	wire _w4476_ ;
	wire _w4475_ ;
	wire _w4474_ ;
	wire _w4473_ ;
	wire _w4472_ ;
	wire _w4471_ ;
	wire _w4470_ ;
	wire _w4469_ ;
	wire _w4468_ ;
	wire _w4467_ ;
	wire _w4466_ ;
	wire _w4465_ ;
	wire _w4464_ ;
	wire _w4463_ ;
	wire _w4462_ ;
	wire _w4461_ ;
	wire _w4460_ ;
	wire _w4459_ ;
	wire _w4458_ ;
	wire _w4457_ ;
	wire _w4456_ ;
	wire _w4455_ ;
	wire _w4454_ ;
	wire _w4453_ ;
	wire _w4452_ ;
	wire _w4451_ ;
	wire _w4450_ ;
	wire _w4449_ ;
	wire _w4448_ ;
	wire _w4447_ ;
	wire _w4446_ ;
	wire _w4445_ ;
	wire _w4444_ ;
	wire _w4443_ ;
	wire _w4442_ ;
	wire _w4441_ ;
	wire _w4440_ ;
	wire _w4439_ ;
	wire _w4438_ ;
	wire _w4437_ ;
	wire _w4436_ ;
	wire _w4435_ ;
	wire _w4434_ ;
	wire _w4433_ ;
	wire _w4432_ ;
	wire _w4431_ ;
	wire _w4430_ ;
	wire _w4429_ ;
	wire _w4428_ ;
	wire _w4427_ ;
	wire _w4426_ ;
	wire _w4425_ ;
	wire _w4424_ ;
	wire _w4423_ ;
	wire _w4422_ ;
	wire _w4421_ ;
	wire _w4420_ ;
	wire _w4419_ ;
	wire _w4418_ ;
	wire _w4417_ ;
	wire _w4416_ ;
	wire _w4415_ ;
	wire _w4414_ ;
	wire _w4413_ ;
	wire _w4412_ ;
	wire _w4411_ ;
	wire _w4410_ ;
	wire _w4409_ ;
	wire _w4408_ ;
	wire _w4407_ ;
	wire _w4406_ ;
	wire _w4405_ ;
	wire _w4404_ ;
	wire _w4403_ ;
	wire _w4402_ ;
	wire _w4401_ ;
	wire _w4400_ ;
	wire _w4399_ ;
	wire _w4398_ ;
	wire _w4397_ ;
	wire _w4396_ ;
	wire _w4395_ ;
	wire _w4394_ ;
	wire _w4393_ ;
	wire _w4392_ ;
	wire _w4391_ ;
	wire _w4390_ ;
	wire _w4389_ ;
	wire _w4388_ ;
	wire _w4387_ ;
	wire _w4386_ ;
	wire _w4385_ ;
	wire _w4384_ ;
	wire _w4383_ ;
	wire _w4382_ ;
	wire _w4381_ ;
	wire _w4380_ ;
	wire _w4379_ ;
	wire _w4378_ ;
	wire _w4377_ ;
	wire _w4376_ ;
	wire _w4375_ ;
	wire _w4374_ ;
	wire _w4373_ ;
	wire _w4372_ ;
	wire _w4371_ ;
	wire _w4370_ ;
	wire _w4369_ ;
	wire _w4368_ ;
	wire _w4367_ ;
	wire _w4366_ ;
	wire _w4365_ ;
	wire _w4364_ ;
	wire _w4363_ ;
	wire _w4362_ ;
	wire _w4361_ ;
	wire _w4360_ ;
	wire _w4359_ ;
	wire _w4358_ ;
	wire _w4357_ ;
	wire _w4356_ ;
	wire _w4355_ ;
	wire _w4354_ ;
	wire _w4353_ ;
	wire _w4352_ ;
	wire _w4351_ ;
	wire _w4350_ ;
	wire _w4349_ ;
	wire _w4348_ ;
	wire _w4347_ ;
	wire _w4346_ ;
	wire _w4345_ ;
	wire _w4344_ ;
	wire _w4343_ ;
	wire _w4342_ ;
	wire _w4341_ ;
	wire _w4340_ ;
	wire _w4339_ ;
	wire _w4338_ ;
	wire _w4337_ ;
	wire _w4336_ ;
	wire _w4335_ ;
	wire _w4334_ ;
	wire _w4333_ ;
	wire _w4332_ ;
	wire _w4331_ ;
	wire _w4330_ ;
	wire _w4329_ ;
	wire _w4328_ ;
	wire _w4327_ ;
	wire _w4326_ ;
	wire _w4325_ ;
	wire _w4324_ ;
	wire _w4323_ ;
	wire _w4322_ ;
	wire _w4321_ ;
	wire _w4320_ ;
	wire _w4319_ ;
	wire _w4318_ ;
	wire _w4317_ ;
	wire _w4316_ ;
	wire _w4315_ ;
	wire _w4314_ ;
	wire _w4313_ ;
	wire _w4312_ ;
	wire _w4311_ ;
	wire _w4310_ ;
	wire _w4309_ ;
	wire _w4308_ ;
	wire _w4307_ ;
	wire _w4306_ ;
	wire _w4305_ ;
	wire _w4304_ ;
	wire _w4303_ ;
	wire _w4302_ ;
	wire _w4301_ ;
	wire _w4300_ ;
	wire _w4299_ ;
	wire _w4298_ ;
	wire _w4297_ ;
	wire _w4296_ ;
	wire _w4295_ ;
	wire _w4294_ ;
	wire _w4293_ ;
	wire _w4292_ ;
	wire _w4291_ ;
	wire _w4290_ ;
	wire _w4289_ ;
	wire _w4288_ ;
	wire _w4287_ ;
	wire _w4286_ ;
	wire _w4285_ ;
	wire _w4284_ ;
	wire _w4283_ ;
	wire _w4282_ ;
	wire _w4281_ ;
	wire _w4280_ ;
	wire _w4279_ ;
	wire _w4278_ ;
	wire _w4277_ ;
	wire _w4276_ ;
	wire _w4275_ ;
	wire _w4274_ ;
	wire _w4273_ ;
	wire _w4272_ ;
	wire _w4271_ ;
	wire _w4270_ ;
	wire _w4269_ ;
	wire _w4268_ ;
	wire _w4267_ ;
	wire _w4266_ ;
	wire _w4265_ ;
	wire _w4264_ ;
	wire _w4263_ ;
	wire _w4262_ ;
	wire _w4261_ ;
	wire _w4260_ ;
	wire _w4259_ ;
	wire _w4258_ ;
	wire _w4257_ ;
	wire _w4256_ ;
	wire _w4255_ ;
	wire _w4254_ ;
	wire _w4253_ ;
	wire _w4252_ ;
	wire _w4251_ ;
	wire _w4250_ ;
	wire _w4249_ ;
	wire _w4248_ ;
	wire _w4247_ ;
	wire _w4246_ ;
	wire _w4245_ ;
	wire _w4244_ ;
	wire _w4243_ ;
	wire _w4242_ ;
	wire _w4241_ ;
	wire _w4240_ ;
	wire _w4239_ ;
	wire _w4238_ ;
	wire _w4237_ ;
	wire _w4236_ ;
	wire _w4235_ ;
	wire _w4234_ ;
	wire _w4233_ ;
	wire _w4232_ ;
	wire _w4231_ ;
	wire _w4230_ ;
	wire _w4229_ ;
	wire _w4228_ ;
	wire _w4227_ ;
	wire _w4226_ ;
	wire _w4225_ ;
	wire _w4224_ ;
	wire _w4223_ ;
	wire _w4222_ ;
	wire _w4221_ ;
	wire _w4220_ ;
	wire _w4219_ ;
	wire _w4218_ ;
	wire _w4217_ ;
	wire _w4216_ ;
	wire _w4215_ ;
	wire _w4214_ ;
	wire _w4213_ ;
	wire _w4212_ ;
	wire _w4211_ ;
	wire _w4210_ ;
	wire _w4209_ ;
	wire _w4208_ ;
	wire _w4207_ ;
	wire _w4206_ ;
	wire _w4205_ ;
	wire _w4204_ ;
	wire _w4203_ ;
	wire _w4202_ ;
	wire _w4201_ ;
	wire _w4200_ ;
	wire _w4199_ ;
	wire _w4198_ ;
	wire _w4197_ ;
	wire _w4196_ ;
	wire _w4195_ ;
	wire _w4194_ ;
	wire _w4193_ ;
	wire _w4192_ ;
	wire _w4191_ ;
	wire _w4190_ ;
	wire _w4189_ ;
	wire _w4188_ ;
	wire _w4187_ ;
	wire _w4186_ ;
	wire _w4185_ ;
	wire _w4184_ ;
	wire _w4183_ ;
	wire _w4182_ ;
	wire _w4181_ ;
	wire _w4180_ ;
	wire _w4179_ ;
	wire _w4178_ ;
	wire _w4177_ ;
	wire _w4176_ ;
	wire _w4175_ ;
	wire _w4174_ ;
	wire _w4173_ ;
	wire _w4172_ ;
	wire _w4171_ ;
	wire _w4170_ ;
	wire _w4169_ ;
	wire _w4168_ ;
	wire _w4167_ ;
	wire _w4166_ ;
	wire _w4165_ ;
	wire _w4164_ ;
	wire _w4163_ ;
	wire _w4162_ ;
	wire _w4161_ ;
	wire _w4160_ ;
	wire _w4159_ ;
	wire _w4158_ ;
	wire _w4157_ ;
	wire _w4156_ ;
	wire _w4155_ ;
	wire _w4154_ ;
	wire _w4153_ ;
	wire _w4152_ ;
	wire _w4151_ ;
	wire _w4150_ ;
	wire _w4149_ ;
	wire _w4148_ ;
	wire _w4147_ ;
	wire _w4146_ ;
	wire _w4145_ ;
	wire _w4144_ ;
	wire _w4143_ ;
	wire _w4142_ ;
	wire _w4141_ ;
	wire _w4140_ ;
	wire _w4139_ ;
	wire _w4138_ ;
	wire _w4137_ ;
	wire _w4136_ ;
	wire _w4135_ ;
	wire _w4134_ ;
	wire _w4133_ ;
	wire _w4132_ ;
	wire _w4131_ ;
	wire _w4130_ ;
	wire _w4129_ ;
	wire _w4128_ ;
	wire _w4127_ ;
	wire _w4126_ ;
	wire _w4125_ ;
	wire _w4124_ ;
	wire _w4123_ ;
	wire _w4122_ ;
	wire _w4121_ ;
	wire _w4120_ ;
	wire _w4119_ ;
	wire _w4118_ ;
	wire _w4117_ ;
	wire _w4116_ ;
	wire _w4115_ ;
	wire _w4114_ ;
	wire _w4113_ ;
	wire _w4112_ ;
	wire _w4111_ ;
	wire _w4110_ ;
	wire _w4109_ ;
	wire _w4108_ ;
	wire _w4107_ ;
	wire _w4106_ ;
	wire _w4105_ ;
	wire _w4104_ ;
	wire _w4103_ ;
	wire _w4102_ ;
	wire _w4101_ ;
	wire _w4100_ ;
	wire _w4099_ ;
	wire _w4098_ ;
	wire _w4097_ ;
	wire _w4096_ ;
	wire _w4095_ ;
	wire _w4094_ ;
	wire _w4093_ ;
	wire _w4092_ ;
	wire _w4091_ ;
	wire _w4090_ ;
	wire _w4089_ ;
	wire _w4088_ ;
	wire _w4087_ ;
	wire _w4086_ ;
	wire _w4085_ ;
	wire _w4084_ ;
	wire _w4083_ ;
	wire _w4082_ ;
	wire _w4081_ ;
	wire _w4080_ ;
	wire _w4079_ ;
	wire _w4078_ ;
	wire _w4077_ ;
	wire _w4076_ ;
	wire _w4075_ ;
	wire _w4074_ ;
	wire _w4073_ ;
	wire _w4072_ ;
	wire _w4071_ ;
	wire _w4070_ ;
	wire _w4069_ ;
	wire _w4068_ ;
	wire _w4067_ ;
	wire _w4066_ ;
	wire _w4065_ ;
	wire _w4064_ ;
	wire _w4063_ ;
	wire _w4062_ ;
	wire _w4061_ ;
	wire _w4060_ ;
	wire _w4059_ ;
	wire _w4058_ ;
	wire _w4057_ ;
	wire _w4056_ ;
	wire _w4055_ ;
	wire _w4054_ ;
	wire _w4053_ ;
	wire _w4052_ ;
	wire _w4051_ ;
	wire _w4050_ ;
	wire _w4049_ ;
	wire _w4048_ ;
	wire _w4047_ ;
	wire _w4046_ ;
	wire _w4045_ ;
	wire _w4044_ ;
	wire _w4043_ ;
	wire _w4042_ ;
	wire _w4041_ ;
	wire _w4040_ ;
	wire _w4039_ ;
	wire _w4038_ ;
	wire _w4037_ ;
	wire _w4036_ ;
	wire _w4035_ ;
	wire _w4034_ ;
	wire _w4033_ ;
	wire _w4032_ ;
	wire _w4031_ ;
	wire _w4030_ ;
	wire _w4029_ ;
	wire _w4028_ ;
	wire _w4027_ ;
	wire _w4026_ ;
	wire _w4025_ ;
	wire _w4024_ ;
	wire _w4023_ ;
	wire _w4022_ ;
	wire _w4021_ ;
	wire _w4020_ ;
	wire _w4019_ ;
	wire _w4018_ ;
	wire _w4017_ ;
	wire _w4016_ ;
	wire _w4015_ ;
	wire _w4014_ ;
	wire _w4013_ ;
	wire _w4012_ ;
	wire _w4011_ ;
	wire _w4010_ ;
	wire _w4009_ ;
	wire _w4008_ ;
	wire _w4007_ ;
	wire _w4006_ ;
	wire _w4005_ ;
	wire _w4004_ ;
	wire _w4003_ ;
	wire _w4002_ ;
	wire _w4001_ ;
	wire _w4000_ ;
	wire _w3999_ ;
	wire _w3998_ ;
	wire _w3997_ ;
	wire _w3996_ ;
	wire _w3995_ ;
	wire _w3994_ ;
	wire _w3993_ ;
	wire _w3992_ ;
	wire _w3991_ ;
	wire _w3990_ ;
	wire _w3989_ ;
	wire _w3988_ ;
	wire _w3987_ ;
	wire _w3986_ ;
	wire _w3985_ ;
	wire _w3984_ ;
	wire _w3983_ ;
	wire _w3982_ ;
	wire _w3981_ ;
	wire _w3980_ ;
	wire _w3979_ ;
	wire _w3978_ ;
	wire _w3977_ ;
	wire _w3976_ ;
	wire _w3975_ ;
	wire _w3974_ ;
	wire _w3973_ ;
	wire _w3972_ ;
	wire _w3971_ ;
	wire _w3970_ ;
	wire _w3969_ ;
	wire _w3968_ ;
	wire _w3967_ ;
	wire _w3966_ ;
	wire _w3965_ ;
	wire _w3964_ ;
	wire _w3963_ ;
	wire _w3962_ ;
	wire _w3961_ ;
	wire _w3960_ ;
	wire _w3959_ ;
	wire _w3958_ ;
	wire _w3957_ ;
	wire _w3956_ ;
	wire _w3955_ ;
	wire _w3954_ ;
	wire _w3953_ ;
	wire _w3952_ ;
	wire _w3951_ ;
	wire _w3950_ ;
	wire _w3949_ ;
	wire _w3948_ ;
	wire _w3947_ ;
	wire _w3946_ ;
	wire _w3945_ ;
	wire _w3944_ ;
	wire _w3943_ ;
	wire _w3942_ ;
	wire _w3941_ ;
	wire _w3940_ ;
	wire _w3939_ ;
	wire _w3938_ ;
	wire _w3937_ ;
	wire _w3936_ ;
	wire _w3935_ ;
	wire _w3934_ ;
	wire _w3933_ ;
	wire _w3932_ ;
	wire _w3931_ ;
	wire _w3930_ ;
	wire _w3929_ ;
	wire _w3928_ ;
	wire _w3927_ ;
	wire _w3926_ ;
	wire _w3925_ ;
	wire _w3924_ ;
	wire _w3923_ ;
	wire _w3922_ ;
	wire _w3921_ ;
	wire _w3920_ ;
	wire _w3919_ ;
	wire _w3918_ ;
	wire _w3917_ ;
	wire _w3916_ ;
	wire _w3915_ ;
	wire _w3914_ ;
	wire _w3913_ ;
	wire _w3912_ ;
	wire _w3911_ ;
	wire _w3910_ ;
	wire _w3909_ ;
	wire _w3908_ ;
	wire _w3907_ ;
	wire _w3906_ ;
	wire _w3905_ ;
	wire _w3904_ ;
	wire _w3903_ ;
	wire _w3902_ ;
	wire _w3901_ ;
	wire _w3900_ ;
	wire _w3899_ ;
	wire _w3898_ ;
	wire _w3897_ ;
	wire _w3896_ ;
	wire _w3895_ ;
	wire _w3894_ ;
	wire _w3893_ ;
	wire _w3892_ ;
	wire _w3891_ ;
	wire _w3890_ ;
	wire _w3889_ ;
	wire _w3888_ ;
	wire _w3887_ ;
	wire _w3886_ ;
	wire _w3885_ ;
	wire _w3884_ ;
	wire _w3883_ ;
	wire _w3882_ ;
	wire _w3881_ ;
	wire _w3880_ ;
	wire _w3879_ ;
	wire _w3878_ ;
	wire _w3877_ ;
	wire _w3876_ ;
	wire _w3875_ ;
	wire _w3874_ ;
	wire _w3873_ ;
	wire _w3872_ ;
	wire _w3871_ ;
	wire _w3870_ ;
	wire _w3869_ ;
	wire _w3868_ ;
	wire _w3867_ ;
	wire _w3866_ ;
	wire _w3865_ ;
	wire _w3864_ ;
	wire _w3863_ ;
	wire _w3862_ ;
	wire _w3861_ ;
	wire _w3860_ ;
	wire _w3859_ ;
	wire _w3858_ ;
	wire _w3857_ ;
	wire _w3856_ ;
	wire _w3855_ ;
	wire _w3854_ ;
	wire _w3853_ ;
	wire _w3852_ ;
	wire _w3851_ ;
	wire _w3850_ ;
	wire _w3849_ ;
	wire _w3848_ ;
	wire _w3847_ ;
	wire _w3846_ ;
	wire _w3845_ ;
	wire _w3844_ ;
	wire _w3843_ ;
	wire _w3842_ ;
	wire _w3841_ ;
	wire _w3840_ ;
	wire _w3839_ ;
	wire _w3838_ ;
	wire _w3837_ ;
	wire _w3836_ ;
	wire _w3835_ ;
	wire _w3834_ ;
	wire _w3833_ ;
	wire _w3832_ ;
	wire _w3831_ ;
	wire _w3830_ ;
	wire _w3829_ ;
	wire _w3828_ ;
	wire _w3827_ ;
	wire _w3826_ ;
	wire _w3825_ ;
	wire _w3824_ ;
	wire _w3823_ ;
	wire _w3822_ ;
	wire _w3821_ ;
	wire _w3820_ ;
	wire _w3819_ ;
	wire _w3818_ ;
	wire _w3817_ ;
	wire _w3816_ ;
	wire _w3815_ ;
	wire _w3814_ ;
	wire _w3813_ ;
	wire _w3812_ ;
	wire _w3811_ ;
	wire _w3810_ ;
	wire _w3809_ ;
	wire _w3808_ ;
	wire _w3807_ ;
	wire _w3806_ ;
	wire _w3805_ ;
	wire _w3804_ ;
	wire _w3803_ ;
	wire _w3802_ ;
	wire _w3801_ ;
	wire _w3800_ ;
	wire _w3799_ ;
	wire _w3798_ ;
	wire _w3797_ ;
	wire _w3796_ ;
	wire _w3795_ ;
	wire _w3794_ ;
	wire _w3793_ ;
	wire _w3792_ ;
	wire _w3791_ ;
	wire _w3790_ ;
	wire _w3789_ ;
	wire _w3788_ ;
	wire _w3787_ ;
	wire _w3786_ ;
	wire _w3785_ ;
	wire _w3784_ ;
	wire _w3783_ ;
	wire _w3782_ ;
	wire _w3781_ ;
	wire _w3780_ ;
	wire _w3779_ ;
	wire _w3778_ ;
	wire _w3777_ ;
	wire _w3776_ ;
	wire _w3775_ ;
	wire _w3774_ ;
	wire _w3773_ ;
	wire _w3772_ ;
	wire _w3771_ ;
	wire _w3770_ ;
	wire _w3769_ ;
	wire _w3768_ ;
	wire _w3767_ ;
	wire _w3766_ ;
	wire _w3765_ ;
	wire _w3764_ ;
	wire _w3763_ ;
	wire _w3762_ ;
	wire _w3761_ ;
	wire _w3760_ ;
	wire _w3759_ ;
	wire _w3758_ ;
	wire _w3757_ ;
	wire _w3756_ ;
	wire _w3755_ ;
	wire _w3754_ ;
	wire _w3753_ ;
	wire _w3752_ ;
	wire _w3751_ ;
	wire _w3750_ ;
	wire _w3749_ ;
	wire _w3748_ ;
	wire _w3747_ ;
	wire _w3746_ ;
	wire _w3745_ ;
	wire _w3744_ ;
	wire _w3743_ ;
	wire _w3742_ ;
	wire _w3741_ ;
	wire _w3740_ ;
	wire _w3739_ ;
	wire _w3738_ ;
	wire _w3737_ ;
	wire _w3736_ ;
	wire _w3735_ ;
	wire _w3734_ ;
	wire _w3733_ ;
	wire _w3732_ ;
	wire _w3731_ ;
	wire _w3730_ ;
	wire _w3729_ ;
	wire _w3728_ ;
	wire _w3727_ ;
	wire _w3726_ ;
	wire _w3725_ ;
	wire _w3724_ ;
	wire _w3723_ ;
	wire _w3722_ ;
	wire _w3721_ ;
	wire _w3720_ ;
	wire _w3719_ ;
	wire _w3718_ ;
	wire _w3717_ ;
	wire _w3716_ ;
	wire _w3715_ ;
	wire _w3714_ ;
	wire _w3713_ ;
	wire _w3712_ ;
	wire _w3711_ ;
	wire _w3710_ ;
	wire _w3709_ ;
	wire _w3708_ ;
	wire _w3707_ ;
	wire _w3706_ ;
	wire _w3705_ ;
	wire _w3704_ ;
	wire _w3703_ ;
	wire _w3702_ ;
	wire _w3701_ ;
	wire _w3700_ ;
	wire _w3699_ ;
	wire _w3698_ ;
	wire _w3697_ ;
	wire _w3696_ ;
	wire _w3695_ ;
	wire _w3694_ ;
	wire _w3693_ ;
	wire _w3692_ ;
	wire _w3691_ ;
	wire _w3690_ ;
	wire _w3689_ ;
	wire _w3688_ ;
	wire _w3687_ ;
	wire _w3686_ ;
	wire _w3685_ ;
	wire _w3684_ ;
	wire _w3683_ ;
	wire _w3682_ ;
	wire _w3681_ ;
	wire _w3680_ ;
	wire _w3679_ ;
	wire _w3678_ ;
	wire _w3677_ ;
	wire _w3676_ ;
	wire _w3675_ ;
	wire _w3674_ ;
	wire _w3673_ ;
	wire _w3672_ ;
	wire _w3671_ ;
	wire _w3670_ ;
	wire _w3669_ ;
	wire _w3668_ ;
	wire _w3667_ ;
	wire _w3666_ ;
	wire _w3665_ ;
	wire _w3664_ ;
	wire _w3663_ ;
	wire _w3662_ ;
	wire _w3661_ ;
	wire _w3660_ ;
	wire _w3659_ ;
	wire _w3658_ ;
	wire _w3657_ ;
	wire _w3656_ ;
	wire _w3655_ ;
	wire _w3654_ ;
	wire _w3653_ ;
	wire _w3652_ ;
	wire _w3651_ ;
	wire _w3650_ ;
	wire _w3649_ ;
	wire _w3648_ ;
	wire _w3647_ ;
	wire _w3646_ ;
	wire _w3645_ ;
	wire _w3644_ ;
	wire _w3643_ ;
	wire _w3642_ ;
	wire _w3641_ ;
	wire _w3640_ ;
	wire _w3639_ ;
	wire _w3638_ ;
	wire _w3637_ ;
	wire _w3636_ ;
	wire _w3635_ ;
	wire _w3634_ ;
	wire _w3633_ ;
	wire _w3632_ ;
	wire _w3631_ ;
	wire _w3630_ ;
	wire _w3629_ ;
	wire _w3628_ ;
	wire _w3627_ ;
	wire _w3626_ ;
	wire _w3625_ ;
	wire _w3624_ ;
	wire _w3623_ ;
	wire _w3622_ ;
	wire _w3621_ ;
	wire _w3620_ ;
	wire _w3619_ ;
	wire _w3618_ ;
	wire _w3617_ ;
	wire _w3616_ ;
	wire _w3615_ ;
	wire _w3614_ ;
	wire _w3613_ ;
	wire _w3612_ ;
	wire _w3611_ ;
	wire _w3610_ ;
	wire _w3609_ ;
	wire _w3608_ ;
	wire _w3607_ ;
	wire _w3606_ ;
	wire _w3605_ ;
	wire _w3604_ ;
	wire _w3603_ ;
	wire _w3602_ ;
	wire _w3601_ ;
	wire _w3600_ ;
	wire _w3599_ ;
	wire _w3598_ ;
	wire _w3597_ ;
	wire _w3596_ ;
	wire _w3595_ ;
	wire _w3594_ ;
	wire _w3593_ ;
	wire _w3592_ ;
	wire _w3591_ ;
	wire _w3590_ ;
	wire _w3589_ ;
	wire _w3588_ ;
	wire _w3587_ ;
	wire _w3586_ ;
	wire _w3585_ ;
	wire _w3584_ ;
	wire _w3583_ ;
	wire _w3582_ ;
	wire _w3581_ ;
	wire _w3580_ ;
	wire _w3579_ ;
	wire _w3578_ ;
	wire _w3577_ ;
	wire _w3576_ ;
	wire _w3575_ ;
	wire _w3574_ ;
	wire _w3573_ ;
	wire _w3572_ ;
	wire _w3571_ ;
	wire _w3570_ ;
	wire _w3569_ ;
	wire _w3568_ ;
	wire _w3567_ ;
	wire _w3566_ ;
	wire _w3565_ ;
	wire _w3564_ ;
	wire _w3563_ ;
	wire _w3562_ ;
	wire _w3561_ ;
	wire _w3560_ ;
	wire _w3559_ ;
	wire _w3558_ ;
	wire _w3557_ ;
	wire _w3556_ ;
	wire _w3555_ ;
	wire _w3554_ ;
	wire _w3553_ ;
	wire _w3552_ ;
	wire _w3551_ ;
	wire _w3550_ ;
	wire _w3549_ ;
	wire _w3548_ ;
	wire _w3547_ ;
	wire _w3546_ ;
	wire _w3545_ ;
	wire _w3544_ ;
	wire _w3543_ ;
	wire _w3542_ ;
	wire _w3541_ ;
	wire _w3540_ ;
	wire _w3539_ ;
	wire _w3538_ ;
	wire _w3537_ ;
	wire _w3536_ ;
	wire _w3535_ ;
	wire _w3534_ ;
	wire _w3533_ ;
	wire _w3532_ ;
	wire _w3531_ ;
	wire _w3530_ ;
	wire _w3529_ ;
	wire _w3528_ ;
	wire _w3527_ ;
	wire _w3526_ ;
	wire _w3525_ ;
	wire _w3524_ ;
	wire _w3523_ ;
	wire _w3522_ ;
	wire _w3521_ ;
	wire _w3520_ ;
	wire _w3519_ ;
	wire _w3518_ ;
	wire _w3517_ ;
	wire _w3516_ ;
	wire _w3515_ ;
	wire _w3514_ ;
	wire _w3513_ ;
	wire _w3512_ ;
	wire _w3511_ ;
	wire _w3510_ ;
	wire _w3509_ ;
	wire _w3508_ ;
	wire _w3507_ ;
	wire _w3506_ ;
	wire _w3505_ ;
	wire _w3504_ ;
	wire _w3503_ ;
	wire _w3502_ ;
	wire _w3501_ ;
	wire _w3500_ ;
	wire _w3499_ ;
	wire _w3498_ ;
	wire _w3497_ ;
	wire _w3496_ ;
	wire _w3495_ ;
	wire _w3494_ ;
	wire _w3493_ ;
	wire _w3492_ ;
	wire _w3491_ ;
	wire _w3490_ ;
	wire _w3489_ ;
	wire _w3488_ ;
	wire _w3487_ ;
	wire _w3486_ ;
	wire _w3485_ ;
	wire _w3484_ ;
	wire _w3483_ ;
	wire _w3482_ ;
	wire _w3481_ ;
	wire _w3480_ ;
	wire _w3479_ ;
	wire _w3478_ ;
	wire _w3477_ ;
	wire _w3476_ ;
	wire _w3475_ ;
	wire _w3474_ ;
	wire _w3473_ ;
	wire _w3472_ ;
	wire _w3471_ ;
	wire _w3470_ ;
	wire _w3469_ ;
	wire _w3468_ ;
	wire _w3467_ ;
	wire _w3466_ ;
	wire _w3465_ ;
	wire _w3464_ ;
	wire _w3463_ ;
	wire _w3462_ ;
	wire _w3461_ ;
	wire _w3460_ ;
	wire _w3459_ ;
	wire _w3458_ ;
	wire _w3457_ ;
	wire _w3456_ ;
	wire _w3455_ ;
	wire _w3454_ ;
	wire _w3453_ ;
	wire _w3452_ ;
	wire _w3451_ ;
	wire _w3450_ ;
	wire _w3449_ ;
	wire _w3448_ ;
	wire _w3447_ ;
	wire _w3446_ ;
	wire _w3445_ ;
	wire _w3444_ ;
	wire _w3443_ ;
	wire _w3442_ ;
	wire _w3441_ ;
	wire _w3440_ ;
	wire _w3439_ ;
	wire _w3438_ ;
	wire _w3437_ ;
	wire _w3436_ ;
	wire _w3435_ ;
	wire _w3434_ ;
	wire _w3433_ ;
	wire _w3432_ ;
	wire _w3431_ ;
	wire _w3430_ ;
	wire _w3429_ ;
	wire _w3428_ ;
	wire _w3427_ ;
	wire _w3426_ ;
	wire _w3425_ ;
	wire _w3424_ ;
	wire _w3423_ ;
	wire _w3422_ ;
	wire _w3421_ ;
	wire _w3420_ ;
	wire _w3419_ ;
	wire _w3418_ ;
	wire _w3417_ ;
	wire _w3416_ ;
	wire _w3415_ ;
	wire _w3414_ ;
	wire _w3413_ ;
	wire _w3412_ ;
	wire _w3411_ ;
	wire _w3410_ ;
	wire _w3409_ ;
	wire _w3408_ ;
	wire _w3407_ ;
	wire _w3406_ ;
	wire _w3405_ ;
	wire _w3404_ ;
	wire _w3403_ ;
	wire _w3402_ ;
	wire _w3401_ ;
	wire _w3400_ ;
	wire _w3399_ ;
	wire _w3398_ ;
	wire _w3397_ ;
	wire _w3396_ ;
	wire _w3395_ ;
	wire _w3394_ ;
	wire _w3393_ ;
	wire _w3392_ ;
	wire _w3391_ ;
	wire _w3390_ ;
	wire _w3389_ ;
	wire _w3388_ ;
	wire _w3387_ ;
	wire _w3386_ ;
	wire _w3385_ ;
	wire _w3384_ ;
	wire _w3383_ ;
	wire _w3382_ ;
	wire _w3381_ ;
	wire _w3380_ ;
	wire _w3379_ ;
	wire _w3378_ ;
	wire _w3377_ ;
	wire _w3376_ ;
	wire _w3375_ ;
	wire _w3374_ ;
	wire _w3373_ ;
	wire _w3372_ ;
	wire _w3371_ ;
	wire _w3370_ ;
	wire _w3369_ ;
	wire _w3368_ ;
	wire _w3367_ ;
	wire _w3366_ ;
	wire _w3365_ ;
	wire _w3364_ ;
	wire _w3363_ ;
	wire _w3362_ ;
	wire _w3361_ ;
	wire _w3360_ ;
	wire _w3359_ ;
	wire _w3358_ ;
	wire _w3357_ ;
	wire _w3356_ ;
	wire _w3355_ ;
	wire _w3354_ ;
	wire _w3353_ ;
	wire _w3352_ ;
	wire _w3351_ ;
	wire _w3350_ ;
	wire _w3349_ ;
	wire _w3348_ ;
	wire _w3347_ ;
	wire _w3346_ ;
	wire _w3345_ ;
	wire _w3344_ ;
	wire _w3343_ ;
	wire _w3342_ ;
	wire _w3341_ ;
	wire _w3340_ ;
	wire _w3339_ ;
	wire _w3338_ ;
	wire _w3337_ ;
	wire _w3336_ ;
	wire _w3335_ ;
	wire _w3334_ ;
	wire _w3333_ ;
	wire _w3332_ ;
	wire _w3331_ ;
	wire _w3330_ ;
	wire _w3329_ ;
	wire _w3328_ ;
	wire _w3327_ ;
	wire _w3326_ ;
	wire _w3325_ ;
	wire _w3324_ ;
	wire _w3323_ ;
	wire _w3322_ ;
	wire _w3321_ ;
	wire _w3320_ ;
	wire _w3319_ ;
	wire _w3318_ ;
	wire _w3317_ ;
	wire _w3316_ ;
	wire _w3315_ ;
	wire _w3314_ ;
	wire _w3313_ ;
	wire _w3312_ ;
	wire _w3311_ ;
	wire _w3310_ ;
	wire _w3309_ ;
	wire _w3308_ ;
	wire _w3307_ ;
	wire _w3306_ ;
	wire _w3305_ ;
	wire _w3304_ ;
	wire _w3303_ ;
	wire _w3302_ ;
	wire _w3301_ ;
	wire _w3300_ ;
	wire _w3299_ ;
	wire _w3298_ ;
	wire _w3297_ ;
	wire _w3296_ ;
	wire _w3295_ ;
	wire _w3294_ ;
	wire _w3293_ ;
	wire _w3292_ ;
	wire _w3291_ ;
	wire _w3290_ ;
	wire _w3289_ ;
	wire _w3288_ ;
	wire _w3287_ ;
	wire _w3286_ ;
	wire _w3285_ ;
	wire _w3284_ ;
	wire _w3283_ ;
	wire _w3282_ ;
	wire _w3281_ ;
	wire _w3280_ ;
	wire _w3279_ ;
	wire _w3278_ ;
	wire _w3277_ ;
	wire _w3276_ ;
	wire _w3275_ ;
	wire _w3274_ ;
	wire _w3273_ ;
	wire _w3272_ ;
	wire _w3271_ ;
	wire _w3270_ ;
	wire _w3269_ ;
	wire _w3268_ ;
	wire _w3267_ ;
	wire _w3266_ ;
	wire _w3265_ ;
	wire _w3264_ ;
	wire _w3263_ ;
	wire _w3262_ ;
	wire _w3261_ ;
	wire _w3260_ ;
	wire _w3259_ ;
	wire _w3258_ ;
	wire _w3257_ ;
	wire _w3256_ ;
	wire _w3255_ ;
	wire _w3254_ ;
	wire _w3253_ ;
	wire _w3252_ ;
	wire _w3251_ ;
	wire _w3250_ ;
	wire _w3249_ ;
	wire _w3248_ ;
	wire _w3247_ ;
	wire _w3246_ ;
	wire _w3245_ ;
	wire _w3244_ ;
	wire _w3243_ ;
	wire _w3242_ ;
	wire _w3241_ ;
	wire _w3240_ ;
	wire _w3239_ ;
	wire _w3238_ ;
	wire _w3237_ ;
	wire _w3236_ ;
	wire _w3235_ ;
	wire _w3234_ ;
	wire _w3233_ ;
	wire _w3232_ ;
	wire _w3231_ ;
	wire _w3230_ ;
	wire _w3229_ ;
	wire _w3228_ ;
	wire _w3227_ ;
	wire _w3226_ ;
	wire _w3225_ ;
	wire _w3224_ ;
	wire _w3223_ ;
	wire _w3222_ ;
	wire _w3221_ ;
	wire _w3220_ ;
	wire _w3219_ ;
	wire _w3218_ ;
	wire _w3217_ ;
	wire _w3216_ ;
	wire _w3215_ ;
	wire _w3214_ ;
	wire _w3213_ ;
	wire _w3212_ ;
	wire _w3211_ ;
	wire _w3210_ ;
	wire _w3209_ ;
	wire _w3208_ ;
	wire _w3207_ ;
	wire _w3206_ ;
	wire _w3205_ ;
	wire _w3204_ ;
	wire _w3203_ ;
	wire _w3202_ ;
	wire _w3201_ ;
	wire _w3200_ ;
	wire _w3199_ ;
	wire _w3198_ ;
	wire _w3197_ ;
	wire _w3196_ ;
	wire _w3195_ ;
	wire _w3194_ ;
	wire _w3193_ ;
	wire _w3192_ ;
	wire _w3191_ ;
	wire _w3190_ ;
	wire _w3189_ ;
	wire _w3188_ ;
	wire _w3187_ ;
	wire _w3186_ ;
	wire _w3185_ ;
	wire _w3184_ ;
	wire _w3183_ ;
	wire _w3182_ ;
	wire _w3181_ ;
	wire _w3180_ ;
	wire _w3179_ ;
	wire _w3178_ ;
	wire _w3177_ ;
	wire _w3176_ ;
	wire _w3175_ ;
	wire _w3174_ ;
	wire _w3173_ ;
	wire _w3172_ ;
	wire _w3171_ ;
	wire _w3170_ ;
	wire _w3169_ ;
	wire _w3168_ ;
	wire _w3167_ ;
	wire _w3166_ ;
	wire _w3165_ ;
	wire _w3164_ ;
	wire _w3163_ ;
	wire _w3162_ ;
	wire _w3161_ ;
	wire _w3160_ ;
	wire _w3159_ ;
	wire _w3158_ ;
	wire _w3157_ ;
	wire _w3156_ ;
	wire _w3155_ ;
	wire _w3154_ ;
	wire _w3153_ ;
	wire _w3152_ ;
	wire _w3151_ ;
	wire _w3150_ ;
	wire _w3149_ ;
	wire _w3148_ ;
	wire _w3147_ ;
	wire _w3146_ ;
	wire _w3145_ ;
	wire _w3144_ ;
	wire _w3143_ ;
	wire _w3142_ ;
	wire _w3141_ ;
	wire _w3140_ ;
	wire _w3139_ ;
	wire _w3138_ ;
	wire _w3137_ ;
	wire _w3136_ ;
	wire _w3135_ ;
	wire _w3134_ ;
	wire _w3133_ ;
	wire _w3132_ ;
	wire _w3131_ ;
	wire _w3130_ ;
	wire _w3129_ ;
	wire _w3128_ ;
	wire _w3127_ ;
	wire _w3126_ ;
	wire _w3125_ ;
	wire _w3124_ ;
	wire _w3123_ ;
	wire _w3122_ ;
	wire _w3121_ ;
	wire _w3120_ ;
	wire _w3119_ ;
	wire _w3118_ ;
	wire _w3117_ ;
	wire _w3116_ ;
	wire _w3115_ ;
	wire _w3114_ ;
	wire _w3113_ ;
	wire _w3112_ ;
	wire _w3111_ ;
	wire _w3110_ ;
	wire _w3109_ ;
	wire _w3108_ ;
	wire _w3107_ ;
	wire _w3106_ ;
	wire _w3105_ ;
	wire _w3104_ ;
	wire _w3103_ ;
	wire _w3102_ ;
	wire _w3101_ ;
	wire _w3100_ ;
	wire _w3099_ ;
	wire _w3098_ ;
	wire _w3097_ ;
	wire _w3096_ ;
	wire _w3095_ ;
	wire _w3094_ ;
	wire _w3093_ ;
	wire _w3092_ ;
	wire _w3091_ ;
	wire _w3090_ ;
	wire _w3089_ ;
	wire _w3088_ ;
	wire _w3087_ ;
	wire _w3086_ ;
	wire _w3085_ ;
	wire _w3084_ ;
	wire _w3083_ ;
	wire _w3082_ ;
	wire _w3081_ ;
	wire _w3080_ ;
	wire _w3079_ ;
	wire _w3078_ ;
	wire _w3077_ ;
	wire _w3076_ ;
	wire _w3075_ ;
	wire _w3074_ ;
	wire _w3073_ ;
	wire _w3072_ ;
	wire _w3071_ ;
	wire _w3070_ ;
	wire _w3069_ ;
	wire _w3068_ ;
	wire _w3067_ ;
	wire _w3066_ ;
	wire _w3065_ ;
	wire _w3064_ ;
	wire _w3063_ ;
	wire _w3062_ ;
	wire _w3061_ ;
	wire _w3060_ ;
	wire _w3059_ ;
	wire _w3058_ ;
	wire _w3057_ ;
	wire _w3056_ ;
	wire _w3055_ ;
	wire _w3054_ ;
	wire _w3053_ ;
	wire _w3052_ ;
	wire _w3051_ ;
	wire _w3050_ ;
	wire _w3049_ ;
	wire _w3048_ ;
	wire _w3047_ ;
	wire _w3046_ ;
	wire _w3045_ ;
	wire _w3044_ ;
	wire _w3043_ ;
	wire _w3042_ ;
	wire _w3041_ ;
	wire _w3040_ ;
	wire _w3039_ ;
	wire _w3038_ ;
	wire _w3037_ ;
	wire _w3036_ ;
	wire _w3035_ ;
	wire _w3034_ ;
	wire _w3033_ ;
	wire _w3032_ ;
	wire _w3031_ ;
	wire _w3030_ ;
	wire _w3029_ ;
	wire _w3028_ ;
	wire _w3027_ ;
	wire _w3026_ ;
	wire _w3025_ ;
	wire _w3024_ ;
	wire _w3023_ ;
	wire _w3022_ ;
	wire _w3021_ ;
	wire _w3020_ ;
	wire _w3019_ ;
	wire _w3018_ ;
	wire _w3017_ ;
	wire _w3016_ ;
	wire _w3015_ ;
	wire _w3014_ ;
	wire _w3013_ ;
	wire _w3012_ ;
	wire _w3011_ ;
	wire _w3010_ ;
	wire _w3009_ ;
	wire _w3008_ ;
	wire _w3007_ ;
	wire _w3006_ ;
	wire _w3005_ ;
	wire _w3004_ ;
	wire _w3003_ ;
	wire _w3002_ ;
	wire _w3001_ ;
	wire _w3000_ ;
	wire _w2999_ ;
	wire _w2998_ ;
	wire _w2997_ ;
	wire _w2996_ ;
	wire _w2995_ ;
	wire _w2994_ ;
	wire _w2993_ ;
	wire _w2992_ ;
	wire _w2991_ ;
	wire _w2990_ ;
	wire _w2989_ ;
	wire _w2988_ ;
	wire _w2987_ ;
	wire _w2986_ ;
	wire _w2985_ ;
	wire _w2984_ ;
	wire _w2983_ ;
	wire _w2982_ ;
	wire _w2981_ ;
	wire _w2980_ ;
	wire _w2979_ ;
	wire _w2978_ ;
	wire _w2977_ ;
	wire _w2976_ ;
	wire _w2975_ ;
	wire _w2974_ ;
	wire _w2973_ ;
	wire _w2972_ ;
	wire _w2971_ ;
	wire _w2970_ ;
	wire _w2969_ ;
	wire _w2968_ ;
	wire _w2967_ ;
	wire _w2966_ ;
	wire _w2965_ ;
	wire _w2964_ ;
	wire _w2963_ ;
	wire _w2962_ ;
	wire _w2961_ ;
	wire _w2960_ ;
	wire _w2959_ ;
	wire _w2958_ ;
	wire _w2957_ ;
	wire _w2956_ ;
	wire _w2955_ ;
	wire _w2954_ ;
	wire _w2953_ ;
	wire _w2952_ ;
	wire _w2951_ ;
	wire _w2950_ ;
	wire _w2949_ ;
	wire _w2948_ ;
	wire _w2947_ ;
	wire _w2946_ ;
	wire _w2945_ ;
	wire _w2944_ ;
	wire _w2943_ ;
	wire _w2942_ ;
	wire _w2941_ ;
	wire _w2940_ ;
	wire _w2939_ ;
	wire _w2938_ ;
	wire _w2937_ ;
	wire _w2936_ ;
	wire _w2935_ ;
	wire _w2934_ ;
	wire _w2933_ ;
	wire _w2932_ ;
	wire _w2931_ ;
	wire _w2930_ ;
	wire _w2929_ ;
	wire _w2928_ ;
	wire _w2927_ ;
	wire _w2926_ ;
	wire _w2925_ ;
	wire _w2924_ ;
	wire _w2923_ ;
	wire _w2922_ ;
	wire _w2921_ ;
	wire _w2920_ ;
	wire _w2919_ ;
	wire _w2918_ ;
	wire _w2917_ ;
	wire _w2916_ ;
	wire _w2915_ ;
	wire _w2914_ ;
	wire _w2913_ ;
	wire _w2912_ ;
	wire _w2911_ ;
	wire _w2910_ ;
	wire _w2909_ ;
	wire _w2908_ ;
	wire _w2907_ ;
	wire _w2906_ ;
	wire _w2905_ ;
	wire _w2904_ ;
	wire _w2903_ ;
	wire _w2902_ ;
	wire _w2901_ ;
	wire _w2900_ ;
	wire _w2899_ ;
	wire _w2898_ ;
	wire _w2897_ ;
	wire _w2896_ ;
	wire _w2895_ ;
	wire _w2894_ ;
	wire _w2893_ ;
	wire _w2892_ ;
	wire _w2891_ ;
	wire _w2890_ ;
	wire _w2889_ ;
	wire _w2888_ ;
	wire _w2887_ ;
	wire _w2886_ ;
	wire _w2885_ ;
	wire _w2884_ ;
	wire _w2883_ ;
	wire _w2882_ ;
	wire _w2881_ ;
	wire _w2880_ ;
	wire _w2879_ ;
	wire _w2878_ ;
	wire _w2877_ ;
	wire _w2876_ ;
	wire _w2875_ ;
	wire _w2874_ ;
	wire _w2873_ ;
	wire _w2872_ ;
	wire _w2871_ ;
	wire _w2870_ ;
	wire _w2869_ ;
	wire _w2868_ ;
	wire _w2867_ ;
	wire _w2866_ ;
	wire _w2865_ ;
	wire _w2864_ ;
	wire _w2863_ ;
	wire _w2862_ ;
	wire _w2861_ ;
	wire _w2860_ ;
	wire _w2859_ ;
	wire _w2858_ ;
	wire _w2857_ ;
	wire _w2856_ ;
	wire _w2855_ ;
	wire _w2854_ ;
	wire _w2853_ ;
	wire _w2852_ ;
	wire _w2851_ ;
	wire _w2850_ ;
	wire _w2849_ ;
	wire _w2848_ ;
	wire _w2847_ ;
	wire _w2846_ ;
	wire _w2845_ ;
	wire _w2844_ ;
	wire _w2843_ ;
	wire _w2842_ ;
	wire _w2841_ ;
	wire _w2840_ ;
	wire _w2839_ ;
	wire _w2838_ ;
	wire _w2837_ ;
	wire _w2836_ ;
	wire _w2835_ ;
	wire _w2834_ ;
	wire _w2833_ ;
	wire _w2832_ ;
	wire _w2831_ ;
	wire _w2830_ ;
	wire _w2829_ ;
	wire _w2828_ ;
	wire _w2827_ ;
	wire _w2826_ ;
	wire _w2825_ ;
	wire _w2824_ ;
	wire _w2823_ ;
	wire _w2822_ ;
	wire _w2821_ ;
	wire _w2820_ ;
	wire _w2819_ ;
	wire _w2818_ ;
	wire _w2817_ ;
	wire _w2816_ ;
	wire _w2815_ ;
	wire _w2814_ ;
	wire _w2813_ ;
	wire _w2812_ ;
	wire _w2811_ ;
	wire _w2810_ ;
	wire _w1561_ ;
	wire _w1560_ ;
	wire _w1559_ ;
	wire _w1558_ ;
	wire _w1557_ ;
	wire _w1556_ ;
	wire _w1555_ ;
	wire _w1554_ ;
	wire _w1553_ ;
	wire _w1552_ ;
	wire _w1551_ ;
	wire _w1550_ ;
	wire _w1549_ ;
	wire _w1548_ ;
	wire _w1547_ ;
	wire _w1546_ ;
	wire _w1545_ ;
	wire _w1544_ ;
	wire _w1543_ ;
	wire _w1542_ ;
	wire _w1541_ ;
	wire _w1540_ ;
	wire _w1539_ ;
	wire _w1538_ ;
	wire _w1537_ ;
	wire _w1536_ ;
	wire _w1535_ ;
	wire _w1534_ ;
	wire _w1533_ ;
	wire _w1532_ ;
	wire _w1531_ ;
	wire _w1530_ ;
	wire _w1529_ ;
	wire _w1528_ ;
	wire _w1527_ ;
	wire _w1526_ ;
	wire _w1525_ ;
	wire _w1524_ ;
	wire _w1523_ ;
	wire _w1522_ ;
	wire _w1521_ ;
	wire _w1520_ ;
	wire _w1519_ ;
	wire _w1518_ ;
	wire _w1517_ ;
	wire _w1516_ ;
	wire _w1515_ ;
	wire _w1514_ ;
	wire _w1513_ ;
	wire _w1512_ ;
	wire _w1511_ ;
	wire _w1510_ ;
	wire _w1509_ ;
	wire _w1508_ ;
	wire _w1507_ ;
	wire _w1506_ ;
	wire _w1505_ ;
	wire _w1504_ ;
	wire _w1503_ ;
	wire _w1502_ ;
	wire _w1501_ ;
	wire _w1500_ ;
	wire _w1499_ ;
	wire _w1498_ ;
	wire _w1497_ ;
	wire _w1496_ ;
	wire _w1495_ ;
	wire _w1494_ ;
	wire _w1493_ ;
	wire _w1492_ ;
	wire _w1491_ ;
	wire _w1490_ ;
	wire _w1489_ ;
	wire _w1488_ ;
	wire _w1487_ ;
	wire _w1486_ ;
	wire _w1485_ ;
	wire _w1484_ ;
	wire _w1483_ ;
	wire _w1482_ ;
	wire _w1481_ ;
	wire _w1480_ ;
	wire _w1479_ ;
	wire _w1478_ ;
	wire _w1477_ ;
	wire _w1476_ ;
	wire _w1475_ ;
	wire _w1474_ ;
	wire _w1473_ ;
	wire _w1472_ ;
	wire _w1471_ ;
	wire _w1470_ ;
	wire _w1469_ ;
	wire _w1468_ ;
	wire _w1467_ ;
	wire _w1466_ ;
	wire _w1465_ ;
	wire _w1464_ ;
	wire _w1463_ ;
	wire _w1462_ ;
	wire _w1461_ ;
	wire _w1460_ ;
	wire _w1459_ ;
	wire _w1458_ ;
	wire _w1457_ ;
	wire _w1456_ ;
	wire _w1455_ ;
	wire _w1454_ ;
	wire _w1453_ ;
	wire _w1452_ ;
	wire _w1451_ ;
	wire _w1450_ ;
	wire _w1449_ ;
	wire _w1448_ ;
	wire _w1447_ ;
	wire _w1446_ ;
	wire _w1445_ ;
	wire _w1444_ ;
	wire _w1443_ ;
	wire _w1442_ ;
	wire _w1441_ ;
	wire _w1440_ ;
	wire _w1439_ ;
	wire _w1438_ ;
	wire _w1437_ ;
	wire _w1436_ ;
	wire _w1435_ ;
	wire _w1434_ ;
	wire _w1433_ ;
	wire _w1432_ ;
	wire _w1431_ ;
	wire _w1430_ ;
	wire _w1429_ ;
	wire _w1428_ ;
	wire _w1427_ ;
	wire _w1426_ ;
	wire _w1425_ ;
	wire _w1424_ ;
	wire _w1423_ ;
	wire _w1422_ ;
	wire _w1421_ ;
	wire _w1420_ ;
	wire _w1419_ ;
	wire _w1418_ ;
	wire _w1417_ ;
	wire _w1416_ ;
	wire _w1415_ ;
	wire _w1414_ ;
	wire _w1413_ ;
	wire _w1412_ ;
	wire _w1411_ ;
	wire _w1410_ ;
	wire _w1409_ ;
	wire _w1408_ ;
	wire _w1407_ ;
	wire _w1406_ ;
	wire _w1405_ ;
	wire _w1404_ ;
	wire _w1403_ ;
	wire _w1402_ ;
	wire _w1401_ ;
	wire _w1400_ ;
	wire _w1399_ ;
	wire _w1398_ ;
	wire _w1397_ ;
	wire _w1396_ ;
	wire _w1395_ ;
	wire _w1394_ ;
	wire _w1393_ ;
	wire _w1392_ ;
	wire _w1391_ ;
	wire _w1390_ ;
	wire _w1389_ ;
	wire _w1388_ ;
	wire _w1387_ ;
	wire _w1386_ ;
	wire _w1385_ ;
	wire _w1384_ ;
	wire _w1383_ ;
	wire _w1382_ ;
	wire _w1381_ ;
	wire _w1380_ ;
	wire _w1379_ ;
	wire _w1378_ ;
	wire _w1377_ ;
	wire _w1376_ ;
	wire _w1375_ ;
	wire _w1374_ ;
	wire _w1373_ ;
	wire _w1372_ ;
	wire _w1371_ ;
	wire _w1370_ ;
	wire _w1369_ ;
	wire _w1368_ ;
	wire _w1367_ ;
	wire _w1366_ ;
	wire _w1365_ ;
	wire _w1364_ ;
	wire _w1363_ ;
	wire _w1362_ ;
	wire _w1361_ ;
	wire _w1360_ ;
	wire _w1359_ ;
	wire _w1358_ ;
	wire _w1357_ ;
	wire _w1356_ ;
	wire _w1355_ ;
	wire _w1354_ ;
	wire _w1353_ ;
	wire _w1352_ ;
	wire _w1351_ ;
	wire _w1350_ ;
	wire _w1349_ ;
	wire _w1348_ ;
	wire _w1347_ ;
	wire _w1346_ ;
	wire _w1345_ ;
	wire _w1344_ ;
	wire _w1343_ ;
	wire _w1342_ ;
	wire _w1341_ ;
	wire _w1340_ ;
	wire _w1339_ ;
	wire _w1338_ ;
	wire _w1337_ ;
	wire _w1336_ ;
	wire _w1335_ ;
	wire _w1334_ ;
	wire _w1333_ ;
	wire _w1332_ ;
	wire _w1331_ ;
	wire _w1330_ ;
	wire _w1329_ ;
	wire _w1328_ ;
	wire _w1327_ ;
	wire _w1326_ ;
	wire _w1325_ ;
	wire _w1324_ ;
	wire _w1323_ ;
	wire _w1322_ ;
	wire _w1321_ ;
	wire _w1320_ ;
	wire _w1319_ ;
	wire _w1318_ ;
	wire _w1317_ ;
	wire _w1316_ ;
	wire _w1315_ ;
	wire _w1314_ ;
	wire _w1313_ ;
	wire _w1312_ ;
	wire _w1311_ ;
	wire _w1310_ ;
	wire _w1309_ ;
	wire _w1308_ ;
	wire _w1307_ ;
	wire _w1306_ ;
	wire _w1305_ ;
	wire _w1304_ ;
	wire _w1303_ ;
	wire _w1302_ ;
	wire _w1301_ ;
	wire _w1300_ ;
	wire _w1299_ ;
	wire _w1298_ ;
	wire _w1297_ ;
	wire _w1296_ ;
	wire _w1295_ ;
	wire _w1294_ ;
	wire _w1293_ ;
	wire _w1292_ ;
	wire _w1291_ ;
	wire _w1290_ ;
	wire _w1289_ ;
	wire _w1288_ ;
	wire _w1287_ ;
	wire _w1286_ ;
	wire _w1285_ ;
	wire _w1284_ ;
	wire _w1283_ ;
	wire _w1282_ ;
	wire _w1281_ ;
	wire _w1280_ ;
	wire _w1279_ ;
	wire _w1278_ ;
	wire _w1277_ ;
	wire _w1276_ ;
	wire _w1275_ ;
	wire _w1274_ ;
	wire _w1273_ ;
	wire _w1272_ ;
	wire _w1271_ ;
	wire _w1270_ ;
	wire _w1269_ ;
	wire _w1268_ ;
	wire _w1267_ ;
	wire _w1266_ ;
	wire _w1265_ ;
	wire _w1264_ ;
	wire _w1263_ ;
	wire _w1262_ ;
	wire _w1261_ ;
	wire _w1260_ ;
	wire _w1259_ ;
	wire _w1258_ ;
	wire _w1257_ ;
	wire _w1256_ ;
	wire _w1255_ ;
	wire _w1254_ ;
	wire _w1253_ ;
	wire _w1252_ ;
	wire _w1251_ ;
	wire _w1250_ ;
	wire _w1249_ ;
	wire _w1248_ ;
	wire _w1247_ ;
	wire _w1246_ ;
	wire _w1245_ ;
	wire _w1244_ ;
	wire _w1243_ ;
	wire _w1242_ ;
	wire _w1241_ ;
	wire _w1240_ ;
	wire _w1239_ ;
	wire _w1238_ ;
	wire _w1237_ ;
	wire _w1236_ ;
	wire _w1235_ ;
	wire _w1234_ ;
	wire _w1233_ ;
	wire _w1232_ ;
	wire _w1231_ ;
	wire _w1230_ ;
	wire _w1229_ ;
	wire _w1228_ ;
	wire _w1227_ ;
	wire _w1226_ ;
	wire _w1225_ ;
	wire _w1224_ ;
	wire _w1223_ ;
	wire _w1222_ ;
	wire _w1221_ ;
	wire _w1220_ ;
	wire _w1219_ ;
	wire _w1218_ ;
	wire _w1217_ ;
	wire _w1216_ ;
	wire _w1215_ ;
	wire _w1214_ ;
	wire _w1213_ ;
	wire _w1212_ ;
	wire _w1211_ ;
	wire _w1210_ ;
	wire _w1209_ ;
	wire _w1208_ ;
	wire _w1207_ ;
	wire _w1206_ ;
	wire _w1205_ ;
	wire _w1204_ ;
	wire _w1203_ ;
	wire _w1202_ ;
	wire _w1201_ ;
	wire _w1200_ ;
	wire _w1199_ ;
	wire _w1198_ ;
	wire _w1197_ ;
	wire _w1196_ ;
	wire _w1195_ ;
	wire _w1194_ ;
	wire _w1193_ ;
	wire _w1192_ ;
	wire _w1191_ ;
	wire _w1190_ ;
	wire _w1189_ ;
	wire _w1188_ ;
	wire _w1187_ ;
	wire _w1186_ ;
	wire _w1185_ ;
	wire _w1184_ ;
	wire _w1183_ ;
	wire _w1182_ ;
	wire _w1181_ ;
	wire _w1180_ ;
	wire _w1179_ ;
	wire _w1178_ ;
	wire _w1177_ ;
	wire _w1176_ ;
	wire _w1175_ ;
	wire _w1174_ ;
	wire _w1173_ ;
	wire _w1172_ ;
	wire _w1171_ ;
	wire _w1170_ ;
	wire _w1169_ ;
	wire _w1168_ ;
	wire _w1167_ ;
	wire _w1166_ ;
	wire _w1165_ ;
	wire _w1164_ ;
	wire _w1163_ ;
	wire _w1162_ ;
	wire _w1161_ ;
	wire _w1160_ ;
	wire _w1159_ ;
	wire _w1158_ ;
	wire _w1157_ ;
	wire _w1156_ ;
	wire _w1155_ ;
	wire _w1154_ ;
	wire _w1153_ ;
	wire _w1152_ ;
	wire _w1151_ ;
	wire _w1150_ ;
	wire _w1149_ ;
	wire _w1148_ ;
	wire _w1147_ ;
	wire _w1146_ ;
	wire _w1145_ ;
	wire _w1144_ ;
	wire _w1143_ ;
	wire _w1142_ ;
	wire _w1141_ ;
	wire _w1140_ ;
	wire _w1139_ ;
	wire _w1138_ ;
	wire _w1137_ ;
	wire _w1136_ ;
	wire _w1135_ ;
	wire _w1134_ ;
	wire _w1133_ ;
	wire _w1132_ ;
	wire _w1131_ ;
	wire _w1130_ ;
	wire _w1129_ ;
	wire _w1128_ ;
	wire _w1127_ ;
	wire _w1126_ ;
	wire _w1125_ ;
	wire _w1124_ ;
	wire _w1123_ ;
	wire _w1122_ ;
	wire _w1121_ ;
	wire _w1120_ ;
	wire _w1119_ ;
	wire _w1118_ ;
	wire _w1117_ ;
	wire _w1116_ ;
	wire _w1115_ ;
	wire _w1114_ ;
	wire _w1113_ ;
	wire _w1112_ ;
	wire _w1111_ ;
	wire _w1110_ ;
	wire _w1109_ ;
	wire _w1108_ ;
	wire _w1107_ ;
	wire _w1106_ ;
	wire _w1105_ ;
	wire _w1104_ ;
	wire _w1103_ ;
	wire _w1102_ ;
	wire _w1101_ ;
	wire _w1100_ ;
	wire _w1099_ ;
	wire _w1098_ ;
	wire _w1097_ ;
	wire _w1096_ ;
	wire _w1095_ ;
	wire _w1094_ ;
	wire _w1093_ ;
	wire _w1092_ ;
	wire _w1091_ ;
	wire _w1090_ ;
	wire _w1089_ ;
	wire _w1088_ ;
	wire _w1087_ ;
	wire _w1086_ ;
	wire _w1085_ ;
	wire _w1084_ ;
	wire _w1083_ ;
	wire _w1082_ ;
	wire _w1081_ ;
	wire _w1080_ ;
	wire _w1079_ ;
	wire _w1078_ ;
	wire _w1077_ ;
	wire _w1076_ ;
	wire _w1075_ ;
	wire _w1074_ ;
	wire _w1073_ ;
	wire _w1072_ ;
	wire _w1071_ ;
	wire _w1070_ ;
	wire _w1069_ ;
	wire _w1068_ ;
	wire _w1067_ ;
	wire _w1066_ ;
	wire _w1065_ ;
	wire _w1064_ ;
	wire _w1063_ ;
	wire _w1062_ ;
	wire _w1061_ ;
	wire _w1060_ ;
	wire _w1059_ ;
	wire _w1058_ ;
	wire _w1057_ ;
	wire _w1056_ ;
	wire _w1055_ ;
	wire _w1054_ ;
	wire _w1053_ ;
	wire _w1052_ ;
	wire _w1051_ ;
	wire _w1050_ ;
	wire _w1049_ ;
	wire _w1048_ ;
	wire _w1047_ ;
	wire _w1046_ ;
	wire _w1045_ ;
	wire _w1044_ ;
	wire _w1043_ ;
	wire _w1042_ ;
	wire _w1041_ ;
	wire _w1040_ ;
	wire _w1039_ ;
	wire _w1038_ ;
	wire _w1037_ ;
	wire _w1036_ ;
	wire _w1035_ ;
	wire _w1034_ ;
	wire _w1033_ ;
	wire _w1032_ ;
	wire _w1031_ ;
	wire _w1030_ ;
	wire _w1029_ ;
	wire _w1028_ ;
	wire _w1027_ ;
	wire _w1026_ ;
	wire _w1025_ ;
	wire _w1024_ ;
	wire _w1023_ ;
	wire _w1022_ ;
	wire _w1021_ ;
	wire _w1020_ ;
	wire _w1019_ ;
	wire _w1018_ ;
	wire _w1017_ ;
	wire _w1016_ ;
	wire _w1015_ ;
	wire _w1014_ ;
	wire _w1013_ ;
	wire _w1012_ ;
	wire _w1011_ ;
	wire _w1010_ ;
	wire _w1009_ ;
	wire _w1008_ ;
	wire _w1007_ ;
	wire _w1006_ ;
	wire _w1005_ ;
	wire _w1004_ ;
	wire _w1003_ ;
	wire _w1002_ ;
	wire _w1001_ ;
	wire _w1000_ ;
	wire _w999_ ;
	wire _w998_ ;
	wire _w997_ ;
	wire _w996_ ;
	wire _w995_ ;
	wire _w994_ ;
	wire _w709_ ;
	wire _w708_ ;
	wire _w707_ ;
	wire _w706_ ;
	wire _w705_ ;
	wire _w704_ ;
	wire _w703_ ;
	wire _w702_ ;
	wire _w701_ ;
	wire _w700_ ;
	wire _w699_ ;
	wire _w698_ ;
	wire _w697_ ;
	wire _w696_ ;
	wire _w695_ ;
	wire _w694_ ;
	wire _w693_ ;
	wire _w692_ ;
	wire _w691_ ;
	wire _w690_ ;
	wire _w689_ ;
	wire _w688_ ;
	wire _w687_ ;
	wire _w686_ ;
	wire _w685_ ;
	wire _w684_ ;
	wire _w683_ ;
	wire _w682_ ;
	wire _w681_ ;
	wire _w680_ ;
	wire _w679_ ;
	wire _w678_ ;
	wire _w677_ ;
	wire _w676_ ;
	wire _w675_ ;
	wire _w674_ ;
	wire _w673_ ;
	wire _w672_ ;
	wire _w671_ ;
	wire _w670_ ;
	wire _w669_ ;
	wire _w668_ ;
	wire _w667_ ;
	wire _w666_ ;
	wire _w665_ ;
	wire _w664_ ;
	wire _w663_ ;
	wire _w662_ ;
	wire _w661_ ;
	wire _w660_ ;
	wire _w659_ ;
	wire _w658_ ;
	wire _w657_ ;
	wire _w656_ ;
	wire _w655_ ;
	wire _w654_ ;
	wire _w653_ ;
	wire _w652_ ;
	wire _w651_ ;
	wire _w650_ ;
	wire _w649_ ;
	wire _w648_ ;
	wire _w647_ ;
	wire _w646_ ;
	wire _w645_ ;
	wire _w644_ ;
	wire _w643_ ;
	wire _w642_ ;
	wire _w641_ ;
	wire _w640_ ;
	wire _w639_ ;
	wire _w638_ ;
	wire _w637_ ;
	wire _w636_ ;
	wire _w635_ ;
	wire _w634_ ;
	wire _w633_ ;
	wire _w632_ ;
	wire _w631_ ;
	wire _w630_ ;
	wire _w629_ ;
	wire _w628_ ;
	wire _w627_ ;
	wire _w626_ ;
	wire _w625_ ;
	wire _w624_ ;
	wire _w623_ ;
	wire _w622_ ;
	wire _w621_ ;
	wire _w620_ ;
	wire _w619_ ;
	wire _w618_ ;
	wire _w617_ ;
	wire _w616_ ;
	wire _w615_ ;
	wire _w614_ ;
	wire _w613_ ;
	wire _w612_ ;
	wire _w611_ ;
	wire _w610_ ;
	wire _w609_ ;
	wire _w608_ ;
	wire _w607_ ;
	wire _w606_ ;
	wire _w605_ ;
	wire _w604_ ;
	wire _w603_ ;
	wire _w602_ ;
	wire _w601_ ;
	wire _w600_ ;
	wire _w599_ ;
	wire _w598_ ;
	wire _w597_ ;
	wire _w596_ ;
	wire _w595_ ;
	wire _w594_ ;
	wire _w593_ ;
	wire _w592_ ;
	wire _w591_ ;
	wire _w590_ ;
	wire _w589_ ;
	wire _w588_ ;
	wire _w587_ ;
	wire _w586_ ;
	wire _w585_ ;
	wire _w584_ ;
	wire _w583_ ;
	wire _w582_ ;
	wire _w581_ ;
	wire _w580_ ;
	wire _w511_ ;
	wire _w510_ ;
	wire _w509_ ;
	wire _w508_ ;
	wire _w507_ ;
	wire _w506_ ;
	wire _w505_ ;
	wire _w504_ ;
	wire _w503_ ;
	wire _w502_ ;
	wire _w501_ ;
	wire _w500_ ;
	wire _w499_ ;
	wire _w498_ ;
	wire _w497_ ;
	wire _w496_ ;
	wire _w495_ ;
	wire _w494_ ;
	wire _w493_ ;
	wire _w492_ ;
	wire _w491_ ;
	wire _w490_ ;
	wire _w489_ ;
	wire _w488_ ;
	wire _w487_ ;
	wire _w486_ ;
	wire _w485_ ;
	wire _w484_ ;
	wire _w483_ ;
	wire _w482_ ;
	wire _w465_ ;
	wire _w464_ ;
	wire _w463_ ;
	wire _w462_ ;
	wire _w461_ ;
	wire _w460_ ;
	wire _w459_ ;
	wire _w458_ ;
	wire _w457_ ;
	wire _w456_ ;
	wire _w455_ ;
	wire _w454_ ;
	wire _w453_ ;
	wire _w466_ ;
	wire _w467_ ;
	wire _w468_ ;
	wire _w469_ ;
	wire _w470_ ;
	wire _w471_ ;
	wire _w472_ ;
	wire _w473_ ;
	wire _w474_ ;
	wire _w475_ ;
	wire _w476_ ;
	wire _w477_ ;
	wire _w478_ ;
	wire _w479_ ;
	wire _w480_ ;
	wire _w481_ ;
	wire _w512_ ;
	wire _w513_ ;
	wire _w514_ ;
	wire _w515_ ;
	wire _w516_ ;
	wire _w517_ ;
	wire _w518_ ;
	wire _w519_ ;
	wire _w520_ ;
	wire _w521_ ;
	wire _w522_ ;
	wire _w523_ ;
	wire _w524_ ;
	wire _w525_ ;
	wire _w526_ ;
	wire _w527_ ;
	wire _w528_ ;
	wire _w529_ ;
	wire _w530_ ;
	wire _w531_ ;
	wire _w532_ ;
	wire _w533_ ;
	wire _w534_ ;
	wire _w535_ ;
	wire _w536_ ;
	wire _w537_ ;
	wire _w538_ ;
	wire _w539_ ;
	wire _w540_ ;
	wire _w541_ ;
	wire _w542_ ;
	wire _w543_ ;
	wire _w544_ ;
	wire _w545_ ;
	wire _w546_ ;
	wire _w547_ ;
	wire _w548_ ;
	wire _w549_ ;
	wire _w550_ ;
	wire _w551_ ;
	wire _w552_ ;
	wire _w553_ ;
	wire _w554_ ;
	wire _w555_ ;
	wire _w556_ ;
	wire _w557_ ;
	wire _w558_ ;
	wire _w559_ ;
	wire _w560_ ;
	wire _w561_ ;
	wire _w562_ ;
	wire _w563_ ;
	wire _w564_ ;
	wire _w565_ ;
	wire _w566_ ;
	wire _w567_ ;
	wire _w568_ ;
	wire _w569_ ;
	wire _w570_ ;
	wire _w571_ ;
	wire _w572_ ;
	wire _w573_ ;
	wire _w574_ ;
	wire _w575_ ;
	wire _w576_ ;
	wire _w577_ ;
	wire _w578_ ;
	wire _w579_ ;
	wire _w710_ ;
	wire _w711_ ;
	wire _w712_ ;
	wire _w713_ ;
	wire _w714_ ;
	wire _w715_ ;
	wire _w716_ ;
	wire _w717_ ;
	wire _w718_ ;
	wire _w719_ ;
	wire _w720_ ;
	wire _w721_ ;
	wire _w722_ ;
	wire _w723_ ;
	wire _w724_ ;
	wire _w725_ ;
	wire _w726_ ;
	wire _w727_ ;
	wire _w728_ ;
	wire _w729_ ;
	wire _w730_ ;
	wire _w731_ ;
	wire _w732_ ;
	wire _w733_ ;
	wire _w734_ ;
	wire _w735_ ;
	wire _w736_ ;
	wire _w737_ ;
	wire _w738_ ;
	wire _w739_ ;
	wire _w740_ ;
	wire _w741_ ;
	wire _w742_ ;
	wire _w743_ ;
	wire _w744_ ;
	wire _w745_ ;
	wire _w746_ ;
	wire _w747_ ;
	wire _w748_ ;
	wire _w749_ ;
	wire _w750_ ;
	wire _w751_ ;
	wire _w752_ ;
	wire _w753_ ;
	wire _w754_ ;
	wire _w755_ ;
	wire _w756_ ;
	wire _w757_ ;
	wire _w758_ ;
	wire _w759_ ;
	wire _w760_ ;
	wire _w761_ ;
	wire _w762_ ;
	wire _w763_ ;
	wire _w764_ ;
	wire _w765_ ;
	wire _w766_ ;
	wire _w767_ ;
	wire _w768_ ;
	wire _w769_ ;
	wire _w770_ ;
	wire _w771_ ;
	wire _w772_ ;
	wire _w773_ ;
	wire _w774_ ;
	wire _w775_ ;
	wire _w776_ ;
	wire _w777_ ;
	wire _w778_ ;
	wire _w779_ ;
	wire _w780_ ;
	wire _w781_ ;
	wire _w782_ ;
	wire _w783_ ;
	wire _w784_ ;
	wire _w785_ ;
	wire _w786_ ;
	wire _w787_ ;
	wire _w788_ ;
	wire _w789_ ;
	wire _w790_ ;
	wire _w791_ ;
	wire _w792_ ;
	wire _w793_ ;
	wire _w794_ ;
	wire _w795_ ;
	wire _w796_ ;
	wire _w797_ ;
	wire _w798_ ;
	wire _w799_ ;
	wire _w800_ ;
	wire _w801_ ;
	wire _w802_ ;
	wire _w803_ ;
	wire _w804_ ;
	wire _w805_ ;
	wire _w806_ ;
	wire _w807_ ;
	wire _w808_ ;
	wire _w809_ ;
	wire _w810_ ;
	wire _w811_ ;
	wire _w812_ ;
	wire _w813_ ;
	wire _w814_ ;
	wire _w815_ ;
	wire _w816_ ;
	wire _w817_ ;
	wire _w818_ ;
	wire _w819_ ;
	wire _w820_ ;
	wire _w821_ ;
	wire _w822_ ;
	wire _w823_ ;
	wire _w824_ ;
	wire _w825_ ;
	wire _w826_ ;
	wire _w827_ ;
	wire _w828_ ;
	wire _w829_ ;
	wire _w830_ ;
	wire _w831_ ;
	wire _w832_ ;
	wire _w833_ ;
	wire _w834_ ;
	wire _w835_ ;
	wire _w836_ ;
	wire _w837_ ;
	wire _w838_ ;
	wire _w839_ ;
	wire _w840_ ;
	wire _w841_ ;
	wire _w842_ ;
	wire _w843_ ;
	wire _w844_ ;
	wire _w845_ ;
	wire _w846_ ;
	wire _w847_ ;
	wire _w848_ ;
	wire _w849_ ;
	wire _w850_ ;
	wire _w851_ ;
	wire _w852_ ;
	wire _w853_ ;
	wire _w854_ ;
	wire _w855_ ;
	wire _w856_ ;
	wire _w857_ ;
	wire _w858_ ;
	wire _w859_ ;
	wire _w860_ ;
	wire _w861_ ;
	wire _w862_ ;
	wire _w863_ ;
	wire _w864_ ;
	wire _w865_ ;
	wire _w866_ ;
	wire _w867_ ;
	wire _w868_ ;
	wire _w869_ ;
	wire _w870_ ;
	wire _w871_ ;
	wire _w872_ ;
	wire _w873_ ;
	wire _w874_ ;
	wire _w875_ ;
	wire _w876_ ;
	wire _w877_ ;
	wire _w878_ ;
	wire _w879_ ;
	wire _w880_ ;
	wire _w881_ ;
	wire _w882_ ;
	wire _w883_ ;
	wire _w884_ ;
	wire _w885_ ;
	wire _w886_ ;
	wire _w887_ ;
	wire _w888_ ;
	wire _w889_ ;
	wire _w890_ ;
	wire _w891_ ;
	wire _w892_ ;
	wire _w893_ ;
	wire _w894_ ;
	wire _w895_ ;
	wire _w896_ ;
	wire _w897_ ;
	wire _w898_ ;
	wire _w899_ ;
	wire _w900_ ;
	wire _w901_ ;
	wire _w902_ ;
	wire _w903_ ;
	wire _w904_ ;
	wire _w905_ ;
	wire _w906_ ;
	wire _w907_ ;
	wire _w908_ ;
	wire _w909_ ;
	wire _w910_ ;
	wire _w911_ ;
	wire _w912_ ;
	wire _w913_ ;
	wire _w914_ ;
	wire _w915_ ;
	wire _w916_ ;
	wire _w917_ ;
	wire _w918_ ;
	wire _w919_ ;
	wire _w920_ ;
	wire _w921_ ;
	wire _w922_ ;
	wire _w923_ ;
	wire _w924_ ;
	wire _w925_ ;
	wire _w926_ ;
	wire _w927_ ;
	wire _w928_ ;
	wire _w929_ ;
	wire _w930_ ;
	wire _w931_ ;
	wire _w932_ ;
	wire _w933_ ;
	wire _w934_ ;
	wire _w935_ ;
	wire _w936_ ;
	wire _w937_ ;
	wire _w938_ ;
	wire _w939_ ;
	wire _w940_ ;
	wire _w941_ ;
	wire _w942_ ;
	wire _w943_ ;
	wire _w944_ ;
	wire _w945_ ;
	wire _w946_ ;
	wire _w947_ ;
	wire _w948_ ;
	wire _w949_ ;
	wire _w950_ ;
	wire _w951_ ;
	wire _w952_ ;
	wire _w953_ ;
	wire _w954_ ;
	wire _w955_ ;
	wire _w956_ ;
	wire _w957_ ;
	wire _w958_ ;
	wire _w959_ ;
	wire _w960_ ;
	wire _w961_ ;
	wire _w962_ ;
	wire _w963_ ;
	wire _w964_ ;
	wire _w965_ ;
	wire _w966_ ;
	wire _w967_ ;
	wire _w968_ ;
	wire _w969_ ;
	wire _w970_ ;
	wire _w971_ ;
	wire _w972_ ;
	wire _w973_ ;
	wire _w974_ ;
	wire _w975_ ;
	wire _w976_ ;
	wire _w977_ ;
	wire _w978_ ;
	wire _w979_ ;
	wire _w980_ ;
	wire _w981_ ;
	wire _w982_ ;
	wire _w983_ ;
	wire _w984_ ;
	wire _w985_ ;
	wire _w986_ ;
	wire _w987_ ;
	wire _w988_ ;
	wire _w989_ ;
	wire _w990_ ;
	wire _w991_ ;
	wire _w992_ ;
	wire _w993_ ;
	wire _w1562_ ;
	wire _w1563_ ;
	wire _w1564_ ;
	wire _w1565_ ;
	wire _w1566_ ;
	wire _w1567_ ;
	wire _w1568_ ;
	wire _w1569_ ;
	wire _w1570_ ;
	wire _w1571_ ;
	wire _w1572_ ;
	wire _w1573_ ;
	wire _w1574_ ;
	wire _w1575_ ;
	wire _w1576_ ;
	wire _w1577_ ;
	wire _w1578_ ;
	wire _w1579_ ;
	wire _w1580_ ;
	wire _w1581_ ;
	wire _w1582_ ;
	wire _w1583_ ;
	wire _w1584_ ;
	wire _w1585_ ;
	wire _w1586_ ;
	wire _w1587_ ;
	wire _w1588_ ;
	wire _w1589_ ;
	wire _w1590_ ;
	wire _w1591_ ;
	wire _w1592_ ;
	wire _w1593_ ;
	wire _w1594_ ;
	wire _w1595_ ;
	wire _w1596_ ;
	wire _w1597_ ;
	wire _w1598_ ;
	wire _w1599_ ;
	wire _w1600_ ;
	wire _w1601_ ;
	wire _w1602_ ;
	wire _w1603_ ;
	wire _w1604_ ;
	wire _w1605_ ;
	wire _w1606_ ;
	wire _w1607_ ;
	wire _w1608_ ;
	wire _w1609_ ;
	wire _w1610_ ;
	wire _w1611_ ;
	wire _w1612_ ;
	wire _w1613_ ;
	wire _w1614_ ;
	wire _w1615_ ;
	wire _w1616_ ;
	wire _w1617_ ;
	wire _w1618_ ;
	wire _w1619_ ;
	wire _w1620_ ;
	wire _w1621_ ;
	wire _w1622_ ;
	wire _w1623_ ;
	wire _w1624_ ;
	wire _w1625_ ;
	wire _w1626_ ;
	wire _w1627_ ;
	wire _w1628_ ;
	wire _w1629_ ;
	wire _w1630_ ;
	wire _w1631_ ;
	wire _w1632_ ;
	wire _w1633_ ;
	wire _w1634_ ;
	wire _w1635_ ;
	wire _w1636_ ;
	wire _w1637_ ;
	wire _w1638_ ;
	wire _w1639_ ;
	wire _w1640_ ;
	wire _w1641_ ;
	wire _w1642_ ;
	wire _w1643_ ;
	wire _w1644_ ;
	wire _w1645_ ;
	wire _w1646_ ;
	wire _w1647_ ;
	wire _w1648_ ;
	wire _w1649_ ;
	wire _w1650_ ;
	wire _w1651_ ;
	wire _w1652_ ;
	wire _w1653_ ;
	wire _w1654_ ;
	wire _w1655_ ;
	wire _w1656_ ;
	wire _w1657_ ;
	wire _w1658_ ;
	wire _w1659_ ;
	wire _w1660_ ;
	wire _w1661_ ;
	wire _w1662_ ;
	wire _w1663_ ;
	wire _w1664_ ;
	wire _w1665_ ;
	wire _w1666_ ;
	wire _w1667_ ;
	wire _w1668_ ;
	wire _w1669_ ;
	wire _w1670_ ;
	wire _w1671_ ;
	wire _w1672_ ;
	wire _w1673_ ;
	wire _w1674_ ;
	wire _w1675_ ;
	wire _w1676_ ;
	wire _w1677_ ;
	wire _w1678_ ;
	wire _w1679_ ;
	wire _w1680_ ;
	wire _w1681_ ;
	wire _w1682_ ;
	wire _w1683_ ;
	wire _w1684_ ;
	wire _w1685_ ;
	wire _w1686_ ;
	wire _w1687_ ;
	wire _w1688_ ;
	wire _w1689_ ;
	wire _w1690_ ;
	wire _w1691_ ;
	wire _w1692_ ;
	wire _w1693_ ;
	wire _w1694_ ;
	wire _w1695_ ;
	wire _w1696_ ;
	wire _w1697_ ;
	wire _w1698_ ;
	wire _w1699_ ;
	wire _w1700_ ;
	wire _w1701_ ;
	wire _w1702_ ;
	wire _w1703_ ;
	wire _w1704_ ;
	wire _w1705_ ;
	wire _w1706_ ;
	wire _w1707_ ;
	wire _w1708_ ;
	wire _w1709_ ;
	wire _w1710_ ;
	wire _w1711_ ;
	wire _w1712_ ;
	wire _w1713_ ;
	wire _w1714_ ;
	wire _w1715_ ;
	wire _w1716_ ;
	wire _w1717_ ;
	wire _w1718_ ;
	wire _w1719_ ;
	wire _w1720_ ;
	wire _w1721_ ;
	wire _w1722_ ;
	wire _w1723_ ;
	wire _w1724_ ;
	wire _w1725_ ;
	wire _w1726_ ;
	wire _w1727_ ;
	wire _w1728_ ;
	wire _w1729_ ;
	wire _w1730_ ;
	wire _w1731_ ;
	wire _w1732_ ;
	wire _w1733_ ;
	wire _w1734_ ;
	wire _w1735_ ;
	wire _w1736_ ;
	wire _w1737_ ;
	wire _w1738_ ;
	wire _w1739_ ;
	wire _w1740_ ;
	wire _w1741_ ;
	wire _w1742_ ;
	wire _w1743_ ;
	wire _w1744_ ;
	wire _w1745_ ;
	wire _w1746_ ;
	wire _w1747_ ;
	wire _w1748_ ;
	wire _w1749_ ;
	wire _w1750_ ;
	wire _w1751_ ;
	wire _w1752_ ;
	wire _w1753_ ;
	wire _w1754_ ;
	wire _w1755_ ;
	wire _w1756_ ;
	wire _w1757_ ;
	wire _w1758_ ;
	wire _w1759_ ;
	wire _w1760_ ;
	wire _w1761_ ;
	wire _w1762_ ;
	wire _w1763_ ;
	wire _w1764_ ;
	wire _w1765_ ;
	wire _w1766_ ;
	wire _w1767_ ;
	wire _w1768_ ;
	wire _w1769_ ;
	wire _w1770_ ;
	wire _w1771_ ;
	wire _w1772_ ;
	wire _w1773_ ;
	wire _w1774_ ;
	wire _w1775_ ;
	wire _w1776_ ;
	wire _w1777_ ;
	wire _w1778_ ;
	wire _w1779_ ;
	wire _w1780_ ;
	wire _w1781_ ;
	wire _w1782_ ;
	wire _w1783_ ;
	wire _w1784_ ;
	wire _w1785_ ;
	wire _w1786_ ;
	wire _w1787_ ;
	wire _w1788_ ;
	wire _w1789_ ;
	wire _w1790_ ;
	wire _w1791_ ;
	wire _w1792_ ;
	wire _w1793_ ;
	wire _w1794_ ;
	wire _w1795_ ;
	wire _w1796_ ;
	wire _w1797_ ;
	wire _w1798_ ;
	wire _w1799_ ;
	wire _w1800_ ;
	wire _w1801_ ;
	wire _w1802_ ;
	wire _w1803_ ;
	wire _w1804_ ;
	wire _w1805_ ;
	wire _w1806_ ;
	wire _w1807_ ;
	wire _w1808_ ;
	wire _w1809_ ;
	wire _w1810_ ;
	wire _w1811_ ;
	wire _w1812_ ;
	wire _w1813_ ;
	wire _w1814_ ;
	wire _w1815_ ;
	wire _w1816_ ;
	wire _w1817_ ;
	wire _w1818_ ;
	wire _w1819_ ;
	wire _w1820_ ;
	wire _w1821_ ;
	wire _w1822_ ;
	wire _w1823_ ;
	wire _w1824_ ;
	wire _w1825_ ;
	wire _w1826_ ;
	wire _w1827_ ;
	wire _w1828_ ;
	wire _w1829_ ;
	wire _w1830_ ;
	wire _w1831_ ;
	wire _w1832_ ;
	wire _w1833_ ;
	wire _w1834_ ;
	wire _w1835_ ;
	wire _w1836_ ;
	wire _w1837_ ;
	wire _w1838_ ;
	wire _w1839_ ;
	wire _w1840_ ;
	wire _w1841_ ;
	wire _w1842_ ;
	wire _w1843_ ;
	wire _w1844_ ;
	wire _w1845_ ;
	wire _w1846_ ;
	wire _w1847_ ;
	wire _w1848_ ;
	wire _w1849_ ;
	wire _w1850_ ;
	wire _w1851_ ;
	wire _w1852_ ;
	wire _w1853_ ;
	wire _w1854_ ;
	wire _w1855_ ;
	wire _w1856_ ;
	wire _w1857_ ;
	wire _w1858_ ;
	wire _w1859_ ;
	wire _w1860_ ;
	wire _w1861_ ;
	wire _w1862_ ;
	wire _w1863_ ;
	wire _w1864_ ;
	wire _w1865_ ;
	wire _w1866_ ;
	wire _w1867_ ;
	wire _w1868_ ;
	wire _w1869_ ;
	wire _w1870_ ;
	wire _w1871_ ;
	wire _w1872_ ;
	wire _w1873_ ;
	wire _w1874_ ;
	wire _w1875_ ;
	wire _w1876_ ;
	wire _w1877_ ;
	wire _w1878_ ;
	wire _w1879_ ;
	wire _w1880_ ;
	wire _w1881_ ;
	wire _w1882_ ;
	wire _w1883_ ;
	wire _w1884_ ;
	wire _w1885_ ;
	wire _w1886_ ;
	wire _w1887_ ;
	wire _w1888_ ;
	wire _w1889_ ;
	wire _w1890_ ;
	wire _w1891_ ;
	wire _w1892_ ;
	wire _w1893_ ;
	wire _w1894_ ;
	wire _w1895_ ;
	wire _w1896_ ;
	wire _w1897_ ;
	wire _w1898_ ;
	wire _w1899_ ;
	wire _w1900_ ;
	wire _w1901_ ;
	wire _w1902_ ;
	wire _w1903_ ;
	wire _w1904_ ;
	wire _w1905_ ;
	wire _w1906_ ;
	wire _w1907_ ;
	wire _w1908_ ;
	wire _w1909_ ;
	wire _w1910_ ;
	wire _w1911_ ;
	wire _w1912_ ;
	wire _w1913_ ;
	wire _w1914_ ;
	wire _w1915_ ;
	wire _w1916_ ;
	wire _w1917_ ;
	wire _w1918_ ;
	wire _w1919_ ;
	wire _w1920_ ;
	wire _w1921_ ;
	wire _w1922_ ;
	wire _w1923_ ;
	wire _w1924_ ;
	wire _w1925_ ;
	wire _w1926_ ;
	wire _w1927_ ;
	wire _w1928_ ;
	wire _w1929_ ;
	wire _w1930_ ;
	wire _w1931_ ;
	wire _w1932_ ;
	wire _w1933_ ;
	wire _w1934_ ;
	wire _w1935_ ;
	wire _w1936_ ;
	wire _w1937_ ;
	wire _w1938_ ;
	wire _w1939_ ;
	wire _w1940_ ;
	wire _w1941_ ;
	wire _w1942_ ;
	wire _w1943_ ;
	wire _w1944_ ;
	wire _w1945_ ;
	wire _w1946_ ;
	wire _w1947_ ;
	wire _w1948_ ;
	wire _w1949_ ;
	wire _w1950_ ;
	wire _w1951_ ;
	wire _w1952_ ;
	wire _w1953_ ;
	wire _w1954_ ;
	wire _w1955_ ;
	wire _w1956_ ;
	wire _w1957_ ;
	wire _w1958_ ;
	wire _w1959_ ;
	wire _w1960_ ;
	wire _w1961_ ;
	wire _w1962_ ;
	wire _w1963_ ;
	wire _w1964_ ;
	wire _w1965_ ;
	wire _w1966_ ;
	wire _w1967_ ;
	wire _w1968_ ;
	wire _w1969_ ;
	wire _w1970_ ;
	wire _w1971_ ;
	wire _w1972_ ;
	wire _w1973_ ;
	wire _w1974_ ;
	wire _w1975_ ;
	wire _w1976_ ;
	wire _w1977_ ;
	wire _w1978_ ;
	wire _w1979_ ;
	wire _w1980_ ;
	wire _w1981_ ;
	wire _w1982_ ;
	wire _w1983_ ;
	wire _w1984_ ;
	wire _w1985_ ;
	wire _w1986_ ;
	wire _w1987_ ;
	wire _w1988_ ;
	wire _w1989_ ;
	wire _w1990_ ;
	wire _w1991_ ;
	wire _w1992_ ;
	wire _w1993_ ;
	wire _w1994_ ;
	wire _w1995_ ;
	wire _w1996_ ;
	wire _w1997_ ;
	wire _w1998_ ;
	wire _w1999_ ;
	wire _w2000_ ;
	wire _w2001_ ;
	wire _w2002_ ;
	wire _w2003_ ;
	wire _w2004_ ;
	wire _w2005_ ;
	wire _w2006_ ;
	wire _w2007_ ;
	wire _w2008_ ;
	wire _w2009_ ;
	wire _w2010_ ;
	wire _w2011_ ;
	wire _w2012_ ;
	wire _w2013_ ;
	wire _w2014_ ;
	wire _w2015_ ;
	wire _w2016_ ;
	wire _w2017_ ;
	wire _w2018_ ;
	wire _w2019_ ;
	wire _w2020_ ;
	wire _w2021_ ;
	wire _w2022_ ;
	wire _w2023_ ;
	wire _w2024_ ;
	wire _w2025_ ;
	wire _w2026_ ;
	wire _w2027_ ;
	wire _w2028_ ;
	wire _w2029_ ;
	wire _w2030_ ;
	wire _w2031_ ;
	wire _w2032_ ;
	wire _w2033_ ;
	wire _w2034_ ;
	wire _w2035_ ;
	wire _w2036_ ;
	wire _w2037_ ;
	wire _w2038_ ;
	wire _w2039_ ;
	wire _w2040_ ;
	wire _w2041_ ;
	wire _w2042_ ;
	wire _w2043_ ;
	wire _w2044_ ;
	wire _w2045_ ;
	wire _w2046_ ;
	wire _w2047_ ;
	wire _w2048_ ;
	wire _w2049_ ;
	wire _w2050_ ;
	wire _w2051_ ;
	wire _w2052_ ;
	wire _w2053_ ;
	wire _w2054_ ;
	wire _w2055_ ;
	wire _w2056_ ;
	wire _w2057_ ;
	wire _w2058_ ;
	wire _w2059_ ;
	wire _w2060_ ;
	wire _w2061_ ;
	wire _w2062_ ;
	wire _w2063_ ;
	wire _w2064_ ;
	wire _w2065_ ;
	wire _w2066_ ;
	wire _w2067_ ;
	wire _w2068_ ;
	wire _w2069_ ;
	wire _w2070_ ;
	wire _w2071_ ;
	wire _w2072_ ;
	wire _w2073_ ;
	wire _w2074_ ;
	wire _w2075_ ;
	wire _w2076_ ;
	wire _w2077_ ;
	wire _w2078_ ;
	wire _w2079_ ;
	wire _w2080_ ;
	wire _w2081_ ;
	wire _w2082_ ;
	wire _w2083_ ;
	wire _w2084_ ;
	wire _w2085_ ;
	wire _w2086_ ;
	wire _w2087_ ;
	wire _w2088_ ;
	wire _w2089_ ;
	wire _w2090_ ;
	wire _w2091_ ;
	wire _w2092_ ;
	wire _w2093_ ;
	wire _w2094_ ;
	wire _w2095_ ;
	wire _w2096_ ;
	wire _w2097_ ;
	wire _w2098_ ;
	wire _w2099_ ;
	wire _w2100_ ;
	wire _w2101_ ;
	wire _w2102_ ;
	wire _w2103_ ;
	wire _w2104_ ;
	wire _w2105_ ;
	wire _w2106_ ;
	wire _w2107_ ;
	wire _w2108_ ;
	wire _w2109_ ;
	wire _w2110_ ;
	wire _w2111_ ;
	wire _w2112_ ;
	wire _w2113_ ;
	wire _w2114_ ;
	wire _w2115_ ;
	wire _w2116_ ;
	wire _w2117_ ;
	wire _w2118_ ;
	wire _w2119_ ;
	wire _w2120_ ;
	wire _w2121_ ;
	wire _w2122_ ;
	wire _w2123_ ;
	wire _w2124_ ;
	wire _w2125_ ;
	wire _w2126_ ;
	wire _w2127_ ;
	wire _w2128_ ;
	wire _w2129_ ;
	wire _w2130_ ;
	wire _w2131_ ;
	wire _w2132_ ;
	wire _w2133_ ;
	wire _w2134_ ;
	wire _w2135_ ;
	wire _w2136_ ;
	wire _w2137_ ;
	wire _w2138_ ;
	wire _w2139_ ;
	wire _w2140_ ;
	wire _w2141_ ;
	wire _w2142_ ;
	wire _w2143_ ;
	wire _w2144_ ;
	wire _w2145_ ;
	wire _w2146_ ;
	wire _w2147_ ;
	wire _w2148_ ;
	wire _w2149_ ;
	wire _w2150_ ;
	wire _w2151_ ;
	wire _w2152_ ;
	wire _w2153_ ;
	wire _w2154_ ;
	wire _w2155_ ;
	wire _w2156_ ;
	wire _w2157_ ;
	wire _w2158_ ;
	wire _w2159_ ;
	wire _w2160_ ;
	wire _w2161_ ;
	wire _w2162_ ;
	wire _w2163_ ;
	wire _w2164_ ;
	wire _w2165_ ;
	wire _w2166_ ;
	wire _w2167_ ;
	wire _w2168_ ;
	wire _w2169_ ;
	wire _w2170_ ;
	wire _w2171_ ;
	wire _w2172_ ;
	wire _w2173_ ;
	wire _w2174_ ;
	wire _w2175_ ;
	wire _w2176_ ;
	wire _w2177_ ;
	wire _w2178_ ;
	wire _w2179_ ;
	wire _w2180_ ;
	wire _w2181_ ;
	wire _w2182_ ;
	wire _w2183_ ;
	wire _w2184_ ;
	wire _w2185_ ;
	wire _w2186_ ;
	wire _w2187_ ;
	wire _w2188_ ;
	wire _w2189_ ;
	wire _w2190_ ;
	wire _w2191_ ;
	wire _w2192_ ;
	wire _w2193_ ;
	wire _w2194_ ;
	wire _w2195_ ;
	wire _w2196_ ;
	wire _w2197_ ;
	wire _w2198_ ;
	wire _w2199_ ;
	wire _w2200_ ;
	wire _w2201_ ;
	wire _w2202_ ;
	wire _w2203_ ;
	wire _w2204_ ;
	wire _w2205_ ;
	wire _w2206_ ;
	wire _w2207_ ;
	wire _w2208_ ;
	wire _w2209_ ;
	wire _w2210_ ;
	wire _w2211_ ;
	wire _w2212_ ;
	wire _w2213_ ;
	wire _w2214_ ;
	wire _w2215_ ;
	wire _w2216_ ;
	wire _w2217_ ;
	wire _w2218_ ;
	wire _w2219_ ;
	wire _w2220_ ;
	wire _w2221_ ;
	wire _w2222_ ;
	wire _w2223_ ;
	wire _w2224_ ;
	wire _w2225_ ;
	wire _w2226_ ;
	wire _w2227_ ;
	wire _w2228_ ;
	wire _w2229_ ;
	wire _w2230_ ;
	wire _w2231_ ;
	wire _w2232_ ;
	wire _w2233_ ;
	wire _w2234_ ;
	wire _w2235_ ;
	wire _w2236_ ;
	wire _w2237_ ;
	wire _w2238_ ;
	wire _w2239_ ;
	wire _w2240_ ;
	wire _w2241_ ;
	wire _w2242_ ;
	wire _w2243_ ;
	wire _w2244_ ;
	wire _w2245_ ;
	wire _w2246_ ;
	wire _w2247_ ;
	wire _w2248_ ;
	wire _w2249_ ;
	wire _w2250_ ;
	wire _w2251_ ;
	wire _w2252_ ;
	wire _w2253_ ;
	wire _w2254_ ;
	wire _w2255_ ;
	wire _w2256_ ;
	wire _w2257_ ;
	wire _w2258_ ;
	wire _w2259_ ;
	wire _w2260_ ;
	wire _w2261_ ;
	wire _w2262_ ;
	wire _w2263_ ;
	wire _w2264_ ;
	wire _w2265_ ;
	wire _w2266_ ;
	wire _w2267_ ;
	wire _w2268_ ;
	wire _w2269_ ;
	wire _w2270_ ;
	wire _w2271_ ;
	wire _w2272_ ;
	wire _w2273_ ;
	wire _w2274_ ;
	wire _w2275_ ;
	wire _w2276_ ;
	wire _w2277_ ;
	wire _w2278_ ;
	wire _w2279_ ;
	wire _w2280_ ;
	wire _w2281_ ;
	wire _w2282_ ;
	wire _w2283_ ;
	wire _w2284_ ;
	wire _w2285_ ;
	wire _w2286_ ;
	wire _w2287_ ;
	wire _w2288_ ;
	wire _w2289_ ;
	wire _w2290_ ;
	wire _w2291_ ;
	wire _w2292_ ;
	wire _w2293_ ;
	wire _w2294_ ;
	wire _w2295_ ;
	wire _w2296_ ;
	wire _w2297_ ;
	wire _w2298_ ;
	wire _w2299_ ;
	wire _w2300_ ;
	wire _w2301_ ;
	wire _w2302_ ;
	wire _w2303_ ;
	wire _w2304_ ;
	wire _w2305_ ;
	wire _w2306_ ;
	wire _w2307_ ;
	wire _w2308_ ;
	wire _w2309_ ;
	wire _w2310_ ;
	wire _w2311_ ;
	wire _w2312_ ;
	wire _w2313_ ;
	wire _w2314_ ;
	wire _w2315_ ;
	wire _w2316_ ;
	wire _w2317_ ;
	wire _w2318_ ;
	wire _w2319_ ;
	wire _w2320_ ;
	wire _w2321_ ;
	wire _w2322_ ;
	wire _w2323_ ;
	wire _w2324_ ;
	wire _w2325_ ;
	wire _w2326_ ;
	wire _w2327_ ;
	wire _w2328_ ;
	wire _w2329_ ;
	wire _w2330_ ;
	wire _w2331_ ;
	wire _w2332_ ;
	wire _w2333_ ;
	wire _w2334_ ;
	wire _w2335_ ;
	wire _w2336_ ;
	wire _w2337_ ;
	wire _w2338_ ;
	wire _w2339_ ;
	wire _w2340_ ;
	wire _w2341_ ;
	wire _w2342_ ;
	wire _w2343_ ;
	wire _w2344_ ;
	wire _w2345_ ;
	wire _w2346_ ;
	wire _w2347_ ;
	wire _w2348_ ;
	wire _w2349_ ;
	wire _w2350_ ;
	wire _w2351_ ;
	wire _w2352_ ;
	wire _w2353_ ;
	wire _w2354_ ;
	wire _w2355_ ;
	wire _w2356_ ;
	wire _w2357_ ;
	wire _w2358_ ;
	wire _w2359_ ;
	wire _w2360_ ;
	wire _w2361_ ;
	wire _w2362_ ;
	wire _w2363_ ;
	wire _w2364_ ;
	wire _w2365_ ;
	wire _w2366_ ;
	wire _w2367_ ;
	wire _w2368_ ;
	wire _w2369_ ;
	wire _w2370_ ;
	wire _w2371_ ;
	wire _w2372_ ;
	wire _w2373_ ;
	wire _w2374_ ;
	wire _w2375_ ;
	wire _w2376_ ;
	wire _w2377_ ;
	wire _w2378_ ;
	wire _w2379_ ;
	wire _w2380_ ;
	wire _w2381_ ;
	wire _w2382_ ;
	wire _w2383_ ;
	wire _w2384_ ;
	wire _w2385_ ;
	wire _w2386_ ;
	wire _w2387_ ;
	wire _w2388_ ;
	wire _w2389_ ;
	wire _w2390_ ;
	wire _w2391_ ;
	wire _w2392_ ;
	wire _w2393_ ;
	wire _w2394_ ;
	wire _w2395_ ;
	wire _w2396_ ;
	wire _w2397_ ;
	wire _w2398_ ;
	wire _w2399_ ;
	wire _w2400_ ;
	wire _w2401_ ;
	wire _w2402_ ;
	wire _w2403_ ;
	wire _w2404_ ;
	wire _w2405_ ;
	wire _w2406_ ;
	wire _w2407_ ;
	wire _w2408_ ;
	wire _w2409_ ;
	wire _w2410_ ;
	wire _w2411_ ;
	wire _w2412_ ;
	wire _w2413_ ;
	wire _w2414_ ;
	wire _w2415_ ;
	wire _w2416_ ;
	wire _w2417_ ;
	wire _w2418_ ;
	wire _w2419_ ;
	wire _w2420_ ;
	wire _w2421_ ;
	wire _w2422_ ;
	wire _w2423_ ;
	wire _w2424_ ;
	wire _w2425_ ;
	wire _w2426_ ;
	wire _w2427_ ;
	wire _w2428_ ;
	wire _w2429_ ;
	wire _w2430_ ;
	wire _w2431_ ;
	wire _w2432_ ;
	wire _w2433_ ;
	wire _w2434_ ;
	wire _w2435_ ;
	wire _w2436_ ;
	wire _w2437_ ;
	wire _w2438_ ;
	wire _w2439_ ;
	wire _w2440_ ;
	wire _w2441_ ;
	wire _w2442_ ;
	wire _w2443_ ;
	wire _w2444_ ;
	wire _w2445_ ;
	wire _w2446_ ;
	wire _w2447_ ;
	wire _w2448_ ;
	wire _w2449_ ;
	wire _w2450_ ;
	wire _w2451_ ;
	wire _w2452_ ;
	wire _w2453_ ;
	wire _w2454_ ;
	wire _w2455_ ;
	wire _w2456_ ;
	wire _w2457_ ;
	wire _w2458_ ;
	wire _w2459_ ;
	wire _w2460_ ;
	wire _w2461_ ;
	wire _w2462_ ;
	wire _w2463_ ;
	wire _w2464_ ;
	wire _w2465_ ;
	wire _w2466_ ;
	wire _w2467_ ;
	wire _w2468_ ;
	wire _w2469_ ;
	wire _w2470_ ;
	wire _w2471_ ;
	wire _w2472_ ;
	wire _w2473_ ;
	wire _w2474_ ;
	wire _w2475_ ;
	wire _w2476_ ;
	wire _w2477_ ;
	wire _w2478_ ;
	wire _w2479_ ;
	wire _w2480_ ;
	wire _w2481_ ;
	wire _w2482_ ;
	wire _w2483_ ;
	wire _w2484_ ;
	wire _w2485_ ;
	wire _w2486_ ;
	wire _w2487_ ;
	wire _w2488_ ;
	wire _w2489_ ;
	wire _w2490_ ;
	wire _w2491_ ;
	wire _w2492_ ;
	wire _w2493_ ;
	wire _w2494_ ;
	wire _w2495_ ;
	wire _w2496_ ;
	wire _w2497_ ;
	wire _w2498_ ;
	wire _w2499_ ;
	wire _w2500_ ;
	wire _w2501_ ;
	wire _w2502_ ;
	wire _w2503_ ;
	wire _w2504_ ;
	wire _w2505_ ;
	wire _w2506_ ;
	wire _w2507_ ;
	wire _w2508_ ;
	wire _w2509_ ;
	wire _w2510_ ;
	wire _w2511_ ;
	wire _w2512_ ;
	wire _w2513_ ;
	wire _w2514_ ;
	wire _w2515_ ;
	wire _w2516_ ;
	wire _w2517_ ;
	wire _w2518_ ;
	wire _w2519_ ;
	wire _w2520_ ;
	wire _w2521_ ;
	wire _w2522_ ;
	wire _w2523_ ;
	wire _w2524_ ;
	wire _w2525_ ;
	wire _w2526_ ;
	wire _w2527_ ;
	wire _w2528_ ;
	wire _w2529_ ;
	wire _w2530_ ;
	wire _w2531_ ;
	wire _w2532_ ;
	wire _w2533_ ;
	wire _w2534_ ;
	wire _w2535_ ;
	wire _w2536_ ;
	wire _w2537_ ;
	wire _w2538_ ;
	wire _w2539_ ;
	wire _w2540_ ;
	wire _w2541_ ;
	wire _w2542_ ;
	wire _w2543_ ;
	wire _w2544_ ;
	wire _w2545_ ;
	wire _w2546_ ;
	wire _w2547_ ;
	wire _w2548_ ;
	wire _w2549_ ;
	wire _w2550_ ;
	wire _w2551_ ;
	wire _w2552_ ;
	wire _w2553_ ;
	wire _w2554_ ;
	wire _w2555_ ;
	wire _w2556_ ;
	wire _w2557_ ;
	wire _w2558_ ;
	wire _w2559_ ;
	wire _w2560_ ;
	wire _w2561_ ;
	wire _w2562_ ;
	wire _w2563_ ;
	wire _w2564_ ;
	wire _w2565_ ;
	wire _w2566_ ;
	wire _w2567_ ;
	wire _w2568_ ;
	wire _w2569_ ;
	wire _w2570_ ;
	wire _w2571_ ;
	wire _w2572_ ;
	wire _w2573_ ;
	wire _w2574_ ;
	wire _w2575_ ;
	wire _w2576_ ;
	wire _w2577_ ;
	wire _w2578_ ;
	wire _w2579_ ;
	wire _w2580_ ;
	wire _w2581_ ;
	wire _w2582_ ;
	wire _w2583_ ;
	wire _w2584_ ;
	wire _w2585_ ;
	wire _w2586_ ;
	wire _w2587_ ;
	wire _w2588_ ;
	wire _w2589_ ;
	wire _w2590_ ;
	wire _w2591_ ;
	wire _w2592_ ;
	wire _w2593_ ;
	wire _w2594_ ;
	wire _w2595_ ;
	wire _w2596_ ;
	wire _w2597_ ;
	wire _w2598_ ;
	wire _w2599_ ;
	wire _w2600_ ;
	wire _w2601_ ;
	wire _w2602_ ;
	wire _w2603_ ;
	wire _w2604_ ;
	wire _w2605_ ;
	wire _w2606_ ;
	wire _w2607_ ;
	wire _w2608_ ;
	wire _w2609_ ;
	wire _w2610_ ;
	wire _w2611_ ;
	wire _w2612_ ;
	wire _w2613_ ;
	wire _w2614_ ;
	wire _w2615_ ;
	wire _w2616_ ;
	wire _w2617_ ;
	wire _w2618_ ;
	wire _w2619_ ;
	wire _w2620_ ;
	wire _w2621_ ;
	wire _w2622_ ;
	wire _w2623_ ;
	wire _w2624_ ;
	wire _w2625_ ;
	wire _w2626_ ;
	wire _w2627_ ;
	wire _w2628_ ;
	wire _w2629_ ;
	wire _w2630_ ;
	wire _w2631_ ;
	wire _w2632_ ;
	wire _w2633_ ;
	wire _w2634_ ;
	wire _w2635_ ;
	wire _w2636_ ;
	wire _w2637_ ;
	wire _w2638_ ;
	wire _w2639_ ;
	wire _w2640_ ;
	wire _w2641_ ;
	wire _w2642_ ;
	wire _w2643_ ;
	wire _w2644_ ;
	wire _w2645_ ;
	wire _w2646_ ;
	wire _w2647_ ;
	wire _w2648_ ;
	wire _w2649_ ;
	wire _w2650_ ;
	wire _w2651_ ;
	wire _w2652_ ;
	wire _w2653_ ;
	wire _w2654_ ;
	wire _w2655_ ;
	wire _w2656_ ;
	wire _w2657_ ;
	wire _w2658_ ;
	wire _w2659_ ;
	wire _w2660_ ;
	wire _w2661_ ;
	wire _w2662_ ;
	wire _w2663_ ;
	wire _w2664_ ;
	wire _w2665_ ;
	wire _w2666_ ;
	wire _w2667_ ;
	wire _w2668_ ;
	wire _w2669_ ;
	wire _w2670_ ;
	wire _w2671_ ;
	wire _w2672_ ;
	wire _w2673_ ;
	wire _w2674_ ;
	wire _w2675_ ;
	wire _w2676_ ;
	wire _w2677_ ;
	wire _w2678_ ;
	wire _w2679_ ;
	wire _w2680_ ;
	wire _w2681_ ;
	wire _w2682_ ;
	wire _w2683_ ;
	wire _w2684_ ;
	wire _w2685_ ;
	wire _w2686_ ;
	wire _w2687_ ;
	wire _w2688_ ;
	wire _w2689_ ;
	wire _w2690_ ;
	wire _w2691_ ;
	wire _w2692_ ;
	wire _w2693_ ;
	wire _w2694_ ;
	wire _w2695_ ;
	wire _w2696_ ;
	wire _w2697_ ;
	wire _w2698_ ;
	wire _w2699_ ;
	wire _w2700_ ;
	wire _w2701_ ;
	wire _w2702_ ;
	wire _w2703_ ;
	wire _w2704_ ;
	wire _w2705_ ;
	wire _w2706_ ;
	wire _w2707_ ;
	wire _w2708_ ;
	wire _w2709_ ;
	wire _w2710_ ;
	wire _w2711_ ;
	wire _w2712_ ;
	wire _w2713_ ;
	wire _w2714_ ;
	wire _w2715_ ;
	wire _w2716_ ;
	wire _w2717_ ;
	wire _w2718_ ;
	wire _w2719_ ;
	wire _w2720_ ;
	wire _w2721_ ;
	wire _w2722_ ;
	wire _w2723_ ;
	wire _w2724_ ;
	wire _w2725_ ;
	wire _w2726_ ;
	wire _w2727_ ;
	wire _w2728_ ;
	wire _w2729_ ;
	wire _w2730_ ;
	wire _w2731_ ;
	wire _w2732_ ;
	wire _w2733_ ;
	wire _w2734_ ;
	wire _w2735_ ;
	wire _w2736_ ;
	wire _w2737_ ;
	wire _w2738_ ;
	wire _w2739_ ;
	wire _w2740_ ;
	wire _w2741_ ;
	wire _w2742_ ;
	wire _w2743_ ;
	wire _w2744_ ;
	wire _w2745_ ;
	wire _w2746_ ;
	wire _w2747_ ;
	wire _w2748_ ;
	wire _w2749_ ;
	wire _w2750_ ;
	wire _w2751_ ;
	wire _w2752_ ;
	wire _w2753_ ;
	wire _w2754_ ;
	wire _w2755_ ;
	wire _w2756_ ;
	wire _w2757_ ;
	wire _w2758_ ;
	wire _w2759_ ;
	wire _w2760_ ;
	wire _w2761_ ;
	wire _w2762_ ;
	wire _w2763_ ;
	wire _w2764_ ;
	wire _w2765_ ;
	wire _w2766_ ;
	wire _w2767_ ;
	wire _w2768_ ;
	wire _w2769_ ;
	wire _w2770_ ;
	wire _w2771_ ;
	wire _w2772_ ;
	wire _w2773_ ;
	wire _w2774_ ;
	wire _w2775_ ;
	wire _w2776_ ;
	wire _w2777_ ;
	wire _w2778_ ;
	wire _w2779_ ;
	wire _w2780_ ;
	wire _w2781_ ;
	wire _w2782_ ;
	wire _w2783_ ;
	wire _w2784_ ;
	wire _w2785_ ;
	wire _w2786_ ;
	wire _w2787_ ;
	wire _w2788_ ;
	wire _w2789_ ;
	wire _w2790_ ;
	wire _w2791_ ;
	wire _w2792_ ;
	wire _w2793_ ;
	wire _w2794_ ;
	wire _w2795_ ;
	wire _w2796_ ;
	wire _w2797_ ;
	wire _w2798_ ;
	wire _w2799_ ;
	wire _w2800_ ;
	wire _w2801_ ;
	wire _w2802_ ;
	wire _w2803_ ;
	wire _w2804_ ;
	wire _w2805_ ;
	wire _w2806_ ;
	wire _w2807_ ;
	wire _w2808_ ;
	wire _w2809_ ;
	LUT4 #(
		.INIT('h0002)
	) name0 (
		\InstQueueRd_Addr_reg[0]/NET0131 ,
		\InstQueueRd_Addr_reg[1]/NET0131 ,
		\InstQueueRd_Addr_reg[2]/NET0131 ,
		\InstQueueRd_Addr_reg[3]/NET0131 ,
		_w453_
	);
	LUT4 #(
		.INIT('h0200)
	) name1 (
		\InstQueueRd_Addr_reg[0]/NET0131 ,
		\InstQueueRd_Addr_reg[1]/NET0131 ,
		\InstQueueRd_Addr_reg[2]/NET0131 ,
		\InstQueueRd_Addr_reg[3]/NET0131 ,
		_w454_
	);
	LUT4 #(
		.INIT('h135f)
	) name2 (
		\InstQueue_reg[1][7]/NET0131 ,
		\InstQueue_reg[9][7]/NET0131 ,
		_w453_,
		_w454_,
		_w455_
	);
	LUT4 #(
		.INIT('h2000)
	) name3 (
		\InstQueueRd_Addr_reg[0]/NET0131 ,
		\InstQueueRd_Addr_reg[1]/NET0131 ,
		\InstQueueRd_Addr_reg[2]/NET0131 ,
		\InstQueueRd_Addr_reg[3]/NET0131 ,
		_w456_
	);
	LUT2 #(
		.INIT('h8)
	) name4 (
		\InstQueueRd_Addr_reg[0]/NET0131 ,
		\InstQueueRd_Addr_reg[1]/NET0131 ,
		_w457_
	);
	LUT4 #(
		.INIT('h0800)
	) name5 (
		\InstQueueRd_Addr_reg[0]/NET0131 ,
		\InstQueueRd_Addr_reg[1]/NET0131 ,
		\InstQueueRd_Addr_reg[2]/NET0131 ,
		\InstQueueRd_Addr_reg[3]/NET0131 ,
		_w458_
	);
	LUT4 #(
		.INIT('h153f)
	) name6 (
		\InstQueue_reg[11][7]/NET0131 ,
		\InstQueue_reg[13][7]/NET0131 ,
		_w456_,
		_w458_,
		_w459_
	);
	LUT4 #(
		.INIT('h4000)
	) name7 (
		\InstQueueRd_Addr_reg[0]/NET0131 ,
		\InstQueueRd_Addr_reg[1]/NET0131 ,
		\InstQueueRd_Addr_reg[2]/NET0131 ,
		\InstQueueRd_Addr_reg[3]/NET0131 ,
		_w460_
	);
	LUT4 #(
		.INIT('h0040)
	) name8 (
		\InstQueueRd_Addr_reg[0]/NET0131 ,
		\InstQueueRd_Addr_reg[1]/NET0131 ,
		\InstQueueRd_Addr_reg[2]/NET0131 ,
		\InstQueueRd_Addr_reg[3]/NET0131 ,
		_w461_
	);
	LUT4 #(
		.INIT('h135f)
	) name9 (
		\InstQueue_reg[14][7]/NET0131 ,
		\InstQueue_reg[6][7]/NET0131 ,
		_w460_,
		_w461_,
		_w462_
	);
	LUT4 #(
		.INIT('h0001)
	) name10 (
		\InstQueueRd_Addr_reg[0]/NET0131 ,
		\InstQueueRd_Addr_reg[1]/NET0131 ,
		\InstQueueRd_Addr_reg[2]/NET0131 ,
		\InstQueueRd_Addr_reg[3]/NET0131 ,
		_w463_
	);
	LUT4 #(
		.INIT('h0010)
	) name11 (
		\InstQueueRd_Addr_reg[0]/NET0131 ,
		\InstQueueRd_Addr_reg[1]/NET0131 ,
		\InstQueueRd_Addr_reg[2]/NET0131 ,
		\InstQueueRd_Addr_reg[3]/NET0131 ,
		_w464_
	);
	LUT4 #(
		.INIT('h135f)
	) name12 (
		\InstQueue_reg[0][7]/NET0131 ,
		\InstQueue_reg[4][7]/NET0131 ,
		_w463_,
		_w464_,
		_w465_
	);
	LUT4 #(
		.INIT('h8000)
	) name13 (
		_w462_,
		_w465_,
		_w455_,
		_w459_,
		_w466_
	);
	LUT4 #(
		.INIT('h0020)
	) name14 (
		\InstQueueRd_Addr_reg[0]/NET0131 ,
		\InstQueueRd_Addr_reg[1]/NET0131 ,
		\InstQueueRd_Addr_reg[2]/NET0131 ,
		\InstQueueRd_Addr_reg[3]/NET0131 ,
		_w467_
	);
	LUT4 #(
		.INIT('h0100)
	) name15 (
		\InstQueueRd_Addr_reg[0]/NET0131 ,
		\InstQueueRd_Addr_reg[1]/NET0131 ,
		\InstQueueRd_Addr_reg[2]/NET0131 ,
		\InstQueueRd_Addr_reg[3]/NET0131 ,
		_w468_
	);
	LUT4 #(
		.INIT('h135f)
	) name16 (
		\InstQueue_reg[5][7]/NET0131 ,
		\InstQueue_reg[8][7]/NET0131 ,
		_w467_,
		_w468_,
		_w469_
	);
	LUT4 #(
		.INIT('h1000)
	) name17 (
		\InstQueueRd_Addr_reg[0]/NET0131 ,
		\InstQueueRd_Addr_reg[1]/NET0131 ,
		\InstQueueRd_Addr_reg[2]/NET0131 ,
		\InstQueueRd_Addr_reg[3]/NET0131 ,
		_w470_
	);
	LUT4 #(
		.INIT('h0400)
	) name18 (
		\InstQueueRd_Addr_reg[0]/NET0131 ,
		\InstQueueRd_Addr_reg[1]/NET0131 ,
		\InstQueueRd_Addr_reg[2]/NET0131 ,
		\InstQueueRd_Addr_reg[3]/NET0131 ,
		_w471_
	);
	LUT4 #(
		.INIT('h153f)
	) name19 (
		\InstQueue_reg[10][7]/NET0131 ,
		\InstQueue_reg[12][7]/NET0131 ,
		_w470_,
		_w471_,
		_w472_
	);
	LUT4 #(
		.INIT('h8000)
	) name20 (
		\InstQueueRd_Addr_reg[0]/NET0131 ,
		\InstQueueRd_Addr_reg[1]/NET0131 ,
		\InstQueueRd_Addr_reg[2]/NET0131 ,
		\InstQueueRd_Addr_reg[3]/NET0131 ,
		_w473_
	);
	LUT4 #(
		.INIT('h0004)
	) name21 (
		\InstQueueRd_Addr_reg[0]/NET0131 ,
		\InstQueueRd_Addr_reg[1]/NET0131 ,
		\InstQueueRd_Addr_reg[2]/NET0131 ,
		\InstQueueRd_Addr_reg[3]/NET0131 ,
		_w474_
	);
	LUT4 #(
		.INIT('h135f)
	) name22 (
		\InstQueue_reg[15][7]/NET0131 ,
		\InstQueue_reg[2][7]/NET0131 ,
		_w473_,
		_w474_,
		_w475_
	);
	LUT4 #(
		.INIT('h0008)
	) name23 (
		\InstQueueRd_Addr_reg[0]/NET0131 ,
		\InstQueueRd_Addr_reg[1]/NET0131 ,
		\InstQueueRd_Addr_reg[2]/NET0131 ,
		\InstQueueRd_Addr_reg[3]/NET0131 ,
		_w476_
	);
	LUT4 #(
		.INIT('h0080)
	) name24 (
		\InstQueueRd_Addr_reg[0]/NET0131 ,
		\InstQueueRd_Addr_reg[1]/NET0131 ,
		\InstQueueRd_Addr_reg[2]/NET0131 ,
		\InstQueueRd_Addr_reg[3]/NET0131 ,
		_w477_
	);
	LUT4 #(
		.INIT('h135f)
	) name25 (
		\InstQueue_reg[3][7]/NET0131 ,
		\InstQueue_reg[7][7]/NET0131 ,
		_w476_,
		_w477_,
		_w478_
	);
	LUT4 #(
		.INIT('h8000)
	) name26 (
		_w475_,
		_w478_,
		_w469_,
		_w472_,
		_w479_
	);
	LUT2 #(
		.INIT('h8)
	) name27 (
		_w466_,
		_w479_,
		_w480_
	);
	LUT4 #(
		.INIT('h135f)
	) name28 (
		\InstQueue_reg[0][6]/NET0131 ,
		\InstQueue_reg[1][6]/NET0131 ,
		_w463_,
		_w453_,
		_w481_
	);
	LUT4 #(
		.INIT('h135f)
	) name29 (
		\InstQueue_reg[5][6]/NET0131 ,
		\InstQueue_reg[8][6]/NET0131 ,
		_w467_,
		_w468_,
		_w482_
	);
	LUT4 #(
		.INIT('h153f)
	) name30 (
		\InstQueue_reg[11][6]/NET0131 ,
		\InstQueue_reg[14][6]/NET0131 ,
		_w460_,
		_w458_,
		_w483_
	);
	LUT4 #(
		.INIT('h153f)
	) name31 (
		\InstQueue_reg[3][6]/NET0131 ,
		\InstQueue_reg[6][6]/NET0131 ,
		_w461_,
		_w476_,
		_w484_
	);
	LUT4 #(
		.INIT('h8000)
	) name32 (
		_w483_,
		_w484_,
		_w481_,
		_w482_,
		_w485_
	);
	LUT4 #(
		.INIT('h153f)
	) name33 (
		\InstQueue_reg[2][6]/NET0131 ,
		\InstQueue_reg[9][6]/NET0131 ,
		_w454_,
		_w474_,
		_w486_
	);
	LUT4 #(
		.INIT('h153f)
	) name34 (
		\InstQueue_reg[13][6]/NET0131 ,
		\InstQueue_reg[4][6]/NET0131 ,
		_w464_,
		_w456_,
		_w487_
	);
	LUT4 #(
		.INIT('h153f)
	) name35 (
		\InstQueue_reg[12][6]/NET0131 ,
		\InstQueue_reg[7][6]/NET0131 ,
		_w477_,
		_w470_,
		_w488_
	);
	LUT4 #(
		.INIT('h153f)
	) name36 (
		\InstQueue_reg[10][6]/NET0131 ,
		\InstQueue_reg[15][6]/NET0131 ,
		_w473_,
		_w471_,
		_w489_
	);
	LUT4 #(
		.INIT('h8000)
	) name37 (
		_w488_,
		_w489_,
		_w486_,
		_w487_,
		_w490_
	);
	LUT2 #(
		.INIT('h8)
	) name38 (
		_w485_,
		_w490_,
		_w491_
	);
	LUT4 #(
		.INIT('h0777)
	) name39 (
		_w466_,
		_w479_,
		_w485_,
		_w490_,
		_w492_
	);
	LUT4 #(
		.INIT('h153f)
	) name40 (
		\InstQueue_reg[11][2]/NET0131 ,
		\InstQueue_reg[14][2]/NET0131 ,
		_w460_,
		_w458_,
		_w493_
	);
	LUT4 #(
		.INIT('h135f)
	) name41 (
		\InstQueue_reg[7][2]/NET0131 ,
		\InstQueue_reg[8][2]/NET0131 ,
		_w477_,
		_w468_,
		_w494_
	);
	LUT4 #(
		.INIT('h135f)
	) name42 (
		\InstQueue_reg[13][2]/NET0131 ,
		\InstQueue_reg[2][2]/NET0131 ,
		_w456_,
		_w474_,
		_w495_
	);
	LUT4 #(
		.INIT('h153f)
	) name43 (
		\InstQueue_reg[10][2]/NET0131 ,
		\InstQueue_reg[15][2]/NET0131 ,
		_w473_,
		_w471_,
		_w496_
	);
	LUT4 #(
		.INIT('h8000)
	) name44 (
		_w495_,
		_w496_,
		_w493_,
		_w494_,
		_w497_
	);
	LUT4 #(
		.INIT('h135f)
	) name45 (
		\InstQueue_reg[0][2]/NET0131 ,
		\InstQueue_reg[5][2]/NET0131 ,
		_w463_,
		_w467_,
		_w498_
	);
	LUT4 #(
		.INIT('h153f)
	) name46 (
		\InstQueue_reg[12][2]/NET0131 ,
		\InstQueue_reg[9][2]/NET0131 ,
		_w454_,
		_w470_,
		_w499_
	);
	LUT4 #(
		.INIT('h153f)
	) name47 (
		\InstQueue_reg[3][2]/NET0131 ,
		\InstQueue_reg[4][2]/NET0131 ,
		_w464_,
		_w476_,
		_w500_
	);
	LUT4 #(
		.INIT('h153f)
	) name48 (
		\InstQueue_reg[1][2]/NET0131 ,
		\InstQueue_reg[6][2]/NET0131 ,
		_w461_,
		_w453_,
		_w501_
	);
	LUT4 #(
		.INIT('h8000)
	) name49 (
		_w500_,
		_w501_,
		_w498_,
		_w499_,
		_w502_
	);
	LUT2 #(
		.INIT('h8)
	) name50 (
		_w497_,
		_w502_,
		_w503_
	);
	LUT4 #(
		.INIT('h135f)
	) name51 (
		\InstQueue_reg[14][1]/NET0131 ,
		\InstQueue_reg[5][1]/NET0131 ,
		_w460_,
		_w467_,
		_w504_
	);
	LUT4 #(
		.INIT('h135f)
	) name52 (
		\InstQueue_reg[15][1]/NET0131 ,
		\InstQueue_reg[8][1]/NET0131 ,
		_w473_,
		_w468_,
		_w505_
	);
	LUT4 #(
		.INIT('h135f)
	) name53 (
		\InstQueue_reg[0][1]/NET0131 ,
		\InstQueue_reg[1][1]/NET0131 ,
		_w463_,
		_w453_,
		_w506_
	);
	LUT4 #(
		.INIT('h153f)
	) name54 (
		\InstQueue_reg[12][1]/NET0131 ,
		\InstQueue_reg[7][1]/NET0131 ,
		_w477_,
		_w470_,
		_w507_
	);
	LUT4 #(
		.INIT('h8000)
	) name55 (
		_w506_,
		_w507_,
		_w504_,
		_w505_,
		_w508_
	);
	LUT4 #(
		.INIT('h153f)
	) name56 (
		\InstQueue_reg[2][1]/NET0131 ,
		\InstQueue_reg[9][1]/NET0131 ,
		_w454_,
		_w474_,
		_w509_
	);
	LUT4 #(
		.INIT('h135f)
	) name57 (
		\InstQueue_reg[11][1]/NET0131 ,
		\InstQueue_reg[3][1]/NET0131 ,
		_w458_,
		_w476_,
		_w510_
	);
	LUT4 #(
		.INIT('h153f)
	) name58 (
		\InstQueue_reg[10][1]/NET0131 ,
		\InstQueue_reg[6][1]/NET0131 ,
		_w461_,
		_w471_,
		_w511_
	);
	LUT4 #(
		.INIT('h153f)
	) name59 (
		\InstQueue_reg[13][1]/NET0131 ,
		\InstQueue_reg[4][1]/NET0131 ,
		_w464_,
		_w456_,
		_w512_
	);
	LUT4 #(
		.INIT('h8000)
	) name60 (
		_w511_,
		_w512_,
		_w509_,
		_w510_,
		_w513_
	);
	LUT2 #(
		.INIT('h8)
	) name61 (
		_w508_,
		_w513_,
		_w514_
	);
	LUT4 #(
		.INIT('h8000)
	) name62 (
		_w497_,
		_w502_,
		_w508_,
		_w513_,
		_w515_
	);
	LUT4 #(
		.INIT('h153f)
	) name63 (
		\InstQueue_reg[0][3]/NET0131 ,
		\InstQueue_reg[14][3]/NET0131 ,
		_w460_,
		_w463_,
		_w516_
	);
	LUT4 #(
		.INIT('h153f)
	) name64 (
		\InstQueue_reg[12][3]/NET0131 ,
		\InstQueue_reg[5][3]/NET0131 ,
		_w467_,
		_w470_,
		_w517_
	);
	LUT4 #(
		.INIT('h153f)
	) name65 (
		\InstQueue_reg[10][3]/NET0131 ,
		\InstQueue_reg[15][3]/NET0131 ,
		_w473_,
		_w471_,
		_w518_
	);
	LUT4 #(
		.INIT('h153f)
	) name66 (
		\InstQueue_reg[1][3]/NET0131 ,
		\InstQueue_reg[4][3]/NET0131 ,
		_w464_,
		_w453_,
		_w519_
	);
	LUT4 #(
		.INIT('h8000)
	) name67 (
		_w518_,
		_w519_,
		_w516_,
		_w517_,
		_w520_
	);
	LUT4 #(
		.INIT('h153f)
	) name68 (
		\InstQueue_reg[13][3]/NET0131 ,
		\InstQueue_reg[6][3]/NET0131 ,
		_w461_,
		_w456_,
		_w521_
	);
	LUT4 #(
		.INIT('h135f)
	) name69 (
		\InstQueue_reg[3][3]/NET0131 ,
		\InstQueue_reg[7][3]/NET0131 ,
		_w476_,
		_w477_,
		_w522_
	);
	LUT4 #(
		.INIT('h135f)
	) name70 (
		\InstQueue_reg[11][3]/NET0131 ,
		\InstQueue_reg[2][3]/NET0131 ,
		_w458_,
		_w474_,
		_w523_
	);
	LUT4 #(
		.INIT('h153f)
	) name71 (
		\InstQueue_reg[8][3]/NET0131 ,
		\InstQueue_reg[9][3]/NET0131 ,
		_w454_,
		_w468_,
		_w524_
	);
	LUT4 #(
		.INIT('h8000)
	) name72 (
		_w523_,
		_w524_,
		_w521_,
		_w522_,
		_w525_
	);
	LUT4 #(
		.INIT('h153f)
	) name73 (
		\InstQueue_reg[11][0]/NET0131 ,
		\InstQueue_reg[14][0]/NET0131 ,
		_w460_,
		_w458_,
		_w526_
	);
	LUT4 #(
		.INIT('h135f)
	) name74 (
		\InstQueue_reg[6][0]/NET0131 ,
		\InstQueue_reg[9][0]/NET0131 ,
		_w461_,
		_w454_,
		_w527_
	);
	LUT4 #(
		.INIT('h153f)
	) name75 (
		\InstQueue_reg[10][0]/NET0131 ,
		\InstQueue_reg[13][0]/NET0131 ,
		_w456_,
		_w471_,
		_w528_
	);
	LUT4 #(
		.INIT('h135f)
	) name76 (
		\InstQueue_reg[0][0]/NET0131 ,
		\InstQueue_reg[1][0]/NET0131 ,
		_w463_,
		_w453_,
		_w529_
	);
	LUT4 #(
		.INIT('h8000)
	) name77 (
		_w528_,
		_w529_,
		_w526_,
		_w527_,
		_w530_
	);
	LUT4 #(
		.INIT('h135f)
	) name78 (
		\InstQueue_reg[2][0]/NET0131 ,
		\InstQueue_reg[8][0]/NET0131 ,
		_w474_,
		_w468_,
		_w531_
	);
	LUT4 #(
		.INIT('h153f)
	) name79 (
		\InstQueue_reg[12][0]/NET0131 ,
		\InstQueue_reg[15][0]/NET0131 ,
		_w473_,
		_w470_,
		_w532_
	);
	LUT4 #(
		.INIT('h153f)
	) name80 (
		\InstQueue_reg[3][0]/NET0131 ,
		\InstQueue_reg[4][0]/NET0131 ,
		_w464_,
		_w476_,
		_w533_
	);
	LUT4 #(
		.INIT('h153f)
	) name81 (
		\InstQueue_reg[5][0]/NET0131 ,
		\InstQueue_reg[7][0]/NET0131 ,
		_w477_,
		_w467_,
		_w534_
	);
	LUT4 #(
		.INIT('h8000)
	) name82 (
		_w533_,
		_w534_,
		_w531_,
		_w532_,
		_w535_
	);
	LUT4 #(
		.INIT('h8000)
	) name83 (
		_w520_,
		_w525_,
		_w530_,
		_w535_,
		_w536_
	);
	LUT2 #(
		.INIT('h8)
	) name84 (
		_w515_,
		_w536_,
		_w537_
	);
	LUT4 #(
		.INIT('h135f)
	) name85 (
		\InstQueue_reg[1][5]/NET0131 ,
		\InstQueue_reg[5][5]/NET0131 ,
		_w453_,
		_w467_,
		_w538_
	);
	LUT4 #(
		.INIT('h153f)
	) name86 (
		\InstQueue_reg[12][5]/NET0131 ,
		\InstQueue_reg[15][5]/NET0131 ,
		_w473_,
		_w470_,
		_w539_
	);
	LUT4 #(
		.INIT('h135f)
	) name87 (
		\InstQueue_reg[14][5]/NET0131 ,
		\InstQueue_reg[4][5]/NET0131 ,
		_w460_,
		_w464_,
		_w540_
	);
	LUT4 #(
		.INIT('h153f)
	) name88 (
		\InstQueue_reg[10][5]/NET0131 ,
		\InstQueue_reg[2][5]/NET0131 ,
		_w474_,
		_w471_,
		_w541_
	);
	LUT4 #(
		.INIT('h8000)
	) name89 (
		_w540_,
		_w541_,
		_w538_,
		_w539_,
		_w542_
	);
	LUT4 #(
		.INIT('h135f)
	) name90 (
		\InstQueue_reg[0][5]/NET0131 ,
		\InstQueue_reg[13][5]/NET0131 ,
		_w463_,
		_w456_,
		_w543_
	);
	LUT4 #(
		.INIT('h135f)
	) name91 (
		\InstQueue_reg[11][5]/NET0131 ,
		\InstQueue_reg[7][5]/NET0131 ,
		_w458_,
		_w477_,
		_w544_
	);
	LUT4 #(
		.INIT('h135f)
	) name92 (
		\InstQueue_reg[6][5]/NET0131 ,
		\InstQueue_reg[9][5]/NET0131 ,
		_w461_,
		_w454_,
		_w545_
	);
	LUT4 #(
		.INIT('h135f)
	) name93 (
		\InstQueue_reg[3][5]/NET0131 ,
		\InstQueue_reg[8][5]/NET0131 ,
		_w476_,
		_w468_,
		_w546_
	);
	LUT4 #(
		.INIT('h8000)
	) name94 (
		_w545_,
		_w546_,
		_w543_,
		_w544_,
		_w547_
	);
	LUT2 #(
		.INIT('h8)
	) name95 (
		_w542_,
		_w547_,
		_w548_
	);
	LUT4 #(
		.INIT('h8000)
	) name96 (
		_w492_,
		_w515_,
		_w536_,
		_w548_,
		_w549_
	);
	LUT4 #(
		.INIT('h0777)
	) name97 (
		_w520_,
		_w525_,
		_w530_,
		_w535_,
		_w550_
	);
	LUT4 #(
		.INIT('h0888)
	) name98 (
		_w497_,
		_w502_,
		_w508_,
		_w513_,
		_w551_
	);
	LUT2 #(
		.INIT('h8)
	) name99 (
		_w550_,
		_w551_,
		_w552_
	);
	LUT4 #(
		.INIT('h7000)
	) name100 (
		_w466_,
		_w479_,
		_w485_,
		_w490_,
		_w553_
	);
	LUT4 #(
		.INIT('h135f)
	) name101 (
		\InstQueue_reg[11][4]/NET0131 ,
		\InstQueue_reg[3][4]/NET0131 ,
		_w458_,
		_w476_,
		_w554_
	);
	LUT4 #(
		.INIT('h135f)
	) name102 (
		\InstQueue_reg[15][4]/NET0131 ,
		\InstQueue_reg[8][4]/NET0131 ,
		_w473_,
		_w468_,
		_w555_
	);
	LUT4 #(
		.INIT('h153f)
	) name103 (
		\InstQueue_reg[12][4]/NET0131 ,
		\InstQueue_reg[14][4]/NET0131 ,
		_w460_,
		_w470_,
		_w556_
	);
	LUT4 #(
		.INIT('h135f)
	) name104 (
		\InstQueue_reg[1][4]/NET0131 ,
		\InstQueue_reg[2][4]/NET0131 ,
		_w453_,
		_w474_,
		_w557_
	);
	LUT4 #(
		.INIT('h8000)
	) name105 (
		_w556_,
		_w557_,
		_w554_,
		_w555_,
		_w558_
	);
	LUT4 #(
		.INIT('h135f)
	) name106 (
		\InstQueue_reg[0][4]/NET0131 ,
		\InstQueue_reg[5][4]/NET0131 ,
		_w463_,
		_w467_,
		_w559_
	);
	LUT4 #(
		.INIT('h153f)
	) name107 (
		\InstQueue_reg[10][4]/NET0131 ,
		\InstQueue_reg[7][4]/NET0131 ,
		_w477_,
		_w471_,
		_w560_
	);
	LUT4 #(
		.INIT('h153f)
	) name108 (
		\InstQueue_reg[13][4]/NET0131 ,
		\InstQueue_reg[6][4]/NET0131 ,
		_w461_,
		_w456_,
		_w561_
	);
	LUT4 #(
		.INIT('h135f)
	) name109 (
		\InstQueue_reg[4][4]/NET0131 ,
		\InstQueue_reg[9][4]/NET0131 ,
		_w464_,
		_w454_,
		_w562_
	);
	LUT4 #(
		.INIT('h8000)
	) name110 (
		_w561_,
		_w562_,
		_w559_,
		_w560_,
		_w563_
	);
	LUT2 #(
		.INIT('h8)
	) name111 (
		_w558_,
		_w563_,
		_w564_
	);
	LUT4 #(
		.INIT('h8000)
	) name112 (
		_w542_,
		_w547_,
		_w558_,
		_w563_,
		_w565_
	);
	LUT4 #(
		.INIT('h8000)
	) name113 (
		_w550_,
		_w551_,
		_w553_,
		_w565_,
		_w566_
	);
	LUT4 #(
		.INIT('h7000)
	) name114 (
		_w542_,
		_w547_,
		_w558_,
		_w563_,
		_w567_
	);
	LUT2 #(
		.INIT('h4)
	) name115 (
		_w503_,
		_w536_,
		_w568_
	);
	LUT4 #(
		.INIT('h2000)
	) name116 (
		_w492_,
		_w503_,
		_w536_,
		_w567_,
		_w569_
	);
	LUT4 #(
		.INIT('h8000)
	) name117 (
		_w515_,
		_w550_,
		_w553_,
		_w565_,
		_w570_
	);
	LUT3 #(
		.INIT('h01)
	) name118 (
		_w566_,
		_w569_,
		_w570_,
		_w571_
	);
	LUT4 #(
		.INIT('h0001)
	) name119 (
		_w549_,
		_w566_,
		_w569_,
		_w570_,
		_w572_
	);
	LUT4 #(
		.INIT('h8000)
	) name120 (
		_w492_,
		_w515_,
		_w550_,
		_w567_,
		_w573_
	);
	LUT4 #(
		.INIT('h8000)
	) name121 (
		_w492_,
		_w550_,
		_w551_,
		_w567_,
		_w574_
	);
	LUT2 #(
		.INIT('h1)
	) name122 (
		_w573_,
		_w574_,
		_w575_
	);
	LUT3 #(
		.INIT('h04)
	) name123 (
		_w548_,
		_w553_,
		_w564_,
		_w576_
	);
	LUT2 #(
		.INIT('h8)
	) name124 (
		_w552_,
		_w576_,
		_w577_
	);
	LUT4 #(
		.INIT('h7000)
	) name125 (
		_w520_,
		_w525_,
		_w530_,
		_w535_,
		_w578_
	);
	LUT2 #(
		.INIT('h8)
	) name126 (
		_w515_,
		_w578_,
		_w579_
	);
	LUT2 #(
		.INIT('h8)
	) name127 (
		_w576_,
		_w579_,
		_w580_
	);
	LUT3 #(
		.INIT('h37)
	) name128 (
		_w552_,
		_w576_,
		_w579_,
		_w581_
	);
	LUT3 #(
		.INIT('h80)
	) name129 (
		_w572_,
		_w575_,
		_w581_,
		_w582_
	);
	LUT4 #(
		.INIT('h8000)
	) name130 (
		_w466_,
		_w479_,
		_w485_,
		_w490_,
		_w583_
	);
	LUT3 #(
		.INIT('h80)
	) name131 (
		_w514_,
		_w565_,
		_w583_,
		_w584_
	);
	LUT4 #(
		.INIT('h0888)
	) name132 (
		_w466_,
		_w479_,
		_w485_,
		_w490_,
		_w585_
	);
	LUT3 #(
		.INIT('h40)
	) name133 (
		_w514_,
		_w567_,
		_w585_,
		_w586_
	);
	LUT3 #(
		.INIT('ha8)
	) name134 (
		_w568_,
		_w584_,
		_w586_,
		_w587_
	);
	LUT4 #(
		.INIT('hd9fb)
	) name135 (
		_w480_,
		_w491_,
		_w564_,
		_w565_,
		_w588_
	);
	LUT4 #(
		.INIT('h0888)
	) name136 (
		_w520_,
		_w525_,
		_w530_,
		_w535_,
		_w589_
	);
	LUT4 #(
		.INIT('h8000)
	) name137 (
		_w551_,
		_w565_,
		_w585_,
		_w589_,
		_w590_
	);
	LUT3 #(
		.INIT('h0d)
	) name138 (
		_w537_,
		_w588_,
		_w590_,
		_w591_
	);
	LUT4 #(
		.INIT('h8000)
	) name139 (
		_w492_,
		_w551_,
		_w567_,
		_w578_,
		_w592_
	);
	LUT2 #(
		.INIT('h4)
	) name140 (
		_w503_,
		_w589_,
		_w593_
	);
	LUT3 #(
		.INIT('h13)
	) name141 (
		_w584_,
		_w592_,
		_w593_,
		_w594_
	);
	LUT3 #(
		.INIT('h40)
	) name142 (
		_w587_,
		_w591_,
		_w594_,
		_w595_
	);
	LUT4 #(
		.INIT('h8421)
	) name143 (
		\InstQueueRd_Addr_reg[0]/NET0131 ,
		\InstQueueRd_Addr_reg[1]/NET0131 ,
		\InstQueueWr_Addr_reg[0]/NET0131 ,
		\InstQueueWr_Addr_reg[1]/NET0131 ,
		_w596_
	);
	LUT4 #(
		.INIT('h08ce)
	) name144 (
		\InstQueueRd_Addr_reg[0]/NET0131 ,
		\InstQueueRd_Addr_reg[1]/NET0131 ,
		\InstQueueWr_Addr_reg[0]/NET0131 ,
		\InstQueueWr_Addr_reg[1]/NET0131 ,
		_w597_
	);
	LUT2 #(
		.INIT('h9)
	) name145 (
		\InstQueueRd_Addr_reg[2]/NET0131 ,
		\InstQueueWr_Addr_reg[2]/NET0131 ,
		_w598_
	);
	LUT3 #(
		.INIT('h41)
	) name146 (
		_w596_,
		_w597_,
		_w598_,
		_w599_
	);
	LUT2 #(
		.INIT('h4)
	) name147 (
		\InstQueueRd_Addr_reg[3]/NET0131 ,
		\InstQueueWr_Addr_reg[3]/NET0131 ,
		_w600_
	);
	LUT2 #(
		.INIT('h2)
	) name148 (
		\InstQueueRd_Addr_reg[3]/NET0131 ,
		\InstQueueWr_Addr_reg[3]/NET0131 ,
		_w601_
	);
	LUT2 #(
		.INIT('h9)
	) name149 (
		\InstQueueRd_Addr_reg[3]/NET0131 ,
		\InstQueueWr_Addr_reg[3]/NET0131 ,
		_w602_
	);
	LUT3 #(
		.INIT('hb2)
	) name150 (
		\InstQueueRd_Addr_reg[2]/NET0131 ,
		\InstQueueWr_Addr_reg[2]/NET0131 ,
		_w597_,
		_w603_
	);
	LUT4 #(
		.INIT('h004d)
	) name151 (
		\InstQueueRd_Addr_reg[2]/NET0131 ,
		\InstQueueWr_Addr_reg[2]/NET0131 ,
		_w597_,
		_w601_,
		_w604_
	);
	LUT4 #(
		.INIT('h40d4)
	) name152 (
		\InstQueueRd_Addr_reg[3]/NET0131 ,
		\InstQueueWr_Addr_reg[3]/NET0131 ,
		_w599_,
		_w603_,
		_w605_
	);
	LUT4 #(
		.INIT('hc800)
	) name153 (
		_w552_,
		_w576_,
		_w579_,
		_w605_,
		_w606_
	);
	LUT2 #(
		.INIT('h9)
	) name154 (
		\InstQueueRd_Addr_reg[0]/NET0131 ,
		\InstQueueRd_Addr_reg[1]/NET0131 ,
		_w607_
	);
	LUT4 #(
		.INIT('h00fb)
	) name155 (
		_w582_,
		_w595_,
		_w606_,
		_w607_,
		_w608_
	);
	LUT4 #(
		.INIT('h4920)
	) name156 (
		\InstQueueRd_Addr_reg[2]/NET0131 ,
		\InstQueueWr_Addr_reg[2]/NET0131 ,
		_w597_,
		_w602_,
		_w609_
	);
	LUT4 #(
		.INIT('h39c6)
	) name157 (
		\InstQueueRd_Addr_reg[0]/NET0131 ,
		\InstQueueRd_Addr_reg[1]/NET0131 ,
		\InstQueueWr_Addr_reg[0]/NET0131 ,
		\InstQueueWr_Addr_reg[1]/NET0131 ,
		_w610_
	);
	LUT4 #(
		.INIT('hee0e)
	) name158 (
		_w600_,
		_w604_,
		_w609_,
		_w610_,
		_w611_
	);
	LUT2 #(
		.INIT('h4)
	) name159 (
		READY_n_pad,
		_w611_,
		_w612_
	);
	LUT3 #(
		.INIT('h0b)
	) name160 (
		_w514_,
		_w569_,
		_w570_,
		_w613_
	);
	LUT2 #(
		.INIT('h4)
	) name161 (
		\State_reg[0]/NET0131 ,
		\State_reg[1]/NET0131 ,
		_w614_
	);
	LUT3 #(
		.INIT('h04)
	) name162 (
		\State_reg[0]/NET0131 ,
		\State_reg[1]/NET0131 ,
		\State_reg[2]/NET0131 ,
		_w615_
	);
	LUT3 #(
		.INIT('h10)
	) name163 (
		\State_reg[0]/NET0131 ,
		\State_reg[1]/NET0131 ,
		\State_reg[2]/NET0131 ,
		_w616_
	);
	LUT3 #(
		.INIT('heb)
	) name164 (
		\State_reg[0]/NET0131 ,
		\State_reg[1]/NET0131 ,
		\State_reg[2]/NET0131 ,
		_w617_
	);
	LUT4 #(
		.INIT('h00f4)
	) name165 (
		_w514_,
		_w569_,
		_w570_,
		_w617_,
		_w618_
	);
	LUT3 #(
		.INIT('h13)
	) name166 (
		_w514_,
		_w566_,
		_w569_,
		_w619_
	);
	LUT4 #(
		.INIT('h1511)
	) name167 (
		_w549_,
		_w612_,
		_w618_,
		_w619_,
		_w620_
	);
	LUT4 #(
		.INIT('hf400)
	) name168 (
		_w514_,
		_w569_,
		_w570_,
		_w617_,
		_w621_
	);
	LUT3 #(
		.INIT('h0e)
	) name169 (
		_w569_,
		_w570_,
		_w612_,
		_w622_
	);
	LUT2 #(
		.INIT('h2)
	) name170 (
		_w566_,
		_w612_,
		_w623_
	);
	LUT3 #(
		.INIT('h01)
	) name171 (
		_w621_,
		_w622_,
		_w623_,
		_w624_
	);
	LUT4 #(
		.INIT('h00c8)
	) name172 (
		_w552_,
		_w576_,
		_w579_,
		_w605_,
		_w625_
	);
	LUT2 #(
		.INIT('h2)
	) name173 (
		_w575_,
		_w625_,
		_w626_
	);
	LUT4 #(
		.INIT('h27af)
	) name174 (
		\InstQueueRd_Addr_reg[1]/NET0131 ,
		_w626_,
		_w620_,
		_w624_,
		_w627_
	);
	LUT2 #(
		.INIT('h1)
	) name175 (
		_w608_,
		_w627_,
		_w628_
	);
	LUT4 #(
		.INIT('h0010)
	) name176 (
		\InstQueueRd_Addr_reg[0]/NET0131 ,
		_w582_,
		_w595_,
		_w606_,
		_w629_
	);
	LUT4 #(
		.INIT('h0080)
	) name177 (
		\InstQueueRd_Addr_reg[0]/NET0131 ,
		_w572_,
		_w575_,
		_w625_,
		_w630_
	);
	LUT4 #(
		.INIT('h1113)
	) name178 (
		\InstQueueWr_Addr_reg[0]/NET0131 ,
		\InstQueueWr_Addr_reg[1]/NET0131 ,
		_w629_,
		_w630_,
		_w631_
	);
	LUT2 #(
		.INIT('h2)
	) name179 (
		_w628_,
		_w631_,
		_w632_
	);
	LUT4 #(
		.INIT('h0110)
	) name180 (
		READY_n_pad,
		\State_reg[0]/NET0131 ,
		\State_reg[1]/NET0131 ,
		\State_reg[2]/NET0131 ,
		_w633_
	);
	LUT2 #(
		.INIT('h8)
	) name181 (
		_w611_,
		_w633_,
		_w634_
	);
	LUT3 #(
		.INIT('h08)
	) name182 (
		_w514_,
		_w569_,
		_w612_,
		_w635_
	);
	LUT4 #(
		.INIT('hff13)
	) name183 (
		_w514_,
		_w566_,
		_w569_,
		_w612_,
		_w636_
	);
	LUT3 #(
		.INIT('h13)
	) name184 (
		_w613_,
		_w634_,
		_w636_,
		_w637_
	);
	LUT3 #(
		.INIT('h07)
	) name185 (
		\InstQueueRd_Addr_reg[0]/NET0131 ,
		\InstQueueRd_Addr_reg[1]/NET0131 ,
		\InstQueueRd_Addr_reg[2]/NET0131 ,
		_w638_
	);
	LUT2 #(
		.INIT('h2)
	) name186 (
		_w605_,
		_w638_,
		_w639_
	);
	LUT4 #(
		.INIT('h00c8)
	) name187 (
		_w552_,
		_w576_,
		_w579_,
		_w639_,
		_w640_
	);
	LUT2 #(
		.INIT('h2)
	) name188 (
		_w575_,
		_w640_,
		_w641_
	);
	LUT3 #(
		.INIT('h8a)
	) name189 (
		\InstQueueRd_Addr_reg[3]/NET0131 ,
		_w637_,
		_w641_,
		_w642_
	);
	LUT4 #(
		.INIT('hec00)
	) name190 (
		_w514_,
		_w566_,
		_w569_,
		_w611_,
		_w643_
	);
	LUT4 #(
		.INIT('hf400)
	) name191 (
		_w514_,
		_w569_,
		_w570_,
		_w634_,
		_w644_
	);
	LUT4 #(
		.INIT('h0203)
	) name192 (
		READY_n_pad,
		_w549_,
		_w644_,
		_w643_,
		_w645_
	);
	LUT3 #(
		.INIT('h78)
	) name193 (
		\InstQueueRd_Addr_reg[1]/NET0131 ,
		\InstQueueRd_Addr_reg[2]/NET0131 ,
		\InstQueueRd_Addr_reg[3]/NET0131 ,
		_w646_
	);
	LUT2 #(
		.INIT('h4)
	) name194 (
		_w645_,
		_w646_,
		_w647_
	);
	LUT4 #(
		.INIT('h807f)
	) name195 (
		\InstQueueRd_Addr_reg[0]/NET0131 ,
		\InstQueueRd_Addr_reg[1]/NET0131 ,
		\InstQueueRd_Addr_reg[2]/NET0131 ,
		\InstQueueRd_Addr_reg[3]/NET0131 ,
		_w648_
	);
	LUT3 #(
		.INIT('h04)
	) name196 (
		\InstQueueRd_Addr_reg[3]/NET0131 ,
		_w605_,
		_w638_,
		_w649_
	);
	LUT4 #(
		.INIT('hc800)
	) name197 (
		_w552_,
		_w576_,
		_w579_,
		_w649_,
		_w650_
	);
	LUT4 #(
		.INIT('h00f4)
	) name198 (
		_w582_,
		_w595_,
		_w648_,
		_w650_,
		_w651_
	);
	LUT3 #(
		.INIT('h10)
	) name199 (
		_w647_,
		_w642_,
		_w651_,
		_w652_
	);
	LUT4 #(
		.INIT('h0200)
	) name200 (
		\InstQueueWr_Addr_reg[3]/NET0131 ,
		_w647_,
		_w642_,
		_w651_,
		_w653_
	);
	LUT4 #(
		.INIT('h8880)
	) name201 (
		\InstQueueWr_Addr_reg[0]/NET0131 ,
		\InstQueueWr_Addr_reg[1]/NET0131 ,
		_w629_,
		_w630_,
		_w654_
	);
	LUT3 #(
		.INIT('h78)
	) name202 (
		\InstQueueRd_Addr_reg[0]/NET0131 ,
		\InstQueueRd_Addr_reg[1]/NET0131 ,
		\InstQueueRd_Addr_reg[2]/NET0131 ,
		_w655_
	);
	LUT3 #(
		.INIT('hb0)
	) name203 (
		_w582_,
		_w595_,
		_w655_,
		_w656_
	);
	LUT2 #(
		.INIT('h6)
	) name204 (
		\InstQueueRd_Addr_reg[1]/NET0131 ,
		\InstQueueRd_Addr_reg[2]/NET0131 ,
		_w657_
	);
	LUT3 #(
		.INIT('hc6)
	) name205 (
		\InstQueueRd_Addr_reg[1]/NET0131 ,
		\InstQueueRd_Addr_reg[2]/NET0131 ,
		READY_n_pad,
		_w658_
	);
	LUT2 #(
		.INIT('h2)
	) name206 (
		_w611_,
		_w617_,
		_w659_
	);
	LUT3 #(
		.INIT('h02)
	) name207 (
		_w611_,
		_w617_,
		_w658_,
		_w660_
	);
	LUT3 #(
		.INIT('h51)
	) name208 (
		\InstQueueRd_Addr_reg[2]/NET0131 ,
		_w611_,
		_w617_,
		_w661_
	);
	LUT4 #(
		.INIT('h00f4)
	) name209 (
		_w514_,
		_w569_,
		_w570_,
		_w661_,
		_w662_
	);
	LUT2 #(
		.INIT('h4)
	) name210 (
		_w660_,
		_w662_,
		_w663_
	);
	LUT3 #(
		.INIT('he2)
	) name211 (
		\InstQueueRd_Addr_reg[2]/NET0131 ,
		_w611_,
		_w658_,
		_w664_
	);
	LUT4 #(
		.INIT('hec00)
	) name212 (
		_w514_,
		_w566_,
		_w569_,
		_w664_,
		_w665_
	);
	LUT2 #(
		.INIT('h8)
	) name213 (
		_w549_,
		_w657_,
		_w666_
	);
	LUT3 #(
		.INIT('h2e)
	) name214 (
		\InstQueueRd_Addr_reg[2]/NET0131 ,
		_w605_,
		_w655_,
		_w667_
	);
	LUT4 #(
		.INIT('hc800)
	) name215 (
		_w552_,
		_w576_,
		_w579_,
		_w667_,
		_w668_
	);
	LUT3 #(
		.INIT('ha8)
	) name216 (
		\InstQueueRd_Addr_reg[2]/NET0131 ,
		_w573_,
		_w574_,
		_w669_
	);
	LUT4 #(
		.INIT('h0001)
	) name217 (
		_w665_,
		_w668_,
		_w666_,
		_w669_,
		_w670_
	);
	LUT2 #(
		.INIT('h4)
	) name218 (
		_w663_,
		_w670_,
		_w671_
	);
	LUT3 #(
		.INIT('h20)
	) name219 (
		\InstQueueWr_Addr_reg[2]/NET0131 ,
		_w656_,
		_w671_,
		_w672_
	);
	LUT3 #(
		.INIT('h01)
	) name220 (
		_w654_,
		_w653_,
		_w672_,
		_w673_
	);
	LUT3 #(
		.INIT('h45)
	) name221 (
		\InstQueueWr_Addr_reg[2]/NET0131 ,
		_w656_,
		_w671_,
		_w674_
	);
	LUT2 #(
		.INIT('h4)
	) name222 (
		_w653_,
		_w674_,
		_w675_
	);
	LUT3 #(
		.INIT('h20)
	) name223 (
		\InstQueueWr_Addr_reg[3]/NET0131 ,
		_w656_,
		_w671_,
		_w676_
	);
	LUT2 #(
		.INIT('h2)
	) name224 (
		\More_reg/NET0131 ,
		_w633_,
		_w677_
	);
	LUT2 #(
		.INIT('h2)
	) name225 (
		_w611_,
		_w677_,
		_w678_
	);
	LUT3 #(
		.INIT('h07)
	) name226 (
		_w613_,
		_w636_,
		_w678_,
		_w679_
	);
	LUT4 #(
		.INIT('h1842)
	) name227 (
		\InstQueueRd_Addr_reg[0]/NET0131 ,
		\InstQueueRd_Addr_reg[1]/NET0131 ,
		\InstQueueWr_Addr_reg[0]/NET0131 ,
		\InstQueueWr_Addr_reg[1]/NET0131 ,
		_w680_
	);
	LUT4 #(
		.INIT('hee0e)
	) name228 (
		_w600_,
		_w604_,
		_w609_,
		_w680_,
		_w681_
	);
	LUT2 #(
		.INIT('h2)
	) name229 (
		_w574_,
		_w681_,
		_w682_
	);
	LUT2 #(
		.INIT('h2)
	) name230 (
		_w573_,
		_w605_,
		_w683_
	);
	LUT2 #(
		.INIT('h1)
	) name231 (
		_w625_,
		_w683_,
		_w684_
	);
	LUT3 #(
		.INIT('h01)
	) name232 (
		_w625_,
		_w682_,
		_w683_,
		_w685_
	);
	LUT4 #(
		.INIT('haaa8)
	) name233 (
		READY_n_pad,
		_w566_,
		_w569_,
		_w570_,
		_w686_
	);
	LUT2 #(
		.INIT('h8)
	) name234 (
		\Flush_reg/NET0131 ,
		_w611_,
		_w687_
	);
	LUT2 #(
		.INIT('h8)
	) name235 (
		_w573_,
		_w605_,
		_w688_
	);
	LUT4 #(
		.INIT('h135f)
	) name236 (
		_w573_,
		_w574_,
		_w605_,
		_w681_,
		_w689_
	);
	LUT4 #(
		.INIT('h1f00)
	) name237 (
		_w621_,
		_w686_,
		_w687_,
		_w689_,
		_w690_
	);
	LUT3 #(
		.INIT('h40)
	) name238 (
		_w679_,
		_w685_,
		_w690_,
		_w691_
	);
	LUT3 #(
		.INIT('he0)
	) name239 (
		_w652_,
		_w676_,
		_w691_,
		_w692_
	);
	LUT4 #(
		.INIT('h0b00)
	) name240 (
		_w632_,
		_w673_,
		_w675_,
		_w692_,
		_w693_
	);
	LUT3 #(
		.INIT('h40)
	) name241 (
		\DataWidth_reg[1]/NET0131 ,
		_w570_,
		_w634_,
		_w694_
	);
	LUT4 #(
		.INIT('h0020)
	) name242 (
		\State2_reg[0]/NET0131 ,
		\State2_reg[1]/NET0131 ,
		\State2_reg[2]/NET0131 ,
		\State2_reg[3]/NET0131 ,
		_w695_
	);
	LUT4 #(
		.INIT('h0040)
	) name243 (
		\State2_reg[0]/NET0131 ,
		\State2_reg[1]/NET0131 ,
		\State2_reg[2]/NET0131 ,
		\State2_reg[3]/NET0131 ,
		_w696_
	);
	LUT4 #(
		.INIT('h0008)
	) name244 (
		\State2_reg[0]/NET0131 ,
		\State2_reg[1]/NET0131 ,
		\State2_reg[2]/NET0131 ,
		\State2_reg[3]/NET0131 ,
		_w697_
	);
	LUT4 #(
		.INIT('hffb7)
	) name245 (
		\State2_reg[0]/NET0131 ,
		\State2_reg[1]/NET0131 ,
		\State2_reg[2]/NET0131 ,
		\State2_reg[3]/NET0131 ,
		_w698_
	);
	LUT2 #(
		.INIT('h2)
	) name246 (
		READY_n_pad,
		_w698_,
		_w699_
	);
	LUT4 #(
		.INIT('h0004)
	) name247 (
		\State2_reg[0]/NET0131 ,
		\State2_reg[1]/NET0131 ,
		\State2_reg[2]/NET0131 ,
		\State2_reg[3]/NET0131 ,
		_w700_
	);
	LUT4 #(
		.INIT('h0002)
	) name248 (
		\State2_reg[0]/NET0131 ,
		\State2_reg[1]/NET0131 ,
		\State2_reg[2]/NET0131 ,
		\State2_reg[3]/NET0131 ,
		_w701_
	);
	LUT4 #(
		.INIT('h8caf)
	) name249 (
		\DataWidth_reg[1]/NET0131 ,
		READY_n_pad,
		_w700_,
		_w701_,
		_w702_
	);
	LUT2 #(
		.INIT('h4)
	) name250 (
		_w699_,
		_w702_,
		_w703_
	);
	LUT4 #(
		.INIT('hd0ff)
	) name251 (
		_w693_,
		_w694_,
		_w695_,
		_w703_,
		_w704_
	);
	LUT2 #(
		.INIT('h1)
	) name252 (
		\State2_reg[0]/NET0131 ,
		\State2_reg[3]/NET0131 ,
		_w705_
	);
	LUT4 #(
		.INIT('h0010)
	) name253 (
		\State2_reg[0]/NET0131 ,
		\State2_reg[1]/NET0131 ,
		\State2_reg[2]/NET0131 ,
		\State2_reg[3]/NET0131 ,
		_w706_
	);
	LUT2 #(
		.INIT('h8)
	) name254 (
		\DataWidth_reg[1]/NET0131 ,
		_w700_,
		_w707_
	);
	LUT3 #(
		.INIT('h07)
	) name255 (
		\DataWidth_reg[1]/NET0131 ,
		_w700_,
		_w706_,
		_w708_
	);
	LUT4 #(
		.INIT('hff9f)
	) name256 (
		\State2_reg[0]/NET0131 ,
		\State2_reg[1]/NET0131 ,
		\State2_reg[2]/NET0131 ,
		\State2_reg[3]/NET0131 ,
		_w709_
	);
	LUT3 #(
		.INIT('hb0)
	) name257 (
		READY_n_pad,
		_w697_,
		_w709_,
		_w710_
	);
	LUT2 #(
		.INIT('h7)
	) name258 (
		_w708_,
		_w710_,
		_w711_
	);
	LUT4 #(
		.INIT('h0080)
	) name259 (
		\State2_reg[0]/NET0131 ,
		\State2_reg[1]/NET0131 ,
		\State2_reg[2]/NET0131 ,
		\State2_reg[3]/NET0131 ,
		_w712_
	);
	LUT2 #(
		.INIT('h4)
	) name260 (
		\Flush_reg/NET0131 ,
		\InstQueueRd_Addr_reg[2]/NET0131 ,
		_w713_
	);
	LUT3 #(
		.INIT('he0)
	) name261 (
		\InstQueueRd_Addr_reg[0]/NET0131 ,
		\InstQueueRd_Addr_reg[1]/NET0131 ,
		\InstQueueRd_Addr_reg[3]/NET0131 ,
		_w714_
	);
	LUT3 #(
		.INIT('h2a)
	) name262 (
		_w712_,
		_w713_,
		_w714_,
		_w715_
	);
	LUT4 #(
		.INIT('h0008)
	) name263 (
		READY_n_pad,
		\State2_reg[0]/NET0131 ,
		\State2_reg[2]/NET0131 ,
		\State2_reg[3]/NET0131 ,
		_w716_
	);
	LUT3 #(
		.INIT('h80)
	) name264 (
		READY_n_pad,
		\State2_reg[1]/NET0131 ,
		\State2_reg[2]/NET0131 ,
		_w717_
	);
	LUT4 #(
		.INIT('h0200)
	) name265 (
		\State2_reg[0]/NET0131 ,
		\State2_reg[1]/NET0131 ,
		\State2_reg[2]/NET0131 ,
		\State2_reg[3]/NET0131 ,
		_w718_
	);
	LUT4 #(
		.INIT('h000d)
	) name266 (
		_w705_,
		_w717_,
		_w718_,
		_w716_,
		_w719_
	);
	LUT2 #(
		.INIT('h4)
	) name267 (
		_w715_,
		_w719_,
		_w720_
	);
	LUT4 #(
		.INIT('h70ff)
	) name268 (
		_w693_,
		_w694_,
		_w695_,
		_w720_,
		_w721_
	);
	LUT4 #(
		.INIT('h0100)
	) name269 (
		\State2_reg[0]/NET0131 ,
		\State2_reg[1]/NET0131 ,
		\State2_reg[2]/NET0131 ,
		\State2_reg[3]/NET0131 ,
		_w722_
	);
	LUT4 #(
		.INIT('h0180)
	) name270 (
		\State2_reg[0]/NET0131 ,
		\State2_reg[1]/NET0131 ,
		\State2_reg[2]/NET0131 ,
		\State2_reg[3]/NET0131 ,
		_w723_
	);
	LUT3 #(
		.INIT('h80)
	) name271 (
		\InstAddrPointer_reg[1]/NET0131 ,
		\InstAddrPointer_reg[2]/NET0131 ,
		\InstAddrPointer_reg[3]/NET0131 ,
		_w724_
	);
	LUT4 #(
		.INIT('h8000)
	) name272 (
		\InstAddrPointer_reg[1]/NET0131 ,
		\InstAddrPointer_reg[2]/NET0131 ,
		\InstAddrPointer_reg[3]/NET0131 ,
		\InstAddrPointer_reg[4]/NET0131 ,
		_w725_
	);
	LUT2 #(
		.INIT('h8)
	) name273 (
		\InstAddrPointer_reg[5]/NET0131 ,
		\InstAddrPointer_reg[6]/NET0131 ,
		_w726_
	);
	LUT4 #(
		.INIT('h8000)
	) name274 (
		\InstAddrPointer_reg[7]/NET0131 ,
		\InstAddrPointer_reg[8]/NET0131 ,
		_w725_,
		_w726_,
		_w727_
	);
	LUT3 #(
		.INIT('h80)
	) name275 (
		\InstAddrPointer_reg[10]/NET0131 ,
		\InstAddrPointer_reg[9]/NET0131 ,
		_w727_,
		_w728_
	);
	LUT2 #(
		.INIT('h8)
	) name276 (
		\InstAddrPointer_reg[10]/NET0131 ,
		\InstAddrPointer_reg[11]/NET0131 ,
		_w729_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name277 (
		\InstAddrPointer_reg[10]/NET0131 ,
		\InstAddrPointer_reg[11]/NET0131 ,
		\InstAddrPointer_reg[9]/NET0131 ,
		_w727_,
		_w730_
	);
	LUT2 #(
		.INIT('h8)
	) name278 (
		\InstAddrPointer_reg[12]/NET0131 ,
		_w730_,
		_w731_
	);
	LUT3 #(
		.INIT('h80)
	) name279 (
		\InstAddrPointer_reg[12]/NET0131 ,
		\InstAddrPointer_reg[13]/NET0131 ,
		_w730_,
		_w732_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name280 (
		\InstAddrPointer_reg[7]/NET0131 ,
		\InstAddrPointer_reg[8]/NET0131 ,
		_w725_,
		_w726_,
		_w733_
	);
	LUT2 #(
		.INIT('h8)
	) name281 (
		\InstAddrPointer_reg[9]/NET0131 ,
		_w733_,
		_w734_
	);
	LUT3 #(
		.INIT('h80)
	) name282 (
		\InstAddrPointer_reg[10]/NET0131 ,
		\InstAddrPointer_reg[9]/NET0131 ,
		_w733_,
		_w735_
	);
	LUT4 #(
		.INIT('h8000)
	) name283 (
		\InstAddrPointer_reg[12]/NET0131 ,
		\InstAddrPointer_reg[13]/NET0131 ,
		_w730_,
		_w735_,
		_w736_
	);
	LUT4 #(
		.INIT('h8007)
	) name284 (
		\InstQueueRd_Addr_reg[0]/NET0131 ,
		\InstQueueRd_Addr_reg[1]/NET0131 ,
		\InstQueueRd_Addr_reg[2]/NET0131 ,
		\InstQueueRd_Addr_reg[3]/NET0131 ,
		_w737_
	);
	LUT4 #(
		.INIT('hcdef)
	) name285 (
		\InstQueueRd_Addr_reg[0]/NET0131 ,
		\InstQueueRd_Addr_reg[1]/NET0131 ,
		\InstQueue_reg[1][3]/NET0131 ,
		\InstQueue_reg[2][3]/NET0131 ,
		_w738_
	);
	LUT2 #(
		.INIT('h2)
	) name286 (
		_w737_,
		_w738_,
		_w739_
	);
	LUT4 #(
		.INIT('h135f)
	) name287 (
		\InstQueue_reg[0][3]/NET0131 ,
		\InstQueue_reg[13][3]/NET0131 ,
		_w473_,
		_w470_,
		_w740_
	);
	LUT4 #(
		.INIT('h135f)
	) name288 (
		\InstQueue_reg[4][3]/NET0131 ,
		\InstQueue_reg[9][3]/NET0131 ,
		_w476_,
		_w468_,
		_w741_
	);
	LUT4 #(
		.INIT('h135f)
	) name289 (
		\InstQueue_reg[14][3]/NET0131 ,
		\InstQueue_reg[3][3]/NET0131 ,
		_w456_,
		_w474_,
		_w742_
	);
	LUT3 #(
		.INIT('h80)
	) name290 (
		_w740_,
		_w741_,
		_w742_,
		_w743_
	);
	LUT4 #(
		.INIT('h135f)
	) name291 (
		\InstQueue_reg[5][3]/NET0131 ,
		\InstQueue_reg[8][3]/NET0131 ,
		_w464_,
		_w477_,
		_w744_
	);
	LUT4 #(
		.INIT('h135f)
	) name292 (
		\InstQueue_reg[12][3]/NET0131 ,
		\InstQueue_reg[6][3]/NET0131 ,
		_w458_,
		_w467_,
		_w745_
	);
	LUT4 #(
		.INIT('h153f)
	) name293 (
		\InstQueue_reg[11][3]/NET0131 ,
		\InstQueue_reg[7][3]/NET0131 ,
		_w461_,
		_w471_,
		_w746_
	);
	LUT4 #(
		.INIT('h153f)
	) name294 (
		\InstQueue_reg[10][3]/NET0131 ,
		\InstQueue_reg[15][3]/NET0131 ,
		_w460_,
		_w454_,
		_w747_
	);
	LUT4 #(
		.INIT('h8000)
	) name295 (
		_w746_,
		_w747_,
		_w744_,
		_w745_,
		_w748_
	);
	LUT3 #(
		.INIT('h40)
	) name296 (
		_w739_,
		_w743_,
		_w748_,
		_w749_
	);
	LUT3 #(
		.INIT('h78)
	) name297 (
		\InstAddrPointer_reg[1]/NET0131 ,
		\InstAddrPointer_reg[2]/NET0131 ,
		\InstAddrPointer_reg[3]/NET0131 ,
		_w750_
	);
	LUT4 #(
		.INIT('h0040)
	) name298 (
		_w739_,
		_w743_,
		_w748_,
		_w750_,
		_w751_
	);
	LUT2 #(
		.INIT('h6)
	) name299 (
		\InstAddrPointer_reg[1]/NET0131 ,
		\InstAddrPointer_reg[2]/NET0131 ,
		_w752_
	);
	LUT4 #(
		.INIT('h135f)
	) name300 (
		\InstQueue_reg[10][2]/NET0131 ,
		\InstQueue_reg[6][2]/NET0131 ,
		_w454_,
		_w467_,
		_w753_
	);
	LUT4 #(
		.INIT('h153f)
	) name301 (
		\InstQueue_reg[11][2]/NET0131 ,
		\InstQueue_reg[12][2]/NET0131 ,
		_w458_,
		_w471_,
		_w754_
	);
	LUT4 #(
		.INIT('h153f)
	) name302 (
		\InstQueue_reg[14][2]/NET0131 ,
		\InstQueue_reg[15][2]/NET0131 ,
		_w460_,
		_w456_,
		_w755_
	);
	LUT4 #(
		.INIT('h135f)
	) name303 (
		\InstQueue_reg[2][2]/NET0131 ,
		\InstQueue_reg[9][2]/NET0131 ,
		_w453_,
		_w468_,
		_w756_
	);
	LUT4 #(
		.INIT('h8000)
	) name304 (
		_w755_,
		_w756_,
		_w753_,
		_w754_,
		_w757_
	);
	LUT4 #(
		.INIT('h135f)
	) name305 (
		\InstQueue_reg[3][2]/NET0131 ,
		\InstQueue_reg[8][2]/NET0131 ,
		_w474_,
		_w477_,
		_w758_
	);
	LUT4 #(
		.INIT('h135f)
	) name306 (
		\InstQueue_reg[0][2]/NET0131 ,
		\InstQueue_reg[13][2]/NET0131 ,
		_w473_,
		_w470_,
		_w759_
	);
	LUT4 #(
		.INIT('h135f)
	) name307 (
		\InstQueue_reg[1][2]/NET0131 ,
		\InstQueue_reg[5][2]/NET0131 ,
		_w463_,
		_w464_,
		_w760_
	);
	LUT4 #(
		.INIT('h153f)
	) name308 (
		\InstQueue_reg[4][2]/NET0131 ,
		\InstQueue_reg[7][2]/NET0131 ,
		_w461_,
		_w476_,
		_w761_
	);
	LUT4 #(
		.INIT('h8000)
	) name309 (
		_w760_,
		_w761_,
		_w758_,
		_w759_,
		_w762_
	);
	LUT2 #(
		.INIT('h8)
	) name310 (
		_w757_,
		_w762_,
		_w763_
	);
	LUT3 #(
		.INIT('h40)
	) name311 (
		_w752_,
		_w757_,
		_w762_,
		_w764_
	);
	LUT2 #(
		.INIT('h1)
	) name312 (
		_w751_,
		_w764_,
		_w765_
	);
	LUT4 #(
		.INIT('h153f)
	) name313 (
		\InstQueue_reg[13][1]/NET0131 ,
		\InstQueue_reg[7][1]/NET0131 ,
		_w461_,
		_w470_,
		_w766_
	);
	LUT4 #(
		.INIT('h135f)
	) name314 (
		\InstQueue_reg[1][1]/NET0131 ,
		\InstQueue_reg[6][1]/NET0131 ,
		_w463_,
		_w467_,
		_w767_
	);
	LUT4 #(
		.INIT('h153f)
	) name315 (
		\InstQueue_reg[12][1]/NET0131 ,
		\InstQueue_reg[14][1]/NET0131 ,
		_w456_,
		_w458_,
		_w768_
	);
	LUT4 #(
		.INIT('h153f)
	) name316 (
		\InstQueue_reg[11][1]/NET0131 ,
		\InstQueue_reg[5][1]/NET0131 ,
		_w464_,
		_w471_,
		_w769_
	);
	LUT4 #(
		.INIT('h8000)
	) name317 (
		_w768_,
		_w769_,
		_w766_,
		_w767_,
		_w770_
	);
	LUT4 #(
		.INIT('h7800)
	) name318 (
		\InstQueueRd_Addr_reg[0]/NET0131 ,
		\InstQueueRd_Addr_reg[1]/NET0131 ,
		\InstQueueRd_Addr_reg[2]/NET0131 ,
		\InstQueueRd_Addr_reg[3]/NET0131 ,
		_w771_
	);
	LUT3 #(
		.INIT('h40)
	) name319 (
		\InstQueueRd_Addr_reg[0]/NET0131 ,
		\InstQueueRd_Addr_reg[1]/NET0131 ,
		\InstQueue_reg[15][1]/NET0131 ,
		_w772_
	);
	LUT2 #(
		.INIT('h8)
	) name320 (
		_w771_,
		_w772_,
		_w773_
	);
	LUT4 #(
		.INIT('h135f)
	) name321 (
		\InstQueue_reg[4][1]/NET0131 ,
		\InstQueue_reg[9][1]/NET0131 ,
		_w476_,
		_w468_,
		_w774_
	);
	LUT4 #(
		.INIT('h135f)
	) name322 (
		\InstQueue_reg[0][1]/NET0131 ,
		\InstQueue_reg[8][1]/NET0131 ,
		_w473_,
		_w477_,
		_w775_
	);
	LUT3 #(
		.INIT('h40)
	) name323 (
		_w773_,
		_w774_,
		_w775_,
		_w776_
	);
	LUT3 #(
		.INIT('h20)
	) name324 (
		\InstQueueRd_Addr_reg[0]/NET0131 ,
		\InstQueueRd_Addr_reg[1]/NET0131 ,
		\InstQueue_reg[10][1]/NET0131 ,
		_w777_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name325 (
		\InstQueueRd_Addr_reg[0]/NET0131 ,
		\InstQueueRd_Addr_reg[1]/NET0131 ,
		\InstQueue_reg[2][1]/NET0131 ,
		\InstQueue_reg[3][1]/NET0131 ,
		_w778_
	);
	LUT4 #(
		.INIT('hefcd)
	) name326 (
		_w648_,
		_w655_,
		_w777_,
		_w778_,
		_w779_
	);
	LUT3 #(
		.INIT('h80)
	) name327 (
		_w770_,
		_w776_,
		_w779_,
		_w780_
	);
	LUT4 #(
		.INIT('h1555)
	) name328 (
		\InstAddrPointer_reg[1]/NET0131 ,
		_w770_,
		_w776_,
		_w779_,
		_w781_
	);
	LUT4 #(
		.INIT('h153f)
	) name329 (
		\InstQueue_reg[10][0]/NET0131 ,
		\InstQueue_reg[2][0]/NET0131 ,
		_w453_,
		_w454_,
		_w782_
	);
	LUT4 #(
		.INIT('h153f)
	) name330 (
		\InstQueue_reg[13][0]/NET0131 ,
		\InstQueue_reg[3][0]/NET0131 ,
		_w474_,
		_w470_,
		_w783_
	);
	LUT4 #(
		.INIT('h135f)
	) name331 (
		\InstQueue_reg[15][0]/NET0131 ,
		\InstQueue_reg[9][0]/NET0131 ,
		_w460_,
		_w468_,
		_w784_
	);
	LUT4 #(
		.INIT('h153f)
	) name332 (
		\InstQueue_reg[5][0]/NET0131 ,
		\InstQueue_reg[7][0]/NET0131 ,
		_w461_,
		_w464_,
		_w785_
	);
	LUT4 #(
		.INIT('h8000)
	) name333 (
		_w784_,
		_w785_,
		_w782_,
		_w783_,
		_w786_
	);
	LUT4 #(
		.INIT('h135f)
	) name334 (
		\InstQueue_reg[1][0]/NET0131 ,
		\InstQueue_reg[8][0]/NET0131 ,
		_w463_,
		_w477_,
		_w787_
	);
	LUT4 #(
		.INIT('h135f)
	) name335 (
		\InstQueue_reg[0][0]/NET0131 ,
		\InstQueue_reg[6][0]/NET0131 ,
		_w473_,
		_w467_,
		_w788_
	);
	LUT4 #(
		.INIT('h153f)
	) name336 (
		\InstQueue_reg[11][0]/NET0131 ,
		\InstQueue_reg[14][0]/NET0131 ,
		_w456_,
		_w471_,
		_w789_
	);
	LUT4 #(
		.INIT('h135f)
	) name337 (
		\InstQueue_reg[12][0]/NET0131 ,
		\InstQueue_reg[4][0]/NET0131 ,
		_w458_,
		_w476_,
		_w790_
	);
	LUT4 #(
		.INIT('h8000)
	) name338 (
		_w789_,
		_w790_,
		_w787_,
		_w788_,
		_w791_
	);
	LUT2 #(
		.INIT('h8)
	) name339 (
		_w786_,
		_w791_,
		_w792_
	);
	LUT3 #(
		.INIT('h2a)
	) name340 (
		\InstAddrPointer_reg[0]/NET0131 ,
		_w786_,
		_w791_,
		_w793_
	);
	LUT3 #(
		.INIT('h8e)
	) name341 (
		\InstAddrPointer_reg[1]/NET0131 ,
		_w780_,
		_w793_,
		_w794_
	);
	LUT4 #(
		.INIT('hbf00)
	) name342 (
		_w739_,
		_w743_,
		_w748_,
		_w750_,
		_w795_
	);
	LUT3 #(
		.INIT('h2a)
	) name343 (
		_w752_,
		_w757_,
		_w762_,
		_w796_
	);
	LUT3 #(
		.INIT('h23)
	) name344 (
		_w751_,
		_w795_,
		_w796_,
		_w797_
	);
	LUT2 #(
		.INIT('h8)
	) name345 (
		\InstAddrPointer_reg[5]/NET0131 ,
		_w725_,
		_w798_
	);
	LUT2 #(
		.INIT('h6)
	) name346 (
		\InstAddrPointer_reg[5]/NET0131 ,
		_w725_,
		_w799_
	);
	LUT4 #(
		.INIT('h135f)
	) name347 (
		\InstQueue_reg[15][5]/NET0131 ,
		\InstQueue_reg[4][5]/NET0131 ,
		_w460_,
		_w476_,
		_w800_
	);
	LUT4 #(
		.INIT('h153f)
	) name348 (
		\InstQueue_reg[11][5]/NET0131 ,
		\InstQueue_reg[13][5]/NET0131 ,
		_w470_,
		_w471_,
		_w801_
	);
	LUT4 #(
		.INIT('h135f)
	) name349 (
		\InstQueue_reg[12][5]/NET0131 ,
		\InstQueue_reg[9][5]/NET0131 ,
		_w458_,
		_w468_,
		_w802_
	);
	LUT4 #(
		.INIT('h153f)
	) name350 (
		\InstQueue_reg[0][5]/NET0131 ,
		\InstQueue_reg[2][5]/NET0131 ,
		_w453_,
		_w473_,
		_w803_
	);
	LUT4 #(
		.INIT('h8000)
	) name351 (
		_w802_,
		_w803_,
		_w800_,
		_w801_,
		_w804_
	);
	LUT4 #(
		.INIT('h135f)
	) name352 (
		\InstQueue_reg[1][5]/NET0131 ,
		\InstQueue_reg[6][5]/NET0131 ,
		_w463_,
		_w467_,
		_w805_
	);
	LUT4 #(
		.INIT('h135f)
	) name353 (
		\InstQueue_reg[10][5]/NET0131 ,
		\InstQueue_reg[14][5]/NET0131 ,
		_w454_,
		_w456_,
		_w806_
	);
	LUT4 #(
		.INIT('h135f)
	) name354 (
		\InstQueue_reg[3][5]/NET0131 ,
		\InstQueue_reg[8][5]/NET0131 ,
		_w474_,
		_w477_,
		_w807_
	);
	LUT4 #(
		.INIT('h153f)
	) name355 (
		\InstQueue_reg[5][5]/NET0131 ,
		\InstQueue_reg[7][5]/NET0131 ,
		_w461_,
		_w464_,
		_w808_
	);
	LUT4 #(
		.INIT('h8000)
	) name356 (
		_w807_,
		_w808_,
		_w805_,
		_w806_,
		_w809_
	);
	LUT2 #(
		.INIT('h8)
	) name357 (
		_w804_,
		_w809_,
		_w810_
	);
	LUT3 #(
		.INIT('h40)
	) name358 (
		_w799_,
		_w804_,
		_w809_,
		_w811_
	);
	LUT4 #(
		.INIT('h7f80)
	) name359 (
		\InstAddrPointer_reg[1]/NET0131 ,
		\InstAddrPointer_reg[2]/NET0131 ,
		\InstAddrPointer_reg[3]/NET0131 ,
		\InstAddrPointer_reg[4]/NET0131 ,
		_w812_
	);
	LUT4 #(
		.INIT('h153f)
	) name360 (
		\InstQueue_reg[11][4]/NET0131 ,
		\InstQueue_reg[1][4]/NET0131 ,
		_w463_,
		_w471_,
		_w813_
	);
	LUT4 #(
		.INIT('h135f)
	) name361 (
		\InstQueue_reg[4][4]/NET0131 ,
		\InstQueue_reg[6][4]/NET0131 ,
		_w476_,
		_w467_,
		_w814_
	);
	LUT4 #(
		.INIT('h153f)
	) name362 (
		\InstQueue_reg[2][4]/NET0131 ,
		\InstQueue_reg[5][4]/NET0131 ,
		_w464_,
		_w453_,
		_w815_
	);
	LUT4 #(
		.INIT('h153f)
	) name363 (
		\InstQueue_reg[10][4]/NET0131 ,
		\InstQueue_reg[15][4]/NET0131 ,
		_w460_,
		_w454_,
		_w816_
	);
	LUT4 #(
		.INIT('h8000)
	) name364 (
		_w815_,
		_w816_,
		_w813_,
		_w814_,
		_w817_
	);
	LUT3 #(
		.INIT('h10)
	) name365 (
		\InstQueueRd_Addr_reg[0]/NET0131 ,
		\InstQueueRd_Addr_reg[1]/NET0131 ,
		\InstQueue_reg[13][4]/NET0131 ,
		_w818_
	);
	LUT2 #(
		.INIT('h8)
	) name366 (
		_w771_,
		_w818_,
		_w819_
	);
	LUT2 #(
		.INIT('h8)
	) name367 (
		\InstQueue_reg[9][4]/NET0131 ,
		_w468_,
		_w820_
	);
	LUT4 #(
		.INIT('h153f)
	) name368 (
		\InstQueue_reg[3][4]/NET0131 ,
		\InstQueue_reg[7][4]/NET0131 ,
		_w461_,
		_w474_,
		_w821_
	);
	LUT4 #(
		.INIT('h135f)
	) name369 (
		\InstQueue_reg[12][4]/NET0131 ,
		\InstQueue_reg[8][4]/NET0131 ,
		_w458_,
		_w477_,
		_w822_
	);
	LUT4 #(
		.INIT('h153f)
	) name370 (
		\InstQueue_reg[0][4]/NET0131 ,
		\InstQueue_reg[14][4]/NET0131 ,
		_w456_,
		_w473_,
		_w823_
	);
	LUT4 #(
		.INIT('h4000)
	) name371 (
		_w820_,
		_w822_,
		_w823_,
		_w821_,
		_w824_
	);
	LUT3 #(
		.INIT('h40)
	) name372 (
		_w819_,
		_w817_,
		_w824_,
		_w825_
	);
	LUT4 #(
		.INIT('h1000)
	) name373 (
		_w812_,
		_w819_,
		_w817_,
		_w824_,
		_w826_
	);
	LUT2 #(
		.INIT('h1)
	) name374 (
		_w811_,
		_w826_,
		_w827_
	);
	LUT4 #(
		.INIT('h2f00)
	) name375 (
		_w765_,
		_w794_,
		_w797_,
		_w827_,
		_w828_
	);
	LUT3 #(
		.INIT('h2a)
	) name376 (
		_w799_,
		_w804_,
		_w809_,
		_w829_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name377 (
		_w812_,
		_w819_,
		_w817_,
		_w824_,
		_w830_
	);
	LUT3 #(
		.INIT('h23)
	) name378 (
		_w811_,
		_w829_,
		_w830_,
		_w831_
	);
	LUT3 #(
		.INIT('h6a)
	) name379 (
		\InstAddrPointer_reg[7]/NET0131 ,
		_w725_,
		_w726_,
		_w832_
	);
	LUT4 #(
		.INIT('hff53)
	) name380 (
		\InstQueue_reg[0][7]/NET0131 ,
		\InstQueue_reg[8][7]/NET0131 ,
		_w648_,
		_w655_,
		_w833_
	);
	LUT2 #(
		.INIT('h2)
	) name381 (
		_w457_,
		_w833_,
		_w834_
	);
	LUT4 #(
		.INIT('h135f)
	) name382 (
		\InstQueue_reg[6][7]/NET0131 ,
		\InstQueue_reg[9][7]/NET0131 ,
		_w467_,
		_w468_,
		_w835_
	);
	LUT4 #(
		.INIT('h153f)
	) name383 (
		\InstQueue_reg[13][7]/NET0131 ,
		\InstQueue_reg[14][7]/NET0131 ,
		_w456_,
		_w470_,
		_w836_
	);
	LUT4 #(
		.INIT('h153f)
	) name384 (
		\InstQueue_reg[10][7]/NET0131 ,
		\InstQueue_reg[15][7]/NET0131 ,
		_w460_,
		_w454_,
		_w837_
	);
	LUT3 #(
		.INIT('h80)
	) name385 (
		_w835_,
		_w836_,
		_w837_,
		_w838_
	);
	LUT4 #(
		.INIT('h153f)
	) name386 (
		\InstQueue_reg[11][7]/NET0131 ,
		\InstQueue_reg[1][7]/NET0131 ,
		_w463_,
		_w471_,
		_w839_
	);
	LUT4 #(
		.INIT('h153f)
	) name387 (
		\InstQueue_reg[3][7]/NET0131 ,
		\InstQueue_reg[5][7]/NET0131 ,
		_w464_,
		_w474_,
		_w840_
	);
	LUT4 #(
		.INIT('h153f)
	) name388 (
		\InstQueue_reg[2][7]/NET0131 ,
		\InstQueue_reg[7][7]/NET0131 ,
		_w461_,
		_w453_,
		_w841_
	);
	LUT4 #(
		.INIT('h135f)
	) name389 (
		\InstQueue_reg[12][7]/NET0131 ,
		\InstQueue_reg[4][7]/NET0131 ,
		_w458_,
		_w476_,
		_w842_
	);
	LUT4 #(
		.INIT('h8000)
	) name390 (
		_w841_,
		_w842_,
		_w839_,
		_w840_,
		_w843_
	);
	LUT3 #(
		.INIT('h40)
	) name391 (
		_w834_,
		_w838_,
		_w843_,
		_w844_
	);
	LUT4 #(
		.INIT('h1000)
	) name392 (
		_w832_,
		_w834_,
		_w838_,
		_w843_,
		_w845_
	);
	LUT3 #(
		.INIT('h6c)
	) name393 (
		\InstAddrPointer_reg[5]/NET0131 ,
		\InstAddrPointer_reg[6]/NET0131 ,
		_w725_,
		_w846_
	);
	LUT4 #(
		.INIT('h135f)
	) name394 (
		\InstQueue_reg[15][6]/NET0131 ,
		\InstQueue_reg[9][6]/NET0131 ,
		_w460_,
		_w468_,
		_w847_
	);
	LUT4 #(
		.INIT('h135f)
	) name395 (
		\InstQueue_reg[10][6]/NET0131 ,
		\InstQueue_reg[13][6]/NET0131 ,
		_w454_,
		_w470_,
		_w848_
	);
	LUT4 #(
		.INIT('h153f)
	) name396 (
		\InstQueue_reg[11][6]/NET0131 ,
		\InstQueue_reg[8][6]/NET0131 ,
		_w477_,
		_w471_,
		_w849_
	);
	LUT4 #(
		.INIT('h135f)
	) name397 (
		\InstQueue_reg[3][6]/NET0131 ,
		\InstQueue_reg[6][6]/NET0131 ,
		_w474_,
		_w467_,
		_w850_
	);
	LUT4 #(
		.INIT('h8000)
	) name398 (
		_w849_,
		_w850_,
		_w847_,
		_w848_,
		_w851_
	);
	LUT4 #(
		.INIT('h153f)
	) name399 (
		\InstQueue_reg[12][6]/NET0131 ,
		\InstQueue_reg[1][6]/NET0131 ,
		_w463_,
		_w458_,
		_w852_
	);
	LUT4 #(
		.INIT('h153f)
	) name400 (
		\InstQueue_reg[0][6]/NET0131 ,
		\InstQueue_reg[5][6]/NET0131 ,
		_w464_,
		_w473_,
		_w853_
	);
	LUT4 #(
		.INIT('h153f)
	) name401 (
		\InstQueue_reg[4][6]/NET0131 ,
		\InstQueue_reg[7][6]/NET0131 ,
		_w461_,
		_w476_,
		_w854_
	);
	LUT4 #(
		.INIT('h153f)
	) name402 (
		\InstQueue_reg[14][6]/NET0131 ,
		\InstQueue_reg[2][6]/NET0131 ,
		_w453_,
		_w456_,
		_w855_
	);
	LUT4 #(
		.INIT('h8000)
	) name403 (
		_w854_,
		_w855_,
		_w852_,
		_w853_,
		_w856_
	);
	LUT2 #(
		.INIT('h8)
	) name404 (
		_w851_,
		_w856_,
		_w857_
	);
	LUT3 #(
		.INIT('h40)
	) name405 (
		_w846_,
		_w851_,
		_w856_,
		_w858_
	);
	LUT2 #(
		.INIT('h1)
	) name406 (
		_w845_,
		_w858_,
		_w859_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name407 (
		_w832_,
		_w834_,
		_w838_,
		_w843_,
		_w860_
	);
	LUT3 #(
		.INIT('h2a)
	) name408 (
		_w846_,
		_w851_,
		_w856_,
		_w861_
	);
	LUT3 #(
		.INIT('h23)
	) name409 (
		_w845_,
		_w860_,
		_w861_,
		_w862_
	);
	LUT4 #(
		.INIT('h4f00)
	) name410 (
		_w828_,
		_w831_,
		_w859_,
		_w862_,
		_w863_
	);
	LUT4 #(
		.INIT('h8000)
	) name411 (
		\InstAddrPointer_reg[10]/NET0131 ,
		\InstAddrPointer_reg[11]/NET0131 ,
		\InstAddrPointer_reg[12]/NET0131 ,
		\InstAddrPointer_reg[9]/NET0131 ,
		_w864_
	);
	LUT3 #(
		.INIT('h80)
	) name412 (
		\InstAddrPointer_reg[13]/NET0131 ,
		_w727_,
		_w864_,
		_w865_
	);
	LUT4 #(
		.INIT('h8000)
	) name413 (
		\InstAddrPointer_reg[13]/NET0131 ,
		\InstAddrPointer_reg[14]/NET0131 ,
		_w727_,
		_w864_,
		_w866_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name414 (
		\InstAddrPointer_reg[13]/NET0131 ,
		\InstAddrPointer_reg[14]/NET0131 ,
		_w727_,
		_w864_,
		_w867_
	);
	LUT3 #(
		.INIT('h80)
	) name415 (
		\InstAddrPointer_reg[13]/NET0131 ,
		\InstAddrPointer_reg[14]/NET0131 ,
		\InstAddrPointer_reg[15]/NET0131 ,
		_w868_
	);
	LUT4 #(
		.INIT('h8000)
	) name416 (
		\InstAddrPointer_reg[10]/NET0131 ,
		\InstAddrPointer_reg[11]/NET0131 ,
		\InstAddrPointer_reg[12]/NET0131 ,
		\InstAddrPointer_reg[16]/NET0131 ,
		_w869_
	);
	LUT2 #(
		.INIT('h8)
	) name417 (
		_w868_,
		_w869_,
		_w870_
	);
	LUT3 #(
		.INIT('h80)
	) name418 (
		\InstAddrPointer_reg[9]/NET0131 ,
		_w868_,
		_w869_,
		_w871_
	);
	LUT2 #(
		.INIT('h8)
	) name419 (
		_w727_,
		_w871_,
		_w872_
	);
	LUT2 #(
		.INIT('h8)
	) name420 (
		\InstAddrPointer_reg[18]/NET0131 ,
		\InstAddrPointer_reg[19]/NET0131 ,
		_w873_
	);
	LUT3 #(
		.INIT('h80)
	) name421 (
		\InstAddrPointer_reg[17]/NET0131 ,
		\InstAddrPointer_reg[18]/NET0131 ,
		\InstAddrPointer_reg[19]/NET0131 ,
		_w874_
	);
	LUT3 #(
		.INIT('h80)
	) name422 (
		_w727_,
		_w871_,
		_w874_,
		_w875_
	);
	LUT2 #(
		.INIT('h8)
	) name423 (
		\InstAddrPointer_reg[20]/NET0131 ,
		\InstAddrPointer_reg[21]/NET0131 ,
		_w876_
	);
	LUT3 #(
		.INIT('h80)
	) name424 (
		\InstAddrPointer_reg[20]/NET0131 ,
		\InstAddrPointer_reg[21]/NET0131 ,
		\InstAddrPointer_reg[22]/NET0131 ,
		_w877_
	);
	LUT4 #(
		.INIT('h8000)
	) name425 (
		\InstAddrPointer_reg[20]/NET0131 ,
		\InstAddrPointer_reg[21]/NET0131 ,
		\InstAddrPointer_reg[22]/NET0131 ,
		\InstAddrPointer_reg[23]/NET0131 ,
		_w878_
	);
	LUT2 #(
		.INIT('h8)
	) name426 (
		\InstAddrPointer_reg[24]/NET0131 ,
		_w878_,
		_w879_
	);
	LUT4 #(
		.INIT('h8000)
	) name427 (
		_w727_,
		_w871_,
		_w874_,
		_w879_,
		_w880_
	);
	LUT3 #(
		.INIT('h80)
	) name428 (
		\InstAddrPointer_reg[25]/NET0131 ,
		\InstAddrPointer_reg[26]/NET0131 ,
		_w880_,
		_w881_
	);
	LUT3 #(
		.INIT('h6c)
	) name429 (
		\InstAddrPointer_reg[25]/NET0131 ,
		\InstAddrPointer_reg[26]/NET0131 ,
		_w880_,
		_w882_
	);
	LUT2 #(
		.INIT('h6)
	) name430 (
		\InstAddrPointer_reg[25]/NET0131 ,
		_w880_,
		_w883_
	);
	LUT3 #(
		.INIT('h48)
	) name431 (
		\InstAddrPointer_reg[25]/NET0131 ,
		\InstAddrPointer_reg[26]/NET0131 ,
		_w880_,
		_w884_
	);
	LUT4 #(
		.INIT('h8000)
	) name432 (
		_w727_,
		_w877_,
		_w871_,
		_w874_,
		_w885_
	);
	LUT4 #(
		.INIT('h00ec)
	) name433 (
		\InstAddrPointer_reg[23]/NET0131 ,
		\InstAddrPointer_reg[24]/NET0131 ,
		_w885_,
		_w880_,
		_w886_
	);
	LUT2 #(
		.INIT('h6)
	) name434 (
		\InstAddrPointer_reg[23]/NET0131 ,
		_w885_,
		_w887_
	);
	LUT3 #(
		.INIT('h80)
	) name435 (
		_w884_,
		_w886_,
		_w887_,
		_w888_
	);
	LUT3 #(
		.INIT('h80)
	) name436 (
		\InstAddrPointer_reg[24]/NET0131 ,
		\InstAddrPointer_reg[25]/NET0131 ,
		\InstAddrPointer_reg[26]/NET0131 ,
		_w889_
	);
	LUT4 #(
		.INIT('h8000)
	) name437 (
		\InstAddrPointer_reg[23]/NET0131 ,
		\InstAddrPointer_reg[27]/NET0131 ,
		_w889_,
		_w885_,
		_w890_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name438 (
		\InstAddrPointer_reg[23]/NET0131 ,
		\InstAddrPointer_reg[27]/NET0131 ,
		_w889_,
		_w885_,
		_w891_
	);
	LUT2 #(
		.INIT('h8)
	) name439 (
		\InstAddrPointer_reg[28]/NET0131 ,
		_w891_,
		_w892_
	);
	LUT2 #(
		.INIT('h8)
	) name440 (
		\InstAddrPointer_reg[27]/NET0131 ,
		\InstAddrPointer_reg[28]/NET0131 ,
		_w893_
	);
	LUT4 #(
		.INIT('h8000)
	) name441 (
		\InstAddrPointer_reg[25]/NET0131 ,
		\InstAddrPointer_reg[26]/NET0131 ,
		_w880_,
		_w893_,
		_w894_
	);
	LUT3 #(
		.INIT('h80)
	) name442 (
		\InstAddrPointer_reg[27]/NET0131 ,
		\InstAddrPointer_reg[28]/NET0131 ,
		\InstAddrPointer_reg[29]/NET0131 ,
		_w895_
	);
	LUT4 #(
		.INIT('h8000)
	) name443 (
		\InstAddrPointer_reg[25]/NET0131 ,
		\InstAddrPointer_reg[26]/NET0131 ,
		_w880_,
		_w895_,
		_w896_
	);
	LUT3 #(
		.INIT('h6a)
	) name444 (
		\InstAddrPointer_reg[29]/NET0131 ,
		_w881_,
		_w893_,
		_w897_
	);
	LUT3 #(
		.INIT('h80)
	) name445 (
		_w892_,
		_w888_,
		_w897_,
		_w898_
	);
	LUT4 #(
		.INIT('h8000)
	) name446 (
		\InstAddrPointer_reg[30]/NET0131 ,
		_w892_,
		_w888_,
		_w897_,
		_w899_
	);
	LUT2 #(
		.INIT('h1)
	) name447 (
		\InstAddrPointer_reg[15]/NET0131 ,
		_w866_,
		_w900_
	);
	LUT2 #(
		.INIT('h8)
	) name448 (
		\InstAddrPointer_reg[15]/NET0131 ,
		_w866_,
		_w901_
	);
	LUT2 #(
		.INIT('h6)
	) name449 (
		\InstAddrPointer_reg[15]/NET0131 ,
		_w866_,
		_w902_
	);
	LUT3 #(
		.INIT('h20)
	) name450 (
		\InstAddrPointer_reg[15]/NET0131 ,
		\InstAddrPointer_reg[16]/NET0131 ,
		_w866_,
		_w903_
	);
	LUT3 #(
		.INIT('h93)
	) name451 (
		\InstAddrPointer_reg[15]/NET0131 ,
		\InstAddrPointer_reg[16]/NET0131 ,
		_w866_,
		_w904_
	);
	LUT3 #(
		.INIT('h80)
	) name452 (
		\InstAddrPointer_reg[17]/NET0131 ,
		_w727_,
		_w871_,
		_w905_
	);
	LUT3 #(
		.INIT('h6a)
	) name453 (
		\InstAddrPointer_reg[17]/NET0131 ,
		_w727_,
		_w871_,
		_w906_
	);
	LUT4 #(
		.INIT('h6c00)
	) name454 (
		\InstAddrPointer_reg[15]/NET0131 ,
		\InstAddrPointer_reg[16]/NET0131 ,
		_w866_,
		_w906_,
		_w907_
	);
	LUT4 #(
		.INIT('h8000)
	) name455 (
		\InstAddrPointer_reg[17]/NET0131 ,
		\InstAddrPointer_reg[18]/NET0131 ,
		_w727_,
		_w871_,
		_w908_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name456 (
		\InstAddrPointer_reg[17]/NET0131 ,
		\InstAddrPointer_reg[18]/NET0131 ,
		_w727_,
		_w871_,
		_w909_
	);
	LUT2 #(
		.INIT('h8)
	) name457 (
		\InstAddrPointer_reg[19]/NET0131 ,
		_w909_,
		_w910_
	);
	LUT4 #(
		.INIT('h8000)
	) name458 (
		_w727_,
		_w876_,
		_w871_,
		_w874_,
		_w911_
	);
	LUT3 #(
		.INIT('h32)
	) name459 (
		\InstAddrPointer_reg[22]/NET0131 ,
		_w885_,
		_w911_,
		_w912_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name460 (
		\InstAddrPointer_reg[20]/NET0131 ,
		_w727_,
		_w871_,
		_w874_,
		_w913_
	);
	LUT2 #(
		.INIT('h8)
	) name461 (
		\InstAddrPointer_reg[21]/NET0131 ,
		_w913_,
		_w914_
	);
	LUT4 #(
		.INIT('h4080)
	) name462 (
		\InstAddrPointer_reg[20]/NET0131 ,
		\InstAddrPointer_reg[21]/NET0131 ,
		\InstAddrPointer_reg[22]/NET0131 ,
		_w875_,
		_w915_
	);
	LUT3 #(
		.INIT('h80)
	) name463 (
		_w907_,
		_w910_,
		_w915_,
		_w916_
	);
	LUT4 #(
		.INIT('h8000)
	) name464 (
		_w902_,
		_w907_,
		_w910_,
		_w915_,
		_w917_
	);
	LUT2 #(
		.INIT('h8)
	) name465 (
		_w899_,
		_w917_,
		_w918_
	);
	LUT4 #(
		.INIT('h2000)
	) name466 (
		_w736_,
		_w863_,
		_w867_,
		_w918_,
		_w919_
	);
	LUT4 #(
		.INIT('h8000)
	) name467 (
		\InstAddrPointer_reg[27]/NET0131 ,
		\InstAddrPointer_reg[28]/NET0131 ,
		\InstAddrPointer_reg[29]/NET0131 ,
		\InstAddrPointer_reg[30]/NET0131 ,
		_w920_
	);
	LUT4 #(
		.INIT('h8000)
	) name468 (
		\InstAddrPointer_reg[23]/NET0131 ,
		_w889_,
		_w885_,
		_w920_,
		_w921_
	);
	LUT2 #(
		.INIT('h9)
	) name469 (
		\InstAddrPointer_reg[31]/NET0131 ,
		_w921_,
		_w922_
	);
	LUT4 #(
		.INIT('h008e)
	) name470 (
		\InstAddrPointer_reg[1]/NET0131 ,
		_w780_,
		_w793_,
		_w796_,
		_w923_
	);
	LUT3 #(
		.INIT('h01)
	) name471 (
		_w826_,
		_w751_,
		_w764_,
		_w924_
	);
	LUT3 #(
		.INIT('h0b)
	) name472 (
		_w826_,
		_w795_,
		_w830_,
		_w925_
	);
	LUT2 #(
		.INIT('h1)
	) name473 (
		_w858_,
		_w811_,
		_w926_
	);
	LUT4 #(
		.INIT('h4f00)
	) name474 (
		_w923_,
		_w924_,
		_w925_,
		_w926_,
		_w927_
	);
	LUT3 #(
		.INIT('h0b)
	) name475 (
		_w858_,
		_w829_,
		_w861_,
		_w928_
	);
	LUT4 #(
		.INIT('h004d)
	) name476 (
		_w846_,
		_w857_,
		_w829_,
		_w860_,
		_w929_
	);
	LUT2 #(
		.INIT('h2)
	) name477 (
		_w733_,
		_w845_,
		_w930_
	);
	LUT2 #(
		.INIT('h6)
	) name478 (
		\InstAddrPointer_reg[9]/NET0131 ,
		_w727_,
		_w931_
	);
	LUT3 #(
		.INIT('h28)
	) name479 (
		\InstAddrPointer_reg[10]/NET0131 ,
		\InstAddrPointer_reg[9]/NET0131 ,
		_w727_,
		_w932_
	);
	LUT4 #(
		.INIT('hb000)
	) name480 (
		_w927_,
		_w929_,
		_w930_,
		_w932_,
		_w933_
	);
	LUT2 #(
		.INIT('h8)
	) name481 (
		\InstAddrPointer_reg[15]/NET0131 ,
		_w867_,
		_w934_
	);
	LUT2 #(
		.INIT('h8)
	) name482 (
		_w732_,
		_w934_,
		_w935_
	);
	LUT2 #(
		.INIT('h8)
	) name483 (
		_w916_,
		_w935_,
		_w936_
	);
	LUT2 #(
		.INIT('h2)
	) name484 (
		_w899_,
		_w922_,
		_w937_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name485 (
		_w844_,
		_w933_,
		_w936_,
		_w937_,
		_w938_
	);
	LUT3 #(
		.INIT('hb0)
	) name486 (
		_w919_,
		_w922_,
		_w938_,
		_w939_
	);
	LUT2 #(
		.INIT('h8)
	) name487 (
		\InstAddrPointer_reg[0]/NET0131 ,
		\InstAddrPointer_reg[1]/NET0131 ,
		_w940_
	);
	LUT4 #(
		.INIT('h8000)
	) name488 (
		\InstAddrPointer_reg[0]/NET0131 ,
		\InstAddrPointer_reg[1]/NET0131 ,
		\InstAddrPointer_reg[2]/NET0131 ,
		\InstAddrPointer_reg[3]/NET0131 ,
		_w941_
	);
	LUT4 #(
		.INIT('h8000)
	) name489 (
		\InstAddrPointer_reg[4]/NET0131 ,
		\InstAddrPointer_reg[7]/NET0131 ,
		_w726_,
		_w941_,
		_w942_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name490 (
		\InstAddrPointer_reg[4]/NET0131 ,
		\InstAddrPointer_reg[7]/NET0131 ,
		_w726_,
		_w941_,
		_w943_
	);
	LUT4 #(
		.INIT('h0040)
	) name491 (
		_w834_,
		_w838_,
		_w843_,
		_w943_,
		_w944_
	);
	LUT4 #(
		.INIT('h78f0)
	) name492 (
		\InstAddrPointer_reg[4]/NET0131 ,
		\InstAddrPointer_reg[5]/NET0131 ,
		\InstAddrPointer_reg[6]/NET0131 ,
		_w941_,
		_w945_
	);
	LUT3 #(
		.INIT('h08)
	) name493 (
		_w851_,
		_w856_,
		_w945_,
		_w946_
	);
	LUT3 #(
		.INIT('h6c)
	) name494 (
		\InstAddrPointer_reg[4]/NET0131 ,
		\InstAddrPointer_reg[5]/NET0131 ,
		_w941_,
		_w947_
	);
	LUT3 #(
		.INIT('h08)
	) name495 (
		_w804_,
		_w809_,
		_w947_,
		_w948_
	);
	LUT2 #(
		.INIT('h1)
	) name496 (
		_w946_,
		_w948_,
		_w949_
	);
	LUT3 #(
		.INIT('h78)
	) name497 (
		\InstAddrPointer_reg[0]/NET0131 ,
		\InstAddrPointer_reg[1]/NET0131 ,
		\InstAddrPointer_reg[2]/NET0131 ,
		_w950_
	);
	LUT3 #(
		.INIT('h70)
	) name498 (
		_w757_,
		_w762_,
		_w950_,
		_w951_
	);
	LUT3 #(
		.INIT('h80)
	) name499 (
		\InstAddrPointer_reg[0]/NET0131 ,
		_w786_,
		_w791_,
		_w952_
	);
	LUT3 #(
		.INIT('h08)
	) name500 (
		_w757_,
		_w762_,
		_w950_,
		_w953_
	);
	LUT2 #(
		.INIT('h6)
	) name501 (
		\InstAddrPointer_reg[0]/NET0131 ,
		\InstAddrPointer_reg[1]/NET0131 ,
		_w954_
	);
	LUT4 #(
		.INIT('h0080)
	) name502 (
		_w770_,
		_w776_,
		_w779_,
		_w954_,
		_w955_
	);
	LUT4 #(
		.INIT('h000b)
	) name503 (
		_w781_,
		_w952_,
		_w953_,
		_w955_,
		_w956_
	);
	LUT2 #(
		.INIT('h6)
	) name504 (
		\InstAddrPointer_reg[4]/NET0131 ,
		_w941_,
		_w957_
	);
	LUT4 #(
		.INIT('h0040)
	) name505 (
		_w819_,
		_w817_,
		_w824_,
		_w957_,
		_w958_
	);
	LUT4 #(
		.INIT('h7f80)
	) name506 (
		\InstAddrPointer_reg[0]/NET0131 ,
		\InstAddrPointer_reg[1]/NET0131 ,
		\InstAddrPointer_reg[2]/NET0131 ,
		\InstAddrPointer_reg[3]/NET0131 ,
		_w959_
	);
	LUT4 #(
		.INIT('h0040)
	) name507 (
		_w739_,
		_w743_,
		_w748_,
		_w959_,
		_w960_
	);
	LUT2 #(
		.INIT('h1)
	) name508 (
		_w958_,
		_w960_,
		_w961_
	);
	LUT4 #(
		.INIT('ha800)
	) name509 (
		_w949_,
		_w951_,
		_w956_,
		_w961_,
		_w962_
	);
	LUT4 #(
		.INIT('hbf00)
	) name510 (
		_w819_,
		_w817_,
		_w824_,
		_w957_,
		_w963_
	);
	LUT4 #(
		.INIT('hbf00)
	) name511 (
		_w739_,
		_w743_,
		_w748_,
		_w959_,
		_w964_
	);
	LUT3 #(
		.INIT('h23)
	) name512 (
		_w958_,
		_w963_,
		_w964_,
		_w965_
	);
	LUT3 #(
		.INIT('h70)
	) name513 (
		_w851_,
		_w856_,
		_w945_,
		_w966_
	);
	LUT3 #(
		.INIT('h70)
	) name514 (
		_w804_,
		_w809_,
		_w947_,
		_w967_
	);
	LUT3 #(
		.INIT('h23)
	) name515 (
		_w946_,
		_w966_,
		_w967_,
		_w968_
	);
	LUT3 #(
		.INIT('hd0)
	) name516 (
		_w949_,
		_w965_,
		_w968_,
		_w969_
	);
	LUT3 #(
		.INIT('h80)
	) name517 (
		\InstAddrPointer_reg[0]/NET0131 ,
		\InstAddrPointer_reg[9]/NET0131 ,
		_w727_,
		_w970_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name518 (
		\InstAddrPointer_reg[0]/NET0131 ,
		\InstAddrPointer_reg[10]/NET0131 ,
		\InstAddrPointer_reg[9]/NET0131 ,
		_w727_,
		_w971_
	);
	LUT3 #(
		.INIT('h13)
	) name519 (
		\InstAddrPointer_reg[8]/NET0131 ,
		\InstAddrPointer_reg[9]/NET0131 ,
		_w942_,
		_w972_
	);
	LUT2 #(
		.INIT('h1)
	) name520 (
		_w970_,
		_w972_,
		_w973_
	);
	LUT3 #(
		.INIT('h98)
	) name521 (
		\InstAddrPointer_reg[10]/NET0131 ,
		_w970_,
		_w972_,
		_w974_
	);
	LUT4 #(
		.INIT('hbf00)
	) name522 (
		_w834_,
		_w838_,
		_w843_,
		_w943_,
		_w975_
	);
	LUT2 #(
		.INIT('h6)
	) name523 (
		\InstAddrPointer_reg[8]/NET0131 ,
		_w942_,
		_w976_
	);
	LUT2 #(
		.INIT('h1)
	) name524 (
		_w975_,
		_w976_,
		_w977_
	);
	LUT3 #(
		.INIT('h02)
	) name525 (
		_w974_,
		_w975_,
		_w976_,
		_w978_
	);
	LUT4 #(
		.INIT('hba00)
	) name526 (
		_w944_,
		_w962_,
		_w969_,
		_w978_,
		_w979_
	);
	LUT4 #(
		.INIT('h8000)
	) name527 (
		\InstAddrPointer_reg[0]/NET0131 ,
		\InstAddrPointer_reg[9]/NET0131 ,
		_w727_,
		_w729_,
		_w980_
	);
	LUT3 #(
		.INIT('h80)
	) name528 (
		\InstAddrPointer_reg[8]/NET0131 ,
		_w864_,
		_w942_,
		_w981_
	);
	LUT3 #(
		.INIT('h0e)
	) name529 (
		\InstAddrPointer_reg[12]/NET0131 ,
		_w980_,
		_w981_,
		_w982_
	);
	LUT3 #(
		.INIT('h6c)
	) name530 (
		\InstAddrPointer_reg[10]/NET0131 ,
		\InstAddrPointer_reg[11]/NET0131 ,
		_w970_,
		_w983_
	);
	LUT4 #(
		.INIT('h8000)
	) name531 (
		\InstAddrPointer_reg[13]/NET0131 ,
		\InstAddrPointer_reg[8]/NET0131 ,
		_w864_,
		_w942_,
		_w984_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name532 (
		\InstAddrPointer_reg[13]/NET0131 ,
		\InstAddrPointer_reg[8]/NET0131 ,
		_w864_,
		_w942_,
		_w985_
	);
	LUT4 #(
		.INIT('h7f4c)
	) name533 (
		\InstAddrPointer_reg[0]/NET0131 ,
		\InstAddrPointer_reg[14]/NET0131 ,
		_w865_,
		_w984_,
		_w986_
	);
	LUT4 #(
		.INIT('h0001)
	) name534 (
		_w982_,
		_w983_,
		_w985_,
		_w986_,
		_w987_
	);
	LUT3 #(
		.INIT('h6c)
	) name535 (
		\InstAddrPointer_reg[0]/NET0131 ,
		\InstAddrPointer_reg[15]/NET0131 ,
		_w866_,
		_w988_
	);
	LUT4 #(
		.INIT('h070f)
	) name536 (
		\InstAddrPointer_reg[0]/NET0131 ,
		\InstAddrPointer_reg[15]/NET0131 ,
		\InstAddrPointer_reg[16]/NET0131 ,
		_w866_,
		_w989_
	);
	LUT3 #(
		.INIT('h80)
	) name537 (
		\InstAddrPointer_reg[0]/NET0131 ,
		_w727_,
		_w871_,
		_w990_
	);
	LUT2 #(
		.INIT('h1)
	) name538 (
		_w989_,
		_w990_,
		_w991_
	);
	LUT3 #(
		.INIT('h6c)
	) name539 (
		\InstAddrPointer_reg[0]/NET0131 ,
		\InstAddrPointer_reg[18]/NET0131 ,
		_w905_,
		_w992_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name540 (
		\InstAddrPointer_reg[0]/NET0131 ,
		\InstAddrPointer_reg[17]/NET0131 ,
		_w727_,
		_w871_,
		_w993_
	);
	LUT4 #(
		.INIT('h8103)
	) name541 (
		\InstAddrPointer_reg[0]/NET0131 ,
		\InstAddrPointer_reg[17]/NET0131 ,
		\InstAddrPointer_reg[18]/NET0131 ,
		_w872_,
		_w994_
	);
	LUT3 #(
		.INIT('he0)
	) name542 (
		_w989_,
		_w990_,
		_w994_,
		_w995_
	);
	LUT3 #(
		.INIT('h20)
	) name543 (
		_w987_,
		_w988_,
		_w995_,
		_w996_
	);
	LUT4 #(
		.INIT('h8000)
	) name544 (
		\InstAddrPointer_reg[0]/NET0131 ,
		_w727_,
		_w871_,
		_w874_,
		_w997_
	);
	LUT4 #(
		.INIT('h00ec)
	) name545 (
		\InstAddrPointer_reg[0]/NET0131 ,
		\InstAddrPointer_reg[19]/NET0131 ,
		_w908_,
		_w997_,
		_w998_
	);
	LUT2 #(
		.INIT('h8)
	) name546 (
		_w879_,
		_w997_,
		_w999_
	);
	LUT4 #(
		.INIT('h070f)
	) name547 (
		\InstAddrPointer_reg[0]/NET0131 ,
		\InstAddrPointer_reg[23]/NET0131 ,
		\InstAddrPointer_reg[24]/NET0131 ,
		_w885_,
		_w1000_
	);
	LUT2 #(
		.INIT('h1)
	) name548 (
		_w999_,
		_w1000_,
		_w1001_
	);
	LUT3 #(
		.INIT('h6c)
	) name549 (
		\InstAddrPointer_reg[0]/NET0131 ,
		\InstAddrPointer_reg[23]/NET0131 ,
		_w885_,
		_w1002_
	);
	LUT2 #(
		.INIT('h8)
	) name550 (
		\InstAddrPointer_reg[0]/NET0131 ,
		_w911_,
		_w1003_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name551 (
		\InstAddrPointer_reg[0]/NET0131 ,
		\InstAddrPointer_reg[22]/NET0131 ,
		_w876_,
		_w875_,
		_w1004_
	);
	LUT4 #(
		.INIT('h0302)
	) name552 (
		_w999_,
		_w1002_,
		_w1004_,
		_w1000_,
		_w1005_
	);
	LUT3 #(
		.INIT('h13)
	) name553 (
		\InstAddrPointer_reg[20]/NET0131 ,
		\InstAddrPointer_reg[21]/NET0131 ,
		_w997_,
		_w1006_
	);
	LUT2 #(
		.INIT('h1)
	) name554 (
		_w1006_,
		_w1003_,
		_w1007_
	);
	LUT2 #(
		.INIT('h6)
	) name555 (
		\InstAddrPointer_reg[20]/NET0131 ,
		_w997_,
		_w1008_
	);
	LUT3 #(
		.INIT('h6a)
	) name556 (
		\InstAddrPointer_reg[25]/NET0131 ,
		_w879_,
		_w997_,
		_w1009_
	);
	LUT4 #(
		.INIT('h9333)
	) name557 (
		\InstAddrPointer_reg[25]/NET0131 ,
		\InstAddrPointer_reg[26]/NET0131 ,
		_w879_,
		_w997_,
		_w1010_
	);
	LUT4 #(
		.INIT('h8111)
	) name558 (
		\InstAddrPointer_reg[25]/NET0131 ,
		\InstAddrPointer_reg[26]/NET0131 ,
		_w879_,
		_w997_,
		_w1011_
	);
	LUT4 #(
		.INIT('h0e00)
	) name559 (
		_w1006_,
		_w1003_,
		_w1008_,
		_w1011_,
		_w1012_
	);
	LUT3 #(
		.INIT('h40)
	) name560 (
		_w998_,
		_w1005_,
		_w1012_,
		_w1013_
	);
	LUT4 #(
		.INIT('h870f)
	) name561 (
		\InstAddrPointer_reg[0]/NET0131 ,
		\InstAddrPointer_reg[29]/NET0131 ,
		\InstAddrPointer_reg[30]/NET0131 ,
		_w894_,
		_w1014_
	);
	LUT4 #(
		.INIT('h8000)
	) name562 (
		\InstAddrPointer_reg[0]/NET0131 ,
		\InstAddrPointer_reg[23]/NET0131 ,
		_w889_,
		_w885_,
		_w1015_
	);
	LUT2 #(
		.INIT('h6)
	) name563 (
		\InstAddrPointer_reg[27]/NET0131 ,
		_w1015_,
		_w1016_
	);
	LUT3 #(
		.INIT('h6c)
	) name564 (
		\InstAddrPointer_reg[27]/NET0131 ,
		\InstAddrPointer_reg[28]/NET0131 ,
		_w1015_,
		_w1017_
	);
	LUT3 #(
		.INIT('h81)
	) name565 (
		\InstAddrPointer_reg[27]/NET0131 ,
		\InstAddrPointer_reg[28]/NET0131 ,
		_w1015_,
		_w1018_
	);
	LUT3 #(
		.INIT('h93)
	) name566 (
		\InstAddrPointer_reg[0]/NET0131 ,
		\InstAddrPointer_reg[29]/NET0131 ,
		_w894_,
		_w1019_
	);
	LUT3 #(
		.INIT('h80)
	) name567 (
		_w1014_,
		_w1018_,
		_w1019_,
		_w1020_
	);
	LUT4 #(
		.INIT('h8000)
	) name568 (
		_w979_,
		_w996_,
		_w1013_,
		_w1020_,
		_w1021_
	);
	LUT3 #(
		.INIT('h93)
	) name569 (
		\InstAddrPointer_reg[0]/NET0131 ,
		\InstAddrPointer_reg[31]/NET0131 ,
		_w921_,
		_w1022_
	);
	LUT3 #(
		.INIT('hbe)
	) name570 (
		_w844_,
		_w1021_,
		_w1022_,
		_w1023_
	);
	LUT4 #(
		.INIT('h1d11)
	) name571 (
		\InstAddrPointer_reg[31]/NET0131 ,
		_w681_,
		_w939_,
		_w1023_,
		_w1024_
	);
	LUT4 #(
		.INIT('hf800)
	) name572 (
		\InstAddrPointer_reg[0]/NET0131 ,
		\InstAddrPointer_reg[1]/NET0131 ,
		\InstAddrPointer_reg[2]/NET0131 ,
		\InstAddrPointer_reg[3]/NET0131 ,
		_w1025_
	);
	LUT2 #(
		.INIT('h6)
	) name573 (
		\InstAddrPointer_reg[4]/NET0131 ,
		_w1025_,
		_w1026_
	);
	LUT4 #(
		.INIT('h0040)
	) name574 (
		_w819_,
		_w817_,
		_w824_,
		_w1026_,
		_w1027_
	);
	LUT4 #(
		.INIT('h07f8)
	) name575 (
		\InstAddrPointer_reg[0]/NET0131 ,
		\InstAddrPointer_reg[1]/NET0131 ,
		\InstAddrPointer_reg[2]/NET0131 ,
		\InstAddrPointer_reg[3]/NET0131 ,
		_w1028_
	);
	LUT4 #(
		.INIT('h0040)
	) name576 (
		_w739_,
		_w743_,
		_w748_,
		_w1028_,
		_w1029_
	);
	LUT2 #(
		.INIT('h1)
	) name577 (
		_w1027_,
		_w1029_,
		_w1030_
	);
	LUT3 #(
		.INIT('h80)
	) name578 (
		_w757_,
		_w762_,
		_w950_,
		_w1031_
	);
	LUT3 #(
		.INIT('h07)
	) name579 (
		_w757_,
		_w762_,
		_w950_,
		_w1032_
	);
	LUT3 #(
		.INIT('h15)
	) name580 (
		\InstAddrPointer_reg[0]/NET0131 ,
		_w786_,
		_w791_,
		_w1033_
	);
	LUT4 #(
		.INIT('h020b)
	) name581 (
		_w780_,
		_w954_,
		_w1032_,
		_w1033_,
		_w1034_
	);
	LUT4 #(
		.INIT('hbf00)
	) name582 (
		_w819_,
		_w817_,
		_w824_,
		_w1026_,
		_w1035_
	);
	LUT4 #(
		.INIT('hbf00)
	) name583 (
		_w739_,
		_w743_,
		_w748_,
		_w1028_,
		_w1036_
	);
	LUT3 #(
		.INIT('h23)
	) name584 (
		_w1027_,
		_w1035_,
		_w1036_,
		_w1037_
	);
	LUT4 #(
		.INIT('hfd00)
	) name585 (
		_w1030_,
		_w1031_,
		_w1034_,
		_w1037_,
		_w1038_
	);
	LUT3 #(
		.INIT('h6c)
	) name586 (
		\InstAddrPointer_reg[4]/NET0131 ,
		\InstAddrPointer_reg[5]/NET0131 ,
		_w1025_,
		_w1039_
	);
	LUT3 #(
		.INIT('h08)
	) name587 (
		_w804_,
		_w809_,
		_w1039_,
		_w1040_
	);
	LUT4 #(
		.INIT('h78f0)
	) name588 (
		\InstAddrPointer_reg[4]/NET0131 ,
		\InstAddrPointer_reg[5]/NET0131 ,
		\InstAddrPointer_reg[6]/NET0131 ,
		_w1025_,
		_w1041_
	);
	LUT3 #(
		.INIT('h08)
	) name589 (
		_w851_,
		_w856_,
		_w1041_,
		_w1042_
	);
	LUT2 #(
		.INIT('h1)
	) name590 (
		_w1040_,
		_w1042_,
		_w1043_
	);
	LUT4 #(
		.INIT('h8000)
	) name591 (
		\InstAddrPointer_reg[4]/NET0131 ,
		\InstAddrPointer_reg[7]/NET0131 ,
		_w726_,
		_w1025_,
		_w1044_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name592 (
		\InstAddrPointer_reg[4]/NET0131 ,
		\InstAddrPointer_reg[7]/NET0131 ,
		_w726_,
		_w1025_,
		_w1045_
	);
	LUT4 #(
		.INIT('hbf00)
	) name593 (
		_w834_,
		_w838_,
		_w843_,
		_w1045_,
		_w1046_
	);
	LUT3 #(
		.INIT('h70)
	) name594 (
		_w851_,
		_w856_,
		_w1041_,
		_w1047_
	);
	LUT3 #(
		.INIT('h70)
	) name595 (
		_w804_,
		_w809_,
		_w1039_,
		_w1048_
	);
	LUT3 #(
		.INIT('h23)
	) name596 (
		_w1042_,
		_w1047_,
		_w1048_,
		_w1049_
	);
	LUT4 #(
		.INIT('h020b)
	) name597 (
		_w857_,
		_w1041_,
		_w1046_,
		_w1048_,
		_w1050_
	);
	LUT4 #(
		.INIT('h0040)
	) name598 (
		_w834_,
		_w838_,
		_w843_,
		_w1045_,
		_w1051_
	);
	LUT2 #(
		.INIT('h6)
	) name599 (
		\InstAddrPointer_reg[8]/NET0131 ,
		_w1044_,
		_w1052_
	);
	LUT2 #(
		.INIT('h4)
	) name600 (
		_w1051_,
		_w1052_,
		_w1053_
	);
	LUT4 #(
		.INIT('h4f00)
	) name601 (
		_w1038_,
		_w1043_,
		_w1050_,
		_w1053_,
		_w1054_
	);
	LUT3 #(
		.INIT('h80)
	) name602 (
		\InstAddrPointer_reg[8]/NET0131 ,
		_w864_,
		_w1044_,
		_w1055_
	);
	LUT4 #(
		.INIT('h8000)
	) name603 (
		\InstAddrPointer_reg[13]/NET0131 ,
		\InstAddrPointer_reg[8]/NET0131 ,
		_w864_,
		_w1044_,
		_w1056_
	);
	LUT3 #(
		.INIT('h6c)
	) name604 (
		\InstAddrPointer_reg[14]/NET0131 ,
		\InstAddrPointer_reg[15]/NET0131 ,
		_w1056_,
		_w1057_
	);
	LUT4 #(
		.INIT('h60c0)
	) name605 (
		\InstAddrPointer_reg[14]/NET0131 ,
		\InstAddrPointer_reg[15]/NET0131 ,
		\InstAddrPointer_reg[16]/NET0131 ,
		_w1056_,
		_w1058_
	);
	LUT4 #(
		.INIT('h8000)
	) name606 (
		\InstAddrPointer_reg[10]/NET0131 ,
		\InstAddrPointer_reg[8]/NET0131 ,
		\InstAddrPointer_reg[9]/NET0131 ,
		_w1044_,
		_w1059_
	);
	LUT2 #(
		.INIT('h6)
	) name607 (
		\InstAddrPointer_reg[11]/NET0131 ,
		_w1059_,
		_w1060_
	);
	LUT3 #(
		.INIT('h48)
	) name608 (
		\InstAddrPointer_reg[11]/NET0131 ,
		\InstAddrPointer_reg[12]/NET0131 ,
		_w1059_,
		_w1061_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name609 (
		\InstAddrPointer_reg[13]/NET0131 ,
		\InstAddrPointer_reg[8]/NET0131 ,
		_w864_,
		_w1044_,
		_w1062_
	);
	LUT2 #(
		.INIT('h8)
	) name610 (
		\InstAddrPointer_reg[14]/NET0131 ,
		_w1062_,
		_w1063_
	);
	LUT2 #(
		.INIT('h8)
	) name611 (
		_w1061_,
		_w1063_,
		_w1064_
	);
	LUT3 #(
		.INIT('h6c)
	) name612 (
		\InstAddrPointer_reg[8]/NET0131 ,
		\InstAddrPointer_reg[9]/NET0131 ,
		_w1044_,
		_w1065_
	);
	LUT4 #(
		.INIT('h28a0)
	) name613 (
		\InstAddrPointer_reg[10]/NET0131 ,
		\InstAddrPointer_reg[8]/NET0131 ,
		\InstAddrPointer_reg[9]/NET0131 ,
		_w1044_,
		_w1066_
	);
	LUT4 #(
		.INIT('h8000)
	) name614 (
		_w1061_,
		_w1063_,
		_w1066_,
		_w1058_,
		_w1067_
	);
	LUT4 #(
		.INIT('h8000)
	) name615 (
		\InstAddrPointer_reg[8]/NET0131 ,
		\InstAddrPointer_reg[9]/NET0131 ,
		_w870_,
		_w1044_,
		_w1068_
	);
	LUT2 #(
		.INIT('h6)
	) name616 (
		\InstAddrPointer_reg[17]/NET0131 ,
		_w1068_,
		_w1069_
	);
	LUT3 #(
		.INIT('h48)
	) name617 (
		\InstAddrPointer_reg[17]/NET0131 ,
		_w873_,
		_w1068_,
		_w1070_
	);
	LUT3 #(
		.INIT('h80)
	) name618 (
		\InstAddrPointer_reg[20]/NET0131 ,
		_w874_,
		_w1068_,
		_w1071_
	);
	LUT3 #(
		.INIT('h6a)
	) name619 (
		\InstAddrPointer_reg[20]/NET0131 ,
		_w874_,
		_w1068_,
		_w1072_
	);
	LUT4 #(
		.INIT('h4888)
	) name620 (
		\InstAddrPointer_reg[20]/NET0131 ,
		\InstAddrPointer_reg[21]/NET0131 ,
		_w874_,
		_w1068_,
		_w1073_
	);
	LUT4 #(
		.INIT('h8000)
	) name621 (
		_w1054_,
		_w1067_,
		_w1070_,
		_w1073_,
		_w1074_
	);
	LUT3 #(
		.INIT('h80)
	) name622 (
		_w874_,
		_w878_,
		_w1068_,
		_w1075_
	);
	LUT4 #(
		.INIT('h8000)
	) name623 (
		_w889_,
		_w874_,
		_w878_,
		_w1068_,
		_w1076_
	);
	LUT4 #(
		.INIT('h8000)
	) name624 (
		\InstAddrPointer_reg[29]/NET0131 ,
		\InstAddrPointer_reg[30]/NET0131 ,
		_w893_,
		_w1076_,
		_w1077_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name625 (
		\InstAddrPointer_reg[29]/NET0131 ,
		\InstAddrPointer_reg[30]/NET0131 ,
		_w893_,
		_w1076_,
		_w1078_
	);
	LUT4 #(
		.INIT('h8000)
	) name626 (
		\InstAddrPointer_reg[24]/NET0131 ,
		_w874_,
		_w878_,
		_w1068_,
		_w1079_
	);
	LUT2 #(
		.INIT('h8)
	) name627 (
		\InstAddrPointer_reg[25]/NET0131 ,
		_w1079_,
		_w1080_
	);
	LUT4 #(
		.INIT('h78f0)
	) name628 (
		\InstAddrPointer_reg[24]/NET0131 ,
		\InstAddrPointer_reg[25]/NET0131 ,
		\InstAddrPointer_reg[26]/NET0131 ,
		_w1075_,
		_w1081_
	);
	LUT4 #(
		.INIT('h8000)
	) name629 (
		\InstAddrPointer_reg[22]/NET0131 ,
		_w876_,
		_w874_,
		_w1068_,
		_w1082_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name630 (
		\InstAddrPointer_reg[22]/NET0131 ,
		_w876_,
		_w874_,
		_w1068_,
		_w1083_
	);
	LUT2 #(
		.INIT('h8)
	) name631 (
		\InstAddrPointer_reg[23]/NET0131 ,
		_w1083_,
		_w1084_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name632 (
		\InstAddrPointer_reg[24]/NET0131 ,
		_w874_,
		_w878_,
		_w1068_,
		_w1085_
	);
	LUT3 #(
		.INIT('h80)
	) name633 (
		\InstAddrPointer_reg[23]/NET0131 ,
		_w1083_,
		_w1085_,
		_w1086_
	);
	LUT4 #(
		.INIT('h8000)
	) name634 (
		\InstAddrPointer_reg[23]/NET0131 ,
		\InstAddrPointer_reg[25]/NET0131 ,
		_w1083_,
		_w1085_,
		_w1087_
	);
	LUT2 #(
		.INIT('h8)
	) name635 (
		_w1081_,
		_w1087_,
		_w1088_
	);
	LUT3 #(
		.INIT('h6a)
	) name636 (
		\InstAddrPointer_reg[29]/NET0131 ,
		_w893_,
		_w1076_,
		_w1089_
	);
	LUT3 #(
		.INIT('h6c)
	) name637 (
		\InstAddrPointer_reg[27]/NET0131 ,
		\InstAddrPointer_reg[28]/NET0131 ,
		_w1076_,
		_w1090_
	);
	LUT4 #(
		.INIT('h2080)
	) name638 (
		\InstAddrPointer_reg[27]/NET0131 ,
		\InstAddrPointer_reg[28]/NET0131 ,
		\InstAddrPointer_reg[29]/NET0131 ,
		_w1076_,
		_w1091_
	);
	LUT3 #(
		.INIT('h80)
	) name639 (
		_w1081_,
		_w1087_,
		_w1091_,
		_w1092_
	);
	LUT4 #(
		.INIT('h8000)
	) name640 (
		_w1078_,
		_w1081_,
		_w1087_,
		_w1091_,
		_w1093_
	);
	LUT2 #(
		.INIT('h9)
	) name641 (
		\InstAddrPointer_reg[31]/NET0131 ,
		_w1077_,
		_w1094_
	);
	LUT4 #(
		.INIT('h802a)
	) name642 (
		_w688_,
		_w1074_,
		_w1093_,
		_w1094_,
		_w1095_
	);
	LUT4 #(
		.INIT('h00f4)
	) name643 (
		_w514_,
		_w569_,
		_w570_,
		_w634_,
		_w1096_
	);
	LUT2 #(
		.INIT('h2)
	) name644 (
		_w566_,
		_w611_,
		_w1097_
	);
	LUT3 #(
		.INIT('h01)
	) name645 (
		_w625_,
		_w683_,
		_w1097_,
		_w1098_
	);
	LUT4 #(
		.INIT('h0001)
	) name646 (
		_w625_,
		_w635_,
		_w683_,
		_w1097_,
		_w1099_
	);
	LUT2 #(
		.INIT('h8)
	) name647 (
		_w566_,
		_w611_,
		_w1100_
	);
	LUT3 #(
		.INIT('h80)
	) name648 (
		READY_n_pad,
		_w566_,
		_w611_,
		_w1101_
	);
	LUT4 #(
		.INIT('haa8a)
	) name649 (
		\InstAddrPointer_reg[31]/NET0131 ,
		_w1096_,
		_w1099_,
		_w1101_,
		_w1102_
	);
	LUT2 #(
		.INIT('h2)
	) name650 (
		_w606_,
		_w1094_,
		_w1103_
	);
	LUT3 #(
		.INIT('h0b)
	) name651 (
		_w582_,
		_w595_,
		_w1022_,
		_w1104_
	);
	LUT2 #(
		.INIT('h1)
	) name652 (
		_w645_,
		_w922_,
		_w1105_
	);
	LUT4 #(
		.INIT('h0001)
	) name653 (
		_w1104_,
		_w1102_,
		_w1105_,
		_w1103_,
		_w1106_
	);
	LUT2 #(
		.INIT('h4)
	) name654 (
		_w1095_,
		_w1106_,
		_w1107_
	);
	LUT4 #(
		.INIT('h08cc)
	) name655 (
		_w574_,
		_w695_,
		_w1024_,
		_w1107_,
		_w1108_
	);
	LUT4 #(
		.INIT('h0001)
	) name656 (
		\State2_reg[0]/NET0131 ,
		\State2_reg[1]/NET0131 ,
		\State2_reg[2]/NET0131 ,
		\State2_reg[3]/NET0131 ,
		_w1109_
	);
	LUT4 #(
		.INIT('hfc21)
	) name657 (
		\State2_reg[0]/NET0131 ,
		\State2_reg[1]/NET0131 ,
		\State2_reg[2]/NET0131 ,
		\State2_reg[3]/NET0131 ,
		_w1110_
	);
	LUT4 #(
		.INIT('h3f15)
	) name658 (
		\InstAddrPointer_reg[31]/NET0131 ,
		\rEIP_reg[31]/NET0131 ,
		_w1109_,
		_w1110_,
		_w1111_
	);
	LUT2 #(
		.INIT('hb)
	) name659 (
		_w1108_,
		_w1111_,
		_w1112_
	);
	LUT2 #(
		.INIT('h8)
	) name660 (
		_w736_,
		_w934_,
		_w1113_
	);
	LUT2 #(
		.INIT('h4)
	) name661 (
		_w863_,
		_w1113_,
		_w1114_
	);
	LUT3 #(
		.INIT('h40)
	) name662 (
		_w863_,
		_w916_,
		_w1113_,
		_w1115_
	);
	LUT4 #(
		.INIT('h4000)
	) name663 (
		_w863_,
		_w898_,
		_w916_,
		_w1113_,
		_w1116_
	);
	LUT2 #(
		.INIT('h6)
	) name664 (
		\InstAddrPointer_reg[30]/NET0131 ,
		_w896_,
		_w1117_
	);
	LUT4 #(
		.INIT('h4000)
	) name665 (
		_w863_,
		_w899_,
		_w916_,
		_w1113_,
		_w1118_
	);
	LUT4 #(
		.INIT('h00a8)
	) name666 (
		_w844_,
		_w1116_,
		_w1117_,
		_w1118_,
		_w1119_
	);
	LUT2 #(
		.INIT('h1)
	) name667 (
		_w951_,
		_w964_,
		_w1120_
	);
	LUT3 #(
		.INIT('h01)
	) name668 (
		_w948_,
		_w958_,
		_w960_,
		_w1121_
	);
	LUT3 #(
		.INIT('h0b)
	) name669 (
		_w948_,
		_w963_,
		_w967_,
		_w1122_
	);
	LUT4 #(
		.INIT('h4f00)
	) name670 (
		_w956_,
		_w1120_,
		_w1121_,
		_w1122_,
		_w1123_
	);
	LUT2 #(
		.INIT('h1)
	) name671 (
		_w944_,
		_w946_,
		_w1124_
	);
	LUT3 #(
		.INIT('h54)
	) name672 (
		_w944_,
		_w966_,
		_w975_,
		_w1125_
	);
	LUT3 #(
		.INIT('h0b)
	) name673 (
		_w1123_,
		_w1124_,
		_w1125_,
		_w1126_
	);
	LUT4 #(
		.INIT('h0045)
	) name674 (
		_w976_,
		_w1123_,
		_w1124_,
		_w1125_,
		_w1127_
	);
	LUT3 #(
		.INIT('h02)
	) name675 (
		_w974_,
		_w982_,
		_w983_,
		_w1128_
	);
	LUT4 #(
		.INIT('h0002)
	) name676 (
		_w974_,
		_w982_,
		_w983_,
		_w985_,
		_w1129_
	);
	LUT4 #(
		.INIT('h00e0)
	) name677 (
		_w989_,
		_w990_,
		_w994_,
		_w998_,
		_w1130_
	);
	LUT4 #(
		.INIT('h0054)
	) name678 (
		_w986_,
		_w1006_,
		_w1003_,
		_w1008_,
		_w1131_
	);
	LUT3 #(
		.INIT('h40)
	) name679 (
		_w988_,
		_w1130_,
		_w1131_,
		_w1132_
	);
	LUT2 #(
		.INIT('h4)
	) name680 (
		_w1009_,
		_w1005_,
		_w1133_
	);
	LUT2 #(
		.INIT('h8)
	) name681 (
		_w1132_,
		_w1133_,
		_w1134_
	);
	LUT3 #(
		.INIT('h80)
	) name682 (
		_w1010_,
		_w1018_,
		_w1019_,
		_w1135_
	);
	LUT4 #(
		.INIT('h8000)
	) name683 (
		_w1127_,
		_w1129_,
		_w1134_,
		_w1135_,
		_w1136_
	);
	LUT4 #(
		.INIT('hafae)
	) name684 (
		_w844_,
		_w1014_,
		_w1021_,
		_w1136_,
		_w1137_
	);
	LUT4 #(
		.INIT('h1d11)
	) name685 (
		\InstAddrPointer_reg[30]/NET0131 ,
		_w681_,
		_w1119_,
		_w1137_,
		_w1138_
	);
	LUT3 #(
		.INIT('h48)
	) name686 (
		\InstAddrPointer_reg[8]/NET0131 ,
		\InstAddrPointer_reg[9]/NET0131 ,
		_w1044_,
		_w1139_
	);
	LUT3 #(
		.INIT('h01)
	) name687 (
		_w1040_,
		_w1027_,
		_w1029_,
		_w1140_
	);
	LUT4 #(
		.INIT('hf100)
	) name688 (
		_w1031_,
		_w1034_,
		_w1036_,
		_w1140_,
		_w1141_
	);
	LUT3 #(
		.INIT('h54)
	) name689 (
		_w1040_,
		_w1035_,
		_w1048_,
		_w1142_
	);
	LUT2 #(
		.INIT('h1)
	) name690 (
		_w1042_,
		_w1051_,
		_w1143_
	);
	LUT3 #(
		.INIT('h51)
	) name691 (
		_w1046_,
		_w1047_,
		_w1051_,
		_w1144_
	);
	LUT4 #(
		.INIT('h1f00)
	) name692 (
		_w1141_,
		_w1142_,
		_w1143_,
		_w1144_,
		_w1145_
	);
	LUT4 #(
		.INIT('h4080)
	) name693 (
		\InstAddrPointer_reg[11]/NET0131 ,
		\InstAddrPointer_reg[12]/NET0131 ,
		\InstAddrPointer_reg[13]/NET0131 ,
		_w1059_,
		_w1146_
	);
	LUT2 #(
		.INIT('h6)
	) name694 (
		\InstAddrPointer_reg[14]/NET0131 ,
		_w1056_,
		_w1147_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name695 (
		\InstAddrPointer_reg[10]/NET0131 ,
		\InstAddrPointer_reg[8]/NET0131 ,
		\InstAddrPointer_reg[9]/NET0131 ,
		_w1044_,
		_w1148_
	);
	LUT3 #(
		.INIT('h60)
	) name696 (
		\InstAddrPointer_reg[17]/NET0131 ,
		_w1068_,
		_w1148_,
		_w1149_
	);
	LUT4 #(
		.INIT('h8000)
	) name697 (
		_w1058_,
		_w1146_,
		_w1147_,
		_w1149_,
		_w1150_
	);
	LUT3 #(
		.INIT('h20)
	) name698 (
		_w1139_,
		_w1145_,
		_w1150_,
		_w1151_
	);
	LUT3 #(
		.INIT('h6c)
	) name699 (
		\InstAddrPointer_reg[17]/NET0131 ,
		\InstAddrPointer_reg[18]/NET0131 ,
		_w1068_,
		_w1152_
	);
	LUT4 #(
		.INIT('h60c0)
	) name700 (
		\InstAddrPointer_reg[17]/NET0131 ,
		\InstAddrPointer_reg[18]/NET0131 ,
		\InstAddrPointer_reg[19]/NET0131 ,
		_w1068_,
		_w1153_
	);
	LUT2 #(
		.INIT('h8)
	) name701 (
		_w1073_,
		_w1153_,
		_w1154_
	);
	LUT4 #(
		.INIT('h2000)
	) name702 (
		_w1139_,
		_w1145_,
		_w1150_,
		_w1154_,
		_w1155_
	);
	LUT4 #(
		.INIT('h2888)
	) name703 (
		_w688_,
		_w1078_,
		_w1092_,
		_w1155_,
		_w1156_
	);
	LUT3 #(
		.INIT('h0b)
	) name704 (
		_w582_,
		_w595_,
		_w1014_,
		_w1157_
	);
	LUT3 #(
		.INIT('h01)
	) name705 (
		_w621_,
		_w622_,
		_w1101_,
		_w1158_
	);
	LUT3 #(
		.INIT('h2a)
	) name706 (
		\InstAddrPointer_reg[30]/NET0131 ,
		_w1098_,
		_w1158_,
		_w1159_
	);
	LUT2 #(
		.INIT('h8)
	) name707 (
		_w606_,
		_w1078_,
		_w1160_
	);
	LUT3 #(
		.INIT('h0b)
	) name708 (
		_w620_,
		_w1117_,
		_w1160_,
		_w1161_
	);
	LUT3 #(
		.INIT('h10)
	) name709 (
		_w1157_,
		_w1159_,
		_w1161_,
		_w1162_
	);
	LUT2 #(
		.INIT('h4)
	) name710 (
		_w1156_,
		_w1162_,
		_w1163_
	);
	LUT4 #(
		.INIT('h08cc)
	) name711 (
		_w574_,
		_w695_,
		_w1138_,
		_w1163_,
		_w1164_
	);
	LUT4 #(
		.INIT('h3f15)
	) name712 (
		\InstAddrPointer_reg[30]/NET0131 ,
		\rEIP_reg[30]/NET0131 ,
		_w1109_,
		_w1110_,
		_w1165_
	);
	LUT2 #(
		.INIT('hb)
	) name713 (
		_w1164_,
		_w1165_,
		_w1166_
	);
	LUT2 #(
		.INIT('h2)
	) name714 (
		\InstAddrPointer_reg[28]/NET0131 ,
		_w681_,
		_w1167_
	);
	LUT4 #(
		.INIT('h8000)
	) name715 (
		_w736_,
		_w907_,
		_w910_,
		_w934_,
		_w1168_
	);
	LUT4 #(
		.INIT('h4888)
	) name716 (
		\InstAddrPointer_reg[22]/NET0131 ,
		\InstAddrPointer_reg[23]/NET0131 ,
		_w876_,
		_w875_,
		_w1169_
	);
	LUT2 #(
		.INIT('h8)
	) name717 (
		_w914_,
		_w1169_,
		_w1170_
	);
	LUT3 #(
		.INIT('h40)
	) name718 (
		_w863_,
		_w1168_,
		_w1170_,
		_w1171_
	);
	LUT3 #(
		.INIT('h80)
	) name719 (
		_w891_,
		_w884_,
		_w886_,
		_w1172_
	);
	LUT4 #(
		.INIT('h4000)
	) name720 (
		_w863_,
		_w1168_,
		_w1170_,
		_w1172_,
		_w1173_
	);
	LUT2 #(
		.INIT('h9)
	) name721 (
		\InstAddrPointer_reg[28]/NET0131 ,
		_w890_,
		_w1174_
	);
	LUT3 #(
		.INIT('h28)
	) name722 (
		_w844_,
		_w1173_,
		_w1174_,
		_w1175_
	);
	LUT4 #(
		.INIT('h0020)
	) name723 (
		_w974_,
		_w976_,
		_w987_,
		_w988_,
		_w1176_
	);
	LUT4 #(
		.INIT('h0b00)
	) name724 (
		_w1123_,
		_w1124_,
		_w1125_,
		_w1176_,
		_w1177_
	);
	LUT3 #(
		.INIT('h08)
	) name725 (
		_w1005_,
		_w1012_,
		_w1016_,
		_w1178_
	);
	LUT3 #(
		.INIT('h80)
	) name726 (
		_w1130_,
		_w1177_,
		_w1178_,
		_w1179_
	);
	LUT4 #(
		.INIT('h8aa8)
	) name727 (
		_w681_,
		_w844_,
		_w1017_,
		_w1179_,
		_w1180_
	);
	LUT4 #(
		.INIT('h8a88)
	) name728 (
		_w574_,
		_w1167_,
		_w1175_,
		_w1180_,
		_w1181_
	);
	LUT4 #(
		.INIT('h2080)
	) name729 (
		\InstAddrPointer_reg[11]/NET0131 ,
		\InstAddrPointer_reg[8]/NET0131 ,
		\InstAddrPointer_reg[9]/NET0131 ,
		_w1044_,
		_w1182_
	);
	LUT2 #(
		.INIT('h8)
	) name730 (
		_w1148_,
		_w1182_,
		_w1183_
	);
	LUT4 #(
		.INIT('h0e0c)
	) name731 (
		\InstAddrPointer_reg[11]/NET0131 ,
		\InstAddrPointer_reg[12]/NET0131 ,
		_w1055_,
		_w1059_,
		_w1184_
	);
	LUT2 #(
		.INIT('h8)
	) name732 (
		_w868_,
		_w1184_,
		_w1185_
	);
	LUT3 #(
		.INIT('h40)
	) name733 (
		_w1145_,
		_w1183_,
		_w1185_,
		_w1186_
	);
	LUT4 #(
		.INIT('h070f)
	) name734 (
		\InstAddrPointer_reg[14]/NET0131 ,
		\InstAddrPointer_reg[15]/NET0131 ,
		\InstAddrPointer_reg[16]/NET0131 ,
		_w1056_,
		_w1187_
	);
	LUT2 #(
		.INIT('h1)
	) name735 (
		_w1068_,
		_w1187_,
		_w1188_
	);
	LUT3 #(
		.INIT('h02)
	) name736 (
		_w874_,
		_w1068_,
		_w1187_,
		_w1189_
	);
	LUT4 #(
		.INIT('h4000)
	) name737 (
		_w1145_,
		_w1183_,
		_w1185_,
		_w1189_,
		_w1190_
	);
	LUT2 #(
		.INIT('h6)
	) name738 (
		\InstAddrPointer_reg[27]/NET0131 ,
		_w1076_,
		_w1191_
	);
	LUT3 #(
		.INIT('h48)
	) name739 (
		\InstAddrPointer_reg[27]/NET0131 ,
		_w1073_,
		_w1076_,
		_w1192_
	);
	LUT3 #(
		.INIT('h80)
	) name740 (
		_w1081_,
		_w1087_,
		_w1192_,
		_w1193_
	);
	LUT4 #(
		.INIT('h2888)
	) name741 (
		_w688_,
		_w1090_,
		_w1190_,
		_w1193_,
		_w1194_
	);
	LUT4 #(
		.INIT('h00f4)
	) name742 (
		_w514_,
		_w569_,
		_w570_,
		_w659_,
		_w1195_
	);
	LUT4 #(
		.INIT('h00ec)
	) name743 (
		_w514_,
		_w566_,
		_w569_,
		_w611_,
		_w1196_
	);
	LUT4 #(
		.INIT('h0001)
	) name744 (
		_w625_,
		_w683_,
		_w1195_,
		_w1196_,
		_w1197_
	);
	LUT3 #(
		.INIT('ha2)
	) name745 (
		READY_n_pad,
		_w613_,
		_w643_,
		_w1198_
	);
	LUT3 #(
		.INIT('ha2)
	) name746 (
		\InstAddrPointer_reg[28]/NET0131 ,
		_w1197_,
		_w1198_,
		_w1199_
	);
	LUT4 #(
		.INIT('haa20)
	) name747 (
		\InstAddrPointer_reg[28]/NET0131 ,
		_w514_,
		_w569_,
		_w570_,
		_w1200_
	);
	LUT3 #(
		.INIT('h31)
	) name748 (
		_w620_,
		_w1174_,
		_w1200_,
		_w1201_
	);
	LUT2 #(
		.INIT('h8)
	) name749 (
		_w606_,
		_w1090_,
		_w1202_
	);
	LUT4 #(
		.INIT('h004f)
	) name750 (
		_w582_,
		_w595_,
		_w1017_,
		_w1202_,
		_w1203_
	);
	LUT3 #(
		.INIT('h10)
	) name751 (
		_w1201_,
		_w1199_,
		_w1203_,
		_w1204_
	);
	LUT2 #(
		.INIT('h4)
	) name752 (
		_w1194_,
		_w1204_,
		_w1205_
	);
	LUT4 #(
		.INIT('h3f15)
	) name753 (
		\InstAddrPointer_reg[28]/NET0131 ,
		\rEIP_reg[28]/NET0131 ,
		_w1109_,
		_w1110_,
		_w1206_
	);
	LUT4 #(
		.INIT('h8aff)
	) name754 (
		_w695_,
		_w1181_,
		_w1205_,
		_w1206_,
		_w1207_
	);
	LUT2 #(
		.INIT('h2)
	) name755 (
		\InstAddrPointer_reg[23]/NET0131 ,
		_w681_,
		_w1208_
	);
	LUT4 #(
		.INIT('h000e)
	) name756 (
		_w1006_,
		_w1003_,
		_w1008_,
		_w1004_,
		_w1209_
	);
	LUT2 #(
		.INIT('h8)
	) name757 (
		_w979_,
		_w987_,
		_w1210_
	);
	LUT4 #(
		.INIT('h0800)
	) name758 (
		_w979_,
		_w987_,
		_w988_,
		_w1130_,
		_w1211_
	);
	LUT2 #(
		.INIT('h4)
	) name759 (
		_w1002_,
		_w1209_,
		_w1212_
	);
	LUT4 #(
		.INIT('h4111)
	) name760 (
		_w844_,
		_w1002_,
		_w1209_,
		_w1211_,
		_w1213_
	);
	LUT3 #(
		.INIT('h15)
	) name761 (
		_w887_,
		_w933_,
		_w936_,
		_w1214_
	);
	LUT4 #(
		.INIT('h222a)
	) name762 (
		_w681_,
		_w844_,
		_w1171_,
		_w1214_,
		_w1215_
	);
	LUT4 #(
		.INIT('h8a88)
	) name763 (
		_w574_,
		_w1208_,
		_w1213_,
		_w1215_,
		_w1216_
	);
	LUT3 #(
		.INIT('h80)
	) name764 (
		_w1073_,
		_w1084_,
		_w1190_,
		_w1217_
	);
	LUT3 #(
		.INIT('h32)
	) name765 (
		\InstAddrPointer_reg[23]/NET0131 ,
		_w1075_,
		_w1082_,
		_w1218_
	);
	LUT4 #(
		.INIT('haa80)
	) name766 (
		_w688_,
		_w1074_,
		_w1083_,
		_w1218_,
		_w1219_
	);
	LUT4 #(
		.INIT('h0004)
	) name767 (
		_w625_,
		_w636_,
		_w683_,
		_w1096_,
		_w1220_
	);
	LUT4 #(
		.INIT('h00c8)
	) name768 (
		_w552_,
		_w576_,
		_w579_,
		_w1082_,
		_w1221_
	);
	LUT3 #(
		.INIT('ha2)
	) name769 (
		\InstAddrPointer_reg[23]/NET0131 ,
		_w1220_,
		_w1221_,
		_w1222_
	);
	LUT2 #(
		.INIT('h4)
	) name770 (
		_w620_,
		_w887_,
		_w1223_
	);
	LUT2 #(
		.INIT('h8)
	) name771 (
		_w606_,
		_w1218_,
		_w1224_
	);
	LUT4 #(
		.INIT('h004f)
	) name772 (
		_w582_,
		_w595_,
		_w1002_,
		_w1224_,
		_w1225_
	);
	LUT3 #(
		.INIT('h10)
	) name773 (
		_w1223_,
		_w1222_,
		_w1225_,
		_w1226_
	);
	LUT3 #(
		.INIT('hb0)
	) name774 (
		_w1217_,
		_w1219_,
		_w1226_,
		_w1227_
	);
	LUT2 #(
		.INIT('h8)
	) name775 (
		\rEIP_reg[23]/NET0131 ,
		_w1109_,
		_w1228_
	);
	LUT4 #(
		.INIT('h3f15)
	) name776 (
		\InstAddrPointer_reg[23]/NET0131 ,
		\rEIP_reg[23]/NET0131 ,
		_w1109_,
		_w1110_,
		_w1229_
	);
	LUT4 #(
		.INIT('h8aff)
	) name777 (
		_w695_,
		_w1216_,
		_w1227_,
		_w1229_,
		_w1230_
	);
	LUT4 #(
		.INIT('h1555)
	) name778 (
		_w891_,
		_w888_,
		_w933_,
		_w936_,
		_w1231_
	);
	LUT3 #(
		.INIT('h02)
	) name779 (
		_w844_,
		_w1173_,
		_w1231_,
		_w1232_
	);
	LUT4 #(
		.INIT('h8000)
	) name780 (
		_w979_,
		_w996_,
		_w1013_,
		_w1016_,
		_w1233_
	);
	LUT4 #(
		.INIT('h007f)
	) name781 (
		_w979_,
		_w996_,
		_w1013_,
		_w1016_,
		_w1234_
	);
	LUT3 #(
		.INIT('h01)
	) name782 (
		_w844_,
		_w1234_,
		_w1233_,
		_w1235_
	);
	LUT4 #(
		.INIT('h111d)
	) name783 (
		\InstAddrPointer_reg[27]/NET0131 ,
		_w681_,
		_w1232_,
		_w1235_,
		_w1236_
	);
	LUT3 #(
		.INIT('h07)
	) name784 (
		_w1074_,
		_w1088_,
		_w1191_,
		_w1237_
	);
	LUT4 #(
		.INIT('h8000)
	) name785 (
		_w1054_,
		_w1067_,
		_w1070_,
		_w1193_,
		_w1238_
	);
	LUT2 #(
		.INIT('h2)
	) name786 (
		_w688_,
		_w1238_,
		_w1239_
	);
	LUT4 #(
		.INIT('h00c8)
	) name787 (
		_w552_,
		_w576_,
		_w579_,
		_w1076_,
		_w1240_
	);
	LUT4 #(
		.INIT('haa8a)
	) name788 (
		\InstAddrPointer_reg[27]/NET0131 ,
		_w1096_,
		_w1099_,
		_w1240_,
		_w1241_
	);
	LUT3 #(
		.INIT('h80)
	) name789 (
		\InstAddrPointer_reg[27]/NET0131 ,
		READY_n_pad,
		_w566_,
		_w1242_
	);
	LUT2 #(
		.INIT('h4)
	) name790 (
		READY_n_pad,
		_w891_,
		_w1243_
	);
	LUT4 #(
		.INIT('h040f)
	) name791 (
		_w618_,
		_w619_,
		_w1242_,
		_w1243_,
		_w1244_
	);
	LUT2 #(
		.INIT('h2)
	) name792 (
		_w611_,
		_w1244_,
		_w1245_
	);
	LUT2 #(
		.INIT('h8)
	) name793 (
		_w549_,
		_w891_,
		_w1246_
	);
	LUT3 #(
		.INIT('h07)
	) name794 (
		_w606_,
		_w1191_,
		_w1246_,
		_w1247_
	);
	LUT4 #(
		.INIT('h4f00)
	) name795 (
		_w582_,
		_w595_,
		_w1016_,
		_w1247_,
		_w1248_
	);
	LUT3 #(
		.INIT('h10)
	) name796 (
		_w1241_,
		_w1245_,
		_w1248_,
		_w1249_
	);
	LUT3 #(
		.INIT('hb0)
	) name797 (
		_w1237_,
		_w1239_,
		_w1249_,
		_w1250_
	);
	LUT4 #(
		.INIT('h08cc)
	) name798 (
		_w574_,
		_w695_,
		_w1236_,
		_w1250_,
		_w1251_
	);
	LUT4 #(
		.INIT('h3f15)
	) name799 (
		\InstAddrPointer_reg[27]/NET0131 ,
		\rEIP_reg[27]/NET0131 ,
		_w1109_,
		_w1110_,
		_w1252_
	);
	LUT2 #(
		.INIT('hb)
	) name800 (
		_w1251_,
		_w1252_,
		_w1253_
	);
	LUT4 #(
		.INIT('h1d11)
	) name801 (
		\PhyAddrPointer_reg[31]/NET0131 ,
		_w681_,
		_w939_,
		_w1023_,
		_w1254_
	);
	LUT4 #(
		.INIT('h028a)
	) name802 (
		\PhyAddrPointer_reg[31]/NET0131 ,
		_w573_,
		_w574_,
		_w605_,
		_w1255_
	);
	LUT2 #(
		.INIT('h1)
	) name803 (
		_w1095_,
		_w1255_,
		_w1256_
	);
	LUT4 #(
		.INIT('h08cc)
	) name804 (
		_w574_,
		_w695_,
		_w1254_,
		_w1256_,
		_w1257_
	);
	LUT3 #(
		.INIT('h80)
	) name805 (
		\PhyAddrPointer_reg[2]/NET0131 ,
		\PhyAddrPointer_reg[3]/NET0131 ,
		\PhyAddrPointer_reg[4]/NET0131 ,
		_w1258_
	);
	LUT4 #(
		.INIT('h8000)
	) name806 (
		\PhyAddrPointer_reg[2]/NET0131 ,
		\PhyAddrPointer_reg[3]/NET0131 ,
		\PhyAddrPointer_reg[4]/NET0131 ,
		\PhyAddrPointer_reg[5]/NET0131 ,
		_w1259_
	);
	LUT3 #(
		.INIT('h80)
	) name807 (
		\PhyAddrPointer_reg[6]/NET0131 ,
		\PhyAddrPointer_reg[7]/NET0131 ,
		_w1259_,
		_w1260_
	);
	LUT4 #(
		.INIT('h8000)
	) name808 (
		\PhyAddrPointer_reg[6]/NET0131 ,
		\PhyAddrPointer_reg[7]/NET0131 ,
		\PhyAddrPointer_reg[8]/NET0131 ,
		_w1259_,
		_w1261_
	);
	LUT3 #(
		.INIT('h80)
	) name809 (
		\PhyAddrPointer_reg[10]/NET0131 ,
		\PhyAddrPointer_reg[9]/NET0131 ,
		_w1261_,
		_w1262_
	);
	LUT4 #(
		.INIT('h8000)
	) name810 (
		\PhyAddrPointer_reg[10]/NET0131 ,
		\PhyAddrPointer_reg[11]/NET0131 ,
		\PhyAddrPointer_reg[9]/NET0131 ,
		_w1261_,
		_w1263_
	);
	LUT3 #(
		.INIT('h80)
	) name811 (
		\PhyAddrPointer_reg[12]/NET0131 ,
		\PhyAddrPointer_reg[13]/NET0131 ,
		_w1263_,
		_w1264_
	);
	LUT2 #(
		.INIT('h8)
	) name812 (
		\PhyAddrPointer_reg[14]/NET0131 ,
		\PhyAddrPointer_reg[15]/NET0131 ,
		_w1265_
	);
	LUT3 #(
		.INIT('h80)
	) name813 (
		\PhyAddrPointer_reg[14]/NET0131 ,
		\PhyAddrPointer_reg[15]/NET0131 ,
		\PhyAddrPointer_reg[16]/NET0131 ,
		_w1266_
	);
	LUT4 #(
		.INIT('h8000)
	) name814 (
		\PhyAddrPointer_reg[14]/NET0131 ,
		\PhyAddrPointer_reg[15]/NET0131 ,
		\PhyAddrPointer_reg[16]/NET0131 ,
		\PhyAddrPointer_reg[17]/NET0131 ,
		_w1267_
	);
	LUT2 #(
		.INIT('h8)
	) name815 (
		\PhyAddrPointer_reg[18]/NET0131 ,
		\PhyAddrPointer_reg[19]/NET0131 ,
		_w1268_
	);
	LUT3 #(
		.INIT('h80)
	) name816 (
		\PhyAddrPointer_reg[18]/NET0131 ,
		\PhyAddrPointer_reg[19]/NET0131 ,
		\PhyAddrPointer_reg[20]/NET0131 ,
		_w1269_
	);
	LUT4 #(
		.INIT('h8000)
	) name817 (
		\PhyAddrPointer_reg[18]/NET0131 ,
		\PhyAddrPointer_reg[19]/NET0131 ,
		\PhyAddrPointer_reg[20]/NET0131 ,
		\PhyAddrPointer_reg[21]/NET0131 ,
		_w1270_
	);
	LUT2 #(
		.INIT('h8)
	) name818 (
		_w1267_,
		_w1270_,
		_w1271_
	);
	LUT4 #(
		.INIT('h8000)
	) name819 (
		\PhyAddrPointer_reg[12]/NET0131 ,
		\PhyAddrPointer_reg[13]/NET0131 ,
		_w1263_,
		_w1271_,
		_w1272_
	);
	LUT2 #(
		.INIT('h8)
	) name820 (
		\PhyAddrPointer_reg[22]/NET0131 ,
		\PhyAddrPointer_reg[23]/NET0131 ,
		_w1273_
	);
	LUT3 #(
		.INIT('h80)
	) name821 (
		\PhyAddrPointer_reg[24]/NET0131 ,
		_w1272_,
		_w1273_,
		_w1274_
	);
	LUT2 #(
		.INIT('h8)
	) name822 (
		\PhyAddrPointer_reg[25]/NET0131 ,
		\PhyAddrPointer_reg[26]/NET0131 ,
		_w1275_
	);
	LUT4 #(
		.INIT('h8000)
	) name823 (
		\PhyAddrPointer_reg[24]/NET0131 ,
		_w1272_,
		_w1273_,
		_w1275_,
		_w1276_
	);
	LUT3 #(
		.INIT('h80)
	) name824 (
		\PhyAddrPointer_reg[27]/NET0131 ,
		\PhyAddrPointer_reg[28]/NET0131 ,
		_w1276_,
		_w1277_
	);
	LUT4 #(
		.INIT('h8000)
	) name825 (
		\PhyAddrPointer_reg[27]/NET0131 ,
		\PhyAddrPointer_reg[28]/NET0131 ,
		\PhyAddrPointer_reg[29]/NET0131 ,
		_w1276_,
		_w1278_
	);
	LUT4 #(
		.INIT('h78f0)
	) name826 (
		\PhyAddrPointer_reg[1]/NET0131 ,
		\PhyAddrPointer_reg[30]/NET0131 ,
		\PhyAddrPointer_reg[31]/NET0131 ,
		_w1278_,
		_w1279_
	);
	LUT4 #(
		.INIT('hffeb)
	) name827 (
		\State2_reg[0]/NET0131 ,
		\State2_reg[1]/NET0131 ,
		\State2_reg[2]/NET0131 ,
		\State2_reg[3]/NET0131 ,
		_w1280_
	);
	LUT3 #(
		.INIT('h0d)
	) name828 (
		\DataWidth_reg[1]/NET0131 ,
		_w706_,
		_w1280_,
		_w1281_
	);
	LUT4 #(
		.INIT('h60c0)
	) name829 (
		\PhyAddrPointer_reg[30]/NET0131 ,
		\PhyAddrPointer_reg[31]/NET0131 ,
		_w707_,
		_w1278_,
		_w1282_
	);
	LUT4 #(
		.INIT('hfc35)
	) name830 (
		\State2_reg[0]/NET0131 ,
		\State2_reg[1]/NET0131 ,
		\State2_reg[2]/NET0131 ,
		\State2_reg[3]/NET0131 ,
		_w1283_
	);
	LUT4 #(
		.INIT('h3f15)
	) name831 (
		\PhyAddrPointer_reg[31]/NET0131 ,
		\rEIP_reg[31]/NET0131 ,
		_w1109_,
		_w1283_,
		_w1284_
	);
	LUT4 #(
		.INIT('h0700)
	) name832 (
		_w1279_,
		_w1281_,
		_w1282_,
		_w1284_,
		_w1285_
	);
	LUT2 #(
		.INIT('hb)
	) name833 (
		_w1257_,
		_w1285_,
		_w1286_
	);
	LUT3 #(
		.INIT('h32)
	) name834 (
		\InstAddrPointer_reg[19]/NET0131 ,
		_w875_,
		_w908_,
		_w1287_
	);
	LUT4 #(
		.INIT('h4000)
	) name835 (
		_w863_,
		_w907_,
		_w909_,
		_w1113_,
		_w1288_
	);
	LUT3 #(
		.INIT('h8a)
	) name836 (
		_w844_,
		_w863_,
		_w1168_,
		_w1289_
	);
	LUT3 #(
		.INIT('he0)
	) name837 (
		_w1287_,
		_w1288_,
		_w1289_,
		_w1290_
	);
	LUT3 #(
		.INIT('h70)
	) name838 (
		_w979_,
		_w996_,
		_w998_,
		_w1291_
	);
	LUT3 #(
		.INIT('h54)
	) name839 (
		_w844_,
		_w1211_,
		_w1291_,
		_w1292_
	);
	LUT4 #(
		.INIT('h111d)
	) name840 (
		\InstAddrPointer_reg[19]/NET0131 ,
		_w681_,
		_w1290_,
		_w1292_,
		_w1293_
	);
	LUT4 #(
		.INIT('h78f0)
	) name841 (
		\InstAddrPointer_reg[17]/NET0131 ,
		\InstAddrPointer_reg[18]/NET0131 ,
		\InstAddrPointer_reg[19]/NET0131 ,
		_w1068_,
		_w1294_
	);
	LUT4 #(
		.INIT('h8000)
	) name842 (
		\InstAddrPointer_reg[18]/NET0131 ,
		_w1069_,
		_w1054_,
		_w1067_,
		_w1295_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name843 (
		_w688_,
		_w1054_,
		_w1067_,
		_w1070_,
		_w1296_
	);
	LUT3 #(
		.INIT('he0)
	) name844 (
		_w1294_,
		_w1295_,
		_w1296_,
		_w1297_
	);
	LUT3 #(
		.INIT('h2a)
	) name845 (
		\InstAddrPointer_reg[19]/NET0131 ,
		_w624_,
		_w684_,
		_w1298_
	);
	LUT2 #(
		.INIT('h4)
	) name846 (
		_w620_,
		_w1287_,
		_w1299_
	);
	LUT2 #(
		.INIT('h8)
	) name847 (
		_w606_,
		_w1294_,
		_w1300_
	);
	LUT4 #(
		.INIT('h004f)
	) name848 (
		_w582_,
		_w595_,
		_w998_,
		_w1300_,
		_w1301_
	);
	LUT3 #(
		.INIT('h10)
	) name849 (
		_w1299_,
		_w1298_,
		_w1301_,
		_w1302_
	);
	LUT2 #(
		.INIT('h4)
	) name850 (
		_w1297_,
		_w1302_,
		_w1303_
	);
	LUT4 #(
		.INIT('h08cc)
	) name851 (
		_w574_,
		_w695_,
		_w1293_,
		_w1303_,
		_w1304_
	);
	LUT2 #(
		.INIT('h8)
	) name852 (
		\rEIP_reg[19]/NET0131 ,
		_w1109_,
		_w1305_
	);
	LUT4 #(
		.INIT('h3f15)
	) name853 (
		\InstAddrPointer_reg[19]/NET0131 ,
		\rEIP_reg[19]/NET0131 ,
		_w1109_,
		_w1110_,
		_w1306_
	);
	LUT2 #(
		.INIT('hb)
	) name854 (
		_w1304_,
		_w1306_,
		_w1307_
	);
	LUT4 #(
		.INIT('h4111)
	) name855 (
		_w844_,
		_w1008_,
		_w1130_,
		_w1177_,
		_w1308_
	);
	LUT3 #(
		.INIT('h40)
	) name856 (
		_w863_,
		_w913_,
		_w1168_,
		_w1309_
	);
	LUT4 #(
		.INIT('h280a)
	) name857 (
		_w844_,
		_w863_,
		_w913_,
		_w1168_,
		_w1310_
	);
	LUT4 #(
		.INIT('hddd1)
	) name858 (
		\InstAddrPointer_reg[20]/NET0131 ,
		_w681_,
		_w1310_,
		_w1308_,
		_w1311_
	);
	LUT3 #(
		.INIT('h28)
	) name859 (
		_w688_,
		_w1072_,
		_w1190_,
		_w1312_
	);
	LUT4 #(
		.INIT('ha8a0)
	) name860 (
		\InstAddrPointer_reg[20]/NET0131 ,
		_w514_,
		_w566_,
		_w569_,
		_w1313_
	);
	LUT3 #(
		.INIT('hc4)
	) name861 (
		_w645_,
		_w913_,
		_w1313_,
		_w1314_
	);
	LUT2 #(
		.INIT('h2)
	) name862 (
		\InstAddrPointer_reg[20]/NET0131 ,
		_w1220_,
		_w1315_
	);
	LUT2 #(
		.INIT('h8)
	) name863 (
		_w606_,
		_w1072_,
		_w1316_
	);
	LUT4 #(
		.INIT('h004f)
	) name864 (
		_w582_,
		_w595_,
		_w1008_,
		_w1316_,
		_w1317_
	);
	LUT3 #(
		.INIT('h10)
	) name865 (
		_w1315_,
		_w1314_,
		_w1317_,
		_w1318_
	);
	LUT4 #(
		.INIT('h0d00)
	) name866 (
		_w574_,
		_w1311_,
		_w1312_,
		_w1318_,
		_w1319_
	);
	LUT4 #(
		.INIT('h3f15)
	) name867 (
		\InstAddrPointer_reg[20]/NET0131 ,
		\rEIP_reg[20]/NET0131 ,
		_w1109_,
		_w1110_,
		_w1320_
	);
	LUT3 #(
		.INIT('h2f)
	) name868 (
		_w695_,
		_w1319_,
		_w1320_,
		_w1321_
	);
	LUT2 #(
		.INIT('h2)
	) name869 (
		\InstAddrPointer_reg[22]/NET0131 ,
		_w681_,
		_w1322_
	);
	LUT4 #(
		.INIT('h2333)
	) name870 (
		_w863_,
		_w912_,
		_w914_,
		_w1168_,
		_w1323_
	);
	LUT3 #(
		.INIT('ha8)
	) name871 (
		_w844_,
		_w1115_,
		_w1323_,
		_w1324_
	);
	LUT3 #(
		.INIT('h80)
	) name872 (
		_w1127_,
		_w1129_,
		_w1132_,
		_w1325_
	);
	LUT4 #(
		.INIT('h8aa8)
	) name873 (
		_w681_,
		_w844_,
		_w1004_,
		_w1325_,
		_w1326_
	);
	LUT4 #(
		.INIT('h8a88)
	) name874 (
		_w574_,
		_w1322_,
		_w1324_,
		_w1326_,
		_w1327_
	);
	LUT3 #(
		.INIT('h28)
	) name875 (
		_w688_,
		_w1083_,
		_w1155_,
		_w1328_
	);
	LUT4 #(
		.INIT('ha080)
	) name876 (
		READY_n_pad,
		_w566_,
		_w611_,
		_w618_,
		_w1329_
	);
	LUT4 #(
		.INIT('haaa2)
	) name877 (
		\InstAddrPointer_reg[22]/NET0131 ,
		_w1099_,
		_w1195_,
		_w1329_,
		_w1330_
	);
	LUT2 #(
		.INIT('h4)
	) name878 (
		_w620_,
		_w912_,
		_w1331_
	);
	LUT2 #(
		.INIT('h8)
	) name879 (
		_w606_,
		_w1083_,
		_w1332_
	);
	LUT4 #(
		.INIT('h004f)
	) name880 (
		_w582_,
		_w595_,
		_w1004_,
		_w1332_,
		_w1333_
	);
	LUT3 #(
		.INIT('h10)
	) name881 (
		_w1330_,
		_w1331_,
		_w1333_,
		_w1334_
	);
	LUT2 #(
		.INIT('h4)
	) name882 (
		_w1328_,
		_w1334_,
		_w1335_
	);
	LUT4 #(
		.INIT('h3f15)
	) name883 (
		\InstAddrPointer_reg[22]/NET0131 ,
		\rEIP_reg[22]/NET0131 ,
		_w1109_,
		_w1110_,
		_w1336_
	);
	LUT4 #(
		.INIT('h8aff)
	) name884 (
		_w695_,
		_w1327_,
		_w1335_,
		_w1336_,
		_w1337_
	);
	LUT4 #(
		.INIT('h070f)
	) name885 (
		_w1073_,
		_w1084_,
		_w1085_,
		_w1190_,
		_w1338_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name886 (
		_w688_,
		_w1073_,
		_w1086_,
		_w1190_,
		_w1339_
	);
	LUT2 #(
		.INIT('h4)
	) name887 (
		_w1338_,
		_w1339_,
		_w1340_
	);
	LUT2 #(
		.INIT('h2)
	) name888 (
		\InstAddrPointer_reg[24]/NET0131 ,
		_w681_,
		_w1341_
	);
	LUT4 #(
		.INIT('h9ccc)
	) name889 (
		_w863_,
		_w886_,
		_w1168_,
		_w1170_,
		_w1342_
	);
	LUT2 #(
		.INIT('h2)
	) name890 (
		_w844_,
		_w1342_,
		_w1343_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name891 (
		_w1001_,
		_w1130_,
		_w1177_,
		_w1212_,
		_w1344_
	);
	LUT4 #(
		.INIT('h1f00)
	) name892 (
		_w951_,
		_w956_,
		_w961_,
		_w965_,
		_w1345_
	);
	LUT3 #(
		.INIT('h01)
	) name893 (
		_w944_,
		_w946_,
		_w948_,
		_w1346_
	);
	LUT4 #(
		.INIT('h3110)
	) name894 (
		_w857_,
		_w944_,
		_w945_,
		_w967_,
		_w1347_
	);
	LUT2 #(
		.INIT('h2)
	) name895 (
		_w977_,
		_w1347_,
		_w1348_
	);
	LUT4 #(
		.INIT('h8a00)
	) name896 (
		_w1128_,
		_w1345_,
		_w1346_,
		_w1348_,
		_w1349_
	);
	LUT3 #(
		.INIT('h01)
	) name897 (
		_w985_,
		_w986_,
		_w1008_,
		_w1350_
	);
	LUT3 #(
		.INIT('h40)
	) name898 (
		_w988_,
		_w1130_,
		_w1350_,
		_w1351_
	);
	LUT2 #(
		.INIT('h4)
	) name899 (
		_w1007_,
		_w1005_,
		_w1352_
	);
	LUT3 #(
		.INIT('h80)
	) name900 (
		_w1349_,
		_w1351_,
		_w1352_,
		_w1353_
	);
	LUT4 #(
		.INIT('h1555)
	) name901 (
		_w844_,
		_w1349_,
		_w1351_,
		_w1352_,
		_w1354_
	);
	LUT3 #(
		.INIT('h8a)
	) name902 (
		_w681_,
		_w1344_,
		_w1354_,
		_w1355_
	);
	LUT4 #(
		.INIT('h8a88)
	) name903 (
		_w574_,
		_w1341_,
		_w1343_,
		_w1355_,
		_w1356_
	);
	LUT2 #(
		.INIT('h2)
	) name904 (
		\InstAddrPointer_reg[24]/NET0131 ,
		_w1220_,
		_w1357_
	);
	LUT2 #(
		.INIT('h4)
	) name905 (
		_w645_,
		_w886_,
		_w1358_
	);
	LUT2 #(
		.INIT('h8)
	) name906 (
		_w606_,
		_w1085_,
		_w1359_
	);
	LUT4 #(
		.INIT('h004f)
	) name907 (
		_w582_,
		_w595_,
		_w1001_,
		_w1359_,
		_w1360_
	);
	LUT3 #(
		.INIT('h10)
	) name908 (
		_w1358_,
		_w1357_,
		_w1360_,
		_w1361_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name909 (
		_w695_,
		_w1356_,
		_w1340_,
		_w1361_,
		_w1362_
	);
	LUT2 #(
		.INIT('h8)
	) name910 (
		\rEIP_reg[24]/NET0131 ,
		_w1109_,
		_w1363_
	);
	LUT4 #(
		.INIT('h3f15)
	) name911 (
		\InstAddrPointer_reg[24]/NET0131 ,
		\rEIP_reg[24]/NET0131 ,
		_w1109_,
		_w1110_,
		_w1364_
	);
	LUT2 #(
		.INIT('hb)
	) name912 (
		_w1362_,
		_w1364_,
		_w1365_
	);
	LUT4 #(
		.INIT('h1d11)
	) name913 (
		\PhyAddrPointer_reg[30]/NET0131 ,
		_w681_,
		_w1119_,
		_w1137_,
		_w1366_
	);
	LUT4 #(
		.INIT('h028a)
	) name914 (
		\PhyAddrPointer_reg[30]/NET0131 ,
		_w573_,
		_w574_,
		_w605_,
		_w1367_
	);
	LUT2 #(
		.INIT('h1)
	) name915 (
		_w1156_,
		_w1367_,
		_w1368_
	);
	LUT4 #(
		.INIT('h08cc)
	) name916 (
		_w574_,
		_w695_,
		_w1366_,
		_w1368_,
		_w1369_
	);
	LUT3 #(
		.INIT('h6c)
	) name917 (
		\PhyAddrPointer_reg[1]/NET0131 ,
		\PhyAddrPointer_reg[30]/NET0131 ,
		_w1278_,
		_w1370_
	);
	LUT4 #(
		.INIT('h6c00)
	) name918 (
		\PhyAddrPointer_reg[1]/NET0131 ,
		\PhyAddrPointer_reg[30]/NET0131 ,
		_w1278_,
		_w1281_,
		_w1371_
	);
	LUT4 #(
		.INIT('h3f15)
	) name919 (
		\PhyAddrPointer_reg[30]/NET0131 ,
		\rEIP_reg[30]/NET0131 ,
		_w1109_,
		_w1283_,
		_w1372_
	);
	LUT4 #(
		.INIT('hb700)
	) name920 (
		\PhyAddrPointer_reg[30]/NET0131 ,
		_w707_,
		_w1278_,
		_w1372_,
		_w1373_
	);
	LUT2 #(
		.INIT('h4)
	) name921 (
		_w1371_,
		_w1373_,
		_w1374_
	);
	LUT2 #(
		.INIT('hb)
	) name922 (
		_w1369_,
		_w1374_,
		_w1375_
	);
	LUT2 #(
		.INIT('h2)
	) name923 (
		\InstAddrPointer_reg[11]/NET0131 ,
		_w681_,
		_w1376_
	);
	LUT3 #(
		.INIT('h84)
	) name924 (
		_w730_,
		_w844_,
		_w933_,
		_w1377_
	);
	LUT4 #(
		.INIT('h8aa8)
	) name925 (
		_w681_,
		_w844_,
		_w979_,
		_w983_,
		_w1378_
	);
	LUT4 #(
		.INIT('h8a88)
	) name926 (
		_w574_,
		_w1376_,
		_w1377_,
		_w1378_,
		_w1379_
	);
	LUT4 #(
		.INIT('h28a0)
	) name927 (
		_w688_,
		_w1054_,
		_w1060_,
		_w1066_,
		_w1380_
	);
	LUT4 #(
		.INIT('h1300)
	) name928 (
		_w514_,
		_w566_,
		_w569_,
		_w617_,
		_w1381_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name929 (
		\InstAddrPointer_reg[11]/NET0131 ,
		_w611_,
		_w633_,
		_w728_,
		_w1382_
	);
	LUT4 #(
		.INIT('h00f7)
	) name930 (
		_w612_,
		_w730_,
		_w1381_,
		_w1382_,
		_w1383_
	);
	LUT4 #(
		.INIT('hec00)
	) name931 (
		_w514_,
		_w566_,
		_w569_,
		_w730_,
		_w1384_
	);
	LUT3 #(
		.INIT('h08)
	) name932 (
		_w613_,
		_w636_,
		_w1384_,
		_w1385_
	);
	LUT2 #(
		.INIT('h1)
	) name933 (
		_w1383_,
		_w1385_,
		_w1386_
	);
	LUT3 #(
		.INIT('h84)
	) name934 (
		\InstAddrPointer_reg[11]/NET0131 ,
		_w605_,
		_w1059_,
		_w1387_
	);
	LUT2 #(
		.INIT('h1)
	) name935 (
		\InstAddrPointer_reg[11]/NET0131 ,
		_w605_,
		_w1388_
	);
	LUT4 #(
		.INIT('h00c8)
	) name936 (
		_w552_,
		_w576_,
		_w579_,
		_w1388_,
		_w1389_
	);
	LUT3 #(
		.INIT('h08)
	) name937 (
		\InstAddrPointer_reg[11]/NET0131 ,
		_w573_,
		_w605_,
		_w1390_
	);
	LUT2 #(
		.INIT('h8)
	) name938 (
		_w549_,
		_w730_,
		_w1391_
	);
	LUT4 #(
		.INIT('h000b)
	) name939 (
		_w1387_,
		_w1389_,
		_w1390_,
		_w1391_,
		_w1392_
	);
	LUT4 #(
		.INIT('h4f00)
	) name940 (
		_w582_,
		_w595_,
		_w983_,
		_w1392_,
		_w1393_
	);
	LUT3 #(
		.INIT('h10)
	) name941 (
		_w1386_,
		_w1380_,
		_w1393_,
		_w1394_
	);
	LUT4 #(
		.INIT('h3f15)
	) name942 (
		\InstAddrPointer_reg[11]/NET0131 ,
		\rEIP_reg[11]/NET0131 ,
		_w1109_,
		_w1110_,
		_w1395_
	);
	LUT4 #(
		.INIT('h8aff)
	) name943 (
		_w695_,
		_w1379_,
		_w1394_,
		_w1395_,
		_w1396_
	);
	LUT3 #(
		.INIT('h2a)
	) name944 (
		_w986_,
		_w1127_,
		_w1129_,
		_w1397_
	);
	LUT4 #(
		.INIT('hc408)
	) name945 (
		_w736_,
		_w844_,
		_w863_,
		_w867_,
		_w1398_
	);
	LUT4 #(
		.INIT('h00ab)
	) name946 (
		_w844_,
		_w1210_,
		_w1397_,
		_w1398_,
		_w1399_
	);
	LUT4 #(
		.INIT('h08c8)
	) name947 (
		\InstAddrPointer_reg[14]/NET0131 ,
		_w574_,
		_w681_,
		_w1399_,
		_w1400_
	);
	LUT4 #(
		.INIT('h0800)
	) name948 (
		_w1052_,
		_w1066_,
		_w1145_,
		_w1146_,
		_w1401_
	);
	LUT3 #(
		.INIT('h28)
	) name949 (
		_w688_,
		_w1147_,
		_w1401_,
		_w1402_
	);
	LUT2 #(
		.INIT('h2)
	) name950 (
		\InstAddrPointer_reg[14]/NET0131 ,
		_w1220_,
		_w1403_
	);
	LUT2 #(
		.INIT('h4)
	) name951 (
		_w645_,
		_w867_,
		_w1404_
	);
	LUT2 #(
		.INIT('h8)
	) name952 (
		_w606_,
		_w1147_,
		_w1405_
	);
	LUT4 #(
		.INIT('h004f)
	) name953 (
		_w582_,
		_w595_,
		_w986_,
		_w1405_,
		_w1406_
	);
	LUT3 #(
		.INIT('h10)
	) name954 (
		_w1404_,
		_w1403_,
		_w1406_,
		_w1407_
	);
	LUT2 #(
		.INIT('h4)
	) name955 (
		_w1402_,
		_w1407_,
		_w1408_
	);
	LUT4 #(
		.INIT('h3f15)
	) name956 (
		\InstAddrPointer_reg[14]/NET0131 ,
		\rEIP_reg[14]/NET0131 ,
		_w1109_,
		_w1110_,
		_w1409_
	);
	LUT4 #(
		.INIT('h8aff)
	) name957 (
		_w695_,
		_w1400_,
		_w1408_,
		_w1409_,
		_w1410_
	);
	LUT2 #(
		.INIT('h2)
	) name958 (
		\InstAddrPointer_reg[25]/NET0131 ,
		_w681_,
		_w1411_
	);
	LUT3 #(
		.INIT('h6c)
	) name959 (
		\InstAddrPointer_reg[20]/NET0131 ,
		\InstAddrPointer_reg[21]/NET0131 ,
		_w875_,
		_w1412_
	);
	LUT3 #(
		.INIT('h80)
	) name960 (
		_w886_,
		_w1169_,
		_w1412_,
		_w1413_
	);
	LUT4 #(
		.INIT('h6c00)
	) name961 (
		\InstAddrPointer_reg[15]/NET0131 ,
		\InstAddrPointer_reg[16]/NET0131 ,
		_w866_,
		_w932_,
		_w1414_
	);
	LUT3 #(
		.INIT('h80)
	) name962 (
		_w732_,
		_w934_,
		_w1414_,
		_w1415_
	);
	LUT4 #(
		.INIT('hb000)
	) name963 (
		_w927_,
		_w929_,
		_w930_,
		_w1415_,
		_w1416_
	);
	LUT4 #(
		.INIT('h4888)
	) name964 (
		\InstAddrPointer_reg[17]/NET0131 ,
		\InstAddrPointer_reg[20]/NET0131 ,
		_w727_,
		_w871_,
		_w1417_
	);
	LUT3 #(
		.INIT('h80)
	) name965 (
		\InstAddrPointer_reg[19]/NET0131 ,
		_w909_,
		_w1417_,
		_w1418_
	);
	LUT4 #(
		.INIT('h1555)
	) name966 (
		_w883_,
		_w1413_,
		_w1416_,
		_w1418_,
		_w1419_
	);
	LUT3 #(
		.INIT('h80)
	) name967 (
		\InstAddrPointer_reg[25]/NET0131 ,
		_w886_,
		_w1169_,
		_w1420_
	);
	LUT4 #(
		.INIT('h4000)
	) name968 (
		_w863_,
		_w914_,
		_w1168_,
		_w1420_,
		_w1421_
	);
	LUT3 #(
		.INIT('ha8)
	) name969 (
		_w844_,
		_w1419_,
		_w1421_,
		_w1422_
	);
	LUT4 #(
		.INIT('h8aa8)
	) name970 (
		_w681_,
		_w844_,
		_w1009_,
		_w1353_,
		_w1423_
	);
	LUT4 #(
		.INIT('h8a88)
	) name971 (
		_w574_,
		_w1411_,
		_w1422_,
		_w1423_,
		_w1424_
	);
	LUT2 #(
		.INIT('h6)
	) name972 (
		\InstAddrPointer_reg[25]/NET0131 ,
		_w1079_,
		_w1425_
	);
	LUT4 #(
		.INIT('h2a80)
	) name973 (
		_w688_,
		_w1074_,
		_w1086_,
		_w1425_,
		_w1426_
	);
	LUT4 #(
		.INIT('haaa2)
	) name974 (
		\InstAddrPointer_reg[25]/NET0131 ,
		_w1099_,
		_w1195_,
		_w1329_,
		_w1427_
	);
	LUT4 #(
		.INIT('h5040)
	) name975 (
		READY_n_pad,
		_w566_,
		_w611_,
		_w618_,
		_w1428_
	);
	LUT4 #(
		.INIT('h1333)
	) name976 (
		_w514_,
		_w549_,
		_w569_,
		_w612_,
		_w1429_
	);
	LUT3 #(
		.INIT('h8a)
	) name977 (
		_w883_,
		_w1428_,
		_w1429_,
		_w1430_
	);
	LUT2 #(
		.INIT('h8)
	) name978 (
		_w606_,
		_w1425_,
		_w1431_
	);
	LUT4 #(
		.INIT('h004f)
	) name979 (
		_w582_,
		_w595_,
		_w1009_,
		_w1431_,
		_w1432_
	);
	LUT3 #(
		.INIT('h10)
	) name980 (
		_w1430_,
		_w1427_,
		_w1432_,
		_w1433_
	);
	LUT2 #(
		.INIT('h4)
	) name981 (
		_w1426_,
		_w1433_,
		_w1434_
	);
	LUT4 #(
		.INIT('h3f15)
	) name982 (
		\InstAddrPointer_reg[25]/NET0131 ,
		\rEIP_reg[25]/NET0131 ,
		_w1109_,
		_w1110_,
		_w1435_
	);
	LUT4 #(
		.INIT('h8aff)
	) name983 (
		_w695_,
		_w1424_,
		_w1434_,
		_w1435_,
		_w1436_
	);
	LUT2 #(
		.INIT('h2)
	) name984 (
		\PhyAddrPointer_reg[15]/NET0131 ,
		_w681_,
		_w1437_
	);
	LUT4 #(
		.INIT('h00df)
	) name985 (
		_w736_,
		_w863_,
		_w867_,
		_w902_,
		_w1438_
	);
	LUT3 #(
		.INIT('ha8)
	) name986 (
		_w844_,
		_w1114_,
		_w1438_,
		_w1439_
	);
	LUT4 #(
		.INIT('h4015)
	) name987 (
		_w844_,
		_w979_,
		_w987_,
		_w988_,
		_w1440_
	);
	LUT2 #(
		.INIT('h2)
	) name988 (
		_w681_,
		_w1440_,
		_w1441_
	);
	LUT4 #(
		.INIT('h8a88)
	) name989 (
		_w574_,
		_w1437_,
		_w1439_,
		_w1441_,
		_w1442_
	);
	LUT4 #(
		.INIT('h028a)
	) name990 (
		\PhyAddrPointer_reg[15]/NET0131 ,
		_w573_,
		_w574_,
		_w605_,
		_w1443_
	);
	LUT3 #(
		.INIT('h80)
	) name991 (
		_w1054_,
		_w1064_,
		_w1066_,
		_w1444_
	);
	LUT4 #(
		.INIT('h8000)
	) name992 (
		_w1054_,
		_w1064_,
		_w1066_,
		_w1057_,
		_w1445_
	);
	LUT4 #(
		.INIT('h007f)
	) name993 (
		_w1054_,
		_w1064_,
		_w1066_,
		_w1057_,
		_w1446_
	);
	LUT3 #(
		.INIT('h02)
	) name994 (
		_w688_,
		_w1446_,
		_w1445_,
		_w1447_
	);
	LUT4 #(
		.INIT('h0d07)
	) name995 (
		_w688_,
		_w1057_,
		_w1443_,
		_w1444_,
		_w1448_
	);
	LUT4 #(
		.INIT('h8000)
	) name996 (
		\PhyAddrPointer_reg[12]/NET0131 ,
		\PhyAddrPointer_reg[13]/NET0131 ,
		\PhyAddrPointer_reg[1]/NET0131 ,
		_w1263_,
		_w1449_
	);
	LUT3 #(
		.INIT('h6c)
	) name997 (
		\PhyAddrPointer_reg[14]/NET0131 ,
		\PhyAddrPointer_reg[15]/NET0131 ,
		_w1449_,
		_w1450_
	);
	LUT4 #(
		.INIT('h60c0)
	) name998 (
		\PhyAddrPointer_reg[14]/NET0131 ,
		\PhyAddrPointer_reg[15]/NET0131 ,
		_w706_,
		_w1449_,
		_w1451_
	);
	LUT4 #(
		.INIT('h8000)
	) name999 (
		\PhyAddrPointer_reg[12]/NET0131 ,
		\PhyAddrPointer_reg[13]/NET0131 ,
		\PhyAddrPointer_reg[14]/NET0131 ,
		_w1263_,
		_w1452_
	);
	LUT2 #(
		.INIT('h1)
	) name1000 (
		\DataWidth_reg[1]/NET0131 ,
		\PhyAddrPointer_reg[1]/NET0131 ,
		_w1453_
	);
	LUT4 #(
		.INIT('h8848)
	) name1001 (
		\PhyAddrPointer_reg[15]/NET0131 ,
		_w700_,
		_w1452_,
		_w1453_,
		_w1454_
	);
	LUT4 #(
		.INIT('h3f15)
	) name1002 (
		\PhyAddrPointer_reg[15]/NET0131 ,
		\rEIP_reg[15]/NET0131 ,
		_w1109_,
		_w1283_,
		_w1455_
	);
	LUT3 #(
		.INIT('h10)
	) name1003 (
		_w1454_,
		_w1451_,
		_w1455_,
		_w1456_
	);
	LUT4 #(
		.INIT('h8aff)
	) name1004 (
		_w695_,
		_w1442_,
		_w1448_,
		_w1456_,
		_w1457_
	);
	LUT2 #(
		.INIT('h2)
	) name1005 (
		\PhyAddrPointer_reg[23]/NET0131 ,
		_w681_,
		_w1458_
	);
	LUT4 #(
		.INIT('haa20)
	) name1006 (
		_w574_,
		_w1213_,
		_w1215_,
		_w1458_,
		_w1459_
	);
	LUT4 #(
		.INIT('h028a)
	) name1007 (
		\PhyAddrPointer_reg[23]/NET0131 ,
		_w573_,
		_w574_,
		_w605_,
		_w1460_
	);
	LUT3 #(
		.INIT('h0b)
	) name1008 (
		_w1217_,
		_w1219_,
		_w1460_,
		_w1461_
	);
	LUT2 #(
		.INIT('h8)
	) name1009 (
		\PhyAddrPointer_reg[1]/NET0131 ,
		_w1272_,
		_w1462_
	);
	LUT4 #(
		.INIT('h78f0)
	) name1010 (
		\PhyAddrPointer_reg[1]/NET0131 ,
		\PhyAddrPointer_reg[22]/NET0131 ,
		\PhyAddrPointer_reg[23]/NET0131 ,
		_w1272_,
		_w1463_
	);
	LUT2 #(
		.INIT('h8)
	) name1011 (
		_w1281_,
		_w1463_,
		_w1464_
	);
	LUT4 #(
		.INIT('hc444)
	) name1012 (
		_w707_,
		_w1283_,
		_w1272_,
		_w1273_,
		_w1465_
	);
	LUT2 #(
		.INIT('h8)
	) name1013 (
		\PhyAddrPointer_reg[22]/NET0131 ,
		_w1272_,
		_w1466_
	);
	LUT4 #(
		.INIT('h2000)
	) name1014 (
		\PhyAddrPointer_reg[22]/NET0131 ,
		\PhyAddrPointer_reg[23]/NET0131 ,
		_w707_,
		_w1272_,
		_w1467_
	);
	LUT4 #(
		.INIT('h0031)
	) name1015 (
		\PhyAddrPointer_reg[23]/NET0131 ,
		_w1228_,
		_w1465_,
		_w1467_,
		_w1468_
	);
	LUT2 #(
		.INIT('h4)
	) name1016 (
		_w1464_,
		_w1468_,
		_w1469_
	);
	LUT4 #(
		.INIT('h8aff)
	) name1017 (
		_w695_,
		_w1459_,
		_w1461_,
		_w1469_,
		_w1470_
	);
	LUT4 #(
		.INIT('h111d)
	) name1018 (
		\PhyAddrPointer_reg[27]/NET0131 ,
		_w681_,
		_w1232_,
		_w1235_,
		_w1471_
	);
	LUT4 #(
		.INIT('h028a)
	) name1019 (
		\PhyAddrPointer_reg[27]/NET0131 ,
		_w573_,
		_w574_,
		_w605_,
		_w1472_
	);
	LUT3 #(
		.INIT('h0b)
	) name1020 (
		_w1237_,
		_w1239_,
		_w1472_,
		_w1473_
	);
	LUT4 #(
		.INIT('h08cc)
	) name1021 (
		_w574_,
		_w695_,
		_w1471_,
		_w1473_,
		_w1474_
	);
	LUT4 #(
		.INIT('h8000)
	) name1022 (
		\PhyAddrPointer_reg[1]/NET0131 ,
		\PhyAddrPointer_reg[24]/NET0131 ,
		_w1272_,
		_w1273_,
		_w1475_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name1023 (
		\PhyAddrPointer_reg[1]/NET0131 ,
		\PhyAddrPointer_reg[27]/NET0131 ,
		_w1274_,
		_w1275_,
		_w1476_
	);
	LUT4 #(
		.INIT('h3f15)
	) name1024 (
		\PhyAddrPointer_reg[27]/NET0131 ,
		\rEIP_reg[27]/NET0131 ,
		_w1109_,
		_w1283_,
		_w1477_
	);
	LUT4 #(
		.INIT('hb700)
	) name1025 (
		\PhyAddrPointer_reg[27]/NET0131 ,
		_w707_,
		_w1276_,
		_w1477_,
		_w1478_
	);
	LUT3 #(
		.INIT('h70)
	) name1026 (
		_w1281_,
		_w1476_,
		_w1478_,
		_w1479_
	);
	LUT2 #(
		.INIT('hb)
	) name1027 (
		_w1474_,
		_w1479_,
		_w1480_
	);
	LUT2 #(
		.INIT('h2)
	) name1028 (
		\PhyAddrPointer_reg[28]/NET0131 ,
		_w681_,
		_w1481_
	);
	LUT4 #(
		.INIT('haa20)
	) name1029 (
		_w574_,
		_w1175_,
		_w1180_,
		_w1481_,
		_w1482_
	);
	LUT4 #(
		.INIT('h028a)
	) name1030 (
		\PhyAddrPointer_reg[28]/NET0131 ,
		_w573_,
		_w574_,
		_w605_,
		_w1483_
	);
	LUT2 #(
		.INIT('h1)
	) name1031 (
		_w1194_,
		_w1483_,
		_w1484_
	);
	LUT4 #(
		.INIT('h78f0)
	) name1032 (
		\PhyAddrPointer_reg[1]/NET0131 ,
		\PhyAddrPointer_reg[27]/NET0131 ,
		\PhyAddrPointer_reg[28]/NET0131 ,
		_w1276_,
		_w1485_
	);
	LUT4 #(
		.INIT('h60c0)
	) name1033 (
		\PhyAddrPointer_reg[27]/NET0131 ,
		\PhyAddrPointer_reg[28]/NET0131 ,
		_w707_,
		_w1276_,
		_w1486_
	);
	LUT4 #(
		.INIT('h3f15)
	) name1034 (
		\PhyAddrPointer_reg[28]/NET0131 ,
		\rEIP_reg[28]/NET0131 ,
		_w1109_,
		_w1283_,
		_w1487_
	);
	LUT4 #(
		.INIT('h1300)
	) name1035 (
		_w1281_,
		_w1486_,
		_w1485_,
		_w1487_,
		_w1488_
	);
	LUT4 #(
		.INIT('h8aff)
	) name1036 (
		_w695_,
		_w1482_,
		_w1484_,
		_w1488_,
		_w1489_
	);
	LUT3 #(
		.INIT('h80)
	) name1037 (
		\InstAddrPointer_reg[28]/NET0131 ,
		_w891_,
		_w884_,
		_w1490_
	);
	LUT2 #(
		.INIT('h8)
	) name1038 (
		_w1413_,
		_w1490_,
		_w1491_
	);
	LUT4 #(
		.INIT('h2888)
	) name1039 (
		_w844_,
		_w897_,
		_w1309_,
		_w1491_,
		_w1492_
	);
	LUT4 #(
		.INIT('h8010)
	) name1040 (
		\InstAddrPointer_reg[27]/NET0131 ,
		\InstAddrPointer_reg[28]/NET0131 ,
		_w1011_,
		_w1015_,
		_w1493_
	);
	LUT4 #(
		.INIT('h8000)
	) name1041 (
		_w1349_,
		_w1351_,
		_w1352_,
		_w1493_,
		_w1494_
	);
	LUT3 #(
		.INIT('hbe)
	) name1042 (
		_w844_,
		_w1019_,
		_w1494_,
		_w1495_
	);
	LUT4 #(
		.INIT('h1d11)
	) name1043 (
		\PhyAddrPointer_reg[29]/NET0131 ,
		_w681_,
		_w1492_,
		_w1495_,
		_w1496_
	);
	LUT4 #(
		.INIT('h028a)
	) name1044 (
		\PhyAddrPointer_reg[29]/NET0131 ,
		_w573_,
		_w574_,
		_w605_,
		_w1497_
	);
	LUT3 #(
		.INIT('h13)
	) name1045 (
		_w1090_,
		_w1089_,
		_w1238_,
		_w1498_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name1046 (
		\InstAddrPointer_reg[29]/NET0131 ,
		_w688_,
		_w1090_,
		_w1238_,
		_w1499_
	);
	LUT3 #(
		.INIT('h45)
	) name1047 (
		_w1497_,
		_w1498_,
		_w1499_,
		_w1500_
	);
	LUT4 #(
		.INIT('h08cc)
	) name1048 (
		_w574_,
		_w695_,
		_w1496_,
		_w1500_,
		_w1501_
	);
	LUT3 #(
		.INIT('h6c)
	) name1049 (
		\PhyAddrPointer_reg[1]/NET0131 ,
		\PhyAddrPointer_reg[29]/NET0131 ,
		_w1277_,
		_w1502_
	);
	LUT4 #(
		.INIT('h60c0)
	) name1050 (
		\PhyAddrPointer_reg[1]/NET0131 ,
		\PhyAddrPointer_reg[29]/NET0131 ,
		_w706_,
		_w1277_,
		_w1503_
	);
	LUT4 #(
		.INIT('h0080)
	) name1051 (
		\PhyAddrPointer_reg[27]/NET0131 ,
		\PhyAddrPointer_reg[28]/NET0131 ,
		_w1276_,
		_w1453_,
		_w1504_
	);
	LUT4 #(
		.INIT('h3f15)
	) name1052 (
		\PhyAddrPointer_reg[29]/NET0131 ,
		\rEIP_reg[29]/NET0131 ,
		_w1109_,
		_w1283_,
		_w1505_
	);
	LUT4 #(
		.INIT('hb700)
	) name1053 (
		\PhyAddrPointer_reg[29]/NET0131 ,
		_w700_,
		_w1504_,
		_w1505_,
		_w1506_
	);
	LUT2 #(
		.INIT('h4)
	) name1054 (
		_w1503_,
		_w1506_,
		_w1507_
	);
	LUT2 #(
		.INIT('hb)
	) name1055 (
		_w1501_,
		_w1507_,
		_w1508_
	);
	LUT2 #(
		.INIT('h2)
	) name1056 (
		\InstAddrPointer_reg[8]/NET0131 ,
		_w681_,
		_w1509_
	);
	LUT3 #(
		.INIT('h48)
	) name1057 (
		_w733_,
		_w844_,
		_w863_,
		_w1510_
	);
	LUT4 #(
		.INIT('h8aa8)
	) name1058 (
		_w681_,
		_w844_,
		_w976_,
		_w1126_,
		_w1511_
	);
	LUT4 #(
		.INIT('h8a88)
	) name1059 (
		_w574_,
		_w1509_,
		_w1510_,
		_w1511_,
		_w1512_
	);
	LUT3 #(
		.INIT('h82)
	) name1060 (
		_w688_,
		_w1052_,
		_w1145_,
		_w1513_
	);
	LUT4 #(
		.INIT('h8088)
	) name1061 (
		READY_n_pad,
		_w611_,
		_w618_,
		_w619_,
		_w1514_
	);
	LUT3 #(
		.INIT('ha2)
	) name1062 (
		\InstAddrPointer_reg[8]/NET0131 ,
		_w1197_,
		_w1514_,
		_w1515_
	);
	LUT2 #(
		.INIT('h4)
	) name1063 (
		_w620_,
		_w733_,
		_w1516_
	);
	LUT2 #(
		.INIT('h8)
	) name1064 (
		_w606_,
		_w1052_,
		_w1517_
	);
	LUT4 #(
		.INIT('h004f)
	) name1065 (
		_w582_,
		_w595_,
		_w976_,
		_w1517_,
		_w1518_
	);
	LUT4 #(
		.INIT('h0100)
	) name1066 (
		_w1515_,
		_w1513_,
		_w1516_,
		_w1518_,
		_w1519_
	);
	LUT4 #(
		.INIT('h3f15)
	) name1067 (
		\InstAddrPointer_reg[8]/NET0131 ,
		\rEIP_reg[8]/NET0131 ,
		_w1109_,
		_w1110_,
		_w1520_
	);
	LUT4 #(
		.INIT('h8aff)
	) name1068 (
		_w695_,
		_w1512_,
		_w1519_,
		_w1520_,
		_w1521_
	);
	LUT2 #(
		.INIT('h2)
	) name1069 (
		\InstAddrPointer_reg[12]/NET0131 ,
		_w681_,
		_w1522_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name1070 (
		\InstAddrPointer_reg[12]/NET0131 ,
		\InstAddrPointer_reg[9]/NET0131 ,
		_w727_,
		_w729_,
		_w1523_
	);
	LUT3 #(
		.INIT('h6a)
	) name1071 (
		\InstAddrPointer_reg[10]/NET0131 ,
		\InstAddrPointer_reg[9]/NET0131 ,
		_w727_,
		_w1524_
	);
	LUT4 #(
		.INIT('h0800)
	) name1072 (
		\InstAddrPointer_reg[11]/NET0131 ,
		_w734_,
		_w863_,
		_w1524_,
		_w1525_
	);
	LUT3 #(
		.INIT('h82)
	) name1073 (
		_w844_,
		_w1523_,
		_w1525_,
		_w1526_
	);
	LUT3 #(
		.INIT('h81)
	) name1074 (
		\InstAddrPointer_reg[10]/NET0131 ,
		\InstAddrPointer_reg[11]/NET0131 ,
		_w970_,
		_w1527_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name1075 (
		_w973_,
		_w982_,
		_w1127_,
		_w1527_,
		_w1528_
	);
	LUT3 #(
		.INIT('h15)
	) name1076 (
		_w844_,
		_w1127_,
		_w1128_,
		_w1529_
	);
	LUT3 #(
		.INIT('h8a)
	) name1077 (
		_w681_,
		_w1528_,
		_w1529_,
		_w1530_
	);
	LUT4 #(
		.INIT('h8a88)
	) name1078 (
		_w574_,
		_w1522_,
		_w1526_,
		_w1530_,
		_w1531_
	);
	LUT4 #(
		.INIT('h82a0)
	) name1079 (
		_w688_,
		_w1145_,
		_w1184_,
		_w1183_,
		_w1532_
	);
	LUT4 #(
		.INIT('ha8a0)
	) name1080 (
		\InstAddrPointer_reg[12]/NET0131 ,
		_w514_,
		_w566_,
		_w569_,
		_w1533_
	);
	LUT3 #(
		.INIT('hc4)
	) name1081 (
		_w645_,
		_w1523_,
		_w1533_,
		_w1534_
	);
	LUT3 #(
		.INIT('hb0)
	) name1082 (
		_w582_,
		_w595_,
		_w982_,
		_w1535_
	);
	LUT4 #(
		.INIT('haaa2)
	) name1083 (
		\InstAddrPointer_reg[12]/NET0131 ,
		_w636_,
		_w683_,
		_w1096_,
		_w1536_
	);
	LUT2 #(
		.INIT('h2)
	) name1084 (
		_w605_,
		_w1184_,
		_w1537_
	);
	LUT2 #(
		.INIT('h1)
	) name1085 (
		\InstAddrPointer_reg[12]/NET0131 ,
		_w605_,
		_w1538_
	);
	LUT4 #(
		.INIT('h00c8)
	) name1086 (
		_w552_,
		_w576_,
		_w579_,
		_w1538_,
		_w1539_
	);
	LUT2 #(
		.INIT('h4)
	) name1087 (
		_w1537_,
		_w1539_,
		_w1540_
	);
	LUT2 #(
		.INIT('h1)
	) name1088 (
		_w1536_,
		_w1540_,
		_w1541_
	);
	LUT4 #(
		.INIT('h0100)
	) name1089 (
		_w1532_,
		_w1535_,
		_w1534_,
		_w1541_,
		_w1542_
	);
	LUT4 #(
		.INIT('h3f15)
	) name1090 (
		\InstAddrPointer_reg[12]/NET0131 ,
		\rEIP_reg[12]/NET0131 ,
		_w1109_,
		_w1110_,
		_w1543_
	);
	LUT4 #(
		.INIT('h8aff)
	) name1091 (
		_w695_,
		_w1531_,
		_w1542_,
		_w1543_,
		_w1544_
	);
	LUT2 #(
		.INIT('h2)
	) name1092 (
		\PhyAddrPointer_reg[11]/NET0131 ,
		_w681_,
		_w1545_
	);
	LUT4 #(
		.INIT('haa20)
	) name1093 (
		_w574_,
		_w1377_,
		_w1378_,
		_w1545_,
		_w1546_
	);
	LUT4 #(
		.INIT('h028a)
	) name1094 (
		\PhyAddrPointer_reg[11]/NET0131 ,
		_w573_,
		_w574_,
		_w605_,
		_w1547_
	);
	LUT2 #(
		.INIT('h1)
	) name1095 (
		_w1380_,
		_w1547_,
		_w1548_
	);
	LUT4 #(
		.INIT('h8000)
	) name1096 (
		\PhyAddrPointer_reg[10]/NET0131 ,
		\PhyAddrPointer_reg[1]/NET0131 ,
		\PhyAddrPointer_reg[9]/NET0131 ,
		_w1261_,
		_w1549_
	);
	LUT3 #(
		.INIT('h6a)
	) name1097 (
		\PhyAddrPointer_reg[11]/NET0131 ,
		\PhyAddrPointer_reg[1]/NET0131 ,
		_w1262_,
		_w1550_
	);
	LUT4 #(
		.INIT('h6a00)
	) name1098 (
		\PhyAddrPointer_reg[11]/NET0131 ,
		\PhyAddrPointer_reg[1]/NET0131 ,
		_w1262_,
		_w1281_,
		_w1551_
	);
	LUT4 #(
		.INIT('h3f15)
	) name1099 (
		\PhyAddrPointer_reg[11]/NET0131 ,
		\rEIP_reg[11]/NET0131 ,
		_w1109_,
		_w1283_,
		_w1552_
	);
	LUT4 #(
		.INIT('hb700)
	) name1100 (
		\PhyAddrPointer_reg[11]/NET0131 ,
		_w707_,
		_w1262_,
		_w1552_,
		_w1553_
	);
	LUT2 #(
		.INIT('h4)
	) name1101 (
		_w1551_,
		_w1553_,
		_w1554_
	);
	LUT4 #(
		.INIT('h8aff)
	) name1102 (
		_w695_,
		_w1546_,
		_w1548_,
		_w1554_,
		_w1555_
	);
	LUT4 #(
		.INIT('h08c8)
	) name1103 (
		\PhyAddrPointer_reg[14]/NET0131 ,
		_w574_,
		_w681_,
		_w1399_,
		_w1556_
	);
	LUT4 #(
		.INIT('h028a)
	) name1104 (
		\PhyAddrPointer_reg[14]/NET0131 ,
		_w573_,
		_w574_,
		_w605_,
		_w1557_
	);
	LUT4 #(
		.INIT('h00d7)
	) name1105 (
		_w688_,
		_w1147_,
		_w1401_,
		_w1557_,
		_w1558_
	);
	LUT2 #(
		.INIT('h6)
	) name1106 (
		\PhyAddrPointer_reg[14]/NET0131 ,
		_w1449_,
		_w1559_
	);
	LUT3 #(
		.INIT('h48)
	) name1107 (
		\PhyAddrPointer_reg[14]/NET0131 ,
		_w1281_,
		_w1449_,
		_w1560_
	);
	LUT4 #(
		.INIT('h3f15)
	) name1108 (
		\PhyAddrPointer_reg[14]/NET0131 ,
		\rEIP_reg[14]/NET0131 ,
		_w1109_,
		_w1283_,
		_w1561_
	);
	LUT4 #(
		.INIT('hb700)
	) name1109 (
		\PhyAddrPointer_reg[14]/NET0131 ,
		_w707_,
		_w1264_,
		_w1561_,
		_w1562_
	);
	LUT2 #(
		.INIT('h4)
	) name1110 (
		_w1560_,
		_w1562_,
		_w1563_
	);
	LUT4 #(
		.INIT('h8aff)
	) name1111 (
		_w695_,
		_w1556_,
		_w1558_,
		_w1563_,
		_w1564_
	);
	LUT4 #(
		.INIT('h111d)
	) name1112 (
		\PhyAddrPointer_reg[19]/NET0131 ,
		_w681_,
		_w1290_,
		_w1292_,
		_w1565_
	);
	LUT4 #(
		.INIT('h028a)
	) name1113 (
		\PhyAddrPointer_reg[19]/NET0131 ,
		_w573_,
		_w574_,
		_w605_,
		_w1566_
	);
	LUT4 #(
		.INIT('h001f)
	) name1114 (
		_w1294_,
		_w1295_,
		_w1296_,
		_w1566_,
		_w1567_
	);
	LUT4 #(
		.INIT('h08cc)
	) name1115 (
		_w574_,
		_w695_,
		_w1565_,
		_w1567_,
		_w1568_
	);
	LUT4 #(
		.INIT('h8000)
	) name1116 (
		\PhyAddrPointer_reg[12]/NET0131 ,
		\PhyAddrPointer_reg[13]/NET0131 ,
		_w1263_,
		_w1267_,
		_w1569_
	);
	LUT4 #(
		.INIT('h8000)
	) name1117 (
		\PhyAddrPointer_reg[18]/NET0131 ,
		\PhyAddrPointer_reg[19]/NET0131 ,
		\PhyAddrPointer_reg[1]/NET0131 ,
		_w1569_,
		_w1570_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name1118 (
		\PhyAddrPointer_reg[18]/NET0131 ,
		\PhyAddrPointer_reg[19]/NET0131 ,
		\PhyAddrPointer_reg[1]/NET0131 ,
		_w1569_,
		_w1571_
	);
	LUT2 #(
		.INIT('h8)
	) name1119 (
		_w1281_,
		_w1571_,
		_w1572_
	);
	LUT4 #(
		.INIT('hb030)
	) name1120 (
		\PhyAddrPointer_reg[18]/NET0131 ,
		_w707_,
		_w1283_,
		_w1569_,
		_w1573_
	);
	LUT3 #(
		.INIT('h20)
	) name1121 (
		\DataWidth_reg[1]/NET0131 ,
		\PhyAddrPointer_reg[19]/NET0131 ,
		_w700_,
		_w1574_
	);
	LUT4 #(
		.INIT('h1333)
	) name1122 (
		\PhyAddrPointer_reg[18]/NET0131 ,
		_w1305_,
		_w1569_,
		_w1574_,
		_w1575_
	);
	LUT3 #(
		.INIT('hd0)
	) name1123 (
		\PhyAddrPointer_reg[19]/NET0131 ,
		_w1573_,
		_w1575_,
		_w1576_
	);
	LUT2 #(
		.INIT('h4)
	) name1124 (
		_w1572_,
		_w1576_,
		_w1577_
	);
	LUT2 #(
		.INIT('hb)
	) name1125 (
		_w1568_,
		_w1577_,
		_w1578_
	);
	LUT4 #(
		.INIT('hddd1)
	) name1126 (
		\PhyAddrPointer_reg[20]/NET0131 ,
		_w681_,
		_w1310_,
		_w1308_,
		_w1579_
	);
	LUT4 #(
		.INIT('h028a)
	) name1127 (
		\PhyAddrPointer_reg[20]/NET0131 ,
		_w573_,
		_w574_,
		_w605_,
		_w1580_
	);
	LUT4 #(
		.INIT('h00d7)
	) name1128 (
		_w688_,
		_w1072_,
		_w1190_,
		_w1580_,
		_w1581_
	);
	LUT4 #(
		.INIT('h08cc)
	) name1129 (
		_w574_,
		_w695_,
		_w1579_,
		_w1581_,
		_w1582_
	);
	LUT3 #(
		.INIT('h80)
	) name1130 (
		\PhyAddrPointer_reg[1]/NET0131 ,
		_w1269_,
		_w1569_,
		_w1583_
	);
	LUT3 #(
		.INIT('h0e)
	) name1131 (
		\PhyAddrPointer_reg[20]/NET0131 ,
		_w1570_,
		_w1583_,
		_w1584_
	);
	LUT4 #(
		.INIT('h00c8)
	) name1132 (
		\PhyAddrPointer_reg[20]/NET0131 ,
		_w706_,
		_w1570_,
		_w1583_,
		_w1585_
	);
	LUT3 #(
		.INIT('hc8)
	) name1133 (
		\DataWidth_reg[1]/NET0131 ,
		\PhyAddrPointer_reg[19]/NET0131 ,
		\PhyAddrPointer_reg[1]/NET0131 ,
		_w1586_
	);
	LUT4 #(
		.INIT('h1333)
	) name1134 (
		\PhyAddrPointer_reg[18]/NET0131 ,
		\PhyAddrPointer_reg[20]/NET0131 ,
		_w1569_,
		_w1586_,
		_w1587_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name1135 (
		_w700_,
		_w1269_,
		_w1453_,
		_w1569_,
		_w1588_
	);
	LUT4 #(
		.INIT('h3f15)
	) name1136 (
		\PhyAddrPointer_reg[20]/NET0131 ,
		\rEIP_reg[20]/NET0131 ,
		_w1109_,
		_w1283_,
		_w1589_
	);
	LUT3 #(
		.INIT('hb0)
	) name1137 (
		_w1587_,
		_w1588_,
		_w1589_,
		_w1590_
	);
	LUT2 #(
		.INIT('h4)
	) name1138 (
		_w1585_,
		_w1590_,
		_w1591_
	);
	LUT2 #(
		.INIT('hb)
	) name1139 (
		_w1582_,
		_w1591_,
		_w1592_
	);
	LUT2 #(
		.INIT('h2)
	) name1140 (
		\PhyAddrPointer_reg[22]/NET0131 ,
		_w681_,
		_w1593_
	);
	LUT4 #(
		.INIT('haa20)
	) name1141 (
		_w574_,
		_w1324_,
		_w1326_,
		_w1593_,
		_w1594_
	);
	LUT4 #(
		.INIT('h028a)
	) name1142 (
		\PhyAddrPointer_reg[22]/NET0131 ,
		_w573_,
		_w574_,
		_w605_,
		_w1595_
	);
	LUT4 #(
		.INIT('h00d7)
	) name1143 (
		_w688_,
		_w1083_,
		_w1155_,
		_w1595_,
		_w1596_
	);
	LUT3 #(
		.INIT('h6c)
	) name1144 (
		\PhyAddrPointer_reg[1]/NET0131 ,
		\PhyAddrPointer_reg[22]/NET0131 ,
		_w1272_,
		_w1597_
	);
	LUT4 #(
		.INIT('h60c0)
	) name1145 (
		\PhyAddrPointer_reg[1]/NET0131 ,
		\PhyAddrPointer_reg[22]/NET0131 ,
		_w706_,
		_w1272_,
		_w1598_
	);
	LUT4 #(
		.INIT('h8848)
	) name1146 (
		\PhyAddrPointer_reg[22]/NET0131 ,
		_w700_,
		_w1272_,
		_w1453_,
		_w1599_
	);
	LUT4 #(
		.INIT('h3f15)
	) name1147 (
		\PhyAddrPointer_reg[22]/NET0131 ,
		\rEIP_reg[22]/NET0131 ,
		_w1109_,
		_w1283_,
		_w1600_
	);
	LUT3 #(
		.INIT('h10)
	) name1148 (
		_w1599_,
		_w1598_,
		_w1600_,
		_w1601_
	);
	LUT4 #(
		.INIT('h8aff)
	) name1149 (
		_w695_,
		_w1594_,
		_w1596_,
		_w1601_,
		_w1602_
	);
	LUT2 #(
		.INIT('h2)
	) name1150 (
		\PhyAddrPointer_reg[24]/NET0131 ,
		_w681_,
		_w1603_
	);
	LUT4 #(
		.INIT('haa20)
	) name1151 (
		_w574_,
		_w1343_,
		_w1355_,
		_w1603_,
		_w1604_
	);
	LUT4 #(
		.INIT('h028a)
	) name1152 (
		\PhyAddrPointer_reg[24]/NET0131 ,
		_w573_,
		_w574_,
		_w605_,
		_w1605_
	);
	LUT3 #(
		.INIT('h0b)
	) name1153 (
		_w1338_,
		_w1339_,
		_w1605_,
		_w1606_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name1154 (
		\PhyAddrPointer_reg[1]/NET0131 ,
		\PhyAddrPointer_reg[24]/NET0131 ,
		_w1272_,
		_w1273_,
		_w1607_
	);
	LUT2 #(
		.INIT('h8)
	) name1155 (
		_w1281_,
		_w1607_,
		_w1608_
	);
	LUT3 #(
		.INIT('h20)
	) name1156 (
		\DataWidth_reg[1]/NET0131 ,
		\PhyAddrPointer_reg[24]/NET0131 ,
		_w700_,
		_w1609_
	);
	LUT4 #(
		.INIT('h070f)
	) name1157 (
		_w1272_,
		_w1273_,
		_w1363_,
		_w1609_,
		_w1610_
	);
	LUT3 #(
		.INIT('hd0)
	) name1158 (
		\PhyAddrPointer_reg[24]/NET0131 ,
		_w1465_,
		_w1610_,
		_w1611_
	);
	LUT2 #(
		.INIT('h4)
	) name1159 (
		_w1608_,
		_w1611_,
		_w1612_
	);
	LUT4 #(
		.INIT('h8aff)
	) name1160 (
		_w695_,
		_w1604_,
		_w1606_,
		_w1612_,
		_w1613_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name1161 (
		_w844_,
		_w888_,
		_w933_,
		_w936_,
		_w1614_
	);
	LUT3 #(
		.INIT('he0)
	) name1162 (
		_w882_,
		_w1421_,
		_w1614_,
		_w1615_
	);
	LUT4 #(
		.INIT('h4000)
	) name1163 (
		_w1010_,
		_w1127_,
		_w1129_,
		_w1134_,
		_w1616_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name1164 (
		_w1010_,
		_w1127_,
		_w1129_,
		_w1134_,
		_w1617_
	);
	LUT3 #(
		.INIT('h01)
	) name1165 (
		_w844_,
		_w1617_,
		_w1616_,
		_w1618_
	);
	LUT4 #(
		.INIT('h111d)
	) name1166 (
		\PhyAddrPointer_reg[26]/NET0131 ,
		_w681_,
		_w1615_,
		_w1618_,
		_w1619_
	);
	LUT4 #(
		.INIT('h028a)
	) name1167 (
		\PhyAddrPointer_reg[26]/NET0131 ,
		_w573_,
		_w574_,
		_w605_,
		_w1620_
	);
	LUT4 #(
		.INIT('h2888)
	) name1168 (
		_w688_,
		_w1081_,
		_w1087_,
		_w1155_,
		_w1621_
	);
	LUT2 #(
		.INIT('h1)
	) name1169 (
		_w1620_,
		_w1621_,
		_w1622_
	);
	LUT4 #(
		.INIT('h08cc)
	) name1170 (
		_w574_,
		_w695_,
		_w1619_,
		_w1622_,
		_w1623_
	);
	LUT4 #(
		.INIT('h0080)
	) name1171 (
		\PhyAddrPointer_reg[24]/NET0131 ,
		_w1272_,
		_w1273_,
		_w1453_,
		_w1624_
	);
	LUT4 #(
		.INIT('hb030)
	) name1172 (
		\PhyAddrPointer_reg[25]/NET0131 ,
		_w700_,
		_w1283_,
		_w1624_,
		_w1625_
	);
	LUT3 #(
		.INIT('h6c)
	) name1173 (
		\PhyAddrPointer_reg[25]/NET0131 ,
		\PhyAddrPointer_reg[26]/NET0131 ,
		_w1475_,
		_w1626_
	);
	LUT4 #(
		.INIT('h60c0)
	) name1174 (
		\PhyAddrPointer_reg[25]/NET0131 ,
		\PhyAddrPointer_reg[26]/NET0131 ,
		_w706_,
		_w1475_,
		_w1627_
	);
	LUT2 #(
		.INIT('h4)
	) name1175 (
		\PhyAddrPointer_reg[26]/NET0131 ,
		_w700_,
		_w1628_
	);
	LUT2 #(
		.INIT('h8)
	) name1176 (
		\rEIP_reg[26]/NET0131 ,
		_w1109_,
		_w1629_
	);
	LUT4 #(
		.INIT('h007f)
	) name1177 (
		\PhyAddrPointer_reg[25]/NET0131 ,
		_w1624_,
		_w1628_,
		_w1629_,
		_w1630_
	);
	LUT4 #(
		.INIT('h3100)
	) name1178 (
		\PhyAddrPointer_reg[26]/NET0131 ,
		_w1627_,
		_w1625_,
		_w1630_,
		_w1631_
	);
	LUT2 #(
		.INIT('hb)
	) name1179 (
		_w1623_,
		_w1631_,
		_w1632_
	);
	LUT2 #(
		.INIT('h2)
	) name1180 (
		\InstAddrPointer_reg[9]/NET0131 ,
		_w681_,
		_w1633_
	);
	LUT4 #(
		.INIT('h4fb0)
	) name1181 (
		_w927_,
		_w929_,
		_w930_,
		_w931_,
		_w1634_
	);
	LUT4 #(
		.INIT('h65aa)
	) name1182 (
		_w973_,
		_w1345_,
		_w1346_,
		_w1348_,
		_w1635_
	);
	LUT4 #(
		.INIT('ha820)
	) name1183 (
		_w681_,
		_w844_,
		_w1635_,
		_w1634_,
		_w1636_
	);
	LUT3 #(
		.INIT('ha8)
	) name1184 (
		_w574_,
		_w1633_,
		_w1636_,
		_w1637_
	);
	LUT3 #(
		.INIT('h28)
	) name1185 (
		_w688_,
		_w1054_,
		_w1065_,
		_w1638_
	);
	LUT2 #(
		.INIT('h4)
	) name1186 (
		_w620_,
		_w931_,
		_w1639_
	);
	LUT3 #(
		.INIT('h2a)
	) name1187 (
		\InstAddrPointer_reg[9]/NET0131 ,
		_w624_,
		_w684_,
		_w1640_
	);
	LUT2 #(
		.INIT('h8)
	) name1188 (
		_w606_,
		_w1065_,
		_w1641_
	);
	LUT4 #(
		.INIT('h004f)
	) name1189 (
		_w582_,
		_w595_,
		_w973_,
		_w1641_,
		_w1642_
	);
	LUT4 #(
		.INIT('h0100)
	) name1190 (
		_w1640_,
		_w1638_,
		_w1639_,
		_w1642_,
		_w1643_
	);
	LUT4 #(
		.INIT('h3f15)
	) name1191 (
		\InstAddrPointer_reg[9]/NET0131 ,
		\rEIP_reg[9]/NET0131 ,
		_w1109_,
		_w1110_,
		_w1644_
	);
	LUT4 #(
		.INIT('h8aff)
	) name1192 (
		_w695_,
		_w1637_,
		_w1643_,
		_w1644_,
		_w1645_
	);
	LUT2 #(
		.INIT('h2)
	) name1193 (
		\PhyAddrPointer_reg[16]/NET0131 ,
		_w681_,
		_w1646_
	);
	LUT4 #(
		.INIT('h82a0)
	) name1194 (
		_w844_,
		_w863_,
		_w904_,
		_w1113_,
		_w1647_
	);
	LUT4 #(
		.INIT('h8aa8)
	) name1195 (
		_w681_,
		_w844_,
		_w991_,
		_w1177_,
		_w1648_
	);
	LUT4 #(
		.INIT('h8a88)
	) name1196 (
		_w574_,
		_w1646_,
		_w1647_,
		_w1648_,
		_w1649_
	);
	LUT4 #(
		.INIT('h4000)
	) name1197 (
		_w1145_,
		_w1183_,
		_w1185_,
		_w1188_,
		_w1650_
	);
	LUT4 #(
		.INIT('h00bf)
	) name1198 (
		_w1145_,
		_w1183_,
		_w1185_,
		_w1188_,
		_w1651_
	);
	LUT3 #(
		.INIT('h02)
	) name1199 (
		_w688_,
		_w1651_,
		_w1650_,
		_w1652_
	);
	LUT4 #(
		.INIT('h028a)
	) name1200 (
		\PhyAddrPointer_reg[16]/NET0131 ,
		_w573_,
		_w574_,
		_w605_,
		_w1653_
	);
	LUT4 #(
		.INIT('h00d7)
	) name1201 (
		_w688_,
		_w1186_,
		_w1188_,
		_w1653_,
		_w1654_
	);
	LUT3 #(
		.INIT('h15)
	) name1202 (
		\PhyAddrPointer_reg[16]/NET0131 ,
		_w1265_,
		_w1449_,
		_w1655_
	);
	LUT4 #(
		.INIT('h8000)
	) name1203 (
		\PhyAddrPointer_reg[12]/NET0131 ,
		\PhyAddrPointer_reg[13]/NET0131 ,
		_w1263_,
		_w1266_,
		_w1656_
	);
	LUT2 #(
		.INIT('h8)
	) name1204 (
		\PhyAddrPointer_reg[1]/NET0131 ,
		_w1656_,
		_w1657_
	);
	LUT2 #(
		.INIT('h1)
	) name1205 (
		_w1655_,
		_w1657_,
		_w1658_
	);
	LUT3 #(
		.INIT('h02)
	) name1206 (
		_w1281_,
		_w1655_,
		_w1657_,
		_w1659_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name1207 (
		\PhyAddrPointer_reg[16]/NET0131 ,
		_w707_,
		_w1283_,
		_w1656_,
		_w1660_
	);
	LUT4 #(
		.INIT('h0080)
	) name1208 (
		\PhyAddrPointer_reg[15]/NET0131 ,
		_w707_,
		_w1452_,
		_w1656_,
		_w1661_
	);
	LUT2 #(
		.INIT('h8)
	) name1209 (
		\rEIP_reg[16]/NET0131 ,
		_w1109_,
		_w1662_
	);
	LUT3 #(
		.INIT('h01)
	) name1210 (
		_w1661_,
		_w1660_,
		_w1662_,
		_w1663_
	);
	LUT2 #(
		.INIT('h4)
	) name1211 (
		_w1659_,
		_w1663_,
		_w1664_
	);
	LUT4 #(
		.INIT('h8aff)
	) name1212 (
		_w695_,
		_w1649_,
		_w1654_,
		_w1664_,
		_w1665_
	);
	LUT2 #(
		.INIT('h2)
	) name1213 (
		\PhyAddrPointer_reg[17]/NET0131 ,
		_w681_,
		_w1666_
	);
	LUT3 #(
		.INIT('h82)
	) name1214 (
		_w844_,
		_w906_,
		_w1416_,
		_w1667_
	);
	LUT4 #(
		.INIT('h0008)
	) name1215 (
		_w974_,
		_w987_,
		_w988_,
		_w991_,
		_w1668_
	);
	LUT4 #(
		.INIT('hb000)
	) name1216 (
		_w1345_,
		_w1346_,
		_w1348_,
		_w1668_,
		_w1669_
	);
	LUT4 #(
		.INIT('h8aa8)
	) name1217 (
		_w681_,
		_w844_,
		_w993_,
		_w1669_,
		_w1670_
	);
	LUT4 #(
		.INIT('h8a88)
	) name1218 (
		_w574_,
		_w1666_,
		_w1667_,
		_w1670_,
		_w1671_
	);
	LUT4 #(
		.INIT('h2888)
	) name1219 (
		_w688_,
		_w1069_,
		_w1054_,
		_w1067_,
		_w1672_
	);
	LUT4 #(
		.INIT('h028a)
	) name1220 (
		\PhyAddrPointer_reg[17]/NET0131 ,
		_w573_,
		_w574_,
		_w605_,
		_w1673_
	);
	LUT2 #(
		.INIT('h1)
	) name1221 (
		_w1672_,
		_w1673_,
		_w1674_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name1222 (
		\PhyAddrPointer_reg[17]/NET0131 ,
		\PhyAddrPointer_reg[1]/NET0131 ,
		_w1264_,
		_w1266_,
		_w1675_
	);
	LUT4 #(
		.INIT('h08aa)
	) name1223 (
		\PhyAddrPointer_reg[17]/NET0131 ,
		_w707_,
		_w1656_,
		_w1283_,
		_w1676_
	);
	LUT3 #(
		.INIT('h20)
	) name1224 (
		\DataWidth_reg[1]/NET0131 ,
		\PhyAddrPointer_reg[17]/NET0131 ,
		_w700_,
		_w1677_
	);
	LUT2 #(
		.INIT('h8)
	) name1225 (
		\rEIP_reg[17]/NET0131 ,
		_w1109_,
		_w1678_
	);
	LUT3 #(
		.INIT('h07)
	) name1226 (
		_w1656_,
		_w1677_,
		_w1678_,
		_w1679_
	);
	LUT4 #(
		.INIT('h1300)
	) name1227 (
		_w1281_,
		_w1676_,
		_w1675_,
		_w1679_,
		_w1680_
	);
	LUT4 #(
		.INIT('h8aff)
	) name1228 (
		_w695_,
		_w1671_,
		_w1674_,
		_w1680_,
		_w1681_
	);
	LUT2 #(
		.INIT('h2)
	) name1229 (
		\PhyAddrPointer_reg[18]/NET0131 ,
		_w681_,
		_w1682_
	);
	LUT4 #(
		.INIT('hb4f0)
	) name1230 (
		_w863_,
		_w907_,
		_w909_,
		_w1113_,
		_w1683_
	);
	LUT4 #(
		.INIT('h1411)
	) name1231 (
		_w844_,
		_w992_,
		_w993_,
		_w1669_,
		_w1684_
	);
	LUT4 #(
		.INIT('h0a02)
	) name1232 (
		_w681_,
		_w844_,
		_w1684_,
		_w1683_,
		_w1685_
	);
	LUT4 #(
		.INIT('h028a)
	) name1233 (
		\PhyAddrPointer_reg[18]/NET0131 ,
		_w573_,
		_w574_,
		_w605_,
		_w1686_
	);
	LUT4 #(
		.INIT('h2000)
	) name1234 (
		_w1139_,
		_w1145_,
		_w1150_,
		_w1152_,
		_w1687_
	);
	LUT4 #(
		.INIT('h00df)
	) name1235 (
		_w1139_,
		_w1145_,
		_w1150_,
		_w1152_,
		_w1688_
	);
	LUT3 #(
		.INIT('h02)
	) name1236 (
		_w688_,
		_w1688_,
		_w1687_,
		_w1689_
	);
	LUT4 #(
		.INIT('h00d7)
	) name1237 (
		_w688_,
		_w1151_,
		_w1152_,
		_w1686_,
		_w1690_
	);
	LUT4 #(
		.INIT('h5700)
	) name1238 (
		_w574_,
		_w1682_,
		_w1685_,
		_w1690_,
		_w1691_
	);
	LUT3 #(
		.INIT('h6a)
	) name1239 (
		\PhyAddrPointer_reg[18]/NET0131 ,
		\PhyAddrPointer_reg[1]/NET0131 ,
		_w1569_,
		_w1692_
	);
	LUT4 #(
		.INIT('h60a0)
	) name1240 (
		\PhyAddrPointer_reg[18]/NET0131 ,
		\PhyAddrPointer_reg[1]/NET0131 ,
		_w1281_,
		_w1569_,
		_w1693_
	);
	LUT4 #(
		.INIT('h3f15)
	) name1241 (
		\PhyAddrPointer_reg[18]/NET0131 ,
		\rEIP_reg[18]/NET0131 ,
		_w1109_,
		_w1283_,
		_w1694_
	);
	LUT4 #(
		.INIT('hb700)
	) name1242 (
		\PhyAddrPointer_reg[18]/NET0131 ,
		_w707_,
		_w1569_,
		_w1694_,
		_w1695_
	);
	LUT2 #(
		.INIT('h4)
	) name1243 (
		_w1693_,
		_w1695_,
		_w1696_
	);
	LUT3 #(
		.INIT('h2f)
	) name1244 (
		_w695_,
		_w1691_,
		_w1696_,
		_w1697_
	);
	LUT2 #(
		.INIT('h2)
	) name1245 (
		\PhyAddrPointer_reg[25]/NET0131 ,
		_w681_,
		_w1698_
	);
	LUT4 #(
		.INIT('haa20)
	) name1246 (
		_w574_,
		_w1422_,
		_w1423_,
		_w1698_,
		_w1699_
	);
	LUT4 #(
		.INIT('h028a)
	) name1247 (
		\PhyAddrPointer_reg[25]/NET0131 ,
		_w573_,
		_w574_,
		_w605_,
		_w1700_
	);
	LUT2 #(
		.INIT('h1)
	) name1248 (
		_w1426_,
		_w1700_,
		_w1701_
	);
	LUT3 #(
		.INIT('h48)
	) name1249 (
		\PhyAddrPointer_reg[25]/NET0131 ,
		_w700_,
		_w1624_,
		_w1702_
	);
	LUT2 #(
		.INIT('h6)
	) name1250 (
		\PhyAddrPointer_reg[25]/NET0131 ,
		_w1475_,
		_w1703_
	);
	LUT4 #(
		.INIT('h3f15)
	) name1251 (
		\PhyAddrPointer_reg[25]/NET0131 ,
		\rEIP_reg[25]/NET0131 ,
		_w1109_,
		_w1283_,
		_w1704_
	);
	LUT4 #(
		.INIT('hb700)
	) name1252 (
		\PhyAddrPointer_reg[25]/NET0131 ,
		_w706_,
		_w1475_,
		_w1704_,
		_w1705_
	);
	LUT2 #(
		.INIT('h4)
	) name1253 (
		_w1702_,
		_w1705_,
		_w1706_
	);
	LUT4 #(
		.INIT('h8aff)
	) name1254 (
		_w695_,
		_w1699_,
		_w1701_,
		_w1706_,
		_w1707_
	);
	LUT2 #(
		.INIT('h2)
	) name1255 (
		\PhyAddrPointer_reg[8]/NET0131 ,
		_w681_,
		_w1708_
	);
	LUT4 #(
		.INIT('haa20)
	) name1256 (
		_w574_,
		_w1510_,
		_w1511_,
		_w1708_,
		_w1709_
	);
	LUT4 #(
		.INIT('h028a)
	) name1257 (
		\PhyAddrPointer_reg[8]/NET0131 ,
		_w573_,
		_w574_,
		_w605_,
		_w1710_
	);
	LUT4 #(
		.INIT('h007d)
	) name1258 (
		_w688_,
		_w1052_,
		_w1145_,
		_w1710_,
		_w1711_
	);
	LUT3 #(
		.INIT('h6c)
	) name1259 (
		\PhyAddrPointer_reg[1]/NET0131 ,
		\PhyAddrPointer_reg[8]/NET0131 ,
		_w1260_,
		_w1712_
	);
	LUT4 #(
		.INIT('h4105)
	) name1260 (
		\DataWidth_reg[1]/NET0131 ,
		\PhyAddrPointer_reg[1]/NET0131 ,
		\PhyAddrPointer_reg[8]/NET0131 ,
		_w1260_,
		_w1713_
	);
	LUT4 #(
		.INIT('h78f0)
	) name1261 (
		\PhyAddrPointer_reg[6]/NET0131 ,
		\PhyAddrPointer_reg[7]/NET0131 ,
		\PhyAddrPointer_reg[8]/NET0131 ,
		_w1259_,
		_w1714_
	);
	LUT3 #(
		.INIT('hc4)
	) name1262 (
		\DataWidth_reg[1]/NET0131 ,
		_w700_,
		_w1714_,
		_w1715_
	);
	LUT4 #(
		.INIT('h60c0)
	) name1263 (
		\PhyAddrPointer_reg[1]/NET0131 ,
		\PhyAddrPointer_reg[8]/NET0131 ,
		_w706_,
		_w1260_,
		_w1716_
	);
	LUT4 #(
		.INIT('h3f15)
	) name1264 (
		\PhyAddrPointer_reg[8]/NET0131 ,
		\rEIP_reg[8]/NET0131 ,
		_w1109_,
		_w1283_,
		_w1717_
	);
	LUT4 #(
		.INIT('h4500)
	) name1265 (
		_w1716_,
		_w1713_,
		_w1715_,
		_w1717_,
		_w1718_
	);
	LUT4 #(
		.INIT('h8aff)
	) name1266 (
		_w695_,
		_w1709_,
		_w1711_,
		_w1718_,
		_w1719_
	);
	LUT4 #(
		.INIT('h00ec)
	) name1267 (
		_w514_,
		_w566_,
		_w569_,
		_w724_,
		_w1720_
	);
	LUT4 #(
		.INIT('haa8a)
	) name1268 (
		\InstAddrPointer_reg[4]/NET0131 ,
		_w637_,
		_w684_,
		_w1720_,
		_w1721_
	);
	LUT3 #(
		.INIT('hb0)
	) name1269 (
		_w582_,
		_w595_,
		_w957_,
		_w1722_
	);
	LUT3 #(
		.INIT('h4a)
	) name1270 (
		\InstAddrPointer_reg[4]/NET0131 ,
		_w605_,
		_w1025_,
		_w1723_
	);
	LUT4 #(
		.INIT('hc800)
	) name1271 (
		_w552_,
		_w576_,
		_w579_,
		_w1723_,
		_w1724_
	);
	LUT3 #(
		.INIT('h0b)
	) name1272 (
		_w645_,
		_w812_,
		_w1724_,
		_w1725_
	);
	LUT4 #(
		.INIT('h6555)
	) name1273 (
		_w812_,
		_w819_,
		_w817_,
		_w824_,
		_w1726_
	);
	LUT4 #(
		.INIT('h2fd0)
	) name1274 (
		_w765_,
		_w794_,
		_w797_,
		_w1726_,
		_w1727_
	);
	LUT4 #(
		.INIT('h08c8)
	) name1275 (
		\InstAddrPointer_reg[4]/NET0131 ,
		_w574_,
		_w681_,
		_w1727_,
		_w1728_
	);
	LUT4 #(
		.INIT('h40bf)
	) name1276 (
		_w819_,
		_w817_,
		_w824_,
		_w1026_,
		_w1729_
	);
	LUT4 #(
		.INIT('h5501)
	) name1277 (
		_w1029_,
		_w1031_,
		_w1034_,
		_w1036_,
		_w1730_
	);
	LUT3 #(
		.INIT('h28)
	) name1278 (
		_w688_,
		_w1729_,
		_w1730_,
		_w1731_
	);
	LUT2 #(
		.INIT('h1)
	) name1279 (
		_w1728_,
		_w1731_,
		_w1732_
	);
	LUT4 #(
		.INIT('h1000)
	) name1280 (
		_w1722_,
		_w1721_,
		_w1725_,
		_w1732_,
		_w1733_
	);
	LUT2 #(
		.INIT('h8)
	) name1281 (
		\rEIP_reg[4]/NET0131 ,
		_w1109_,
		_w1734_
	);
	LUT4 #(
		.INIT('h3f15)
	) name1282 (
		\InstAddrPointer_reg[4]/NET0131 ,
		\rEIP_reg[4]/NET0131 ,
		_w1109_,
		_w1110_,
		_w1735_
	);
	LUT3 #(
		.INIT('h2f)
	) name1283 (
		_w695_,
		_w1733_,
		_w1735_,
		_w1736_
	);
	LUT2 #(
		.INIT('h2)
	) name1284 (
		\InstAddrPointer_reg[6]/NET0131 ,
		_w681_,
		_w1737_
	);
	LUT3 #(
		.INIT('h95)
	) name1285 (
		_w846_,
		_w851_,
		_w856_,
		_w1738_
	);
	LUT4 #(
		.INIT('h8a20)
	) name1286 (
		_w844_,
		_w828_,
		_w831_,
		_w1738_,
		_w1739_
	);
	LUT3 #(
		.INIT('h87)
	) name1287 (
		_w851_,
		_w856_,
		_w945_,
		_w1740_
	);
	LUT4 #(
		.INIT('ha88a)
	) name1288 (
		_w681_,
		_w844_,
		_w1123_,
		_w1740_,
		_w1741_
	);
	LUT4 #(
		.INIT('h8a88)
	) name1289 (
		_w574_,
		_w1737_,
		_w1739_,
		_w1741_,
		_w1742_
	);
	LUT3 #(
		.INIT('h87)
	) name1290 (
		_w851_,
		_w856_,
		_w1041_,
		_w1743_
	);
	LUT4 #(
		.INIT('h02a8)
	) name1291 (
		_w688_,
		_w1141_,
		_w1142_,
		_w1743_,
		_w1744_
	);
	LUT4 #(
		.INIT('h008a)
	) name1292 (
		_w611_,
		_w618_,
		_w619_,
		_w798_,
		_w1745_
	);
	LUT3 #(
		.INIT('hc4)
	) name1293 (
		_w620_,
		_w846_,
		_w1745_,
		_w1746_
	);
	LUT3 #(
		.INIT('ha2)
	) name1294 (
		\InstAddrPointer_reg[6]/NET0131 ,
		_w1197_,
		_w1514_,
		_w1747_
	);
	LUT2 #(
		.INIT('h8)
	) name1295 (
		_w606_,
		_w1041_,
		_w1748_
	);
	LUT4 #(
		.INIT('h004f)
	) name1296 (
		_w582_,
		_w595_,
		_w945_,
		_w1748_,
		_w1749_
	);
	LUT4 #(
		.INIT('h0100)
	) name1297 (
		_w1747_,
		_w1746_,
		_w1744_,
		_w1749_,
		_w1750_
	);
	LUT4 #(
		.INIT('h3f15)
	) name1298 (
		\InstAddrPointer_reg[6]/NET0131 ,
		\rEIP_reg[6]/NET0131 ,
		_w1109_,
		_w1110_,
		_w1751_
	);
	LUT4 #(
		.INIT('h8aff)
	) name1299 (
		_w695_,
		_w1742_,
		_w1750_,
		_w1751_,
		_w1752_
	);
	LUT2 #(
		.INIT('h2)
	) name1300 (
		\PhyAddrPointer_reg[10]/NET0131 ,
		_w681_,
		_w1753_
	);
	LUT4 #(
		.INIT('h08c4)
	) name1301 (
		_w734_,
		_w844_,
		_w863_,
		_w1524_,
		_w1754_
	);
	LUT3 #(
		.INIT('h8a)
	) name1302 (
		_w971_,
		_w973_,
		_w1127_,
		_w1755_
	);
	LUT2 #(
		.INIT('h1)
	) name1303 (
		_w844_,
		_w979_,
		_w1756_
	);
	LUT4 #(
		.INIT('h008a)
	) name1304 (
		_w681_,
		_w1755_,
		_w1756_,
		_w1754_,
		_w1757_
	);
	LUT3 #(
		.INIT('h0d)
	) name1305 (
		_w1139_,
		_w1145_,
		_w1148_,
		_w1758_
	);
	LUT4 #(
		.INIT('haa2a)
	) name1306 (
		_w688_,
		_w1052_,
		_w1066_,
		_w1145_,
		_w1759_
	);
	LUT2 #(
		.INIT('h4)
	) name1307 (
		_w1758_,
		_w1759_,
		_w1760_
	);
	LUT4 #(
		.INIT('h028a)
	) name1308 (
		\PhyAddrPointer_reg[10]/NET0131 ,
		_w573_,
		_w574_,
		_w605_,
		_w1761_
	);
	LUT3 #(
		.INIT('h0b)
	) name1309 (
		_w1758_,
		_w1759_,
		_w1761_,
		_w1762_
	);
	LUT4 #(
		.INIT('h5700)
	) name1310 (
		_w574_,
		_w1753_,
		_w1757_,
		_w1762_,
		_w1763_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name1311 (
		\PhyAddrPointer_reg[10]/NET0131 ,
		\PhyAddrPointer_reg[1]/NET0131 ,
		\PhyAddrPointer_reg[9]/NET0131 ,
		_w1261_,
		_w1764_
	);
	LUT3 #(
		.INIT('h6a)
	) name1312 (
		\PhyAddrPointer_reg[10]/NET0131 ,
		\PhyAddrPointer_reg[9]/NET0131 ,
		_w1261_,
		_w1765_
	);
	LUT4 #(
		.INIT('hc840)
	) name1313 (
		\DataWidth_reg[1]/NET0131 ,
		_w700_,
		_w1764_,
		_w1765_,
		_w1766_
	);
	LUT4 #(
		.INIT('h3f15)
	) name1314 (
		\PhyAddrPointer_reg[10]/NET0131 ,
		\rEIP_reg[10]/NET0131 ,
		_w1109_,
		_w1283_,
		_w1767_
	);
	LUT3 #(
		.INIT('h70)
	) name1315 (
		_w706_,
		_w1764_,
		_w1767_,
		_w1768_
	);
	LUT2 #(
		.INIT('h4)
	) name1316 (
		_w1766_,
		_w1768_,
		_w1769_
	);
	LUT3 #(
		.INIT('h2f)
	) name1317 (
		_w695_,
		_w1763_,
		_w1769_,
		_w1770_
	);
	LUT4 #(
		.INIT('h8488)
	) name1318 (
		_w832_,
		_w844_,
		_w927_,
		_w928_,
		_w1771_
	);
	LUT4 #(
		.INIT('h1411)
	) name1319 (
		_w844_,
		_w943_,
		_w962_,
		_w969_,
		_w1772_
	);
	LUT4 #(
		.INIT('hddd1)
	) name1320 (
		\PhyAddrPointer_reg[7]/NET0131 ,
		_w681_,
		_w1772_,
		_w1771_,
		_w1773_
	);
	LUT4 #(
		.INIT('h40bf)
	) name1321 (
		_w834_,
		_w838_,
		_w843_,
		_w1045_,
		_w1774_
	);
	LUT3 #(
		.INIT('hb0)
	) name1322 (
		_w1038_,
		_w1043_,
		_w1049_,
		_w1775_
	);
	LUT4 #(
		.INIT('h4f00)
	) name1323 (
		_w1038_,
		_w1043_,
		_w1049_,
		_w1774_,
		_w1776_
	);
	LUT4 #(
		.INIT('h00b0)
	) name1324 (
		_w1038_,
		_w1043_,
		_w1049_,
		_w1774_,
		_w1777_
	);
	LUT3 #(
		.INIT('h02)
	) name1325 (
		_w688_,
		_w1777_,
		_w1776_,
		_w1778_
	);
	LUT4 #(
		.INIT('h028a)
	) name1326 (
		\PhyAddrPointer_reg[7]/NET0131 ,
		_w573_,
		_w574_,
		_w605_,
		_w1779_
	);
	LUT4 #(
		.INIT('h007d)
	) name1327 (
		_w688_,
		_w1774_,
		_w1775_,
		_w1779_,
		_w1780_
	);
	LUT4 #(
		.INIT('h08cc)
	) name1328 (
		_w574_,
		_w695_,
		_w1773_,
		_w1780_,
		_w1781_
	);
	LUT4 #(
		.INIT('h78f0)
	) name1329 (
		\PhyAddrPointer_reg[1]/NET0131 ,
		\PhyAddrPointer_reg[6]/NET0131 ,
		\PhyAddrPointer_reg[7]/NET0131 ,
		_w1259_,
		_w1782_
	);
	LUT3 #(
		.INIT('h6c)
	) name1330 (
		\PhyAddrPointer_reg[6]/NET0131 ,
		\PhyAddrPointer_reg[7]/NET0131 ,
		_w1259_,
		_w1783_
	);
	LUT4 #(
		.INIT('hc840)
	) name1331 (
		\DataWidth_reg[1]/NET0131 ,
		_w700_,
		_w1782_,
		_w1783_,
		_w1784_
	);
	LUT4 #(
		.INIT('h3f15)
	) name1332 (
		\PhyAddrPointer_reg[7]/NET0131 ,
		\rEIP_reg[7]/NET0131 ,
		_w1109_,
		_w1283_,
		_w1785_
	);
	LUT3 #(
		.INIT('h70)
	) name1333 (
		_w706_,
		_w1782_,
		_w1785_,
		_w1786_
	);
	LUT2 #(
		.INIT('h4)
	) name1334 (
		_w1784_,
		_w1786_,
		_w1787_
	);
	LUT2 #(
		.INIT('hb)
	) name1335 (
		_w1781_,
		_w1787_,
		_w1788_
	);
	LUT2 #(
		.INIT('h2)
	) name1336 (
		\InstAddrPointer_reg[3]/NET0131 ,
		_w681_,
		_w1789_
	);
	LUT4 #(
		.INIT('h40bf)
	) name1337 (
		_w739_,
		_w743_,
		_w748_,
		_w750_,
		_w1790_
	);
	LUT4 #(
		.INIT('h02a8)
	) name1338 (
		_w844_,
		_w764_,
		_w923_,
		_w1790_,
		_w1791_
	);
	LUT3 #(
		.INIT('h10)
	) name1339 (
		_w956_,
		_w960_,
		_w1120_,
		_w1792_
	);
	LUT4 #(
		.INIT('h40bf)
	) name1340 (
		_w739_,
		_w743_,
		_w748_,
		_w959_,
		_w1793_
	);
	LUT4 #(
		.INIT('h5501)
	) name1341 (
		_w844_,
		_w951_,
		_w956_,
		_w1793_,
		_w1794_
	);
	LUT4 #(
		.INIT('h008a)
	) name1342 (
		_w681_,
		_w1792_,
		_w1794_,
		_w1791_,
		_w1795_
	);
	LUT3 #(
		.INIT('ha8)
	) name1343 (
		_w574_,
		_w1789_,
		_w1795_,
		_w1796_
	);
	LUT3 #(
		.INIT('hb0)
	) name1344 (
		_w582_,
		_w595_,
		_w959_,
		_w1797_
	);
	LUT4 #(
		.INIT('h40bf)
	) name1345 (
		_w739_,
		_w743_,
		_w748_,
		_w1028_,
		_w1798_
	);
	LUT3 #(
		.INIT('h0e)
	) name1346 (
		_w1031_,
		_w1034_,
		_w1798_,
		_w1799_
	);
	LUT3 #(
		.INIT('h10)
	) name1347 (
		_w1031_,
		_w1034_,
		_w1798_,
		_w1800_
	);
	LUT3 #(
		.INIT('h02)
	) name1348 (
		_w688_,
		_w1800_,
		_w1799_,
		_w1801_
	);
	LUT2 #(
		.INIT('h8)
	) name1349 (
		_w549_,
		_w750_,
		_w1802_
	);
	LUT3 #(
		.INIT('h07)
	) name1350 (
		_w606_,
		_w1028_,
		_w1802_,
		_w1803_
	);
	LUT2 #(
		.INIT('h4)
	) name1351 (
		_w1801_,
		_w1803_,
		_w1804_
	);
	LUT3 #(
		.INIT('h80)
	) name1352 (
		\InstAddrPointer_reg[3]/NET0131 ,
		_w514_,
		_w569_,
		_w1805_
	);
	LUT4 #(
		.INIT('h0075)
	) name1353 (
		_w611_,
		_w618_,
		_w619_,
		_w1805_,
		_w1806_
	);
	LUT4 #(
		.INIT('hf078)
	) name1354 (
		\InstAddrPointer_reg[1]/NET0131 ,
		\InstAddrPointer_reg[2]/NET0131 ,
		\InstAddrPointer_reg[3]/NET0131 ,
		READY_n_pad,
		_w1807_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name1355 (
		\InstAddrPointer_reg[3]/NET0131 ,
		_w1197_,
		_w1806_,
		_w1807_,
		_w1808_
	);
	LUT4 #(
		.INIT('h1000)
	) name1356 (
		_w1797_,
		_w1796_,
		_w1804_,
		_w1808_,
		_w1809_
	);
	LUT4 #(
		.INIT('h3f15)
	) name1357 (
		\InstAddrPointer_reg[3]/NET0131 ,
		\rEIP_reg[3]/NET0131 ,
		_w1109_,
		_w1110_,
		_w1810_
	);
	LUT3 #(
		.INIT('h2f)
	) name1358 (
		_w695_,
		_w1809_,
		_w1810_,
		_w1811_
	);
	LUT3 #(
		.INIT('h95)
	) name1359 (
		_w799_,
		_w804_,
		_w809_,
		_w1812_
	);
	LUT4 #(
		.INIT('h4fb0)
	) name1360 (
		_w923_,
		_w924_,
		_w925_,
		_w1812_,
		_w1813_
	);
	LUT4 #(
		.INIT('h08c8)
	) name1361 (
		\InstAddrPointer_reg[5]/NET0131 ,
		_w574_,
		_w681_,
		_w1813_,
		_w1814_
	);
	LUT3 #(
		.INIT('h87)
	) name1362 (
		_w804_,
		_w809_,
		_w1039_,
		_w1815_
	);
	LUT3 #(
		.INIT('h82)
	) name1363 (
		_w688_,
		_w1038_,
		_w1815_,
		_w1816_
	);
	LUT3 #(
		.INIT('h8a)
	) name1364 (
		\InstAddrPointer_reg[5]/NET0131 ,
		_w637_,
		_w684_,
		_w1817_
	);
	LUT2 #(
		.INIT('h4)
	) name1365 (
		_w645_,
		_w799_,
		_w1818_
	);
	LUT2 #(
		.INIT('h8)
	) name1366 (
		_w606_,
		_w1039_,
		_w1819_
	);
	LUT4 #(
		.INIT('h004f)
	) name1367 (
		_w582_,
		_w595_,
		_w947_,
		_w1819_,
		_w1820_
	);
	LUT4 #(
		.INIT('h0100)
	) name1368 (
		_w1817_,
		_w1818_,
		_w1816_,
		_w1820_,
		_w1821_
	);
	LUT4 #(
		.INIT('h3f15)
	) name1369 (
		\InstAddrPointer_reg[5]/NET0131 ,
		\rEIP_reg[5]/NET0131 ,
		_w1109_,
		_w1110_,
		_w1822_
	);
	LUT4 #(
		.INIT('h8aff)
	) name1370 (
		_w695_,
		_w1814_,
		_w1821_,
		_w1822_,
		_w1823_
	);
	LUT4 #(
		.INIT('hfc7f)
	) name1371 (
		\State2_reg[0]/NET0131 ,
		\State2_reg[1]/NET0131 ,
		\State2_reg[2]/NET0131 ,
		\State2_reg[3]/NET0131 ,
		_w1824_
	);
	LUT4 #(
		.INIT('hfc20)
	) name1372 (
		\State2_reg[0]/NET0131 ,
		\State2_reg[1]/NET0131 ,
		\State2_reg[2]/NET0131 ,
		\State2_reg[3]/NET0131 ,
		_w1825_
	);
	LUT2 #(
		.INIT('h2)
	) name1373 (
		\EAX_reg[31]/NET0131 ,
		_w1825_,
		_w1826_
	);
	LUT4 #(
		.INIT('h8000)
	) name1374 (
		\EAX_reg[0]/NET0131 ,
		\EAX_reg[1]/NET0131 ,
		\EAX_reg[2]/NET0131 ,
		\EAX_reg[3]/NET0131 ,
		_w1827_
	);
	LUT4 #(
		.INIT('h8000)
	) name1375 (
		\EAX_reg[4]/NET0131 ,
		\EAX_reg[5]/NET0131 ,
		\EAX_reg[6]/NET0131 ,
		_w1827_,
		_w1828_
	);
	LUT4 #(
		.INIT('h8000)
	) name1376 (
		\EAX_reg[7]/NET0131 ,
		\EAX_reg[8]/NET0131 ,
		\EAX_reg[9]/NET0131 ,
		_w1828_,
		_w1829_
	);
	LUT2 #(
		.INIT('h8)
	) name1377 (
		\EAX_reg[10]/NET0131 ,
		_w1829_,
		_w1830_
	);
	LUT3 #(
		.INIT('h80)
	) name1378 (
		\EAX_reg[10]/NET0131 ,
		\EAX_reg[11]/NET0131 ,
		_w1829_,
		_w1831_
	);
	LUT4 #(
		.INIT('h8000)
	) name1379 (
		\EAX_reg[10]/NET0131 ,
		\EAX_reg[11]/NET0131 ,
		\EAX_reg[12]/NET0131 ,
		_w1829_,
		_w1832_
	);
	LUT2 #(
		.INIT('h8)
	) name1380 (
		\EAX_reg[13]/NET0131 ,
		_w1832_,
		_w1833_
	);
	LUT3 #(
		.INIT('h80)
	) name1381 (
		\EAX_reg[13]/NET0131 ,
		\EAX_reg[14]/NET0131 ,
		_w1832_,
		_w1834_
	);
	LUT4 #(
		.INIT('h8000)
	) name1382 (
		\EAX_reg[13]/NET0131 ,
		\EAX_reg[14]/NET0131 ,
		\EAX_reg[15]/NET0131 ,
		_w1832_,
		_w1835_
	);
	LUT3 #(
		.INIT('h80)
	) name1383 (
		\EAX_reg[16]/NET0131 ,
		\EAX_reg[17]/NET0131 ,
		_w1835_,
		_w1836_
	);
	LUT4 #(
		.INIT('h8000)
	) name1384 (
		\EAX_reg[16]/NET0131 ,
		\EAX_reg[17]/NET0131 ,
		\EAX_reg[18]/NET0131 ,
		_w1835_,
		_w1837_
	);
	LUT2 #(
		.INIT('h8)
	) name1385 (
		\EAX_reg[20]/NET0131 ,
		\EAX_reg[21]/NET0131 ,
		_w1838_
	);
	LUT3 #(
		.INIT('h80)
	) name1386 (
		\EAX_reg[20]/NET0131 ,
		\EAX_reg[21]/NET0131 ,
		\EAX_reg[22]/NET0131 ,
		_w1839_
	);
	LUT3 #(
		.INIT('h80)
	) name1387 (
		\EAX_reg[19]/NET0131 ,
		_w1837_,
		_w1839_,
		_w1840_
	);
	LUT2 #(
		.INIT('h8)
	) name1388 (
		\EAX_reg[23]/NET0131 ,
		\EAX_reg[24]/NET0131 ,
		_w1841_
	);
	LUT3 #(
		.INIT('h80)
	) name1389 (
		\EAX_reg[23]/NET0131 ,
		\EAX_reg[24]/NET0131 ,
		\EAX_reg[25]/NET0131 ,
		_w1842_
	);
	LUT2 #(
		.INIT('h8)
	) name1390 (
		\EAX_reg[26]/NET0131 ,
		\EAX_reg[27]/NET0131 ,
		_w1843_
	);
	LUT2 #(
		.INIT('h8)
	) name1391 (
		_w1842_,
		_w1843_,
		_w1844_
	);
	LUT4 #(
		.INIT('h8000)
	) name1392 (
		\EAX_reg[19]/NET0131 ,
		_w1837_,
		_w1839_,
		_w1844_,
		_w1845_
	);
	LUT2 #(
		.INIT('h8)
	) name1393 (
		\EAX_reg[28]/NET0131 ,
		\EAX_reg[29]/NET0131 ,
		_w1846_
	);
	LUT3 #(
		.INIT('h80)
	) name1394 (
		\EAX_reg[30]/NET0131 ,
		_w1845_,
		_w1846_,
		_w1847_
	);
	LUT4 #(
		.INIT('h8000)
	) name1395 (
		_w515_,
		_w536_,
		_w565_,
		_w585_,
		_w1848_
	);
	LUT3 #(
		.INIT('h80)
	) name1396 (
		_w576_,
		_w579_,
		_w605_,
		_w1849_
	);
	LUT4 #(
		.INIT('h0013)
	) name1397 (
		_w514_,
		_w566_,
		_w569_,
		_w1848_,
		_w1850_
	);
	LUT3 #(
		.INIT('h32)
	) name1398 (
		_w580_,
		_w1849_,
		_w1850_,
		_w1851_
	);
	LUT4 #(
		.INIT('h080d)
	) name1399 (
		_w580_,
		_w605_,
		_w623_,
		_w1850_,
		_w1852_
	);
	LUT4 #(
		.INIT('h135f)
	) name1400 (
		\InstQueue_reg[0][7]/NET0131 ,
		\InstQueue_reg[14][7]/NET0131 ,
		_w456_,
		_w458_,
		_w1853_
	);
	LUT4 #(
		.INIT('h153f)
	) name1401 (
		\InstQueue_reg[2][7]/NET0131 ,
		\InstQueue_reg[9][7]/NET0131 ,
		_w461_,
		_w473_,
		_w1854_
	);
	LUT4 #(
		.INIT('h153f)
	) name1402 (
		\InstQueue_reg[11][7]/NET0131 ,
		\InstQueue_reg[5][7]/NET0131 ,
		_w474_,
		_w468_,
		_w1855_
	);
	LUT4 #(
		.INIT('h135f)
	) name1403 (
		\InstQueue_reg[4][7]/NET0131 ,
		\InstQueue_reg[8][7]/NET0131 ,
		_w453_,
		_w467_,
		_w1856_
	);
	LUT4 #(
		.INIT('h8000)
	) name1404 (
		_w1855_,
		_w1856_,
		_w1853_,
		_w1854_,
		_w1857_
	);
	LUT4 #(
		.INIT('h135f)
	) name1405 (
		\InstQueue_reg[10][7]/NET0131 ,
		\InstQueue_reg[15][7]/NET0131 ,
		_w477_,
		_w470_,
		_w1858_
	);
	LUT4 #(
		.INIT('h153f)
	) name1406 (
		\InstQueue_reg[13][7]/NET0131 ,
		\InstQueue_reg[6][7]/NET0131 ,
		_w476_,
		_w471_,
		_w1859_
	);
	LUT4 #(
		.INIT('h135f)
	) name1407 (
		\InstQueue_reg[1][7]/NET0131 ,
		\InstQueue_reg[3][7]/NET0131 ,
		_w460_,
		_w463_,
		_w1860_
	);
	LUT4 #(
		.INIT('h153f)
	) name1408 (
		\InstQueue_reg[12][7]/NET0131 ,
		\InstQueue_reg[7][7]/NET0131 ,
		_w464_,
		_w454_,
		_w1861_
	);
	LUT4 #(
		.INIT('h8000)
	) name1409 (
		_w1860_,
		_w1861_,
		_w1858_,
		_w1859_,
		_w1862_
	);
	LUT4 #(
		.INIT('h135f)
	) name1410 (
		\InstQueue_reg[15][0]/NET0131 ,
		\InstQueue_reg[7][0]/NET0131 ,
		_w458_,
		_w476_,
		_w1863_
	);
	LUT4 #(
		.INIT('h153f)
	) name1411 (
		\InstQueue_reg[3][0]/NET0131 ,
		\InstQueue_reg[4][0]/NET0131 ,
		_w463_,
		_w473_,
		_w1864_
	);
	LUT4 #(
		.INIT('h153f)
	) name1412 (
		\InstQueue_reg[0][0]/NET0131 ,
		\InstQueue_reg[10][0]/NET0131 ,
		_w461_,
		_w470_,
		_w1865_
	);
	LUT4 #(
		.INIT('h135f)
	) name1413 (
		\InstQueue_reg[8][0]/NET0131 ,
		\InstQueue_reg[9][0]/NET0131 ,
		_w464_,
		_w467_,
		_w1866_
	);
	LUT4 #(
		.INIT('h8000)
	) name1414 (
		_w1865_,
		_w1866_,
		_w1863_,
		_w1864_,
		_w1867_
	);
	LUT4 #(
		.INIT('h153f)
	) name1415 (
		\InstQueue_reg[11][0]/NET0131 ,
		\InstQueue_reg[5][0]/NET0131 ,
		_w453_,
		_w477_,
		_w1868_
	);
	LUT4 #(
		.INIT('h135f)
	) name1416 (
		\InstQueue_reg[13][0]/NET0131 ,
		\InstQueue_reg[6][0]/NET0131 ,
		_w454_,
		_w474_,
		_w1869_
	);
	LUT4 #(
		.INIT('h153f)
	) name1417 (
		\InstQueue_reg[12][0]/NET0131 ,
		\InstQueue_reg[2][0]/NET0131 ,
		_w460_,
		_w468_,
		_w1870_
	);
	LUT4 #(
		.INIT('h153f)
	) name1418 (
		\InstQueue_reg[14][0]/NET0131 ,
		\InstQueue_reg[1][0]/NET0131 ,
		_w456_,
		_w471_,
		_w1871_
	);
	LUT4 #(
		.INIT('h8000)
	) name1419 (
		_w1870_,
		_w1871_,
		_w1868_,
		_w1869_,
		_w1872_
	);
	LUT4 #(
		.INIT('h0777)
	) name1420 (
		_w1857_,
		_w1862_,
		_w1867_,
		_w1872_,
		_w1873_
	);
	LUT4 #(
		.INIT('h135f)
	) name1421 (
		\InstQueue_reg[11][1]/NET0131 ,
		\InstQueue_reg[9][1]/NET0131 ,
		_w477_,
		_w467_,
		_w1874_
	);
	LUT4 #(
		.INIT('h153f)
	) name1422 (
		\InstQueue_reg[15][1]/NET0131 ,
		\InstQueue_reg[4][1]/NET0131 ,
		_w463_,
		_w458_,
		_w1875_
	);
	LUT4 #(
		.INIT('h153f)
	) name1423 (
		\InstQueue_reg[1][1]/NET0131 ,
		\InstQueue_reg[8][1]/NET0131 ,
		_w464_,
		_w456_,
		_w1876_
	);
	LUT4 #(
		.INIT('h153f)
	) name1424 (
		\InstQueue_reg[0][1]/NET0131 ,
		\InstQueue_reg[6][1]/NET0131 ,
		_w474_,
		_w470_,
		_w1877_
	);
	LUT4 #(
		.INIT('h8000)
	) name1425 (
		_w1876_,
		_w1877_,
		_w1874_,
		_w1875_,
		_w1878_
	);
	LUT4 #(
		.INIT('h135f)
	) name1426 (
		\InstQueue_reg[3][1]/NET0131 ,
		\InstQueue_reg[7][1]/NET0131 ,
		_w473_,
		_w476_,
		_w1879_
	);
	LUT4 #(
		.INIT('h135f)
	) name1427 (
		\InstQueue_reg[13][1]/NET0131 ,
		\InstQueue_reg[14][1]/NET0131 ,
		_w454_,
		_w471_,
		_w1880_
	);
	LUT4 #(
		.INIT('h153f)
	) name1428 (
		\InstQueue_reg[12][1]/NET0131 ,
		\InstQueue_reg[2][1]/NET0131 ,
		_w460_,
		_w468_,
		_w1881_
	);
	LUT4 #(
		.INIT('h135f)
	) name1429 (
		\InstQueue_reg[10][1]/NET0131 ,
		\InstQueue_reg[5][1]/NET0131 ,
		_w461_,
		_w453_,
		_w1882_
	);
	LUT4 #(
		.INIT('h8000)
	) name1430 (
		_w1881_,
		_w1882_,
		_w1879_,
		_w1880_,
		_w1883_
	);
	LUT2 #(
		.INIT('h8)
	) name1431 (
		_w1878_,
		_w1883_,
		_w1884_
	);
	LUT4 #(
		.INIT('h153f)
	) name1432 (
		\InstQueue_reg[3][2]/NET0131 ,
		\InstQueue_reg[5][2]/NET0131 ,
		_w453_,
		_w473_,
		_w1885_
	);
	LUT4 #(
		.INIT('h153f)
	) name1433 (
		\InstQueue_reg[14][2]/NET0131 ,
		\InstQueue_reg[8][2]/NET0131 ,
		_w464_,
		_w471_,
		_w1886_
	);
	LUT4 #(
		.INIT('h153f)
	) name1434 (
		\InstQueue_reg[15][2]/NET0131 ,
		\InstQueue_reg[1][2]/NET0131 ,
		_w456_,
		_w458_,
		_w1887_
	);
	LUT4 #(
		.INIT('h153f)
	) name1435 (
		\InstQueue_reg[13][2]/NET0131 ,
		\InstQueue_reg[4][2]/NET0131 ,
		_w463_,
		_w454_,
		_w1888_
	);
	LUT4 #(
		.INIT('h8000)
	) name1436 (
		_w1887_,
		_w1888_,
		_w1885_,
		_w1886_,
		_w1889_
	);
	LUT4 #(
		.INIT('h135f)
	) name1437 (
		\InstQueue_reg[11][2]/NET0131 ,
		\InstQueue_reg[9][2]/NET0131 ,
		_w477_,
		_w467_,
		_w1890_
	);
	LUT4 #(
		.INIT('h135f)
	) name1438 (
		\InstQueue_reg[10][2]/NET0131 ,
		\InstQueue_reg[7][2]/NET0131 ,
		_w461_,
		_w476_,
		_w1891_
	);
	LUT4 #(
		.INIT('h135f)
	) name1439 (
		\InstQueue_reg[2][2]/NET0131 ,
		\InstQueue_reg[6][2]/NET0131 ,
		_w460_,
		_w474_,
		_w1892_
	);
	LUT4 #(
		.INIT('h153f)
	) name1440 (
		\InstQueue_reg[0][2]/NET0131 ,
		\InstQueue_reg[12][2]/NET0131 ,
		_w468_,
		_w470_,
		_w1893_
	);
	LUT4 #(
		.INIT('h8000)
	) name1441 (
		_w1892_,
		_w1893_,
		_w1890_,
		_w1891_,
		_w1894_
	);
	LUT2 #(
		.INIT('h8)
	) name1442 (
		_w1889_,
		_w1894_,
		_w1895_
	);
	LUT4 #(
		.INIT('h153f)
	) name1443 (
		\InstQueue_reg[3][3]/NET0131 ,
		\InstQueue_reg[5][3]/NET0131 ,
		_w453_,
		_w473_,
		_w1896_
	);
	LUT4 #(
		.INIT('h153f)
	) name1444 (
		\InstQueue_reg[14][3]/NET0131 ,
		\InstQueue_reg[8][3]/NET0131 ,
		_w464_,
		_w471_,
		_w1897_
	);
	LUT4 #(
		.INIT('h153f)
	) name1445 (
		\InstQueue_reg[15][3]/NET0131 ,
		\InstQueue_reg[1][3]/NET0131 ,
		_w456_,
		_w458_,
		_w1898_
	);
	LUT4 #(
		.INIT('h153f)
	) name1446 (
		\InstQueue_reg[13][3]/NET0131 ,
		\InstQueue_reg[4][3]/NET0131 ,
		_w463_,
		_w454_,
		_w1899_
	);
	LUT4 #(
		.INIT('h8000)
	) name1447 (
		_w1898_,
		_w1899_,
		_w1896_,
		_w1897_,
		_w1900_
	);
	LUT4 #(
		.INIT('h135f)
	) name1448 (
		\InstQueue_reg[11][3]/NET0131 ,
		\InstQueue_reg[9][3]/NET0131 ,
		_w477_,
		_w467_,
		_w1901_
	);
	LUT4 #(
		.INIT('h135f)
	) name1449 (
		\InstQueue_reg[10][3]/NET0131 ,
		\InstQueue_reg[7][3]/NET0131 ,
		_w461_,
		_w476_,
		_w1902_
	);
	LUT4 #(
		.INIT('h135f)
	) name1450 (
		\InstQueue_reg[2][3]/NET0131 ,
		\InstQueue_reg[6][3]/NET0131 ,
		_w460_,
		_w474_,
		_w1903_
	);
	LUT4 #(
		.INIT('h153f)
	) name1451 (
		\InstQueue_reg[0][3]/NET0131 ,
		\InstQueue_reg[12][3]/NET0131 ,
		_w468_,
		_w470_,
		_w1904_
	);
	LUT4 #(
		.INIT('h8000)
	) name1452 (
		_w1903_,
		_w1904_,
		_w1901_,
		_w1902_,
		_w1905_
	);
	LUT2 #(
		.INIT('h8)
	) name1453 (
		_w1900_,
		_w1905_,
		_w1906_
	);
	LUT4 #(
		.INIT('h0002)
	) name1454 (
		_w1873_,
		_w1884_,
		_w1895_,
		_w1906_,
		_w1907_
	);
	LUT4 #(
		.INIT('h135f)
	) name1455 (
		\InstQueue_reg[11][4]/NET0131 ,
		\InstQueue_reg[9][4]/NET0131 ,
		_w477_,
		_w467_,
		_w1908_
	);
	LUT4 #(
		.INIT('h153f)
	) name1456 (
		\InstQueue_reg[15][4]/NET0131 ,
		\InstQueue_reg[4][4]/NET0131 ,
		_w463_,
		_w458_,
		_w1909_
	);
	LUT4 #(
		.INIT('h153f)
	) name1457 (
		\InstQueue_reg[1][4]/NET0131 ,
		\InstQueue_reg[8][4]/NET0131 ,
		_w464_,
		_w456_,
		_w1910_
	);
	LUT4 #(
		.INIT('h153f)
	) name1458 (
		\InstQueue_reg[0][4]/NET0131 ,
		\InstQueue_reg[6][4]/NET0131 ,
		_w474_,
		_w470_,
		_w1911_
	);
	LUT4 #(
		.INIT('h8000)
	) name1459 (
		_w1910_,
		_w1911_,
		_w1908_,
		_w1909_,
		_w1912_
	);
	LUT4 #(
		.INIT('h135f)
	) name1460 (
		\InstQueue_reg[3][4]/NET0131 ,
		\InstQueue_reg[7][4]/NET0131 ,
		_w473_,
		_w476_,
		_w1913_
	);
	LUT4 #(
		.INIT('h135f)
	) name1461 (
		\InstQueue_reg[13][4]/NET0131 ,
		\InstQueue_reg[14][4]/NET0131 ,
		_w454_,
		_w471_,
		_w1914_
	);
	LUT4 #(
		.INIT('h153f)
	) name1462 (
		\InstQueue_reg[12][4]/NET0131 ,
		\InstQueue_reg[2][4]/NET0131 ,
		_w460_,
		_w468_,
		_w1915_
	);
	LUT4 #(
		.INIT('h135f)
	) name1463 (
		\InstQueue_reg[10][4]/NET0131 ,
		\InstQueue_reg[5][4]/NET0131 ,
		_w461_,
		_w453_,
		_w1916_
	);
	LUT4 #(
		.INIT('h8000)
	) name1464 (
		_w1915_,
		_w1916_,
		_w1913_,
		_w1914_,
		_w1917_
	);
	LUT2 #(
		.INIT('h8)
	) name1465 (
		_w1912_,
		_w1917_,
		_w1918_
	);
	LUT4 #(
		.INIT('h135f)
	) name1466 (
		\InstQueue_reg[3][5]/NET0131 ,
		\InstQueue_reg[9][5]/NET0131 ,
		_w473_,
		_w467_,
		_w1919_
	);
	LUT4 #(
		.INIT('h153f)
	) name1467 (
		\InstQueue_reg[14][5]/NET0131 ,
		\InstQueue_reg[6][5]/NET0131 ,
		_w474_,
		_w471_,
		_w1920_
	);
	LUT4 #(
		.INIT('h135f)
	) name1468 (
		\InstQueue_reg[10][5]/NET0131 ,
		\InstQueue_reg[12][5]/NET0131 ,
		_w461_,
		_w468_,
		_w1921_
	);
	LUT4 #(
		.INIT('h153f)
	) name1469 (
		\InstQueue_reg[13][5]/NET0131 ,
		\InstQueue_reg[4][5]/NET0131 ,
		_w463_,
		_w454_,
		_w1922_
	);
	LUT4 #(
		.INIT('h8000)
	) name1470 (
		_w1921_,
		_w1922_,
		_w1919_,
		_w1920_,
		_w1923_
	);
	LUT4 #(
		.INIT('h153f)
	) name1471 (
		\InstQueue_reg[11][5]/NET0131 ,
		\InstQueue_reg[5][5]/NET0131 ,
		_w453_,
		_w477_,
		_w1924_
	);
	LUT4 #(
		.INIT('h153f)
	) name1472 (
		\InstQueue_reg[1][5]/NET0131 ,
		\InstQueue_reg[8][5]/NET0131 ,
		_w464_,
		_w456_,
		_w1925_
	);
	LUT4 #(
		.INIT('h153f)
	) name1473 (
		\InstQueue_reg[0][5]/NET0131 ,
		\InstQueue_reg[2][5]/NET0131 ,
		_w460_,
		_w470_,
		_w1926_
	);
	LUT4 #(
		.INIT('h135f)
	) name1474 (
		\InstQueue_reg[15][5]/NET0131 ,
		\InstQueue_reg[7][5]/NET0131 ,
		_w458_,
		_w476_,
		_w1927_
	);
	LUT4 #(
		.INIT('h8000)
	) name1475 (
		_w1926_,
		_w1927_,
		_w1924_,
		_w1925_,
		_w1928_
	);
	LUT2 #(
		.INIT('h8)
	) name1476 (
		_w1923_,
		_w1928_,
		_w1929_
	);
	LUT4 #(
		.INIT('h135f)
	) name1477 (
		\InstQueue_reg[15][6]/NET0131 ,
		\InstQueue_reg[3][6]/NET0131 ,
		_w458_,
		_w473_,
		_w1930_
	);
	LUT4 #(
		.INIT('h135f)
	) name1478 (
		\InstQueue_reg[10][6]/NET0131 ,
		\InstQueue_reg[9][6]/NET0131 ,
		_w461_,
		_w467_,
		_w1931_
	);
	LUT4 #(
		.INIT('h153f)
	) name1479 (
		\InstQueue_reg[14][6]/NET0131 ,
		\InstQueue_reg[1][6]/NET0131 ,
		_w456_,
		_w471_,
		_w1932_
	);
	LUT4 #(
		.INIT('h153f)
	) name1480 (
		\InstQueue_reg[0][6]/NET0131 ,
		\InstQueue_reg[8][6]/NET0131 ,
		_w464_,
		_w470_,
		_w1933_
	);
	LUT4 #(
		.INIT('h8000)
	) name1481 (
		_w1932_,
		_w1933_,
		_w1930_,
		_w1931_,
		_w1934_
	);
	LUT4 #(
		.INIT('h153f)
	) name1482 (
		\InstQueue_reg[11][6]/NET0131 ,
		\InstQueue_reg[5][6]/NET0131 ,
		_w453_,
		_w477_,
		_w1935_
	);
	LUT4 #(
		.INIT('h135f)
	) name1483 (
		\InstQueue_reg[4][6]/NET0131 ,
		\InstQueue_reg[6][6]/NET0131 ,
		_w463_,
		_w474_,
		_w1936_
	);
	LUT4 #(
		.INIT('h153f)
	) name1484 (
		\InstQueue_reg[12][6]/NET0131 ,
		\InstQueue_reg[2][6]/NET0131 ,
		_w460_,
		_w468_,
		_w1937_
	);
	LUT4 #(
		.INIT('h135f)
	) name1485 (
		\InstQueue_reg[13][6]/NET0131 ,
		\InstQueue_reg[7][6]/NET0131 ,
		_w454_,
		_w476_,
		_w1938_
	);
	LUT4 #(
		.INIT('h8000)
	) name1486 (
		_w1937_,
		_w1938_,
		_w1935_,
		_w1936_,
		_w1939_
	);
	LUT2 #(
		.INIT('h8)
	) name1487 (
		_w1934_,
		_w1939_,
		_w1940_
	);
	LUT4 #(
		.INIT('h0002)
	) name1488 (
		_w1907_,
		_w1918_,
		_w1929_,
		_w1940_,
		_w1941_
	);
	LUT4 #(
		.INIT('h153f)
	) name1489 (
		\InstQueue_reg[3][7]/NET0131 ,
		\InstQueue_reg[5][7]/NET0131 ,
		_w453_,
		_w473_,
		_w1942_
	);
	LUT4 #(
		.INIT('h153f)
	) name1490 (
		\InstQueue_reg[14][7]/NET0131 ,
		\InstQueue_reg[8][7]/NET0131 ,
		_w464_,
		_w471_,
		_w1943_
	);
	LUT4 #(
		.INIT('h153f)
	) name1491 (
		\InstQueue_reg[15][7]/NET0131 ,
		\InstQueue_reg[1][7]/NET0131 ,
		_w456_,
		_w458_,
		_w1944_
	);
	LUT4 #(
		.INIT('h153f)
	) name1492 (
		\InstQueue_reg[13][7]/NET0131 ,
		\InstQueue_reg[4][7]/NET0131 ,
		_w463_,
		_w454_,
		_w1945_
	);
	LUT4 #(
		.INIT('h8000)
	) name1493 (
		_w1944_,
		_w1945_,
		_w1942_,
		_w1943_,
		_w1946_
	);
	LUT4 #(
		.INIT('h135f)
	) name1494 (
		\InstQueue_reg[11][7]/NET0131 ,
		\InstQueue_reg[9][7]/NET0131 ,
		_w477_,
		_w467_,
		_w1947_
	);
	LUT4 #(
		.INIT('h135f)
	) name1495 (
		\InstQueue_reg[10][7]/NET0131 ,
		\InstQueue_reg[7][7]/NET0131 ,
		_w461_,
		_w476_,
		_w1948_
	);
	LUT4 #(
		.INIT('h135f)
	) name1496 (
		\InstQueue_reg[2][7]/NET0131 ,
		\InstQueue_reg[6][7]/NET0131 ,
		_w460_,
		_w474_,
		_w1949_
	);
	LUT4 #(
		.INIT('h153f)
	) name1497 (
		\InstQueue_reg[0][7]/NET0131 ,
		\InstQueue_reg[12][7]/NET0131 ,
		_w468_,
		_w470_,
		_w1950_
	);
	LUT4 #(
		.INIT('h8000)
	) name1498 (
		_w1949_,
		_w1950_,
		_w1947_,
		_w1948_,
		_w1951_
	);
	LUT2 #(
		.INIT('h8)
	) name1499 (
		_w1946_,
		_w1951_,
		_w1952_
	);
	LUT4 #(
		.INIT('h8000)
	) name1500 (
		\Datai[31]_pad ,
		_w514_,
		_w569_,
		_w612_,
		_w1953_
	);
	LUT4 #(
		.INIT('h00f7)
	) name1501 (
		_w1849_,
		_w1941_,
		_w1952_,
		_w1953_,
		_w1954_
	);
	LUT4 #(
		.INIT('h7500)
	) name1502 (
		\EAX_reg[31]/NET0131 ,
		_w635_,
		_w1852_,
		_w1954_,
		_w1955_
	);
	LUT4 #(
		.INIT('hb700)
	) name1503 (
		\EAX_reg[31]/NET0131 ,
		_w1848_,
		_w1847_,
		_w1955_,
		_w1956_
	);
	LUT3 #(
		.INIT('hce)
	) name1504 (
		_w695_,
		_w1826_,
		_w1956_,
		_w1957_
	);
	LUT2 #(
		.INIT('h8)
	) name1505 (
		\EBX_reg[25]/NET0131 ,
		\EBX_reg[26]/NET0131 ,
		_w1958_
	);
	LUT2 #(
		.INIT('h8)
	) name1506 (
		\EBX_reg[21]/NET0131 ,
		\EBX_reg[22]/NET0131 ,
		_w1959_
	);
	LUT4 #(
		.INIT('h8000)
	) name1507 (
		\EBX_reg[0]/NET0131 ,
		\EBX_reg[1]/NET0131 ,
		\EBX_reg[2]/NET0131 ,
		\EBX_reg[3]/NET0131 ,
		_w1960_
	);
	LUT4 #(
		.INIT('h8000)
	) name1508 (
		\EBX_reg[4]/NET0131 ,
		\EBX_reg[5]/NET0131 ,
		\EBX_reg[6]/NET0131 ,
		_w1960_,
		_w1961_
	);
	LUT4 #(
		.INIT('h8000)
	) name1509 (
		\EBX_reg[7]/NET0131 ,
		\EBX_reg[8]/NET0131 ,
		\EBX_reg[9]/NET0131 ,
		_w1961_,
		_w1962_
	);
	LUT2 #(
		.INIT('h8)
	) name1510 (
		\EBX_reg[10]/NET0131 ,
		_w1962_,
		_w1963_
	);
	LUT3 #(
		.INIT('h80)
	) name1511 (
		\EBX_reg[10]/NET0131 ,
		\EBX_reg[11]/NET0131 ,
		_w1962_,
		_w1964_
	);
	LUT4 #(
		.INIT('h8000)
	) name1512 (
		\EBX_reg[10]/NET0131 ,
		\EBX_reg[11]/NET0131 ,
		\EBX_reg[12]/NET0131 ,
		_w1962_,
		_w1965_
	);
	LUT2 #(
		.INIT('h8)
	) name1513 (
		\EBX_reg[13]/NET0131 ,
		_w1965_,
		_w1966_
	);
	LUT3 #(
		.INIT('h80)
	) name1514 (
		\EBX_reg[13]/NET0131 ,
		\EBX_reg[14]/NET0131 ,
		_w1965_,
		_w1967_
	);
	LUT4 #(
		.INIT('h8000)
	) name1515 (
		\EBX_reg[13]/NET0131 ,
		\EBX_reg[14]/NET0131 ,
		\EBX_reg[15]/NET0131 ,
		_w1965_,
		_w1968_
	);
	LUT3 #(
		.INIT('h80)
	) name1516 (
		\EBX_reg[16]/NET0131 ,
		\EBX_reg[17]/NET0131 ,
		_w1968_,
		_w1969_
	);
	LUT3 #(
		.INIT('h80)
	) name1517 (
		\EBX_reg[18]/NET0131 ,
		\EBX_reg[19]/NET0131 ,
		\EBX_reg[20]/NET0131 ,
		_w1970_
	);
	LUT4 #(
		.INIT('h8000)
	) name1518 (
		\EBX_reg[16]/NET0131 ,
		\EBX_reg[17]/NET0131 ,
		_w1968_,
		_w1970_,
		_w1971_
	);
	LUT4 #(
		.INIT('h8000)
	) name1519 (
		\EBX_reg[23]/NET0131 ,
		\EBX_reg[24]/NET0131 ,
		_w1959_,
		_w1971_,
		_w1972_
	);
	LUT3 #(
		.INIT('h80)
	) name1520 (
		_w552_,
		_w576_,
		_w605_,
		_w1973_
	);
	LUT3 #(
		.INIT('h70)
	) name1521 (
		_w552_,
		_w576_,
		_w590_,
		_w1974_
	);
	LUT4 #(
		.INIT('h078f)
	) name1522 (
		_w552_,
		_w576_,
		_w590_,
		_w605_,
		_w1975_
	);
	LUT4 #(
		.INIT('h00d5)
	) name1523 (
		_w590_,
		_w1958_,
		_w1972_,
		_w1975_,
		_w1976_
	);
	LUT2 #(
		.INIT('h9)
	) name1524 (
		_w1907_,
		_w1918_,
		_w1977_
	);
	LUT2 #(
		.INIT('h8)
	) name1525 (
		_w1973_,
		_w1977_,
		_w1978_
	);
	LUT2 #(
		.INIT('h4)
	) name1526 (
		\EBX_reg[27]/NET0131 ,
		_w590_,
		_w1979_
	);
	LUT4 #(
		.INIT('h1555)
	) name1527 (
		_w1978_,
		_w1958_,
		_w1972_,
		_w1979_,
		_w1980_
	);
	LUT4 #(
		.INIT('h08cc)
	) name1528 (
		\EBX_reg[27]/NET0131 ,
		_w695_,
		_w1976_,
		_w1980_,
		_w1981_
	);
	LUT2 #(
		.INIT('h2)
	) name1529 (
		\EBX_reg[27]/NET0131 ,
		_w1825_,
		_w1982_
	);
	LUT2 #(
		.INIT('he)
	) name1530 (
		_w1981_,
		_w1982_,
		_w1983_
	);
	LUT4 #(
		.INIT('he420)
	) name1531 (
		_w573_,
		_w574_,
		_w605_,
		_w681_,
		_w1984_
	);
	LUT2 #(
		.INIT('h2)
	) name1532 (
		\PhyAddrPointer_reg[4]/NET0131 ,
		_w1984_,
		_w1985_
	);
	LUT3 #(
		.INIT('h08)
	) name1533 (
		_w574_,
		_w681_,
		_w1727_,
		_w1986_
	);
	LUT4 #(
		.INIT('haaa8)
	) name1534 (
		_w695_,
		_w1731_,
		_w1985_,
		_w1986_,
		_w1987_
	);
	LUT4 #(
		.INIT('h8000)
	) name1535 (
		\PhyAddrPointer_reg[1]/NET0131 ,
		\PhyAddrPointer_reg[2]/NET0131 ,
		\PhyAddrPointer_reg[3]/NET0131 ,
		\PhyAddrPointer_reg[4]/NET0131 ,
		_w1988_
	);
	LUT4 #(
		.INIT('h7f80)
	) name1536 (
		\PhyAddrPointer_reg[1]/NET0131 ,
		\PhyAddrPointer_reg[2]/NET0131 ,
		\PhyAddrPointer_reg[3]/NET0131 ,
		\PhyAddrPointer_reg[4]/NET0131 ,
		_w1989_
	);
	LUT4 #(
		.INIT('hf400)
	) name1537 (
		\DataWidth_reg[1]/NET0131 ,
		_w700_,
		_w706_,
		_w1989_,
		_w1990_
	);
	LUT2 #(
		.INIT('h2)
	) name1538 (
		\PhyAddrPointer_reg[4]/NET0131 ,
		_w1283_,
		_w1991_
	);
	LUT3 #(
		.INIT('h78)
	) name1539 (
		\PhyAddrPointer_reg[2]/NET0131 ,
		\PhyAddrPointer_reg[3]/NET0131 ,
		\PhyAddrPointer_reg[4]/NET0131 ,
		_w1992_
	);
	LUT3 #(
		.INIT('h80)
	) name1540 (
		\DataWidth_reg[1]/NET0131 ,
		_w700_,
		_w1992_,
		_w1993_
	);
	LUT4 #(
		.INIT('h0001)
	) name1541 (
		_w1734_,
		_w1993_,
		_w1991_,
		_w1990_,
		_w1994_
	);
	LUT2 #(
		.INIT('hb)
	) name1542 (
		_w1987_,
		_w1994_,
		_w1995_
	);
	LUT3 #(
		.INIT('h09)
	) name1543 (
		\InstAddrPointer_reg[1]/NET0131 ,
		\InstAddrPointer_reg[2]/NET0131 ,
		READY_n_pad,
		_w1996_
	);
	LUT2 #(
		.INIT('h2)
	) name1544 (
		_w643_,
		_w1996_,
		_w1997_
	);
	LUT4 #(
		.INIT('h0001)
	) name1545 (
		_w682_,
		_w683_,
		_w1096_,
		_w1196_,
		_w1998_
	);
	LUT3 #(
		.INIT('h8a)
	) name1546 (
		\InstAddrPointer_reg[2]/NET0131 ,
		_w1997_,
		_w1998_,
		_w1999_
	);
	LUT3 #(
		.INIT('hb0)
	) name1547 (
		_w582_,
		_w595_,
		_w950_,
		_w2000_
	);
	LUT3 #(
		.INIT('ha6)
	) name1548 (
		\InstAddrPointer_reg[2]/NET0131 ,
		_w605_,
		_w940_,
		_w2001_
	);
	LUT4 #(
		.INIT('hc800)
	) name1549 (
		_w552_,
		_w576_,
		_w579_,
		_w2001_,
		_w2002_
	);
	LUT3 #(
		.INIT('h87)
	) name1550 (
		_w757_,
		_w762_,
		_w950_,
		_w2003_
	);
	LUT4 #(
		.INIT('h00d4)
	) name1551 (
		_w780_,
		_w954_,
		_w1033_,
		_w2003_,
		_w2004_
	);
	LUT4 #(
		.INIT('h2b00)
	) name1552 (
		_w780_,
		_w954_,
		_w1033_,
		_w2003_,
		_w2005_
	);
	LUT4 #(
		.INIT('h0008)
	) name1553 (
		_w573_,
		_w605_,
		_w2005_,
		_w2004_,
		_w2006_
	);
	LUT3 #(
		.INIT('h95)
	) name1554 (
		_w752_,
		_w757_,
		_w762_,
		_w2007_
	);
	LUT4 #(
		.INIT('h008e)
	) name1555 (
		\InstAddrPointer_reg[1]/NET0131 ,
		_w780_,
		_w793_,
		_w2007_,
		_w2008_
	);
	LUT4 #(
		.INIT('h7100)
	) name1556 (
		\InstAddrPointer_reg[1]/NET0131 ,
		_w780_,
		_w793_,
		_w2007_,
		_w2009_
	);
	LUT4 #(
		.INIT('h0008)
	) name1557 (
		_w574_,
		_w681_,
		_w2009_,
		_w2008_,
		_w2010_
	);
	LUT3 #(
		.INIT('h01)
	) name1558 (
		_w2002_,
		_w2006_,
		_w2010_,
		_w2011_
	);
	LUT3 #(
		.INIT('hb0)
	) name1559 (
		_w645_,
		_w752_,
		_w2011_,
		_w2012_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name1560 (
		_w695_,
		_w1999_,
		_w2000_,
		_w2012_,
		_w2013_
	);
	LUT2 #(
		.INIT('h8)
	) name1561 (
		\rEIP_reg[2]/NET0131 ,
		_w1109_,
		_w2014_
	);
	LUT4 #(
		.INIT('h3f15)
	) name1562 (
		\InstAddrPointer_reg[2]/NET0131 ,
		\rEIP_reg[2]/NET0131 ,
		_w1109_,
		_w1110_,
		_w2015_
	);
	LUT2 #(
		.INIT('hb)
	) name1563 (
		_w2013_,
		_w2015_,
		_w2016_
	);
	LUT3 #(
		.INIT('h6a)
	) name1564 (
		\InstAddrPointer_reg[0]/NET0131 ,
		_w786_,
		_w791_,
		_w2017_
	);
	LUT3 #(
		.INIT('h08)
	) name1565 (
		_w574_,
		_w681_,
		_w2017_,
		_w2018_
	);
	LUT3 #(
		.INIT('h80)
	) name1566 (
		_w573_,
		_w605_,
		_w2017_,
		_w2019_
	);
	LUT2 #(
		.INIT('h1)
	) name1567 (
		_w2018_,
		_w2019_,
		_w2020_
	);
	LUT4 #(
		.INIT('h0010)
	) name1568 (
		\InstAddrPointer_reg[0]/NET0131 ,
		_w582_,
		_w595_,
		_w606_,
		_w2021_
	);
	LUT2 #(
		.INIT('h8)
	) name1569 (
		\InstAddrPointer_reg[0]/NET0131 ,
		_w572_,
		_w2022_
	);
	LUT2 #(
		.INIT('h8)
	) name1570 (
		_w685_,
		_w2022_,
		_w2023_
	);
	LUT4 #(
		.INIT('h222a)
	) name1571 (
		_w695_,
		_w2020_,
		_w2021_,
		_w2023_,
		_w2024_
	);
	LUT2 #(
		.INIT('h8)
	) name1572 (
		\rEIP_reg[0]/NET0131 ,
		_w1109_,
		_w2025_
	);
	LUT4 #(
		.INIT('h3f15)
	) name1573 (
		\InstAddrPointer_reg[0]/NET0131 ,
		\rEIP_reg[0]/NET0131 ,
		_w1109_,
		_w1110_,
		_w2026_
	);
	LUT2 #(
		.INIT('hb)
	) name1574 (
		_w2024_,
		_w2026_,
		_w2027_
	);
	LUT2 #(
		.INIT('h2)
	) name1575 (
		\EAX_reg[26]/NET0131 ,
		_w1825_,
		_w2028_
	);
	LUT4 #(
		.INIT('h8000)
	) name1576 (
		\EAX_reg[19]/NET0131 ,
		_w1837_,
		_w1839_,
		_w1842_,
		_w2029_
	);
	LUT3 #(
		.INIT('h48)
	) name1577 (
		\EAX_reg[26]/NET0131 ,
		_w1848_,
		_w2029_,
		_w2030_
	);
	LUT4 #(
		.INIT('h8000)
	) name1578 (
		\Datai[26]_pad ,
		_w514_,
		_w569_,
		_w612_,
		_w2031_
	);
	LUT2 #(
		.INIT('h2)
	) name1579 (
		\Datai[10]_pad ,
		READY_n_pad,
		_w2032_
	);
	LUT3 #(
		.INIT('h80)
	) name1580 (
		_w566_,
		_w611_,
		_w2032_,
		_w2033_
	);
	LUT4 #(
		.INIT('h02fd)
	) name1581 (
		_w1873_,
		_w1884_,
		_w1895_,
		_w1906_,
		_w2034_
	);
	LUT4 #(
		.INIT('h8000)
	) name1582 (
		_w576_,
		_w579_,
		_w605_,
		_w2034_,
		_w2035_
	);
	LUT3 #(
		.INIT('h01)
	) name1583 (
		_w2033_,
		_w2035_,
		_w2031_,
		_w2036_
	);
	LUT4 #(
		.INIT('h7500)
	) name1584 (
		\EAX_reg[26]/NET0131 ,
		_w635_,
		_w1852_,
		_w2036_,
		_w2037_
	);
	LUT4 #(
		.INIT('hecee)
	) name1585 (
		_w695_,
		_w2028_,
		_w2030_,
		_w2037_,
		_w2038_
	);
	LUT4 #(
		.INIT('hfffc)
	) name1586 (
		\State2_reg[0]/NET0131 ,
		\State2_reg[1]/NET0131 ,
		\State2_reg[2]/NET0131 ,
		\State2_reg[3]/NET0131 ,
		_w2039_
	);
	LUT4 #(
		.INIT('hfc23)
	) name1587 (
		\State2_reg[0]/NET0131 ,
		\State2_reg[1]/NET0131 ,
		\State2_reg[2]/NET0131 ,
		\State2_reg[3]/NET0131 ,
		_w2040_
	);
	LUT2 #(
		.INIT('h2)
	) name1588 (
		\uWord_reg[12]/NET0131 ,
		_w1825_,
		_w2041_
	);
	LUT4 #(
		.INIT('h0001)
	) name1589 (
		\EAX_reg[13]/NET0131 ,
		\EAX_reg[14]/NET0131 ,
		\EAX_reg[15]/NET0131 ,
		\EAX_reg[1]/NET0131 ,
		_w2042_
	);
	LUT4 #(
		.INIT('h0001)
	) name1590 (
		\EAX_reg[0]/NET0131 ,
		\EAX_reg[10]/NET0131 ,
		\EAX_reg[11]/NET0131 ,
		\EAX_reg[12]/NET0131 ,
		_w2043_
	);
	LUT4 #(
		.INIT('h0001)
	) name1591 (
		\EAX_reg[6]/NET0131 ,
		\EAX_reg[7]/NET0131 ,
		\EAX_reg[8]/NET0131 ,
		\EAX_reg[9]/NET0131 ,
		_w2044_
	);
	LUT4 #(
		.INIT('h0001)
	) name1592 (
		\EAX_reg[2]/NET0131 ,
		\EAX_reg[3]/NET0131 ,
		\EAX_reg[4]/NET0131 ,
		\EAX_reg[5]/NET0131 ,
		_w2045_
	);
	LUT4 #(
		.INIT('h8000)
	) name1593 (
		_w2044_,
		_w2045_,
		_w2042_,
		_w2043_,
		_w2046_
	);
	LUT4 #(
		.INIT('h0080)
	) name1594 (
		\EAX_reg[16]/NET0131 ,
		\EAX_reg[17]/NET0131 ,
		\EAX_reg[31]/NET0131 ,
		_w2046_,
		_w2047_
	);
	LUT4 #(
		.INIT('h8000)
	) name1595 (
		\EAX_reg[18]/NET0131 ,
		\EAX_reg[19]/NET0131 ,
		_w1839_,
		_w2047_,
		_w2048_
	);
	LUT2 #(
		.INIT('h8)
	) name1596 (
		_w1841_,
		_w2048_,
		_w2049_
	);
	LUT3 #(
		.INIT('h80)
	) name1597 (
		\EAX_reg[25]/NET0131 ,
		_w1841_,
		_w2048_,
		_w2050_
	);
	LUT4 #(
		.INIT('h8000)
	) name1598 (
		\EAX_reg[25]/NET0131 ,
		\EAX_reg[26]/NET0131 ,
		_w1841_,
		_w2048_,
		_w2051_
	);
	LUT3 #(
		.INIT('h80)
	) name1599 (
		\EAX_reg[27]/NET0131 ,
		\EAX_reg[28]/NET0131 ,
		_w2051_,
		_w2052_
	);
	LUT4 #(
		.INIT('h60c0)
	) name1600 (
		\EAX_reg[27]/NET0131 ,
		\EAX_reg[28]/NET0131 ,
		_w570_,
		_w2051_,
		_w2053_
	);
	LUT2 #(
		.INIT('h8)
	) name1601 (
		\Datai[12]_pad ,
		_w566_,
		_w2054_
	);
	LUT3 #(
		.INIT('h20)
	) name1602 (
		\Datai[12]_pad ,
		READY_n_pad,
		_w566_,
		_w2055_
	);
	LUT3 #(
		.INIT('ha8)
	) name1603 (
		_w611_,
		_w2053_,
		_w2055_,
		_w2056_
	);
	LUT3 #(
		.INIT('he0)
	) name1604 (
		_w566_,
		_w570_,
		_w611_,
		_w2057_
	);
	LUT4 #(
		.INIT('h7400)
	) name1605 (
		READY_n_pad,
		_w566_,
		_w570_,
		_w611_,
		_w2058_
	);
	LUT2 #(
		.INIT('h2)
	) name1606 (
		\uWord_reg[12]/NET0131 ,
		_w2058_,
		_w2059_
	);
	LUT4 #(
		.INIT('heeec)
	) name1607 (
		_w695_,
		_w2041_,
		_w2056_,
		_w2059_,
		_w2060_
	);
	LUT4 #(
		.INIT('hfda0)
	) name1608 (
		\State2_reg[0]/NET0131 ,
		\State2_reg[1]/NET0131 ,
		\State2_reg[2]/NET0131 ,
		\State2_reg[3]/NET0131 ,
		_w2061_
	);
	LUT2 #(
		.INIT('h2)
	) name1609 (
		\InstQueueRd_Addr_reg[0]/NET0131 ,
		_w2061_,
		_w2062_
	);
	LUT3 #(
		.INIT('h72)
	) name1610 (
		\Flush_reg/NET0131 ,
		\InstAddrPointer_reg[0]/NET0131 ,
		\InstQueueRd_Addr_reg[0]/NET0131 ,
		_w2063_
	);
	LUT4 #(
		.INIT('h23af)
	) name1611 (
		\InstQueueRd_Addr_reg[0]/NET0131 ,
		_w712_,
		_w722_,
		_w2063_,
		_w2064_
	);
	LUT2 #(
		.INIT('h4)
	) name1612 (
		_w2062_,
		_w2064_,
		_w2065_
	);
	LUT4 #(
		.INIT('h10ff)
	) name1613 (
		_w629_,
		_w630_,
		_w695_,
		_w2065_,
		_w2066_
	);
	LUT4 #(
		.INIT('h0880)
	) name1614 (
		\Flush_reg/NET0131 ,
		\InstAddrPointer_reg[0]/NET0131 ,
		\InstAddrPointer_reg[1]/NET0131 ,
		\InstAddrPointer_reg[31]/NET0131 ,
		_w2067_
	);
	LUT3 #(
		.INIT('ha8)
	) name1615 (
		_w712_,
		_w713_,
		_w2067_,
		_w2068_
	);
	LUT4 #(
		.INIT('h3f15)
	) name1616 (
		\InstQueueRd_Addr_reg[2]/NET0131 ,
		_w655_,
		_w722_,
		_w2061_,
		_w2069_
	);
	LUT2 #(
		.INIT('h4)
	) name1617 (
		_w2068_,
		_w2069_,
		_w2070_
	);
	LUT4 #(
		.INIT('hb0ff)
	) name1618 (
		_w656_,
		_w671_,
		_w695_,
		_w2070_,
		_w2071_
	);
	LUT2 #(
		.INIT('h2)
	) name1619 (
		\PhyAddrPointer_reg[3]/NET0131 ,
		_w681_,
		_w2072_
	);
	LUT4 #(
		.INIT('h028a)
	) name1620 (
		\PhyAddrPointer_reg[3]/NET0131 ,
		_w573_,
		_w574_,
		_w605_,
		_w2073_
	);
	LUT4 #(
		.INIT('h00fd)
	) name1621 (
		_w688_,
		_w1800_,
		_w1799_,
		_w2073_,
		_w2074_
	);
	LUT4 #(
		.INIT('h5700)
	) name1622 (
		_w574_,
		_w1795_,
		_w2072_,
		_w2074_,
		_w2075_
	);
	LUT3 #(
		.INIT('he0)
	) name1623 (
		\DataWidth_reg[1]/NET0131 ,
		\PhyAddrPointer_reg[1]/NET0131 ,
		\PhyAddrPointer_reg[2]/NET0131 ,
		_w2076_
	);
	LUT4 #(
		.INIT('hfe35)
	) name1624 (
		\State2_reg[0]/NET0131 ,
		\State2_reg[1]/NET0131 ,
		\State2_reg[2]/NET0131 ,
		\State2_reg[3]/NET0131 ,
		_w2077_
	);
	LUT4 #(
		.INIT('h48ea)
	) name1625 (
		\PhyAddrPointer_reg[3]/NET0131 ,
		_w700_,
		_w2076_,
		_w2077_,
		_w2078_
	);
	LUT3 #(
		.INIT('h78)
	) name1626 (
		\PhyAddrPointer_reg[1]/NET0131 ,
		\PhyAddrPointer_reg[2]/NET0131 ,
		\PhyAddrPointer_reg[3]/NET0131 ,
		_w2079_
	);
	LUT2 #(
		.INIT('h8)
	) name1627 (
		_w706_,
		_w2079_,
		_w2080_
	);
	LUT4 #(
		.INIT('h135f)
	) name1628 (
		\PhyAddrPointer_reg[3]/NET0131 ,
		\rEIP_reg[3]/NET0131 ,
		_w718_,
		_w1109_,
		_w2081_
	);
	LUT3 #(
		.INIT('h10)
	) name1629 (
		_w2078_,
		_w2080_,
		_w2081_,
		_w2082_
	);
	LUT3 #(
		.INIT('h2f)
	) name1630 (
		_w695_,
		_w2075_,
		_w2082_,
		_w2083_
	);
	LUT4 #(
		.INIT('h08c8)
	) name1631 (
		\PhyAddrPointer_reg[5]/NET0131 ,
		_w574_,
		_w681_,
		_w1813_,
		_w2084_
	);
	LUT4 #(
		.INIT('h028a)
	) name1632 (
		\PhyAddrPointer_reg[5]/NET0131 ,
		_w573_,
		_w574_,
		_w605_,
		_w2085_
	);
	LUT4 #(
		.INIT('h007d)
	) name1633 (
		_w688_,
		_w1038_,
		_w1815_,
		_w2085_,
		_w2086_
	);
	LUT4 #(
		.INIT('h7f4c)
	) name1634 (
		\PhyAddrPointer_reg[1]/NET0131 ,
		\PhyAddrPointer_reg[5]/NET0131 ,
		_w1258_,
		_w1988_,
		_w2087_
	);
	LUT4 #(
		.INIT('h7f80)
	) name1635 (
		\PhyAddrPointer_reg[2]/NET0131 ,
		\PhyAddrPointer_reg[3]/NET0131 ,
		\PhyAddrPointer_reg[4]/NET0131 ,
		\PhyAddrPointer_reg[5]/NET0131 ,
		_w2088_
	);
	LUT3 #(
		.INIT('hc4)
	) name1636 (
		\DataWidth_reg[1]/NET0131 ,
		_w700_,
		_w2088_,
		_w2089_
	);
	LUT3 #(
		.INIT('he0)
	) name1637 (
		\DataWidth_reg[1]/NET0131 ,
		_w2087_,
		_w2089_,
		_w2090_
	);
	LUT4 #(
		.INIT('h3f15)
	) name1638 (
		\PhyAddrPointer_reg[5]/NET0131 ,
		\rEIP_reg[5]/NET0131 ,
		_w1109_,
		_w1283_,
		_w2091_
	);
	LUT3 #(
		.INIT('h70)
	) name1639 (
		_w706_,
		_w2087_,
		_w2091_,
		_w2092_
	);
	LUT2 #(
		.INIT('h4)
	) name1640 (
		_w2090_,
		_w2092_,
		_w2093_
	);
	LUT4 #(
		.INIT('h8aff)
	) name1641 (
		_w695_,
		_w2084_,
		_w2086_,
		_w2093_,
		_w2094_
	);
	LUT2 #(
		.INIT('h2)
	) name1642 (
		\PhyAddrPointer_reg[6]/NET0131 ,
		_w681_,
		_w2095_
	);
	LUT4 #(
		.INIT('haa20)
	) name1643 (
		_w574_,
		_w1739_,
		_w1741_,
		_w2095_,
		_w2096_
	);
	LUT4 #(
		.INIT('h028a)
	) name1644 (
		\PhyAddrPointer_reg[6]/NET0131 ,
		_w573_,
		_w574_,
		_w605_,
		_w2097_
	);
	LUT2 #(
		.INIT('h1)
	) name1645 (
		_w1744_,
		_w2097_,
		_w2098_
	);
	LUT4 #(
		.INIT('h8848)
	) name1646 (
		\PhyAddrPointer_reg[6]/NET0131 ,
		_w700_,
		_w1259_,
		_w1453_,
		_w2099_
	);
	LUT3 #(
		.INIT('h6c)
	) name1647 (
		\PhyAddrPointer_reg[1]/NET0131 ,
		\PhyAddrPointer_reg[6]/NET0131 ,
		_w1259_,
		_w2100_
	);
	LUT4 #(
		.INIT('h60c0)
	) name1648 (
		\PhyAddrPointer_reg[1]/NET0131 ,
		\PhyAddrPointer_reg[6]/NET0131 ,
		_w706_,
		_w1259_,
		_w2101_
	);
	LUT4 #(
		.INIT('h3f15)
	) name1649 (
		\PhyAddrPointer_reg[6]/NET0131 ,
		\rEIP_reg[6]/NET0131 ,
		_w1109_,
		_w1283_,
		_w2102_
	);
	LUT3 #(
		.INIT('h10)
	) name1650 (
		_w2101_,
		_w2099_,
		_w2102_,
		_w2103_
	);
	LUT4 #(
		.INIT('h8aff)
	) name1651 (
		_w695_,
		_w2096_,
		_w2098_,
		_w2103_,
		_w2104_
	);
	LUT3 #(
		.INIT('h8a)
	) name1652 (
		\InstAddrPointer_reg[1]/NET0131 ,
		_w682_,
		_w1220_,
		_w2105_
	);
	LUT4 #(
		.INIT('hfb00)
	) name1653 (
		_w582_,
		_w595_,
		_w606_,
		_w954_,
		_w2106_
	);
	LUT4 #(
		.INIT('h807f)
	) name1654 (
		_w770_,
		_w776_,
		_w779_,
		_w954_,
		_w2107_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name1655 (
		\InstAddrPointer_reg[1]/NET0131 ,
		_w770_,
		_w776_,
		_w779_,
		_w2108_
	);
	LUT4 #(
		.INIT('h4051)
	) name1656 (
		_w844_,
		_w952_,
		_w2108_,
		_w2107_,
		_w2109_
	);
	LUT3 #(
		.INIT('h28)
	) name1657 (
		_w844_,
		_w793_,
		_w2108_,
		_w2110_
	);
	LUT4 #(
		.INIT('h8880)
	) name1658 (
		_w574_,
		_w681_,
		_w2109_,
		_w2110_,
		_w2111_
	);
	LUT2 #(
		.INIT('h2)
	) name1659 (
		_w1033_,
		_w2108_,
		_w2112_
	);
	LUT2 #(
		.INIT('h1)
	) name1660 (
		_w1033_,
		_w2107_,
		_w2113_
	);
	LUT4 #(
		.INIT('h0008)
	) name1661 (
		_w573_,
		_w605_,
		_w2113_,
		_w2112_,
		_w2114_
	);
	LUT2 #(
		.INIT('h1)
	) name1662 (
		_w2111_,
		_w2114_,
		_w2115_
	);
	LUT3 #(
		.INIT('he0)
	) name1663 (
		\InstAddrPointer_reg[1]/NET0131 ,
		_w645_,
		_w2115_,
		_w2116_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name1664 (
		_w695_,
		_w2106_,
		_w2105_,
		_w2116_,
		_w2117_
	);
	LUT2 #(
		.INIT('h8)
	) name1665 (
		\rEIP_reg[1]/NET0131 ,
		_w1109_,
		_w2118_
	);
	LUT4 #(
		.INIT('h3f15)
	) name1666 (
		\InstAddrPointer_reg[1]/NET0131 ,
		\rEIP_reg[1]/NET0131 ,
		_w1109_,
		_w1110_,
		_w2119_
	);
	LUT2 #(
		.INIT('hb)
	) name1667 (
		_w2117_,
		_w2119_,
		_w2120_
	);
	LUT2 #(
		.INIT('h4)
	) name1668 (
		\Flush_reg/NET0131 ,
		\InstQueueRd_Addr_reg[1]/NET0131 ,
		_w2121_
	);
	LUT4 #(
		.INIT('h8008)
	) name1669 (
		\Flush_reg/NET0131 ,
		\InstAddrPointer_reg[0]/NET0131 ,
		\InstAddrPointer_reg[1]/NET0131 ,
		\InstAddrPointer_reg[31]/NET0131 ,
		_w2122_
	);
	LUT3 #(
		.INIT('ha8)
	) name1670 (
		_w712_,
		_w2121_,
		_w2122_,
		_w2123_
	);
	LUT4 #(
		.INIT('h9f13)
	) name1671 (
		\InstQueueRd_Addr_reg[0]/NET0131 ,
		\InstQueueRd_Addr_reg[1]/NET0131 ,
		_w722_,
		_w2061_,
		_w2124_
	);
	LUT2 #(
		.INIT('h4)
	) name1672 (
		_w2123_,
		_w2124_,
		_w2125_
	);
	LUT4 #(
		.INIT('he0ff)
	) name1673 (
		_w608_,
		_w627_,
		_w695_,
		_w2125_,
		_w2126_
	);
	LUT2 #(
		.INIT('h2)
	) name1674 (
		\EAX_reg[29]/NET0131 ,
		_w1825_,
		_w2127_
	);
	LUT4 #(
		.INIT('hb300)
	) name1675 (
		\EAX_reg[28]/NET0131 ,
		_w1848_,
		_w1845_,
		_w1852_,
		_w2128_
	);
	LUT2 #(
		.INIT('h4)
	) name1676 (
		\EAX_reg[29]/NET0131 ,
		_w1848_,
		_w2129_
	);
	LUT4 #(
		.INIT('h02fd)
	) name1677 (
		_w1907_,
		_w1918_,
		_w1929_,
		_w1940_,
		_w2130_
	);
	LUT3 #(
		.INIT('h20)
	) name1678 (
		\Datai[13]_pad ,
		READY_n_pad,
		_w611_,
		_w2131_
	);
	LUT2 #(
		.INIT('h8)
	) name1679 (
		_w566_,
		_w2131_,
		_w2132_
	);
	LUT3 #(
		.INIT('h10)
	) name1680 (
		\Datai[29]_pad ,
		READY_n_pad,
		_w611_,
		_w2133_
	);
	LUT3 #(
		.INIT('h45)
	) name1681 (
		\EAX_reg[29]/NET0131 ,
		READY_n_pad,
		_w611_,
		_w2134_
	);
	LUT4 #(
		.INIT('h0008)
	) name1682 (
		_w514_,
		_w569_,
		_w2134_,
		_w2133_,
		_w2135_
	);
	LUT4 #(
		.INIT('h0007)
	) name1683 (
		_w1849_,
		_w2130_,
		_w2132_,
		_w2135_,
		_w2136_
	);
	LUT4 #(
		.INIT('h7f00)
	) name1684 (
		\EAX_reg[28]/NET0131 ,
		_w1845_,
		_w2129_,
		_w2136_,
		_w2137_
	);
	LUT4 #(
		.INIT('h08cc)
	) name1685 (
		\EAX_reg[29]/NET0131 ,
		_w695_,
		_w2128_,
		_w2137_,
		_w2138_
	);
	LUT2 #(
		.INIT('he)
	) name1686 (
		_w2127_,
		_w2138_,
		_w2139_
	);
	LUT4 #(
		.INIT('h8000)
	) name1687 (
		\EBX_reg[16]/NET0131 ,
		\EBX_reg[17]/NET0131 ,
		\EBX_reg[18]/NET0131 ,
		_w1968_,
		_w2140_
	);
	LUT4 #(
		.INIT('h8000)
	) name1688 (
		\EBX_reg[20]/NET0131 ,
		\EBX_reg[21]/NET0131 ,
		\EBX_reg[22]/NET0131 ,
		\EBX_reg[23]/NET0131 ,
		_w2141_
	);
	LUT3 #(
		.INIT('h80)
	) name1689 (
		\EBX_reg[19]/NET0131 ,
		_w2140_,
		_w2141_,
		_w2142_
	);
	LUT4 #(
		.INIT('h8000)
	) name1690 (
		\EBX_reg[19]/NET0131 ,
		\EBX_reg[24]/NET0131 ,
		_w2140_,
		_w2141_,
		_w2143_
	);
	LUT4 #(
		.INIT('h60c0)
	) name1691 (
		\EBX_reg[25]/NET0131 ,
		\EBX_reg[26]/NET0131 ,
		_w590_,
		_w2143_,
		_w2144_
	);
	LUT4 #(
		.INIT('h8000)
	) name1692 (
		_w552_,
		_w576_,
		_w605_,
		_w2034_,
		_w2145_
	);
	LUT3 #(
		.INIT('h07)
	) name1693 (
		\EBX_reg[26]/NET0131 ,
		_w1975_,
		_w2145_,
		_w2146_
	);
	LUT2 #(
		.INIT('h2)
	) name1694 (
		\EBX_reg[26]/NET0131 ,
		_w1825_,
		_w2147_
	);
	LUT4 #(
		.INIT('hff8a)
	) name1695 (
		_w695_,
		_w2144_,
		_w2146_,
		_w2147_,
		_w2148_
	);
	LUT2 #(
		.INIT('h8)
	) name1696 (
		_w570_,
		_w611_,
		_w2149_
	);
	LUT3 #(
		.INIT('h6c)
	) name1697 (
		\EAX_reg[23]/NET0131 ,
		\EAX_reg[24]/NET0131 ,
		_w2048_,
		_w2150_
	);
	LUT4 #(
		.INIT('h0903)
	) name1698 (
		\EAX_reg[23]/NET0131 ,
		\EAX_reg[24]/NET0131 ,
		_w617_,
		_w2048_,
		_w2151_
	);
	LUT3 #(
		.INIT('h08)
	) name1699 (
		_w570_,
		_w611_,
		_w2151_,
		_w2152_
	);
	LUT4 #(
		.INIT('hf400)
	) name1700 (
		_w514_,
		_w569_,
		_w570_,
		_w611_,
		_w2153_
	);
	LUT3 #(
		.INIT('h40)
	) name1701 (
		_w514_,
		_w569_,
		_w617_,
		_w2154_
	);
	LUT2 #(
		.INIT('h2)
	) name1702 (
		_w2153_,
		_w2154_,
		_w2155_
	);
	LUT4 #(
		.INIT('haa8a)
	) name1703 (
		\Datao[24]_pad ,
		_w2152_,
		_w2153_,
		_w2154_,
		_w2156_
	);
	LUT2 #(
		.INIT('h8)
	) name1704 (
		_w570_,
		_w2150_,
		_w2157_
	);
	LUT3 #(
		.INIT('h80)
	) name1705 (
		_w570_,
		_w659_,
		_w2150_,
		_w2158_
	);
	LUT4 #(
		.INIT('hfc60)
	) name1706 (
		\State2_reg[0]/NET0131 ,
		\State2_reg[1]/NET0131 ,
		\State2_reg[2]/NET0131 ,
		\State2_reg[3]/NET0131 ,
		_w2159_
	);
	LUT4 #(
		.INIT('h3f15)
	) name1707 (
		\Datao[24]_pad ,
		\uWord_reg[8]/NET0131 ,
		_w696_,
		_w2159_,
		_w2160_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name1708 (
		_w695_,
		_w2156_,
		_w2158_,
		_w2160_,
		_w2161_
	);
	LUT4 #(
		.INIT('h0903)
	) name1709 (
		\EAX_reg[27]/NET0131 ,
		\EAX_reg[28]/NET0131 ,
		_w617_,
		_w2051_,
		_w2162_
	);
	LUT4 #(
		.INIT('h0c04)
	) name1710 (
		_w2149_,
		_w2153_,
		_w2154_,
		_w2162_,
		_w2163_
	);
	LUT2 #(
		.INIT('h8)
	) name1711 (
		_w659_,
		_w2053_,
		_w2164_
	);
	LUT4 #(
		.INIT('hcc08)
	) name1712 (
		\Datao[28]_pad ,
		_w695_,
		_w2163_,
		_w2164_,
		_w2165_
	);
	LUT4 #(
		.INIT('h3f15)
	) name1713 (
		\Datao[28]_pad ,
		\uWord_reg[12]/NET0131 ,
		_w696_,
		_w2159_,
		_w2166_
	);
	LUT2 #(
		.INIT('hb)
	) name1714 (
		_w2165_,
		_w2166_,
		_w2167_
	);
	LUT4 #(
		.INIT('hef00)
	) name1715 (
		_w647_,
		_w642_,
		_w651_,
		_w695_,
		_w2168_
	);
	LUT2 #(
		.INIT('h4)
	) name1716 (
		\Flush_reg/NET0131 ,
		\InstQueueRd_Addr_reg[3]/NET0131 ,
		_w2169_
	);
	LUT3 #(
		.INIT('ha8)
	) name1717 (
		_w712_,
		_w2067_,
		_w2169_,
		_w2170_
	);
	LUT4 #(
		.INIT('hcf45)
	) name1718 (
		\InstQueueRd_Addr_reg[3]/NET0131 ,
		_w648_,
		_w722_,
		_w2061_,
		_w2171_
	);
	LUT2 #(
		.INIT('h4)
	) name1719 (
		_w2170_,
		_w2171_,
		_w2172_
	);
	LUT2 #(
		.INIT('hb)
	) name1720 (
		_w2168_,
		_w2172_,
		_w2173_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name1721 (
		\uWord_reg[8]/NET0131 ,
		_w695_,
		_w1825_,
		_w2058_,
		_w2174_
	);
	LUT2 #(
		.INIT('h8)
	) name1722 (
		_w611_,
		_w695_,
		_w2175_
	);
	LUT2 #(
		.INIT('h8)
	) name1723 (
		\Datai[8]_pad ,
		_w566_,
		_w2176_
	);
	LUT3 #(
		.INIT('h20)
	) name1724 (
		\Datai[8]_pad ,
		READY_n_pad,
		_w566_,
		_w2177_
	);
	LUT3 #(
		.INIT('hc8)
	) name1725 (
		_w2157_,
		_w2175_,
		_w2177_,
		_w2178_
	);
	LUT2 #(
		.INIT('he)
	) name1726 (
		_w2174_,
		_w2178_,
		_w2179_
	);
	LUT2 #(
		.INIT('h8)
	) name1727 (
		\EBX_reg[27]/NET0131 ,
		\EBX_reg[28]/NET0131 ,
		_w2180_
	);
	LUT3 #(
		.INIT('h80)
	) name1728 (
		_w1958_,
		_w1972_,
		_w2180_,
		_w2181_
	);
	LUT4 #(
		.INIT('h31fd)
	) name1729 (
		\EBX_reg[29]/NET0131 ,
		_w1973_,
		_w1974_,
		_w2130_,
		_w2182_
	);
	LUT4 #(
		.INIT('hb700)
	) name1730 (
		\EBX_reg[29]/NET0131 ,
		_w590_,
		_w2181_,
		_w2182_,
		_w2183_
	);
	LUT2 #(
		.INIT('h2)
	) name1731 (
		\EBX_reg[29]/NET0131 ,
		_w1825_,
		_w2184_
	);
	LUT3 #(
		.INIT('hf2)
	) name1732 (
		_w695_,
		_w2183_,
		_w2184_,
		_w2185_
	);
	LUT3 #(
		.INIT('h20)
	) name1733 (
		\InstQueueWr_Addr_reg[0]/NET0131 ,
		\InstQueueWr_Addr_reg[1]/NET0131 ,
		\InstQueueWr_Addr_reg[2]/NET0131 ,
		_w2186_
	);
	LUT4 #(
		.INIT('h2000)
	) name1734 (
		\InstQueueWr_Addr_reg[0]/NET0131 ,
		\InstQueueWr_Addr_reg[1]/NET0131 ,
		\InstQueueWr_Addr_reg[2]/NET0131 ,
		\InstQueueWr_Addr_reg[3]/NET0131 ,
		_w2187_
	);
	LUT4 #(
		.INIT('h0001)
	) name1735 (
		\Datai[13]_pad ,
		\Datai[14]_pad ,
		\Datai[15]_pad ,
		\Datai[1]_pad ,
		_w2188_
	);
	LUT4 #(
		.INIT('h0001)
	) name1736 (
		\Datai[0]_pad ,
		\Datai[10]_pad ,
		\Datai[11]_pad ,
		\Datai[12]_pad ,
		_w2189_
	);
	LUT4 #(
		.INIT('h0001)
	) name1737 (
		\Datai[6]_pad ,
		\Datai[7]_pad ,
		\Datai[8]_pad ,
		\Datai[9]_pad ,
		_w2190_
	);
	LUT4 #(
		.INIT('h0001)
	) name1738 (
		\Datai[2]_pad ,
		\Datai[3]_pad ,
		\Datai[4]_pad ,
		\Datai[5]_pad ,
		_w2191_
	);
	LUT4 #(
		.INIT('h8000)
	) name1739 (
		_w2190_,
		_w2191_,
		_w2188_,
		_w2189_,
		_w2192_
	);
	LUT4 #(
		.INIT('h0001)
	) name1740 (
		\Datai[20]_pad ,
		\Datai[21]_pad ,
		\Datai[22]_pad ,
		\Datai[23]_pad ,
		_w2193_
	);
	LUT4 #(
		.INIT('h0001)
	) name1741 (
		\Datai[16]_pad ,
		\Datai[17]_pad ,
		\Datai[18]_pad ,
		\Datai[19]_pad ,
		_w2194_
	);
	LUT2 #(
		.INIT('h8)
	) name1742 (
		_w2193_,
		_w2194_,
		_w2195_
	);
	LUT4 #(
		.INIT('h0888)
	) name1743 (
		\Datai[24]_pad ,
		\Datai[31]_pad ,
		_w2192_,
		_w2195_,
		_w2196_
	);
	LUT4 #(
		.INIT('h8000)
	) name1744 (
		\Datai[25]_pad ,
		\Datai[26]_pad ,
		\Datai[27]_pad ,
		_w2196_,
		_w2197_
	);
	LUT3 #(
		.INIT('h48)
	) name1745 (
		\Datai[28]_pad ,
		_w2187_,
		_w2197_,
		_w2198_
	);
	LUT4 #(
		.INIT('h0080)
	) name1746 (
		\Datai[16]_pad ,
		\Datai[17]_pad ,
		\Datai[31]_pad ,
		_w2192_,
		_w2199_
	);
	LUT4 #(
		.INIT('h8000)
	) name1747 (
		\Datai[18]_pad ,
		\Datai[19]_pad ,
		\Datai[20]_pad ,
		_w2199_,
		_w2200_
	);
	LUT4 #(
		.INIT('h78f0)
	) name1748 (
		\Datai[18]_pad ,
		\Datai[19]_pad ,
		\Datai[20]_pad ,
		_w2199_,
		_w2201_
	);
	LUT2 #(
		.INIT('h4)
	) name1749 (
		\InstQueueWr_Addr_reg[0]/NET0131 ,
		\InstQueueWr_Addr_reg[1]/NET0131 ,
		_w2202_
	);
	LUT4 #(
		.INIT('h4000)
	) name1750 (
		\InstQueueWr_Addr_reg[0]/NET0131 ,
		\InstQueueWr_Addr_reg[1]/NET0131 ,
		\InstQueueWr_Addr_reg[2]/NET0131 ,
		\InstQueueWr_Addr_reg[3]/NET0131 ,
		_w2203_
	);
	LUT2 #(
		.INIT('h8)
	) name1751 (
		_w2201_,
		_w2203_,
		_w2204_
	);
	LUT4 #(
		.INIT('h0001)
	) name1752 (
		\InstQueueWr_Addr_reg[0]/NET0131 ,
		\InstQueueWr_Addr_reg[1]/NET0131 ,
		\InstQueueWr_Addr_reg[2]/NET0131 ,
		\InstQueueWr_Addr_reg[3]/NET0131 ,
		_w2205_
	);
	LUT3 #(
		.INIT('h80)
	) name1753 (
		\InstQueueWr_Addr_reg[0]/NET0131 ,
		\InstQueueWr_Addr_reg[1]/NET0131 ,
		\InstQueueWr_Addr_reg[2]/NET0131 ,
		_w2206_
	);
	LUT4 #(
		.INIT('h8000)
	) name1754 (
		\InstQueueWr_Addr_reg[0]/NET0131 ,
		\InstQueueWr_Addr_reg[1]/NET0131 ,
		\InstQueueWr_Addr_reg[2]/NET0131 ,
		\InstQueueWr_Addr_reg[3]/NET0131 ,
		_w2207_
	);
	LUT4 #(
		.INIT('h7ffe)
	) name1755 (
		\InstQueueWr_Addr_reg[0]/NET0131 ,
		\InstQueueWr_Addr_reg[1]/NET0131 ,
		\InstQueueWr_Addr_reg[2]/NET0131 ,
		\InstQueueWr_Addr_reg[3]/NET0131 ,
		_w2208_
	);
	LUT4 #(
		.INIT('h5553)
	) name1756 (
		\Datai[4]_pad ,
		\InstQueue_reg[0][4]/NET0131 ,
		_w2205_,
		_w2207_,
		_w2209_
	);
	LUT4 #(
		.INIT('h9fff)
	) name1757 (
		\InstQueueWr_Addr_reg[0]/NET0131 ,
		\InstQueueWr_Addr_reg[1]/NET0131 ,
		\InstQueueWr_Addr_reg[2]/NET0131 ,
		\InstQueueWr_Addr_reg[3]/NET0131 ,
		_w2210_
	);
	LUT2 #(
		.INIT('h2)
	) name1758 (
		\DataWidth_reg[1]/NET0131 ,
		_w2210_,
		_w2211_
	);
	LUT2 #(
		.INIT('h1)
	) name1759 (
		_w2209_,
		_w2211_,
		_w2212_
	);
	LUT4 #(
		.INIT('h0057)
	) name1760 (
		\DataWidth_reg[1]/NET0131 ,
		_w2198_,
		_w2204_,
		_w2212_,
		_w2213_
	);
	LUT4 #(
		.INIT('hc055)
	) name1761 (
		\InstQueue_reg[0][4]/NET0131 ,
		_w558_,
		_w563_,
		_w2205_,
		_w2214_
	);
	LUT4 #(
		.INIT('hfd14)
	) name1762 (
		\State2_reg[0]/NET0131 ,
		\State2_reg[1]/NET0131 ,
		\State2_reg[2]/NET0131 ,
		\State2_reg[3]/NET0131 ,
		_w2215_
	);
	LUT2 #(
		.INIT('h2)
	) name1763 (
		\InstQueue_reg[0][4]/NET0131 ,
		_w2215_,
		_w2216_
	);
	LUT3 #(
		.INIT('h0d)
	) name1764 (
		_w706_,
		_w2209_,
		_w2216_,
		_w2217_
	);
	LUT3 #(
		.INIT('hd0)
	) name1765 (
		_w722_,
		_w2214_,
		_w2217_,
		_w2218_
	);
	LUT3 #(
		.INIT('h2f)
	) name1766 (
		_w700_,
		_w2213_,
		_w2218_,
		_w2219_
	);
	LUT4 #(
		.INIT('h0080)
	) name1767 (
		\InstQueueWr_Addr_reg[0]/NET0131 ,
		\InstQueueWr_Addr_reg[1]/NET0131 ,
		\InstQueueWr_Addr_reg[2]/NET0131 ,
		\InstQueueWr_Addr_reg[3]/NET0131 ,
		_w2220_
	);
	LUT3 #(
		.INIT('h60)
	) name1768 (
		\Datai[28]_pad ,
		_w2197_,
		_w2220_,
		_w2221_
	);
	LUT4 #(
		.INIT('h0100)
	) name1769 (
		\InstQueueWr_Addr_reg[0]/NET0131 ,
		\InstQueueWr_Addr_reg[1]/NET0131 ,
		\InstQueueWr_Addr_reg[2]/NET0131 ,
		\InstQueueWr_Addr_reg[3]/NET0131 ,
		_w2222_
	);
	LUT2 #(
		.INIT('h8)
	) name1770 (
		_w2201_,
		_w2222_,
		_w2223_
	);
	LUT4 #(
		.INIT('h0400)
	) name1771 (
		\InstQueueWr_Addr_reg[0]/NET0131 ,
		\InstQueueWr_Addr_reg[1]/NET0131 ,
		\InstQueueWr_Addr_reg[2]/NET0131 ,
		\InstQueueWr_Addr_reg[3]/NET0131 ,
		_w2224_
	);
	LUT4 #(
		.INIT('h0200)
	) name1772 (
		\InstQueueWr_Addr_reg[0]/NET0131 ,
		\InstQueueWr_Addr_reg[1]/NET0131 ,
		\InstQueueWr_Addr_reg[2]/NET0131 ,
		\InstQueueWr_Addr_reg[3]/NET0131 ,
		_w2225_
	);
	LUT4 #(
		.INIT('hf9ff)
	) name1773 (
		\InstQueueWr_Addr_reg[0]/NET0131 ,
		\InstQueueWr_Addr_reg[1]/NET0131 ,
		\InstQueueWr_Addr_reg[2]/NET0131 ,
		\InstQueueWr_Addr_reg[3]/NET0131 ,
		_w2226_
	);
	LUT4 #(
		.INIT('h5553)
	) name1774 (
		\Datai[4]_pad ,
		\InstQueue_reg[10][4]/NET0131 ,
		_w2224_,
		_w2225_,
		_w2227_
	);
	LUT4 #(
		.INIT('hfe7f)
	) name1775 (
		\InstQueueWr_Addr_reg[0]/NET0131 ,
		\InstQueueWr_Addr_reg[1]/NET0131 ,
		\InstQueueWr_Addr_reg[2]/NET0131 ,
		\InstQueueWr_Addr_reg[3]/NET0131 ,
		_w2228_
	);
	LUT2 #(
		.INIT('h2)
	) name1776 (
		\DataWidth_reg[1]/NET0131 ,
		_w2228_,
		_w2229_
	);
	LUT2 #(
		.INIT('h1)
	) name1777 (
		_w2227_,
		_w2229_,
		_w2230_
	);
	LUT4 #(
		.INIT('h0057)
	) name1778 (
		\DataWidth_reg[1]/NET0131 ,
		_w2221_,
		_w2223_,
		_w2230_,
		_w2231_
	);
	LUT4 #(
		.INIT('hc055)
	) name1779 (
		\InstQueue_reg[10][4]/NET0131 ,
		_w558_,
		_w563_,
		_w2224_,
		_w2232_
	);
	LUT2 #(
		.INIT('h2)
	) name1780 (
		\InstQueue_reg[10][4]/NET0131 ,
		_w2215_,
		_w2233_
	);
	LUT3 #(
		.INIT('h0d)
	) name1781 (
		_w706_,
		_w2227_,
		_w2233_,
		_w2234_
	);
	LUT3 #(
		.INIT('hd0)
	) name1782 (
		_w722_,
		_w2232_,
		_w2234_,
		_w2235_
	);
	LUT3 #(
		.INIT('h2f)
	) name1783 (
		_w700_,
		_w2231_,
		_w2235_,
		_w2236_
	);
	LUT3 #(
		.INIT('h60)
	) name1784 (
		\Datai[28]_pad ,
		_w2197_,
		_w2222_,
		_w2237_
	);
	LUT2 #(
		.INIT('h8)
	) name1785 (
		_w2201_,
		_w2225_,
		_w2238_
	);
	LUT4 #(
		.INIT('h0800)
	) name1786 (
		\InstQueueWr_Addr_reg[0]/NET0131 ,
		\InstQueueWr_Addr_reg[1]/NET0131 ,
		\InstQueueWr_Addr_reg[2]/NET0131 ,
		\InstQueueWr_Addr_reg[3]/NET0131 ,
		_w2239_
	);
	LUT4 #(
		.INIT('hf3ff)
	) name1787 (
		\InstQueueWr_Addr_reg[0]/NET0131 ,
		\InstQueueWr_Addr_reg[1]/NET0131 ,
		\InstQueueWr_Addr_reg[2]/NET0131 ,
		\InstQueueWr_Addr_reg[3]/NET0131 ,
		_w2240_
	);
	LUT4 #(
		.INIT('h5553)
	) name1788 (
		\Datai[4]_pad ,
		\InstQueue_reg[11][4]/NET0131 ,
		_w2224_,
		_w2239_,
		_w2241_
	);
	LUT4 #(
		.INIT('hfcff)
	) name1789 (
		\InstQueueWr_Addr_reg[0]/NET0131 ,
		\InstQueueWr_Addr_reg[1]/NET0131 ,
		\InstQueueWr_Addr_reg[2]/NET0131 ,
		\InstQueueWr_Addr_reg[3]/NET0131 ,
		_w2242_
	);
	LUT2 #(
		.INIT('h2)
	) name1790 (
		\DataWidth_reg[1]/NET0131 ,
		_w2242_,
		_w2243_
	);
	LUT2 #(
		.INIT('h1)
	) name1791 (
		_w2241_,
		_w2243_,
		_w2244_
	);
	LUT4 #(
		.INIT('h0057)
	) name1792 (
		\DataWidth_reg[1]/NET0131 ,
		_w2237_,
		_w2238_,
		_w2244_,
		_w2245_
	);
	LUT4 #(
		.INIT('hc055)
	) name1793 (
		\InstQueue_reg[11][4]/NET0131 ,
		_w558_,
		_w563_,
		_w2239_,
		_w2246_
	);
	LUT2 #(
		.INIT('h2)
	) name1794 (
		\InstQueue_reg[11][4]/NET0131 ,
		_w2215_,
		_w2247_
	);
	LUT3 #(
		.INIT('h0d)
	) name1795 (
		_w706_,
		_w2241_,
		_w2247_,
		_w2248_
	);
	LUT3 #(
		.INIT('hd0)
	) name1796 (
		_w722_,
		_w2246_,
		_w2248_,
		_w2249_
	);
	LUT3 #(
		.INIT('h2f)
	) name1797 (
		_w700_,
		_w2245_,
		_w2249_,
		_w2250_
	);
	LUT3 #(
		.INIT('h60)
	) name1798 (
		\Datai[28]_pad ,
		_w2197_,
		_w2225_,
		_w2251_
	);
	LUT2 #(
		.INIT('h8)
	) name1799 (
		_w2201_,
		_w2224_,
		_w2252_
	);
	LUT4 #(
		.INIT('h1000)
	) name1800 (
		\InstQueueWr_Addr_reg[0]/NET0131 ,
		\InstQueueWr_Addr_reg[1]/NET0131 ,
		\InstQueueWr_Addr_reg[2]/NET0131 ,
		\InstQueueWr_Addr_reg[3]/NET0131 ,
		_w2253_
	);
	LUT4 #(
		.INIT('he7ff)
	) name1801 (
		\InstQueueWr_Addr_reg[0]/NET0131 ,
		\InstQueueWr_Addr_reg[1]/NET0131 ,
		\InstQueueWr_Addr_reg[2]/NET0131 ,
		\InstQueueWr_Addr_reg[3]/NET0131 ,
		_w2254_
	);
	LUT4 #(
		.INIT('h5553)
	) name1802 (
		\Datai[4]_pad ,
		\InstQueue_reg[12][4]/NET0131 ,
		_w2239_,
		_w2253_,
		_w2255_
	);
	LUT2 #(
		.INIT('h2)
	) name1803 (
		\DataWidth_reg[1]/NET0131 ,
		_w2226_,
		_w2256_
	);
	LUT2 #(
		.INIT('h1)
	) name1804 (
		_w2255_,
		_w2256_,
		_w2257_
	);
	LUT4 #(
		.INIT('h0057)
	) name1805 (
		\DataWidth_reg[1]/NET0131 ,
		_w2251_,
		_w2252_,
		_w2257_,
		_w2258_
	);
	LUT4 #(
		.INIT('hc055)
	) name1806 (
		\InstQueue_reg[12][4]/NET0131 ,
		_w558_,
		_w563_,
		_w2253_,
		_w2259_
	);
	LUT2 #(
		.INIT('h2)
	) name1807 (
		\InstQueue_reg[12][4]/NET0131 ,
		_w2215_,
		_w2260_
	);
	LUT3 #(
		.INIT('h0d)
	) name1808 (
		_w706_,
		_w2255_,
		_w2260_,
		_w2261_
	);
	LUT3 #(
		.INIT('hd0)
	) name1809 (
		_w722_,
		_w2259_,
		_w2261_,
		_w2262_
	);
	LUT3 #(
		.INIT('h2f)
	) name1810 (
		_w700_,
		_w2258_,
		_w2262_,
		_w2263_
	);
	LUT3 #(
		.INIT('h60)
	) name1811 (
		\Datai[28]_pad ,
		_w2197_,
		_w2224_,
		_w2264_
	);
	LUT2 #(
		.INIT('h8)
	) name1812 (
		_w2201_,
		_w2239_,
		_w2265_
	);
	LUT4 #(
		.INIT('hcfff)
	) name1813 (
		\InstQueueWr_Addr_reg[0]/NET0131 ,
		\InstQueueWr_Addr_reg[1]/NET0131 ,
		\InstQueueWr_Addr_reg[2]/NET0131 ,
		\InstQueueWr_Addr_reg[3]/NET0131 ,
		_w2266_
	);
	LUT4 #(
		.INIT('h5553)
	) name1814 (
		\Datai[4]_pad ,
		\InstQueue_reg[13][4]/NET0131 ,
		_w2187_,
		_w2253_,
		_w2267_
	);
	LUT2 #(
		.INIT('h2)
	) name1815 (
		\DataWidth_reg[1]/NET0131 ,
		_w2240_,
		_w2268_
	);
	LUT2 #(
		.INIT('h1)
	) name1816 (
		_w2267_,
		_w2268_,
		_w2269_
	);
	LUT4 #(
		.INIT('h0057)
	) name1817 (
		\DataWidth_reg[1]/NET0131 ,
		_w2264_,
		_w2265_,
		_w2269_,
		_w2270_
	);
	LUT4 #(
		.INIT('hc055)
	) name1818 (
		\InstQueue_reg[13][4]/NET0131 ,
		_w558_,
		_w563_,
		_w2187_,
		_w2271_
	);
	LUT2 #(
		.INIT('h2)
	) name1819 (
		\InstQueue_reg[13][4]/NET0131 ,
		_w2215_,
		_w2272_
	);
	LUT3 #(
		.INIT('h0d)
	) name1820 (
		_w706_,
		_w2267_,
		_w2272_,
		_w2273_
	);
	LUT3 #(
		.INIT('hd0)
	) name1821 (
		_w722_,
		_w2271_,
		_w2273_,
		_w2274_
	);
	LUT3 #(
		.INIT('h2f)
	) name1822 (
		_w700_,
		_w2270_,
		_w2274_,
		_w2275_
	);
	LUT3 #(
		.INIT('h60)
	) name1823 (
		\Datai[28]_pad ,
		_w2197_,
		_w2239_,
		_w2276_
	);
	LUT2 #(
		.INIT('h8)
	) name1824 (
		_w2201_,
		_w2253_,
		_w2277_
	);
	LUT4 #(
		.INIT('h5553)
	) name1825 (
		\Datai[4]_pad ,
		\InstQueue_reg[14][4]/NET0131 ,
		_w2187_,
		_w2203_,
		_w2278_
	);
	LUT2 #(
		.INIT('h2)
	) name1826 (
		\DataWidth_reg[1]/NET0131 ,
		_w2254_,
		_w2279_
	);
	LUT2 #(
		.INIT('h1)
	) name1827 (
		_w2278_,
		_w2279_,
		_w2280_
	);
	LUT4 #(
		.INIT('h0057)
	) name1828 (
		\DataWidth_reg[1]/NET0131 ,
		_w2276_,
		_w2277_,
		_w2280_,
		_w2281_
	);
	LUT4 #(
		.INIT('hc055)
	) name1829 (
		\InstQueue_reg[14][4]/NET0131 ,
		_w558_,
		_w563_,
		_w2203_,
		_w2282_
	);
	LUT2 #(
		.INIT('h2)
	) name1830 (
		\InstQueue_reg[14][4]/NET0131 ,
		_w2215_,
		_w2283_
	);
	LUT3 #(
		.INIT('h0d)
	) name1831 (
		_w706_,
		_w2278_,
		_w2283_,
		_w2284_
	);
	LUT3 #(
		.INIT('hd0)
	) name1832 (
		_w722_,
		_w2282_,
		_w2284_,
		_w2285_
	);
	LUT3 #(
		.INIT('h2f)
	) name1833 (
		_w700_,
		_w2281_,
		_w2285_,
		_w2286_
	);
	LUT3 #(
		.INIT('h60)
	) name1834 (
		\Datai[28]_pad ,
		_w2197_,
		_w2253_,
		_w2287_
	);
	LUT2 #(
		.INIT('h8)
	) name1835 (
		_w2187_,
		_w2201_,
		_w2288_
	);
	LUT4 #(
		.INIT('h3fff)
	) name1836 (
		\InstQueueWr_Addr_reg[0]/NET0131 ,
		\InstQueueWr_Addr_reg[1]/NET0131 ,
		\InstQueueWr_Addr_reg[2]/NET0131 ,
		\InstQueueWr_Addr_reg[3]/NET0131 ,
		_w2289_
	);
	LUT4 #(
		.INIT('h5553)
	) name1837 (
		\Datai[4]_pad ,
		\InstQueue_reg[15][4]/NET0131 ,
		_w2207_,
		_w2203_,
		_w2290_
	);
	LUT2 #(
		.INIT('h2)
	) name1838 (
		\DataWidth_reg[1]/NET0131 ,
		_w2266_,
		_w2291_
	);
	LUT2 #(
		.INIT('h1)
	) name1839 (
		_w2290_,
		_w2291_,
		_w2292_
	);
	LUT4 #(
		.INIT('h0057)
	) name1840 (
		\DataWidth_reg[1]/NET0131 ,
		_w2287_,
		_w2288_,
		_w2292_,
		_w2293_
	);
	LUT4 #(
		.INIT('hc055)
	) name1841 (
		\InstQueue_reg[15][4]/NET0131 ,
		_w558_,
		_w563_,
		_w2207_,
		_w2294_
	);
	LUT2 #(
		.INIT('h2)
	) name1842 (
		\InstQueue_reg[15][4]/NET0131 ,
		_w2215_,
		_w2295_
	);
	LUT3 #(
		.INIT('h0d)
	) name1843 (
		_w706_,
		_w2290_,
		_w2295_,
		_w2296_
	);
	LUT3 #(
		.INIT('hd0)
	) name1844 (
		_w722_,
		_w2294_,
		_w2296_,
		_w2297_
	);
	LUT3 #(
		.INIT('h2f)
	) name1845 (
		_w700_,
		_w2293_,
		_w2297_,
		_w2298_
	);
	LUT3 #(
		.INIT('h60)
	) name1846 (
		\Datai[28]_pad ,
		_w2197_,
		_w2203_,
		_w2299_
	);
	LUT2 #(
		.INIT('h8)
	) name1847 (
		_w2207_,
		_w2201_,
		_w2300_
	);
	LUT4 #(
		.INIT('h0002)
	) name1848 (
		\InstQueueWr_Addr_reg[0]/NET0131 ,
		\InstQueueWr_Addr_reg[1]/NET0131 ,
		\InstQueueWr_Addr_reg[2]/NET0131 ,
		\InstQueueWr_Addr_reg[3]/NET0131 ,
		_w2301_
	);
	LUT4 #(
		.INIT('hfffc)
	) name1849 (
		\InstQueueWr_Addr_reg[0]/NET0131 ,
		\InstQueueWr_Addr_reg[1]/NET0131 ,
		\InstQueueWr_Addr_reg[2]/NET0131 ,
		\InstQueueWr_Addr_reg[3]/NET0131 ,
		_w2302_
	);
	LUT4 #(
		.INIT('h5553)
	) name1850 (
		\Datai[4]_pad ,
		\InstQueue_reg[1][4]/NET0131 ,
		_w2205_,
		_w2301_,
		_w2303_
	);
	LUT2 #(
		.INIT('h2)
	) name1851 (
		\DataWidth_reg[1]/NET0131 ,
		_w2289_,
		_w2304_
	);
	LUT2 #(
		.INIT('h1)
	) name1852 (
		_w2303_,
		_w2304_,
		_w2305_
	);
	LUT4 #(
		.INIT('h0057)
	) name1853 (
		\DataWidth_reg[1]/NET0131 ,
		_w2299_,
		_w2300_,
		_w2305_,
		_w2306_
	);
	LUT4 #(
		.INIT('hc055)
	) name1854 (
		\InstQueue_reg[1][4]/NET0131 ,
		_w558_,
		_w563_,
		_w2301_,
		_w2307_
	);
	LUT2 #(
		.INIT('h2)
	) name1855 (
		\InstQueue_reg[1][4]/NET0131 ,
		_w2215_,
		_w2308_
	);
	LUT3 #(
		.INIT('h0d)
	) name1856 (
		_w706_,
		_w2303_,
		_w2308_,
		_w2309_
	);
	LUT3 #(
		.INIT('hd0)
	) name1857 (
		_w722_,
		_w2307_,
		_w2309_,
		_w2310_
	);
	LUT3 #(
		.INIT('h2f)
	) name1858 (
		_w700_,
		_w2306_,
		_w2310_,
		_w2311_
	);
	LUT2 #(
		.INIT('h8)
	) name1859 (
		_w2205_,
		_w2201_,
		_w2312_
	);
	LUT3 #(
		.INIT('h48)
	) name1860 (
		\Datai[28]_pad ,
		_w2207_,
		_w2197_,
		_w2313_
	);
	LUT4 #(
		.INIT('h0004)
	) name1861 (
		\InstQueueWr_Addr_reg[0]/NET0131 ,
		\InstQueueWr_Addr_reg[1]/NET0131 ,
		\InstQueueWr_Addr_reg[2]/NET0131 ,
		\InstQueueWr_Addr_reg[3]/NET0131 ,
		_w2314_
	);
	LUT4 #(
		.INIT('hfff9)
	) name1862 (
		\InstQueueWr_Addr_reg[0]/NET0131 ,
		\InstQueueWr_Addr_reg[1]/NET0131 ,
		\InstQueueWr_Addr_reg[2]/NET0131 ,
		\InstQueueWr_Addr_reg[3]/NET0131 ,
		_w2315_
	);
	LUT4 #(
		.INIT('h5553)
	) name1863 (
		\Datai[4]_pad ,
		\InstQueue_reg[2][4]/NET0131 ,
		_w2301_,
		_w2314_,
		_w2316_
	);
	LUT2 #(
		.INIT('h2)
	) name1864 (
		\DataWidth_reg[1]/NET0131 ,
		_w2208_,
		_w2317_
	);
	LUT2 #(
		.INIT('h1)
	) name1865 (
		_w2316_,
		_w2317_,
		_w2318_
	);
	LUT4 #(
		.INIT('h0057)
	) name1866 (
		\DataWidth_reg[1]/NET0131 ,
		_w2312_,
		_w2313_,
		_w2318_,
		_w2319_
	);
	LUT4 #(
		.INIT('hc055)
	) name1867 (
		\InstQueue_reg[2][4]/NET0131 ,
		_w558_,
		_w563_,
		_w2314_,
		_w2320_
	);
	LUT2 #(
		.INIT('h2)
	) name1868 (
		\InstQueue_reg[2][4]/NET0131 ,
		_w2215_,
		_w2321_
	);
	LUT3 #(
		.INIT('h0d)
	) name1869 (
		_w706_,
		_w2316_,
		_w2321_,
		_w2322_
	);
	LUT3 #(
		.INIT('hd0)
	) name1870 (
		_w722_,
		_w2320_,
		_w2322_,
		_w2323_
	);
	LUT3 #(
		.INIT('h2f)
	) name1871 (
		_w700_,
		_w2319_,
		_w2323_,
		_w2324_
	);
	LUT3 #(
		.INIT('h48)
	) name1872 (
		\Datai[28]_pad ,
		_w2205_,
		_w2197_,
		_w2325_
	);
	LUT2 #(
		.INIT('h8)
	) name1873 (
		_w2201_,
		_w2301_,
		_w2326_
	);
	LUT4 #(
		.INIT('h0008)
	) name1874 (
		\InstQueueWr_Addr_reg[0]/NET0131 ,
		\InstQueueWr_Addr_reg[1]/NET0131 ,
		\InstQueueWr_Addr_reg[2]/NET0131 ,
		\InstQueueWr_Addr_reg[3]/NET0131 ,
		_w2327_
	);
	LUT4 #(
		.INIT('hfff3)
	) name1875 (
		\InstQueueWr_Addr_reg[0]/NET0131 ,
		\InstQueueWr_Addr_reg[1]/NET0131 ,
		\InstQueueWr_Addr_reg[2]/NET0131 ,
		\InstQueueWr_Addr_reg[3]/NET0131 ,
		_w2328_
	);
	LUT4 #(
		.INIT('h5553)
	) name1876 (
		\Datai[4]_pad ,
		\InstQueue_reg[3][4]/NET0131 ,
		_w2314_,
		_w2327_,
		_w2329_
	);
	LUT2 #(
		.INIT('h2)
	) name1877 (
		\DataWidth_reg[1]/NET0131 ,
		_w2302_,
		_w2330_
	);
	LUT2 #(
		.INIT('h1)
	) name1878 (
		_w2329_,
		_w2330_,
		_w2331_
	);
	LUT4 #(
		.INIT('h0057)
	) name1879 (
		\DataWidth_reg[1]/NET0131 ,
		_w2325_,
		_w2326_,
		_w2331_,
		_w2332_
	);
	LUT4 #(
		.INIT('hc055)
	) name1880 (
		\InstQueue_reg[3][4]/NET0131 ,
		_w558_,
		_w563_,
		_w2327_,
		_w2333_
	);
	LUT2 #(
		.INIT('h2)
	) name1881 (
		\InstQueue_reg[3][4]/NET0131 ,
		_w2215_,
		_w2334_
	);
	LUT3 #(
		.INIT('h0d)
	) name1882 (
		_w706_,
		_w2329_,
		_w2334_,
		_w2335_
	);
	LUT3 #(
		.INIT('hd0)
	) name1883 (
		_w722_,
		_w2333_,
		_w2335_,
		_w2336_
	);
	LUT3 #(
		.INIT('h2f)
	) name1884 (
		_w700_,
		_w2332_,
		_w2336_,
		_w2337_
	);
	LUT3 #(
		.INIT('h60)
	) name1885 (
		\Datai[28]_pad ,
		_w2197_,
		_w2301_,
		_w2338_
	);
	LUT2 #(
		.INIT('h8)
	) name1886 (
		_w2201_,
		_w2314_,
		_w2339_
	);
	LUT4 #(
		.INIT('h0010)
	) name1887 (
		\InstQueueWr_Addr_reg[0]/NET0131 ,
		\InstQueueWr_Addr_reg[1]/NET0131 ,
		\InstQueueWr_Addr_reg[2]/NET0131 ,
		\InstQueueWr_Addr_reg[3]/NET0131 ,
		_w2340_
	);
	LUT4 #(
		.INIT('hffe7)
	) name1888 (
		\InstQueueWr_Addr_reg[0]/NET0131 ,
		\InstQueueWr_Addr_reg[1]/NET0131 ,
		\InstQueueWr_Addr_reg[2]/NET0131 ,
		\InstQueueWr_Addr_reg[3]/NET0131 ,
		_w2341_
	);
	LUT4 #(
		.INIT('h5553)
	) name1889 (
		\Datai[4]_pad ,
		\InstQueue_reg[4][4]/NET0131 ,
		_w2327_,
		_w2340_,
		_w2342_
	);
	LUT2 #(
		.INIT('h2)
	) name1890 (
		\DataWidth_reg[1]/NET0131 ,
		_w2315_,
		_w2343_
	);
	LUT2 #(
		.INIT('h1)
	) name1891 (
		_w2342_,
		_w2343_,
		_w2344_
	);
	LUT4 #(
		.INIT('h0057)
	) name1892 (
		\DataWidth_reg[1]/NET0131 ,
		_w2338_,
		_w2339_,
		_w2344_,
		_w2345_
	);
	LUT4 #(
		.INIT('hc055)
	) name1893 (
		\InstQueue_reg[4][4]/NET0131 ,
		_w558_,
		_w563_,
		_w2340_,
		_w2346_
	);
	LUT2 #(
		.INIT('h2)
	) name1894 (
		\InstQueue_reg[4][4]/NET0131 ,
		_w2215_,
		_w2347_
	);
	LUT3 #(
		.INIT('h0d)
	) name1895 (
		_w706_,
		_w2342_,
		_w2347_,
		_w2348_
	);
	LUT3 #(
		.INIT('hd0)
	) name1896 (
		_w722_,
		_w2346_,
		_w2348_,
		_w2349_
	);
	LUT3 #(
		.INIT('h2f)
	) name1897 (
		_w700_,
		_w2345_,
		_w2349_,
		_w2350_
	);
	LUT3 #(
		.INIT('h60)
	) name1898 (
		\Datai[28]_pad ,
		_w2197_,
		_w2314_,
		_w2351_
	);
	LUT2 #(
		.INIT('h8)
	) name1899 (
		_w2201_,
		_w2327_,
		_w2352_
	);
	LUT4 #(
		.INIT('h0020)
	) name1900 (
		\InstQueueWr_Addr_reg[0]/NET0131 ,
		\InstQueueWr_Addr_reg[1]/NET0131 ,
		\InstQueueWr_Addr_reg[2]/NET0131 ,
		\InstQueueWr_Addr_reg[3]/NET0131 ,
		_w2353_
	);
	LUT4 #(
		.INIT('hffcf)
	) name1901 (
		\InstQueueWr_Addr_reg[0]/NET0131 ,
		\InstQueueWr_Addr_reg[1]/NET0131 ,
		\InstQueueWr_Addr_reg[2]/NET0131 ,
		\InstQueueWr_Addr_reg[3]/NET0131 ,
		_w2354_
	);
	LUT4 #(
		.INIT('h5553)
	) name1902 (
		\Datai[4]_pad ,
		\InstQueue_reg[5][4]/NET0131 ,
		_w2340_,
		_w2353_,
		_w2355_
	);
	LUT2 #(
		.INIT('h2)
	) name1903 (
		\DataWidth_reg[1]/NET0131 ,
		_w2328_,
		_w2356_
	);
	LUT2 #(
		.INIT('h1)
	) name1904 (
		_w2355_,
		_w2356_,
		_w2357_
	);
	LUT4 #(
		.INIT('h0057)
	) name1905 (
		\DataWidth_reg[1]/NET0131 ,
		_w2351_,
		_w2352_,
		_w2357_,
		_w2358_
	);
	LUT4 #(
		.INIT('hc055)
	) name1906 (
		\InstQueue_reg[5][4]/NET0131 ,
		_w558_,
		_w563_,
		_w2353_,
		_w2359_
	);
	LUT2 #(
		.INIT('h2)
	) name1907 (
		\InstQueue_reg[5][4]/NET0131 ,
		_w2215_,
		_w2360_
	);
	LUT3 #(
		.INIT('h0d)
	) name1908 (
		_w706_,
		_w2355_,
		_w2360_,
		_w2361_
	);
	LUT3 #(
		.INIT('hd0)
	) name1909 (
		_w722_,
		_w2359_,
		_w2361_,
		_w2362_
	);
	LUT3 #(
		.INIT('h2f)
	) name1910 (
		_w700_,
		_w2358_,
		_w2362_,
		_w2363_
	);
	LUT3 #(
		.INIT('h60)
	) name1911 (
		\Datai[28]_pad ,
		_w2197_,
		_w2327_,
		_w2364_
	);
	LUT2 #(
		.INIT('h8)
	) name1912 (
		_w2201_,
		_w2340_,
		_w2365_
	);
	LUT4 #(
		.INIT('h0040)
	) name1913 (
		\InstQueueWr_Addr_reg[0]/NET0131 ,
		\InstQueueWr_Addr_reg[1]/NET0131 ,
		\InstQueueWr_Addr_reg[2]/NET0131 ,
		\InstQueueWr_Addr_reg[3]/NET0131 ,
		_w2366_
	);
	LUT4 #(
		.INIT('hff9f)
	) name1914 (
		\InstQueueWr_Addr_reg[0]/NET0131 ,
		\InstQueueWr_Addr_reg[1]/NET0131 ,
		\InstQueueWr_Addr_reg[2]/NET0131 ,
		\InstQueueWr_Addr_reg[3]/NET0131 ,
		_w2367_
	);
	LUT4 #(
		.INIT('h5553)
	) name1915 (
		\Datai[4]_pad ,
		\InstQueue_reg[6][4]/NET0131 ,
		_w2353_,
		_w2366_,
		_w2368_
	);
	LUT2 #(
		.INIT('h2)
	) name1916 (
		\DataWidth_reg[1]/NET0131 ,
		_w2341_,
		_w2369_
	);
	LUT2 #(
		.INIT('h1)
	) name1917 (
		_w2368_,
		_w2369_,
		_w2370_
	);
	LUT4 #(
		.INIT('h0057)
	) name1918 (
		\DataWidth_reg[1]/NET0131 ,
		_w2364_,
		_w2365_,
		_w2370_,
		_w2371_
	);
	LUT4 #(
		.INIT('hc055)
	) name1919 (
		\InstQueue_reg[6][4]/NET0131 ,
		_w558_,
		_w563_,
		_w2366_,
		_w2372_
	);
	LUT2 #(
		.INIT('h2)
	) name1920 (
		\InstQueue_reg[6][4]/NET0131 ,
		_w2215_,
		_w2373_
	);
	LUT3 #(
		.INIT('h0d)
	) name1921 (
		_w706_,
		_w2368_,
		_w2373_,
		_w2374_
	);
	LUT3 #(
		.INIT('hd0)
	) name1922 (
		_w722_,
		_w2372_,
		_w2374_,
		_w2375_
	);
	LUT3 #(
		.INIT('h2f)
	) name1923 (
		_w700_,
		_w2371_,
		_w2375_,
		_w2376_
	);
	LUT3 #(
		.INIT('h60)
	) name1924 (
		\Datai[28]_pad ,
		_w2197_,
		_w2340_,
		_w2377_
	);
	LUT2 #(
		.INIT('h8)
	) name1925 (
		_w2201_,
		_w2353_,
		_w2378_
	);
	LUT4 #(
		.INIT('hff3f)
	) name1926 (
		\InstQueueWr_Addr_reg[0]/NET0131 ,
		\InstQueueWr_Addr_reg[1]/NET0131 ,
		\InstQueueWr_Addr_reg[2]/NET0131 ,
		\InstQueueWr_Addr_reg[3]/NET0131 ,
		_w2379_
	);
	LUT4 #(
		.INIT('h5553)
	) name1927 (
		\Datai[4]_pad ,
		\InstQueue_reg[7][4]/NET0131 ,
		_w2220_,
		_w2366_,
		_w2380_
	);
	LUT2 #(
		.INIT('h2)
	) name1928 (
		\DataWidth_reg[1]/NET0131 ,
		_w2354_,
		_w2381_
	);
	LUT2 #(
		.INIT('h1)
	) name1929 (
		_w2380_,
		_w2381_,
		_w2382_
	);
	LUT4 #(
		.INIT('h0057)
	) name1930 (
		\DataWidth_reg[1]/NET0131 ,
		_w2377_,
		_w2378_,
		_w2382_,
		_w2383_
	);
	LUT4 #(
		.INIT('hc055)
	) name1931 (
		\InstQueue_reg[7][4]/NET0131 ,
		_w558_,
		_w563_,
		_w2220_,
		_w2384_
	);
	LUT2 #(
		.INIT('h2)
	) name1932 (
		\InstQueue_reg[7][4]/NET0131 ,
		_w2215_,
		_w2385_
	);
	LUT3 #(
		.INIT('h0d)
	) name1933 (
		_w706_,
		_w2380_,
		_w2385_,
		_w2386_
	);
	LUT3 #(
		.INIT('hd0)
	) name1934 (
		_w722_,
		_w2384_,
		_w2386_,
		_w2387_
	);
	LUT3 #(
		.INIT('h2f)
	) name1935 (
		_w700_,
		_w2383_,
		_w2387_,
		_w2388_
	);
	LUT3 #(
		.INIT('h60)
	) name1936 (
		\Datai[28]_pad ,
		_w2197_,
		_w2353_,
		_w2389_
	);
	LUT2 #(
		.INIT('h8)
	) name1937 (
		_w2201_,
		_w2366_,
		_w2390_
	);
	LUT4 #(
		.INIT('h5553)
	) name1938 (
		\Datai[4]_pad ,
		\InstQueue_reg[8][4]/NET0131 ,
		_w2220_,
		_w2222_,
		_w2391_
	);
	LUT2 #(
		.INIT('h2)
	) name1939 (
		\DataWidth_reg[1]/NET0131 ,
		_w2367_,
		_w2392_
	);
	LUT2 #(
		.INIT('h1)
	) name1940 (
		_w2391_,
		_w2392_,
		_w2393_
	);
	LUT4 #(
		.INIT('h0057)
	) name1941 (
		\DataWidth_reg[1]/NET0131 ,
		_w2389_,
		_w2390_,
		_w2393_,
		_w2394_
	);
	LUT4 #(
		.INIT('hc055)
	) name1942 (
		\InstQueue_reg[8][4]/NET0131 ,
		_w558_,
		_w563_,
		_w2222_,
		_w2395_
	);
	LUT2 #(
		.INIT('h2)
	) name1943 (
		\InstQueue_reg[8][4]/NET0131 ,
		_w2215_,
		_w2396_
	);
	LUT3 #(
		.INIT('h0d)
	) name1944 (
		_w706_,
		_w2391_,
		_w2396_,
		_w2397_
	);
	LUT3 #(
		.INIT('hd0)
	) name1945 (
		_w722_,
		_w2395_,
		_w2397_,
		_w2398_
	);
	LUT3 #(
		.INIT('h2f)
	) name1946 (
		_w700_,
		_w2394_,
		_w2398_,
		_w2399_
	);
	LUT3 #(
		.INIT('h60)
	) name1947 (
		\Datai[28]_pad ,
		_w2197_,
		_w2366_,
		_w2400_
	);
	LUT2 #(
		.INIT('h8)
	) name1948 (
		_w2201_,
		_w2220_,
		_w2401_
	);
	LUT4 #(
		.INIT('h5553)
	) name1949 (
		\Datai[4]_pad ,
		\InstQueue_reg[9][4]/NET0131 ,
		_w2225_,
		_w2222_,
		_w2402_
	);
	LUT2 #(
		.INIT('h2)
	) name1950 (
		\DataWidth_reg[1]/NET0131 ,
		_w2379_,
		_w2403_
	);
	LUT2 #(
		.INIT('h1)
	) name1951 (
		_w2402_,
		_w2403_,
		_w2404_
	);
	LUT4 #(
		.INIT('h0057)
	) name1952 (
		\DataWidth_reg[1]/NET0131 ,
		_w2400_,
		_w2401_,
		_w2404_,
		_w2405_
	);
	LUT4 #(
		.INIT('hc055)
	) name1953 (
		\InstQueue_reg[9][4]/NET0131 ,
		_w558_,
		_w563_,
		_w2225_,
		_w2406_
	);
	LUT2 #(
		.INIT('h2)
	) name1954 (
		\InstQueue_reg[9][4]/NET0131 ,
		_w2215_,
		_w2407_
	);
	LUT3 #(
		.INIT('h0d)
	) name1955 (
		_w706_,
		_w2402_,
		_w2407_,
		_w2408_
	);
	LUT3 #(
		.INIT('hd0)
	) name1956 (
		_w722_,
		_w2406_,
		_w2408_,
		_w2409_
	);
	LUT3 #(
		.INIT('h2f)
	) name1957 (
		_w700_,
		_w2405_,
		_w2409_,
		_w2410_
	);
	LUT4 #(
		.INIT('h000d)
	) name1958 (
		\PhyAddrPointer_reg[2]/NET0131 ,
		_w1984_,
		_w2006_,
		_w2010_,
		_w2411_
	);
	LUT2 #(
		.INIT('h2)
	) name1959 (
		\PhyAddrPointer_reg[2]/NET0131 ,
		_w1283_,
		_w2412_
	);
	LUT2 #(
		.INIT('h6)
	) name1960 (
		\PhyAddrPointer_reg[1]/NET0131 ,
		\PhyAddrPointer_reg[2]/NET0131 ,
		_w2413_
	);
	LUT4 #(
		.INIT('hf400)
	) name1961 (
		\DataWidth_reg[1]/NET0131 ,
		_w700_,
		_w706_,
		_w2413_,
		_w2414_
	);
	LUT3 #(
		.INIT('h20)
	) name1962 (
		\DataWidth_reg[1]/NET0131 ,
		\PhyAddrPointer_reg[2]/NET0131 ,
		_w700_,
		_w2415_
	);
	LUT4 #(
		.INIT('h0001)
	) name1963 (
		_w2014_,
		_w2414_,
		_w2412_,
		_w2415_,
		_w2416_
	);
	LUT3 #(
		.INIT('h2f)
	) name1964 (
		_w695_,
		_w2411_,
		_w2416_,
		_w2417_
	);
	LUT4 #(
		.INIT('h8000)
	) name1965 (
		\EAX_reg[18]/NET0131 ,
		\EAX_reg[19]/NET0131 ,
		\EAX_reg[20]/NET0131 ,
		_w2047_,
		_w2418_
	);
	LUT4 #(
		.INIT('h78f0)
	) name1966 (
		\EAX_reg[18]/NET0131 ,
		\EAX_reg[19]/NET0131 ,
		\EAX_reg[20]/NET0131 ,
		_w2047_,
		_w2419_
	);
	LUT3 #(
		.INIT('h80)
	) name1967 (
		_w570_,
		_w611_,
		_w2419_,
		_w2420_
	);
	LUT4 #(
		.INIT('h0800)
	) name1968 (
		_w570_,
		_w611_,
		_w617_,
		_w2419_,
		_w2421_
	);
	LUT4 #(
		.INIT('hf400)
	) name1969 (
		_w514_,
		_w569_,
		_w570_,
		_w659_,
		_w2422_
	);
	LUT4 #(
		.INIT('hc0c8)
	) name1970 (
		\Datao[20]_pad ,
		_w695_,
		_w2421_,
		_w2422_,
		_w2423_
	);
	LUT4 #(
		.INIT('h3f15)
	) name1971 (
		\Datao[20]_pad ,
		\uWord_reg[4]/NET0131 ,
		_w696_,
		_w2159_,
		_w2424_
	);
	LUT2 #(
		.INIT('hb)
	) name1972 (
		_w2423_,
		_w2424_,
		_w2425_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name1973 (
		\uWord_reg[4]/NET0131 ,
		_w695_,
		_w1825_,
		_w2058_,
		_w2426_
	);
	LUT2 #(
		.INIT('h8)
	) name1974 (
		\Datai[4]_pad ,
		_w566_,
		_w2427_
	);
	LUT3 #(
		.INIT('h80)
	) name1975 (
		\Datai[4]_pad ,
		_w566_,
		_w612_,
		_w2428_
	);
	LUT3 #(
		.INIT('ha8)
	) name1976 (
		_w695_,
		_w2420_,
		_w2428_,
		_w2429_
	);
	LUT2 #(
		.INIT('he)
	) name1977 (
		_w2426_,
		_w2429_,
		_w2430_
	);
	LUT2 #(
		.INIT('h2)
	) name1978 (
		\EAX_reg[25]/NET0131 ,
		_w1825_,
		_w2431_
	);
	LUT4 #(
		.INIT('h8000)
	) name1979 (
		\EAX_reg[19]/NET0131 ,
		\EAX_reg[23]/NET0131 ,
		_w1837_,
		_w1839_,
		_w2432_
	);
	LUT3 #(
		.INIT('h13)
	) name1980 (
		\EAX_reg[24]/NET0131 ,
		\EAX_reg[25]/NET0131 ,
		_w2432_,
		_w2433_
	);
	LUT2 #(
		.INIT('h2)
	) name1981 (
		_w1848_,
		_w2029_,
		_w2434_
	);
	LUT4 #(
		.INIT('h08a2)
	) name1982 (
		_w605_,
		_w1873_,
		_w1884_,
		_w1895_,
		_w2435_
	);
	LUT3 #(
		.INIT('h80)
	) name1983 (
		_w576_,
		_w579_,
		_w2435_,
		_w2436_
	);
	LUT3 #(
		.INIT('h80)
	) name1984 (
		\Datai[25]_pad ,
		_w514_,
		_w569_,
		_w2437_
	);
	LUT2 #(
		.INIT('h8)
	) name1985 (
		\Datai[9]_pad ,
		_w566_,
		_w2438_
	);
	LUT4 #(
		.INIT('h1113)
	) name1986 (
		_w612_,
		_w2436_,
		_w2437_,
		_w2438_,
		_w2439_
	);
	LUT4 #(
		.INIT('h7500)
	) name1987 (
		\EAX_reg[25]/NET0131 ,
		_w635_,
		_w1852_,
		_w2439_,
		_w2440_
	);
	LUT4 #(
		.INIT('h20aa)
	) name1988 (
		_w695_,
		_w2433_,
		_w2434_,
		_w2440_,
		_w2441_
	);
	LUT2 #(
		.INIT('he)
	) name1989 (
		_w2431_,
		_w2441_,
		_w2442_
	);
	LUT4 #(
		.INIT('h8000)
	) name1990 (
		\Datai[28]_pad ,
		\Datai[29]_pad ,
		\Datai[30]_pad ,
		_w2197_,
		_w2443_
	);
	LUT3 #(
		.INIT('h08)
	) name1991 (
		\Datai[31]_pad ,
		_w2187_,
		_w2443_,
		_w2444_
	);
	LUT4 #(
		.INIT('h78f0)
	) name1992 (
		\Datai[21]_pad ,
		\Datai[22]_pad ,
		\Datai[23]_pad ,
		_w2200_,
		_w2445_
	);
	LUT2 #(
		.INIT('h8)
	) name1993 (
		_w2203_,
		_w2445_,
		_w2446_
	);
	LUT4 #(
		.INIT('h5553)
	) name1994 (
		\Datai[7]_pad ,
		\InstQueue_reg[0][7]/NET0131 ,
		_w2205_,
		_w2207_,
		_w2447_
	);
	LUT2 #(
		.INIT('h1)
	) name1995 (
		_w2211_,
		_w2447_,
		_w2448_
	);
	LUT4 #(
		.INIT('h0057)
	) name1996 (
		\DataWidth_reg[1]/NET0131 ,
		_w2444_,
		_w2446_,
		_w2448_,
		_w2449_
	);
	LUT4 #(
		.INIT('hc055)
	) name1997 (
		\InstQueue_reg[0][7]/NET0131 ,
		_w466_,
		_w479_,
		_w2205_,
		_w2450_
	);
	LUT2 #(
		.INIT('h2)
	) name1998 (
		\InstQueue_reg[0][7]/NET0131 ,
		_w2215_,
		_w2451_
	);
	LUT3 #(
		.INIT('h0d)
	) name1999 (
		_w706_,
		_w2447_,
		_w2451_,
		_w2452_
	);
	LUT3 #(
		.INIT('hd0)
	) name2000 (
		_w722_,
		_w2450_,
		_w2452_,
		_w2453_
	);
	LUT3 #(
		.INIT('h2f)
	) name2001 (
		_w700_,
		_w2449_,
		_w2453_,
		_w2454_
	);
	LUT3 #(
		.INIT('h08)
	) name2002 (
		\Datai[31]_pad ,
		_w2220_,
		_w2443_,
		_w2455_
	);
	LUT2 #(
		.INIT('h8)
	) name2003 (
		_w2222_,
		_w2445_,
		_w2456_
	);
	LUT4 #(
		.INIT('h5553)
	) name2004 (
		\Datai[7]_pad ,
		\InstQueue_reg[10][7]/NET0131 ,
		_w2224_,
		_w2225_,
		_w2457_
	);
	LUT2 #(
		.INIT('h1)
	) name2005 (
		_w2229_,
		_w2457_,
		_w2458_
	);
	LUT4 #(
		.INIT('h0057)
	) name2006 (
		\DataWidth_reg[1]/NET0131 ,
		_w2455_,
		_w2456_,
		_w2458_,
		_w2459_
	);
	LUT4 #(
		.INIT('hc055)
	) name2007 (
		\InstQueue_reg[10][7]/NET0131 ,
		_w466_,
		_w479_,
		_w2224_,
		_w2460_
	);
	LUT2 #(
		.INIT('h2)
	) name2008 (
		\InstQueue_reg[10][7]/NET0131 ,
		_w2215_,
		_w2461_
	);
	LUT3 #(
		.INIT('h0d)
	) name2009 (
		_w706_,
		_w2457_,
		_w2461_,
		_w2462_
	);
	LUT3 #(
		.INIT('hd0)
	) name2010 (
		_w722_,
		_w2460_,
		_w2462_,
		_w2463_
	);
	LUT3 #(
		.INIT('h2f)
	) name2011 (
		_w700_,
		_w2459_,
		_w2463_,
		_w2464_
	);
	LUT3 #(
		.INIT('h08)
	) name2012 (
		\Datai[31]_pad ,
		_w2222_,
		_w2443_,
		_w2465_
	);
	LUT2 #(
		.INIT('h8)
	) name2013 (
		_w2225_,
		_w2445_,
		_w2466_
	);
	LUT4 #(
		.INIT('h5553)
	) name2014 (
		\Datai[7]_pad ,
		\InstQueue_reg[11][7]/NET0131 ,
		_w2224_,
		_w2239_,
		_w2467_
	);
	LUT2 #(
		.INIT('h1)
	) name2015 (
		_w2243_,
		_w2467_,
		_w2468_
	);
	LUT4 #(
		.INIT('h0057)
	) name2016 (
		\DataWidth_reg[1]/NET0131 ,
		_w2465_,
		_w2466_,
		_w2468_,
		_w2469_
	);
	LUT4 #(
		.INIT('hc055)
	) name2017 (
		\InstQueue_reg[11][7]/NET0131 ,
		_w466_,
		_w479_,
		_w2239_,
		_w2470_
	);
	LUT2 #(
		.INIT('h2)
	) name2018 (
		\InstQueue_reg[11][7]/NET0131 ,
		_w2215_,
		_w2471_
	);
	LUT3 #(
		.INIT('h0d)
	) name2019 (
		_w706_,
		_w2467_,
		_w2471_,
		_w2472_
	);
	LUT3 #(
		.INIT('hd0)
	) name2020 (
		_w722_,
		_w2470_,
		_w2472_,
		_w2473_
	);
	LUT3 #(
		.INIT('h2f)
	) name2021 (
		_w700_,
		_w2469_,
		_w2473_,
		_w2474_
	);
	LUT3 #(
		.INIT('h08)
	) name2022 (
		\Datai[31]_pad ,
		_w2225_,
		_w2443_,
		_w2475_
	);
	LUT2 #(
		.INIT('h8)
	) name2023 (
		_w2224_,
		_w2445_,
		_w2476_
	);
	LUT4 #(
		.INIT('h5553)
	) name2024 (
		\Datai[7]_pad ,
		\InstQueue_reg[12][7]/NET0131 ,
		_w2239_,
		_w2253_,
		_w2477_
	);
	LUT2 #(
		.INIT('h1)
	) name2025 (
		_w2256_,
		_w2477_,
		_w2478_
	);
	LUT4 #(
		.INIT('h0057)
	) name2026 (
		\DataWidth_reg[1]/NET0131 ,
		_w2475_,
		_w2476_,
		_w2478_,
		_w2479_
	);
	LUT4 #(
		.INIT('hc055)
	) name2027 (
		\InstQueue_reg[12][7]/NET0131 ,
		_w466_,
		_w479_,
		_w2253_,
		_w2480_
	);
	LUT2 #(
		.INIT('h2)
	) name2028 (
		\InstQueue_reg[12][7]/NET0131 ,
		_w2215_,
		_w2481_
	);
	LUT3 #(
		.INIT('h0d)
	) name2029 (
		_w706_,
		_w2477_,
		_w2481_,
		_w2482_
	);
	LUT3 #(
		.INIT('hd0)
	) name2030 (
		_w722_,
		_w2480_,
		_w2482_,
		_w2483_
	);
	LUT3 #(
		.INIT('h2f)
	) name2031 (
		_w700_,
		_w2479_,
		_w2483_,
		_w2484_
	);
	LUT3 #(
		.INIT('h08)
	) name2032 (
		\Datai[31]_pad ,
		_w2224_,
		_w2443_,
		_w2485_
	);
	LUT2 #(
		.INIT('h8)
	) name2033 (
		_w2239_,
		_w2445_,
		_w2486_
	);
	LUT4 #(
		.INIT('h5553)
	) name2034 (
		\Datai[7]_pad ,
		\InstQueue_reg[13][7]/NET0131 ,
		_w2187_,
		_w2253_,
		_w2487_
	);
	LUT2 #(
		.INIT('h1)
	) name2035 (
		_w2268_,
		_w2487_,
		_w2488_
	);
	LUT4 #(
		.INIT('h0057)
	) name2036 (
		\DataWidth_reg[1]/NET0131 ,
		_w2485_,
		_w2486_,
		_w2488_,
		_w2489_
	);
	LUT4 #(
		.INIT('hc055)
	) name2037 (
		\InstQueue_reg[13][7]/NET0131 ,
		_w466_,
		_w479_,
		_w2187_,
		_w2490_
	);
	LUT2 #(
		.INIT('h2)
	) name2038 (
		\InstQueue_reg[13][7]/NET0131 ,
		_w2215_,
		_w2491_
	);
	LUT3 #(
		.INIT('h0d)
	) name2039 (
		_w706_,
		_w2487_,
		_w2491_,
		_w2492_
	);
	LUT3 #(
		.INIT('hd0)
	) name2040 (
		_w722_,
		_w2490_,
		_w2492_,
		_w2493_
	);
	LUT3 #(
		.INIT('h2f)
	) name2041 (
		_w700_,
		_w2489_,
		_w2493_,
		_w2494_
	);
	LUT3 #(
		.INIT('h08)
	) name2042 (
		\Datai[31]_pad ,
		_w2239_,
		_w2443_,
		_w2495_
	);
	LUT2 #(
		.INIT('h8)
	) name2043 (
		_w2253_,
		_w2445_,
		_w2496_
	);
	LUT4 #(
		.INIT('h5553)
	) name2044 (
		\Datai[7]_pad ,
		\InstQueue_reg[14][7]/NET0131 ,
		_w2187_,
		_w2203_,
		_w2497_
	);
	LUT2 #(
		.INIT('h1)
	) name2045 (
		_w2279_,
		_w2497_,
		_w2498_
	);
	LUT4 #(
		.INIT('h0057)
	) name2046 (
		\DataWidth_reg[1]/NET0131 ,
		_w2495_,
		_w2496_,
		_w2498_,
		_w2499_
	);
	LUT4 #(
		.INIT('hc055)
	) name2047 (
		\InstQueue_reg[14][7]/NET0131 ,
		_w466_,
		_w479_,
		_w2203_,
		_w2500_
	);
	LUT2 #(
		.INIT('h2)
	) name2048 (
		\InstQueue_reg[14][7]/NET0131 ,
		_w2215_,
		_w2501_
	);
	LUT3 #(
		.INIT('h0d)
	) name2049 (
		_w706_,
		_w2497_,
		_w2501_,
		_w2502_
	);
	LUT3 #(
		.INIT('hd0)
	) name2050 (
		_w722_,
		_w2500_,
		_w2502_,
		_w2503_
	);
	LUT3 #(
		.INIT('h2f)
	) name2051 (
		_w700_,
		_w2499_,
		_w2503_,
		_w2504_
	);
	LUT3 #(
		.INIT('h08)
	) name2052 (
		\Datai[31]_pad ,
		_w2253_,
		_w2443_,
		_w2505_
	);
	LUT2 #(
		.INIT('h8)
	) name2053 (
		_w2187_,
		_w2445_,
		_w2506_
	);
	LUT4 #(
		.INIT('h5553)
	) name2054 (
		\Datai[7]_pad ,
		\InstQueue_reg[15][7]/NET0131 ,
		_w2207_,
		_w2203_,
		_w2507_
	);
	LUT2 #(
		.INIT('h1)
	) name2055 (
		_w2291_,
		_w2507_,
		_w2508_
	);
	LUT4 #(
		.INIT('h0057)
	) name2056 (
		\DataWidth_reg[1]/NET0131 ,
		_w2505_,
		_w2506_,
		_w2508_,
		_w2509_
	);
	LUT4 #(
		.INIT('hc055)
	) name2057 (
		\InstQueue_reg[15][7]/NET0131 ,
		_w466_,
		_w479_,
		_w2207_,
		_w2510_
	);
	LUT2 #(
		.INIT('h2)
	) name2058 (
		\InstQueue_reg[15][7]/NET0131 ,
		_w2215_,
		_w2511_
	);
	LUT3 #(
		.INIT('h0d)
	) name2059 (
		_w706_,
		_w2507_,
		_w2511_,
		_w2512_
	);
	LUT3 #(
		.INIT('hd0)
	) name2060 (
		_w722_,
		_w2510_,
		_w2512_,
		_w2513_
	);
	LUT3 #(
		.INIT('h2f)
	) name2061 (
		_w700_,
		_w2509_,
		_w2513_,
		_w2514_
	);
	LUT3 #(
		.INIT('h08)
	) name2062 (
		\Datai[31]_pad ,
		_w2203_,
		_w2443_,
		_w2515_
	);
	LUT2 #(
		.INIT('h8)
	) name2063 (
		_w2207_,
		_w2445_,
		_w2516_
	);
	LUT4 #(
		.INIT('h5553)
	) name2064 (
		\Datai[7]_pad ,
		\InstQueue_reg[1][7]/NET0131 ,
		_w2205_,
		_w2301_,
		_w2517_
	);
	LUT2 #(
		.INIT('h1)
	) name2065 (
		_w2304_,
		_w2517_,
		_w2518_
	);
	LUT4 #(
		.INIT('h0057)
	) name2066 (
		\DataWidth_reg[1]/NET0131 ,
		_w2515_,
		_w2516_,
		_w2518_,
		_w2519_
	);
	LUT4 #(
		.INIT('hc055)
	) name2067 (
		\InstQueue_reg[1][7]/NET0131 ,
		_w466_,
		_w479_,
		_w2301_,
		_w2520_
	);
	LUT2 #(
		.INIT('h2)
	) name2068 (
		\InstQueue_reg[1][7]/NET0131 ,
		_w2215_,
		_w2521_
	);
	LUT3 #(
		.INIT('h0d)
	) name2069 (
		_w706_,
		_w2517_,
		_w2521_,
		_w2522_
	);
	LUT3 #(
		.INIT('hd0)
	) name2070 (
		_w722_,
		_w2520_,
		_w2522_,
		_w2523_
	);
	LUT3 #(
		.INIT('h2f)
	) name2071 (
		_w700_,
		_w2519_,
		_w2523_,
		_w2524_
	);
	LUT2 #(
		.INIT('h8)
	) name2072 (
		_w2205_,
		_w2445_,
		_w2525_
	);
	LUT3 #(
		.INIT('h08)
	) name2073 (
		\Datai[31]_pad ,
		_w2207_,
		_w2443_,
		_w2526_
	);
	LUT4 #(
		.INIT('h5553)
	) name2074 (
		\Datai[7]_pad ,
		\InstQueue_reg[2][7]/NET0131 ,
		_w2301_,
		_w2314_,
		_w2527_
	);
	LUT2 #(
		.INIT('h1)
	) name2075 (
		_w2317_,
		_w2527_,
		_w2528_
	);
	LUT4 #(
		.INIT('h0057)
	) name2076 (
		\DataWidth_reg[1]/NET0131 ,
		_w2525_,
		_w2526_,
		_w2528_,
		_w2529_
	);
	LUT4 #(
		.INIT('hc055)
	) name2077 (
		\InstQueue_reg[2][7]/NET0131 ,
		_w466_,
		_w479_,
		_w2314_,
		_w2530_
	);
	LUT2 #(
		.INIT('h2)
	) name2078 (
		\InstQueue_reg[2][7]/NET0131 ,
		_w2215_,
		_w2531_
	);
	LUT3 #(
		.INIT('h0d)
	) name2079 (
		_w706_,
		_w2527_,
		_w2531_,
		_w2532_
	);
	LUT3 #(
		.INIT('hd0)
	) name2080 (
		_w722_,
		_w2530_,
		_w2532_,
		_w2533_
	);
	LUT3 #(
		.INIT('h2f)
	) name2081 (
		_w700_,
		_w2529_,
		_w2533_,
		_w2534_
	);
	LUT3 #(
		.INIT('h08)
	) name2082 (
		\Datai[31]_pad ,
		_w2205_,
		_w2443_,
		_w2535_
	);
	LUT2 #(
		.INIT('h8)
	) name2083 (
		_w2301_,
		_w2445_,
		_w2536_
	);
	LUT4 #(
		.INIT('h5553)
	) name2084 (
		\Datai[7]_pad ,
		\InstQueue_reg[3][7]/NET0131 ,
		_w2314_,
		_w2327_,
		_w2537_
	);
	LUT2 #(
		.INIT('h1)
	) name2085 (
		_w2330_,
		_w2537_,
		_w2538_
	);
	LUT4 #(
		.INIT('h0057)
	) name2086 (
		\DataWidth_reg[1]/NET0131 ,
		_w2535_,
		_w2536_,
		_w2538_,
		_w2539_
	);
	LUT4 #(
		.INIT('hc055)
	) name2087 (
		\InstQueue_reg[3][7]/NET0131 ,
		_w466_,
		_w479_,
		_w2327_,
		_w2540_
	);
	LUT2 #(
		.INIT('h2)
	) name2088 (
		\InstQueue_reg[3][7]/NET0131 ,
		_w2215_,
		_w2541_
	);
	LUT3 #(
		.INIT('h0d)
	) name2089 (
		_w706_,
		_w2537_,
		_w2541_,
		_w2542_
	);
	LUT3 #(
		.INIT('hd0)
	) name2090 (
		_w722_,
		_w2540_,
		_w2542_,
		_w2543_
	);
	LUT3 #(
		.INIT('h2f)
	) name2091 (
		_w700_,
		_w2539_,
		_w2543_,
		_w2544_
	);
	LUT3 #(
		.INIT('h08)
	) name2092 (
		\Datai[31]_pad ,
		_w2301_,
		_w2443_,
		_w2545_
	);
	LUT2 #(
		.INIT('h8)
	) name2093 (
		_w2314_,
		_w2445_,
		_w2546_
	);
	LUT4 #(
		.INIT('h5553)
	) name2094 (
		\Datai[7]_pad ,
		\InstQueue_reg[4][7]/NET0131 ,
		_w2327_,
		_w2340_,
		_w2547_
	);
	LUT2 #(
		.INIT('h1)
	) name2095 (
		_w2343_,
		_w2547_,
		_w2548_
	);
	LUT4 #(
		.INIT('h0057)
	) name2096 (
		\DataWidth_reg[1]/NET0131 ,
		_w2545_,
		_w2546_,
		_w2548_,
		_w2549_
	);
	LUT4 #(
		.INIT('hc055)
	) name2097 (
		\InstQueue_reg[4][7]/NET0131 ,
		_w466_,
		_w479_,
		_w2340_,
		_w2550_
	);
	LUT2 #(
		.INIT('h2)
	) name2098 (
		\InstQueue_reg[4][7]/NET0131 ,
		_w2215_,
		_w2551_
	);
	LUT3 #(
		.INIT('h0d)
	) name2099 (
		_w706_,
		_w2547_,
		_w2551_,
		_w2552_
	);
	LUT3 #(
		.INIT('hd0)
	) name2100 (
		_w722_,
		_w2550_,
		_w2552_,
		_w2553_
	);
	LUT3 #(
		.INIT('h2f)
	) name2101 (
		_w700_,
		_w2549_,
		_w2553_,
		_w2554_
	);
	LUT3 #(
		.INIT('h08)
	) name2102 (
		\Datai[31]_pad ,
		_w2314_,
		_w2443_,
		_w2555_
	);
	LUT2 #(
		.INIT('h8)
	) name2103 (
		_w2327_,
		_w2445_,
		_w2556_
	);
	LUT4 #(
		.INIT('h5553)
	) name2104 (
		\Datai[7]_pad ,
		\InstQueue_reg[5][7]/NET0131 ,
		_w2340_,
		_w2353_,
		_w2557_
	);
	LUT2 #(
		.INIT('h1)
	) name2105 (
		_w2356_,
		_w2557_,
		_w2558_
	);
	LUT4 #(
		.INIT('h0057)
	) name2106 (
		\DataWidth_reg[1]/NET0131 ,
		_w2555_,
		_w2556_,
		_w2558_,
		_w2559_
	);
	LUT4 #(
		.INIT('hc055)
	) name2107 (
		\InstQueue_reg[5][7]/NET0131 ,
		_w466_,
		_w479_,
		_w2353_,
		_w2560_
	);
	LUT2 #(
		.INIT('h2)
	) name2108 (
		\InstQueue_reg[5][7]/NET0131 ,
		_w2215_,
		_w2561_
	);
	LUT3 #(
		.INIT('h0d)
	) name2109 (
		_w706_,
		_w2557_,
		_w2561_,
		_w2562_
	);
	LUT3 #(
		.INIT('hd0)
	) name2110 (
		_w722_,
		_w2560_,
		_w2562_,
		_w2563_
	);
	LUT3 #(
		.INIT('h2f)
	) name2111 (
		_w700_,
		_w2559_,
		_w2563_,
		_w2564_
	);
	LUT3 #(
		.INIT('h08)
	) name2112 (
		\Datai[31]_pad ,
		_w2327_,
		_w2443_,
		_w2565_
	);
	LUT2 #(
		.INIT('h8)
	) name2113 (
		_w2340_,
		_w2445_,
		_w2566_
	);
	LUT4 #(
		.INIT('h5553)
	) name2114 (
		\Datai[7]_pad ,
		\InstQueue_reg[6][7]/NET0131 ,
		_w2353_,
		_w2366_,
		_w2567_
	);
	LUT2 #(
		.INIT('h1)
	) name2115 (
		_w2369_,
		_w2567_,
		_w2568_
	);
	LUT4 #(
		.INIT('h0057)
	) name2116 (
		\DataWidth_reg[1]/NET0131 ,
		_w2565_,
		_w2566_,
		_w2568_,
		_w2569_
	);
	LUT4 #(
		.INIT('hc055)
	) name2117 (
		\InstQueue_reg[6][7]/NET0131 ,
		_w466_,
		_w479_,
		_w2366_,
		_w2570_
	);
	LUT2 #(
		.INIT('h2)
	) name2118 (
		\InstQueue_reg[6][7]/NET0131 ,
		_w2215_,
		_w2571_
	);
	LUT3 #(
		.INIT('h0d)
	) name2119 (
		_w706_,
		_w2567_,
		_w2571_,
		_w2572_
	);
	LUT3 #(
		.INIT('hd0)
	) name2120 (
		_w722_,
		_w2570_,
		_w2572_,
		_w2573_
	);
	LUT3 #(
		.INIT('h2f)
	) name2121 (
		_w700_,
		_w2569_,
		_w2573_,
		_w2574_
	);
	LUT3 #(
		.INIT('h08)
	) name2122 (
		\Datai[31]_pad ,
		_w2340_,
		_w2443_,
		_w2575_
	);
	LUT2 #(
		.INIT('h8)
	) name2123 (
		_w2353_,
		_w2445_,
		_w2576_
	);
	LUT4 #(
		.INIT('h5553)
	) name2124 (
		\Datai[7]_pad ,
		\InstQueue_reg[7][7]/NET0131 ,
		_w2220_,
		_w2366_,
		_w2577_
	);
	LUT2 #(
		.INIT('h1)
	) name2125 (
		_w2381_,
		_w2577_,
		_w2578_
	);
	LUT4 #(
		.INIT('h0057)
	) name2126 (
		\DataWidth_reg[1]/NET0131 ,
		_w2575_,
		_w2576_,
		_w2578_,
		_w2579_
	);
	LUT4 #(
		.INIT('hc055)
	) name2127 (
		\InstQueue_reg[7][7]/NET0131 ,
		_w466_,
		_w479_,
		_w2220_,
		_w2580_
	);
	LUT2 #(
		.INIT('h2)
	) name2128 (
		\InstQueue_reg[7][7]/NET0131 ,
		_w2215_,
		_w2581_
	);
	LUT3 #(
		.INIT('h0d)
	) name2129 (
		_w706_,
		_w2577_,
		_w2581_,
		_w2582_
	);
	LUT3 #(
		.INIT('hd0)
	) name2130 (
		_w722_,
		_w2580_,
		_w2582_,
		_w2583_
	);
	LUT3 #(
		.INIT('h2f)
	) name2131 (
		_w700_,
		_w2579_,
		_w2583_,
		_w2584_
	);
	LUT3 #(
		.INIT('h08)
	) name2132 (
		\Datai[31]_pad ,
		_w2353_,
		_w2443_,
		_w2585_
	);
	LUT2 #(
		.INIT('h8)
	) name2133 (
		_w2366_,
		_w2445_,
		_w2586_
	);
	LUT4 #(
		.INIT('h5553)
	) name2134 (
		\Datai[7]_pad ,
		\InstQueue_reg[8][7]/NET0131 ,
		_w2220_,
		_w2222_,
		_w2587_
	);
	LUT2 #(
		.INIT('h1)
	) name2135 (
		_w2392_,
		_w2587_,
		_w2588_
	);
	LUT4 #(
		.INIT('h0057)
	) name2136 (
		\DataWidth_reg[1]/NET0131 ,
		_w2585_,
		_w2586_,
		_w2588_,
		_w2589_
	);
	LUT4 #(
		.INIT('hc055)
	) name2137 (
		\InstQueue_reg[8][7]/NET0131 ,
		_w466_,
		_w479_,
		_w2222_,
		_w2590_
	);
	LUT2 #(
		.INIT('h2)
	) name2138 (
		\InstQueue_reg[8][7]/NET0131 ,
		_w2215_,
		_w2591_
	);
	LUT3 #(
		.INIT('h0d)
	) name2139 (
		_w706_,
		_w2587_,
		_w2591_,
		_w2592_
	);
	LUT3 #(
		.INIT('hd0)
	) name2140 (
		_w722_,
		_w2590_,
		_w2592_,
		_w2593_
	);
	LUT3 #(
		.INIT('h2f)
	) name2141 (
		_w700_,
		_w2589_,
		_w2593_,
		_w2594_
	);
	LUT3 #(
		.INIT('h08)
	) name2142 (
		\Datai[31]_pad ,
		_w2366_,
		_w2443_,
		_w2595_
	);
	LUT2 #(
		.INIT('h8)
	) name2143 (
		_w2220_,
		_w2445_,
		_w2596_
	);
	LUT4 #(
		.INIT('h5553)
	) name2144 (
		\Datai[7]_pad ,
		\InstQueue_reg[9][7]/NET0131 ,
		_w2225_,
		_w2222_,
		_w2597_
	);
	LUT2 #(
		.INIT('h1)
	) name2145 (
		_w2403_,
		_w2597_,
		_w2598_
	);
	LUT4 #(
		.INIT('h0057)
	) name2146 (
		\DataWidth_reg[1]/NET0131 ,
		_w2595_,
		_w2596_,
		_w2598_,
		_w2599_
	);
	LUT4 #(
		.INIT('hc055)
	) name2147 (
		\InstQueue_reg[9][7]/NET0131 ,
		_w466_,
		_w479_,
		_w2225_,
		_w2600_
	);
	LUT2 #(
		.INIT('h2)
	) name2148 (
		\InstQueue_reg[9][7]/NET0131 ,
		_w2215_,
		_w2601_
	);
	LUT3 #(
		.INIT('h0d)
	) name2149 (
		_w706_,
		_w2597_,
		_w2601_,
		_w2602_
	);
	LUT3 #(
		.INIT('hd0)
	) name2150 (
		_w722_,
		_w2600_,
		_w2602_,
		_w2603_
	);
	LUT3 #(
		.INIT('h2f)
	) name2151 (
		_w700_,
		_w2599_,
		_w2603_,
		_w2604_
	);
	LUT2 #(
		.INIT('h8)
	) name2152 (
		\rEIP_reg[22]/NET0131 ,
		\rEIP_reg[23]/NET0131 ,
		_w2605_
	);
	LUT4 #(
		.INIT('h8000)
	) name2153 (
		\rEIP_reg[1]/NET0131 ,
		\rEIP_reg[2]/NET0131 ,
		\rEIP_reg[3]/NET0131 ,
		\rEIP_reg[4]/NET0131 ,
		_w2606_
	);
	LUT4 #(
		.INIT('h8000)
	) name2154 (
		\rEIP_reg[5]/NET0131 ,
		\rEIP_reg[6]/NET0131 ,
		\rEIP_reg[7]/NET0131 ,
		_w2606_,
		_w2607_
	);
	LUT4 #(
		.INIT('h8000)
	) name2155 (
		\rEIP_reg[10]/NET0131 ,
		\rEIP_reg[8]/NET0131 ,
		\rEIP_reg[9]/NET0131 ,
		_w2607_,
		_w2608_
	);
	LUT3 #(
		.INIT('h80)
	) name2156 (
		\rEIP_reg[11]/NET0131 ,
		\rEIP_reg[12]/NET0131 ,
		_w2608_,
		_w2609_
	);
	LUT4 #(
		.INIT('h8000)
	) name2157 (
		\rEIP_reg[11]/NET0131 ,
		\rEIP_reg[12]/NET0131 ,
		\rEIP_reg[13]/NET0131 ,
		_w2608_,
		_w2610_
	);
	LUT4 #(
		.INIT('h8000)
	) name2158 (
		\rEIP_reg[14]/NET0131 ,
		\rEIP_reg[15]/NET0131 ,
		\rEIP_reg[16]/NET0131 ,
		_w2610_,
		_w2611_
	);
	LUT2 #(
		.INIT('h8)
	) name2159 (
		\rEIP_reg[17]/NET0131 ,
		\rEIP_reg[18]/NET0131 ,
		_w2612_
	);
	LUT3 #(
		.INIT('h80)
	) name2160 (
		\rEIP_reg[17]/NET0131 ,
		\rEIP_reg[18]/NET0131 ,
		\rEIP_reg[19]/NET0131 ,
		_w2613_
	);
	LUT2 #(
		.INIT('h8)
	) name2161 (
		\rEIP_reg[20]/NET0131 ,
		\rEIP_reg[21]/NET0131 ,
		_w2614_
	);
	LUT2 #(
		.INIT('h8)
	) name2162 (
		_w2613_,
		_w2614_,
		_w2615_
	);
	LUT3 #(
		.INIT('h80)
	) name2163 (
		_w2605_,
		_w2611_,
		_w2615_,
		_w2616_
	);
	LUT2 #(
		.INIT('h8)
	) name2164 (
		\rEIP_reg[24]/NET0131 ,
		\rEIP_reg[25]/NET0131 ,
		_w2617_
	);
	LUT3 #(
		.INIT('h80)
	) name2165 (
		\rEIP_reg[24]/NET0131 ,
		\rEIP_reg[25]/NET0131 ,
		\rEIP_reg[26]/NET0131 ,
		_w2618_
	);
	LUT4 #(
		.INIT('h8000)
	) name2166 (
		_w2605_,
		_w2611_,
		_w2615_,
		_w2618_,
		_w2619_
	);
	LUT2 #(
		.INIT('h8)
	) name2167 (
		\rEIP_reg[27]/NET0131 ,
		\rEIP_reg[28]/NET0131 ,
		_w2620_
	);
	LUT3 #(
		.INIT('h80)
	) name2168 (
		\rEIP_reg[27]/NET0131 ,
		\rEIP_reg[28]/NET0131 ,
		\rEIP_reg[29]/NET0131 ,
		_w2621_
	);
	LUT4 #(
		.INIT('h8000)
	) name2169 (
		\rEIP_reg[27]/NET0131 ,
		\rEIP_reg[28]/NET0131 ,
		\rEIP_reg[29]/NET0131 ,
		\rEIP_reg[30]/NET0131 ,
		_w2622_
	);
	LUT2 #(
		.INIT('h1)
	) name2170 (
		\DataWidth_reg[1]/NET0131 ,
		READY_n_pad,
		_w2623_
	);
	LUT4 #(
		.INIT('h6a00)
	) name2171 (
		\rEIP_reg[31]/NET0131 ,
		_w2619_,
		_w2622_,
		_w2623_,
		_w2624_
	);
	LUT4 #(
		.INIT('h0001)
	) name2172 (
		\EBX_reg[0]/NET0131 ,
		\EBX_reg[1]/NET0131 ,
		\EBX_reg[2]/NET0131 ,
		\EBX_reg[3]/NET0131 ,
		_w2625_
	);
	LUT4 #(
		.INIT('h0100)
	) name2173 (
		\EBX_reg[4]/NET0131 ,
		\EBX_reg[5]/NET0131 ,
		\EBX_reg[6]/NET0131 ,
		_w2625_,
		_w2626_
	);
	LUT4 #(
		.INIT('h0100)
	) name2174 (
		\EBX_reg[7]/NET0131 ,
		\EBX_reg[8]/NET0131 ,
		\EBX_reg[9]/NET0131 ,
		_w2626_,
		_w2627_
	);
	LUT3 #(
		.INIT('h01)
	) name2175 (
		\EBX_reg[10]/NET0131 ,
		\EBX_reg[11]/NET0131 ,
		\EBX_reg[12]/NET0131 ,
		_w2628_
	);
	LUT4 #(
		.INIT('h1000)
	) name2176 (
		\EBX_reg[13]/NET0131 ,
		\EBX_reg[14]/NET0131 ,
		_w2627_,
		_w2628_,
		_w2629_
	);
	LUT4 #(
		.INIT('h0100)
	) name2177 (
		\EBX_reg[15]/NET0131 ,
		\EBX_reg[16]/NET0131 ,
		\EBX_reg[17]/NET0131 ,
		_w2629_,
		_w2630_
	);
	LUT4 #(
		.INIT('h0001)
	) name2178 (
		\EBX_reg[20]/NET0131 ,
		\EBX_reg[21]/NET0131 ,
		\EBX_reg[22]/NET0131 ,
		\EBX_reg[23]/NET0131 ,
		_w2631_
	);
	LUT4 #(
		.INIT('h1000)
	) name2179 (
		\EBX_reg[18]/NET0131 ,
		\EBX_reg[19]/NET0131 ,
		_w2630_,
		_w2631_,
		_w2632_
	);
	LUT2 #(
		.INIT('h1)
	) name2180 (
		\EBX_reg[24]/NET0131 ,
		\EBX_reg[25]/NET0131 ,
		_w2633_
	);
	LUT3 #(
		.INIT('h01)
	) name2181 (
		\EBX_reg[24]/NET0131 ,
		\EBX_reg[25]/NET0131 ,
		\EBX_reg[26]/NET0131 ,
		_w2634_
	);
	LUT3 #(
		.INIT('h32)
	) name2182 (
		\DataWidth_reg[1]/NET0131 ,
		\EBX_reg[29]/NET0131 ,
		READY_n_pad,
		_w2635_
	);
	LUT4 #(
		.INIT('h0100)
	) name2183 (
		\EBX_reg[27]/NET0131 ,
		\EBX_reg[28]/NET0131 ,
		\EBX_reg[30]/NET0131 ,
		\EBX_reg[31]/NET0131 ,
		_w2636_
	);
	LUT2 #(
		.INIT('h8)
	) name2184 (
		_w2635_,
		_w2636_,
		_w2637_
	);
	LUT3 #(
		.INIT('h80)
	) name2185 (
		_w2632_,
		_w2634_,
		_w2637_,
		_w2638_
	);
	LUT3 #(
		.INIT('ha8)
	) name2186 (
		_w1100_,
		_w2624_,
		_w2638_,
		_w2639_
	);
	LUT4 #(
		.INIT('hfe00)
	) name2187 (
		_w566_,
		_w569_,
		_w570_,
		_w611_,
		_w2640_
	);
	LUT2 #(
		.INIT('h2)
	) name2188 (
		\rEIP_reg[31]/NET0131 ,
		_w2640_,
		_w2641_
	);
	LUT2 #(
		.INIT('h4)
	) name2189 (
		\DataWidth_reg[1]/NET0131 ,
		_w633_,
		_w2642_
	);
	LUT4 #(
		.INIT('h9500)
	) name2190 (
		\rEIP_reg[31]/NET0131 ,
		_w2619_,
		_w2622_,
		_w2642_,
		_w2643_
	);
	LUT3 #(
		.INIT('h23)
	) name2191 (
		\DataWidth_reg[1]/NET0131 ,
		\EBX_reg[31]/NET0131 ,
		_w633_,
		_w2644_
	);
	LUT3 #(
		.INIT('h08)
	) name2192 (
		_w570_,
		_w611_,
		_w2644_,
		_w2645_
	);
	LUT3 #(
		.INIT('h45)
	) name2193 (
		_w2641_,
		_w2643_,
		_w2645_,
		_w2646_
	);
	LUT3 #(
		.INIT('h8a)
	) name2194 (
		_w695_,
		_w2639_,
		_w2646_,
		_w2647_
	);
	LUT2 #(
		.INIT('h8)
	) name2195 (
		\DataWidth_reg[1]/NET0131 ,
		\rEIP_reg[31]/NET0131 ,
		_w2648_
	);
	LUT2 #(
		.INIT('h1)
	) name2196 (
		_w1476_,
		_w1485_,
		_w2649_
	);
	LUT2 #(
		.INIT('h1)
	) name2197 (
		_w1463_,
		_w1607_,
		_w2650_
	);
	LUT3 #(
		.INIT('h40)
	) name2198 (
		\PhyAddrPointer_reg[0]/NET0131 ,
		\PhyAddrPointer_reg[1]/NET0131 ,
		_w1569_,
		_w2651_
	);
	LUT4 #(
		.INIT('h4000)
	) name2199 (
		\PhyAddrPointer_reg[0]/NET0131 ,
		\PhyAddrPointer_reg[1]/NET0131 ,
		_w1271_,
		_w1569_,
		_w2652_
	);
	LUT2 #(
		.INIT('h8)
	) name2200 (
		\PhyAddrPointer_reg[22]/NET0131 ,
		_w2652_,
		_w2653_
	);
	LUT4 #(
		.INIT('h8200)
	) name2201 (
		\PhyAddrPointer_reg[22]/NET0131 ,
		\PhyAddrPointer_reg[25]/NET0131 ,
		_w1475_,
		_w2652_,
		_w2654_
	);
	LUT2 #(
		.INIT('h8)
	) name2202 (
		_w2650_,
		_w2654_,
		_w2655_
	);
	LUT3 #(
		.INIT('h40)
	) name2203 (
		_w1626_,
		_w2650_,
		_w2654_,
		_w2656_
	);
	LUT3 #(
		.INIT('h40)
	) name2204 (
		_w1502_,
		_w2656_,
		_w2649_,
		_w2657_
	);
	LUT4 #(
		.INIT('h4105)
	) name2205 (
		\DataWidth_reg[1]/NET0131 ,
		\PhyAddrPointer_reg[1]/NET0131 ,
		\PhyAddrPointer_reg[30]/NET0131 ,
		_w1278_,
		_w2658_
	);
	LUT2 #(
		.INIT('h8)
	) name2206 (
		_w1279_,
		_w2658_,
		_w2659_
	);
	LUT4 #(
		.INIT('ha888)
	) name2207 (
		_w700_,
		_w2648_,
		_w2657_,
		_w2659_,
		_w2660_
	);
	LUT4 #(
		.INIT('hfe25)
	) name2208 (
		\State2_reg[0]/NET0131 ,
		\State2_reg[1]/NET0131 ,
		\State2_reg[2]/NET0131 ,
		\State2_reg[3]/NET0131 ,
		_w2661_
	);
	LUT4 #(
		.INIT('h5f13)
	) name2209 (
		\PhyAddrPointer_reg[31]/NET0131 ,
		\rEIP_reg[31]/NET0131 ,
		_w718_,
		_w2661_,
		_w2662_
	);
	LUT3 #(
		.INIT('hef)
	) name2210 (
		_w2660_,
		_w2647_,
		_w2662_,
		_w2663_
	);
	LUT4 #(
		.INIT('h4080)
	) name2211 (
		\EAX_reg[27]/NET0131 ,
		_w570_,
		_w611_,
		_w2051_,
		_w2664_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name2212 (
		\Datao[27]_pad ,
		_w617_,
		_w2422_,
		_w2664_,
		_w2665_
	);
	LUT4 #(
		.INIT('h3f15)
	) name2213 (
		\Datao[27]_pad ,
		\uWord_reg[11]/NET0131 ,
		_w696_,
		_w2159_,
		_w2666_
	);
	LUT3 #(
		.INIT('h2f)
	) name2214 (
		_w695_,
		_w2665_,
		_w2666_,
		_w2667_
	);
	LUT4 #(
		.INIT('h7030)
	) name2215 (
		_w635_,
		_w695_,
		_w1825_,
		_w1852_,
		_w2668_
	);
	LUT3 #(
		.INIT('h20)
	) name2216 (
		\Datai[2]_pad ,
		READY_n_pad,
		_w611_,
		_w2669_
	);
	LUT4 #(
		.INIT('hec00)
	) name2217 (
		_w514_,
		_w566_,
		_w569_,
		_w2669_,
		_w2670_
	);
	LUT4 #(
		.INIT('h0080)
	) name2218 (
		_w576_,
		_w579_,
		_w605_,
		_w763_,
		_w2671_
	);
	LUT3 #(
		.INIT('h78)
	) name2219 (
		\EAX_reg[0]/NET0131 ,
		\EAX_reg[1]/NET0131 ,
		\EAX_reg[2]/NET0131 ,
		_w2672_
	);
	LUT2 #(
		.INIT('h8)
	) name2220 (
		_w1848_,
		_w2672_,
		_w2673_
	);
	LUT4 #(
		.INIT('haaa8)
	) name2221 (
		_w695_,
		_w2671_,
		_w2670_,
		_w2673_,
		_w2674_
	);
	LUT3 #(
		.INIT('hf2)
	) name2222 (
		\EAX_reg[2]/NET0131 ,
		_w2668_,
		_w2674_,
		_w2675_
	);
	LUT2 #(
		.INIT('h2)
	) name2223 (
		\uWord_reg[11]/NET0131 ,
		_w1825_,
		_w2676_
	);
	LUT3 #(
		.INIT('h20)
	) name2224 (
		\Datai[11]_pad ,
		READY_n_pad,
		_w611_,
		_w2677_
	);
	LUT2 #(
		.INIT('h8)
	) name2225 (
		_w566_,
		_w2677_,
		_w2678_
	);
	LUT4 #(
		.INIT('h000d)
	) name2226 (
		\uWord_reg[11]/NET0131 ,
		_w2058_,
		_w2664_,
		_w2678_,
		_w2679_
	);
	LUT3 #(
		.INIT('hce)
	) name2227 (
		_w695_,
		_w2676_,
		_w2679_,
		_w2680_
	);
	LUT3 #(
		.INIT('h20)
	) name2228 (
		\Datai[3]_pad ,
		READY_n_pad,
		_w611_,
		_w2681_
	);
	LUT4 #(
		.INIT('hec00)
	) name2229 (
		_w514_,
		_w566_,
		_w569_,
		_w2681_,
		_w2682_
	);
	LUT4 #(
		.INIT('h0080)
	) name2230 (
		_w576_,
		_w579_,
		_w605_,
		_w749_,
		_w2683_
	);
	LUT4 #(
		.INIT('h7f80)
	) name2231 (
		\EAX_reg[0]/NET0131 ,
		\EAX_reg[1]/NET0131 ,
		\EAX_reg[2]/NET0131 ,
		\EAX_reg[3]/NET0131 ,
		_w2684_
	);
	LUT2 #(
		.INIT('h8)
	) name2232 (
		_w1848_,
		_w2684_,
		_w2685_
	);
	LUT4 #(
		.INIT('haaa8)
	) name2233 (
		_w695_,
		_w2683_,
		_w2682_,
		_w2685_,
		_w2686_
	);
	LUT3 #(
		.INIT('hf2)
	) name2234 (
		\EAX_reg[3]/NET0131 ,
		_w2668_,
		_w2686_,
		_w2687_
	);
	LUT3 #(
		.INIT('h20)
	) name2235 (
		\Datai[4]_pad ,
		READY_n_pad,
		_w643_,
		_w2688_
	);
	LUT4 #(
		.INIT('h0080)
	) name2236 (
		_w576_,
		_w579_,
		_w605_,
		_w825_,
		_w2689_
	);
	LUT2 #(
		.INIT('h6)
	) name2237 (
		\EAX_reg[4]/NET0131 ,
		_w1827_,
		_w2690_
	);
	LUT2 #(
		.INIT('h8)
	) name2238 (
		_w1848_,
		_w2690_,
		_w2691_
	);
	LUT2 #(
		.INIT('h1)
	) name2239 (
		_w2689_,
		_w2691_,
		_w2692_
	);
	LUT3 #(
		.INIT('h8a)
	) name2240 (
		_w695_,
		_w2688_,
		_w2692_,
		_w2693_
	);
	LUT3 #(
		.INIT('hf2)
	) name2241 (
		\EAX_reg[4]/NET0131 ,
		_w2668_,
		_w2693_,
		_w2694_
	);
	LUT3 #(
		.INIT('h20)
	) name2242 (
		\Datai[5]_pad ,
		READY_n_pad,
		_w643_,
		_w2695_
	);
	LUT4 #(
		.INIT('h0080)
	) name2243 (
		_w576_,
		_w579_,
		_w605_,
		_w810_,
		_w2696_
	);
	LUT3 #(
		.INIT('h6c)
	) name2244 (
		\EAX_reg[4]/NET0131 ,
		\EAX_reg[5]/NET0131 ,
		_w1827_,
		_w2697_
	);
	LUT2 #(
		.INIT('h8)
	) name2245 (
		_w1848_,
		_w2697_,
		_w2698_
	);
	LUT2 #(
		.INIT('h1)
	) name2246 (
		_w2696_,
		_w2698_,
		_w2699_
	);
	LUT3 #(
		.INIT('h8a)
	) name2247 (
		_w695_,
		_w2695_,
		_w2699_,
		_w2700_
	);
	LUT3 #(
		.INIT('hf2)
	) name2248 (
		\EAX_reg[5]/NET0131 ,
		_w2668_,
		_w2700_,
		_w2701_
	);
	LUT3 #(
		.INIT('h20)
	) name2249 (
		\Datai[6]_pad ,
		READY_n_pad,
		_w643_,
		_w2702_
	);
	LUT4 #(
		.INIT('h0080)
	) name2250 (
		_w576_,
		_w579_,
		_w605_,
		_w857_,
		_w2703_
	);
	LUT4 #(
		.INIT('h78f0)
	) name2251 (
		\EAX_reg[4]/NET0131 ,
		\EAX_reg[5]/NET0131 ,
		\EAX_reg[6]/NET0131 ,
		_w1827_,
		_w2704_
	);
	LUT2 #(
		.INIT('h8)
	) name2252 (
		_w1848_,
		_w2704_,
		_w2705_
	);
	LUT2 #(
		.INIT('h1)
	) name2253 (
		_w2703_,
		_w2705_,
		_w2706_
	);
	LUT3 #(
		.INIT('h8a)
	) name2254 (
		_w695_,
		_w2702_,
		_w2706_,
		_w2707_
	);
	LUT3 #(
		.INIT('hf2)
	) name2255 (
		\EAX_reg[6]/NET0131 ,
		_w2668_,
		_w2707_,
		_w2708_
	);
	LUT3 #(
		.INIT('h20)
	) name2256 (
		\Datai[7]_pad ,
		READY_n_pad,
		_w643_,
		_w2709_
	);
	LUT4 #(
		.INIT('h0080)
	) name2257 (
		_w576_,
		_w579_,
		_w605_,
		_w844_,
		_w2710_
	);
	LUT2 #(
		.INIT('h6)
	) name2258 (
		\EAX_reg[7]/NET0131 ,
		_w1828_,
		_w2711_
	);
	LUT2 #(
		.INIT('h8)
	) name2259 (
		_w1848_,
		_w2711_,
		_w2712_
	);
	LUT2 #(
		.INIT('h1)
	) name2260 (
		_w2710_,
		_w2712_,
		_w2713_
	);
	LUT3 #(
		.INIT('h8a)
	) name2261 (
		_w695_,
		_w2709_,
		_w2713_,
		_w2714_
	);
	LUT3 #(
		.INIT('hf2)
	) name2262 (
		\EAX_reg[7]/NET0131 ,
		_w2668_,
		_w2714_,
		_w2715_
	);
	LUT3 #(
		.INIT('h20)
	) name2263 (
		\Datai[9]_pad ,
		READY_n_pad,
		_w643_,
		_w2716_
	);
	LUT4 #(
		.INIT('h135f)
	) name2264 (
		\InstQueue_reg[4][1]/NET0131 ,
		\InstQueue_reg[7][1]/NET0131 ,
		_w474_,
		_w467_,
		_w2717_
	);
	LUT4 #(
		.INIT('h153f)
	) name2265 (
		\InstQueue_reg[12][1]/NET0131 ,
		\InstQueue_reg[8][1]/NET0131 ,
		_w461_,
		_w471_,
		_w2718_
	);
	LUT4 #(
		.INIT('h153f)
	) name2266 (
		\InstQueue_reg[10][1]/NET0131 ,
		\InstQueue_reg[13][1]/NET0131 ,
		_w458_,
		_w468_,
		_w2719_
	);
	LUT4 #(
		.INIT('h135f)
	) name2267 (
		\InstQueue_reg[1][1]/NET0131 ,
		\InstQueue_reg[9][1]/NET0131 ,
		_w473_,
		_w477_,
		_w2720_
	);
	LUT4 #(
		.INIT('h8000)
	) name2268 (
		_w2719_,
		_w2720_,
		_w2717_,
		_w2718_,
		_w2721_
	);
	LUT4 #(
		.INIT('h153f)
	) name2269 (
		\InstQueue_reg[14][1]/NET0131 ,
		\InstQueue_reg[15][1]/NET0131 ,
		_w456_,
		_w470_,
		_w2722_
	);
	LUT4 #(
		.INIT('h135f)
	) name2270 (
		\InstQueue_reg[3][1]/NET0131 ,
		\InstQueue_reg[5][1]/NET0131 ,
		_w453_,
		_w476_,
		_w2723_
	);
	LUT4 #(
		.INIT('h135f)
	) name2271 (
		\InstQueue_reg[0][1]/NET0131 ,
		\InstQueue_reg[11][1]/NET0131 ,
		_w460_,
		_w454_,
		_w2724_
	);
	LUT4 #(
		.INIT('h135f)
	) name2272 (
		\InstQueue_reg[2][1]/NET0131 ,
		\InstQueue_reg[6][1]/NET0131 ,
		_w463_,
		_w464_,
		_w2725_
	);
	LUT4 #(
		.INIT('h8000)
	) name2273 (
		_w2724_,
		_w2725_,
		_w2722_,
		_w2723_,
		_w2726_
	);
	LUT2 #(
		.INIT('h8)
	) name2274 (
		_w2721_,
		_w2726_,
		_w2727_
	);
	LUT4 #(
		.INIT('h0080)
	) name2275 (
		_w576_,
		_w579_,
		_w605_,
		_w2727_,
		_w2728_
	);
	LUT4 #(
		.INIT('h78f0)
	) name2276 (
		\EAX_reg[7]/NET0131 ,
		\EAX_reg[8]/NET0131 ,
		\EAX_reg[9]/NET0131 ,
		_w1828_,
		_w2729_
	);
	LUT2 #(
		.INIT('h8)
	) name2277 (
		_w1848_,
		_w2729_,
		_w2730_
	);
	LUT2 #(
		.INIT('h1)
	) name2278 (
		_w2728_,
		_w2730_,
		_w2731_
	);
	LUT3 #(
		.INIT('h8a)
	) name2279 (
		_w695_,
		_w2716_,
		_w2731_,
		_w2732_
	);
	LUT3 #(
		.INIT('hf2)
	) name2280 (
		\EAX_reg[9]/NET0131 ,
		_w2668_,
		_w2732_,
		_w2733_
	);
	LUT3 #(
		.INIT('h20)
	) name2281 (
		\Datai[8]_pad ,
		READY_n_pad,
		_w643_,
		_w2734_
	);
	LUT4 #(
		.INIT('h153f)
	) name2282 (
		\InstQueue_reg[14][0]/NET0131 ,
		\InstQueue_reg[6][0]/NET0131 ,
		_w464_,
		_w470_,
		_w2735_
	);
	LUT4 #(
		.INIT('h153f)
	) name2283 (
		\InstQueue_reg[13][0]/NET0131 ,
		\InstQueue_reg[2][0]/NET0131 ,
		_w463_,
		_w458_,
		_w2736_
	);
	LUT4 #(
		.INIT('h153f)
	) name2284 (
		\InstQueue_reg[10][0]/NET0131 ,
		\InstQueue_reg[8][0]/NET0131 ,
		_w461_,
		_w468_,
		_w2737_
	);
	LUT4 #(
		.INIT('h135f)
	) name2285 (
		\InstQueue_reg[1][0]/NET0131 ,
		\InstQueue_reg[9][0]/NET0131 ,
		_w473_,
		_w477_,
		_w2738_
	);
	LUT4 #(
		.INIT('h8000)
	) name2286 (
		_w2737_,
		_w2738_,
		_w2735_,
		_w2736_,
		_w2739_
	);
	LUT4 #(
		.INIT('h135f)
	) name2287 (
		\InstQueue_reg[11][0]/NET0131 ,
		\InstQueue_reg[15][0]/NET0131 ,
		_w454_,
		_w456_,
		_w2740_
	);
	LUT4 #(
		.INIT('h135f)
	) name2288 (
		\InstQueue_reg[4][0]/NET0131 ,
		\InstQueue_reg[7][0]/NET0131 ,
		_w474_,
		_w467_,
		_w2741_
	);
	LUT4 #(
		.INIT('h135f)
	) name2289 (
		\InstQueue_reg[0][0]/NET0131 ,
		\InstQueue_reg[5][0]/NET0131 ,
		_w460_,
		_w476_,
		_w2742_
	);
	LUT4 #(
		.INIT('h153f)
	) name2290 (
		\InstQueue_reg[12][0]/NET0131 ,
		\InstQueue_reg[3][0]/NET0131 ,
		_w453_,
		_w471_,
		_w2743_
	);
	LUT4 #(
		.INIT('h8000)
	) name2291 (
		_w2742_,
		_w2743_,
		_w2740_,
		_w2741_,
		_w2744_
	);
	LUT2 #(
		.INIT('h8)
	) name2292 (
		_w2739_,
		_w2744_,
		_w2745_
	);
	LUT4 #(
		.INIT('h0080)
	) name2293 (
		_w576_,
		_w579_,
		_w605_,
		_w2745_,
		_w2746_
	);
	LUT3 #(
		.INIT('h6c)
	) name2294 (
		\EAX_reg[7]/NET0131 ,
		\EAX_reg[8]/NET0131 ,
		_w1828_,
		_w2747_
	);
	LUT2 #(
		.INIT('h8)
	) name2295 (
		_w1848_,
		_w2747_,
		_w2748_
	);
	LUT2 #(
		.INIT('h1)
	) name2296 (
		_w2746_,
		_w2748_,
		_w2749_
	);
	LUT3 #(
		.INIT('h8a)
	) name2297 (
		_w695_,
		_w2734_,
		_w2749_,
		_w2750_
	);
	LUT3 #(
		.INIT('hf2)
	) name2298 (
		\EAX_reg[8]/NET0131 ,
		_w2668_,
		_w2750_,
		_w2751_
	);
	LUT4 #(
		.INIT('hec00)
	) name2299 (
		_w514_,
		_w566_,
		_w569_,
		_w2677_,
		_w2752_
	);
	LUT2 #(
		.INIT('h2)
	) name2300 (
		_w1848_,
		_w1831_,
		_w2753_
	);
	LUT3 #(
		.INIT('h48)
	) name2301 (
		\EAX_reg[11]/NET0131 ,
		_w1848_,
		_w1830_,
		_w2754_
	);
	LUT4 #(
		.INIT('h135f)
	) name2302 (
		\InstQueue_reg[13][3]/NET0131 ,
		\InstQueue_reg[7][3]/NET0131 ,
		_w458_,
		_w467_,
		_w2755_
	);
	LUT4 #(
		.INIT('h135f)
	) name2303 (
		\InstQueue_reg[10][3]/NET0131 ,
		\InstQueue_reg[12][3]/NET0131 ,
		_w468_,
		_w471_,
		_w2756_
	);
	LUT4 #(
		.INIT('h135f)
	) name2304 (
		\InstQueue_reg[2][3]/NET0131 ,
		\InstQueue_reg[3][3]/NET0131 ,
		_w463_,
		_w453_,
		_w2757_
	);
	LUT4 #(
		.INIT('h135f)
	) name2305 (
		\InstQueue_reg[1][3]/NET0131 ,
		\InstQueue_reg[9][3]/NET0131 ,
		_w473_,
		_w477_,
		_w2758_
	);
	LUT4 #(
		.INIT('h8000)
	) name2306 (
		_w2757_,
		_w2758_,
		_w2755_,
		_w2756_,
		_w2759_
	);
	LUT4 #(
		.INIT('h135f)
	) name2307 (
		\InstQueue_reg[11][3]/NET0131 ,
		\InstQueue_reg[4][3]/NET0131 ,
		_w454_,
		_w474_,
		_w2760_
	);
	LUT4 #(
		.INIT('h153f)
	) name2308 (
		\InstQueue_reg[6][3]/NET0131 ,
		\InstQueue_reg[8][3]/NET0131 ,
		_w461_,
		_w464_,
		_w2761_
	);
	LUT4 #(
		.INIT('h135f)
	) name2309 (
		\InstQueue_reg[0][3]/NET0131 ,
		\InstQueue_reg[15][3]/NET0131 ,
		_w460_,
		_w456_,
		_w2762_
	);
	LUT4 #(
		.INIT('h153f)
	) name2310 (
		\InstQueue_reg[14][3]/NET0131 ,
		\InstQueue_reg[5][3]/NET0131 ,
		_w476_,
		_w470_,
		_w2763_
	);
	LUT4 #(
		.INIT('h8000)
	) name2311 (
		_w2762_,
		_w2763_,
		_w2760_,
		_w2761_,
		_w2764_
	);
	LUT2 #(
		.INIT('h8)
	) name2312 (
		_w2759_,
		_w2764_,
		_w2765_
	);
	LUT4 #(
		.INIT('h0080)
	) name2313 (
		_w576_,
		_w579_,
		_w605_,
		_w2765_,
		_w2766_
	);
	LUT4 #(
		.INIT('haaa8)
	) name2314 (
		_w695_,
		_w2754_,
		_w2766_,
		_w2752_,
		_w2767_
	);
	LUT3 #(
		.INIT('hf2)
	) name2315 (
		\EAX_reg[11]/NET0131 ,
		_w2668_,
		_w2767_,
		_w2768_
	);
	LUT3 #(
		.INIT('h80)
	) name2316 (
		_w552_,
		_w576_,
		_w2435_,
		_w2769_
	);
	LUT3 #(
		.INIT('h07)
	) name2317 (
		\EBX_reg[25]/NET0131 ,
		_w1975_,
		_w2769_,
		_w2770_
	);
	LUT4 #(
		.INIT('hb700)
	) name2318 (
		\EBX_reg[25]/NET0131 ,
		_w590_,
		_w1972_,
		_w2770_,
		_w2771_
	);
	LUT2 #(
		.INIT('h2)
	) name2319 (
		\EBX_reg[25]/NET0131 ,
		_w1825_,
		_w2772_
	);
	LUT3 #(
		.INIT('hf2)
	) name2320 (
		_w695_,
		_w2771_,
		_w2772_,
		_w2773_
	);
	LUT4 #(
		.INIT('h135f)
	) name2321 (
		\InstQueue_reg[4][2]/NET0131 ,
		\InstQueue_reg[7][2]/NET0131 ,
		_w474_,
		_w467_,
		_w2774_
	);
	LUT4 #(
		.INIT('h153f)
	) name2322 (
		\InstQueue_reg[12][2]/NET0131 ,
		\InstQueue_reg[8][2]/NET0131 ,
		_w461_,
		_w471_,
		_w2775_
	);
	LUT4 #(
		.INIT('h153f)
	) name2323 (
		\InstQueue_reg[10][2]/NET0131 ,
		\InstQueue_reg[13][2]/NET0131 ,
		_w458_,
		_w468_,
		_w2776_
	);
	LUT4 #(
		.INIT('h135f)
	) name2324 (
		\InstQueue_reg[1][2]/NET0131 ,
		\InstQueue_reg[9][2]/NET0131 ,
		_w473_,
		_w477_,
		_w2777_
	);
	LUT4 #(
		.INIT('h8000)
	) name2325 (
		_w2776_,
		_w2777_,
		_w2774_,
		_w2775_,
		_w2778_
	);
	LUT4 #(
		.INIT('h153f)
	) name2326 (
		\InstQueue_reg[14][2]/NET0131 ,
		\InstQueue_reg[15][2]/NET0131 ,
		_w456_,
		_w470_,
		_w2779_
	);
	LUT4 #(
		.INIT('h135f)
	) name2327 (
		\InstQueue_reg[3][2]/NET0131 ,
		\InstQueue_reg[5][2]/NET0131 ,
		_w453_,
		_w476_,
		_w2780_
	);
	LUT4 #(
		.INIT('h135f)
	) name2328 (
		\InstQueue_reg[0][2]/NET0131 ,
		\InstQueue_reg[11][2]/NET0131 ,
		_w460_,
		_w454_,
		_w2781_
	);
	LUT4 #(
		.INIT('h135f)
	) name2329 (
		\InstQueue_reg[2][2]/NET0131 ,
		\InstQueue_reg[6][2]/NET0131 ,
		_w463_,
		_w464_,
		_w2782_
	);
	LUT4 #(
		.INIT('h8000)
	) name2330 (
		_w2781_,
		_w2782_,
		_w2779_,
		_w2780_,
		_w2783_
	);
	LUT2 #(
		.INIT('h8)
	) name2331 (
		_w2778_,
		_w2783_,
		_w2784_
	);
	LUT4 #(
		.INIT('h0080)
	) name2332 (
		_w576_,
		_w579_,
		_w605_,
		_w2784_,
		_w2785_
	);
	LUT3 #(
		.INIT('h48)
	) name2333 (
		\EAX_reg[10]/NET0131 ,
		_w1848_,
		_w1829_,
		_w2786_
	);
	LUT4 #(
		.INIT('h0007)
	) name2334 (
		_w643_,
		_w2032_,
		_w2785_,
		_w2786_,
		_w2787_
	);
	LUT2 #(
		.INIT('h2)
	) name2335 (
		_w695_,
		_w2787_,
		_w2788_
	);
	LUT3 #(
		.INIT('hf2)
	) name2336 (
		\EAX_reg[10]/NET0131 ,
		_w2668_,
		_w2788_,
		_w2789_
	);
	LUT2 #(
		.INIT('h2)
	) name2337 (
		\EAX_reg[12]/NET0131 ,
		_w1825_,
		_w2790_
	);
	LUT4 #(
		.INIT('haa8a)
	) name2338 (
		\EAX_reg[12]/NET0131 ,
		_w635_,
		_w1852_,
		_w2753_,
		_w2791_
	);
	LUT3 #(
		.INIT('h20)
	) name2339 (
		\Datai[12]_pad ,
		READY_n_pad,
		_w643_,
		_w2792_
	);
	LUT2 #(
		.INIT('h2)
	) name2340 (
		_w1848_,
		_w1832_,
		_w2793_
	);
	LUT3 #(
		.INIT('h40)
	) name2341 (
		\EAX_reg[12]/NET0131 ,
		_w1848_,
		_w1831_,
		_w2794_
	);
	LUT4 #(
		.INIT('h135f)
	) name2342 (
		\InstQueue_reg[4][4]/NET0131 ,
		\InstQueue_reg[7][4]/NET0131 ,
		_w474_,
		_w467_,
		_w2795_
	);
	LUT4 #(
		.INIT('h153f)
	) name2343 (
		\InstQueue_reg[12][4]/NET0131 ,
		\InstQueue_reg[6][4]/NET0131 ,
		_w464_,
		_w471_,
		_w2796_
	);
	LUT4 #(
		.INIT('h135f)
	) name2344 (
		\InstQueue_reg[2][4]/NET0131 ,
		\InstQueue_reg[3][4]/NET0131 ,
		_w463_,
		_w453_,
		_w2797_
	);
	LUT4 #(
		.INIT('h153f)
	) name2345 (
		\InstQueue_reg[10][4]/NET0131 ,
		\InstQueue_reg[1][4]/NET0131 ,
		_w473_,
		_w468_,
		_w2798_
	);
	LUT4 #(
		.INIT('h8000)
	) name2346 (
		_w2797_,
		_w2798_,
		_w2795_,
		_w2796_,
		_w2799_
	);
	LUT4 #(
		.INIT('h153f)
	) name2347 (
		\InstQueue_reg[14][4]/NET0131 ,
		\InstQueue_reg[9][4]/NET0131 ,
		_w477_,
		_w470_,
		_w2800_
	);
	LUT4 #(
		.INIT('h153f)
	) name2348 (
		\InstQueue_reg[13][4]/NET0131 ,
		\InstQueue_reg[15][4]/NET0131 ,
		_w456_,
		_w458_,
		_w2801_
	);
	LUT4 #(
		.INIT('h135f)
	) name2349 (
		\InstQueue_reg[0][4]/NET0131 ,
		\InstQueue_reg[11][4]/NET0131 ,
		_w460_,
		_w454_,
		_w2802_
	);
	LUT4 #(
		.INIT('h153f)
	) name2350 (
		\InstQueue_reg[5][4]/NET0131 ,
		\InstQueue_reg[8][4]/NET0131 ,
		_w461_,
		_w476_,
		_w2803_
	);
	LUT4 #(
		.INIT('h8000)
	) name2351 (
		_w2802_,
		_w2803_,
		_w2800_,
		_w2801_,
		_w2804_
	);
	LUT2 #(
		.INIT('h8)
	) name2352 (
		_w2799_,
		_w2804_,
		_w2805_
	);
	LUT4 #(
		.INIT('h0080)
	) name2353 (
		_w576_,
		_w579_,
		_w605_,
		_w2805_,
		_w2806_
	);
	LUT2 #(
		.INIT('h1)
	) name2354 (
		_w2794_,
		_w2806_,
		_w2807_
	);
	LUT2 #(
		.INIT('h4)
	) name2355 (
		_w2792_,
		_w2807_,
		_w2808_
	);
	LUT4 #(
		.INIT('hecee)
	) name2356 (
		_w695_,
		_w2790_,
		_w2791_,
		_w2808_,
		_w2809_
	);
	LUT2 #(
		.INIT('h2)
	) name2357 (
		\EAX_reg[13]/NET0131 ,
		_w1825_,
		_w2810_
	);
	LUT4 #(
		.INIT('h008d)
	) name2358 (
		_w580_,
		_w605_,
		_w1850_,
		_w2793_,
		_w2811_
	);
	LUT4 #(
		.INIT('h3533)
	) name2359 (
		\Datai[13]_pad ,
		\EAX_reg[13]/NET0131 ,
		READY_n_pad,
		_w611_,
		_w2812_
	);
	LUT4 #(
		.INIT('h00ec)
	) name2360 (
		_w514_,
		_w566_,
		_w569_,
		_w2812_,
		_w2813_
	);
	LUT3 #(
		.INIT('h40)
	) name2361 (
		\EAX_reg[13]/NET0131 ,
		_w1848_,
		_w1832_,
		_w2814_
	);
	LUT4 #(
		.INIT('h135f)
	) name2362 (
		\InstQueue_reg[4][5]/NET0131 ,
		\InstQueue_reg[7][5]/NET0131 ,
		_w474_,
		_w467_,
		_w2815_
	);
	LUT4 #(
		.INIT('h153f)
	) name2363 (
		\InstQueue_reg[12][5]/NET0131 ,
		\InstQueue_reg[8][5]/NET0131 ,
		_w461_,
		_w471_,
		_w2816_
	);
	LUT4 #(
		.INIT('h153f)
	) name2364 (
		\InstQueue_reg[10][5]/NET0131 ,
		\InstQueue_reg[13][5]/NET0131 ,
		_w458_,
		_w468_,
		_w2817_
	);
	LUT4 #(
		.INIT('h135f)
	) name2365 (
		\InstQueue_reg[1][5]/NET0131 ,
		\InstQueue_reg[9][5]/NET0131 ,
		_w473_,
		_w477_,
		_w2818_
	);
	LUT4 #(
		.INIT('h8000)
	) name2366 (
		_w2817_,
		_w2818_,
		_w2815_,
		_w2816_,
		_w2819_
	);
	LUT4 #(
		.INIT('h153f)
	) name2367 (
		\InstQueue_reg[14][5]/NET0131 ,
		\InstQueue_reg[15][5]/NET0131 ,
		_w456_,
		_w470_,
		_w2820_
	);
	LUT4 #(
		.INIT('h135f)
	) name2368 (
		\InstQueue_reg[3][5]/NET0131 ,
		\InstQueue_reg[5][5]/NET0131 ,
		_w453_,
		_w476_,
		_w2821_
	);
	LUT4 #(
		.INIT('h135f)
	) name2369 (
		\InstQueue_reg[0][5]/NET0131 ,
		\InstQueue_reg[11][5]/NET0131 ,
		_w460_,
		_w454_,
		_w2822_
	);
	LUT4 #(
		.INIT('h135f)
	) name2370 (
		\InstQueue_reg[2][5]/NET0131 ,
		\InstQueue_reg[6][5]/NET0131 ,
		_w463_,
		_w464_,
		_w2823_
	);
	LUT4 #(
		.INIT('h8000)
	) name2371 (
		_w2822_,
		_w2823_,
		_w2820_,
		_w2821_,
		_w2824_
	);
	LUT2 #(
		.INIT('h8)
	) name2372 (
		_w2819_,
		_w2824_,
		_w2825_
	);
	LUT4 #(
		.INIT('h0080)
	) name2373 (
		_w576_,
		_w579_,
		_w605_,
		_w2825_,
		_w2826_
	);
	LUT3 #(
		.INIT('h01)
	) name2374 (
		_w2814_,
		_w2826_,
		_w2813_,
		_w2827_
	);
	LUT4 #(
		.INIT('h08cc)
	) name2375 (
		\EAX_reg[13]/NET0131 ,
		_w695_,
		_w2811_,
		_w2827_,
		_w2828_
	);
	LUT2 #(
		.INIT('he)
	) name2376 (
		_w2810_,
		_w2828_,
		_w2829_
	);
	LUT2 #(
		.INIT('h2)
	) name2377 (
		\EAX_reg[14]/NET0131 ,
		_w1825_,
		_w2830_
	);
	LUT2 #(
		.INIT('h2)
	) name2378 (
		_w1848_,
		_w1833_,
		_w2831_
	);
	LUT4 #(
		.INIT('haa8a)
	) name2379 (
		\EAX_reg[14]/NET0131 ,
		_w635_,
		_w1852_,
		_w2831_,
		_w2832_
	);
	LUT3 #(
		.INIT('h20)
	) name2380 (
		\Datai[14]_pad ,
		READY_n_pad,
		_w643_,
		_w2833_
	);
	LUT4 #(
		.INIT('h135f)
	) name2381 (
		\InstQueue_reg[6][6]/NET0131 ,
		\InstQueue_reg[7][6]/NET0131 ,
		_w464_,
		_w467_,
		_w2834_
	);
	LUT4 #(
		.INIT('h153f)
	) name2382 (
		\InstQueue_reg[12][6]/NET0131 ,
		\InstQueue_reg[15][6]/NET0131 ,
		_w456_,
		_w471_,
		_w2835_
	);
	LUT4 #(
		.INIT('h135f)
	) name2383 (
		\InstQueue_reg[2][6]/NET0131 ,
		\InstQueue_reg[3][6]/NET0131 ,
		_w463_,
		_w453_,
		_w2836_
	);
	LUT4 #(
		.INIT('h135f)
	) name2384 (
		\InstQueue_reg[1][6]/NET0131 ,
		\InstQueue_reg[9][6]/NET0131 ,
		_w473_,
		_w477_,
		_w2837_
	);
	LUT4 #(
		.INIT('h8000)
	) name2385 (
		_w2836_,
		_w2837_,
		_w2834_,
		_w2835_,
		_w2838_
	);
	LUT4 #(
		.INIT('h135f)
	) name2386 (
		\InstQueue_reg[11][6]/NET0131 ,
		\InstQueue_reg[4][6]/NET0131 ,
		_w454_,
		_w474_,
		_w2839_
	);
	LUT4 #(
		.INIT('h153f)
	) name2387 (
		\InstQueue_reg[13][6]/NET0131 ,
		\InstQueue_reg[8][6]/NET0131 ,
		_w461_,
		_w458_,
		_w2840_
	);
	LUT4 #(
		.INIT('h135f)
	) name2388 (
		\InstQueue_reg[0][6]/NET0131 ,
		\InstQueue_reg[10][6]/NET0131 ,
		_w460_,
		_w468_,
		_w2841_
	);
	LUT4 #(
		.INIT('h153f)
	) name2389 (
		\InstQueue_reg[14][6]/NET0131 ,
		\InstQueue_reg[5][6]/NET0131 ,
		_w476_,
		_w470_,
		_w2842_
	);
	LUT4 #(
		.INIT('h8000)
	) name2390 (
		_w2841_,
		_w2842_,
		_w2839_,
		_w2840_,
		_w2843_
	);
	LUT2 #(
		.INIT('h8)
	) name2391 (
		_w2838_,
		_w2843_,
		_w2844_
	);
	LUT4 #(
		.INIT('h0080)
	) name2392 (
		_w576_,
		_w579_,
		_w605_,
		_w2844_,
		_w2845_
	);
	LUT3 #(
		.INIT('h40)
	) name2393 (
		\EAX_reg[14]/NET0131 ,
		_w1848_,
		_w1833_,
		_w2846_
	);
	LUT2 #(
		.INIT('h1)
	) name2394 (
		_w2845_,
		_w2846_,
		_w2847_
	);
	LUT2 #(
		.INIT('h4)
	) name2395 (
		_w2833_,
		_w2847_,
		_w2848_
	);
	LUT4 #(
		.INIT('hecee)
	) name2396 (
		_w695_,
		_w2830_,
		_w2832_,
		_w2848_,
		_w2849_
	);
	LUT2 #(
		.INIT('h2)
	) name2397 (
		\EAX_reg[15]/NET0131 ,
		_w1825_,
		_w2850_
	);
	LUT2 #(
		.INIT('h2)
	) name2398 (
		_w1848_,
		_w1834_,
		_w2851_
	);
	LUT4 #(
		.INIT('haa8a)
	) name2399 (
		\EAX_reg[15]/NET0131 ,
		_w635_,
		_w1852_,
		_w2851_,
		_w2852_
	);
	LUT3 #(
		.INIT('h40)
	) name2400 (
		\EAX_reg[15]/NET0131 ,
		_w1848_,
		_w1834_,
		_w2853_
	);
	LUT4 #(
		.INIT('h135f)
	) name2401 (
		\InstQueue_reg[6][7]/NET0131 ,
		\InstQueue_reg[7][7]/NET0131 ,
		_w464_,
		_w467_,
		_w2854_
	);
	LUT4 #(
		.INIT('h153f)
	) name2402 (
		\InstQueue_reg[15][7]/NET0131 ,
		\InstQueue_reg[3][7]/NET0131 ,
		_w453_,
		_w456_,
		_w2855_
	);
	LUT4 #(
		.INIT('h153f)
	) name2403 (
		\InstQueue_reg[2][7]/NET0131 ,
		\InstQueue_reg[8][7]/NET0131 ,
		_w461_,
		_w463_,
		_w2856_
	);
	LUT4 #(
		.INIT('h135f)
	) name2404 (
		\InstQueue_reg[1][7]/NET0131 ,
		\InstQueue_reg[9][7]/NET0131 ,
		_w473_,
		_w477_,
		_w2857_
	);
	LUT4 #(
		.INIT('h8000)
	) name2405 (
		_w2856_,
		_w2857_,
		_w2854_,
		_w2855_,
		_w2858_
	);
	LUT4 #(
		.INIT('h153f)
	) name2406 (
		\InstQueue_reg[14][7]/NET0131 ,
		\InstQueue_reg[4][7]/NET0131 ,
		_w474_,
		_w470_,
		_w2859_
	);
	LUT4 #(
		.INIT('h153f)
	) name2407 (
		\InstQueue_reg[12][7]/NET0131 ,
		\InstQueue_reg[13][7]/NET0131 ,
		_w458_,
		_w471_,
		_w2860_
	);
	LUT4 #(
		.INIT('h135f)
	) name2408 (
		\InstQueue_reg[0][7]/NET0131 ,
		\InstQueue_reg[10][7]/NET0131 ,
		_w460_,
		_w468_,
		_w2861_
	);
	LUT4 #(
		.INIT('h135f)
	) name2409 (
		\InstQueue_reg[11][7]/NET0131 ,
		\InstQueue_reg[5][7]/NET0131 ,
		_w454_,
		_w476_,
		_w2862_
	);
	LUT4 #(
		.INIT('h8000)
	) name2410 (
		_w2861_,
		_w2862_,
		_w2859_,
		_w2860_,
		_w2863_
	);
	LUT2 #(
		.INIT('h8)
	) name2411 (
		_w2858_,
		_w2863_,
		_w2864_
	);
	LUT4 #(
		.INIT('h0080)
	) name2412 (
		_w576_,
		_w579_,
		_w605_,
		_w2864_,
		_w2865_
	);
	LUT4 #(
		.INIT('h00df)
	) name2413 (
		\Datai[15]_pad ,
		READY_n_pad,
		_w643_,
		_w2865_,
		_w2866_
	);
	LUT2 #(
		.INIT('h4)
	) name2414 (
		_w2853_,
		_w2866_,
		_w2867_
	);
	LUT4 #(
		.INIT('hecee)
	) name2415 (
		_w695_,
		_w2850_,
		_w2852_,
		_w2867_,
		_w2868_
	);
	LUT3 #(
		.INIT('h20)
	) name2416 (
		\Datai[1]_pad ,
		READY_n_pad,
		_w611_,
		_w2869_
	);
	LUT4 #(
		.INIT('hec00)
	) name2417 (
		_w514_,
		_w566_,
		_w569_,
		_w2869_,
		_w2870_
	);
	LUT4 #(
		.INIT('h0080)
	) name2418 (
		_w576_,
		_w579_,
		_w605_,
		_w780_,
		_w2871_
	);
	LUT2 #(
		.INIT('h6)
	) name2419 (
		\EAX_reg[0]/NET0131 ,
		\EAX_reg[1]/NET0131 ,
		_w2872_
	);
	LUT2 #(
		.INIT('h8)
	) name2420 (
		_w1848_,
		_w2872_,
		_w2873_
	);
	LUT4 #(
		.INIT('haaa8)
	) name2421 (
		_w695_,
		_w2871_,
		_w2870_,
		_w2873_,
		_w2874_
	);
	LUT3 #(
		.INIT('hf2)
	) name2422 (
		\EAX_reg[1]/NET0131 ,
		_w2668_,
		_w2874_,
		_w2875_
	);
	LUT4 #(
		.INIT('h78f0)
	) name2423 (
		\Datai[25]_pad ,
		\Datai[26]_pad ,
		\Datai[27]_pad ,
		_w2196_,
		_w2876_
	);
	LUT4 #(
		.INIT('h6c00)
	) name2424 (
		\Datai[18]_pad ,
		\Datai[19]_pad ,
		_w2199_,
		_w2203_,
		_w2877_
	);
	LUT4 #(
		.INIT('haa80)
	) name2425 (
		\DataWidth_reg[1]/NET0131 ,
		_w2187_,
		_w2876_,
		_w2877_,
		_w2878_
	);
	LUT4 #(
		.INIT('h5553)
	) name2426 (
		\Datai[3]_pad ,
		\InstQueue_reg[0][3]/NET0131 ,
		_w2205_,
		_w2207_,
		_w2879_
	);
	LUT2 #(
		.INIT('h1)
	) name2427 (
		_w2211_,
		_w2879_,
		_w2880_
	);
	LUT4 #(
		.INIT('hc055)
	) name2428 (
		\InstQueue_reg[0][3]/NET0131 ,
		_w520_,
		_w525_,
		_w2205_,
		_w2881_
	);
	LUT2 #(
		.INIT('h2)
	) name2429 (
		\InstQueue_reg[0][3]/NET0131 ,
		_w2215_,
		_w2882_
	);
	LUT3 #(
		.INIT('h0d)
	) name2430 (
		_w706_,
		_w2879_,
		_w2882_,
		_w2883_
	);
	LUT3 #(
		.INIT('hd0)
	) name2431 (
		_w722_,
		_w2881_,
		_w2883_,
		_w2884_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name2432 (
		_w700_,
		_w2878_,
		_w2880_,
		_w2884_,
		_w2885_
	);
	LUT4 #(
		.INIT('h78f0)
	) name2433 (
		\Datai[28]_pad ,
		\Datai[29]_pad ,
		\Datai[30]_pad ,
		_w2197_,
		_w2886_
	);
	LUT4 #(
		.INIT('h6c00)
	) name2434 (
		\Datai[21]_pad ,
		\Datai[22]_pad ,
		_w2200_,
		_w2203_,
		_w2887_
	);
	LUT4 #(
		.INIT('haa80)
	) name2435 (
		\DataWidth_reg[1]/NET0131 ,
		_w2187_,
		_w2886_,
		_w2887_,
		_w2888_
	);
	LUT4 #(
		.INIT('h5553)
	) name2436 (
		\Datai[6]_pad ,
		\InstQueue_reg[0][6]/NET0131 ,
		_w2205_,
		_w2207_,
		_w2889_
	);
	LUT2 #(
		.INIT('h1)
	) name2437 (
		_w2211_,
		_w2889_,
		_w2890_
	);
	LUT4 #(
		.INIT('hc055)
	) name2438 (
		\InstQueue_reg[0][6]/NET0131 ,
		_w485_,
		_w490_,
		_w2205_,
		_w2891_
	);
	LUT2 #(
		.INIT('h2)
	) name2439 (
		\InstQueue_reg[0][6]/NET0131 ,
		_w2215_,
		_w2892_
	);
	LUT3 #(
		.INIT('h0d)
	) name2440 (
		_w706_,
		_w2889_,
		_w2892_,
		_w2893_
	);
	LUT3 #(
		.INIT('hd0)
	) name2441 (
		_w722_,
		_w2891_,
		_w2893_,
		_w2894_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name2442 (
		_w700_,
		_w2888_,
		_w2890_,
		_w2894_,
		_w2895_
	);
	LUT4 #(
		.INIT('h6c00)
	) name2443 (
		\Datai[18]_pad ,
		\Datai[19]_pad ,
		_w2199_,
		_w2222_,
		_w2896_
	);
	LUT4 #(
		.INIT('haa80)
	) name2444 (
		\DataWidth_reg[1]/NET0131 ,
		_w2220_,
		_w2876_,
		_w2896_,
		_w2897_
	);
	LUT4 #(
		.INIT('h5553)
	) name2445 (
		\Datai[3]_pad ,
		\InstQueue_reg[10][3]/NET0131 ,
		_w2224_,
		_w2225_,
		_w2898_
	);
	LUT2 #(
		.INIT('h1)
	) name2446 (
		_w2229_,
		_w2898_,
		_w2899_
	);
	LUT4 #(
		.INIT('hc055)
	) name2447 (
		\InstQueue_reg[10][3]/NET0131 ,
		_w520_,
		_w525_,
		_w2224_,
		_w2900_
	);
	LUT2 #(
		.INIT('h2)
	) name2448 (
		\InstQueue_reg[10][3]/NET0131 ,
		_w2215_,
		_w2901_
	);
	LUT3 #(
		.INIT('h0d)
	) name2449 (
		_w706_,
		_w2898_,
		_w2901_,
		_w2902_
	);
	LUT3 #(
		.INIT('hd0)
	) name2450 (
		_w722_,
		_w2900_,
		_w2902_,
		_w2903_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name2451 (
		_w700_,
		_w2897_,
		_w2899_,
		_w2903_,
		_w2904_
	);
	LUT4 #(
		.INIT('h6c00)
	) name2452 (
		\Datai[21]_pad ,
		\Datai[22]_pad ,
		_w2200_,
		_w2222_,
		_w2905_
	);
	LUT4 #(
		.INIT('haa80)
	) name2453 (
		\DataWidth_reg[1]/NET0131 ,
		_w2220_,
		_w2886_,
		_w2905_,
		_w2906_
	);
	LUT4 #(
		.INIT('h5553)
	) name2454 (
		\Datai[6]_pad ,
		\InstQueue_reg[10][6]/NET0131 ,
		_w2224_,
		_w2225_,
		_w2907_
	);
	LUT2 #(
		.INIT('h1)
	) name2455 (
		_w2229_,
		_w2907_,
		_w2908_
	);
	LUT4 #(
		.INIT('hc055)
	) name2456 (
		\InstQueue_reg[10][6]/NET0131 ,
		_w485_,
		_w490_,
		_w2224_,
		_w2909_
	);
	LUT2 #(
		.INIT('h2)
	) name2457 (
		\InstQueue_reg[10][6]/NET0131 ,
		_w2215_,
		_w2910_
	);
	LUT3 #(
		.INIT('h0d)
	) name2458 (
		_w706_,
		_w2907_,
		_w2910_,
		_w2911_
	);
	LUT3 #(
		.INIT('hd0)
	) name2459 (
		_w722_,
		_w2909_,
		_w2911_,
		_w2912_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name2460 (
		_w700_,
		_w2906_,
		_w2908_,
		_w2912_,
		_w2913_
	);
	LUT4 #(
		.INIT('h6c00)
	) name2461 (
		\Datai[18]_pad ,
		\Datai[19]_pad ,
		_w2199_,
		_w2225_,
		_w2914_
	);
	LUT4 #(
		.INIT('haa80)
	) name2462 (
		\DataWidth_reg[1]/NET0131 ,
		_w2222_,
		_w2876_,
		_w2914_,
		_w2915_
	);
	LUT4 #(
		.INIT('h5553)
	) name2463 (
		\Datai[3]_pad ,
		\InstQueue_reg[11][3]/NET0131 ,
		_w2224_,
		_w2239_,
		_w2916_
	);
	LUT2 #(
		.INIT('h1)
	) name2464 (
		_w2243_,
		_w2916_,
		_w2917_
	);
	LUT4 #(
		.INIT('hc055)
	) name2465 (
		\InstQueue_reg[11][3]/NET0131 ,
		_w520_,
		_w525_,
		_w2239_,
		_w2918_
	);
	LUT2 #(
		.INIT('h2)
	) name2466 (
		\InstQueue_reg[11][3]/NET0131 ,
		_w2215_,
		_w2919_
	);
	LUT3 #(
		.INIT('h0d)
	) name2467 (
		_w706_,
		_w2916_,
		_w2919_,
		_w2920_
	);
	LUT3 #(
		.INIT('hd0)
	) name2468 (
		_w722_,
		_w2918_,
		_w2920_,
		_w2921_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name2469 (
		_w700_,
		_w2915_,
		_w2917_,
		_w2921_,
		_w2922_
	);
	LUT4 #(
		.INIT('h6c00)
	) name2470 (
		\Datai[21]_pad ,
		\Datai[22]_pad ,
		_w2200_,
		_w2225_,
		_w2923_
	);
	LUT4 #(
		.INIT('haa80)
	) name2471 (
		\DataWidth_reg[1]/NET0131 ,
		_w2222_,
		_w2886_,
		_w2923_,
		_w2924_
	);
	LUT4 #(
		.INIT('h5553)
	) name2472 (
		\Datai[6]_pad ,
		\InstQueue_reg[11][6]/NET0131 ,
		_w2224_,
		_w2239_,
		_w2925_
	);
	LUT2 #(
		.INIT('h1)
	) name2473 (
		_w2243_,
		_w2925_,
		_w2926_
	);
	LUT4 #(
		.INIT('hc055)
	) name2474 (
		\InstQueue_reg[11][6]/NET0131 ,
		_w485_,
		_w490_,
		_w2239_,
		_w2927_
	);
	LUT2 #(
		.INIT('h2)
	) name2475 (
		\InstQueue_reg[11][6]/NET0131 ,
		_w2215_,
		_w2928_
	);
	LUT3 #(
		.INIT('h0d)
	) name2476 (
		_w706_,
		_w2925_,
		_w2928_,
		_w2929_
	);
	LUT3 #(
		.INIT('hd0)
	) name2477 (
		_w722_,
		_w2927_,
		_w2929_,
		_w2930_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name2478 (
		_w700_,
		_w2924_,
		_w2926_,
		_w2930_,
		_w2931_
	);
	LUT4 #(
		.INIT('h6c00)
	) name2479 (
		\Datai[18]_pad ,
		\Datai[19]_pad ,
		_w2199_,
		_w2224_,
		_w2932_
	);
	LUT4 #(
		.INIT('haa80)
	) name2480 (
		\DataWidth_reg[1]/NET0131 ,
		_w2225_,
		_w2876_,
		_w2932_,
		_w2933_
	);
	LUT4 #(
		.INIT('h5553)
	) name2481 (
		\Datai[3]_pad ,
		\InstQueue_reg[12][3]/NET0131 ,
		_w2239_,
		_w2253_,
		_w2934_
	);
	LUT2 #(
		.INIT('h1)
	) name2482 (
		_w2256_,
		_w2934_,
		_w2935_
	);
	LUT4 #(
		.INIT('hc055)
	) name2483 (
		\InstQueue_reg[12][3]/NET0131 ,
		_w520_,
		_w525_,
		_w2253_,
		_w2936_
	);
	LUT2 #(
		.INIT('h2)
	) name2484 (
		\InstQueue_reg[12][3]/NET0131 ,
		_w2215_,
		_w2937_
	);
	LUT3 #(
		.INIT('h0d)
	) name2485 (
		_w706_,
		_w2934_,
		_w2937_,
		_w2938_
	);
	LUT3 #(
		.INIT('hd0)
	) name2486 (
		_w722_,
		_w2936_,
		_w2938_,
		_w2939_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name2487 (
		_w700_,
		_w2933_,
		_w2935_,
		_w2939_,
		_w2940_
	);
	LUT4 #(
		.INIT('h6c00)
	) name2488 (
		\Datai[21]_pad ,
		\Datai[22]_pad ,
		_w2200_,
		_w2224_,
		_w2941_
	);
	LUT4 #(
		.INIT('haa80)
	) name2489 (
		\DataWidth_reg[1]/NET0131 ,
		_w2225_,
		_w2886_,
		_w2941_,
		_w2942_
	);
	LUT4 #(
		.INIT('h5553)
	) name2490 (
		\Datai[6]_pad ,
		\InstQueue_reg[12][6]/NET0131 ,
		_w2239_,
		_w2253_,
		_w2943_
	);
	LUT2 #(
		.INIT('h1)
	) name2491 (
		_w2256_,
		_w2943_,
		_w2944_
	);
	LUT4 #(
		.INIT('hc055)
	) name2492 (
		\InstQueue_reg[12][6]/NET0131 ,
		_w485_,
		_w490_,
		_w2253_,
		_w2945_
	);
	LUT2 #(
		.INIT('h2)
	) name2493 (
		\InstQueue_reg[12][6]/NET0131 ,
		_w2215_,
		_w2946_
	);
	LUT3 #(
		.INIT('h0d)
	) name2494 (
		_w706_,
		_w2943_,
		_w2946_,
		_w2947_
	);
	LUT3 #(
		.INIT('hd0)
	) name2495 (
		_w722_,
		_w2945_,
		_w2947_,
		_w2948_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name2496 (
		_w700_,
		_w2942_,
		_w2944_,
		_w2948_,
		_w2949_
	);
	LUT4 #(
		.INIT('h6c00)
	) name2497 (
		\Datai[18]_pad ,
		\Datai[19]_pad ,
		_w2199_,
		_w2239_,
		_w2950_
	);
	LUT4 #(
		.INIT('haa80)
	) name2498 (
		\DataWidth_reg[1]/NET0131 ,
		_w2224_,
		_w2876_,
		_w2950_,
		_w2951_
	);
	LUT4 #(
		.INIT('h5553)
	) name2499 (
		\Datai[3]_pad ,
		\InstQueue_reg[13][3]/NET0131 ,
		_w2187_,
		_w2253_,
		_w2952_
	);
	LUT2 #(
		.INIT('h1)
	) name2500 (
		_w2268_,
		_w2952_,
		_w2953_
	);
	LUT4 #(
		.INIT('hc055)
	) name2501 (
		\InstQueue_reg[13][3]/NET0131 ,
		_w520_,
		_w525_,
		_w2187_,
		_w2954_
	);
	LUT2 #(
		.INIT('h2)
	) name2502 (
		\InstQueue_reg[13][3]/NET0131 ,
		_w2215_,
		_w2955_
	);
	LUT3 #(
		.INIT('h0d)
	) name2503 (
		_w706_,
		_w2952_,
		_w2955_,
		_w2956_
	);
	LUT3 #(
		.INIT('hd0)
	) name2504 (
		_w722_,
		_w2954_,
		_w2956_,
		_w2957_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name2505 (
		_w700_,
		_w2951_,
		_w2953_,
		_w2957_,
		_w2958_
	);
	LUT4 #(
		.INIT('h6c00)
	) name2506 (
		\Datai[21]_pad ,
		\Datai[22]_pad ,
		_w2200_,
		_w2239_,
		_w2959_
	);
	LUT4 #(
		.INIT('haa80)
	) name2507 (
		\DataWidth_reg[1]/NET0131 ,
		_w2224_,
		_w2886_,
		_w2959_,
		_w2960_
	);
	LUT4 #(
		.INIT('h5553)
	) name2508 (
		\Datai[6]_pad ,
		\InstQueue_reg[13][6]/NET0131 ,
		_w2187_,
		_w2253_,
		_w2961_
	);
	LUT2 #(
		.INIT('h1)
	) name2509 (
		_w2268_,
		_w2961_,
		_w2962_
	);
	LUT4 #(
		.INIT('hc055)
	) name2510 (
		\InstQueue_reg[13][6]/NET0131 ,
		_w485_,
		_w490_,
		_w2187_,
		_w2963_
	);
	LUT2 #(
		.INIT('h2)
	) name2511 (
		\InstQueue_reg[13][6]/NET0131 ,
		_w2215_,
		_w2964_
	);
	LUT3 #(
		.INIT('h0d)
	) name2512 (
		_w706_,
		_w2961_,
		_w2964_,
		_w2965_
	);
	LUT3 #(
		.INIT('hd0)
	) name2513 (
		_w722_,
		_w2963_,
		_w2965_,
		_w2966_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name2514 (
		_w700_,
		_w2960_,
		_w2962_,
		_w2966_,
		_w2967_
	);
	LUT4 #(
		.INIT('h6c00)
	) name2515 (
		\Datai[18]_pad ,
		\Datai[19]_pad ,
		_w2199_,
		_w2253_,
		_w2968_
	);
	LUT4 #(
		.INIT('haa80)
	) name2516 (
		\DataWidth_reg[1]/NET0131 ,
		_w2239_,
		_w2876_,
		_w2968_,
		_w2969_
	);
	LUT4 #(
		.INIT('h5553)
	) name2517 (
		\Datai[3]_pad ,
		\InstQueue_reg[14][3]/NET0131 ,
		_w2187_,
		_w2203_,
		_w2970_
	);
	LUT2 #(
		.INIT('h1)
	) name2518 (
		_w2279_,
		_w2970_,
		_w2971_
	);
	LUT4 #(
		.INIT('hc055)
	) name2519 (
		\InstQueue_reg[14][3]/NET0131 ,
		_w520_,
		_w525_,
		_w2203_,
		_w2972_
	);
	LUT2 #(
		.INIT('h2)
	) name2520 (
		\InstQueue_reg[14][3]/NET0131 ,
		_w2215_,
		_w2973_
	);
	LUT3 #(
		.INIT('h0d)
	) name2521 (
		_w706_,
		_w2970_,
		_w2973_,
		_w2974_
	);
	LUT3 #(
		.INIT('hd0)
	) name2522 (
		_w722_,
		_w2972_,
		_w2974_,
		_w2975_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name2523 (
		_w700_,
		_w2969_,
		_w2971_,
		_w2975_,
		_w2976_
	);
	LUT4 #(
		.INIT('h6c00)
	) name2524 (
		\Datai[21]_pad ,
		\Datai[22]_pad ,
		_w2200_,
		_w2253_,
		_w2977_
	);
	LUT4 #(
		.INIT('haa80)
	) name2525 (
		\DataWidth_reg[1]/NET0131 ,
		_w2239_,
		_w2886_,
		_w2977_,
		_w2978_
	);
	LUT4 #(
		.INIT('h5553)
	) name2526 (
		\Datai[6]_pad ,
		\InstQueue_reg[14][6]/NET0131 ,
		_w2187_,
		_w2203_,
		_w2979_
	);
	LUT2 #(
		.INIT('h1)
	) name2527 (
		_w2279_,
		_w2979_,
		_w2980_
	);
	LUT4 #(
		.INIT('hc055)
	) name2528 (
		\InstQueue_reg[14][6]/NET0131 ,
		_w485_,
		_w490_,
		_w2203_,
		_w2981_
	);
	LUT2 #(
		.INIT('h2)
	) name2529 (
		\InstQueue_reg[14][6]/NET0131 ,
		_w2215_,
		_w2982_
	);
	LUT3 #(
		.INIT('h0d)
	) name2530 (
		_w706_,
		_w2979_,
		_w2982_,
		_w2983_
	);
	LUT3 #(
		.INIT('hd0)
	) name2531 (
		_w722_,
		_w2981_,
		_w2983_,
		_w2984_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name2532 (
		_w700_,
		_w2978_,
		_w2980_,
		_w2984_,
		_w2985_
	);
	LUT4 #(
		.INIT('h60c0)
	) name2533 (
		\Datai[18]_pad ,
		\Datai[19]_pad ,
		_w2187_,
		_w2199_,
		_w2986_
	);
	LUT4 #(
		.INIT('haa80)
	) name2534 (
		\DataWidth_reg[1]/NET0131 ,
		_w2253_,
		_w2876_,
		_w2986_,
		_w2987_
	);
	LUT4 #(
		.INIT('h5553)
	) name2535 (
		\Datai[3]_pad ,
		\InstQueue_reg[15][3]/NET0131 ,
		_w2207_,
		_w2203_,
		_w2988_
	);
	LUT2 #(
		.INIT('h1)
	) name2536 (
		_w2291_,
		_w2988_,
		_w2989_
	);
	LUT4 #(
		.INIT('hc055)
	) name2537 (
		\InstQueue_reg[15][3]/NET0131 ,
		_w520_,
		_w525_,
		_w2207_,
		_w2990_
	);
	LUT2 #(
		.INIT('h2)
	) name2538 (
		\InstQueue_reg[15][3]/NET0131 ,
		_w2215_,
		_w2991_
	);
	LUT3 #(
		.INIT('h0d)
	) name2539 (
		_w706_,
		_w2988_,
		_w2991_,
		_w2992_
	);
	LUT3 #(
		.INIT('hd0)
	) name2540 (
		_w722_,
		_w2990_,
		_w2992_,
		_w2993_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name2541 (
		_w700_,
		_w2987_,
		_w2989_,
		_w2993_,
		_w2994_
	);
	LUT4 #(
		.INIT('h60c0)
	) name2542 (
		\Datai[21]_pad ,
		\Datai[22]_pad ,
		_w2187_,
		_w2200_,
		_w2995_
	);
	LUT4 #(
		.INIT('haa80)
	) name2543 (
		\DataWidth_reg[1]/NET0131 ,
		_w2253_,
		_w2886_,
		_w2995_,
		_w2996_
	);
	LUT4 #(
		.INIT('h5553)
	) name2544 (
		\Datai[6]_pad ,
		\InstQueue_reg[15][6]/NET0131 ,
		_w2207_,
		_w2203_,
		_w2997_
	);
	LUT2 #(
		.INIT('h1)
	) name2545 (
		_w2291_,
		_w2997_,
		_w2998_
	);
	LUT4 #(
		.INIT('hc055)
	) name2546 (
		\InstQueue_reg[15][6]/NET0131 ,
		_w485_,
		_w490_,
		_w2207_,
		_w2999_
	);
	LUT2 #(
		.INIT('h2)
	) name2547 (
		\InstQueue_reg[15][6]/NET0131 ,
		_w2215_,
		_w3000_
	);
	LUT3 #(
		.INIT('h0d)
	) name2548 (
		_w706_,
		_w2997_,
		_w3000_,
		_w3001_
	);
	LUT3 #(
		.INIT('hd0)
	) name2549 (
		_w722_,
		_w2999_,
		_w3001_,
		_w3002_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name2550 (
		_w700_,
		_w2996_,
		_w2998_,
		_w3002_,
		_w3003_
	);
	LUT4 #(
		.INIT('h60c0)
	) name2551 (
		\Datai[18]_pad ,
		\Datai[19]_pad ,
		_w2207_,
		_w2199_,
		_w3004_
	);
	LUT4 #(
		.INIT('haa80)
	) name2552 (
		\DataWidth_reg[1]/NET0131 ,
		_w2203_,
		_w2876_,
		_w3004_,
		_w3005_
	);
	LUT4 #(
		.INIT('h5553)
	) name2553 (
		\Datai[3]_pad ,
		\InstQueue_reg[1][3]/NET0131 ,
		_w2205_,
		_w2301_,
		_w3006_
	);
	LUT2 #(
		.INIT('h1)
	) name2554 (
		_w2304_,
		_w3006_,
		_w3007_
	);
	LUT4 #(
		.INIT('hc055)
	) name2555 (
		\InstQueue_reg[1][3]/NET0131 ,
		_w520_,
		_w525_,
		_w2301_,
		_w3008_
	);
	LUT2 #(
		.INIT('h2)
	) name2556 (
		\InstQueue_reg[1][3]/NET0131 ,
		_w2215_,
		_w3009_
	);
	LUT3 #(
		.INIT('h0d)
	) name2557 (
		_w706_,
		_w3006_,
		_w3009_,
		_w3010_
	);
	LUT3 #(
		.INIT('hd0)
	) name2558 (
		_w722_,
		_w3008_,
		_w3010_,
		_w3011_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name2559 (
		_w700_,
		_w3005_,
		_w3007_,
		_w3011_,
		_w3012_
	);
	LUT4 #(
		.INIT('h60c0)
	) name2560 (
		\Datai[21]_pad ,
		\Datai[22]_pad ,
		_w2207_,
		_w2200_,
		_w3013_
	);
	LUT4 #(
		.INIT('haa80)
	) name2561 (
		\DataWidth_reg[1]/NET0131 ,
		_w2203_,
		_w2886_,
		_w3013_,
		_w3014_
	);
	LUT4 #(
		.INIT('h5553)
	) name2562 (
		\Datai[6]_pad ,
		\InstQueue_reg[1][6]/NET0131 ,
		_w2205_,
		_w2301_,
		_w3015_
	);
	LUT2 #(
		.INIT('h1)
	) name2563 (
		_w2304_,
		_w3015_,
		_w3016_
	);
	LUT4 #(
		.INIT('hc055)
	) name2564 (
		\InstQueue_reg[1][6]/NET0131 ,
		_w485_,
		_w490_,
		_w2301_,
		_w3017_
	);
	LUT2 #(
		.INIT('h2)
	) name2565 (
		\InstQueue_reg[1][6]/NET0131 ,
		_w2215_,
		_w3018_
	);
	LUT3 #(
		.INIT('h0d)
	) name2566 (
		_w706_,
		_w3015_,
		_w3018_,
		_w3019_
	);
	LUT3 #(
		.INIT('hd0)
	) name2567 (
		_w722_,
		_w3017_,
		_w3019_,
		_w3020_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name2568 (
		_w700_,
		_w3014_,
		_w3016_,
		_w3020_,
		_w3021_
	);
	LUT4 #(
		.INIT('h60c0)
	) name2569 (
		\Datai[18]_pad ,
		\Datai[19]_pad ,
		_w2205_,
		_w2199_,
		_w3022_
	);
	LUT4 #(
		.INIT('haa80)
	) name2570 (
		\DataWidth_reg[1]/NET0131 ,
		_w2207_,
		_w2876_,
		_w3022_,
		_w3023_
	);
	LUT4 #(
		.INIT('h5553)
	) name2571 (
		\Datai[3]_pad ,
		\InstQueue_reg[2][3]/NET0131 ,
		_w2301_,
		_w2314_,
		_w3024_
	);
	LUT2 #(
		.INIT('h1)
	) name2572 (
		_w2317_,
		_w3024_,
		_w3025_
	);
	LUT4 #(
		.INIT('hc055)
	) name2573 (
		\InstQueue_reg[2][3]/NET0131 ,
		_w520_,
		_w525_,
		_w2314_,
		_w3026_
	);
	LUT2 #(
		.INIT('h2)
	) name2574 (
		\InstQueue_reg[2][3]/NET0131 ,
		_w2215_,
		_w3027_
	);
	LUT3 #(
		.INIT('h0d)
	) name2575 (
		_w706_,
		_w3024_,
		_w3027_,
		_w3028_
	);
	LUT3 #(
		.INIT('hd0)
	) name2576 (
		_w722_,
		_w3026_,
		_w3028_,
		_w3029_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name2577 (
		_w700_,
		_w3023_,
		_w3025_,
		_w3029_,
		_w3030_
	);
	LUT4 #(
		.INIT('h60c0)
	) name2578 (
		\Datai[21]_pad ,
		\Datai[22]_pad ,
		_w2205_,
		_w2200_,
		_w3031_
	);
	LUT4 #(
		.INIT('haa80)
	) name2579 (
		\DataWidth_reg[1]/NET0131 ,
		_w2207_,
		_w2886_,
		_w3031_,
		_w3032_
	);
	LUT4 #(
		.INIT('h5553)
	) name2580 (
		\Datai[6]_pad ,
		\InstQueue_reg[2][6]/NET0131 ,
		_w2301_,
		_w2314_,
		_w3033_
	);
	LUT2 #(
		.INIT('h1)
	) name2581 (
		_w2317_,
		_w3033_,
		_w3034_
	);
	LUT4 #(
		.INIT('hc055)
	) name2582 (
		\InstQueue_reg[2][6]/NET0131 ,
		_w485_,
		_w490_,
		_w2314_,
		_w3035_
	);
	LUT2 #(
		.INIT('h2)
	) name2583 (
		\InstQueue_reg[2][6]/NET0131 ,
		_w2215_,
		_w3036_
	);
	LUT3 #(
		.INIT('h0d)
	) name2584 (
		_w706_,
		_w3033_,
		_w3036_,
		_w3037_
	);
	LUT3 #(
		.INIT('hd0)
	) name2585 (
		_w722_,
		_w3035_,
		_w3037_,
		_w3038_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name2586 (
		_w700_,
		_w3032_,
		_w3034_,
		_w3038_,
		_w3039_
	);
	LUT4 #(
		.INIT('h6c00)
	) name2587 (
		\Datai[18]_pad ,
		\Datai[19]_pad ,
		_w2199_,
		_w2301_,
		_w3040_
	);
	LUT4 #(
		.INIT('haa80)
	) name2588 (
		\DataWidth_reg[1]/NET0131 ,
		_w2205_,
		_w2876_,
		_w3040_,
		_w3041_
	);
	LUT4 #(
		.INIT('h5553)
	) name2589 (
		\Datai[3]_pad ,
		\InstQueue_reg[3][3]/NET0131 ,
		_w2314_,
		_w2327_,
		_w3042_
	);
	LUT2 #(
		.INIT('h1)
	) name2590 (
		_w2330_,
		_w3042_,
		_w3043_
	);
	LUT4 #(
		.INIT('hc055)
	) name2591 (
		\InstQueue_reg[3][3]/NET0131 ,
		_w520_,
		_w525_,
		_w2327_,
		_w3044_
	);
	LUT2 #(
		.INIT('h2)
	) name2592 (
		\InstQueue_reg[3][3]/NET0131 ,
		_w2215_,
		_w3045_
	);
	LUT3 #(
		.INIT('h0d)
	) name2593 (
		_w706_,
		_w3042_,
		_w3045_,
		_w3046_
	);
	LUT3 #(
		.INIT('hd0)
	) name2594 (
		_w722_,
		_w3044_,
		_w3046_,
		_w3047_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name2595 (
		_w700_,
		_w3041_,
		_w3043_,
		_w3047_,
		_w3048_
	);
	LUT4 #(
		.INIT('h6c00)
	) name2596 (
		\Datai[21]_pad ,
		\Datai[22]_pad ,
		_w2200_,
		_w2301_,
		_w3049_
	);
	LUT4 #(
		.INIT('haa80)
	) name2597 (
		\DataWidth_reg[1]/NET0131 ,
		_w2205_,
		_w2886_,
		_w3049_,
		_w3050_
	);
	LUT4 #(
		.INIT('h5553)
	) name2598 (
		\Datai[6]_pad ,
		\InstQueue_reg[3][6]/NET0131 ,
		_w2314_,
		_w2327_,
		_w3051_
	);
	LUT2 #(
		.INIT('h1)
	) name2599 (
		_w2330_,
		_w3051_,
		_w3052_
	);
	LUT4 #(
		.INIT('hc055)
	) name2600 (
		\InstQueue_reg[3][6]/NET0131 ,
		_w485_,
		_w490_,
		_w2327_,
		_w3053_
	);
	LUT2 #(
		.INIT('h2)
	) name2601 (
		\InstQueue_reg[3][6]/NET0131 ,
		_w2215_,
		_w3054_
	);
	LUT3 #(
		.INIT('h0d)
	) name2602 (
		_w706_,
		_w3051_,
		_w3054_,
		_w3055_
	);
	LUT3 #(
		.INIT('hd0)
	) name2603 (
		_w722_,
		_w3053_,
		_w3055_,
		_w3056_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name2604 (
		_w700_,
		_w3050_,
		_w3052_,
		_w3056_,
		_w3057_
	);
	LUT4 #(
		.INIT('h6c00)
	) name2605 (
		\Datai[18]_pad ,
		\Datai[19]_pad ,
		_w2199_,
		_w2314_,
		_w3058_
	);
	LUT4 #(
		.INIT('haa80)
	) name2606 (
		\DataWidth_reg[1]/NET0131 ,
		_w2301_,
		_w2876_,
		_w3058_,
		_w3059_
	);
	LUT4 #(
		.INIT('h5553)
	) name2607 (
		\Datai[3]_pad ,
		\InstQueue_reg[4][3]/NET0131 ,
		_w2327_,
		_w2340_,
		_w3060_
	);
	LUT2 #(
		.INIT('h1)
	) name2608 (
		_w2343_,
		_w3060_,
		_w3061_
	);
	LUT4 #(
		.INIT('hc055)
	) name2609 (
		\InstQueue_reg[4][3]/NET0131 ,
		_w520_,
		_w525_,
		_w2340_,
		_w3062_
	);
	LUT2 #(
		.INIT('h2)
	) name2610 (
		\InstQueue_reg[4][3]/NET0131 ,
		_w2215_,
		_w3063_
	);
	LUT3 #(
		.INIT('h0d)
	) name2611 (
		_w706_,
		_w3060_,
		_w3063_,
		_w3064_
	);
	LUT3 #(
		.INIT('hd0)
	) name2612 (
		_w722_,
		_w3062_,
		_w3064_,
		_w3065_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name2613 (
		_w700_,
		_w3059_,
		_w3061_,
		_w3065_,
		_w3066_
	);
	LUT4 #(
		.INIT('h6c00)
	) name2614 (
		\Datai[21]_pad ,
		\Datai[22]_pad ,
		_w2200_,
		_w2314_,
		_w3067_
	);
	LUT4 #(
		.INIT('haa80)
	) name2615 (
		\DataWidth_reg[1]/NET0131 ,
		_w2301_,
		_w2886_,
		_w3067_,
		_w3068_
	);
	LUT4 #(
		.INIT('h5553)
	) name2616 (
		\Datai[6]_pad ,
		\InstQueue_reg[4][6]/NET0131 ,
		_w2327_,
		_w2340_,
		_w3069_
	);
	LUT2 #(
		.INIT('h1)
	) name2617 (
		_w2343_,
		_w3069_,
		_w3070_
	);
	LUT4 #(
		.INIT('hc055)
	) name2618 (
		\InstQueue_reg[4][6]/NET0131 ,
		_w485_,
		_w490_,
		_w2340_,
		_w3071_
	);
	LUT2 #(
		.INIT('h2)
	) name2619 (
		\InstQueue_reg[4][6]/NET0131 ,
		_w2215_,
		_w3072_
	);
	LUT3 #(
		.INIT('h0d)
	) name2620 (
		_w706_,
		_w3069_,
		_w3072_,
		_w3073_
	);
	LUT3 #(
		.INIT('hd0)
	) name2621 (
		_w722_,
		_w3071_,
		_w3073_,
		_w3074_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name2622 (
		_w700_,
		_w3068_,
		_w3070_,
		_w3074_,
		_w3075_
	);
	LUT4 #(
		.INIT('h6c00)
	) name2623 (
		\Datai[18]_pad ,
		\Datai[19]_pad ,
		_w2199_,
		_w2327_,
		_w3076_
	);
	LUT4 #(
		.INIT('haa80)
	) name2624 (
		\DataWidth_reg[1]/NET0131 ,
		_w2314_,
		_w2876_,
		_w3076_,
		_w3077_
	);
	LUT4 #(
		.INIT('h5553)
	) name2625 (
		\Datai[3]_pad ,
		\InstQueue_reg[5][3]/NET0131 ,
		_w2340_,
		_w2353_,
		_w3078_
	);
	LUT2 #(
		.INIT('h1)
	) name2626 (
		_w2356_,
		_w3078_,
		_w3079_
	);
	LUT4 #(
		.INIT('hc055)
	) name2627 (
		\InstQueue_reg[5][3]/NET0131 ,
		_w520_,
		_w525_,
		_w2353_,
		_w3080_
	);
	LUT2 #(
		.INIT('h2)
	) name2628 (
		\InstQueue_reg[5][3]/NET0131 ,
		_w2215_,
		_w3081_
	);
	LUT3 #(
		.INIT('h0d)
	) name2629 (
		_w706_,
		_w3078_,
		_w3081_,
		_w3082_
	);
	LUT3 #(
		.INIT('hd0)
	) name2630 (
		_w722_,
		_w3080_,
		_w3082_,
		_w3083_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name2631 (
		_w700_,
		_w3077_,
		_w3079_,
		_w3083_,
		_w3084_
	);
	LUT4 #(
		.INIT('h6c00)
	) name2632 (
		\Datai[21]_pad ,
		\Datai[22]_pad ,
		_w2200_,
		_w2327_,
		_w3085_
	);
	LUT4 #(
		.INIT('haa80)
	) name2633 (
		\DataWidth_reg[1]/NET0131 ,
		_w2314_,
		_w2886_,
		_w3085_,
		_w3086_
	);
	LUT4 #(
		.INIT('h5553)
	) name2634 (
		\Datai[6]_pad ,
		\InstQueue_reg[5][6]/NET0131 ,
		_w2340_,
		_w2353_,
		_w3087_
	);
	LUT2 #(
		.INIT('h1)
	) name2635 (
		_w2356_,
		_w3087_,
		_w3088_
	);
	LUT4 #(
		.INIT('hc055)
	) name2636 (
		\InstQueue_reg[5][6]/NET0131 ,
		_w485_,
		_w490_,
		_w2353_,
		_w3089_
	);
	LUT2 #(
		.INIT('h2)
	) name2637 (
		\InstQueue_reg[5][6]/NET0131 ,
		_w2215_,
		_w3090_
	);
	LUT3 #(
		.INIT('h0d)
	) name2638 (
		_w706_,
		_w3087_,
		_w3090_,
		_w3091_
	);
	LUT3 #(
		.INIT('hd0)
	) name2639 (
		_w722_,
		_w3089_,
		_w3091_,
		_w3092_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name2640 (
		_w700_,
		_w3086_,
		_w3088_,
		_w3092_,
		_w3093_
	);
	LUT4 #(
		.INIT('h6c00)
	) name2641 (
		\Datai[18]_pad ,
		\Datai[19]_pad ,
		_w2199_,
		_w2340_,
		_w3094_
	);
	LUT4 #(
		.INIT('haa80)
	) name2642 (
		\DataWidth_reg[1]/NET0131 ,
		_w2327_,
		_w2876_,
		_w3094_,
		_w3095_
	);
	LUT4 #(
		.INIT('h5553)
	) name2643 (
		\Datai[3]_pad ,
		\InstQueue_reg[6][3]/NET0131 ,
		_w2353_,
		_w2366_,
		_w3096_
	);
	LUT2 #(
		.INIT('h1)
	) name2644 (
		_w2369_,
		_w3096_,
		_w3097_
	);
	LUT4 #(
		.INIT('hc055)
	) name2645 (
		\InstQueue_reg[6][3]/NET0131 ,
		_w520_,
		_w525_,
		_w2366_,
		_w3098_
	);
	LUT2 #(
		.INIT('h2)
	) name2646 (
		\InstQueue_reg[6][3]/NET0131 ,
		_w2215_,
		_w3099_
	);
	LUT3 #(
		.INIT('h0d)
	) name2647 (
		_w706_,
		_w3096_,
		_w3099_,
		_w3100_
	);
	LUT3 #(
		.INIT('hd0)
	) name2648 (
		_w722_,
		_w3098_,
		_w3100_,
		_w3101_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name2649 (
		_w700_,
		_w3095_,
		_w3097_,
		_w3101_,
		_w3102_
	);
	LUT4 #(
		.INIT('h6c00)
	) name2650 (
		\Datai[21]_pad ,
		\Datai[22]_pad ,
		_w2200_,
		_w2340_,
		_w3103_
	);
	LUT4 #(
		.INIT('haa80)
	) name2651 (
		\DataWidth_reg[1]/NET0131 ,
		_w2327_,
		_w2886_,
		_w3103_,
		_w3104_
	);
	LUT4 #(
		.INIT('h5553)
	) name2652 (
		\Datai[6]_pad ,
		\InstQueue_reg[6][6]/NET0131 ,
		_w2353_,
		_w2366_,
		_w3105_
	);
	LUT2 #(
		.INIT('h1)
	) name2653 (
		_w2369_,
		_w3105_,
		_w3106_
	);
	LUT4 #(
		.INIT('hc055)
	) name2654 (
		\InstQueue_reg[6][6]/NET0131 ,
		_w485_,
		_w490_,
		_w2366_,
		_w3107_
	);
	LUT2 #(
		.INIT('h2)
	) name2655 (
		\InstQueue_reg[6][6]/NET0131 ,
		_w2215_,
		_w3108_
	);
	LUT3 #(
		.INIT('h0d)
	) name2656 (
		_w706_,
		_w3105_,
		_w3108_,
		_w3109_
	);
	LUT3 #(
		.INIT('hd0)
	) name2657 (
		_w722_,
		_w3107_,
		_w3109_,
		_w3110_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name2658 (
		_w700_,
		_w3104_,
		_w3106_,
		_w3110_,
		_w3111_
	);
	LUT4 #(
		.INIT('h6c00)
	) name2659 (
		\Datai[18]_pad ,
		\Datai[19]_pad ,
		_w2199_,
		_w2353_,
		_w3112_
	);
	LUT4 #(
		.INIT('haa80)
	) name2660 (
		\DataWidth_reg[1]/NET0131 ,
		_w2340_,
		_w2876_,
		_w3112_,
		_w3113_
	);
	LUT4 #(
		.INIT('h5553)
	) name2661 (
		\Datai[3]_pad ,
		\InstQueue_reg[7][3]/NET0131 ,
		_w2220_,
		_w2366_,
		_w3114_
	);
	LUT2 #(
		.INIT('h1)
	) name2662 (
		_w2381_,
		_w3114_,
		_w3115_
	);
	LUT4 #(
		.INIT('hc055)
	) name2663 (
		\InstQueue_reg[7][3]/NET0131 ,
		_w520_,
		_w525_,
		_w2220_,
		_w3116_
	);
	LUT2 #(
		.INIT('h2)
	) name2664 (
		\InstQueue_reg[7][3]/NET0131 ,
		_w2215_,
		_w3117_
	);
	LUT3 #(
		.INIT('h0d)
	) name2665 (
		_w706_,
		_w3114_,
		_w3117_,
		_w3118_
	);
	LUT3 #(
		.INIT('hd0)
	) name2666 (
		_w722_,
		_w3116_,
		_w3118_,
		_w3119_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name2667 (
		_w700_,
		_w3113_,
		_w3115_,
		_w3119_,
		_w3120_
	);
	LUT4 #(
		.INIT('h6c00)
	) name2668 (
		\Datai[21]_pad ,
		\Datai[22]_pad ,
		_w2200_,
		_w2353_,
		_w3121_
	);
	LUT4 #(
		.INIT('haa80)
	) name2669 (
		\DataWidth_reg[1]/NET0131 ,
		_w2340_,
		_w2886_,
		_w3121_,
		_w3122_
	);
	LUT4 #(
		.INIT('h5553)
	) name2670 (
		\Datai[6]_pad ,
		\InstQueue_reg[7][6]/NET0131 ,
		_w2220_,
		_w2366_,
		_w3123_
	);
	LUT2 #(
		.INIT('h1)
	) name2671 (
		_w2381_,
		_w3123_,
		_w3124_
	);
	LUT4 #(
		.INIT('hc055)
	) name2672 (
		\InstQueue_reg[7][6]/NET0131 ,
		_w485_,
		_w490_,
		_w2220_,
		_w3125_
	);
	LUT2 #(
		.INIT('h2)
	) name2673 (
		\InstQueue_reg[7][6]/NET0131 ,
		_w2215_,
		_w3126_
	);
	LUT3 #(
		.INIT('h0d)
	) name2674 (
		_w706_,
		_w3123_,
		_w3126_,
		_w3127_
	);
	LUT3 #(
		.INIT('hd0)
	) name2675 (
		_w722_,
		_w3125_,
		_w3127_,
		_w3128_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name2676 (
		_w700_,
		_w3122_,
		_w3124_,
		_w3128_,
		_w3129_
	);
	LUT4 #(
		.INIT('h6c00)
	) name2677 (
		\Datai[18]_pad ,
		\Datai[19]_pad ,
		_w2199_,
		_w2366_,
		_w3130_
	);
	LUT4 #(
		.INIT('haa80)
	) name2678 (
		\DataWidth_reg[1]/NET0131 ,
		_w2353_,
		_w2876_,
		_w3130_,
		_w3131_
	);
	LUT4 #(
		.INIT('h5553)
	) name2679 (
		\Datai[3]_pad ,
		\InstQueue_reg[8][3]/NET0131 ,
		_w2220_,
		_w2222_,
		_w3132_
	);
	LUT2 #(
		.INIT('h1)
	) name2680 (
		_w2392_,
		_w3132_,
		_w3133_
	);
	LUT4 #(
		.INIT('hc055)
	) name2681 (
		\InstQueue_reg[8][3]/NET0131 ,
		_w520_,
		_w525_,
		_w2222_,
		_w3134_
	);
	LUT2 #(
		.INIT('h2)
	) name2682 (
		\InstQueue_reg[8][3]/NET0131 ,
		_w2215_,
		_w3135_
	);
	LUT3 #(
		.INIT('h0d)
	) name2683 (
		_w706_,
		_w3132_,
		_w3135_,
		_w3136_
	);
	LUT3 #(
		.INIT('hd0)
	) name2684 (
		_w722_,
		_w3134_,
		_w3136_,
		_w3137_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name2685 (
		_w700_,
		_w3131_,
		_w3133_,
		_w3137_,
		_w3138_
	);
	LUT4 #(
		.INIT('h6c00)
	) name2686 (
		\Datai[21]_pad ,
		\Datai[22]_pad ,
		_w2200_,
		_w2366_,
		_w3139_
	);
	LUT4 #(
		.INIT('haa80)
	) name2687 (
		\DataWidth_reg[1]/NET0131 ,
		_w2353_,
		_w2886_,
		_w3139_,
		_w3140_
	);
	LUT4 #(
		.INIT('h5553)
	) name2688 (
		\Datai[6]_pad ,
		\InstQueue_reg[8][6]/NET0131 ,
		_w2220_,
		_w2222_,
		_w3141_
	);
	LUT2 #(
		.INIT('h1)
	) name2689 (
		_w2392_,
		_w3141_,
		_w3142_
	);
	LUT4 #(
		.INIT('hc055)
	) name2690 (
		\InstQueue_reg[8][6]/NET0131 ,
		_w485_,
		_w490_,
		_w2222_,
		_w3143_
	);
	LUT2 #(
		.INIT('h2)
	) name2691 (
		\InstQueue_reg[8][6]/NET0131 ,
		_w2215_,
		_w3144_
	);
	LUT3 #(
		.INIT('h0d)
	) name2692 (
		_w706_,
		_w3141_,
		_w3144_,
		_w3145_
	);
	LUT3 #(
		.INIT('hd0)
	) name2693 (
		_w722_,
		_w3143_,
		_w3145_,
		_w3146_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name2694 (
		_w700_,
		_w3140_,
		_w3142_,
		_w3146_,
		_w3147_
	);
	LUT4 #(
		.INIT('h6c00)
	) name2695 (
		\Datai[18]_pad ,
		\Datai[19]_pad ,
		_w2199_,
		_w2220_,
		_w3148_
	);
	LUT4 #(
		.INIT('haa80)
	) name2696 (
		\DataWidth_reg[1]/NET0131 ,
		_w2366_,
		_w2876_,
		_w3148_,
		_w3149_
	);
	LUT4 #(
		.INIT('h5553)
	) name2697 (
		\Datai[3]_pad ,
		\InstQueue_reg[9][3]/NET0131 ,
		_w2225_,
		_w2222_,
		_w3150_
	);
	LUT2 #(
		.INIT('h1)
	) name2698 (
		_w2403_,
		_w3150_,
		_w3151_
	);
	LUT4 #(
		.INIT('hc055)
	) name2699 (
		\InstQueue_reg[9][3]/NET0131 ,
		_w520_,
		_w525_,
		_w2225_,
		_w3152_
	);
	LUT2 #(
		.INIT('h2)
	) name2700 (
		\InstQueue_reg[9][3]/NET0131 ,
		_w2215_,
		_w3153_
	);
	LUT3 #(
		.INIT('h0d)
	) name2701 (
		_w706_,
		_w3150_,
		_w3153_,
		_w3154_
	);
	LUT3 #(
		.INIT('hd0)
	) name2702 (
		_w722_,
		_w3152_,
		_w3154_,
		_w3155_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name2703 (
		_w700_,
		_w3149_,
		_w3151_,
		_w3155_,
		_w3156_
	);
	LUT4 #(
		.INIT('h6c00)
	) name2704 (
		\Datai[21]_pad ,
		\Datai[22]_pad ,
		_w2200_,
		_w2220_,
		_w3157_
	);
	LUT4 #(
		.INIT('haa80)
	) name2705 (
		\DataWidth_reg[1]/NET0131 ,
		_w2366_,
		_w2886_,
		_w3157_,
		_w3158_
	);
	LUT4 #(
		.INIT('h5553)
	) name2706 (
		\Datai[6]_pad ,
		\InstQueue_reg[9][6]/NET0131 ,
		_w2225_,
		_w2222_,
		_w3159_
	);
	LUT2 #(
		.INIT('h1)
	) name2707 (
		_w2403_,
		_w3159_,
		_w3160_
	);
	LUT4 #(
		.INIT('hc055)
	) name2708 (
		\InstQueue_reg[9][6]/NET0131 ,
		_w485_,
		_w490_,
		_w2225_,
		_w3161_
	);
	LUT2 #(
		.INIT('h2)
	) name2709 (
		\InstQueue_reg[9][6]/NET0131 ,
		_w2215_,
		_w3162_
	);
	LUT3 #(
		.INIT('h0d)
	) name2710 (
		_w706_,
		_w3159_,
		_w3162_,
		_w3163_
	);
	LUT3 #(
		.INIT('hd0)
	) name2711 (
		_w722_,
		_w3161_,
		_w3163_,
		_w3164_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name2712 (
		_w700_,
		_w3158_,
		_w3160_,
		_w3164_,
		_w3165_
	);
	LUT4 #(
		.INIT('h08aa)
	) name2713 (
		\PhyAddrPointer_reg[0]/NET0131 ,
		_w695_,
		_w1984_,
		_w1110_,
		_w3166_
	);
	LUT4 #(
		.INIT('h0057)
	) name2714 (
		_w695_,
		_w2018_,
		_w2019_,
		_w2025_,
		_w3167_
	);
	LUT2 #(
		.INIT('hb)
	) name2715 (
		_w3166_,
		_w3167_,
		_w3168_
	);
	LUT4 #(
		.INIT('h1450)
	) name2716 (
		\DataWidth_reg[1]/NET0131 ,
		\PhyAddrPointer_reg[0]/NET0131 ,
		\PhyAddrPointer_reg[1]/NET0131 ,
		_w1279_,
		_w3169_
	);
	LUT2 #(
		.INIT('h2)
	) name2717 (
		\DataWidth_reg[1]/NET0131 ,
		\rEIP_reg[1]/NET0131 ,
		_w3170_
	);
	LUT2 #(
		.INIT('h2)
	) name2718 (
		_w700_,
		_w3170_,
		_w3171_
	);
	LUT2 #(
		.INIT('h2)
	) name2719 (
		\rEIP_reg[1]/NET0131 ,
		_w2640_,
		_w3172_
	);
	LUT3 #(
		.INIT('h23)
	) name2720 (
		\DataWidth_reg[1]/NET0131 ,
		\EBX_reg[1]/NET0131 ,
		_w633_,
		_w3173_
	);
	LUT2 #(
		.INIT('h6)
	) name2721 (
		\EBX_reg[0]/NET0131 ,
		\EBX_reg[1]/NET0131 ,
		_w3174_
	);
	LUT3 #(
		.INIT('h60)
	) name2722 (
		\EBX_reg[0]/NET0131 ,
		\EBX_reg[1]/NET0131 ,
		\EBX_reg[31]/NET0131 ,
		_w3175_
	);
	LUT4 #(
		.INIT('hf3a2)
	) name2723 (
		\DataWidth_reg[1]/NET0131 ,
		\EBX_reg[1]/NET0131 ,
		\EBX_reg[31]/NET0131 ,
		READY_n_pad,
		_w3176_
	);
	LUT2 #(
		.INIT('h4)
	) name2724 (
		_w3175_,
		_w3176_,
		_w3177_
	);
	LUT4 #(
		.INIT('hf351)
	) name2725 (
		_w566_,
		_w570_,
		_w3173_,
		_w3177_,
		_w3178_
	);
	LUT3 #(
		.INIT('h10)
	) name2726 (
		\DataWidth_reg[1]/NET0131 ,
		READY_n_pad,
		\rEIP_reg[1]/NET0131 ,
		_w3179_
	);
	LUT3 #(
		.INIT('h08)
	) name2727 (
		_w570_,
		_w617_,
		_w3173_,
		_w3180_
	);
	LUT2 #(
		.INIT('h2)
	) name2728 (
		_w569_,
		_w607_,
		_w3181_
	);
	LUT4 #(
		.INIT('h1110)
	) name2729 (
		_w3180_,
		_w3181_,
		_w3178_,
		_w3179_,
		_w3182_
	);
	LUT4 #(
		.INIT('hc0c8)
	) name2730 (
		_w611_,
		_w695_,
		_w3172_,
		_w3182_,
		_w3183_
	);
	LUT4 #(
		.INIT('h5f13)
	) name2731 (
		\PhyAddrPointer_reg[1]/NET0131 ,
		\rEIP_reg[1]/NET0131 ,
		_w718_,
		_w2661_,
		_w3184_
	);
	LUT4 #(
		.INIT('hbaff)
	) name2732 (
		_w3183_,
		_w3169_,
		_w3171_,
		_w3184_,
		_w3185_
	);
	LUT4 #(
		.INIT('h4000)
	) name2733 (
		\PhyAddrPointer_reg[0]/NET0131 ,
		\PhyAddrPointer_reg[1]/NET0131 ,
		_w1268_,
		_w1569_,
		_w3186_
	);
	LUT4 #(
		.INIT('h0541)
	) name2734 (
		\DataWidth_reg[1]/NET0131 ,
		_w1279_,
		_w1584_,
		_w3186_,
		_w3187_
	);
	LUT2 #(
		.INIT('h2)
	) name2735 (
		\DataWidth_reg[1]/NET0131 ,
		\rEIP_reg[20]/NET0131 ,
		_w3188_
	);
	LUT2 #(
		.INIT('h2)
	) name2736 (
		_w700_,
		_w3188_,
		_w3189_
	);
	LUT2 #(
		.INIT('h4)
	) name2737 (
		_w3187_,
		_w3189_,
		_w3190_
	);
	LUT2 #(
		.INIT('h2)
	) name2738 (
		\rEIP_reg[20]/NET0131 ,
		_w2640_,
		_w3191_
	);
	LUT3 #(
		.INIT('h23)
	) name2739 (
		\DataWidth_reg[1]/NET0131 ,
		\EBX_reg[20]/NET0131 ,
		_w633_,
		_w3192_
	);
	LUT2 #(
		.INIT('h2)
	) name2740 (
		_w570_,
		_w3192_,
		_w3193_
	);
	LUT4 #(
		.INIT('he0f0)
	) name2741 (
		\EBX_reg[18]/NET0131 ,
		\EBX_reg[19]/NET0131 ,
		\EBX_reg[31]/NET0131 ,
		_w2630_,
		_w3194_
	);
	LUT4 #(
		.INIT('hc4c8)
	) name2742 (
		\EBX_reg[20]/NET0131 ,
		_w566_,
		_w2623_,
		_w3194_,
		_w3195_
	);
	LUT3 #(
		.INIT('h6a)
	) name2743 (
		\rEIP_reg[20]/NET0131 ,
		_w2611_,
		_w2613_,
		_w3196_
	);
	LUT4 #(
		.INIT('hf070)
	) name2744 (
		_w570_,
		_w617_,
		_w2623_,
		_w3192_,
		_w3197_
	);
	LUT3 #(
		.INIT('h8a)
	) name2745 (
		_w611_,
		_w3196_,
		_w3197_,
		_w3198_
	);
	LUT4 #(
		.INIT('h0155)
	) name2746 (
		_w3191_,
		_w3193_,
		_w3195_,
		_w3198_,
		_w3199_
	);
	LUT4 #(
		.INIT('h5f13)
	) name2747 (
		\PhyAddrPointer_reg[20]/NET0131 ,
		\rEIP_reg[20]/NET0131 ,
		_w718_,
		_w2661_,
		_w3200_
	);
	LUT3 #(
		.INIT('hd0)
	) name2748 (
		_w695_,
		_w3199_,
		_w3200_,
		_w3201_
	);
	LUT2 #(
		.INIT('hb)
	) name2749 (
		_w3190_,
		_w3201_,
		_w3202_
	);
	LUT4 #(
		.INIT('h1333)
	) name2750 (
		\PhyAddrPointer_reg[1]/NET0131 ,
		\PhyAddrPointer_reg[21]/NET0131 ,
		_w1269_,
		_w1569_,
		_w3203_
	);
	LUT2 #(
		.INIT('h1)
	) name2751 (
		_w1462_,
		_w3203_,
		_w3204_
	);
	LUT2 #(
		.INIT('h4)
	) name2752 (
		\PhyAddrPointer_reg[0]/NET0131 ,
		\PhyAddrPointer_reg[1]/NET0131 ,
		_w3205_
	);
	LUT4 #(
		.INIT('h4000)
	) name2753 (
		\PhyAddrPointer_reg[0]/NET0131 ,
		\PhyAddrPointer_reg[1]/NET0131 ,
		\PhyAddrPointer_reg[2]/NET0131 ,
		\PhyAddrPointer_reg[3]/NET0131 ,
		_w3206_
	);
	LUT2 #(
		.INIT('h8)
	) name2754 (
		\PhyAddrPointer_reg[4]/NET0131 ,
		_w3206_,
		_w3207_
	);
	LUT2 #(
		.INIT('h8)
	) name2755 (
		_w1261_,
		_w3207_,
		_w3208_
	);
	LUT4 #(
		.INIT('h8000)
	) name2756 (
		\PhyAddrPointer_reg[1]/NET0131 ,
		_w1269_,
		_w1569_,
		_w3208_,
		_w3209_
	);
	LUT4 #(
		.INIT('h0541)
	) name2757 (
		\DataWidth_reg[1]/NET0131 ,
		_w1279_,
		_w3204_,
		_w3209_,
		_w3210_
	);
	LUT2 #(
		.INIT('h2)
	) name2758 (
		\DataWidth_reg[1]/NET0131 ,
		\rEIP_reg[21]/NET0131 ,
		_w3211_
	);
	LUT2 #(
		.INIT('h2)
	) name2759 (
		_w700_,
		_w3211_,
		_w3212_
	);
	LUT2 #(
		.INIT('h4)
	) name2760 (
		_w3210_,
		_w3212_,
		_w3213_
	);
	LUT4 #(
		.INIT('h0100)
	) name2761 (
		\EBX_reg[18]/NET0131 ,
		\EBX_reg[19]/NET0131 ,
		\EBX_reg[20]/NET0131 ,
		_w2630_,
		_w3214_
	);
	LUT4 #(
		.INIT('h0509)
	) name2762 (
		\EBX_reg[21]/NET0131 ,
		\EBX_reg[31]/NET0131 ,
		_w2623_,
		_w3214_,
		_w3215_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name2763 (
		\rEIP_reg[20]/NET0131 ,
		\rEIP_reg[21]/NET0131 ,
		_w2611_,
		_w2613_,
		_w3216_
	);
	LUT3 #(
		.INIT('ha2)
	) name2764 (
		_w1100_,
		_w2623_,
		_w3216_,
		_w3217_
	);
	LUT2 #(
		.INIT('h2)
	) name2765 (
		\rEIP_reg[21]/NET0131 ,
		_w2640_,
		_w3218_
	);
	LUT3 #(
		.INIT('h23)
	) name2766 (
		\DataWidth_reg[1]/NET0131 ,
		\EBX_reg[21]/NET0131 ,
		_w633_,
		_w3219_
	);
	LUT3 #(
		.INIT('h08)
	) name2767 (
		_w570_,
		_w611_,
		_w3219_,
		_w3220_
	);
	LUT4 #(
		.INIT('hfb00)
	) name2768 (
		_w617_,
		_w2623_,
		_w3216_,
		_w3220_,
		_w3221_
	);
	LUT4 #(
		.INIT('h000b)
	) name2769 (
		_w3215_,
		_w3217_,
		_w3218_,
		_w3221_,
		_w3222_
	);
	LUT4 #(
		.INIT('h5f13)
	) name2770 (
		\PhyAddrPointer_reg[21]/NET0131 ,
		\rEIP_reg[21]/NET0131 ,
		_w718_,
		_w2661_,
		_w3223_
	);
	LUT3 #(
		.INIT('hd0)
	) name2771 (
		_w695_,
		_w3222_,
		_w3223_,
		_w3224_
	);
	LUT2 #(
		.INIT('hb)
	) name2772 (
		_w3213_,
		_w3224_,
		_w3225_
	);
	LUT4 #(
		.INIT('h0541)
	) name2773 (
		\DataWidth_reg[1]/NET0131 ,
		_w1279_,
		_w1597_,
		_w2652_,
		_w3226_
	);
	LUT2 #(
		.INIT('h2)
	) name2774 (
		\DataWidth_reg[1]/NET0131 ,
		\rEIP_reg[22]/NET0131 ,
		_w3227_
	);
	LUT2 #(
		.INIT('h2)
	) name2775 (
		_w700_,
		_w3227_,
		_w3228_
	);
	LUT2 #(
		.INIT('h4)
	) name2776 (
		_w3226_,
		_w3228_,
		_w3229_
	);
	LUT3 #(
		.INIT('h8c)
	) name2777 (
		\EBX_reg[21]/NET0131 ,
		\EBX_reg[31]/NET0131 ,
		_w3214_,
		_w3230_
	);
	LUT4 #(
		.INIT('h9500)
	) name2778 (
		\rEIP_reg[22]/NET0131 ,
		_w2611_,
		_w2615_,
		_w2623_,
		_w3231_
	);
	LUT2 #(
		.INIT('h2)
	) name2779 (
		_w1100_,
		_w3231_,
		_w3232_
	);
	LUT4 #(
		.INIT('hde00)
	) name2780 (
		\EBX_reg[22]/NET0131 ,
		_w2623_,
		_w3230_,
		_w3232_,
		_w3233_
	);
	LUT4 #(
		.INIT('h9500)
	) name2781 (
		\rEIP_reg[22]/NET0131 ,
		_w2611_,
		_w2615_,
		_w2642_,
		_w3234_
	);
	LUT3 #(
		.INIT('h23)
	) name2782 (
		\DataWidth_reg[1]/NET0131 ,
		\EBX_reg[22]/NET0131 ,
		_w633_,
		_w3235_
	);
	LUT3 #(
		.INIT('h08)
	) name2783 (
		_w570_,
		_w611_,
		_w3235_,
		_w3236_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name2784 (
		\rEIP_reg[22]/NET0131 ,
		_w2640_,
		_w3234_,
		_w3236_,
		_w3237_
	);
	LUT4 #(
		.INIT('h5f13)
	) name2785 (
		\PhyAddrPointer_reg[22]/NET0131 ,
		\rEIP_reg[22]/NET0131 ,
		_w718_,
		_w2661_,
		_w3238_
	);
	LUT4 #(
		.INIT('h7500)
	) name2786 (
		_w695_,
		_w3233_,
		_w3237_,
		_w3238_,
		_w3239_
	);
	LUT2 #(
		.INIT('hb)
	) name2787 (
		_w3229_,
		_w3239_,
		_w3240_
	);
	LUT4 #(
		.INIT('h0541)
	) name2788 (
		\DataWidth_reg[1]/NET0131 ,
		_w1279_,
		_w1463_,
		_w2653_,
		_w3241_
	);
	LUT2 #(
		.INIT('h2)
	) name2789 (
		\DataWidth_reg[1]/NET0131 ,
		\rEIP_reg[23]/NET0131 ,
		_w3242_
	);
	LUT2 #(
		.INIT('h2)
	) name2790 (
		_w700_,
		_w3242_,
		_w3243_
	);
	LUT2 #(
		.INIT('h4)
	) name2791 (
		_w3241_,
		_w3243_,
		_w3244_
	);
	LUT4 #(
		.INIT('he0f0)
	) name2792 (
		\EBX_reg[21]/NET0131 ,
		\EBX_reg[22]/NET0131 ,
		\EBX_reg[31]/NET0131 ,
		_w3214_,
		_w3245_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name2793 (
		\rEIP_reg[22]/NET0131 ,
		\rEIP_reg[23]/NET0131 ,
		_w2611_,
		_w2615_,
		_w3246_
	);
	LUT3 #(
		.INIT('ha2)
	) name2794 (
		_w1100_,
		_w2623_,
		_w3246_,
		_w3247_
	);
	LUT4 #(
		.INIT('hde00)
	) name2795 (
		\EBX_reg[23]/NET0131 ,
		_w2623_,
		_w3245_,
		_w3247_,
		_w3248_
	);
	LUT2 #(
		.INIT('h2)
	) name2796 (
		\rEIP_reg[23]/NET0131 ,
		_w2640_,
		_w3249_
	);
	LUT3 #(
		.INIT('h23)
	) name2797 (
		\DataWidth_reg[1]/NET0131 ,
		\EBX_reg[23]/NET0131 ,
		_w633_,
		_w3250_
	);
	LUT3 #(
		.INIT('h08)
	) name2798 (
		_w570_,
		_w611_,
		_w3250_,
		_w3251_
	);
	LUT3 #(
		.INIT('hd0)
	) name2799 (
		_w2642_,
		_w3246_,
		_w3251_,
		_w3252_
	);
	LUT2 #(
		.INIT('h1)
	) name2800 (
		_w3249_,
		_w3252_,
		_w3253_
	);
	LUT4 #(
		.INIT('h5f13)
	) name2801 (
		\PhyAddrPointer_reg[23]/NET0131 ,
		\rEIP_reg[23]/NET0131 ,
		_w718_,
		_w2661_,
		_w3254_
	);
	LUT4 #(
		.INIT('h7500)
	) name2802 (
		_w695_,
		_w3248_,
		_w3253_,
		_w3254_,
		_w3255_
	);
	LUT2 #(
		.INIT('hb)
	) name2803 (
		_w3244_,
		_w3255_,
		_w3256_
	);
	LUT3 #(
		.INIT('h20)
	) name2804 (
		\PhyAddrPointer_reg[22]/NET0131 ,
		_w1463_,
		_w2652_,
		_w3257_
	);
	LUT4 #(
		.INIT('h0541)
	) name2805 (
		\DataWidth_reg[1]/NET0131 ,
		_w1279_,
		_w1607_,
		_w3257_,
		_w3258_
	);
	LUT2 #(
		.INIT('h2)
	) name2806 (
		\DataWidth_reg[1]/NET0131 ,
		\rEIP_reg[24]/NET0131 ,
		_w3259_
	);
	LUT2 #(
		.INIT('h2)
	) name2807 (
		_w700_,
		_w3259_,
		_w3260_
	);
	LUT2 #(
		.INIT('h4)
	) name2808 (
		_w3258_,
		_w3260_,
		_w3261_
	);
	LUT4 #(
		.INIT('h0509)
	) name2809 (
		\EBX_reg[24]/NET0131 ,
		\EBX_reg[31]/NET0131 ,
		_w2623_,
		_w2632_,
		_w3262_
	);
	LUT4 #(
		.INIT('h8000)
	) name2810 (
		\rEIP_reg[24]/NET0131 ,
		_w2605_,
		_w2611_,
		_w2615_,
		_w3263_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name2811 (
		\rEIP_reg[24]/NET0131 ,
		_w2605_,
		_w2611_,
		_w2615_,
		_w3264_
	);
	LUT3 #(
		.INIT('ha2)
	) name2812 (
		_w1100_,
		_w2623_,
		_w3264_,
		_w3265_
	);
	LUT2 #(
		.INIT('h4)
	) name2813 (
		_w3262_,
		_w3265_,
		_w3266_
	);
	LUT3 #(
		.INIT('h32)
	) name2814 (
		\DataWidth_reg[1]/NET0131 ,
		\EBX_reg[24]/NET0131 ,
		READY_n_pad,
		_w3267_
	);
	LUT3 #(
		.INIT('h02)
	) name2815 (
		_w611_,
		_w617_,
		_w3267_,
		_w3268_
	);
	LUT4 #(
		.INIT('h53f3)
	) name2816 (
		\EBX_reg[24]/NET0131 ,
		\rEIP_reg[24]/NET0131 ,
		_w611_,
		_w617_,
		_w3269_
	);
	LUT4 #(
		.INIT('h2f00)
	) name2817 (
		_w2623_,
		_w3264_,
		_w3268_,
		_w3269_,
		_w3270_
	);
	LUT4 #(
		.INIT('h01cf)
	) name2818 (
		_w566_,
		_w569_,
		_w570_,
		_w611_,
		_w3271_
	);
	LUT2 #(
		.INIT('h8)
	) name2819 (
		\rEIP_reg[24]/NET0131 ,
		_w3271_,
		_w3272_
	);
	LUT3 #(
		.INIT('h0d)
	) name2820 (
		_w570_,
		_w3270_,
		_w3272_,
		_w3273_
	);
	LUT4 #(
		.INIT('h5f13)
	) name2821 (
		\PhyAddrPointer_reg[24]/NET0131 ,
		\rEIP_reg[24]/NET0131 ,
		_w718_,
		_w2661_,
		_w3274_
	);
	LUT4 #(
		.INIT('h7500)
	) name2822 (
		_w695_,
		_w3266_,
		_w3273_,
		_w3274_,
		_w3275_
	);
	LUT2 #(
		.INIT('hb)
	) name2823 (
		_w3261_,
		_w3275_,
		_w3276_
	);
	LUT4 #(
		.INIT('h0400)
	) name2824 (
		_w1463_,
		_w1466_,
		_w1607_,
		_w3209_,
		_w3277_
	);
	LUT4 #(
		.INIT('h0541)
	) name2825 (
		\DataWidth_reg[1]/NET0131 ,
		_w1279_,
		_w1703_,
		_w3277_,
		_w3278_
	);
	LUT2 #(
		.INIT('h2)
	) name2826 (
		\DataWidth_reg[1]/NET0131 ,
		\rEIP_reg[25]/NET0131 ,
		_w3279_
	);
	LUT2 #(
		.INIT('h2)
	) name2827 (
		_w700_,
		_w3279_,
		_w3280_
	);
	LUT2 #(
		.INIT('h4)
	) name2828 (
		_w3278_,
		_w3280_,
		_w3281_
	);
	LUT3 #(
		.INIT('h8c)
	) name2829 (
		\EBX_reg[24]/NET0131 ,
		\EBX_reg[31]/NET0131 ,
		_w2632_,
		_w3282_
	);
	LUT4 #(
		.INIT('h4c8c)
	) name2830 (
		\rEIP_reg[25]/NET0131 ,
		_w1100_,
		_w2623_,
		_w3263_,
		_w3283_
	);
	LUT4 #(
		.INIT('hde00)
	) name2831 (
		\EBX_reg[25]/NET0131 ,
		_w2623_,
		_w3282_,
		_w3283_,
		_w3284_
	);
	LUT2 #(
		.INIT('h2)
	) name2832 (
		\rEIP_reg[25]/NET0131 ,
		_w2640_,
		_w3285_
	);
	LUT3 #(
		.INIT('h23)
	) name2833 (
		\DataWidth_reg[1]/NET0131 ,
		\EBX_reg[25]/NET0131 ,
		_w633_,
		_w3286_
	);
	LUT3 #(
		.INIT('h08)
	) name2834 (
		_w570_,
		_w611_,
		_w3286_,
		_w3287_
	);
	LUT4 #(
		.INIT('h7b00)
	) name2835 (
		\rEIP_reg[25]/NET0131 ,
		_w2642_,
		_w3263_,
		_w3287_,
		_w3288_
	);
	LUT2 #(
		.INIT('h1)
	) name2836 (
		_w3285_,
		_w3288_,
		_w3289_
	);
	LUT4 #(
		.INIT('h5f13)
	) name2837 (
		\PhyAddrPointer_reg[25]/NET0131 ,
		\rEIP_reg[25]/NET0131 ,
		_w718_,
		_w2661_,
		_w3290_
	);
	LUT4 #(
		.INIT('h7500)
	) name2838 (
		_w695_,
		_w3284_,
		_w3289_,
		_w3290_,
		_w3291_
	);
	LUT2 #(
		.INIT('hb)
	) name2839 (
		_w3281_,
		_w3291_,
		_w3292_
	);
	LUT4 #(
		.INIT('h0541)
	) name2840 (
		\DataWidth_reg[1]/NET0131 ,
		_w1279_,
		_w1626_,
		_w2655_,
		_w3293_
	);
	LUT2 #(
		.INIT('h2)
	) name2841 (
		\DataWidth_reg[1]/NET0131 ,
		\rEIP_reg[26]/NET0131 ,
		_w3294_
	);
	LUT2 #(
		.INIT('h2)
	) name2842 (
		_w700_,
		_w3294_,
		_w3295_
	);
	LUT2 #(
		.INIT('h4)
	) name2843 (
		_w3293_,
		_w3295_,
		_w3296_
	);
	LUT3 #(
		.INIT('h2a)
	) name2844 (
		\EBX_reg[31]/NET0131 ,
		_w2633_,
		_w2632_,
		_w3297_
	);
	LUT3 #(
		.INIT('h21)
	) name2845 (
		\EBX_reg[26]/NET0131 ,
		_w2623_,
		_w3297_,
		_w3298_
	);
	LUT4 #(
		.INIT('h78f0)
	) name2846 (
		\rEIP_reg[24]/NET0131 ,
		\rEIP_reg[25]/NET0131 ,
		\rEIP_reg[26]/NET0131 ,
		_w2616_,
		_w3299_
	);
	LUT3 #(
		.INIT('ha2)
	) name2847 (
		_w1100_,
		_w2623_,
		_w3299_,
		_w3300_
	);
	LUT2 #(
		.INIT('h2)
	) name2848 (
		\rEIP_reg[26]/NET0131 ,
		_w2640_,
		_w3301_
	);
	LUT3 #(
		.INIT('h23)
	) name2849 (
		\DataWidth_reg[1]/NET0131 ,
		\EBX_reg[26]/NET0131 ,
		_w633_,
		_w3302_
	);
	LUT3 #(
		.INIT('h08)
	) name2850 (
		_w570_,
		_w611_,
		_w3302_,
		_w3303_
	);
	LUT4 #(
		.INIT('h0233)
	) name2851 (
		_w2642_,
		_w3301_,
		_w3299_,
		_w3303_,
		_w3304_
	);
	LUT4 #(
		.INIT('h20aa)
	) name2852 (
		_w695_,
		_w3298_,
		_w3300_,
		_w3304_,
		_w3305_
	);
	LUT4 #(
		.INIT('h5f13)
	) name2853 (
		\PhyAddrPointer_reg[26]/NET0131 ,
		\rEIP_reg[26]/NET0131 ,
		_w718_,
		_w2661_,
		_w3306_
	);
	LUT3 #(
		.INIT('hef)
	) name2854 (
		_w3305_,
		_w3296_,
		_w3306_,
		_w3307_
	);
	LUT4 #(
		.INIT('h0541)
	) name2855 (
		\DataWidth_reg[1]/NET0131 ,
		_w1279_,
		_w1476_,
		_w2656_,
		_w3308_
	);
	LUT2 #(
		.INIT('h2)
	) name2856 (
		\DataWidth_reg[1]/NET0131 ,
		\rEIP_reg[27]/NET0131 ,
		_w3309_
	);
	LUT2 #(
		.INIT('h2)
	) name2857 (
		_w700_,
		_w3309_,
		_w3310_
	);
	LUT2 #(
		.INIT('h4)
	) name2858 (
		_w3308_,
		_w3310_,
		_w3311_
	);
	LUT3 #(
		.INIT('h2a)
	) name2859 (
		\EBX_reg[31]/NET0131 ,
		_w2632_,
		_w2634_,
		_w3312_
	);
	LUT4 #(
		.INIT('h48cc)
	) name2860 (
		\rEIP_reg[27]/NET0131 ,
		_w1100_,
		_w2619_,
		_w2623_,
		_w3313_
	);
	LUT4 #(
		.INIT('hde00)
	) name2861 (
		\EBX_reg[27]/NET0131 ,
		_w2623_,
		_w3312_,
		_w3313_,
		_w3314_
	);
	LUT2 #(
		.INIT('h2)
	) name2862 (
		\rEIP_reg[27]/NET0131 ,
		_w2640_,
		_w3315_
	);
	LUT4 #(
		.INIT('h2100)
	) name2863 (
		\rEIP_reg[27]/NET0131 ,
		_w617_,
		_w2619_,
		_w2623_,
		_w3316_
	);
	LUT3 #(
		.INIT('h23)
	) name2864 (
		\DataWidth_reg[1]/NET0131 ,
		\EBX_reg[27]/NET0131 ,
		_w633_,
		_w3317_
	);
	LUT3 #(
		.INIT('h08)
	) name2865 (
		_w570_,
		_w611_,
		_w3317_,
		_w3318_
	);
	LUT3 #(
		.INIT('h45)
	) name2866 (
		_w3315_,
		_w3316_,
		_w3318_,
		_w3319_
	);
	LUT4 #(
		.INIT('h5f13)
	) name2867 (
		\PhyAddrPointer_reg[27]/NET0131 ,
		\rEIP_reg[27]/NET0131 ,
		_w718_,
		_w2661_,
		_w3320_
	);
	LUT4 #(
		.INIT('h7500)
	) name2868 (
		_w695_,
		_w3314_,
		_w3319_,
		_w3320_,
		_w3321_
	);
	LUT2 #(
		.INIT('hb)
	) name2869 (
		_w3311_,
		_w3321_,
		_w3322_
	);
	LUT4 #(
		.INIT('h1000)
	) name2870 (
		_w1476_,
		_w1626_,
		_w2650_,
		_w2654_,
		_w3323_
	);
	LUT4 #(
		.INIT('h0541)
	) name2871 (
		\DataWidth_reg[1]/NET0131 ,
		_w1279_,
		_w1485_,
		_w3323_,
		_w3324_
	);
	LUT2 #(
		.INIT('h2)
	) name2872 (
		\DataWidth_reg[1]/NET0131 ,
		\rEIP_reg[28]/NET0131 ,
		_w3325_
	);
	LUT2 #(
		.INIT('h2)
	) name2873 (
		_w700_,
		_w3325_,
		_w3326_
	);
	LUT2 #(
		.INIT('h4)
	) name2874 (
		_w3324_,
		_w3326_,
		_w3327_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name2875 (
		\EBX_reg[27]/NET0131 ,
		\EBX_reg[31]/NET0131 ,
		_w2632_,
		_w2634_,
		_w3328_
	);
	LUT3 #(
		.INIT('h21)
	) name2876 (
		\EBX_reg[28]/NET0131 ,
		_w2623_,
		_w3328_,
		_w3329_
	);
	LUT4 #(
		.INIT('h9300)
	) name2877 (
		\rEIP_reg[27]/NET0131 ,
		\rEIP_reg[28]/NET0131 ,
		_w2619_,
		_w2623_,
		_w3330_
	);
	LUT2 #(
		.INIT('h2)
	) name2878 (
		_w1100_,
		_w3330_,
		_w3331_
	);
	LUT2 #(
		.INIT('h2)
	) name2879 (
		\rEIP_reg[28]/NET0131 ,
		_w2640_,
		_w3332_
	);
	LUT4 #(
		.INIT('h9300)
	) name2880 (
		\rEIP_reg[27]/NET0131 ,
		\rEIP_reg[28]/NET0131 ,
		_w2619_,
		_w2642_,
		_w3333_
	);
	LUT3 #(
		.INIT('h23)
	) name2881 (
		\DataWidth_reg[1]/NET0131 ,
		\EBX_reg[28]/NET0131 ,
		_w633_,
		_w3334_
	);
	LUT3 #(
		.INIT('h08)
	) name2882 (
		_w570_,
		_w611_,
		_w3334_,
		_w3335_
	);
	LUT3 #(
		.INIT('h45)
	) name2883 (
		_w3332_,
		_w3333_,
		_w3335_,
		_w3336_
	);
	LUT4 #(
		.INIT('h20aa)
	) name2884 (
		_w695_,
		_w3329_,
		_w3331_,
		_w3336_,
		_w3337_
	);
	LUT4 #(
		.INIT('h5f13)
	) name2885 (
		\PhyAddrPointer_reg[28]/NET0131 ,
		\rEIP_reg[28]/NET0131 ,
		_w718_,
		_w2661_,
		_w3338_
	);
	LUT3 #(
		.INIT('hef)
	) name2886 (
		_w3337_,
		_w3327_,
		_w3338_,
		_w3339_
	);
	LUT4 #(
		.INIT('h1000)
	) name2887 (
		\EBX_reg[27]/NET0131 ,
		\EBX_reg[28]/NET0131 ,
		_w2632_,
		_w2634_,
		_w3340_
	);
	LUT4 #(
		.INIT('h0509)
	) name2888 (
		\EBX_reg[29]/NET0131 ,
		\EBX_reg[31]/NET0131 ,
		_w2623_,
		_w3340_,
		_w3341_
	);
	LUT4 #(
		.INIT('h9500)
	) name2889 (
		\rEIP_reg[29]/NET0131 ,
		_w2619_,
		_w2620_,
		_w2623_,
		_w3342_
	);
	LUT2 #(
		.INIT('h2)
	) name2890 (
		_w1100_,
		_w3342_,
		_w3343_
	);
	LUT2 #(
		.INIT('h8)
	) name2891 (
		\rEIP_reg[29]/NET0131 ,
		_w3271_,
		_w3344_
	);
	LUT3 #(
		.INIT('h02)
	) name2892 (
		_w611_,
		_w617_,
		_w2635_,
		_w3345_
	);
	LUT4 #(
		.INIT('h53f3)
	) name2893 (
		\EBX_reg[29]/NET0131 ,
		\rEIP_reg[29]/NET0131 ,
		_w611_,
		_w617_,
		_w3346_
	);
	LUT4 #(
		.INIT('h20aa)
	) name2894 (
		_w570_,
		_w3342_,
		_w3345_,
		_w3346_,
		_w3347_
	);
	LUT4 #(
		.INIT('h1011)
	) name2895 (
		_w3344_,
		_w3347_,
		_w3341_,
		_w3343_,
		_w3348_
	);
	LUT3 #(
		.INIT('h81)
	) name2896 (
		\PhyAddrPointer_reg[25]/NET0131 ,
		\PhyAddrPointer_reg[26]/NET0131 ,
		_w1475_,
		_w3349_
	);
	LUT4 #(
		.INIT('h1000)
	) name2897 (
		_w1476_,
		_w1485_,
		_w3277_,
		_w3349_,
		_w3350_
	);
	LUT4 #(
		.INIT('h0541)
	) name2898 (
		\DataWidth_reg[1]/NET0131 ,
		_w1279_,
		_w1502_,
		_w3350_,
		_w3351_
	);
	LUT2 #(
		.INIT('h2)
	) name2899 (
		\DataWidth_reg[1]/NET0131 ,
		\rEIP_reg[29]/NET0131 ,
		_w3352_
	);
	LUT2 #(
		.INIT('h2)
	) name2900 (
		_w700_,
		_w3352_,
		_w3353_
	);
	LUT4 #(
		.INIT('h5f13)
	) name2901 (
		\PhyAddrPointer_reg[29]/NET0131 ,
		\rEIP_reg[29]/NET0131 ,
		_w718_,
		_w2661_,
		_w3354_
	);
	LUT3 #(
		.INIT('hb0)
	) name2902 (
		_w3351_,
		_w3353_,
		_w3354_,
		_w3355_
	);
	LUT3 #(
		.INIT('h2f)
	) name2903 (
		_w695_,
		_w3348_,
		_w3355_,
		_w3356_
	);
	LUT4 #(
		.INIT('h0541)
	) name2904 (
		\DataWidth_reg[1]/NET0131 ,
		_w1279_,
		_w2413_,
		_w3205_,
		_w3357_
	);
	LUT2 #(
		.INIT('h2)
	) name2905 (
		\DataWidth_reg[1]/NET0131 ,
		\rEIP_reg[2]/NET0131 ,
		_w3358_
	);
	LUT2 #(
		.INIT('h2)
	) name2906 (
		_w700_,
		_w3358_,
		_w3359_
	);
	LUT2 #(
		.INIT('h2)
	) name2907 (
		\rEIP_reg[2]/NET0131 ,
		_w2640_,
		_w3360_
	);
	LUT3 #(
		.INIT('h14)
	) name2908 (
		\DataWidth_reg[1]/NET0131 ,
		\rEIP_reg[1]/NET0131 ,
		\rEIP_reg[2]/NET0131 ,
		_w3361_
	);
	LUT4 #(
		.INIT('h0373)
	) name2909 (
		\DataWidth_reg[1]/NET0131 ,
		\EBX_reg[2]/NET0131 ,
		_w633_,
		_w3361_,
		_w3362_
	);
	LUT2 #(
		.INIT('h2)
	) name2910 (
		_w570_,
		_w3362_,
		_w3363_
	);
	LUT4 #(
		.INIT('h0110)
	) name2911 (
		\DataWidth_reg[1]/NET0131 ,
		READY_n_pad,
		\rEIP_reg[1]/NET0131 ,
		\rEIP_reg[2]/NET0131 ,
		_w3364_
	);
	LUT3 #(
		.INIT('he0)
	) name2912 (
		\EBX_reg[0]/NET0131 ,
		\EBX_reg[1]/NET0131 ,
		\EBX_reg[31]/NET0131 ,
		_w3365_
	);
	LUT4 #(
		.INIT('h0e0d)
	) name2913 (
		\EBX_reg[2]/NET0131 ,
		_w2623_,
		_w3364_,
		_w3365_,
		_w3366_
	);
	LUT4 #(
		.INIT('h3f15)
	) name2914 (
		_w566_,
		_w569_,
		_w655_,
		_w3366_,
		_w3367_
	);
	LUT3 #(
		.INIT('h8a)
	) name2915 (
		_w611_,
		_w3363_,
		_w3367_,
		_w3368_
	);
	LUT4 #(
		.INIT('h5f13)
	) name2916 (
		\PhyAddrPointer_reg[2]/NET0131 ,
		\rEIP_reg[2]/NET0131 ,
		_w718_,
		_w2661_,
		_w3369_
	);
	LUT4 #(
		.INIT('h5700)
	) name2917 (
		_w695_,
		_w3360_,
		_w3368_,
		_w3369_,
		_w3370_
	);
	LUT3 #(
		.INIT('h4f)
	) name2918 (
		_w3357_,
		_w3359_,
		_w3370_,
		_w3371_
	);
	LUT4 #(
		.INIT('h6a00)
	) name2919 (
		\rEIP_reg[30]/NET0131 ,
		_w2619_,
		_w2621_,
		_w2623_,
		_w3372_
	);
	LUT4 #(
		.INIT('h0001)
	) name2920 (
		\EBX_reg[26]/NET0131 ,
		\EBX_reg[27]/NET0131 ,
		\EBX_reg[28]/NET0131 ,
		\EBX_reg[29]/NET0131 ,
		_w3373_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name2921 (
		\EBX_reg[31]/NET0131 ,
		_w2633_,
		_w2632_,
		_w3373_,
		_w3374_
	);
	LUT4 #(
		.INIT('h0e0d)
	) name2922 (
		\EBX_reg[30]/NET0131 ,
		_w2623_,
		_w3372_,
		_w3374_,
		_w3375_
	);
	LUT2 #(
		.INIT('h2)
	) name2923 (
		_w1100_,
		_w3375_,
		_w3376_
	);
	LUT2 #(
		.INIT('h8)
	) name2924 (
		\rEIP_reg[30]/NET0131 ,
		_w3271_,
		_w3377_
	);
	LUT3 #(
		.INIT('hc8)
	) name2925 (
		\DataWidth_reg[1]/NET0131 ,
		\EBX_reg[30]/NET0131 ,
		READY_n_pad,
		_w3378_
	);
	LUT4 #(
		.INIT('h53f3)
	) name2926 (
		\EBX_reg[30]/NET0131 ,
		\rEIP_reg[30]/NET0131 ,
		_w611_,
		_w617_,
		_w3379_
	);
	LUT4 #(
		.INIT('h5700)
	) name2927 (
		_w659_,
		_w3372_,
		_w3378_,
		_w3379_,
		_w3380_
	);
	LUT3 #(
		.INIT('h31)
	) name2928 (
		_w570_,
		_w3377_,
		_w3380_,
		_w3381_
	);
	LUT3 #(
		.INIT('h8a)
	) name2929 (
		_w695_,
		_w3376_,
		_w3381_,
		_w3382_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name2930 (
		_w1279_,
		_w1502_,
		_w2656_,
		_w2649_,
		_w3383_
	);
	LUT2 #(
		.INIT('h2)
	) name2931 (
		\DataWidth_reg[1]/NET0131 ,
		\rEIP_reg[30]/NET0131 ,
		_w3384_
	);
	LUT2 #(
		.INIT('h2)
	) name2932 (
		_w700_,
		_w3384_,
		_w3385_
	);
	LUT4 #(
		.INIT('hbe00)
	) name2933 (
		\DataWidth_reg[1]/NET0131 ,
		_w1370_,
		_w3383_,
		_w3385_,
		_w3386_
	);
	LUT4 #(
		.INIT('h5f13)
	) name2934 (
		\PhyAddrPointer_reg[30]/NET0131 ,
		\rEIP_reg[30]/NET0131 ,
		_w718_,
		_w2661_,
		_w3387_
	);
	LUT2 #(
		.INIT('h4)
	) name2935 (
		_w3386_,
		_w3387_,
		_w3388_
	);
	LUT2 #(
		.INIT('hb)
	) name2936 (
		_w3382_,
		_w3388_,
		_w3389_
	);
	LUT3 #(
		.INIT('h40)
	) name2937 (
		\PhyAddrPointer_reg[0]/NET0131 ,
		\PhyAddrPointer_reg[1]/NET0131 ,
		\PhyAddrPointer_reg[2]/NET0131 ,
		_w3390_
	);
	LUT4 #(
		.INIT('h0541)
	) name2938 (
		\DataWidth_reg[1]/NET0131 ,
		_w1279_,
		_w2079_,
		_w3390_,
		_w3391_
	);
	LUT2 #(
		.INIT('h2)
	) name2939 (
		\DataWidth_reg[1]/NET0131 ,
		\rEIP_reg[3]/NET0131 ,
		_w3392_
	);
	LUT2 #(
		.INIT('h2)
	) name2940 (
		_w700_,
		_w3392_,
		_w3393_
	);
	LUT2 #(
		.INIT('h2)
	) name2941 (
		\rEIP_reg[3]/NET0131 ,
		_w2640_,
		_w3394_
	);
	LUT4 #(
		.INIT('hfe00)
	) name2942 (
		\EBX_reg[0]/NET0131 ,
		\EBX_reg[1]/NET0131 ,
		\EBX_reg[2]/NET0131 ,
		\EBX_reg[31]/NET0131 ,
		_w3395_
	);
	LUT3 #(
		.INIT('h12)
	) name2943 (
		\EBX_reg[3]/NET0131 ,
		_w2623_,
		_w3395_,
		_w3396_
	);
	LUT4 #(
		.INIT('h1540)
	) name2944 (
		\DataWidth_reg[1]/NET0131 ,
		\rEIP_reg[1]/NET0131 ,
		\rEIP_reg[2]/NET0131 ,
		\rEIP_reg[3]/NET0131 ,
		_w3397_
	);
	LUT2 #(
		.INIT('h4)
	) name2945 (
		READY_n_pad,
		_w3397_,
		_w3398_
	);
	LUT2 #(
		.INIT('h1)
	) name2946 (
		_w3396_,
		_w3398_,
		_w3399_
	);
	LUT2 #(
		.INIT('h2)
	) name2947 (
		_w566_,
		_w3399_,
		_w3400_
	);
	LUT4 #(
		.INIT('h0373)
	) name2948 (
		\DataWidth_reg[1]/NET0131 ,
		\EBX_reg[3]/NET0131 ,
		_w633_,
		_w3397_,
		_w3401_
	);
	LUT4 #(
		.INIT('hf531)
	) name2949 (
		_w569_,
		_w570_,
		_w648_,
		_w3401_,
		_w3402_
	);
	LUT3 #(
		.INIT('h8a)
	) name2950 (
		_w611_,
		_w3400_,
		_w3402_,
		_w3403_
	);
	LUT4 #(
		.INIT('h5f13)
	) name2951 (
		\PhyAddrPointer_reg[3]/NET0131 ,
		\rEIP_reg[3]/NET0131 ,
		_w718_,
		_w2661_,
		_w3404_
	);
	LUT4 #(
		.INIT('h5700)
	) name2952 (
		_w695_,
		_w3394_,
		_w3403_,
		_w3404_,
		_w3405_
	);
	LUT3 #(
		.INIT('h4f)
	) name2953 (
		_w3391_,
		_w3393_,
		_w3405_,
		_w3406_
	);
	LUT4 #(
		.INIT('h0541)
	) name2954 (
		\DataWidth_reg[1]/NET0131 ,
		_w1279_,
		_w1989_,
		_w3206_,
		_w3407_
	);
	LUT2 #(
		.INIT('h2)
	) name2955 (
		\DataWidth_reg[1]/NET0131 ,
		\rEIP_reg[4]/NET0131 ,
		_w3408_
	);
	LUT2 #(
		.INIT('h2)
	) name2956 (
		_w700_,
		_w3408_,
		_w3409_
	);
	LUT4 #(
		.INIT('h0309)
	) name2957 (
		\EBX_reg[31]/NET0131 ,
		\EBX_reg[4]/NET0131 ,
		_w2623_,
		_w2625_,
		_w3410_
	);
	LUT4 #(
		.INIT('h7f80)
	) name2958 (
		\rEIP_reg[1]/NET0131 ,
		\rEIP_reg[2]/NET0131 ,
		\rEIP_reg[3]/NET0131 ,
		\rEIP_reg[4]/NET0131 ,
		_w3411_
	);
	LUT2 #(
		.INIT('h2)
	) name2959 (
		_w2623_,
		_w3411_,
		_w3412_
	);
	LUT2 #(
		.INIT('h1)
	) name2960 (
		_w3410_,
		_w3412_,
		_w3413_
	);
	LUT3 #(
		.INIT('h80)
	) name2961 (
		_w566_,
		_w611_,
		_w3413_,
		_w3414_
	);
	LUT4 #(
		.INIT('hdc8c)
	) name2962 (
		\DataWidth_reg[1]/NET0131 ,
		\EBX_reg[4]/NET0131 ,
		_w633_,
		_w3411_,
		_w3415_
	);
	LUT3 #(
		.INIT('h80)
	) name2963 (
		_w570_,
		_w611_,
		_w3415_,
		_w3416_
	);
	LUT4 #(
		.INIT('h000d)
	) name2964 (
		\rEIP_reg[4]/NET0131 ,
		_w2640_,
		_w3414_,
		_w3416_,
		_w3417_
	);
	LUT2 #(
		.INIT('h2)
	) name2965 (
		\rEIP_reg[4]/NET0131 ,
		_w2661_,
		_w3418_
	);
	LUT3 #(
		.INIT('h07)
	) name2966 (
		\PhyAddrPointer_reg[4]/NET0131 ,
		_w718_,
		_w1109_,
		_w3419_
	);
	LUT2 #(
		.INIT('h4)
	) name2967 (
		_w3418_,
		_w3419_,
		_w3420_
	);
	LUT3 #(
		.INIT('hd0)
	) name2968 (
		_w695_,
		_w3417_,
		_w3420_,
		_w3421_
	);
	LUT3 #(
		.INIT('h4f)
	) name2969 (
		_w3407_,
		_w3409_,
		_w3421_,
		_w3422_
	);
	LUT4 #(
		.INIT('h0541)
	) name2970 (
		\DataWidth_reg[1]/NET0131 ,
		_w1279_,
		_w2087_,
		_w3207_,
		_w3423_
	);
	LUT2 #(
		.INIT('h2)
	) name2971 (
		\DataWidth_reg[1]/NET0131 ,
		\rEIP_reg[5]/NET0131 ,
		_w3424_
	);
	LUT2 #(
		.INIT('h2)
	) name2972 (
		_w700_,
		_w3424_,
		_w3425_
	);
	LUT3 #(
		.INIT('h8a)
	) name2973 (
		\EBX_reg[31]/NET0131 ,
		\EBX_reg[4]/NET0131 ,
		_w2625_,
		_w3426_
	);
	LUT3 #(
		.INIT('h90)
	) name2974 (
		\rEIP_reg[5]/NET0131 ,
		_w2606_,
		_w2623_,
		_w3427_
	);
	LUT4 #(
		.INIT('h00de)
	) name2975 (
		\EBX_reg[5]/NET0131 ,
		_w2623_,
		_w3426_,
		_w3427_,
		_w3428_
	);
	LUT3 #(
		.INIT('h80)
	) name2976 (
		_w566_,
		_w611_,
		_w3428_,
		_w3429_
	);
	LUT3 #(
		.INIT('h23)
	) name2977 (
		\DataWidth_reg[1]/NET0131 ,
		\EBX_reg[5]/NET0131 ,
		_w633_,
		_w3430_
	);
	LUT4 #(
		.INIT('h4010)
	) name2978 (
		\DataWidth_reg[1]/NET0131 ,
		\rEIP_reg[5]/NET0131 ,
		_w633_,
		_w2606_,
		_w3431_
	);
	LUT2 #(
		.INIT('h1)
	) name2979 (
		_w3430_,
		_w3431_,
		_w3432_
	);
	LUT3 #(
		.INIT('h80)
	) name2980 (
		_w570_,
		_w611_,
		_w3432_,
		_w3433_
	);
	LUT4 #(
		.INIT('h000d)
	) name2981 (
		\rEIP_reg[5]/NET0131 ,
		_w2640_,
		_w3429_,
		_w3433_,
		_w3434_
	);
	LUT2 #(
		.INIT('h2)
	) name2982 (
		\rEIP_reg[5]/NET0131 ,
		_w2661_,
		_w3435_
	);
	LUT3 #(
		.INIT('h07)
	) name2983 (
		\PhyAddrPointer_reg[5]/NET0131 ,
		_w718_,
		_w1109_,
		_w3436_
	);
	LUT2 #(
		.INIT('h4)
	) name2984 (
		_w3435_,
		_w3436_,
		_w3437_
	);
	LUT3 #(
		.INIT('hd0)
	) name2985 (
		_w695_,
		_w3434_,
		_w3437_,
		_w3438_
	);
	LUT3 #(
		.INIT('h4f)
	) name2986 (
		_w3423_,
		_w3425_,
		_w3438_,
		_w3439_
	);
	LUT3 #(
		.INIT('h40)
	) name2987 (
		\PhyAddrPointer_reg[0]/NET0131 ,
		\PhyAddrPointer_reg[1]/NET0131 ,
		_w1259_,
		_w3440_
	);
	LUT4 #(
		.INIT('h0541)
	) name2988 (
		\DataWidth_reg[1]/NET0131 ,
		_w1279_,
		_w2100_,
		_w3440_,
		_w3441_
	);
	LUT2 #(
		.INIT('h2)
	) name2989 (
		\DataWidth_reg[1]/NET0131 ,
		\rEIP_reg[6]/NET0131 ,
		_w3442_
	);
	LUT2 #(
		.INIT('h2)
	) name2990 (
		_w700_,
		_w3442_,
		_w3443_
	);
	LUT3 #(
		.INIT('h6c)
	) name2991 (
		\rEIP_reg[5]/NET0131 ,
		\rEIP_reg[6]/NET0131 ,
		_w2606_,
		_w3444_
	);
	LUT3 #(
		.INIT('he2)
	) name2992 (
		\EBX_reg[6]/NET0131 ,
		_w2642_,
		_w3444_,
		_w3445_
	);
	LUT4 #(
		.INIT('h9300)
	) name2993 (
		\rEIP_reg[5]/NET0131 ,
		\rEIP_reg[6]/NET0131 ,
		_w2606_,
		_w2623_,
		_w3446_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name2994 (
		\EBX_reg[31]/NET0131 ,
		\EBX_reg[4]/NET0131 ,
		\EBX_reg[5]/NET0131 ,
		_w2625_,
		_w3447_
	);
	LUT4 #(
		.INIT('h0d0e)
	) name2995 (
		\EBX_reg[6]/NET0131 ,
		_w2623_,
		_w3446_,
		_w3447_,
		_w3448_
	);
	LUT4 #(
		.INIT('h153f)
	) name2996 (
		_w566_,
		_w570_,
		_w3445_,
		_w3448_,
		_w3449_
	);
	LUT4 #(
		.INIT('h7505)
	) name2997 (
		\rEIP_reg[6]/NET0131 ,
		_w571_,
		_w611_,
		_w3449_,
		_w3450_
	);
	LUT2 #(
		.INIT('h2)
	) name2998 (
		\rEIP_reg[6]/NET0131 ,
		_w2661_,
		_w3451_
	);
	LUT3 #(
		.INIT('h07)
	) name2999 (
		\PhyAddrPointer_reg[6]/NET0131 ,
		_w718_,
		_w1109_,
		_w3452_
	);
	LUT2 #(
		.INIT('h4)
	) name3000 (
		_w3451_,
		_w3452_,
		_w3453_
	);
	LUT3 #(
		.INIT('hd0)
	) name3001 (
		_w695_,
		_w3450_,
		_w3453_,
		_w3454_
	);
	LUT3 #(
		.INIT('h4f)
	) name3002 (
		_w3441_,
		_w3443_,
		_w3454_,
		_w3455_
	);
	LUT4 #(
		.INIT('h4000)
	) name3003 (
		\PhyAddrPointer_reg[0]/NET0131 ,
		\PhyAddrPointer_reg[1]/NET0131 ,
		\PhyAddrPointer_reg[6]/NET0131 ,
		_w1259_,
		_w3456_
	);
	LUT4 #(
		.INIT('h0541)
	) name3004 (
		\DataWidth_reg[1]/NET0131 ,
		_w1279_,
		_w1782_,
		_w3456_,
		_w3457_
	);
	LUT2 #(
		.INIT('h2)
	) name3005 (
		\DataWidth_reg[1]/NET0131 ,
		\rEIP_reg[7]/NET0131 ,
		_w3458_
	);
	LUT2 #(
		.INIT('h2)
	) name3006 (
		_w700_,
		_w3458_,
		_w3459_
	);
	LUT4 #(
		.INIT('h78f0)
	) name3007 (
		\rEIP_reg[5]/NET0131 ,
		\rEIP_reg[6]/NET0131 ,
		\rEIP_reg[7]/NET0131 ,
		_w2606_,
		_w3460_
	);
	LUT3 #(
		.INIT('he2)
	) name3008 (
		\EBX_reg[7]/NET0131 ,
		_w2642_,
		_w3460_,
		_w3461_
	);
	LUT3 #(
		.INIT('h80)
	) name3009 (
		_w570_,
		_w611_,
		_w3461_,
		_w3462_
	);
	LUT2 #(
		.INIT('h2)
	) name3010 (
		_w2623_,
		_w3460_,
		_w3463_
	);
	LUT4 #(
		.INIT('h0309)
	) name3011 (
		\EBX_reg[31]/NET0131 ,
		\EBX_reg[7]/NET0131 ,
		_w2623_,
		_w2626_,
		_w3464_
	);
	LUT2 #(
		.INIT('h1)
	) name3012 (
		_w3463_,
		_w3464_,
		_w3465_
	);
	LUT3 #(
		.INIT('h80)
	) name3013 (
		_w566_,
		_w611_,
		_w3465_,
		_w3466_
	);
	LUT4 #(
		.INIT('h000d)
	) name3014 (
		\rEIP_reg[7]/NET0131 ,
		_w2640_,
		_w3462_,
		_w3466_,
		_w3467_
	);
	LUT2 #(
		.INIT('h2)
	) name3015 (
		\rEIP_reg[7]/NET0131 ,
		_w2661_,
		_w3468_
	);
	LUT3 #(
		.INIT('h07)
	) name3016 (
		\PhyAddrPointer_reg[7]/NET0131 ,
		_w718_,
		_w1109_,
		_w3469_
	);
	LUT2 #(
		.INIT('h4)
	) name3017 (
		_w3468_,
		_w3469_,
		_w3470_
	);
	LUT3 #(
		.INIT('hd0)
	) name3018 (
		_w695_,
		_w3467_,
		_w3470_,
		_w3471_
	);
	LUT3 #(
		.INIT('h4f)
	) name3019 (
		_w3457_,
		_w3459_,
		_w3471_,
		_w3472_
	);
	LUT2 #(
		.INIT('h8)
	) name3020 (
		\PhyAddrPointer_reg[7]/NET0131 ,
		_w3456_,
		_w3473_
	);
	LUT4 #(
		.INIT('h0541)
	) name3021 (
		\DataWidth_reg[1]/NET0131 ,
		_w1279_,
		_w1712_,
		_w3473_,
		_w3474_
	);
	LUT2 #(
		.INIT('h2)
	) name3022 (
		\DataWidth_reg[1]/NET0131 ,
		\rEIP_reg[8]/NET0131 ,
		_w3475_
	);
	LUT2 #(
		.INIT('h2)
	) name3023 (
		_w700_,
		_w3475_,
		_w3476_
	);
	LUT2 #(
		.INIT('h2)
	) name3024 (
		\rEIP_reg[8]/NET0131 ,
		_w2640_,
		_w3477_
	);
	LUT4 #(
		.INIT('h3caa)
	) name3025 (
		\EBX_reg[8]/NET0131 ,
		\rEIP_reg[8]/NET0131 ,
		_w2607_,
		_w2642_,
		_w3478_
	);
	LUT2 #(
		.INIT('h8)
	) name3026 (
		_w570_,
		_w3478_,
		_w3479_
	);
	LUT3 #(
		.INIT('h8a)
	) name3027 (
		\EBX_reg[31]/NET0131 ,
		\EBX_reg[7]/NET0131 ,
		_w2626_,
		_w3480_
	);
	LUT3 #(
		.INIT('h21)
	) name3028 (
		\EBX_reg[8]/NET0131 ,
		_w2623_,
		_w3480_,
		_w3481_
	);
	LUT3 #(
		.INIT('h90)
	) name3029 (
		\rEIP_reg[8]/NET0131 ,
		_w2607_,
		_w2623_,
		_w3482_
	);
	LUT3 #(
		.INIT('h02)
	) name3030 (
		_w566_,
		_w3482_,
		_w3481_,
		_w3483_
	);
	LUT3 #(
		.INIT('ha8)
	) name3031 (
		_w611_,
		_w3479_,
		_w3483_,
		_w3484_
	);
	LUT2 #(
		.INIT('h2)
	) name3032 (
		\rEIP_reg[8]/NET0131 ,
		_w2661_,
		_w3485_
	);
	LUT3 #(
		.INIT('h07)
	) name3033 (
		\PhyAddrPointer_reg[8]/NET0131 ,
		_w718_,
		_w1109_,
		_w3486_
	);
	LUT2 #(
		.INIT('h4)
	) name3034 (
		_w3485_,
		_w3486_,
		_w3487_
	);
	LUT4 #(
		.INIT('h5700)
	) name3035 (
		_w695_,
		_w3477_,
		_w3484_,
		_w3487_,
		_w3488_
	);
	LUT3 #(
		.INIT('h4f)
	) name3036 (
		_w3474_,
		_w3476_,
		_w3488_,
		_w3489_
	);
	LUT3 #(
		.INIT('h6c)
	) name3037 (
		\PhyAddrPointer_reg[1]/NET0131 ,
		\PhyAddrPointer_reg[9]/NET0131 ,
		_w1261_,
		_w3490_
	);
	LUT4 #(
		.INIT('h0451)
	) name3038 (
		\DataWidth_reg[1]/NET0131 ,
		_w1279_,
		_w3208_,
		_w3490_,
		_w3491_
	);
	LUT2 #(
		.INIT('h2)
	) name3039 (
		\DataWidth_reg[1]/NET0131 ,
		\rEIP_reg[9]/NET0131 ,
		_w3492_
	);
	LUT2 #(
		.INIT('h2)
	) name3040 (
		_w700_,
		_w3492_,
		_w3493_
	);
	LUT2 #(
		.INIT('h2)
	) name3041 (
		\rEIP_reg[9]/NET0131 ,
		_w2640_,
		_w3494_
	);
	LUT4 #(
		.INIT('h9300)
	) name3042 (
		\rEIP_reg[8]/NET0131 ,
		\rEIP_reg[9]/NET0131 ,
		_w2607_,
		_w2642_,
		_w3495_
	);
	LUT3 #(
		.INIT('h23)
	) name3043 (
		\DataWidth_reg[1]/NET0131 ,
		\EBX_reg[9]/NET0131 ,
		_w633_,
		_w3496_
	);
	LUT3 #(
		.INIT('h02)
	) name3044 (
		_w570_,
		_w3496_,
		_w3495_,
		_w3497_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name3045 (
		\EBX_reg[31]/NET0131 ,
		\EBX_reg[7]/NET0131 ,
		\EBX_reg[8]/NET0131 ,
		_w2626_,
		_w3498_
	);
	LUT3 #(
		.INIT('h21)
	) name3046 (
		\EBX_reg[9]/NET0131 ,
		_w2623_,
		_w3498_,
		_w3499_
	);
	LUT4 #(
		.INIT('h9300)
	) name3047 (
		\rEIP_reg[8]/NET0131 ,
		\rEIP_reg[9]/NET0131 ,
		_w2607_,
		_w2623_,
		_w3500_
	);
	LUT3 #(
		.INIT('h02)
	) name3048 (
		_w566_,
		_w3500_,
		_w3499_,
		_w3501_
	);
	LUT3 #(
		.INIT('ha8)
	) name3049 (
		_w611_,
		_w3497_,
		_w3501_,
		_w3502_
	);
	LUT2 #(
		.INIT('h2)
	) name3050 (
		\rEIP_reg[9]/NET0131 ,
		_w2661_,
		_w3503_
	);
	LUT3 #(
		.INIT('h07)
	) name3051 (
		\PhyAddrPointer_reg[9]/NET0131 ,
		_w718_,
		_w1109_,
		_w3504_
	);
	LUT2 #(
		.INIT('h4)
	) name3052 (
		_w3503_,
		_w3504_,
		_w3505_
	);
	LUT4 #(
		.INIT('h5700)
	) name3053 (
		_w695_,
		_w3494_,
		_w3502_,
		_w3505_,
		_w3506_
	);
	LUT3 #(
		.INIT('h4f)
	) name3054 (
		_w3491_,
		_w3493_,
		_w3506_,
		_w3507_
	);
	LUT4 #(
		.INIT('h000d)
	) name3055 (
		\PhyAddrPointer_reg[1]/NET0131 ,
		_w1984_,
		_w2111_,
		_w2114_,
		_w3508_
	);
	LUT4 #(
		.INIT('h80cc)
	) name3056 (
		\DataWidth_reg[1]/NET0131 ,
		\PhyAddrPointer_reg[1]/NET0131 ,
		_w700_,
		_w1283_,
		_w3509_
	);
	LUT4 #(
		.INIT('h3310)
	) name3057 (
		\DataWidth_reg[1]/NET0131 ,
		\PhyAddrPointer_reg[1]/NET0131 ,
		_w700_,
		_w706_,
		_w3510_
	);
	LUT3 #(
		.INIT('h01)
	) name3058 (
		_w2118_,
		_w3510_,
		_w3509_,
		_w3511_
	);
	LUT3 #(
		.INIT('h2f)
	) name3059 (
		_w695_,
		_w3508_,
		_w3511_,
		_w3512_
	);
	LUT3 #(
		.INIT('h80)
	) name3060 (
		\PhyAddrPointer_reg[9]/NET0131 ,
		_w1261_,
		_w3205_,
		_w3513_
	);
	LUT4 #(
		.INIT('h0541)
	) name3061 (
		\DataWidth_reg[1]/NET0131 ,
		_w1279_,
		_w1764_,
		_w3513_,
		_w3514_
	);
	LUT2 #(
		.INIT('h2)
	) name3062 (
		\DataWidth_reg[1]/NET0131 ,
		\rEIP_reg[10]/NET0131 ,
		_w3515_
	);
	LUT2 #(
		.INIT('h2)
	) name3063 (
		_w700_,
		_w3515_,
		_w3516_
	);
	LUT2 #(
		.INIT('h2)
	) name3064 (
		\rEIP_reg[10]/NET0131 ,
		_w2640_,
		_w3517_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name3065 (
		\rEIP_reg[10]/NET0131 ,
		\rEIP_reg[8]/NET0131 ,
		\rEIP_reg[9]/NET0131 ,
		_w2607_,
		_w3518_
	);
	LUT2 #(
		.INIT('h2)
	) name3066 (
		_w2623_,
		_w3518_,
		_w3519_
	);
	LUT3 #(
		.INIT('h23)
	) name3067 (
		\DataWidth_reg[1]/NET0131 ,
		\EBX_reg[10]/NET0131 ,
		_w633_,
		_w3520_
	);
	LUT4 #(
		.INIT('h0509)
	) name3068 (
		\EBX_reg[10]/NET0131 ,
		\EBX_reg[31]/NET0131 ,
		_w2623_,
		_w2627_,
		_w3521_
	);
	LUT4 #(
		.INIT('hf351)
	) name3069 (
		_w566_,
		_w570_,
		_w3520_,
		_w3521_,
		_w3522_
	);
	LUT3 #(
		.INIT('h08)
	) name3070 (
		_w570_,
		_w617_,
		_w3520_,
		_w3523_
	);
	LUT4 #(
		.INIT('haa02)
	) name3071 (
		_w611_,
		_w3519_,
		_w3522_,
		_w3523_,
		_w3524_
	);
	LUT2 #(
		.INIT('h2)
	) name3072 (
		\rEIP_reg[10]/NET0131 ,
		_w2661_,
		_w3525_
	);
	LUT3 #(
		.INIT('h07)
	) name3073 (
		\PhyAddrPointer_reg[10]/NET0131 ,
		_w718_,
		_w1109_,
		_w3526_
	);
	LUT2 #(
		.INIT('h4)
	) name3074 (
		_w3525_,
		_w3526_,
		_w3527_
	);
	LUT4 #(
		.INIT('h5700)
	) name3075 (
		_w695_,
		_w3517_,
		_w3524_,
		_w3527_,
		_w3528_
	);
	LUT3 #(
		.INIT('h4f)
	) name3076 (
		_w3514_,
		_w3516_,
		_w3528_,
		_w3529_
	);
	LUT2 #(
		.INIT('h4)
	) name3077 (
		\PhyAddrPointer_reg[0]/NET0131 ,
		_w1549_,
		_w3530_
	);
	LUT4 #(
		.INIT('h0541)
	) name3078 (
		\DataWidth_reg[1]/NET0131 ,
		_w1279_,
		_w1550_,
		_w3530_,
		_w3531_
	);
	LUT2 #(
		.INIT('h2)
	) name3079 (
		\DataWidth_reg[1]/NET0131 ,
		\rEIP_reg[11]/NET0131 ,
		_w3532_
	);
	LUT2 #(
		.INIT('h2)
	) name3080 (
		_w700_,
		_w3532_,
		_w3533_
	);
	LUT2 #(
		.INIT('h2)
	) name3081 (
		\rEIP_reg[11]/NET0131 ,
		_w2640_,
		_w3534_
	);
	LUT3 #(
		.INIT('h90)
	) name3082 (
		\rEIP_reg[11]/NET0131 ,
		_w2608_,
		_w2623_,
		_w3535_
	);
	LUT3 #(
		.INIT('h23)
	) name3083 (
		\DataWidth_reg[1]/NET0131 ,
		\EBX_reg[11]/NET0131 ,
		_w633_,
		_w3536_
	);
	LUT3 #(
		.INIT('h8c)
	) name3084 (
		\EBX_reg[10]/NET0131 ,
		\EBX_reg[31]/NET0131 ,
		_w2627_,
		_w3537_
	);
	LUT3 #(
		.INIT('h21)
	) name3085 (
		\EBX_reg[11]/NET0131 ,
		_w2623_,
		_w3537_,
		_w3538_
	);
	LUT4 #(
		.INIT('hf351)
	) name3086 (
		_w566_,
		_w570_,
		_w3536_,
		_w3538_,
		_w3539_
	);
	LUT3 #(
		.INIT('h08)
	) name3087 (
		_w570_,
		_w617_,
		_w3536_,
		_w3540_
	);
	LUT4 #(
		.INIT('haa02)
	) name3088 (
		_w611_,
		_w3535_,
		_w3539_,
		_w3540_,
		_w3541_
	);
	LUT2 #(
		.INIT('h2)
	) name3089 (
		\rEIP_reg[11]/NET0131 ,
		_w2661_,
		_w3542_
	);
	LUT3 #(
		.INIT('h07)
	) name3090 (
		\PhyAddrPointer_reg[11]/NET0131 ,
		_w718_,
		_w1109_,
		_w3543_
	);
	LUT2 #(
		.INIT('h4)
	) name3091 (
		_w3542_,
		_w3543_,
		_w3544_
	);
	LUT4 #(
		.INIT('h5700)
	) name3092 (
		_w695_,
		_w3534_,
		_w3541_,
		_w3544_,
		_w3545_
	);
	LUT3 #(
		.INIT('h4f)
	) name3093 (
		_w3531_,
		_w3533_,
		_w3545_,
		_w3546_
	);
	LUT3 #(
		.INIT('h6a)
	) name3094 (
		\PhyAddrPointer_reg[12]/NET0131 ,
		\PhyAddrPointer_reg[1]/NET0131 ,
		_w1263_,
		_w3547_
	);
	LUT2 #(
		.INIT('h8)
	) name3095 (
		_w1263_,
		_w3205_,
		_w3548_
	);
	LUT4 #(
		.INIT('h0541)
	) name3096 (
		\DataWidth_reg[1]/NET0131 ,
		_w1279_,
		_w3547_,
		_w3548_,
		_w3549_
	);
	LUT2 #(
		.INIT('h2)
	) name3097 (
		\DataWidth_reg[1]/NET0131 ,
		\rEIP_reg[12]/NET0131 ,
		_w3550_
	);
	LUT2 #(
		.INIT('h2)
	) name3098 (
		_w700_,
		_w3550_,
		_w3551_
	);
	LUT2 #(
		.INIT('h2)
	) name3099 (
		\rEIP_reg[12]/NET0131 ,
		_w2640_,
		_w3552_
	);
	LUT4 #(
		.INIT('h9300)
	) name3100 (
		\rEIP_reg[11]/NET0131 ,
		\rEIP_reg[12]/NET0131 ,
		_w2608_,
		_w2623_,
		_w3553_
	);
	LUT3 #(
		.INIT('h23)
	) name3101 (
		\DataWidth_reg[1]/NET0131 ,
		\EBX_reg[12]/NET0131 ,
		_w633_,
		_w3554_
	);
	LUT4 #(
		.INIT('he0f0)
	) name3102 (
		\EBX_reg[10]/NET0131 ,
		\EBX_reg[11]/NET0131 ,
		\EBX_reg[31]/NET0131 ,
		_w2627_,
		_w3555_
	);
	LUT3 #(
		.INIT('h21)
	) name3103 (
		\EBX_reg[12]/NET0131 ,
		_w2623_,
		_w3555_,
		_w3556_
	);
	LUT4 #(
		.INIT('hf351)
	) name3104 (
		_w566_,
		_w570_,
		_w3554_,
		_w3556_,
		_w3557_
	);
	LUT3 #(
		.INIT('h08)
	) name3105 (
		_w570_,
		_w617_,
		_w3554_,
		_w3558_
	);
	LUT4 #(
		.INIT('haa02)
	) name3106 (
		_w611_,
		_w3553_,
		_w3557_,
		_w3558_,
		_w3559_
	);
	LUT2 #(
		.INIT('h2)
	) name3107 (
		\rEIP_reg[12]/NET0131 ,
		_w2661_,
		_w3560_
	);
	LUT3 #(
		.INIT('h07)
	) name3108 (
		\PhyAddrPointer_reg[12]/NET0131 ,
		_w718_,
		_w1109_,
		_w3561_
	);
	LUT2 #(
		.INIT('h4)
	) name3109 (
		_w3560_,
		_w3561_,
		_w3562_
	);
	LUT4 #(
		.INIT('h5700)
	) name3110 (
		_w695_,
		_w3552_,
		_w3559_,
		_w3562_,
		_w3563_
	);
	LUT3 #(
		.INIT('h4f)
	) name3111 (
		_w3549_,
		_w3551_,
		_w3563_,
		_w3564_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name3112 (
		\PhyAddrPointer_reg[12]/NET0131 ,
		\PhyAddrPointer_reg[13]/NET0131 ,
		\PhyAddrPointer_reg[1]/NET0131 ,
		_w1263_,
		_w3565_
	);
	LUT4 #(
		.INIT('h8000)
	) name3113 (
		\PhyAddrPointer_reg[12]/NET0131 ,
		\PhyAddrPointer_reg[1]/NET0131 ,
		_w1263_,
		_w3208_,
		_w3566_
	);
	LUT4 #(
		.INIT('h0541)
	) name3114 (
		\DataWidth_reg[1]/NET0131 ,
		_w1279_,
		_w3565_,
		_w3566_,
		_w3567_
	);
	LUT2 #(
		.INIT('h2)
	) name3115 (
		\DataWidth_reg[1]/NET0131 ,
		\rEIP_reg[13]/NET0131 ,
		_w3568_
	);
	LUT2 #(
		.INIT('h2)
	) name3116 (
		_w700_,
		_w3568_,
		_w3569_
	);
	LUT2 #(
		.INIT('h2)
	) name3117 (
		\rEIP_reg[13]/NET0131 ,
		_w2640_,
		_w3570_
	);
	LUT4 #(
		.INIT('h78f0)
	) name3118 (
		\rEIP_reg[11]/NET0131 ,
		\rEIP_reg[12]/NET0131 ,
		\rEIP_reg[13]/NET0131 ,
		_w2608_,
		_w3571_
	);
	LUT2 #(
		.INIT('h2)
	) name3119 (
		_w2642_,
		_w3571_,
		_w3572_
	);
	LUT3 #(
		.INIT('h23)
	) name3120 (
		\DataWidth_reg[1]/NET0131 ,
		\EBX_reg[13]/NET0131 ,
		_w633_,
		_w3573_
	);
	LUT3 #(
		.INIT('h02)
	) name3121 (
		_w570_,
		_w3573_,
		_w3572_,
		_w3574_
	);
	LUT3 #(
		.INIT('h2a)
	) name3122 (
		\EBX_reg[31]/NET0131 ,
		_w2627_,
		_w2628_,
		_w3575_
	);
	LUT3 #(
		.INIT('h21)
	) name3123 (
		\EBX_reg[13]/NET0131 ,
		_w2623_,
		_w3575_,
		_w3576_
	);
	LUT2 #(
		.INIT('h2)
	) name3124 (
		_w2623_,
		_w3571_,
		_w3577_
	);
	LUT3 #(
		.INIT('h02)
	) name3125 (
		_w566_,
		_w3577_,
		_w3576_,
		_w3578_
	);
	LUT3 #(
		.INIT('ha8)
	) name3126 (
		_w611_,
		_w3574_,
		_w3578_,
		_w3579_
	);
	LUT2 #(
		.INIT('h2)
	) name3127 (
		\rEIP_reg[13]/NET0131 ,
		_w2661_,
		_w3580_
	);
	LUT3 #(
		.INIT('h07)
	) name3128 (
		\PhyAddrPointer_reg[13]/NET0131 ,
		_w718_,
		_w1109_,
		_w3581_
	);
	LUT2 #(
		.INIT('h4)
	) name3129 (
		_w3580_,
		_w3581_,
		_w3582_
	);
	LUT4 #(
		.INIT('h5700)
	) name3130 (
		_w695_,
		_w3570_,
		_w3579_,
		_w3582_,
		_w3583_
	);
	LUT3 #(
		.INIT('h4f)
	) name3131 (
		_w3567_,
		_w3569_,
		_w3583_,
		_w3584_
	);
	LUT2 #(
		.INIT('h4)
	) name3132 (
		\PhyAddrPointer_reg[0]/NET0131 ,
		_w1449_,
		_w3585_
	);
	LUT4 #(
		.INIT('h0541)
	) name3133 (
		\DataWidth_reg[1]/NET0131 ,
		_w1279_,
		_w1559_,
		_w3585_,
		_w3586_
	);
	LUT2 #(
		.INIT('h2)
	) name3134 (
		\DataWidth_reg[1]/NET0131 ,
		\rEIP_reg[14]/NET0131 ,
		_w3587_
	);
	LUT2 #(
		.INIT('h2)
	) name3135 (
		_w700_,
		_w3587_,
		_w3588_
	);
	LUT2 #(
		.INIT('h2)
	) name3136 (
		\rEIP_reg[14]/NET0131 ,
		_w2640_,
		_w3589_
	);
	LUT3 #(
		.INIT('h90)
	) name3137 (
		\rEIP_reg[14]/NET0131 ,
		_w2610_,
		_w2642_,
		_w3590_
	);
	LUT3 #(
		.INIT('h23)
	) name3138 (
		\DataWidth_reg[1]/NET0131 ,
		\EBX_reg[14]/NET0131 ,
		_w633_,
		_w3591_
	);
	LUT3 #(
		.INIT('h02)
	) name3139 (
		_w570_,
		_w3591_,
		_w3590_,
		_w3592_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name3140 (
		\EBX_reg[13]/NET0131 ,
		\EBX_reg[31]/NET0131 ,
		_w2627_,
		_w2628_,
		_w3593_
	);
	LUT3 #(
		.INIT('h21)
	) name3141 (
		\EBX_reg[14]/NET0131 ,
		_w2623_,
		_w3593_,
		_w3594_
	);
	LUT3 #(
		.INIT('h90)
	) name3142 (
		\rEIP_reg[14]/NET0131 ,
		_w2610_,
		_w2623_,
		_w3595_
	);
	LUT3 #(
		.INIT('h02)
	) name3143 (
		_w566_,
		_w3595_,
		_w3594_,
		_w3596_
	);
	LUT3 #(
		.INIT('ha8)
	) name3144 (
		_w611_,
		_w3592_,
		_w3596_,
		_w3597_
	);
	LUT2 #(
		.INIT('h2)
	) name3145 (
		\rEIP_reg[14]/NET0131 ,
		_w2661_,
		_w3598_
	);
	LUT3 #(
		.INIT('h07)
	) name3146 (
		\PhyAddrPointer_reg[14]/NET0131 ,
		_w718_,
		_w1109_,
		_w3599_
	);
	LUT2 #(
		.INIT('h4)
	) name3147 (
		_w3598_,
		_w3599_,
		_w3600_
	);
	LUT4 #(
		.INIT('h5700)
	) name3148 (
		_w695_,
		_w3589_,
		_w3597_,
		_w3600_,
		_w3601_
	);
	LUT3 #(
		.INIT('h4f)
	) name3149 (
		_w3586_,
		_w3588_,
		_w3601_,
		_w3602_
	);
	LUT3 #(
		.INIT('h40)
	) name3150 (
		\PhyAddrPointer_reg[0]/NET0131 ,
		\PhyAddrPointer_reg[14]/NET0131 ,
		_w1449_,
		_w3603_
	);
	LUT4 #(
		.INIT('h0541)
	) name3151 (
		\DataWidth_reg[1]/NET0131 ,
		_w1279_,
		_w1450_,
		_w3603_,
		_w3604_
	);
	LUT2 #(
		.INIT('h2)
	) name3152 (
		\DataWidth_reg[1]/NET0131 ,
		\rEIP_reg[15]/NET0131 ,
		_w3605_
	);
	LUT2 #(
		.INIT('h2)
	) name3153 (
		_w700_,
		_w3605_,
		_w3606_
	);
	LUT2 #(
		.INIT('h2)
	) name3154 (
		\rEIP_reg[15]/NET0131 ,
		_w2640_,
		_w3607_
	);
	LUT3 #(
		.INIT('h23)
	) name3155 (
		\DataWidth_reg[1]/NET0131 ,
		\EBX_reg[15]/NET0131 ,
		_w633_,
		_w3608_
	);
	LUT4 #(
		.INIT('h0509)
	) name3156 (
		\EBX_reg[15]/NET0131 ,
		\EBX_reg[31]/NET0131 ,
		_w2623_,
		_w2629_,
		_w3609_
	);
	LUT4 #(
		.INIT('hf351)
	) name3157 (
		_w566_,
		_w570_,
		_w3608_,
		_w3609_,
		_w3610_
	);
	LUT3 #(
		.INIT('h6c)
	) name3158 (
		\rEIP_reg[14]/NET0131 ,
		\rEIP_reg[15]/NET0131 ,
		_w2610_,
		_w3611_
	);
	LUT4 #(
		.INIT('hf070)
	) name3159 (
		_w570_,
		_w617_,
		_w2623_,
		_w3608_,
		_w3612_
	);
	LUT4 #(
		.INIT('h008a)
	) name3160 (
		_w611_,
		_w3611_,
		_w3612_,
		_w3610_,
		_w3613_
	);
	LUT2 #(
		.INIT('h2)
	) name3161 (
		\rEIP_reg[15]/NET0131 ,
		_w2661_,
		_w3614_
	);
	LUT3 #(
		.INIT('h07)
	) name3162 (
		\PhyAddrPointer_reg[15]/NET0131 ,
		_w718_,
		_w1109_,
		_w3615_
	);
	LUT2 #(
		.INIT('h4)
	) name3163 (
		_w3614_,
		_w3615_,
		_w3616_
	);
	LUT4 #(
		.INIT('h5700)
	) name3164 (
		_w695_,
		_w3607_,
		_w3613_,
		_w3616_,
		_w3617_
	);
	LUT3 #(
		.INIT('h4f)
	) name3165 (
		_w3604_,
		_w3606_,
		_w3617_,
		_w3618_
	);
	LUT3 #(
		.INIT('h80)
	) name3166 (
		\PhyAddrPointer_reg[15]/NET0131 ,
		_w1452_,
		_w3205_,
		_w3619_
	);
	LUT4 #(
		.INIT('h0541)
	) name3167 (
		\DataWidth_reg[1]/NET0131 ,
		_w1279_,
		_w1658_,
		_w3619_,
		_w3620_
	);
	LUT2 #(
		.INIT('h2)
	) name3168 (
		\DataWidth_reg[1]/NET0131 ,
		\rEIP_reg[16]/NET0131 ,
		_w3621_
	);
	LUT2 #(
		.INIT('h2)
	) name3169 (
		_w700_,
		_w3621_,
		_w3622_
	);
	LUT4 #(
		.INIT('h78f0)
	) name3170 (
		\rEIP_reg[14]/NET0131 ,
		\rEIP_reg[15]/NET0131 ,
		\rEIP_reg[16]/NET0131 ,
		_w2610_,
		_w3623_
	);
	LUT3 #(
		.INIT('h04)
	) name3171 (
		_w617_,
		_w2623_,
		_w3623_,
		_w3624_
	);
	LUT3 #(
		.INIT('h23)
	) name3172 (
		\DataWidth_reg[1]/NET0131 ,
		\EBX_reg[16]/NET0131 ,
		_w633_,
		_w3625_
	);
	LUT3 #(
		.INIT('h08)
	) name3173 (
		_w570_,
		_w611_,
		_w3625_,
		_w3626_
	);
	LUT2 #(
		.INIT('h4)
	) name3174 (
		_w3624_,
		_w3626_,
		_w3627_
	);
	LUT3 #(
		.INIT('h8c)
	) name3175 (
		\EBX_reg[15]/NET0131 ,
		\EBX_reg[31]/NET0131 ,
		_w2629_,
		_w3628_
	);
	LUT3 #(
		.INIT('h21)
	) name3176 (
		\EBX_reg[16]/NET0131 ,
		_w2623_,
		_w3628_,
		_w3629_
	);
	LUT4 #(
		.INIT('h8808)
	) name3177 (
		_w566_,
		_w611_,
		_w2623_,
		_w3623_,
		_w3630_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name3178 (
		\rEIP_reg[16]/NET0131 ,
		_w2640_,
		_w3629_,
		_w3630_,
		_w3631_
	);
	LUT2 #(
		.INIT('h2)
	) name3179 (
		\rEIP_reg[16]/NET0131 ,
		_w2661_,
		_w3632_
	);
	LUT3 #(
		.INIT('h07)
	) name3180 (
		\PhyAddrPointer_reg[16]/NET0131 ,
		_w718_,
		_w1109_,
		_w3633_
	);
	LUT2 #(
		.INIT('h4)
	) name3181 (
		_w3632_,
		_w3633_,
		_w3634_
	);
	LUT4 #(
		.INIT('h7500)
	) name3182 (
		_w695_,
		_w3627_,
		_w3631_,
		_w3634_,
		_w3635_
	);
	LUT3 #(
		.INIT('h4f)
	) name3183 (
		_w3620_,
		_w3622_,
		_w3635_,
		_w3636_
	);
	LUT3 #(
		.INIT('h80)
	) name3184 (
		\PhyAddrPointer_reg[1]/NET0131 ,
		_w1656_,
		_w3208_,
		_w3637_
	);
	LUT4 #(
		.INIT('h0541)
	) name3185 (
		\DataWidth_reg[1]/NET0131 ,
		_w1279_,
		_w1675_,
		_w3637_,
		_w3638_
	);
	LUT2 #(
		.INIT('h2)
	) name3186 (
		\DataWidth_reg[1]/NET0131 ,
		\rEIP_reg[17]/NET0131 ,
		_w3639_
	);
	LUT2 #(
		.INIT('h2)
	) name3187 (
		_w700_,
		_w3639_,
		_w3640_
	);
	LUT3 #(
		.INIT('h60)
	) name3188 (
		\rEIP_reg[17]/NET0131 ,
		_w2611_,
		_w2623_,
		_w3641_
	);
	LUT4 #(
		.INIT('hc355)
	) name3189 (
		\EBX_reg[17]/NET0131 ,
		\rEIP_reg[17]/NET0131 ,
		_w2611_,
		_w2623_,
		_w3642_
	);
	LUT4 #(
		.INIT('h53f3)
	) name3190 (
		\EBX_reg[17]/NET0131 ,
		\rEIP_reg[17]/NET0131 ,
		_w611_,
		_w617_,
		_w3643_
	);
	LUT4 #(
		.INIT('h08aa)
	) name3191 (
		_w570_,
		_w659_,
		_w3642_,
		_w3643_,
		_w3644_
	);
	LUT2 #(
		.INIT('h8)
	) name3192 (
		\rEIP_reg[17]/NET0131 ,
		_w3271_,
		_w3645_
	);
	LUT4 #(
		.INIT('he0f0)
	) name3193 (
		\EBX_reg[15]/NET0131 ,
		\EBX_reg[16]/NET0131 ,
		\EBX_reg[31]/NET0131 ,
		_w2629_,
		_w3646_
	);
	LUT3 #(
		.INIT('h12)
	) name3194 (
		\EBX_reg[17]/NET0131 ,
		_w2623_,
		_w3646_,
		_w3647_
	);
	LUT3 #(
		.INIT('ha8)
	) name3195 (
		_w1100_,
		_w3641_,
		_w3647_,
		_w3648_
	);
	LUT4 #(
		.INIT('haaa8)
	) name3196 (
		_w695_,
		_w3645_,
		_w3648_,
		_w3644_,
		_w3649_
	);
	LUT2 #(
		.INIT('h2)
	) name3197 (
		\rEIP_reg[17]/NET0131 ,
		_w2661_,
		_w3650_
	);
	LUT3 #(
		.INIT('h07)
	) name3198 (
		\PhyAddrPointer_reg[17]/NET0131 ,
		_w718_,
		_w1109_,
		_w3651_
	);
	LUT2 #(
		.INIT('h4)
	) name3199 (
		_w3650_,
		_w3651_,
		_w3652_
	);
	LUT4 #(
		.INIT('hf4ff)
	) name3200 (
		_w3638_,
		_w3640_,
		_w3649_,
		_w3652_,
		_w3653_
	);
	LUT4 #(
		.INIT('h0541)
	) name3201 (
		\DataWidth_reg[1]/NET0131 ,
		_w1279_,
		_w1692_,
		_w2651_,
		_w3654_
	);
	LUT2 #(
		.INIT('h2)
	) name3202 (
		\DataWidth_reg[1]/NET0131 ,
		\rEIP_reg[18]/NET0131 ,
		_w3655_
	);
	LUT2 #(
		.INIT('h2)
	) name3203 (
		_w700_,
		_w3655_,
		_w3656_
	);
	LUT4 #(
		.INIT('h0509)
	) name3204 (
		\EBX_reg[18]/NET0131 ,
		\EBX_reg[31]/NET0131 ,
		_w2623_,
		_w2630_,
		_w3657_
	);
	LUT4 #(
		.INIT('h9300)
	) name3205 (
		\rEIP_reg[17]/NET0131 ,
		\rEIP_reg[18]/NET0131 ,
		_w2611_,
		_w2623_,
		_w3658_
	);
	LUT3 #(
		.INIT('h02)
	) name3206 (
		_w1100_,
		_w3658_,
		_w3657_,
		_w3659_
	);
	LUT4 #(
		.INIT('h9300)
	) name3207 (
		\rEIP_reg[17]/NET0131 ,
		\rEIP_reg[18]/NET0131 ,
		_w2611_,
		_w2642_,
		_w3660_
	);
	LUT3 #(
		.INIT('h23)
	) name3208 (
		\DataWidth_reg[1]/NET0131 ,
		\EBX_reg[18]/NET0131 ,
		_w633_,
		_w3661_
	);
	LUT3 #(
		.INIT('h08)
	) name3209 (
		_w570_,
		_w611_,
		_w3661_,
		_w3662_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name3210 (
		\rEIP_reg[18]/NET0131 ,
		_w2640_,
		_w3660_,
		_w3662_,
		_w3663_
	);
	LUT2 #(
		.INIT('h2)
	) name3211 (
		\rEIP_reg[18]/NET0131 ,
		_w2661_,
		_w3664_
	);
	LUT3 #(
		.INIT('h07)
	) name3212 (
		\PhyAddrPointer_reg[18]/NET0131 ,
		_w718_,
		_w1109_,
		_w3665_
	);
	LUT2 #(
		.INIT('h4)
	) name3213 (
		_w3664_,
		_w3665_,
		_w3666_
	);
	LUT4 #(
		.INIT('h7500)
	) name3214 (
		_w695_,
		_w3659_,
		_w3663_,
		_w3666_,
		_w3667_
	);
	LUT3 #(
		.INIT('h4f)
	) name3215 (
		_w3654_,
		_w3656_,
		_w3667_,
		_w3668_
	);
	LUT4 #(
		.INIT('h4000)
	) name3216 (
		\PhyAddrPointer_reg[0]/NET0131 ,
		\PhyAddrPointer_reg[18]/NET0131 ,
		\PhyAddrPointer_reg[1]/NET0131 ,
		_w1569_,
		_w3669_
	);
	LUT4 #(
		.INIT('h0541)
	) name3217 (
		\DataWidth_reg[1]/NET0131 ,
		_w1279_,
		_w1571_,
		_w3669_,
		_w3670_
	);
	LUT2 #(
		.INIT('h2)
	) name3218 (
		\DataWidth_reg[1]/NET0131 ,
		\rEIP_reg[19]/NET0131 ,
		_w3671_
	);
	LUT2 #(
		.INIT('h2)
	) name3219 (
		_w700_,
		_w3671_,
		_w3672_
	);
	LUT2 #(
		.INIT('h4)
	) name3220 (
		_w3670_,
		_w3672_,
		_w3673_
	);
	LUT4 #(
		.INIT('h78f0)
	) name3221 (
		\rEIP_reg[17]/NET0131 ,
		\rEIP_reg[18]/NET0131 ,
		\rEIP_reg[19]/NET0131 ,
		_w2611_,
		_w3674_
	);
	LUT3 #(
		.INIT('h23)
	) name3222 (
		\DataWidth_reg[1]/NET0131 ,
		\EBX_reg[19]/NET0131 ,
		_w633_,
		_w3675_
	);
	LUT3 #(
		.INIT('h08)
	) name3223 (
		_w570_,
		_w611_,
		_w3675_,
		_w3676_
	);
	LUT4 #(
		.INIT('hfb00)
	) name3224 (
		_w617_,
		_w2623_,
		_w3674_,
		_w3676_,
		_w3677_
	);
	LUT3 #(
		.INIT('h8c)
	) name3225 (
		\EBX_reg[18]/NET0131 ,
		\EBX_reg[31]/NET0131 ,
		_w2630_,
		_w3678_
	);
	LUT3 #(
		.INIT('h21)
	) name3226 (
		\EBX_reg[19]/NET0131 ,
		_w2623_,
		_w3678_,
		_w3679_
	);
	LUT3 #(
		.INIT('ha2)
	) name3227 (
		_w1100_,
		_w2623_,
		_w3674_,
		_w3680_
	);
	LUT2 #(
		.INIT('h2)
	) name3228 (
		\rEIP_reg[19]/NET0131 ,
		_w2640_,
		_w3681_
	);
	LUT4 #(
		.INIT('h000b)
	) name3229 (
		_w3679_,
		_w3680_,
		_w3681_,
		_w3677_,
		_w3682_
	);
	LUT2 #(
		.INIT('h2)
	) name3230 (
		\rEIP_reg[19]/NET0131 ,
		_w2661_,
		_w3683_
	);
	LUT3 #(
		.INIT('h07)
	) name3231 (
		\PhyAddrPointer_reg[19]/NET0131 ,
		_w718_,
		_w1109_,
		_w3684_
	);
	LUT2 #(
		.INIT('h4)
	) name3232 (
		_w3683_,
		_w3684_,
		_w3685_
	);
	LUT3 #(
		.INIT('hd0)
	) name3233 (
		_w695_,
		_w3682_,
		_w3685_,
		_w3686_
	);
	LUT2 #(
		.INIT('hb)
	) name3234 (
		_w3673_,
		_w3686_,
		_w3687_
	);
	LUT3 #(
		.INIT('h23)
	) name3235 (
		\DataWidth_reg[1]/NET0131 ,
		READY_n_pad,
		_w570_,
		_w3688_
	);
	LUT3 #(
		.INIT('h40)
	) name3236 (
		_w621_,
		_w2640_,
		_w3688_,
		_w3689_
	);
	LUT3 #(
		.INIT('hc8)
	) name3237 (
		\RequestPending_reg/NET0131 ,
		_w695_,
		_w2640_,
		_w3690_
	);
	LUT4 #(
		.INIT('hfff4)
	) name3238 (
		\State2_reg[0]/NET0131 ,
		\State2_reg[1]/NET0131 ,
		\State2_reg[2]/NET0131 ,
		\State2_reg[3]/NET0131 ,
		_w3691_
	);
	LUT4 #(
		.INIT('h80aa)
	) name3239 (
		\RequestPending_reg/NET0131 ,
		_w705_,
		_w717_,
		_w1824_,
		_w3692_
	);
	LUT2 #(
		.INIT('h2)
	) name3240 (
		_w3691_,
		_w3692_,
		_w3693_
	);
	LUT3 #(
		.INIT('h4f)
	) name3241 (
		_w3689_,
		_w3690_,
		_w3693_,
		_w3694_
	);
	LUT2 #(
		.INIT('h6)
	) name3242 (
		\EAX_reg[23]/NET0131 ,
		_w2048_,
		_w3695_
	);
	LUT3 #(
		.INIT('h21)
	) name3243 (
		\EAX_reg[23]/NET0131 ,
		_w617_,
		_w2048_,
		_w3696_
	);
	LUT3 #(
		.INIT('h08)
	) name3244 (
		_w570_,
		_w611_,
		_w3696_,
		_w3697_
	);
	LUT4 #(
		.INIT('haaa2)
	) name3245 (
		\Datao[23]_pad ,
		_w2153_,
		_w2154_,
		_w3697_,
		_w3698_
	);
	LUT2 #(
		.INIT('h8)
	) name3246 (
		_w570_,
		_w3695_,
		_w3699_
	);
	LUT3 #(
		.INIT('h80)
	) name3247 (
		_w570_,
		_w659_,
		_w3695_,
		_w3700_
	);
	LUT4 #(
		.INIT('h3f15)
	) name3248 (
		\Datao[23]_pad ,
		\uWord_reg[7]/NET0131 ,
		_w696_,
		_w2159_,
		_w3701_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name3249 (
		_w695_,
		_w3698_,
		_w3700_,
		_w3701_,
		_w3702_
	);
	LUT3 #(
		.INIT('h6c)
	) name3250 (
		\EAX_reg[18]/NET0131 ,
		\EAX_reg[19]/NET0131 ,
		_w2047_,
		_w3703_
	);
	LUT4 #(
		.INIT('h0903)
	) name3251 (
		\EAX_reg[18]/NET0131 ,
		\EAX_reg[19]/NET0131 ,
		_w617_,
		_w2047_,
		_w3704_
	);
	LUT3 #(
		.INIT('h08)
	) name3252 (
		_w570_,
		_w611_,
		_w3704_,
		_w3705_
	);
	LUT4 #(
		.INIT('haaa2)
	) name3253 (
		\Datao[19]_pad ,
		_w2153_,
		_w2154_,
		_w3705_,
		_w3706_
	);
	LUT3 #(
		.INIT('h80)
	) name3254 (
		_w570_,
		_w611_,
		_w3703_,
		_w3707_
	);
	LUT4 #(
		.INIT('h0800)
	) name3255 (
		_w570_,
		_w611_,
		_w617_,
		_w3703_,
		_w3708_
	);
	LUT4 #(
		.INIT('h3f15)
	) name3256 (
		\Datao[19]_pad ,
		\uWord_reg[3]/NET0131 ,
		_w696_,
		_w2159_,
		_w3709_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name3257 (
		_w695_,
		_w3706_,
		_w3708_,
		_w3709_,
		_w3710_
	);
	LUT2 #(
		.INIT('h2)
	) name3258 (
		\uWord_reg[3]/NET0131 ,
		_w1825_,
		_w3711_
	);
	LUT4 #(
		.INIT('h1d3f)
	) name3259 (
		\Datai[3]_pad ,
		READY_n_pad,
		\uWord_reg[3]/NET0131 ,
		_w611_,
		_w3712_
	);
	LUT2 #(
		.INIT('h2)
	) name3260 (
		_w566_,
		_w3712_,
		_w3713_
	);
	LUT4 #(
		.INIT('h02aa)
	) name3261 (
		\uWord_reg[3]/NET0131 ,
		_w566_,
		_w570_,
		_w611_,
		_w3714_
	);
	LUT4 #(
		.INIT('haaa8)
	) name3262 (
		_w695_,
		_w3707_,
		_w3713_,
		_w3714_,
		_w3715_
	);
	LUT2 #(
		.INIT('he)
	) name3263 (
		_w3711_,
		_w3715_,
		_w3716_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name3264 (
		\uWord_reg[7]/NET0131 ,
		_w695_,
		_w1825_,
		_w2058_,
		_w3717_
	);
	LUT2 #(
		.INIT('h8)
	) name3265 (
		\Datai[7]_pad ,
		_w566_,
		_w3718_
	);
	LUT3 #(
		.INIT('h20)
	) name3266 (
		\Datai[7]_pad ,
		READY_n_pad,
		_w566_,
		_w3719_
	);
	LUT3 #(
		.INIT('ha8)
	) name3267 (
		_w2175_,
		_w3699_,
		_w3719_,
		_w3720_
	);
	LUT2 #(
		.INIT('he)
	) name3268 (
		_w3717_,
		_w3720_,
		_w3721_
	);
	LUT3 #(
		.INIT('h2a)
	) name3269 (
		\MemoryFetch_reg/NET0131 ,
		_w569_,
		_w611_,
		_w3722_
	);
	LUT3 #(
		.INIT('hc4)
	) name3270 (
		\MemoryFetch_reg/NET0131 ,
		_w2039_,
		_w2040_,
		_w3723_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name3271 (
		_w695_,
		_w2057_,
		_w3722_,
		_w3723_,
		_w3724_
	);
	LUT4 #(
		.INIT('hc0e0)
	) name3272 (
		\ReadRequest_reg/NET0131 ,
		_w643_,
		_w695_,
		_w2153_,
		_w3725_
	);
	LUT3 #(
		.INIT('hc4)
	) name3273 (
		\ReadRequest_reg/NET0131 ,
		_w2039_,
		_w2040_,
		_w3726_
	);
	LUT2 #(
		.INIT('hb)
	) name3274 (
		_w3725_,
		_w3726_,
		_w3727_
	);
	LUT4 #(
		.INIT('h5445)
	) name3275 (
		\EBX_reg[0]/NET0131 ,
		\State_reg[0]/NET0131 ,
		\State_reg[1]/NET0131 ,
		\State_reg[2]/NET0131 ,
		_w3728_
	);
	LUT4 #(
		.INIT('h5f1f)
	) name3276 (
		_w566_,
		_w570_,
		_w611_,
		_w3728_,
		_w3729_
	);
	LUT3 #(
		.INIT('h32)
	) name3277 (
		\DataWidth_reg[1]/NET0131 ,
		\EBX_reg[0]/NET0131 ,
		READY_n_pad,
		_w3730_
	);
	LUT4 #(
		.INIT('h222a)
	) name3278 (
		\rEIP_reg[0]/NET0131 ,
		_w2640_,
		_w3729_,
		_w3730_,
		_w3731_
	);
	LUT2 #(
		.INIT('h4)
	) name3279 (
		\InstQueueRd_Addr_reg[0]/NET0131 ,
		_w569_,
		_w3732_
	);
	LUT4 #(
		.INIT('h3f11)
	) name3280 (
		_w566_,
		_w570_,
		_w617_,
		_w2623_,
		_w3733_
	);
	LUT4 #(
		.INIT('hc0c8)
	) name3281 (
		\EBX_reg[0]/NET0131 ,
		_w611_,
		_w3732_,
		_w3733_,
		_w3734_
	);
	LUT4 #(
		.INIT('hcc40)
	) name3282 (
		\DataWidth_reg[1]/NET0131 ,
		\PhyAddrPointer_reg[0]/NET0131 ,
		_w700_,
		_w718_,
		_w3735_
	);
	LUT4 #(
		.INIT('h0700)
	) name3283 (
		\DataWidth_reg[1]/NET0131 ,
		_w700_,
		_w706_,
		_w2077_,
		_w3736_
	);
	LUT3 #(
		.INIT('h31)
	) name3284 (
		\rEIP_reg[0]/NET0131 ,
		_w3735_,
		_w3736_,
		_w3737_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name3285 (
		_w695_,
		_w3731_,
		_w3734_,
		_w3737_,
		_w3738_
	);
	LUT4 #(
		.INIT('h8000)
	) name3286 (
		\EAX_reg[27]/NET0131 ,
		\EAX_reg[28]/NET0131 ,
		\EAX_reg[29]/NET0131 ,
		_w2051_,
		_w3739_
	);
	LUT4 #(
		.INIT('hd0e0)
	) name3287 (
		\EAX_reg[30]/NET0131 ,
		_w617_,
		_w2149_,
		_w3739_,
		_w3740_
	);
	LUT4 #(
		.INIT('h4080)
	) name3288 (
		\EAX_reg[30]/NET0131 ,
		_w570_,
		_w659_,
		_w3739_,
		_w3741_
	);
	LUT4 #(
		.INIT('h005d)
	) name3289 (
		\Datao[30]_pad ,
		_w2155_,
		_w3740_,
		_w3741_,
		_w3742_
	);
	LUT4 #(
		.INIT('h3f15)
	) name3290 (
		\Datao[30]_pad ,
		\uWord_reg[14]/NET0131 ,
		_w696_,
		_w2159_,
		_w3743_
	);
	LUT3 #(
		.INIT('h2f)
	) name3291 (
		_w695_,
		_w3742_,
		_w3743_,
		_w3744_
	);
	LUT3 #(
		.INIT('h48)
	) name3292 (
		\EAX_reg[28]/NET0131 ,
		_w1848_,
		_w1845_,
		_w3745_
	);
	LUT3 #(
		.INIT('h8a)
	) name3293 (
		\EAX_reg[28]/NET0131 ,
		_w635_,
		_w1852_,
		_w3746_
	);
	LUT4 #(
		.INIT('h08a2)
	) name3294 (
		_w605_,
		_w1907_,
		_w1918_,
		_w1929_,
		_w3747_
	);
	LUT2 #(
		.INIT('h8)
	) name3295 (
		_w580_,
		_w3747_,
		_w3748_
	);
	LUT3 #(
		.INIT('h80)
	) name3296 (
		\Datai[28]_pad ,
		_w514_,
		_w569_,
		_w3749_
	);
	LUT3 #(
		.INIT('ha8)
	) name3297 (
		_w612_,
		_w2054_,
		_w3749_,
		_w3750_
	);
	LUT2 #(
		.INIT('h1)
	) name3298 (
		_w3748_,
		_w3750_,
		_w3751_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name3299 (
		_w695_,
		_w3745_,
		_w3746_,
		_w3751_,
		_w3752_
	);
	LUT2 #(
		.INIT('h2)
	) name3300 (
		\EAX_reg[28]/NET0131 ,
		_w1825_,
		_w3753_
	);
	LUT2 #(
		.INIT('he)
	) name3301 (
		_w3752_,
		_w3753_,
		_w3754_
	);
	LUT2 #(
		.INIT('h2)
	) name3302 (
		\uWord_reg[14]/NET0131 ,
		_w1825_,
		_w3755_
	);
	LUT2 #(
		.INIT('h8)
	) name3303 (
		\Datai[14]_pad ,
		_w566_,
		_w3756_
	);
	LUT3 #(
		.INIT('h20)
	) name3304 (
		\Datai[14]_pad ,
		READY_n_pad,
		_w566_,
		_w3757_
	);
	LUT4 #(
		.INIT('h00b7)
	) name3305 (
		\EAX_reg[30]/NET0131 ,
		_w570_,
		_w3739_,
		_w3757_,
		_w3758_
	);
	LUT2 #(
		.INIT('h2)
	) name3306 (
		\uWord_reg[14]/NET0131 ,
		_w2058_,
		_w3759_
	);
	LUT4 #(
		.INIT('hcc08)
	) name3307 (
		_w611_,
		_w695_,
		_w3758_,
		_w3759_,
		_w3760_
	);
	LUT2 #(
		.INIT('he)
	) name3308 (
		_w3755_,
		_w3760_,
		_w3761_
	);
	LUT3 #(
		.INIT('h20)
	) name3309 (
		\Datai[0]_pad ,
		READY_n_pad,
		_w643_,
		_w3762_
	);
	LUT4 #(
		.INIT('h0080)
	) name3310 (
		_w576_,
		_w579_,
		_w605_,
		_w792_,
		_w3763_
	);
	LUT2 #(
		.INIT('h4)
	) name3311 (
		\EAX_reg[0]/NET0131 ,
		_w1848_,
		_w3764_
	);
	LUT2 #(
		.INIT('h1)
	) name3312 (
		_w3763_,
		_w3764_,
		_w3765_
	);
	LUT3 #(
		.INIT('h8a)
	) name3313 (
		_w695_,
		_w3762_,
		_w3765_,
		_w3766_
	);
	LUT3 #(
		.INIT('hf2)
	) name3314 (
		\EAX_reg[0]/NET0131 ,
		_w2668_,
		_w3766_,
		_w3767_
	);
	LUT4 #(
		.INIT('h1333)
	) name3315 (
		\EBX_reg[27]/NET0131 ,
		\EBX_reg[28]/NET0131 ,
		_w1958_,
		_w2143_,
		_w3768_
	);
	LUT3 #(
		.INIT('h80)
	) name3316 (
		_w1958_,
		_w2143_,
		_w2180_,
		_w3769_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name3317 (
		_w590_,
		_w1958_,
		_w2143_,
		_w2180_,
		_w3770_
	);
	LUT4 #(
		.INIT('h135f)
	) name3318 (
		\EBX_reg[28]/NET0131 ,
		_w577_,
		_w1975_,
		_w3747_,
		_w3771_
	);
	LUT4 #(
		.INIT('h20aa)
	) name3319 (
		_w695_,
		_w3768_,
		_w3770_,
		_w3771_,
		_w3772_
	);
	LUT2 #(
		.INIT('h2)
	) name3320 (
		\EBX_reg[28]/NET0131 ,
		_w1825_,
		_w3773_
	);
	LUT2 #(
		.INIT('he)
	) name3321 (
		_w3772_,
		_w3773_,
		_w3774_
	);
	LUT3 #(
		.INIT('h8a)
	) name3322 (
		\EAX_reg[16]/NET0131 ,
		_w635_,
		_w1852_,
		_w3775_
	);
	LUT3 #(
		.INIT('h48)
	) name3323 (
		\EAX_reg[16]/NET0131 ,
		_w1848_,
		_w1835_,
		_w3776_
	);
	LUT4 #(
		.INIT('h153f)
	) name3324 (
		\InstQueue_reg[12][0]/NET0131 ,
		\InstQueue_reg[1][0]/NET0131 ,
		_w460_,
		_w454_,
		_w3777_
	);
	LUT4 #(
		.INIT('h153f)
	) name3325 (
		\InstQueue_reg[13][0]/NET0131 ,
		\InstQueue_reg[15][0]/NET0131 ,
		_w470_,
		_w471_,
		_w3778_
	);
	LUT4 #(
		.INIT('h135f)
	) name3326 (
		\InstQueue_reg[2][0]/NET0131 ,
		\InstQueue_reg[6][0]/NET0131 ,
		_w473_,
		_w476_,
		_w3779_
	);
	LUT4 #(
		.INIT('h153f)
	) name3327 (
		\InstQueue_reg[5][0]/NET0131 ,
		\InstQueue_reg[7][0]/NET0131 ,
		_w464_,
		_w474_,
		_w3780_
	);
	LUT4 #(
		.INIT('h8000)
	) name3328 (
		_w3779_,
		_w3780_,
		_w3777_,
		_w3778_,
		_w3781_
	);
	LUT4 #(
		.INIT('h153f)
	) name3329 (
		\InstQueue_reg[11][0]/NET0131 ,
		\InstQueue_reg[9][0]/NET0131 ,
		_w461_,
		_w468_,
		_w3782_
	);
	LUT4 #(
		.INIT('h153f)
	) name3330 (
		\InstQueue_reg[10][0]/NET0131 ,
		\InstQueue_reg[3][0]/NET0131 ,
		_w463_,
		_w477_,
		_w3783_
	);
	LUT4 #(
		.INIT('h135f)
	) name3331 (
		\InstQueue_reg[0][0]/NET0131 ,
		\InstQueue_reg[8][0]/NET0131 ,
		_w456_,
		_w467_,
		_w3784_
	);
	LUT4 #(
		.INIT('h153f)
	) name3332 (
		\InstQueue_reg[14][0]/NET0131 ,
		\InstQueue_reg[4][0]/NET0131 ,
		_w453_,
		_w458_,
		_w3785_
	);
	LUT4 #(
		.INIT('h8000)
	) name3333 (
		_w3784_,
		_w3785_,
		_w3782_,
		_w3783_,
		_w3786_
	);
	LUT2 #(
		.INIT('h8)
	) name3334 (
		_w3781_,
		_w3786_,
		_w3787_
	);
	LUT4 #(
		.INIT('h0080)
	) name3335 (
		_w576_,
		_w579_,
		_w605_,
		_w3787_,
		_w3788_
	);
	LUT3 #(
		.INIT('h80)
	) name3336 (
		\Datai[16]_pad ,
		_w514_,
		_w569_,
		_w3789_
	);
	LUT2 #(
		.INIT('h8)
	) name3337 (
		\Datai[0]_pad ,
		_w566_,
		_w3790_
	);
	LUT4 #(
		.INIT('h1113)
	) name3338 (
		_w612_,
		_w3788_,
		_w3789_,
		_w3790_,
		_w3791_
	);
	LUT2 #(
		.INIT('h4)
	) name3339 (
		_w3776_,
		_w3791_,
		_w3792_
	);
	LUT2 #(
		.INIT('h2)
	) name3340 (
		\EAX_reg[16]/NET0131 ,
		_w1825_,
		_w3793_
	);
	LUT4 #(
		.INIT('hff8a)
	) name3341 (
		_w695_,
		_w3775_,
		_w3792_,
		_w3793_,
		_w3794_
	);
	LUT4 #(
		.INIT('h70f0)
	) name3342 (
		\EAX_reg[16]/NET0131 ,
		\EAX_reg[17]/NET0131 ,
		_w1848_,
		_w1835_,
		_w3795_
	);
	LUT4 #(
		.INIT('h60c0)
	) name3343 (
		\EAX_reg[16]/NET0131 ,
		\EAX_reg[17]/NET0131 ,
		_w1848_,
		_w1835_,
		_w3796_
	);
	LUT4 #(
		.INIT('h153f)
	) name3344 (
		\InstQueue_reg[12][1]/NET0131 ,
		\InstQueue_reg[1][1]/NET0131 ,
		_w460_,
		_w454_,
		_w3797_
	);
	LUT4 #(
		.INIT('h153f)
	) name3345 (
		\InstQueue_reg[15][1]/NET0131 ,
		\InstQueue_reg[8][1]/NET0131 ,
		_w467_,
		_w470_,
		_w3798_
	);
	LUT4 #(
		.INIT('h135f)
	) name3346 (
		\InstQueue_reg[2][1]/NET0131 ,
		\InstQueue_reg[6][1]/NET0131 ,
		_w473_,
		_w476_,
		_w3799_
	);
	LUT4 #(
		.INIT('h153f)
	) name3347 (
		\InstQueue_reg[5][1]/NET0131 ,
		\InstQueue_reg[7][1]/NET0131 ,
		_w464_,
		_w474_,
		_w3800_
	);
	LUT4 #(
		.INIT('h8000)
	) name3348 (
		_w3799_,
		_w3800_,
		_w3797_,
		_w3798_,
		_w3801_
	);
	LUT4 #(
		.INIT('h153f)
	) name3349 (
		\InstQueue_reg[11][1]/NET0131 ,
		\InstQueue_reg[9][1]/NET0131 ,
		_w461_,
		_w468_,
		_w3802_
	);
	LUT4 #(
		.INIT('h135f)
	) name3350 (
		\InstQueue_reg[10][1]/NET0131 ,
		\InstQueue_reg[13][1]/NET0131 ,
		_w477_,
		_w471_,
		_w3803_
	);
	LUT4 #(
		.INIT('h153f)
	) name3351 (
		\InstQueue_reg[0][1]/NET0131 ,
		\InstQueue_reg[3][1]/NET0131 ,
		_w463_,
		_w456_,
		_w3804_
	);
	LUT4 #(
		.INIT('h153f)
	) name3352 (
		\InstQueue_reg[14][1]/NET0131 ,
		\InstQueue_reg[4][1]/NET0131 ,
		_w453_,
		_w458_,
		_w3805_
	);
	LUT4 #(
		.INIT('h8000)
	) name3353 (
		_w3804_,
		_w3805_,
		_w3802_,
		_w3803_,
		_w3806_
	);
	LUT2 #(
		.INIT('h8)
	) name3354 (
		_w3801_,
		_w3806_,
		_w3807_
	);
	LUT4 #(
		.INIT('h0080)
	) name3355 (
		_w576_,
		_w579_,
		_w605_,
		_w3807_,
		_w3808_
	);
	LUT3 #(
		.INIT('h80)
	) name3356 (
		\Datai[17]_pad ,
		_w514_,
		_w569_,
		_w3809_
	);
	LUT2 #(
		.INIT('h8)
	) name3357 (
		\Datai[1]_pad ,
		_w566_,
		_w3810_
	);
	LUT4 #(
		.INIT('h1113)
	) name3358 (
		_w612_,
		_w3808_,
		_w3809_,
		_w3810_,
		_w3811_
	);
	LUT4 #(
		.INIT('h7500)
	) name3359 (
		\EAX_reg[17]/NET0131 ,
		_w635_,
		_w1852_,
		_w3811_,
		_w3812_
	);
	LUT2 #(
		.INIT('h2)
	) name3360 (
		\EAX_reg[17]/NET0131 ,
		_w1825_,
		_w3813_
	);
	LUT4 #(
		.INIT('hff8a)
	) name3361 (
		_w695_,
		_w3796_,
		_w3812_,
		_w3813_,
		_w3814_
	);
	LUT2 #(
		.INIT('h2)
	) name3362 (
		\EAX_reg[18]/NET0131 ,
		_w1825_,
		_w3815_
	);
	LUT4 #(
		.INIT('h008d)
	) name3363 (
		_w580_,
		_w605_,
		_w1850_,
		_w3795_,
		_w3816_
	);
	LUT2 #(
		.INIT('h4)
	) name3364 (
		\EAX_reg[18]/NET0131 ,
		_w1848_,
		_w3817_
	);
	LUT2 #(
		.INIT('h8)
	) name3365 (
		_w1836_,
		_w3817_,
		_w3818_
	);
	LUT4 #(
		.INIT('h3533)
	) name3366 (
		\Datai[18]_pad ,
		\EAX_reg[18]/NET0131 ,
		READY_n_pad,
		_w611_,
		_w3819_
	);
	LUT3 #(
		.INIT('h08)
	) name3367 (
		_w514_,
		_w569_,
		_w3819_,
		_w3820_
	);
	LUT4 #(
		.INIT('h153f)
	) name3368 (
		\InstQueue_reg[0][2]/NET0131 ,
		\InstQueue_reg[9][2]/NET0131 ,
		_w461_,
		_w456_,
		_w3821_
	);
	LUT4 #(
		.INIT('h135f)
	) name3369 (
		\InstQueue_reg[11][2]/NET0131 ,
		\InstQueue_reg[13][2]/NET0131 ,
		_w468_,
		_w471_,
		_w3822_
	);
	LUT4 #(
		.INIT('h153f)
	) name3370 (
		\InstQueue_reg[15][2]/NET0131 ,
		\InstQueue_reg[3][2]/NET0131 ,
		_w463_,
		_w470_,
		_w3823_
	);
	LUT4 #(
		.INIT('h153f)
	) name3371 (
		\InstQueue_reg[10][2]/NET0131 ,
		\InstQueue_reg[2][2]/NET0131 ,
		_w473_,
		_w477_,
		_w3824_
	);
	LUT4 #(
		.INIT('h8000)
	) name3372 (
		_w3823_,
		_w3824_,
		_w3821_,
		_w3822_,
		_w3825_
	);
	LUT4 #(
		.INIT('h135f)
	) name3373 (
		\InstQueue_reg[12][2]/NET0131 ,
		\InstQueue_reg[5][2]/NET0131 ,
		_w454_,
		_w474_,
		_w3826_
	);
	LUT4 #(
		.INIT('h135f)
	) name3374 (
		\InstQueue_reg[4][2]/NET0131 ,
		\InstQueue_reg[8][2]/NET0131 ,
		_w453_,
		_w467_,
		_w3827_
	);
	LUT4 #(
		.INIT('h135f)
	) name3375 (
		\InstQueue_reg[1][2]/NET0131 ,
		\InstQueue_reg[6][2]/NET0131 ,
		_w460_,
		_w476_,
		_w3828_
	);
	LUT4 #(
		.INIT('h153f)
	) name3376 (
		\InstQueue_reg[14][2]/NET0131 ,
		\InstQueue_reg[7][2]/NET0131 ,
		_w464_,
		_w458_,
		_w3829_
	);
	LUT4 #(
		.INIT('h8000)
	) name3377 (
		_w3828_,
		_w3829_,
		_w3826_,
		_w3827_,
		_w3830_
	);
	LUT2 #(
		.INIT('h8)
	) name3378 (
		_w3825_,
		_w3830_,
		_w3831_
	);
	LUT4 #(
		.INIT('h0080)
	) name3379 (
		_w576_,
		_w579_,
		_w605_,
		_w3831_,
		_w3832_
	);
	LUT4 #(
		.INIT('h3533)
	) name3380 (
		\Datai[2]_pad ,
		\EAX_reg[18]/NET0131 ,
		READY_n_pad,
		_w611_,
		_w3833_
	);
	LUT2 #(
		.INIT('h2)
	) name3381 (
		_w566_,
		_w3833_,
		_w3834_
	);
	LUT3 #(
		.INIT('h01)
	) name3382 (
		_w3832_,
		_w3834_,
		_w3820_,
		_w3835_
	);
	LUT4 #(
		.INIT('h0d00)
	) name3383 (
		\EAX_reg[18]/NET0131 ,
		_w3816_,
		_w3818_,
		_w3835_,
		_w3836_
	);
	LUT3 #(
		.INIT('hce)
	) name3384 (
		_w695_,
		_w3815_,
		_w3836_,
		_w3837_
	);
	LUT3 #(
		.INIT('h48)
	) name3385 (
		\EAX_reg[19]/NET0131 ,
		_w1848_,
		_w1837_,
		_w3838_
	);
	LUT4 #(
		.INIT('h135f)
	) name3386 (
		\InstQueue_reg[1][3]/NET0131 ,
		\InstQueue_reg[6][3]/NET0131 ,
		_w460_,
		_w476_,
		_w3839_
	);
	LUT4 #(
		.INIT('h153f)
	) name3387 (
		\InstQueue_reg[0][3]/NET0131 ,
		\InstQueue_reg[3][3]/NET0131 ,
		_w463_,
		_w456_,
		_w3840_
	);
	LUT4 #(
		.INIT('h135f)
	) name3388 (
		\InstQueue_reg[2][3]/NET0131 ,
		\InstQueue_reg[8][3]/NET0131 ,
		_w473_,
		_w467_,
		_w3841_
	);
	LUT4 #(
		.INIT('h153f)
	) name3389 (
		\InstQueue_reg[11][3]/NET0131 ,
		\InstQueue_reg[4][3]/NET0131 ,
		_w453_,
		_w468_,
		_w3842_
	);
	LUT4 #(
		.INIT('h8000)
	) name3390 (
		_w3841_,
		_w3842_,
		_w3839_,
		_w3840_,
		_w3843_
	);
	LUT4 #(
		.INIT('h135f)
	) name3391 (
		\InstQueue_reg[12][3]/NET0131 ,
		\InstQueue_reg[15][3]/NET0131 ,
		_w454_,
		_w470_,
		_w3844_
	);
	LUT4 #(
		.INIT('h153f)
	) name3392 (
		\InstQueue_reg[10][3]/NET0131 ,
		\InstQueue_reg[5][3]/NET0131 ,
		_w474_,
		_w477_,
		_w3845_
	);
	LUT4 #(
		.INIT('h153f)
	) name3393 (
		\InstQueue_reg[14][3]/NET0131 ,
		\InstQueue_reg[9][3]/NET0131 ,
		_w461_,
		_w458_,
		_w3846_
	);
	LUT4 #(
		.INIT('h153f)
	) name3394 (
		\InstQueue_reg[13][3]/NET0131 ,
		\InstQueue_reg[7][3]/NET0131 ,
		_w464_,
		_w471_,
		_w3847_
	);
	LUT4 #(
		.INIT('h8000)
	) name3395 (
		_w3846_,
		_w3847_,
		_w3844_,
		_w3845_,
		_w3848_
	);
	LUT2 #(
		.INIT('h8)
	) name3396 (
		_w3843_,
		_w3848_,
		_w3849_
	);
	LUT4 #(
		.INIT('h0080)
	) name3397 (
		_w576_,
		_w579_,
		_w605_,
		_w3849_,
		_w3850_
	);
	LUT3 #(
		.INIT('h80)
	) name3398 (
		\Datai[19]_pad ,
		_w514_,
		_w569_,
		_w3851_
	);
	LUT2 #(
		.INIT('h8)
	) name3399 (
		\Datai[3]_pad ,
		_w566_,
		_w3852_
	);
	LUT4 #(
		.INIT('h1113)
	) name3400 (
		_w612_,
		_w3850_,
		_w3851_,
		_w3852_,
		_w3853_
	);
	LUT4 #(
		.INIT('h7500)
	) name3401 (
		\EAX_reg[19]/NET0131 ,
		_w635_,
		_w1852_,
		_w3853_,
		_w3854_
	);
	LUT2 #(
		.INIT('h2)
	) name3402 (
		\EAX_reg[19]/NET0131 ,
		_w1825_,
		_w3855_
	);
	LUT4 #(
		.INIT('hff8a)
	) name3403 (
		_w695_,
		_w3838_,
		_w3854_,
		_w3855_,
		_w3856_
	);
	LUT2 #(
		.INIT('h2)
	) name3404 (
		\More_reg/NET0131 ,
		_w1825_,
		_w3857_
	);
	LUT4 #(
		.INIT('hffb0)
	) name3405 (
		_w679_,
		_w685_,
		_w695_,
		_w3857_,
		_w3858_
	);
	LUT3 #(
		.INIT('h80)
	) name3406 (
		\EAX_reg[19]/NET0131 ,
		\EAX_reg[20]/NET0131 ,
		_w1837_,
		_w3859_
	);
	LUT4 #(
		.INIT('h60c0)
	) name3407 (
		\EAX_reg[19]/NET0131 ,
		\EAX_reg[20]/NET0131 ,
		_w1848_,
		_w1837_,
		_w3860_
	);
	LUT4 #(
		.INIT('h135f)
	) name3408 (
		\InstQueue_reg[1][4]/NET0131 ,
		\InstQueue_reg[6][4]/NET0131 ,
		_w460_,
		_w476_,
		_w3861_
	);
	LUT4 #(
		.INIT('h153f)
	) name3409 (
		\InstQueue_reg[15][4]/NET0131 ,
		\InstQueue_reg[3][4]/NET0131 ,
		_w463_,
		_w470_,
		_w3862_
	);
	LUT4 #(
		.INIT('h135f)
	) name3410 (
		\InstQueue_reg[2][4]/NET0131 ,
		\InstQueue_reg[8][4]/NET0131 ,
		_w473_,
		_w467_,
		_w3863_
	);
	LUT4 #(
		.INIT('h153f)
	) name3411 (
		\InstQueue_reg[11][4]/NET0131 ,
		\InstQueue_reg[7][4]/NET0131 ,
		_w464_,
		_w468_,
		_w3864_
	);
	LUT4 #(
		.INIT('h8000)
	) name3412 (
		_w3863_,
		_w3864_,
		_w3861_,
		_w3862_,
		_w3865_
	);
	LUT4 #(
		.INIT('h153f)
	) name3413 (
		\InstQueue_reg[12][4]/NET0131 ,
		\InstQueue_reg[9][4]/NET0131 ,
		_w461_,
		_w454_,
		_w3866_
	);
	LUT4 #(
		.INIT('h153f)
	) name3414 (
		\InstQueue_reg[10][4]/NET0131 ,
		\InstQueue_reg[5][4]/NET0131 ,
		_w474_,
		_w477_,
		_w3867_
	);
	LUT4 #(
		.INIT('h135f)
	) name3415 (
		\InstQueue_reg[0][4]/NET0131 ,
		\InstQueue_reg[14][4]/NET0131 ,
		_w456_,
		_w458_,
		_w3868_
	);
	LUT4 #(
		.INIT('h153f)
	) name3416 (
		\InstQueue_reg[13][4]/NET0131 ,
		\InstQueue_reg[4][4]/NET0131 ,
		_w453_,
		_w471_,
		_w3869_
	);
	LUT4 #(
		.INIT('h8000)
	) name3417 (
		_w3868_,
		_w3869_,
		_w3866_,
		_w3867_,
		_w3870_
	);
	LUT2 #(
		.INIT('h8)
	) name3418 (
		_w3865_,
		_w3870_,
		_w3871_
	);
	LUT4 #(
		.INIT('h0080)
	) name3419 (
		_w576_,
		_w579_,
		_w605_,
		_w3871_,
		_w3872_
	);
	LUT3 #(
		.INIT('h80)
	) name3420 (
		\Datai[20]_pad ,
		_w514_,
		_w569_,
		_w3873_
	);
	LUT4 #(
		.INIT('h0507)
	) name3421 (
		_w612_,
		_w2427_,
		_w3872_,
		_w3873_,
		_w3874_
	);
	LUT4 #(
		.INIT('h7500)
	) name3422 (
		\EAX_reg[20]/NET0131 ,
		_w635_,
		_w1852_,
		_w3874_,
		_w3875_
	);
	LUT2 #(
		.INIT('h2)
	) name3423 (
		\EAX_reg[20]/NET0131 ,
		_w1825_,
		_w3876_
	);
	LUT4 #(
		.INIT('hff8a)
	) name3424 (
		_w695_,
		_w3860_,
		_w3875_,
		_w3876_,
		_w3877_
	);
	LUT4 #(
		.INIT('h8000)
	) name3425 (
		\EAX_reg[19]/NET0131 ,
		\EAX_reg[20]/NET0131 ,
		\EAX_reg[21]/NET0131 ,
		_w1837_,
		_w3878_
	);
	LUT3 #(
		.INIT('h48)
	) name3426 (
		\EAX_reg[21]/NET0131 ,
		_w1848_,
		_w3859_,
		_w3879_
	);
	LUT4 #(
		.INIT('h153f)
	) name3427 (
		\InstQueue_reg[0][5]/NET0131 ,
		\InstQueue_reg[1][5]/NET0131 ,
		_w460_,
		_w456_,
		_w3880_
	);
	LUT4 #(
		.INIT('h135f)
	) name3428 (
		\InstQueue_reg[3][5]/NET0131 ,
		\InstQueue_reg[6][5]/NET0131 ,
		_w463_,
		_w476_,
		_w3881_
	);
	LUT4 #(
		.INIT('h135f)
	) name3429 (
		\InstQueue_reg[2][5]/NET0131 ,
		\InstQueue_reg[8][5]/NET0131 ,
		_w473_,
		_w467_,
		_w3882_
	);
	LUT4 #(
		.INIT('h153f)
	) name3430 (
		\InstQueue_reg[10][5]/NET0131 ,
		\InstQueue_reg[7][5]/NET0131 ,
		_w464_,
		_w477_,
		_w3883_
	);
	LUT4 #(
		.INIT('h8000)
	) name3431 (
		_w3882_,
		_w3883_,
		_w3880_,
		_w3881_,
		_w3884_
	);
	LUT4 #(
		.INIT('h153f)
	) name3432 (
		\InstQueue_reg[13][5]/NET0131 ,
		\InstQueue_reg[5][5]/NET0131 ,
		_w474_,
		_w471_,
		_w3885_
	);
	LUT4 #(
		.INIT('h135f)
	) name3433 (
		\InstQueue_reg[11][5]/NET0131 ,
		\InstQueue_reg[15][5]/NET0131 ,
		_w468_,
		_w470_,
		_w3886_
	);
	LUT4 #(
		.INIT('h153f)
	) name3434 (
		\InstQueue_reg[14][5]/NET0131 ,
		\InstQueue_reg[4][5]/NET0131 ,
		_w453_,
		_w458_,
		_w3887_
	);
	LUT4 #(
		.INIT('h153f)
	) name3435 (
		\InstQueue_reg[12][5]/NET0131 ,
		\InstQueue_reg[9][5]/NET0131 ,
		_w461_,
		_w454_,
		_w3888_
	);
	LUT4 #(
		.INIT('h8000)
	) name3436 (
		_w3887_,
		_w3888_,
		_w3885_,
		_w3886_,
		_w3889_
	);
	LUT2 #(
		.INIT('h8)
	) name3437 (
		_w3884_,
		_w3889_,
		_w3890_
	);
	LUT4 #(
		.INIT('h0080)
	) name3438 (
		_w576_,
		_w579_,
		_w605_,
		_w3890_,
		_w3891_
	);
	LUT2 #(
		.INIT('h8)
	) name3439 (
		\Datai[5]_pad ,
		_w566_,
		_w3892_
	);
	LUT3 #(
		.INIT('h80)
	) name3440 (
		\Datai[21]_pad ,
		_w514_,
		_w569_,
		_w3893_
	);
	LUT4 #(
		.INIT('h1113)
	) name3441 (
		_w612_,
		_w3891_,
		_w3892_,
		_w3893_,
		_w3894_
	);
	LUT4 #(
		.INIT('h7500)
	) name3442 (
		\EAX_reg[21]/NET0131 ,
		_w635_,
		_w1852_,
		_w3894_,
		_w3895_
	);
	LUT2 #(
		.INIT('h2)
	) name3443 (
		\EAX_reg[21]/NET0131 ,
		_w1825_,
		_w3896_
	);
	LUT4 #(
		.INIT('hff8a)
	) name3444 (
		_w695_,
		_w3879_,
		_w3895_,
		_w3896_,
		_w3897_
	);
	LUT2 #(
		.INIT('h2)
	) name3445 (
		\EAX_reg[22]/NET0131 ,
		_w1825_,
		_w3898_
	);
	LUT4 #(
		.INIT('h5010)
	) name3446 (
		_w635_,
		_w1848_,
		_w1852_,
		_w3878_,
		_w3899_
	);
	LUT2 #(
		.INIT('h4)
	) name3447 (
		\EAX_reg[22]/NET0131 ,
		_w1848_,
		_w3900_
	);
	LUT4 #(
		.INIT('h135f)
	) name3448 (
		\InstQueue_reg[5][6]/NET0131 ,
		\InstQueue_reg[6][6]/NET0131 ,
		_w474_,
		_w476_,
		_w3901_
	);
	LUT4 #(
		.INIT('h135f)
	) name3449 (
		\InstQueue_reg[12][6]/NET0131 ,
		\InstQueue_reg[13][6]/NET0131 ,
		_w454_,
		_w471_,
		_w3902_
	);
	LUT4 #(
		.INIT('h135f)
	) name3450 (
		\InstQueue_reg[14][6]/NET0131 ,
		\InstQueue_reg[15][6]/NET0131 ,
		_w458_,
		_w470_,
		_w3903_
	);
	LUT4 #(
		.INIT('h153f)
	) name3451 (
		\InstQueue_reg[10][6]/NET0131 ,
		\InstQueue_reg[2][6]/NET0131 ,
		_w473_,
		_w477_,
		_w3904_
	);
	LUT4 #(
		.INIT('h8000)
	) name3452 (
		_w3903_,
		_w3904_,
		_w3901_,
		_w3902_,
		_w3905_
	);
	LUT4 #(
		.INIT('h135f)
	) name3453 (
		\InstQueue_reg[0][6]/NET0131 ,
		\InstQueue_reg[11][6]/NET0131 ,
		_w456_,
		_w468_,
		_w3906_
	);
	LUT4 #(
		.INIT('h135f)
	) name3454 (
		\InstQueue_reg[3][6]/NET0131 ,
		\InstQueue_reg[8][6]/NET0131 ,
		_w463_,
		_w467_,
		_w3907_
	);
	LUT4 #(
		.INIT('h135f)
	) name3455 (
		\InstQueue_reg[1][6]/NET0131 ,
		\InstQueue_reg[9][6]/NET0131 ,
		_w460_,
		_w461_,
		_w3908_
	);
	LUT4 #(
		.INIT('h153f)
	) name3456 (
		\InstQueue_reg[4][6]/NET0131 ,
		\InstQueue_reg[7][6]/NET0131 ,
		_w464_,
		_w453_,
		_w3909_
	);
	LUT4 #(
		.INIT('h8000)
	) name3457 (
		_w3908_,
		_w3909_,
		_w3906_,
		_w3907_,
		_w3910_
	);
	LUT2 #(
		.INIT('h8)
	) name3458 (
		_w3905_,
		_w3910_,
		_w3911_
	);
	LUT4 #(
		.INIT('h0080)
	) name3459 (
		_w576_,
		_w579_,
		_w605_,
		_w3911_,
		_w3912_
	);
	LUT2 #(
		.INIT('h8)
	) name3460 (
		\Datai[6]_pad ,
		_w566_,
		_w3913_
	);
	LUT3 #(
		.INIT('h80)
	) name3461 (
		\Datai[22]_pad ,
		_w514_,
		_w569_,
		_w3914_
	);
	LUT4 #(
		.INIT('h1113)
	) name3462 (
		_w612_,
		_w3912_,
		_w3913_,
		_w3914_,
		_w3915_
	);
	LUT3 #(
		.INIT('h70)
	) name3463 (
		_w3878_,
		_w3900_,
		_w3915_,
		_w3916_
	);
	LUT4 #(
		.INIT('h08cc)
	) name3464 (
		\EAX_reg[22]/NET0131 ,
		_w695_,
		_w3899_,
		_w3916_,
		_w3917_
	);
	LUT2 #(
		.INIT('he)
	) name3465 (
		_w3898_,
		_w3917_,
		_w3918_
	);
	LUT3 #(
		.INIT('h48)
	) name3466 (
		\EAX_reg[23]/NET0131 ,
		_w1848_,
		_w1840_,
		_w3919_
	);
	LUT4 #(
		.INIT('h7888)
	) name3467 (
		_w1857_,
		_w1862_,
		_w1867_,
		_w1872_,
		_w3920_
	);
	LUT4 #(
		.INIT('h8000)
	) name3468 (
		_w576_,
		_w579_,
		_w605_,
		_w3920_,
		_w3921_
	);
	LUT3 #(
		.INIT('h80)
	) name3469 (
		\Datai[23]_pad ,
		_w514_,
		_w569_,
		_w3922_
	);
	LUT4 #(
		.INIT('h0507)
	) name3470 (
		_w612_,
		_w3718_,
		_w3921_,
		_w3922_,
		_w3923_
	);
	LUT4 #(
		.INIT('h7500)
	) name3471 (
		\EAX_reg[23]/NET0131 ,
		_w635_,
		_w1852_,
		_w3923_,
		_w3924_
	);
	LUT2 #(
		.INIT('h2)
	) name3472 (
		\EAX_reg[23]/NET0131 ,
		_w1825_,
		_w3925_
	);
	LUT4 #(
		.INIT('hff8a)
	) name3473 (
		_w695_,
		_w3919_,
		_w3924_,
		_w3925_,
		_w3926_
	);
	LUT2 #(
		.INIT('h2)
	) name3474 (
		\EAX_reg[24]/NET0131 ,
		_w1825_,
		_w3927_
	);
	LUT4 #(
		.INIT('h5010)
	) name3475 (
		_w635_,
		_w1848_,
		_w1852_,
		_w2432_,
		_w3928_
	);
	LUT2 #(
		.INIT('h4)
	) name3476 (
		\EAX_reg[24]/NET0131 ,
		_w1848_,
		_w3929_
	);
	LUT2 #(
		.INIT('h9)
	) name3477 (
		_w1873_,
		_w1884_,
		_w3930_
	);
	LUT4 #(
		.INIT('h8000)
	) name3478 (
		_w576_,
		_w579_,
		_w605_,
		_w3930_,
		_w3931_
	);
	LUT3 #(
		.INIT('h80)
	) name3479 (
		\Datai[24]_pad ,
		_w514_,
		_w569_,
		_w3932_
	);
	LUT4 #(
		.INIT('h0507)
	) name3480 (
		_w612_,
		_w2176_,
		_w3931_,
		_w3932_,
		_w3933_
	);
	LUT3 #(
		.INIT('h70)
	) name3481 (
		_w2432_,
		_w3929_,
		_w3933_,
		_w3934_
	);
	LUT4 #(
		.INIT('h08cc)
	) name3482 (
		\EAX_reg[24]/NET0131 ,
		_w695_,
		_w3928_,
		_w3934_,
		_w3935_
	);
	LUT2 #(
		.INIT('he)
	) name3483 (
		_w3927_,
		_w3935_,
		_w3936_
	);
	LUT3 #(
		.INIT('h48)
	) name3484 (
		\EAX_reg[26]/NET0131 ,
		_w570_,
		_w2050_,
		_w3937_
	);
	LUT4 #(
		.INIT('h4080)
	) name3485 (
		\EAX_reg[26]/NET0131 ,
		_w570_,
		_w659_,
		_w2050_,
		_w3938_
	);
	LUT4 #(
		.INIT('hcc08)
	) name3486 (
		\Datao[26]_pad ,
		_w695_,
		_w2422_,
		_w3938_,
		_w3939_
	);
	LUT4 #(
		.INIT('h3f15)
	) name3487 (
		\Datao[26]_pad ,
		\uWord_reg[10]/NET0131 ,
		_w696_,
		_w2159_,
		_w3940_
	);
	LUT2 #(
		.INIT('hb)
	) name3488 (
		_w3939_,
		_w3940_,
		_w3941_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name3489 (
		\uWord_reg[0]/NET0131 ,
		_w695_,
		_w1825_,
		_w2058_,
		_w3942_
	);
	LUT3 #(
		.INIT('ha6)
	) name3490 (
		\EAX_reg[16]/NET0131 ,
		\EAX_reg[31]/NET0131 ,
		_w2046_,
		_w3943_
	);
	LUT3 #(
		.INIT('h80)
	) name3491 (
		_w570_,
		_w611_,
		_w3943_,
		_w3944_
	);
	LUT3 #(
		.INIT('h80)
	) name3492 (
		\Datai[0]_pad ,
		_w566_,
		_w612_,
		_w3945_
	);
	LUT3 #(
		.INIT('ha8)
	) name3493 (
		_w695_,
		_w3944_,
		_w3945_,
		_w3946_
	);
	LUT2 #(
		.INIT('he)
	) name3494 (
		_w3942_,
		_w3946_,
		_w3947_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name3495 (
		\uWord_reg[10]/NET0131 ,
		_w695_,
		_w1825_,
		_w2058_,
		_w3948_
	);
	LUT2 #(
		.INIT('h8)
	) name3496 (
		_w566_,
		_w2032_,
		_w3949_
	);
	LUT3 #(
		.INIT('ha8)
	) name3497 (
		_w2175_,
		_w3937_,
		_w3949_,
		_w3950_
	);
	LUT2 #(
		.INIT('he)
	) name3498 (
		_w3948_,
		_w3950_,
		_w3951_
	);
	LUT2 #(
		.INIT('h2)
	) name3499 (
		\uWord_reg[13]/NET0131 ,
		_w1825_,
		_w3952_
	);
	LUT3 #(
		.INIT('h60)
	) name3500 (
		\EAX_reg[29]/NET0131 ,
		_w2052_,
		_w2149_,
		_w3953_
	);
	LUT3 #(
		.INIT('h0d)
	) name3501 (
		\uWord_reg[13]/NET0131 ,
		_w2058_,
		_w2132_,
		_w3954_
	);
	LUT4 #(
		.INIT('hecee)
	) name3502 (
		_w695_,
		_w3952_,
		_w3953_,
		_w3954_,
		_w3955_
	);
	LUT2 #(
		.INIT('h2)
	) name3503 (
		\uWord_reg[1]/NET0131 ,
		_w1825_,
		_w3956_
	);
	LUT4 #(
		.INIT('h1d3f)
	) name3504 (
		\Datai[1]_pad ,
		READY_n_pad,
		\uWord_reg[1]/NET0131 ,
		_w611_,
		_w3957_
	);
	LUT2 #(
		.INIT('h2)
	) name3505 (
		_w566_,
		_w3957_,
		_w3958_
	);
	LUT4 #(
		.INIT('h02aa)
	) name3506 (
		\uWord_reg[1]/NET0131 ,
		_w566_,
		_w570_,
		_w611_,
		_w3959_
	);
	LUT4 #(
		.INIT('hcc6c)
	) name3507 (
		\EAX_reg[16]/NET0131 ,
		\EAX_reg[17]/NET0131 ,
		\EAX_reg[31]/NET0131 ,
		_w2046_,
		_w3960_
	);
	LUT3 #(
		.INIT('h80)
	) name3508 (
		_w570_,
		_w611_,
		_w3960_,
		_w3961_
	);
	LUT4 #(
		.INIT('haaa8)
	) name3509 (
		_w695_,
		_w3959_,
		_w3958_,
		_w3961_,
		_w3962_
	);
	LUT2 #(
		.INIT('he)
	) name3510 (
		_w3956_,
		_w3962_,
		_w3963_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name3511 (
		\uWord_reg[2]/NET0131 ,
		_w695_,
		_w1825_,
		_w2058_,
		_w3964_
	);
	LUT2 #(
		.INIT('h8)
	) name3512 (
		_w566_,
		_w2669_,
		_w3965_
	);
	LUT2 #(
		.INIT('h6)
	) name3513 (
		\EAX_reg[18]/NET0131 ,
		_w2047_,
		_w3966_
	);
	LUT3 #(
		.INIT('h80)
	) name3514 (
		_w570_,
		_w611_,
		_w3966_,
		_w3967_
	);
	LUT3 #(
		.INIT('ha8)
	) name3515 (
		_w695_,
		_w3965_,
		_w3967_,
		_w3968_
	);
	LUT2 #(
		.INIT('he)
	) name3516 (
		_w3964_,
		_w3968_,
		_w3969_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name3517 (
		\uWord_reg[5]/NET0131 ,
		_w695_,
		_w1825_,
		_w2058_,
		_w3970_
	);
	LUT3 #(
		.INIT('h20)
	) name3518 (
		\Datai[5]_pad ,
		READY_n_pad,
		_w566_,
		_w3971_
	);
	LUT2 #(
		.INIT('h1)
	) name3519 (
		\EAX_reg[21]/NET0131 ,
		_w2418_,
		_w3972_
	);
	LUT4 #(
		.INIT('h8000)
	) name3520 (
		\EAX_reg[18]/NET0131 ,
		\EAX_reg[19]/NET0131 ,
		_w1838_,
		_w2047_,
		_w3973_
	);
	LUT3 #(
		.INIT('h02)
	) name3521 (
		_w570_,
		_w3973_,
		_w3972_,
		_w3974_
	);
	LUT3 #(
		.INIT('ha8)
	) name3522 (
		_w2175_,
		_w3971_,
		_w3974_,
		_w3975_
	);
	LUT2 #(
		.INIT('he)
	) name3523 (
		_w3970_,
		_w3975_,
		_w3976_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name3524 (
		\uWord_reg[6]/NET0131 ,
		_w695_,
		_w1825_,
		_w2058_,
		_w3977_
	);
	LUT3 #(
		.INIT('h20)
	) name3525 (
		\Datai[6]_pad ,
		READY_n_pad,
		_w566_,
		_w3978_
	);
	LUT2 #(
		.INIT('h1)
	) name3526 (
		\EAX_reg[22]/NET0131 ,
		_w3973_,
		_w3979_
	);
	LUT3 #(
		.INIT('h02)
	) name3527 (
		_w570_,
		_w2048_,
		_w3979_,
		_w3980_
	);
	LUT3 #(
		.INIT('ha8)
	) name3528 (
		_w2175_,
		_w3978_,
		_w3980_,
		_w3981_
	);
	LUT2 #(
		.INIT('he)
	) name3529 (
		_w3977_,
		_w3981_,
		_w3982_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name3530 (
		\uWord_reg[9]/NET0131 ,
		_w695_,
		_w1825_,
		_w2058_,
		_w3983_
	);
	LUT3 #(
		.INIT('h80)
	) name3531 (
		\Datai[9]_pad ,
		_w566_,
		_w612_,
		_w3984_
	);
	LUT4 #(
		.INIT('h4080)
	) name3532 (
		\EAX_reg[25]/NET0131 ,
		_w570_,
		_w611_,
		_w2049_,
		_w3985_
	);
	LUT3 #(
		.INIT('ha8)
	) name3533 (
		_w695_,
		_w3984_,
		_w3985_,
		_w3986_
	);
	LUT2 #(
		.INIT('he)
	) name3534 (
		_w3983_,
		_w3986_,
		_w3987_
	);
	LUT4 #(
		.INIT('h8a0a)
	) name3535 (
		\EBX_reg[0]/NET0131 ,
		_w695_,
		_w1825_,
		_w1975_,
		_w3988_
	);
	LUT2 #(
		.INIT('h4)
	) name3536 (
		\EBX_reg[0]/NET0131 ,
		_w590_,
		_w3989_
	);
	LUT4 #(
		.INIT('h0080)
	) name3537 (
		_w552_,
		_w576_,
		_w605_,
		_w792_,
		_w3990_
	);
	LUT3 #(
		.INIT('ha8)
	) name3538 (
		_w695_,
		_w3989_,
		_w3990_,
		_w3991_
	);
	LUT2 #(
		.INIT('he)
	) name3539 (
		_w3988_,
		_w3991_,
		_w3992_
	);
	LUT4 #(
		.INIT('h0080)
	) name3540 (
		_w552_,
		_w576_,
		_w605_,
		_w2784_,
		_w3993_
	);
	LUT2 #(
		.INIT('h2)
	) name3541 (
		_w590_,
		_w1963_,
		_w3994_
	);
	LUT3 #(
		.INIT('h48)
	) name3542 (
		\EBX_reg[10]/NET0131 ,
		_w590_,
		_w1962_,
		_w3995_
	);
	LUT4 #(
		.INIT('h0007)
	) name3543 (
		\EBX_reg[10]/NET0131 ,
		_w1975_,
		_w3993_,
		_w3995_,
		_w3996_
	);
	LUT2 #(
		.INIT('h2)
	) name3544 (
		\EBX_reg[10]/NET0131 ,
		_w1825_,
		_w3997_
	);
	LUT3 #(
		.INIT('hf2)
	) name3545 (
		_w695_,
		_w3996_,
		_w3997_,
		_w3998_
	);
	LUT3 #(
		.INIT('ha8)
	) name3546 (
		\EBX_reg[11]/NET0131 ,
		_w1975_,
		_w3994_,
		_w3999_
	);
	LUT4 #(
		.INIT('h0080)
	) name3547 (
		_w552_,
		_w576_,
		_w605_,
		_w2765_,
		_w4000_
	);
	LUT3 #(
		.INIT('h40)
	) name3548 (
		\EBX_reg[11]/NET0131 ,
		_w590_,
		_w1963_,
		_w4001_
	);
	LUT2 #(
		.INIT('h1)
	) name3549 (
		_w4000_,
		_w4001_,
		_w4002_
	);
	LUT2 #(
		.INIT('h2)
	) name3550 (
		\EBX_reg[11]/NET0131 ,
		_w1825_,
		_w4003_
	);
	LUT4 #(
		.INIT('hff8a)
	) name3551 (
		_w695_,
		_w3999_,
		_w4002_,
		_w4003_,
		_w4004_
	);
	LUT3 #(
		.INIT('h48)
	) name3552 (
		\EBX_reg[12]/NET0131 ,
		_w590_,
		_w1964_,
		_w4005_
	);
	LUT4 #(
		.INIT('h0080)
	) name3553 (
		_w552_,
		_w576_,
		_w605_,
		_w2805_,
		_w4006_
	);
	LUT4 #(
		.INIT('h0007)
	) name3554 (
		\EBX_reg[12]/NET0131 ,
		_w1975_,
		_w4006_,
		_w4005_,
		_w4007_
	);
	LUT2 #(
		.INIT('h2)
	) name3555 (
		\EBX_reg[12]/NET0131 ,
		_w1825_,
		_w4008_
	);
	LUT3 #(
		.INIT('hf2)
	) name3556 (
		_w695_,
		_w4007_,
		_w4008_,
		_w4009_
	);
	LUT2 #(
		.INIT('h2)
	) name3557 (
		\EBX_reg[14]/NET0131 ,
		_w1825_,
		_w4010_
	);
	LUT2 #(
		.INIT('h2)
	) name3558 (
		_w590_,
		_w1966_,
		_w4011_
	);
	LUT3 #(
		.INIT('ha8)
	) name3559 (
		\EBX_reg[14]/NET0131 ,
		_w1975_,
		_w4011_,
		_w4012_
	);
	LUT4 #(
		.INIT('h0080)
	) name3560 (
		_w552_,
		_w576_,
		_w605_,
		_w2844_,
		_w4013_
	);
	LUT3 #(
		.INIT('h40)
	) name3561 (
		\EBX_reg[14]/NET0131 ,
		_w590_,
		_w1966_,
		_w4014_
	);
	LUT2 #(
		.INIT('h1)
	) name3562 (
		_w4013_,
		_w4014_,
		_w4015_
	);
	LUT4 #(
		.INIT('hecee)
	) name3563 (
		_w695_,
		_w4010_,
		_w4012_,
		_w4015_,
		_w4016_
	);
	LUT3 #(
		.INIT('h48)
	) name3564 (
		\EBX_reg[13]/NET0131 ,
		_w590_,
		_w1965_,
		_w4017_
	);
	LUT4 #(
		.INIT('h0080)
	) name3565 (
		_w552_,
		_w576_,
		_w605_,
		_w2825_,
		_w4018_
	);
	LUT4 #(
		.INIT('h0007)
	) name3566 (
		\EBX_reg[13]/NET0131 ,
		_w1975_,
		_w4017_,
		_w4018_,
		_w4019_
	);
	LUT2 #(
		.INIT('h2)
	) name3567 (
		\EBX_reg[13]/NET0131 ,
		_w1825_,
		_w4020_
	);
	LUT3 #(
		.INIT('hf2)
	) name3568 (
		_w695_,
		_w4019_,
		_w4020_,
		_w4021_
	);
	LUT3 #(
		.INIT('h48)
	) name3569 (
		\EBX_reg[15]/NET0131 ,
		_w590_,
		_w1967_,
		_w4022_
	);
	LUT4 #(
		.INIT('h0080)
	) name3570 (
		_w552_,
		_w576_,
		_w605_,
		_w2864_,
		_w4023_
	);
	LUT4 #(
		.INIT('h0007)
	) name3571 (
		\EBX_reg[15]/NET0131 ,
		_w1975_,
		_w4023_,
		_w4022_,
		_w4024_
	);
	LUT2 #(
		.INIT('h2)
	) name3572 (
		\EBX_reg[15]/NET0131 ,
		_w1825_,
		_w4025_
	);
	LUT3 #(
		.INIT('hf2)
	) name3573 (
		_w695_,
		_w4024_,
		_w4025_,
		_w4026_
	);
	LUT3 #(
		.INIT('h48)
	) name3574 (
		\EBX_reg[16]/NET0131 ,
		_w590_,
		_w1968_,
		_w4027_
	);
	LUT4 #(
		.INIT('h0080)
	) name3575 (
		_w552_,
		_w576_,
		_w605_,
		_w3787_,
		_w4028_
	);
	LUT4 #(
		.INIT('h0007)
	) name3576 (
		\EBX_reg[16]/NET0131 ,
		_w1975_,
		_w4028_,
		_w4027_,
		_w4029_
	);
	LUT2 #(
		.INIT('h2)
	) name3577 (
		\EBX_reg[16]/NET0131 ,
		_w1825_,
		_w4030_
	);
	LUT3 #(
		.INIT('hf2)
	) name3578 (
		_w695_,
		_w4029_,
		_w4030_,
		_w4031_
	);
	LUT4 #(
		.INIT('h60c0)
	) name3579 (
		\EBX_reg[16]/NET0131 ,
		\EBX_reg[17]/NET0131 ,
		_w590_,
		_w1968_,
		_w4032_
	);
	LUT4 #(
		.INIT('h0080)
	) name3580 (
		_w552_,
		_w576_,
		_w605_,
		_w3807_,
		_w4033_
	);
	LUT4 #(
		.INIT('h0007)
	) name3581 (
		\EBX_reg[17]/NET0131 ,
		_w1975_,
		_w4033_,
		_w4032_,
		_w4034_
	);
	LUT2 #(
		.INIT('h2)
	) name3582 (
		\EBX_reg[17]/NET0131 ,
		_w1825_,
		_w4035_
	);
	LUT3 #(
		.INIT('hf2)
	) name3583 (
		_w695_,
		_w4034_,
		_w4035_,
		_w4036_
	);
	LUT3 #(
		.INIT('h48)
	) name3584 (
		\EBX_reg[18]/NET0131 ,
		_w590_,
		_w1969_,
		_w4037_
	);
	LUT4 #(
		.INIT('h0080)
	) name3585 (
		_w552_,
		_w576_,
		_w605_,
		_w3831_,
		_w4038_
	);
	LUT3 #(
		.INIT('h07)
	) name3586 (
		\EBX_reg[18]/NET0131 ,
		_w1975_,
		_w4038_,
		_w4039_
	);
	LUT2 #(
		.INIT('h2)
	) name3587 (
		\EBX_reg[18]/NET0131 ,
		_w1825_,
		_w4040_
	);
	LUT4 #(
		.INIT('hff8a)
	) name3588 (
		_w695_,
		_w4037_,
		_w4039_,
		_w4040_,
		_w4041_
	);
	LUT3 #(
		.INIT('h48)
	) name3589 (
		\EBX_reg[19]/NET0131 ,
		_w590_,
		_w2140_,
		_w4042_
	);
	LUT4 #(
		.INIT('h0080)
	) name3590 (
		_w552_,
		_w576_,
		_w605_,
		_w3849_,
		_w4043_
	);
	LUT3 #(
		.INIT('h07)
	) name3591 (
		\EBX_reg[19]/NET0131 ,
		_w1975_,
		_w4043_,
		_w4044_
	);
	LUT2 #(
		.INIT('h2)
	) name3592 (
		\EBX_reg[19]/NET0131 ,
		_w1825_,
		_w4045_
	);
	LUT4 #(
		.INIT('hff8a)
	) name3593 (
		_w695_,
		_w4042_,
		_w4044_,
		_w4045_,
		_w4046_
	);
	LUT4 #(
		.INIT('h0080)
	) name3594 (
		_w552_,
		_w576_,
		_w605_,
		_w780_,
		_w4047_
	);
	LUT2 #(
		.INIT('h8)
	) name3595 (
		_w590_,
		_w3174_,
		_w4048_
	);
	LUT4 #(
		.INIT('h0007)
	) name3596 (
		\EBX_reg[1]/NET0131 ,
		_w1975_,
		_w4047_,
		_w4048_,
		_w4049_
	);
	LUT2 #(
		.INIT('h2)
	) name3597 (
		\EBX_reg[1]/NET0131 ,
		_w1825_,
		_w4050_
	);
	LUT3 #(
		.INIT('hf2)
	) name3598 (
		_w695_,
		_w4049_,
		_w4050_,
		_w4051_
	);
	LUT3 #(
		.INIT('h13)
	) name3599 (
		\EBX_reg[19]/NET0131 ,
		\EBX_reg[20]/NET0131 ,
		_w2140_,
		_w4052_
	);
	LUT2 #(
		.INIT('h2)
	) name3600 (
		_w590_,
		_w1971_,
		_w4053_
	);
	LUT4 #(
		.INIT('h0080)
	) name3601 (
		_w552_,
		_w576_,
		_w605_,
		_w3871_,
		_w4054_
	);
	LUT3 #(
		.INIT('h07)
	) name3602 (
		\EBX_reg[20]/NET0131 ,
		_w1975_,
		_w4054_,
		_w4055_
	);
	LUT4 #(
		.INIT('h20aa)
	) name3603 (
		_w695_,
		_w4052_,
		_w4053_,
		_w4055_,
		_w4056_
	);
	LUT2 #(
		.INIT('h2)
	) name3604 (
		\EBX_reg[20]/NET0131 ,
		_w1825_,
		_w4057_
	);
	LUT2 #(
		.INIT('he)
	) name3605 (
		_w4056_,
		_w4057_,
		_w4058_
	);
	LUT3 #(
		.INIT('h48)
	) name3606 (
		\EBX_reg[21]/NET0131 ,
		_w590_,
		_w1971_,
		_w4059_
	);
	LUT4 #(
		.INIT('h0080)
	) name3607 (
		_w552_,
		_w576_,
		_w605_,
		_w3890_,
		_w4060_
	);
	LUT3 #(
		.INIT('h07)
	) name3608 (
		\EBX_reg[21]/NET0131 ,
		_w1975_,
		_w4060_,
		_w4061_
	);
	LUT2 #(
		.INIT('h2)
	) name3609 (
		\EBX_reg[21]/NET0131 ,
		_w1825_,
		_w4062_
	);
	LUT4 #(
		.INIT('hff8a)
	) name3610 (
		_w695_,
		_w4059_,
		_w4061_,
		_w4062_,
		_w4063_
	);
	LUT4 #(
		.INIT('h60c0)
	) name3611 (
		\EBX_reg[21]/NET0131 ,
		\EBX_reg[22]/NET0131 ,
		_w590_,
		_w1971_,
		_w4064_
	);
	LUT4 #(
		.INIT('h0080)
	) name3612 (
		_w552_,
		_w576_,
		_w605_,
		_w3911_,
		_w4065_
	);
	LUT3 #(
		.INIT('h07)
	) name3613 (
		\EBX_reg[22]/NET0131 ,
		_w1975_,
		_w4065_,
		_w4066_
	);
	LUT2 #(
		.INIT('h2)
	) name3614 (
		\EBX_reg[22]/NET0131 ,
		_w1825_,
		_w4067_
	);
	LUT4 #(
		.INIT('hff8a)
	) name3615 (
		_w695_,
		_w4064_,
		_w4066_,
		_w4067_,
		_w4068_
	);
	LUT4 #(
		.INIT('h4888)
	) name3616 (
		\EBX_reg[23]/NET0131 ,
		_w590_,
		_w1959_,
		_w1971_,
		_w4069_
	);
	LUT4 #(
		.INIT('h8000)
	) name3617 (
		_w552_,
		_w576_,
		_w605_,
		_w3920_,
		_w4070_
	);
	LUT3 #(
		.INIT('h07)
	) name3618 (
		\EBX_reg[23]/NET0131 ,
		_w1975_,
		_w4070_,
		_w4071_
	);
	LUT2 #(
		.INIT('h2)
	) name3619 (
		\EBX_reg[23]/NET0131 ,
		_w1825_,
		_w4072_
	);
	LUT4 #(
		.INIT('hff8a)
	) name3620 (
		_w695_,
		_w4069_,
		_w4071_,
		_w4072_,
		_w4073_
	);
	LUT4 #(
		.INIT('h8000)
	) name3621 (
		_w552_,
		_w576_,
		_w605_,
		_w3930_,
		_w4074_
	);
	LUT3 #(
		.INIT('h07)
	) name3622 (
		\EBX_reg[24]/NET0131 ,
		_w1975_,
		_w4074_,
		_w4075_
	);
	LUT4 #(
		.INIT('hb700)
	) name3623 (
		\EBX_reg[24]/NET0131 ,
		_w590_,
		_w2142_,
		_w4075_,
		_w4076_
	);
	LUT2 #(
		.INIT('h2)
	) name3624 (
		\EBX_reg[24]/NET0131 ,
		_w1825_,
		_w4077_
	);
	LUT3 #(
		.INIT('hf2)
	) name3625 (
		_w695_,
		_w4076_,
		_w4077_,
		_w4078_
	);
	LUT4 #(
		.INIT('h0080)
	) name3626 (
		_w552_,
		_w576_,
		_w605_,
		_w763_,
		_w4079_
	);
	LUT3 #(
		.INIT('h78)
	) name3627 (
		\EBX_reg[0]/NET0131 ,
		\EBX_reg[1]/NET0131 ,
		\EBX_reg[2]/NET0131 ,
		_w4080_
	);
	LUT2 #(
		.INIT('h8)
	) name3628 (
		_w590_,
		_w4080_,
		_w4081_
	);
	LUT4 #(
		.INIT('h0007)
	) name3629 (
		\EBX_reg[2]/NET0131 ,
		_w1975_,
		_w4079_,
		_w4081_,
		_w4082_
	);
	LUT2 #(
		.INIT('h2)
	) name3630 (
		\EBX_reg[2]/NET0131 ,
		_w1825_,
		_w4083_
	);
	LUT3 #(
		.INIT('hf2)
	) name3631 (
		_w695_,
		_w4082_,
		_w4083_,
		_w4084_
	);
	LUT4 #(
		.INIT('h0080)
	) name3632 (
		_w552_,
		_w576_,
		_w605_,
		_w749_,
		_w4085_
	);
	LUT4 #(
		.INIT('h7f80)
	) name3633 (
		\EBX_reg[0]/NET0131 ,
		\EBX_reg[1]/NET0131 ,
		\EBX_reg[2]/NET0131 ,
		\EBX_reg[3]/NET0131 ,
		_w4086_
	);
	LUT2 #(
		.INIT('h8)
	) name3634 (
		_w590_,
		_w4086_,
		_w4087_
	);
	LUT4 #(
		.INIT('h0007)
	) name3635 (
		\EBX_reg[3]/NET0131 ,
		_w1975_,
		_w4085_,
		_w4087_,
		_w4088_
	);
	LUT2 #(
		.INIT('h2)
	) name3636 (
		\EBX_reg[3]/NET0131 ,
		_w1825_,
		_w4089_
	);
	LUT3 #(
		.INIT('hf2)
	) name3637 (
		_w695_,
		_w4088_,
		_w4089_,
		_w4090_
	);
	LUT4 #(
		.INIT('h0080)
	) name3638 (
		_w552_,
		_w576_,
		_w605_,
		_w825_,
		_w4091_
	);
	LUT2 #(
		.INIT('h6)
	) name3639 (
		\EBX_reg[4]/NET0131 ,
		_w1960_,
		_w4092_
	);
	LUT2 #(
		.INIT('h8)
	) name3640 (
		_w590_,
		_w4092_,
		_w4093_
	);
	LUT4 #(
		.INIT('h0007)
	) name3641 (
		\EBX_reg[4]/NET0131 ,
		_w1975_,
		_w4091_,
		_w4093_,
		_w4094_
	);
	LUT2 #(
		.INIT('h2)
	) name3642 (
		\EBX_reg[4]/NET0131 ,
		_w1825_,
		_w4095_
	);
	LUT3 #(
		.INIT('hf2)
	) name3643 (
		_w695_,
		_w4094_,
		_w4095_,
		_w4096_
	);
	LUT4 #(
		.INIT('h0080)
	) name3644 (
		_w552_,
		_w576_,
		_w605_,
		_w810_,
		_w4097_
	);
	LUT3 #(
		.INIT('h6c)
	) name3645 (
		\EBX_reg[4]/NET0131 ,
		\EBX_reg[5]/NET0131 ,
		_w1960_,
		_w4098_
	);
	LUT2 #(
		.INIT('h8)
	) name3646 (
		_w590_,
		_w4098_,
		_w4099_
	);
	LUT4 #(
		.INIT('h0007)
	) name3647 (
		\EBX_reg[5]/NET0131 ,
		_w1975_,
		_w4097_,
		_w4099_,
		_w4100_
	);
	LUT2 #(
		.INIT('h2)
	) name3648 (
		\EBX_reg[5]/NET0131 ,
		_w1825_,
		_w4101_
	);
	LUT3 #(
		.INIT('hf2)
	) name3649 (
		_w695_,
		_w4100_,
		_w4101_,
		_w4102_
	);
	LUT4 #(
		.INIT('h0080)
	) name3650 (
		_w552_,
		_w576_,
		_w605_,
		_w857_,
		_w4103_
	);
	LUT4 #(
		.INIT('h78f0)
	) name3651 (
		\EBX_reg[4]/NET0131 ,
		\EBX_reg[5]/NET0131 ,
		\EBX_reg[6]/NET0131 ,
		_w1960_,
		_w4104_
	);
	LUT2 #(
		.INIT('h8)
	) name3652 (
		_w590_,
		_w4104_,
		_w4105_
	);
	LUT4 #(
		.INIT('h0007)
	) name3653 (
		\EBX_reg[6]/NET0131 ,
		_w1975_,
		_w4103_,
		_w4105_,
		_w4106_
	);
	LUT2 #(
		.INIT('h2)
	) name3654 (
		\EBX_reg[6]/NET0131 ,
		_w1825_,
		_w4107_
	);
	LUT3 #(
		.INIT('hf2)
	) name3655 (
		_w695_,
		_w4106_,
		_w4107_,
		_w4108_
	);
	LUT4 #(
		.INIT('h0080)
	) name3656 (
		_w552_,
		_w576_,
		_w605_,
		_w844_,
		_w4109_
	);
	LUT2 #(
		.INIT('h6)
	) name3657 (
		\EBX_reg[7]/NET0131 ,
		_w1961_,
		_w4110_
	);
	LUT2 #(
		.INIT('h8)
	) name3658 (
		_w590_,
		_w4110_,
		_w4111_
	);
	LUT4 #(
		.INIT('h0007)
	) name3659 (
		\EBX_reg[7]/NET0131 ,
		_w1975_,
		_w4109_,
		_w4111_,
		_w4112_
	);
	LUT2 #(
		.INIT('h2)
	) name3660 (
		\EBX_reg[7]/NET0131 ,
		_w1825_,
		_w4113_
	);
	LUT3 #(
		.INIT('hf2)
	) name3661 (
		_w695_,
		_w4112_,
		_w4113_,
		_w4114_
	);
	LUT4 #(
		.INIT('h0080)
	) name3662 (
		_w552_,
		_w576_,
		_w605_,
		_w2745_,
		_w4115_
	);
	LUT3 #(
		.INIT('h6c)
	) name3663 (
		\EBX_reg[7]/NET0131 ,
		\EBX_reg[8]/NET0131 ,
		_w1961_,
		_w4116_
	);
	LUT2 #(
		.INIT('h8)
	) name3664 (
		_w590_,
		_w4116_,
		_w4117_
	);
	LUT4 #(
		.INIT('h0007)
	) name3665 (
		\EBX_reg[8]/NET0131 ,
		_w1975_,
		_w4115_,
		_w4117_,
		_w4118_
	);
	LUT2 #(
		.INIT('h2)
	) name3666 (
		\EBX_reg[8]/NET0131 ,
		_w1825_,
		_w4119_
	);
	LUT3 #(
		.INIT('hf2)
	) name3667 (
		_w695_,
		_w4118_,
		_w4119_,
		_w4120_
	);
	LUT4 #(
		.INIT('h0080)
	) name3668 (
		_w552_,
		_w576_,
		_w605_,
		_w2727_,
		_w4121_
	);
	LUT4 #(
		.INIT('h78f0)
	) name3669 (
		\EBX_reg[7]/NET0131 ,
		\EBX_reg[8]/NET0131 ,
		\EBX_reg[9]/NET0131 ,
		_w1961_,
		_w4122_
	);
	LUT2 #(
		.INIT('h8)
	) name3670 (
		_w590_,
		_w4122_,
		_w4123_
	);
	LUT4 #(
		.INIT('h0007)
	) name3671 (
		\EBX_reg[9]/NET0131 ,
		_w1975_,
		_w4121_,
		_w4123_,
		_w4124_
	);
	LUT2 #(
		.INIT('h2)
	) name3672 (
		\EBX_reg[9]/NET0131 ,
		_w1825_,
		_w4125_
	);
	LUT3 #(
		.INIT('hf2)
	) name3673 (
		_w695_,
		_w4124_,
		_w4125_,
		_w4126_
	);
	LUT2 #(
		.INIT('h2)
	) name3674 (
		\Flush_reg/NET0131 ,
		_w1825_,
		_w4127_
	);
	LUT3 #(
		.INIT('hf4)
	) name3675 (
		_w690_,
		_w695_,
		_w4127_,
		_w4128_
	);
	LUT4 #(
		.INIT('h60c0)
	) name3676 (
		\Datai[25]_pad ,
		\Datai[26]_pad ,
		_w2187_,
		_w2196_,
		_w4129_
	);
	LUT3 #(
		.INIT('h60)
	) name3677 (
		\Datai[18]_pad ,
		_w2199_,
		_w2203_,
		_w4130_
	);
	LUT4 #(
		.INIT('h5553)
	) name3678 (
		\Datai[2]_pad ,
		\InstQueue_reg[0][2]/NET0131 ,
		_w2205_,
		_w2207_,
		_w4131_
	);
	LUT2 #(
		.INIT('h1)
	) name3679 (
		_w2211_,
		_w4131_,
		_w4132_
	);
	LUT4 #(
		.INIT('h0057)
	) name3680 (
		\DataWidth_reg[1]/NET0131 ,
		_w4129_,
		_w4130_,
		_w4132_,
		_w4133_
	);
	LUT4 #(
		.INIT('hc055)
	) name3681 (
		\InstQueue_reg[0][2]/NET0131 ,
		_w497_,
		_w502_,
		_w2205_,
		_w4134_
	);
	LUT2 #(
		.INIT('h2)
	) name3682 (
		\InstQueue_reg[0][2]/NET0131 ,
		_w2215_,
		_w4135_
	);
	LUT3 #(
		.INIT('h0d)
	) name3683 (
		_w706_,
		_w4131_,
		_w4135_,
		_w4136_
	);
	LUT3 #(
		.INIT('hd0)
	) name3684 (
		_w722_,
		_w4134_,
		_w4136_,
		_w4137_
	);
	LUT3 #(
		.INIT('h2f)
	) name3685 (
		_w700_,
		_w4133_,
		_w4137_,
		_w4138_
	);
	LUT4 #(
		.INIT('h6c00)
	) name3686 (
		\Datai[25]_pad ,
		\Datai[26]_pad ,
		_w2196_,
		_w2220_,
		_w4139_
	);
	LUT3 #(
		.INIT('h60)
	) name3687 (
		\Datai[18]_pad ,
		_w2199_,
		_w2222_,
		_w4140_
	);
	LUT4 #(
		.INIT('h5553)
	) name3688 (
		\Datai[2]_pad ,
		\InstQueue_reg[10][2]/NET0131 ,
		_w2224_,
		_w2225_,
		_w4141_
	);
	LUT2 #(
		.INIT('h1)
	) name3689 (
		_w2229_,
		_w4141_,
		_w4142_
	);
	LUT4 #(
		.INIT('h0057)
	) name3690 (
		\DataWidth_reg[1]/NET0131 ,
		_w4139_,
		_w4140_,
		_w4142_,
		_w4143_
	);
	LUT4 #(
		.INIT('hc055)
	) name3691 (
		\InstQueue_reg[10][2]/NET0131 ,
		_w497_,
		_w502_,
		_w2224_,
		_w4144_
	);
	LUT2 #(
		.INIT('h2)
	) name3692 (
		\InstQueue_reg[10][2]/NET0131 ,
		_w2215_,
		_w4145_
	);
	LUT3 #(
		.INIT('h0d)
	) name3693 (
		_w706_,
		_w4141_,
		_w4145_,
		_w4146_
	);
	LUT3 #(
		.INIT('hd0)
	) name3694 (
		_w722_,
		_w4144_,
		_w4146_,
		_w4147_
	);
	LUT3 #(
		.INIT('h2f)
	) name3695 (
		_w700_,
		_w4143_,
		_w4147_,
		_w4148_
	);
	LUT4 #(
		.INIT('h6c00)
	) name3696 (
		\Datai[25]_pad ,
		\Datai[26]_pad ,
		_w2196_,
		_w2222_,
		_w4149_
	);
	LUT3 #(
		.INIT('h60)
	) name3697 (
		\Datai[18]_pad ,
		_w2199_,
		_w2225_,
		_w4150_
	);
	LUT4 #(
		.INIT('h5553)
	) name3698 (
		\Datai[2]_pad ,
		\InstQueue_reg[11][2]/NET0131 ,
		_w2224_,
		_w2239_,
		_w4151_
	);
	LUT2 #(
		.INIT('h1)
	) name3699 (
		_w2243_,
		_w4151_,
		_w4152_
	);
	LUT4 #(
		.INIT('h0057)
	) name3700 (
		\DataWidth_reg[1]/NET0131 ,
		_w4149_,
		_w4150_,
		_w4152_,
		_w4153_
	);
	LUT4 #(
		.INIT('hc055)
	) name3701 (
		\InstQueue_reg[11][2]/NET0131 ,
		_w497_,
		_w502_,
		_w2239_,
		_w4154_
	);
	LUT2 #(
		.INIT('h2)
	) name3702 (
		\InstQueue_reg[11][2]/NET0131 ,
		_w2215_,
		_w4155_
	);
	LUT3 #(
		.INIT('h0d)
	) name3703 (
		_w706_,
		_w4151_,
		_w4155_,
		_w4156_
	);
	LUT3 #(
		.INIT('hd0)
	) name3704 (
		_w722_,
		_w4154_,
		_w4156_,
		_w4157_
	);
	LUT3 #(
		.INIT('h2f)
	) name3705 (
		_w700_,
		_w4153_,
		_w4157_,
		_w4158_
	);
	LUT4 #(
		.INIT('h6c00)
	) name3706 (
		\Datai[25]_pad ,
		\Datai[26]_pad ,
		_w2196_,
		_w2225_,
		_w4159_
	);
	LUT3 #(
		.INIT('h60)
	) name3707 (
		\Datai[18]_pad ,
		_w2199_,
		_w2224_,
		_w4160_
	);
	LUT4 #(
		.INIT('h5553)
	) name3708 (
		\Datai[2]_pad ,
		\InstQueue_reg[12][2]/NET0131 ,
		_w2239_,
		_w2253_,
		_w4161_
	);
	LUT2 #(
		.INIT('h1)
	) name3709 (
		_w2256_,
		_w4161_,
		_w4162_
	);
	LUT4 #(
		.INIT('h0057)
	) name3710 (
		\DataWidth_reg[1]/NET0131 ,
		_w4159_,
		_w4160_,
		_w4162_,
		_w4163_
	);
	LUT4 #(
		.INIT('hc055)
	) name3711 (
		\InstQueue_reg[12][2]/NET0131 ,
		_w497_,
		_w502_,
		_w2253_,
		_w4164_
	);
	LUT2 #(
		.INIT('h2)
	) name3712 (
		\InstQueue_reg[12][2]/NET0131 ,
		_w2215_,
		_w4165_
	);
	LUT3 #(
		.INIT('h0d)
	) name3713 (
		_w706_,
		_w4161_,
		_w4165_,
		_w4166_
	);
	LUT3 #(
		.INIT('hd0)
	) name3714 (
		_w722_,
		_w4164_,
		_w4166_,
		_w4167_
	);
	LUT3 #(
		.INIT('h2f)
	) name3715 (
		_w700_,
		_w4163_,
		_w4167_,
		_w4168_
	);
	LUT4 #(
		.INIT('h6c00)
	) name3716 (
		\Datai[25]_pad ,
		\Datai[26]_pad ,
		_w2196_,
		_w2224_,
		_w4169_
	);
	LUT3 #(
		.INIT('h60)
	) name3717 (
		\Datai[18]_pad ,
		_w2199_,
		_w2239_,
		_w4170_
	);
	LUT4 #(
		.INIT('h5553)
	) name3718 (
		\Datai[2]_pad ,
		\InstQueue_reg[13][2]/NET0131 ,
		_w2187_,
		_w2253_,
		_w4171_
	);
	LUT2 #(
		.INIT('h1)
	) name3719 (
		_w2268_,
		_w4171_,
		_w4172_
	);
	LUT4 #(
		.INIT('h0057)
	) name3720 (
		\DataWidth_reg[1]/NET0131 ,
		_w4169_,
		_w4170_,
		_w4172_,
		_w4173_
	);
	LUT4 #(
		.INIT('hc055)
	) name3721 (
		\InstQueue_reg[13][2]/NET0131 ,
		_w497_,
		_w502_,
		_w2187_,
		_w4174_
	);
	LUT2 #(
		.INIT('h2)
	) name3722 (
		\InstQueue_reg[13][2]/NET0131 ,
		_w2215_,
		_w4175_
	);
	LUT3 #(
		.INIT('h0d)
	) name3723 (
		_w706_,
		_w4171_,
		_w4175_,
		_w4176_
	);
	LUT3 #(
		.INIT('hd0)
	) name3724 (
		_w722_,
		_w4174_,
		_w4176_,
		_w4177_
	);
	LUT3 #(
		.INIT('h2f)
	) name3725 (
		_w700_,
		_w4173_,
		_w4177_,
		_w4178_
	);
	LUT4 #(
		.INIT('h6c00)
	) name3726 (
		\Datai[25]_pad ,
		\Datai[26]_pad ,
		_w2196_,
		_w2239_,
		_w4179_
	);
	LUT3 #(
		.INIT('h60)
	) name3727 (
		\Datai[18]_pad ,
		_w2199_,
		_w2253_,
		_w4180_
	);
	LUT4 #(
		.INIT('h5553)
	) name3728 (
		\Datai[2]_pad ,
		\InstQueue_reg[14][2]/NET0131 ,
		_w2187_,
		_w2203_,
		_w4181_
	);
	LUT2 #(
		.INIT('h1)
	) name3729 (
		_w2279_,
		_w4181_,
		_w4182_
	);
	LUT4 #(
		.INIT('h0057)
	) name3730 (
		\DataWidth_reg[1]/NET0131 ,
		_w4179_,
		_w4180_,
		_w4182_,
		_w4183_
	);
	LUT4 #(
		.INIT('hc055)
	) name3731 (
		\InstQueue_reg[14][2]/NET0131 ,
		_w497_,
		_w502_,
		_w2203_,
		_w4184_
	);
	LUT2 #(
		.INIT('h2)
	) name3732 (
		\InstQueue_reg[14][2]/NET0131 ,
		_w2215_,
		_w4185_
	);
	LUT3 #(
		.INIT('h0d)
	) name3733 (
		_w706_,
		_w4181_,
		_w4185_,
		_w4186_
	);
	LUT3 #(
		.INIT('hd0)
	) name3734 (
		_w722_,
		_w4184_,
		_w4186_,
		_w4187_
	);
	LUT3 #(
		.INIT('h2f)
	) name3735 (
		_w700_,
		_w4183_,
		_w4187_,
		_w4188_
	);
	LUT4 #(
		.INIT('h6c00)
	) name3736 (
		\Datai[25]_pad ,
		\Datai[26]_pad ,
		_w2196_,
		_w2253_,
		_w4189_
	);
	LUT3 #(
		.INIT('h48)
	) name3737 (
		\Datai[18]_pad ,
		_w2187_,
		_w2199_,
		_w4190_
	);
	LUT4 #(
		.INIT('h5553)
	) name3738 (
		\Datai[2]_pad ,
		\InstQueue_reg[15][2]/NET0131 ,
		_w2207_,
		_w2203_,
		_w4191_
	);
	LUT2 #(
		.INIT('h1)
	) name3739 (
		_w2291_,
		_w4191_,
		_w4192_
	);
	LUT4 #(
		.INIT('h0057)
	) name3740 (
		\DataWidth_reg[1]/NET0131 ,
		_w4189_,
		_w4190_,
		_w4192_,
		_w4193_
	);
	LUT4 #(
		.INIT('hc055)
	) name3741 (
		\InstQueue_reg[15][2]/NET0131 ,
		_w497_,
		_w502_,
		_w2207_,
		_w4194_
	);
	LUT2 #(
		.INIT('h2)
	) name3742 (
		\InstQueue_reg[15][2]/NET0131 ,
		_w2215_,
		_w4195_
	);
	LUT3 #(
		.INIT('h0d)
	) name3743 (
		_w706_,
		_w4191_,
		_w4195_,
		_w4196_
	);
	LUT3 #(
		.INIT('hd0)
	) name3744 (
		_w722_,
		_w4194_,
		_w4196_,
		_w4197_
	);
	LUT3 #(
		.INIT('h2f)
	) name3745 (
		_w700_,
		_w4193_,
		_w4197_,
		_w4198_
	);
	LUT4 #(
		.INIT('h6c00)
	) name3746 (
		\Datai[25]_pad ,
		\Datai[26]_pad ,
		_w2196_,
		_w2203_,
		_w4199_
	);
	LUT3 #(
		.INIT('h48)
	) name3747 (
		\Datai[18]_pad ,
		_w2207_,
		_w2199_,
		_w4200_
	);
	LUT4 #(
		.INIT('h5553)
	) name3748 (
		\Datai[2]_pad ,
		\InstQueue_reg[1][2]/NET0131 ,
		_w2205_,
		_w2301_,
		_w4201_
	);
	LUT2 #(
		.INIT('h1)
	) name3749 (
		_w2304_,
		_w4201_,
		_w4202_
	);
	LUT4 #(
		.INIT('h0057)
	) name3750 (
		\DataWidth_reg[1]/NET0131 ,
		_w4199_,
		_w4200_,
		_w4202_,
		_w4203_
	);
	LUT4 #(
		.INIT('hc055)
	) name3751 (
		\InstQueue_reg[1][2]/NET0131 ,
		_w497_,
		_w502_,
		_w2301_,
		_w4204_
	);
	LUT2 #(
		.INIT('h2)
	) name3752 (
		\InstQueue_reg[1][2]/NET0131 ,
		_w2215_,
		_w4205_
	);
	LUT3 #(
		.INIT('h0d)
	) name3753 (
		_w706_,
		_w4201_,
		_w4205_,
		_w4206_
	);
	LUT3 #(
		.INIT('hd0)
	) name3754 (
		_w722_,
		_w4204_,
		_w4206_,
		_w4207_
	);
	LUT3 #(
		.INIT('h2f)
	) name3755 (
		_w700_,
		_w4203_,
		_w4207_,
		_w4208_
	);
	LUT3 #(
		.INIT('h48)
	) name3756 (
		\Datai[18]_pad ,
		_w2205_,
		_w2199_,
		_w4209_
	);
	LUT4 #(
		.INIT('h60c0)
	) name3757 (
		\Datai[25]_pad ,
		\Datai[26]_pad ,
		_w2207_,
		_w2196_,
		_w4210_
	);
	LUT4 #(
		.INIT('h5553)
	) name3758 (
		\Datai[2]_pad ,
		\InstQueue_reg[2][2]/NET0131 ,
		_w2301_,
		_w2314_,
		_w4211_
	);
	LUT2 #(
		.INIT('h1)
	) name3759 (
		_w2317_,
		_w4211_,
		_w4212_
	);
	LUT4 #(
		.INIT('h0057)
	) name3760 (
		\DataWidth_reg[1]/NET0131 ,
		_w4209_,
		_w4210_,
		_w4212_,
		_w4213_
	);
	LUT4 #(
		.INIT('hc055)
	) name3761 (
		\InstQueue_reg[2][2]/NET0131 ,
		_w497_,
		_w502_,
		_w2314_,
		_w4214_
	);
	LUT2 #(
		.INIT('h2)
	) name3762 (
		\InstQueue_reg[2][2]/NET0131 ,
		_w2215_,
		_w4215_
	);
	LUT3 #(
		.INIT('h0d)
	) name3763 (
		_w706_,
		_w4211_,
		_w4215_,
		_w4216_
	);
	LUT3 #(
		.INIT('hd0)
	) name3764 (
		_w722_,
		_w4214_,
		_w4216_,
		_w4217_
	);
	LUT3 #(
		.INIT('h2f)
	) name3765 (
		_w700_,
		_w4213_,
		_w4217_,
		_w4218_
	);
	LUT4 #(
		.INIT('h60c0)
	) name3766 (
		\Datai[25]_pad ,
		\Datai[26]_pad ,
		_w2205_,
		_w2196_,
		_w4219_
	);
	LUT3 #(
		.INIT('h60)
	) name3767 (
		\Datai[18]_pad ,
		_w2199_,
		_w2301_,
		_w4220_
	);
	LUT4 #(
		.INIT('h5553)
	) name3768 (
		\Datai[2]_pad ,
		\InstQueue_reg[3][2]/NET0131 ,
		_w2314_,
		_w2327_,
		_w4221_
	);
	LUT2 #(
		.INIT('h1)
	) name3769 (
		_w2330_,
		_w4221_,
		_w4222_
	);
	LUT4 #(
		.INIT('h0057)
	) name3770 (
		\DataWidth_reg[1]/NET0131 ,
		_w4219_,
		_w4220_,
		_w4222_,
		_w4223_
	);
	LUT4 #(
		.INIT('hc055)
	) name3771 (
		\InstQueue_reg[3][2]/NET0131 ,
		_w497_,
		_w502_,
		_w2327_,
		_w4224_
	);
	LUT2 #(
		.INIT('h2)
	) name3772 (
		\InstQueue_reg[3][2]/NET0131 ,
		_w2215_,
		_w4225_
	);
	LUT3 #(
		.INIT('h0d)
	) name3773 (
		_w706_,
		_w4221_,
		_w4225_,
		_w4226_
	);
	LUT3 #(
		.INIT('hd0)
	) name3774 (
		_w722_,
		_w4224_,
		_w4226_,
		_w4227_
	);
	LUT3 #(
		.INIT('h2f)
	) name3775 (
		_w700_,
		_w4223_,
		_w4227_,
		_w4228_
	);
	LUT4 #(
		.INIT('h6c00)
	) name3776 (
		\Datai[25]_pad ,
		\Datai[26]_pad ,
		_w2196_,
		_w2301_,
		_w4229_
	);
	LUT3 #(
		.INIT('h60)
	) name3777 (
		\Datai[18]_pad ,
		_w2199_,
		_w2314_,
		_w4230_
	);
	LUT4 #(
		.INIT('h5553)
	) name3778 (
		\Datai[2]_pad ,
		\InstQueue_reg[4][2]/NET0131 ,
		_w2327_,
		_w2340_,
		_w4231_
	);
	LUT2 #(
		.INIT('h1)
	) name3779 (
		_w2343_,
		_w4231_,
		_w4232_
	);
	LUT4 #(
		.INIT('h0057)
	) name3780 (
		\DataWidth_reg[1]/NET0131 ,
		_w4229_,
		_w4230_,
		_w4232_,
		_w4233_
	);
	LUT4 #(
		.INIT('hc055)
	) name3781 (
		\InstQueue_reg[4][2]/NET0131 ,
		_w497_,
		_w502_,
		_w2340_,
		_w4234_
	);
	LUT2 #(
		.INIT('h2)
	) name3782 (
		\InstQueue_reg[4][2]/NET0131 ,
		_w2215_,
		_w4235_
	);
	LUT3 #(
		.INIT('h0d)
	) name3783 (
		_w706_,
		_w4231_,
		_w4235_,
		_w4236_
	);
	LUT3 #(
		.INIT('hd0)
	) name3784 (
		_w722_,
		_w4234_,
		_w4236_,
		_w4237_
	);
	LUT3 #(
		.INIT('h2f)
	) name3785 (
		_w700_,
		_w4233_,
		_w4237_,
		_w4238_
	);
	LUT4 #(
		.INIT('h6c00)
	) name3786 (
		\Datai[25]_pad ,
		\Datai[26]_pad ,
		_w2196_,
		_w2314_,
		_w4239_
	);
	LUT3 #(
		.INIT('h60)
	) name3787 (
		\Datai[18]_pad ,
		_w2199_,
		_w2327_,
		_w4240_
	);
	LUT4 #(
		.INIT('h5553)
	) name3788 (
		\Datai[2]_pad ,
		\InstQueue_reg[5][2]/NET0131 ,
		_w2340_,
		_w2353_,
		_w4241_
	);
	LUT2 #(
		.INIT('h1)
	) name3789 (
		_w2356_,
		_w4241_,
		_w4242_
	);
	LUT4 #(
		.INIT('h0057)
	) name3790 (
		\DataWidth_reg[1]/NET0131 ,
		_w4239_,
		_w4240_,
		_w4242_,
		_w4243_
	);
	LUT4 #(
		.INIT('hc055)
	) name3791 (
		\InstQueue_reg[5][2]/NET0131 ,
		_w497_,
		_w502_,
		_w2353_,
		_w4244_
	);
	LUT2 #(
		.INIT('h2)
	) name3792 (
		\InstQueue_reg[5][2]/NET0131 ,
		_w2215_,
		_w4245_
	);
	LUT3 #(
		.INIT('h0d)
	) name3793 (
		_w706_,
		_w4241_,
		_w4245_,
		_w4246_
	);
	LUT3 #(
		.INIT('hd0)
	) name3794 (
		_w722_,
		_w4244_,
		_w4246_,
		_w4247_
	);
	LUT3 #(
		.INIT('h2f)
	) name3795 (
		_w700_,
		_w4243_,
		_w4247_,
		_w4248_
	);
	LUT4 #(
		.INIT('h6c00)
	) name3796 (
		\Datai[25]_pad ,
		\Datai[26]_pad ,
		_w2196_,
		_w2327_,
		_w4249_
	);
	LUT3 #(
		.INIT('h60)
	) name3797 (
		\Datai[18]_pad ,
		_w2199_,
		_w2340_,
		_w4250_
	);
	LUT4 #(
		.INIT('h5553)
	) name3798 (
		\Datai[2]_pad ,
		\InstQueue_reg[6][2]/NET0131 ,
		_w2353_,
		_w2366_,
		_w4251_
	);
	LUT2 #(
		.INIT('h1)
	) name3799 (
		_w2369_,
		_w4251_,
		_w4252_
	);
	LUT4 #(
		.INIT('h0057)
	) name3800 (
		\DataWidth_reg[1]/NET0131 ,
		_w4249_,
		_w4250_,
		_w4252_,
		_w4253_
	);
	LUT4 #(
		.INIT('hc055)
	) name3801 (
		\InstQueue_reg[6][2]/NET0131 ,
		_w497_,
		_w502_,
		_w2366_,
		_w4254_
	);
	LUT2 #(
		.INIT('h2)
	) name3802 (
		\InstQueue_reg[6][2]/NET0131 ,
		_w2215_,
		_w4255_
	);
	LUT3 #(
		.INIT('h0d)
	) name3803 (
		_w706_,
		_w4251_,
		_w4255_,
		_w4256_
	);
	LUT3 #(
		.INIT('hd0)
	) name3804 (
		_w722_,
		_w4254_,
		_w4256_,
		_w4257_
	);
	LUT3 #(
		.INIT('h2f)
	) name3805 (
		_w700_,
		_w4253_,
		_w4257_,
		_w4258_
	);
	LUT4 #(
		.INIT('h6c00)
	) name3806 (
		\Datai[25]_pad ,
		\Datai[26]_pad ,
		_w2196_,
		_w2340_,
		_w4259_
	);
	LUT3 #(
		.INIT('h60)
	) name3807 (
		\Datai[18]_pad ,
		_w2199_,
		_w2353_,
		_w4260_
	);
	LUT4 #(
		.INIT('h5553)
	) name3808 (
		\Datai[2]_pad ,
		\InstQueue_reg[7][2]/NET0131 ,
		_w2220_,
		_w2366_,
		_w4261_
	);
	LUT2 #(
		.INIT('h1)
	) name3809 (
		_w2381_,
		_w4261_,
		_w4262_
	);
	LUT4 #(
		.INIT('h0057)
	) name3810 (
		\DataWidth_reg[1]/NET0131 ,
		_w4259_,
		_w4260_,
		_w4262_,
		_w4263_
	);
	LUT4 #(
		.INIT('hc055)
	) name3811 (
		\InstQueue_reg[7][2]/NET0131 ,
		_w497_,
		_w502_,
		_w2220_,
		_w4264_
	);
	LUT2 #(
		.INIT('h2)
	) name3812 (
		\InstQueue_reg[7][2]/NET0131 ,
		_w2215_,
		_w4265_
	);
	LUT3 #(
		.INIT('h0d)
	) name3813 (
		_w706_,
		_w4261_,
		_w4265_,
		_w4266_
	);
	LUT3 #(
		.INIT('hd0)
	) name3814 (
		_w722_,
		_w4264_,
		_w4266_,
		_w4267_
	);
	LUT3 #(
		.INIT('h2f)
	) name3815 (
		_w700_,
		_w4263_,
		_w4267_,
		_w4268_
	);
	LUT4 #(
		.INIT('h6c00)
	) name3816 (
		\Datai[25]_pad ,
		\Datai[26]_pad ,
		_w2196_,
		_w2353_,
		_w4269_
	);
	LUT3 #(
		.INIT('h60)
	) name3817 (
		\Datai[18]_pad ,
		_w2199_,
		_w2366_,
		_w4270_
	);
	LUT4 #(
		.INIT('h5553)
	) name3818 (
		\Datai[2]_pad ,
		\InstQueue_reg[8][2]/NET0131 ,
		_w2220_,
		_w2222_,
		_w4271_
	);
	LUT2 #(
		.INIT('h1)
	) name3819 (
		_w2392_,
		_w4271_,
		_w4272_
	);
	LUT4 #(
		.INIT('h0057)
	) name3820 (
		\DataWidth_reg[1]/NET0131 ,
		_w4269_,
		_w4270_,
		_w4272_,
		_w4273_
	);
	LUT4 #(
		.INIT('hc055)
	) name3821 (
		\InstQueue_reg[8][2]/NET0131 ,
		_w497_,
		_w502_,
		_w2222_,
		_w4274_
	);
	LUT2 #(
		.INIT('h2)
	) name3822 (
		\InstQueue_reg[8][2]/NET0131 ,
		_w2215_,
		_w4275_
	);
	LUT3 #(
		.INIT('h0d)
	) name3823 (
		_w706_,
		_w4271_,
		_w4275_,
		_w4276_
	);
	LUT3 #(
		.INIT('hd0)
	) name3824 (
		_w722_,
		_w4274_,
		_w4276_,
		_w4277_
	);
	LUT3 #(
		.INIT('h2f)
	) name3825 (
		_w700_,
		_w4273_,
		_w4277_,
		_w4278_
	);
	LUT4 #(
		.INIT('h6c00)
	) name3826 (
		\Datai[25]_pad ,
		\Datai[26]_pad ,
		_w2196_,
		_w2366_,
		_w4279_
	);
	LUT3 #(
		.INIT('h60)
	) name3827 (
		\Datai[18]_pad ,
		_w2199_,
		_w2220_,
		_w4280_
	);
	LUT4 #(
		.INIT('h5553)
	) name3828 (
		\Datai[2]_pad ,
		\InstQueue_reg[9][2]/NET0131 ,
		_w2225_,
		_w2222_,
		_w4281_
	);
	LUT2 #(
		.INIT('h1)
	) name3829 (
		_w2403_,
		_w4281_,
		_w4282_
	);
	LUT4 #(
		.INIT('h0057)
	) name3830 (
		\DataWidth_reg[1]/NET0131 ,
		_w4279_,
		_w4280_,
		_w4282_,
		_w4283_
	);
	LUT4 #(
		.INIT('hc055)
	) name3831 (
		\InstQueue_reg[9][2]/NET0131 ,
		_w497_,
		_w502_,
		_w2225_,
		_w4284_
	);
	LUT2 #(
		.INIT('h2)
	) name3832 (
		\InstQueue_reg[9][2]/NET0131 ,
		_w2215_,
		_w4285_
	);
	LUT3 #(
		.INIT('h0d)
	) name3833 (
		_w706_,
		_w4281_,
		_w4285_,
		_w4286_
	);
	LUT3 #(
		.INIT('hd0)
	) name3834 (
		_w722_,
		_w4284_,
		_w4286_,
		_w4287_
	);
	LUT3 #(
		.INIT('h2f)
	) name3835 (
		_w700_,
		_w4283_,
		_w4287_,
		_w4288_
	);
	LUT2 #(
		.INIT('h2)
	) name3836 (
		\Datao[29]_pad ,
		_w2422_,
		_w4289_
	);
	LUT4 #(
		.INIT('h1200)
	) name3837 (
		\EAX_reg[29]/NET0131 ,
		_w617_,
		_w2052_,
		_w2149_,
		_w4290_
	);
	LUT4 #(
		.INIT('h3f15)
	) name3838 (
		\Datao[29]_pad ,
		\uWord_reg[13]/NET0131 ,
		_w696_,
		_w2159_,
		_w4291_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name3839 (
		_w695_,
		_w4289_,
		_w4290_,
		_w4291_,
		_w4292_
	);
	LUT2 #(
		.INIT('h8)
	) name3840 (
		\CodeFetch_reg/NET0131 ,
		_w695_,
		_w4293_
	);
	LUT3 #(
		.INIT('h31)
	) name3841 (
		\CodeFetch_reg/NET0131 ,
		_w701_,
		_w1825_,
		_w4294_
	);
	LUT3 #(
		.INIT('h4f)
	) name3842 (
		_w2640_,
		_w4293_,
		_w4294_,
		_w4295_
	);
	LUT4 #(
		.INIT('h0800)
	) name3843 (
		_w570_,
		_w611_,
		_w617_,
		_w3966_,
		_w4296_
	);
	LUT4 #(
		.INIT('hcc08)
	) name3844 (
		\Datao[18]_pad ,
		_w695_,
		_w2422_,
		_w4296_,
		_w4297_
	);
	LUT4 #(
		.INIT('h3f15)
	) name3845 (
		\Datao[18]_pad ,
		\uWord_reg[2]/NET0131 ,
		_w696_,
		_w2159_,
		_w4298_
	);
	LUT2 #(
		.INIT('hb)
	) name3846 (
		_w4297_,
		_w4298_,
		_w4299_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name3847 (
		\lWord_reg[0]/NET0131 ,
		_w695_,
		_w1825_,
		_w2058_,
		_w4300_
	);
	LUT3 #(
		.INIT('h80)
	) name3848 (
		\EAX_reg[0]/NET0131 ,
		_w570_,
		_w611_,
		_w4301_
	);
	LUT3 #(
		.INIT('ha8)
	) name3849 (
		_w695_,
		_w3945_,
		_w4301_,
		_w4302_
	);
	LUT2 #(
		.INIT('he)
	) name3850 (
		_w4300_,
		_w4302_,
		_w4303_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name3851 (
		\lWord_reg[10]/NET0131 ,
		_w695_,
		_w1825_,
		_w2058_,
		_w4304_
	);
	LUT4 #(
		.INIT('h135f)
	) name3852 (
		\EAX_reg[10]/NET0131 ,
		_w566_,
		_w570_,
		_w2032_,
		_w4305_
	);
	LUT2 #(
		.INIT('h2)
	) name3853 (
		_w2175_,
		_w4305_,
		_w4306_
	);
	LUT2 #(
		.INIT('he)
	) name3854 (
		_w4304_,
		_w4306_,
		_w4307_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name3855 (
		\lWord_reg[11]/NET0131 ,
		_w695_,
		_w1825_,
		_w2058_,
		_w4308_
	);
	LUT3 #(
		.INIT('h80)
	) name3856 (
		\EAX_reg[11]/NET0131 ,
		_w570_,
		_w611_,
		_w4309_
	);
	LUT3 #(
		.INIT('ha8)
	) name3857 (
		_w695_,
		_w2678_,
		_w4309_,
		_w4310_
	);
	LUT2 #(
		.INIT('he)
	) name3858 (
		_w4308_,
		_w4310_,
		_w4311_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name3859 (
		\lWord_reg[12]/NET0131 ,
		_w695_,
		_w1825_,
		_w2058_,
		_w4312_
	);
	LUT3 #(
		.INIT('h80)
	) name3860 (
		\EAX_reg[12]/NET0131 ,
		_w570_,
		_w611_,
		_w4313_
	);
	LUT3 #(
		.INIT('h80)
	) name3861 (
		\Datai[12]_pad ,
		_w566_,
		_w612_,
		_w4314_
	);
	LUT3 #(
		.INIT('ha8)
	) name3862 (
		_w695_,
		_w4313_,
		_w4314_,
		_w4315_
	);
	LUT2 #(
		.INIT('he)
	) name3863 (
		_w4312_,
		_w4315_,
		_w4316_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name3864 (
		\lWord_reg[13]/NET0131 ,
		_w695_,
		_w1825_,
		_w2058_,
		_w4317_
	);
	LUT3 #(
		.INIT('h80)
	) name3865 (
		\EAX_reg[13]/NET0131 ,
		_w570_,
		_w611_,
		_w4318_
	);
	LUT3 #(
		.INIT('ha8)
	) name3866 (
		_w695_,
		_w2132_,
		_w4318_,
		_w4319_
	);
	LUT2 #(
		.INIT('he)
	) name3867 (
		_w4317_,
		_w4319_,
		_w4320_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name3868 (
		\lWord_reg[14]/NET0131 ,
		_w695_,
		_w1825_,
		_w2058_,
		_w4321_
	);
	LUT3 #(
		.INIT('h80)
	) name3869 (
		\EAX_reg[14]/NET0131 ,
		_w570_,
		_w611_,
		_w4322_
	);
	LUT3 #(
		.INIT('h80)
	) name3870 (
		\Datai[14]_pad ,
		_w566_,
		_w612_,
		_w4323_
	);
	LUT3 #(
		.INIT('ha8)
	) name3871 (
		_w695_,
		_w4322_,
		_w4323_,
		_w4324_
	);
	LUT2 #(
		.INIT('he)
	) name3872 (
		_w4321_,
		_w4324_,
		_w4325_
	);
	LUT4 #(
		.INIT('h1d3f)
	) name3873 (
		\Datai[15]_pad ,
		READY_n_pad,
		\lWord_reg[15]/NET0131 ,
		_w611_,
		_w4326_
	);
	LUT2 #(
		.INIT('h2)
	) name3874 (
		_w566_,
		_w4326_,
		_w4327_
	);
	LUT4 #(
		.INIT('h02aa)
	) name3875 (
		\lWord_reg[15]/NET0131 ,
		_w566_,
		_w570_,
		_w611_,
		_w4328_
	);
	LUT3 #(
		.INIT('h80)
	) name3876 (
		\EAX_reg[15]/NET0131 ,
		_w570_,
		_w611_,
		_w4329_
	);
	LUT4 #(
		.INIT('haaa8)
	) name3877 (
		_w695_,
		_w4328_,
		_w4327_,
		_w4329_,
		_w4330_
	);
	LUT2 #(
		.INIT('h2)
	) name3878 (
		\lWord_reg[15]/NET0131 ,
		_w1825_,
		_w4331_
	);
	LUT2 #(
		.INIT('he)
	) name3879 (
		_w4330_,
		_w4331_,
		_w4332_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name3880 (
		\lWord_reg[1]/NET0131 ,
		_w695_,
		_w1825_,
		_w2058_,
		_w4333_
	);
	LUT3 #(
		.INIT('h80)
	) name3881 (
		\EAX_reg[1]/NET0131 ,
		_w570_,
		_w611_,
		_w4334_
	);
	LUT2 #(
		.INIT('h8)
	) name3882 (
		_w566_,
		_w2869_,
		_w4335_
	);
	LUT3 #(
		.INIT('ha8)
	) name3883 (
		_w695_,
		_w4334_,
		_w4335_,
		_w4336_
	);
	LUT2 #(
		.INIT('he)
	) name3884 (
		_w4333_,
		_w4336_,
		_w4337_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name3885 (
		\lWord_reg[2]/NET0131 ,
		_w695_,
		_w1825_,
		_w2058_,
		_w4338_
	);
	LUT3 #(
		.INIT('h80)
	) name3886 (
		\EAX_reg[2]/NET0131 ,
		_w570_,
		_w611_,
		_w4339_
	);
	LUT3 #(
		.INIT('ha8)
	) name3887 (
		_w695_,
		_w3965_,
		_w4339_,
		_w4340_
	);
	LUT2 #(
		.INIT('he)
	) name3888 (
		_w4338_,
		_w4340_,
		_w4341_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name3889 (
		\lWord_reg[3]/NET0131 ,
		_w695_,
		_w1825_,
		_w2058_,
		_w4342_
	);
	LUT3 #(
		.INIT('h80)
	) name3890 (
		\EAX_reg[3]/NET0131 ,
		_w570_,
		_w611_,
		_w4343_
	);
	LUT2 #(
		.INIT('h8)
	) name3891 (
		_w566_,
		_w2681_,
		_w4344_
	);
	LUT3 #(
		.INIT('ha8)
	) name3892 (
		_w695_,
		_w4343_,
		_w4344_,
		_w4345_
	);
	LUT2 #(
		.INIT('he)
	) name3893 (
		_w4342_,
		_w4345_,
		_w4346_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name3894 (
		\lWord_reg[4]/NET0131 ,
		_w695_,
		_w1825_,
		_w2058_,
		_w4347_
	);
	LUT3 #(
		.INIT('h80)
	) name3895 (
		\EAX_reg[4]/NET0131 ,
		_w570_,
		_w611_,
		_w4348_
	);
	LUT3 #(
		.INIT('ha8)
	) name3896 (
		_w695_,
		_w2428_,
		_w4348_,
		_w4349_
	);
	LUT2 #(
		.INIT('he)
	) name3897 (
		_w4347_,
		_w4349_,
		_w4350_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name3898 (
		\lWord_reg[5]/NET0131 ,
		_w695_,
		_w1825_,
		_w2058_,
		_w4351_
	);
	LUT3 #(
		.INIT('h80)
	) name3899 (
		\EAX_reg[5]/NET0131 ,
		_w570_,
		_w611_,
		_w4352_
	);
	LUT3 #(
		.INIT('h80)
	) name3900 (
		\Datai[5]_pad ,
		_w566_,
		_w612_,
		_w4353_
	);
	LUT3 #(
		.INIT('ha8)
	) name3901 (
		_w695_,
		_w4352_,
		_w4353_,
		_w4354_
	);
	LUT2 #(
		.INIT('he)
	) name3902 (
		_w4351_,
		_w4354_,
		_w4355_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name3903 (
		\lWord_reg[6]/NET0131 ,
		_w695_,
		_w1825_,
		_w2058_,
		_w4356_
	);
	LUT3 #(
		.INIT('h80)
	) name3904 (
		\EAX_reg[6]/NET0131 ,
		_w570_,
		_w611_,
		_w4357_
	);
	LUT3 #(
		.INIT('h80)
	) name3905 (
		\Datai[6]_pad ,
		_w566_,
		_w612_,
		_w4358_
	);
	LUT3 #(
		.INIT('ha8)
	) name3906 (
		_w695_,
		_w4357_,
		_w4358_,
		_w4359_
	);
	LUT2 #(
		.INIT('he)
	) name3907 (
		_w4356_,
		_w4359_,
		_w4360_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name3908 (
		\lWord_reg[7]/NET0131 ,
		_w695_,
		_w1825_,
		_w2058_,
		_w4361_
	);
	LUT3 #(
		.INIT('h80)
	) name3909 (
		\EAX_reg[7]/NET0131 ,
		_w570_,
		_w611_,
		_w4362_
	);
	LUT3 #(
		.INIT('h80)
	) name3910 (
		\Datai[7]_pad ,
		_w566_,
		_w612_,
		_w4363_
	);
	LUT3 #(
		.INIT('ha8)
	) name3911 (
		_w695_,
		_w4362_,
		_w4363_,
		_w4364_
	);
	LUT2 #(
		.INIT('he)
	) name3912 (
		_w4361_,
		_w4364_,
		_w4365_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name3913 (
		\lWord_reg[8]/NET0131 ,
		_w695_,
		_w1825_,
		_w2058_,
		_w4366_
	);
	LUT3 #(
		.INIT('h80)
	) name3914 (
		\EAX_reg[8]/NET0131 ,
		_w570_,
		_w611_,
		_w4367_
	);
	LUT3 #(
		.INIT('h80)
	) name3915 (
		\Datai[8]_pad ,
		_w566_,
		_w612_,
		_w4368_
	);
	LUT3 #(
		.INIT('ha8)
	) name3916 (
		_w695_,
		_w4367_,
		_w4368_,
		_w4369_
	);
	LUT2 #(
		.INIT('he)
	) name3917 (
		_w4366_,
		_w4369_,
		_w4370_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name3918 (
		\lWord_reg[9]/NET0131 ,
		_w695_,
		_w1825_,
		_w2058_,
		_w4371_
	);
	LUT3 #(
		.INIT('h80)
	) name3919 (
		\EAX_reg[9]/NET0131 ,
		_w570_,
		_w611_,
		_w4372_
	);
	LUT3 #(
		.INIT('ha8)
	) name3920 (
		_w695_,
		_w3984_,
		_w4372_,
		_w4373_
	);
	LUT2 #(
		.INIT('he)
	) name3921 (
		_w4371_,
		_w4373_,
		_w4374_
	);
	LUT4 #(
		.INIT('h1d11)
	) name3922 (
		\InstAddrPointer_reg[29]/NET0131 ,
		_w681_,
		_w1492_,
		_w1495_,
		_w4375_
	);
	LUT3 #(
		.INIT('h2a)
	) name3923 (
		\InstAddrPointer_reg[29]/NET0131 ,
		_w624_,
		_w684_,
		_w4376_
	);
	LUT2 #(
		.INIT('h4)
	) name3924 (
		_w620_,
		_w897_,
		_w4377_
	);
	LUT2 #(
		.INIT('h8)
	) name3925 (
		_w606_,
		_w1089_,
		_w4378_
	);
	LUT4 #(
		.INIT('h00f4)
	) name3926 (
		_w582_,
		_w595_,
		_w1019_,
		_w4378_,
		_w4379_
	);
	LUT3 #(
		.INIT('h10)
	) name3927 (
		_w4377_,
		_w4376_,
		_w4379_,
		_w4380_
	);
	LUT3 #(
		.INIT('hb0)
	) name3928 (
		_w1498_,
		_w1499_,
		_w4380_,
		_w4381_
	);
	LUT4 #(
		.INIT('h08cc)
	) name3929 (
		_w574_,
		_w695_,
		_w4375_,
		_w4381_,
		_w4382_
	);
	LUT4 #(
		.INIT('h3f15)
	) name3930 (
		\InstAddrPointer_reg[29]/NET0131 ,
		\rEIP_reg[29]/NET0131 ,
		_w1109_,
		_w1110_,
		_w4383_
	);
	LUT2 #(
		.INIT('hb)
	) name3931 (
		_w4382_,
		_w4383_,
		_w4384_
	);
	LUT4 #(
		.INIT('h60c0)
	) name3932 (
		\Datai[28]_pad ,
		\Datai[29]_pad ,
		_w2187_,
		_w2197_,
		_w4385_
	);
	LUT3 #(
		.INIT('h60)
	) name3933 (
		\Datai[21]_pad ,
		_w2200_,
		_w2203_,
		_w4386_
	);
	LUT4 #(
		.INIT('h5553)
	) name3934 (
		\Datai[5]_pad ,
		\InstQueue_reg[0][5]/NET0131 ,
		_w2205_,
		_w2207_,
		_w4387_
	);
	LUT2 #(
		.INIT('h1)
	) name3935 (
		_w2211_,
		_w4387_,
		_w4388_
	);
	LUT4 #(
		.INIT('h0057)
	) name3936 (
		\DataWidth_reg[1]/NET0131 ,
		_w4385_,
		_w4386_,
		_w4388_,
		_w4389_
	);
	LUT4 #(
		.INIT('hc055)
	) name3937 (
		\InstQueue_reg[0][5]/NET0131 ,
		_w542_,
		_w547_,
		_w2205_,
		_w4390_
	);
	LUT2 #(
		.INIT('h2)
	) name3938 (
		\InstQueue_reg[0][5]/NET0131 ,
		_w2215_,
		_w4391_
	);
	LUT3 #(
		.INIT('h0d)
	) name3939 (
		_w706_,
		_w4387_,
		_w4391_,
		_w4392_
	);
	LUT3 #(
		.INIT('hd0)
	) name3940 (
		_w722_,
		_w4390_,
		_w4392_,
		_w4393_
	);
	LUT3 #(
		.INIT('h2f)
	) name3941 (
		_w700_,
		_w4389_,
		_w4393_,
		_w4394_
	);
	LUT4 #(
		.INIT('h6c00)
	) name3942 (
		\Datai[28]_pad ,
		\Datai[29]_pad ,
		_w2197_,
		_w2220_,
		_w4395_
	);
	LUT3 #(
		.INIT('h60)
	) name3943 (
		\Datai[21]_pad ,
		_w2200_,
		_w2222_,
		_w4396_
	);
	LUT4 #(
		.INIT('h5553)
	) name3944 (
		\Datai[5]_pad ,
		\InstQueue_reg[10][5]/NET0131 ,
		_w2224_,
		_w2225_,
		_w4397_
	);
	LUT2 #(
		.INIT('h1)
	) name3945 (
		_w2229_,
		_w4397_,
		_w4398_
	);
	LUT4 #(
		.INIT('h0057)
	) name3946 (
		\DataWidth_reg[1]/NET0131 ,
		_w4395_,
		_w4396_,
		_w4398_,
		_w4399_
	);
	LUT4 #(
		.INIT('hc055)
	) name3947 (
		\InstQueue_reg[10][5]/NET0131 ,
		_w542_,
		_w547_,
		_w2224_,
		_w4400_
	);
	LUT2 #(
		.INIT('h2)
	) name3948 (
		\InstQueue_reg[10][5]/NET0131 ,
		_w2215_,
		_w4401_
	);
	LUT3 #(
		.INIT('h0d)
	) name3949 (
		_w706_,
		_w4397_,
		_w4401_,
		_w4402_
	);
	LUT3 #(
		.INIT('hd0)
	) name3950 (
		_w722_,
		_w4400_,
		_w4402_,
		_w4403_
	);
	LUT3 #(
		.INIT('h2f)
	) name3951 (
		_w700_,
		_w4399_,
		_w4403_,
		_w4404_
	);
	LUT4 #(
		.INIT('h6c00)
	) name3952 (
		\Datai[28]_pad ,
		\Datai[29]_pad ,
		_w2197_,
		_w2222_,
		_w4405_
	);
	LUT3 #(
		.INIT('h60)
	) name3953 (
		\Datai[21]_pad ,
		_w2200_,
		_w2225_,
		_w4406_
	);
	LUT4 #(
		.INIT('h5553)
	) name3954 (
		\Datai[5]_pad ,
		\InstQueue_reg[11][5]/NET0131 ,
		_w2224_,
		_w2239_,
		_w4407_
	);
	LUT2 #(
		.INIT('h1)
	) name3955 (
		_w2243_,
		_w4407_,
		_w4408_
	);
	LUT4 #(
		.INIT('h0057)
	) name3956 (
		\DataWidth_reg[1]/NET0131 ,
		_w4405_,
		_w4406_,
		_w4408_,
		_w4409_
	);
	LUT4 #(
		.INIT('hc055)
	) name3957 (
		\InstQueue_reg[11][5]/NET0131 ,
		_w542_,
		_w547_,
		_w2239_,
		_w4410_
	);
	LUT2 #(
		.INIT('h2)
	) name3958 (
		\InstQueue_reg[11][5]/NET0131 ,
		_w2215_,
		_w4411_
	);
	LUT3 #(
		.INIT('h0d)
	) name3959 (
		_w706_,
		_w4407_,
		_w4411_,
		_w4412_
	);
	LUT3 #(
		.INIT('hd0)
	) name3960 (
		_w722_,
		_w4410_,
		_w4412_,
		_w4413_
	);
	LUT3 #(
		.INIT('h2f)
	) name3961 (
		_w700_,
		_w4409_,
		_w4413_,
		_w4414_
	);
	LUT4 #(
		.INIT('h6c00)
	) name3962 (
		\Datai[28]_pad ,
		\Datai[29]_pad ,
		_w2197_,
		_w2225_,
		_w4415_
	);
	LUT3 #(
		.INIT('h60)
	) name3963 (
		\Datai[21]_pad ,
		_w2200_,
		_w2224_,
		_w4416_
	);
	LUT4 #(
		.INIT('h5553)
	) name3964 (
		\Datai[5]_pad ,
		\InstQueue_reg[12][5]/NET0131 ,
		_w2239_,
		_w2253_,
		_w4417_
	);
	LUT2 #(
		.INIT('h1)
	) name3965 (
		_w2256_,
		_w4417_,
		_w4418_
	);
	LUT4 #(
		.INIT('h0057)
	) name3966 (
		\DataWidth_reg[1]/NET0131 ,
		_w4415_,
		_w4416_,
		_w4418_,
		_w4419_
	);
	LUT4 #(
		.INIT('hc055)
	) name3967 (
		\InstQueue_reg[12][5]/NET0131 ,
		_w542_,
		_w547_,
		_w2253_,
		_w4420_
	);
	LUT2 #(
		.INIT('h2)
	) name3968 (
		\InstQueue_reg[12][5]/NET0131 ,
		_w2215_,
		_w4421_
	);
	LUT3 #(
		.INIT('h0d)
	) name3969 (
		_w706_,
		_w4417_,
		_w4421_,
		_w4422_
	);
	LUT3 #(
		.INIT('hd0)
	) name3970 (
		_w722_,
		_w4420_,
		_w4422_,
		_w4423_
	);
	LUT3 #(
		.INIT('h2f)
	) name3971 (
		_w700_,
		_w4419_,
		_w4423_,
		_w4424_
	);
	LUT4 #(
		.INIT('h6c00)
	) name3972 (
		\Datai[28]_pad ,
		\Datai[29]_pad ,
		_w2197_,
		_w2224_,
		_w4425_
	);
	LUT3 #(
		.INIT('h60)
	) name3973 (
		\Datai[21]_pad ,
		_w2200_,
		_w2239_,
		_w4426_
	);
	LUT4 #(
		.INIT('h5553)
	) name3974 (
		\Datai[5]_pad ,
		\InstQueue_reg[13][5]/NET0131 ,
		_w2187_,
		_w2253_,
		_w4427_
	);
	LUT2 #(
		.INIT('h1)
	) name3975 (
		_w2268_,
		_w4427_,
		_w4428_
	);
	LUT4 #(
		.INIT('h0057)
	) name3976 (
		\DataWidth_reg[1]/NET0131 ,
		_w4425_,
		_w4426_,
		_w4428_,
		_w4429_
	);
	LUT4 #(
		.INIT('hc055)
	) name3977 (
		\InstQueue_reg[13][5]/NET0131 ,
		_w542_,
		_w547_,
		_w2187_,
		_w4430_
	);
	LUT2 #(
		.INIT('h2)
	) name3978 (
		\InstQueue_reg[13][5]/NET0131 ,
		_w2215_,
		_w4431_
	);
	LUT3 #(
		.INIT('h0d)
	) name3979 (
		_w706_,
		_w4427_,
		_w4431_,
		_w4432_
	);
	LUT3 #(
		.INIT('hd0)
	) name3980 (
		_w722_,
		_w4430_,
		_w4432_,
		_w4433_
	);
	LUT3 #(
		.INIT('h2f)
	) name3981 (
		_w700_,
		_w4429_,
		_w4433_,
		_w4434_
	);
	LUT4 #(
		.INIT('h6c00)
	) name3982 (
		\Datai[28]_pad ,
		\Datai[29]_pad ,
		_w2197_,
		_w2239_,
		_w4435_
	);
	LUT3 #(
		.INIT('h60)
	) name3983 (
		\Datai[21]_pad ,
		_w2200_,
		_w2253_,
		_w4436_
	);
	LUT4 #(
		.INIT('h5553)
	) name3984 (
		\Datai[5]_pad ,
		\InstQueue_reg[14][5]/NET0131 ,
		_w2187_,
		_w2203_,
		_w4437_
	);
	LUT2 #(
		.INIT('h1)
	) name3985 (
		_w2279_,
		_w4437_,
		_w4438_
	);
	LUT4 #(
		.INIT('h0057)
	) name3986 (
		\DataWidth_reg[1]/NET0131 ,
		_w4435_,
		_w4436_,
		_w4438_,
		_w4439_
	);
	LUT4 #(
		.INIT('hc055)
	) name3987 (
		\InstQueue_reg[14][5]/NET0131 ,
		_w542_,
		_w547_,
		_w2203_,
		_w4440_
	);
	LUT2 #(
		.INIT('h2)
	) name3988 (
		\InstQueue_reg[14][5]/NET0131 ,
		_w2215_,
		_w4441_
	);
	LUT3 #(
		.INIT('h0d)
	) name3989 (
		_w706_,
		_w4437_,
		_w4441_,
		_w4442_
	);
	LUT3 #(
		.INIT('hd0)
	) name3990 (
		_w722_,
		_w4440_,
		_w4442_,
		_w4443_
	);
	LUT3 #(
		.INIT('h2f)
	) name3991 (
		_w700_,
		_w4439_,
		_w4443_,
		_w4444_
	);
	LUT4 #(
		.INIT('h6c00)
	) name3992 (
		\Datai[28]_pad ,
		\Datai[29]_pad ,
		_w2197_,
		_w2253_,
		_w4445_
	);
	LUT3 #(
		.INIT('h48)
	) name3993 (
		\Datai[21]_pad ,
		_w2187_,
		_w2200_,
		_w4446_
	);
	LUT4 #(
		.INIT('h5553)
	) name3994 (
		\Datai[5]_pad ,
		\InstQueue_reg[15][5]/NET0131 ,
		_w2207_,
		_w2203_,
		_w4447_
	);
	LUT2 #(
		.INIT('h1)
	) name3995 (
		_w2291_,
		_w4447_,
		_w4448_
	);
	LUT4 #(
		.INIT('h0057)
	) name3996 (
		\DataWidth_reg[1]/NET0131 ,
		_w4445_,
		_w4446_,
		_w4448_,
		_w4449_
	);
	LUT4 #(
		.INIT('hc055)
	) name3997 (
		\InstQueue_reg[15][5]/NET0131 ,
		_w542_,
		_w547_,
		_w2207_,
		_w4450_
	);
	LUT2 #(
		.INIT('h2)
	) name3998 (
		\InstQueue_reg[15][5]/NET0131 ,
		_w2215_,
		_w4451_
	);
	LUT3 #(
		.INIT('h0d)
	) name3999 (
		_w706_,
		_w4447_,
		_w4451_,
		_w4452_
	);
	LUT3 #(
		.INIT('hd0)
	) name4000 (
		_w722_,
		_w4450_,
		_w4452_,
		_w4453_
	);
	LUT3 #(
		.INIT('h2f)
	) name4001 (
		_w700_,
		_w4449_,
		_w4453_,
		_w4454_
	);
	LUT4 #(
		.INIT('h6c00)
	) name4002 (
		\Datai[28]_pad ,
		\Datai[29]_pad ,
		_w2197_,
		_w2203_,
		_w4455_
	);
	LUT3 #(
		.INIT('h48)
	) name4003 (
		\Datai[21]_pad ,
		_w2207_,
		_w2200_,
		_w4456_
	);
	LUT4 #(
		.INIT('h5553)
	) name4004 (
		\Datai[5]_pad ,
		\InstQueue_reg[1][5]/NET0131 ,
		_w2205_,
		_w2301_,
		_w4457_
	);
	LUT2 #(
		.INIT('h1)
	) name4005 (
		_w2304_,
		_w4457_,
		_w4458_
	);
	LUT4 #(
		.INIT('h0057)
	) name4006 (
		\DataWidth_reg[1]/NET0131 ,
		_w4455_,
		_w4456_,
		_w4458_,
		_w4459_
	);
	LUT4 #(
		.INIT('hc055)
	) name4007 (
		\InstQueue_reg[1][5]/NET0131 ,
		_w542_,
		_w547_,
		_w2301_,
		_w4460_
	);
	LUT2 #(
		.INIT('h2)
	) name4008 (
		\InstQueue_reg[1][5]/NET0131 ,
		_w2215_,
		_w4461_
	);
	LUT3 #(
		.INIT('h0d)
	) name4009 (
		_w706_,
		_w4457_,
		_w4461_,
		_w4462_
	);
	LUT3 #(
		.INIT('hd0)
	) name4010 (
		_w722_,
		_w4460_,
		_w4462_,
		_w4463_
	);
	LUT3 #(
		.INIT('h2f)
	) name4011 (
		_w700_,
		_w4459_,
		_w4463_,
		_w4464_
	);
	LUT3 #(
		.INIT('h48)
	) name4012 (
		\Datai[21]_pad ,
		_w2205_,
		_w2200_,
		_w4465_
	);
	LUT4 #(
		.INIT('h60c0)
	) name4013 (
		\Datai[28]_pad ,
		\Datai[29]_pad ,
		_w2207_,
		_w2197_,
		_w4466_
	);
	LUT4 #(
		.INIT('h5553)
	) name4014 (
		\Datai[5]_pad ,
		\InstQueue_reg[2][5]/NET0131 ,
		_w2301_,
		_w2314_,
		_w4467_
	);
	LUT2 #(
		.INIT('h1)
	) name4015 (
		_w2317_,
		_w4467_,
		_w4468_
	);
	LUT4 #(
		.INIT('h0057)
	) name4016 (
		\DataWidth_reg[1]/NET0131 ,
		_w4465_,
		_w4466_,
		_w4468_,
		_w4469_
	);
	LUT4 #(
		.INIT('hc055)
	) name4017 (
		\InstQueue_reg[2][5]/NET0131 ,
		_w542_,
		_w547_,
		_w2314_,
		_w4470_
	);
	LUT2 #(
		.INIT('h2)
	) name4018 (
		\InstQueue_reg[2][5]/NET0131 ,
		_w2215_,
		_w4471_
	);
	LUT3 #(
		.INIT('h0d)
	) name4019 (
		_w706_,
		_w4467_,
		_w4471_,
		_w4472_
	);
	LUT3 #(
		.INIT('hd0)
	) name4020 (
		_w722_,
		_w4470_,
		_w4472_,
		_w4473_
	);
	LUT3 #(
		.INIT('h2f)
	) name4021 (
		_w700_,
		_w4469_,
		_w4473_,
		_w4474_
	);
	LUT4 #(
		.INIT('h60c0)
	) name4022 (
		\Datai[28]_pad ,
		\Datai[29]_pad ,
		_w2205_,
		_w2197_,
		_w4475_
	);
	LUT3 #(
		.INIT('h60)
	) name4023 (
		\Datai[21]_pad ,
		_w2200_,
		_w2301_,
		_w4476_
	);
	LUT4 #(
		.INIT('h5553)
	) name4024 (
		\Datai[5]_pad ,
		\InstQueue_reg[3][5]/NET0131 ,
		_w2314_,
		_w2327_,
		_w4477_
	);
	LUT2 #(
		.INIT('h1)
	) name4025 (
		_w2330_,
		_w4477_,
		_w4478_
	);
	LUT4 #(
		.INIT('h0057)
	) name4026 (
		\DataWidth_reg[1]/NET0131 ,
		_w4475_,
		_w4476_,
		_w4478_,
		_w4479_
	);
	LUT4 #(
		.INIT('hc055)
	) name4027 (
		\InstQueue_reg[3][5]/NET0131 ,
		_w542_,
		_w547_,
		_w2327_,
		_w4480_
	);
	LUT2 #(
		.INIT('h2)
	) name4028 (
		\InstQueue_reg[3][5]/NET0131 ,
		_w2215_,
		_w4481_
	);
	LUT3 #(
		.INIT('h0d)
	) name4029 (
		_w706_,
		_w4477_,
		_w4481_,
		_w4482_
	);
	LUT3 #(
		.INIT('hd0)
	) name4030 (
		_w722_,
		_w4480_,
		_w4482_,
		_w4483_
	);
	LUT3 #(
		.INIT('h2f)
	) name4031 (
		_w700_,
		_w4479_,
		_w4483_,
		_w4484_
	);
	LUT4 #(
		.INIT('h6c00)
	) name4032 (
		\Datai[28]_pad ,
		\Datai[29]_pad ,
		_w2197_,
		_w2301_,
		_w4485_
	);
	LUT3 #(
		.INIT('h60)
	) name4033 (
		\Datai[21]_pad ,
		_w2200_,
		_w2314_,
		_w4486_
	);
	LUT4 #(
		.INIT('h5553)
	) name4034 (
		\Datai[5]_pad ,
		\InstQueue_reg[4][5]/NET0131 ,
		_w2327_,
		_w2340_,
		_w4487_
	);
	LUT2 #(
		.INIT('h1)
	) name4035 (
		_w2343_,
		_w4487_,
		_w4488_
	);
	LUT4 #(
		.INIT('h0057)
	) name4036 (
		\DataWidth_reg[1]/NET0131 ,
		_w4485_,
		_w4486_,
		_w4488_,
		_w4489_
	);
	LUT4 #(
		.INIT('hc055)
	) name4037 (
		\InstQueue_reg[4][5]/NET0131 ,
		_w542_,
		_w547_,
		_w2340_,
		_w4490_
	);
	LUT2 #(
		.INIT('h2)
	) name4038 (
		\InstQueue_reg[4][5]/NET0131 ,
		_w2215_,
		_w4491_
	);
	LUT3 #(
		.INIT('h0d)
	) name4039 (
		_w706_,
		_w4487_,
		_w4491_,
		_w4492_
	);
	LUT3 #(
		.INIT('hd0)
	) name4040 (
		_w722_,
		_w4490_,
		_w4492_,
		_w4493_
	);
	LUT3 #(
		.INIT('h2f)
	) name4041 (
		_w700_,
		_w4489_,
		_w4493_,
		_w4494_
	);
	LUT4 #(
		.INIT('h6c00)
	) name4042 (
		\Datai[28]_pad ,
		\Datai[29]_pad ,
		_w2197_,
		_w2314_,
		_w4495_
	);
	LUT3 #(
		.INIT('h60)
	) name4043 (
		\Datai[21]_pad ,
		_w2200_,
		_w2327_,
		_w4496_
	);
	LUT4 #(
		.INIT('h5553)
	) name4044 (
		\Datai[5]_pad ,
		\InstQueue_reg[5][5]/NET0131 ,
		_w2340_,
		_w2353_,
		_w4497_
	);
	LUT2 #(
		.INIT('h1)
	) name4045 (
		_w2356_,
		_w4497_,
		_w4498_
	);
	LUT4 #(
		.INIT('h0057)
	) name4046 (
		\DataWidth_reg[1]/NET0131 ,
		_w4495_,
		_w4496_,
		_w4498_,
		_w4499_
	);
	LUT4 #(
		.INIT('hc055)
	) name4047 (
		\InstQueue_reg[5][5]/NET0131 ,
		_w542_,
		_w547_,
		_w2353_,
		_w4500_
	);
	LUT2 #(
		.INIT('h2)
	) name4048 (
		\InstQueue_reg[5][5]/NET0131 ,
		_w2215_,
		_w4501_
	);
	LUT3 #(
		.INIT('h0d)
	) name4049 (
		_w706_,
		_w4497_,
		_w4501_,
		_w4502_
	);
	LUT3 #(
		.INIT('hd0)
	) name4050 (
		_w722_,
		_w4500_,
		_w4502_,
		_w4503_
	);
	LUT3 #(
		.INIT('h2f)
	) name4051 (
		_w700_,
		_w4499_,
		_w4503_,
		_w4504_
	);
	LUT4 #(
		.INIT('h6c00)
	) name4052 (
		\Datai[28]_pad ,
		\Datai[29]_pad ,
		_w2197_,
		_w2327_,
		_w4505_
	);
	LUT3 #(
		.INIT('h60)
	) name4053 (
		\Datai[21]_pad ,
		_w2200_,
		_w2340_,
		_w4506_
	);
	LUT4 #(
		.INIT('h5553)
	) name4054 (
		\Datai[5]_pad ,
		\InstQueue_reg[6][5]/NET0131 ,
		_w2353_,
		_w2366_,
		_w4507_
	);
	LUT2 #(
		.INIT('h1)
	) name4055 (
		_w2369_,
		_w4507_,
		_w4508_
	);
	LUT4 #(
		.INIT('h0057)
	) name4056 (
		\DataWidth_reg[1]/NET0131 ,
		_w4505_,
		_w4506_,
		_w4508_,
		_w4509_
	);
	LUT4 #(
		.INIT('hc055)
	) name4057 (
		\InstQueue_reg[6][5]/NET0131 ,
		_w542_,
		_w547_,
		_w2366_,
		_w4510_
	);
	LUT2 #(
		.INIT('h2)
	) name4058 (
		\InstQueue_reg[6][5]/NET0131 ,
		_w2215_,
		_w4511_
	);
	LUT3 #(
		.INIT('h0d)
	) name4059 (
		_w706_,
		_w4507_,
		_w4511_,
		_w4512_
	);
	LUT3 #(
		.INIT('hd0)
	) name4060 (
		_w722_,
		_w4510_,
		_w4512_,
		_w4513_
	);
	LUT3 #(
		.INIT('h2f)
	) name4061 (
		_w700_,
		_w4509_,
		_w4513_,
		_w4514_
	);
	LUT4 #(
		.INIT('h6c00)
	) name4062 (
		\Datai[28]_pad ,
		\Datai[29]_pad ,
		_w2197_,
		_w2340_,
		_w4515_
	);
	LUT3 #(
		.INIT('h60)
	) name4063 (
		\Datai[21]_pad ,
		_w2200_,
		_w2353_,
		_w4516_
	);
	LUT4 #(
		.INIT('h5553)
	) name4064 (
		\Datai[5]_pad ,
		\InstQueue_reg[7][5]/NET0131 ,
		_w2220_,
		_w2366_,
		_w4517_
	);
	LUT2 #(
		.INIT('h1)
	) name4065 (
		_w2381_,
		_w4517_,
		_w4518_
	);
	LUT4 #(
		.INIT('h0057)
	) name4066 (
		\DataWidth_reg[1]/NET0131 ,
		_w4515_,
		_w4516_,
		_w4518_,
		_w4519_
	);
	LUT4 #(
		.INIT('hc055)
	) name4067 (
		\InstQueue_reg[7][5]/NET0131 ,
		_w542_,
		_w547_,
		_w2220_,
		_w4520_
	);
	LUT2 #(
		.INIT('h2)
	) name4068 (
		\InstQueue_reg[7][5]/NET0131 ,
		_w2215_,
		_w4521_
	);
	LUT3 #(
		.INIT('h0d)
	) name4069 (
		_w706_,
		_w4517_,
		_w4521_,
		_w4522_
	);
	LUT3 #(
		.INIT('hd0)
	) name4070 (
		_w722_,
		_w4520_,
		_w4522_,
		_w4523_
	);
	LUT3 #(
		.INIT('h2f)
	) name4071 (
		_w700_,
		_w4519_,
		_w4523_,
		_w4524_
	);
	LUT4 #(
		.INIT('h6c00)
	) name4072 (
		\Datai[28]_pad ,
		\Datai[29]_pad ,
		_w2197_,
		_w2353_,
		_w4525_
	);
	LUT3 #(
		.INIT('h60)
	) name4073 (
		\Datai[21]_pad ,
		_w2200_,
		_w2366_,
		_w4526_
	);
	LUT4 #(
		.INIT('h5553)
	) name4074 (
		\Datai[5]_pad ,
		\InstQueue_reg[8][5]/NET0131 ,
		_w2220_,
		_w2222_,
		_w4527_
	);
	LUT2 #(
		.INIT('h1)
	) name4075 (
		_w2392_,
		_w4527_,
		_w4528_
	);
	LUT4 #(
		.INIT('h0057)
	) name4076 (
		\DataWidth_reg[1]/NET0131 ,
		_w4525_,
		_w4526_,
		_w4528_,
		_w4529_
	);
	LUT4 #(
		.INIT('hc055)
	) name4077 (
		\InstQueue_reg[8][5]/NET0131 ,
		_w542_,
		_w547_,
		_w2222_,
		_w4530_
	);
	LUT2 #(
		.INIT('h2)
	) name4078 (
		\InstQueue_reg[8][5]/NET0131 ,
		_w2215_,
		_w4531_
	);
	LUT3 #(
		.INIT('h0d)
	) name4079 (
		_w706_,
		_w4527_,
		_w4531_,
		_w4532_
	);
	LUT3 #(
		.INIT('hd0)
	) name4080 (
		_w722_,
		_w4530_,
		_w4532_,
		_w4533_
	);
	LUT3 #(
		.INIT('h2f)
	) name4081 (
		_w700_,
		_w4529_,
		_w4533_,
		_w4534_
	);
	LUT4 #(
		.INIT('h6c00)
	) name4082 (
		\Datai[28]_pad ,
		\Datai[29]_pad ,
		_w2197_,
		_w2366_,
		_w4535_
	);
	LUT3 #(
		.INIT('h60)
	) name4083 (
		\Datai[21]_pad ,
		_w2200_,
		_w2220_,
		_w4536_
	);
	LUT4 #(
		.INIT('h5553)
	) name4084 (
		\Datai[5]_pad ,
		\InstQueue_reg[9][5]/NET0131 ,
		_w2225_,
		_w2222_,
		_w4537_
	);
	LUT2 #(
		.INIT('h1)
	) name4085 (
		_w2403_,
		_w4537_,
		_w4538_
	);
	LUT4 #(
		.INIT('h0057)
	) name4086 (
		\DataWidth_reg[1]/NET0131 ,
		_w4535_,
		_w4536_,
		_w4538_,
		_w4539_
	);
	LUT4 #(
		.INIT('hc055)
	) name4087 (
		\InstQueue_reg[9][5]/NET0131 ,
		_w542_,
		_w547_,
		_w2225_,
		_w4540_
	);
	LUT2 #(
		.INIT('h2)
	) name4088 (
		\InstQueue_reg[9][5]/NET0131 ,
		_w2215_,
		_w4541_
	);
	LUT3 #(
		.INIT('h0d)
	) name4089 (
		_w706_,
		_w4537_,
		_w4541_,
		_w4542_
	);
	LUT3 #(
		.INIT('hd0)
	) name4090 (
		_w722_,
		_w4540_,
		_w4542_,
		_w4543_
	);
	LUT3 #(
		.INIT('h2f)
	) name4091 (
		_w700_,
		_w4539_,
		_w4543_,
		_w4544_
	);
	LUT2 #(
		.INIT('he)
	) name4092 (
		\rEIP_reg[0]/NET0131 ,
		\rEIP_reg[1]/NET0131 ,
		_w4545_
	);
	LUT3 #(
		.INIT('he0)
	) name4093 (
		\rEIP_reg[0]/NET0131 ,
		\rEIP_reg[1]/NET0131 ,
		\rEIP_reg[31]/NET0131 ,
		_w4546_
	);
	LUT4 #(
		.INIT('he000)
	) name4094 (
		\rEIP_reg[0]/NET0131 ,
		\rEIP_reg[1]/NET0131 ,
		\rEIP_reg[2]/NET0131 ,
		\rEIP_reg[31]/NET0131 ,
		_w4547_
	);
	LUT3 #(
		.INIT('h80)
	) name4095 (
		\rEIP_reg[3]/NET0131 ,
		\rEIP_reg[4]/NET0131 ,
		_w4547_,
		_w4548_
	);
	LUT4 #(
		.INIT('h8000)
	) name4096 (
		\rEIP_reg[3]/NET0131 ,
		\rEIP_reg[4]/NET0131 ,
		\rEIP_reg[5]/NET0131 ,
		_w4547_,
		_w4549_
	);
	LUT3 #(
		.INIT('h80)
	) name4097 (
		\rEIP_reg[6]/NET0131 ,
		\rEIP_reg[7]/NET0131 ,
		_w4549_,
		_w4550_
	);
	LUT4 #(
		.INIT('h8000)
	) name4098 (
		\rEIP_reg[6]/NET0131 ,
		\rEIP_reg[7]/NET0131 ,
		\rEIP_reg[8]/NET0131 ,
		_w4549_,
		_w4551_
	);
	LUT3 #(
		.INIT('h80)
	) name4099 (
		\rEIP_reg[10]/NET0131 ,
		\rEIP_reg[9]/NET0131 ,
		_w4551_,
		_w4552_
	);
	LUT4 #(
		.INIT('h8000)
	) name4100 (
		\rEIP_reg[10]/NET0131 ,
		\rEIP_reg[11]/NET0131 ,
		\rEIP_reg[9]/NET0131 ,
		_w4551_,
		_w4553_
	);
	LUT3 #(
		.INIT('h80)
	) name4101 (
		\rEIP_reg[12]/NET0131 ,
		\rEIP_reg[13]/NET0131 ,
		_w4553_,
		_w4554_
	);
	LUT4 #(
		.INIT('h8000)
	) name4102 (
		\rEIP_reg[12]/NET0131 ,
		\rEIP_reg[13]/NET0131 ,
		\rEIP_reg[14]/NET0131 ,
		_w4553_,
		_w4555_
	);
	LUT3 #(
		.INIT('h80)
	) name4103 (
		\rEIP_reg[15]/NET0131 ,
		\rEIP_reg[16]/NET0131 ,
		_w4555_,
		_w4556_
	);
	LUT4 #(
		.INIT('h8000)
	) name4104 (
		\rEIP_reg[15]/NET0131 ,
		\rEIP_reg[16]/NET0131 ,
		_w2615_,
		_w4555_,
		_w4557_
	);
	LUT3 #(
		.INIT('h80)
	) name4105 (
		_w2605_,
		_w2617_,
		_w4557_,
		_w4558_
	);
	LUT4 #(
		.INIT('h8000)
	) name4106 (
		\rEIP_reg[26]/NET0131 ,
		_w2605_,
		_w2617_,
		_w4557_,
		_w4559_
	);
	LUT4 #(
		.INIT('h4888)
	) name4107 (
		\rEIP_reg[30]/NET0131 ,
		_w615_,
		_w2621_,
		_w4559_,
		_w4560_
	);
	LUT3 #(
		.INIT('h8a)
	) name4108 (
		\Address[28]_pad ,
		\State_reg[0]/NET0131 ,
		\State_reg[1]/NET0131 ,
		_w4561_
	);
	LUT2 #(
		.INIT('h8)
	) name4109 (
		\rEIP_reg[0]/NET0131 ,
		\rEIP_reg[31]/NET0131 ,
		_w4562_
	);
	LUT4 #(
		.INIT('h8000)
	) name4110 (
		_w2605_,
		_w2611_,
		_w2615_,
		_w4562_,
		_w4563_
	);
	LUT4 #(
		.INIT('h1555)
	) name4111 (
		\rEIP_reg[29]/NET0131 ,
		_w2618_,
		_w2620_,
		_w4563_,
		_w4564_
	);
	LUT3 #(
		.INIT('h40)
	) name4112 (
		\State_reg[0]/NET0131 ,
		\State_reg[1]/NET0131 ,
		\State_reg[2]/NET0131 ,
		_w4565_
	);
	LUT4 #(
		.INIT('h70f0)
	) name4113 (
		_w2618_,
		_w2621_,
		_w4565_,
		_w4563_,
		_w4566_
	);
	LUT3 #(
		.INIT('h45)
	) name4114 (
		_w4561_,
		_w4564_,
		_w4566_,
		_w4567_
	);
	LUT2 #(
		.INIT('hb)
	) name4115 (
		_w4560_,
		_w4567_,
		_w4568_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name4116 (
		\Datao[25]_pad ,
		_w617_,
		_w2422_,
		_w3985_,
		_w4569_
	);
	LUT4 #(
		.INIT('h3f15)
	) name4117 (
		\Datao[25]_pad ,
		\uWord_reg[9]/NET0131 ,
		_w696_,
		_w2159_,
		_w4570_
	);
	LUT3 #(
		.INIT('h2f)
	) name4118 (
		_w695_,
		_w4569_,
		_w4570_,
		_w4571_
	);
	LUT2 #(
		.INIT('h1)
	) name4119 (
		_w617_,
		_w3960_,
		_w4572_
	);
	LUT3 #(
		.INIT('h08)
	) name4120 (
		_w570_,
		_w611_,
		_w4572_,
		_w4573_
	);
	LUT4 #(
		.INIT('haaa2)
	) name4121 (
		\Datao[17]_pad ,
		_w2153_,
		_w2154_,
		_w4573_,
		_w4574_
	);
	LUT4 #(
		.INIT('h0800)
	) name4122 (
		_w570_,
		_w611_,
		_w617_,
		_w3960_,
		_w4575_
	);
	LUT4 #(
		.INIT('h3f15)
	) name4123 (
		\Datao[17]_pad ,
		\uWord_reg[1]/NET0131 ,
		_w696_,
		_w2159_,
		_w4576_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name4124 (
		_w695_,
		_w4574_,
		_w4575_,
		_w4576_,
		_w4577_
	);
	LUT4 #(
		.INIT('h0509)
	) name4125 (
		\EAX_reg[16]/NET0131 ,
		\EAX_reg[31]/NET0131 ,
		_w617_,
		_w2046_,
		_w4578_
	);
	LUT3 #(
		.INIT('h08)
	) name4126 (
		_w570_,
		_w611_,
		_w4578_,
		_w4579_
	);
	LUT4 #(
		.INIT('haaa2)
	) name4127 (
		\Datao[16]_pad ,
		_w2153_,
		_w2154_,
		_w4579_,
		_w4580_
	);
	LUT4 #(
		.INIT('h0800)
	) name4128 (
		_w570_,
		_w611_,
		_w617_,
		_w3943_,
		_w4581_
	);
	LUT4 #(
		.INIT('h3f15)
	) name4129 (
		\Datao[16]_pad ,
		\uWord_reg[0]/NET0131 ,
		_w696_,
		_w2159_,
		_w4582_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name4130 (
		_w695_,
		_w4580_,
		_w4581_,
		_w4582_,
		_w4583_
	);
	LUT4 #(
		.INIT('h0008)
	) name4131 (
		_w570_,
		_w659_,
		_w3973_,
		_w3972_,
		_w4584_
	);
	LUT4 #(
		.INIT('hcc08)
	) name4132 (
		\Datao[21]_pad ,
		_w695_,
		_w2422_,
		_w4584_,
		_w4585_
	);
	LUT4 #(
		.INIT('h3f15)
	) name4133 (
		\Datao[21]_pad ,
		\uWord_reg[5]/NET0131 ,
		_w696_,
		_w2159_,
		_w4586_
	);
	LUT2 #(
		.INIT('hb)
	) name4134 (
		_w4585_,
		_w4586_,
		_w4587_
	);
	LUT4 #(
		.INIT('h1050)
	) name4135 (
		\Flush_reg/NET0131 ,
		\InstQueueRd_Addr_reg[2]/NET0131 ,
		_w712_,
		_w714_,
		_w4588_
	);
	LUT4 #(
		.INIT('hfd9f)
	) name4136 (
		\State2_reg[0]/NET0131 ,
		\State2_reg[1]/NET0131 ,
		\State2_reg[2]/NET0131 ,
		\State2_reg[3]/NET0131 ,
		_w4589_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name4137 (
		\InstQueueWr_Addr_reg[2]/NET0131 ,
		_w3691_,
		_w4588_,
		_w4589_,
		_w4590_
	);
	LUT4 #(
		.INIT('hcc08)
	) name4138 (
		\DataWidth_reg[1]/NET0131 ,
		\InstQueueWr_Addr_reg[2]/NET0131 ,
		_w706_,
		_w2202_,
		_w4591_
	);
	LUT3 #(
		.INIT('h54)
	) name4139 (
		_w722_,
		_w1280_,
		_w4591_,
		_w4592_
	);
	LUT2 #(
		.INIT('h4)
	) name4140 (
		_w1280_,
		_w2202_,
		_w4593_
	);
	LUT3 #(
		.INIT('h07)
	) name4141 (
		\InstQueueWr_Addr_reg[0]/NET0131 ,
		\InstQueueWr_Addr_reg[1]/NET0131 ,
		\InstQueueWr_Addr_reg[2]/NET0131 ,
		_w4594_
	);
	LUT3 #(
		.INIT('h70)
	) name4142 (
		\DataWidth_reg[1]/NET0131 ,
		_w700_,
		_w4594_,
		_w4595_
	);
	LUT3 #(
		.INIT('h45)
	) name4143 (
		_w2206_,
		_w4593_,
		_w4595_,
		_w4596_
	);
	LUT3 #(
		.INIT('hba)
	) name4144 (
		_w4590_,
		_w4592_,
		_w4596_,
		_w4597_
	);
	LUT4 #(
		.INIT('h8000)
	) name4145 (
		\rEIP_reg[15]/NET0131 ,
		\rEIP_reg[16]/NET0131 ,
		_w2612_,
		_w4555_,
		_w4598_
	);
	LUT4 #(
		.INIT('h60c0)
	) name4146 (
		\rEIP_reg[17]/NET0131 ,
		\rEIP_reg[18]/NET0131 ,
		_w615_,
		_w4556_,
		_w4599_
	);
	LUT3 #(
		.INIT('h8a)
	) name4147 (
		\Address[16]_pad ,
		\State_reg[0]/NET0131 ,
		\State_reg[1]/NET0131 ,
		_w4600_
	);
	LUT3 #(
		.INIT('h80)
	) name4148 (
		\rEIP_reg[14]/NET0131 ,
		_w2610_,
		_w4562_,
		_w4601_
	);
	LUT4 #(
		.INIT('h8000)
	) name4149 (
		\rEIP_reg[14]/NET0131 ,
		\rEIP_reg[15]/NET0131 ,
		_w2610_,
		_w4562_,
		_w4602_
	);
	LUT3 #(
		.INIT('h80)
	) name4150 (
		\rEIP_reg[16]/NET0131 ,
		\rEIP_reg[17]/NET0131 ,
		_w4602_,
		_w4603_
	);
	LUT4 #(
		.INIT('h60c0)
	) name4151 (
		\rEIP_reg[16]/NET0131 ,
		\rEIP_reg[17]/NET0131 ,
		_w4565_,
		_w4602_,
		_w4604_
	);
	LUT2 #(
		.INIT('h1)
	) name4152 (
		_w4600_,
		_w4604_,
		_w4605_
	);
	LUT2 #(
		.INIT('hb)
	) name4153 (
		_w4599_,
		_w4605_,
		_w4606_
	);
	LUT4 #(
		.INIT('hc0a0)
	) name4154 (
		\Datao[2]_pad ,
		\EAX_reg[2]/NET0131 ,
		_w695_,
		_w2422_,
		_w4607_
	);
	LUT4 #(
		.INIT('h3f15)
	) name4155 (
		\Datao[2]_pad ,
		\lWord_reg[2]/NET0131 ,
		_w696_,
		_w2159_,
		_w4608_
	);
	LUT2 #(
		.INIT('hb)
	) name4156 (
		_w4607_,
		_w4608_,
		_w4609_
	);
	LUT4 #(
		.INIT('hc0a0)
	) name4157 (
		\Datao[3]_pad ,
		\EAX_reg[3]/NET0131 ,
		_w695_,
		_w2422_,
		_w4610_
	);
	LUT4 #(
		.INIT('h3f15)
	) name4158 (
		\Datao[3]_pad ,
		\lWord_reg[3]/NET0131 ,
		_w696_,
		_w2159_,
		_w4611_
	);
	LUT2 #(
		.INIT('hb)
	) name4159 (
		_w4610_,
		_w4611_,
		_w4612_
	);
	LUT4 #(
		.INIT('hc0a0)
	) name4160 (
		\Datao[4]_pad ,
		\EAX_reg[4]/NET0131 ,
		_w695_,
		_w2422_,
		_w4613_
	);
	LUT4 #(
		.INIT('h3f15)
	) name4161 (
		\Datao[4]_pad ,
		\lWord_reg[4]/NET0131 ,
		_w696_,
		_w2159_,
		_w4614_
	);
	LUT2 #(
		.INIT('hb)
	) name4162 (
		_w4613_,
		_w4614_,
		_w4615_
	);
	LUT4 #(
		.INIT('hc0a0)
	) name4163 (
		\Datao[5]_pad ,
		\EAX_reg[5]/NET0131 ,
		_w695_,
		_w2422_,
		_w4616_
	);
	LUT4 #(
		.INIT('h3f15)
	) name4164 (
		\Datao[5]_pad ,
		\lWord_reg[5]/NET0131 ,
		_w696_,
		_w2159_,
		_w4617_
	);
	LUT2 #(
		.INIT('hb)
	) name4165 (
		_w4616_,
		_w4617_,
		_w4618_
	);
	LUT4 #(
		.INIT('hc0a0)
	) name4166 (
		\Datao[6]_pad ,
		\EAX_reg[6]/NET0131 ,
		_w695_,
		_w2422_,
		_w4619_
	);
	LUT4 #(
		.INIT('h3f15)
	) name4167 (
		\Datao[6]_pad ,
		\lWord_reg[6]/NET0131 ,
		_w696_,
		_w2159_,
		_w4620_
	);
	LUT2 #(
		.INIT('hb)
	) name4168 (
		_w4619_,
		_w4620_,
		_w4621_
	);
	LUT4 #(
		.INIT('hc0a0)
	) name4169 (
		\Datao[7]_pad ,
		\EAX_reg[7]/NET0131 ,
		_w695_,
		_w2422_,
		_w4622_
	);
	LUT4 #(
		.INIT('h3f15)
	) name4170 (
		\Datao[7]_pad ,
		\lWord_reg[7]/NET0131 ,
		_w696_,
		_w2159_,
		_w4623_
	);
	LUT2 #(
		.INIT('hb)
	) name4171 (
		_w4622_,
		_w4623_,
		_w4624_
	);
	LUT4 #(
		.INIT('hc0a0)
	) name4172 (
		\Datao[8]_pad ,
		\EAX_reg[8]/NET0131 ,
		_w695_,
		_w2422_,
		_w4625_
	);
	LUT4 #(
		.INIT('h3f15)
	) name4173 (
		\Datao[8]_pad ,
		\lWord_reg[8]/NET0131 ,
		_w696_,
		_w2159_,
		_w4626_
	);
	LUT2 #(
		.INIT('hb)
	) name4174 (
		_w4625_,
		_w4626_,
		_w4627_
	);
	LUT4 #(
		.INIT('hc0a0)
	) name4175 (
		\Datao[9]_pad ,
		\EAX_reg[9]/NET0131 ,
		_w695_,
		_w2422_,
		_w4628_
	);
	LUT4 #(
		.INIT('h3f15)
	) name4176 (
		\Datao[9]_pad ,
		\lWord_reg[9]/NET0131 ,
		_w696_,
		_w2159_,
		_w4629_
	);
	LUT2 #(
		.INIT('hb)
	) name4177 (
		_w4628_,
		_w4629_,
		_w4630_
	);
	LUT4 #(
		.INIT('hc0a0)
	) name4178 (
		\Datao[0]_pad ,
		\EAX_reg[0]/NET0131 ,
		_w695_,
		_w2422_,
		_w4631_
	);
	LUT4 #(
		.INIT('h3f15)
	) name4179 (
		\Datao[0]_pad ,
		\lWord_reg[0]/NET0131 ,
		_w696_,
		_w2159_,
		_w4632_
	);
	LUT2 #(
		.INIT('hb)
	) name4180 (
		_w4631_,
		_w4632_,
		_w4633_
	);
	LUT4 #(
		.INIT('hc0a0)
	) name4181 (
		\Datao[10]_pad ,
		\EAX_reg[10]/NET0131 ,
		_w695_,
		_w2422_,
		_w4634_
	);
	LUT4 #(
		.INIT('h3f15)
	) name4182 (
		\Datao[10]_pad ,
		\lWord_reg[10]/NET0131 ,
		_w696_,
		_w2159_,
		_w4635_
	);
	LUT2 #(
		.INIT('hb)
	) name4183 (
		_w4634_,
		_w4635_,
		_w4636_
	);
	LUT4 #(
		.INIT('hc0a0)
	) name4184 (
		\Datao[12]_pad ,
		\EAX_reg[12]/NET0131 ,
		_w695_,
		_w2422_,
		_w4637_
	);
	LUT4 #(
		.INIT('h3f15)
	) name4185 (
		\Datao[12]_pad ,
		\lWord_reg[12]/NET0131 ,
		_w696_,
		_w2159_,
		_w4638_
	);
	LUT2 #(
		.INIT('hb)
	) name4186 (
		_w4637_,
		_w4638_,
		_w4639_
	);
	LUT4 #(
		.INIT('hc0a0)
	) name4187 (
		\Datao[11]_pad ,
		\EAX_reg[11]/NET0131 ,
		_w695_,
		_w2422_,
		_w4640_
	);
	LUT4 #(
		.INIT('h3f15)
	) name4188 (
		\Datao[11]_pad ,
		\lWord_reg[11]/NET0131 ,
		_w696_,
		_w2159_,
		_w4641_
	);
	LUT2 #(
		.INIT('hb)
	) name4189 (
		_w4640_,
		_w4641_,
		_w4642_
	);
	LUT4 #(
		.INIT('hc0a0)
	) name4190 (
		\Datao[13]_pad ,
		\EAX_reg[13]/NET0131 ,
		_w695_,
		_w2422_,
		_w4643_
	);
	LUT4 #(
		.INIT('h3f15)
	) name4191 (
		\Datao[13]_pad ,
		\lWord_reg[13]/NET0131 ,
		_w696_,
		_w2159_,
		_w4644_
	);
	LUT2 #(
		.INIT('hb)
	) name4192 (
		_w4643_,
		_w4644_,
		_w4645_
	);
	LUT4 #(
		.INIT('hc0a0)
	) name4193 (
		\Datao[14]_pad ,
		\EAX_reg[14]/NET0131 ,
		_w695_,
		_w2422_,
		_w4646_
	);
	LUT4 #(
		.INIT('h3f15)
	) name4194 (
		\Datao[14]_pad ,
		\lWord_reg[14]/NET0131 ,
		_w696_,
		_w2159_,
		_w4647_
	);
	LUT2 #(
		.INIT('hb)
	) name4195 (
		_w4646_,
		_w4647_,
		_w4648_
	);
	LUT4 #(
		.INIT('hc0a0)
	) name4196 (
		\Datao[15]_pad ,
		\EAX_reg[15]/NET0131 ,
		_w695_,
		_w2422_,
		_w4649_
	);
	LUT4 #(
		.INIT('h3f15)
	) name4197 (
		\Datao[15]_pad ,
		\lWord_reg[15]/NET0131 ,
		_w696_,
		_w2159_,
		_w4650_
	);
	LUT2 #(
		.INIT('hb)
	) name4198 (
		_w4649_,
		_w4650_,
		_w4651_
	);
	LUT4 #(
		.INIT('hc0a0)
	) name4199 (
		\Datao[1]_pad ,
		\EAX_reg[1]/NET0131 ,
		_w695_,
		_w2422_,
		_w4652_
	);
	LUT4 #(
		.INIT('h3f15)
	) name4200 (
		\Datao[1]_pad ,
		\lWord_reg[1]/NET0131 ,
		_w696_,
		_w2159_,
		_w4653_
	);
	LUT2 #(
		.INIT('hb)
	) name4201 (
		_w4652_,
		_w4653_,
		_w4654_
	);
	LUT4 #(
		.INIT('h0008)
	) name4202 (
		\DataWidth_reg[1]/NET0131 ,
		_w700_,
		_w2186_,
		_w2253_,
		_w4655_
	);
	LUT4 #(
		.INIT('h807f)
	) name4203 (
		\InstQueueWr_Addr_reg[0]/NET0131 ,
		\InstQueueWr_Addr_reg[1]/NET0131 ,
		\InstQueueWr_Addr_reg[2]/NET0131 ,
		\InstQueueWr_Addr_reg[3]/NET0131 ,
		_w4656_
	);
	LUT4 #(
		.INIT('h3fc0)
	) name4204 (
		\InstQueueWr_Addr_reg[0]/NET0131 ,
		\InstQueueWr_Addr_reg[1]/NET0131 ,
		\InstQueueWr_Addr_reg[2]/NET0131 ,
		\InstQueueWr_Addr_reg[3]/NET0131 ,
		_w4657_
	);
	LUT3 #(
		.INIT('he0)
	) name4205 (
		_w1281_,
		_w4655_,
		_w4657_,
		_w4658_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name4206 (
		\InstQueueWr_Addr_reg[3]/NET0131 ,
		_w3691_,
		_w4588_,
		_w4589_,
		_w4659_
	);
	LUT2 #(
		.INIT('h2)
	) name4207 (
		_w722_,
		_w4656_,
		_w4660_
	);
	LUT4 #(
		.INIT('hefcf)
	) name4208 (
		\InstQueueWr_Addr_reg[0]/NET0131 ,
		\InstQueueWr_Addr_reg[1]/NET0131 ,
		\InstQueueWr_Addr_reg[2]/NET0131 ,
		\InstQueueWr_Addr_reg[3]/NET0131 ,
		_w4661_
	);
	LUT4 #(
		.INIT('h0008)
	) name4209 (
		\DataWidth_reg[1]/NET0131 ,
		_w700_,
		_w2253_,
		_w4661_,
		_w4662_
	);
	LUT2 #(
		.INIT('h1)
	) name4210 (
		_w4660_,
		_w4662_,
		_w4663_
	);
	LUT3 #(
		.INIT('hef)
	) name4211 (
		_w4659_,
		_w4658_,
		_w4663_,
		_w4664_
	);
	LUT3 #(
		.INIT('h8a)
	) name4212 (
		\InstQueueWr_Addr_reg[1]/NET0131 ,
		_w4588_,
		_w4589_,
		_w4665_
	);
	LUT2 #(
		.INIT('h4)
	) name4213 (
		\InstQueueWr_Addr_reg[0]/NET0131 ,
		_w722_,
		_w4666_
	);
	LUT4 #(
		.INIT('h4c00)
	) name4214 (
		\DataWidth_reg[1]/NET0131 ,
		\InstQueueWr_Addr_reg[1]/NET0131 ,
		_w700_,
		_w3691_,
		_w4667_
	);
	LUT3 #(
		.INIT('h13)
	) name4215 (
		\InstQueueWr_Addr_reg[0]/NET0131 ,
		\InstQueueWr_Addr_reg[1]/NET0131 ,
		_w722_,
		_w4668_
	);
	LUT4 #(
		.INIT('h8acf)
	) name4216 (
		_w1281_,
		_w4666_,
		_w4667_,
		_w4668_,
		_w4669_
	);
	LUT2 #(
		.INIT('he)
	) name4217 (
		_w4665_,
		_w4669_,
		_w4670_
	);
	LUT4 #(
		.INIT('hfd80)
	) name4218 (
		\State2_reg[0]/NET0131 ,
		\State2_reg[1]/NET0131 ,
		\State2_reg[2]/NET0131 ,
		\State2_reg[3]/NET0131 ,
		_w4671_
	);
	LUT2 #(
		.INIT('h2)
	) name4219 (
		\InstQueueWr_Addr_reg[0]/NET0131 ,
		_w4671_,
		_w4672_
	);
	LUT2 #(
		.INIT('h1)
	) name4220 (
		\Flush_reg/NET0131 ,
		\InstQueueWr_Addr_reg[0]/NET0131 ,
		_w4673_
	);
	LUT4 #(
		.INIT('h002a)
	) name4221 (
		_w712_,
		_w713_,
		_w714_,
		_w4673_,
		_w4674_
	);
	LUT3 #(
		.INIT('hfe)
	) name4222 (
		_w4666_,
		_w4674_,
		_w4672_,
		_w4675_
	);
	LUT3 #(
		.INIT('h48)
	) name4223 (
		\Datai[25]_pad ,
		_w2187_,
		_w2196_,
		_w4676_
	);
	LUT4 #(
		.INIT('hcc6c)
	) name4224 (
		\Datai[16]_pad ,
		\Datai[17]_pad ,
		\Datai[31]_pad ,
		_w2192_,
		_w4677_
	);
	LUT2 #(
		.INIT('h8)
	) name4225 (
		_w2203_,
		_w4677_,
		_w4678_
	);
	LUT4 #(
		.INIT('h5553)
	) name4226 (
		\Datai[1]_pad ,
		\InstQueue_reg[0][1]/NET0131 ,
		_w2205_,
		_w2207_,
		_w4679_
	);
	LUT2 #(
		.INIT('h1)
	) name4227 (
		_w2211_,
		_w4679_,
		_w4680_
	);
	LUT4 #(
		.INIT('h0057)
	) name4228 (
		\DataWidth_reg[1]/NET0131 ,
		_w4676_,
		_w4678_,
		_w4680_,
		_w4681_
	);
	LUT4 #(
		.INIT('hc055)
	) name4229 (
		\InstQueue_reg[0][1]/NET0131 ,
		_w508_,
		_w513_,
		_w2205_,
		_w4682_
	);
	LUT2 #(
		.INIT('h2)
	) name4230 (
		\InstQueue_reg[0][1]/NET0131 ,
		_w2215_,
		_w4683_
	);
	LUT3 #(
		.INIT('h0d)
	) name4231 (
		_w706_,
		_w4679_,
		_w4683_,
		_w4684_
	);
	LUT3 #(
		.INIT('hd0)
	) name4232 (
		_w722_,
		_w4682_,
		_w4684_,
		_w4685_
	);
	LUT3 #(
		.INIT('h2f)
	) name4233 (
		_w700_,
		_w4681_,
		_w4685_,
		_w4686_
	);
	LUT3 #(
		.INIT('h60)
	) name4234 (
		\Datai[25]_pad ,
		_w2196_,
		_w2220_,
		_w4687_
	);
	LUT2 #(
		.INIT('h8)
	) name4235 (
		_w2222_,
		_w4677_,
		_w4688_
	);
	LUT4 #(
		.INIT('h5553)
	) name4236 (
		\Datai[1]_pad ,
		\InstQueue_reg[10][1]/NET0131 ,
		_w2224_,
		_w2225_,
		_w4689_
	);
	LUT2 #(
		.INIT('h1)
	) name4237 (
		_w2229_,
		_w4689_,
		_w4690_
	);
	LUT4 #(
		.INIT('h0057)
	) name4238 (
		\DataWidth_reg[1]/NET0131 ,
		_w4687_,
		_w4688_,
		_w4690_,
		_w4691_
	);
	LUT4 #(
		.INIT('hc055)
	) name4239 (
		\InstQueue_reg[10][1]/NET0131 ,
		_w508_,
		_w513_,
		_w2224_,
		_w4692_
	);
	LUT2 #(
		.INIT('h2)
	) name4240 (
		\InstQueue_reg[10][1]/NET0131 ,
		_w2215_,
		_w4693_
	);
	LUT3 #(
		.INIT('h0d)
	) name4241 (
		_w706_,
		_w4689_,
		_w4693_,
		_w4694_
	);
	LUT3 #(
		.INIT('hd0)
	) name4242 (
		_w722_,
		_w4692_,
		_w4694_,
		_w4695_
	);
	LUT3 #(
		.INIT('h2f)
	) name4243 (
		_w700_,
		_w4691_,
		_w4695_,
		_w4696_
	);
	LUT4 #(
		.INIT('ha666)
	) name4244 (
		\Datai[24]_pad ,
		\Datai[31]_pad ,
		_w2192_,
		_w2195_,
		_w4697_
	);
	LUT4 #(
		.INIT('ha600)
	) name4245 (
		\Datai[16]_pad ,
		\Datai[31]_pad ,
		_w2192_,
		_w2225_,
		_w4698_
	);
	LUT4 #(
		.INIT('haa80)
	) name4246 (
		\DataWidth_reg[1]/NET0131 ,
		_w2222_,
		_w4697_,
		_w4698_,
		_w4699_
	);
	LUT4 #(
		.INIT('h5553)
	) name4247 (
		\Datai[0]_pad ,
		\InstQueue_reg[11][0]/NET0131 ,
		_w2224_,
		_w2239_,
		_w4700_
	);
	LUT2 #(
		.INIT('h1)
	) name4248 (
		_w2243_,
		_w4700_,
		_w4701_
	);
	LUT3 #(
		.INIT('ha8)
	) name4249 (
		_w700_,
		_w4699_,
		_w4701_,
		_w4702_
	);
	LUT4 #(
		.INIT('hc055)
	) name4250 (
		\InstQueue_reg[11][0]/NET0131 ,
		_w530_,
		_w535_,
		_w2239_,
		_w4703_
	);
	LUT2 #(
		.INIT('h2)
	) name4251 (
		\InstQueue_reg[11][0]/NET0131 ,
		_w2215_,
		_w4704_
	);
	LUT3 #(
		.INIT('h0d)
	) name4252 (
		_w706_,
		_w4700_,
		_w4704_,
		_w4705_
	);
	LUT3 #(
		.INIT('hd0)
	) name4253 (
		_w722_,
		_w4703_,
		_w4705_,
		_w4706_
	);
	LUT2 #(
		.INIT('hb)
	) name4254 (
		_w4702_,
		_w4706_,
		_w4707_
	);
	LUT3 #(
		.INIT('h60)
	) name4255 (
		\Datai[25]_pad ,
		_w2196_,
		_w2222_,
		_w4708_
	);
	LUT2 #(
		.INIT('h8)
	) name4256 (
		_w2225_,
		_w4677_,
		_w4709_
	);
	LUT4 #(
		.INIT('h5553)
	) name4257 (
		\Datai[1]_pad ,
		\InstQueue_reg[11][1]/NET0131 ,
		_w2224_,
		_w2239_,
		_w4710_
	);
	LUT2 #(
		.INIT('h1)
	) name4258 (
		_w2243_,
		_w4710_,
		_w4711_
	);
	LUT4 #(
		.INIT('h0057)
	) name4259 (
		\DataWidth_reg[1]/NET0131 ,
		_w4708_,
		_w4709_,
		_w4711_,
		_w4712_
	);
	LUT4 #(
		.INIT('hc055)
	) name4260 (
		\InstQueue_reg[11][1]/NET0131 ,
		_w508_,
		_w513_,
		_w2239_,
		_w4713_
	);
	LUT2 #(
		.INIT('h2)
	) name4261 (
		\InstQueue_reg[11][1]/NET0131 ,
		_w2215_,
		_w4714_
	);
	LUT3 #(
		.INIT('h0d)
	) name4262 (
		_w706_,
		_w4710_,
		_w4714_,
		_w4715_
	);
	LUT3 #(
		.INIT('hd0)
	) name4263 (
		_w722_,
		_w4713_,
		_w4715_,
		_w4716_
	);
	LUT3 #(
		.INIT('h2f)
	) name4264 (
		_w700_,
		_w4712_,
		_w4716_,
		_w4717_
	);
	LUT3 #(
		.INIT('h60)
	) name4265 (
		\Datai[25]_pad ,
		_w2196_,
		_w2225_,
		_w4718_
	);
	LUT2 #(
		.INIT('h8)
	) name4266 (
		_w2224_,
		_w4677_,
		_w4719_
	);
	LUT4 #(
		.INIT('h5553)
	) name4267 (
		\Datai[1]_pad ,
		\InstQueue_reg[12][1]/NET0131 ,
		_w2239_,
		_w2253_,
		_w4720_
	);
	LUT2 #(
		.INIT('h1)
	) name4268 (
		_w2256_,
		_w4720_,
		_w4721_
	);
	LUT4 #(
		.INIT('h0057)
	) name4269 (
		\DataWidth_reg[1]/NET0131 ,
		_w4718_,
		_w4719_,
		_w4721_,
		_w4722_
	);
	LUT4 #(
		.INIT('hc055)
	) name4270 (
		\InstQueue_reg[12][1]/NET0131 ,
		_w508_,
		_w513_,
		_w2253_,
		_w4723_
	);
	LUT2 #(
		.INIT('h2)
	) name4271 (
		\InstQueue_reg[12][1]/NET0131 ,
		_w2215_,
		_w4724_
	);
	LUT3 #(
		.INIT('h0d)
	) name4272 (
		_w706_,
		_w4720_,
		_w4724_,
		_w4725_
	);
	LUT3 #(
		.INIT('hd0)
	) name4273 (
		_w722_,
		_w4723_,
		_w4725_,
		_w4726_
	);
	LUT3 #(
		.INIT('h2f)
	) name4274 (
		_w700_,
		_w4722_,
		_w4726_,
		_w4727_
	);
	LUT3 #(
		.INIT('h60)
	) name4275 (
		\Datai[25]_pad ,
		_w2196_,
		_w2224_,
		_w4728_
	);
	LUT2 #(
		.INIT('h8)
	) name4276 (
		_w2239_,
		_w4677_,
		_w4729_
	);
	LUT4 #(
		.INIT('h5553)
	) name4277 (
		\Datai[1]_pad ,
		\InstQueue_reg[13][1]/NET0131 ,
		_w2187_,
		_w2253_,
		_w4730_
	);
	LUT2 #(
		.INIT('h1)
	) name4278 (
		_w2268_,
		_w4730_,
		_w4731_
	);
	LUT4 #(
		.INIT('h0057)
	) name4279 (
		\DataWidth_reg[1]/NET0131 ,
		_w4728_,
		_w4729_,
		_w4731_,
		_w4732_
	);
	LUT4 #(
		.INIT('hc055)
	) name4280 (
		\InstQueue_reg[13][1]/NET0131 ,
		_w508_,
		_w513_,
		_w2187_,
		_w4733_
	);
	LUT2 #(
		.INIT('h2)
	) name4281 (
		\InstQueue_reg[13][1]/NET0131 ,
		_w2215_,
		_w4734_
	);
	LUT3 #(
		.INIT('h0d)
	) name4282 (
		_w706_,
		_w4730_,
		_w4734_,
		_w4735_
	);
	LUT3 #(
		.INIT('hd0)
	) name4283 (
		_w722_,
		_w4733_,
		_w4735_,
		_w4736_
	);
	LUT3 #(
		.INIT('h2f)
	) name4284 (
		_w700_,
		_w4732_,
		_w4736_,
		_w4737_
	);
	LUT3 #(
		.INIT('h60)
	) name4285 (
		\Datai[25]_pad ,
		_w2196_,
		_w2239_,
		_w4738_
	);
	LUT2 #(
		.INIT('h8)
	) name4286 (
		_w2253_,
		_w4677_,
		_w4739_
	);
	LUT4 #(
		.INIT('h5553)
	) name4287 (
		\Datai[1]_pad ,
		\InstQueue_reg[14][1]/NET0131 ,
		_w2187_,
		_w2203_,
		_w4740_
	);
	LUT2 #(
		.INIT('h1)
	) name4288 (
		_w2279_,
		_w4740_,
		_w4741_
	);
	LUT4 #(
		.INIT('h0057)
	) name4289 (
		\DataWidth_reg[1]/NET0131 ,
		_w4738_,
		_w4739_,
		_w4741_,
		_w4742_
	);
	LUT4 #(
		.INIT('hc055)
	) name4290 (
		\InstQueue_reg[14][1]/NET0131 ,
		_w508_,
		_w513_,
		_w2203_,
		_w4743_
	);
	LUT2 #(
		.INIT('h2)
	) name4291 (
		\InstQueue_reg[14][1]/NET0131 ,
		_w2215_,
		_w4744_
	);
	LUT3 #(
		.INIT('h0d)
	) name4292 (
		_w706_,
		_w4740_,
		_w4744_,
		_w4745_
	);
	LUT3 #(
		.INIT('hd0)
	) name4293 (
		_w722_,
		_w4743_,
		_w4745_,
		_w4746_
	);
	LUT3 #(
		.INIT('h2f)
	) name4294 (
		_w700_,
		_w4742_,
		_w4746_,
		_w4747_
	);
	LUT3 #(
		.INIT('h60)
	) name4295 (
		\Datai[25]_pad ,
		_w2196_,
		_w2253_,
		_w4748_
	);
	LUT2 #(
		.INIT('h8)
	) name4296 (
		_w2187_,
		_w4677_,
		_w4749_
	);
	LUT4 #(
		.INIT('h5553)
	) name4297 (
		\Datai[1]_pad ,
		\InstQueue_reg[15][1]/NET0131 ,
		_w2207_,
		_w2203_,
		_w4750_
	);
	LUT2 #(
		.INIT('h1)
	) name4298 (
		_w2291_,
		_w4750_,
		_w4751_
	);
	LUT4 #(
		.INIT('h0057)
	) name4299 (
		\DataWidth_reg[1]/NET0131 ,
		_w4748_,
		_w4749_,
		_w4751_,
		_w4752_
	);
	LUT4 #(
		.INIT('hc055)
	) name4300 (
		\InstQueue_reg[15][1]/NET0131 ,
		_w508_,
		_w513_,
		_w2207_,
		_w4753_
	);
	LUT2 #(
		.INIT('h2)
	) name4301 (
		\InstQueue_reg[15][1]/NET0131 ,
		_w2215_,
		_w4754_
	);
	LUT3 #(
		.INIT('h0d)
	) name4302 (
		_w706_,
		_w4750_,
		_w4754_,
		_w4755_
	);
	LUT3 #(
		.INIT('hd0)
	) name4303 (
		_w722_,
		_w4753_,
		_w4755_,
		_w4756_
	);
	LUT3 #(
		.INIT('h2f)
	) name4304 (
		_w700_,
		_w4752_,
		_w4756_,
		_w4757_
	);
	LUT3 #(
		.INIT('h60)
	) name4305 (
		\Datai[25]_pad ,
		_w2196_,
		_w2203_,
		_w4758_
	);
	LUT2 #(
		.INIT('h8)
	) name4306 (
		_w2207_,
		_w4677_,
		_w4759_
	);
	LUT4 #(
		.INIT('h5553)
	) name4307 (
		\Datai[1]_pad ,
		\InstQueue_reg[1][1]/NET0131 ,
		_w2205_,
		_w2301_,
		_w4760_
	);
	LUT2 #(
		.INIT('h1)
	) name4308 (
		_w2304_,
		_w4760_,
		_w4761_
	);
	LUT4 #(
		.INIT('h0057)
	) name4309 (
		\DataWidth_reg[1]/NET0131 ,
		_w4758_,
		_w4759_,
		_w4761_,
		_w4762_
	);
	LUT4 #(
		.INIT('hc055)
	) name4310 (
		\InstQueue_reg[1][1]/NET0131 ,
		_w508_,
		_w513_,
		_w2301_,
		_w4763_
	);
	LUT2 #(
		.INIT('h2)
	) name4311 (
		\InstQueue_reg[1][1]/NET0131 ,
		_w2215_,
		_w4764_
	);
	LUT3 #(
		.INIT('h0d)
	) name4312 (
		_w706_,
		_w4760_,
		_w4764_,
		_w4765_
	);
	LUT3 #(
		.INIT('hd0)
	) name4313 (
		_w722_,
		_w4763_,
		_w4765_,
		_w4766_
	);
	LUT3 #(
		.INIT('h2f)
	) name4314 (
		_w700_,
		_w4762_,
		_w4766_,
		_w4767_
	);
	LUT2 #(
		.INIT('h8)
	) name4315 (
		_w2205_,
		_w4677_,
		_w4768_
	);
	LUT3 #(
		.INIT('h48)
	) name4316 (
		\Datai[25]_pad ,
		_w2207_,
		_w2196_,
		_w4769_
	);
	LUT4 #(
		.INIT('h5553)
	) name4317 (
		\Datai[1]_pad ,
		\InstQueue_reg[2][1]/NET0131 ,
		_w2301_,
		_w2314_,
		_w4770_
	);
	LUT2 #(
		.INIT('h1)
	) name4318 (
		_w2317_,
		_w4770_,
		_w4771_
	);
	LUT4 #(
		.INIT('h0057)
	) name4319 (
		\DataWidth_reg[1]/NET0131 ,
		_w4768_,
		_w4769_,
		_w4771_,
		_w4772_
	);
	LUT4 #(
		.INIT('hc055)
	) name4320 (
		\InstQueue_reg[2][1]/NET0131 ,
		_w508_,
		_w513_,
		_w2314_,
		_w4773_
	);
	LUT2 #(
		.INIT('h2)
	) name4321 (
		\InstQueue_reg[2][1]/NET0131 ,
		_w2215_,
		_w4774_
	);
	LUT3 #(
		.INIT('h0d)
	) name4322 (
		_w706_,
		_w4770_,
		_w4774_,
		_w4775_
	);
	LUT3 #(
		.INIT('hd0)
	) name4323 (
		_w722_,
		_w4773_,
		_w4775_,
		_w4776_
	);
	LUT3 #(
		.INIT('h2f)
	) name4324 (
		_w700_,
		_w4772_,
		_w4776_,
		_w4777_
	);
	LUT4 #(
		.INIT('ha600)
	) name4325 (
		\Datai[16]_pad ,
		\Datai[31]_pad ,
		_w2192_,
		_w2301_,
		_w4778_
	);
	LUT4 #(
		.INIT('haa80)
	) name4326 (
		\DataWidth_reg[1]/NET0131 ,
		_w2205_,
		_w4697_,
		_w4778_,
		_w4779_
	);
	LUT4 #(
		.INIT('h5553)
	) name4327 (
		\Datai[0]_pad ,
		\InstQueue_reg[3][0]/NET0131 ,
		_w2314_,
		_w2327_,
		_w4780_
	);
	LUT2 #(
		.INIT('h1)
	) name4328 (
		_w2330_,
		_w4780_,
		_w4781_
	);
	LUT3 #(
		.INIT('ha8)
	) name4329 (
		_w700_,
		_w4779_,
		_w4781_,
		_w4782_
	);
	LUT4 #(
		.INIT('hc055)
	) name4330 (
		\InstQueue_reg[3][0]/NET0131 ,
		_w530_,
		_w535_,
		_w2327_,
		_w4783_
	);
	LUT2 #(
		.INIT('h2)
	) name4331 (
		\InstQueue_reg[3][0]/NET0131 ,
		_w2215_,
		_w4784_
	);
	LUT3 #(
		.INIT('h0d)
	) name4332 (
		_w706_,
		_w4780_,
		_w4784_,
		_w4785_
	);
	LUT3 #(
		.INIT('hd0)
	) name4333 (
		_w722_,
		_w4783_,
		_w4785_,
		_w4786_
	);
	LUT2 #(
		.INIT('hb)
	) name4334 (
		_w4782_,
		_w4786_,
		_w4787_
	);
	LUT3 #(
		.INIT('h48)
	) name4335 (
		\Datai[25]_pad ,
		_w2205_,
		_w2196_,
		_w4788_
	);
	LUT2 #(
		.INIT('h8)
	) name4336 (
		_w2301_,
		_w4677_,
		_w4789_
	);
	LUT4 #(
		.INIT('h5553)
	) name4337 (
		\Datai[1]_pad ,
		\InstQueue_reg[3][1]/NET0131 ,
		_w2314_,
		_w2327_,
		_w4790_
	);
	LUT2 #(
		.INIT('h1)
	) name4338 (
		_w2330_,
		_w4790_,
		_w4791_
	);
	LUT4 #(
		.INIT('h0057)
	) name4339 (
		\DataWidth_reg[1]/NET0131 ,
		_w4788_,
		_w4789_,
		_w4791_,
		_w4792_
	);
	LUT4 #(
		.INIT('hc055)
	) name4340 (
		\InstQueue_reg[3][1]/NET0131 ,
		_w508_,
		_w513_,
		_w2327_,
		_w4793_
	);
	LUT2 #(
		.INIT('h2)
	) name4341 (
		\InstQueue_reg[3][1]/NET0131 ,
		_w2215_,
		_w4794_
	);
	LUT3 #(
		.INIT('h0d)
	) name4342 (
		_w706_,
		_w4790_,
		_w4794_,
		_w4795_
	);
	LUT3 #(
		.INIT('hd0)
	) name4343 (
		_w722_,
		_w4793_,
		_w4795_,
		_w4796_
	);
	LUT3 #(
		.INIT('h2f)
	) name4344 (
		_w700_,
		_w4792_,
		_w4796_,
		_w4797_
	);
	LUT3 #(
		.INIT('h60)
	) name4345 (
		\Datai[25]_pad ,
		_w2196_,
		_w2301_,
		_w4798_
	);
	LUT2 #(
		.INIT('h8)
	) name4346 (
		_w2314_,
		_w4677_,
		_w4799_
	);
	LUT4 #(
		.INIT('h5553)
	) name4347 (
		\Datai[1]_pad ,
		\InstQueue_reg[4][1]/NET0131 ,
		_w2327_,
		_w2340_,
		_w4800_
	);
	LUT2 #(
		.INIT('h1)
	) name4348 (
		_w2343_,
		_w4800_,
		_w4801_
	);
	LUT4 #(
		.INIT('h0057)
	) name4349 (
		\DataWidth_reg[1]/NET0131 ,
		_w4798_,
		_w4799_,
		_w4801_,
		_w4802_
	);
	LUT4 #(
		.INIT('hc055)
	) name4350 (
		\InstQueue_reg[4][1]/NET0131 ,
		_w508_,
		_w513_,
		_w2340_,
		_w4803_
	);
	LUT2 #(
		.INIT('h2)
	) name4351 (
		\InstQueue_reg[4][1]/NET0131 ,
		_w2215_,
		_w4804_
	);
	LUT3 #(
		.INIT('h0d)
	) name4352 (
		_w706_,
		_w4800_,
		_w4804_,
		_w4805_
	);
	LUT3 #(
		.INIT('hd0)
	) name4353 (
		_w722_,
		_w4803_,
		_w4805_,
		_w4806_
	);
	LUT3 #(
		.INIT('h2f)
	) name4354 (
		_w700_,
		_w4802_,
		_w4806_,
		_w4807_
	);
	LUT3 #(
		.INIT('h60)
	) name4355 (
		\Datai[25]_pad ,
		_w2196_,
		_w2314_,
		_w4808_
	);
	LUT2 #(
		.INIT('h8)
	) name4356 (
		_w2327_,
		_w4677_,
		_w4809_
	);
	LUT4 #(
		.INIT('h5553)
	) name4357 (
		\Datai[1]_pad ,
		\InstQueue_reg[5][1]/NET0131 ,
		_w2340_,
		_w2353_,
		_w4810_
	);
	LUT2 #(
		.INIT('h1)
	) name4358 (
		_w2356_,
		_w4810_,
		_w4811_
	);
	LUT4 #(
		.INIT('h0057)
	) name4359 (
		\DataWidth_reg[1]/NET0131 ,
		_w4808_,
		_w4809_,
		_w4811_,
		_w4812_
	);
	LUT4 #(
		.INIT('hc055)
	) name4360 (
		\InstQueue_reg[5][1]/NET0131 ,
		_w508_,
		_w513_,
		_w2353_,
		_w4813_
	);
	LUT2 #(
		.INIT('h2)
	) name4361 (
		\InstQueue_reg[5][1]/NET0131 ,
		_w2215_,
		_w4814_
	);
	LUT3 #(
		.INIT('h0d)
	) name4362 (
		_w706_,
		_w4810_,
		_w4814_,
		_w4815_
	);
	LUT3 #(
		.INIT('hd0)
	) name4363 (
		_w722_,
		_w4813_,
		_w4815_,
		_w4816_
	);
	LUT3 #(
		.INIT('h2f)
	) name4364 (
		_w700_,
		_w4812_,
		_w4816_,
		_w4817_
	);
	LUT3 #(
		.INIT('h60)
	) name4365 (
		\Datai[25]_pad ,
		_w2196_,
		_w2327_,
		_w4818_
	);
	LUT2 #(
		.INIT('h8)
	) name4366 (
		_w2340_,
		_w4677_,
		_w4819_
	);
	LUT4 #(
		.INIT('h5553)
	) name4367 (
		\Datai[1]_pad ,
		\InstQueue_reg[6][1]/NET0131 ,
		_w2353_,
		_w2366_,
		_w4820_
	);
	LUT2 #(
		.INIT('h1)
	) name4368 (
		_w2369_,
		_w4820_,
		_w4821_
	);
	LUT4 #(
		.INIT('h0057)
	) name4369 (
		\DataWidth_reg[1]/NET0131 ,
		_w4818_,
		_w4819_,
		_w4821_,
		_w4822_
	);
	LUT4 #(
		.INIT('hc055)
	) name4370 (
		\InstQueue_reg[6][1]/NET0131 ,
		_w508_,
		_w513_,
		_w2366_,
		_w4823_
	);
	LUT2 #(
		.INIT('h2)
	) name4371 (
		\InstQueue_reg[6][1]/NET0131 ,
		_w2215_,
		_w4824_
	);
	LUT3 #(
		.INIT('h0d)
	) name4372 (
		_w706_,
		_w4820_,
		_w4824_,
		_w4825_
	);
	LUT3 #(
		.INIT('hd0)
	) name4373 (
		_w722_,
		_w4823_,
		_w4825_,
		_w4826_
	);
	LUT3 #(
		.INIT('h2f)
	) name4374 (
		_w700_,
		_w4822_,
		_w4826_,
		_w4827_
	);
	LUT4 #(
		.INIT('ha600)
	) name4375 (
		\Datai[16]_pad ,
		\Datai[31]_pad ,
		_w2192_,
		_w2353_,
		_w4828_
	);
	LUT4 #(
		.INIT('haa80)
	) name4376 (
		\DataWidth_reg[1]/NET0131 ,
		_w2340_,
		_w4697_,
		_w4828_,
		_w4829_
	);
	LUT4 #(
		.INIT('h5553)
	) name4377 (
		\Datai[0]_pad ,
		\InstQueue_reg[7][0]/NET0131 ,
		_w2220_,
		_w2366_,
		_w4830_
	);
	LUT2 #(
		.INIT('h1)
	) name4378 (
		_w2381_,
		_w4830_,
		_w4831_
	);
	LUT3 #(
		.INIT('ha8)
	) name4379 (
		_w700_,
		_w4829_,
		_w4831_,
		_w4832_
	);
	LUT4 #(
		.INIT('hc055)
	) name4380 (
		\InstQueue_reg[7][0]/NET0131 ,
		_w530_,
		_w535_,
		_w2220_,
		_w4833_
	);
	LUT2 #(
		.INIT('h2)
	) name4381 (
		\InstQueue_reg[7][0]/NET0131 ,
		_w2215_,
		_w4834_
	);
	LUT3 #(
		.INIT('h0d)
	) name4382 (
		_w706_,
		_w4830_,
		_w4834_,
		_w4835_
	);
	LUT3 #(
		.INIT('hd0)
	) name4383 (
		_w722_,
		_w4833_,
		_w4835_,
		_w4836_
	);
	LUT2 #(
		.INIT('hb)
	) name4384 (
		_w4832_,
		_w4836_,
		_w4837_
	);
	LUT3 #(
		.INIT('h60)
	) name4385 (
		\Datai[25]_pad ,
		_w2196_,
		_w2340_,
		_w4838_
	);
	LUT2 #(
		.INIT('h8)
	) name4386 (
		_w2353_,
		_w4677_,
		_w4839_
	);
	LUT4 #(
		.INIT('h5553)
	) name4387 (
		\Datai[1]_pad ,
		\InstQueue_reg[7][1]/NET0131 ,
		_w2220_,
		_w2366_,
		_w4840_
	);
	LUT2 #(
		.INIT('h1)
	) name4388 (
		_w2381_,
		_w4840_,
		_w4841_
	);
	LUT4 #(
		.INIT('h0057)
	) name4389 (
		\DataWidth_reg[1]/NET0131 ,
		_w4838_,
		_w4839_,
		_w4841_,
		_w4842_
	);
	LUT4 #(
		.INIT('hc055)
	) name4390 (
		\InstQueue_reg[7][1]/NET0131 ,
		_w508_,
		_w513_,
		_w2220_,
		_w4843_
	);
	LUT2 #(
		.INIT('h2)
	) name4391 (
		\InstQueue_reg[7][1]/NET0131 ,
		_w2215_,
		_w4844_
	);
	LUT3 #(
		.INIT('h0d)
	) name4392 (
		_w706_,
		_w4840_,
		_w4844_,
		_w4845_
	);
	LUT3 #(
		.INIT('hd0)
	) name4393 (
		_w722_,
		_w4843_,
		_w4845_,
		_w4846_
	);
	LUT3 #(
		.INIT('h2f)
	) name4394 (
		_w700_,
		_w4842_,
		_w4846_,
		_w4847_
	);
	LUT3 #(
		.INIT('h60)
	) name4395 (
		\Datai[25]_pad ,
		_w2196_,
		_w2353_,
		_w4848_
	);
	LUT2 #(
		.INIT('h8)
	) name4396 (
		_w2366_,
		_w4677_,
		_w4849_
	);
	LUT4 #(
		.INIT('h5553)
	) name4397 (
		\Datai[1]_pad ,
		\InstQueue_reg[8][1]/NET0131 ,
		_w2220_,
		_w2222_,
		_w4850_
	);
	LUT2 #(
		.INIT('h1)
	) name4398 (
		_w2392_,
		_w4850_,
		_w4851_
	);
	LUT4 #(
		.INIT('h0057)
	) name4399 (
		\DataWidth_reg[1]/NET0131 ,
		_w4848_,
		_w4849_,
		_w4851_,
		_w4852_
	);
	LUT4 #(
		.INIT('hc055)
	) name4400 (
		\InstQueue_reg[8][1]/NET0131 ,
		_w508_,
		_w513_,
		_w2222_,
		_w4853_
	);
	LUT2 #(
		.INIT('h2)
	) name4401 (
		\InstQueue_reg[8][1]/NET0131 ,
		_w2215_,
		_w4854_
	);
	LUT3 #(
		.INIT('h0d)
	) name4402 (
		_w706_,
		_w4850_,
		_w4854_,
		_w4855_
	);
	LUT3 #(
		.INIT('hd0)
	) name4403 (
		_w722_,
		_w4853_,
		_w4855_,
		_w4856_
	);
	LUT3 #(
		.INIT('h2f)
	) name4404 (
		_w700_,
		_w4852_,
		_w4856_,
		_w4857_
	);
	LUT3 #(
		.INIT('h60)
	) name4405 (
		\Datai[25]_pad ,
		_w2196_,
		_w2366_,
		_w4858_
	);
	LUT2 #(
		.INIT('h8)
	) name4406 (
		_w2220_,
		_w4677_,
		_w4859_
	);
	LUT4 #(
		.INIT('h5553)
	) name4407 (
		\Datai[1]_pad ,
		\InstQueue_reg[9][1]/NET0131 ,
		_w2225_,
		_w2222_,
		_w4860_
	);
	LUT2 #(
		.INIT('h1)
	) name4408 (
		_w2403_,
		_w4860_,
		_w4861_
	);
	LUT4 #(
		.INIT('h0057)
	) name4409 (
		\DataWidth_reg[1]/NET0131 ,
		_w4858_,
		_w4859_,
		_w4861_,
		_w4862_
	);
	LUT4 #(
		.INIT('hc055)
	) name4410 (
		\InstQueue_reg[9][1]/NET0131 ,
		_w508_,
		_w513_,
		_w2225_,
		_w4863_
	);
	LUT2 #(
		.INIT('h2)
	) name4411 (
		\InstQueue_reg[9][1]/NET0131 ,
		_w2215_,
		_w4864_
	);
	LUT3 #(
		.INIT('h0d)
	) name4412 (
		_w706_,
		_w4860_,
		_w4864_,
		_w4865_
	);
	LUT3 #(
		.INIT('hd0)
	) name4413 (
		_w722_,
		_w4863_,
		_w4865_,
		_w4866_
	);
	LUT3 #(
		.INIT('h2f)
	) name4414 (
		_w700_,
		_w4862_,
		_w4866_,
		_w4867_
	);
	LUT3 #(
		.INIT('h48)
	) name4415 (
		\rEIP_reg[26]/NET0131 ,
		_w615_,
		_w4558_,
		_w4868_
	);
	LUT3 #(
		.INIT('h8a)
	) name4416 (
		\Address[24]_pad ,
		\State_reg[0]/NET0131 ,
		\State_reg[1]/NET0131 ,
		_w4869_
	);
	LUT4 #(
		.INIT('h60a0)
	) name4417 (
		\rEIP_reg[25]/NET0131 ,
		_w3263_,
		_w4565_,
		_w4562_,
		_w4870_
	);
	LUT2 #(
		.INIT('h1)
	) name4418 (
		_w4869_,
		_w4870_,
		_w4871_
	);
	LUT2 #(
		.INIT('hb)
	) name4419 (
		_w4868_,
		_w4871_,
		_w4872_
	);
	LUT3 #(
		.INIT('h48)
	) name4420 (
		\rEIP_reg[14]/NET0131 ,
		_w615_,
		_w4554_,
		_w4873_
	);
	LUT3 #(
		.INIT('h8a)
	) name4421 (
		\Address[12]_pad ,
		\State_reg[0]/NET0131 ,
		\State_reg[1]/NET0131 ,
		_w4874_
	);
	LUT4 #(
		.INIT('h60a0)
	) name4422 (
		\rEIP_reg[13]/NET0131 ,
		_w2609_,
		_w4565_,
		_w4562_,
		_w4875_
	);
	LUT2 #(
		.INIT('h1)
	) name4423 (
		_w4874_,
		_w4875_,
		_w4876_
	);
	LUT2 #(
		.INIT('hb)
	) name4424 (
		_w4873_,
		_w4876_,
		_w4877_
	);
	LUT3 #(
		.INIT('h48)
	) name4425 (
		\rEIP_reg[22]/NET0131 ,
		_w615_,
		_w4557_,
		_w4878_
	);
	LUT3 #(
		.INIT('h8a)
	) name4426 (
		\Address[20]_pad ,
		\State_reg[0]/NET0131 ,
		\State_reg[1]/NET0131 ,
		_w4879_
	);
	LUT3 #(
		.INIT('h80)
	) name4427 (
		_w2611_,
		_w2613_,
		_w4562_,
		_w4880_
	);
	LUT4 #(
		.INIT('h8000)
	) name4428 (
		\rEIP_reg[20]/NET0131 ,
		_w2611_,
		_w2613_,
		_w4562_,
		_w4881_
	);
	LUT4 #(
		.INIT('h70f0)
	) name4429 (
		_w2611_,
		_w2615_,
		_w4565_,
		_w4562_,
		_w4882_
	);
	LUT4 #(
		.INIT('h0133)
	) name4430 (
		\rEIP_reg[21]/NET0131 ,
		_w4879_,
		_w4881_,
		_w4882_,
		_w4883_
	);
	LUT2 #(
		.INIT('hb)
	) name4431 (
		_w4878_,
		_w4883_,
		_w4884_
	);
	LUT4 #(
		.INIT('h60a0)
	) name4432 (
		\rEIP_reg[10]/NET0131 ,
		\rEIP_reg[9]/NET0131 ,
		_w615_,
		_w4551_,
		_w4885_
	);
	LUT3 #(
		.INIT('h8a)
	) name4433 (
		\Address[8]_pad ,
		\State_reg[0]/NET0131 ,
		\State_reg[1]/NET0131 ,
		_w4886_
	);
	LUT4 #(
		.INIT('h8000)
	) name4434 (
		\rEIP_reg[5]/NET0131 ,
		\rEIP_reg[6]/NET0131 ,
		_w2606_,
		_w4562_,
		_w4887_
	);
	LUT3 #(
		.INIT('h80)
	) name4435 (
		\rEIP_reg[7]/NET0131 ,
		\rEIP_reg[8]/NET0131 ,
		_w4887_,
		_w4888_
	);
	LUT4 #(
		.INIT('h8000)
	) name4436 (
		\rEIP_reg[7]/NET0131 ,
		\rEIP_reg[8]/NET0131 ,
		\rEIP_reg[9]/NET0131 ,
		_w4887_,
		_w4889_
	);
	LUT4 #(
		.INIT('h0b07)
	) name4437 (
		\rEIP_reg[9]/NET0131 ,
		_w4565_,
		_w4886_,
		_w4888_,
		_w4890_
	);
	LUT2 #(
		.INIT('hb)
	) name4438 (
		_w4885_,
		_w4890_,
		_w4891_
	);
	LUT4 #(
		.INIT('ha600)
	) name4439 (
		\Datai[16]_pad ,
		\Datai[31]_pad ,
		_w2192_,
		_w2203_,
		_w4892_
	);
	LUT4 #(
		.INIT('haa80)
	) name4440 (
		\DataWidth_reg[1]/NET0131 ,
		_w2187_,
		_w4697_,
		_w4892_,
		_w4893_
	);
	LUT4 #(
		.INIT('h5553)
	) name4441 (
		\Datai[0]_pad ,
		\InstQueue_reg[0][0]/NET0131 ,
		_w2205_,
		_w2207_,
		_w4894_
	);
	LUT2 #(
		.INIT('h1)
	) name4442 (
		_w2211_,
		_w4894_,
		_w4895_
	);
	LUT3 #(
		.INIT('ha8)
	) name4443 (
		_w700_,
		_w4893_,
		_w4895_,
		_w4896_
	);
	LUT4 #(
		.INIT('hc055)
	) name4444 (
		\InstQueue_reg[0][0]/NET0131 ,
		_w530_,
		_w535_,
		_w2205_,
		_w4897_
	);
	LUT2 #(
		.INIT('h2)
	) name4445 (
		\InstQueue_reg[0][0]/NET0131 ,
		_w2215_,
		_w4898_
	);
	LUT3 #(
		.INIT('h0d)
	) name4446 (
		_w706_,
		_w4894_,
		_w4898_,
		_w4899_
	);
	LUT3 #(
		.INIT('hd0)
	) name4447 (
		_w722_,
		_w4897_,
		_w4899_,
		_w4900_
	);
	LUT2 #(
		.INIT('hb)
	) name4448 (
		_w4896_,
		_w4900_,
		_w4901_
	);
	LUT4 #(
		.INIT('ha600)
	) name4449 (
		\Datai[16]_pad ,
		\Datai[31]_pad ,
		_w2192_,
		_w2222_,
		_w4902_
	);
	LUT4 #(
		.INIT('haa80)
	) name4450 (
		\DataWidth_reg[1]/NET0131 ,
		_w2220_,
		_w4697_,
		_w4902_,
		_w4903_
	);
	LUT4 #(
		.INIT('h5553)
	) name4451 (
		\Datai[0]_pad ,
		\InstQueue_reg[10][0]/NET0131 ,
		_w2224_,
		_w2225_,
		_w4904_
	);
	LUT2 #(
		.INIT('h1)
	) name4452 (
		_w2229_,
		_w4904_,
		_w4905_
	);
	LUT3 #(
		.INIT('ha8)
	) name4453 (
		_w700_,
		_w4903_,
		_w4905_,
		_w4906_
	);
	LUT4 #(
		.INIT('hc055)
	) name4454 (
		\InstQueue_reg[10][0]/NET0131 ,
		_w530_,
		_w535_,
		_w2224_,
		_w4907_
	);
	LUT2 #(
		.INIT('h2)
	) name4455 (
		\InstQueue_reg[10][0]/NET0131 ,
		_w2215_,
		_w4908_
	);
	LUT3 #(
		.INIT('h0d)
	) name4456 (
		_w706_,
		_w4904_,
		_w4908_,
		_w4909_
	);
	LUT3 #(
		.INIT('hd0)
	) name4457 (
		_w722_,
		_w4907_,
		_w4909_,
		_w4910_
	);
	LUT2 #(
		.INIT('hb)
	) name4458 (
		_w4906_,
		_w4910_,
		_w4911_
	);
	LUT4 #(
		.INIT('ha600)
	) name4459 (
		\Datai[16]_pad ,
		\Datai[31]_pad ,
		_w2192_,
		_w2224_,
		_w4912_
	);
	LUT4 #(
		.INIT('haa80)
	) name4460 (
		\DataWidth_reg[1]/NET0131 ,
		_w2225_,
		_w4697_,
		_w4912_,
		_w4913_
	);
	LUT4 #(
		.INIT('h5553)
	) name4461 (
		\Datai[0]_pad ,
		\InstQueue_reg[12][0]/NET0131 ,
		_w2239_,
		_w2253_,
		_w4914_
	);
	LUT2 #(
		.INIT('h1)
	) name4462 (
		_w2256_,
		_w4914_,
		_w4915_
	);
	LUT3 #(
		.INIT('ha8)
	) name4463 (
		_w700_,
		_w4913_,
		_w4915_,
		_w4916_
	);
	LUT4 #(
		.INIT('hc055)
	) name4464 (
		\InstQueue_reg[12][0]/NET0131 ,
		_w530_,
		_w535_,
		_w2253_,
		_w4917_
	);
	LUT2 #(
		.INIT('h2)
	) name4465 (
		\InstQueue_reg[12][0]/NET0131 ,
		_w2215_,
		_w4918_
	);
	LUT3 #(
		.INIT('h0d)
	) name4466 (
		_w706_,
		_w4914_,
		_w4918_,
		_w4919_
	);
	LUT3 #(
		.INIT('hd0)
	) name4467 (
		_w722_,
		_w4917_,
		_w4919_,
		_w4920_
	);
	LUT2 #(
		.INIT('hb)
	) name4468 (
		_w4916_,
		_w4920_,
		_w4921_
	);
	LUT4 #(
		.INIT('ha600)
	) name4469 (
		\Datai[16]_pad ,
		\Datai[31]_pad ,
		_w2192_,
		_w2239_,
		_w4922_
	);
	LUT4 #(
		.INIT('haa80)
	) name4470 (
		\DataWidth_reg[1]/NET0131 ,
		_w2224_,
		_w4697_,
		_w4922_,
		_w4923_
	);
	LUT4 #(
		.INIT('h5553)
	) name4471 (
		\Datai[0]_pad ,
		\InstQueue_reg[13][0]/NET0131 ,
		_w2187_,
		_w2253_,
		_w4924_
	);
	LUT2 #(
		.INIT('h1)
	) name4472 (
		_w2268_,
		_w4924_,
		_w4925_
	);
	LUT3 #(
		.INIT('ha8)
	) name4473 (
		_w700_,
		_w4923_,
		_w4925_,
		_w4926_
	);
	LUT4 #(
		.INIT('hc055)
	) name4474 (
		\InstQueue_reg[13][0]/NET0131 ,
		_w530_,
		_w535_,
		_w2187_,
		_w4927_
	);
	LUT2 #(
		.INIT('h2)
	) name4475 (
		\InstQueue_reg[13][0]/NET0131 ,
		_w2215_,
		_w4928_
	);
	LUT3 #(
		.INIT('h0d)
	) name4476 (
		_w706_,
		_w4924_,
		_w4928_,
		_w4929_
	);
	LUT3 #(
		.INIT('hd0)
	) name4477 (
		_w722_,
		_w4927_,
		_w4929_,
		_w4930_
	);
	LUT2 #(
		.INIT('hb)
	) name4478 (
		_w4926_,
		_w4930_,
		_w4931_
	);
	LUT4 #(
		.INIT('ha600)
	) name4479 (
		\Datai[16]_pad ,
		\Datai[31]_pad ,
		_w2192_,
		_w2253_,
		_w4932_
	);
	LUT4 #(
		.INIT('haa80)
	) name4480 (
		\DataWidth_reg[1]/NET0131 ,
		_w2239_,
		_w4697_,
		_w4932_,
		_w4933_
	);
	LUT4 #(
		.INIT('h5553)
	) name4481 (
		\Datai[0]_pad ,
		\InstQueue_reg[14][0]/NET0131 ,
		_w2187_,
		_w2203_,
		_w4934_
	);
	LUT2 #(
		.INIT('h1)
	) name4482 (
		_w2279_,
		_w4934_,
		_w4935_
	);
	LUT3 #(
		.INIT('ha8)
	) name4483 (
		_w700_,
		_w4933_,
		_w4935_,
		_w4936_
	);
	LUT4 #(
		.INIT('hc055)
	) name4484 (
		\InstQueue_reg[14][0]/NET0131 ,
		_w530_,
		_w535_,
		_w2203_,
		_w4937_
	);
	LUT2 #(
		.INIT('h2)
	) name4485 (
		\InstQueue_reg[14][0]/NET0131 ,
		_w2215_,
		_w4938_
	);
	LUT3 #(
		.INIT('h0d)
	) name4486 (
		_w706_,
		_w4934_,
		_w4938_,
		_w4939_
	);
	LUT3 #(
		.INIT('hd0)
	) name4487 (
		_w722_,
		_w4937_,
		_w4939_,
		_w4940_
	);
	LUT2 #(
		.INIT('hb)
	) name4488 (
		_w4936_,
		_w4940_,
		_w4941_
	);
	LUT4 #(
		.INIT('ha060)
	) name4489 (
		\Datai[16]_pad ,
		\Datai[31]_pad ,
		_w2187_,
		_w2192_,
		_w4942_
	);
	LUT4 #(
		.INIT('haa80)
	) name4490 (
		\DataWidth_reg[1]/NET0131 ,
		_w2253_,
		_w4697_,
		_w4942_,
		_w4943_
	);
	LUT4 #(
		.INIT('h5553)
	) name4491 (
		\Datai[0]_pad ,
		\InstQueue_reg[15][0]/NET0131 ,
		_w2207_,
		_w2203_,
		_w4944_
	);
	LUT2 #(
		.INIT('h1)
	) name4492 (
		_w2291_,
		_w4944_,
		_w4945_
	);
	LUT3 #(
		.INIT('ha8)
	) name4493 (
		_w700_,
		_w4943_,
		_w4945_,
		_w4946_
	);
	LUT4 #(
		.INIT('hc055)
	) name4494 (
		\InstQueue_reg[15][0]/NET0131 ,
		_w530_,
		_w535_,
		_w2207_,
		_w4947_
	);
	LUT2 #(
		.INIT('h2)
	) name4495 (
		\InstQueue_reg[15][0]/NET0131 ,
		_w2215_,
		_w4948_
	);
	LUT3 #(
		.INIT('h0d)
	) name4496 (
		_w706_,
		_w4944_,
		_w4948_,
		_w4949_
	);
	LUT3 #(
		.INIT('hd0)
	) name4497 (
		_w722_,
		_w4947_,
		_w4949_,
		_w4950_
	);
	LUT2 #(
		.INIT('hb)
	) name4498 (
		_w4946_,
		_w4950_,
		_w4951_
	);
	LUT4 #(
		.INIT('ha060)
	) name4499 (
		\Datai[16]_pad ,
		\Datai[31]_pad ,
		_w2207_,
		_w2192_,
		_w4952_
	);
	LUT4 #(
		.INIT('haa80)
	) name4500 (
		\DataWidth_reg[1]/NET0131 ,
		_w2203_,
		_w4697_,
		_w4952_,
		_w4953_
	);
	LUT4 #(
		.INIT('h5553)
	) name4501 (
		\Datai[0]_pad ,
		\InstQueue_reg[1][0]/NET0131 ,
		_w2205_,
		_w2301_,
		_w4954_
	);
	LUT2 #(
		.INIT('h1)
	) name4502 (
		_w2304_,
		_w4954_,
		_w4955_
	);
	LUT3 #(
		.INIT('ha8)
	) name4503 (
		_w700_,
		_w4953_,
		_w4955_,
		_w4956_
	);
	LUT4 #(
		.INIT('hc055)
	) name4504 (
		\InstQueue_reg[1][0]/NET0131 ,
		_w530_,
		_w535_,
		_w2301_,
		_w4957_
	);
	LUT2 #(
		.INIT('h2)
	) name4505 (
		\InstQueue_reg[1][0]/NET0131 ,
		_w2215_,
		_w4958_
	);
	LUT3 #(
		.INIT('h0d)
	) name4506 (
		_w706_,
		_w4954_,
		_w4958_,
		_w4959_
	);
	LUT3 #(
		.INIT('hd0)
	) name4507 (
		_w722_,
		_w4957_,
		_w4959_,
		_w4960_
	);
	LUT2 #(
		.INIT('hb)
	) name4508 (
		_w4956_,
		_w4960_,
		_w4961_
	);
	LUT4 #(
		.INIT('ha060)
	) name4509 (
		\Datai[16]_pad ,
		\Datai[31]_pad ,
		_w2205_,
		_w2192_,
		_w4962_
	);
	LUT4 #(
		.INIT('haa80)
	) name4510 (
		\DataWidth_reg[1]/NET0131 ,
		_w2207_,
		_w4697_,
		_w4962_,
		_w4963_
	);
	LUT4 #(
		.INIT('h5553)
	) name4511 (
		\Datai[0]_pad ,
		\InstQueue_reg[2][0]/NET0131 ,
		_w2301_,
		_w2314_,
		_w4964_
	);
	LUT2 #(
		.INIT('h1)
	) name4512 (
		_w2317_,
		_w4964_,
		_w4965_
	);
	LUT3 #(
		.INIT('ha8)
	) name4513 (
		_w700_,
		_w4963_,
		_w4965_,
		_w4966_
	);
	LUT4 #(
		.INIT('hc055)
	) name4514 (
		\InstQueue_reg[2][0]/NET0131 ,
		_w530_,
		_w535_,
		_w2314_,
		_w4967_
	);
	LUT2 #(
		.INIT('h2)
	) name4515 (
		\InstQueue_reg[2][0]/NET0131 ,
		_w2215_,
		_w4968_
	);
	LUT3 #(
		.INIT('h0d)
	) name4516 (
		_w706_,
		_w4964_,
		_w4968_,
		_w4969_
	);
	LUT3 #(
		.INIT('hd0)
	) name4517 (
		_w722_,
		_w4967_,
		_w4969_,
		_w4970_
	);
	LUT2 #(
		.INIT('hb)
	) name4518 (
		_w4966_,
		_w4970_,
		_w4971_
	);
	LUT4 #(
		.INIT('ha600)
	) name4519 (
		\Datai[16]_pad ,
		\Datai[31]_pad ,
		_w2192_,
		_w2314_,
		_w4972_
	);
	LUT4 #(
		.INIT('haa80)
	) name4520 (
		\DataWidth_reg[1]/NET0131 ,
		_w2301_,
		_w4697_,
		_w4972_,
		_w4973_
	);
	LUT4 #(
		.INIT('h5553)
	) name4521 (
		\Datai[0]_pad ,
		\InstQueue_reg[4][0]/NET0131 ,
		_w2327_,
		_w2340_,
		_w4974_
	);
	LUT2 #(
		.INIT('h1)
	) name4522 (
		_w2343_,
		_w4974_,
		_w4975_
	);
	LUT3 #(
		.INIT('ha8)
	) name4523 (
		_w700_,
		_w4973_,
		_w4975_,
		_w4976_
	);
	LUT4 #(
		.INIT('hc055)
	) name4524 (
		\InstQueue_reg[4][0]/NET0131 ,
		_w530_,
		_w535_,
		_w2340_,
		_w4977_
	);
	LUT2 #(
		.INIT('h2)
	) name4525 (
		\InstQueue_reg[4][0]/NET0131 ,
		_w2215_,
		_w4978_
	);
	LUT3 #(
		.INIT('h0d)
	) name4526 (
		_w706_,
		_w4974_,
		_w4978_,
		_w4979_
	);
	LUT3 #(
		.INIT('hd0)
	) name4527 (
		_w722_,
		_w4977_,
		_w4979_,
		_w4980_
	);
	LUT2 #(
		.INIT('hb)
	) name4528 (
		_w4976_,
		_w4980_,
		_w4981_
	);
	LUT4 #(
		.INIT('ha600)
	) name4529 (
		\Datai[16]_pad ,
		\Datai[31]_pad ,
		_w2192_,
		_w2327_,
		_w4982_
	);
	LUT4 #(
		.INIT('haa80)
	) name4530 (
		\DataWidth_reg[1]/NET0131 ,
		_w2314_,
		_w4697_,
		_w4982_,
		_w4983_
	);
	LUT4 #(
		.INIT('h5553)
	) name4531 (
		\Datai[0]_pad ,
		\InstQueue_reg[5][0]/NET0131 ,
		_w2340_,
		_w2353_,
		_w4984_
	);
	LUT2 #(
		.INIT('h1)
	) name4532 (
		_w2356_,
		_w4984_,
		_w4985_
	);
	LUT3 #(
		.INIT('ha8)
	) name4533 (
		_w700_,
		_w4983_,
		_w4985_,
		_w4986_
	);
	LUT4 #(
		.INIT('hc055)
	) name4534 (
		\InstQueue_reg[5][0]/NET0131 ,
		_w530_,
		_w535_,
		_w2353_,
		_w4987_
	);
	LUT2 #(
		.INIT('h2)
	) name4535 (
		\InstQueue_reg[5][0]/NET0131 ,
		_w2215_,
		_w4988_
	);
	LUT3 #(
		.INIT('h0d)
	) name4536 (
		_w706_,
		_w4984_,
		_w4988_,
		_w4989_
	);
	LUT3 #(
		.INIT('hd0)
	) name4537 (
		_w722_,
		_w4987_,
		_w4989_,
		_w4990_
	);
	LUT2 #(
		.INIT('hb)
	) name4538 (
		_w4986_,
		_w4990_,
		_w4991_
	);
	LUT4 #(
		.INIT('ha600)
	) name4539 (
		\Datai[16]_pad ,
		\Datai[31]_pad ,
		_w2192_,
		_w2340_,
		_w4992_
	);
	LUT4 #(
		.INIT('haa80)
	) name4540 (
		\DataWidth_reg[1]/NET0131 ,
		_w2327_,
		_w4697_,
		_w4992_,
		_w4993_
	);
	LUT4 #(
		.INIT('h5553)
	) name4541 (
		\Datai[0]_pad ,
		\InstQueue_reg[6][0]/NET0131 ,
		_w2353_,
		_w2366_,
		_w4994_
	);
	LUT2 #(
		.INIT('h1)
	) name4542 (
		_w2369_,
		_w4994_,
		_w4995_
	);
	LUT3 #(
		.INIT('ha8)
	) name4543 (
		_w700_,
		_w4993_,
		_w4995_,
		_w4996_
	);
	LUT4 #(
		.INIT('hc055)
	) name4544 (
		\InstQueue_reg[6][0]/NET0131 ,
		_w530_,
		_w535_,
		_w2366_,
		_w4997_
	);
	LUT2 #(
		.INIT('h2)
	) name4545 (
		\InstQueue_reg[6][0]/NET0131 ,
		_w2215_,
		_w4998_
	);
	LUT3 #(
		.INIT('h0d)
	) name4546 (
		_w706_,
		_w4994_,
		_w4998_,
		_w4999_
	);
	LUT3 #(
		.INIT('hd0)
	) name4547 (
		_w722_,
		_w4997_,
		_w4999_,
		_w5000_
	);
	LUT2 #(
		.INIT('hb)
	) name4548 (
		_w4996_,
		_w5000_,
		_w5001_
	);
	LUT4 #(
		.INIT('ha600)
	) name4549 (
		\Datai[16]_pad ,
		\Datai[31]_pad ,
		_w2192_,
		_w2366_,
		_w5002_
	);
	LUT4 #(
		.INIT('haa80)
	) name4550 (
		\DataWidth_reg[1]/NET0131 ,
		_w2353_,
		_w4697_,
		_w5002_,
		_w5003_
	);
	LUT4 #(
		.INIT('h5553)
	) name4551 (
		\Datai[0]_pad ,
		\InstQueue_reg[8][0]/NET0131 ,
		_w2220_,
		_w2222_,
		_w5004_
	);
	LUT2 #(
		.INIT('h1)
	) name4552 (
		_w2392_,
		_w5004_,
		_w5005_
	);
	LUT3 #(
		.INIT('ha8)
	) name4553 (
		_w700_,
		_w5003_,
		_w5005_,
		_w5006_
	);
	LUT4 #(
		.INIT('hc055)
	) name4554 (
		\InstQueue_reg[8][0]/NET0131 ,
		_w530_,
		_w535_,
		_w2222_,
		_w5007_
	);
	LUT2 #(
		.INIT('h2)
	) name4555 (
		\InstQueue_reg[8][0]/NET0131 ,
		_w2215_,
		_w5008_
	);
	LUT3 #(
		.INIT('h0d)
	) name4556 (
		_w706_,
		_w5004_,
		_w5008_,
		_w5009_
	);
	LUT3 #(
		.INIT('hd0)
	) name4557 (
		_w722_,
		_w5007_,
		_w5009_,
		_w5010_
	);
	LUT2 #(
		.INIT('hb)
	) name4558 (
		_w5006_,
		_w5010_,
		_w5011_
	);
	LUT4 #(
		.INIT('ha600)
	) name4559 (
		\Datai[16]_pad ,
		\Datai[31]_pad ,
		_w2192_,
		_w2220_,
		_w5012_
	);
	LUT4 #(
		.INIT('haa80)
	) name4560 (
		\DataWidth_reg[1]/NET0131 ,
		_w2366_,
		_w4697_,
		_w5012_,
		_w5013_
	);
	LUT4 #(
		.INIT('h5553)
	) name4561 (
		\Datai[0]_pad ,
		\InstQueue_reg[9][0]/NET0131 ,
		_w2225_,
		_w2222_,
		_w5014_
	);
	LUT2 #(
		.INIT('h1)
	) name4562 (
		_w2403_,
		_w5014_,
		_w5015_
	);
	LUT3 #(
		.INIT('ha8)
	) name4563 (
		_w700_,
		_w5013_,
		_w5015_,
		_w5016_
	);
	LUT4 #(
		.INIT('hc055)
	) name4564 (
		\InstQueue_reg[9][0]/NET0131 ,
		_w530_,
		_w535_,
		_w2225_,
		_w5017_
	);
	LUT2 #(
		.INIT('h2)
	) name4565 (
		\InstQueue_reg[9][0]/NET0131 ,
		_w2215_,
		_w5018_
	);
	LUT3 #(
		.INIT('h0d)
	) name4566 (
		_w706_,
		_w5014_,
		_w5018_,
		_w5019_
	);
	LUT3 #(
		.INIT('hd0)
	) name4567 (
		_w722_,
		_w5017_,
		_w5019_,
		_w5020_
	);
	LUT2 #(
		.INIT('hb)
	) name4568 (
		_w5016_,
		_w5020_,
		_w5021_
	);
	LUT3 #(
		.INIT('h48)
	) name4569 (
		\rEIP_reg[6]/NET0131 ,
		_w615_,
		_w4549_,
		_w5022_
	);
	LUT3 #(
		.INIT('h8a)
	) name4570 (
		\Address[4]_pad ,
		\State_reg[0]/NET0131 ,
		\State_reg[1]/NET0131 ,
		_w5023_
	);
	LUT3 #(
		.INIT('h80)
	) name4571 (
		\rEIP_reg[0]/NET0131 ,
		\rEIP_reg[1]/NET0131 ,
		\rEIP_reg[31]/NET0131 ,
		_w5024_
	);
	LUT4 #(
		.INIT('h8000)
	) name4572 (
		\rEIP_reg[0]/NET0131 ,
		\rEIP_reg[1]/NET0131 ,
		\rEIP_reg[2]/NET0131 ,
		\rEIP_reg[31]/NET0131 ,
		_w5025_
	);
	LUT3 #(
		.INIT('h80)
	) name4573 (
		\rEIP_reg[3]/NET0131 ,
		\rEIP_reg[4]/NET0131 ,
		_w5025_,
		_w5026_
	);
	LUT4 #(
		.INIT('h8000)
	) name4574 (
		\rEIP_reg[3]/NET0131 ,
		\rEIP_reg[4]/NET0131 ,
		\rEIP_reg[5]/NET0131 ,
		_w5025_,
		_w5027_
	);
	LUT4 #(
		.INIT('h0b07)
	) name4575 (
		\rEIP_reg[5]/NET0131 ,
		_w4565_,
		_w5023_,
		_w5026_,
		_w5028_
	);
	LUT2 #(
		.INIT('hb)
	) name4576 (
		_w5022_,
		_w5028_,
		_w5029_
	);
	LUT4 #(
		.INIT('h4888)
	) name4577 (
		\rEIP_reg[29]/NET0131 ,
		_w615_,
		_w2620_,
		_w4559_,
		_w5030_
	);
	LUT3 #(
		.INIT('h8a)
	) name4578 (
		\Address[27]_pad ,
		\State_reg[0]/NET0131 ,
		\State_reg[1]/NET0131 ,
		_w5031_
	);
	LUT4 #(
		.INIT('h1333)
	) name4579 (
		\rEIP_reg[27]/NET0131 ,
		\rEIP_reg[28]/NET0131 ,
		_w2618_,
		_w4563_,
		_w5032_
	);
	LUT4 #(
		.INIT('h70f0)
	) name4580 (
		_w2618_,
		_w2620_,
		_w4565_,
		_w4563_,
		_w5033_
	);
	LUT3 #(
		.INIT('h45)
	) name4581 (
		_w5031_,
		_w5032_,
		_w5033_,
		_w5034_
	);
	LUT2 #(
		.INIT('hb)
	) name4582 (
		_w5030_,
		_w5034_,
		_w5035_
	);
	LUT3 #(
		.INIT('h45)
	) name4583 (
		\Address[15]_pad ,
		\State_reg[0]/NET0131 ,
		\State_reg[1]/NET0131 ,
		_w5036_
	);
	LUT4 #(
		.INIT('hd070)
	) name4584 (
		\State_reg[2]/NET0131 ,
		\rEIP_reg[16]/NET0131 ,
		_w614_,
		_w4602_,
		_w5037_
	);
	LUT4 #(
		.INIT('heb00)
	) name4585 (
		\State_reg[2]/NET0131 ,
		\rEIP_reg[17]/NET0131 ,
		_w4556_,
		_w5037_,
		_w5038_
	);
	LUT2 #(
		.INIT('h1)
	) name4586 (
		_w5036_,
		_w5038_,
		_w5039_
	);
	LUT4 #(
		.INIT('h1333)
	) name4587 (
		\rEIP_reg[24]/NET0131 ,
		\rEIP_reg[25]/NET0131 ,
		_w2605_,
		_w4557_,
		_w5040_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name4588 (
		_w615_,
		_w2605_,
		_w2617_,
		_w4557_,
		_w5041_
	);
	LUT3 #(
		.INIT('h8a)
	) name4589 (
		\Address[23]_pad ,
		\State_reg[0]/NET0131 ,
		\State_reg[1]/NET0131 ,
		_w5042_
	);
	LUT4 #(
		.INIT('h60a0)
	) name4590 (
		\rEIP_reg[24]/NET0131 ,
		_w2616_,
		_w4565_,
		_w4562_,
		_w5043_
	);
	LUT4 #(
		.INIT('hefee)
	) name4591 (
		_w5042_,
		_w5043_,
		_w5040_,
		_w5041_,
		_w5044_
	);
	LUT4 #(
		.INIT('h60c0)
	) name4592 (
		\rEIP_reg[12]/NET0131 ,
		\rEIP_reg[13]/NET0131 ,
		_w615_,
		_w4553_,
		_w5045_
	);
	LUT3 #(
		.INIT('h8a)
	) name4593 (
		\Address[11]_pad ,
		\State_reg[0]/NET0131 ,
		\State_reg[1]/NET0131 ,
		_w5046_
	);
	LUT4 #(
		.INIT('h9300)
	) name4594 (
		\rEIP_reg[11]/NET0131 ,
		\rEIP_reg[12]/NET0131 ,
		_w2608_,
		_w4562_,
		_w5047_
	);
	LUT3 #(
		.INIT('h13)
	) name4595 (
		\rEIP_reg[0]/NET0131 ,
		\rEIP_reg[12]/NET0131 ,
		\rEIP_reg[31]/NET0131 ,
		_w5048_
	);
	LUT2 #(
		.INIT('h2)
	) name4596 (
		_w4565_,
		_w5048_,
		_w5049_
	);
	LUT3 #(
		.INIT('h45)
	) name4597 (
		_w5046_,
		_w5047_,
		_w5049_,
		_w5050_
	);
	LUT2 #(
		.INIT('hb)
	) name4598 (
		_w5045_,
		_w5050_,
		_w5051_
	);
	LUT3 #(
		.INIT('h48)
	) name4599 (
		\rEIP_reg[5]/NET0131 ,
		_w615_,
		_w4548_,
		_w5052_
	);
	LUT3 #(
		.INIT('h8a)
	) name4600 (
		\Address[3]_pad ,
		\State_reg[0]/NET0131 ,
		\State_reg[1]/NET0131 ,
		_w5053_
	);
	LUT4 #(
		.INIT('h60c0)
	) name4601 (
		\rEIP_reg[3]/NET0131 ,
		\rEIP_reg[4]/NET0131 ,
		_w4565_,
		_w5025_,
		_w5054_
	);
	LUT2 #(
		.INIT('h1)
	) name4602 (
		_w5053_,
		_w5054_,
		_w5055_
	);
	LUT2 #(
		.INIT('hb)
	) name4603 (
		_w5052_,
		_w5055_,
		_w5056_
	);
	LUT4 #(
		.INIT('h070f)
	) name4604 (
		\rEIP_reg[19]/NET0131 ,
		\rEIP_reg[20]/NET0131 ,
		\rEIP_reg[21]/NET0131 ,
		_w4598_,
		_w5057_
	);
	LUT2 #(
		.INIT('h2)
	) name4605 (
		_w615_,
		_w4557_,
		_w5058_
	);
	LUT3 #(
		.INIT('h8a)
	) name4606 (
		\Address[19]_pad ,
		\State_reg[0]/NET0131 ,
		\State_reg[1]/NET0131 ,
		_w5059_
	);
	LUT4 #(
		.INIT('h00b7)
	) name4607 (
		\rEIP_reg[20]/NET0131 ,
		_w4565_,
		_w4880_,
		_w5059_,
		_w5060_
	);
	LUT3 #(
		.INIT('h4f)
	) name4608 (
		_w5057_,
		_w5058_,
		_w5060_,
		_w5061_
	);
	LUT3 #(
		.INIT('h48)
	) name4609 (
		\rEIP_reg[9]/NET0131 ,
		_w615_,
		_w4551_,
		_w5062_
	);
	LUT3 #(
		.INIT('h8a)
	) name4610 (
		\Address[7]_pad ,
		\State_reg[0]/NET0131 ,
		\State_reg[1]/NET0131 ,
		_w5063_
	);
	LUT4 #(
		.INIT('h60c0)
	) name4611 (
		\rEIP_reg[7]/NET0131 ,
		\rEIP_reg[8]/NET0131 ,
		_w4565_,
		_w4887_,
		_w5064_
	);
	LUT2 #(
		.INIT('h1)
	) name4612 (
		_w5063_,
		_w5064_,
		_w5065_
	);
	LUT2 #(
		.INIT('hb)
	) name4613 (
		_w5062_,
		_w5065_,
		_w5066_
	);
	LUT4 #(
		.INIT('h60c0)
	) name4614 (
		\rEIP_reg[15]/NET0131 ,
		\rEIP_reg[16]/NET0131 ,
		_w615_,
		_w4555_,
		_w5067_
	);
	LUT3 #(
		.INIT('h8a)
	) name4615 (
		\Address[14]_pad ,
		\State_reg[0]/NET0131 ,
		\State_reg[1]/NET0131 ,
		_w5068_
	);
	LUT4 #(
		.INIT('h00b7)
	) name4616 (
		\rEIP_reg[15]/NET0131 ,
		_w4565_,
		_w4601_,
		_w5068_,
		_w5069_
	);
	LUT2 #(
		.INIT('hb)
	) name4617 (
		_w5067_,
		_w5069_,
		_w5070_
	);
	LUT4 #(
		.INIT('h60c0)
	) name4618 (
		\rEIP_reg[27]/NET0131 ,
		\rEIP_reg[28]/NET0131 ,
		_w615_,
		_w4559_,
		_w5071_
	);
	LUT3 #(
		.INIT('h8a)
	) name4619 (
		\Address[26]_pad ,
		\State_reg[0]/NET0131 ,
		\State_reg[1]/NET0131 ,
		_w5072_
	);
	LUT4 #(
		.INIT('h60a0)
	) name4620 (
		\rEIP_reg[27]/NET0131 ,
		_w2618_,
		_w4565_,
		_w4563_,
		_w5073_
	);
	LUT2 #(
		.INIT('h1)
	) name4621 (
		_w5072_,
		_w5073_,
		_w5074_
	);
	LUT2 #(
		.INIT('hb)
	) name4622 (
		_w5071_,
		_w5074_,
		_w5075_
	);
	LUT4 #(
		.INIT('h4888)
	) name4623 (
		\rEIP_reg[24]/NET0131 ,
		_w615_,
		_w2605_,
		_w4557_,
		_w5076_
	);
	LUT3 #(
		.INIT('h8a)
	) name4624 (
		\Address[22]_pad ,
		\State_reg[0]/NET0131 ,
		\State_reg[1]/NET0131 ,
		_w5077_
	);
	LUT4 #(
		.INIT('h8000)
	) name4625 (
		\rEIP_reg[22]/NET0131 ,
		_w2611_,
		_w2615_,
		_w4562_,
		_w5078_
	);
	LUT4 #(
		.INIT('h0c08)
	) name4626 (
		\rEIP_reg[23]/NET0131 ,
		_w4565_,
		_w4563_,
		_w5078_,
		_w5079_
	);
	LUT3 #(
		.INIT('hfe)
	) name4627 (
		_w5077_,
		_w5079_,
		_w5076_,
		_w5080_
	);
	LUT3 #(
		.INIT('h48)
	) name4628 (
		\rEIP_reg[12]/NET0131 ,
		_w615_,
		_w4553_,
		_w5081_
	);
	LUT3 #(
		.INIT('h8a)
	) name4629 (
		\Address[10]_pad ,
		\State_reg[0]/NET0131 ,
		\State_reg[1]/NET0131 ,
		_w5082_
	);
	LUT3 #(
		.INIT('h13)
	) name4630 (
		\rEIP_reg[0]/NET0131 ,
		\rEIP_reg[11]/NET0131 ,
		\rEIP_reg[31]/NET0131 ,
		_w5083_
	);
	LUT2 #(
		.INIT('h2)
	) name4631 (
		_w4565_,
		_w5083_,
		_w5084_
	);
	LUT4 #(
		.INIT('h6f00)
	) name4632 (
		\rEIP_reg[11]/NET0131 ,
		_w2608_,
		_w4562_,
		_w5084_,
		_w5085_
	);
	LUT2 #(
		.INIT('h1)
	) name4633 (
		_w5082_,
		_w5085_,
		_w5086_
	);
	LUT2 #(
		.INIT('hb)
	) name4634 (
		_w5081_,
		_w5086_,
		_w5087_
	);
	LUT4 #(
		.INIT('h60c0)
	) name4635 (
		\rEIP_reg[3]/NET0131 ,
		\rEIP_reg[4]/NET0131 ,
		_w615_,
		_w4547_,
		_w5088_
	);
	LUT3 #(
		.INIT('h8a)
	) name4636 (
		\Address[2]_pad ,
		\State_reg[0]/NET0131 ,
		\State_reg[1]/NET0131 ,
		_w5089_
	);
	LUT4 #(
		.INIT('h00b7)
	) name4637 (
		\rEIP_reg[3]/NET0131 ,
		_w4565_,
		_w5025_,
		_w5089_,
		_w5090_
	);
	LUT2 #(
		.INIT('hb)
	) name4638 (
		_w5088_,
		_w5090_,
		_w5091_
	);
	LUT4 #(
		.INIT('h60c0)
	) name4639 (
		\rEIP_reg[19]/NET0131 ,
		\rEIP_reg[20]/NET0131 ,
		_w615_,
		_w4598_,
		_w5092_
	);
	LUT3 #(
		.INIT('h8a)
	) name4640 (
		\Address[18]_pad ,
		\State_reg[0]/NET0131 ,
		\State_reg[1]/NET0131 ,
		_w5093_
	);
	LUT4 #(
		.INIT('h8000)
	) name4641 (
		\rEIP_reg[16]/NET0131 ,
		\rEIP_reg[17]/NET0131 ,
		\rEIP_reg[18]/NET0131 ,
		_w4602_,
		_w5094_
	);
	LUT4 #(
		.INIT('h70f0)
	) name4642 (
		_w2611_,
		_w2613_,
		_w4565_,
		_w4562_,
		_w5095_
	);
	LUT4 #(
		.INIT('h0133)
	) name4643 (
		\rEIP_reg[19]/NET0131 ,
		_w5093_,
		_w5094_,
		_w5095_,
		_w5096_
	);
	LUT2 #(
		.INIT('hb)
	) name4644 (
		_w5092_,
		_w5096_,
		_w5097_
	);
	LUT3 #(
		.INIT('h8a)
	) name4645 (
		\Address[6]_pad ,
		\State_reg[0]/NET0131 ,
		\State_reg[1]/NET0131 ,
		_w5098_
	);
	LUT4 #(
		.INIT('h00b7)
	) name4646 (
		\rEIP_reg[7]/NET0131 ,
		_w4565_,
		_w4887_,
		_w5098_,
		_w5099_
	);
	LUT4 #(
		.INIT('h48ff)
	) name4647 (
		\rEIP_reg[8]/NET0131 ,
		_w615_,
		_w4550_,
		_w5099_,
		_w5100_
	);
	LUT3 #(
		.INIT('h48)
	) name4648 (
		\rEIP_reg[27]/NET0131 ,
		_w615_,
		_w4559_,
		_w5101_
	);
	LUT3 #(
		.INIT('h8a)
	) name4649 (
		\Address[25]_pad ,
		\State_reg[0]/NET0131 ,
		\State_reg[1]/NET0131 ,
		_w5102_
	);
	LUT4 #(
		.INIT('h1333)
	) name4650 (
		\rEIP_reg[25]/NET0131 ,
		\rEIP_reg[26]/NET0131 ,
		_w3263_,
		_w4562_,
		_w5103_
	);
	LUT3 #(
		.INIT('h4c)
	) name4651 (
		_w2618_,
		_w4565_,
		_w4563_,
		_w5104_
	);
	LUT3 #(
		.INIT('h45)
	) name4652 (
		_w5102_,
		_w5103_,
		_w5104_,
		_w5105_
	);
	LUT2 #(
		.INIT('hb)
	) name4653 (
		_w5101_,
		_w5105_,
		_w5106_
	);
	LUT4 #(
		.INIT('h4888)
	) name4654 (
		\rEIP_reg[31]/NET0131 ,
		_w615_,
		_w2622_,
		_w4559_,
		_w5107_
	);
	LUT3 #(
		.INIT('h8a)
	) name4655 (
		\Address[29]_pad ,
		\State_reg[0]/NET0131 ,
		\State_reg[1]/NET0131 ,
		_w5108_
	);
	LUT4 #(
		.INIT('h8000)
	) name4656 (
		\rEIP_reg[0]/NET0131 ,
		\rEIP_reg[31]/NET0131 ,
		_w2619_,
		_w2622_,
		_w5109_
	);
	LUT4 #(
		.INIT('h1555)
	) name4657 (
		\rEIP_reg[30]/NET0131 ,
		_w2618_,
		_w2621_,
		_w4563_,
		_w5110_
	);
	LUT4 #(
		.INIT('h3331)
	) name4658 (
		_w4565_,
		_w5108_,
		_w5110_,
		_w5109_,
		_w5111_
	);
	LUT2 #(
		.INIT('hb)
	) name4659 (
		_w5107_,
		_w5111_,
		_w5112_
	);
	LUT3 #(
		.INIT('h48)
	) name4660 (
		\rEIP_reg[15]/NET0131 ,
		_w615_,
		_w4555_,
		_w5113_
	);
	LUT3 #(
		.INIT('h8a)
	) name4661 (
		\Address[13]_pad ,
		\State_reg[0]/NET0131 ,
		\State_reg[1]/NET0131 ,
		_w5114_
	);
	LUT4 #(
		.INIT('h60a0)
	) name4662 (
		\rEIP_reg[14]/NET0131 ,
		_w2610_,
		_w4565_,
		_w4562_,
		_w5115_
	);
	LUT2 #(
		.INIT('h1)
	) name4663 (
		_w5114_,
		_w5115_,
		_w5116_
	);
	LUT2 #(
		.INIT('hb)
	) name4664 (
		_w5113_,
		_w5116_,
		_w5117_
	);
	LUT3 #(
		.INIT('h8a)
	) name4665 (
		\Address[9]_pad ,
		\State_reg[0]/NET0131 ,
		\State_reg[1]/NET0131 ,
		_w5118_
	);
	LUT4 #(
		.INIT('h00b7)
	) name4666 (
		\rEIP_reg[10]/NET0131 ,
		_w4565_,
		_w4889_,
		_w5118_,
		_w5119_
	);
	LUT4 #(
		.INIT('h48ff)
	) name4667 (
		\rEIP_reg[11]/NET0131 ,
		_w615_,
		_w4552_,
		_w5119_,
		_w5120_
	);
	LUT4 #(
		.INIT('h60c0)
	) name4668 (
		\rEIP_reg[22]/NET0131 ,
		\rEIP_reg[23]/NET0131 ,
		_w615_,
		_w4557_,
		_w5121_
	);
	LUT3 #(
		.INIT('h8a)
	) name4669 (
		\Address[21]_pad ,
		\State_reg[0]/NET0131 ,
		\State_reg[1]/NET0131 ,
		_w5122_
	);
	LUT4 #(
		.INIT('h1555)
	) name4670 (
		\rEIP_reg[22]/NET0131 ,
		_w2611_,
		_w2615_,
		_w4562_,
		_w5123_
	);
	LUT4 #(
		.INIT('h0f0d)
	) name4671 (
		_w4565_,
		_w5078_,
		_w5122_,
		_w5123_,
		_w5124_
	);
	LUT2 #(
		.INIT('hb)
	) name4672 (
		_w5121_,
		_w5124_,
		_w5125_
	);
	LUT2 #(
		.INIT('h7)
	) name4673 (
		\DataWidth_reg[0]/NET0131 ,
		\DataWidth_reg[1]/NET0131 ,
		_w5126_
	);
	LUT3 #(
		.INIT('h80)
	) name4674 (
		\ByteEnable_reg[2]/NET0131 ,
		\DataWidth_reg[0]/NET0131 ,
		\DataWidth_reg[1]/NET0131 ,
		_w5127_
	);
	LUT4 #(
		.INIT('h7013)
	) name4675 (
		\DataWidth_reg[0]/NET0131 ,
		\DataWidth_reg[1]/NET0131 ,
		\rEIP_reg[0]/NET0131 ,
		\rEIP_reg[1]/NET0131 ,
		_w5128_
	);
	LUT2 #(
		.INIT('he)
	) name4676 (
		_w5127_,
		_w5128_,
		_w5129_
	);
	LUT4 #(
		.INIT('h3310)
	) name4677 (
		HOLD_pad,
		READY_n_pad,
		\State_reg[0]/NET0131 ,
		\State_reg[2]/NET0131 ,
		_w5130_
	);
	LUT4 #(
		.INIT('h40c0)
	) name4678 (
		HOLD_pad,
		\RequestPending_reg/NET0131 ,
		\State_reg[0]/NET0131 ,
		\State_reg[2]/NET0131 ,
		_w5131_
	);
	LUT4 #(
		.INIT('hfcfe)
	) name4679 (
		\State_reg[1]/NET0131 ,
		_w616_,
		_w5131_,
		_w5130_,
		_w5132_
	);
	LUT3 #(
		.INIT('h01)
	) name4680 (
		\DataWidth_reg[0]/NET0131 ,
		\DataWidth_reg[1]/NET0131 ,
		\rEIP_reg[0]/NET0131 ,
		_w5133_
	);
	LUT4 #(
		.INIT('h407f)
	) name4681 (
		\ByteEnable_reg[1]/NET0131 ,
		\DataWidth_reg[0]/NET0131 ,
		\DataWidth_reg[1]/NET0131 ,
		\rEIP_reg[1]/NET0131 ,
		_w5134_
	);
	LUT2 #(
		.INIT('hb)
	) name4682 (
		_w5133_,
		_w5134_,
		_w5135_
	);
	LUT4 #(
		.INIT('h0acf)
	) name4683 (
		NA_n_pad,
		READY_n_pad,
		\State_reg[0]/NET0131 ,
		\State_reg[2]/NET0131 ,
		_w5136_
	);
	LUT3 #(
		.INIT('h02)
	) name4684 (
		\State_reg[0]/NET0131 ,
		\State_reg[1]/NET0131 ,
		\State_reg[2]/NET0131 ,
		_w5137_
	);
	LUT4 #(
		.INIT('hcc04)
	) name4685 (
		HOLD_pad,
		\RequestPending_reg/NET0131 ,
		_w5136_,
		_w5137_,
		_w5138_
	);
	LUT2 #(
		.INIT('h1)
	) name4686 (
		_w4565_,
		_w5138_,
		_w5139_
	);
	LUT3 #(
		.INIT('h48)
	) name4687 (
		\rEIP_reg[3]/NET0131 ,
		_w615_,
		_w4547_,
		_w5140_
	);
	LUT3 #(
		.INIT('h8a)
	) name4688 (
		\Address[1]_pad ,
		\State_reg[0]/NET0131 ,
		\State_reg[1]/NET0131 ,
		_w5141_
	);
	LUT4 #(
		.INIT('h00b7)
	) name4689 (
		\rEIP_reg[2]/NET0131 ,
		_w4565_,
		_w5024_,
		_w5141_,
		_w5142_
	);
	LUT2 #(
		.INIT('hb)
	) name4690 (
		_w5140_,
		_w5142_,
		_w5143_
	);
	LUT3 #(
		.INIT('h48)
	) name4691 (
		\rEIP_reg[19]/NET0131 ,
		_w615_,
		_w4598_,
		_w5144_
	);
	LUT3 #(
		.INIT('h8a)
	) name4692 (
		\Address[17]_pad ,
		\State_reg[0]/NET0131 ,
		\State_reg[1]/NET0131 ,
		_w5145_
	);
	LUT4 #(
		.INIT('h00b7)
	) name4693 (
		\rEIP_reg[18]/NET0131 ,
		_w4565_,
		_w4603_,
		_w5145_,
		_w5146_
	);
	LUT2 #(
		.INIT('hb)
	) name4694 (
		_w5144_,
		_w5146_,
		_w5147_
	);
	LUT4 #(
		.INIT('h60c0)
	) name4695 (
		\rEIP_reg[6]/NET0131 ,
		\rEIP_reg[7]/NET0131 ,
		_w615_,
		_w4549_,
		_w5148_
	);
	LUT3 #(
		.INIT('h8a)
	) name4696 (
		\Address[5]_pad ,
		\State_reg[0]/NET0131 ,
		\State_reg[1]/NET0131 ,
		_w5149_
	);
	LUT4 #(
		.INIT('h0c08)
	) name4697 (
		\rEIP_reg[6]/NET0131 ,
		_w4565_,
		_w4887_,
		_w5027_,
		_w5150_
	);
	LUT3 #(
		.INIT('hfe)
	) name4698 (
		_w5149_,
		_w5150_,
		_w5148_,
		_w5151_
	);
	LUT3 #(
		.INIT('h08)
	) name4699 (
		\State_reg[0]/NET0131 ,
		\State_reg[1]/NET0131 ,
		\State_reg[2]/NET0131 ,
		_w5152_
	);
	LUT3 #(
		.INIT('hc8)
	) name4700 (
		HOLD_pad,
		READY_n_pad,
		\RequestPending_reg/NET0131 ,
		_w5153_
	);
	LUT4 #(
		.INIT('h5444)
	) name4701 (
		NA_n_pad,
		_w616_,
		_w5152_,
		_w5153_,
		_w5154_
	);
	LUT3 #(
		.INIT('h0e)
	) name4702 (
		\RequestPending_reg/NET0131 ,
		\State_reg[1]/NET0131 ,
		\State_reg[2]/NET0131 ,
		_w5155_
	);
	LUT2 #(
		.INIT('h8)
	) name4703 (
		HOLD_pad,
		\State_reg[0]/NET0131 ,
		_w5156_
	);
	LUT4 #(
		.INIT('hb000)
	) name4704 (
		READY_n_pad,
		\State_reg[0]/NET0131 ,
		\State_reg[1]/NET0131 ,
		\State_reg[2]/NET0131 ,
		_w5157_
	);
	LUT3 #(
		.INIT('h0b)
	) name4705 (
		_w5155_,
		_w5156_,
		_w5157_,
		_w5158_
	);
	LUT2 #(
		.INIT('hb)
	) name4706 (
		_w5154_,
		_w5158_,
		_w5159_
	);
	LUT3 #(
		.INIT('h80)
	) name4707 (
		\ByteEnable_reg[3]/NET0131 ,
		\DataWidth_reg[0]/NET0131 ,
		\DataWidth_reg[1]/NET0131 ,
		_w5160_
	);
	LUT4 #(
		.INIT('h0133)
	) name4708 (
		\DataWidth_reg[0]/NET0131 ,
		\DataWidth_reg[1]/NET0131 ,
		\rEIP_reg[0]/NET0131 ,
		\rEIP_reg[1]/NET0131 ,
		_w5161_
	);
	LUT2 #(
		.INIT('he)
	) name4709 (
		_w5160_,
		_w5161_,
		_w5162_
	);
	LUT3 #(
		.INIT('h48)
	) name4710 (
		\rEIP_reg[2]/NET0131 ,
		_w615_,
		_w4546_,
		_w5163_
	);
	LUT3 #(
		.INIT('h8a)
	) name4711 (
		\Address[0]_pad ,
		\State_reg[0]/NET0131 ,
		\State_reg[1]/NET0131 ,
		_w5164_
	);
	LUT4 #(
		.INIT('h00b7)
	) name4712 (
		\rEIP_reg[1]/NET0131 ,
		_w4565_,
		_w4562_,
		_w5164_,
		_w5165_
	);
	LUT2 #(
		.INIT('hb)
	) name4713 (
		_w5163_,
		_w5165_,
		_w5166_
	);
	LUT4 #(
		.INIT('h5414)
	) name4714 (
		\DataWidth_reg[1]/NET0131 ,
		\State_reg[0]/NET0131 ,
		\State_reg[1]/NET0131 ,
		\State_reg[2]/NET0131 ,
		_w5167_
	);
	LUT4 #(
		.INIT('h0140)
	) name4715 (
		\BS16_n_pad ,
		\State_reg[0]/NET0131 ,
		\State_reg[1]/NET0131 ,
		\State_reg[2]/NET0131 ,
		_w5168_
	);
	LUT2 #(
		.INIT('h1)
	) name4716 (
		_w5167_,
		_w5168_,
		_w5169_
	);
	LUT4 #(
		.INIT('h8bcb)
	) name4717 (
		ADS_n_pad,
		\State_reg[0]/NET0131 ,
		\State_reg[1]/NET0131 ,
		\State_reg[2]/NET0131 ,
		_w5170_
	);
	LUT4 #(
		.INIT('hacaa)
	) name4718 (
		\BE_n[2]_pad ,
		\ByteEnable_reg[2]/NET0131 ,
		\State_reg[0]/NET0131 ,
		\State_reg[1]/NET0131 ,
		_w5171_
	);
	LUT4 #(
		.INIT('hacaa)
	) name4719 (
		\BE_n[0]_pad ,
		\ByteEnable_reg[0]/NET0131 ,
		\State_reg[0]/NET0131 ,
		\State_reg[1]/NET0131 ,
		_w5172_
	);
	LUT4 #(
		.INIT('hacaa)
	) name4720 (
		\BE_n[1]_pad ,
		\ByteEnable_reg[1]/NET0131 ,
		\State_reg[0]/NET0131 ,
		\State_reg[1]/NET0131 ,
		_w5173_
	);
	LUT4 #(
		.INIT('hacaa)
	) name4721 (
		\BE_n[3]_pad ,
		\ByteEnable_reg[3]/NET0131 ,
		\State_reg[0]/NET0131 ,
		\State_reg[1]/NET0131 ,
		_w5174_
	);
	LUT4 #(
		.INIT('hdf10)
	) name4722 (
		\ReadRequest_reg/NET0131 ,
		\State_reg[0]/NET0131 ,
		\State_reg[1]/NET0131 ,
		W_R_n_pad,
		_w5175_
	);
	LUT4 #(
		.INIT('hacaa)
	) name4723 (
		M_IO_n_pad,
		\MemoryFetch_reg/NET0131 ,
		\State_reg[0]/NET0131 ,
		\State_reg[1]/NET0131 ,
		_w5176_
	);
	LUT4 #(
		.INIT('h4544)
	) name4724 (
		D_C_n_pad,
		\State_reg[0]/NET0131 ,
		\State_reg[1]/NET0131 ,
		\State_reg[2]/NET0131 ,
		_w5177_
	);
	LUT3 #(
		.INIT('h20)
	) name4725 (
		\CodeFetch_reg/NET0131 ,
		\State_reg[0]/NET0131 ,
		\State_reg[1]/NET0131 ,
		_w5178_
	);
	LUT2 #(
		.INIT('h1)
	) name4726 (
		_w5177_,
		_w5178_,
		_w5179_
	);
	LUT4 #(
		.INIT('ha828)
	) name4727 (
		\DataWidth_reg[0]/NET0131 ,
		\State_reg[0]/NET0131 ,
		\State_reg[1]/NET0131 ,
		\State_reg[2]/NET0131 ,
		_w5180_
	);
	LUT2 #(
		.INIT('he)
	) name4728 (
		_w5168_,
		_w5180_,
		_w5181_
	);
	LUT2 #(
		.INIT('h2)
	) name4729 (
		\InstAddrPointer_reg[13]/NET0131 ,
		_w681_,
		_w5182_
	);
	LUT3 #(
		.INIT('h6a)
	) name4730 (
		\InstAddrPointer_reg[13]/NET0131 ,
		_w727_,
		_w864_,
		_w5183_
	);
	LUT3 #(
		.INIT('h70)
	) name4731 (
		_w731_,
		_w933_,
		_w5183_,
		_w5184_
	);
	LUT4 #(
		.INIT('hb0f0)
	) name4732 (
		\InstAddrPointer_reg[13]/NET0131 ,
		_w731_,
		_w844_,
		_w933_,
		_w5185_
	);
	LUT2 #(
		.INIT('h4)
	) name4733 (
		_w5184_,
		_w5185_,
		_w5186_
	);
	LUT2 #(
		.INIT('h2)
	) name4734 (
		_w985_,
		_w1349_,
		_w5187_
	);
	LUT3 #(
		.INIT('h15)
	) name4735 (
		_w844_,
		_w1127_,
		_w1129_,
		_w5188_
	);
	LUT3 #(
		.INIT('h8a)
	) name4736 (
		_w681_,
		_w5187_,
		_w5188_,
		_w5189_
	);
	LUT4 #(
		.INIT('h8a88)
	) name4737 (
		_w574_,
		_w5182_,
		_w5186_,
		_w5189_,
		_w5190_
	);
	LUT3 #(
		.INIT('h80)
	) name4738 (
		_w1054_,
		_w1061_,
		_w1066_,
		_w5191_
	);
	LUT4 #(
		.INIT('h8000)
	) name4739 (
		_w1054_,
		_w1062_,
		_w1061_,
		_w1066_,
		_w5192_
	);
	LUT4 #(
		.INIT('h1333)
	) name4740 (
		_w1054_,
		_w1062_,
		_w1061_,
		_w1066_,
		_w5193_
	);
	LUT3 #(
		.INIT('h02)
	) name4741 (
		_w688_,
		_w5193_,
		_w5192_,
		_w5194_
	);
	LUT2 #(
		.INIT('h2)
	) name4742 (
		\InstAddrPointer_reg[13]/NET0131 ,
		_w1220_,
		_w5195_
	);
	LUT2 #(
		.INIT('h4)
	) name4743 (
		_w645_,
		_w5183_,
		_w5196_
	);
	LUT2 #(
		.INIT('h8)
	) name4744 (
		_w606_,
		_w1062_,
		_w5197_
	);
	LUT4 #(
		.INIT('h004f)
	) name4745 (
		_w582_,
		_w595_,
		_w985_,
		_w5197_,
		_w5198_
	);
	LUT3 #(
		.INIT('h10)
	) name4746 (
		_w5195_,
		_w5196_,
		_w5198_,
		_w5199_
	);
	LUT2 #(
		.INIT('h4)
	) name4747 (
		_w5194_,
		_w5199_,
		_w5200_
	);
	LUT2 #(
		.INIT('h8)
	) name4748 (
		\rEIP_reg[13]/NET0131 ,
		_w1109_,
		_w5201_
	);
	LUT4 #(
		.INIT('h3f15)
	) name4749 (
		\InstAddrPointer_reg[13]/NET0131 ,
		\rEIP_reg[13]/NET0131 ,
		_w1109_,
		_w1110_,
		_w5202_
	);
	LUT4 #(
		.INIT('h8aff)
	) name4750 (
		_w695_,
		_w5190_,
		_w5200_,
		_w5202_,
		_w5203_
	);
	LUT2 #(
		.INIT('h2)
	) name4751 (
		\InstAddrPointer_reg[16]/NET0131 ,
		_w681_,
		_w5204_
	);
	LUT4 #(
		.INIT('haa20)
	) name4752 (
		_w574_,
		_w1647_,
		_w1648_,
		_w5204_,
		_w5205_
	);
	LUT4 #(
		.INIT('h00ec)
	) name4753 (
		_w514_,
		_w566_,
		_w569_,
		_w904_,
		_w5206_
	);
	LUT3 #(
		.INIT('h08)
	) name4754 (
		_w613_,
		_w636_,
		_w5206_,
		_w5207_
	);
	LUT4 #(
		.INIT('h8000)
	) name4755 (
		\InstAddrPointer_reg[15]/NET0131 ,
		_w611_,
		_w633_,
		_w866_,
		_w5208_
	);
	LUT2 #(
		.INIT('h2)
	) name4756 (
		\InstAddrPointer_reg[16]/NET0131 ,
		_w5208_,
		_w5209_
	);
	LUT4 #(
		.INIT('h00f7)
	) name4757 (
		_w612_,
		_w903_,
		_w1381_,
		_w5209_,
		_w5210_
	);
	LUT2 #(
		.INIT('h1)
	) name4758 (
		_w5207_,
		_w5210_,
		_w5211_
	);
	LUT3 #(
		.INIT('hb0)
	) name4759 (
		_w582_,
		_w595_,
		_w991_,
		_w5212_
	);
	LUT2 #(
		.INIT('h2)
	) name4760 (
		_w549_,
		_w904_,
		_w5213_
	);
	LUT2 #(
		.INIT('h1)
	) name4761 (
		\InstAddrPointer_reg[16]/NET0131 ,
		_w605_,
		_w5214_
	);
	LUT4 #(
		.INIT('hc800)
	) name4762 (
		_w552_,
		_w576_,
		_w579_,
		_w1188_,
		_w5215_
	);
	LUT4 #(
		.INIT('h0f0e)
	) name4763 (
		_w625_,
		_w683_,
		_w5214_,
		_w5215_,
		_w5216_
	);
	LUT2 #(
		.INIT('h1)
	) name4764 (
		_w5213_,
		_w5216_,
		_w5217_
	);
	LUT3 #(
		.INIT('h10)
	) name4765 (
		_w5212_,
		_w5211_,
		_w5217_,
		_w5218_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name4766 (
		_w695_,
		_w1652_,
		_w5205_,
		_w5218_,
		_w5219_
	);
	LUT4 #(
		.INIT('h3f15)
	) name4767 (
		\InstAddrPointer_reg[16]/NET0131 ,
		\rEIP_reg[16]/NET0131 ,
		_w1109_,
		_w1110_,
		_w5220_
	);
	LUT2 #(
		.INIT('hb)
	) name4768 (
		_w5219_,
		_w5220_,
		_w5221_
	);
	LUT2 #(
		.INIT('h2)
	) name4769 (
		\InstAddrPointer_reg[17]/NET0131 ,
		_w681_,
		_w5222_
	);
	LUT4 #(
		.INIT('haa20)
	) name4770 (
		_w574_,
		_w1667_,
		_w1670_,
		_w5222_,
		_w5223_
	);
	LUT4 #(
		.INIT('h2111)
	) name4771 (
		\InstAddrPointer_reg[17]/NET0131 ,
		READY_n_pad,
		_w727_,
		_w871_,
		_w5224_
	);
	LUT4 #(
		.INIT('h00f4)
	) name4772 (
		_w514_,
		_w569_,
		_w570_,
		_w5224_,
		_w5225_
	);
	LUT4 #(
		.INIT('h0001)
	) name4773 (
		_w683_,
		_w1195_,
		_w1196_,
		_w5225_,
		_w5226_
	);
	LUT2 #(
		.INIT('h2)
	) name4774 (
		\InstAddrPointer_reg[17]/NET0131 ,
		_w5226_,
		_w5227_
	);
	LUT3 #(
		.INIT('hb0)
	) name4775 (
		_w582_,
		_w595_,
		_w993_,
		_w5228_
	);
	LUT4 #(
		.INIT('h9aaa)
	) name4776 (
		\InstAddrPointer_reg[17]/NET0131 ,
		READY_n_pad,
		_w727_,
		_w871_,
		_w5229_
	);
	LUT4 #(
		.INIT('h8a00)
	) name4777 (
		_w611_,
		_w618_,
		_w619_,
		_w5229_,
		_w5230_
	);
	LUT2 #(
		.INIT('h8)
	) name4778 (
		_w549_,
		_w906_,
		_w5231_
	);
	LUT3 #(
		.INIT('h84)
	) name4779 (
		\InstAddrPointer_reg[17]/NET0131 ,
		_w605_,
		_w1068_,
		_w5232_
	);
	LUT2 #(
		.INIT('h1)
	) name4780 (
		\InstAddrPointer_reg[17]/NET0131 ,
		_w605_,
		_w5233_
	);
	LUT4 #(
		.INIT('h00c8)
	) name4781 (
		_w552_,
		_w576_,
		_w579_,
		_w5233_,
		_w5234_
	);
	LUT3 #(
		.INIT('h45)
	) name4782 (
		_w5231_,
		_w5232_,
		_w5234_,
		_w5235_
	);
	LUT2 #(
		.INIT('h4)
	) name4783 (
		_w5230_,
		_w5235_,
		_w5236_
	);
	LUT4 #(
		.INIT('h0100)
	) name4784 (
		_w1672_,
		_w5227_,
		_w5228_,
		_w5236_,
		_w5237_
	);
	LUT4 #(
		.INIT('h3f15)
	) name4785 (
		\InstAddrPointer_reg[17]/NET0131 ,
		\rEIP_reg[17]/NET0131 ,
		_w1109_,
		_w1110_,
		_w5238_
	);
	LUT4 #(
		.INIT('h8aff)
	) name4786 (
		_w695_,
		_w5223_,
		_w5237_,
		_w5238_,
		_w5239_
	);
	LUT2 #(
		.INIT('h2)
	) name4787 (
		\InstAddrPointer_reg[10]/NET0131 ,
		_w681_,
		_w5240_
	);
	LUT3 #(
		.INIT('ha8)
	) name4788 (
		_w574_,
		_w1757_,
		_w5240_,
		_w5241_
	);
	LUT4 #(
		.INIT('h8088)
	) name4789 (
		\InstAddrPointer_reg[10]/NET0131 ,
		_w611_,
		_w618_,
		_w619_,
		_w5242_
	);
	LUT3 #(
		.INIT('hc4)
	) name4790 (
		_w620_,
		_w1524_,
		_w5242_,
		_w5243_
	);
	LUT3 #(
		.INIT('ha2)
	) name4791 (
		\InstAddrPointer_reg[10]/NET0131 ,
		_w1197_,
		_w1514_,
		_w5244_
	);
	LUT2 #(
		.INIT('h8)
	) name4792 (
		_w606_,
		_w1148_,
		_w5245_
	);
	LUT4 #(
		.INIT('h004f)
	) name4793 (
		_w582_,
		_w595_,
		_w971_,
		_w5245_,
		_w5246_
	);
	LUT3 #(
		.INIT('h10)
	) name4794 (
		_w5244_,
		_w5243_,
		_w5246_,
		_w5247_
	);
	LUT2 #(
		.INIT('h4)
	) name4795 (
		_w1760_,
		_w5247_,
		_w5248_
	);
	LUT4 #(
		.INIT('h3f15)
	) name4796 (
		\InstAddrPointer_reg[10]/NET0131 ,
		\rEIP_reg[10]/NET0131 ,
		_w1109_,
		_w1110_,
		_w5249_
	);
	LUT4 #(
		.INIT('h8aff)
	) name4797 (
		_w695_,
		_w5241_,
		_w5248_,
		_w5249_,
		_w5250_
	);
	LUT4 #(
		.INIT('h60c0)
	) name4798 (
		\EBX_reg[29]/NET0131 ,
		\EBX_reg[30]/NET0131 ,
		_w590_,
		_w3769_,
		_w5251_
	);
	LUT2 #(
		.INIT('h8)
	) name4799 (
		\EBX_reg[30]/NET0131 ,
		_w1975_,
		_w5252_
	);
	LUT3 #(
		.INIT('h90)
	) name4800 (
		_w1941_,
		_w1952_,
		_w1973_,
		_w5253_
	);
	LUT2 #(
		.INIT('h1)
	) name4801 (
		_w5252_,
		_w5253_,
		_w5254_
	);
	LUT2 #(
		.INIT('h2)
	) name4802 (
		\EBX_reg[30]/NET0131 ,
		_w1825_,
		_w5255_
	);
	LUT4 #(
		.INIT('hff8a)
	) name4803 (
		_w695_,
		_w5251_,
		_w5254_,
		_w5255_,
		_w5256_
	);
	LUT4 #(
		.INIT('h111d)
	) name4804 (
		\InstAddrPointer_reg[26]/NET0131 ,
		_w681_,
		_w1615_,
		_w1618_,
		_w5257_
	);
	LUT4 #(
		.INIT('h00c8)
	) name4805 (
		_w552_,
		_w576_,
		_w579_,
		_w1080_,
		_w5258_
	);
	LUT4 #(
		.INIT('haa2a)
	) name4806 (
		\InstAddrPointer_reg[26]/NET0131 ,
		_w624_,
		_w684_,
		_w5258_,
		_w5259_
	);
	LUT2 #(
		.INIT('h4)
	) name4807 (
		_w620_,
		_w882_,
		_w5260_
	);
	LUT2 #(
		.INIT('h8)
	) name4808 (
		_w606_,
		_w1081_,
		_w5261_
	);
	LUT4 #(
		.INIT('h00f4)
	) name4809 (
		_w582_,
		_w595_,
		_w1010_,
		_w5261_,
		_w5262_
	);
	LUT3 #(
		.INIT('h10)
	) name4810 (
		_w5259_,
		_w5260_,
		_w5262_,
		_w5263_
	);
	LUT2 #(
		.INIT('h4)
	) name4811 (
		_w1621_,
		_w5263_,
		_w5264_
	);
	LUT4 #(
		.INIT('h08cc)
	) name4812 (
		_w574_,
		_w695_,
		_w5257_,
		_w5264_,
		_w5265_
	);
	LUT4 #(
		.INIT('h3f15)
	) name4813 (
		\InstAddrPointer_reg[26]/NET0131 ,
		\rEIP_reg[26]/NET0131 ,
		_w1109_,
		_w1110_,
		_w5266_
	);
	LUT2 #(
		.INIT('hb)
	) name4814 (
		_w5265_,
		_w5266_,
		_w5267_
	);
	LUT4 #(
		.INIT('h4888)
	) name4815 (
		\EAX_reg[30]/NET0131 ,
		_w1848_,
		_w1845_,
		_w1846_,
		_w5268_
	);
	LUT3 #(
		.INIT('h8a)
	) name4816 (
		\EAX_reg[30]/NET0131 ,
		_w635_,
		_w1852_,
		_w5269_
	);
	LUT3 #(
		.INIT('h82)
	) name4817 (
		_w1849_,
		_w1941_,
		_w1952_,
		_w5270_
	);
	LUT3 #(
		.INIT('h80)
	) name4818 (
		\Datai[30]_pad ,
		_w514_,
		_w569_,
		_w5271_
	);
	LUT3 #(
		.INIT('ha8)
	) name4819 (
		_w612_,
		_w3756_,
		_w5271_,
		_w5272_
	);
	LUT2 #(
		.INIT('h1)
	) name4820 (
		_w5270_,
		_w5272_,
		_w5273_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name4821 (
		_w695_,
		_w5268_,
		_w5269_,
		_w5273_,
		_w5274_
	);
	LUT2 #(
		.INIT('h2)
	) name4822 (
		\EAX_reg[30]/NET0131 ,
		_w1825_,
		_w5275_
	);
	LUT2 #(
		.INIT('he)
	) name4823 (
		_w5274_,
		_w5275_,
		_w5276_
	);
	LUT4 #(
		.INIT('h8000)
	) name4824 (
		\EBX_reg[27]/NET0131 ,
		\EBX_reg[28]/NET0131 ,
		\EBX_reg[29]/NET0131 ,
		\EBX_reg[30]/NET0131 ,
		_w5277_
	);
	LUT3 #(
		.INIT('h80)
	) name4825 (
		_w1958_,
		_w1972_,
		_w5277_,
		_w5278_
	);
	LUT2 #(
		.INIT('h8)
	) name4826 (
		\EBX_reg[31]/NET0131 ,
		_w1975_,
		_w5279_
	);
	LUT3 #(
		.INIT('h20)
	) name4827 (
		_w1941_,
		_w1952_,
		_w1973_,
		_w5280_
	);
	LUT2 #(
		.INIT('h1)
	) name4828 (
		_w5279_,
		_w5280_,
		_w5281_
	);
	LUT4 #(
		.INIT('hb700)
	) name4829 (
		\EBX_reg[31]/NET0131 ,
		_w590_,
		_w5278_,
		_w5281_,
		_w5282_
	);
	LUT2 #(
		.INIT('h2)
	) name4830 (
		\EBX_reg[31]/NET0131 ,
		_w1825_,
		_w5283_
	);
	LUT3 #(
		.INIT('hf2)
	) name4831 (
		_w695_,
		_w5282_,
		_w5283_,
		_w5284_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name4832 (
		\Datao_reg[22]/NET0131 ,
		_w695_,
		_w2159_,
		_w2422_,
		_w5285_
	);
	LUT2 #(
		.INIT('h8)
	) name4833 (
		\uWord_reg[6]/NET0131 ,
		_w696_,
		_w5286_
	);
	LUT3 #(
		.INIT('h20)
	) name4834 (
		_w611_,
		_w617_,
		_w695_,
		_w5287_
	);
	LUT4 #(
		.INIT('h0200)
	) name4835 (
		_w570_,
		_w2048_,
		_w3979_,
		_w5287_,
		_w5288_
	);
	LUT2 #(
		.INIT('h1)
	) name4836 (
		_w5286_,
		_w5288_,
		_w5289_
	);
	LUT2 #(
		.INIT('hb)
	) name4837 (
		_w5285_,
		_w5289_,
		_w5290_
	);
	LUT4 #(
		.INIT('hddd1)
	) name4838 (
		\InstAddrPointer_reg[7]/NET0131 ,
		_w681_,
		_w1772_,
		_w1771_,
		_w5291_
	);
	LUT2 #(
		.INIT('h2)
	) name4839 (
		_w574_,
		_w5291_,
		_w5292_
	);
	LUT2 #(
		.INIT('h2)
	) name4840 (
		\InstAddrPointer_reg[7]/NET0131 ,
		_w1220_,
		_w5293_
	);
	LUT2 #(
		.INIT('h4)
	) name4841 (
		_w645_,
		_w832_,
		_w5294_
	);
	LUT2 #(
		.INIT('h8)
	) name4842 (
		_w606_,
		_w1045_,
		_w5295_
	);
	LUT4 #(
		.INIT('h004f)
	) name4843 (
		_w582_,
		_w595_,
		_w943_,
		_w5295_,
		_w5296_
	);
	LUT4 #(
		.INIT('h0100)
	) name4844 (
		_w1778_,
		_w5294_,
		_w5293_,
		_w5296_,
		_w5297_
	);
	LUT4 #(
		.INIT('h3f15)
	) name4845 (
		\InstAddrPointer_reg[7]/NET0131 ,
		\rEIP_reg[7]/NET0131 ,
		_w1109_,
		_w1110_,
		_w5298_
	);
	LUT4 #(
		.INIT('h8aff)
	) name4846 (
		_w695_,
		_w5292_,
		_w5297_,
		_w5298_,
		_w5299_
	);
	LUT4 #(
		.INIT('h8222)
	) name4847 (
		_w844_,
		_w1412_,
		_w1416_,
		_w1418_,
		_w5300_
	);
	LUT4 #(
		.INIT('h4111)
	) name4848 (
		_w844_,
		_w1007_,
		_w1349_,
		_w1351_,
		_w5301_
	);
	LUT4 #(
		.INIT('hddd1)
	) name4849 (
		\PhyAddrPointer_reg[21]/NET0131 ,
		_w681_,
		_w5301_,
		_w5300_,
		_w5302_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name4850 (
		\InstAddrPointer_reg[20]/NET0131 ,
		\InstAddrPointer_reg[21]/NET0131 ,
		_w874_,
		_w1068_,
		_w5303_
	);
	LUT4 #(
		.INIT('h8000)
	) name4851 (
		_w1054_,
		_w1067_,
		_w1070_,
		_w1072_,
		_w5304_
	);
	LUT4 #(
		.INIT('h2220)
	) name4852 (
		_w688_,
		_w1074_,
		_w5303_,
		_w5304_,
		_w5305_
	);
	LUT4 #(
		.INIT('h028a)
	) name4853 (
		\PhyAddrPointer_reg[21]/NET0131 ,
		_w573_,
		_w574_,
		_w605_,
		_w5306_
	);
	LUT4 #(
		.INIT('h0031)
	) name4854 (
		_w574_,
		_w5305_,
		_w5302_,
		_w5306_,
		_w5307_
	);
	LUT3 #(
		.INIT('h02)
	) name4855 (
		_w1281_,
		_w1462_,
		_w3203_,
		_w5308_
	);
	LUT4 #(
		.INIT('hc444)
	) name4856 (
		_w707_,
		_w1283_,
		_w1269_,
		_w1569_,
		_w5309_
	);
	LUT3 #(
		.INIT('h20)
	) name4857 (
		\DataWidth_reg[1]/NET0131 ,
		\PhyAddrPointer_reg[21]/NET0131 ,
		_w700_,
		_w5310_
	);
	LUT2 #(
		.INIT('h8)
	) name4858 (
		\rEIP_reg[21]/NET0131 ,
		_w1109_,
		_w5311_
	);
	LUT4 #(
		.INIT('h007f)
	) name4859 (
		_w1269_,
		_w1569_,
		_w5310_,
		_w5311_,
		_w5312_
	);
	LUT3 #(
		.INIT('hd0)
	) name4860 (
		\PhyAddrPointer_reg[21]/NET0131 ,
		_w5309_,
		_w5312_,
		_w5313_
	);
	LUT2 #(
		.INIT('h4)
	) name4861 (
		_w5308_,
		_w5313_,
		_w5314_
	);
	LUT3 #(
		.INIT('h2f)
	) name4862 (
		_w695_,
		_w5307_,
		_w5314_,
		_w5315_
	);
	LUT2 #(
		.INIT('h2)
	) name4863 (
		\InstAddrPointer_reg[15]/NET0131 ,
		_w681_,
		_w5316_
	);
	LUT4 #(
		.INIT('haa20)
	) name4864 (
		_w574_,
		_w1439_,
		_w1441_,
		_w5316_,
		_w5317_
	);
	LUT4 #(
		.INIT('h1511)
	) name4865 (
		\InstAddrPointer_reg[15]/NET0131 ,
		_w612_,
		_w618_,
		_w619_,
		_w5318_
	);
	LUT4 #(
		.INIT('h8000)
	) name4866 (
		_w492_,
		_w515_,
		_w536_,
		_w565_,
		_w5319_
	);
	LUT3 #(
		.INIT('h0e)
	) name4867 (
		_w571_,
		_w5318_,
		_w5319_,
		_w5320_
	);
	LUT4 #(
		.INIT('hec00)
	) name4868 (
		_w613_,
		_w634_,
		_w636_,
		_w901_,
		_w5321_
	);
	LUT2 #(
		.INIT('h1)
	) name4869 (
		_w900_,
		_w5321_,
		_w5322_
	);
	LUT2 #(
		.INIT('h2)
	) name4870 (
		\InstAddrPointer_reg[15]/NET0131 ,
		_w605_,
		_w5323_
	);
	LUT4 #(
		.INIT('h9333)
	) name4871 (
		\InstAddrPointer_reg[14]/NET0131 ,
		\InstAddrPointer_reg[15]/NET0131 ,
		_w605_,
		_w1056_,
		_w5324_
	);
	LUT4 #(
		.INIT('h00c8)
	) name4872 (
		_w552_,
		_w576_,
		_w579_,
		_w5324_,
		_w5325_
	);
	LUT2 #(
		.INIT('h8)
	) name4873 (
		_w573_,
		_w5323_,
		_w5326_
	);
	LUT3 #(
		.INIT('h20)
	) name4874 (
		_w549_,
		_w564_,
		_w902_,
		_w5327_
	);
	LUT3 #(
		.INIT('h01)
	) name4875 (
		_w5326_,
		_w5325_,
		_w5327_,
		_w5328_
	);
	LUT4 #(
		.INIT('h4f00)
	) name4876 (
		_w582_,
		_w595_,
		_w988_,
		_w5328_,
		_w5329_
	);
	LUT3 #(
		.INIT('hb0)
	) name4877 (
		_w5320_,
		_w5322_,
		_w5329_,
		_w5330_
	);
	LUT2 #(
		.INIT('h4)
	) name4878 (
		_w1447_,
		_w5330_,
		_w5331_
	);
	LUT4 #(
		.INIT('h3f15)
	) name4879 (
		\InstAddrPointer_reg[15]/NET0131 ,
		\rEIP_reg[15]/NET0131 ,
		_w1109_,
		_w1110_,
		_w5332_
	);
	LUT4 #(
		.INIT('h8aff)
	) name4880 (
		_w695_,
		_w5317_,
		_w5331_,
		_w5332_,
		_w5333_
	);
	LUT2 #(
		.INIT('h2)
	) name4881 (
		\PhyAddrPointer_reg[13]/NET0131 ,
		_w681_,
		_w5334_
	);
	LUT4 #(
		.INIT('haa20)
	) name4882 (
		_w574_,
		_w5186_,
		_w5189_,
		_w5334_,
		_w5335_
	);
	LUT4 #(
		.INIT('h028a)
	) name4883 (
		\PhyAddrPointer_reg[13]/NET0131 ,
		_w573_,
		_w574_,
		_w605_,
		_w5336_
	);
	LUT4 #(
		.INIT('h00d7)
	) name4884 (
		_w688_,
		_w1062_,
		_w5191_,
		_w5336_,
		_w5337_
	);
	LUT2 #(
		.INIT('h8)
	) name4885 (
		_w1281_,
		_w3565_,
		_w5338_
	);
	LUT4 #(
		.INIT('hb030)
	) name4886 (
		\PhyAddrPointer_reg[12]/NET0131 ,
		_w707_,
		_w1283_,
		_w1263_,
		_w5339_
	);
	LUT3 #(
		.INIT('h20)
	) name4887 (
		\DataWidth_reg[1]/NET0131 ,
		\PhyAddrPointer_reg[13]/NET0131 ,
		_w700_,
		_w5340_
	);
	LUT4 #(
		.INIT('h070f)
	) name4888 (
		\PhyAddrPointer_reg[12]/NET0131 ,
		_w1263_,
		_w5201_,
		_w5340_,
		_w5341_
	);
	LUT3 #(
		.INIT('hd0)
	) name4889 (
		\PhyAddrPointer_reg[13]/NET0131 ,
		_w5339_,
		_w5341_,
		_w5342_
	);
	LUT2 #(
		.INIT('h4)
	) name4890 (
		_w5338_,
		_w5342_,
		_w5343_
	);
	LUT4 #(
		.INIT('h8aff)
	) name4891 (
		_w695_,
		_w5335_,
		_w5337_,
		_w5343_,
		_w5344_
	);
	LUT2 #(
		.INIT('h2)
	) name4892 (
		\EAX_reg[27]/NET0131 ,
		_w1825_,
		_w5345_
	);
	LUT4 #(
		.INIT('h0b03)
	) name4893 (
		\EAX_reg[26]/NET0131 ,
		_w1848_,
		_w1851_,
		_w2029_,
		_w5346_
	);
	LUT2 #(
		.INIT('h4)
	) name4894 (
		\EAX_reg[27]/NET0131 ,
		_w1848_,
		_w5347_
	);
	LUT4 #(
		.INIT('h3533)
	) name4895 (
		\Datai[27]_pad ,
		\EAX_reg[27]/NET0131 ,
		READY_n_pad,
		_w611_,
		_w5348_
	);
	LUT3 #(
		.INIT('h08)
	) name4896 (
		_w514_,
		_w569_,
		_w5348_,
		_w5349_
	);
	LUT4 #(
		.INIT('h3533)
	) name4897 (
		\Datai[11]_pad ,
		\EAX_reg[27]/NET0131 ,
		READY_n_pad,
		_w611_,
		_w5350_
	);
	LUT2 #(
		.INIT('h2)
	) name4898 (
		_w566_,
		_w5350_,
		_w5351_
	);
	LUT4 #(
		.INIT('h0007)
	) name4899 (
		_w1849_,
		_w1977_,
		_w5351_,
		_w5349_,
		_w5352_
	);
	LUT4 #(
		.INIT('h7f00)
	) name4900 (
		\EAX_reg[26]/NET0131 ,
		_w2029_,
		_w5347_,
		_w5352_,
		_w5353_
	);
	LUT4 #(
		.INIT('h08cc)
	) name4901 (
		\EAX_reg[27]/NET0131 ,
		_w695_,
		_w5346_,
		_w5353_,
		_w5354_
	);
	LUT2 #(
		.INIT('he)
	) name4902 (
		_w5345_,
		_w5354_,
		_w5355_
	);
	LUT2 #(
		.INIT('h2)
	) name4903 (
		\PhyAddrPointer_reg[9]/NET0131 ,
		_w681_,
		_w5356_
	);
	LUT4 #(
		.INIT('h028a)
	) name4904 (
		\PhyAddrPointer_reg[9]/NET0131 ,
		_w573_,
		_w574_,
		_w605_,
		_w5357_
	);
	LUT4 #(
		.INIT('h00d7)
	) name4905 (
		_w688_,
		_w1054_,
		_w1065_,
		_w5357_,
		_w5358_
	);
	LUT4 #(
		.INIT('h5700)
	) name4906 (
		_w574_,
		_w1636_,
		_w5356_,
		_w5358_,
		_w5359_
	);
	LUT4 #(
		.INIT('h6c00)
	) name4907 (
		\PhyAddrPointer_reg[1]/NET0131 ,
		\PhyAddrPointer_reg[9]/NET0131 ,
		_w1261_,
		_w1281_,
		_w5360_
	);
	LUT4 #(
		.INIT('h3f15)
	) name4908 (
		\PhyAddrPointer_reg[9]/NET0131 ,
		\rEIP_reg[9]/NET0131 ,
		_w1109_,
		_w1283_,
		_w5361_
	);
	LUT4 #(
		.INIT('hb700)
	) name4909 (
		\PhyAddrPointer_reg[9]/NET0131 ,
		_w707_,
		_w1261_,
		_w5361_,
		_w5362_
	);
	LUT2 #(
		.INIT('h4)
	) name4910 (
		_w5360_,
		_w5362_,
		_w5363_
	);
	LUT3 #(
		.INIT('h2f)
	) name4911 (
		_w695_,
		_w5359_,
		_w5363_,
		_w5364_
	);
	LUT2 #(
		.INIT('h2)
	) name4912 (
		\PhyAddrPointer_reg[12]/NET0131 ,
		_w681_,
		_w5365_
	);
	LUT4 #(
		.INIT('haa20)
	) name4913 (
		_w574_,
		_w1526_,
		_w1530_,
		_w5365_,
		_w5366_
	);
	LUT4 #(
		.INIT('h028a)
	) name4914 (
		\PhyAddrPointer_reg[12]/NET0131 ,
		_w573_,
		_w574_,
		_w605_,
		_w5367_
	);
	LUT2 #(
		.INIT('h1)
	) name4915 (
		_w1532_,
		_w5367_,
		_w5368_
	);
	LUT4 #(
		.INIT('h4111)
	) name4916 (
		\DataWidth_reg[1]/NET0131 ,
		\PhyAddrPointer_reg[12]/NET0131 ,
		\PhyAddrPointer_reg[1]/NET0131 ,
		_w1263_,
		_w5369_
	);
	LUT4 #(
		.INIT('h70d0)
	) name4917 (
		\DataWidth_reg[1]/NET0131 ,
		\PhyAddrPointer_reg[12]/NET0131 ,
		_w700_,
		_w1263_,
		_w5370_
	);
	LUT4 #(
		.INIT('h60a0)
	) name4918 (
		\PhyAddrPointer_reg[12]/NET0131 ,
		\PhyAddrPointer_reg[1]/NET0131 ,
		_w706_,
		_w1263_,
		_w5371_
	);
	LUT4 #(
		.INIT('h3f15)
	) name4919 (
		\PhyAddrPointer_reg[12]/NET0131 ,
		\rEIP_reg[12]/NET0131 ,
		_w1109_,
		_w1283_,
		_w5372_
	);
	LUT4 #(
		.INIT('h4500)
	) name4920 (
		_w5371_,
		_w5369_,
		_w5370_,
		_w5372_,
		_w5373_
	);
	LUT4 #(
		.INIT('h8aff)
	) name4921 (
		_w695_,
		_w5366_,
		_w5368_,
		_w5373_,
		_w5374_
	);
	LUT2 #(
		.INIT('h2)
	) name4922 (
		\InstAddrPointer_reg[18]/NET0131 ,
		_w681_,
		_w5375_
	);
	LUT3 #(
		.INIT('ha8)
	) name4923 (
		_w574_,
		_w1685_,
		_w5375_,
		_w5376_
	);
	LUT3 #(
		.INIT('h8a)
	) name4924 (
		\InstAddrPointer_reg[18]/NET0131 ,
		_w637_,
		_w684_,
		_w5377_
	);
	LUT2 #(
		.INIT('h4)
	) name4925 (
		_w645_,
		_w909_,
		_w5378_
	);
	LUT2 #(
		.INIT('h8)
	) name4926 (
		_w606_,
		_w1152_,
		_w5379_
	);
	LUT4 #(
		.INIT('h004f)
	) name4927 (
		_w582_,
		_w595_,
		_w992_,
		_w5379_,
		_w5380_
	);
	LUT3 #(
		.INIT('h10)
	) name4928 (
		_w5377_,
		_w5378_,
		_w5380_,
		_w5381_
	);
	LUT2 #(
		.INIT('h4)
	) name4929 (
		_w1689_,
		_w5381_,
		_w5382_
	);
	LUT4 #(
		.INIT('h3f15)
	) name4930 (
		\InstAddrPointer_reg[18]/NET0131 ,
		\rEIP_reg[18]/NET0131 ,
		_w1109_,
		_w1110_,
		_w5383_
	);
	LUT4 #(
		.INIT('h8aff)
	) name4931 (
		_w695_,
		_w5376_,
		_w5382_,
		_w5383_,
		_w5384_
	);
	LUT4 #(
		.INIT('hddd1)
	) name4932 (
		\InstAddrPointer_reg[21]/NET0131 ,
		_w681_,
		_w5301_,
		_w5300_,
		_w5385_
	);
	LUT4 #(
		.INIT('h00c8)
	) name4933 (
		_w552_,
		_w576_,
		_w579_,
		_w1071_,
		_w5386_
	);
	LUT4 #(
		.INIT('haa8a)
	) name4934 (
		\InstAddrPointer_reg[21]/NET0131 ,
		_w637_,
		_w684_,
		_w5386_,
		_w5387_
	);
	LUT3 #(
		.INIT('hb0)
	) name4935 (
		_w582_,
		_w595_,
		_w1007_,
		_w5388_
	);
	LUT2 #(
		.INIT('h8)
	) name4936 (
		_w606_,
		_w5303_,
		_w5389_
	);
	LUT3 #(
		.INIT('h0b)
	) name4937 (
		_w645_,
		_w1412_,
		_w5389_,
		_w5390_
	);
	LUT3 #(
		.INIT('h10)
	) name4938 (
		_w5387_,
		_w5388_,
		_w5390_,
		_w5391_
	);
	LUT4 #(
		.INIT('h3100)
	) name4939 (
		_w574_,
		_w5305_,
		_w5385_,
		_w5391_,
		_w5392_
	);
	LUT4 #(
		.INIT('h3f15)
	) name4940 (
		\InstAddrPointer_reg[21]/NET0131 ,
		\rEIP_reg[21]/NET0131 ,
		_w1109_,
		_w1110_,
		_w5393_
	);
	LUT3 #(
		.INIT('h2f)
	) name4941 (
		_w695_,
		_w5392_,
		_w5393_,
		_w5394_
	);
	assign \_al_n0  = 1'b0;
	assign \_al_n1  = 1'b1;
	assign \g47521/_2_  = _w704_ ;
	assign \g47523/_0_  = _w711_ ;
	assign \g47526/_0_  = _w721_ ;
	assign \g47529/_0_  = _w723_ ;
	assign \g47533/_0_  = _w1112_ ;
	assign \g47540/_0_  = _w1166_ ;
	assign \g47551/_0_  = _w1207_ ;
	assign \g47552/_0_  = _w1230_ ;
	assign \g47553/_0_  = _w1253_ ;
	assign \g47563/_2_  = _w1286_ ;
	assign \g47566/_0_  = _w1307_ ;
	assign \g47567/_0_  = _w1321_ ;
	assign \g47568/_0_  = _w1337_ ;
	assign \g47569/_0_  = _w1365_ ;
	assign \g47583/_2_  = _w1375_ ;
	assign \g47584/_0_  = _w1396_ ;
	assign \g47585/_0_  = _w1410_ ;
	assign \g47589/_0_  = _w1436_ ;
	assign \g47602/_0_  = _w1457_ ;
	assign \g47603/_0_  = _w1470_ ;
	assign \g47604/_2_  = _w1480_ ;
	assign \g47605/_0_  = _w1489_ ;
	assign \g47606/_2_  = _w1508_ ;
	assign \g47609/_0_  = _w1521_ ;
	assign \g47611/_0_  = _w1544_ ;
	assign \g47631/_0_  = _w1555_ ;
	assign \g47632/_0_  = _w1564_ ;
	assign \g47633/_0_  = _w1578_ ;
	assign \g47635/_0_  = _w1592_ ;
	assign \g47636/_0_  = _w1602_ ;
	assign \g47637/_0_  = _w1613_ ;
	assign \g47638/_2_  = _w1632_ ;
	assign \g47643/_0_  = _w1645_ ;
	assign \g47665/_2_  = _w1665_ ;
	assign \g47666/_0_  = _w1681_ ;
	assign \g47667/_0_  = _w1697_ ;
	assign \g47670/_0_  = _w1707_ ;
	assign \g47672/_0_  = _w1719_ ;
	assign \g47677/_0_  = _w1736_ ;
	assign \g47678/_0_  = _w1752_ ;
	assign \g47706/_0_  = _w1770_ ;
	assign \g47711/_0_  = _w1788_ ;
	assign \g47717/_0_  = _w1811_ ;
	assign \g47718/_0_  = _w1823_ ;
	assign \g47721/_0_  = _w1957_ ;
	assign \g47722/_0_  = _w1983_ ;
	assign \g47751/_0_  = _w1995_ ;
	assign \g47755/_0_  = _w2016_ ;
	assign \g47756/_0_  = _w2027_ ;
	assign \g47757/_0_  = _w2038_ ;
	assign \g47759/_0_  = _w2060_ ;
	assign \g47789/_0_  = _w2066_ ;
	assign \g47793/_0_  = _w2071_ ;
	assign \g47797/_0_  = _w2083_ ;
	assign \g47798/_0_  = _w2094_ ;
	assign \g47799/_0_  = _w2104_ ;
	assign \g47802/_0_  = _w2120_ ;
	assign \g47804/_0_  = _w2126_ ;
	assign \g47807/_0_  = _w2139_ ;
	assign \g47809/_0_  = _w2148_ ;
	assign \g47862/_0_  = _w2161_ ;
	assign \g47863/_0_  = _w2167_ ;
	assign \g47864/_0_  = _w2173_ ;
	assign \g47869/_0_  = _w2179_ ;
	assign \g47870/_0_  = _w2185_ ;
	assign \g47924/_0_  = _w2219_ ;
	assign \g47925/_0_  = _w2236_ ;
	assign \g47926/_0_  = _w2250_ ;
	assign \g47927/_0_  = _w2263_ ;
	assign \g47928/_0_  = _w2275_ ;
	assign \g47930/_0_  = _w2286_ ;
	assign \g47932/_0_  = _w2298_ ;
	assign \g47933/_0_  = _w2311_ ;
	assign \g47934/_0_  = _w2324_ ;
	assign \g47935/_0_  = _w2337_ ;
	assign \g47936/_0_  = _w2350_ ;
	assign \g47937/_0_  = _w2363_ ;
	assign \g47938/_0_  = _w2376_ ;
	assign \g47939/_0_  = _w2388_ ;
	assign \g47940/_0_  = _w2399_ ;
	assign \g47941/_0_  = _w2410_ ;
	assign \g47957/_0_  = _w2417_ ;
	assign \g47970/_0_  = _w2425_ ;
	assign \g47973/_0_  = _w2430_ ;
	assign \g47975/_0_  = _w2442_ ;
	assign \g48058/_0_  = _w2454_ ;
	assign \g48059/_0_  = _w2464_ ;
	assign \g48060/_0_  = _w2474_ ;
	assign \g48061/_0_  = _w2484_ ;
	assign \g48062/_0_  = _w2494_ ;
	assign \g48064/_0_  = _w2504_ ;
	assign \g48065/_0_  = _w2514_ ;
	assign \g48066/_0_  = _w2524_ ;
	assign \g48067/_0_  = _w2534_ ;
	assign \g48068/_0_  = _w2544_ ;
	assign \g48069/_0_  = _w2554_ ;
	assign \g48070/_0_  = _w2564_ ;
	assign \g48071/_0_  = _w2574_ ;
	assign \g48072/_0_  = _w2584_ ;
	assign \g48073/_0_  = _w2594_ ;
	assign \g48074/_0_  = _w2604_ ;
	assign \g48087/_0_  = _w2663_ ;
	assign \g48110/_0_  = _w2667_ ;
	assign \g48117/_0_  = _w2675_ ;
	assign \g48118/_0_  = _w2680_ ;
	assign \g48119/_0_  = _w2687_ ;
	assign \g48120/_0_  = _w2694_ ;
	assign \g48121/_0_  = _w2701_ ;
	assign \g48122/_0_  = _w2708_ ;
	assign \g48124/_0_  = _w2715_ ;
	assign \g48125/_0_  = _w2733_ ;
	assign \g48126/_0_  = _w2751_ ;
	assign \g48127/_0_  = _w2768_ ;
	assign \g48128/_0_  = _w2773_ ;
	assign \g48129/_0_  = _w2789_ ;
	assign \g48130/_0_  = _w2809_ ;
	assign \g48131/_0_  = _w2829_ ;
	assign \g48132/_0_  = _w2849_ ;
	assign \g48133/_0_  = _w2868_ ;
	assign \g48134/_0_  = _w2875_ ;
	assign \g48168/_0_  = _w2885_ ;
	assign \g48169/_0_  = _w2895_ ;
	assign \g48170/_0_  = _w2904_ ;
	assign \g48171/_0_  = _w2913_ ;
	assign \g48172/_0_  = _w2922_ ;
	assign \g48173/_0_  = _w2931_ ;
	assign \g48174/_0_  = _w2940_ ;
	assign \g48175/_0_  = _w2949_ ;
	assign \g48177/_0_  = _w2958_ ;
	assign \g48178/_0_  = _w2967_ ;
	assign \g48179/_0_  = _w2976_ ;
	assign \g48180/_0_  = _w2985_ ;
	assign \g48181/_0_  = _w2994_ ;
	assign \g48182/_0_  = _w3003_ ;
	assign \g48183/_0_  = _w3012_ ;
	assign \g48184/_0_  = _w3021_ ;
	assign \g48185/_0_  = _w3030_ ;
	assign \g48186/_0_  = _w3039_ ;
	assign \g48187/_0_  = _w3048_ ;
	assign \g48188/_0_  = _w3057_ ;
	assign \g48189/_0_  = _w3066_ ;
	assign \g48192/_0_  = _w3075_ ;
	assign \g48193/_0_  = _w3084_ ;
	assign \g48194/_0_  = _w3093_ ;
	assign \g48195/_0_  = _w3102_ ;
	assign \g48196/_0_  = _w3111_ ;
	assign \g48197/_0_  = _w3120_ ;
	assign \g48198/_0_  = _w3129_ ;
	assign \g48199/_0_  = _w3138_ ;
	assign \g48200/_0_  = _w3147_ ;
	assign \g48201/_0_  = _w3156_ ;
	assign \g48202/_0_  = _w3165_ ;
	assign \g48203/_0_  = _w3168_ ;
	assign \g48213/_0_  = _w3185_ ;
	assign \g48214/_0_  = _w3202_ ;
	assign \g48215/_0_  = _w3225_ ;
	assign \g48216/_0_  = _w3240_ ;
	assign \g48217/_0_  = _w3256_ ;
	assign \g48218/_0_  = _w3276_ ;
	assign \g48219/_0_  = _w3292_ ;
	assign \g48220/_0_  = _w3307_ ;
	assign \g48221/_0_  = _w3322_ ;
	assign \g48222/_0_  = _w3339_ ;
	assign \g48223/_0_  = _w3356_ ;
	assign \g48224/_0_  = _w3371_ ;
	assign \g48225/_0_  = _w3389_ ;
	assign \g48226/_0_  = _w3406_ ;
	assign \g48227/_0_  = _w3422_ ;
	assign \g48228/_0_  = _w3439_ ;
	assign \g48229/_0_  = _w3455_ ;
	assign \g48230/_0_  = _w3472_ ;
	assign \g48231/_0_  = _w3489_ ;
	assign \g48232/_0_  = _w3507_ ;
	assign \g48234/_0_  = _w3512_ ;
	assign \g48236/_0_  = _w3529_ ;
	assign \g48237/_0_  = _w3546_ ;
	assign \g48238/_0_  = _w3564_ ;
	assign \g48239/_0_  = _w3584_ ;
	assign \g48240/_0_  = _w3602_ ;
	assign \g48241/_0_  = _w3618_ ;
	assign \g48243/_0_  = _w3636_ ;
	assign \g48244/_0_  = _w3653_ ;
	assign \g48245/_0_  = _w3668_ ;
	assign \g48246/_0_  = _w3687_ ;
	assign \g48263/_0_  = _w3694_ ;
	assign \g48270/_0_  = _w3702_ ;
	assign \g48273/_0_  = _w3710_ ;
	assign \g48276/_0_  = _w3716_ ;
	assign \g48277/_0_  = _w3721_ ;
	assign \g48370/_0_  = _w3724_ ;
	assign \g48377/_0_  = _w3727_ ;
	assign \g48391/_0_  = _w3738_ ;
	assign \g48423/_0_  = _w3744_ ;
	assign \g48428/_0_  = _w3754_ ;
	assign \g48429/_0_  = _w3761_ ;
	assign \g48431/_0_  = _w3767_ ;
	assign \g48433/_0_  = _w3774_ ;
	assign \g48434/_0_  = _w3794_ ;
	assign \g48435/_0_  = _w3814_ ;
	assign \g48436/_0_  = _w3837_ ;
	assign \g48437/_0_  = _w3856_ ;
	assign \g48438/_0_  = _w3858_ ;
	assign \g48439/_0_  = _w3877_ ;
	assign \g48440/_0_  = _w3897_ ;
	assign \g48441/_0_  = _w3918_ ;
	assign \g48442/_0_  = _w3926_ ;
	assign \g48443/_0_  = _w3936_ ;
	assign \g48610/_0_  = _w3941_ ;
	assign \g48634/_0_  = _w3947_ ;
	assign \g48635/_0_  = _w3951_ ;
	assign \g48636/_0_  = _w3955_ ;
	assign \g48637/_0_  = _w3963_ ;
	assign \g48638/_0_  = _w3969_ ;
	assign \g48639/_0_  = _w3976_ ;
	assign \g48640/_0_  = _w3982_ ;
	assign \g48642/_0_  = _w3987_ ;
	assign \g48643/_0_  = _w3992_ ;
	assign \g48644/_0_  = _w3998_ ;
	assign \g48645/_0_  = _w4004_ ;
	assign \g48646/_0_  = _w4009_ ;
	assign \g48647/_0_  = _w4016_ ;
	assign \g48648/_0_  = _w4021_ ;
	assign \g48649/_0_  = _w4026_ ;
	assign \g48650/_0_  = _w4031_ ;
	assign \g48651/_0_  = _w4036_ ;
	assign \g48652/_0_  = _w4041_ ;
	assign \g48653/_0_  = _w4046_ ;
	assign \g48654/_0_  = _w4051_ ;
	assign \g48655/_0_  = _w4058_ ;
	assign \g48656/_0_  = _w4063_ ;
	assign \g48657/_0_  = _w4068_ ;
	assign \g48658/_0_  = _w4073_ ;
	assign \g48659/_0_  = _w4078_ ;
	assign \g48660/_0_  = _w4084_ ;
	assign \g48662/_0_  = _w4090_ ;
	assign \g48663/_0_  = _w4096_ ;
	assign \g48664/_0_  = _w4102_ ;
	assign \g48665/_0_  = _w4108_ ;
	assign \g48666/_0_  = _w4114_ ;
	assign \g48667/_0_  = _w4120_ ;
	assign \g48668/_0_  = _w4126_ ;
	assign \g48669/_0_  = _w4128_ ;
	assign \g48750/_0_  = _w4138_ ;
	assign \g48753/_0_  = _w4148_ ;
	assign \g48756/_0_  = _w4158_ ;
	assign \g48759/_0_  = _w4168_ ;
	assign \g48763/_0_  = _w4178_ ;
	assign \g48766/_0_  = _w4188_ ;
	assign \g48769/_0_  = _w4198_ ;
	assign \g48772/_0_  = _w4208_ ;
	assign \g48775/_0_  = _w4218_ ;
	assign \g48778/_0_  = _w4228_ ;
	assign \g48781/_0_  = _w4238_ ;
	assign \g48785/_0_  = _w4248_ ;
	assign \g48789/_0_  = _w4258_ ;
	assign \g48792/_0_  = _w4268_ ;
	assign \g48796/_0_  = _w4278_ ;
	assign \g48799/_0_  = _w4288_ ;
	assign \g48937/_0_  = _w4292_ ;
	assign \g48958/_0_  = _w4295_ ;
	assign \g48959/_0_  = _w4299_ ;
	assign \g48964/_0_  = _w4303_ ;
	assign \g48965/_0_  = _w4307_ ;
	assign \g48966/_0_  = _w4311_ ;
	assign \g48967/_0_  = _w4316_ ;
	assign \g48968/_0_  = _w4320_ ;
	assign \g48969/_0_  = _w4325_ ;
	assign \g48970/_0_  = _w4332_ ;
	assign \g48971/_0_  = _w4337_ ;
	assign \g48972/_0_  = _w4341_ ;
	assign \g48973/_0_  = _w4346_ ;
	assign \g48974/_0_  = _w4350_ ;
	assign \g48975/_0_  = _w4355_ ;
	assign \g48976/_0_  = _w4360_ ;
	assign \g48977/_0_  = _w4365_ ;
	assign \g48978/_0_  = _w4370_ ;
	assign \g48979/_0_  = _w4374_ ;
	assign \g49/_0_  = _w4384_ ;
	assign \g49069/_0_  = _w4394_ ;
	assign \g49070/_0_  = _w4404_ ;
	assign \g49071/_0_  = _w4414_ ;
	assign \g49073/_0_  = _w4424_ ;
	assign \g49074/_0_  = _w4434_ ;
	assign \g49076/_0_  = _w4444_ ;
	assign \g49078/_0_  = _w4454_ ;
	assign \g49081/_0_  = _w4464_ ;
	assign \g49083/_0_  = _w4474_ ;
	assign \g49085/_0_  = _w4484_ ;
	assign \g49087/_0_  = _w4494_ ;
	assign \g49088/_0_  = _w4504_ ;
	assign \g49090/_0_  = _w4514_ ;
	assign \g49092/_0_  = _w4524_ ;
	assign \g49095/_0_  = _w4534_ ;
	assign \g49098/_0_  = _w4544_ ;
	assign \g49125/_0_  = _w4568_ ;
	assign \g49162/_0_  = _w4571_ ;
	assign \g49202/_0_  = _w4577_ ;
	assign \g49203/_0_  = _w4583_ ;
	assign \g49206/_0_  = _w4587_ ;
	assign \g49340/_0_  = _w4597_ ;
	assign \g49457/_0_  = _w4606_ ;
	assign \g49512/_0_  = _w4609_ ;
	assign \g49513/_0_  = _w4612_ ;
	assign \g49514/_0_  = _w4615_ ;
	assign \g49515/_0_  = _w4618_ ;
	assign \g49516/_0_  = _w4621_ ;
	assign \g49517/_0_  = _w4624_ ;
	assign \g49518/_0_  = _w4627_ ;
	assign \g49519/_0_  = _w4630_ ;
	assign \g49520/_0_  = _w4633_ ;
	assign \g49521/_0_  = _w4636_ ;
	assign \g49522/_0_  = _w4639_ ;
	assign \g49523/_0_  = _w4642_ ;
	assign \g49524/_0_  = _w4645_ ;
	assign \g49525/_0_  = _w4648_ ;
	assign \g49526/_0_  = _w4651_ ;
	assign \g49527/_0_  = _w4654_ ;
	assign \g49534/_0_  = _w4664_ ;
	assign \g49551/_0_  = _w4670_ ;
	assign \g49573/_0_  = _w4675_ ;
	assign \g49574/_0_  = _w4686_ ;
	assign \g49578/_0_  = _w4696_ ;
	assign \g49582/_0_  = _w4707_ ;
	assign \g49584/_0_  = _w4717_ ;
	assign \g49592/_0_  = _w4727_ ;
	assign \g49600/_0_  = _w4737_ ;
	assign \g49604/_0_  = _w4747_ ;
	assign \g49608/_0_  = _w4757_ ;
	assign \g49612/_0_  = _w4767_ ;
	assign \g49616/_0_  = _w4777_ ;
	assign \g49619/_0_  = _w4787_ ;
	assign \g49620/_0_  = _w4797_ ;
	assign \g49623/_0_  = _w4807_ ;
	assign \g49627/_0_  = _w4817_ ;
	assign \g49630/_0_  = _w4827_ ;
	assign \g49634/_0_  = _w4837_ ;
	assign \g49635/_0_  = _w4847_ ;
	assign \g49639/_0_  = _w4857_ ;
	assign \g49645/_0_  = _w4867_ ;
	assign \g49744/_0_  = _w4872_ ;
	assign \g49766/_0_  = _w4877_ ;
	assign \g50098/_0_  = _w4884_ ;
	assign \g50124/_0_  = _w4891_ ;
	assign \g50195/_0_  = _w4901_ ;
	assign \g50198/_0_  = _w4911_ ;
	assign \g50201/_0_  = _w4921_ ;
	assign \g50203/_0_  = _w4931_ ;
	assign \g50205/_0_  = _w4941_ ;
	assign \g50207/_0_  = _w4951_ ;
	assign \g50209/_0_  = _w4961_ ;
	assign \g50213/_0_  = _w4971_ ;
	assign \g50222/_0_  = _w4981_ ;
	assign \g50228/_0_  = _w4991_ ;
	assign \g50231/_0_  = _w5001_ ;
	assign \g50237/_0_  = _w5011_ ;
	assign \g50240/_0_  = _w5021_ ;
	assign \g50335/_0_  = _w5029_ ;
	assign \g50477/_0_  = _w5035_ ;
	assign \g50478/_0_  = _w5039_ ;
	assign \g50671/_0_  = _w5044_ ;
	assign \g50757/_0_  = _w5051_ ;
	assign \g50938/_0_  = _w5056_ ;
	assign \g50998/_0_  = _w5061_ ;
	assign \g51008/_0_  = _w5066_ ;
	assign \g51579/_0_  = _w5070_ ;
	assign \g51637/_0_  = _w5075_ ;
	assign \g51662/_0_  = _w5080_ ;
	assign \g52424/_0_  = _w5087_ ;
	assign \g53184/_0_  = _w5091_ ;
	assign \g53206/_0_  = _w5097_ ;
	assign \g53270/_0_  = _w5100_ ;
	assign \g53730/_0_  = _w5106_ ;
	assign \g53754/_0_  = _w5112_ ;
	assign \g54176/_0_  = _w5117_ ;
	assign \g54214/_0_  = _w5120_ ;
	assign \g54229/_0_  = _w5125_ ;
	assign \g54392/_0_  = _w5129_ ;
	assign \g54400/_0_  = _w5132_ ;
	assign \g54415/_0_  = _w5135_ ;
	assign \g54421/_0_  = _w5139_ ;
	assign \g54604/_0_  = _w5143_ ;
	assign \g54607/_0_  = _w5147_ ;
	assign \g54638/_0_  = _w5151_ ;
	assign \g54694/_0_  = _w5159_ ;
	assign \g54759/_0_  = _w5162_ ;
	assign \g55607/_0_  = _w5166_ ;
	assign \g55863/_1_  = _w5126_ ;
	assign \g56073/_0_  = _w5169_ ;
	assign \g56292/_0_  = _w5170_ ;
	assign \g56320/_0_  = _w5171_ ;
	assign \g56527/_0_  = _w5172_ ;
	assign \g56531/_0_  = _w5173_ ;
	assign \g56533/_0_  = _w5174_ ;
	assign \g56562/_0_  = _w5175_ ;
	assign \g56615/_0_  = _w5176_ ;
	assign \g56720/_0_  = _w5179_ ;
	assign \g57044/_0_  = _w5181_ ;
	assign \g60635/_1_  = _w4545_ ;
	assign \g62873/_0_  = _w5203_ ;
	assign \g62886/_0_  = _w5221_ ;
	assign \g63001/_0_  = _w5239_ ;
	assign \g63101/_0_  = _w5250_ ;
	assign \g63129/_0_  = _w5256_ ;
	assign \g63198/_0_  = _w5267_ ;
	assign \g63449/_0_  = _w5276_ ;
	assign \g63471/_0_  = _w5284_ ;
	assign \g63493/_0_  = _w5290_ ;
	assign \g63626/_0_  = _w5299_ ;
	assign \g63688/_0_  = _w5315_ ;
	assign \g63800/_0_  = _w5333_ ;
	assign \g63934/_0_  = _w5344_ ;
	assign \g63954/_0_  = _w5355_ ;
	assign \g64060/_0_  = _w5364_ ;
	assign \g64375/_0_  = _w5374_ ;
	assign \g65/_0_  = _w5384_ ;
	assign \g67/_0_  = _w5394_ ;
endmodule;