module top (\priority[0] , \priority[1] , \priority[2] , \priority[3] , \priority[4] , \priority[5] , \priority[6] , \priority[7] , \priority[8] , \priority[9] , \priority[10] , \priority[11] , \priority[12] , \priority[13] , \priority[14] , \priority[15] , \priority[16] , \priority[17] , \priority[18] , \priority[19] , \priority[20] , \priority[21] , \priority[22] , \priority[23] , \priority[24] , \priority[25] , \priority[26] , \priority[27] , \priority[28] , \priority[29] , \priority[30] , \priority[31] , \priority[32] , \priority[33] , \priority[34] , \priority[35] , \priority[36] , \priority[37] , \priority[38] , \priority[39] , \priority[40] , \priority[41] , \priority[42] , \priority[43] , \priority[44] , \priority[45] , \priority[46] , \priority[47] , \priority[48] , \priority[49] , \priority[50] , \priority[51] , \priority[52] , \priority[53] , \priority[54] , \priority[55] , \priority[56] , \priority[57] , \priority[58] , \priority[59] , \priority[60] , \priority[61] , \priority[62] , \priority[63] , \priority[64] , \priority[65] , \priority[66] , \priority[67] , \priority[68] , \priority[69] , \priority[70] , \priority[71] , \priority[72] , \priority[73] , \priority[74] , \priority[75] , \priority[76] , \priority[77] , \priority[78] , \priority[79] , \priority[80] , \priority[81] , \priority[82] , \priority[83] , \priority[84] , \priority[85] , \priority[86] , \priority[87] , \priority[88] , \priority[89] , \priority[90] , \priority[91] , \priority[92] , \priority[93] , \priority[94] , \priority[95] , \priority[96] , \priority[97] , \priority[98] , \priority[99] , \priority[100] , \priority[101] , \priority[102] , \priority[103] , \priority[104] , \priority[105] , \priority[106] , \priority[107] , \priority[108] , \priority[109] , \priority[110] , \priority[111] , \priority[112] , \priority[113] , \priority[114] , \priority[115] , \priority[116] , \priority[117] , \priority[118] , \priority[119] , \priority[120] , \priority[121] , \priority[122] , \priority[123] , \priority[124] , \priority[125] , \priority[126] , \priority[127] , \req[0] , \req[1] , \req[2] , \req[3] , \req[4] , \req[5] , \req[6] , \req[7] , \req[8] , \req[9] , \req[10] , \req[11] , \req[12] , \req[13] , \req[14] , \req[15] , \req[16] , \req[17] , \req[18] , \req[19] , \req[20] , \req[21] , \req[22] , \req[23] , \req[24] , \req[25] , \req[26] , \req[27] , \req[28] , \req[29] , \req[30] , \req[31] , \req[32] , \req[33] , \req[34] , \req[35] , \req[36] , \req[37] , \req[38] , \req[39] , \req[40] , \req[41] , \req[42] , \req[43] , \req[44] , \req[45] , \req[46] , \req[47] , \req[48] , \req[49] , \req[50] , \req[51] , \req[52] , \req[53] , \req[54] , \req[55] , \req[56] , \req[57] , \req[58] , \req[59] , \req[60] , \req[61] , \req[62] , \req[63] , \req[64] , \req[65] , \req[66] , \req[67] , \req[68] , \req[69] , \req[70] , \req[71] , \req[72] , \req[73] , \req[74] , \req[75] , \req[76] , \req[77] , \req[78] , \req[79] , \req[80] , \req[81] , \req[82] , \req[83] , \req[84] , \req[85] , \req[86] , \req[87] , \req[88] , \req[89] , \req[90] , \req[91] , \req[92] , \req[93] , \req[94] , \req[95] , \req[96] , \req[97] , \req[98] , \req[99] , \req[100] , \req[101] , \req[102] , \req[103] , \req[104] , \req[105] , \req[106] , \req[107] , \req[108] , \req[109] , \req[110] , \req[111] , \req[112] , \req[113] , \req[114] , \req[115] , \req[116] , \req[117] , \req[118] , \req[119] , \req[120] , \req[121] , \req[122] , \req[123] , \req[124] , \req[125] , \req[126] , \req[127] , \grant[0] , \grant[1] , \grant[2] , \grant[3] , \grant[4] , \grant[5] , \grant[6] , \grant[7] , \grant[8] , \grant[9] , \grant[10] , \grant[11] , \grant[12] , \grant[13] , \grant[14] , \grant[15] , \grant[16] , \grant[17] , \grant[18] , \grant[19] , \grant[20] , \grant[21] , \grant[22] , \grant[23] , \grant[24] , \grant[25] , \grant[26] , \grant[27] , \grant[28] , \grant[29] , \grant[30] , \grant[31] , \grant[32] , \grant[33] , \grant[34] , \grant[35] , \grant[36] , \grant[37] , \grant[38] , \grant[39] , \grant[40] , \grant[41] , \grant[42] , \grant[43] , \grant[44] , \grant[45] , \grant[46] , \grant[47] , \grant[48] , \grant[49] , \grant[50] , \grant[51] , \grant[52] , \grant[53] , \grant[54] , \grant[55] , \grant[56] , \grant[57] , \grant[58] , \grant[59] , \grant[60] , \grant[61] , \grant[62] , \grant[63] , \grant[64] , \grant[65] , \grant[66] , \grant[67] , \grant[68] , \grant[69] , \grant[70] , \grant[71] , \grant[72] , \grant[73] , \grant[74] , \grant[75] , \grant[76] , \grant[77] , \grant[78] , \grant[79] , \grant[80] , \grant[81] , \grant[82] , \grant[83] , \grant[84] , \grant[85] , \grant[86] , \grant[87] , \grant[88] , \grant[89] , \grant[90] , \grant[91] , \grant[92] , \grant[93] , \grant[94] , \grant[95] , \grant[96] , \grant[97] , \grant[98] , \grant[99] , \grant[100] , \grant[101] , \grant[102] , \grant[103] , \grant[104] , \grant[105] , \grant[106] , \grant[107] , \grant[108] , \grant[109] , \grant[110] , \grant[111] , \grant[112] , \grant[113] , \grant[114] , \grant[115] , \grant[116] , \grant[117] , \grant[118] , \grant[119] , \grant[120] , \grant[121] , \grant[122] , \grant[123] , \grant[124] , \grant[125] , \grant[126] , \grant[127] , anyGrant);
	input \priority[0]  ;
	input \priority[1]  ;
	input \priority[2]  ;
	input \priority[3]  ;
	input \priority[4]  ;
	input \priority[5]  ;
	input \priority[6]  ;
	input \priority[7]  ;
	input \priority[8]  ;
	input \priority[9]  ;
	input \priority[10]  ;
	input \priority[11]  ;
	input \priority[12]  ;
	input \priority[13]  ;
	input \priority[14]  ;
	input \priority[15]  ;
	input \priority[16]  ;
	input \priority[17]  ;
	input \priority[18]  ;
	input \priority[19]  ;
	input \priority[20]  ;
	input \priority[21]  ;
	input \priority[22]  ;
	input \priority[23]  ;
	input \priority[24]  ;
	input \priority[25]  ;
	input \priority[26]  ;
	input \priority[27]  ;
	input \priority[28]  ;
	input \priority[29]  ;
	input \priority[30]  ;
	input \priority[31]  ;
	input \priority[32]  ;
	input \priority[33]  ;
	input \priority[34]  ;
	input \priority[35]  ;
	input \priority[36]  ;
	input \priority[37]  ;
	input \priority[38]  ;
	input \priority[39]  ;
	input \priority[40]  ;
	input \priority[41]  ;
	input \priority[42]  ;
	input \priority[43]  ;
	input \priority[44]  ;
	input \priority[45]  ;
	input \priority[46]  ;
	input \priority[47]  ;
	input \priority[48]  ;
	input \priority[49]  ;
	input \priority[50]  ;
	input \priority[51]  ;
	input \priority[52]  ;
	input \priority[53]  ;
	input \priority[54]  ;
	input \priority[55]  ;
	input \priority[56]  ;
	input \priority[57]  ;
	input \priority[58]  ;
	input \priority[59]  ;
	input \priority[60]  ;
	input \priority[61]  ;
	input \priority[62]  ;
	input \priority[63]  ;
	input \priority[64]  ;
	input \priority[65]  ;
	input \priority[66]  ;
	input \priority[67]  ;
	input \priority[68]  ;
	input \priority[69]  ;
	input \priority[70]  ;
	input \priority[71]  ;
	input \priority[72]  ;
	input \priority[73]  ;
	input \priority[74]  ;
	input \priority[75]  ;
	input \priority[76]  ;
	input \priority[77]  ;
	input \priority[78]  ;
	input \priority[79]  ;
	input \priority[80]  ;
	input \priority[81]  ;
	input \priority[82]  ;
	input \priority[83]  ;
	input \priority[84]  ;
	input \priority[85]  ;
	input \priority[86]  ;
	input \priority[87]  ;
	input \priority[88]  ;
	input \priority[89]  ;
	input \priority[90]  ;
	input \priority[91]  ;
	input \priority[92]  ;
	input \priority[93]  ;
	input \priority[94]  ;
	input \priority[95]  ;
	input \priority[96]  ;
	input \priority[97]  ;
	input \priority[98]  ;
	input \priority[99]  ;
	input \priority[100]  ;
	input \priority[101]  ;
	input \priority[102]  ;
	input \priority[103]  ;
	input \priority[104]  ;
	input \priority[105]  ;
	input \priority[106]  ;
	input \priority[107]  ;
	input \priority[108]  ;
	input \priority[109]  ;
	input \priority[110]  ;
	input \priority[111]  ;
	input \priority[112]  ;
	input \priority[113]  ;
	input \priority[114]  ;
	input \priority[115]  ;
	input \priority[116]  ;
	input \priority[117]  ;
	input \priority[118]  ;
	input \priority[119]  ;
	input \priority[120]  ;
	input \priority[121]  ;
	input \priority[122]  ;
	input \priority[123]  ;
	input \priority[124]  ;
	input \priority[125]  ;
	input \priority[126]  ;
	input \priority[127]  ;
	input \req[0]  ;
	input \req[1]  ;
	input \req[2]  ;
	input \req[3]  ;
	input \req[4]  ;
	input \req[5]  ;
	input \req[6]  ;
	input \req[7]  ;
	input \req[8]  ;
	input \req[9]  ;
	input \req[10]  ;
	input \req[11]  ;
	input \req[12]  ;
	input \req[13]  ;
	input \req[14]  ;
	input \req[15]  ;
	input \req[16]  ;
	input \req[17]  ;
	input \req[18]  ;
	input \req[19]  ;
	input \req[20]  ;
	input \req[21]  ;
	input \req[22]  ;
	input \req[23]  ;
	input \req[24]  ;
	input \req[25]  ;
	input \req[26]  ;
	input \req[27]  ;
	input \req[28]  ;
	input \req[29]  ;
	input \req[30]  ;
	input \req[31]  ;
	input \req[32]  ;
	input \req[33]  ;
	input \req[34]  ;
	input \req[35]  ;
	input \req[36]  ;
	input \req[37]  ;
	input \req[38]  ;
	input \req[39]  ;
	input \req[40]  ;
	input \req[41]  ;
	input \req[42]  ;
	input \req[43]  ;
	input \req[44]  ;
	input \req[45]  ;
	input \req[46]  ;
	input \req[47]  ;
	input \req[48]  ;
	input \req[49]  ;
	input \req[50]  ;
	input \req[51]  ;
	input \req[52]  ;
	input \req[53]  ;
	input \req[54]  ;
	input \req[55]  ;
	input \req[56]  ;
	input \req[57]  ;
	input \req[58]  ;
	input \req[59]  ;
	input \req[60]  ;
	input \req[61]  ;
	input \req[62]  ;
	input \req[63]  ;
	input \req[64]  ;
	input \req[65]  ;
	input \req[66]  ;
	input \req[67]  ;
	input \req[68]  ;
	input \req[69]  ;
	input \req[70]  ;
	input \req[71]  ;
	input \req[72]  ;
	input \req[73]  ;
	input \req[74]  ;
	input \req[75]  ;
	input \req[76]  ;
	input \req[77]  ;
	input \req[78]  ;
	input \req[79]  ;
	input \req[80]  ;
	input \req[81]  ;
	input \req[82]  ;
	input \req[83]  ;
	input \req[84]  ;
	input \req[85]  ;
	input \req[86]  ;
	input \req[87]  ;
	input \req[88]  ;
	input \req[89]  ;
	input \req[90]  ;
	input \req[91]  ;
	input \req[92]  ;
	input \req[93]  ;
	input \req[94]  ;
	input \req[95]  ;
	input \req[96]  ;
	input \req[97]  ;
	input \req[98]  ;
	input \req[99]  ;
	input \req[100]  ;
	input \req[101]  ;
	input \req[102]  ;
	input \req[103]  ;
	input \req[104]  ;
	input \req[105]  ;
	input \req[106]  ;
	input \req[107]  ;
	input \req[108]  ;
	input \req[109]  ;
	input \req[110]  ;
	input \req[111]  ;
	input \req[112]  ;
	input \req[113]  ;
	input \req[114]  ;
	input \req[115]  ;
	input \req[116]  ;
	input \req[117]  ;
	input \req[118]  ;
	input \req[119]  ;
	input \req[120]  ;
	input \req[121]  ;
	input \req[122]  ;
	input \req[123]  ;
	input \req[124]  ;
	input \req[125]  ;
	input \req[126]  ;
	input \req[127]  ;
	output \grant[0]  ;
	output \grant[1]  ;
	output \grant[2]  ;
	output \grant[3]  ;
	output \grant[4]  ;
	output \grant[5]  ;
	output \grant[6]  ;
	output \grant[7]  ;
	output \grant[8]  ;
	output \grant[9]  ;
	output \grant[10]  ;
	output \grant[11]  ;
	output \grant[12]  ;
	output \grant[13]  ;
	output \grant[14]  ;
	output \grant[15]  ;
	output \grant[16]  ;
	output \grant[17]  ;
	output \grant[18]  ;
	output \grant[19]  ;
	output \grant[20]  ;
	output \grant[21]  ;
	output \grant[22]  ;
	output \grant[23]  ;
	output \grant[24]  ;
	output \grant[25]  ;
	output \grant[26]  ;
	output \grant[27]  ;
	output \grant[28]  ;
	output \grant[29]  ;
	output \grant[30]  ;
	output \grant[31]  ;
	output \grant[32]  ;
	output \grant[33]  ;
	output \grant[34]  ;
	output \grant[35]  ;
	output \grant[36]  ;
	output \grant[37]  ;
	output \grant[38]  ;
	output \grant[39]  ;
	output \grant[40]  ;
	output \grant[41]  ;
	output \grant[42]  ;
	output \grant[43]  ;
	output \grant[44]  ;
	output \grant[45]  ;
	output \grant[46]  ;
	output \grant[47]  ;
	output \grant[48]  ;
	output \grant[49]  ;
	output \grant[50]  ;
	output \grant[51]  ;
	output \grant[52]  ;
	output \grant[53]  ;
	output \grant[54]  ;
	output \grant[55]  ;
	output \grant[56]  ;
	output \grant[57]  ;
	output \grant[58]  ;
	output \grant[59]  ;
	output \grant[60]  ;
	output \grant[61]  ;
	output \grant[62]  ;
	output \grant[63]  ;
	output \grant[64]  ;
	output \grant[65]  ;
	output \grant[66]  ;
	output \grant[67]  ;
	output \grant[68]  ;
	output \grant[69]  ;
	output \grant[70]  ;
	output \grant[71]  ;
	output \grant[72]  ;
	output \grant[73]  ;
	output \grant[74]  ;
	output \grant[75]  ;
	output \grant[76]  ;
	output \grant[77]  ;
	output \grant[78]  ;
	output \grant[79]  ;
	output \grant[80]  ;
	output \grant[81]  ;
	output \grant[82]  ;
	output \grant[83]  ;
	output \grant[84]  ;
	output \grant[85]  ;
	output \grant[86]  ;
	output \grant[87]  ;
	output \grant[88]  ;
	output \grant[89]  ;
	output \grant[90]  ;
	output \grant[91]  ;
	output \grant[92]  ;
	output \grant[93]  ;
	output \grant[94]  ;
	output \grant[95]  ;
	output \grant[96]  ;
	output \grant[97]  ;
	output \grant[98]  ;
	output \grant[99]  ;
	output \grant[100]  ;
	output \grant[101]  ;
	output \grant[102]  ;
	output \grant[103]  ;
	output \grant[104]  ;
	output \grant[105]  ;
	output \grant[106]  ;
	output \grant[107]  ;
	output \grant[108]  ;
	output \grant[109]  ;
	output \grant[110]  ;
	output \grant[111]  ;
	output \grant[112]  ;
	output \grant[113]  ;
	output \grant[114]  ;
	output \grant[115]  ;
	output \grant[116]  ;
	output \grant[117]  ;
	output \grant[118]  ;
	output \grant[119]  ;
	output \grant[120]  ;
	output \grant[121]  ;
	output \grant[122]  ;
	output \grant[123]  ;
	output \grant[124]  ;
	output \grant[125]  ;
	output \grant[126]  ;
	output \grant[127]  ;
	output anyGrant ;
	wire _w2860_ ;
	wire _w2859_ ;
	wire _w2858_ ;
	wire _w2857_ ;
	wire _w2856_ ;
	wire _w2855_ ;
	wire _w2854_ ;
	wire _w2853_ ;
	wire _w2852_ ;
	wire _w2851_ ;
	wire _w2850_ ;
	wire _w2849_ ;
	wire _w2848_ ;
	wire _w2847_ ;
	wire _w2846_ ;
	wire _w2845_ ;
	wire _w2844_ ;
	wire _w2843_ ;
	wire _w2842_ ;
	wire _w2841_ ;
	wire _w2840_ ;
	wire _w2839_ ;
	wire _w2838_ ;
	wire _w2837_ ;
	wire _w2836_ ;
	wire _w2835_ ;
	wire _w2834_ ;
	wire _w2833_ ;
	wire _w2832_ ;
	wire _w2831_ ;
	wire _w2830_ ;
	wire _w2829_ ;
	wire _w2828_ ;
	wire _w2827_ ;
	wire _w2826_ ;
	wire _w2825_ ;
	wire _w2824_ ;
	wire _w2823_ ;
	wire _w2822_ ;
	wire _w2821_ ;
	wire _w2820_ ;
	wire _w2819_ ;
	wire _w2818_ ;
	wire _w2817_ ;
	wire _w2816_ ;
	wire _w2815_ ;
	wire _w2814_ ;
	wire _w2813_ ;
	wire _w2812_ ;
	wire _w2811_ ;
	wire _w2810_ ;
	wire _w2809_ ;
	wire _w2808_ ;
	wire _w2807_ ;
	wire _w2806_ ;
	wire _w2805_ ;
	wire _w2804_ ;
	wire _w2803_ ;
	wire _w2802_ ;
	wire _w2801_ ;
	wire _w2800_ ;
	wire _w2799_ ;
	wire _w2798_ ;
	wire _w2797_ ;
	wire _w2796_ ;
	wire _w2795_ ;
	wire _w2794_ ;
	wire _w2793_ ;
	wire _w2792_ ;
	wire _w2791_ ;
	wire _w2790_ ;
	wire _w2789_ ;
	wire _w2788_ ;
	wire _w2787_ ;
	wire _w2786_ ;
	wire _w2785_ ;
	wire _w2784_ ;
	wire _w2783_ ;
	wire _w2782_ ;
	wire _w2781_ ;
	wire _w2780_ ;
	wire _w2779_ ;
	wire _w2778_ ;
	wire _w2777_ ;
	wire _w2776_ ;
	wire _w2775_ ;
	wire _w2774_ ;
	wire _w2773_ ;
	wire _w2772_ ;
	wire _w2771_ ;
	wire _w2770_ ;
	wire _w2769_ ;
	wire _w2768_ ;
	wire _w2767_ ;
	wire _w2766_ ;
	wire _w2765_ ;
	wire _w2764_ ;
	wire _w2763_ ;
	wire _w2762_ ;
	wire _w2761_ ;
	wire _w2760_ ;
	wire _w2759_ ;
	wire _w2758_ ;
	wire _w2757_ ;
	wire _w2756_ ;
	wire _w2755_ ;
	wire _w2754_ ;
	wire _w2753_ ;
	wire _w2752_ ;
	wire _w2751_ ;
	wire _w2750_ ;
	wire _w2749_ ;
	wire _w2748_ ;
	wire _w2747_ ;
	wire _w2746_ ;
	wire _w2745_ ;
	wire _w2744_ ;
	wire _w2743_ ;
	wire _w2742_ ;
	wire _w2741_ ;
	wire _w2740_ ;
	wire _w2739_ ;
	wire _w2738_ ;
	wire _w2737_ ;
	wire _w2736_ ;
	wire _w2735_ ;
	wire _w2734_ ;
	wire _w2733_ ;
	wire _w2732_ ;
	wire _w2731_ ;
	wire _w2730_ ;
	wire _w2729_ ;
	wire _w2728_ ;
	wire _w2727_ ;
	wire _w2726_ ;
	wire _w2725_ ;
	wire _w2724_ ;
	wire _w2723_ ;
	wire _w2722_ ;
	wire _w2721_ ;
	wire _w2720_ ;
	wire _w2719_ ;
	wire _w2718_ ;
	wire _w2717_ ;
	wire _w2716_ ;
	wire _w2715_ ;
	wire _w2714_ ;
	wire _w2713_ ;
	wire _w2712_ ;
	wire _w2711_ ;
	wire _w2710_ ;
	wire _w2709_ ;
	wire _w2708_ ;
	wire _w2707_ ;
	wire _w2706_ ;
	wire _w2705_ ;
	wire _w2704_ ;
	wire _w2703_ ;
	wire _w2702_ ;
	wire _w2701_ ;
	wire _w2700_ ;
	wire _w2699_ ;
	wire _w2698_ ;
	wire _w2697_ ;
	wire _w2696_ ;
	wire _w2695_ ;
	wire _w2694_ ;
	wire _w2693_ ;
	wire _w2692_ ;
	wire _w2691_ ;
	wire _w2690_ ;
	wire _w2689_ ;
	wire _w2688_ ;
	wire _w2687_ ;
	wire _w2686_ ;
	wire _w2685_ ;
	wire _w2684_ ;
	wire _w2683_ ;
	wire _w2682_ ;
	wire _w2681_ ;
	wire _w2680_ ;
	wire _w2679_ ;
	wire _w2678_ ;
	wire _w2677_ ;
	wire _w2676_ ;
	wire _w2675_ ;
	wire _w2674_ ;
	wire _w2673_ ;
	wire _w2672_ ;
	wire _w2671_ ;
	wire _w2670_ ;
	wire _w2669_ ;
	wire _w2668_ ;
	wire _w2667_ ;
	wire _w2666_ ;
	wire _w2665_ ;
	wire _w2664_ ;
	wire _w2663_ ;
	wire _w2662_ ;
	wire _w2661_ ;
	wire _w2660_ ;
	wire _w2659_ ;
	wire _w2658_ ;
	wire _w2657_ ;
	wire _w2656_ ;
	wire _w2655_ ;
	wire _w2654_ ;
	wire _w2653_ ;
	wire _w2652_ ;
	wire _w2651_ ;
	wire _w2650_ ;
	wire _w2649_ ;
	wire _w2648_ ;
	wire _w2647_ ;
	wire _w2646_ ;
	wire _w2645_ ;
	wire _w2644_ ;
	wire _w2643_ ;
	wire _w2642_ ;
	wire _w2641_ ;
	wire _w2640_ ;
	wire _w2639_ ;
	wire _w2638_ ;
	wire _w2637_ ;
	wire _w2636_ ;
	wire _w2635_ ;
	wire _w2634_ ;
	wire _w2633_ ;
	wire _w2632_ ;
	wire _w2631_ ;
	wire _w2630_ ;
	wire _w2629_ ;
	wire _w2628_ ;
	wire _w2627_ ;
	wire _w2626_ ;
	wire _w2625_ ;
	wire _w2624_ ;
	wire _w2623_ ;
	wire _w2622_ ;
	wire _w2621_ ;
	wire _w2620_ ;
	wire _w2619_ ;
	wire _w2618_ ;
	wire _w2617_ ;
	wire _w2616_ ;
	wire _w2615_ ;
	wire _w1366_ ;
	wire _w1365_ ;
	wire _w1364_ ;
	wire _w1363_ ;
	wire _w1362_ ;
	wire _w1361_ ;
	wire _w1360_ ;
	wire _w1359_ ;
	wire _w1358_ ;
	wire _w1357_ ;
	wire _w1356_ ;
	wire _w1355_ ;
	wire _w1354_ ;
	wire _w1353_ ;
	wire _w1352_ ;
	wire _w1351_ ;
	wire _w1350_ ;
	wire _w1349_ ;
	wire _w1348_ ;
	wire _w1347_ ;
	wire _w1346_ ;
	wire _w1345_ ;
	wire _w1344_ ;
	wire _w1343_ ;
	wire _w1342_ ;
	wire _w1341_ ;
	wire _w1340_ ;
	wire _w1339_ ;
	wire _w1338_ ;
	wire _w1337_ ;
	wire _w1336_ ;
	wire _w1335_ ;
	wire _w1334_ ;
	wire _w1333_ ;
	wire _w1332_ ;
	wire _w1331_ ;
	wire _w1330_ ;
	wire _w1329_ ;
	wire _w1328_ ;
	wire _w1327_ ;
	wire _w1326_ ;
	wire _w1325_ ;
	wire _w1324_ ;
	wire _w1323_ ;
	wire _w1322_ ;
	wire _w1321_ ;
	wire _w1320_ ;
	wire _w1319_ ;
	wire _w1318_ ;
	wire _w1317_ ;
	wire _w1316_ ;
	wire _w1315_ ;
	wire _w1314_ ;
	wire _w1313_ ;
	wire _w1312_ ;
	wire _w1311_ ;
	wire _w1310_ ;
	wire _w1309_ ;
	wire _w1308_ ;
	wire _w1307_ ;
	wire _w1306_ ;
	wire _w1305_ ;
	wire _w1304_ ;
	wire _w1303_ ;
	wire _w1302_ ;
	wire _w1301_ ;
	wire _w1300_ ;
	wire _w1299_ ;
	wire _w1298_ ;
	wire _w1297_ ;
	wire _w1296_ ;
	wire _w1295_ ;
	wire _w1294_ ;
	wire _w1293_ ;
	wire _w1292_ ;
	wire _w1291_ ;
	wire _w1290_ ;
	wire _w1289_ ;
	wire _w1288_ ;
	wire _w1287_ ;
	wire _w1286_ ;
	wire _w1285_ ;
	wire _w1284_ ;
	wire _w1283_ ;
	wire _w1282_ ;
	wire _w1281_ ;
	wire _w1280_ ;
	wire _w1279_ ;
	wire _w1278_ ;
	wire _w1277_ ;
	wire _w1276_ ;
	wire _w1275_ ;
	wire _w1274_ ;
	wire _w1273_ ;
	wire _w1272_ ;
	wire _w1271_ ;
	wire _w1270_ ;
	wire _w1269_ ;
	wire _w1268_ ;
	wire _w1267_ ;
	wire _w1266_ ;
	wire _w1265_ ;
	wire _w1264_ ;
	wire _w1263_ ;
	wire _w1262_ ;
	wire _w1261_ ;
	wire _w1260_ ;
	wire _w1259_ ;
	wire _w1258_ ;
	wire _w1257_ ;
	wire _w1256_ ;
	wire _w1255_ ;
	wire _w1254_ ;
	wire _w1253_ ;
	wire _w1252_ ;
	wire _w1251_ ;
	wire _w1250_ ;
	wire _w1249_ ;
	wire _w1248_ ;
	wire _w1247_ ;
	wire _w1246_ ;
	wire _w1245_ ;
	wire _w1244_ ;
	wire _w1243_ ;
	wire _w1242_ ;
	wire _w1241_ ;
	wire _w1240_ ;
	wire _w1239_ ;
	wire _w1238_ ;
	wire _w1237_ ;
	wire _w1236_ ;
	wire _w1235_ ;
	wire _w1234_ ;
	wire _w1233_ ;
	wire _w1232_ ;
	wire _w1231_ ;
	wire _w1230_ ;
	wire _w1229_ ;
	wire _w1228_ ;
	wire _w1227_ ;
	wire _w1226_ ;
	wire _w1225_ ;
	wire _w1224_ ;
	wire _w1223_ ;
	wire _w1222_ ;
	wire _w1221_ ;
	wire _w1220_ ;
	wire _w1219_ ;
	wire _w1218_ ;
	wire _w1217_ ;
	wire _w1216_ ;
	wire _w1215_ ;
	wire _w1214_ ;
	wire _w1213_ ;
	wire _w1212_ ;
	wire _w1211_ ;
	wire _w1210_ ;
	wire _w1209_ ;
	wire _w1208_ ;
	wire _w1207_ ;
	wire _w1206_ ;
	wire _w1205_ ;
	wire _w1204_ ;
	wire _w1203_ ;
	wire _w1202_ ;
	wire _w1201_ ;
	wire _w1200_ ;
	wire _w1199_ ;
	wire _w1198_ ;
	wire _w1197_ ;
	wire _w1196_ ;
	wire _w1195_ ;
	wire _w1194_ ;
	wire _w1193_ ;
	wire _w1192_ ;
	wire _w1191_ ;
	wire _w1190_ ;
	wire _w1189_ ;
	wire _w1188_ ;
	wire _w1187_ ;
	wire _w1186_ ;
	wire _w1185_ ;
	wire _w1184_ ;
	wire _w1183_ ;
	wire _w1182_ ;
	wire _w1181_ ;
	wire _w1180_ ;
	wire _w1179_ ;
	wire _w1178_ ;
	wire _w1177_ ;
	wire _w1176_ ;
	wire _w1175_ ;
	wire _w1174_ ;
	wire _w1173_ ;
	wire _w1172_ ;
	wire _w1171_ ;
	wire _w1170_ ;
	wire _w1169_ ;
	wire _w1168_ ;
	wire _w1167_ ;
	wire _w1166_ ;
	wire _w1165_ ;
	wire _w1164_ ;
	wire _w1163_ ;
	wire _w1162_ ;
	wire _w1161_ ;
	wire _w1160_ ;
	wire _w1159_ ;
	wire _w1158_ ;
	wire _w1157_ ;
	wire _w1156_ ;
	wire _w1155_ ;
	wire _w1154_ ;
	wire _w1153_ ;
	wire _w1152_ ;
	wire _w1151_ ;
	wire _w1150_ ;
	wire _w1149_ ;
	wire _w1148_ ;
	wire _w1147_ ;
	wire _w1146_ ;
	wire _w1145_ ;
	wire _w1144_ ;
	wire _w1143_ ;
	wire _w1142_ ;
	wire _w1141_ ;
	wire _w1140_ ;
	wire _w1139_ ;
	wire _w1138_ ;
	wire _w1137_ ;
	wire _w1136_ ;
	wire _w1135_ ;
	wire _w1134_ ;
	wire _w1133_ ;
	wire _w1132_ ;
	wire _w1131_ ;
	wire _w1130_ ;
	wire _w1129_ ;
	wire _w1128_ ;
	wire _w1127_ ;
	wire _w1126_ ;
	wire _w1125_ ;
	wire _w1124_ ;
	wire _w1123_ ;
	wire _w1122_ ;
	wire _w1121_ ;
	wire _w1120_ ;
	wire _w1119_ ;
	wire _w1118_ ;
	wire _w1117_ ;
	wire _w1116_ ;
	wire _w1115_ ;
	wire _w1114_ ;
	wire _w1113_ ;
	wire _w1112_ ;
	wire _w1111_ ;
	wire _w1110_ ;
	wire _w1109_ ;
	wire _w1108_ ;
	wire _w1107_ ;
	wire _w1106_ ;
	wire _w1105_ ;
	wire _w1104_ ;
	wire _w1103_ ;
	wire _w1102_ ;
	wire _w1101_ ;
	wire _w1100_ ;
	wire _w1099_ ;
	wire _w1098_ ;
	wire _w1097_ ;
	wire _w1096_ ;
	wire _w1095_ ;
	wire _w1094_ ;
	wire _w1093_ ;
	wire _w1092_ ;
	wire _w1091_ ;
	wire _w1090_ ;
	wire _w1089_ ;
	wire _w1088_ ;
	wire _w1087_ ;
	wire _w1086_ ;
	wire _w1085_ ;
	wire _w1084_ ;
	wire _w1083_ ;
	wire _w1082_ ;
	wire _w1081_ ;
	wire _w1080_ ;
	wire _w1079_ ;
	wire _w1078_ ;
	wire _w1077_ ;
	wire _w1076_ ;
	wire _w1075_ ;
	wire _w1074_ ;
	wire _w1073_ ;
	wire _w1072_ ;
	wire _w1071_ ;
	wire _w1070_ ;
	wire _w1069_ ;
	wire _w1068_ ;
	wire _w1067_ ;
	wire _w1066_ ;
	wire _w1065_ ;
	wire _w1064_ ;
	wire _w1063_ ;
	wire _w1062_ ;
	wire _w1061_ ;
	wire _w1060_ ;
	wire _w1059_ ;
	wire _w1058_ ;
	wire _w1057_ ;
	wire _w1056_ ;
	wire _w1055_ ;
	wire _w1054_ ;
	wire _w1053_ ;
	wire _w1052_ ;
	wire _w1051_ ;
	wire _w1050_ ;
	wire _w1049_ ;
	wire _w1048_ ;
	wire _w1047_ ;
	wire _w1046_ ;
	wire _w1045_ ;
	wire _w1044_ ;
	wire _w1043_ ;
	wire _w1042_ ;
	wire _w1041_ ;
	wire _w1040_ ;
	wire _w1039_ ;
	wire _w1038_ ;
	wire _w1037_ ;
	wire _w1036_ ;
	wire _w1035_ ;
	wire _w1034_ ;
	wire _w1033_ ;
	wire _w1032_ ;
	wire _w1031_ ;
	wire _w1030_ ;
	wire _w1029_ ;
	wire _w1028_ ;
	wire _w1027_ ;
	wire _w1026_ ;
	wire _w1025_ ;
	wire _w1024_ ;
	wire _w1023_ ;
	wire _w1022_ ;
	wire _w1021_ ;
	wire _w1020_ ;
	wire _w1019_ ;
	wire _w1018_ ;
	wire _w1017_ ;
	wire _w1016_ ;
	wire _w1015_ ;
	wire _w1014_ ;
	wire _w1013_ ;
	wire _w1012_ ;
	wire _w1011_ ;
	wire _w1010_ ;
	wire _w1009_ ;
	wire _w1008_ ;
	wire _w1007_ ;
	wire _w1006_ ;
	wire _w1005_ ;
	wire _w1004_ ;
	wire _w1003_ ;
	wire _w1002_ ;
	wire _w1001_ ;
	wire _w1000_ ;
	wire _w999_ ;
	wire _w998_ ;
	wire _w997_ ;
	wire _w996_ ;
	wire _w995_ ;
	wire _w994_ ;
	wire _w993_ ;
	wire _w992_ ;
	wire _w991_ ;
	wire _w990_ ;
	wire _w989_ ;
	wire _w988_ ;
	wire _w987_ ;
	wire _w986_ ;
	wire _w985_ ;
	wire _w984_ ;
	wire _w983_ ;
	wire _w982_ ;
	wire _w981_ ;
	wire _w980_ ;
	wire _w979_ ;
	wire _w978_ ;
	wire _w977_ ;
	wire _w976_ ;
	wire _w975_ ;
	wire _w974_ ;
	wire _w973_ ;
	wire _w972_ ;
	wire _w971_ ;
	wire _w970_ ;
	wire _w969_ ;
	wire _w968_ ;
	wire _w967_ ;
	wire _w966_ ;
	wire _w965_ ;
	wire _w964_ ;
	wire _w963_ ;
	wire _w962_ ;
	wire _w961_ ;
	wire _w960_ ;
	wire _w959_ ;
	wire _w958_ ;
	wire _w957_ ;
	wire _w956_ ;
	wire _w955_ ;
	wire _w954_ ;
	wire _w953_ ;
	wire _w952_ ;
	wire _w951_ ;
	wire _w950_ ;
	wire _w949_ ;
	wire _w948_ ;
	wire _w947_ ;
	wire _w946_ ;
	wire _w945_ ;
	wire _w944_ ;
	wire _w943_ ;
	wire _w942_ ;
	wire _w941_ ;
	wire _w940_ ;
	wire _w939_ ;
	wire _w938_ ;
	wire _w937_ ;
	wire _w936_ ;
	wire _w935_ ;
	wire _w934_ ;
	wire _w933_ ;
	wire _w932_ ;
	wire _w931_ ;
	wire _w930_ ;
	wire _w929_ ;
	wire _w928_ ;
	wire _w927_ ;
	wire _w926_ ;
	wire _w925_ ;
	wire _w924_ ;
	wire _w923_ ;
	wire _w922_ ;
	wire _w921_ ;
	wire _w920_ ;
	wire _w919_ ;
	wire _w918_ ;
	wire _w917_ ;
	wire _w916_ ;
	wire _w915_ ;
	wire _w914_ ;
	wire _w913_ ;
	wire _w912_ ;
	wire _w911_ ;
	wire _w910_ ;
	wire _w909_ ;
	wire _w908_ ;
	wire _w907_ ;
	wire _w906_ ;
	wire _w905_ ;
	wire _w904_ ;
	wire _w903_ ;
	wire _w902_ ;
	wire _w901_ ;
	wire _w900_ ;
	wire _w899_ ;
	wire _w898_ ;
	wire _w897_ ;
	wire _w896_ ;
	wire _w895_ ;
	wire _w894_ ;
	wire _w893_ ;
	wire _w892_ ;
	wire _w891_ ;
	wire _w890_ ;
	wire _w889_ ;
	wire _w888_ ;
	wire _w887_ ;
	wire _w886_ ;
	wire _w885_ ;
	wire _w884_ ;
	wire _w883_ ;
	wire _w882_ ;
	wire _w881_ ;
	wire _w880_ ;
	wire _w879_ ;
	wire _w878_ ;
	wire _w877_ ;
	wire _w876_ ;
	wire _w875_ ;
	wire _w874_ ;
	wire _w873_ ;
	wire _w872_ ;
	wire _w871_ ;
	wire _w870_ ;
	wire _w869_ ;
	wire _w868_ ;
	wire _w867_ ;
	wire _w866_ ;
	wire _w865_ ;
	wire _w864_ ;
	wire _w863_ ;
	wire _w862_ ;
	wire _w861_ ;
	wire _w860_ ;
	wire _w859_ ;
	wire _w858_ ;
	wire _w857_ ;
	wire _w856_ ;
	wire _w855_ ;
	wire _w854_ ;
	wire _w853_ ;
	wire _w852_ ;
	wire _w851_ ;
	wire _w850_ ;
	wire _w849_ ;
	wire _w848_ ;
	wire _w847_ ;
	wire _w846_ ;
	wire _w845_ ;
	wire _w844_ ;
	wire _w843_ ;
	wire _w842_ ;
	wire _w841_ ;
	wire _w840_ ;
	wire _w839_ ;
	wire _w838_ ;
	wire _w837_ ;
	wire _w836_ ;
	wire _w835_ ;
	wire _w834_ ;
	wire _w833_ ;
	wire _w832_ ;
	wire _w831_ ;
	wire _w830_ ;
	wire _w829_ ;
	wire _w828_ ;
	wire _w827_ ;
	wire _w826_ ;
	wire _w825_ ;
	wire _w824_ ;
	wire _w823_ ;
	wire _w822_ ;
	wire _w821_ ;
	wire _w820_ ;
	wire _w819_ ;
	wire _w818_ ;
	wire _w817_ ;
	wire _w816_ ;
	wire _w815_ ;
	wire _w814_ ;
	wire _w813_ ;
	wire _w812_ ;
	wire _w811_ ;
	wire _w810_ ;
	wire _w809_ ;
	wire _w808_ ;
	wire _w807_ ;
	wire _w806_ ;
	wire _w805_ ;
	wire _w804_ ;
	wire _w803_ ;
	wire _w802_ ;
	wire _w801_ ;
	wire _w800_ ;
	wire _w799_ ;
	wire _w514_ ;
	wire _w513_ ;
	wire _w512_ ;
	wire _w511_ ;
	wire _w510_ ;
	wire _w509_ ;
	wire _w508_ ;
	wire _w507_ ;
	wire _w506_ ;
	wire _w505_ ;
	wire _w504_ ;
	wire _w503_ ;
	wire _w502_ ;
	wire _w501_ ;
	wire _w500_ ;
	wire _w499_ ;
	wire _w498_ ;
	wire _w497_ ;
	wire _w496_ ;
	wire _w495_ ;
	wire _w494_ ;
	wire _w493_ ;
	wire _w492_ ;
	wire _w491_ ;
	wire _w490_ ;
	wire _w489_ ;
	wire _w488_ ;
	wire _w487_ ;
	wire _w486_ ;
	wire _w485_ ;
	wire _w484_ ;
	wire _w483_ ;
	wire _w482_ ;
	wire _w481_ ;
	wire _w480_ ;
	wire _w479_ ;
	wire _w478_ ;
	wire _w477_ ;
	wire _w476_ ;
	wire _w475_ ;
	wire _w474_ ;
	wire _w473_ ;
	wire _w472_ ;
	wire _w471_ ;
	wire _w470_ ;
	wire _w469_ ;
	wire _w468_ ;
	wire _w467_ ;
	wire _w466_ ;
	wire _w465_ ;
	wire _w464_ ;
	wire _w463_ ;
	wire _w462_ ;
	wire _w461_ ;
	wire _w460_ ;
	wire _w459_ ;
	wire _w458_ ;
	wire _w457_ ;
	wire _w456_ ;
	wire _w455_ ;
	wire _w454_ ;
	wire _w453_ ;
	wire _w452_ ;
	wire _w451_ ;
	wire _w450_ ;
	wire _w449_ ;
	wire _w448_ ;
	wire _w447_ ;
	wire _w446_ ;
	wire _w445_ ;
	wire _w444_ ;
	wire _w443_ ;
	wire _w442_ ;
	wire _w441_ ;
	wire _w440_ ;
	wire _w439_ ;
	wire _w438_ ;
	wire _w437_ ;
	wire _w436_ ;
	wire _w435_ ;
	wire _w434_ ;
	wire _w433_ ;
	wire _w432_ ;
	wire _w431_ ;
	wire _w430_ ;
	wire _w429_ ;
	wire _w428_ ;
	wire _w427_ ;
	wire _w426_ ;
	wire _w425_ ;
	wire _w424_ ;
	wire _w423_ ;
	wire _w422_ ;
	wire _w421_ ;
	wire _w420_ ;
	wire _w419_ ;
	wire _w418_ ;
	wire _w417_ ;
	wire _w416_ ;
	wire _w415_ ;
	wire _w414_ ;
	wire _w413_ ;
	wire _w412_ ;
	wire _w411_ ;
	wire _w410_ ;
	wire _w409_ ;
	wire _w408_ ;
	wire _w407_ ;
	wire _w406_ ;
	wire _w405_ ;
	wire _w404_ ;
	wire _w403_ ;
	wire _w402_ ;
	wire _w401_ ;
	wire _w400_ ;
	wire _w399_ ;
	wire _w398_ ;
	wire _w397_ ;
	wire _w396_ ;
	wire _w395_ ;
	wire _w394_ ;
	wire _w393_ ;
	wire _w392_ ;
	wire _w391_ ;
	wire _w390_ ;
	wire _w389_ ;
	wire _w388_ ;
	wire _w387_ ;
	wire _w386_ ;
	wire _w385_ ;
	wire _w316_ ;
	wire _w315_ ;
	wire _w314_ ;
	wire _w313_ ;
	wire _w312_ ;
	wire _w311_ ;
	wire _w310_ ;
	wire _w309_ ;
	wire _w308_ ;
	wire _w307_ ;
	wire _w306_ ;
	wire _w305_ ;
	wire _w304_ ;
	wire _w303_ ;
	wire _w302_ ;
	wire _w301_ ;
	wire _w300_ ;
	wire _w299_ ;
	wire _w298_ ;
	wire _w297_ ;
	wire _w296_ ;
	wire _w295_ ;
	wire _w294_ ;
	wire _w293_ ;
	wire _w292_ ;
	wire _w291_ ;
	wire _w290_ ;
	wire _w289_ ;
	wire _w288_ ;
	wire _w287_ ;
	wire _w270_ ;
	wire _w269_ ;
	wire _w268_ ;
	wire _w267_ ;
	wire _w266_ ;
	wire _w265_ ;
	wire _w264_ ;
	wire _w263_ ;
	wire _w262_ ;
	wire _w261_ ;
	wire _w260_ ;
	wire _w259_ ;
	wire _w258_ ;
	wire _w271_ ;
	wire _w272_ ;
	wire _w273_ ;
	wire _w274_ ;
	wire _w275_ ;
	wire _w276_ ;
	wire _w277_ ;
	wire _w278_ ;
	wire _w279_ ;
	wire _w280_ ;
	wire _w281_ ;
	wire _w282_ ;
	wire _w283_ ;
	wire _w284_ ;
	wire _w285_ ;
	wire _w286_ ;
	wire _w317_ ;
	wire _w318_ ;
	wire _w319_ ;
	wire _w320_ ;
	wire _w321_ ;
	wire _w322_ ;
	wire _w323_ ;
	wire _w324_ ;
	wire _w325_ ;
	wire _w326_ ;
	wire _w327_ ;
	wire _w328_ ;
	wire _w329_ ;
	wire _w330_ ;
	wire _w331_ ;
	wire _w332_ ;
	wire _w333_ ;
	wire _w334_ ;
	wire _w335_ ;
	wire _w336_ ;
	wire _w337_ ;
	wire _w338_ ;
	wire _w339_ ;
	wire _w340_ ;
	wire _w341_ ;
	wire _w342_ ;
	wire _w343_ ;
	wire _w344_ ;
	wire _w345_ ;
	wire _w346_ ;
	wire _w347_ ;
	wire _w348_ ;
	wire _w349_ ;
	wire _w350_ ;
	wire _w351_ ;
	wire _w352_ ;
	wire _w353_ ;
	wire _w354_ ;
	wire _w355_ ;
	wire _w356_ ;
	wire _w357_ ;
	wire _w358_ ;
	wire _w359_ ;
	wire _w360_ ;
	wire _w361_ ;
	wire _w362_ ;
	wire _w363_ ;
	wire _w364_ ;
	wire _w365_ ;
	wire _w366_ ;
	wire _w367_ ;
	wire _w368_ ;
	wire _w369_ ;
	wire _w370_ ;
	wire _w371_ ;
	wire _w372_ ;
	wire _w373_ ;
	wire _w374_ ;
	wire _w375_ ;
	wire _w376_ ;
	wire _w377_ ;
	wire _w378_ ;
	wire _w379_ ;
	wire _w380_ ;
	wire _w381_ ;
	wire _w382_ ;
	wire _w383_ ;
	wire _w384_ ;
	wire _w515_ ;
	wire _w516_ ;
	wire _w517_ ;
	wire _w518_ ;
	wire _w519_ ;
	wire _w520_ ;
	wire _w521_ ;
	wire _w522_ ;
	wire _w523_ ;
	wire _w524_ ;
	wire _w525_ ;
	wire _w526_ ;
	wire _w527_ ;
	wire _w528_ ;
	wire _w529_ ;
	wire _w530_ ;
	wire _w531_ ;
	wire _w532_ ;
	wire _w533_ ;
	wire _w534_ ;
	wire _w535_ ;
	wire _w536_ ;
	wire _w537_ ;
	wire _w538_ ;
	wire _w539_ ;
	wire _w540_ ;
	wire _w541_ ;
	wire _w542_ ;
	wire _w543_ ;
	wire _w544_ ;
	wire _w545_ ;
	wire _w546_ ;
	wire _w547_ ;
	wire _w548_ ;
	wire _w549_ ;
	wire _w550_ ;
	wire _w551_ ;
	wire _w552_ ;
	wire _w553_ ;
	wire _w554_ ;
	wire _w555_ ;
	wire _w556_ ;
	wire _w557_ ;
	wire _w558_ ;
	wire _w559_ ;
	wire _w560_ ;
	wire _w561_ ;
	wire _w562_ ;
	wire _w563_ ;
	wire _w564_ ;
	wire _w565_ ;
	wire _w566_ ;
	wire _w567_ ;
	wire _w568_ ;
	wire _w569_ ;
	wire _w570_ ;
	wire _w571_ ;
	wire _w572_ ;
	wire _w573_ ;
	wire _w574_ ;
	wire _w575_ ;
	wire _w576_ ;
	wire _w577_ ;
	wire _w578_ ;
	wire _w579_ ;
	wire _w580_ ;
	wire _w581_ ;
	wire _w582_ ;
	wire _w583_ ;
	wire _w584_ ;
	wire _w585_ ;
	wire _w586_ ;
	wire _w587_ ;
	wire _w588_ ;
	wire _w589_ ;
	wire _w590_ ;
	wire _w591_ ;
	wire _w592_ ;
	wire _w593_ ;
	wire _w594_ ;
	wire _w595_ ;
	wire _w596_ ;
	wire _w597_ ;
	wire _w598_ ;
	wire _w599_ ;
	wire _w600_ ;
	wire _w601_ ;
	wire _w602_ ;
	wire _w603_ ;
	wire _w604_ ;
	wire _w605_ ;
	wire _w606_ ;
	wire _w607_ ;
	wire _w608_ ;
	wire _w609_ ;
	wire _w610_ ;
	wire _w611_ ;
	wire _w612_ ;
	wire _w613_ ;
	wire _w614_ ;
	wire _w615_ ;
	wire _w616_ ;
	wire _w617_ ;
	wire _w618_ ;
	wire _w619_ ;
	wire _w620_ ;
	wire _w621_ ;
	wire _w622_ ;
	wire _w623_ ;
	wire _w624_ ;
	wire _w625_ ;
	wire _w626_ ;
	wire _w627_ ;
	wire _w628_ ;
	wire _w629_ ;
	wire _w630_ ;
	wire _w631_ ;
	wire _w632_ ;
	wire _w633_ ;
	wire _w634_ ;
	wire _w635_ ;
	wire _w636_ ;
	wire _w637_ ;
	wire _w638_ ;
	wire _w639_ ;
	wire _w640_ ;
	wire _w641_ ;
	wire _w642_ ;
	wire _w643_ ;
	wire _w644_ ;
	wire _w645_ ;
	wire _w646_ ;
	wire _w647_ ;
	wire _w648_ ;
	wire _w649_ ;
	wire _w650_ ;
	wire _w651_ ;
	wire _w652_ ;
	wire _w653_ ;
	wire _w654_ ;
	wire _w655_ ;
	wire _w656_ ;
	wire _w657_ ;
	wire _w658_ ;
	wire _w659_ ;
	wire _w660_ ;
	wire _w661_ ;
	wire _w662_ ;
	wire _w663_ ;
	wire _w664_ ;
	wire _w665_ ;
	wire _w666_ ;
	wire _w667_ ;
	wire _w668_ ;
	wire _w669_ ;
	wire _w670_ ;
	wire _w671_ ;
	wire _w672_ ;
	wire _w673_ ;
	wire _w674_ ;
	wire _w675_ ;
	wire _w676_ ;
	wire _w677_ ;
	wire _w678_ ;
	wire _w679_ ;
	wire _w680_ ;
	wire _w681_ ;
	wire _w682_ ;
	wire _w683_ ;
	wire _w684_ ;
	wire _w685_ ;
	wire _w686_ ;
	wire _w687_ ;
	wire _w688_ ;
	wire _w689_ ;
	wire _w690_ ;
	wire _w691_ ;
	wire _w692_ ;
	wire _w693_ ;
	wire _w694_ ;
	wire _w695_ ;
	wire _w696_ ;
	wire _w697_ ;
	wire _w698_ ;
	wire _w699_ ;
	wire _w700_ ;
	wire _w701_ ;
	wire _w702_ ;
	wire _w703_ ;
	wire _w704_ ;
	wire _w705_ ;
	wire _w706_ ;
	wire _w707_ ;
	wire _w708_ ;
	wire _w709_ ;
	wire _w710_ ;
	wire _w711_ ;
	wire _w712_ ;
	wire _w713_ ;
	wire _w714_ ;
	wire _w715_ ;
	wire _w716_ ;
	wire _w717_ ;
	wire _w718_ ;
	wire _w719_ ;
	wire _w720_ ;
	wire _w721_ ;
	wire _w722_ ;
	wire _w723_ ;
	wire _w724_ ;
	wire _w725_ ;
	wire _w726_ ;
	wire _w727_ ;
	wire _w728_ ;
	wire _w729_ ;
	wire _w730_ ;
	wire _w731_ ;
	wire _w732_ ;
	wire _w733_ ;
	wire _w734_ ;
	wire _w735_ ;
	wire _w736_ ;
	wire _w737_ ;
	wire _w738_ ;
	wire _w739_ ;
	wire _w740_ ;
	wire _w741_ ;
	wire _w742_ ;
	wire _w743_ ;
	wire _w744_ ;
	wire _w745_ ;
	wire _w746_ ;
	wire _w747_ ;
	wire _w748_ ;
	wire _w749_ ;
	wire _w750_ ;
	wire _w751_ ;
	wire _w752_ ;
	wire _w753_ ;
	wire _w754_ ;
	wire _w755_ ;
	wire _w756_ ;
	wire _w757_ ;
	wire _w758_ ;
	wire _w759_ ;
	wire _w760_ ;
	wire _w761_ ;
	wire _w762_ ;
	wire _w763_ ;
	wire _w764_ ;
	wire _w765_ ;
	wire _w766_ ;
	wire _w767_ ;
	wire _w768_ ;
	wire _w769_ ;
	wire _w770_ ;
	wire _w771_ ;
	wire _w772_ ;
	wire _w773_ ;
	wire _w774_ ;
	wire _w775_ ;
	wire _w776_ ;
	wire _w777_ ;
	wire _w778_ ;
	wire _w779_ ;
	wire _w780_ ;
	wire _w781_ ;
	wire _w782_ ;
	wire _w783_ ;
	wire _w784_ ;
	wire _w785_ ;
	wire _w786_ ;
	wire _w787_ ;
	wire _w788_ ;
	wire _w789_ ;
	wire _w790_ ;
	wire _w791_ ;
	wire _w792_ ;
	wire _w793_ ;
	wire _w794_ ;
	wire _w795_ ;
	wire _w796_ ;
	wire _w797_ ;
	wire _w798_ ;
	wire _w1367_ ;
	wire _w1368_ ;
	wire _w1369_ ;
	wire _w1370_ ;
	wire _w1371_ ;
	wire _w1372_ ;
	wire _w1373_ ;
	wire _w1374_ ;
	wire _w1375_ ;
	wire _w1376_ ;
	wire _w1377_ ;
	wire _w1378_ ;
	wire _w1379_ ;
	wire _w1380_ ;
	wire _w1381_ ;
	wire _w1382_ ;
	wire _w1383_ ;
	wire _w1384_ ;
	wire _w1385_ ;
	wire _w1386_ ;
	wire _w1387_ ;
	wire _w1388_ ;
	wire _w1389_ ;
	wire _w1390_ ;
	wire _w1391_ ;
	wire _w1392_ ;
	wire _w1393_ ;
	wire _w1394_ ;
	wire _w1395_ ;
	wire _w1396_ ;
	wire _w1397_ ;
	wire _w1398_ ;
	wire _w1399_ ;
	wire _w1400_ ;
	wire _w1401_ ;
	wire _w1402_ ;
	wire _w1403_ ;
	wire _w1404_ ;
	wire _w1405_ ;
	wire _w1406_ ;
	wire _w1407_ ;
	wire _w1408_ ;
	wire _w1409_ ;
	wire _w1410_ ;
	wire _w1411_ ;
	wire _w1412_ ;
	wire _w1413_ ;
	wire _w1414_ ;
	wire _w1415_ ;
	wire _w1416_ ;
	wire _w1417_ ;
	wire _w1418_ ;
	wire _w1419_ ;
	wire _w1420_ ;
	wire _w1421_ ;
	wire _w1422_ ;
	wire _w1423_ ;
	wire _w1424_ ;
	wire _w1425_ ;
	wire _w1426_ ;
	wire _w1427_ ;
	wire _w1428_ ;
	wire _w1429_ ;
	wire _w1430_ ;
	wire _w1431_ ;
	wire _w1432_ ;
	wire _w1433_ ;
	wire _w1434_ ;
	wire _w1435_ ;
	wire _w1436_ ;
	wire _w1437_ ;
	wire _w1438_ ;
	wire _w1439_ ;
	wire _w1440_ ;
	wire _w1441_ ;
	wire _w1442_ ;
	wire _w1443_ ;
	wire _w1444_ ;
	wire _w1445_ ;
	wire _w1446_ ;
	wire _w1447_ ;
	wire _w1448_ ;
	wire _w1449_ ;
	wire _w1450_ ;
	wire _w1451_ ;
	wire _w1452_ ;
	wire _w1453_ ;
	wire _w1454_ ;
	wire _w1455_ ;
	wire _w1456_ ;
	wire _w1457_ ;
	wire _w1458_ ;
	wire _w1459_ ;
	wire _w1460_ ;
	wire _w1461_ ;
	wire _w1462_ ;
	wire _w1463_ ;
	wire _w1464_ ;
	wire _w1465_ ;
	wire _w1466_ ;
	wire _w1467_ ;
	wire _w1468_ ;
	wire _w1469_ ;
	wire _w1470_ ;
	wire _w1471_ ;
	wire _w1472_ ;
	wire _w1473_ ;
	wire _w1474_ ;
	wire _w1475_ ;
	wire _w1476_ ;
	wire _w1477_ ;
	wire _w1478_ ;
	wire _w1479_ ;
	wire _w1480_ ;
	wire _w1481_ ;
	wire _w1482_ ;
	wire _w1483_ ;
	wire _w1484_ ;
	wire _w1485_ ;
	wire _w1486_ ;
	wire _w1487_ ;
	wire _w1488_ ;
	wire _w1489_ ;
	wire _w1490_ ;
	wire _w1491_ ;
	wire _w1492_ ;
	wire _w1493_ ;
	wire _w1494_ ;
	wire _w1495_ ;
	wire _w1496_ ;
	wire _w1497_ ;
	wire _w1498_ ;
	wire _w1499_ ;
	wire _w1500_ ;
	wire _w1501_ ;
	wire _w1502_ ;
	wire _w1503_ ;
	wire _w1504_ ;
	wire _w1505_ ;
	wire _w1506_ ;
	wire _w1507_ ;
	wire _w1508_ ;
	wire _w1509_ ;
	wire _w1510_ ;
	wire _w1511_ ;
	wire _w1512_ ;
	wire _w1513_ ;
	wire _w1514_ ;
	wire _w1515_ ;
	wire _w1516_ ;
	wire _w1517_ ;
	wire _w1518_ ;
	wire _w1519_ ;
	wire _w1520_ ;
	wire _w1521_ ;
	wire _w1522_ ;
	wire _w1523_ ;
	wire _w1524_ ;
	wire _w1525_ ;
	wire _w1526_ ;
	wire _w1527_ ;
	wire _w1528_ ;
	wire _w1529_ ;
	wire _w1530_ ;
	wire _w1531_ ;
	wire _w1532_ ;
	wire _w1533_ ;
	wire _w1534_ ;
	wire _w1535_ ;
	wire _w1536_ ;
	wire _w1537_ ;
	wire _w1538_ ;
	wire _w1539_ ;
	wire _w1540_ ;
	wire _w1541_ ;
	wire _w1542_ ;
	wire _w1543_ ;
	wire _w1544_ ;
	wire _w1545_ ;
	wire _w1546_ ;
	wire _w1547_ ;
	wire _w1548_ ;
	wire _w1549_ ;
	wire _w1550_ ;
	wire _w1551_ ;
	wire _w1552_ ;
	wire _w1553_ ;
	wire _w1554_ ;
	wire _w1555_ ;
	wire _w1556_ ;
	wire _w1557_ ;
	wire _w1558_ ;
	wire _w1559_ ;
	wire _w1560_ ;
	wire _w1561_ ;
	wire _w1562_ ;
	wire _w1563_ ;
	wire _w1564_ ;
	wire _w1565_ ;
	wire _w1566_ ;
	wire _w1567_ ;
	wire _w1568_ ;
	wire _w1569_ ;
	wire _w1570_ ;
	wire _w1571_ ;
	wire _w1572_ ;
	wire _w1573_ ;
	wire _w1574_ ;
	wire _w1575_ ;
	wire _w1576_ ;
	wire _w1577_ ;
	wire _w1578_ ;
	wire _w1579_ ;
	wire _w1580_ ;
	wire _w1581_ ;
	wire _w1582_ ;
	wire _w1583_ ;
	wire _w1584_ ;
	wire _w1585_ ;
	wire _w1586_ ;
	wire _w1587_ ;
	wire _w1588_ ;
	wire _w1589_ ;
	wire _w1590_ ;
	wire _w1591_ ;
	wire _w1592_ ;
	wire _w1593_ ;
	wire _w1594_ ;
	wire _w1595_ ;
	wire _w1596_ ;
	wire _w1597_ ;
	wire _w1598_ ;
	wire _w1599_ ;
	wire _w1600_ ;
	wire _w1601_ ;
	wire _w1602_ ;
	wire _w1603_ ;
	wire _w1604_ ;
	wire _w1605_ ;
	wire _w1606_ ;
	wire _w1607_ ;
	wire _w1608_ ;
	wire _w1609_ ;
	wire _w1610_ ;
	wire _w1611_ ;
	wire _w1612_ ;
	wire _w1613_ ;
	wire _w1614_ ;
	wire _w1615_ ;
	wire _w1616_ ;
	wire _w1617_ ;
	wire _w1618_ ;
	wire _w1619_ ;
	wire _w1620_ ;
	wire _w1621_ ;
	wire _w1622_ ;
	wire _w1623_ ;
	wire _w1624_ ;
	wire _w1625_ ;
	wire _w1626_ ;
	wire _w1627_ ;
	wire _w1628_ ;
	wire _w1629_ ;
	wire _w1630_ ;
	wire _w1631_ ;
	wire _w1632_ ;
	wire _w1633_ ;
	wire _w1634_ ;
	wire _w1635_ ;
	wire _w1636_ ;
	wire _w1637_ ;
	wire _w1638_ ;
	wire _w1639_ ;
	wire _w1640_ ;
	wire _w1641_ ;
	wire _w1642_ ;
	wire _w1643_ ;
	wire _w1644_ ;
	wire _w1645_ ;
	wire _w1646_ ;
	wire _w1647_ ;
	wire _w1648_ ;
	wire _w1649_ ;
	wire _w1650_ ;
	wire _w1651_ ;
	wire _w1652_ ;
	wire _w1653_ ;
	wire _w1654_ ;
	wire _w1655_ ;
	wire _w1656_ ;
	wire _w1657_ ;
	wire _w1658_ ;
	wire _w1659_ ;
	wire _w1660_ ;
	wire _w1661_ ;
	wire _w1662_ ;
	wire _w1663_ ;
	wire _w1664_ ;
	wire _w1665_ ;
	wire _w1666_ ;
	wire _w1667_ ;
	wire _w1668_ ;
	wire _w1669_ ;
	wire _w1670_ ;
	wire _w1671_ ;
	wire _w1672_ ;
	wire _w1673_ ;
	wire _w1674_ ;
	wire _w1675_ ;
	wire _w1676_ ;
	wire _w1677_ ;
	wire _w1678_ ;
	wire _w1679_ ;
	wire _w1680_ ;
	wire _w1681_ ;
	wire _w1682_ ;
	wire _w1683_ ;
	wire _w1684_ ;
	wire _w1685_ ;
	wire _w1686_ ;
	wire _w1687_ ;
	wire _w1688_ ;
	wire _w1689_ ;
	wire _w1690_ ;
	wire _w1691_ ;
	wire _w1692_ ;
	wire _w1693_ ;
	wire _w1694_ ;
	wire _w1695_ ;
	wire _w1696_ ;
	wire _w1697_ ;
	wire _w1698_ ;
	wire _w1699_ ;
	wire _w1700_ ;
	wire _w1701_ ;
	wire _w1702_ ;
	wire _w1703_ ;
	wire _w1704_ ;
	wire _w1705_ ;
	wire _w1706_ ;
	wire _w1707_ ;
	wire _w1708_ ;
	wire _w1709_ ;
	wire _w1710_ ;
	wire _w1711_ ;
	wire _w1712_ ;
	wire _w1713_ ;
	wire _w1714_ ;
	wire _w1715_ ;
	wire _w1716_ ;
	wire _w1717_ ;
	wire _w1718_ ;
	wire _w1719_ ;
	wire _w1720_ ;
	wire _w1721_ ;
	wire _w1722_ ;
	wire _w1723_ ;
	wire _w1724_ ;
	wire _w1725_ ;
	wire _w1726_ ;
	wire _w1727_ ;
	wire _w1728_ ;
	wire _w1729_ ;
	wire _w1730_ ;
	wire _w1731_ ;
	wire _w1732_ ;
	wire _w1733_ ;
	wire _w1734_ ;
	wire _w1735_ ;
	wire _w1736_ ;
	wire _w1737_ ;
	wire _w1738_ ;
	wire _w1739_ ;
	wire _w1740_ ;
	wire _w1741_ ;
	wire _w1742_ ;
	wire _w1743_ ;
	wire _w1744_ ;
	wire _w1745_ ;
	wire _w1746_ ;
	wire _w1747_ ;
	wire _w1748_ ;
	wire _w1749_ ;
	wire _w1750_ ;
	wire _w1751_ ;
	wire _w1752_ ;
	wire _w1753_ ;
	wire _w1754_ ;
	wire _w1755_ ;
	wire _w1756_ ;
	wire _w1757_ ;
	wire _w1758_ ;
	wire _w1759_ ;
	wire _w1760_ ;
	wire _w1761_ ;
	wire _w1762_ ;
	wire _w1763_ ;
	wire _w1764_ ;
	wire _w1765_ ;
	wire _w1766_ ;
	wire _w1767_ ;
	wire _w1768_ ;
	wire _w1769_ ;
	wire _w1770_ ;
	wire _w1771_ ;
	wire _w1772_ ;
	wire _w1773_ ;
	wire _w1774_ ;
	wire _w1775_ ;
	wire _w1776_ ;
	wire _w1777_ ;
	wire _w1778_ ;
	wire _w1779_ ;
	wire _w1780_ ;
	wire _w1781_ ;
	wire _w1782_ ;
	wire _w1783_ ;
	wire _w1784_ ;
	wire _w1785_ ;
	wire _w1786_ ;
	wire _w1787_ ;
	wire _w1788_ ;
	wire _w1789_ ;
	wire _w1790_ ;
	wire _w1791_ ;
	wire _w1792_ ;
	wire _w1793_ ;
	wire _w1794_ ;
	wire _w1795_ ;
	wire _w1796_ ;
	wire _w1797_ ;
	wire _w1798_ ;
	wire _w1799_ ;
	wire _w1800_ ;
	wire _w1801_ ;
	wire _w1802_ ;
	wire _w1803_ ;
	wire _w1804_ ;
	wire _w1805_ ;
	wire _w1806_ ;
	wire _w1807_ ;
	wire _w1808_ ;
	wire _w1809_ ;
	wire _w1810_ ;
	wire _w1811_ ;
	wire _w1812_ ;
	wire _w1813_ ;
	wire _w1814_ ;
	wire _w1815_ ;
	wire _w1816_ ;
	wire _w1817_ ;
	wire _w1818_ ;
	wire _w1819_ ;
	wire _w1820_ ;
	wire _w1821_ ;
	wire _w1822_ ;
	wire _w1823_ ;
	wire _w1824_ ;
	wire _w1825_ ;
	wire _w1826_ ;
	wire _w1827_ ;
	wire _w1828_ ;
	wire _w1829_ ;
	wire _w1830_ ;
	wire _w1831_ ;
	wire _w1832_ ;
	wire _w1833_ ;
	wire _w1834_ ;
	wire _w1835_ ;
	wire _w1836_ ;
	wire _w1837_ ;
	wire _w1838_ ;
	wire _w1839_ ;
	wire _w1840_ ;
	wire _w1841_ ;
	wire _w1842_ ;
	wire _w1843_ ;
	wire _w1844_ ;
	wire _w1845_ ;
	wire _w1846_ ;
	wire _w1847_ ;
	wire _w1848_ ;
	wire _w1849_ ;
	wire _w1850_ ;
	wire _w1851_ ;
	wire _w1852_ ;
	wire _w1853_ ;
	wire _w1854_ ;
	wire _w1855_ ;
	wire _w1856_ ;
	wire _w1857_ ;
	wire _w1858_ ;
	wire _w1859_ ;
	wire _w1860_ ;
	wire _w1861_ ;
	wire _w1862_ ;
	wire _w1863_ ;
	wire _w1864_ ;
	wire _w1865_ ;
	wire _w1866_ ;
	wire _w1867_ ;
	wire _w1868_ ;
	wire _w1869_ ;
	wire _w1870_ ;
	wire _w1871_ ;
	wire _w1872_ ;
	wire _w1873_ ;
	wire _w1874_ ;
	wire _w1875_ ;
	wire _w1876_ ;
	wire _w1877_ ;
	wire _w1878_ ;
	wire _w1879_ ;
	wire _w1880_ ;
	wire _w1881_ ;
	wire _w1882_ ;
	wire _w1883_ ;
	wire _w1884_ ;
	wire _w1885_ ;
	wire _w1886_ ;
	wire _w1887_ ;
	wire _w1888_ ;
	wire _w1889_ ;
	wire _w1890_ ;
	wire _w1891_ ;
	wire _w1892_ ;
	wire _w1893_ ;
	wire _w1894_ ;
	wire _w1895_ ;
	wire _w1896_ ;
	wire _w1897_ ;
	wire _w1898_ ;
	wire _w1899_ ;
	wire _w1900_ ;
	wire _w1901_ ;
	wire _w1902_ ;
	wire _w1903_ ;
	wire _w1904_ ;
	wire _w1905_ ;
	wire _w1906_ ;
	wire _w1907_ ;
	wire _w1908_ ;
	wire _w1909_ ;
	wire _w1910_ ;
	wire _w1911_ ;
	wire _w1912_ ;
	wire _w1913_ ;
	wire _w1914_ ;
	wire _w1915_ ;
	wire _w1916_ ;
	wire _w1917_ ;
	wire _w1918_ ;
	wire _w1919_ ;
	wire _w1920_ ;
	wire _w1921_ ;
	wire _w1922_ ;
	wire _w1923_ ;
	wire _w1924_ ;
	wire _w1925_ ;
	wire _w1926_ ;
	wire _w1927_ ;
	wire _w1928_ ;
	wire _w1929_ ;
	wire _w1930_ ;
	wire _w1931_ ;
	wire _w1932_ ;
	wire _w1933_ ;
	wire _w1934_ ;
	wire _w1935_ ;
	wire _w1936_ ;
	wire _w1937_ ;
	wire _w1938_ ;
	wire _w1939_ ;
	wire _w1940_ ;
	wire _w1941_ ;
	wire _w1942_ ;
	wire _w1943_ ;
	wire _w1944_ ;
	wire _w1945_ ;
	wire _w1946_ ;
	wire _w1947_ ;
	wire _w1948_ ;
	wire _w1949_ ;
	wire _w1950_ ;
	wire _w1951_ ;
	wire _w1952_ ;
	wire _w1953_ ;
	wire _w1954_ ;
	wire _w1955_ ;
	wire _w1956_ ;
	wire _w1957_ ;
	wire _w1958_ ;
	wire _w1959_ ;
	wire _w1960_ ;
	wire _w1961_ ;
	wire _w1962_ ;
	wire _w1963_ ;
	wire _w1964_ ;
	wire _w1965_ ;
	wire _w1966_ ;
	wire _w1967_ ;
	wire _w1968_ ;
	wire _w1969_ ;
	wire _w1970_ ;
	wire _w1971_ ;
	wire _w1972_ ;
	wire _w1973_ ;
	wire _w1974_ ;
	wire _w1975_ ;
	wire _w1976_ ;
	wire _w1977_ ;
	wire _w1978_ ;
	wire _w1979_ ;
	wire _w1980_ ;
	wire _w1981_ ;
	wire _w1982_ ;
	wire _w1983_ ;
	wire _w1984_ ;
	wire _w1985_ ;
	wire _w1986_ ;
	wire _w1987_ ;
	wire _w1988_ ;
	wire _w1989_ ;
	wire _w1990_ ;
	wire _w1991_ ;
	wire _w1992_ ;
	wire _w1993_ ;
	wire _w1994_ ;
	wire _w1995_ ;
	wire _w1996_ ;
	wire _w1997_ ;
	wire _w1998_ ;
	wire _w1999_ ;
	wire _w2000_ ;
	wire _w2001_ ;
	wire _w2002_ ;
	wire _w2003_ ;
	wire _w2004_ ;
	wire _w2005_ ;
	wire _w2006_ ;
	wire _w2007_ ;
	wire _w2008_ ;
	wire _w2009_ ;
	wire _w2010_ ;
	wire _w2011_ ;
	wire _w2012_ ;
	wire _w2013_ ;
	wire _w2014_ ;
	wire _w2015_ ;
	wire _w2016_ ;
	wire _w2017_ ;
	wire _w2018_ ;
	wire _w2019_ ;
	wire _w2020_ ;
	wire _w2021_ ;
	wire _w2022_ ;
	wire _w2023_ ;
	wire _w2024_ ;
	wire _w2025_ ;
	wire _w2026_ ;
	wire _w2027_ ;
	wire _w2028_ ;
	wire _w2029_ ;
	wire _w2030_ ;
	wire _w2031_ ;
	wire _w2032_ ;
	wire _w2033_ ;
	wire _w2034_ ;
	wire _w2035_ ;
	wire _w2036_ ;
	wire _w2037_ ;
	wire _w2038_ ;
	wire _w2039_ ;
	wire _w2040_ ;
	wire _w2041_ ;
	wire _w2042_ ;
	wire _w2043_ ;
	wire _w2044_ ;
	wire _w2045_ ;
	wire _w2046_ ;
	wire _w2047_ ;
	wire _w2048_ ;
	wire _w2049_ ;
	wire _w2050_ ;
	wire _w2051_ ;
	wire _w2052_ ;
	wire _w2053_ ;
	wire _w2054_ ;
	wire _w2055_ ;
	wire _w2056_ ;
	wire _w2057_ ;
	wire _w2058_ ;
	wire _w2059_ ;
	wire _w2060_ ;
	wire _w2061_ ;
	wire _w2062_ ;
	wire _w2063_ ;
	wire _w2064_ ;
	wire _w2065_ ;
	wire _w2066_ ;
	wire _w2067_ ;
	wire _w2068_ ;
	wire _w2069_ ;
	wire _w2070_ ;
	wire _w2071_ ;
	wire _w2072_ ;
	wire _w2073_ ;
	wire _w2074_ ;
	wire _w2075_ ;
	wire _w2076_ ;
	wire _w2077_ ;
	wire _w2078_ ;
	wire _w2079_ ;
	wire _w2080_ ;
	wire _w2081_ ;
	wire _w2082_ ;
	wire _w2083_ ;
	wire _w2084_ ;
	wire _w2085_ ;
	wire _w2086_ ;
	wire _w2087_ ;
	wire _w2088_ ;
	wire _w2089_ ;
	wire _w2090_ ;
	wire _w2091_ ;
	wire _w2092_ ;
	wire _w2093_ ;
	wire _w2094_ ;
	wire _w2095_ ;
	wire _w2096_ ;
	wire _w2097_ ;
	wire _w2098_ ;
	wire _w2099_ ;
	wire _w2100_ ;
	wire _w2101_ ;
	wire _w2102_ ;
	wire _w2103_ ;
	wire _w2104_ ;
	wire _w2105_ ;
	wire _w2106_ ;
	wire _w2107_ ;
	wire _w2108_ ;
	wire _w2109_ ;
	wire _w2110_ ;
	wire _w2111_ ;
	wire _w2112_ ;
	wire _w2113_ ;
	wire _w2114_ ;
	wire _w2115_ ;
	wire _w2116_ ;
	wire _w2117_ ;
	wire _w2118_ ;
	wire _w2119_ ;
	wire _w2120_ ;
	wire _w2121_ ;
	wire _w2122_ ;
	wire _w2123_ ;
	wire _w2124_ ;
	wire _w2125_ ;
	wire _w2126_ ;
	wire _w2127_ ;
	wire _w2128_ ;
	wire _w2129_ ;
	wire _w2130_ ;
	wire _w2131_ ;
	wire _w2132_ ;
	wire _w2133_ ;
	wire _w2134_ ;
	wire _w2135_ ;
	wire _w2136_ ;
	wire _w2137_ ;
	wire _w2138_ ;
	wire _w2139_ ;
	wire _w2140_ ;
	wire _w2141_ ;
	wire _w2142_ ;
	wire _w2143_ ;
	wire _w2144_ ;
	wire _w2145_ ;
	wire _w2146_ ;
	wire _w2147_ ;
	wire _w2148_ ;
	wire _w2149_ ;
	wire _w2150_ ;
	wire _w2151_ ;
	wire _w2152_ ;
	wire _w2153_ ;
	wire _w2154_ ;
	wire _w2155_ ;
	wire _w2156_ ;
	wire _w2157_ ;
	wire _w2158_ ;
	wire _w2159_ ;
	wire _w2160_ ;
	wire _w2161_ ;
	wire _w2162_ ;
	wire _w2163_ ;
	wire _w2164_ ;
	wire _w2165_ ;
	wire _w2166_ ;
	wire _w2167_ ;
	wire _w2168_ ;
	wire _w2169_ ;
	wire _w2170_ ;
	wire _w2171_ ;
	wire _w2172_ ;
	wire _w2173_ ;
	wire _w2174_ ;
	wire _w2175_ ;
	wire _w2176_ ;
	wire _w2177_ ;
	wire _w2178_ ;
	wire _w2179_ ;
	wire _w2180_ ;
	wire _w2181_ ;
	wire _w2182_ ;
	wire _w2183_ ;
	wire _w2184_ ;
	wire _w2185_ ;
	wire _w2186_ ;
	wire _w2187_ ;
	wire _w2188_ ;
	wire _w2189_ ;
	wire _w2190_ ;
	wire _w2191_ ;
	wire _w2192_ ;
	wire _w2193_ ;
	wire _w2194_ ;
	wire _w2195_ ;
	wire _w2196_ ;
	wire _w2197_ ;
	wire _w2198_ ;
	wire _w2199_ ;
	wire _w2200_ ;
	wire _w2201_ ;
	wire _w2202_ ;
	wire _w2203_ ;
	wire _w2204_ ;
	wire _w2205_ ;
	wire _w2206_ ;
	wire _w2207_ ;
	wire _w2208_ ;
	wire _w2209_ ;
	wire _w2210_ ;
	wire _w2211_ ;
	wire _w2212_ ;
	wire _w2213_ ;
	wire _w2214_ ;
	wire _w2215_ ;
	wire _w2216_ ;
	wire _w2217_ ;
	wire _w2218_ ;
	wire _w2219_ ;
	wire _w2220_ ;
	wire _w2221_ ;
	wire _w2222_ ;
	wire _w2223_ ;
	wire _w2224_ ;
	wire _w2225_ ;
	wire _w2226_ ;
	wire _w2227_ ;
	wire _w2228_ ;
	wire _w2229_ ;
	wire _w2230_ ;
	wire _w2231_ ;
	wire _w2232_ ;
	wire _w2233_ ;
	wire _w2234_ ;
	wire _w2235_ ;
	wire _w2236_ ;
	wire _w2237_ ;
	wire _w2238_ ;
	wire _w2239_ ;
	wire _w2240_ ;
	wire _w2241_ ;
	wire _w2242_ ;
	wire _w2243_ ;
	wire _w2244_ ;
	wire _w2245_ ;
	wire _w2246_ ;
	wire _w2247_ ;
	wire _w2248_ ;
	wire _w2249_ ;
	wire _w2250_ ;
	wire _w2251_ ;
	wire _w2252_ ;
	wire _w2253_ ;
	wire _w2254_ ;
	wire _w2255_ ;
	wire _w2256_ ;
	wire _w2257_ ;
	wire _w2258_ ;
	wire _w2259_ ;
	wire _w2260_ ;
	wire _w2261_ ;
	wire _w2262_ ;
	wire _w2263_ ;
	wire _w2264_ ;
	wire _w2265_ ;
	wire _w2266_ ;
	wire _w2267_ ;
	wire _w2268_ ;
	wire _w2269_ ;
	wire _w2270_ ;
	wire _w2271_ ;
	wire _w2272_ ;
	wire _w2273_ ;
	wire _w2274_ ;
	wire _w2275_ ;
	wire _w2276_ ;
	wire _w2277_ ;
	wire _w2278_ ;
	wire _w2279_ ;
	wire _w2280_ ;
	wire _w2281_ ;
	wire _w2282_ ;
	wire _w2283_ ;
	wire _w2284_ ;
	wire _w2285_ ;
	wire _w2286_ ;
	wire _w2287_ ;
	wire _w2288_ ;
	wire _w2289_ ;
	wire _w2290_ ;
	wire _w2291_ ;
	wire _w2292_ ;
	wire _w2293_ ;
	wire _w2294_ ;
	wire _w2295_ ;
	wire _w2296_ ;
	wire _w2297_ ;
	wire _w2298_ ;
	wire _w2299_ ;
	wire _w2300_ ;
	wire _w2301_ ;
	wire _w2302_ ;
	wire _w2303_ ;
	wire _w2304_ ;
	wire _w2305_ ;
	wire _w2306_ ;
	wire _w2307_ ;
	wire _w2308_ ;
	wire _w2309_ ;
	wire _w2310_ ;
	wire _w2311_ ;
	wire _w2312_ ;
	wire _w2313_ ;
	wire _w2314_ ;
	wire _w2315_ ;
	wire _w2316_ ;
	wire _w2317_ ;
	wire _w2318_ ;
	wire _w2319_ ;
	wire _w2320_ ;
	wire _w2321_ ;
	wire _w2322_ ;
	wire _w2323_ ;
	wire _w2324_ ;
	wire _w2325_ ;
	wire _w2326_ ;
	wire _w2327_ ;
	wire _w2328_ ;
	wire _w2329_ ;
	wire _w2330_ ;
	wire _w2331_ ;
	wire _w2332_ ;
	wire _w2333_ ;
	wire _w2334_ ;
	wire _w2335_ ;
	wire _w2336_ ;
	wire _w2337_ ;
	wire _w2338_ ;
	wire _w2339_ ;
	wire _w2340_ ;
	wire _w2341_ ;
	wire _w2342_ ;
	wire _w2343_ ;
	wire _w2344_ ;
	wire _w2345_ ;
	wire _w2346_ ;
	wire _w2347_ ;
	wire _w2348_ ;
	wire _w2349_ ;
	wire _w2350_ ;
	wire _w2351_ ;
	wire _w2352_ ;
	wire _w2353_ ;
	wire _w2354_ ;
	wire _w2355_ ;
	wire _w2356_ ;
	wire _w2357_ ;
	wire _w2358_ ;
	wire _w2359_ ;
	wire _w2360_ ;
	wire _w2361_ ;
	wire _w2362_ ;
	wire _w2363_ ;
	wire _w2364_ ;
	wire _w2365_ ;
	wire _w2366_ ;
	wire _w2367_ ;
	wire _w2368_ ;
	wire _w2369_ ;
	wire _w2370_ ;
	wire _w2371_ ;
	wire _w2372_ ;
	wire _w2373_ ;
	wire _w2374_ ;
	wire _w2375_ ;
	wire _w2376_ ;
	wire _w2377_ ;
	wire _w2378_ ;
	wire _w2379_ ;
	wire _w2380_ ;
	wire _w2381_ ;
	wire _w2382_ ;
	wire _w2383_ ;
	wire _w2384_ ;
	wire _w2385_ ;
	wire _w2386_ ;
	wire _w2387_ ;
	wire _w2388_ ;
	wire _w2389_ ;
	wire _w2390_ ;
	wire _w2391_ ;
	wire _w2392_ ;
	wire _w2393_ ;
	wire _w2394_ ;
	wire _w2395_ ;
	wire _w2396_ ;
	wire _w2397_ ;
	wire _w2398_ ;
	wire _w2399_ ;
	wire _w2400_ ;
	wire _w2401_ ;
	wire _w2402_ ;
	wire _w2403_ ;
	wire _w2404_ ;
	wire _w2405_ ;
	wire _w2406_ ;
	wire _w2407_ ;
	wire _w2408_ ;
	wire _w2409_ ;
	wire _w2410_ ;
	wire _w2411_ ;
	wire _w2412_ ;
	wire _w2413_ ;
	wire _w2414_ ;
	wire _w2415_ ;
	wire _w2416_ ;
	wire _w2417_ ;
	wire _w2418_ ;
	wire _w2419_ ;
	wire _w2420_ ;
	wire _w2421_ ;
	wire _w2422_ ;
	wire _w2423_ ;
	wire _w2424_ ;
	wire _w2425_ ;
	wire _w2426_ ;
	wire _w2427_ ;
	wire _w2428_ ;
	wire _w2429_ ;
	wire _w2430_ ;
	wire _w2431_ ;
	wire _w2432_ ;
	wire _w2433_ ;
	wire _w2434_ ;
	wire _w2435_ ;
	wire _w2436_ ;
	wire _w2437_ ;
	wire _w2438_ ;
	wire _w2439_ ;
	wire _w2440_ ;
	wire _w2441_ ;
	wire _w2442_ ;
	wire _w2443_ ;
	wire _w2444_ ;
	wire _w2445_ ;
	wire _w2446_ ;
	wire _w2447_ ;
	wire _w2448_ ;
	wire _w2449_ ;
	wire _w2450_ ;
	wire _w2451_ ;
	wire _w2452_ ;
	wire _w2453_ ;
	wire _w2454_ ;
	wire _w2455_ ;
	wire _w2456_ ;
	wire _w2457_ ;
	wire _w2458_ ;
	wire _w2459_ ;
	wire _w2460_ ;
	wire _w2461_ ;
	wire _w2462_ ;
	wire _w2463_ ;
	wire _w2464_ ;
	wire _w2465_ ;
	wire _w2466_ ;
	wire _w2467_ ;
	wire _w2468_ ;
	wire _w2469_ ;
	wire _w2470_ ;
	wire _w2471_ ;
	wire _w2472_ ;
	wire _w2473_ ;
	wire _w2474_ ;
	wire _w2475_ ;
	wire _w2476_ ;
	wire _w2477_ ;
	wire _w2478_ ;
	wire _w2479_ ;
	wire _w2480_ ;
	wire _w2481_ ;
	wire _w2482_ ;
	wire _w2483_ ;
	wire _w2484_ ;
	wire _w2485_ ;
	wire _w2486_ ;
	wire _w2487_ ;
	wire _w2488_ ;
	wire _w2489_ ;
	wire _w2490_ ;
	wire _w2491_ ;
	wire _w2492_ ;
	wire _w2493_ ;
	wire _w2494_ ;
	wire _w2495_ ;
	wire _w2496_ ;
	wire _w2497_ ;
	wire _w2498_ ;
	wire _w2499_ ;
	wire _w2500_ ;
	wire _w2501_ ;
	wire _w2502_ ;
	wire _w2503_ ;
	wire _w2504_ ;
	wire _w2505_ ;
	wire _w2506_ ;
	wire _w2507_ ;
	wire _w2508_ ;
	wire _w2509_ ;
	wire _w2510_ ;
	wire _w2511_ ;
	wire _w2512_ ;
	wire _w2513_ ;
	wire _w2514_ ;
	wire _w2515_ ;
	wire _w2516_ ;
	wire _w2517_ ;
	wire _w2518_ ;
	wire _w2519_ ;
	wire _w2520_ ;
	wire _w2521_ ;
	wire _w2522_ ;
	wire _w2523_ ;
	wire _w2524_ ;
	wire _w2525_ ;
	wire _w2526_ ;
	wire _w2527_ ;
	wire _w2528_ ;
	wire _w2529_ ;
	wire _w2530_ ;
	wire _w2531_ ;
	wire _w2532_ ;
	wire _w2533_ ;
	wire _w2534_ ;
	wire _w2535_ ;
	wire _w2536_ ;
	wire _w2537_ ;
	wire _w2538_ ;
	wire _w2539_ ;
	wire _w2540_ ;
	wire _w2541_ ;
	wire _w2542_ ;
	wire _w2543_ ;
	wire _w2544_ ;
	wire _w2545_ ;
	wire _w2546_ ;
	wire _w2547_ ;
	wire _w2548_ ;
	wire _w2549_ ;
	wire _w2550_ ;
	wire _w2551_ ;
	wire _w2552_ ;
	wire _w2553_ ;
	wire _w2554_ ;
	wire _w2555_ ;
	wire _w2556_ ;
	wire _w2557_ ;
	wire _w2558_ ;
	wire _w2559_ ;
	wire _w2560_ ;
	wire _w2561_ ;
	wire _w2562_ ;
	wire _w2563_ ;
	wire _w2564_ ;
	wire _w2565_ ;
	wire _w2566_ ;
	wire _w2567_ ;
	wire _w2568_ ;
	wire _w2569_ ;
	wire _w2570_ ;
	wire _w2571_ ;
	wire _w2572_ ;
	wire _w2573_ ;
	wire _w2574_ ;
	wire _w2575_ ;
	wire _w2576_ ;
	wire _w2577_ ;
	wire _w2578_ ;
	wire _w2579_ ;
	wire _w2580_ ;
	wire _w2581_ ;
	wire _w2582_ ;
	wire _w2583_ ;
	wire _w2584_ ;
	wire _w2585_ ;
	wire _w2586_ ;
	wire _w2587_ ;
	wire _w2588_ ;
	wire _w2589_ ;
	wire _w2590_ ;
	wire _w2591_ ;
	wire _w2592_ ;
	wire _w2593_ ;
	wire _w2594_ ;
	wire _w2595_ ;
	wire _w2596_ ;
	wire _w2597_ ;
	wire _w2598_ ;
	wire _w2599_ ;
	wire _w2600_ ;
	wire _w2601_ ;
	wire _w2602_ ;
	wire _w2603_ ;
	wire _w2604_ ;
	wire _w2605_ ;
	wire _w2606_ ;
	wire _w2607_ ;
	wire _w2608_ ;
	wire _w2609_ ;
	wire _w2610_ ;
	wire _w2611_ ;
	wire _w2612_ ;
	wire _w2613_ ;
	wire _w2614_ ;
	LUT4 #(
		.INIT('h0501)
	) name0 (
		\priority[0] ,
		\priority[126] ,
		\priority[127] ,
		\req[126] ,
		_w258_
	);
	LUT3 #(
		.INIT('h8c)
	) name1 (
		\priority[0] ,
		\req[0] ,
		\req[127] ,
		_w259_
	);
	LUT2 #(
		.INIT('h4)
	) name2 (
		_w258_,
		_w259_,
		_w260_
	);
	LUT3 #(
		.INIT('h31)
	) name3 (
		\priority[1] ,
		\priority[2] ,
		\req[1] ,
		_w261_
	);
	LUT2 #(
		.INIT('h1)
	) name4 (
		\req[2] ,
		\req[3] ,
		_w262_
	);
	LUT4 #(
		.INIT('h0301)
	) name5 (
		\priority[6] ,
		\priority[7] ,
		\priority[8] ,
		\req[6] ,
		_w263_
	);
	LUT4 #(
		.INIT('h0301)
	) name6 (
		\priority[3] ,
		\priority[4] ,
		\priority[5] ,
		\req[3] ,
		_w264_
	);
	LUT4 #(
		.INIT('hb000)
	) name7 (
		_w261_,
		_w262_,
		_w263_,
		_w264_,
		_w265_
	);
	LUT2 #(
		.INIT('h1)
	) name8 (
		\req[5] ,
		\req[6] ,
		_w266_
	);
	LUT4 #(
		.INIT('h000b)
	) name9 (
		\priority[5] ,
		\req[4] ,
		\req[5] ,
		\req[6] ,
		_w267_
	);
	LUT2 #(
		.INIT('h1)
	) name10 (
		\req[11] ,
		\req[12] ,
		_w268_
	);
	LUT4 #(
		.INIT('h000b)
	) name11 (
		\priority[11] ,
		\req[10] ,
		\req[11] ,
		\req[12] ,
		_w269_
	);
	LUT2 #(
		.INIT('h1)
	) name12 (
		\req[8] ,
		\req[9] ,
		_w270_
	);
	LUT4 #(
		.INIT('h000b)
	) name13 (
		\priority[8] ,
		\req[7] ,
		\req[8] ,
		\req[9] ,
		_w271_
	);
	LUT4 #(
		.INIT('hd000)
	) name14 (
		_w263_,
		_w267_,
		_w269_,
		_w271_,
		_w272_
	);
	LUT4 #(
		.INIT('h0301)
	) name15 (
		\priority[9] ,
		\priority[10] ,
		\priority[11] ,
		\req[9] ,
		_w273_
	);
	LUT4 #(
		.INIT('h0301)
	) name16 (
		\priority[15] ,
		\priority[16] ,
		\priority[17] ,
		\req[15] ,
		_w274_
	);
	LUT4 #(
		.INIT('h0301)
	) name17 (
		\priority[12] ,
		\priority[13] ,
		\priority[14] ,
		\req[12] ,
		_w275_
	);
	LUT4 #(
		.INIT('hd000)
	) name18 (
		_w269_,
		_w273_,
		_w274_,
		_w275_,
		_w276_
	);
	LUT2 #(
		.INIT('h1)
	) name19 (
		\req[14] ,
		\req[15] ,
		_w277_
	);
	LUT4 #(
		.INIT('h000b)
	) name20 (
		\priority[14] ,
		\req[13] ,
		\req[14] ,
		\req[15] ,
		_w278_
	);
	LUT2 #(
		.INIT('h1)
	) name21 (
		\req[20] ,
		\req[21] ,
		_w279_
	);
	LUT4 #(
		.INIT('h000b)
	) name22 (
		\priority[20] ,
		\req[19] ,
		\req[20] ,
		\req[21] ,
		_w280_
	);
	LUT2 #(
		.INIT('h1)
	) name23 (
		\req[17] ,
		\req[18] ,
		_w281_
	);
	LUT4 #(
		.INIT('h000b)
	) name24 (
		\priority[17] ,
		\req[16] ,
		\req[17] ,
		\req[18] ,
		_w282_
	);
	LUT4 #(
		.INIT('hd000)
	) name25 (
		_w274_,
		_w278_,
		_w280_,
		_w282_,
		_w283_
	);
	LUT4 #(
		.INIT('h4f00)
	) name26 (
		_w265_,
		_w272_,
		_w276_,
		_w283_,
		_w284_
	);
	LUT4 #(
		.INIT('h0301)
	) name27 (
		\priority[18] ,
		\priority[19] ,
		\priority[20] ,
		\req[18] ,
		_w285_
	);
	LUT4 #(
		.INIT('h0301)
	) name28 (
		\priority[24] ,
		\priority[25] ,
		\priority[26] ,
		\req[24] ,
		_w286_
	);
	LUT4 #(
		.INIT('h0301)
	) name29 (
		\priority[21] ,
		\priority[22] ,
		\priority[23] ,
		\req[21] ,
		_w287_
	);
	LUT4 #(
		.INIT('hd000)
	) name30 (
		_w280_,
		_w285_,
		_w286_,
		_w287_,
		_w288_
	);
	LUT2 #(
		.INIT('h1)
	) name31 (
		\req[23] ,
		\req[24] ,
		_w289_
	);
	LUT4 #(
		.INIT('h000b)
	) name32 (
		\priority[23] ,
		\req[22] ,
		\req[23] ,
		\req[24] ,
		_w290_
	);
	LUT2 #(
		.INIT('h1)
	) name33 (
		\req[29] ,
		\req[30] ,
		_w291_
	);
	LUT4 #(
		.INIT('h000b)
	) name34 (
		\priority[29] ,
		\req[28] ,
		\req[29] ,
		\req[30] ,
		_w292_
	);
	LUT2 #(
		.INIT('h1)
	) name35 (
		\req[26] ,
		\req[27] ,
		_w293_
	);
	LUT4 #(
		.INIT('h000b)
	) name36 (
		\priority[26] ,
		\req[25] ,
		\req[26] ,
		\req[27] ,
		_w294_
	);
	LUT4 #(
		.INIT('hd000)
	) name37 (
		_w286_,
		_w290_,
		_w292_,
		_w294_,
		_w295_
	);
	LUT4 #(
		.INIT('h0301)
	) name38 (
		\priority[27] ,
		\priority[28] ,
		\priority[29] ,
		\req[27] ,
		_w296_
	);
	LUT4 #(
		.INIT('h0301)
	) name39 (
		\priority[33] ,
		\priority[34] ,
		\priority[35] ,
		\req[33] ,
		_w297_
	);
	LUT4 #(
		.INIT('h0301)
	) name40 (
		\priority[30] ,
		\priority[31] ,
		\priority[32] ,
		\req[30] ,
		_w298_
	);
	LUT4 #(
		.INIT('hd000)
	) name41 (
		_w292_,
		_w296_,
		_w297_,
		_w298_,
		_w299_
	);
	LUT4 #(
		.INIT('h4f00)
	) name42 (
		_w284_,
		_w288_,
		_w295_,
		_w299_,
		_w300_
	);
	LUT2 #(
		.INIT('h1)
	) name43 (
		\req[32] ,
		\req[33] ,
		_w301_
	);
	LUT4 #(
		.INIT('h000b)
	) name44 (
		\priority[32] ,
		\req[31] ,
		\req[32] ,
		\req[33] ,
		_w302_
	);
	LUT2 #(
		.INIT('h1)
	) name45 (
		\req[38] ,
		\req[39] ,
		_w303_
	);
	LUT4 #(
		.INIT('h000b)
	) name46 (
		\priority[38] ,
		\req[37] ,
		\req[38] ,
		\req[39] ,
		_w304_
	);
	LUT2 #(
		.INIT('h1)
	) name47 (
		\req[35] ,
		\req[36] ,
		_w305_
	);
	LUT4 #(
		.INIT('h000b)
	) name48 (
		\priority[35] ,
		\req[34] ,
		\req[35] ,
		\req[36] ,
		_w306_
	);
	LUT4 #(
		.INIT('hd000)
	) name49 (
		_w297_,
		_w302_,
		_w304_,
		_w306_,
		_w307_
	);
	LUT4 #(
		.INIT('h0301)
	) name50 (
		\priority[36] ,
		\priority[37] ,
		\priority[38] ,
		\req[36] ,
		_w308_
	);
	LUT4 #(
		.INIT('h0301)
	) name51 (
		\priority[42] ,
		\priority[43] ,
		\priority[44] ,
		\req[42] ,
		_w309_
	);
	LUT4 #(
		.INIT('h0301)
	) name52 (
		\priority[39] ,
		\priority[40] ,
		\priority[41] ,
		\req[39] ,
		_w310_
	);
	LUT4 #(
		.INIT('hd000)
	) name53 (
		_w304_,
		_w308_,
		_w309_,
		_w310_,
		_w311_
	);
	LUT2 #(
		.INIT('h1)
	) name54 (
		\req[41] ,
		\req[42] ,
		_w312_
	);
	LUT4 #(
		.INIT('h000b)
	) name55 (
		\priority[41] ,
		\req[40] ,
		\req[41] ,
		\req[42] ,
		_w313_
	);
	LUT2 #(
		.INIT('h1)
	) name56 (
		\req[47] ,
		\req[48] ,
		_w314_
	);
	LUT4 #(
		.INIT('h000b)
	) name57 (
		\priority[47] ,
		\req[46] ,
		\req[47] ,
		\req[48] ,
		_w315_
	);
	LUT2 #(
		.INIT('h1)
	) name58 (
		\req[44] ,
		\req[45] ,
		_w316_
	);
	LUT4 #(
		.INIT('h000b)
	) name59 (
		\priority[44] ,
		\req[43] ,
		\req[44] ,
		\req[45] ,
		_w317_
	);
	LUT4 #(
		.INIT('hd000)
	) name60 (
		_w309_,
		_w313_,
		_w315_,
		_w317_,
		_w318_
	);
	LUT4 #(
		.INIT('h4f00)
	) name61 (
		_w300_,
		_w307_,
		_w311_,
		_w318_,
		_w319_
	);
	LUT4 #(
		.INIT('h0301)
	) name62 (
		\priority[45] ,
		\priority[46] ,
		\priority[47] ,
		\req[45] ,
		_w320_
	);
	LUT4 #(
		.INIT('h0301)
	) name63 (
		\priority[51] ,
		\priority[52] ,
		\priority[53] ,
		\req[51] ,
		_w321_
	);
	LUT4 #(
		.INIT('h0301)
	) name64 (
		\priority[48] ,
		\priority[49] ,
		\priority[50] ,
		\req[48] ,
		_w322_
	);
	LUT4 #(
		.INIT('hd000)
	) name65 (
		_w315_,
		_w320_,
		_w321_,
		_w322_,
		_w323_
	);
	LUT2 #(
		.INIT('h1)
	) name66 (
		\req[50] ,
		\req[51] ,
		_w324_
	);
	LUT4 #(
		.INIT('h000b)
	) name67 (
		\priority[50] ,
		\req[49] ,
		\req[50] ,
		\req[51] ,
		_w325_
	);
	LUT2 #(
		.INIT('h1)
	) name68 (
		\req[56] ,
		\req[57] ,
		_w326_
	);
	LUT4 #(
		.INIT('h000b)
	) name69 (
		\priority[56] ,
		\req[55] ,
		\req[56] ,
		\req[57] ,
		_w327_
	);
	LUT2 #(
		.INIT('h1)
	) name70 (
		\req[53] ,
		\req[54] ,
		_w328_
	);
	LUT4 #(
		.INIT('h000b)
	) name71 (
		\priority[53] ,
		\req[52] ,
		\req[53] ,
		\req[54] ,
		_w329_
	);
	LUT4 #(
		.INIT('hd000)
	) name72 (
		_w321_,
		_w325_,
		_w327_,
		_w329_,
		_w330_
	);
	LUT4 #(
		.INIT('h0301)
	) name73 (
		\priority[54] ,
		\priority[55] ,
		\priority[56] ,
		\req[54] ,
		_w331_
	);
	LUT4 #(
		.INIT('h0301)
	) name74 (
		\priority[60] ,
		\priority[61] ,
		\priority[62] ,
		\req[60] ,
		_w332_
	);
	LUT4 #(
		.INIT('h0301)
	) name75 (
		\priority[57] ,
		\priority[58] ,
		\priority[59] ,
		\req[57] ,
		_w333_
	);
	LUT4 #(
		.INIT('hd000)
	) name76 (
		_w327_,
		_w331_,
		_w332_,
		_w333_,
		_w334_
	);
	LUT4 #(
		.INIT('h4f00)
	) name77 (
		_w319_,
		_w323_,
		_w330_,
		_w334_,
		_w335_
	);
	LUT2 #(
		.INIT('h1)
	) name78 (
		\req[59] ,
		\req[60] ,
		_w336_
	);
	LUT4 #(
		.INIT('h000b)
	) name79 (
		\priority[59] ,
		\req[58] ,
		\req[59] ,
		\req[60] ,
		_w337_
	);
	LUT2 #(
		.INIT('h1)
	) name80 (
		\req[65] ,
		\req[66] ,
		_w338_
	);
	LUT4 #(
		.INIT('h000b)
	) name81 (
		\priority[65] ,
		\req[64] ,
		\req[65] ,
		\req[66] ,
		_w339_
	);
	LUT2 #(
		.INIT('h1)
	) name82 (
		\req[62] ,
		\req[63] ,
		_w340_
	);
	LUT4 #(
		.INIT('h000b)
	) name83 (
		\priority[62] ,
		\req[61] ,
		\req[62] ,
		\req[63] ,
		_w341_
	);
	LUT4 #(
		.INIT('hd000)
	) name84 (
		_w332_,
		_w337_,
		_w339_,
		_w341_,
		_w342_
	);
	LUT4 #(
		.INIT('h0301)
	) name85 (
		\priority[63] ,
		\priority[64] ,
		\priority[65] ,
		\req[63] ,
		_w343_
	);
	LUT4 #(
		.INIT('h0301)
	) name86 (
		\priority[69] ,
		\priority[70] ,
		\priority[71] ,
		\req[69] ,
		_w344_
	);
	LUT4 #(
		.INIT('h0301)
	) name87 (
		\priority[66] ,
		\priority[67] ,
		\priority[68] ,
		\req[66] ,
		_w345_
	);
	LUT4 #(
		.INIT('hd000)
	) name88 (
		_w339_,
		_w343_,
		_w344_,
		_w345_,
		_w346_
	);
	LUT2 #(
		.INIT('h1)
	) name89 (
		\req[68] ,
		\req[69] ,
		_w347_
	);
	LUT4 #(
		.INIT('h000b)
	) name90 (
		\priority[68] ,
		\req[67] ,
		\req[68] ,
		\req[69] ,
		_w348_
	);
	LUT2 #(
		.INIT('h1)
	) name91 (
		\req[74] ,
		\req[75] ,
		_w349_
	);
	LUT4 #(
		.INIT('h000b)
	) name92 (
		\priority[74] ,
		\req[73] ,
		\req[74] ,
		\req[75] ,
		_w350_
	);
	LUT2 #(
		.INIT('h1)
	) name93 (
		\req[71] ,
		\req[72] ,
		_w351_
	);
	LUT4 #(
		.INIT('h000b)
	) name94 (
		\priority[71] ,
		\req[70] ,
		\req[71] ,
		\req[72] ,
		_w352_
	);
	LUT4 #(
		.INIT('hd000)
	) name95 (
		_w344_,
		_w348_,
		_w350_,
		_w352_,
		_w353_
	);
	LUT4 #(
		.INIT('h4f00)
	) name96 (
		_w335_,
		_w342_,
		_w346_,
		_w353_,
		_w354_
	);
	LUT4 #(
		.INIT('h0301)
	) name97 (
		\priority[72] ,
		\priority[73] ,
		\priority[74] ,
		\req[72] ,
		_w355_
	);
	LUT4 #(
		.INIT('h0301)
	) name98 (
		\priority[78] ,
		\priority[79] ,
		\priority[80] ,
		\req[78] ,
		_w356_
	);
	LUT4 #(
		.INIT('h0301)
	) name99 (
		\priority[75] ,
		\priority[76] ,
		\priority[77] ,
		\req[75] ,
		_w357_
	);
	LUT4 #(
		.INIT('hd000)
	) name100 (
		_w350_,
		_w355_,
		_w356_,
		_w357_,
		_w358_
	);
	LUT2 #(
		.INIT('h1)
	) name101 (
		\req[77] ,
		\req[78] ,
		_w359_
	);
	LUT4 #(
		.INIT('h000b)
	) name102 (
		\priority[77] ,
		\req[76] ,
		\req[77] ,
		\req[78] ,
		_w360_
	);
	LUT2 #(
		.INIT('h1)
	) name103 (
		\req[83] ,
		\req[84] ,
		_w361_
	);
	LUT4 #(
		.INIT('h000b)
	) name104 (
		\priority[83] ,
		\req[82] ,
		\req[83] ,
		\req[84] ,
		_w362_
	);
	LUT2 #(
		.INIT('h1)
	) name105 (
		\req[80] ,
		\req[81] ,
		_w363_
	);
	LUT4 #(
		.INIT('h000b)
	) name106 (
		\priority[80] ,
		\req[79] ,
		\req[80] ,
		\req[81] ,
		_w364_
	);
	LUT4 #(
		.INIT('hd000)
	) name107 (
		_w356_,
		_w360_,
		_w362_,
		_w364_,
		_w365_
	);
	LUT4 #(
		.INIT('h0301)
	) name108 (
		\priority[81] ,
		\priority[82] ,
		\priority[83] ,
		\req[81] ,
		_w366_
	);
	LUT4 #(
		.INIT('h0301)
	) name109 (
		\priority[87] ,
		\priority[88] ,
		\priority[89] ,
		\req[87] ,
		_w367_
	);
	LUT4 #(
		.INIT('h0301)
	) name110 (
		\priority[84] ,
		\priority[85] ,
		\priority[86] ,
		\req[84] ,
		_w368_
	);
	LUT4 #(
		.INIT('hd000)
	) name111 (
		_w362_,
		_w366_,
		_w367_,
		_w368_,
		_w369_
	);
	LUT4 #(
		.INIT('h4f00)
	) name112 (
		_w354_,
		_w358_,
		_w365_,
		_w369_,
		_w370_
	);
	LUT2 #(
		.INIT('h1)
	) name113 (
		\req[86] ,
		\req[87] ,
		_w371_
	);
	LUT4 #(
		.INIT('h000b)
	) name114 (
		\priority[86] ,
		\req[85] ,
		\req[86] ,
		\req[87] ,
		_w372_
	);
	LUT2 #(
		.INIT('h1)
	) name115 (
		\req[92] ,
		\req[93] ,
		_w373_
	);
	LUT4 #(
		.INIT('h000b)
	) name116 (
		\priority[92] ,
		\req[91] ,
		\req[92] ,
		\req[93] ,
		_w374_
	);
	LUT2 #(
		.INIT('h1)
	) name117 (
		\req[89] ,
		\req[90] ,
		_w375_
	);
	LUT4 #(
		.INIT('h000b)
	) name118 (
		\priority[89] ,
		\req[88] ,
		\req[89] ,
		\req[90] ,
		_w376_
	);
	LUT4 #(
		.INIT('hd000)
	) name119 (
		_w367_,
		_w372_,
		_w374_,
		_w376_,
		_w377_
	);
	LUT4 #(
		.INIT('h0301)
	) name120 (
		\priority[90] ,
		\priority[91] ,
		\priority[92] ,
		\req[90] ,
		_w378_
	);
	LUT4 #(
		.INIT('h0301)
	) name121 (
		\priority[96] ,
		\priority[97] ,
		\priority[98] ,
		\req[96] ,
		_w379_
	);
	LUT4 #(
		.INIT('h0301)
	) name122 (
		\priority[93] ,
		\priority[94] ,
		\priority[95] ,
		\req[93] ,
		_w380_
	);
	LUT4 #(
		.INIT('hd000)
	) name123 (
		_w374_,
		_w378_,
		_w379_,
		_w380_,
		_w381_
	);
	LUT2 #(
		.INIT('h1)
	) name124 (
		\req[95] ,
		\req[96] ,
		_w382_
	);
	LUT4 #(
		.INIT('h000b)
	) name125 (
		\priority[95] ,
		\req[94] ,
		\req[95] ,
		\req[96] ,
		_w383_
	);
	LUT2 #(
		.INIT('h1)
	) name126 (
		\req[101] ,
		\req[102] ,
		_w384_
	);
	LUT4 #(
		.INIT('h000b)
	) name127 (
		\priority[101] ,
		\req[100] ,
		\req[101] ,
		\req[102] ,
		_w385_
	);
	LUT2 #(
		.INIT('h1)
	) name128 (
		\req[98] ,
		\req[99] ,
		_w386_
	);
	LUT4 #(
		.INIT('h000b)
	) name129 (
		\priority[98] ,
		\req[97] ,
		\req[98] ,
		\req[99] ,
		_w387_
	);
	LUT4 #(
		.INIT('hd000)
	) name130 (
		_w379_,
		_w383_,
		_w385_,
		_w387_,
		_w388_
	);
	LUT4 #(
		.INIT('h4f00)
	) name131 (
		_w370_,
		_w377_,
		_w381_,
		_w388_,
		_w389_
	);
	LUT4 #(
		.INIT('h0301)
	) name132 (
		\priority[99] ,
		\priority[100] ,
		\priority[101] ,
		\req[99] ,
		_w390_
	);
	LUT4 #(
		.INIT('h0301)
	) name133 (
		\priority[105] ,
		\priority[106] ,
		\priority[107] ,
		\req[105] ,
		_w391_
	);
	LUT4 #(
		.INIT('h0301)
	) name134 (
		\priority[102] ,
		\priority[103] ,
		\priority[104] ,
		\req[102] ,
		_w392_
	);
	LUT4 #(
		.INIT('hd000)
	) name135 (
		_w385_,
		_w390_,
		_w391_,
		_w392_,
		_w393_
	);
	LUT2 #(
		.INIT('h1)
	) name136 (
		\req[104] ,
		\req[105] ,
		_w394_
	);
	LUT4 #(
		.INIT('h000b)
	) name137 (
		\priority[104] ,
		\req[103] ,
		\req[104] ,
		\req[105] ,
		_w395_
	);
	LUT2 #(
		.INIT('h1)
	) name138 (
		\req[110] ,
		\req[111] ,
		_w396_
	);
	LUT4 #(
		.INIT('h000b)
	) name139 (
		\priority[110] ,
		\req[109] ,
		\req[110] ,
		\req[111] ,
		_w397_
	);
	LUT2 #(
		.INIT('h1)
	) name140 (
		\req[107] ,
		\req[108] ,
		_w398_
	);
	LUT4 #(
		.INIT('h000b)
	) name141 (
		\priority[107] ,
		\req[106] ,
		\req[107] ,
		\req[108] ,
		_w399_
	);
	LUT4 #(
		.INIT('hd000)
	) name142 (
		_w391_,
		_w395_,
		_w397_,
		_w399_,
		_w400_
	);
	LUT4 #(
		.INIT('h0301)
	) name143 (
		\priority[108] ,
		\priority[109] ,
		\priority[110] ,
		\req[108] ,
		_w401_
	);
	LUT4 #(
		.INIT('h0301)
	) name144 (
		\priority[114] ,
		\priority[115] ,
		\priority[116] ,
		\req[114] ,
		_w402_
	);
	LUT4 #(
		.INIT('h0301)
	) name145 (
		\priority[111] ,
		\priority[112] ,
		\priority[113] ,
		\req[111] ,
		_w403_
	);
	LUT4 #(
		.INIT('hd000)
	) name146 (
		_w397_,
		_w401_,
		_w402_,
		_w403_,
		_w404_
	);
	LUT4 #(
		.INIT('h4f00)
	) name147 (
		_w389_,
		_w393_,
		_w400_,
		_w404_,
		_w405_
	);
	LUT2 #(
		.INIT('h1)
	) name148 (
		\req[113] ,
		\req[114] ,
		_w406_
	);
	LUT4 #(
		.INIT('h000b)
	) name149 (
		\priority[113] ,
		\req[112] ,
		\req[113] ,
		\req[114] ,
		_w407_
	);
	LUT2 #(
		.INIT('h1)
	) name150 (
		\req[119] ,
		\req[120] ,
		_w408_
	);
	LUT4 #(
		.INIT('h000b)
	) name151 (
		\priority[119] ,
		\req[118] ,
		\req[119] ,
		\req[120] ,
		_w409_
	);
	LUT2 #(
		.INIT('h1)
	) name152 (
		\req[116] ,
		\req[117] ,
		_w410_
	);
	LUT4 #(
		.INIT('h000b)
	) name153 (
		\priority[116] ,
		\req[115] ,
		\req[116] ,
		\req[117] ,
		_w411_
	);
	LUT4 #(
		.INIT('hd000)
	) name154 (
		_w402_,
		_w407_,
		_w409_,
		_w411_,
		_w412_
	);
	LUT4 #(
		.INIT('h0301)
	) name155 (
		\priority[117] ,
		\priority[118] ,
		\priority[119] ,
		\req[117] ,
		_w413_
	);
	LUT4 #(
		.INIT('h0301)
	) name156 (
		\priority[123] ,
		\priority[124] ,
		\priority[125] ,
		\req[123] ,
		_w414_
	);
	LUT4 #(
		.INIT('h0301)
	) name157 (
		\priority[120] ,
		\priority[121] ,
		\priority[122] ,
		\req[120] ,
		_w415_
	);
	LUT4 #(
		.INIT('hd000)
	) name158 (
		_w409_,
		_w413_,
		_w414_,
		_w415_,
		_w416_
	);
	LUT2 #(
		.INIT('h1)
	) name159 (
		\req[122] ,
		\req[123] ,
		_w417_
	);
	LUT4 #(
		.INIT('h000b)
	) name160 (
		\priority[122] ,
		\req[121] ,
		\req[122] ,
		\req[123] ,
		_w418_
	);
	LUT2 #(
		.INIT('h1)
	) name161 (
		\req[125] ,
		\req[126] ,
		_w419_
	);
	LUT4 #(
		.INIT('h000b)
	) name162 (
		\priority[125] ,
		\req[124] ,
		\req[125] ,
		\req[126] ,
		_w420_
	);
	LUT4 #(
		.INIT('ha200)
	) name163 (
		_w259_,
		_w414_,
		_w418_,
		_w420_,
		_w421_
	);
	LUT4 #(
		.INIT('h4f00)
	) name164 (
		_w405_,
		_w412_,
		_w416_,
		_w421_,
		_w422_
	);
	LUT2 #(
		.INIT('he)
	) name165 (
		_w260_,
		_w422_,
		_w423_
	);
	LUT4 #(
		.INIT('h1101)
	) name166 (
		\priority[0] ,
		\priority[1] ,
		\priority[127] ,
		\req[127] ,
		_w424_
	);
	LUT3 #(
		.INIT('hb0)
	) name167 (
		\priority[1] ,
		\req[0] ,
		\req[1] ,
		_w425_
	);
	LUT2 #(
		.INIT('h4)
	) name168 (
		_w424_,
		_w425_,
		_w426_
	);
	LUT3 #(
		.INIT('h31)
	) name169 (
		\priority[2] ,
		\priority[3] ,
		\req[2] ,
		_w427_
	);
	LUT2 #(
		.INIT('h1)
	) name170 (
		\req[3] ,
		\req[4] ,
		_w428_
	);
	LUT4 #(
		.INIT('h0301)
	) name171 (
		\priority[7] ,
		\priority[8] ,
		\priority[9] ,
		\req[7] ,
		_w429_
	);
	LUT4 #(
		.INIT('h0301)
	) name172 (
		\priority[4] ,
		\priority[5] ,
		\priority[6] ,
		\req[4] ,
		_w430_
	);
	LUT4 #(
		.INIT('hb000)
	) name173 (
		_w427_,
		_w428_,
		_w429_,
		_w430_,
		_w431_
	);
	LUT2 #(
		.INIT('h1)
	) name174 (
		\req[6] ,
		\req[7] ,
		_w432_
	);
	LUT4 #(
		.INIT('h000b)
	) name175 (
		\priority[6] ,
		\req[5] ,
		\req[6] ,
		\req[7] ,
		_w433_
	);
	LUT2 #(
		.INIT('h1)
	) name176 (
		\req[12] ,
		\req[13] ,
		_w434_
	);
	LUT4 #(
		.INIT('h000b)
	) name177 (
		\priority[12] ,
		\req[11] ,
		\req[12] ,
		\req[13] ,
		_w435_
	);
	LUT2 #(
		.INIT('h1)
	) name178 (
		\req[9] ,
		\req[10] ,
		_w436_
	);
	LUT4 #(
		.INIT('h000b)
	) name179 (
		\priority[9] ,
		\req[8] ,
		\req[9] ,
		\req[10] ,
		_w437_
	);
	LUT4 #(
		.INIT('hd000)
	) name180 (
		_w429_,
		_w433_,
		_w435_,
		_w437_,
		_w438_
	);
	LUT4 #(
		.INIT('h0301)
	) name181 (
		\priority[10] ,
		\priority[11] ,
		\priority[12] ,
		\req[10] ,
		_w439_
	);
	LUT4 #(
		.INIT('h0301)
	) name182 (
		\priority[16] ,
		\priority[17] ,
		\priority[18] ,
		\req[16] ,
		_w440_
	);
	LUT4 #(
		.INIT('h0301)
	) name183 (
		\priority[13] ,
		\priority[14] ,
		\priority[15] ,
		\req[13] ,
		_w441_
	);
	LUT4 #(
		.INIT('hd000)
	) name184 (
		_w435_,
		_w439_,
		_w440_,
		_w441_,
		_w442_
	);
	LUT2 #(
		.INIT('h1)
	) name185 (
		\req[15] ,
		\req[16] ,
		_w443_
	);
	LUT4 #(
		.INIT('h000b)
	) name186 (
		\priority[15] ,
		\req[14] ,
		\req[15] ,
		\req[16] ,
		_w444_
	);
	LUT2 #(
		.INIT('h1)
	) name187 (
		\req[21] ,
		\req[22] ,
		_w445_
	);
	LUT4 #(
		.INIT('h000b)
	) name188 (
		\priority[21] ,
		\req[20] ,
		\req[21] ,
		\req[22] ,
		_w446_
	);
	LUT2 #(
		.INIT('h1)
	) name189 (
		\req[18] ,
		\req[19] ,
		_w447_
	);
	LUT4 #(
		.INIT('h000b)
	) name190 (
		\priority[18] ,
		\req[17] ,
		\req[18] ,
		\req[19] ,
		_w448_
	);
	LUT4 #(
		.INIT('hd000)
	) name191 (
		_w440_,
		_w444_,
		_w446_,
		_w448_,
		_w449_
	);
	LUT4 #(
		.INIT('h4f00)
	) name192 (
		_w431_,
		_w438_,
		_w442_,
		_w449_,
		_w450_
	);
	LUT4 #(
		.INIT('h0301)
	) name193 (
		\priority[19] ,
		\priority[20] ,
		\priority[21] ,
		\req[19] ,
		_w451_
	);
	LUT4 #(
		.INIT('h0301)
	) name194 (
		\priority[25] ,
		\priority[26] ,
		\priority[27] ,
		\req[25] ,
		_w452_
	);
	LUT4 #(
		.INIT('h0301)
	) name195 (
		\priority[22] ,
		\priority[23] ,
		\priority[24] ,
		\req[22] ,
		_w453_
	);
	LUT4 #(
		.INIT('hd000)
	) name196 (
		_w446_,
		_w451_,
		_w452_,
		_w453_,
		_w454_
	);
	LUT2 #(
		.INIT('h1)
	) name197 (
		\req[24] ,
		\req[25] ,
		_w455_
	);
	LUT4 #(
		.INIT('h000b)
	) name198 (
		\priority[24] ,
		\req[23] ,
		\req[24] ,
		\req[25] ,
		_w456_
	);
	LUT2 #(
		.INIT('h1)
	) name199 (
		\req[30] ,
		\req[31] ,
		_w457_
	);
	LUT4 #(
		.INIT('h000b)
	) name200 (
		\priority[30] ,
		\req[29] ,
		\req[30] ,
		\req[31] ,
		_w458_
	);
	LUT2 #(
		.INIT('h1)
	) name201 (
		\req[27] ,
		\req[28] ,
		_w459_
	);
	LUT4 #(
		.INIT('h000b)
	) name202 (
		\priority[27] ,
		\req[26] ,
		\req[27] ,
		\req[28] ,
		_w460_
	);
	LUT4 #(
		.INIT('hd000)
	) name203 (
		_w452_,
		_w456_,
		_w458_,
		_w460_,
		_w461_
	);
	LUT4 #(
		.INIT('h0301)
	) name204 (
		\priority[28] ,
		\priority[29] ,
		\priority[30] ,
		\req[28] ,
		_w462_
	);
	LUT4 #(
		.INIT('h0301)
	) name205 (
		\priority[34] ,
		\priority[35] ,
		\priority[36] ,
		\req[34] ,
		_w463_
	);
	LUT4 #(
		.INIT('h0301)
	) name206 (
		\priority[31] ,
		\priority[32] ,
		\priority[33] ,
		\req[31] ,
		_w464_
	);
	LUT4 #(
		.INIT('hd000)
	) name207 (
		_w458_,
		_w462_,
		_w463_,
		_w464_,
		_w465_
	);
	LUT4 #(
		.INIT('h4f00)
	) name208 (
		_w450_,
		_w454_,
		_w461_,
		_w465_,
		_w466_
	);
	LUT2 #(
		.INIT('h1)
	) name209 (
		\req[33] ,
		\req[34] ,
		_w467_
	);
	LUT4 #(
		.INIT('h000b)
	) name210 (
		\priority[33] ,
		\req[32] ,
		\req[33] ,
		\req[34] ,
		_w468_
	);
	LUT2 #(
		.INIT('h1)
	) name211 (
		\req[39] ,
		\req[40] ,
		_w469_
	);
	LUT4 #(
		.INIT('h000b)
	) name212 (
		\priority[39] ,
		\req[38] ,
		\req[39] ,
		\req[40] ,
		_w470_
	);
	LUT2 #(
		.INIT('h1)
	) name213 (
		\req[36] ,
		\req[37] ,
		_w471_
	);
	LUT4 #(
		.INIT('h000b)
	) name214 (
		\priority[36] ,
		\req[35] ,
		\req[36] ,
		\req[37] ,
		_w472_
	);
	LUT4 #(
		.INIT('hd000)
	) name215 (
		_w463_,
		_w468_,
		_w470_,
		_w472_,
		_w473_
	);
	LUT4 #(
		.INIT('h0301)
	) name216 (
		\priority[37] ,
		\priority[38] ,
		\priority[39] ,
		\req[37] ,
		_w474_
	);
	LUT4 #(
		.INIT('h0301)
	) name217 (
		\priority[43] ,
		\priority[44] ,
		\priority[45] ,
		\req[43] ,
		_w475_
	);
	LUT4 #(
		.INIT('h0301)
	) name218 (
		\priority[40] ,
		\priority[41] ,
		\priority[42] ,
		\req[40] ,
		_w476_
	);
	LUT4 #(
		.INIT('hd000)
	) name219 (
		_w470_,
		_w474_,
		_w475_,
		_w476_,
		_w477_
	);
	LUT2 #(
		.INIT('h1)
	) name220 (
		\req[42] ,
		\req[43] ,
		_w478_
	);
	LUT4 #(
		.INIT('h000b)
	) name221 (
		\priority[42] ,
		\req[41] ,
		\req[42] ,
		\req[43] ,
		_w479_
	);
	LUT2 #(
		.INIT('h1)
	) name222 (
		\req[48] ,
		\req[49] ,
		_w480_
	);
	LUT4 #(
		.INIT('h000b)
	) name223 (
		\priority[48] ,
		\req[47] ,
		\req[48] ,
		\req[49] ,
		_w481_
	);
	LUT2 #(
		.INIT('h1)
	) name224 (
		\req[45] ,
		\req[46] ,
		_w482_
	);
	LUT4 #(
		.INIT('h000b)
	) name225 (
		\priority[45] ,
		\req[44] ,
		\req[45] ,
		\req[46] ,
		_w483_
	);
	LUT4 #(
		.INIT('hd000)
	) name226 (
		_w475_,
		_w479_,
		_w481_,
		_w483_,
		_w484_
	);
	LUT4 #(
		.INIT('h4f00)
	) name227 (
		_w466_,
		_w473_,
		_w477_,
		_w484_,
		_w485_
	);
	LUT4 #(
		.INIT('h0301)
	) name228 (
		\priority[46] ,
		\priority[47] ,
		\priority[48] ,
		\req[46] ,
		_w486_
	);
	LUT4 #(
		.INIT('h0301)
	) name229 (
		\priority[52] ,
		\priority[53] ,
		\priority[54] ,
		\req[52] ,
		_w487_
	);
	LUT4 #(
		.INIT('h0301)
	) name230 (
		\priority[49] ,
		\priority[50] ,
		\priority[51] ,
		\req[49] ,
		_w488_
	);
	LUT4 #(
		.INIT('hd000)
	) name231 (
		_w481_,
		_w486_,
		_w487_,
		_w488_,
		_w489_
	);
	LUT2 #(
		.INIT('h1)
	) name232 (
		\req[51] ,
		\req[52] ,
		_w490_
	);
	LUT4 #(
		.INIT('h000b)
	) name233 (
		\priority[51] ,
		\req[50] ,
		\req[51] ,
		\req[52] ,
		_w491_
	);
	LUT2 #(
		.INIT('h1)
	) name234 (
		\req[57] ,
		\req[58] ,
		_w492_
	);
	LUT4 #(
		.INIT('h000b)
	) name235 (
		\priority[57] ,
		\req[56] ,
		\req[57] ,
		\req[58] ,
		_w493_
	);
	LUT2 #(
		.INIT('h1)
	) name236 (
		\req[54] ,
		\req[55] ,
		_w494_
	);
	LUT4 #(
		.INIT('h000b)
	) name237 (
		\priority[54] ,
		\req[53] ,
		\req[54] ,
		\req[55] ,
		_w495_
	);
	LUT4 #(
		.INIT('hd000)
	) name238 (
		_w487_,
		_w491_,
		_w493_,
		_w495_,
		_w496_
	);
	LUT4 #(
		.INIT('h0301)
	) name239 (
		\priority[55] ,
		\priority[56] ,
		\priority[57] ,
		\req[55] ,
		_w497_
	);
	LUT4 #(
		.INIT('h0301)
	) name240 (
		\priority[61] ,
		\priority[62] ,
		\priority[63] ,
		\req[61] ,
		_w498_
	);
	LUT4 #(
		.INIT('h0301)
	) name241 (
		\priority[58] ,
		\priority[59] ,
		\priority[60] ,
		\req[58] ,
		_w499_
	);
	LUT4 #(
		.INIT('hd000)
	) name242 (
		_w493_,
		_w497_,
		_w498_,
		_w499_,
		_w500_
	);
	LUT4 #(
		.INIT('h4f00)
	) name243 (
		_w485_,
		_w489_,
		_w496_,
		_w500_,
		_w501_
	);
	LUT2 #(
		.INIT('h1)
	) name244 (
		\req[60] ,
		\req[61] ,
		_w502_
	);
	LUT4 #(
		.INIT('h000b)
	) name245 (
		\priority[60] ,
		\req[59] ,
		\req[60] ,
		\req[61] ,
		_w503_
	);
	LUT2 #(
		.INIT('h1)
	) name246 (
		\req[66] ,
		\req[67] ,
		_w504_
	);
	LUT4 #(
		.INIT('h000b)
	) name247 (
		\priority[66] ,
		\req[65] ,
		\req[66] ,
		\req[67] ,
		_w505_
	);
	LUT2 #(
		.INIT('h1)
	) name248 (
		\req[63] ,
		\req[64] ,
		_w506_
	);
	LUT4 #(
		.INIT('h000b)
	) name249 (
		\priority[63] ,
		\req[62] ,
		\req[63] ,
		\req[64] ,
		_w507_
	);
	LUT4 #(
		.INIT('hd000)
	) name250 (
		_w498_,
		_w503_,
		_w505_,
		_w507_,
		_w508_
	);
	LUT4 #(
		.INIT('h0301)
	) name251 (
		\priority[64] ,
		\priority[65] ,
		\priority[66] ,
		\req[64] ,
		_w509_
	);
	LUT4 #(
		.INIT('h0301)
	) name252 (
		\priority[70] ,
		\priority[71] ,
		\priority[72] ,
		\req[70] ,
		_w510_
	);
	LUT4 #(
		.INIT('h0301)
	) name253 (
		\priority[67] ,
		\priority[68] ,
		\priority[69] ,
		\req[67] ,
		_w511_
	);
	LUT4 #(
		.INIT('hd000)
	) name254 (
		_w505_,
		_w509_,
		_w510_,
		_w511_,
		_w512_
	);
	LUT2 #(
		.INIT('h1)
	) name255 (
		\req[69] ,
		\req[70] ,
		_w513_
	);
	LUT4 #(
		.INIT('h000b)
	) name256 (
		\priority[69] ,
		\req[68] ,
		\req[69] ,
		\req[70] ,
		_w514_
	);
	LUT2 #(
		.INIT('h1)
	) name257 (
		\req[75] ,
		\req[76] ,
		_w515_
	);
	LUT4 #(
		.INIT('h000b)
	) name258 (
		\priority[75] ,
		\req[74] ,
		\req[75] ,
		\req[76] ,
		_w516_
	);
	LUT2 #(
		.INIT('h1)
	) name259 (
		\req[72] ,
		\req[73] ,
		_w517_
	);
	LUT4 #(
		.INIT('h000b)
	) name260 (
		\priority[72] ,
		\req[71] ,
		\req[72] ,
		\req[73] ,
		_w518_
	);
	LUT4 #(
		.INIT('hd000)
	) name261 (
		_w510_,
		_w514_,
		_w516_,
		_w518_,
		_w519_
	);
	LUT4 #(
		.INIT('h4f00)
	) name262 (
		_w501_,
		_w508_,
		_w512_,
		_w519_,
		_w520_
	);
	LUT4 #(
		.INIT('h0301)
	) name263 (
		\priority[73] ,
		\priority[74] ,
		\priority[75] ,
		\req[73] ,
		_w521_
	);
	LUT4 #(
		.INIT('h0301)
	) name264 (
		\priority[79] ,
		\priority[80] ,
		\priority[81] ,
		\req[79] ,
		_w522_
	);
	LUT4 #(
		.INIT('h0301)
	) name265 (
		\priority[76] ,
		\priority[77] ,
		\priority[78] ,
		\req[76] ,
		_w523_
	);
	LUT4 #(
		.INIT('hd000)
	) name266 (
		_w516_,
		_w521_,
		_w522_,
		_w523_,
		_w524_
	);
	LUT2 #(
		.INIT('h1)
	) name267 (
		\req[78] ,
		\req[79] ,
		_w525_
	);
	LUT4 #(
		.INIT('h000b)
	) name268 (
		\priority[78] ,
		\req[77] ,
		\req[78] ,
		\req[79] ,
		_w526_
	);
	LUT2 #(
		.INIT('h1)
	) name269 (
		\req[84] ,
		\req[85] ,
		_w527_
	);
	LUT4 #(
		.INIT('h000b)
	) name270 (
		\priority[84] ,
		\req[83] ,
		\req[84] ,
		\req[85] ,
		_w528_
	);
	LUT2 #(
		.INIT('h1)
	) name271 (
		\req[81] ,
		\req[82] ,
		_w529_
	);
	LUT4 #(
		.INIT('h000b)
	) name272 (
		\priority[81] ,
		\req[80] ,
		\req[81] ,
		\req[82] ,
		_w530_
	);
	LUT4 #(
		.INIT('hd000)
	) name273 (
		_w522_,
		_w526_,
		_w528_,
		_w530_,
		_w531_
	);
	LUT4 #(
		.INIT('h0301)
	) name274 (
		\priority[82] ,
		\priority[83] ,
		\priority[84] ,
		\req[82] ,
		_w532_
	);
	LUT4 #(
		.INIT('h0301)
	) name275 (
		\priority[88] ,
		\priority[89] ,
		\priority[90] ,
		\req[88] ,
		_w533_
	);
	LUT4 #(
		.INIT('h0301)
	) name276 (
		\priority[85] ,
		\priority[86] ,
		\priority[87] ,
		\req[85] ,
		_w534_
	);
	LUT4 #(
		.INIT('hd000)
	) name277 (
		_w528_,
		_w532_,
		_w533_,
		_w534_,
		_w535_
	);
	LUT4 #(
		.INIT('h4f00)
	) name278 (
		_w520_,
		_w524_,
		_w531_,
		_w535_,
		_w536_
	);
	LUT2 #(
		.INIT('h1)
	) name279 (
		\req[87] ,
		\req[88] ,
		_w537_
	);
	LUT4 #(
		.INIT('h000b)
	) name280 (
		\priority[87] ,
		\req[86] ,
		\req[87] ,
		\req[88] ,
		_w538_
	);
	LUT2 #(
		.INIT('h1)
	) name281 (
		\req[93] ,
		\req[94] ,
		_w539_
	);
	LUT4 #(
		.INIT('h000b)
	) name282 (
		\priority[93] ,
		\req[92] ,
		\req[93] ,
		\req[94] ,
		_w540_
	);
	LUT2 #(
		.INIT('h1)
	) name283 (
		\req[90] ,
		\req[91] ,
		_w541_
	);
	LUT4 #(
		.INIT('h000b)
	) name284 (
		\priority[90] ,
		\req[89] ,
		\req[90] ,
		\req[91] ,
		_w542_
	);
	LUT4 #(
		.INIT('hd000)
	) name285 (
		_w533_,
		_w538_,
		_w540_,
		_w542_,
		_w543_
	);
	LUT4 #(
		.INIT('h0301)
	) name286 (
		\priority[91] ,
		\priority[92] ,
		\priority[93] ,
		\req[91] ,
		_w544_
	);
	LUT4 #(
		.INIT('h0301)
	) name287 (
		\priority[97] ,
		\priority[98] ,
		\priority[99] ,
		\req[97] ,
		_w545_
	);
	LUT4 #(
		.INIT('h0301)
	) name288 (
		\priority[94] ,
		\priority[95] ,
		\priority[96] ,
		\req[94] ,
		_w546_
	);
	LUT4 #(
		.INIT('hd000)
	) name289 (
		_w540_,
		_w544_,
		_w545_,
		_w546_,
		_w547_
	);
	LUT2 #(
		.INIT('h1)
	) name290 (
		\req[96] ,
		\req[97] ,
		_w548_
	);
	LUT4 #(
		.INIT('h000b)
	) name291 (
		\priority[96] ,
		\req[95] ,
		\req[96] ,
		\req[97] ,
		_w549_
	);
	LUT2 #(
		.INIT('h1)
	) name292 (
		\req[102] ,
		\req[103] ,
		_w550_
	);
	LUT4 #(
		.INIT('h000b)
	) name293 (
		\priority[102] ,
		\req[101] ,
		\req[102] ,
		\req[103] ,
		_w551_
	);
	LUT2 #(
		.INIT('h1)
	) name294 (
		\req[99] ,
		\req[100] ,
		_w552_
	);
	LUT4 #(
		.INIT('h000b)
	) name295 (
		\priority[99] ,
		\req[98] ,
		\req[99] ,
		\req[100] ,
		_w553_
	);
	LUT4 #(
		.INIT('hd000)
	) name296 (
		_w545_,
		_w549_,
		_w551_,
		_w553_,
		_w554_
	);
	LUT4 #(
		.INIT('h4f00)
	) name297 (
		_w536_,
		_w543_,
		_w547_,
		_w554_,
		_w555_
	);
	LUT4 #(
		.INIT('h0301)
	) name298 (
		\priority[100] ,
		\priority[101] ,
		\priority[102] ,
		\req[100] ,
		_w556_
	);
	LUT4 #(
		.INIT('h0301)
	) name299 (
		\priority[106] ,
		\priority[107] ,
		\priority[108] ,
		\req[106] ,
		_w557_
	);
	LUT4 #(
		.INIT('h0301)
	) name300 (
		\priority[103] ,
		\priority[104] ,
		\priority[105] ,
		\req[103] ,
		_w558_
	);
	LUT4 #(
		.INIT('hd000)
	) name301 (
		_w551_,
		_w556_,
		_w557_,
		_w558_,
		_w559_
	);
	LUT2 #(
		.INIT('h1)
	) name302 (
		\req[105] ,
		\req[106] ,
		_w560_
	);
	LUT4 #(
		.INIT('h000b)
	) name303 (
		\priority[105] ,
		\req[104] ,
		\req[105] ,
		\req[106] ,
		_w561_
	);
	LUT2 #(
		.INIT('h1)
	) name304 (
		\req[111] ,
		\req[112] ,
		_w562_
	);
	LUT4 #(
		.INIT('h000b)
	) name305 (
		\priority[111] ,
		\req[110] ,
		\req[111] ,
		\req[112] ,
		_w563_
	);
	LUT2 #(
		.INIT('h1)
	) name306 (
		\req[108] ,
		\req[109] ,
		_w564_
	);
	LUT4 #(
		.INIT('h000b)
	) name307 (
		\priority[108] ,
		\req[107] ,
		\req[108] ,
		\req[109] ,
		_w565_
	);
	LUT4 #(
		.INIT('hd000)
	) name308 (
		_w557_,
		_w561_,
		_w563_,
		_w565_,
		_w566_
	);
	LUT4 #(
		.INIT('h0301)
	) name309 (
		\priority[109] ,
		\priority[110] ,
		\priority[111] ,
		\req[109] ,
		_w567_
	);
	LUT4 #(
		.INIT('h0301)
	) name310 (
		\priority[115] ,
		\priority[116] ,
		\priority[117] ,
		\req[115] ,
		_w568_
	);
	LUT4 #(
		.INIT('h0301)
	) name311 (
		\priority[112] ,
		\priority[113] ,
		\priority[114] ,
		\req[112] ,
		_w569_
	);
	LUT4 #(
		.INIT('hd000)
	) name312 (
		_w563_,
		_w567_,
		_w568_,
		_w569_,
		_w570_
	);
	LUT4 #(
		.INIT('h4f00)
	) name313 (
		_w555_,
		_w559_,
		_w566_,
		_w570_,
		_w571_
	);
	LUT2 #(
		.INIT('h1)
	) name314 (
		\req[114] ,
		\req[115] ,
		_w572_
	);
	LUT4 #(
		.INIT('h000b)
	) name315 (
		\priority[114] ,
		\req[113] ,
		\req[114] ,
		\req[115] ,
		_w573_
	);
	LUT2 #(
		.INIT('h1)
	) name316 (
		\req[120] ,
		\req[121] ,
		_w574_
	);
	LUT4 #(
		.INIT('h000b)
	) name317 (
		\priority[120] ,
		\req[119] ,
		\req[120] ,
		\req[121] ,
		_w575_
	);
	LUT2 #(
		.INIT('h1)
	) name318 (
		\req[117] ,
		\req[118] ,
		_w576_
	);
	LUT4 #(
		.INIT('h000b)
	) name319 (
		\priority[117] ,
		\req[116] ,
		\req[117] ,
		\req[118] ,
		_w577_
	);
	LUT4 #(
		.INIT('hd000)
	) name320 (
		_w568_,
		_w573_,
		_w575_,
		_w577_,
		_w578_
	);
	LUT4 #(
		.INIT('h0301)
	) name321 (
		\priority[118] ,
		\priority[119] ,
		\priority[120] ,
		\req[118] ,
		_w579_
	);
	LUT4 #(
		.INIT('h0301)
	) name322 (
		\priority[124] ,
		\priority[125] ,
		\priority[126] ,
		\req[124] ,
		_w580_
	);
	LUT4 #(
		.INIT('h0301)
	) name323 (
		\priority[121] ,
		\priority[122] ,
		\priority[123] ,
		\req[121] ,
		_w581_
	);
	LUT4 #(
		.INIT('hd000)
	) name324 (
		_w575_,
		_w579_,
		_w580_,
		_w581_,
		_w582_
	);
	LUT2 #(
		.INIT('h1)
	) name325 (
		\req[123] ,
		\req[124] ,
		_w583_
	);
	LUT4 #(
		.INIT('h000b)
	) name326 (
		\priority[123] ,
		\req[122] ,
		\req[123] ,
		\req[124] ,
		_w584_
	);
	LUT2 #(
		.INIT('h1)
	) name327 (
		\req[126] ,
		\req[127] ,
		_w585_
	);
	LUT4 #(
		.INIT('h000b)
	) name328 (
		\priority[126] ,
		\req[125] ,
		\req[126] ,
		\req[127] ,
		_w586_
	);
	LUT4 #(
		.INIT('ha200)
	) name329 (
		_w425_,
		_w580_,
		_w584_,
		_w586_,
		_w587_
	);
	LUT4 #(
		.INIT('h4f00)
	) name330 (
		_w571_,
		_w578_,
		_w582_,
		_w587_,
		_w588_
	);
	LUT2 #(
		.INIT('he)
	) name331 (
		_w426_,
		_w588_,
		_w589_
	);
	LUT4 #(
		.INIT('h0301)
	) name332 (
		\priority[0] ,
		\priority[1] ,
		\priority[2] ,
		\req[0] ,
		_w590_
	);
	LUT3 #(
		.INIT('hb0)
	) name333 (
		\priority[2] ,
		\req[1] ,
		\req[2] ,
		_w591_
	);
	LUT2 #(
		.INIT('h4)
	) name334 (
		_w590_,
		_w591_,
		_w592_
	);
	LUT3 #(
		.INIT('h31)
	) name335 (
		\priority[3] ,
		\priority[4] ,
		\req[3] ,
		_w593_
	);
	LUT2 #(
		.INIT('h1)
	) name336 (
		\req[4] ,
		\req[5] ,
		_w594_
	);
	LUT4 #(
		.INIT('h0301)
	) name337 (
		\priority[8] ,
		\priority[9] ,
		\priority[10] ,
		\req[8] ,
		_w595_
	);
	LUT4 #(
		.INIT('h0301)
	) name338 (
		\priority[5] ,
		\priority[6] ,
		\priority[7] ,
		\req[5] ,
		_w596_
	);
	LUT4 #(
		.INIT('hb000)
	) name339 (
		_w593_,
		_w594_,
		_w595_,
		_w596_,
		_w597_
	);
	LUT2 #(
		.INIT('h1)
	) name340 (
		\req[7] ,
		\req[8] ,
		_w598_
	);
	LUT4 #(
		.INIT('h000b)
	) name341 (
		\priority[7] ,
		\req[6] ,
		\req[7] ,
		\req[8] ,
		_w599_
	);
	LUT2 #(
		.INIT('h1)
	) name342 (
		\req[13] ,
		\req[14] ,
		_w600_
	);
	LUT4 #(
		.INIT('h000b)
	) name343 (
		\priority[13] ,
		\req[12] ,
		\req[13] ,
		\req[14] ,
		_w601_
	);
	LUT2 #(
		.INIT('h1)
	) name344 (
		\req[10] ,
		\req[11] ,
		_w602_
	);
	LUT4 #(
		.INIT('h000b)
	) name345 (
		\priority[10] ,
		\req[9] ,
		\req[10] ,
		\req[11] ,
		_w603_
	);
	LUT4 #(
		.INIT('hd000)
	) name346 (
		_w595_,
		_w599_,
		_w601_,
		_w603_,
		_w604_
	);
	LUT4 #(
		.INIT('h0301)
	) name347 (
		\priority[11] ,
		\priority[12] ,
		\priority[13] ,
		\req[11] ,
		_w605_
	);
	LUT4 #(
		.INIT('h0301)
	) name348 (
		\priority[17] ,
		\priority[18] ,
		\priority[19] ,
		\req[17] ,
		_w606_
	);
	LUT4 #(
		.INIT('h0301)
	) name349 (
		\priority[14] ,
		\priority[15] ,
		\priority[16] ,
		\req[14] ,
		_w607_
	);
	LUT4 #(
		.INIT('hd000)
	) name350 (
		_w601_,
		_w605_,
		_w606_,
		_w607_,
		_w608_
	);
	LUT2 #(
		.INIT('h1)
	) name351 (
		\req[16] ,
		\req[17] ,
		_w609_
	);
	LUT4 #(
		.INIT('h000b)
	) name352 (
		\priority[16] ,
		\req[15] ,
		\req[16] ,
		\req[17] ,
		_w610_
	);
	LUT2 #(
		.INIT('h1)
	) name353 (
		\req[22] ,
		\req[23] ,
		_w611_
	);
	LUT4 #(
		.INIT('h000b)
	) name354 (
		\priority[22] ,
		\req[21] ,
		\req[22] ,
		\req[23] ,
		_w612_
	);
	LUT2 #(
		.INIT('h1)
	) name355 (
		\req[19] ,
		\req[20] ,
		_w613_
	);
	LUT4 #(
		.INIT('h000b)
	) name356 (
		\priority[19] ,
		\req[18] ,
		\req[19] ,
		\req[20] ,
		_w614_
	);
	LUT4 #(
		.INIT('hd000)
	) name357 (
		_w606_,
		_w610_,
		_w612_,
		_w614_,
		_w615_
	);
	LUT4 #(
		.INIT('h4f00)
	) name358 (
		_w597_,
		_w604_,
		_w608_,
		_w615_,
		_w616_
	);
	LUT4 #(
		.INIT('h0301)
	) name359 (
		\priority[20] ,
		\priority[21] ,
		\priority[22] ,
		\req[20] ,
		_w617_
	);
	LUT4 #(
		.INIT('h0301)
	) name360 (
		\priority[26] ,
		\priority[27] ,
		\priority[28] ,
		\req[26] ,
		_w618_
	);
	LUT4 #(
		.INIT('h0301)
	) name361 (
		\priority[23] ,
		\priority[24] ,
		\priority[25] ,
		\req[23] ,
		_w619_
	);
	LUT4 #(
		.INIT('hd000)
	) name362 (
		_w612_,
		_w617_,
		_w618_,
		_w619_,
		_w620_
	);
	LUT2 #(
		.INIT('h1)
	) name363 (
		\req[25] ,
		\req[26] ,
		_w621_
	);
	LUT4 #(
		.INIT('h000b)
	) name364 (
		\priority[25] ,
		\req[24] ,
		\req[25] ,
		\req[26] ,
		_w622_
	);
	LUT2 #(
		.INIT('h1)
	) name365 (
		\req[31] ,
		\req[32] ,
		_w623_
	);
	LUT4 #(
		.INIT('h000b)
	) name366 (
		\priority[31] ,
		\req[30] ,
		\req[31] ,
		\req[32] ,
		_w624_
	);
	LUT2 #(
		.INIT('h1)
	) name367 (
		\req[28] ,
		\req[29] ,
		_w625_
	);
	LUT4 #(
		.INIT('h000b)
	) name368 (
		\priority[28] ,
		\req[27] ,
		\req[28] ,
		\req[29] ,
		_w626_
	);
	LUT4 #(
		.INIT('hd000)
	) name369 (
		_w618_,
		_w622_,
		_w624_,
		_w626_,
		_w627_
	);
	LUT4 #(
		.INIT('h0301)
	) name370 (
		\priority[29] ,
		\priority[30] ,
		\priority[31] ,
		\req[29] ,
		_w628_
	);
	LUT4 #(
		.INIT('h0301)
	) name371 (
		\priority[35] ,
		\priority[36] ,
		\priority[37] ,
		\req[35] ,
		_w629_
	);
	LUT4 #(
		.INIT('h0301)
	) name372 (
		\priority[32] ,
		\priority[33] ,
		\priority[34] ,
		\req[32] ,
		_w630_
	);
	LUT4 #(
		.INIT('hd000)
	) name373 (
		_w624_,
		_w628_,
		_w629_,
		_w630_,
		_w631_
	);
	LUT4 #(
		.INIT('h4f00)
	) name374 (
		_w616_,
		_w620_,
		_w627_,
		_w631_,
		_w632_
	);
	LUT2 #(
		.INIT('h1)
	) name375 (
		\req[34] ,
		\req[35] ,
		_w633_
	);
	LUT4 #(
		.INIT('h000b)
	) name376 (
		\priority[34] ,
		\req[33] ,
		\req[34] ,
		\req[35] ,
		_w634_
	);
	LUT2 #(
		.INIT('h1)
	) name377 (
		\req[40] ,
		\req[41] ,
		_w635_
	);
	LUT4 #(
		.INIT('h000b)
	) name378 (
		\priority[40] ,
		\req[39] ,
		\req[40] ,
		\req[41] ,
		_w636_
	);
	LUT2 #(
		.INIT('h1)
	) name379 (
		\req[37] ,
		\req[38] ,
		_w637_
	);
	LUT4 #(
		.INIT('h000b)
	) name380 (
		\priority[37] ,
		\req[36] ,
		\req[37] ,
		\req[38] ,
		_w638_
	);
	LUT4 #(
		.INIT('hd000)
	) name381 (
		_w629_,
		_w634_,
		_w636_,
		_w638_,
		_w639_
	);
	LUT4 #(
		.INIT('h0301)
	) name382 (
		\priority[38] ,
		\priority[39] ,
		\priority[40] ,
		\req[38] ,
		_w640_
	);
	LUT4 #(
		.INIT('h0301)
	) name383 (
		\priority[44] ,
		\priority[45] ,
		\priority[46] ,
		\req[44] ,
		_w641_
	);
	LUT4 #(
		.INIT('h0301)
	) name384 (
		\priority[41] ,
		\priority[42] ,
		\priority[43] ,
		\req[41] ,
		_w642_
	);
	LUT4 #(
		.INIT('hd000)
	) name385 (
		_w636_,
		_w640_,
		_w641_,
		_w642_,
		_w643_
	);
	LUT2 #(
		.INIT('h1)
	) name386 (
		\req[43] ,
		\req[44] ,
		_w644_
	);
	LUT4 #(
		.INIT('h000b)
	) name387 (
		\priority[43] ,
		\req[42] ,
		\req[43] ,
		\req[44] ,
		_w645_
	);
	LUT2 #(
		.INIT('h1)
	) name388 (
		\req[49] ,
		\req[50] ,
		_w646_
	);
	LUT4 #(
		.INIT('h000b)
	) name389 (
		\priority[49] ,
		\req[48] ,
		\req[49] ,
		\req[50] ,
		_w647_
	);
	LUT2 #(
		.INIT('h1)
	) name390 (
		\req[46] ,
		\req[47] ,
		_w648_
	);
	LUT4 #(
		.INIT('h000b)
	) name391 (
		\priority[46] ,
		\req[45] ,
		\req[46] ,
		\req[47] ,
		_w649_
	);
	LUT4 #(
		.INIT('hd000)
	) name392 (
		_w641_,
		_w645_,
		_w647_,
		_w649_,
		_w650_
	);
	LUT4 #(
		.INIT('h4f00)
	) name393 (
		_w632_,
		_w639_,
		_w643_,
		_w650_,
		_w651_
	);
	LUT4 #(
		.INIT('h0301)
	) name394 (
		\priority[47] ,
		\priority[48] ,
		\priority[49] ,
		\req[47] ,
		_w652_
	);
	LUT4 #(
		.INIT('h0301)
	) name395 (
		\priority[53] ,
		\priority[54] ,
		\priority[55] ,
		\req[53] ,
		_w653_
	);
	LUT4 #(
		.INIT('h0301)
	) name396 (
		\priority[50] ,
		\priority[51] ,
		\priority[52] ,
		\req[50] ,
		_w654_
	);
	LUT4 #(
		.INIT('hd000)
	) name397 (
		_w647_,
		_w652_,
		_w653_,
		_w654_,
		_w655_
	);
	LUT2 #(
		.INIT('h1)
	) name398 (
		\req[52] ,
		\req[53] ,
		_w656_
	);
	LUT4 #(
		.INIT('h000b)
	) name399 (
		\priority[52] ,
		\req[51] ,
		\req[52] ,
		\req[53] ,
		_w657_
	);
	LUT2 #(
		.INIT('h1)
	) name400 (
		\req[58] ,
		\req[59] ,
		_w658_
	);
	LUT4 #(
		.INIT('h000b)
	) name401 (
		\priority[58] ,
		\req[57] ,
		\req[58] ,
		\req[59] ,
		_w659_
	);
	LUT2 #(
		.INIT('h1)
	) name402 (
		\req[55] ,
		\req[56] ,
		_w660_
	);
	LUT4 #(
		.INIT('h000b)
	) name403 (
		\priority[55] ,
		\req[54] ,
		\req[55] ,
		\req[56] ,
		_w661_
	);
	LUT4 #(
		.INIT('hd000)
	) name404 (
		_w653_,
		_w657_,
		_w659_,
		_w661_,
		_w662_
	);
	LUT4 #(
		.INIT('h0301)
	) name405 (
		\priority[56] ,
		\priority[57] ,
		\priority[58] ,
		\req[56] ,
		_w663_
	);
	LUT4 #(
		.INIT('h0301)
	) name406 (
		\priority[62] ,
		\priority[63] ,
		\priority[64] ,
		\req[62] ,
		_w664_
	);
	LUT4 #(
		.INIT('h0301)
	) name407 (
		\priority[59] ,
		\priority[60] ,
		\priority[61] ,
		\req[59] ,
		_w665_
	);
	LUT4 #(
		.INIT('hd000)
	) name408 (
		_w659_,
		_w663_,
		_w664_,
		_w665_,
		_w666_
	);
	LUT4 #(
		.INIT('h4f00)
	) name409 (
		_w651_,
		_w655_,
		_w662_,
		_w666_,
		_w667_
	);
	LUT2 #(
		.INIT('h1)
	) name410 (
		\req[61] ,
		\req[62] ,
		_w668_
	);
	LUT4 #(
		.INIT('h000b)
	) name411 (
		\priority[61] ,
		\req[60] ,
		\req[61] ,
		\req[62] ,
		_w669_
	);
	LUT2 #(
		.INIT('h1)
	) name412 (
		\req[67] ,
		\req[68] ,
		_w670_
	);
	LUT4 #(
		.INIT('h000b)
	) name413 (
		\priority[67] ,
		\req[66] ,
		\req[67] ,
		\req[68] ,
		_w671_
	);
	LUT2 #(
		.INIT('h1)
	) name414 (
		\req[64] ,
		\req[65] ,
		_w672_
	);
	LUT4 #(
		.INIT('h000b)
	) name415 (
		\priority[64] ,
		\req[63] ,
		\req[64] ,
		\req[65] ,
		_w673_
	);
	LUT4 #(
		.INIT('hd000)
	) name416 (
		_w664_,
		_w669_,
		_w671_,
		_w673_,
		_w674_
	);
	LUT4 #(
		.INIT('h0301)
	) name417 (
		\priority[65] ,
		\priority[66] ,
		\priority[67] ,
		\req[65] ,
		_w675_
	);
	LUT4 #(
		.INIT('h0301)
	) name418 (
		\priority[71] ,
		\priority[72] ,
		\priority[73] ,
		\req[71] ,
		_w676_
	);
	LUT4 #(
		.INIT('h0301)
	) name419 (
		\priority[68] ,
		\priority[69] ,
		\priority[70] ,
		\req[68] ,
		_w677_
	);
	LUT4 #(
		.INIT('hd000)
	) name420 (
		_w671_,
		_w675_,
		_w676_,
		_w677_,
		_w678_
	);
	LUT2 #(
		.INIT('h1)
	) name421 (
		\req[70] ,
		\req[71] ,
		_w679_
	);
	LUT4 #(
		.INIT('h000b)
	) name422 (
		\priority[70] ,
		\req[69] ,
		\req[70] ,
		\req[71] ,
		_w680_
	);
	LUT2 #(
		.INIT('h1)
	) name423 (
		\req[76] ,
		\req[77] ,
		_w681_
	);
	LUT4 #(
		.INIT('h000b)
	) name424 (
		\priority[76] ,
		\req[75] ,
		\req[76] ,
		\req[77] ,
		_w682_
	);
	LUT2 #(
		.INIT('h1)
	) name425 (
		\req[73] ,
		\req[74] ,
		_w683_
	);
	LUT4 #(
		.INIT('h000b)
	) name426 (
		\priority[73] ,
		\req[72] ,
		\req[73] ,
		\req[74] ,
		_w684_
	);
	LUT4 #(
		.INIT('hd000)
	) name427 (
		_w676_,
		_w680_,
		_w682_,
		_w684_,
		_w685_
	);
	LUT4 #(
		.INIT('h4f00)
	) name428 (
		_w667_,
		_w674_,
		_w678_,
		_w685_,
		_w686_
	);
	LUT4 #(
		.INIT('h0301)
	) name429 (
		\priority[74] ,
		\priority[75] ,
		\priority[76] ,
		\req[74] ,
		_w687_
	);
	LUT4 #(
		.INIT('h0301)
	) name430 (
		\priority[80] ,
		\priority[81] ,
		\priority[82] ,
		\req[80] ,
		_w688_
	);
	LUT4 #(
		.INIT('h0301)
	) name431 (
		\priority[77] ,
		\priority[78] ,
		\priority[79] ,
		\req[77] ,
		_w689_
	);
	LUT4 #(
		.INIT('hd000)
	) name432 (
		_w682_,
		_w687_,
		_w688_,
		_w689_,
		_w690_
	);
	LUT2 #(
		.INIT('h1)
	) name433 (
		\req[79] ,
		\req[80] ,
		_w691_
	);
	LUT4 #(
		.INIT('h000b)
	) name434 (
		\priority[79] ,
		\req[78] ,
		\req[79] ,
		\req[80] ,
		_w692_
	);
	LUT2 #(
		.INIT('h1)
	) name435 (
		\req[85] ,
		\req[86] ,
		_w693_
	);
	LUT4 #(
		.INIT('h000b)
	) name436 (
		\priority[85] ,
		\req[84] ,
		\req[85] ,
		\req[86] ,
		_w694_
	);
	LUT2 #(
		.INIT('h1)
	) name437 (
		\req[82] ,
		\req[83] ,
		_w695_
	);
	LUT4 #(
		.INIT('h000b)
	) name438 (
		\priority[82] ,
		\req[81] ,
		\req[82] ,
		\req[83] ,
		_w696_
	);
	LUT4 #(
		.INIT('hd000)
	) name439 (
		_w688_,
		_w692_,
		_w694_,
		_w696_,
		_w697_
	);
	LUT4 #(
		.INIT('h0301)
	) name440 (
		\priority[83] ,
		\priority[84] ,
		\priority[85] ,
		\req[83] ,
		_w698_
	);
	LUT4 #(
		.INIT('h0301)
	) name441 (
		\priority[89] ,
		\priority[90] ,
		\priority[91] ,
		\req[89] ,
		_w699_
	);
	LUT4 #(
		.INIT('h0301)
	) name442 (
		\priority[86] ,
		\priority[87] ,
		\priority[88] ,
		\req[86] ,
		_w700_
	);
	LUT4 #(
		.INIT('hd000)
	) name443 (
		_w694_,
		_w698_,
		_w699_,
		_w700_,
		_w701_
	);
	LUT4 #(
		.INIT('h4f00)
	) name444 (
		_w686_,
		_w690_,
		_w697_,
		_w701_,
		_w702_
	);
	LUT2 #(
		.INIT('h1)
	) name445 (
		\req[88] ,
		\req[89] ,
		_w703_
	);
	LUT4 #(
		.INIT('h000b)
	) name446 (
		\priority[88] ,
		\req[87] ,
		\req[88] ,
		\req[89] ,
		_w704_
	);
	LUT2 #(
		.INIT('h1)
	) name447 (
		\req[94] ,
		\req[95] ,
		_w705_
	);
	LUT4 #(
		.INIT('h000b)
	) name448 (
		\priority[94] ,
		\req[93] ,
		\req[94] ,
		\req[95] ,
		_w706_
	);
	LUT2 #(
		.INIT('h1)
	) name449 (
		\req[91] ,
		\req[92] ,
		_w707_
	);
	LUT4 #(
		.INIT('h000b)
	) name450 (
		\priority[91] ,
		\req[90] ,
		\req[91] ,
		\req[92] ,
		_w708_
	);
	LUT4 #(
		.INIT('hd000)
	) name451 (
		_w699_,
		_w704_,
		_w706_,
		_w708_,
		_w709_
	);
	LUT4 #(
		.INIT('h0301)
	) name452 (
		\priority[92] ,
		\priority[93] ,
		\priority[94] ,
		\req[92] ,
		_w710_
	);
	LUT4 #(
		.INIT('h0301)
	) name453 (
		\priority[98] ,
		\priority[99] ,
		\priority[100] ,
		\req[98] ,
		_w711_
	);
	LUT4 #(
		.INIT('h0301)
	) name454 (
		\priority[95] ,
		\priority[96] ,
		\priority[97] ,
		\req[95] ,
		_w712_
	);
	LUT4 #(
		.INIT('hd000)
	) name455 (
		_w706_,
		_w710_,
		_w711_,
		_w712_,
		_w713_
	);
	LUT2 #(
		.INIT('h1)
	) name456 (
		\req[97] ,
		\req[98] ,
		_w714_
	);
	LUT4 #(
		.INIT('h000b)
	) name457 (
		\priority[97] ,
		\req[96] ,
		\req[97] ,
		\req[98] ,
		_w715_
	);
	LUT2 #(
		.INIT('h1)
	) name458 (
		\req[103] ,
		\req[104] ,
		_w716_
	);
	LUT4 #(
		.INIT('h000b)
	) name459 (
		\priority[103] ,
		\req[102] ,
		\req[103] ,
		\req[104] ,
		_w717_
	);
	LUT2 #(
		.INIT('h1)
	) name460 (
		\req[100] ,
		\req[101] ,
		_w718_
	);
	LUT4 #(
		.INIT('h000b)
	) name461 (
		\priority[100] ,
		\req[99] ,
		\req[100] ,
		\req[101] ,
		_w719_
	);
	LUT4 #(
		.INIT('hd000)
	) name462 (
		_w711_,
		_w715_,
		_w717_,
		_w719_,
		_w720_
	);
	LUT4 #(
		.INIT('h4f00)
	) name463 (
		_w702_,
		_w709_,
		_w713_,
		_w720_,
		_w721_
	);
	LUT4 #(
		.INIT('h0301)
	) name464 (
		\priority[101] ,
		\priority[102] ,
		\priority[103] ,
		\req[101] ,
		_w722_
	);
	LUT4 #(
		.INIT('h0301)
	) name465 (
		\priority[107] ,
		\priority[108] ,
		\priority[109] ,
		\req[107] ,
		_w723_
	);
	LUT4 #(
		.INIT('h0301)
	) name466 (
		\priority[104] ,
		\priority[105] ,
		\priority[106] ,
		\req[104] ,
		_w724_
	);
	LUT4 #(
		.INIT('hd000)
	) name467 (
		_w717_,
		_w722_,
		_w723_,
		_w724_,
		_w725_
	);
	LUT2 #(
		.INIT('h1)
	) name468 (
		\req[106] ,
		\req[107] ,
		_w726_
	);
	LUT4 #(
		.INIT('h000b)
	) name469 (
		\priority[106] ,
		\req[105] ,
		\req[106] ,
		\req[107] ,
		_w727_
	);
	LUT2 #(
		.INIT('h1)
	) name470 (
		\req[112] ,
		\req[113] ,
		_w728_
	);
	LUT4 #(
		.INIT('h000b)
	) name471 (
		\priority[112] ,
		\req[111] ,
		\req[112] ,
		\req[113] ,
		_w729_
	);
	LUT2 #(
		.INIT('h1)
	) name472 (
		\req[109] ,
		\req[110] ,
		_w730_
	);
	LUT4 #(
		.INIT('h000b)
	) name473 (
		\priority[109] ,
		\req[108] ,
		\req[109] ,
		\req[110] ,
		_w731_
	);
	LUT4 #(
		.INIT('hd000)
	) name474 (
		_w723_,
		_w727_,
		_w729_,
		_w731_,
		_w732_
	);
	LUT4 #(
		.INIT('h0301)
	) name475 (
		\priority[110] ,
		\priority[111] ,
		\priority[112] ,
		\req[110] ,
		_w733_
	);
	LUT4 #(
		.INIT('h0301)
	) name476 (
		\priority[116] ,
		\priority[117] ,
		\priority[118] ,
		\req[116] ,
		_w734_
	);
	LUT4 #(
		.INIT('h0301)
	) name477 (
		\priority[113] ,
		\priority[114] ,
		\priority[115] ,
		\req[113] ,
		_w735_
	);
	LUT4 #(
		.INIT('hd000)
	) name478 (
		_w729_,
		_w733_,
		_w734_,
		_w735_,
		_w736_
	);
	LUT4 #(
		.INIT('h4f00)
	) name479 (
		_w721_,
		_w725_,
		_w732_,
		_w736_,
		_w737_
	);
	LUT2 #(
		.INIT('h1)
	) name480 (
		\req[115] ,
		\req[116] ,
		_w738_
	);
	LUT4 #(
		.INIT('h000b)
	) name481 (
		\priority[115] ,
		\req[114] ,
		\req[115] ,
		\req[116] ,
		_w739_
	);
	LUT2 #(
		.INIT('h1)
	) name482 (
		\req[121] ,
		\req[122] ,
		_w740_
	);
	LUT4 #(
		.INIT('h000b)
	) name483 (
		\priority[121] ,
		\req[120] ,
		\req[121] ,
		\req[122] ,
		_w741_
	);
	LUT2 #(
		.INIT('h1)
	) name484 (
		\req[118] ,
		\req[119] ,
		_w742_
	);
	LUT4 #(
		.INIT('h000b)
	) name485 (
		\priority[118] ,
		\req[117] ,
		\req[118] ,
		\req[119] ,
		_w743_
	);
	LUT4 #(
		.INIT('hd000)
	) name486 (
		_w734_,
		_w739_,
		_w741_,
		_w743_,
		_w744_
	);
	LUT4 #(
		.INIT('h0301)
	) name487 (
		\priority[119] ,
		\priority[120] ,
		\priority[121] ,
		\req[119] ,
		_w745_
	);
	LUT4 #(
		.INIT('h0301)
	) name488 (
		\priority[125] ,
		\priority[126] ,
		\priority[127] ,
		\req[125] ,
		_w746_
	);
	LUT4 #(
		.INIT('h0301)
	) name489 (
		\priority[122] ,
		\priority[123] ,
		\priority[124] ,
		\req[122] ,
		_w747_
	);
	LUT4 #(
		.INIT('hd000)
	) name490 (
		_w741_,
		_w745_,
		_w746_,
		_w747_,
		_w748_
	);
	LUT2 #(
		.INIT('h1)
	) name491 (
		\req[124] ,
		\req[125] ,
		_w749_
	);
	LUT4 #(
		.INIT('h000b)
	) name492 (
		\priority[124] ,
		\req[123] ,
		\req[124] ,
		\req[125] ,
		_w750_
	);
	LUT2 #(
		.INIT('h1)
	) name493 (
		\req[0] ,
		\req[127] ,
		_w751_
	);
	LUT4 #(
		.INIT('h0023)
	) name494 (
		\priority[127] ,
		\req[0] ,
		\req[126] ,
		\req[127] ,
		_w752_
	);
	LUT4 #(
		.INIT('ha200)
	) name495 (
		_w591_,
		_w746_,
		_w750_,
		_w752_,
		_w753_
	);
	LUT4 #(
		.INIT('h4f00)
	) name496 (
		_w737_,
		_w744_,
		_w748_,
		_w753_,
		_w754_
	);
	LUT2 #(
		.INIT('he)
	) name497 (
		_w592_,
		_w754_,
		_w755_
	);
	LUT4 #(
		.INIT('h0301)
	) name498 (
		\priority[1] ,
		\priority[2] ,
		\priority[3] ,
		\req[1] ,
		_w756_
	);
	LUT3 #(
		.INIT('hb0)
	) name499 (
		\priority[3] ,
		\req[2] ,
		\req[3] ,
		_w757_
	);
	LUT2 #(
		.INIT('h4)
	) name500 (
		_w756_,
		_w757_,
		_w758_
	);
	LUT3 #(
		.INIT('h31)
	) name501 (
		\priority[4] ,
		\priority[5] ,
		\req[4] ,
		_w759_
	);
	LUT4 #(
		.INIT('ha020)
	) name502 (
		_w263_,
		_w266_,
		_w273_,
		_w759_,
		_w760_
	);
	LUT4 #(
		.INIT('h8a00)
	) name503 (
		_w269_,
		_w271_,
		_w273_,
		_w278_,
		_w761_
	);
	LUT4 #(
		.INIT('h8a00)
	) name504 (
		_w274_,
		_w275_,
		_w278_,
		_w285_,
		_w762_
	);
	LUT4 #(
		.INIT('h8a00)
	) name505 (
		_w280_,
		_w282_,
		_w285_,
		_w290_,
		_w763_
	);
	LUT4 #(
		.INIT('h4f00)
	) name506 (
		_w760_,
		_w761_,
		_w762_,
		_w763_,
		_w764_
	);
	LUT4 #(
		.INIT('h8a00)
	) name507 (
		_w286_,
		_w287_,
		_w290_,
		_w296_,
		_w765_
	);
	LUT4 #(
		.INIT('h8a00)
	) name508 (
		_w292_,
		_w294_,
		_w296_,
		_w302_,
		_w766_
	);
	LUT4 #(
		.INIT('h8a00)
	) name509 (
		_w297_,
		_w298_,
		_w302_,
		_w308_,
		_w767_
	);
	LUT4 #(
		.INIT('h4f00)
	) name510 (
		_w764_,
		_w765_,
		_w766_,
		_w767_,
		_w768_
	);
	LUT4 #(
		.INIT('h8a00)
	) name511 (
		_w304_,
		_w306_,
		_w308_,
		_w313_,
		_w769_
	);
	LUT4 #(
		.INIT('h8a00)
	) name512 (
		_w309_,
		_w310_,
		_w313_,
		_w320_,
		_w770_
	);
	LUT4 #(
		.INIT('h8a00)
	) name513 (
		_w315_,
		_w317_,
		_w320_,
		_w325_,
		_w771_
	);
	LUT4 #(
		.INIT('h4f00)
	) name514 (
		_w768_,
		_w769_,
		_w770_,
		_w771_,
		_w772_
	);
	LUT4 #(
		.INIT('h8a00)
	) name515 (
		_w321_,
		_w322_,
		_w325_,
		_w331_,
		_w773_
	);
	LUT4 #(
		.INIT('h8a00)
	) name516 (
		_w327_,
		_w329_,
		_w331_,
		_w337_,
		_w774_
	);
	LUT4 #(
		.INIT('h8a00)
	) name517 (
		_w332_,
		_w333_,
		_w337_,
		_w343_,
		_w775_
	);
	LUT4 #(
		.INIT('h4f00)
	) name518 (
		_w772_,
		_w773_,
		_w774_,
		_w775_,
		_w776_
	);
	LUT4 #(
		.INIT('h8a00)
	) name519 (
		_w339_,
		_w341_,
		_w343_,
		_w348_,
		_w777_
	);
	LUT4 #(
		.INIT('h8a00)
	) name520 (
		_w344_,
		_w345_,
		_w348_,
		_w355_,
		_w778_
	);
	LUT4 #(
		.INIT('h8a00)
	) name521 (
		_w350_,
		_w352_,
		_w355_,
		_w360_,
		_w779_
	);
	LUT4 #(
		.INIT('h4f00)
	) name522 (
		_w776_,
		_w777_,
		_w778_,
		_w779_,
		_w780_
	);
	LUT4 #(
		.INIT('h8a00)
	) name523 (
		_w356_,
		_w357_,
		_w360_,
		_w366_,
		_w781_
	);
	LUT4 #(
		.INIT('h8a00)
	) name524 (
		_w362_,
		_w364_,
		_w366_,
		_w372_,
		_w782_
	);
	LUT4 #(
		.INIT('h8a00)
	) name525 (
		_w367_,
		_w368_,
		_w372_,
		_w378_,
		_w783_
	);
	LUT4 #(
		.INIT('h4f00)
	) name526 (
		_w780_,
		_w781_,
		_w782_,
		_w783_,
		_w784_
	);
	LUT4 #(
		.INIT('h8a00)
	) name527 (
		_w374_,
		_w376_,
		_w378_,
		_w383_,
		_w785_
	);
	LUT4 #(
		.INIT('h8a00)
	) name528 (
		_w379_,
		_w380_,
		_w383_,
		_w390_,
		_w786_
	);
	LUT4 #(
		.INIT('h8a00)
	) name529 (
		_w385_,
		_w387_,
		_w390_,
		_w395_,
		_w787_
	);
	LUT4 #(
		.INIT('h4f00)
	) name530 (
		_w784_,
		_w785_,
		_w786_,
		_w787_,
		_w788_
	);
	LUT4 #(
		.INIT('h8a00)
	) name531 (
		_w391_,
		_w392_,
		_w395_,
		_w401_,
		_w789_
	);
	LUT4 #(
		.INIT('h8a00)
	) name532 (
		_w397_,
		_w399_,
		_w401_,
		_w407_,
		_w790_
	);
	LUT4 #(
		.INIT('h8a00)
	) name533 (
		_w402_,
		_w403_,
		_w407_,
		_w413_,
		_w791_
	);
	LUT4 #(
		.INIT('h4f00)
	) name534 (
		_w788_,
		_w789_,
		_w790_,
		_w791_,
		_w792_
	);
	LUT4 #(
		.INIT('h8a00)
	) name535 (
		_w409_,
		_w411_,
		_w413_,
		_w418_,
		_w793_
	);
	LUT4 #(
		.INIT('h8088)
	) name536 (
		_w258_,
		_w414_,
		_w415_,
		_w418_,
		_w794_
	);
	LUT2 #(
		.INIT('h1)
	) name537 (
		\req[0] ,
		\req[1] ,
		_w795_
	);
	LUT4 #(
		.INIT('h0203)
	) name538 (
		\priority[0] ,
		\req[0] ,
		\req[1] ,
		\req[127] ,
		_w796_
	);
	LUT4 #(
		.INIT('hd000)
	) name539 (
		_w258_,
		_w420_,
		_w757_,
		_w796_,
		_w797_
	);
	LUT4 #(
		.INIT('h4f00)
	) name540 (
		_w792_,
		_w793_,
		_w794_,
		_w797_,
		_w798_
	);
	LUT2 #(
		.INIT('he)
	) name541 (
		_w758_,
		_w798_,
		_w799_
	);
	LUT4 #(
		.INIT('h0301)
	) name542 (
		\priority[2] ,
		\priority[3] ,
		\priority[4] ,
		\req[2] ,
		_w800_
	);
	LUT3 #(
		.INIT('hb0)
	) name543 (
		\priority[4] ,
		\req[3] ,
		\req[4] ,
		_w801_
	);
	LUT2 #(
		.INIT('h4)
	) name544 (
		_w800_,
		_w801_,
		_w802_
	);
	LUT3 #(
		.INIT('h31)
	) name545 (
		\priority[5] ,
		\priority[6] ,
		\req[5] ,
		_w803_
	);
	LUT4 #(
		.INIT('ha020)
	) name546 (
		_w429_,
		_w432_,
		_w439_,
		_w803_,
		_w804_
	);
	LUT4 #(
		.INIT('h8a00)
	) name547 (
		_w435_,
		_w437_,
		_w439_,
		_w444_,
		_w805_
	);
	LUT4 #(
		.INIT('h8a00)
	) name548 (
		_w440_,
		_w441_,
		_w444_,
		_w451_,
		_w806_
	);
	LUT4 #(
		.INIT('h8a00)
	) name549 (
		_w446_,
		_w448_,
		_w451_,
		_w456_,
		_w807_
	);
	LUT4 #(
		.INIT('h4f00)
	) name550 (
		_w804_,
		_w805_,
		_w806_,
		_w807_,
		_w808_
	);
	LUT4 #(
		.INIT('h8a00)
	) name551 (
		_w452_,
		_w453_,
		_w456_,
		_w462_,
		_w809_
	);
	LUT4 #(
		.INIT('h8a00)
	) name552 (
		_w458_,
		_w460_,
		_w462_,
		_w468_,
		_w810_
	);
	LUT4 #(
		.INIT('h8a00)
	) name553 (
		_w463_,
		_w464_,
		_w468_,
		_w474_,
		_w811_
	);
	LUT4 #(
		.INIT('h4f00)
	) name554 (
		_w808_,
		_w809_,
		_w810_,
		_w811_,
		_w812_
	);
	LUT4 #(
		.INIT('h8a00)
	) name555 (
		_w470_,
		_w472_,
		_w474_,
		_w479_,
		_w813_
	);
	LUT4 #(
		.INIT('h8a00)
	) name556 (
		_w475_,
		_w476_,
		_w479_,
		_w486_,
		_w814_
	);
	LUT4 #(
		.INIT('h8a00)
	) name557 (
		_w481_,
		_w483_,
		_w486_,
		_w491_,
		_w815_
	);
	LUT4 #(
		.INIT('h4f00)
	) name558 (
		_w812_,
		_w813_,
		_w814_,
		_w815_,
		_w816_
	);
	LUT4 #(
		.INIT('h8a00)
	) name559 (
		_w487_,
		_w488_,
		_w491_,
		_w497_,
		_w817_
	);
	LUT4 #(
		.INIT('h8a00)
	) name560 (
		_w493_,
		_w495_,
		_w497_,
		_w503_,
		_w818_
	);
	LUT4 #(
		.INIT('h8a00)
	) name561 (
		_w498_,
		_w499_,
		_w503_,
		_w509_,
		_w819_
	);
	LUT4 #(
		.INIT('h4f00)
	) name562 (
		_w816_,
		_w817_,
		_w818_,
		_w819_,
		_w820_
	);
	LUT4 #(
		.INIT('h8a00)
	) name563 (
		_w505_,
		_w507_,
		_w509_,
		_w514_,
		_w821_
	);
	LUT4 #(
		.INIT('h8a00)
	) name564 (
		_w510_,
		_w511_,
		_w514_,
		_w521_,
		_w822_
	);
	LUT4 #(
		.INIT('h8a00)
	) name565 (
		_w516_,
		_w518_,
		_w521_,
		_w526_,
		_w823_
	);
	LUT4 #(
		.INIT('h4f00)
	) name566 (
		_w820_,
		_w821_,
		_w822_,
		_w823_,
		_w824_
	);
	LUT4 #(
		.INIT('h8a00)
	) name567 (
		_w522_,
		_w523_,
		_w526_,
		_w532_,
		_w825_
	);
	LUT4 #(
		.INIT('h8a00)
	) name568 (
		_w528_,
		_w530_,
		_w532_,
		_w538_,
		_w826_
	);
	LUT4 #(
		.INIT('h8a00)
	) name569 (
		_w533_,
		_w534_,
		_w538_,
		_w544_,
		_w827_
	);
	LUT4 #(
		.INIT('h4f00)
	) name570 (
		_w824_,
		_w825_,
		_w826_,
		_w827_,
		_w828_
	);
	LUT4 #(
		.INIT('h8a00)
	) name571 (
		_w540_,
		_w542_,
		_w544_,
		_w549_,
		_w829_
	);
	LUT4 #(
		.INIT('h8a00)
	) name572 (
		_w545_,
		_w546_,
		_w549_,
		_w556_,
		_w830_
	);
	LUT4 #(
		.INIT('h8a00)
	) name573 (
		_w551_,
		_w553_,
		_w556_,
		_w561_,
		_w831_
	);
	LUT4 #(
		.INIT('h4f00)
	) name574 (
		_w828_,
		_w829_,
		_w830_,
		_w831_,
		_w832_
	);
	LUT4 #(
		.INIT('h8a00)
	) name575 (
		_w557_,
		_w558_,
		_w561_,
		_w567_,
		_w833_
	);
	LUT4 #(
		.INIT('h8a00)
	) name576 (
		_w563_,
		_w565_,
		_w567_,
		_w573_,
		_w834_
	);
	LUT4 #(
		.INIT('h8a00)
	) name577 (
		_w568_,
		_w569_,
		_w573_,
		_w579_,
		_w835_
	);
	LUT4 #(
		.INIT('h4f00)
	) name578 (
		_w832_,
		_w833_,
		_w834_,
		_w835_,
		_w836_
	);
	LUT4 #(
		.INIT('h8a00)
	) name579 (
		_w575_,
		_w577_,
		_w579_,
		_w584_,
		_w837_
	);
	LUT4 #(
		.INIT('h8088)
	) name580 (
		_w424_,
		_w580_,
		_w581_,
		_w584_,
		_w838_
	);
	LUT2 #(
		.INIT('h1)
	) name581 (
		\req[1] ,
		\req[2] ,
		_w839_
	);
	LUT4 #(
		.INIT('h000b)
	) name582 (
		\priority[1] ,
		\req[0] ,
		\req[1] ,
		\req[2] ,
		_w840_
	);
	LUT4 #(
		.INIT('hd000)
	) name583 (
		_w424_,
		_w586_,
		_w801_,
		_w840_,
		_w841_
	);
	LUT4 #(
		.INIT('h4f00)
	) name584 (
		_w836_,
		_w837_,
		_w838_,
		_w841_,
		_w842_
	);
	LUT2 #(
		.INIT('he)
	) name585 (
		_w802_,
		_w842_,
		_w843_
	);
	LUT3 #(
		.INIT('hb0)
	) name586 (
		\priority[5] ,
		\req[4] ,
		\req[5] ,
		_w844_
	);
	LUT2 #(
		.INIT('h4)
	) name587 (
		_w264_,
		_w844_,
		_w845_
	);
	LUT3 #(
		.INIT('h31)
	) name588 (
		\priority[6] ,
		\priority[7] ,
		\req[6] ,
		_w846_
	);
	LUT4 #(
		.INIT('ha020)
	) name589 (
		_w595_,
		_w598_,
		_w605_,
		_w846_,
		_w847_
	);
	LUT4 #(
		.INIT('h8a00)
	) name590 (
		_w601_,
		_w603_,
		_w605_,
		_w610_,
		_w848_
	);
	LUT4 #(
		.INIT('h8a00)
	) name591 (
		_w606_,
		_w607_,
		_w610_,
		_w617_,
		_w849_
	);
	LUT4 #(
		.INIT('h8a00)
	) name592 (
		_w612_,
		_w614_,
		_w617_,
		_w622_,
		_w850_
	);
	LUT4 #(
		.INIT('h4f00)
	) name593 (
		_w847_,
		_w848_,
		_w849_,
		_w850_,
		_w851_
	);
	LUT4 #(
		.INIT('h8a00)
	) name594 (
		_w618_,
		_w619_,
		_w622_,
		_w628_,
		_w852_
	);
	LUT4 #(
		.INIT('h8a00)
	) name595 (
		_w624_,
		_w626_,
		_w628_,
		_w634_,
		_w853_
	);
	LUT4 #(
		.INIT('h8a00)
	) name596 (
		_w629_,
		_w630_,
		_w634_,
		_w640_,
		_w854_
	);
	LUT4 #(
		.INIT('h4f00)
	) name597 (
		_w851_,
		_w852_,
		_w853_,
		_w854_,
		_w855_
	);
	LUT4 #(
		.INIT('h8a00)
	) name598 (
		_w636_,
		_w638_,
		_w640_,
		_w645_,
		_w856_
	);
	LUT4 #(
		.INIT('h8a00)
	) name599 (
		_w641_,
		_w642_,
		_w645_,
		_w652_,
		_w857_
	);
	LUT4 #(
		.INIT('h8a00)
	) name600 (
		_w647_,
		_w649_,
		_w652_,
		_w657_,
		_w858_
	);
	LUT4 #(
		.INIT('h4f00)
	) name601 (
		_w855_,
		_w856_,
		_w857_,
		_w858_,
		_w859_
	);
	LUT4 #(
		.INIT('h8a00)
	) name602 (
		_w653_,
		_w654_,
		_w657_,
		_w663_,
		_w860_
	);
	LUT4 #(
		.INIT('h8a00)
	) name603 (
		_w659_,
		_w661_,
		_w663_,
		_w669_,
		_w861_
	);
	LUT4 #(
		.INIT('h8a00)
	) name604 (
		_w664_,
		_w665_,
		_w669_,
		_w675_,
		_w862_
	);
	LUT4 #(
		.INIT('h4f00)
	) name605 (
		_w859_,
		_w860_,
		_w861_,
		_w862_,
		_w863_
	);
	LUT4 #(
		.INIT('h8a00)
	) name606 (
		_w671_,
		_w673_,
		_w675_,
		_w680_,
		_w864_
	);
	LUT4 #(
		.INIT('h8a00)
	) name607 (
		_w676_,
		_w677_,
		_w680_,
		_w687_,
		_w865_
	);
	LUT4 #(
		.INIT('h8a00)
	) name608 (
		_w682_,
		_w684_,
		_w687_,
		_w692_,
		_w866_
	);
	LUT4 #(
		.INIT('h4f00)
	) name609 (
		_w863_,
		_w864_,
		_w865_,
		_w866_,
		_w867_
	);
	LUT4 #(
		.INIT('h8a00)
	) name610 (
		_w688_,
		_w689_,
		_w692_,
		_w698_,
		_w868_
	);
	LUT4 #(
		.INIT('h8a00)
	) name611 (
		_w694_,
		_w696_,
		_w698_,
		_w704_,
		_w869_
	);
	LUT4 #(
		.INIT('h8a00)
	) name612 (
		_w699_,
		_w700_,
		_w704_,
		_w710_,
		_w870_
	);
	LUT4 #(
		.INIT('h4f00)
	) name613 (
		_w867_,
		_w868_,
		_w869_,
		_w870_,
		_w871_
	);
	LUT4 #(
		.INIT('h8a00)
	) name614 (
		_w706_,
		_w708_,
		_w710_,
		_w715_,
		_w872_
	);
	LUT4 #(
		.INIT('h8a00)
	) name615 (
		_w711_,
		_w712_,
		_w715_,
		_w722_,
		_w873_
	);
	LUT4 #(
		.INIT('h8a00)
	) name616 (
		_w717_,
		_w719_,
		_w722_,
		_w727_,
		_w874_
	);
	LUT4 #(
		.INIT('h4f00)
	) name617 (
		_w871_,
		_w872_,
		_w873_,
		_w874_,
		_w875_
	);
	LUT4 #(
		.INIT('h8a00)
	) name618 (
		_w723_,
		_w724_,
		_w727_,
		_w733_,
		_w876_
	);
	LUT4 #(
		.INIT('h8a00)
	) name619 (
		_w729_,
		_w731_,
		_w733_,
		_w739_,
		_w877_
	);
	LUT4 #(
		.INIT('h8a00)
	) name620 (
		_w734_,
		_w735_,
		_w739_,
		_w745_,
		_w878_
	);
	LUT4 #(
		.INIT('h4f00)
	) name621 (
		_w875_,
		_w876_,
		_w877_,
		_w878_,
		_w879_
	);
	LUT4 #(
		.INIT('h8a00)
	) name622 (
		_w741_,
		_w743_,
		_w745_,
		_w750_,
		_w880_
	);
	LUT4 #(
		.INIT('h8088)
	) name623 (
		_w590_,
		_w746_,
		_w747_,
		_w750_,
		_w881_
	);
	LUT4 #(
		.INIT('h000b)
	) name624 (
		\priority[2] ,
		\req[1] ,
		\req[2] ,
		\req[3] ,
		_w882_
	);
	LUT4 #(
		.INIT('hd000)
	) name625 (
		_w590_,
		_w752_,
		_w844_,
		_w882_,
		_w883_
	);
	LUT4 #(
		.INIT('h4f00)
	) name626 (
		_w879_,
		_w880_,
		_w881_,
		_w883_,
		_w884_
	);
	LUT2 #(
		.INIT('he)
	) name627 (
		_w845_,
		_w884_,
		_w885_
	);
	LUT3 #(
		.INIT('hb0)
	) name628 (
		\priority[6] ,
		\req[5] ,
		\req[6] ,
		_w886_
	);
	LUT2 #(
		.INIT('h4)
	) name629 (
		_w430_,
		_w886_,
		_w887_
	);
	LUT3 #(
		.INIT('h31)
	) name630 (
		\priority[7] ,
		\priority[8] ,
		\req[7] ,
		_w888_
	);
	LUT4 #(
		.INIT('hc040)
	) name631 (
		_w270_,
		_w273_,
		_w275_,
		_w888_,
		_w889_
	);
	LUT4 #(
		.INIT('hb000)
	) name632 (
		_w269_,
		_w275_,
		_w278_,
		_w282_,
		_w890_
	);
	LUT4 #(
		.INIT('hb000)
	) name633 (
		_w274_,
		_w282_,
		_w285_,
		_w287_,
		_w891_
	);
	LUT4 #(
		.INIT('hb000)
	) name634 (
		_w280_,
		_w287_,
		_w290_,
		_w294_,
		_w892_
	);
	LUT4 #(
		.INIT('h4f00)
	) name635 (
		_w889_,
		_w890_,
		_w891_,
		_w892_,
		_w893_
	);
	LUT4 #(
		.INIT('hb000)
	) name636 (
		_w286_,
		_w294_,
		_w296_,
		_w298_,
		_w894_
	);
	LUT4 #(
		.INIT('hb000)
	) name637 (
		_w292_,
		_w298_,
		_w302_,
		_w306_,
		_w895_
	);
	LUT4 #(
		.INIT('hb000)
	) name638 (
		_w297_,
		_w306_,
		_w308_,
		_w310_,
		_w896_
	);
	LUT4 #(
		.INIT('h4f00)
	) name639 (
		_w893_,
		_w894_,
		_w895_,
		_w896_,
		_w897_
	);
	LUT4 #(
		.INIT('hb000)
	) name640 (
		_w304_,
		_w310_,
		_w313_,
		_w317_,
		_w898_
	);
	LUT4 #(
		.INIT('hb000)
	) name641 (
		_w309_,
		_w317_,
		_w320_,
		_w322_,
		_w899_
	);
	LUT4 #(
		.INIT('hb000)
	) name642 (
		_w315_,
		_w322_,
		_w325_,
		_w329_,
		_w900_
	);
	LUT4 #(
		.INIT('h4f00)
	) name643 (
		_w897_,
		_w898_,
		_w899_,
		_w900_,
		_w901_
	);
	LUT4 #(
		.INIT('hb000)
	) name644 (
		_w321_,
		_w329_,
		_w331_,
		_w333_,
		_w902_
	);
	LUT4 #(
		.INIT('hb000)
	) name645 (
		_w327_,
		_w333_,
		_w337_,
		_w341_,
		_w903_
	);
	LUT4 #(
		.INIT('hb000)
	) name646 (
		_w332_,
		_w341_,
		_w343_,
		_w345_,
		_w904_
	);
	LUT4 #(
		.INIT('h4f00)
	) name647 (
		_w901_,
		_w902_,
		_w903_,
		_w904_,
		_w905_
	);
	LUT4 #(
		.INIT('hb000)
	) name648 (
		_w339_,
		_w345_,
		_w348_,
		_w352_,
		_w906_
	);
	LUT4 #(
		.INIT('hb000)
	) name649 (
		_w344_,
		_w352_,
		_w355_,
		_w357_,
		_w907_
	);
	LUT4 #(
		.INIT('hb000)
	) name650 (
		_w350_,
		_w357_,
		_w360_,
		_w364_,
		_w908_
	);
	LUT4 #(
		.INIT('h4f00)
	) name651 (
		_w905_,
		_w906_,
		_w907_,
		_w908_,
		_w909_
	);
	LUT4 #(
		.INIT('hb000)
	) name652 (
		_w356_,
		_w364_,
		_w366_,
		_w368_,
		_w910_
	);
	LUT4 #(
		.INIT('hb000)
	) name653 (
		_w362_,
		_w368_,
		_w372_,
		_w376_,
		_w911_
	);
	LUT4 #(
		.INIT('hb000)
	) name654 (
		_w367_,
		_w376_,
		_w378_,
		_w380_,
		_w912_
	);
	LUT4 #(
		.INIT('h4f00)
	) name655 (
		_w909_,
		_w910_,
		_w911_,
		_w912_,
		_w913_
	);
	LUT4 #(
		.INIT('hb000)
	) name656 (
		_w374_,
		_w380_,
		_w383_,
		_w387_,
		_w914_
	);
	LUT4 #(
		.INIT('hb000)
	) name657 (
		_w379_,
		_w387_,
		_w390_,
		_w392_,
		_w915_
	);
	LUT4 #(
		.INIT('hb000)
	) name658 (
		_w385_,
		_w392_,
		_w395_,
		_w399_,
		_w916_
	);
	LUT4 #(
		.INIT('h4f00)
	) name659 (
		_w913_,
		_w914_,
		_w915_,
		_w916_,
		_w917_
	);
	LUT4 #(
		.INIT('hb000)
	) name660 (
		_w391_,
		_w399_,
		_w401_,
		_w403_,
		_w918_
	);
	LUT4 #(
		.INIT('hb000)
	) name661 (
		_w397_,
		_w403_,
		_w407_,
		_w411_,
		_w919_
	);
	LUT4 #(
		.INIT('hb000)
	) name662 (
		_w402_,
		_w411_,
		_w413_,
		_w415_,
		_w920_
	);
	LUT4 #(
		.INIT('h4f00)
	) name663 (
		_w917_,
		_w918_,
		_w919_,
		_w920_,
		_w921_
	);
	LUT4 #(
		.INIT('hb000)
	) name664 (
		_w409_,
		_w415_,
		_w418_,
		_w420_,
		_w922_
	);
	LUT4 #(
		.INIT('h8a00)
	) name665 (
		_w258_,
		_w414_,
		_w420_,
		_w756_,
		_w923_
	);
	LUT4 #(
		.INIT('h000b)
	) name666 (
		\priority[3] ,
		\req[2] ,
		\req[3] ,
		\req[4] ,
		_w924_
	);
	LUT4 #(
		.INIT('hd000)
	) name667 (
		_w756_,
		_w796_,
		_w886_,
		_w924_,
		_w925_
	);
	LUT4 #(
		.INIT('h4f00)
	) name668 (
		_w921_,
		_w922_,
		_w923_,
		_w925_,
		_w926_
	);
	LUT2 #(
		.INIT('he)
	) name669 (
		_w887_,
		_w926_,
		_w927_
	);
	LUT3 #(
		.INIT('hb0)
	) name670 (
		\priority[7] ,
		\req[6] ,
		\req[7] ,
		_w928_
	);
	LUT2 #(
		.INIT('h4)
	) name671 (
		_w596_,
		_w928_,
		_w929_
	);
	LUT3 #(
		.INIT('h31)
	) name672 (
		\priority[8] ,
		\priority[9] ,
		\req[8] ,
		_w930_
	);
	LUT4 #(
		.INIT('hc040)
	) name673 (
		_w436_,
		_w439_,
		_w441_,
		_w930_,
		_w931_
	);
	LUT4 #(
		.INIT('hb000)
	) name674 (
		_w435_,
		_w441_,
		_w444_,
		_w448_,
		_w932_
	);
	LUT4 #(
		.INIT('hb000)
	) name675 (
		_w440_,
		_w448_,
		_w451_,
		_w453_,
		_w933_
	);
	LUT4 #(
		.INIT('hb000)
	) name676 (
		_w446_,
		_w453_,
		_w456_,
		_w460_,
		_w934_
	);
	LUT4 #(
		.INIT('h4f00)
	) name677 (
		_w931_,
		_w932_,
		_w933_,
		_w934_,
		_w935_
	);
	LUT4 #(
		.INIT('hb000)
	) name678 (
		_w452_,
		_w460_,
		_w462_,
		_w464_,
		_w936_
	);
	LUT4 #(
		.INIT('hb000)
	) name679 (
		_w458_,
		_w464_,
		_w468_,
		_w472_,
		_w937_
	);
	LUT4 #(
		.INIT('hb000)
	) name680 (
		_w463_,
		_w472_,
		_w474_,
		_w476_,
		_w938_
	);
	LUT4 #(
		.INIT('h4f00)
	) name681 (
		_w935_,
		_w936_,
		_w937_,
		_w938_,
		_w939_
	);
	LUT4 #(
		.INIT('hb000)
	) name682 (
		_w470_,
		_w476_,
		_w479_,
		_w483_,
		_w940_
	);
	LUT4 #(
		.INIT('hb000)
	) name683 (
		_w475_,
		_w483_,
		_w486_,
		_w488_,
		_w941_
	);
	LUT4 #(
		.INIT('hb000)
	) name684 (
		_w481_,
		_w488_,
		_w491_,
		_w495_,
		_w942_
	);
	LUT4 #(
		.INIT('h4f00)
	) name685 (
		_w939_,
		_w940_,
		_w941_,
		_w942_,
		_w943_
	);
	LUT4 #(
		.INIT('hb000)
	) name686 (
		_w487_,
		_w495_,
		_w497_,
		_w499_,
		_w944_
	);
	LUT4 #(
		.INIT('hb000)
	) name687 (
		_w493_,
		_w499_,
		_w503_,
		_w507_,
		_w945_
	);
	LUT4 #(
		.INIT('hb000)
	) name688 (
		_w498_,
		_w507_,
		_w509_,
		_w511_,
		_w946_
	);
	LUT4 #(
		.INIT('h4f00)
	) name689 (
		_w943_,
		_w944_,
		_w945_,
		_w946_,
		_w947_
	);
	LUT4 #(
		.INIT('hb000)
	) name690 (
		_w505_,
		_w511_,
		_w514_,
		_w518_,
		_w948_
	);
	LUT4 #(
		.INIT('hb000)
	) name691 (
		_w510_,
		_w518_,
		_w521_,
		_w523_,
		_w949_
	);
	LUT4 #(
		.INIT('hb000)
	) name692 (
		_w516_,
		_w523_,
		_w526_,
		_w530_,
		_w950_
	);
	LUT4 #(
		.INIT('h4f00)
	) name693 (
		_w947_,
		_w948_,
		_w949_,
		_w950_,
		_w951_
	);
	LUT4 #(
		.INIT('hb000)
	) name694 (
		_w522_,
		_w530_,
		_w532_,
		_w534_,
		_w952_
	);
	LUT4 #(
		.INIT('hb000)
	) name695 (
		_w528_,
		_w534_,
		_w538_,
		_w542_,
		_w953_
	);
	LUT4 #(
		.INIT('hb000)
	) name696 (
		_w533_,
		_w542_,
		_w544_,
		_w546_,
		_w954_
	);
	LUT4 #(
		.INIT('h4f00)
	) name697 (
		_w951_,
		_w952_,
		_w953_,
		_w954_,
		_w955_
	);
	LUT4 #(
		.INIT('hb000)
	) name698 (
		_w540_,
		_w546_,
		_w549_,
		_w553_,
		_w956_
	);
	LUT4 #(
		.INIT('hb000)
	) name699 (
		_w545_,
		_w553_,
		_w556_,
		_w558_,
		_w957_
	);
	LUT4 #(
		.INIT('hb000)
	) name700 (
		_w551_,
		_w558_,
		_w561_,
		_w565_,
		_w958_
	);
	LUT4 #(
		.INIT('h4f00)
	) name701 (
		_w955_,
		_w956_,
		_w957_,
		_w958_,
		_w959_
	);
	LUT4 #(
		.INIT('hb000)
	) name702 (
		_w557_,
		_w565_,
		_w567_,
		_w569_,
		_w960_
	);
	LUT4 #(
		.INIT('hb000)
	) name703 (
		_w563_,
		_w569_,
		_w573_,
		_w577_,
		_w961_
	);
	LUT4 #(
		.INIT('hb000)
	) name704 (
		_w568_,
		_w577_,
		_w579_,
		_w581_,
		_w962_
	);
	LUT4 #(
		.INIT('h4f00)
	) name705 (
		_w959_,
		_w960_,
		_w961_,
		_w962_,
		_w963_
	);
	LUT4 #(
		.INIT('hb000)
	) name706 (
		_w575_,
		_w581_,
		_w584_,
		_w586_,
		_w964_
	);
	LUT4 #(
		.INIT('h8a00)
	) name707 (
		_w424_,
		_w580_,
		_w586_,
		_w800_,
		_w965_
	);
	LUT4 #(
		.INIT('h000b)
	) name708 (
		\priority[4] ,
		\req[3] ,
		\req[4] ,
		\req[5] ,
		_w966_
	);
	LUT4 #(
		.INIT('hd000)
	) name709 (
		_w800_,
		_w840_,
		_w928_,
		_w966_,
		_w967_
	);
	LUT4 #(
		.INIT('h4f00)
	) name710 (
		_w963_,
		_w964_,
		_w965_,
		_w967_,
		_w968_
	);
	LUT2 #(
		.INIT('he)
	) name711 (
		_w929_,
		_w968_,
		_w969_
	);
	LUT3 #(
		.INIT('hb0)
	) name712 (
		\priority[8] ,
		\req[7] ,
		\req[8] ,
		_w970_
	);
	LUT2 #(
		.INIT('h4)
	) name713 (
		_w263_,
		_w970_,
		_w971_
	);
	LUT3 #(
		.INIT('h31)
	) name714 (
		\priority[9] ,
		\priority[10] ,
		\req[9] ,
		_w972_
	);
	LUT4 #(
		.INIT('hc040)
	) name715 (
		_w602_,
		_w605_,
		_w607_,
		_w972_,
		_w973_
	);
	LUT4 #(
		.INIT('hb000)
	) name716 (
		_w601_,
		_w607_,
		_w610_,
		_w614_,
		_w974_
	);
	LUT4 #(
		.INIT('hb000)
	) name717 (
		_w606_,
		_w614_,
		_w617_,
		_w619_,
		_w975_
	);
	LUT4 #(
		.INIT('hb000)
	) name718 (
		_w612_,
		_w619_,
		_w622_,
		_w626_,
		_w976_
	);
	LUT4 #(
		.INIT('h4f00)
	) name719 (
		_w973_,
		_w974_,
		_w975_,
		_w976_,
		_w977_
	);
	LUT4 #(
		.INIT('hb000)
	) name720 (
		_w618_,
		_w626_,
		_w628_,
		_w630_,
		_w978_
	);
	LUT4 #(
		.INIT('hb000)
	) name721 (
		_w624_,
		_w630_,
		_w634_,
		_w638_,
		_w979_
	);
	LUT4 #(
		.INIT('hb000)
	) name722 (
		_w629_,
		_w638_,
		_w640_,
		_w642_,
		_w980_
	);
	LUT4 #(
		.INIT('h4f00)
	) name723 (
		_w977_,
		_w978_,
		_w979_,
		_w980_,
		_w981_
	);
	LUT4 #(
		.INIT('hb000)
	) name724 (
		_w636_,
		_w642_,
		_w645_,
		_w649_,
		_w982_
	);
	LUT4 #(
		.INIT('hb000)
	) name725 (
		_w641_,
		_w649_,
		_w652_,
		_w654_,
		_w983_
	);
	LUT4 #(
		.INIT('hb000)
	) name726 (
		_w647_,
		_w654_,
		_w657_,
		_w661_,
		_w984_
	);
	LUT4 #(
		.INIT('h4f00)
	) name727 (
		_w981_,
		_w982_,
		_w983_,
		_w984_,
		_w985_
	);
	LUT4 #(
		.INIT('hb000)
	) name728 (
		_w653_,
		_w661_,
		_w663_,
		_w665_,
		_w986_
	);
	LUT4 #(
		.INIT('hb000)
	) name729 (
		_w659_,
		_w665_,
		_w669_,
		_w673_,
		_w987_
	);
	LUT4 #(
		.INIT('hb000)
	) name730 (
		_w664_,
		_w673_,
		_w675_,
		_w677_,
		_w988_
	);
	LUT4 #(
		.INIT('h4f00)
	) name731 (
		_w985_,
		_w986_,
		_w987_,
		_w988_,
		_w989_
	);
	LUT4 #(
		.INIT('hb000)
	) name732 (
		_w671_,
		_w677_,
		_w680_,
		_w684_,
		_w990_
	);
	LUT4 #(
		.INIT('hb000)
	) name733 (
		_w676_,
		_w684_,
		_w687_,
		_w689_,
		_w991_
	);
	LUT4 #(
		.INIT('hb000)
	) name734 (
		_w682_,
		_w689_,
		_w692_,
		_w696_,
		_w992_
	);
	LUT4 #(
		.INIT('h4f00)
	) name735 (
		_w989_,
		_w990_,
		_w991_,
		_w992_,
		_w993_
	);
	LUT4 #(
		.INIT('hb000)
	) name736 (
		_w688_,
		_w696_,
		_w698_,
		_w700_,
		_w994_
	);
	LUT4 #(
		.INIT('hb000)
	) name737 (
		_w694_,
		_w700_,
		_w704_,
		_w708_,
		_w995_
	);
	LUT4 #(
		.INIT('hb000)
	) name738 (
		_w699_,
		_w708_,
		_w710_,
		_w712_,
		_w996_
	);
	LUT4 #(
		.INIT('h4f00)
	) name739 (
		_w993_,
		_w994_,
		_w995_,
		_w996_,
		_w997_
	);
	LUT4 #(
		.INIT('hb000)
	) name740 (
		_w706_,
		_w712_,
		_w715_,
		_w719_,
		_w998_
	);
	LUT4 #(
		.INIT('hb000)
	) name741 (
		_w711_,
		_w719_,
		_w722_,
		_w724_,
		_w999_
	);
	LUT4 #(
		.INIT('hb000)
	) name742 (
		_w717_,
		_w724_,
		_w727_,
		_w731_,
		_w1000_
	);
	LUT4 #(
		.INIT('h4f00)
	) name743 (
		_w997_,
		_w998_,
		_w999_,
		_w1000_,
		_w1001_
	);
	LUT4 #(
		.INIT('hb000)
	) name744 (
		_w723_,
		_w731_,
		_w733_,
		_w735_,
		_w1002_
	);
	LUT4 #(
		.INIT('hb000)
	) name745 (
		_w729_,
		_w735_,
		_w739_,
		_w743_,
		_w1003_
	);
	LUT4 #(
		.INIT('hb000)
	) name746 (
		_w734_,
		_w743_,
		_w745_,
		_w747_,
		_w1004_
	);
	LUT4 #(
		.INIT('h4f00)
	) name747 (
		_w1001_,
		_w1002_,
		_w1003_,
		_w1004_,
		_w1005_
	);
	LUT4 #(
		.INIT('hb000)
	) name748 (
		_w741_,
		_w747_,
		_w750_,
		_w752_,
		_w1006_
	);
	LUT4 #(
		.INIT('h8088)
	) name749 (
		_w264_,
		_w590_,
		_w746_,
		_w752_,
		_w1007_
	);
	LUT4 #(
		.INIT('hc400)
	) name750 (
		_w264_,
		_w267_,
		_w882_,
		_w970_,
		_w1008_
	);
	LUT4 #(
		.INIT('h4f00)
	) name751 (
		_w1005_,
		_w1006_,
		_w1007_,
		_w1008_,
		_w1009_
	);
	LUT2 #(
		.INIT('he)
	) name752 (
		_w971_,
		_w1009_,
		_w1010_
	);
	LUT3 #(
		.INIT('hb0)
	) name753 (
		\priority[9] ,
		\req[8] ,
		\req[9] ,
		_w1011_
	);
	LUT2 #(
		.INIT('h4)
	) name754 (
		_w429_,
		_w1011_,
		_w1012_
	);
	LUT3 #(
		.INIT('h31)
	) name755 (
		\priority[10] ,
		\priority[11] ,
		\req[10] ,
		_w1013_
	);
	LUT4 #(
		.INIT('hc040)
	) name756 (
		_w268_,
		_w274_,
		_w275_,
		_w1013_,
		_w1014_
	);
	LUT4 #(
		.INIT('h30b0)
	) name757 (
		_w283_,
		_w288_,
		_w295_,
		_w1014_,
		_w1015_
	);
	LUT4 #(
		.INIT('h30b0)
	) name758 (
		_w299_,
		_w307_,
		_w311_,
		_w1015_,
		_w1016_
	);
	LUT4 #(
		.INIT('h30b0)
	) name759 (
		_w318_,
		_w323_,
		_w330_,
		_w1016_,
		_w1017_
	);
	LUT4 #(
		.INIT('h30b0)
	) name760 (
		_w334_,
		_w342_,
		_w346_,
		_w1017_,
		_w1018_
	);
	LUT4 #(
		.INIT('h30b0)
	) name761 (
		_w353_,
		_w358_,
		_w365_,
		_w1018_,
		_w1019_
	);
	LUT4 #(
		.INIT('h30b0)
	) name762 (
		_w369_,
		_w377_,
		_w381_,
		_w1019_,
		_w1020_
	);
	LUT4 #(
		.INIT('h30b0)
	) name763 (
		_w388_,
		_w393_,
		_w400_,
		_w1020_,
		_w1021_
	);
	LUT4 #(
		.INIT('h30b0)
	) name764 (
		_w404_,
		_w412_,
		_w416_,
		_w1021_,
		_w1022_
	);
	LUT4 #(
		.INIT('hd000)
	) name765 (
		_w414_,
		_w418_,
		_w420_,
		_w796_,
		_w1023_
	);
	LUT4 #(
		.INIT('h80c0)
	) name766 (
		_w258_,
		_w430_,
		_w756_,
		_w796_,
		_w1024_
	);
	LUT4 #(
		.INIT('hc400)
	) name767 (
		_w430_,
		_w433_,
		_w924_,
		_w1011_,
		_w1025_
	);
	LUT4 #(
		.INIT('h4f00)
	) name768 (
		_w1022_,
		_w1023_,
		_w1024_,
		_w1025_,
		_w1026_
	);
	LUT2 #(
		.INIT('he)
	) name769 (
		_w1012_,
		_w1026_,
		_w1027_
	);
	LUT3 #(
		.INIT('hb0)
	) name770 (
		\priority[10] ,
		\req[9] ,
		\req[10] ,
		_w1028_
	);
	LUT2 #(
		.INIT('h4)
	) name771 (
		_w595_,
		_w1028_,
		_w1029_
	);
	LUT3 #(
		.INIT('h31)
	) name772 (
		\priority[11] ,
		\priority[12] ,
		\req[11] ,
		_w1030_
	);
	LUT4 #(
		.INIT('hc040)
	) name773 (
		_w434_,
		_w440_,
		_w441_,
		_w1030_,
		_w1031_
	);
	LUT4 #(
		.INIT('h30b0)
	) name774 (
		_w449_,
		_w454_,
		_w461_,
		_w1031_,
		_w1032_
	);
	LUT4 #(
		.INIT('h30b0)
	) name775 (
		_w465_,
		_w473_,
		_w477_,
		_w1032_,
		_w1033_
	);
	LUT4 #(
		.INIT('h30b0)
	) name776 (
		_w484_,
		_w489_,
		_w496_,
		_w1033_,
		_w1034_
	);
	LUT4 #(
		.INIT('h3b00)
	) name777 (
		_w500_,
		_w508_,
		_w1034_,
		_w512_,
		_w1035_
	);
	LUT4 #(
		.INIT('h30b0)
	) name778 (
		_w519_,
		_w524_,
		_w531_,
		_w1035_,
		_w1036_
	);
	LUT4 #(
		.INIT('h30b0)
	) name779 (
		_w535_,
		_w543_,
		_w547_,
		_w1036_,
		_w1037_
	);
	LUT4 #(
		.INIT('h30b0)
	) name780 (
		_w554_,
		_w559_,
		_w566_,
		_w1037_,
		_w1038_
	);
	LUT4 #(
		.INIT('h30b0)
	) name781 (
		_w570_,
		_w578_,
		_w582_,
		_w1038_,
		_w1039_
	);
	LUT4 #(
		.INIT('hd000)
	) name782 (
		_w580_,
		_w584_,
		_w586_,
		_w840_,
		_w1040_
	);
	LUT4 #(
		.INIT('h80c0)
	) name783 (
		_w424_,
		_w596_,
		_w800_,
		_w840_,
		_w1041_
	);
	LUT4 #(
		.INIT('hc400)
	) name784 (
		_w596_,
		_w599_,
		_w966_,
		_w1028_,
		_w1042_
	);
	LUT4 #(
		.INIT('h4f00)
	) name785 (
		_w1039_,
		_w1040_,
		_w1041_,
		_w1042_,
		_w1043_
	);
	LUT2 #(
		.INIT('he)
	) name786 (
		_w1029_,
		_w1043_,
		_w1044_
	);
	LUT3 #(
		.INIT('hb0)
	) name787 (
		\priority[11] ,
		\req[10] ,
		\req[11] ,
		_w1045_
	);
	LUT2 #(
		.INIT('h4)
	) name788 (
		_w273_,
		_w1045_,
		_w1046_
	);
	LUT3 #(
		.INIT('h31)
	) name789 (
		\priority[12] ,
		\priority[13] ,
		\req[12] ,
		_w1047_
	);
	LUT4 #(
		.INIT('hc040)
	) name790 (
		_w600_,
		_w606_,
		_w607_,
		_w1047_,
		_w1048_
	);
	LUT4 #(
		.INIT('h30b0)
	) name791 (
		_w615_,
		_w620_,
		_w627_,
		_w1048_,
		_w1049_
	);
	LUT4 #(
		.INIT('h30b0)
	) name792 (
		_w631_,
		_w639_,
		_w643_,
		_w1049_,
		_w1050_
	);
	LUT4 #(
		.INIT('h30b0)
	) name793 (
		_w650_,
		_w655_,
		_w662_,
		_w1050_,
		_w1051_
	);
	LUT4 #(
		.INIT('h30b0)
	) name794 (
		_w666_,
		_w674_,
		_w678_,
		_w1051_,
		_w1052_
	);
	LUT4 #(
		.INIT('h30b0)
	) name795 (
		_w685_,
		_w690_,
		_w697_,
		_w1052_,
		_w1053_
	);
	LUT4 #(
		.INIT('h30b0)
	) name796 (
		_w701_,
		_w709_,
		_w713_,
		_w1053_,
		_w1054_
	);
	LUT4 #(
		.INIT('h30b0)
	) name797 (
		_w720_,
		_w725_,
		_w732_,
		_w1054_,
		_w1055_
	);
	LUT4 #(
		.INIT('h30b0)
	) name798 (
		_w736_,
		_w744_,
		_w748_,
		_w1055_,
		_w1056_
	);
	LUT4 #(
		.INIT('hd000)
	) name799 (
		_w746_,
		_w750_,
		_w752_,
		_w882_,
		_w1057_
	);
	LUT4 #(
		.INIT('h8088)
	) name800 (
		_w263_,
		_w264_,
		_w590_,
		_w882_,
		_w1058_
	);
	LUT4 #(
		.INIT('hd000)
	) name801 (
		_w263_,
		_w267_,
		_w271_,
		_w1045_,
		_w1059_
	);
	LUT4 #(
		.INIT('h4f00)
	) name802 (
		_w1056_,
		_w1057_,
		_w1058_,
		_w1059_,
		_w1060_
	);
	LUT2 #(
		.INIT('he)
	) name803 (
		_w1046_,
		_w1060_,
		_w1061_
	);
	LUT3 #(
		.INIT('hb0)
	) name804 (
		\priority[12] ,
		\req[11] ,
		\req[12] ,
		_w1062_
	);
	LUT2 #(
		.INIT('h4)
	) name805 (
		_w439_,
		_w1062_,
		_w1063_
	);
	LUT3 #(
		.INIT('h31)
	) name806 (
		\priority[13] ,
		\priority[14] ,
		\req[13] ,
		_w1064_
	);
	LUT4 #(
		.INIT('ha020)
	) name807 (
		_w274_,
		_w277_,
		_w285_,
		_w1064_,
		_w1065_
	);
	LUT4 #(
		.INIT('h30b0)
	) name808 (
		_w763_,
		_w765_,
		_w766_,
		_w1065_,
		_w1066_
	);
	LUT4 #(
		.INIT('h30b0)
	) name809 (
		_w767_,
		_w769_,
		_w770_,
		_w1066_,
		_w1067_
	);
	LUT4 #(
		.INIT('h30b0)
	) name810 (
		_w771_,
		_w773_,
		_w774_,
		_w1067_,
		_w1068_
	);
	LUT4 #(
		.INIT('h30b0)
	) name811 (
		_w775_,
		_w777_,
		_w778_,
		_w1068_,
		_w1069_
	);
	LUT4 #(
		.INIT('h30b0)
	) name812 (
		_w779_,
		_w781_,
		_w782_,
		_w1069_,
		_w1070_
	);
	LUT4 #(
		.INIT('h30b0)
	) name813 (
		_w783_,
		_w785_,
		_w786_,
		_w1070_,
		_w1071_
	);
	LUT4 #(
		.INIT('h30b0)
	) name814 (
		_w787_,
		_w789_,
		_w790_,
		_w1071_,
		_w1072_
	);
	LUT4 #(
		.INIT('h30b0)
	) name815 (
		_w791_,
		_w793_,
		_w794_,
		_w1072_,
		_w1073_
	);
	LUT4 #(
		.INIT('hd000)
	) name816 (
		_w258_,
		_w420_,
		_w796_,
		_w924_,
		_w1074_
	);
	LUT4 #(
		.INIT('h8088)
	) name817 (
		_w429_,
		_w430_,
		_w756_,
		_w924_,
		_w1075_
	);
	LUT4 #(
		.INIT('hd000)
	) name818 (
		_w429_,
		_w433_,
		_w437_,
		_w1062_,
		_w1076_
	);
	LUT4 #(
		.INIT('h4f00)
	) name819 (
		_w1073_,
		_w1074_,
		_w1075_,
		_w1076_,
		_w1077_
	);
	LUT2 #(
		.INIT('he)
	) name820 (
		_w1063_,
		_w1077_,
		_w1078_
	);
	LUT3 #(
		.INIT('hb0)
	) name821 (
		\priority[13] ,
		\req[12] ,
		\req[13] ,
		_w1079_
	);
	LUT2 #(
		.INIT('h4)
	) name822 (
		_w605_,
		_w1079_,
		_w1080_
	);
	LUT3 #(
		.INIT('h31)
	) name823 (
		\priority[14] ,
		\priority[15] ,
		\req[14] ,
		_w1081_
	);
	LUT4 #(
		.INIT('ha020)
	) name824 (
		_w440_,
		_w443_,
		_w451_,
		_w1081_,
		_w1082_
	);
	LUT4 #(
		.INIT('h30b0)
	) name825 (
		_w807_,
		_w809_,
		_w810_,
		_w1082_,
		_w1083_
	);
	LUT4 #(
		.INIT('h4c44)
	) name826 (
		_w813_,
		_w814_,
		_w1083_,
		_w811_,
		_w1084_
	);
	LUT4 #(
		.INIT('h30b0)
	) name827 (
		_w815_,
		_w817_,
		_w818_,
		_w1084_,
		_w1085_
	);
	LUT4 #(
		.INIT('h30b0)
	) name828 (
		_w819_,
		_w821_,
		_w822_,
		_w1085_,
		_w1086_
	);
	LUT4 #(
		.INIT('h30b0)
	) name829 (
		_w823_,
		_w825_,
		_w826_,
		_w1086_,
		_w1087_
	);
	LUT4 #(
		.INIT('h30b0)
	) name830 (
		_w827_,
		_w829_,
		_w830_,
		_w1087_,
		_w1088_
	);
	LUT4 #(
		.INIT('h30b0)
	) name831 (
		_w831_,
		_w833_,
		_w834_,
		_w1088_,
		_w1089_
	);
	LUT4 #(
		.INIT('h30b0)
	) name832 (
		_w835_,
		_w837_,
		_w838_,
		_w1089_,
		_w1090_
	);
	LUT4 #(
		.INIT('hd000)
	) name833 (
		_w424_,
		_w586_,
		_w840_,
		_w966_,
		_w1091_
	);
	LUT4 #(
		.INIT('h8088)
	) name834 (
		_w595_,
		_w596_,
		_w800_,
		_w966_,
		_w1092_
	);
	LUT4 #(
		.INIT('hd000)
	) name835 (
		_w595_,
		_w599_,
		_w603_,
		_w1079_,
		_w1093_
	);
	LUT4 #(
		.INIT('h4f00)
	) name836 (
		_w1090_,
		_w1091_,
		_w1092_,
		_w1093_,
		_w1094_
	);
	LUT2 #(
		.INIT('he)
	) name837 (
		_w1080_,
		_w1094_,
		_w1095_
	);
	LUT3 #(
		.INIT('hb0)
	) name838 (
		\priority[14] ,
		\req[13] ,
		\req[14] ,
		_w1096_
	);
	LUT2 #(
		.INIT('h4)
	) name839 (
		_w275_,
		_w1096_,
		_w1097_
	);
	LUT3 #(
		.INIT('h31)
	) name840 (
		\priority[15] ,
		\priority[16] ,
		\req[15] ,
		_w1098_
	);
	LUT4 #(
		.INIT('ha020)
	) name841 (
		_w606_,
		_w609_,
		_w617_,
		_w1098_,
		_w1099_
	);
	LUT4 #(
		.INIT('h30b0)
	) name842 (
		_w850_,
		_w852_,
		_w853_,
		_w1099_,
		_w1100_
	);
	LUT4 #(
		.INIT('h30b0)
	) name843 (
		_w854_,
		_w856_,
		_w857_,
		_w1100_,
		_w1101_
	);
	LUT4 #(
		.INIT('h30b0)
	) name844 (
		_w858_,
		_w860_,
		_w861_,
		_w1101_,
		_w1102_
	);
	LUT4 #(
		.INIT('h30b0)
	) name845 (
		_w862_,
		_w864_,
		_w865_,
		_w1102_,
		_w1103_
	);
	LUT4 #(
		.INIT('h30b0)
	) name846 (
		_w866_,
		_w868_,
		_w869_,
		_w1103_,
		_w1104_
	);
	LUT4 #(
		.INIT('h30b0)
	) name847 (
		_w870_,
		_w872_,
		_w873_,
		_w1104_,
		_w1105_
	);
	LUT4 #(
		.INIT('h30b0)
	) name848 (
		_w874_,
		_w876_,
		_w877_,
		_w1105_,
		_w1106_
	);
	LUT4 #(
		.INIT('h30b0)
	) name849 (
		_w878_,
		_w880_,
		_w881_,
		_w1106_,
		_w1107_
	);
	LUT4 #(
		.INIT('ha200)
	) name850 (
		_w267_,
		_w590_,
		_w752_,
		_w882_,
		_w1108_
	);
	LUT4 #(
		.INIT('h8a00)
	) name851 (
		_w263_,
		_w264_,
		_w267_,
		_w273_,
		_w1109_
	);
	LUT4 #(
		.INIT('h8a00)
	) name852 (
		_w269_,
		_w271_,
		_w273_,
		_w1096_,
		_w1110_
	);
	LUT4 #(
		.INIT('h4f00)
	) name853 (
		_w1107_,
		_w1108_,
		_w1109_,
		_w1110_,
		_w1111_
	);
	LUT2 #(
		.INIT('he)
	) name854 (
		_w1097_,
		_w1111_,
		_w1112_
	);
	LUT3 #(
		.INIT('hb0)
	) name855 (
		\priority[15] ,
		\req[14] ,
		\req[15] ,
		_w1113_
	);
	LUT2 #(
		.INIT('h4)
	) name856 (
		_w441_,
		_w1113_,
		_w1114_
	);
	LUT3 #(
		.INIT('h31)
	) name857 (
		\priority[16] ,
		\priority[17] ,
		\req[16] ,
		_w1115_
	);
	LUT4 #(
		.INIT('hc040)
	) name858 (
		_w281_,
		_w285_,
		_w287_,
		_w1115_,
		_w1116_
	);
	LUT4 #(
		.INIT('h30b0)
	) name859 (
		_w892_,
		_w894_,
		_w895_,
		_w1116_,
		_w1117_
	);
	LUT4 #(
		.INIT('h30b0)
	) name860 (
		_w896_,
		_w898_,
		_w899_,
		_w1117_,
		_w1118_
	);
	LUT4 #(
		.INIT('h30b0)
	) name861 (
		_w900_,
		_w902_,
		_w903_,
		_w1118_,
		_w1119_
	);
	LUT4 #(
		.INIT('h30b0)
	) name862 (
		_w904_,
		_w906_,
		_w907_,
		_w1119_,
		_w1120_
	);
	LUT4 #(
		.INIT('h30b0)
	) name863 (
		_w908_,
		_w910_,
		_w911_,
		_w1120_,
		_w1121_
	);
	LUT4 #(
		.INIT('h30b0)
	) name864 (
		_w912_,
		_w914_,
		_w915_,
		_w1121_,
		_w1122_
	);
	LUT4 #(
		.INIT('h30b0)
	) name865 (
		_w916_,
		_w918_,
		_w919_,
		_w1122_,
		_w1123_
	);
	LUT4 #(
		.INIT('h30b0)
	) name866 (
		_w920_,
		_w922_,
		_w923_,
		_w1123_,
		_w1124_
	);
	LUT4 #(
		.INIT('ha200)
	) name867 (
		_w433_,
		_w756_,
		_w796_,
		_w924_,
		_w1125_
	);
	LUT4 #(
		.INIT('h8a00)
	) name868 (
		_w429_,
		_w430_,
		_w433_,
		_w439_,
		_w1126_
	);
	LUT4 #(
		.INIT('h8a00)
	) name869 (
		_w435_,
		_w437_,
		_w439_,
		_w1113_,
		_w1127_
	);
	LUT4 #(
		.INIT('h4f00)
	) name870 (
		_w1124_,
		_w1125_,
		_w1126_,
		_w1127_,
		_w1128_
	);
	LUT2 #(
		.INIT('he)
	) name871 (
		_w1114_,
		_w1128_,
		_w1129_
	);
	LUT3 #(
		.INIT('hb0)
	) name872 (
		\priority[16] ,
		\req[15] ,
		\req[16] ,
		_w1130_
	);
	LUT2 #(
		.INIT('h4)
	) name873 (
		_w607_,
		_w1130_,
		_w1131_
	);
	LUT3 #(
		.INIT('h31)
	) name874 (
		\priority[17] ,
		\priority[18] ,
		\req[17] ,
		_w1132_
	);
	LUT4 #(
		.INIT('hc040)
	) name875 (
		_w447_,
		_w451_,
		_w453_,
		_w1132_,
		_w1133_
	);
	LUT4 #(
		.INIT('h30b0)
	) name876 (
		_w934_,
		_w936_,
		_w937_,
		_w1133_,
		_w1134_
	);
	LUT4 #(
		.INIT('h30b0)
	) name877 (
		_w938_,
		_w940_,
		_w941_,
		_w1134_,
		_w1135_
	);
	LUT4 #(
		.INIT('h30b0)
	) name878 (
		_w942_,
		_w944_,
		_w945_,
		_w1135_,
		_w1136_
	);
	LUT4 #(
		.INIT('h30b0)
	) name879 (
		_w946_,
		_w948_,
		_w949_,
		_w1136_,
		_w1137_
	);
	LUT4 #(
		.INIT('h30b0)
	) name880 (
		_w950_,
		_w952_,
		_w953_,
		_w1137_,
		_w1138_
	);
	LUT4 #(
		.INIT('h30b0)
	) name881 (
		_w954_,
		_w956_,
		_w957_,
		_w1138_,
		_w1139_
	);
	LUT4 #(
		.INIT('h30b0)
	) name882 (
		_w958_,
		_w960_,
		_w961_,
		_w1139_,
		_w1140_
	);
	LUT4 #(
		.INIT('h30b0)
	) name883 (
		_w962_,
		_w964_,
		_w965_,
		_w1140_,
		_w1141_
	);
	LUT4 #(
		.INIT('ha200)
	) name884 (
		_w599_,
		_w800_,
		_w840_,
		_w966_,
		_w1142_
	);
	LUT4 #(
		.INIT('h8a00)
	) name885 (
		_w595_,
		_w596_,
		_w599_,
		_w605_,
		_w1143_
	);
	LUT4 #(
		.INIT('h8a00)
	) name886 (
		_w601_,
		_w603_,
		_w605_,
		_w1130_,
		_w1144_
	);
	LUT4 #(
		.INIT('h4f00)
	) name887 (
		_w1141_,
		_w1142_,
		_w1143_,
		_w1144_,
		_w1145_
	);
	LUT2 #(
		.INIT('he)
	) name888 (
		_w1131_,
		_w1145_,
		_w1146_
	);
	LUT3 #(
		.INIT('hb0)
	) name889 (
		\priority[17] ,
		\req[16] ,
		\req[17] ,
		_w1147_
	);
	LUT2 #(
		.INIT('h4)
	) name890 (
		_w274_,
		_w1147_,
		_w1148_
	);
	LUT3 #(
		.INIT('h31)
	) name891 (
		\priority[18] ,
		\priority[19] ,
		\req[18] ,
		_w1149_
	);
	LUT4 #(
		.INIT('hc040)
	) name892 (
		_w613_,
		_w617_,
		_w619_,
		_w1149_,
		_w1150_
	);
	LUT4 #(
		.INIT('h30b0)
	) name893 (
		_w976_,
		_w978_,
		_w979_,
		_w1150_,
		_w1151_
	);
	LUT4 #(
		.INIT('h30b0)
	) name894 (
		_w980_,
		_w982_,
		_w983_,
		_w1151_,
		_w1152_
	);
	LUT4 #(
		.INIT('h30b0)
	) name895 (
		_w984_,
		_w986_,
		_w987_,
		_w1152_,
		_w1153_
	);
	LUT4 #(
		.INIT('h30b0)
	) name896 (
		_w988_,
		_w990_,
		_w991_,
		_w1153_,
		_w1154_
	);
	LUT4 #(
		.INIT('h30b0)
	) name897 (
		_w992_,
		_w994_,
		_w995_,
		_w1154_,
		_w1155_
	);
	LUT4 #(
		.INIT('h30b0)
	) name898 (
		_w996_,
		_w998_,
		_w999_,
		_w1155_,
		_w1156_
	);
	LUT4 #(
		.INIT('h30b0)
	) name899 (
		_w1000_,
		_w1002_,
		_w1003_,
		_w1156_,
		_w1157_
	);
	LUT4 #(
		.INIT('h30b0)
	) name900 (
		_w1004_,
		_w1006_,
		_w1007_,
		_w1157_,
		_w1158_
	);
	LUT4 #(
		.INIT('hc040)
	) name901 (
		_w264_,
		_w267_,
		_w271_,
		_w882_,
		_w1159_
	);
	LUT4 #(
		.INIT('hb000)
	) name902 (
		_w263_,
		_w271_,
		_w273_,
		_w275_,
		_w1160_
	);
	LUT4 #(
		.INIT('hb000)
	) name903 (
		_w269_,
		_w275_,
		_w278_,
		_w1147_,
		_w1161_
	);
	LUT4 #(
		.INIT('h4f00)
	) name904 (
		_w1158_,
		_w1159_,
		_w1160_,
		_w1161_,
		_w1162_
	);
	LUT2 #(
		.INIT('he)
	) name905 (
		_w1148_,
		_w1162_,
		_w1163_
	);
	LUT3 #(
		.INIT('hb0)
	) name906 (
		\priority[18] ,
		\req[17] ,
		\req[18] ,
		_w1164_
	);
	LUT2 #(
		.INIT('h4)
	) name907 (
		_w440_,
		_w1164_,
		_w1165_
	);
	LUT3 #(
		.INIT('h31)
	) name908 (
		\priority[19] ,
		\priority[20] ,
		\req[19] ,
		_w1166_
	);
	LUT4 #(
		.INIT('hc040)
	) name909 (
		_w279_,
		_w286_,
		_w287_,
		_w1166_,
		_w1167_
	);
	LUT4 #(
		.INIT('h30b0)
	) name910 (
		_w295_,
		_w299_,
		_w307_,
		_w1167_,
		_w1168_
	);
	LUT4 #(
		.INIT('h30b0)
	) name911 (
		_w311_,
		_w318_,
		_w323_,
		_w1168_,
		_w1169_
	);
	LUT4 #(
		.INIT('h30b0)
	) name912 (
		_w330_,
		_w334_,
		_w342_,
		_w1169_,
		_w1170_
	);
	LUT4 #(
		.INIT('h30b0)
	) name913 (
		_w346_,
		_w353_,
		_w358_,
		_w1170_,
		_w1171_
	);
	LUT4 #(
		.INIT('h30b0)
	) name914 (
		_w365_,
		_w369_,
		_w377_,
		_w1171_,
		_w1172_
	);
	LUT4 #(
		.INIT('h30b0)
	) name915 (
		_w381_,
		_w388_,
		_w393_,
		_w1172_,
		_w1173_
	);
	LUT4 #(
		.INIT('h30b0)
	) name916 (
		_w400_,
		_w404_,
		_w412_,
		_w1173_,
		_w1174_
	);
	LUT4 #(
		.INIT('h30b0)
	) name917 (
		_w416_,
		_w1023_,
		_w1024_,
		_w1174_,
		_w1175_
	);
	LUT4 #(
		.INIT('hc040)
	) name918 (
		_w430_,
		_w433_,
		_w437_,
		_w924_,
		_w1176_
	);
	LUT4 #(
		.INIT('hb000)
	) name919 (
		_w429_,
		_w437_,
		_w439_,
		_w441_,
		_w1177_
	);
	LUT4 #(
		.INIT('hb000)
	) name920 (
		_w435_,
		_w441_,
		_w444_,
		_w1164_,
		_w1178_
	);
	LUT4 #(
		.INIT('h4f00)
	) name921 (
		_w1175_,
		_w1176_,
		_w1177_,
		_w1178_,
		_w1179_
	);
	LUT2 #(
		.INIT('he)
	) name922 (
		_w1165_,
		_w1179_,
		_w1180_
	);
	LUT3 #(
		.INIT('hb0)
	) name923 (
		\priority[19] ,
		\req[18] ,
		\req[19] ,
		_w1181_
	);
	LUT2 #(
		.INIT('h4)
	) name924 (
		_w606_,
		_w1181_,
		_w1182_
	);
	LUT3 #(
		.INIT('h31)
	) name925 (
		\priority[20] ,
		\priority[21] ,
		\req[20] ,
		_w1183_
	);
	LUT4 #(
		.INIT('hc040)
	) name926 (
		_w445_,
		_w452_,
		_w453_,
		_w1183_,
		_w1184_
	);
	LUT4 #(
		.INIT('h30b0)
	) name927 (
		_w461_,
		_w465_,
		_w473_,
		_w1184_,
		_w1185_
	);
	LUT4 #(
		.INIT('h08cc)
	) name928 (
		_w477_,
		_w489_,
		_w1185_,
		_w484_,
		_w1186_
	);
	LUT4 #(
		.INIT('h30b0)
	) name929 (
		_w496_,
		_w500_,
		_w508_,
		_w1186_,
		_w1187_
	);
	LUT4 #(
		.INIT('h44c4)
	) name930 (
		_w519_,
		_w524_,
		_w512_,
		_w1187_,
		_w1188_
	);
	LUT4 #(
		.INIT('h30b0)
	) name931 (
		_w531_,
		_w535_,
		_w543_,
		_w1188_,
		_w1189_
	);
	LUT4 #(
		.INIT('h30b0)
	) name932 (
		_w547_,
		_w554_,
		_w559_,
		_w1189_,
		_w1190_
	);
	LUT4 #(
		.INIT('h30b0)
	) name933 (
		_w566_,
		_w570_,
		_w578_,
		_w1190_,
		_w1191_
	);
	LUT4 #(
		.INIT('h30b0)
	) name934 (
		_w582_,
		_w1040_,
		_w1041_,
		_w1191_,
		_w1192_
	);
	LUT4 #(
		.INIT('hc040)
	) name935 (
		_w596_,
		_w599_,
		_w603_,
		_w966_,
		_w1193_
	);
	LUT4 #(
		.INIT('hb000)
	) name936 (
		_w595_,
		_w603_,
		_w605_,
		_w607_,
		_w1194_
	);
	LUT4 #(
		.INIT('hb000)
	) name937 (
		_w601_,
		_w607_,
		_w610_,
		_w1181_,
		_w1195_
	);
	LUT4 #(
		.INIT('h4f00)
	) name938 (
		_w1192_,
		_w1193_,
		_w1194_,
		_w1195_,
		_w1196_
	);
	LUT2 #(
		.INIT('he)
	) name939 (
		_w1182_,
		_w1196_,
		_w1197_
	);
	LUT3 #(
		.INIT('hb0)
	) name940 (
		\priority[20] ,
		\req[19] ,
		\req[20] ,
		_w1198_
	);
	LUT2 #(
		.INIT('h4)
	) name941 (
		_w285_,
		_w1198_,
		_w1199_
	);
	LUT3 #(
		.INIT('h31)
	) name942 (
		\priority[21] ,
		\priority[22] ,
		\req[21] ,
		_w1200_
	);
	LUT4 #(
		.INIT('hc040)
	) name943 (
		_w611_,
		_w618_,
		_w619_,
		_w1200_,
		_w1201_
	);
	LUT4 #(
		.INIT('h30b0)
	) name944 (
		_w627_,
		_w631_,
		_w639_,
		_w1201_,
		_w1202_
	);
	LUT4 #(
		.INIT('h30b0)
	) name945 (
		_w643_,
		_w650_,
		_w655_,
		_w1202_,
		_w1203_
	);
	LUT4 #(
		.INIT('h30b0)
	) name946 (
		_w662_,
		_w666_,
		_w674_,
		_w1203_,
		_w1204_
	);
	LUT4 #(
		.INIT('h30b0)
	) name947 (
		_w678_,
		_w685_,
		_w690_,
		_w1204_,
		_w1205_
	);
	LUT4 #(
		.INIT('h30b0)
	) name948 (
		_w697_,
		_w701_,
		_w709_,
		_w1205_,
		_w1206_
	);
	LUT4 #(
		.INIT('h30b0)
	) name949 (
		_w713_,
		_w720_,
		_w725_,
		_w1206_,
		_w1207_
	);
	LUT4 #(
		.INIT('h30b0)
	) name950 (
		_w732_,
		_w736_,
		_w744_,
		_w1207_,
		_w1208_
	);
	LUT4 #(
		.INIT('h30b0)
	) name951 (
		_w748_,
		_w1057_,
		_w1058_,
		_w1208_,
		_w1209_
	);
	LUT4 #(
		.INIT('hd000)
	) name952 (
		_w274_,
		_w278_,
		_w282_,
		_w1198_,
		_w1210_
	);
	LUT4 #(
		.INIT('h3b00)
	) name953 (
		_w272_,
		_w276_,
		_w1209_,
		_w1210_,
		_w1211_
	);
	LUT2 #(
		.INIT('he)
	) name954 (
		_w1199_,
		_w1211_,
		_w1212_
	);
	LUT3 #(
		.INIT('hb0)
	) name955 (
		\priority[21] ,
		\req[20] ,
		\req[21] ,
		_w1213_
	);
	LUT2 #(
		.INIT('h4)
	) name956 (
		_w451_,
		_w1213_,
		_w1214_
	);
	LUT3 #(
		.INIT('h31)
	) name957 (
		\priority[22] ,
		\priority[23] ,
		\req[22] ,
		_w1215_
	);
	LUT4 #(
		.INIT('ha020)
	) name958 (
		_w286_,
		_w289_,
		_w296_,
		_w1215_,
		_w1216_
	);
	LUT4 #(
		.INIT('h30b0)
	) name959 (
		_w766_,
		_w767_,
		_w769_,
		_w1216_,
		_w1217_
	);
	LUT4 #(
		.INIT('h30b0)
	) name960 (
		_w770_,
		_w771_,
		_w773_,
		_w1217_,
		_w1218_
	);
	LUT4 #(
		.INIT('h30b0)
	) name961 (
		_w774_,
		_w775_,
		_w777_,
		_w1218_,
		_w1219_
	);
	LUT4 #(
		.INIT('h30b0)
	) name962 (
		_w778_,
		_w779_,
		_w781_,
		_w1219_,
		_w1220_
	);
	LUT4 #(
		.INIT('h30b0)
	) name963 (
		_w782_,
		_w783_,
		_w785_,
		_w1220_,
		_w1221_
	);
	LUT4 #(
		.INIT('h30b0)
	) name964 (
		_w786_,
		_w787_,
		_w789_,
		_w1221_,
		_w1222_
	);
	LUT4 #(
		.INIT('h30b0)
	) name965 (
		_w790_,
		_w791_,
		_w793_,
		_w1222_,
		_w1223_
	);
	LUT4 #(
		.INIT('h30b0)
	) name966 (
		_w794_,
		_w1074_,
		_w1075_,
		_w1223_,
		_w1224_
	);
	LUT4 #(
		.INIT('hd000)
	) name967 (
		_w440_,
		_w444_,
		_w448_,
		_w1213_,
		_w1225_
	);
	LUT4 #(
		.INIT('h3b00)
	) name968 (
		_w438_,
		_w442_,
		_w1224_,
		_w1225_,
		_w1226_
	);
	LUT2 #(
		.INIT('he)
	) name969 (
		_w1214_,
		_w1226_,
		_w1227_
	);
	LUT3 #(
		.INIT('hb0)
	) name970 (
		\priority[22] ,
		\req[21] ,
		\req[22] ,
		_w1228_
	);
	LUT2 #(
		.INIT('h4)
	) name971 (
		_w617_,
		_w1228_,
		_w1229_
	);
	LUT3 #(
		.INIT('h31)
	) name972 (
		\priority[23] ,
		\priority[24] ,
		\req[23] ,
		_w1230_
	);
	LUT4 #(
		.INIT('ha020)
	) name973 (
		_w452_,
		_w455_,
		_w462_,
		_w1230_,
		_w1231_
	);
	LUT4 #(
		.INIT('h0c8c)
	) name974 (
		_w810_,
		_w813_,
		_w811_,
		_w1231_,
		_w1232_
	);
	LUT4 #(
		.INIT('h30b0)
	) name975 (
		_w814_,
		_w815_,
		_w817_,
		_w1232_,
		_w1233_
	);
	LUT4 #(
		.INIT('h30b0)
	) name976 (
		_w818_,
		_w819_,
		_w821_,
		_w1233_,
		_w1234_
	);
	LUT4 #(
		.INIT('h30b0)
	) name977 (
		_w822_,
		_w823_,
		_w825_,
		_w1234_,
		_w1235_
	);
	LUT4 #(
		.INIT('h30b0)
	) name978 (
		_w826_,
		_w827_,
		_w829_,
		_w1235_,
		_w1236_
	);
	LUT4 #(
		.INIT('h30b0)
	) name979 (
		_w830_,
		_w831_,
		_w833_,
		_w1236_,
		_w1237_
	);
	LUT4 #(
		.INIT('h30b0)
	) name980 (
		_w834_,
		_w835_,
		_w837_,
		_w1237_,
		_w1238_
	);
	LUT4 #(
		.INIT('h30b0)
	) name981 (
		_w838_,
		_w1091_,
		_w1092_,
		_w1238_,
		_w1239_
	);
	LUT4 #(
		.INIT('hd000)
	) name982 (
		_w606_,
		_w610_,
		_w614_,
		_w1228_,
		_w1240_
	);
	LUT4 #(
		.INIT('h3b00)
	) name983 (
		_w604_,
		_w608_,
		_w1239_,
		_w1240_,
		_w1241_
	);
	LUT2 #(
		.INIT('he)
	) name984 (
		_w1229_,
		_w1241_,
		_w1242_
	);
	LUT3 #(
		.INIT('hb0)
	) name985 (
		\priority[23] ,
		\req[22] ,
		\req[23] ,
		_w1243_
	);
	LUT2 #(
		.INIT('h4)
	) name986 (
		_w287_,
		_w1243_,
		_w1244_
	);
	LUT3 #(
		.INIT('h31)
	) name987 (
		\priority[24] ,
		\priority[25] ,
		\req[24] ,
		_w1245_
	);
	LUT4 #(
		.INIT('ha020)
	) name988 (
		_w618_,
		_w621_,
		_w628_,
		_w1245_,
		_w1246_
	);
	LUT4 #(
		.INIT('h30b0)
	) name989 (
		_w853_,
		_w854_,
		_w856_,
		_w1246_,
		_w1247_
	);
	LUT4 #(
		.INIT('h30b0)
	) name990 (
		_w857_,
		_w858_,
		_w860_,
		_w1247_,
		_w1248_
	);
	LUT4 #(
		.INIT('h30b0)
	) name991 (
		_w861_,
		_w862_,
		_w864_,
		_w1248_,
		_w1249_
	);
	LUT4 #(
		.INIT('h30b0)
	) name992 (
		_w865_,
		_w866_,
		_w868_,
		_w1249_,
		_w1250_
	);
	LUT4 #(
		.INIT('h30b0)
	) name993 (
		_w869_,
		_w870_,
		_w872_,
		_w1250_,
		_w1251_
	);
	LUT4 #(
		.INIT('h30b0)
	) name994 (
		_w873_,
		_w874_,
		_w876_,
		_w1251_,
		_w1252_
	);
	LUT4 #(
		.INIT('h30b0)
	) name995 (
		_w877_,
		_w878_,
		_w880_,
		_w1252_,
		_w1253_
	);
	LUT4 #(
		.INIT('h30b0)
	) name996 (
		_w881_,
		_w1108_,
		_w1109_,
		_w1253_,
		_w1254_
	);
	LUT4 #(
		.INIT('h8a00)
	) name997 (
		_w280_,
		_w282_,
		_w285_,
		_w1243_,
		_w1255_
	);
	LUT4 #(
		.INIT('h3b00)
	) name998 (
		_w761_,
		_w762_,
		_w1254_,
		_w1255_,
		_w1256_
	);
	LUT2 #(
		.INIT('he)
	) name999 (
		_w1244_,
		_w1256_,
		_w1257_
	);
	LUT3 #(
		.INIT('hb0)
	) name1000 (
		\priority[24] ,
		\req[23] ,
		\req[24] ,
		_w1258_
	);
	LUT2 #(
		.INIT('h4)
	) name1001 (
		_w453_,
		_w1258_,
		_w1259_
	);
	LUT3 #(
		.INIT('h31)
	) name1002 (
		\priority[25] ,
		\priority[26] ,
		\req[25] ,
		_w1260_
	);
	LUT4 #(
		.INIT('hc040)
	) name1003 (
		_w293_,
		_w296_,
		_w298_,
		_w1260_,
		_w1261_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1004 (
		_w895_,
		_w896_,
		_w898_,
		_w1261_,
		_w1262_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1005 (
		_w899_,
		_w900_,
		_w902_,
		_w1262_,
		_w1263_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1006 (
		_w903_,
		_w904_,
		_w906_,
		_w1263_,
		_w1264_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1007 (
		_w907_,
		_w908_,
		_w910_,
		_w1264_,
		_w1265_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1008 (
		_w911_,
		_w912_,
		_w914_,
		_w1265_,
		_w1266_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1009 (
		_w915_,
		_w916_,
		_w918_,
		_w1266_,
		_w1267_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1010 (
		_w919_,
		_w920_,
		_w922_,
		_w1267_,
		_w1268_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1011 (
		_w923_,
		_w1125_,
		_w1126_,
		_w1268_,
		_w1269_
	);
	LUT4 #(
		.INIT('h8a00)
	) name1012 (
		_w446_,
		_w448_,
		_w451_,
		_w1258_,
		_w1270_
	);
	LUT4 #(
		.INIT('h3b00)
	) name1013 (
		_w805_,
		_w806_,
		_w1269_,
		_w1270_,
		_w1271_
	);
	LUT2 #(
		.INIT('he)
	) name1014 (
		_w1259_,
		_w1271_,
		_w1272_
	);
	LUT3 #(
		.INIT('hb0)
	) name1015 (
		\priority[25] ,
		\req[24] ,
		\req[25] ,
		_w1273_
	);
	LUT2 #(
		.INIT('h4)
	) name1016 (
		_w619_,
		_w1273_,
		_w1274_
	);
	LUT3 #(
		.INIT('h31)
	) name1017 (
		\priority[26] ,
		\priority[27] ,
		\req[26] ,
		_w1275_
	);
	LUT4 #(
		.INIT('hc040)
	) name1018 (
		_w459_,
		_w462_,
		_w464_,
		_w1275_,
		_w1276_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1019 (
		_w937_,
		_w938_,
		_w940_,
		_w1276_,
		_w1277_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1020 (
		_w941_,
		_w942_,
		_w944_,
		_w1277_,
		_w1278_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1021 (
		_w945_,
		_w946_,
		_w948_,
		_w1278_,
		_w1279_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1022 (
		_w949_,
		_w950_,
		_w952_,
		_w1279_,
		_w1280_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1023 (
		_w953_,
		_w954_,
		_w956_,
		_w1280_,
		_w1281_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1024 (
		_w957_,
		_w958_,
		_w960_,
		_w1281_,
		_w1282_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1025 (
		_w961_,
		_w962_,
		_w964_,
		_w1282_,
		_w1283_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1026 (
		_w965_,
		_w1142_,
		_w1143_,
		_w1283_,
		_w1284_
	);
	LUT4 #(
		.INIT('h8a00)
	) name1027 (
		_w612_,
		_w614_,
		_w617_,
		_w1273_,
		_w1285_
	);
	LUT4 #(
		.INIT('h3b00)
	) name1028 (
		_w848_,
		_w849_,
		_w1284_,
		_w1285_,
		_w1286_
	);
	LUT2 #(
		.INIT('he)
	) name1029 (
		_w1274_,
		_w1286_,
		_w1287_
	);
	LUT3 #(
		.INIT('hb0)
	) name1030 (
		\priority[26] ,
		\req[25] ,
		\req[26] ,
		_w1288_
	);
	LUT2 #(
		.INIT('h4)
	) name1031 (
		_w286_,
		_w1288_,
		_w1289_
	);
	LUT3 #(
		.INIT('h31)
	) name1032 (
		\priority[27] ,
		\priority[28] ,
		\req[27] ,
		_w1290_
	);
	LUT4 #(
		.INIT('hc040)
	) name1033 (
		_w625_,
		_w628_,
		_w630_,
		_w1290_,
		_w1291_
	);
	LUT4 #(
		.INIT('h3b00)
	) name1034 (
		_w979_,
		_w980_,
		_w1291_,
		_w982_,
		_w1292_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1035 (
		_w983_,
		_w984_,
		_w986_,
		_w1292_,
		_w1293_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1036 (
		_w987_,
		_w988_,
		_w990_,
		_w1293_,
		_w1294_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1037 (
		_w991_,
		_w992_,
		_w994_,
		_w1294_,
		_w1295_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1038 (
		_w995_,
		_w996_,
		_w998_,
		_w1295_,
		_w1296_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1039 (
		_w999_,
		_w1000_,
		_w1002_,
		_w1296_,
		_w1297_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1040 (
		_w1003_,
		_w1004_,
		_w1006_,
		_w1297_,
		_w1298_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1041 (
		_w1007_,
		_w1159_,
		_w1160_,
		_w1298_,
		_w1299_
	);
	LUT4 #(
		.INIT('hb000)
	) name1042 (
		_w280_,
		_w287_,
		_w290_,
		_w1288_,
		_w1300_
	);
	LUT4 #(
		.INIT('h3b00)
	) name1043 (
		_w890_,
		_w891_,
		_w1299_,
		_w1300_,
		_w1301_
	);
	LUT2 #(
		.INIT('he)
	) name1044 (
		_w1289_,
		_w1301_,
		_w1302_
	);
	LUT3 #(
		.INIT('hb0)
	) name1045 (
		\priority[27] ,
		\req[26] ,
		\req[27] ,
		_w1303_
	);
	LUT2 #(
		.INIT('h4)
	) name1046 (
		_w452_,
		_w1303_,
		_w1304_
	);
	LUT3 #(
		.INIT('h31)
	) name1047 (
		\priority[28] ,
		\priority[29] ,
		\req[28] ,
		_w1305_
	);
	LUT4 #(
		.INIT('hc040)
	) name1048 (
		_w291_,
		_w297_,
		_w298_,
		_w1305_,
		_w1306_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1049 (
		_w307_,
		_w311_,
		_w318_,
		_w1306_,
		_w1307_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1050 (
		_w323_,
		_w330_,
		_w334_,
		_w1307_,
		_w1308_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1051 (
		_w342_,
		_w346_,
		_w353_,
		_w1308_,
		_w1309_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1052 (
		_w358_,
		_w365_,
		_w369_,
		_w1309_,
		_w1310_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1053 (
		_w377_,
		_w381_,
		_w388_,
		_w1310_,
		_w1311_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1054 (
		_w393_,
		_w400_,
		_w404_,
		_w1311_,
		_w1312_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1055 (
		_w412_,
		_w416_,
		_w1023_,
		_w1312_,
		_w1313_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1056 (
		_w1024_,
		_w1176_,
		_w1177_,
		_w1313_,
		_w1314_
	);
	LUT4 #(
		.INIT('hb000)
	) name1057 (
		_w446_,
		_w453_,
		_w456_,
		_w1303_,
		_w1315_
	);
	LUT4 #(
		.INIT('h3b00)
	) name1058 (
		_w932_,
		_w933_,
		_w1314_,
		_w1315_,
		_w1316_
	);
	LUT2 #(
		.INIT('he)
	) name1059 (
		_w1304_,
		_w1316_,
		_w1317_
	);
	LUT3 #(
		.INIT('hb0)
	) name1060 (
		\priority[28] ,
		\req[27] ,
		\req[28] ,
		_w1318_
	);
	LUT2 #(
		.INIT('h4)
	) name1061 (
		_w618_,
		_w1318_,
		_w1319_
	);
	LUT3 #(
		.INIT('h31)
	) name1062 (
		\priority[29] ,
		\priority[30] ,
		\req[29] ,
		_w1320_
	);
	LUT4 #(
		.INIT('hc040)
	) name1063 (
		_w457_,
		_w463_,
		_w464_,
		_w1320_,
		_w1321_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1064 (
		_w473_,
		_w477_,
		_w484_,
		_w1321_,
		_w1322_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1065 (
		_w489_,
		_w496_,
		_w500_,
		_w1322_,
		_w1323_
	);
	LUT4 #(
		.INIT('h0c8c)
	) name1066 (
		_w508_,
		_w519_,
		_w512_,
		_w1323_,
		_w1324_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1067 (
		_w524_,
		_w531_,
		_w535_,
		_w1324_,
		_w1325_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1068 (
		_w543_,
		_w547_,
		_w554_,
		_w1325_,
		_w1326_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1069 (
		_w559_,
		_w566_,
		_w570_,
		_w1326_,
		_w1327_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1070 (
		_w578_,
		_w582_,
		_w1040_,
		_w1327_,
		_w1328_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1071 (
		_w1041_,
		_w1193_,
		_w1194_,
		_w1328_,
		_w1329_
	);
	LUT4 #(
		.INIT('hb000)
	) name1072 (
		_w612_,
		_w619_,
		_w622_,
		_w1318_,
		_w1330_
	);
	LUT4 #(
		.INIT('h3b00)
	) name1073 (
		_w974_,
		_w975_,
		_w1329_,
		_w1330_,
		_w1331_
	);
	LUT2 #(
		.INIT('he)
	) name1074 (
		_w1319_,
		_w1331_,
		_w1332_
	);
	LUT3 #(
		.INIT('hb0)
	) name1075 (
		\priority[29] ,
		\req[28] ,
		\req[29] ,
		_w1333_
	);
	LUT2 #(
		.INIT('h4)
	) name1076 (
		_w296_,
		_w1333_,
		_w1334_
	);
	LUT3 #(
		.INIT('h31)
	) name1077 (
		\priority[30] ,
		\priority[31] ,
		\req[30] ,
		_w1335_
	);
	LUT4 #(
		.INIT('hc040)
	) name1078 (
		_w623_,
		_w629_,
		_w630_,
		_w1335_,
		_w1336_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1079 (
		_w639_,
		_w643_,
		_w650_,
		_w1336_,
		_w1337_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1080 (
		_w655_,
		_w662_,
		_w666_,
		_w1337_,
		_w1338_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1081 (
		_w674_,
		_w678_,
		_w685_,
		_w1338_,
		_w1339_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1082 (
		_w690_,
		_w697_,
		_w701_,
		_w1339_,
		_w1340_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1083 (
		_w709_,
		_w713_,
		_w720_,
		_w1340_,
		_w1341_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1084 (
		_w725_,
		_w732_,
		_w736_,
		_w1341_,
		_w1342_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1085 (
		_w744_,
		_w748_,
		_w1057_,
		_w1342_,
		_w1343_
	);
	LUT4 #(
		.INIT('h44c4)
	) name1086 (
		_w272_,
		_w276_,
		_w1058_,
		_w1343_,
		_w1344_
	);
	LUT4 #(
		.INIT('hd000)
	) name1087 (
		_w286_,
		_w290_,
		_w294_,
		_w1333_,
		_w1345_
	);
	LUT4 #(
		.INIT('h3b00)
	) name1088 (
		_w283_,
		_w288_,
		_w1344_,
		_w1345_,
		_w1346_
	);
	LUT2 #(
		.INIT('he)
	) name1089 (
		_w1334_,
		_w1346_,
		_w1347_
	);
	LUT3 #(
		.INIT('hb0)
	) name1090 (
		\priority[30] ,
		\req[29] ,
		\req[30] ,
		_w1348_
	);
	LUT2 #(
		.INIT('h4)
	) name1091 (
		_w462_,
		_w1348_,
		_w1349_
	);
	LUT3 #(
		.INIT('h31)
	) name1092 (
		\priority[31] ,
		\priority[32] ,
		\req[31] ,
		_w1350_
	);
	LUT4 #(
		.INIT('ha020)
	) name1093 (
		_w297_,
		_w301_,
		_w308_,
		_w1350_,
		_w1351_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1094 (
		_w769_,
		_w770_,
		_w771_,
		_w1351_,
		_w1352_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1095 (
		_w773_,
		_w774_,
		_w775_,
		_w1352_,
		_w1353_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1096 (
		_w777_,
		_w778_,
		_w779_,
		_w1353_,
		_w1354_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1097 (
		_w781_,
		_w782_,
		_w783_,
		_w1354_,
		_w1355_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1098 (
		_w785_,
		_w786_,
		_w787_,
		_w1355_,
		_w1356_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1099 (
		_w789_,
		_w790_,
		_w791_,
		_w1356_,
		_w1357_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1100 (
		_w793_,
		_w794_,
		_w1074_,
		_w1357_,
		_w1358_
	);
	LUT4 #(
		.INIT('h44c4)
	) name1101 (
		_w438_,
		_w442_,
		_w1075_,
		_w1358_,
		_w1359_
	);
	LUT4 #(
		.INIT('hd000)
	) name1102 (
		_w452_,
		_w456_,
		_w460_,
		_w1348_,
		_w1360_
	);
	LUT4 #(
		.INIT('h3b00)
	) name1103 (
		_w449_,
		_w454_,
		_w1359_,
		_w1360_,
		_w1361_
	);
	LUT2 #(
		.INIT('he)
	) name1104 (
		_w1349_,
		_w1361_,
		_w1362_
	);
	LUT3 #(
		.INIT('hb0)
	) name1105 (
		\priority[31] ,
		\req[30] ,
		\req[31] ,
		_w1363_
	);
	LUT2 #(
		.INIT('h4)
	) name1106 (
		_w628_,
		_w1363_,
		_w1364_
	);
	LUT3 #(
		.INIT('h31)
	) name1107 (
		\priority[32] ,
		\priority[33] ,
		\req[32] ,
		_w1365_
	);
	LUT4 #(
		.INIT('ha020)
	) name1108 (
		_w463_,
		_w467_,
		_w474_,
		_w1365_,
		_w1366_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1109 (
		_w813_,
		_w814_,
		_w815_,
		_w1366_,
		_w1367_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1110 (
		_w817_,
		_w818_,
		_w819_,
		_w1367_,
		_w1368_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1111 (
		_w821_,
		_w822_,
		_w823_,
		_w1368_,
		_w1369_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1112 (
		_w825_,
		_w826_,
		_w827_,
		_w1369_,
		_w1370_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1113 (
		_w829_,
		_w830_,
		_w831_,
		_w1370_,
		_w1371_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1114 (
		_w833_,
		_w834_,
		_w835_,
		_w1371_,
		_w1372_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1115 (
		_w837_,
		_w838_,
		_w1091_,
		_w1372_,
		_w1373_
	);
	LUT4 #(
		.INIT('h44c4)
	) name1116 (
		_w604_,
		_w608_,
		_w1092_,
		_w1373_,
		_w1374_
	);
	LUT4 #(
		.INIT('hd000)
	) name1117 (
		_w618_,
		_w622_,
		_w626_,
		_w1363_,
		_w1375_
	);
	LUT4 #(
		.INIT('h3b00)
	) name1118 (
		_w615_,
		_w620_,
		_w1374_,
		_w1375_,
		_w1376_
	);
	LUT2 #(
		.INIT('he)
	) name1119 (
		_w1364_,
		_w1376_,
		_w1377_
	);
	LUT3 #(
		.INIT('hb0)
	) name1120 (
		\priority[32] ,
		\req[31] ,
		\req[32] ,
		_w1378_
	);
	LUT2 #(
		.INIT('h4)
	) name1121 (
		_w298_,
		_w1378_,
		_w1379_
	);
	LUT3 #(
		.INIT('h31)
	) name1122 (
		\priority[33] ,
		\priority[34] ,
		\req[33] ,
		_w1380_
	);
	LUT4 #(
		.INIT('ha020)
	) name1123 (
		_w629_,
		_w633_,
		_w640_,
		_w1380_,
		_w1381_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1124 (
		_w856_,
		_w857_,
		_w858_,
		_w1381_,
		_w1382_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1125 (
		_w860_,
		_w861_,
		_w862_,
		_w1382_,
		_w1383_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1126 (
		_w864_,
		_w865_,
		_w866_,
		_w1383_,
		_w1384_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1127 (
		_w868_,
		_w869_,
		_w870_,
		_w1384_,
		_w1385_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1128 (
		_w872_,
		_w873_,
		_w874_,
		_w1385_,
		_w1386_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1129 (
		_w876_,
		_w877_,
		_w878_,
		_w1386_,
		_w1387_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1130 (
		_w880_,
		_w881_,
		_w1108_,
		_w1387_,
		_w1388_
	);
	LUT4 #(
		.INIT('h44c4)
	) name1131 (
		_w761_,
		_w762_,
		_w1109_,
		_w1388_,
		_w1389_
	);
	LUT4 #(
		.INIT('h8a00)
	) name1132 (
		_w292_,
		_w294_,
		_w296_,
		_w1378_,
		_w1390_
	);
	LUT4 #(
		.INIT('h3b00)
	) name1133 (
		_w763_,
		_w765_,
		_w1389_,
		_w1390_,
		_w1391_
	);
	LUT2 #(
		.INIT('he)
	) name1134 (
		_w1379_,
		_w1391_,
		_w1392_
	);
	LUT3 #(
		.INIT('hb0)
	) name1135 (
		\priority[33] ,
		\req[32] ,
		\req[33] ,
		_w1393_
	);
	LUT2 #(
		.INIT('h4)
	) name1136 (
		_w464_,
		_w1393_,
		_w1394_
	);
	LUT3 #(
		.INIT('h31)
	) name1137 (
		\priority[34] ,
		\priority[35] ,
		\req[34] ,
		_w1395_
	);
	LUT4 #(
		.INIT('hc040)
	) name1138 (
		_w305_,
		_w308_,
		_w310_,
		_w1395_,
		_w1396_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1139 (
		_w898_,
		_w899_,
		_w900_,
		_w1396_,
		_w1397_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1140 (
		_w902_,
		_w903_,
		_w904_,
		_w1397_,
		_w1398_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1141 (
		_w906_,
		_w907_,
		_w908_,
		_w1398_,
		_w1399_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1142 (
		_w910_,
		_w911_,
		_w912_,
		_w1399_,
		_w1400_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1143 (
		_w914_,
		_w915_,
		_w916_,
		_w1400_,
		_w1401_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1144 (
		_w918_,
		_w919_,
		_w920_,
		_w1401_,
		_w1402_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1145 (
		_w922_,
		_w923_,
		_w1125_,
		_w1402_,
		_w1403_
	);
	LUT4 #(
		.INIT('h44c4)
	) name1146 (
		_w805_,
		_w806_,
		_w1126_,
		_w1403_,
		_w1404_
	);
	LUT4 #(
		.INIT('h8a00)
	) name1147 (
		_w458_,
		_w460_,
		_w462_,
		_w1393_,
		_w1405_
	);
	LUT4 #(
		.INIT('h3b00)
	) name1148 (
		_w807_,
		_w809_,
		_w1404_,
		_w1405_,
		_w1406_
	);
	LUT2 #(
		.INIT('he)
	) name1149 (
		_w1394_,
		_w1406_,
		_w1407_
	);
	LUT3 #(
		.INIT('hb0)
	) name1150 (
		\priority[34] ,
		\req[33] ,
		\req[34] ,
		_w1408_
	);
	LUT2 #(
		.INIT('h4)
	) name1151 (
		_w630_,
		_w1408_,
		_w1409_
	);
	LUT3 #(
		.INIT('h31)
	) name1152 (
		\priority[35] ,
		\priority[36] ,
		\req[35] ,
		_w1410_
	);
	LUT4 #(
		.INIT('hc040)
	) name1153 (
		_w471_,
		_w474_,
		_w476_,
		_w1410_,
		_w1411_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1154 (
		_w940_,
		_w941_,
		_w942_,
		_w1411_,
		_w1412_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1155 (
		_w944_,
		_w945_,
		_w946_,
		_w1412_,
		_w1413_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1156 (
		_w948_,
		_w949_,
		_w950_,
		_w1413_,
		_w1414_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1157 (
		_w952_,
		_w953_,
		_w954_,
		_w1414_,
		_w1415_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1158 (
		_w956_,
		_w957_,
		_w958_,
		_w1415_,
		_w1416_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1159 (
		_w960_,
		_w961_,
		_w962_,
		_w1416_,
		_w1417_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1160 (
		_w964_,
		_w965_,
		_w1142_,
		_w1417_,
		_w1418_
	);
	LUT4 #(
		.INIT('h44c4)
	) name1161 (
		_w848_,
		_w849_,
		_w1143_,
		_w1418_,
		_w1419_
	);
	LUT4 #(
		.INIT('h8a00)
	) name1162 (
		_w624_,
		_w626_,
		_w628_,
		_w1408_,
		_w1420_
	);
	LUT4 #(
		.INIT('h3b00)
	) name1163 (
		_w850_,
		_w852_,
		_w1419_,
		_w1420_,
		_w1421_
	);
	LUT2 #(
		.INIT('he)
	) name1164 (
		_w1409_,
		_w1421_,
		_w1422_
	);
	LUT3 #(
		.INIT('hb0)
	) name1165 (
		\priority[35] ,
		\req[34] ,
		\req[35] ,
		_w1423_
	);
	LUT2 #(
		.INIT('h4)
	) name1166 (
		_w297_,
		_w1423_,
		_w1424_
	);
	LUT3 #(
		.INIT('h31)
	) name1167 (
		\priority[36] ,
		\priority[37] ,
		\req[36] ,
		_w1425_
	);
	LUT4 #(
		.INIT('hc040)
	) name1168 (
		_w637_,
		_w640_,
		_w642_,
		_w1425_,
		_w1426_
	);
	LUT4 #(
		.INIT('h44c4)
	) name1169 (
		_w983_,
		_w984_,
		_w982_,
		_w1426_,
		_w1427_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1170 (
		_w986_,
		_w987_,
		_w988_,
		_w1427_,
		_w1428_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1171 (
		_w990_,
		_w991_,
		_w992_,
		_w1428_,
		_w1429_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1172 (
		_w994_,
		_w995_,
		_w996_,
		_w1429_,
		_w1430_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1173 (
		_w998_,
		_w999_,
		_w1000_,
		_w1430_,
		_w1431_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1174 (
		_w1002_,
		_w1003_,
		_w1004_,
		_w1431_,
		_w1432_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1175 (
		_w1006_,
		_w1007_,
		_w1159_,
		_w1432_,
		_w1433_
	);
	LUT4 #(
		.INIT('h44c4)
	) name1176 (
		_w890_,
		_w891_,
		_w1160_,
		_w1433_,
		_w1434_
	);
	LUT4 #(
		.INIT('hb000)
	) name1177 (
		_w292_,
		_w298_,
		_w302_,
		_w1423_,
		_w1435_
	);
	LUT4 #(
		.INIT('h3b00)
	) name1178 (
		_w892_,
		_w894_,
		_w1434_,
		_w1435_,
		_w1436_
	);
	LUT2 #(
		.INIT('he)
	) name1179 (
		_w1424_,
		_w1436_,
		_w1437_
	);
	LUT3 #(
		.INIT('hb0)
	) name1180 (
		\priority[36] ,
		\req[35] ,
		\req[36] ,
		_w1438_
	);
	LUT2 #(
		.INIT('h4)
	) name1181 (
		_w463_,
		_w1438_,
		_w1439_
	);
	LUT3 #(
		.INIT('h31)
	) name1182 (
		\priority[37] ,
		\priority[38] ,
		\req[37] ,
		_w1440_
	);
	LUT4 #(
		.INIT('hc040)
	) name1183 (
		_w303_,
		_w309_,
		_w310_,
		_w1440_,
		_w1441_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1184 (
		_w318_,
		_w323_,
		_w330_,
		_w1441_,
		_w1442_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1185 (
		_w334_,
		_w342_,
		_w346_,
		_w1442_,
		_w1443_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1186 (
		_w353_,
		_w358_,
		_w365_,
		_w1443_,
		_w1444_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1187 (
		_w369_,
		_w377_,
		_w381_,
		_w1444_,
		_w1445_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1188 (
		_w388_,
		_w393_,
		_w400_,
		_w1445_,
		_w1446_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1189 (
		_w404_,
		_w412_,
		_w416_,
		_w1446_,
		_w1447_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1190 (
		_w1023_,
		_w1024_,
		_w1176_,
		_w1447_,
		_w1448_
	);
	LUT4 #(
		.INIT('h44c4)
	) name1191 (
		_w932_,
		_w933_,
		_w1177_,
		_w1448_,
		_w1449_
	);
	LUT4 #(
		.INIT('hb000)
	) name1192 (
		_w458_,
		_w464_,
		_w468_,
		_w1438_,
		_w1450_
	);
	LUT4 #(
		.INIT('h3b00)
	) name1193 (
		_w934_,
		_w936_,
		_w1449_,
		_w1450_,
		_w1451_
	);
	LUT2 #(
		.INIT('he)
	) name1194 (
		_w1439_,
		_w1451_,
		_w1452_
	);
	LUT3 #(
		.INIT('hb0)
	) name1195 (
		\priority[37] ,
		\req[36] ,
		\req[37] ,
		_w1453_
	);
	LUT2 #(
		.INIT('h4)
	) name1196 (
		_w629_,
		_w1453_,
		_w1454_
	);
	LUT3 #(
		.INIT('h31)
	) name1197 (
		\priority[38] ,
		\priority[39] ,
		\req[38] ,
		_w1455_
	);
	LUT4 #(
		.INIT('hc040)
	) name1198 (
		_w469_,
		_w475_,
		_w476_,
		_w1455_,
		_w1456_
	);
	LUT4 #(
		.INIT('h5d00)
	) name1199 (
		_w489_,
		_w484_,
		_w1456_,
		_w496_,
		_w1457_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1200 (
		_w500_,
		_w508_,
		_w512_,
		_w1457_,
		_w1458_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1201 (
		_w519_,
		_w524_,
		_w531_,
		_w1458_,
		_w1459_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1202 (
		_w535_,
		_w543_,
		_w547_,
		_w1459_,
		_w1460_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1203 (
		_w554_,
		_w559_,
		_w566_,
		_w1460_,
		_w1461_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1204 (
		_w570_,
		_w578_,
		_w582_,
		_w1461_,
		_w1462_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1205 (
		_w1040_,
		_w1041_,
		_w1193_,
		_w1462_,
		_w1463_
	);
	LUT4 #(
		.INIT('h44c4)
	) name1206 (
		_w974_,
		_w975_,
		_w1194_,
		_w1463_,
		_w1464_
	);
	LUT4 #(
		.INIT('hb000)
	) name1207 (
		_w624_,
		_w630_,
		_w634_,
		_w1453_,
		_w1465_
	);
	LUT4 #(
		.INIT('h3b00)
	) name1208 (
		_w976_,
		_w978_,
		_w1464_,
		_w1465_,
		_w1466_
	);
	LUT2 #(
		.INIT('he)
	) name1209 (
		_w1454_,
		_w1466_,
		_w1467_
	);
	LUT3 #(
		.INIT('hb0)
	) name1210 (
		\priority[38] ,
		\req[37] ,
		\req[38] ,
		_w1468_
	);
	LUT2 #(
		.INIT('h4)
	) name1211 (
		_w308_,
		_w1468_,
		_w1469_
	);
	LUT3 #(
		.INIT('h31)
	) name1212 (
		\priority[39] ,
		\priority[40] ,
		\req[39] ,
		_w1470_
	);
	LUT4 #(
		.INIT('hc040)
	) name1213 (
		_w635_,
		_w641_,
		_w642_,
		_w1470_,
		_w1471_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1214 (
		_w650_,
		_w655_,
		_w662_,
		_w1471_,
		_w1472_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1215 (
		_w666_,
		_w674_,
		_w678_,
		_w1472_,
		_w1473_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1216 (
		_w685_,
		_w690_,
		_w697_,
		_w1473_,
		_w1474_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1217 (
		_w701_,
		_w709_,
		_w713_,
		_w1474_,
		_w1475_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1218 (
		_w720_,
		_w725_,
		_w732_,
		_w1475_,
		_w1476_
	);
	LUT4 #(
		.INIT('h4c44)
	) name1219 (
		_w744_,
		_w748_,
		_w1476_,
		_w736_,
		_w1477_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name1220 (
		_w272_,
		_w1057_,
		_w1058_,
		_w1477_,
		_w1478_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1221 (
		_w276_,
		_w283_,
		_w288_,
		_w1478_,
		_w1479_
	);
	LUT4 #(
		.INIT('hd000)
	) name1222 (
		_w297_,
		_w302_,
		_w306_,
		_w1468_,
		_w1480_
	);
	LUT4 #(
		.INIT('h3b00)
	) name1223 (
		_w295_,
		_w299_,
		_w1479_,
		_w1480_,
		_w1481_
	);
	LUT2 #(
		.INIT('he)
	) name1224 (
		_w1469_,
		_w1481_,
		_w1482_
	);
	LUT3 #(
		.INIT('hb0)
	) name1225 (
		\priority[39] ,
		\req[38] ,
		\req[39] ,
		_w1483_
	);
	LUT2 #(
		.INIT('h4)
	) name1226 (
		_w474_,
		_w1483_,
		_w1484_
	);
	LUT3 #(
		.INIT('h31)
	) name1227 (
		\priority[40] ,
		\priority[41] ,
		\req[40] ,
		_w1485_
	);
	LUT4 #(
		.INIT('ha020)
	) name1228 (
		_w309_,
		_w312_,
		_w320_,
		_w1485_,
		_w1486_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1229 (
		_w771_,
		_w773_,
		_w774_,
		_w1486_,
		_w1487_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1230 (
		_w775_,
		_w777_,
		_w778_,
		_w1487_,
		_w1488_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1231 (
		_w779_,
		_w781_,
		_w782_,
		_w1488_,
		_w1489_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1232 (
		_w783_,
		_w785_,
		_w786_,
		_w1489_,
		_w1490_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1233 (
		_w787_,
		_w789_,
		_w790_,
		_w1490_,
		_w1491_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1234 (
		_w791_,
		_w793_,
		_w794_,
		_w1491_,
		_w1492_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name1235 (
		_w438_,
		_w1074_,
		_w1075_,
		_w1492_,
		_w1493_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1236 (
		_w442_,
		_w449_,
		_w454_,
		_w1493_,
		_w1494_
	);
	LUT4 #(
		.INIT('hd000)
	) name1237 (
		_w463_,
		_w468_,
		_w472_,
		_w1483_,
		_w1495_
	);
	LUT4 #(
		.INIT('h3b00)
	) name1238 (
		_w461_,
		_w465_,
		_w1494_,
		_w1495_,
		_w1496_
	);
	LUT2 #(
		.INIT('he)
	) name1239 (
		_w1484_,
		_w1496_,
		_w1497_
	);
	LUT3 #(
		.INIT('hb0)
	) name1240 (
		\priority[40] ,
		\req[39] ,
		\req[40] ,
		_w1498_
	);
	LUT2 #(
		.INIT('h4)
	) name1241 (
		_w640_,
		_w1498_,
		_w1499_
	);
	LUT3 #(
		.INIT('h31)
	) name1242 (
		\priority[41] ,
		\priority[42] ,
		\req[41] ,
		_w1500_
	);
	LUT4 #(
		.INIT('ha020)
	) name1243 (
		_w475_,
		_w478_,
		_w486_,
		_w1500_,
		_w1501_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1244 (
		_w815_,
		_w817_,
		_w818_,
		_w1501_,
		_w1502_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1245 (
		_w819_,
		_w821_,
		_w822_,
		_w1502_,
		_w1503_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1246 (
		_w823_,
		_w825_,
		_w826_,
		_w1503_,
		_w1504_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1247 (
		_w827_,
		_w829_,
		_w830_,
		_w1504_,
		_w1505_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1248 (
		_w831_,
		_w833_,
		_w834_,
		_w1505_,
		_w1506_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1249 (
		_w835_,
		_w837_,
		_w838_,
		_w1506_,
		_w1507_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name1250 (
		_w604_,
		_w1091_,
		_w1092_,
		_w1507_,
		_w1508_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1251 (
		_w608_,
		_w615_,
		_w620_,
		_w1508_,
		_w1509_
	);
	LUT4 #(
		.INIT('hd000)
	) name1252 (
		_w629_,
		_w634_,
		_w638_,
		_w1498_,
		_w1510_
	);
	LUT4 #(
		.INIT('h3b00)
	) name1253 (
		_w627_,
		_w631_,
		_w1509_,
		_w1510_,
		_w1511_
	);
	LUT2 #(
		.INIT('he)
	) name1254 (
		_w1499_,
		_w1511_,
		_w1512_
	);
	LUT3 #(
		.INIT('hb0)
	) name1255 (
		\priority[41] ,
		\req[40] ,
		\req[41] ,
		_w1513_
	);
	LUT2 #(
		.INIT('h4)
	) name1256 (
		_w310_,
		_w1513_,
		_w1514_
	);
	LUT3 #(
		.INIT('h31)
	) name1257 (
		\priority[42] ,
		\priority[43] ,
		\req[42] ,
		_w1515_
	);
	LUT4 #(
		.INIT('ha020)
	) name1258 (
		_w641_,
		_w644_,
		_w652_,
		_w1515_,
		_w1516_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1259 (
		_w858_,
		_w860_,
		_w861_,
		_w1516_,
		_w1517_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1260 (
		_w862_,
		_w864_,
		_w865_,
		_w1517_,
		_w1518_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1261 (
		_w866_,
		_w868_,
		_w869_,
		_w1518_,
		_w1519_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1262 (
		_w870_,
		_w872_,
		_w873_,
		_w1519_,
		_w1520_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1263 (
		_w874_,
		_w876_,
		_w877_,
		_w1520_,
		_w1521_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1264 (
		_w878_,
		_w880_,
		_w881_,
		_w1521_,
		_w1522_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name1265 (
		_w761_,
		_w1108_,
		_w1109_,
		_w1522_,
		_w1523_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1266 (
		_w762_,
		_w763_,
		_w765_,
		_w1523_,
		_w1524_
	);
	LUT4 #(
		.INIT('h8a00)
	) name1267 (
		_w304_,
		_w306_,
		_w308_,
		_w1513_,
		_w1525_
	);
	LUT4 #(
		.INIT('h3b00)
	) name1268 (
		_w766_,
		_w767_,
		_w1524_,
		_w1525_,
		_w1526_
	);
	LUT2 #(
		.INIT('he)
	) name1269 (
		_w1514_,
		_w1526_,
		_w1527_
	);
	LUT3 #(
		.INIT('hb0)
	) name1270 (
		\priority[42] ,
		\req[41] ,
		\req[42] ,
		_w1528_
	);
	LUT2 #(
		.INIT('h4)
	) name1271 (
		_w476_,
		_w1528_,
		_w1529_
	);
	LUT3 #(
		.INIT('h31)
	) name1272 (
		\priority[43] ,
		\priority[44] ,
		\req[43] ,
		_w1530_
	);
	LUT4 #(
		.INIT('hc040)
	) name1273 (
		_w316_,
		_w320_,
		_w322_,
		_w1530_,
		_w1531_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1274 (
		_w900_,
		_w902_,
		_w903_,
		_w1531_,
		_w1532_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1275 (
		_w904_,
		_w906_,
		_w907_,
		_w1532_,
		_w1533_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1276 (
		_w908_,
		_w910_,
		_w911_,
		_w1533_,
		_w1534_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1277 (
		_w912_,
		_w914_,
		_w915_,
		_w1534_,
		_w1535_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1278 (
		_w916_,
		_w918_,
		_w919_,
		_w1535_,
		_w1536_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1279 (
		_w920_,
		_w922_,
		_w923_,
		_w1536_,
		_w1537_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name1280 (
		_w805_,
		_w1125_,
		_w1126_,
		_w1537_,
		_w1538_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1281 (
		_w806_,
		_w807_,
		_w809_,
		_w1538_,
		_w1539_
	);
	LUT4 #(
		.INIT('h8a00)
	) name1282 (
		_w470_,
		_w472_,
		_w474_,
		_w1528_,
		_w1540_
	);
	LUT4 #(
		.INIT('h3b00)
	) name1283 (
		_w810_,
		_w811_,
		_w1539_,
		_w1540_,
		_w1541_
	);
	LUT2 #(
		.INIT('he)
	) name1284 (
		_w1529_,
		_w1541_,
		_w1542_
	);
	LUT3 #(
		.INIT('hb0)
	) name1285 (
		\priority[43] ,
		\req[42] ,
		\req[43] ,
		_w1543_
	);
	LUT2 #(
		.INIT('h4)
	) name1286 (
		_w642_,
		_w1543_,
		_w1544_
	);
	LUT3 #(
		.INIT('h31)
	) name1287 (
		\priority[44] ,
		\priority[45] ,
		\req[44] ,
		_w1545_
	);
	LUT4 #(
		.INIT('hc040)
	) name1288 (
		_w482_,
		_w486_,
		_w488_,
		_w1545_,
		_w1546_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1289 (
		_w942_,
		_w944_,
		_w945_,
		_w1546_,
		_w1547_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1290 (
		_w946_,
		_w948_,
		_w949_,
		_w1547_,
		_w1548_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1291 (
		_w950_,
		_w952_,
		_w953_,
		_w1548_,
		_w1549_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1292 (
		_w954_,
		_w956_,
		_w957_,
		_w1549_,
		_w1550_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1293 (
		_w958_,
		_w960_,
		_w961_,
		_w1550_,
		_w1551_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1294 (
		_w962_,
		_w964_,
		_w965_,
		_w1551_,
		_w1552_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name1295 (
		_w848_,
		_w1142_,
		_w1143_,
		_w1552_,
		_w1553_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1296 (
		_w849_,
		_w850_,
		_w852_,
		_w1553_,
		_w1554_
	);
	LUT4 #(
		.INIT('h8a00)
	) name1297 (
		_w636_,
		_w638_,
		_w640_,
		_w1543_,
		_w1555_
	);
	LUT4 #(
		.INIT('h3b00)
	) name1298 (
		_w853_,
		_w854_,
		_w1554_,
		_w1555_,
		_w1556_
	);
	LUT2 #(
		.INIT('he)
	) name1299 (
		_w1544_,
		_w1556_,
		_w1557_
	);
	LUT3 #(
		.INIT('hb0)
	) name1300 (
		\priority[44] ,
		\req[43] ,
		\req[44] ,
		_w1558_
	);
	LUT2 #(
		.INIT('h4)
	) name1301 (
		_w309_,
		_w1558_,
		_w1559_
	);
	LUT3 #(
		.INIT('h31)
	) name1302 (
		\priority[45] ,
		\priority[46] ,
		\req[45] ,
		_w1560_
	);
	LUT4 #(
		.INIT('hc040)
	) name1303 (
		_w648_,
		_w652_,
		_w654_,
		_w1560_,
		_w1561_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1304 (
		_w984_,
		_w986_,
		_w987_,
		_w1561_,
		_w1562_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1305 (
		_w988_,
		_w990_,
		_w991_,
		_w1562_,
		_w1563_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1306 (
		_w992_,
		_w994_,
		_w995_,
		_w1563_,
		_w1564_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1307 (
		_w996_,
		_w998_,
		_w999_,
		_w1564_,
		_w1565_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1308 (
		_w1000_,
		_w1002_,
		_w1003_,
		_w1565_,
		_w1566_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1309 (
		_w1004_,
		_w1006_,
		_w1007_,
		_w1566_,
		_w1567_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name1310 (
		_w890_,
		_w1159_,
		_w1160_,
		_w1567_,
		_w1568_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1311 (
		_w891_,
		_w892_,
		_w894_,
		_w1568_,
		_w1569_
	);
	LUT4 #(
		.INIT('hb000)
	) name1312 (
		_w304_,
		_w310_,
		_w313_,
		_w1558_,
		_w1570_
	);
	LUT4 #(
		.INIT('h3b00)
	) name1313 (
		_w895_,
		_w896_,
		_w1569_,
		_w1570_,
		_w1571_
	);
	LUT2 #(
		.INIT('he)
	) name1314 (
		_w1559_,
		_w1571_,
		_w1572_
	);
	LUT3 #(
		.INIT('hb0)
	) name1315 (
		\priority[45] ,
		\req[44] ,
		\req[45] ,
		_w1573_
	);
	LUT2 #(
		.INIT('h4)
	) name1316 (
		_w475_,
		_w1573_,
		_w1574_
	);
	LUT3 #(
		.INIT('h31)
	) name1317 (
		\priority[46] ,
		\priority[47] ,
		\req[46] ,
		_w1575_
	);
	LUT4 #(
		.INIT('hc040)
	) name1318 (
		_w314_,
		_w321_,
		_w322_,
		_w1575_,
		_w1576_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1319 (
		_w330_,
		_w334_,
		_w342_,
		_w1576_,
		_w1577_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1320 (
		_w346_,
		_w353_,
		_w358_,
		_w1577_,
		_w1578_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1321 (
		_w365_,
		_w369_,
		_w377_,
		_w1578_,
		_w1579_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1322 (
		_w381_,
		_w388_,
		_w393_,
		_w1579_,
		_w1580_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1323 (
		_w400_,
		_w404_,
		_w412_,
		_w1580_,
		_w1581_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1324 (
		_w416_,
		_w1023_,
		_w1024_,
		_w1581_,
		_w1582_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name1325 (
		_w932_,
		_w1176_,
		_w1177_,
		_w1582_,
		_w1583_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1326 (
		_w933_,
		_w934_,
		_w936_,
		_w1583_,
		_w1584_
	);
	LUT4 #(
		.INIT('hb000)
	) name1327 (
		_w470_,
		_w476_,
		_w479_,
		_w1573_,
		_w1585_
	);
	LUT4 #(
		.INIT('h3b00)
	) name1328 (
		_w937_,
		_w938_,
		_w1584_,
		_w1585_,
		_w1586_
	);
	LUT2 #(
		.INIT('he)
	) name1329 (
		_w1574_,
		_w1586_,
		_w1587_
	);
	LUT3 #(
		.INIT('hb0)
	) name1330 (
		\priority[46] ,
		\req[45] ,
		\req[46] ,
		_w1588_
	);
	LUT2 #(
		.INIT('h4)
	) name1331 (
		_w641_,
		_w1588_,
		_w1589_
	);
	LUT3 #(
		.INIT('h31)
	) name1332 (
		\priority[47] ,
		\priority[48] ,
		\req[47] ,
		_w1590_
	);
	LUT4 #(
		.INIT('hc040)
	) name1333 (
		_w480_,
		_w487_,
		_w488_,
		_w1590_,
		_w1591_
	);
	LUT4 #(
		.INIT('h44c4)
	) name1334 (
		_w500_,
		_w508_,
		_w496_,
		_w1591_,
		_w1592_
	);
	LUT4 #(
		.INIT('h44c4)
	) name1335 (
		_w519_,
		_w524_,
		_w512_,
		_w1592_,
		_w1593_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1336 (
		_w531_,
		_w535_,
		_w543_,
		_w1593_,
		_w1594_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1337 (
		_w547_,
		_w554_,
		_w559_,
		_w1594_,
		_w1595_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1338 (
		_w566_,
		_w570_,
		_w578_,
		_w1595_,
		_w1596_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1339 (
		_w582_,
		_w1040_,
		_w1041_,
		_w1596_,
		_w1597_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name1340 (
		_w974_,
		_w1193_,
		_w1194_,
		_w1597_,
		_w1598_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1341 (
		_w975_,
		_w976_,
		_w978_,
		_w1598_,
		_w1599_
	);
	LUT4 #(
		.INIT('hb000)
	) name1342 (
		_w636_,
		_w642_,
		_w645_,
		_w1588_,
		_w1600_
	);
	LUT4 #(
		.INIT('h3b00)
	) name1343 (
		_w979_,
		_w980_,
		_w1599_,
		_w1600_,
		_w1601_
	);
	LUT2 #(
		.INIT('he)
	) name1344 (
		_w1589_,
		_w1601_,
		_w1602_
	);
	LUT3 #(
		.INIT('hb0)
	) name1345 (
		\priority[47] ,
		\req[46] ,
		\req[47] ,
		_w1603_
	);
	LUT2 #(
		.INIT('h4)
	) name1346 (
		_w320_,
		_w1603_,
		_w1604_
	);
	LUT3 #(
		.INIT('h31)
	) name1347 (
		\priority[48] ,
		\priority[49] ,
		\req[48] ,
		_w1605_
	);
	LUT4 #(
		.INIT('hc040)
	) name1348 (
		_w646_,
		_w653_,
		_w654_,
		_w1605_,
		_w1606_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1349 (
		_w662_,
		_w666_,
		_w674_,
		_w1606_,
		_w1607_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1350 (
		_w678_,
		_w685_,
		_w690_,
		_w1607_,
		_w1608_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1351 (
		_w697_,
		_w701_,
		_w709_,
		_w1608_,
		_w1609_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1352 (
		_w713_,
		_w720_,
		_w725_,
		_w1609_,
		_w1610_
	);
	LUT4 #(
		.INIT('h0c8c)
	) name1353 (
		_w732_,
		_w744_,
		_w736_,
		_w1610_,
		_w1611_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1354 (
		_w748_,
		_w1057_,
		_w1058_,
		_w1611_,
		_w1612_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1355 (
		_w272_,
		_w276_,
		_w283_,
		_w1612_,
		_w1613_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1356 (
		_w288_,
		_w295_,
		_w299_,
		_w1613_,
		_w1614_
	);
	LUT4 #(
		.INIT('hd000)
	) name1357 (
		_w309_,
		_w313_,
		_w317_,
		_w1603_,
		_w1615_
	);
	LUT4 #(
		.INIT('h3b00)
	) name1358 (
		_w307_,
		_w311_,
		_w1614_,
		_w1615_,
		_w1616_
	);
	LUT2 #(
		.INIT('he)
	) name1359 (
		_w1604_,
		_w1616_,
		_w1617_
	);
	LUT3 #(
		.INIT('hb0)
	) name1360 (
		\priority[48] ,
		\req[47] ,
		\req[48] ,
		_w1618_
	);
	LUT2 #(
		.INIT('h4)
	) name1361 (
		_w486_,
		_w1618_,
		_w1619_
	);
	LUT3 #(
		.INIT('h31)
	) name1362 (
		\priority[49] ,
		\priority[50] ,
		\req[49] ,
		_w1620_
	);
	LUT4 #(
		.INIT('ha020)
	) name1363 (
		_w321_,
		_w324_,
		_w331_,
		_w1620_,
		_w1621_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1364 (
		_w774_,
		_w775_,
		_w777_,
		_w1621_,
		_w1622_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1365 (
		_w778_,
		_w779_,
		_w781_,
		_w1622_,
		_w1623_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1366 (
		_w782_,
		_w783_,
		_w785_,
		_w1623_,
		_w1624_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1367 (
		_w786_,
		_w787_,
		_w789_,
		_w1624_,
		_w1625_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1368 (
		_w790_,
		_w791_,
		_w793_,
		_w1625_,
		_w1626_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1369 (
		_w794_,
		_w1074_,
		_w1075_,
		_w1626_,
		_w1627_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1370 (
		_w438_,
		_w442_,
		_w449_,
		_w1627_,
		_w1628_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1371 (
		_w454_,
		_w461_,
		_w465_,
		_w1628_,
		_w1629_
	);
	LUT4 #(
		.INIT('hd000)
	) name1372 (
		_w475_,
		_w479_,
		_w483_,
		_w1618_,
		_w1630_
	);
	LUT4 #(
		.INIT('h3b00)
	) name1373 (
		_w473_,
		_w477_,
		_w1629_,
		_w1630_,
		_w1631_
	);
	LUT2 #(
		.INIT('he)
	) name1374 (
		_w1619_,
		_w1631_,
		_w1632_
	);
	LUT3 #(
		.INIT('hb0)
	) name1375 (
		\priority[49] ,
		\req[48] ,
		\req[49] ,
		_w1633_
	);
	LUT2 #(
		.INIT('h4)
	) name1376 (
		_w652_,
		_w1633_,
		_w1634_
	);
	LUT3 #(
		.INIT('h31)
	) name1377 (
		\priority[50] ,
		\priority[51] ,
		\req[50] ,
		_w1635_
	);
	LUT4 #(
		.INIT('ha020)
	) name1378 (
		_w487_,
		_w490_,
		_w497_,
		_w1635_,
		_w1636_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1379 (
		_w818_,
		_w819_,
		_w821_,
		_w1636_,
		_w1637_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1380 (
		_w822_,
		_w823_,
		_w825_,
		_w1637_,
		_w1638_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1381 (
		_w826_,
		_w827_,
		_w829_,
		_w1638_,
		_w1639_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1382 (
		_w830_,
		_w831_,
		_w833_,
		_w1639_,
		_w1640_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1383 (
		_w834_,
		_w835_,
		_w837_,
		_w1640_,
		_w1641_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1384 (
		_w838_,
		_w1091_,
		_w1092_,
		_w1641_,
		_w1642_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1385 (
		_w604_,
		_w608_,
		_w615_,
		_w1642_,
		_w1643_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1386 (
		_w620_,
		_w627_,
		_w631_,
		_w1643_,
		_w1644_
	);
	LUT4 #(
		.INIT('hd000)
	) name1387 (
		_w641_,
		_w645_,
		_w649_,
		_w1633_,
		_w1645_
	);
	LUT4 #(
		.INIT('h3b00)
	) name1388 (
		_w639_,
		_w643_,
		_w1644_,
		_w1645_,
		_w1646_
	);
	LUT2 #(
		.INIT('he)
	) name1389 (
		_w1634_,
		_w1646_,
		_w1647_
	);
	LUT3 #(
		.INIT('hb0)
	) name1390 (
		\priority[50] ,
		\req[49] ,
		\req[50] ,
		_w1648_
	);
	LUT2 #(
		.INIT('h4)
	) name1391 (
		_w322_,
		_w1648_,
		_w1649_
	);
	LUT3 #(
		.INIT('h31)
	) name1392 (
		\priority[51] ,
		\priority[52] ,
		\req[51] ,
		_w1650_
	);
	LUT4 #(
		.INIT('ha020)
	) name1393 (
		_w653_,
		_w656_,
		_w663_,
		_w1650_,
		_w1651_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1394 (
		_w861_,
		_w862_,
		_w864_,
		_w1651_,
		_w1652_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1395 (
		_w865_,
		_w866_,
		_w868_,
		_w1652_,
		_w1653_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1396 (
		_w869_,
		_w870_,
		_w872_,
		_w1653_,
		_w1654_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1397 (
		_w873_,
		_w874_,
		_w876_,
		_w1654_,
		_w1655_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1398 (
		_w877_,
		_w878_,
		_w880_,
		_w1655_,
		_w1656_
	);
	LUT4 #(
		.INIT('h4c44)
	) name1399 (
		_w1108_,
		_w1109_,
		_w1656_,
		_w881_,
		_w1657_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1400 (
		_w761_,
		_w762_,
		_w763_,
		_w1657_,
		_w1658_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1401 (
		_w765_,
		_w766_,
		_w767_,
		_w1658_,
		_w1659_
	);
	LUT4 #(
		.INIT('h8a00)
	) name1402 (
		_w315_,
		_w317_,
		_w320_,
		_w1648_,
		_w1660_
	);
	LUT4 #(
		.INIT('h3b00)
	) name1403 (
		_w769_,
		_w770_,
		_w1659_,
		_w1660_,
		_w1661_
	);
	LUT2 #(
		.INIT('he)
	) name1404 (
		_w1649_,
		_w1661_,
		_w1662_
	);
	LUT3 #(
		.INIT('hb0)
	) name1405 (
		\priority[51] ,
		\req[50] ,
		\req[51] ,
		_w1663_
	);
	LUT2 #(
		.INIT('h4)
	) name1406 (
		_w488_,
		_w1663_,
		_w1664_
	);
	LUT3 #(
		.INIT('h31)
	) name1407 (
		\priority[52] ,
		\priority[53] ,
		\req[52] ,
		_w1665_
	);
	LUT4 #(
		.INIT('hc040)
	) name1408 (
		_w328_,
		_w331_,
		_w333_,
		_w1665_,
		_w1666_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1409 (
		_w903_,
		_w904_,
		_w906_,
		_w1666_,
		_w1667_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1410 (
		_w907_,
		_w908_,
		_w910_,
		_w1667_,
		_w1668_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1411 (
		_w911_,
		_w912_,
		_w914_,
		_w1668_,
		_w1669_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1412 (
		_w915_,
		_w916_,
		_w918_,
		_w1669_,
		_w1670_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1413 (
		_w919_,
		_w920_,
		_w922_,
		_w1670_,
		_w1671_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1414 (
		_w923_,
		_w1125_,
		_w1126_,
		_w1671_,
		_w1672_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1415 (
		_w805_,
		_w806_,
		_w807_,
		_w1672_,
		_w1673_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1416 (
		_w809_,
		_w810_,
		_w811_,
		_w1673_,
		_w1674_
	);
	LUT4 #(
		.INIT('h8a00)
	) name1417 (
		_w481_,
		_w483_,
		_w486_,
		_w1663_,
		_w1675_
	);
	LUT4 #(
		.INIT('h3b00)
	) name1418 (
		_w813_,
		_w814_,
		_w1674_,
		_w1675_,
		_w1676_
	);
	LUT2 #(
		.INIT('he)
	) name1419 (
		_w1664_,
		_w1676_,
		_w1677_
	);
	LUT3 #(
		.INIT('hb0)
	) name1420 (
		\priority[52] ,
		\req[51] ,
		\req[52] ,
		_w1678_
	);
	LUT2 #(
		.INIT('h4)
	) name1421 (
		_w654_,
		_w1678_,
		_w1679_
	);
	LUT3 #(
		.INIT('h31)
	) name1422 (
		\priority[53] ,
		\priority[54] ,
		\req[53] ,
		_w1680_
	);
	LUT4 #(
		.INIT('hc040)
	) name1423 (
		_w494_,
		_w497_,
		_w499_,
		_w1680_,
		_w1681_
	);
	LUT4 #(
		.INIT('h08cc)
	) name1424 (
		_w945_,
		_w948_,
		_w1681_,
		_w946_,
		_w1682_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1425 (
		_w949_,
		_w950_,
		_w952_,
		_w1682_,
		_w1683_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1426 (
		_w953_,
		_w954_,
		_w956_,
		_w1683_,
		_w1684_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1427 (
		_w957_,
		_w958_,
		_w960_,
		_w1684_,
		_w1685_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1428 (
		_w961_,
		_w962_,
		_w964_,
		_w1685_,
		_w1686_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1429 (
		_w965_,
		_w1142_,
		_w1143_,
		_w1686_,
		_w1687_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1430 (
		_w848_,
		_w849_,
		_w850_,
		_w1687_,
		_w1688_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1431 (
		_w852_,
		_w853_,
		_w854_,
		_w1688_,
		_w1689_
	);
	LUT4 #(
		.INIT('h8a00)
	) name1432 (
		_w647_,
		_w649_,
		_w652_,
		_w1678_,
		_w1690_
	);
	LUT4 #(
		.INIT('h3b00)
	) name1433 (
		_w856_,
		_w857_,
		_w1689_,
		_w1690_,
		_w1691_
	);
	LUT2 #(
		.INIT('he)
	) name1434 (
		_w1679_,
		_w1691_,
		_w1692_
	);
	LUT3 #(
		.INIT('hb0)
	) name1435 (
		\priority[53] ,
		\req[52] ,
		\req[53] ,
		_w1693_
	);
	LUT2 #(
		.INIT('h4)
	) name1436 (
		_w321_,
		_w1693_,
		_w1694_
	);
	LUT3 #(
		.INIT('h31)
	) name1437 (
		\priority[54] ,
		\priority[55] ,
		\req[54] ,
		_w1695_
	);
	LUT4 #(
		.INIT('hc040)
	) name1438 (
		_w660_,
		_w663_,
		_w665_,
		_w1695_,
		_w1696_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1439 (
		_w987_,
		_w988_,
		_w990_,
		_w1696_,
		_w1697_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1440 (
		_w991_,
		_w992_,
		_w994_,
		_w1697_,
		_w1698_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1441 (
		_w995_,
		_w996_,
		_w998_,
		_w1698_,
		_w1699_
	);
	LUT4 #(
		.INIT('h4c44)
	) name1442 (
		_w1000_,
		_w1002_,
		_w1699_,
		_w999_,
		_w1700_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1443 (
		_w1003_,
		_w1004_,
		_w1006_,
		_w1700_,
		_w1701_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1444 (
		_w1007_,
		_w1159_,
		_w1160_,
		_w1701_,
		_w1702_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1445 (
		_w890_,
		_w891_,
		_w892_,
		_w1702_,
		_w1703_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1446 (
		_w894_,
		_w895_,
		_w896_,
		_w1703_,
		_w1704_
	);
	LUT4 #(
		.INIT('hb000)
	) name1447 (
		_w315_,
		_w322_,
		_w325_,
		_w1693_,
		_w1705_
	);
	LUT4 #(
		.INIT('h3b00)
	) name1448 (
		_w898_,
		_w899_,
		_w1704_,
		_w1705_,
		_w1706_
	);
	LUT2 #(
		.INIT('he)
	) name1449 (
		_w1694_,
		_w1706_,
		_w1707_
	);
	LUT3 #(
		.INIT('hb0)
	) name1450 (
		\priority[54] ,
		\req[53] ,
		\req[54] ,
		_w1708_
	);
	LUT2 #(
		.INIT('h4)
	) name1451 (
		_w487_,
		_w1708_,
		_w1709_
	);
	LUT3 #(
		.INIT('h31)
	) name1452 (
		\priority[55] ,
		\priority[56] ,
		\req[55] ,
		_w1710_
	);
	LUT4 #(
		.INIT('hc040)
	) name1453 (
		_w326_,
		_w332_,
		_w333_,
		_w1710_,
		_w1711_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1454 (
		_w342_,
		_w346_,
		_w353_,
		_w1711_,
		_w1712_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1455 (
		_w358_,
		_w365_,
		_w369_,
		_w1712_,
		_w1713_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1456 (
		_w377_,
		_w381_,
		_w388_,
		_w1713_,
		_w1714_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1457 (
		_w393_,
		_w400_,
		_w404_,
		_w1714_,
		_w1715_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1458 (
		_w412_,
		_w416_,
		_w1023_,
		_w1715_,
		_w1716_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1459 (
		_w1024_,
		_w1176_,
		_w1177_,
		_w1716_,
		_w1717_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1460 (
		_w932_,
		_w933_,
		_w934_,
		_w1717_,
		_w1718_
	);
	LUT4 #(
		.INIT('h08cc)
	) name1461 (
		_w936_,
		_w938_,
		_w1718_,
		_w937_,
		_w1719_
	);
	LUT4 #(
		.INIT('hb000)
	) name1462 (
		_w481_,
		_w488_,
		_w491_,
		_w1708_,
		_w1720_
	);
	LUT4 #(
		.INIT('h3b00)
	) name1463 (
		_w940_,
		_w941_,
		_w1719_,
		_w1720_,
		_w1721_
	);
	LUT2 #(
		.INIT('he)
	) name1464 (
		_w1709_,
		_w1721_,
		_w1722_
	);
	LUT3 #(
		.INIT('hb0)
	) name1465 (
		\priority[55] ,
		\req[54] ,
		\req[55] ,
		_w1723_
	);
	LUT2 #(
		.INIT('h4)
	) name1466 (
		_w653_,
		_w1723_,
		_w1724_
	);
	LUT3 #(
		.INIT('h31)
	) name1467 (
		\priority[56] ,
		\priority[57] ,
		\req[56] ,
		_w1725_
	);
	LUT4 #(
		.INIT('hc040)
	) name1468 (
		_w492_,
		_w498_,
		_w499_,
		_w1725_,
		_w1726_
	);
	LUT4 #(
		.INIT('h0c8c)
	) name1469 (
		_w508_,
		_w519_,
		_w512_,
		_w1726_,
		_w1727_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1470 (
		_w524_,
		_w531_,
		_w535_,
		_w1727_,
		_w1728_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1471 (
		_w543_,
		_w547_,
		_w554_,
		_w1728_,
		_w1729_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1472 (
		_w559_,
		_w566_,
		_w570_,
		_w1729_,
		_w1730_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1473 (
		_w578_,
		_w582_,
		_w1040_,
		_w1730_,
		_w1731_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1474 (
		_w1041_,
		_w1193_,
		_w1194_,
		_w1731_,
		_w1732_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1475 (
		_w974_,
		_w975_,
		_w976_,
		_w1732_,
		_w1733_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1476 (
		_w978_,
		_w979_,
		_w980_,
		_w1733_,
		_w1734_
	);
	LUT4 #(
		.INIT('hb000)
	) name1477 (
		_w647_,
		_w654_,
		_w657_,
		_w1723_,
		_w1735_
	);
	LUT4 #(
		.INIT('h5d00)
	) name1478 (
		_w983_,
		_w982_,
		_w1734_,
		_w1735_,
		_w1736_
	);
	LUT2 #(
		.INIT('he)
	) name1479 (
		_w1724_,
		_w1736_,
		_w1737_
	);
	LUT3 #(
		.INIT('hb0)
	) name1480 (
		\priority[56] ,
		\req[55] ,
		\req[56] ,
		_w1738_
	);
	LUT2 #(
		.INIT('h4)
	) name1481 (
		_w331_,
		_w1738_,
		_w1739_
	);
	LUT3 #(
		.INIT('h31)
	) name1482 (
		\priority[57] ,
		\priority[58] ,
		\req[57] ,
		_w1740_
	);
	LUT4 #(
		.INIT('hc040)
	) name1483 (
		_w658_,
		_w664_,
		_w665_,
		_w1740_,
		_w1741_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1484 (
		_w674_,
		_w678_,
		_w685_,
		_w1741_,
		_w1742_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1485 (
		_w690_,
		_w697_,
		_w701_,
		_w1742_,
		_w1743_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1486 (
		_w709_,
		_w713_,
		_w720_,
		_w1743_,
		_w1744_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1487 (
		_w725_,
		_w732_,
		_w736_,
		_w1744_,
		_w1745_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1488 (
		_w744_,
		_w748_,
		_w1057_,
		_w1745_,
		_w1746_
	);
	LUT4 #(
		.INIT('h44c4)
	) name1489 (
		_w272_,
		_w276_,
		_w1058_,
		_w1746_,
		_w1747_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1490 (
		_w283_,
		_w288_,
		_w295_,
		_w1747_,
		_w1748_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1491 (
		_w299_,
		_w307_,
		_w311_,
		_w1748_,
		_w1749_
	);
	LUT4 #(
		.INIT('hd000)
	) name1492 (
		_w321_,
		_w325_,
		_w329_,
		_w1738_,
		_w1750_
	);
	LUT4 #(
		.INIT('h3b00)
	) name1493 (
		_w318_,
		_w323_,
		_w1749_,
		_w1750_,
		_w1751_
	);
	LUT2 #(
		.INIT('he)
	) name1494 (
		_w1739_,
		_w1751_,
		_w1752_
	);
	LUT3 #(
		.INIT('hb0)
	) name1495 (
		\priority[57] ,
		\req[56] ,
		\req[57] ,
		_w1753_
	);
	LUT2 #(
		.INIT('h4)
	) name1496 (
		_w497_,
		_w1753_,
		_w1754_
	);
	LUT3 #(
		.INIT('h31)
	) name1497 (
		\priority[58] ,
		\priority[59] ,
		\req[58] ,
		_w1755_
	);
	LUT4 #(
		.INIT('ha020)
	) name1498 (
		_w332_,
		_w336_,
		_w343_,
		_w1755_,
		_w1756_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1499 (
		_w777_,
		_w778_,
		_w779_,
		_w1756_,
		_w1757_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1500 (
		_w781_,
		_w782_,
		_w783_,
		_w1757_,
		_w1758_
	);
	LUT4 #(
		.INIT('h08cc)
	) name1501 (
		_w785_,
		_w787_,
		_w1758_,
		_w786_,
		_w1759_
	);
	LUT4 #(
		.INIT('h3b00)
	) name1502 (
		_w789_,
		_w790_,
		_w1759_,
		_w791_,
		_w1760_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1503 (
		_w793_,
		_w794_,
		_w1074_,
		_w1760_,
		_w1761_
	);
	LUT4 #(
		.INIT('h44c4)
	) name1504 (
		_w438_,
		_w442_,
		_w1075_,
		_w1761_,
		_w1762_
	);
	LUT4 #(
		.INIT('h08cc)
	) name1505 (
		_w449_,
		_w461_,
		_w1762_,
		_w454_,
		_w1763_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1506 (
		_w465_,
		_w473_,
		_w477_,
		_w1763_,
		_w1764_
	);
	LUT4 #(
		.INIT('hd000)
	) name1507 (
		_w487_,
		_w491_,
		_w495_,
		_w1753_,
		_w1765_
	);
	LUT4 #(
		.INIT('h5d00)
	) name1508 (
		_w489_,
		_w484_,
		_w1764_,
		_w1765_,
		_w1766_
	);
	LUT2 #(
		.INIT('he)
	) name1509 (
		_w1754_,
		_w1766_,
		_w1767_
	);
	LUT3 #(
		.INIT('hb0)
	) name1510 (
		\priority[58] ,
		\req[57] ,
		\req[58] ,
		_w1768_
	);
	LUT2 #(
		.INIT('h4)
	) name1511 (
		_w663_,
		_w1768_,
		_w1769_
	);
	LUT3 #(
		.INIT('h31)
	) name1512 (
		\priority[59] ,
		\priority[60] ,
		\req[59] ,
		_w1770_
	);
	LUT4 #(
		.INIT('ha020)
	) name1513 (
		_w498_,
		_w502_,
		_w509_,
		_w1770_,
		_w1771_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1514 (
		_w821_,
		_w822_,
		_w823_,
		_w1771_,
		_w1772_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1515 (
		_w825_,
		_w826_,
		_w827_,
		_w1772_,
		_w1773_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1516 (
		_w829_,
		_w830_,
		_w831_,
		_w1773_,
		_w1774_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1517 (
		_w833_,
		_w834_,
		_w835_,
		_w1774_,
		_w1775_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1518 (
		_w837_,
		_w838_,
		_w1091_,
		_w1775_,
		_w1776_
	);
	LUT4 #(
		.INIT('h44c4)
	) name1519 (
		_w604_,
		_w608_,
		_w1092_,
		_w1776_,
		_w1777_
	);
	LUT4 #(
		.INIT('h4c44)
	) name1520 (
		_w620_,
		_w627_,
		_w1777_,
		_w615_,
		_w1778_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1521 (
		_w631_,
		_w639_,
		_w643_,
		_w1778_,
		_w1779_
	);
	LUT4 #(
		.INIT('hd000)
	) name1522 (
		_w653_,
		_w657_,
		_w661_,
		_w1768_,
		_w1780_
	);
	LUT4 #(
		.INIT('h3b00)
	) name1523 (
		_w650_,
		_w655_,
		_w1779_,
		_w1780_,
		_w1781_
	);
	LUT2 #(
		.INIT('he)
	) name1524 (
		_w1769_,
		_w1781_,
		_w1782_
	);
	LUT3 #(
		.INIT('hb0)
	) name1525 (
		\priority[59] ,
		\req[58] ,
		\req[59] ,
		_w1783_
	);
	LUT2 #(
		.INIT('h4)
	) name1526 (
		_w333_,
		_w1783_,
		_w1784_
	);
	LUT3 #(
		.INIT('h31)
	) name1527 (
		\priority[60] ,
		\priority[61] ,
		\req[60] ,
		_w1785_
	);
	LUT4 #(
		.INIT('ha020)
	) name1528 (
		_w664_,
		_w668_,
		_w675_,
		_w1785_,
		_w1786_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1529 (
		_w864_,
		_w865_,
		_w866_,
		_w1786_,
		_w1787_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1530 (
		_w868_,
		_w869_,
		_w870_,
		_w1787_,
		_w1788_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1531 (
		_w872_,
		_w873_,
		_w874_,
		_w1788_,
		_w1789_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1532 (
		_w876_,
		_w877_,
		_w878_,
		_w1789_,
		_w1790_
	);
	LUT4 #(
		.INIT('h0c8c)
	) name1533 (
		_w880_,
		_w1108_,
		_w881_,
		_w1790_,
		_w1791_
	);
	LUT4 #(
		.INIT('h44c4)
	) name1534 (
		_w761_,
		_w762_,
		_w1109_,
		_w1791_,
		_w1792_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1535 (
		_w763_,
		_w765_,
		_w766_,
		_w1792_,
		_w1793_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1536 (
		_w767_,
		_w769_,
		_w770_,
		_w1793_,
		_w1794_
	);
	LUT4 #(
		.INIT('h8a00)
	) name1537 (
		_w327_,
		_w329_,
		_w331_,
		_w1783_,
		_w1795_
	);
	LUT4 #(
		.INIT('h3b00)
	) name1538 (
		_w771_,
		_w773_,
		_w1794_,
		_w1795_,
		_w1796_
	);
	LUT2 #(
		.INIT('he)
	) name1539 (
		_w1784_,
		_w1796_,
		_w1797_
	);
	LUT3 #(
		.INIT('hb0)
	) name1540 (
		\priority[60] ,
		\req[59] ,
		\req[60] ,
		_w1798_
	);
	LUT2 #(
		.INIT('h4)
	) name1541 (
		_w499_,
		_w1798_,
		_w1799_
	);
	LUT3 #(
		.INIT('h31)
	) name1542 (
		\priority[61] ,
		\priority[62] ,
		\req[61] ,
		_w1800_
	);
	LUT4 #(
		.INIT('hc040)
	) name1543 (
		_w340_,
		_w343_,
		_w345_,
		_w1800_,
		_w1801_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1544 (
		_w906_,
		_w907_,
		_w908_,
		_w1801_,
		_w1802_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1545 (
		_w910_,
		_w911_,
		_w912_,
		_w1802_,
		_w1803_
	);
	LUT4 #(
		.INIT('h4c44)
	) name1546 (
		_w915_,
		_w916_,
		_w1803_,
		_w914_,
		_w1804_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1547 (
		_w918_,
		_w919_,
		_w920_,
		_w1804_,
		_w1805_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1548 (
		_w922_,
		_w923_,
		_w1125_,
		_w1805_,
		_w1806_
	);
	LUT4 #(
		.INIT('h44c4)
	) name1549 (
		_w805_,
		_w806_,
		_w1126_,
		_w1806_,
		_w1807_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1550 (
		_w807_,
		_w809_,
		_w810_,
		_w1807_,
		_w1808_
	);
	LUT4 #(
		.INIT('h44c4)
	) name1551 (
		_w813_,
		_w814_,
		_w811_,
		_w1808_,
		_w1809_
	);
	LUT4 #(
		.INIT('h8a00)
	) name1552 (
		_w493_,
		_w495_,
		_w497_,
		_w1798_,
		_w1810_
	);
	LUT4 #(
		.INIT('h3b00)
	) name1553 (
		_w815_,
		_w817_,
		_w1809_,
		_w1810_,
		_w1811_
	);
	LUT2 #(
		.INIT('he)
	) name1554 (
		_w1799_,
		_w1811_,
		_w1812_
	);
	LUT3 #(
		.INIT('hb0)
	) name1555 (
		\priority[61] ,
		\req[60] ,
		\req[61] ,
		_w1813_
	);
	LUT2 #(
		.INIT('h4)
	) name1556 (
		_w665_,
		_w1813_,
		_w1814_
	);
	LUT3 #(
		.INIT('h31)
	) name1557 (
		\priority[62] ,
		\priority[63] ,
		\req[62] ,
		_w1815_
	);
	LUT4 #(
		.INIT('hc040)
	) name1558 (
		_w506_,
		_w509_,
		_w511_,
		_w1815_,
		_w1816_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1559 (
		_w948_,
		_w949_,
		_w950_,
		_w1816_,
		_w1817_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1560 (
		_w952_,
		_w953_,
		_w954_,
		_w1817_,
		_w1818_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1561 (
		_w956_,
		_w957_,
		_w958_,
		_w1818_,
		_w1819_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1562 (
		_w960_,
		_w961_,
		_w962_,
		_w1819_,
		_w1820_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1563 (
		_w964_,
		_w965_,
		_w1142_,
		_w1820_,
		_w1821_
	);
	LUT4 #(
		.INIT('h44c4)
	) name1564 (
		_w848_,
		_w849_,
		_w1143_,
		_w1821_,
		_w1822_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1565 (
		_w850_,
		_w852_,
		_w853_,
		_w1822_,
		_w1823_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1566 (
		_w854_,
		_w856_,
		_w857_,
		_w1823_,
		_w1824_
	);
	LUT4 #(
		.INIT('h8a00)
	) name1567 (
		_w659_,
		_w661_,
		_w663_,
		_w1813_,
		_w1825_
	);
	LUT4 #(
		.INIT('h3b00)
	) name1568 (
		_w858_,
		_w860_,
		_w1824_,
		_w1825_,
		_w1826_
	);
	LUT2 #(
		.INIT('he)
	) name1569 (
		_w1814_,
		_w1826_,
		_w1827_
	);
	LUT3 #(
		.INIT('hb0)
	) name1570 (
		\priority[62] ,
		\req[61] ,
		\req[62] ,
		_w1828_
	);
	LUT2 #(
		.INIT('h4)
	) name1571 (
		_w332_,
		_w1828_,
		_w1829_
	);
	LUT3 #(
		.INIT('h31)
	) name1572 (
		\priority[63] ,
		\priority[64] ,
		\req[63] ,
		_w1830_
	);
	LUT4 #(
		.INIT('hc040)
	) name1573 (
		_w672_,
		_w675_,
		_w677_,
		_w1830_,
		_w1831_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1574 (
		_w990_,
		_w991_,
		_w992_,
		_w1831_,
		_w1832_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1575 (
		_w994_,
		_w995_,
		_w996_,
		_w1832_,
		_w1833_
	);
	LUT4 #(
		.INIT('h0c8c)
	) name1576 (
		_w998_,
		_w1000_,
		_w999_,
		_w1833_,
		_w1834_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1577 (
		_w1002_,
		_w1003_,
		_w1004_,
		_w1834_,
		_w1835_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1578 (
		_w1006_,
		_w1007_,
		_w1159_,
		_w1835_,
		_w1836_
	);
	LUT4 #(
		.INIT('h44c4)
	) name1579 (
		_w890_,
		_w891_,
		_w1160_,
		_w1836_,
		_w1837_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1580 (
		_w892_,
		_w894_,
		_w895_,
		_w1837_,
		_w1838_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1581 (
		_w896_,
		_w898_,
		_w899_,
		_w1838_,
		_w1839_
	);
	LUT4 #(
		.INIT('hb000)
	) name1582 (
		_w327_,
		_w333_,
		_w337_,
		_w1828_,
		_w1840_
	);
	LUT4 #(
		.INIT('h3b00)
	) name1583 (
		_w900_,
		_w902_,
		_w1839_,
		_w1840_,
		_w1841_
	);
	LUT2 #(
		.INIT('he)
	) name1584 (
		_w1829_,
		_w1841_,
		_w1842_
	);
	LUT3 #(
		.INIT('hb0)
	) name1585 (
		\priority[63] ,
		\req[62] ,
		\req[63] ,
		_w1843_
	);
	LUT2 #(
		.INIT('h4)
	) name1586 (
		_w498_,
		_w1843_,
		_w1844_
	);
	LUT3 #(
		.INIT('h31)
	) name1587 (
		\priority[64] ,
		\priority[65] ,
		\req[64] ,
		_w1845_
	);
	LUT4 #(
		.INIT('hc040)
	) name1588 (
		_w338_,
		_w344_,
		_w345_,
		_w1845_,
		_w1846_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1589 (
		_w353_,
		_w358_,
		_w365_,
		_w1846_,
		_w1847_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1590 (
		_w369_,
		_w377_,
		_w381_,
		_w1847_,
		_w1848_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1591 (
		_w388_,
		_w393_,
		_w400_,
		_w1848_,
		_w1849_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1592 (
		_w404_,
		_w412_,
		_w416_,
		_w1849_,
		_w1850_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1593 (
		_w1023_,
		_w1024_,
		_w1176_,
		_w1850_,
		_w1851_
	);
	LUT4 #(
		.INIT('h44c4)
	) name1594 (
		_w932_,
		_w933_,
		_w1177_,
		_w1851_,
		_w1852_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1595 (
		_w934_,
		_w936_,
		_w937_,
		_w1852_,
		_w1853_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1596 (
		_w938_,
		_w940_,
		_w941_,
		_w1853_,
		_w1854_
	);
	LUT4 #(
		.INIT('hb000)
	) name1597 (
		_w493_,
		_w499_,
		_w503_,
		_w1843_,
		_w1855_
	);
	LUT4 #(
		.INIT('h3b00)
	) name1598 (
		_w942_,
		_w944_,
		_w1854_,
		_w1855_,
		_w1856_
	);
	LUT2 #(
		.INIT('he)
	) name1599 (
		_w1844_,
		_w1856_,
		_w1857_
	);
	LUT3 #(
		.INIT('hb0)
	) name1600 (
		\priority[64] ,
		\req[63] ,
		\req[64] ,
		_w1858_
	);
	LUT2 #(
		.INIT('h4)
	) name1601 (
		_w664_,
		_w1858_,
		_w1859_
	);
	LUT3 #(
		.INIT('h31)
	) name1602 (
		\priority[65] ,
		\priority[66] ,
		\req[65] ,
		_w1860_
	);
	LUT4 #(
		.INIT('hc040)
	) name1603 (
		_w504_,
		_w510_,
		_w511_,
		_w1860_,
		_w1861_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1604 (
		_w519_,
		_w524_,
		_w531_,
		_w1861_,
		_w1862_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1605 (
		_w535_,
		_w543_,
		_w547_,
		_w1862_,
		_w1863_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1606 (
		_w554_,
		_w559_,
		_w566_,
		_w1863_,
		_w1864_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1607 (
		_w570_,
		_w578_,
		_w582_,
		_w1864_,
		_w1865_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1608 (
		_w1040_,
		_w1041_,
		_w1193_,
		_w1865_,
		_w1866_
	);
	LUT4 #(
		.INIT('h44c4)
	) name1609 (
		_w974_,
		_w975_,
		_w1194_,
		_w1866_,
		_w1867_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1610 (
		_w976_,
		_w978_,
		_w979_,
		_w1867_,
		_w1868_
	);
	LUT4 #(
		.INIT('h0c8c)
	) name1611 (
		_w980_,
		_w983_,
		_w982_,
		_w1868_,
		_w1869_
	);
	LUT4 #(
		.INIT('hb000)
	) name1612 (
		_w659_,
		_w665_,
		_w669_,
		_w1858_,
		_w1870_
	);
	LUT4 #(
		.INIT('h3b00)
	) name1613 (
		_w984_,
		_w986_,
		_w1869_,
		_w1870_,
		_w1871_
	);
	LUT2 #(
		.INIT('he)
	) name1614 (
		_w1859_,
		_w1871_,
		_w1872_
	);
	LUT3 #(
		.INIT('hb0)
	) name1615 (
		\priority[65] ,
		\req[64] ,
		\req[65] ,
		_w1873_
	);
	LUT2 #(
		.INIT('h4)
	) name1616 (
		_w343_,
		_w1873_,
		_w1874_
	);
	LUT3 #(
		.INIT('h31)
	) name1617 (
		\priority[66] ,
		\priority[67] ,
		\req[66] ,
		_w1875_
	);
	LUT4 #(
		.INIT('hc040)
	) name1618 (
		_w670_,
		_w676_,
		_w677_,
		_w1875_,
		_w1876_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1619 (
		_w685_,
		_w690_,
		_w697_,
		_w1876_,
		_w1877_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1620 (
		_w701_,
		_w709_,
		_w713_,
		_w1877_,
		_w1878_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1621 (
		_w720_,
		_w725_,
		_w732_,
		_w1878_,
		_w1879_
	);
	LUT4 #(
		.INIT('h44c4)
	) name1622 (
		_w744_,
		_w748_,
		_w736_,
		_w1879_,
		_w1880_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name1623 (
		_w272_,
		_w1057_,
		_w1058_,
		_w1880_,
		_w1881_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1624 (
		_w276_,
		_w283_,
		_w288_,
		_w1881_,
		_w1882_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1625 (
		_w295_,
		_w299_,
		_w307_,
		_w1882_,
		_w1883_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1626 (
		_w311_,
		_w318_,
		_w323_,
		_w1883_,
		_w1884_
	);
	LUT4 #(
		.INIT('hd000)
	) name1627 (
		_w332_,
		_w337_,
		_w341_,
		_w1873_,
		_w1885_
	);
	LUT4 #(
		.INIT('h2f00)
	) name1628 (
		_w330_,
		_w1884_,
		_w334_,
		_w1885_,
		_w1886_
	);
	LUT2 #(
		.INIT('he)
	) name1629 (
		_w1874_,
		_w1886_,
		_w1887_
	);
	LUT3 #(
		.INIT('hb0)
	) name1630 (
		\priority[66] ,
		\req[65] ,
		\req[66] ,
		_w1888_
	);
	LUT2 #(
		.INIT('h4)
	) name1631 (
		_w509_,
		_w1888_,
		_w1889_
	);
	LUT3 #(
		.INIT('h31)
	) name1632 (
		\priority[67] ,
		\priority[68] ,
		\req[67] ,
		_w1890_
	);
	LUT4 #(
		.INIT('ha020)
	) name1633 (
		_w344_,
		_w347_,
		_w355_,
		_w1890_,
		_w1891_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1634 (
		_w779_,
		_w781_,
		_w782_,
		_w1891_,
		_w1892_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1635 (
		_w783_,
		_w785_,
		_w786_,
		_w1892_,
		_w1893_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1636 (
		_w787_,
		_w789_,
		_w790_,
		_w1893_,
		_w1894_
	);
	LUT4 #(
		.INIT('h44c4)
	) name1637 (
		_w793_,
		_w794_,
		_w791_,
		_w1894_,
		_w1895_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name1638 (
		_w438_,
		_w1074_,
		_w1075_,
		_w1895_,
		_w1896_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1639 (
		_w442_,
		_w449_,
		_w454_,
		_w1896_,
		_w1897_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1640 (
		_w461_,
		_w465_,
		_w473_,
		_w1897_,
		_w1898_
	);
	LUT4 #(
		.INIT('h0c8c)
	) name1641 (
		_w477_,
		_w489_,
		_w484_,
		_w1898_,
		_w1899_
	);
	LUT4 #(
		.INIT('hd000)
	) name1642 (
		_w498_,
		_w503_,
		_w507_,
		_w1888_,
		_w1900_
	);
	LUT4 #(
		.INIT('h5d00)
	) name1643 (
		_w500_,
		_w496_,
		_w1899_,
		_w1900_,
		_w1901_
	);
	LUT2 #(
		.INIT('he)
	) name1644 (
		_w1889_,
		_w1901_,
		_w1902_
	);
	LUT3 #(
		.INIT('hb0)
	) name1645 (
		\priority[67] ,
		\req[66] ,
		\req[67] ,
		_w1903_
	);
	LUT2 #(
		.INIT('h4)
	) name1646 (
		_w675_,
		_w1903_,
		_w1904_
	);
	LUT3 #(
		.INIT('h31)
	) name1647 (
		\priority[68] ,
		\priority[69] ,
		\req[68] ,
		_w1905_
	);
	LUT4 #(
		.INIT('ha020)
	) name1648 (
		_w510_,
		_w513_,
		_w521_,
		_w1905_,
		_w1906_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1649 (
		_w823_,
		_w825_,
		_w826_,
		_w1906_,
		_w1907_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1650 (
		_w827_,
		_w829_,
		_w830_,
		_w1907_,
		_w1908_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1651 (
		_w831_,
		_w833_,
		_w834_,
		_w1908_,
		_w1909_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1652 (
		_w835_,
		_w837_,
		_w838_,
		_w1909_,
		_w1910_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name1653 (
		_w604_,
		_w1091_,
		_w1092_,
		_w1910_,
		_w1911_
	);
	LUT4 #(
		.INIT('h0c8c)
	) name1654 (
		_w608_,
		_w620_,
		_w615_,
		_w1911_,
		_w1912_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1655 (
		_w627_,
		_w631_,
		_w639_,
		_w1912_,
		_w1913_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1656 (
		_w643_,
		_w650_,
		_w655_,
		_w1913_,
		_w1914_
	);
	LUT4 #(
		.INIT('hd000)
	) name1657 (
		_w664_,
		_w669_,
		_w673_,
		_w1903_,
		_w1915_
	);
	LUT4 #(
		.INIT('h3b00)
	) name1658 (
		_w662_,
		_w666_,
		_w1914_,
		_w1915_,
		_w1916_
	);
	LUT2 #(
		.INIT('he)
	) name1659 (
		_w1904_,
		_w1916_,
		_w1917_
	);
	LUT3 #(
		.INIT('hb0)
	) name1660 (
		\priority[68] ,
		\req[67] ,
		\req[68] ,
		_w1918_
	);
	LUT2 #(
		.INIT('h4)
	) name1661 (
		_w345_,
		_w1918_,
		_w1919_
	);
	LUT3 #(
		.INIT('h31)
	) name1662 (
		\priority[69] ,
		\priority[70] ,
		\req[69] ,
		_w1920_
	);
	LUT4 #(
		.INIT('ha020)
	) name1663 (
		_w676_,
		_w679_,
		_w687_,
		_w1920_,
		_w1921_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1664 (
		_w866_,
		_w868_,
		_w869_,
		_w1921_,
		_w1922_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1665 (
		_w870_,
		_w872_,
		_w873_,
		_w1922_,
		_w1923_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1666 (
		_w874_,
		_w876_,
		_w877_,
		_w1923_,
		_w1924_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1667 (
		_w878_,
		_w880_,
		_w881_,
		_w1924_,
		_w1925_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name1668 (
		_w761_,
		_w1108_,
		_w1109_,
		_w1925_,
		_w1926_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1669 (
		_w762_,
		_w763_,
		_w765_,
		_w1926_,
		_w1927_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1670 (
		_w766_,
		_w767_,
		_w769_,
		_w1927_,
		_w1928_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1671 (
		_w770_,
		_w771_,
		_w773_,
		_w1928_,
		_w1929_
	);
	LUT4 #(
		.INIT('h8a00)
	) name1672 (
		_w339_,
		_w341_,
		_w343_,
		_w1918_,
		_w1930_
	);
	LUT4 #(
		.INIT('h3b00)
	) name1673 (
		_w774_,
		_w775_,
		_w1929_,
		_w1930_,
		_w1931_
	);
	LUT2 #(
		.INIT('he)
	) name1674 (
		_w1919_,
		_w1931_,
		_w1932_
	);
	LUT3 #(
		.INIT('hb0)
	) name1675 (
		\priority[69] ,
		\req[68] ,
		\req[69] ,
		_w1933_
	);
	LUT2 #(
		.INIT('h4)
	) name1676 (
		_w511_,
		_w1933_,
		_w1934_
	);
	LUT3 #(
		.INIT('h31)
	) name1677 (
		\priority[70] ,
		\priority[71] ,
		\req[70] ,
		_w1935_
	);
	LUT4 #(
		.INIT('hc040)
	) name1678 (
		_w351_,
		_w355_,
		_w357_,
		_w1935_,
		_w1936_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1679 (
		_w908_,
		_w910_,
		_w911_,
		_w1936_,
		_w1937_
	);
	LUT4 #(
		.INIT('h0c8c)
	) name1680 (
		_w912_,
		_w915_,
		_w914_,
		_w1937_,
		_w1938_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1681 (
		_w916_,
		_w918_,
		_w919_,
		_w1938_,
		_w1939_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1682 (
		_w920_,
		_w922_,
		_w923_,
		_w1939_,
		_w1940_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name1683 (
		_w805_,
		_w1125_,
		_w1126_,
		_w1940_,
		_w1941_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1684 (
		_w806_,
		_w807_,
		_w809_,
		_w1941_,
		_w1942_
	);
	LUT4 #(
		.INIT('h0c8c)
	) name1685 (
		_w810_,
		_w813_,
		_w811_,
		_w1942_,
		_w1943_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1686 (
		_w814_,
		_w815_,
		_w817_,
		_w1943_,
		_w1944_
	);
	LUT4 #(
		.INIT('h8a00)
	) name1687 (
		_w505_,
		_w507_,
		_w509_,
		_w1933_,
		_w1945_
	);
	LUT4 #(
		.INIT('h3b00)
	) name1688 (
		_w818_,
		_w819_,
		_w1944_,
		_w1945_,
		_w1946_
	);
	LUT2 #(
		.INIT('he)
	) name1689 (
		_w1934_,
		_w1946_,
		_w1947_
	);
	LUT3 #(
		.INIT('hb0)
	) name1690 (
		\priority[70] ,
		\req[69] ,
		\req[70] ,
		_w1948_
	);
	LUT2 #(
		.INIT('h4)
	) name1691 (
		_w677_,
		_w1948_,
		_w1949_
	);
	LUT3 #(
		.INIT('h31)
	) name1692 (
		\priority[71] ,
		\priority[72] ,
		\req[71] ,
		_w1950_
	);
	LUT4 #(
		.INIT('hc040)
	) name1693 (
		_w517_,
		_w521_,
		_w523_,
		_w1950_,
		_w1951_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1694 (
		_w950_,
		_w952_,
		_w953_,
		_w1951_,
		_w1952_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1695 (
		_w954_,
		_w956_,
		_w957_,
		_w1952_,
		_w1953_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1696 (
		_w958_,
		_w960_,
		_w961_,
		_w1953_,
		_w1954_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1697 (
		_w962_,
		_w964_,
		_w965_,
		_w1954_,
		_w1955_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name1698 (
		_w848_,
		_w1142_,
		_w1143_,
		_w1955_,
		_w1956_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1699 (
		_w849_,
		_w850_,
		_w852_,
		_w1956_,
		_w1957_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1700 (
		_w853_,
		_w854_,
		_w856_,
		_w1957_,
		_w1958_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1701 (
		_w857_,
		_w858_,
		_w860_,
		_w1958_,
		_w1959_
	);
	LUT4 #(
		.INIT('h8a00)
	) name1702 (
		_w671_,
		_w673_,
		_w675_,
		_w1948_,
		_w1960_
	);
	LUT4 #(
		.INIT('h3b00)
	) name1703 (
		_w861_,
		_w862_,
		_w1959_,
		_w1960_,
		_w1961_
	);
	LUT2 #(
		.INIT('he)
	) name1704 (
		_w1949_,
		_w1961_,
		_w1962_
	);
	LUT3 #(
		.INIT('hb0)
	) name1705 (
		\priority[71] ,
		\req[70] ,
		\req[71] ,
		_w1963_
	);
	LUT2 #(
		.INIT('h4)
	) name1706 (
		_w344_,
		_w1963_,
		_w1964_
	);
	LUT3 #(
		.INIT('h31)
	) name1707 (
		\priority[72] ,
		\priority[73] ,
		\req[72] ,
		_w1965_
	);
	LUT4 #(
		.INIT('hc040)
	) name1708 (
		_w683_,
		_w687_,
		_w689_,
		_w1965_,
		_w1966_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1709 (
		_w992_,
		_w994_,
		_w995_,
		_w1966_,
		_w1967_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1710 (
		_w996_,
		_w998_,
		_w999_,
		_w1967_,
		_w1968_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1711 (
		_w1000_,
		_w1002_,
		_w1003_,
		_w1968_,
		_w1969_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1712 (
		_w1004_,
		_w1006_,
		_w1007_,
		_w1969_,
		_w1970_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name1713 (
		_w890_,
		_w1159_,
		_w1160_,
		_w1970_,
		_w1971_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1714 (
		_w891_,
		_w892_,
		_w894_,
		_w1971_,
		_w1972_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1715 (
		_w895_,
		_w896_,
		_w898_,
		_w1972_,
		_w1973_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1716 (
		_w899_,
		_w900_,
		_w902_,
		_w1973_,
		_w1974_
	);
	LUT4 #(
		.INIT('hb000)
	) name1717 (
		_w339_,
		_w345_,
		_w348_,
		_w1963_,
		_w1975_
	);
	LUT4 #(
		.INIT('h3b00)
	) name1718 (
		_w903_,
		_w904_,
		_w1974_,
		_w1975_,
		_w1976_
	);
	LUT2 #(
		.INIT('he)
	) name1719 (
		_w1964_,
		_w1976_,
		_w1977_
	);
	LUT3 #(
		.INIT('hb0)
	) name1720 (
		\priority[72] ,
		\req[71] ,
		\req[72] ,
		_w1978_
	);
	LUT2 #(
		.INIT('h4)
	) name1721 (
		_w510_,
		_w1978_,
		_w1979_
	);
	LUT3 #(
		.INIT('h31)
	) name1722 (
		\priority[73] ,
		\priority[74] ,
		\req[73] ,
		_w1980_
	);
	LUT4 #(
		.INIT('hc040)
	) name1723 (
		_w349_,
		_w356_,
		_w357_,
		_w1980_,
		_w1981_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1724 (
		_w365_,
		_w369_,
		_w377_,
		_w1981_,
		_w1982_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1725 (
		_w381_,
		_w388_,
		_w393_,
		_w1982_,
		_w1983_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1726 (
		_w400_,
		_w404_,
		_w412_,
		_w1983_,
		_w1984_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1727 (
		_w416_,
		_w1023_,
		_w1024_,
		_w1984_,
		_w1985_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name1728 (
		_w932_,
		_w1176_,
		_w1177_,
		_w1985_,
		_w1986_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1729 (
		_w933_,
		_w934_,
		_w936_,
		_w1986_,
		_w1987_
	);
	LUT4 #(
		.INIT('h44c4)
	) name1730 (
		_w938_,
		_w940_,
		_w937_,
		_w1987_,
		_w1988_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1731 (
		_w941_,
		_w942_,
		_w944_,
		_w1988_,
		_w1989_
	);
	LUT4 #(
		.INIT('hb000)
	) name1732 (
		_w505_,
		_w511_,
		_w514_,
		_w1978_,
		_w1990_
	);
	LUT4 #(
		.INIT('h3b00)
	) name1733 (
		_w945_,
		_w946_,
		_w1989_,
		_w1990_,
		_w1991_
	);
	LUT2 #(
		.INIT('he)
	) name1734 (
		_w1979_,
		_w1991_,
		_w1992_
	);
	LUT3 #(
		.INIT('hb0)
	) name1735 (
		\priority[73] ,
		\req[72] ,
		\req[73] ,
		_w1993_
	);
	LUT2 #(
		.INIT('h4)
	) name1736 (
		_w676_,
		_w1993_,
		_w1994_
	);
	LUT3 #(
		.INIT('h31)
	) name1737 (
		\priority[74] ,
		\priority[75] ,
		\req[74] ,
		_w1995_
	);
	LUT4 #(
		.INIT('hc040)
	) name1738 (
		_w515_,
		_w522_,
		_w523_,
		_w1995_,
		_w1996_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1739 (
		_w531_,
		_w535_,
		_w543_,
		_w1996_,
		_w1997_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1740 (
		_w547_,
		_w554_,
		_w559_,
		_w1997_,
		_w1998_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1741 (
		_w566_,
		_w570_,
		_w578_,
		_w1998_,
		_w1999_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1742 (
		_w582_,
		_w1040_,
		_w1041_,
		_w1999_,
		_w2000_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name1743 (
		_w974_,
		_w1193_,
		_w1194_,
		_w2000_,
		_w2001_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1744 (
		_w975_,
		_w976_,
		_w978_,
		_w2001_,
		_w2002_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1745 (
		_w979_,
		_w980_,
		_w982_,
		_w2002_,
		_w2003_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1746 (
		_w983_,
		_w984_,
		_w986_,
		_w2003_,
		_w2004_
	);
	LUT4 #(
		.INIT('hb000)
	) name1747 (
		_w671_,
		_w677_,
		_w680_,
		_w1993_,
		_w2005_
	);
	LUT4 #(
		.INIT('h3b00)
	) name1748 (
		_w987_,
		_w988_,
		_w2004_,
		_w2005_,
		_w2006_
	);
	LUT2 #(
		.INIT('he)
	) name1749 (
		_w1994_,
		_w2006_,
		_w2007_
	);
	LUT3 #(
		.INIT('hb0)
	) name1750 (
		\priority[74] ,
		\req[73] ,
		\req[74] ,
		_w2008_
	);
	LUT2 #(
		.INIT('h4)
	) name1751 (
		_w355_,
		_w2008_,
		_w2009_
	);
	LUT3 #(
		.INIT('h31)
	) name1752 (
		\priority[75] ,
		\priority[76] ,
		\req[75] ,
		_w2010_
	);
	LUT4 #(
		.INIT('hc040)
	) name1753 (
		_w681_,
		_w688_,
		_w689_,
		_w2010_,
		_w2011_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1754 (
		_w697_,
		_w701_,
		_w709_,
		_w2011_,
		_w2012_
	);
	LUT4 #(
		.INIT('h4c44)
	) name1755 (
		_w720_,
		_w725_,
		_w2012_,
		_w713_,
		_w2013_
	);
	LUT4 #(
		.INIT('h0c8c)
	) name1756 (
		_w732_,
		_w744_,
		_w736_,
		_w2013_,
		_w2014_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1757 (
		_w748_,
		_w1057_,
		_w1058_,
		_w2014_,
		_w2015_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1758 (
		_w272_,
		_w276_,
		_w283_,
		_w2015_,
		_w2016_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1759 (
		_w288_,
		_w295_,
		_w299_,
		_w2016_,
		_w2017_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1760 (
		_w307_,
		_w311_,
		_w318_,
		_w2017_,
		_w2018_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1761 (
		_w323_,
		_w330_,
		_w334_,
		_w2018_,
		_w2019_
	);
	LUT4 #(
		.INIT('hd000)
	) name1762 (
		_w344_,
		_w348_,
		_w352_,
		_w2008_,
		_w2020_
	);
	LUT4 #(
		.INIT('h3b00)
	) name1763 (
		_w342_,
		_w346_,
		_w2019_,
		_w2020_,
		_w2021_
	);
	LUT2 #(
		.INIT('he)
	) name1764 (
		_w2009_,
		_w2021_,
		_w2022_
	);
	LUT3 #(
		.INIT('hb0)
	) name1765 (
		\priority[75] ,
		\req[74] ,
		\req[75] ,
		_w2023_
	);
	LUT2 #(
		.INIT('h4)
	) name1766 (
		_w521_,
		_w2023_,
		_w2024_
	);
	LUT3 #(
		.INIT('h31)
	) name1767 (
		\priority[76] ,
		\priority[77] ,
		\req[76] ,
		_w2025_
	);
	LUT4 #(
		.INIT('ha020)
	) name1768 (
		_w356_,
		_w359_,
		_w366_,
		_w2025_,
		_w2026_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1769 (
		_w782_,
		_w783_,
		_w785_,
		_w2026_,
		_w2027_
	);
	LUT4 #(
		.INIT('h44c4)
	) name1770 (
		_w787_,
		_w789_,
		_w786_,
		_w2027_,
		_w2028_
	);
	LUT4 #(
		.INIT('h0c8c)
	) name1771 (
		_w790_,
		_w793_,
		_w791_,
		_w2028_,
		_w2029_
	);
	LUT4 #(
		.INIT('h3b00)
	) name1772 (
		_w794_,
		_w1074_,
		_w2029_,
		_w1075_,
		_w2030_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1773 (
		_w438_,
		_w442_,
		_w449_,
		_w2030_,
		_w2031_
	);
	LUT4 #(
		.INIT('h08aa)
	) name1774 (
		_w465_,
		_w454_,
		_w2031_,
		_w461_,
		_w2032_
	);
	LUT4 #(
		.INIT('h08cc)
	) name1775 (
		_w473_,
		_w484_,
		_w2032_,
		_w477_,
		_w2033_
	);
	LUT4 #(
		.INIT('h0c8c)
	) name1776 (
		_w489_,
		_w500_,
		_w496_,
		_w2033_,
		_w2034_
	);
	LUT4 #(
		.INIT('hd000)
	) name1777 (
		_w510_,
		_w514_,
		_w518_,
		_w2023_,
		_w2035_
	);
	LUT4 #(
		.INIT('h3b00)
	) name1778 (
		_w508_,
		_w512_,
		_w2034_,
		_w2035_,
		_w2036_
	);
	LUT2 #(
		.INIT('he)
	) name1779 (
		_w2024_,
		_w2036_,
		_w2037_
	);
	LUT3 #(
		.INIT('hb0)
	) name1780 (
		\priority[76] ,
		\req[75] ,
		\req[76] ,
		_w2038_
	);
	LUT2 #(
		.INIT('h4)
	) name1781 (
		_w687_,
		_w2038_,
		_w2039_
	);
	LUT3 #(
		.INIT('h31)
	) name1782 (
		\priority[77] ,
		\priority[78] ,
		\req[77] ,
		_w2040_
	);
	LUT4 #(
		.INIT('ha020)
	) name1783 (
		_w522_,
		_w525_,
		_w532_,
		_w2040_,
		_w2041_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1784 (
		_w826_,
		_w827_,
		_w829_,
		_w2041_,
		_w2042_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1785 (
		_w830_,
		_w831_,
		_w833_,
		_w2042_,
		_w2043_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1786 (
		_w834_,
		_w835_,
		_w837_,
		_w2043_,
		_w2044_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1787 (
		_w838_,
		_w1091_,
		_w1092_,
		_w2044_,
		_w2045_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1788 (
		_w604_,
		_w608_,
		_w615_,
		_w2045_,
		_w2046_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1789 (
		_w620_,
		_w627_,
		_w631_,
		_w2046_,
		_w2047_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1790 (
		_w639_,
		_w643_,
		_w650_,
		_w2047_,
		_w2048_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1791 (
		_w655_,
		_w662_,
		_w666_,
		_w2048_,
		_w2049_
	);
	LUT4 #(
		.INIT('hd000)
	) name1792 (
		_w676_,
		_w680_,
		_w684_,
		_w2038_,
		_w2050_
	);
	LUT4 #(
		.INIT('h3b00)
	) name1793 (
		_w674_,
		_w678_,
		_w2049_,
		_w2050_,
		_w2051_
	);
	LUT2 #(
		.INIT('he)
	) name1794 (
		_w2039_,
		_w2051_,
		_w2052_
	);
	LUT3 #(
		.INIT('hb0)
	) name1795 (
		\priority[77] ,
		\req[76] ,
		\req[77] ,
		_w2053_
	);
	LUT2 #(
		.INIT('h4)
	) name1796 (
		_w357_,
		_w2053_,
		_w2054_
	);
	LUT3 #(
		.INIT('h31)
	) name1797 (
		\priority[78] ,
		\priority[79] ,
		\req[78] ,
		_w2055_
	);
	LUT4 #(
		.INIT('ha020)
	) name1798 (
		_w688_,
		_w691_,
		_w698_,
		_w2055_,
		_w2056_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1799 (
		_w869_,
		_w870_,
		_w872_,
		_w2056_,
		_w2057_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1800 (
		_w873_,
		_w874_,
		_w876_,
		_w2057_,
		_w2058_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1801 (
		_w877_,
		_w878_,
		_w880_,
		_w2058_,
		_w2059_
	);
	LUT4 #(
		.INIT('h44c4)
	) name1802 (
		_w1108_,
		_w1109_,
		_w881_,
		_w2059_,
		_w2060_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1803 (
		_w761_,
		_w762_,
		_w763_,
		_w2060_,
		_w2061_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1804 (
		_w765_,
		_w766_,
		_w767_,
		_w2061_,
		_w2062_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1805 (
		_w769_,
		_w770_,
		_w771_,
		_w2062_,
		_w2063_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1806 (
		_w773_,
		_w774_,
		_w775_,
		_w2063_,
		_w2064_
	);
	LUT4 #(
		.INIT('h8a00)
	) name1807 (
		_w350_,
		_w352_,
		_w355_,
		_w2053_,
		_w2065_
	);
	LUT4 #(
		.INIT('h3b00)
	) name1808 (
		_w777_,
		_w778_,
		_w2064_,
		_w2065_,
		_w2066_
	);
	LUT2 #(
		.INIT('he)
	) name1809 (
		_w2054_,
		_w2066_,
		_w2067_
	);
	LUT3 #(
		.INIT('hb0)
	) name1810 (
		\priority[78] ,
		\req[77] ,
		\req[78] ,
		_w2068_
	);
	LUT2 #(
		.INIT('h4)
	) name1811 (
		_w523_,
		_w2068_,
		_w2069_
	);
	LUT3 #(
		.INIT('h31)
	) name1812 (
		\priority[79] ,
		\priority[80] ,
		\req[79] ,
		_w2070_
	);
	LUT4 #(
		.INIT('hc040)
	) name1813 (
		_w363_,
		_w366_,
		_w368_,
		_w2070_,
		_w2071_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1814 (
		_w911_,
		_w912_,
		_w914_,
		_w2071_,
		_w2072_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1815 (
		_w915_,
		_w916_,
		_w918_,
		_w2072_,
		_w2073_
	);
	LUT4 #(
		.INIT('h4c44)
	) name1816 (
		_w920_,
		_w922_,
		_w2073_,
		_w919_,
		_w2074_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1817 (
		_w923_,
		_w1125_,
		_w1126_,
		_w2074_,
		_w2075_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1818 (
		_w805_,
		_w806_,
		_w807_,
		_w2075_,
		_w2076_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1819 (
		_w809_,
		_w810_,
		_w811_,
		_w2076_,
		_w2077_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1820 (
		_w813_,
		_w814_,
		_w815_,
		_w2077_,
		_w2078_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1821 (
		_w817_,
		_w818_,
		_w819_,
		_w2078_,
		_w2079_
	);
	LUT4 #(
		.INIT('h8a00)
	) name1822 (
		_w516_,
		_w518_,
		_w521_,
		_w2068_,
		_w2080_
	);
	LUT4 #(
		.INIT('h3b00)
	) name1823 (
		_w821_,
		_w822_,
		_w2079_,
		_w2080_,
		_w2081_
	);
	LUT2 #(
		.INIT('he)
	) name1824 (
		_w2069_,
		_w2081_,
		_w2082_
	);
	LUT3 #(
		.INIT('hb0)
	) name1825 (
		\priority[79] ,
		\req[78] ,
		\req[79] ,
		_w2083_
	);
	LUT2 #(
		.INIT('h4)
	) name1826 (
		_w689_,
		_w2083_,
		_w2084_
	);
	LUT3 #(
		.INIT('h31)
	) name1827 (
		\priority[80] ,
		\priority[81] ,
		\req[80] ,
		_w2085_
	);
	LUT4 #(
		.INIT('hc040)
	) name1828 (
		_w529_,
		_w532_,
		_w534_,
		_w2085_,
		_w2086_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1829 (
		_w953_,
		_w954_,
		_w956_,
		_w2086_,
		_w2087_
	);
	LUT4 #(
		.INIT('h4c44)
	) name1830 (
		_w958_,
		_w960_,
		_w2087_,
		_w957_,
		_w2088_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1831 (
		_w961_,
		_w962_,
		_w964_,
		_w2088_,
		_w2089_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1832 (
		_w965_,
		_w1142_,
		_w1143_,
		_w2089_,
		_w2090_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1833 (
		_w848_,
		_w849_,
		_w850_,
		_w2090_,
		_w2091_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1834 (
		_w852_,
		_w853_,
		_w854_,
		_w2091_,
		_w2092_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1835 (
		_w856_,
		_w857_,
		_w858_,
		_w2092_,
		_w2093_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1836 (
		_w860_,
		_w861_,
		_w862_,
		_w2093_,
		_w2094_
	);
	LUT4 #(
		.INIT('h8a00)
	) name1837 (
		_w682_,
		_w684_,
		_w687_,
		_w2083_,
		_w2095_
	);
	LUT4 #(
		.INIT('h7500)
	) name1838 (
		_w865_,
		_w2094_,
		_w864_,
		_w2095_,
		_w2096_
	);
	LUT2 #(
		.INIT('he)
	) name1839 (
		_w2084_,
		_w2096_,
		_w2097_
	);
	LUT3 #(
		.INIT('hb0)
	) name1840 (
		\priority[80] ,
		\req[79] ,
		\req[80] ,
		_w2098_
	);
	LUT2 #(
		.INIT('h4)
	) name1841 (
		_w356_,
		_w2098_,
		_w2099_
	);
	LUT3 #(
		.INIT('h31)
	) name1842 (
		\priority[81] ,
		\priority[82] ,
		\req[81] ,
		_w2100_
	);
	LUT4 #(
		.INIT('hc040)
	) name1843 (
		_w695_,
		_w698_,
		_w700_,
		_w2100_,
		_w2101_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1844 (
		_w995_,
		_w996_,
		_w998_,
		_w2101_,
		_w2102_
	);
	LUT4 #(
		.INIT('h44c4)
	) name1845 (
		_w1000_,
		_w1002_,
		_w999_,
		_w2102_,
		_w2103_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1846 (
		_w1003_,
		_w1004_,
		_w1006_,
		_w2103_,
		_w2104_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1847 (
		_w1007_,
		_w1159_,
		_w1160_,
		_w2104_,
		_w2105_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1848 (
		_w890_,
		_w891_,
		_w892_,
		_w2105_,
		_w2106_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1849 (
		_w894_,
		_w895_,
		_w896_,
		_w2106_,
		_w2107_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1850 (
		_w898_,
		_w899_,
		_w900_,
		_w2107_,
		_w2108_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1851 (
		_w902_,
		_w903_,
		_w904_,
		_w2108_,
		_w2109_
	);
	LUT4 #(
		.INIT('hb000)
	) name1852 (
		_w350_,
		_w357_,
		_w360_,
		_w2098_,
		_w2110_
	);
	LUT4 #(
		.INIT('h3b00)
	) name1853 (
		_w906_,
		_w907_,
		_w2109_,
		_w2110_,
		_w2111_
	);
	LUT2 #(
		.INIT('he)
	) name1854 (
		_w2099_,
		_w2111_,
		_w2112_
	);
	LUT3 #(
		.INIT('hb0)
	) name1855 (
		\priority[81] ,
		\req[80] ,
		\req[81] ,
		_w2113_
	);
	LUT2 #(
		.INIT('h4)
	) name1856 (
		_w522_,
		_w2113_,
		_w2114_
	);
	LUT3 #(
		.INIT('h31)
	) name1857 (
		\priority[82] ,
		\priority[83] ,
		\req[82] ,
		_w2115_
	);
	LUT4 #(
		.INIT('hc040)
	) name1858 (
		_w361_,
		_w367_,
		_w368_,
		_w2115_,
		_w2116_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1859 (
		_w377_,
		_w381_,
		_w388_,
		_w2116_,
		_w2117_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1860 (
		_w393_,
		_w400_,
		_w404_,
		_w2117_,
		_w2118_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1861 (
		_w412_,
		_w416_,
		_w1023_,
		_w2118_,
		_w2119_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1862 (
		_w1024_,
		_w1176_,
		_w1177_,
		_w2119_,
		_w2120_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1863 (
		_w932_,
		_w933_,
		_w934_,
		_w2120_,
		_w2121_
	);
	LUT4 #(
		.INIT('h0c8c)
	) name1864 (
		_w936_,
		_w938_,
		_w937_,
		_w2121_,
		_w2122_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1865 (
		_w940_,
		_w941_,
		_w942_,
		_w2122_,
		_w2123_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1866 (
		_w944_,
		_w945_,
		_w946_,
		_w2123_,
		_w2124_
	);
	LUT4 #(
		.INIT('hb000)
	) name1867 (
		_w516_,
		_w523_,
		_w526_,
		_w2113_,
		_w2125_
	);
	LUT4 #(
		.INIT('h3b00)
	) name1868 (
		_w948_,
		_w949_,
		_w2124_,
		_w2125_,
		_w2126_
	);
	LUT2 #(
		.INIT('he)
	) name1869 (
		_w2114_,
		_w2126_,
		_w2127_
	);
	LUT3 #(
		.INIT('hb0)
	) name1870 (
		\priority[82] ,
		\req[81] ,
		\req[82] ,
		_w2128_
	);
	LUT2 #(
		.INIT('h4)
	) name1871 (
		_w688_,
		_w2128_,
		_w2129_
	);
	LUT3 #(
		.INIT('h31)
	) name1872 (
		\priority[83] ,
		\priority[84] ,
		\req[83] ,
		_w2130_
	);
	LUT4 #(
		.INIT('hc040)
	) name1873 (
		_w527_,
		_w533_,
		_w534_,
		_w2130_,
		_w2131_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1874 (
		_w543_,
		_w547_,
		_w554_,
		_w2131_,
		_w2132_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1875 (
		_w559_,
		_w566_,
		_w570_,
		_w2132_,
		_w2133_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1876 (
		_w578_,
		_w582_,
		_w1040_,
		_w2133_,
		_w2134_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1877 (
		_w1041_,
		_w1193_,
		_w1194_,
		_w2134_,
		_w2135_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1878 (
		_w974_,
		_w975_,
		_w976_,
		_w2135_,
		_w2136_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1879 (
		_w978_,
		_w979_,
		_w980_,
		_w2136_,
		_w2137_
	);
	LUT4 #(
		.INIT('h44c4)
	) name1880 (
		_w983_,
		_w984_,
		_w982_,
		_w2137_,
		_w2138_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1881 (
		_w986_,
		_w987_,
		_w988_,
		_w2138_,
		_w2139_
	);
	LUT4 #(
		.INIT('hb000)
	) name1882 (
		_w682_,
		_w689_,
		_w692_,
		_w2128_,
		_w2140_
	);
	LUT4 #(
		.INIT('h3b00)
	) name1883 (
		_w990_,
		_w991_,
		_w2139_,
		_w2140_,
		_w2141_
	);
	LUT2 #(
		.INIT('he)
	) name1884 (
		_w2129_,
		_w2141_,
		_w2142_
	);
	LUT3 #(
		.INIT('hb0)
	) name1885 (
		\priority[83] ,
		\req[82] ,
		\req[83] ,
		_w2143_
	);
	LUT2 #(
		.INIT('h4)
	) name1886 (
		_w366_,
		_w2143_,
		_w2144_
	);
	LUT3 #(
		.INIT('h31)
	) name1887 (
		\priority[84] ,
		\priority[85] ,
		\req[84] ,
		_w2145_
	);
	LUT4 #(
		.INIT('hc040)
	) name1888 (
		_w693_,
		_w699_,
		_w700_,
		_w2145_,
		_w2146_
	);
	LUT4 #(
		.INIT('h0c8c)
	) name1889 (
		_w709_,
		_w720_,
		_w713_,
		_w2146_,
		_w2147_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1890 (
		_w725_,
		_w732_,
		_w736_,
		_w2147_,
		_w2148_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1891 (
		_w744_,
		_w748_,
		_w1057_,
		_w2148_,
		_w2149_
	);
	LUT4 #(
		.INIT('h44c4)
	) name1892 (
		_w272_,
		_w276_,
		_w1058_,
		_w2149_,
		_w2150_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1893 (
		_w283_,
		_w288_,
		_w295_,
		_w2150_,
		_w2151_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1894 (
		_w299_,
		_w307_,
		_w311_,
		_w2151_,
		_w2152_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1895 (
		_w318_,
		_w323_,
		_w330_,
		_w2152_,
		_w2153_
	);
	LUT4 #(
		.INIT('h44c4)
	) name1896 (
		_w342_,
		_w346_,
		_w334_,
		_w2153_,
		_w2154_
	);
	LUT4 #(
		.INIT('hd000)
	) name1897 (
		_w356_,
		_w360_,
		_w364_,
		_w2143_,
		_w2155_
	);
	LUT4 #(
		.INIT('h3b00)
	) name1898 (
		_w353_,
		_w358_,
		_w2154_,
		_w2155_,
		_w2156_
	);
	LUT2 #(
		.INIT('he)
	) name1899 (
		_w2144_,
		_w2156_,
		_w2157_
	);
	LUT3 #(
		.INIT('hb0)
	) name1900 (
		\priority[84] ,
		\req[83] ,
		\req[84] ,
		_w2158_
	);
	LUT2 #(
		.INIT('h4)
	) name1901 (
		_w532_,
		_w2158_,
		_w2159_
	);
	LUT3 #(
		.INIT('h31)
	) name1902 (
		\priority[85] ,
		\priority[86] ,
		\req[85] ,
		_w2160_
	);
	LUT4 #(
		.INIT('ha020)
	) name1903 (
		_w367_,
		_w371_,
		_w378_,
		_w2160_,
		_w2161_
	);
	LUT4 #(
		.INIT('h0c8c)
	) name1904 (
		_w785_,
		_w787_,
		_w786_,
		_w2161_,
		_w2162_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1905 (
		_w789_,
		_w790_,
		_w791_,
		_w2162_,
		_w2163_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1906 (
		_w793_,
		_w794_,
		_w1074_,
		_w2163_,
		_w2164_
	);
	LUT4 #(
		.INIT('h44c4)
	) name1907 (
		_w438_,
		_w442_,
		_w1075_,
		_w2164_,
		_w2165_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1908 (
		_w449_,
		_w454_,
		_w461_,
		_w2165_,
		_w2166_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1909 (
		_w465_,
		_w473_,
		_w477_,
		_w2166_,
		_w2167_
	);
	LUT4 #(
		.INIT('h50d0)
	) name1910 (
		_w489_,
		_w484_,
		_w496_,
		_w2167_,
		_w2168_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1911 (
		_w500_,
		_w508_,
		_w512_,
		_w2168_,
		_w2169_
	);
	LUT4 #(
		.INIT('hd000)
	) name1912 (
		_w522_,
		_w526_,
		_w530_,
		_w2158_,
		_w2170_
	);
	LUT4 #(
		.INIT('h3b00)
	) name1913 (
		_w519_,
		_w524_,
		_w2169_,
		_w2170_,
		_w2171_
	);
	LUT2 #(
		.INIT('he)
	) name1914 (
		_w2159_,
		_w2171_,
		_w2172_
	);
	LUT3 #(
		.INIT('hb0)
	) name1915 (
		\priority[85] ,
		\req[84] ,
		\req[85] ,
		_w2173_
	);
	LUT2 #(
		.INIT('h4)
	) name1916 (
		_w698_,
		_w2173_,
		_w2174_
	);
	LUT3 #(
		.INIT('h31)
	) name1917 (
		\priority[86] ,
		\priority[87] ,
		\req[86] ,
		_w2175_
	);
	LUT4 #(
		.INIT('ha020)
	) name1918 (
		_w533_,
		_w537_,
		_w544_,
		_w2175_,
		_w2176_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1919 (
		_w829_,
		_w830_,
		_w831_,
		_w2176_,
		_w2177_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1920 (
		_w833_,
		_w834_,
		_w835_,
		_w2177_,
		_w2178_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1921 (
		_w837_,
		_w838_,
		_w1091_,
		_w2178_,
		_w2179_
	);
	LUT4 #(
		.INIT('h44c4)
	) name1922 (
		_w604_,
		_w608_,
		_w1092_,
		_w2179_,
		_w2180_
	);
	LUT4 #(
		.INIT('h44c4)
	) name1923 (
		_w620_,
		_w627_,
		_w615_,
		_w2180_,
		_w2181_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1924 (
		_w631_,
		_w639_,
		_w643_,
		_w2181_,
		_w2182_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1925 (
		_w650_,
		_w655_,
		_w662_,
		_w2182_,
		_w2183_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1926 (
		_w666_,
		_w674_,
		_w678_,
		_w2183_,
		_w2184_
	);
	LUT4 #(
		.INIT('hd000)
	) name1927 (
		_w688_,
		_w692_,
		_w696_,
		_w2173_,
		_w2185_
	);
	LUT4 #(
		.INIT('h3b00)
	) name1928 (
		_w685_,
		_w690_,
		_w2184_,
		_w2185_,
		_w2186_
	);
	LUT2 #(
		.INIT('he)
	) name1929 (
		_w2174_,
		_w2186_,
		_w2187_
	);
	LUT3 #(
		.INIT('hb0)
	) name1930 (
		\priority[86] ,
		\req[85] ,
		\req[86] ,
		_w2188_
	);
	LUT2 #(
		.INIT('h4)
	) name1931 (
		_w368_,
		_w2188_,
		_w2189_
	);
	LUT3 #(
		.INIT('h31)
	) name1932 (
		\priority[87] ,
		\priority[88] ,
		\req[87] ,
		_w2190_
	);
	LUT4 #(
		.INIT('ha020)
	) name1933 (
		_w699_,
		_w703_,
		_w710_,
		_w2190_,
		_w2191_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1934 (
		_w872_,
		_w873_,
		_w874_,
		_w2191_,
		_w2192_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1935 (
		_w876_,
		_w877_,
		_w878_,
		_w2192_,
		_w2193_
	);
	LUT4 #(
		.INIT('h0c8c)
	) name1936 (
		_w880_,
		_w1108_,
		_w881_,
		_w2193_,
		_w2194_
	);
	LUT4 #(
		.INIT('h44c4)
	) name1937 (
		_w761_,
		_w762_,
		_w1109_,
		_w2194_,
		_w2195_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1938 (
		_w763_,
		_w765_,
		_w766_,
		_w2195_,
		_w2196_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1939 (
		_w767_,
		_w769_,
		_w770_,
		_w2196_,
		_w2197_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1940 (
		_w771_,
		_w773_,
		_w774_,
		_w2197_,
		_w2198_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1941 (
		_w775_,
		_w777_,
		_w778_,
		_w2198_,
		_w2199_
	);
	LUT4 #(
		.INIT('h8a00)
	) name1942 (
		_w362_,
		_w364_,
		_w366_,
		_w2188_,
		_w2200_
	);
	LUT4 #(
		.INIT('h3b00)
	) name1943 (
		_w779_,
		_w781_,
		_w2199_,
		_w2200_,
		_w2201_
	);
	LUT2 #(
		.INIT('he)
	) name1944 (
		_w2189_,
		_w2201_,
		_w2202_
	);
	LUT3 #(
		.INIT('hb0)
	) name1945 (
		\priority[87] ,
		\req[86] ,
		\req[87] ,
		_w2203_
	);
	LUT2 #(
		.INIT('h4)
	) name1946 (
		_w534_,
		_w2203_,
		_w2204_
	);
	LUT3 #(
		.INIT('h31)
	) name1947 (
		\priority[88] ,
		\priority[89] ,
		\req[88] ,
		_w2205_
	);
	LUT4 #(
		.INIT('hc040)
	) name1948 (
		_w375_,
		_w378_,
		_w380_,
		_w2205_,
		_w2206_
	);
	LUT4 #(
		.INIT('h44c4)
	) name1949 (
		_w915_,
		_w916_,
		_w914_,
		_w2206_,
		_w2207_
	);
	LUT4 #(
		.INIT('h0c8c)
	) name1950 (
		_w918_,
		_w920_,
		_w919_,
		_w2207_,
		_w2208_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1951 (
		_w922_,
		_w923_,
		_w1125_,
		_w2208_,
		_w2209_
	);
	LUT4 #(
		.INIT('h44c4)
	) name1952 (
		_w805_,
		_w806_,
		_w1126_,
		_w2209_,
		_w2210_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1953 (
		_w807_,
		_w809_,
		_w810_,
		_w2210_,
		_w2211_
	);
	LUT4 #(
		.INIT('h44c4)
	) name1954 (
		_w813_,
		_w814_,
		_w811_,
		_w2211_,
		_w2212_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1955 (
		_w815_,
		_w817_,
		_w818_,
		_w2212_,
		_w2213_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1956 (
		_w819_,
		_w821_,
		_w822_,
		_w2213_,
		_w2214_
	);
	LUT4 #(
		.INIT('h8a00)
	) name1957 (
		_w528_,
		_w530_,
		_w532_,
		_w2203_,
		_w2215_
	);
	LUT4 #(
		.INIT('h3b00)
	) name1958 (
		_w823_,
		_w825_,
		_w2214_,
		_w2215_,
		_w2216_
	);
	LUT2 #(
		.INIT('he)
	) name1959 (
		_w2204_,
		_w2216_,
		_w2217_
	);
	LUT3 #(
		.INIT('hb0)
	) name1960 (
		\priority[88] ,
		\req[87] ,
		\req[88] ,
		_w2218_
	);
	LUT2 #(
		.INIT('h4)
	) name1961 (
		_w700_,
		_w2218_,
		_w2219_
	);
	LUT3 #(
		.INIT('h31)
	) name1962 (
		\priority[89] ,
		\priority[90] ,
		\req[89] ,
		_w2220_
	);
	LUT4 #(
		.INIT('hc040)
	) name1963 (
		_w541_,
		_w544_,
		_w546_,
		_w2220_,
		_w2221_
	);
	LUT4 #(
		.INIT('h0c8c)
	) name1964 (
		_w956_,
		_w958_,
		_w957_,
		_w2221_,
		_w2222_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1965 (
		_w960_,
		_w961_,
		_w962_,
		_w2222_,
		_w2223_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1966 (
		_w964_,
		_w965_,
		_w1142_,
		_w2223_,
		_w2224_
	);
	LUT4 #(
		.INIT('h44c4)
	) name1967 (
		_w848_,
		_w849_,
		_w1143_,
		_w2224_,
		_w2225_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1968 (
		_w850_,
		_w852_,
		_w853_,
		_w2225_,
		_w2226_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1969 (
		_w854_,
		_w856_,
		_w857_,
		_w2226_,
		_w2227_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1970 (
		_w858_,
		_w860_,
		_w861_,
		_w2227_,
		_w2228_
	);
	LUT4 #(
		.INIT('h0c8c)
	) name1971 (
		_w862_,
		_w865_,
		_w864_,
		_w2228_,
		_w2229_
	);
	LUT4 #(
		.INIT('h8a00)
	) name1972 (
		_w694_,
		_w696_,
		_w698_,
		_w2218_,
		_w2230_
	);
	LUT4 #(
		.INIT('h7500)
	) name1973 (
		_w868_,
		_w2229_,
		_w866_,
		_w2230_,
		_w2231_
	);
	LUT2 #(
		.INIT('he)
	) name1974 (
		_w2219_,
		_w2231_,
		_w2232_
	);
	LUT3 #(
		.INIT('hb0)
	) name1975 (
		\priority[89] ,
		\req[88] ,
		\req[89] ,
		_w2233_
	);
	LUT2 #(
		.INIT('h4)
	) name1976 (
		_w367_,
		_w2233_,
		_w2234_
	);
	LUT3 #(
		.INIT('h31)
	) name1977 (
		\priority[90] ,
		\priority[91] ,
		\req[90] ,
		_w2235_
	);
	LUT4 #(
		.INIT('hc040)
	) name1978 (
		_w707_,
		_w710_,
		_w712_,
		_w2235_,
		_w2236_
	);
	LUT4 #(
		.INIT('h0c8c)
	) name1979 (
		_w998_,
		_w1000_,
		_w999_,
		_w2236_,
		_w2237_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1980 (
		_w1002_,
		_w1003_,
		_w1004_,
		_w2237_,
		_w2238_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1981 (
		_w1006_,
		_w1007_,
		_w1159_,
		_w2238_,
		_w2239_
	);
	LUT4 #(
		.INIT('h44c4)
	) name1982 (
		_w890_,
		_w891_,
		_w1160_,
		_w2239_,
		_w2240_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1983 (
		_w892_,
		_w894_,
		_w895_,
		_w2240_,
		_w2241_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1984 (
		_w896_,
		_w898_,
		_w899_,
		_w2241_,
		_w2242_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1985 (
		_w900_,
		_w902_,
		_w903_,
		_w2242_,
		_w2243_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1986 (
		_w904_,
		_w906_,
		_w907_,
		_w2243_,
		_w2244_
	);
	LUT4 #(
		.INIT('hb000)
	) name1987 (
		_w362_,
		_w368_,
		_w372_,
		_w2233_,
		_w2245_
	);
	LUT4 #(
		.INIT('h3b00)
	) name1988 (
		_w908_,
		_w910_,
		_w2244_,
		_w2245_,
		_w2246_
	);
	LUT2 #(
		.INIT('he)
	) name1989 (
		_w2234_,
		_w2246_,
		_w2247_
	);
	LUT3 #(
		.INIT('hb0)
	) name1990 (
		\priority[90] ,
		\req[89] ,
		\req[90] ,
		_w2248_
	);
	LUT2 #(
		.INIT('h4)
	) name1991 (
		_w533_,
		_w2248_,
		_w2249_
	);
	LUT3 #(
		.INIT('h31)
	) name1992 (
		\priority[91] ,
		\priority[92] ,
		\req[91] ,
		_w2250_
	);
	LUT4 #(
		.INIT('hc040)
	) name1993 (
		_w373_,
		_w379_,
		_w380_,
		_w2250_,
		_w2251_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1994 (
		_w388_,
		_w393_,
		_w400_,
		_w2251_,
		_w2252_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1995 (
		_w404_,
		_w412_,
		_w416_,
		_w2252_,
		_w2253_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1996 (
		_w1023_,
		_w1024_,
		_w1176_,
		_w2253_,
		_w2254_
	);
	LUT4 #(
		.INIT('h44c4)
	) name1997 (
		_w932_,
		_w933_,
		_w1177_,
		_w2254_,
		_w2255_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1998 (
		_w934_,
		_w936_,
		_w937_,
		_w2255_,
		_w2256_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1999 (
		_w938_,
		_w940_,
		_w941_,
		_w2256_,
		_w2257_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2000 (
		_w942_,
		_w944_,
		_w945_,
		_w2257_,
		_w2258_
	);
	LUT4 #(
		.INIT('h44c4)
	) name2001 (
		_w948_,
		_w949_,
		_w946_,
		_w2258_,
		_w2259_
	);
	LUT4 #(
		.INIT('hb000)
	) name2002 (
		_w528_,
		_w534_,
		_w538_,
		_w2248_,
		_w2260_
	);
	LUT4 #(
		.INIT('h3b00)
	) name2003 (
		_w950_,
		_w952_,
		_w2259_,
		_w2260_,
		_w2261_
	);
	LUT2 #(
		.INIT('he)
	) name2004 (
		_w2249_,
		_w2261_,
		_w2262_
	);
	LUT3 #(
		.INIT('hb0)
	) name2005 (
		\priority[91] ,
		\req[90] ,
		\req[91] ,
		_w2263_
	);
	LUT2 #(
		.INIT('h4)
	) name2006 (
		_w699_,
		_w2263_,
		_w2264_
	);
	LUT3 #(
		.INIT('h31)
	) name2007 (
		\priority[92] ,
		\priority[93] ,
		\req[92] ,
		_w2265_
	);
	LUT4 #(
		.INIT('hc040)
	) name2008 (
		_w539_,
		_w545_,
		_w546_,
		_w2265_,
		_w2266_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2009 (
		_w554_,
		_w559_,
		_w566_,
		_w2266_,
		_w2267_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2010 (
		_w570_,
		_w578_,
		_w582_,
		_w2267_,
		_w2268_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2011 (
		_w1040_,
		_w1041_,
		_w1193_,
		_w2268_,
		_w2269_
	);
	LUT4 #(
		.INIT('h44c4)
	) name2012 (
		_w974_,
		_w975_,
		_w1194_,
		_w2269_,
		_w2270_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2013 (
		_w976_,
		_w978_,
		_w979_,
		_w2270_,
		_w2271_
	);
	LUT4 #(
		.INIT('h0c8c)
	) name2014 (
		_w980_,
		_w983_,
		_w982_,
		_w2271_,
		_w2272_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2015 (
		_w984_,
		_w986_,
		_w987_,
		_w2272_,
		_w2273_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2016 (
		_w988_,
		_w990_,
		_w991_,
		_w2273_,
		_w2274_
	);
	LUT4 #(
		.INIT('hb000)
	) name2017 (
		_w694_,
		_w700_,
		_w704_,
		_w2263_,
		_w2275_
	);
	LUT4 #(
		.INIT('h3b00)
	) name2018 (
		_w992_,
		_w994_,
		_w2274_,
		_w2275_,
		_w2276_
	);
	LUT2 #(
		.INIT('he)
	) name2019 (
		_w2264_,
		_w2276_,
		_w2277_
	);
	LUT3 #(
		.INIT('hb0)
	) name2020 (
		\priority[92] ,
		\req[91] ,
		\req[92] ,
		_w2278_
	);
	LUT2 #(
		.INIT('h4)
	) name2021 (
		_w378_,
		_w2278_,
		_w2279_
	);
	LUT3 #(
		.INIT('h31)
	) name2022 (
		\priority[93] ,
		\priority[94] ,
		\req[93] ,
		_w2280_
	);
	LUT4 #(
		.INIT('hc040)
	) name2023 (
		_w705_,
		_w711_,
		_w712_,
		_w2280_,
		_w2281_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2024 (
		_w720_,
		_w725_,
		_w732_,
		_w2281_,
		_w2282_
	);
	LUT4 #(
		.INIT('h44c4)
	) name2025 (
		_w744_,
		_w748_,
		_w736_,
		_w2282_,
		_w2283_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name2026 (
		_w272_,
		_w1057_,
		_w1058_,
		_w2283_,
		_w2284_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2027 (
		_w276_,
		_w283_,
		_w288_,
		_w2284_,
		_w2285_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2028 (
		_w295_,
		_w299_,
		_w307_,
		_w2285_,
		_w2286_
	);
	LUT4 #(
		.INIT('h3b00)
	) name2029 (
		_w311_,
		_w318_,
		_w2286_,
		_w323_,
		_w2287_
	);
	LUT4 #(
		.INIT('h0c8c)
	) name2030 (
		_w330_,
		_w342_,
		_w334_,
		_w2287_,
		_w2288_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2031 (
		_w346_,
		_w353_,
		_w358_,
		_w2288_,
		_w2289_
	);
	LUT4 #(
		.INIT('hd000)
	) name2032 (
		_w367_,
		_w372_,
		_w376_,
		_w2278_,
		_w2290_
	);
	LUT4 #(
		.INIT('h3b00)
	) name2033 (
		_w365_,
		_w369_,
		_w2289_,
		_w2290_,
		_w2291_
	);
	LUT2 #(
		.INIT('he)
	) name2034 (
		_w2279_,
		_w2291_,
		_w2292_
	);
	LUT3 #(
		.INIT('hb0)
	) name2035 (
		\priority[93] ,
		\req[92] ,
		\req[93] ,
		_w2293_
	);
	LUT2 #(
		.INIT('h4)
	) name2036 (
		_w544_,
		_w2293_,
		_w2294_
	);
	LUT3 #(
		.INIT('h31)
	) name2037 (
		\priority[94] ,
		\priority[95] ,
		\req[94] ,
		_w2295_
	);
	LUT4 #(
		.INIT('ha020)
	) name2038 (
		_w379_,
		_w382_,
		_w390_,
		_w2295_,
		_w2296_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2039 (
		_w787_,
		_w789_,
		_w790_,
		_w2296_,
		_w2297_
	);
	LUT4 #(
		.INIT('h44c4)
	) name2040 (
		_w793_,
		_w794_,
		_w791_,
		_w2297_,
		_w2298_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name2041 (
		_w438_,
		_w1074_,
		_w1075_,
		_w2298_,
		_w2299_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2042 (
		_w442_,
		_w449_,
		_w454_,
		_w2299_,
		_w2300_
	);
	LUT4 #(
		.INIT('h44c4)
	) name2043 (
		_w465_,
		_w473_,
		_w461_,
		_w2300_,
		_w2301_
	);
	LUT4 #(
		.INIT('h22a2)
	) name2044 (
		_w489_,
		_w484_,
		_w477_,
		_w2301_,
		_w2302_
	);
	LUT4 #(
		.INIT('h44c4)
	) name2045 (
		_w500_,
		_w508_,
		_w496_,
		_w2302_,
		_w2303_
	);
	LUT4 #(
		.INIT('h44c4)
	) name2046 (
		_w519_,
		_w524_,
		_w512_,
		_w2303_,
		_w2304_
	);
	LUT4 #(
		.INIT('hd000)
	) name2047 (
		_w533_,
		_w538_,
		_w542_,
		_w2293_,
		_w2305_
	);
	LUT4 #(
		.INIT('h7500)
	) name2048 (
		_w535_,
		_w2304_,
		_w531_,
		_w2305_,
		_w2306_
	);
	LUT2 #(
		.INIT('he)
	) name2049 (
		_w2294_,
		_w2306_,
		_w2307_
	);
	LUT3 #(
		.INIT('hb0)
	) name2050 (
		\priority[94] ,
		\req[93] ,
		\req[94] ,
		_w2308_
	);
	LUT2 #(
		.INIT('h4)
	) name2051 (
		_w710_,
		_w2308_,
		_w2309_
	);
	LUT3 #(
		.INIT('h31)
	) name2052 (
		\priority[95] ,
		\priority[96] ,
		\req[95] ,
		_w2310_
	);
	LUT4 #(
		.INIT('ha020)
	) name2053 (
		_w545_,
		_w548_,
		_w556_,
		_w2310_,
		_w2311_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2054 (
		_w831_,
		_w833_,
		_w834_,
		_w2311_,
		_w2312_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2055 (
		_w835_,
		_w837_,
		_w838_,
		_w2312_,
		_w2313_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name2056 (
		_w604_,
		_w1091_,
		_w1092_,
		_w2313_,
		_w2314_
	);
	LUT4 #(
		.INIT('h0c8c)
	) name2057 (
		_w608_,
		_w620_,
		_w615_,
		_w2314_,
		_w2315_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2058 (
		_w627_,
		_w631_,
		_w639_,
		_w2315_,
		_w2316_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2059 (
		_w643_,
		_w650_,
		_w655_,
		_w2316_,
		_w2317_
	);
	LUT4 #(
		.INIT('h4c44)
	) name2060 (
		_w666_,
		_w674_,
		_w2317_,
		_w662_,
		_w2318_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2061 (
		_w678_,
		_w685_,
		_w690_,
		_w2318_,
		_w2319_
	);
	LUT4 #(
		.INIT('hd000)
	) name2062 (
		_w699_,
		_w704_,
		_w708_,
		_w2308_,
		_w2320_
	);
	LUT4 #(
		.INIT('h3b00)
	) name2063 (
		_w697_,
		_w701_,
		_w2319_,
		_w2320_,
		_w2321_
	);
	LUT2 #(
		.INIT('he)
	) name2064 (
		_w2309_,
		_w2321_,
		_w2322_
	);
	LUT3 #(
		.INIT('hb0)
	) name2065 (
		\priority[95] ,
		\req[94] ,
		\req[95] ,
		_w2323_
	);
	LUT2 #(
		.INIT('h4)
	) name2066 (
		_w380_,
		_w2323_,
		_w2324_
	);
	LUT3 #(
		.INIT('h31)
	) name2067 (
		\priority[96] ,
		\priority[97] ,
		\req[96] ,
		_w2325_
	);
	LUT4 #(
		.INIT('ha020)
	) name2068 (
		_w711_,
		_w714_,
		_w722_,
		_w2325_,
		_w2326_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2069 (
		_w874_,
		_w876_,
		_w877_,
		_w2326_,
		_w2327_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2070 (
		_w878_,
		_w880_,
		_w881_,
		_w2327_,
		_w2328_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name2071 (
		_w761_,
		_w1108_,
		_w1109_,
		_w2328_,
		_w2329_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2072 (
		_w762_,
		_w763_,
		_w765_,
		_w2329_,
		_w2330_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2073 (
		_w766_,
		_w767_,
		_w769_,
		_w2330_,
		_w2331_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2074 (
		_w770_,
		_w771_,
		_w773_,
		_w2331_,
		_w2332_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2075 (
		_w774_,
		_w775_,
		_w777_,
		_w2332_,
		_w2333_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2076 (
		_w778_,
		_w779_,
		_w781_,
		_w2333_,
		_w2334_
	);
	LUT4 #(
		.INIT('h8a00)
	) name2077 (
		_w374_,
		_w376_,
		_w378_,
		_w2323_,
		_w2335_
	);
	LUT4 #(
		.INIT('h3b00)
	) name2078 (
		_w782_,
		_w783_,
		_w2334_,
		_w2335_,
		_w2336_
	);
	LUT2 #(
		.INIT('he)
	) name2079 (
		_w2324_,
		_w2336_,
		_w2337_
	);
	LUT3 #(
		.INIT('hb0)
	) name2080 (
		\priority[96] ,
		\req[95] ,
		\req[96] ,
		_w2338_
	);
	LUT2 #(
		.INIT('h4)
	) name2081 (
		_w546_,
		_w2338_,
		_w2339_
	);
	LUT3 #(
		.INIT('h31)
	) name2082 (
		\priority[97] ,
		\priority[98] ,
		\req[97] ,
		_w2340_
	);
	LUT4 #(
		.INIT('hc040)
	) name2083 (
		_w386_,
		_w390_,
		_w392_,
		_w2340_,
		_w2341_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2084 (
		_w916_,
		_w918_,
		_w919_,
		_w2341_,
		_w2342_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2085 (
		_w920_,
		_w922_,
		_w923_,
		_w2342_,
		_w2343_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name2086 (
		_w805_,
		_w1125_,
		_w1126_,
		_w2343_,
		_w2344_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2087 (
		_w806_,
		_w807_,
		_w809_,
		_w2344_,
		_w2345_
	);
	LUT4 #(
		.INIT('h0c8c)
	) name2088 (
		_w810_,
		_w813_,
		_w811_,
		_w2345_,
		_w2346_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2089 (
		_w814_,
		_w815_,
		_w817_,
		_w2346_,
		_w2347_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2090 (
		_w818_,
		_w819_,
		_w821_,
		_w2347_,
		_w2348_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2091 (
		_w822_,
		_w823_,
		_w825_,
		_w2348_,
		_w2349_
	);
	LUT4 #(
		.INIT('h8a00)
	) name2092 (
		_w540_,
		_w542_,
		_w544_,
		_w2338_,
		_w2350_
	);
	LUT4 #(
		.INIT('h3b00)
	) name2093 (
		_w826_,
		_w827_,
		_w2349_,
		_w2350_,
		_w2351_
	);
	LUT2 #(
		.INIT('he)
	) name2094 (
		_w2339_,
		_w2351_,
		_w2352_
	);
	LUT3 #(
		.INIT('hb0)
	) name2095 (
		\priority[97] ,
		\req[96] ,
		\req[97] ,
		_w2353_
	);
	LUT2 #(
		.INIT('h4)
	) name2096 (
		_w712_,
		_w2353_,
		_w2354_
	);
	LUT3 #(
		.INIT('h31)
	) name2097 (
		\priority[98] ,
		\priority[99] ,
		\req[98] ,
		_w2355_
	);
	LUT4 #(
		.INIT('hc040)
	) name2098 (
		_w552_,
		_w556_,
		_w558_,
		_w2355_,
		_w2356_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2099 (
		_w958_,
		_w960_,
		_w961_,
		_w2356_,
		_w2357_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2100 (
		_w962_,
		_w964_,
		_w965_,
		_w2357_,
		_w2358_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name2101 (
		_w848_,
		_w1142_,
		_w1143_,
		_w2358_,
		_w2359_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2102 (
		_w849_,
		_w850_,
		_w852_,
		_w2359_,
		_w2360_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2103 (
		_w853_,
		_w854_,
		_w856_,
		_w2360_,
		_w2361_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2104 (
		_w857_,
		_w858_,
		_w860_,
		_w2361_,
		_w2362_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2105 (
		_w861_,
		_w862_,
		_w864_,
		_w2362_,
		_w2363_
	);
	LUT4 #(
		.INIT('h0c8c)
	) name2106 (
		_w865_,
		_w868_,
		_w866_,
		_w2363_,
		_w2364_
	);
	LUT4 #(
		.INIT('h8a00)
	) name2107 (
		_w706_,
		_w708_,
		_w710_,
		_w2353_,
		_w2365_
	);
	LUT4 #(
		.INIT('h3b00)
	) name2108 (
		_w869_,
		_w870_,
		_w2364_,
		_w2365_,
		_w2366_
	);
	LUT2 #(
		.INIT('he)
	) name2109 (
		_w2354_,
		_w2366_,
		_w2367_
	);
	LUT3 #(
		.INIT('hb0)
	) name2110 (
		\priority[98] ,
		\req[97] ,
		\req[98] ,
		_w2368_
	);
	LUT2 #(
		.INIT('h4)
	) name2111 (
		_w379_,
		_w2368_,
		_w2369_
	);
	LUT3 #(
		.INIT('h31)
	) name2112 (
		\priority[99] ,
		\priority[100] ,
		\req[99] ,
		_w2370_
	);
	LUT4 #(
		.INIT('hc040)
	) name2113 (
		_w718_,
		_w722_,
		_w724_,
		_w2370_,
		_w2371_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2114 (
		_w1000_,
		_w1002_,
		_w1003_,
		_w2371_,
		_w2372_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2115 (
		_w1004_,
		_w1006_,
		_w1007_,
		_w2372_,
		_w2373_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name2116 (
		_w890_,
		_w1159_,
		_w1160_,
		_w2373_,
		_w2374_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2117 (
		_w891_,
		_w892_,
		_w894_,
		_w2374_,
		_w2375_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2118 (
		_w895_,
		_w896_,
		_w898_,
		_w2375_,
		_w2376_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2119 (
		_w899_,
		_w900_,
		_w902_,
		_w2376_,
		_w2377_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2120 (
		_w903_,
		_w904_,
		_w906_,
		_w2377_,
		_w2378_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2121 (
		_w907_,
		_w908_,
		_w910_,
		_w2378_,
		_w2379_
	);
	LUT4 #(
		.INIT('hb000)
	) name2122 (
		_w374_,
		_w380_,
		_w383_,
		_w2368_,
		_w2380_
	);
	LUT4 #(
		.INIT('h3b00)
	) name2123 (
		_w911_,
		_w912_,
		_w2379_,
		_w2380_,
		_w2381_
	);
	LUT2 #(
		.INIT('he)
	) name2124 (
		_w2369_,
		_w2381_,
		_w2382_
	);
	LUT3 #(
		.INIT('hb0)
	) name2125 (
		\priority[99] ,
		\req[98] ,
		\req[99] ,
		_w2383_
	);
	LUT2 #(
		.INIT('h4)
	) name2126 (
		_w545_,
		_w2383_,
		_w2384_
	);
	LUT3 #(
		.INIT('h31)
	) name2127 (
		\priority[100] ,
		\priority[101] ,
		\req[100] ,
		_w2385_
	);
	LUT4 #(
		.INIT('hc040)
	) name2128 (
		_w384_,
		_w391_,
		_w392_,
		_w2385_,
		_w2386_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2129 (
		_w400_,
		_w404_,
		_w412_,
		_w2386_,
		_w2387_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2130 (
		_w416_,
		_w1023_,
		_w1024_,
		_w2387_,
		_w2388_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name2131 (
		_w932_,
		_w1176_,
		_w1177_,
		_w2388_,
		_w2389_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2132 (
		_w933_,
		_w934_,
		_w936_,
		_w2389_,
		_w2390_
	);
	LUT4 #(
		.INIT('h44c4)
	) name2133 (
		_w938_,
		_w940_,
		_w937_,
		_w2390_,
		_w2391_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2134 (
		_w941_,
		_w942_,
		_w944_,
		_w2391_,
		_w2392_
	);
	LUT4 #(
		.INIT('h0c8c)
	) name2135 (
		_w945_,
		_w948_,
		_w946_,
		_w2392_,
		_w2393_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2136 (
		_w949_,
		_w950_,
		_w952_,
		_w2393_,
		_w2394_
	);
	LUT4 #(
		.INIT('hb000)
	) name2137 (
		_w540_,
		_w546_,
		_w549_,
		_w2383_,
		_w2395_
	);
	LUT4 #(
		.INIT('h3b00)
	) name2138 (
		_w953_,
		_w954_,
		_w2394_,
		_w2395_,
		_w2396_
	);
	LUT2 #(
		.INIT('he)
	) name2139 (
		_w2384_,
		_w2396_,
		_w2397_
	);
	LUT3 #(
		.INIT('hb0)
	) name2140 (
		\priority[100] ,
		\req[99] ,
		\req[100] ,
		_w2398_
	);
	LUT2 #(
		.INIT('h4)
	) name2141 (
		_w711_,
		_w2398_,
		_w2399_
	);
	LUT3 #(
		.INIT('h31)
	) name2142 (
		\priority[101] ,
		\priority[102] ,
		\req[101] ,
		_w2400_
	);
	LUT4 #(
		.INIT('hc040)
	) name2143 (
		_w550_,
		_w557_,
		_w558_,
		_w2400_,
		_w2401_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2144 (
		_w566_,
		_w570_,
		_w578_,
		_w2401_,
		_w2402_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2145 (
		_w582_,
		_w1040_,
		_w1041_,
		_w2402_,
		_w2403_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name2146 (
		_w974_,
		_w1193_,
		_w1194_,
		_w2403_,
		_w2404_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2147 (
		_w975_,
		_w976_,
		_w978_,
		_w2404_,
		_w2405_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2148 (
		_w979_,
		_w980_,
		_w982_,
		_w2405_,
		_w2406_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2149 (
		_w983_,
		_w984_,
		_w986_,
		_w2406_,
		_w2407_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2150 (
		_w987_,
		_w988_,
		_w990_,
		_w2407_,
		_w2408_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2151 (
		_w991_,
		_w992_,
		_w994_,
		_w2408_,
		_w2409_
	);
	LUT4 #(
		.INIT('hb000)
	) name2152 (
		_w706_,
		_w712_,
		_w715_,
		_w2398_,
		_w2410_
	);
	LUT4 #(
		.INIT('h3b00)
	) name2153 (
		_w995_,
		_w996_,
		_w2409_,
		_w2410_,
		_w2411_
	);
	LUT2 #(
		.INIT('he)
	) name2154 (
		_w2399_,
		_w2411_,
		_w2412_
	);
	LUT3 #(
		.INIT('hb0)
	) name2155 (
		\priority[101] ,
		\req[100] ,
		\req[101] ,
		_w2413_
	);
	LUT2 #(
		.INIT('h4)
	) name2156 (
		_w390_,
		_w2413_,
		_w2414_
	);
	LUT3 #(
		.INIT('h31)
	) name2157 (
		\priority[102] ,
		\priority[103] ,
		\req[102] ,
		_w2415_
	);
	LUT4 #(
		.INIT('hc040)
	) name2158 (
		_w716_,
		_w723_,
		_w724_,
		_w2415_,
		_w2416_
	);
	LUT4 #(
		.INIT('h0c8c)
	) name2159 (
		_w732_,
		_w744_,
		_w736_,
		_w2416_,
		_w2417_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2160 (
		_w748_,
		_w1057_,
		_w1058_,
		_w2417_,
		_w2418_
	);
	LUT4 #(
		.INIT('h08cc)
	) name2161 (
		_w272_,
		_w283_,
		_w2418_,
		_w276_,
		_w2419_
	);
	LUT4 #(
		.INIT('h3b00)
	) name2162 (
		_w288_,
		_w295_,
		_w2419_,
		_w299_,
		_w2420_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2163 (
		_w307_,
		_w311_,
		_w318_,
		_w2420_,
		_w2421_
	);
	LUT4 #(
		.INIT('h44c4)
	) name2164 (
		_w330_,
		_w334_,
		_w323_,
		_w2421_,
		_w2422_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2165 (
		_w342_,
		_w346_,
		_w353_,
		_w2422_,
		_w2423_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2166 (
		_w358_,
		_w365_,
		_w369_,
		_w2423_,
		_w2424_
	);
	LUT4 #(
		.INIT('hd000)
	) name2167 (
		_w379_,
		_w383_,
		_w387_,
		_w2413_,
		_w2425_
	);
	LUT4 #(
		.INIT('h3b00)
	) name2168 (
		_w377_,
		_w381_,
		_w2424_,
		_w2425_,
		_w2426_
	);
	LUT2 #(
		.INIT('he)
	) name2169 (
		_w2414_,
		_w2426_,
		_w2427_
	);
	LUT3 #(
		.INIT('hb0)
	) name2170 (
		\priority[102] ,
		\req[101] ,
		\req[102] ,
		_w2428_
	);
	LUT2 #(
		.INIT('h4)
	) name2171 (
		_w556_,
		_w2428_,
		_w2429_
	);
	LUT3 #(
		.INIT('h31)
	) name2172 (
		\priority[103] ,
		\priority[104] ,
		\req[103] ,
		_w2430_
	);
	LUT4 #(
		.INIT('ha020)
	) name2173 (
		_w391_,
		_w394_,
		_w401_,
		_w2430_,
		_w2431_
	);
	LUT4 #(
		.INIT('h0c8c)
	) name2174 (
		_w790_,
		_w793_,
		_w791_,
		_w2431_,
		_w2432_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2175 (
		_w794_,
		_w1074_,
		_w1075_,
		_w2432_,
		_w2433_
	);
	LUT4 #(
		.INIT('h4c44)
	) name2176 (
		_w442_,
		_w449_,
		_w2433_,
		_w438_,
		_w2434_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name2177 (
		_w465_,
		_w454_,
		_w461_,
		_w2434_,
		_w2435_
	);
	LUT4 #(
		.INIT('h0c8c)
	) name2178 (
		_w473_,
		_w484_,
		_w477_,
		_w2435_,
		_w2436_
	);
	LUT4 #(
		.INIT('h0c8c)
	) name2179 (
		_w489_,
		_w500_,
		_w496_,
		_w2436_,
		_w2437_
	);
	LUT4 #(
		.INIT('h0c8c)
	) name2180 (
		_w508_,
		_w519_,
		_w512_,
		_w2437_,
		_w2438_
	);
	LUT4 #(
		.INIT('h0c8c)
	) name2181 (
		_w524_,
		_w535_,
		_w531_,
		_w2438_,
		_w2439_
	);
	LUT4 #(
		.INIT('hd000)
	) name2182 (
		_w545_,
		_w549_,
		_w553_,
		_w2428_,
		_w2440_
	);
	LUT4 #(
		.INIT('h3b00)
	) name2183 (
		_w543_,
		_w547_,
		_w2439_,
		_w2440_,
		_w2441_
	);
	LUT2 #(
		.INIT('he)
	) name2184 (
		_w2429_,
		_w2441_,
		_w2442_
	);
	LUT3 #(
		.INIT('hb0)
	) name2185 (
		\priority[103] ,
		\req[102] ,
		\req[103] ,
		_w2443_
	);
	LUT2 #(
		.INIT('h4)
	) name2186 (
		_w722_,
		_w2443_,
		_w2444_
	);
	LUT3 #(
		.INIT('h31)
	) name2187 (
		\priority[104] ,
		\priority[105] ,
		\req[104] ,
		_w2445_
	);
	LUT4 #(
		.INIT('ha020)
	) name2188 (
		_w557_,
		_w560_,
		_w567_,
		_w2445_,
		_w2446_
	);
	LUT4 #(
		.INIT('h4c44)
	) name2189 (
		_w835_,
		_w837_,
		_w2446_,
		_w834_,
		_w2447_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2190 (
		_w838_,
		_w1091_,
		_w1092_,
		_w2447_,
		_w2448_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2191 (
		_w604_,
		_w608_,
		_w615_,
		_w2448_,
		_w2449_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2192 (
		_w620_,
		_w627_,
		_w631_,
		_w2449_,
		_w2450_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2193 (
		_w639_,
		_w643_,
		_w650_,
		_w2450_,
		_w2451_
	);
	LUT4 #(
		.INIT('h0c8c)
	) name2194 (
		_w655_,
		_w666_,
		_w662_,
		_w2451_,
		_w2452_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2195 (
		_w674_,
		_w678_,
		_w685_,
		_w2452_,
		_w2453_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2196 (
		_w690_,
		_w697_,
		_w701_,
		_w2453_,
		_w2454_
	);
	LUT4 #(
		.INIT('hd000)
	) name2197 (
		_w711_,
		_w715_,
		_w719_,
		_w2443_,
		_w2455_
	);
	LUT4 #(
		.INIT('h3b00)
	) name2198 (
		_w709_,
		_w713_,
		_w2454_,
		_w2455_,
		_w2456_
	);
	LUT2 #(
		.INIT('he)
	) name2199 (
		_w2444_,
		_w2456_,
		_w2457_
	);
	LUT3 #(
		.INIT('hb0)
	) name2200 (
		\priority[104] ,
		\req[103] ,
		\req[104] ,
		_w2458_
	);
	LUT2 #(
		.INIT('h4)
	) name2201 (
		_w392_,
		_w2458_,
		_w2459_
	);
	LUT3 #(
		.INIT('h31)
	) name2202 (
		\priority[105] ,
		\priority[106] ,
		\req[105] ,
		_w2460_
	);
	LUT4 #(
		.INIT('ha020)
	) name2203 (
		_w723_,
		_w726_,
		_w733_,
		_w2460_,
		_w2461_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2204 (
		_w877_,
		_w878_,
		_w880_,
		_w2461_,
		_w2462_
	);
	LUT4 #(
		.INIT('h44c4)
	) name2205 (
		_w1108_,
		_w1109_,
		_w881_,
		_w2462_,
		_w2463_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2206 (
		_w761_,
		_w762_,
		_w763_,
		_w2463_,
		_w2464_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2207 (
		_w765_,
		_w766_,
		_w767_,
		_w2464_,
		_w2465_
	);
	LUT4 #(
		.INIT('h3b00)
	) name2208 (
		_w769_,
		_w770_,
		_w2465_,
		_w771_,
		_w2466_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2209 (
		_w773_,
		_w774_,
		_w775_,
		_w2466_,
		_w2467_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2210 (
		_w777_,
		_w778_,
		_w779_,
		_w2467_,
		_w2468_
	);
	LUT4 #(
		.INIT('h3b00)
	) name2211 (
		_w781_,
		_w782_,
		_w2468_,
		_w783_,
		_w2469_
	);
	LUT4 #(
		.INIT('h8a00)
	) name2212 (
		_w385_,
		_w387_,
		_w390_,
		_w2458_,
		_w2470_
	);
	LUT4 #(
		.INIT('h3b00)
	) name2213 (
		_w785_,
		_w786_,
		_w2469_,
		_w2470_,
		_w2471_
	);
	LUT2 #(
		.INIT('he)
	) name2214 (
		_w2459_,
		_w2471_,
		_w2472_
	);
	LUT3 #(
		.INIT('hb0)
	) name2215 (
		\priority[105] ,
		\req[104] ,
		\req[105] ,
		_w2473_
	);
	LUT2 #(
		.INIT('h4)
	) name2216 (
		_w558_,
		_w2473_,
		_w2474_
	);
	LUT3 #(
		.INIT('h31)
	) name2217 (
		\priority[106] ,
		\priority[107] ,
		\req[106] ,
		_w2475_
	);
	LUT4 #(
		.INIT('hc040)
	) name2218 (
		_w398_,
		_w401_,
		_w403_,
		_w2475_,
		_w2476_
	);
	LUT4 #(
		.INIT('h44c4)
	) name2219 (
		_w920_,
		_w922_,
		_w919_,
		_w2476_,
		_w2477_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2220 (
		_w923_,
		_w1125_,
		_w1126_,
		_w2477_,
		_w2478_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2221 (
		_w805_,
		_w806_,
		_w807_,
		_w2478_,
		_w2479_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2222 (
		_w809_,
		_w810_,
		_w811_,
		_w2479_,
		_w2480_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2223 (
		_w813_,
		_w814_,
		_w815_,
		_w2480_,
		_w2481_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2224 (
		_w817_,
		_w818_,
		_w819_,
		_w2481_,
		_w2482_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2225 (
		_w821_,
		_w822_,
		_w823_,
		_w2482_,
		_w2483_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2226 (
		_w825_,
		_w826_,
		_w827_,
		_w2483_,
		_w2484_
	);
	LUT4 #(
		.INIT('h8a00)
	) name2227 (
		_w551_,
		_w553_,
		_w556_,
		_w2473_,
		_w2485_
	);
	LUT4 #(
		.INIT('h7500)
	) name2228 (
		_w830_,
		_w2484_,
		_w829_,
		_w2485_,
		_w2486_
	);
	LUT2 #(
		.INIT('he)
	) name2229 (
		_w2474_,
		_w2486_,
		_w2487_
	);
	LUT3 #(
		.INIT('hb0)
	) name2230 (
		\priority[106] ,
		\req[105] ,
		\req[106] ,
		_w2488_
	);
	LUT2 #(
		.INIT('h4)
	) name2231 (
		_w724_,
		_w2488_,
		_w2489_
	);
	LUT3 #(
		.INIT('h31)
	) name2232 (
		\priority[107] ,
		\priority[108] ,
		\req[107] ,
		_w2490_
	);
	LUT4 #(
		.INIT('hc040)
	) name2233 (
		_w564_,
		_w567_,
		_w569_,
		_w2490_,
		_w2491_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2234 (
		_w961_,
		_w962_,
		_w964_,
		_w2491_,
		_w2492_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2235 (
		_w965_,
		_w1142_,
		_w1143_,
		_w2492_,
		_w2493_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2236 (
		_w848_,
		_w849_,
		_w850_,
		_w2493_,
		_w2494_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2237 (
		_w852_,
		_w853_,
		_w854_,
		_w2494_,
		_w2495_
	);
	LUT4 #(
		.INIT('h3b00)
	) name2238 (
		_w856_,
		_w857_,
		_w2495_,
		_w858_,
		_w2496_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2239 (
		_w860_,
		_w861_,
		_w862_,
		_w2496_,
		_w2497_
	);
	LUT4 #(
		.INIT('h50d0)
	) name2240 (
		_w865_,
		_w864_,
		_w866_,
		_w2497_,
		_w2498_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2241 (
		_w868_,
		_w869_,
		_w870_,
		_w2498_,
		_w2499_
	);
	LUT4 #(
		.INIT('h8a00)
	) name2242 (
		_w717_,
		_w719_,
		_w722_,
		_w2488_,
		_w2500_
	);
	LUT4 #(
		.INIT('h3b00)
	) name2243 (
		_w872_,
		_w873_,
		_w2499_,
		_w2500_,
		_w2501_
	);
	LUT2 #(
		.INIT('he)
	) name2244 (
		_w2489_,
		_w2501_,
		_w2502_
	);
	LUT3 #(
		.INIT('hb0)
	) name2245 (
		\priority[107] ,
		\req[106] ,
		\req[107] ,
		_w2503_
	);
	LUT2 #(
		.INIT('h4)
	) name2246 (
		_w391_,
		_w2503_,
		_w2504_
	);
	LUT3 #(
		.INIT('h31)
	) name2247 (
		\priority[108] ,
		\priority[109] ,
		\req[108] ,
		_w2505_
	);
	LUT4 #(
		.INIT('hc040)
	) name2248 (
		_w730_,
		_w733_,
		_w735_,
		_w2505_,
		_w2506_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2249 (
		_w1003_,
		_w1004_,
		_w1006_,
		_w2506_,
		_w2507_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2250 (
		_w1007_,
		_w1159_,
		_w1160_,
		_w2507_,
		_w2508_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2251 (
		_w890_,
		_w891_,
		_w892_,
		_w2508_,
		_w2509_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2252 (
		_w894_,
		_w895_,
		_w896_,
		_w2509_,
		_w2510_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2253 (
		_w898_,
		_w899_,
		_w900_,
		_w2510_,
		_w2511_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2254 (
		_w902_,
		_w903_,
		_w904_,
		_w2511_,
		_w2512_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2255 (
		_w906_,
		_w907_,
		_w908_,
		_w2512_,
		_w2513_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2256 (
		_w910_,
		_w911_,
		_w912_,
		_w2513_,
		_w2514_
	);
	LUT4 #(
		.INIT('hb000)
	) name2257 (
		_w385_,
		_w392_,
		_w395_,
		_w2503_,
		_w2515_
	);
	LUT4 #(
		.INIT('h5d00)
	) name2258 (
		_w915_,
		_w914_,
		_w2514_,
		_w2515_,
		_w2516_
	);
	LUT2 #(
		.INIT('he)
	) name2259 (
		_w2504_,
		_w2516_,
		_w2517_
	);
	LUT3 #(
		.INIT('hb0)
	) name2260 (
		\priority[108] ,
		\req[107] ,
		\req[108] ,
		_w2518_
	);
	LUT2 #(
		.INIT('h4)
	) name2261 (
		_w557_,
		_w2518_,
		_w2519_
	);
	LUT3 #(
		.INIT('h31)
	) name2262 (
		\priority[109] ,
		\priority[110] ,
		\req[109] ,
		_w2520_
	);
	LUT4 #(
		.INIT('hc040)
	) name2263 (
		_w396_,
		_w402_,
		_w403_,
		_w2520_,
		_w2521_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2264 (
		_w412_,
		_w416_,
		_w1023_,
		_w2521_,
		_w2522_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2265 (
		_w1024_,
		_w1176_,
		_w1177_,
		_w2522_,
		_w2523_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2266 (
		_w932_,
		_w933_,
		_w934_,
		_w2523_,
		_w2524_
	);
	LUT4 #(
		.INIT('h0c8c)
	) name2267 (
		_w936_,
		_w938_,
		_w937_,
		_w2524_,
		_w2525_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2268 (
		_w940_,
		_w941_,
		_w942_,
		_w2525_,
		_w2526_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2269 (
		_w944_,
		_w945_,
		_w946_,
		_w2526_,
		_w2527_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2270 (
		_w948_,
		_w949_,
		_w950_,
		_w2527_,
		_w2528_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2271 (
		_w952_,
		_w953_,
		_w954_,
		_w2528_,
		_w2529_
	);
	LUT4 #(
		.INIT('hb000)
	) name2272 (
		_w551_,
		_w558_,
		_w561_,
		_w2518_,
		_w2530_
	);
	LUT4 #(
		.INIT('h3b00)
	) name2273 (
		_w956_,
		_w957_,
		_w2529_,
		_w2530_,
		_w2531_
	);
	LUT2 #(
		.INIT('he)
	) name2274 (
		_w2519_,
		_w2531_,
		_w2532_
	);
	LUT3 #(
		.INIT('hb0)
	) name2275 (
		\priority[109] ,
		\req[108] ,
		\req[109] ,
		_w2533_
	);
	LUT2 #(
		.INIT('h4)
	) name2276 (
		_w723_,
		_w2533_,
		_w2534_
	);
	LUT3 #(
		.INIT('h31)
	) name2277 (
		\priority[110] ,
		\priority[111] ,
		\req[110] ,
		_w2535_
	);
	LUT4 #(
		.INIT('hc040)
	) name2278 (
		_w562_,
		_w568_,
		_w569_,
		_w2535_,
		_w2536_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2279 (
		_w578_,
		_w582_,
		_w1040_,
		_w2536_,
		_w2537_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2280 (
		_w1041_,
		_w1193_,
		_w1194_,
		_w2537_,
		_w2538_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2281 (
		_w974_,
		_w975_,
		_w976_,
		_w2538_,
		_w2539_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2282 (
		_w978_,
		_w979_,
		_w980_,
		_w2539_,
		_w2540_
	);
	LUT4 #(
		.INIT('h44c4)
	) name2283 (
		_w983_,
		_w984_,
		_w982_,
		_w2540_,
		_w2541_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2284 (
		_w986_,
		_w987_,
		_w988_,
		_w2541_,
		_w2542_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2285 (
		_w990_,
		_w991_,
		_w992_,
		_w2542_,
		_w2543_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2286 (
		_w994_,
		_w995_,
		_w996_,
		_w2543_,
		_w2544_
	);
	LUT4 #(
		.INIT('hb000)
	) name2287 (
		_w717_,
		_w724_,
		_w727_,
		_w2533_,
		_w2545_
	);
	LUT4 #(
		.INIT('h3b00)
	) name2288 (
		_w998_,
		_w999_,
		_w2544_,
		_w2545_,
		_w2546_
	);
	LUT2 #(
		.INIT('he)
	) name2289 (
		_w2534_,
		_w2546_,
		_w2547_
	);
	LUT3 #(
		.INIT('hb0)
	) name2290 (
		\priority[110] ,
		\req[109] ,
		\req[110] ,
		_w2548_
	);
	LUT2 #(
		.INIT('h4)
	) name2291 (
		_w401_,
		_w2548_,
		_w2549_
	);
	LUT3 #(
		.INIT('h31)
	) name2292 (
		\priority[111] ,
		\priority[112] ,
		\req[111] ,
		_w2550_
	);
	LUT4 #(
		.INIT('hc040)
	) name2293 (
		_w728_,
		_w734_,
		_w735_,
		_w2550_,
		_w2551_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2294 (
		_w744_,
		_w748_,
		_w1057_,
		_w2551_,
		_w2552_
	);
	LUT4 #(
		.INIT('h50d0)
	) name2295 (
		_w272_,
		_w1058_,
		_w276_,
		_w2552_,
		_w2553_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2296 (
		_w283_,
		_w288_,
		_w295_,
		_w2553_,
		_w2554_
	);
	LUT4 #(
		.INIT('h44c4)
	) name2297 (
		_w307_,
		_w311_,
		_w299_,
		_w2554_,
		_w2555_
	);
	LUT4 #(
		.INIT('h08cc)
	) name2298 (
		_w318_,
		_w330_,
		_w2555_,
		_w323_,
		_w2556_
	);
	LUT4 #(
		.INIT('h44c4)
	) name2299 (
		_w342_,
		_w346_,
		_w334_,
		_w2556_,
		_w2557_
	);
	LUT4 #(
		.INIT('h08cc)
	) name2300 (
		_w353_,
		_w365_,
		_w2557_,
		_w358_,
		_w2558_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2301 (
		_w369_,
		_w377_,
		_w381_,
		_w2558_,
		_w2559_
	);
	LUT4 #(
		.INIT('hd000)
	) name2302 (
		_w391_,
		_w395_,
		_w399_,
		_w2548_,
		_w2560_
	);
	LUT4 #(
		.INIT('h3b00)
	) name2303 (
		_w388_,
		_w393_,
		_w2559_,
		_w2560_,
		_w2561_
	);
	LUT2 #(
		.INIT('he)
	) name2304 (
		_w2549_,
		_w2561_,
		_w2562_
	);
	LUT3 #(
		.INIT('hb0)
	) name2305 (
		\priority[111] ,
		\req[110] ,
		\req[111] ,
		_w2563_
	);
	LUT2 #(
		.INIT('h4)
	) name2306 (
		_w567_,
		_w2563_,
		_w2564_
	);
	LUT3 #(
		.INIT('h31)
	) name2307 (
		\priority[112] ,
		\priority[113] ,
		\req[112] ,
		_w2565_
	);
	LUT4 #(
		.INIT('ha020)
	) name2308 (
		_w402_,
		_w406_,
		_w413_,
		_w2565_,
		_w2566_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2309 (
		_w793_,
		_w794_,
		_w1074_,
		_w2566_,
		_w2567_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name2310 (
		_w442_,
		_w1075_,
		_w438_,
		_w2567_,
		_w2568_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2311 (
		_w449_,
		_w454_,
		_w461_,
		_w2568_,
		_w2569_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2312 (
		_w465_,
		_w473_,
		_w477_,
		_w2569_,
		_w2570_
	);
	LUT4 #(
		.INIT('h50d0)
	) name2313 (
		_w489_,
		_w484_,
		_w496_,
		_w2570_,
		_w2571_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2314 (
		_w500_,
		_w508_,
		_w512_,
		_w2571_,
		_w2572_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2315 (
		_w519_,
		_w524_,
		_w531_,
		_w2572_,
		_w2573_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2316 (
		_w535_,
		_w543_,
		_w547_,
		_w2573_,
		_w2574_
	);
	LUT4 #(
		.INIT('hd000)
	) name2317 (
		_w557_,
		_w561_,
		_w565_,
		_w2563_,
		_w2575_
	);
	LUT4 #(
		.INIT('h3b00)
	) name2318 (
		_w554_,
		_w559_,
		_w2574_,
		_w2575_,
		_w2576_
	);
	LUT2 #(
		.INIT('he)
	) name2319 (
		_w2564_,
		_w2576_,
		_w2577_
	);
	LUT3 #(
		.INIT('hb0)
	) name2320 (
		\priority[112] ,
		\req[111] ,
		\req[112] ,
		_w2578_
	);
	LUT2 #(
		.INIT('h4)
	) name2321 (
		_w733_,
		_w2578_,
		_w2579_
	);
	LUT3 #(
		.INIT('h31)
	) name2322 (
		\priority[113] ,
		\priority[114] ,
		\req[113] ,
		_w2580_
	);
	LUT4 #(
		.INIT('ha020)
	) name2323 (
		_w568_,
		_w572_,
		_w579_,
		_w2580_,
		_w2581_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2324 (
		_w837_,
		_w838_,
		_w1091_,
		_w2581_,
		_w2582_
	);
	LUT4 #(
		.INIT('h44c4)
	) name2325 (
		_w604_,
		_w608_,
		_w1092_,
		_w2582_,
		_w2583_
	);
	LUT4 #(
		.INIT('h44c4)
	) name2326 (
		_w620_,
		_w627_,
		_w615_,
		_w2583_,
		_w2584_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2327 (
		_w631_,
		_w639_,
		_w643_,
		_w2584_,
		_w2585_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2328 (
		_w650_,
		_w655_,
		_w662_,
		_w2585_,
		_w2586_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2329 (
		_w666_,
		_w674_,
		_w678_,
		_w2586_,
		_w2587_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2330 (
		_w685_,
		_w690_,
		_w697_,
		_w2587_,
		_w2588_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2331 (
		_w701_,
		_w709_,
		_w713_,
		_w2588_,
		_w2589_
	);
	LUT4 #(
		.INIT('hd000)
	) name2332 (
		_w723_,
		_w727_,
		_w731_,
		_w2578_,
		_w2590_
	);
	LUT4 #(
		.INIT('h3b00)
	) name2333 (
		_w720_,
		_w725_,
		_w2589_,
		_w2590_,
		_w2591_
	);
	LUT2 #(
		.INIT('he)
	) name2334 (
		_w2579_,
		_w2591_,
		_w2592_
	);
	LUT3 #(
		.INIT('hb0)
	) name2335 (
		\priority[113] ,
		\req[112] ,
		\req[113] ,
		_w2593_
	);
	LUT2 #(
		.INIT('h4)
	) name2336 (
		_w403_,
		_w2593_,
		_w2594_
	);
	LUT3 #(
		.INIT('h31)
	) name2337 (
		\priority[114] ,
		\priority[115] ,
		\req[114] ,
		_w2595_
	);
	LUT4 #(
		.INIT('ha020)
	) name2338 (
		_w734_,
		_w738_,
		_w745_,
		_w2595_,
		_w2596_
	);
	LUT4 #(
		.INIT('h0c8c)
	) name2339 (
		_w880_,
		_w1108_,
		_w881_,
		_w2596_,
		_w2597_
	);
	LUT4 #(
		.INIT('h44c4)
	) name2340 (
		_w761_,
		_w762_,
		_w1109_,
		_w2597_,
		_w2598_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2341 (
		_w763_,
		_w765_,
		_w766_,
		_w2598_,
		_w2599_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2342 (
		_w767_,
		_w769_,
		_w770_,
		_w2599_,
		_w2600_
	);
	LUT4 #(
		.INIT('h44c4)
	) name2343 (
		_w773_,
		_w774_,
		_w771_,
		_w2600_,
		_w2601_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2344 (
		_w775_,
		_w777_,
		_w778_,
		_w2601_,
		_w2602_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2345 (
		_w779_,
		_w781_,
		_w782_,
		_w2602_,
		_w2603_
	);
	LUT4 #(
		.INIT('h44c4)
	) name2346 (
		_w785_,
		_w786_,
		_w783_,
		_w2603_,
		_w2604_
	);
	LUT4 #(
		.INIT('h8a00)
	) name2347 (
		_w397_,
		_w399_,
		_w401_,
		_w2593_,
		_w2605_
	);
	LUT4 #(
		.INIT('h3b00)
	) name2348 (
		_w787_,
		_w789_,
		_w2604_,
		_w2605_,
		_w2606_
	);
	LUT2 #(
		.INIT('he)
	) name2349 (
		_w2594_,
		_w2606_,
		_w2607_
	);
	LUT3 #(
		.INIT('hb0)
	) name2350 (
		\priority[114] ,
		\req[113] ,
		\req[114] ,
		_w2608_
	);
	LUT2 #(
		.INIT('h4)
	) name2351 (
		_w569_,
		_w2608_,
		_w2609_
	);
	LUT3 #(
		.INIT('h31)
	) name2352 (
		\priority[115] ,
		\priority[116] ,
		\req[115] ,
		_w2610_
	);
	LUT4 #(
		.INIT('hc040)
	) name2353 (
		_w410_,
		_w413_,
		_w415_,
		_w2610_,
		_w2611_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2354 (
		_w922_,
		_w923_,
		_w1125_,
		_w2611_,
		_w2612_
	);
	LUT4 #(
		.INIT('h44c4)
	) name2355 (
		_w805_,
		_w806_,
		_w1126_,
		_w2612_,
		_w2613_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2356 (
		_w807_,
		_w809_,
		_w810_,
		_w2613_,
		_w2614_
	);
	LUT4 #(
		.INIT('h44c4)
	) name2357 (
		_w813_,
		_w814_,
		_w811_,
		_w2614_,
		_w2615_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2358 (
		_w815_,
		_w817_,
		_w818_,
		_w2615_,
		_w2616_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2359 (
		_w819_,
		_w821_,
		_w822_,
		_w2616_,
		_w2617_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2360 (
		_w823_,
		_w825_,
		_w826_,
		_w2617_,
		_w2618_
	);
	LUT4 #(
		.INIT('h0c8c)
	) name2361 (
		_w827_,
		_w830_,
		_w829_,
		_w2618_,
		_w2619_
	);
	LUT4 #(
		.INIT('h8a00)
	) name2362 (
		_w563_,
		_w565_,
		_w567_,
		_w2608_,
		_w2620_
	);
	LUT4 #(
		.INIT('h2f00)
	) name2363 (
		_w831_,
		_w2619_,
		_w833_,
		_w2620_,
		_w2621_
	);
	LUT2 #(
		.INIT('he)
	) name2364 (
		_w2609_,
		_w2621_,
		_w2622_
	);
	LUT3 #(
		.INIT('hb0)
	) name2365 (
		\priority[115] ,
		\req[114] ,
		\req[115] ,
		_w2623_
	);
	LUT2 #(
		.INIT('h4)
	) name2366 (
		_w735_,
		_w2623_,
		_w2624_
	);
	LUT3 #(
		.INIT('h31)
	) name2367 (
		\priority[116] ,
		\priority[117] ,
		\req[116] ,
		_w2625_
	);
	LUT4 #(
		.INIT('hc040)
	) name2368 (
		_w576_,
		_w579_,
		_w581_,
		_w2625_,
		_w2626_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2369 (
		_w964_,
		_w965_,
		_w1142_,
		_w2626_,
		_w2627_
	);
	LUT4 #(
		.INIT('h44c4)
	) name2370 (
		_w848_,
		_w849_,
		_w1143_,
		_w2627_,
		_w2628_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2371 (
		_w850_,
		_w852_,
		_w853_,
		_w2628_,
		_w2629_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2372 (
		_w854_,
		_w856_,
		_w857_,
		_w2629_,
		_w2630_
	);
	LUT4 #(
		.INIT('h44c4)
	) name2373 (
		_w860_,
		_w861_,
		_w858_,
		_w2630_,
		_w2631_
	);
	LUT4 #(
		.INIT('h0c8c)
	) name2374 (
		_w862_,
		_w865_,
		_w864_,
		_w2631_,
		_w2632_
	);
	LUT4 #(
		.INIT('h44c4)
	) name2375 (
		_w868_,
		_w869_,
		_w866_,
		_w2632_,
		_w2633_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2376 (
		_w870_,
		_w872_,
		_w873_,
		_w2633_,
		_w2634_
	);
	LUT4 #(
		.INIT('h8a00)
	) name2377 (
		_w729_,
		_w731_,
		_w733_,
		_w2623_,
		_w2635_
	);
	LUT4 #(
		.INIT('h3b00)
	) name2378 (
		_w874_,
		_w876_,
		_w2634_,
		_w2635_,
		_w2636_
	);
	LUT2 #(
		.INIT('he)
	) name2379 (
		_w2624_,
		_w2636_,
		_w2637_
	);
	LUT3 #(
		.INIT('hb0)
	) name2380 (
		\priority[116] ,
		\req[115] ,
		\req[116] ,
		_w2638_
	);
	LUT2 #(
		.INIT('h4)
	) name2381 (
		_w402_,
		_w2638_,
		_w2639_
	);
	LUT3 #(
		.INIT('h31)
	) name2382 (
		\priority[117] ,
		\priority[118] ,
		\req[117] ,
		_w2640_
	);
	LUT4 #(
		.INIT('hc040)
	) name2383 (
		_w742_,
		_w745_,
		_w747_,
		_w2640_,
		_w2641_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2384 (
		_w1006_,
		_w1007_,
		_w1159_,
		_w2641_,
		_w2642_
	);
	LUT4 #(
		.INIT('h44c4)
	) name2385 (
		_w890_,
		_w891_,
		_w1160_,
		_w2642_,
		_w2643_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2386 (
		_w892_,
		_w894_,
		_w895_,
		_w2643_,
		_w2644_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2387 (
		_w896_,
		_w898_,
		_w899_,
		_w2644_,
		_w2645_
	);
	LUT4 #(
		.INIT('h3b00)
	) name2388 (
		_w900_,
		_w902_,
		_w2645_,
		_w903_,
		_w2646_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2389 (
		_w904_,
		_w906_,
		_w907_,
		_w2646_,
		_w2647_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2390 (
		_w908_,
		_w910_,
		_w911_,
		_w2647_,
		_w2648_
	);
	LUT4 #(
		.INIT('h2a22)
	) name2391 (
		_w915_,
		_w914_,
		_w2648_,
		_w912_,
		_w2649_
	);
	LUT4 #(
		.INIT('hb000)
	) name2392 (
		_w397_,
		_w403_,
		_w407_,
		_w2638_,
		_w2650_
	);
	LUT4 #(
		.INIT('h3b00)
	) name2393 (
		_w916_,
		_w918_,
		_w2649_,
		_w2650_,
		_w2651_
	);
	LUT2 #(
		.INIT('he)
	) name2394 (
		_w2639_,
		_w2651_,
		_w2652_
	);
	LUT3 #(
		.INIT('hb0)
	) name2395 (
		\priority[117] ,
		\req[116] ,
		\req[117] ,
		_w2653_
	);
	LUT2 #(
		.INIT('h4)
	) name2396 (
		_w568_,
		_w2653_,
		_w2654_
	);
	LUT3 #(
		.INIT('h31)
	) name2397 (
		\priority[118] ,
		\priority[119] ,
		\req[118] ,
		_w2655_
	);
	LUT4 #(
		.INIT('hc040)
	) name2398 (
		_w408_,
		_w414_,
		_w415_,
		_w2655_,
		_w2656_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2399 (
		_w1023_,
		_w1024_,
		_w1176_,
		_w2656_,
		_w2657_
	);
	LUT4 #(
		.INIT('h44c4)
	) name2400 (
		_w932_,
		_w933_,
		_w1177_,
		_w2657_,
		_w2658_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2401 (
		_w934_,
		_w936_,
		_w937_,
		_w2658_,
		_w2659_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2402 (
		_w938_,
		_w940_,
		_w941_,
		_w2659_,
		_w2660_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2403 (
		_w942_,
		_w944_,
		_w945_,
		_w2660_,
		_w2661_
	);
	LUT4 #(
		.INIT('h44c4)
	) name2404 (
		_w948_,
		_w949_,
		_w946_,
		_w2661_,
		_w2662_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2405 (
		_w950_,
		_w952_,
		_w953_,
		_w2662_,
		_w2663_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2406 (
		_w954_,
		_w956_,
		_w957_,
		_w2663_,
		_w2664_
	);
	LUT4 #(
		.INIT('hb000)
	) name2407 (
		_w563_,
		_w569_,
		_w573_,
		_w2653_,
		_w2665_
	);
	LUT4 #(
		.INIT('h7500)
	) name2408 (
		_w960_,
		_w2664_,
		_w958_,
		_w2665_,
		_w2666_
	);
	LUT2 #(
		.INIT('he)
	) name2409 (
		_w2654_,
		_w2666_,
		_w2667_
	);
	LUT3 #(
		.INIT('hb0)
	) name2410 (
		\priority[118] ,
		\req[117] ,
		\req[118] ,
		_w2668_
	);
	LUT2 #(
		.INIT('h4)
	) name2411 (
		_w734_,
		_w2668_,
		_w2669_
	);
	LUT3 #(
		.INIT('h31)
	) name2412 (
		\priority[119] ,
		\priority[120] ,
		\req[119] ,
		_w2670_
	);
	LUT4 #(
		.INIT('hc040)
	) name2413 (
		_w574_,
		_w580_,
		_w581_,
		_w2670_,
		_w2671_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2414 (
		_w1040_,
		_w1041_,
		_w1193_,
		_w2671_,
		_w2672_
	);
	LUT4 #(
		.INIT('h44c4)
	) name2415 (
		_w974_,
		_w975_,
		_w1194_,
		_w2672_,
		_w2673_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2416 (
		_w976_,
		_w978_,
		_w979_,
		_w2673_,
		_w2674_
	);
	LUT4 #(
		.INIT('h0c8c)
	) name2417 (
		_w980_,
		_w983_,
		_w982_,
		_w2674_,
		_w2675_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2418 (
		_w984_,
		_w986_,
		_w987_,
		_w2675_,
		_w2676_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2419 (
		_w988_,
		_w990_,
		_w991_,
		_w2676_,
		_w2677_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2420 (
		_w992_,
		_w994_,
		_w995_,
		_w2677_,
		_w2678_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2421 (
		_w996_,
		_w998_,
		_w999_,
		_w2678_,
		_w2679_
	);
	LUT4 #(
		.INIT('hb000)
	) name2422 (
		_w729_,
		_w735_,
		_w739_,
		_w2668_,
		_w2680_
	);
	LUT4 #(
		.INIT('h3b00)
	) name2423 (
		_w1000_,
		_w1002_,
		_w2679_,
		_w2680_,
		_w2681_
	);
	LUT2 #(
		.INIT('he)
	) name2424 (
		_w2669_,
		_w2681_,
		_w2682_
	);
	LUT3 #(
		.INIT('hb0)
	) name2425 (
		\priority[119] ,
		\req[118] ,
		\req[119] ,
		_w2683_
	);
	LUT2 #(
		.INIT('h4)
	) name2426 (
		_w413_,
		_w2683_,
		_w2684_
	);
	LUT3 #(
		.INIT('h31)
	) name2427 (
		\priority[120] ,
		\priority[121] ,
		\req[120] ,
		_w2685_
	);
	LUT4 #(
		.INIT('hc040)
	) name2428 (
		_w740_,
		_w746_,
		_w747_,
		_w2685_,
		_w2686_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name2429 (
		_w272_,
		_w1057_,
		_w1058_,
		_w2686_,
		_w2687_
	);
	LUT4 #(
		.INIT('h44c4)
	) name2430 (
		_w283_,
		_w288_,
		_w276_,
		_w2687_,
		_w2688_
	);
	LUT4 #(
		.INIT('h0c8c)
	) name2431 (
		_w295_,
		_w307_,
		_w299_,
		_w2688_,
		_w2689_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2432 (
		_w311_,
		_w318_,
		_w323_,
		_w2689_,
		_w2690_
	);
	LUT4 #(
		.INIT('h3b00)
	) name2433 (
		_w330_,
		_w334_,
		_w2690_,
		_w342_,
		_w2691_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2434 (
		_w346_,
		_w353_,
		_w358_,
		_w2691_,
		_w2692_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2435 (
		_w365_,
		_w369_,
		_w377_,
		_w2692_,
		_w2693_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2436 (
		_w381_,
		_w388_,
		_w393_,
		_w2693_,
		_w2694_
	);
	LUT4 #(
		.INIT('hd000)
	) name2437 (
		_w402_,
		_w407_,
		_w411_,
		_w2683_,
		_w2695_
	);
	LUT4 #(
		.INIT('h3b00)
	) name2438 (
		_w400_,
		_w404_,
		_w2694_,
		_w2695_,
		_w2696_
	);
	LUT2 #(
		.INIT('he)
	) name2439 (
		_w2684_,
		_w2696_,
		_w2697_
	);
	LUT3 #(
		.INIT('hb0)
	) name2440 (
		\priority[120] ,
		\req[119] ,
		\req[120] ,
		_w2698_
	);
	LUT2 #(
		.INIT('h4)
	) name2441 (
		_w579_,
		_w2698_,
		_w2699_
	);
	LUT3 #(
		.INIT('h31)
	) name2442 (
		\priority[121] ,
		\priority[122] ,
		\req[121] ,
		_w2700_
	);
	LUT4 #(
		.INIT('h8808)
	) name2443 (
		_w258_,
		_w414_,
		_w417_,
		_w2700_,
		_w2701_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2444 (
		_w1074_,
		_w1075_,
		_w438_,
		_w2701_,
		_w2702_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2445 (
		_w442_,
		_w449_,
		_w454_,
		_w2702_,
		_w2703_
	);
	LUT4 #(
		.INIT('h44c4)
	) name2446 (
		_w465_,
		_w473_,
		_w461_,
		_w2703_,
		_w2704_
	);
	LUT4 #(
		.INIT('h22a2)
	) name2447 (
		_w489_,
		_w484_,
		_w477_,
		_w2704_,
		_w2705_
	);
	LUT4 #(
		.INIT('h44c4)
	) name2448 (
		_w500_,
		_w508_,
		_w496_,
		_w2705_,
		_w2706_
	);
	LUT4 #(
		.INIT('h44c4)
	) name2449 (
		_w519_,
		_w524_,
		_w512_,
		_w2706_,
		_w2707_
	);
	LUT4 #(
		.INIT('h5d00)
	) name2450 (
		_w535_,
		_w531_,
		_w2707_,
		_w543_,
		_w2708_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2451 (
		_w547_,
		_w554_,
		_w559_,
		_w2708_,
		_w2709_
	);
	LUT4 #(
		.INIT('hd000)
	) name2452 (
		_w568_,
		_w573_,
		_w577_,
		_w2698_,
		_w2710_
	);
	LUT4 #(
		.INIT('h3b00)
	) name2453 (
		_w566_,
		_w570_,
		_w2709_,
		_w2710_,
		_w2711_
	);
	LUT2 #(
		.INIT('he)
	) name2454 (
		_w2699_,
		_w2711_,
		_w2712_
	);
	LUT3 #(
		.INIT('hb0)
	) name2455 (
		\priority[121] ,
		\req[120] ,
		\req[121] ,
		_w2713_
	);
	LUT2 #(
		.INIT('h4)
	) name2456 (
		_w745_,
		_w2713_,
		_w2714_
	);
	LUT3 #(
		.INIT('h31)
	) name2457 (
		\priority[122] ,
		\priority[123] ,
		\req[122] ,
		_w2715_
	);
	LUT4 #(
		.INIT('h8808)
	) name2458 (
		_w424_,
		_w580_,
		_w583_,
		_w2715_,
		_w2716_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name2459 (
		_w604_,
		_w1091_,
		_w1092_,
		_w2716_,
		_w2717_
	);
	LUT4 #(
		.INIT('h0c8c)
	) name2460 (
		_w608_,
		_w620_,
		_w615_,
		_w2717_,
		_w2718_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2461 (
		_w627_,
		_w631_,
		_w639_,
		_w2718_,
		_w2719_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2462 (
		_w643_,
		_w650_,
		_w655_,
		_w2719_,
		_w2720_
	);
	LUT4 #(
		.INIT('h44c4)
	) name2463 (
		_w666_,
		_w674_,
		_w662_,
		_w2720_,
		_w2721_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2464 (
		_w678_,
		_w685_,
		_w690_,
		_w2721_,
		_w2722_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2465 (
		_w697_,
		_w701_,
		_w709_,
		_w2722_,
		_w2723_
	);
	LUT4 #(
		.INIT('h44c4)
	) name2466 (
		_w720_,
		_w725_,
		_w713_,
		_w2723_,
		_w2724_
	);
	LUT4 #(
		.INIT('hd000)
	) name2467 (
		_w734_,
		_w739_,
		_w743_,
		_w2713_,
		_w2725_
	);
	LUT4 #(
		.INIT('h3b00)
	) name2468 (
		_w732_,
		_w736_,
		_w2724_,
		_w2725_,
		_w2726_
	);
	LUT2 #(
		.INIT('he)
	) name2469 (
		_w2714_,
		_w2726_,
		_w2727_
	);
	LUT3 #(
		.INIT('hb0)
	) name2470 (
		\priority[122] ,
		\req[121] ,
		\req[122] ,
		_w2728_
	);
	LUT2 #(
		.INIT('h4)
	) name2471 (
		_w415_,
		_w2728_,
		_w2729_
	);
	LUT3 #(
		.INIT('h31)
	) name2472 (
		\priority[123] ,
		\priority[124] ,
		\req[123] ,
		_w2730_
	);
	LUT4 #(
		.INIT('h8808)
	) name2473 (
		_w590_,
		_w746_,
		_w749_,
		_w2730_,
		_w2731_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name2474 (
		_w761_,
		_w1108_,
		_w1109_,
		_w2731_,
		_w2732_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2475 (
		_w762_,
		_w763_,
		_w765_,
		_w2732_,
		_w2733_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2476 (
		_w766_,
		_w767_,
		_w769_,
		_w2733_,
		_w2734_
	);
	LUT4 #(
		.INIT('h0c8c)
	) name2477 (
		_w770_,
		_w773_,
		_w771_,
		_w2734_,
		_w2735_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2478 (
		_w774_,
		_w775_,
		_w777_,
		_w2735_,
		_w2736_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2479 (
		_w778_,
		_w779_,
		_w781_,
		_w2736_,
		_w2737_
	);
	LUT4 #(
		.INIT('h0c8c)
	) name2480 (
		_w782_,
		_w785_,
		_w783_,
		_w2737_,
		_w2738_
	);
	LUT4 #(
		.INIT('h44c4)
	) name2481 (
		_w787_,
		_w789_,
		_w786_,
		_w2738_,
		_w2739_
	);
	LUT4 #(
		.INIT('h8a00)
	) name2482 (
		_w409_,
		_w411_,
		_w413_,
		_w2728_,
		_w2740_
	);
	LUT4 #(
		.INIT('h3b00)
	) name2483 (
		_w790_,
		_w791_,
		_w2739_,
		_w2740_,
		_w2741_
	);
	LUT2 #(
		.INIT('he)
	) name2484 (
		_w2729_,
		_w2741_,
		_w2742_
	);
	LUT3 #(
		.INIT('hb0)
	) name2485 (
		\priority[123] ,
		\req[122] ,
		\req[123] ,
		_w2743_
	);
	LUT2 #(
		.INIT('h4)
	) name2486 (
		_w581_,
		_w2743_,
		_w2744_
	);
	LUT3 #(
		.INIT('h31)
	) name2487 (
		\priority[124] ,
		\priority[125] ,
		\req[124] ,
		_w2745_
	);
	LUT4 #(
		.INIT('ha020)
	) name2488 (
		_w258_,
		_w419_,
		_w756_,
		_w2745_,
		_w2746_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name2489 (
		_w805_,
		_w1125_,
		_w1126_,
		_w2746_,
		_w2747_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2490 (
		_w806_,
		_w807_,
		_w809_,
		_w2747_,
		_w2748_
	);
	LUT4 #(
		.INIT('h0c8c)
	) name2491 (
		_w810_,
		_w813_,
		_w811_,
		_w2748_,
		_w2749_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2492 (
		_w814_,
		_w815_,
		_w817_,
		_w2749_,
		_w2750_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2493 (
		_w818_,
		_w819_,
		_w821_,
		_w2750_,
		_w2751_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2494 (
		_w822_,
		_w823_,
		_w825_,
		_w2751_,
		_w2752_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2495 (
		_w826_,
		_w827_,
		_w829_,
		_w2752_,
		_w2753_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2496 (
		_w830_,
		_w831_,
		_w833_,
		_w2753_,
		_w2754_
	);
	LUT4 #(
		.INIT('h8a00)
	) name2497 (
		_w575_,
		_w577_,
		_w579_,
		_w2743_,
		_w2755_
	);
	LUT4 #(
		.INIT('h5d00)
	) name2498 (
		_w835_,
		_w834_,
		_w2754_,
		_w2755_,
		_w2756_
	);
	LUT2 #(
		.INIT('he)
	) name2499 (
		_w2744_,
		_w2756_,
		_w2757_
	);
	LUT3 #(
		.INIT('hb0)
	) name2500 (
		\priority[124] ,
		\req[123] ,
		\req[124] ,
		_w2758_
	);
	LUT2 #(
		.INIT('h4)
	) name2501 (
		_w747_,
		_w2758_,
		_w2759_
	);
	LUT3 #(
		.INIT('h31)
	) name2502 (
		\priority[125] ,
		\priority[126] ,
		\req[125] ,
		_w2760_
	);
	LUT4 #(
		.INIT('ha020)
	) name2503 (
		_w424_,
		_w585_,
		_w800_,
		_w2760_,
		_w2761_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name2504 (
		_w848_,
		_w1142_,
		_w1143_,
		_w2761_,
		_w2762_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2505 (
		_w849_,
		_w850_,
		_w852_,
		_w2762_,
		_w2763_
	);
	LUT4 #(
		.INIT('h4c44)
	) name2506 (
		_w854_,
		_w856_,
		_w2763_,
		_w853_,
		_w2764_
	);
	LUT4 #(
		.INIT('h0c8c)
	) name2507 (
		_w857_,
		_w860_,
		_w858_,
		_w2764_,
		_w2765_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2508 (
		_w861_,
		_w862_,
		_w864_,
		_w2765_,
		_w2766_
	);
	LUT4 #(
		.INIT('h0c8c)
	) name2509 (
		_w865_,
		_w868_,
		_w866_,
		_w2766_,
		_w2767_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2510 (
		_w869_,
		_w870_,
		_w872_,
		_w2767_,
		_w2768_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2511 (
		_w873_,
		_w874_,
		_w876_,
		_w2768_,
		_w2769_
	);
	LUT4 #(
		.INIT('h8a00)
	) name2512 (
		_w741_,
		_w743_,
		_w745_,
		_w2758_,
		_w2770_
	);
	LUT4 #(
		.INIT('h3b00)
	) name2513 (
		_w877_,
		_w878_,
		_w2769_,
		_w2770_,
		_w2771_
	);
	LUT2 #(
		.INIT('he)
	) name2514 (
		_w2759_,
		_w2771_,
		_w2772_
	);
	LUT3 #(
		.INIT('hb0)
	) name2515 (
		\priority[125] ,
		\req[124] ,
		\req[125] ,
		_w2773_
	);
	LUT2 #(
		.INIT('h4)
	) name2516 (
		_w414_,
		_w2773_,
		_w2774_
	);
	LUT3 #(
		.INIT('h31)
	) name2517 (
		\priority[126] ,
		\priority[127] ,
		\req[126] ,
		_w2775_
	);
	LUT4 #(
		.INIT('h8808)
	) name2518 (
		_w264_,
		_w590_,
		_w751_,
		_w2775_,
		_w2776_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name2519 (
		_w890_,
		_w1159_,
		_w1160_,
		_w2776_,
		_w2777_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2520 (
		_w891_,
		_w892_,
		_w894_,
		_w2777_,
		_w2778_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2521 (
		_w895_,
		_w896_,
		_w898_,
		_w2778_,
		_w2779_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2522 (
		_w899_,
		_w900_,
		_w902_,
		_w2779_,
		_w2780_
	);
	LUT4 #(
		.INIT('h44c4)
	) name2523 (
		_w904_,
		_w906_,
		_w903_,
		_w2780_,
		_w2781_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2524 (
		_w907_,
		_w908_,
		_w910_,
		_w2781_,
		_w2782_
	);
	LUT4 #(
		.INIT('h0c8c)
	) name2525 (
		_w911_,
		_w914_,
		_w912_,
		_w2782_,
		_w2783_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2526 (
		_w915_,
		_w916_,
		_w918_,
		_w2783_,
		_w2784_
	);
	LUT4 #(
		.INIT('hb000)
	) name2527 (
		_w409_,
		_w415_,
		_w418_,
		_w2773_,
		_w2785_
	);
	LUT4 #(
		.INIT('h5d00)
	) name2528 (
		_w920_,
		_w919_,
		_w2784_,
		_w2785_,
		_w2786_
	);
	LUT2 #(
		.INIT('he)
	) name2529 (
		_w2774_,
		_w2786_,
		_w2787_
	);
	LUT3 #(
		.INIT('hb0)
	) name2530 (
		\priority[126] ,
		\req[125] ,
		\req[126] ,
		_w2788_
	);
	LUT2 #(
		.INIT('h4)
	) name2531 (
		_w580_,
		_w2788_,
		_w2789_
	);
	LUT3 #(
		.INIT('h51)
	) name2532 (
		\priority[0] ,
		\priority[127] ,
		\req[127] ,
		_w2790_
	);
	LUT4 #(
		.INIT('h8808)
	) name2533 (
		_w430_,
		_w756_,
		_w795_,
		_w2790_,
		_w2791_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name2534 (
		_w932_,
		_w1176_,
		_w1177_,
		_w2791_,
		_w2792_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2535 (
		_w933_,
		_w934_,
		_w936_,
		_w2792_,
		_w2793_
	);
	LUT4 #(
		.INIT('h44c4)
	) name2536 (
		_w938_,
		_w940_,
		_w937_,
		_w2793_,
		_w2794_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2537 (
		_w941_,
		_w942_,
		_w944_,
		_w2794_,
		_w2795_
	);
	LUT4 #(
		.INIT('h0c8c)
	) name2538 (
		_w945_,
		_w948_,
		_w946_,
		_w2795_,
		_w2796_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2539 (
		_w949_,
		_w950_,
		_w952_,
		_w2796_,
		_w2797_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2540 (
		_w953_,
		_w954_,
		_w956_,
		_w2797_,
		_w2798_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name2541 (
		_w960_,
		_w957_,
		_w958_,
		_w2798_,
		_w2799_
	);
	LUT4 #(
		.INIT('hb000)
	) name2542 (
		_w575_,
		_w581_,
		_w584_,
		_w2788_,
		_w2800_
	);
	LUT4 #(
		.INIT('h3b00)
	) name2543 (
		_w961_,
		_w962_,
		_w2799_,
		_w2800_,
		_w2801_
	);
	LUT2 #(
		.INIT('he)
	) name2544 (
		_w2789_,
		_w2801_,
		_w2802_
	);
	LUT3 #(
		.INIT('hb0)
	) name2545 (
		\priority[127] ,
		\req[126] ,
		\req[127] ,
		_w2803_
	);
	LUT2 #(
		.INIT('h4)
	) name2546 (
		_w746_,
		_w2803_,
		_w2804_
	);
	LUT3 #(
		.INIT('h31)
	) name2547 (
		\priority[0] ,
		\priority[1] ,
		\req[0] ,
		_w2805_
	);
	LUT4 #(
		.INIT('h8808)
	) name2548 (
		_w596_,
		_w800_,
		_w839_,
		_w2805_,
		_w2806_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name2549 (
		_w974_,
		_w1193_,
		_w1194_,
		_w2806_,
		_w2807_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2550 (
		_w975_,
		_w976_,
		_w978_,
		_w2807_,
		_w2808_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2551 (
		_w979_,
		_w980_,
		_w982_,
		_w2808_,
		_w2809_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2552 (
		_w983_,
		_w984_,
		_w986_,
		_w2809_,
		_w2810_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2553 (
		_w987_,
		_w988_,
		_w990_,
		_w2810_,
		_w2811_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2554 (
		_w991_,
		_w992_,
		_w994_,
		_w2811_,
		_w2812_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2555 (
		_w995_,
		_w996_,
		_w998_,
		_w2812_,
		_w2813_
	);
	LUT4 #(
		.INIT('h44c4)
	) name2556 (
		_w1000_,
		_w1002_,
		_w999_,
		_w2813_,
		_w2814_
	);
	LUT4 #(
		.INIT('hb000)
	) name2557 (
		_w741_,
		_w747_,
		_w750_,
		_w2803_,
		_w2815_
	);
	LUT4 #(
		.INIT('h3b00)
	) name2558 (
		_w1003_,
		_w1004_,
		_w2814_,
		_w2815_,
		_w2816_
	);
	LUT2 #(
		.INIT('he)
	) name2559 (
		_w2804_,
		_w2816_,
		_w2817_
	);
	LUT4 #(
		.INIT('h0001)
	) name2560 (
		\req[6] ,
		\req[7] ,
		\req[122] ,
		\req[123] ,
		_w2818_
	);
	LUT4 #(
		.INIT('h0001)
	) name2561 (
		\req[12] ,
		\req[13] ,
		\req[18] ,
		\req[19] ,
		_w2819_
	);
	LUT4 #(
		.INIT('h0001)
	) name2562 (
		\req[98] ,
		\req[99] ,
		\req[104] ,
		\req[105] ,
		_w2820_
	);
	LUT4 #(
		.INIT('h0001)
	) name2563 (
		\req[110] ,
		\req[111] ,
		\req[116] ,
		\req[117] ,
		_w2821_
	);
	LUT4 #(
		.INIT('h8000)
	) name2564 (
		_w2818_,
		_w2819_,
		_w2820_,
		_w2821_,
		_w2822_
	);
	LUT4 #(
		.INIT('h0001)
	) name2565 (
		\req[48] ,
		\req[49] ,
		\req[54] ,
		\req[55] ,
		_w2823_
	);
	LUT4 #(
		.INIT('h0001)
	) name2566 (
		\req[60] ,
		\req[61] ,
		\req[66] ,
		\req[67] ,
		_w2824_
	);
	LUT4 #(
		.INIT('h0001)
	) name2567 (
		\req[24] ,
		\req[25] ,
		\req[30] ,
		\req[31] ,
		_w2825_
	);
	LUT4 #(
		.INIT('h0001)
	) name2568 (
		\req[36] ,
		\req[37] ,
		\req[42] ,
		\req[43] ,
		_w2826_
	);
	LUT4 #(
		.INIT('h8000)
	) name2569 (
		_w2823_,
		_w2824_,
		_w2825_,
		_w2826_,
		_w2827_
	);
	LUT4 #(
		.INIT('h0001)
	) name2570 (
		\req[26] ,
		\req[27] ,
		\req[32] ,
		\req[33] ,
		_w2828_
	);
	LUT4 #(
		.INIT('h0001)
	) name2571 (
		\req[38] ,
		\req[39] ,
		\req[44] ,
		\req[45] ,
		_w2829_
	);
	LUT4 #(
		.INIT('h0001)
	) name2572 (
		\req[2] ,
		\req[3] ,
		\req[8] ,
		\req[9] ,
		_w2830_
	);
	LUT4 #(
		.INIT('h0001)
	) name2573 (
		\req[14] ,
		\req[15] ,
		\req[20] ,
		\req[21] ,
		_w2831_
	);
	LUT4 #(
		.INIT('h8000)
	) name2574 (
		_w2828_,
		_w2829_,
		_w2830_,
		_w2831_,
		_w2832_
	);
	LUT4 #(
		.INIT('h0001)
	) name2575 (
		\req[74] ,
		\req[75] ,
		\req[80] ,
		\req[81] ,
		_w2833_
	);
	LUT4 #(
		.INIT('h0001)
	) name2576 (
		\req[86] ,
		\req[87] ,
		\req[92] ,
		\req[93] ,
		_w2834_
	);
	LUT4 #(
		.INIT('h0001)
	) name2577 (
		\req[50] ,
		\req[51] ,
		\req[56] ,
		\req[57] ,
		_w2835_
	);
	LUT4 #(
		.INIT('h0001)
	) name2578 (
		\req[62] ,
		\req[63] ,
		\req[68] ,
		\req[69] ,
		_w2836_
	);
	LUT4 #(
		.INIT('h8000)
	) name2579 (
		_w2833_,
		_w2834_,
		_w2835_,
		_w2836_,
		_w2837_
	);
	LUT4 #(
		.INIT('h8000)
	) name2580 (
		_w2822_,
		_w2827_,
		_w2832_,
		_w2837_,
		_w2838_
	);
	LUT4 #(
		.INIT('h0001)
	) name2581 (
		\req[64] ,
		\req[65] ,
		\req[70] ,
		\req[71] ,
		_w2839_
	);
	LUT4 #(
		.INIT('h0001)
	) name2582 (
		\req[76] ,
		\req[77] ,
		\req[82] ,
		\req[83] ,
		_w2840_
	);
	LUT4 #(
		.INIT('h0001)
	) name2583 (
		\req[40] ,
		\req[41] ,
		\req[46] ,
		\req[47] ,
		_w2841_
	);
	LUT4 #(
		.INIT('h0001)
	) name2584 (
		\req[52] ,
		\req[53] ,
		\req[58] ,
		\req[59] ,
		_w2842_
	);
	LUT4 #(
		.INIT('h8000)
	) name2585 (
		_w2839_,
		_w2840_,
		_w2841_,
		_w2842_,
		_w2843_
	);
	LUT4 #(
		.INIT('h0001)
	) name2586 (
		\req[112] ,
		\req[113] ,
		\req[118] ,
		\req[119] ,
		_w2844_
	);
	LUT4 #(
		.INIT('h0001)
	) name2587 (
		\req[0] ,
		\req[1] ,
		\req[124] ,
		\req[125] ,
		_w2845_
	);
	LUT4 #(
		.INIT('h0001)
	) name2588 (
		\req[88] ,
		\req[89] ,
		\req[94] ,
		\req[95] ,
		_w2846_
	);
	LUT4 #(
		.INIT('h0001)
	) name2589 (
		\req[100] ,
		\req[101] ,
		\req[106] ,
		\req[107] ,
		_w2847_
	);
	LUT4 #(
		.INIT('h8000)
	) name2590 (
		_w2844_,
		_w2845_,
		_w2846_,
		_w2847_,
		_w2848_
	);
	LUT4 #(
		.INIT('h0001)
	) name2591 (
		\req[96] ,
		\req[97] ,
		\req[102] ,
		\req[103] ,
		_w2849_
	);
	LUT4 #(
		.INIT('h0001)
	) name2592 (
		\req[108] ,
		\req[109] ,
		\req[114] ,
		\req[115] ,
		_w2850_
	);
	LUT4 #(
		.INIT('h0001)
	) name2593 (
		\req[72] ,
		\req[73] ,
		\req[78] ,
		\req[79] ,
		_w2851_
	);
	LUT4 #(
		.INIT('h0001)
	) name2594 (
		\req[84] ,
		\req[85] ,
		\req[90] ,
		\req[91] ,
		_w2852_
	);
	LUT4 #(
		.INIT('h8000)
	) name2595 (
		_w2849_,
		_w2850_,
		_w2851_,
		_w2852_,
		_w2853_
	);
	LUT4 #(
		.INIT('h0001)
	) name2596 (
		\req[16] ,
		\req[17] ,
		\req[22] ,
		\req[23] ,
		_w2854_
	);
	LUT4 #(
		.INIT('h0001)
	) name2597 (
		\req[28] ,
		\req[29] ,
		\req[34] ,
		\req[35] ,
		_w2855_
	);
	LUT4 #(
		.INIT('h0001)
	) name2598 (
		\req[120] ,
		\req[121] ,
		\req[126] ,
		\req[127] ,
		_w2856_
	);
	LUT4 #(
		.INIT('h0001)
	) name2599 (
		\req[4] ,
		\req[5] ,
		\req[10] ,
		\req[11] ,
		_w2857_
	);
	LUT4 #(
		.INIT('h8000)
	) name2600 (
		_w2854_,
		_w2855_,
		_w2856_,
		_w2857_,
		_w2858_
	);
	LUT4 #(
		.INIT('h8000)
	) name2601 (
		_w2843_,
		_w2848_,
		_w2853_,
		_w2858_,
		_w2859_
	);
	LUT2 #(
		.INIT('h7)
	) name2602 (
		_w2838_,
		_w2859_,
		_w2860_
	);
	assign \grant[0]  = _w423_ ;
	assign \grant[1]  = _w589_ ;
	assign \grant[2]  = _w755_ ;
	assign \grant[3]  = _w799_ ;
	assign \grant[4]  = _w843_ ;
	assign \grant[5]  = _w885_ ;
	assign \grant[6]  = _w927_ ;
	assign \grant[7]  = _w969_ ;
	assign \grant[8]  = _w1010_ ;
	assign \grant[9]  = _w1027_ ;
	assign \grant[10]  = _w1044_ ;
	assign \grant[11]  = _w1061_ ;
	assign \grant[12]  = _w1078_ ;
	assign \grant[13]  = _w1095_ ;
	assign \grant[14]  = _w1112_ ;
	assign \grant[15]  = _w1129_ ;
	assign \grant[16]  = _w1146_ ;
	assign \grant[17]  = _w1163_ ;
	assign \grant[18]  = _w1180_ ;
	assign \grant[19]  = _w1197_ ;
	assign \grant[20]  = _w1212_ ;
	assign \grant[21]  = _w1227_ ;
	assign \grant[22]  = _w1242_ ;
	assign \grant[23]  = _w1257_ ;
	assign \grant[24]  = _w1272_ ;
	assign \grant[25]  = _w1287_ ;
	assign \grant[26]  = _w1302_ ;
	assign \grant[27]  = _w1317_ ;
	assign \grant[28]  = _w1332_ ;
	assign \grant[29]  = _w1347_ ;
	assign \grant[30]  = _w1362_ ;
	assign \grant[31]  = _w1377_ ;
	assign \grant[32]  = _w1392_ ;
	assign \grant[33]  = _w1407_ ;
	assign \grant[34]  = _w1422_ ;
	assign \grant[35]  = _w1437_ ;
	assign \grant[36]  = _w1452_ ;
	assign \grant[37]  = _w1467_ ;
	assign \grant[38]  = _w1482_ ;
	assign \grant[39]  = _w1497_ ;
	assign \grant[40]  = _w1512_ ;
	assign \grant[41]  = _w1527_ ;
	assign \grant[42]  = _w1542_ ;
	assign \grant[43]  = _w1557_ ;
	assign \grant[44]  = _w1572_ ;
	assign \grant[45]  = _w1587_ ;
	assign \grant[46]  = _w1602_ ;
	assign \grant[47]  = _w1617_ ;
	assign \grant[48]  = _w1632_ ;
	assign \grant[49]  = _w1647_ ;
	assign \grant[50]  = _w1662_ ;
	assign \grant[51]  = _w1677_ ;
	assign \grant[52]  = _w1692_ ;
	assign \grant[53]  = _w1707_ ;
	assign \grant[54]  = _w1722_ ;
	assign \grant[55]  = _w1737_ ;
	assign \grant[56]  = _w1752_ ;
	assign \grant[57]  = _w1767_ ;
	assign \grant[58]  = _w1782_ ;
	assign \grant[59]  = _w1797_ ;
	assign \grant[60]  = _w1812_ ;
	assign \grant[61]  = _w1827_ ;
	assign \grant[62]  = _w1842_ ;
	assign \grant[63]  = _w1857_ ;
	assign \grant[64]  = _w1872_ ;
	assign \grant[65]  = _w1887_ ;
	assign \grant[66]  = _w1902_ ;
	assign \grant[67]  = _w1917_ ;
	assign \grant[68]  = _w1932_ ;
	assign \grant[69]  = _w1947_ ;
	assign \grant[70]  = _w1962_ ;
	assign \grant[71]  = _w1977_ ;
	assign \grant[72]  = _w1992_ ;
	assign \grant[73]  = _w2007_ ;
	assign \grant[74]  = _w2022_ ;
	assign \grant[75]  = _w2037_ ;
	assign \grant[76]  = _w2052_ ;
	assign \grant[77]  = _w2067_ ;
	assign \grant[78]  = _w2082_ ;
	assign \grant[79]  = _w2097_ ;
	assign \grant[80]  = _w2112_ ;
	assign \grant[81]  = _w2127_ ;
	assign \grant[82]  = _w2142_ ;
	assign \grant[83]  = _w2157_ ;
	assign \grant[84]  = _w2172_ ;
	assign \grant[85]  = _w2187_ ;
	assign \grant[86]  = _w2202_ ;
	assign \grant[87]  = _w2217_ ;
	assign \grant[88]  = _w2232_ ;
	assign \grant[89]  = _w2247_ ;
	assign \grant[90]  = _w2262_ ;
	assign \grant[91]  = _w2277_ ;
	assign \grant[92]  = _w2292_ ;
	assign \grant[93]  = _w2307_ ;
	assign \grant[94]  = _w2322_ ;
	assign \grant[95]  = _w2337_ ;
	assign \grant[96]  = _w2352_ ;
	assign \grant[97]  = _w2367_ ;
	assign \grant[98]  = _w2382_ ;
	assign \grant[99]  = _w2397_ ;
	assign \grant[100]  = _w2412_ ;
	assign \grant[101]  = _w2427_ ;
	assign \grant[102]  = _w2442_ ;
	assign \grant[103]  = _w2457_ ;
	assign \grant[104]  = _w2472_ ;
	assign \grant[105]  = _w2487_ ;
	assign \grant[106]  = _w2502_ ;
	assign \grant[107]  = _w2517_ ;
	assign \grant[108]  = _w2532_ ;
	assign \grant[109]  = _w2547_ ;
	assign \grant[110]  = _w2562_ ;
	assign \grant[111]  = _w2577_ ;
	assign \grant[112]  = _w2592_ ;
	assign \grant[113]  = _w2607_ ;
	assign \grant[114]  = _w2622_ ;
	assign \grant[115]  = _w2637_ ;
	assign \grant[116]  = _w2652_ ;
	assign \grant[117]  = _w2667_ ;
	assign \grant[118]  = _w2682_ ;
	assign \grant[119]  = _w2697_ ;
	assign \grant[120]  = _w2712_ ;
	assign \grant[121]  = _w2727_ ;
	assign \grant[122]  = _w2742_ ;
	assign \grant[123]  = _w2757_ ;
	assign \grant[124]  = _w2772_ ;
	assign \grant[125]  = _w2787_ ;
	assign \grant[126]  = _w2802_ ;
	assign \grant[127]  = _w2817_ ;
	assign anyGrant = _w2860_ ;
endmodule;