module top (a_pad, b_pad, c_pad, d_pad, e_pad, f_pad, g_pad, h_pad, i_pad, j_pad, k_pad, l_pad);
	input a_pad ;
	input b_pad ;
	input c_pad ;
	input d_pad ;
	input e_pad ;
	input f_pad ;
	input g_pad ;
	input h_pad ;
	input i_pad ;
	input j_pad ;
	input k_pad ;
	output l_pad ;
	wire _w32_ ;
	wire _w31_ ;
	wire _w30_ ;
	wire _w29_ ;
	wire _w28_ ;
	wire _w27_ ;
	wire _w26_ ;
	wire _w25_ ;
	wire _w12_ ;
	wire _w13_ ;
	wire _w14_ ;
	wire _w15_ ;
	wire _w16_ ;
	wire _w17_ ;
	wire _w18_ ;
	wire _w19_ ;
	wire _w20_ ;
	wire _w21_ ;
	wire _w22_ ;
	wire _w23_ ;
	wire _w24_ ;
	LUT2 #(
		.INIT('h1)
	) name0 (
		e_pad,
		j_pad,
		_w12_
	);
	LUT2 #(
		.INIT('h4)
	) name1 (
		g_pad,
		j_pad,
		_w13_
	);
	LUT2 #(
		.INIT('h1)
	) name2 (
		i_pad,
		_w12_,
		_w14_
	);
	LUT2 #(
		.INIT('h4)
	) name3 (
		_w13_,
		_w14_,
		_w15_
	);
	LUT2 #(
		.INIT('h1)
	) name4 (
		f_pad,
		j_pad,
		_w16_
	);
	LUT2 #(
		.INIT('h4)
	) name5 (
		h_pad,
		j_pad,
		_w17_
	);
	LUT2 #(
		.INIT('h2)
	) name6 (
		i_pad,
		_w16_,
		_w18_
	);
	LUT2 #(
		.INIT('h4)
	) name7 (
		_w17_,
		_w18_,
		_w19_
	);
	LUT2 #(
		.INIT('h1)
	) name8 (
		_w15_,
		_w19_,
		_w20_
	);
	LUT2 #(
		.INIT('h2)
	) name9 (
		k_pad,
		_w20_,
		_w21_
	);
	LUT2 #(
		.INIT('h1)
	) name10 (
		a_pad,
		j_pad,
		_w22_
	);
	LUT2 #(
		.INIT('h4)
	) name11 (
		c_pad,
		j_pad,
		_w23_
	);
	LUT2 #(
		.INIT('h1)
	) name12 (
		i_pad,
		_w22_,
		_w24_
	);
	LUT2 #(
		.INIT('h4)
	) name13 (
		_w23_,
		_w24_,
		_w25_
	);
	LUT2 #(
		.INIT('h4)
	) name14 (
		d_pad,
		j_pad,
		_w26_
	);
	LUT2 #(
		.INIT('h1)
	) name15 (
		b_pad,
		j_pad,
		_w27_
	);
	LUT2 #(
		.INIT('h2)
	) name16 (
		i_pad,
		_w26_,
		_w28_
	);
	LUT2 #(
		.INIT('h4)
	) name17 (
		_w27_,
		_w28_,
		_w29_
	);
	LUT2 #(
		.INIT('h1)
	) name18 (
		_w25_,
		_w29_,
		_w30_
	);
	LUT2 #(
		.INIT('h1)
	) name19 (
		k_pad,
		_w30_,
		_w31_
	);
	LUT2 #(
		.INIT('h1)
	) name20 (
		_w21_,
		_w31_,
		_w32_
	);
	assign l_pad = _w32_ ;
endmodule;