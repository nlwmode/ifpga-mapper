module top (a_pad, \b0_pad , b_pad, \c0_pad , c_pad, \d0_pad , d_pad, \e0_pad , e_pad, f_pad, g_pad, \h0_pad , h_pad, i_pad, j_pad, k_pad, l_pad, m_pad, o_pad, t_pad, v_pad, \a0_pad , \f0_pad , \g0_pad , \i0_pad , \j0_pad , \k0_pad , \l0_pad , \m0_pad , \n0_pad , \o0_pad , \p0_pad , w_pad, x_pad, y_pad, z_pad);
	input a_pad ;
	input \b0_pad  ;
	input b_pad ;
	input \c0_pad  ;
	input c_pad ;
	input \d0_pad  ;
	input d_pad ;
	input \e0_pad  ;
	input e_pad ;
	input f_pad ;
	input g_pad ;
	input \h0_pad  ;
	input h_pad ;
	input i_pad ;
	input j_pad ;
	input k_pad ;
	input l_pad ;
	input m_pad ;
	input o_pad ;
	input t_pad ;
	input v_pad ;
	output \a0_pad  ;
	output \f0_pad  ;
	output \g0_pad  ;
	output \i0_pad  ;
	output \j0_pad  ;
	output \k0_pad  ;
	output \l0_pad  ;
	output \m0_pad  ;
	output \n0_pad  ;
	output \o0_pad  ;
	output \p0_pad  ;
	output w_pad ;
	output x_pad ;
	output y_pad ;
	output z_pad ;
	wire _w64_ ;
	wire _w63_ ;
	wire _w62_ ;
	wire _w61_ ;
	wire _w60_ ;
	wire _w59_ ;
	wire _w58_ ;
	wire _w57_ ;
	wire _w56_ ;
	wire _w55_ ;
	wire _w54_ ;
	wire _w53_ ;
	wire _w52_ ;
	wire _w51_ ;
	wire _w34_ ;
	wire _w33_ ;
	wire _w32_ ;
	wire _w31_ ;
	wire _w30_ ;
	wire _w29_ ;
	wire _w28_ ;
	wire _w27_ ;
	wire _w26_ ;
	wire _w25_ ;
	wire _w24_ ;
	wire _w23_ ;
	wire _w22_ ;
	wire _w35_ ;
	wire _w36_ ;
	wire _w37_ ;
	wire _w38_ ;
	wire _w39_ ;
	wire _w40_ ;
	wire _w41_ ;
	wire _w42_ ;
	wire _w43_ ;
	wire _w44_ ;
	wire _w45_ ;
	wire _w46_ ;
	wire _w47_ ;
	wire _w48_ ;
	wire _w49_ ;
	wire _w50_ ;
	LUT2 #(
		.INIT('h8)
	) name0 (
		i_pad,
		j_pad,
		_w22_
	);
	LUT2 #(
		.INIT('h8)
	) name1 (
		i_pad,
		k_pad,
		_w23_
	);
	LUT2 #(
		.INIT('h4)
	) name2 (
		\c0_pad ,
		_w23_,
		_w24_
	);
	LUT2 #(
		.INIT('h1)
	) name3 (
		o_pad,
		_w24_,
		_w25_
	);
	LUT2 #(
		.INIT('h4)
	) name4 (
		a_pad,
		_w24_,
		_w26_
	);
	LUT2 #(
		.INIT('h2)
	) name5 (
		m_pad,
		_w25_,
		_w27_
	);
	LUT2 #(
		.INIT('h4)
	) name6 (
		_w26_,
		_w27_,
		_w28_
	);
	LUT2 #(
		.INIT('h8)
	) name7 (
		\c0_pad ,
		_w23_,
		_w29_
	);
	LUT2 #(
		.INIT('h1)
	) name8 (
		\h0_pad ,
		_w29_,
		_w30_
	);
	LUT2 #(
		.INIT('h8)
	) name9 (
		b_pad,
		_w24_,
		_w31_
	);
	LUT2 #(
		.INIT('h2)
	) name10 (
		m_pad,
		_w30_,
		_w32_
	);
	LUT2 #(
		.INIT('h4)
	) name11 (
		_w31_,
		_w32_,
		_w33_
	);
	LUT2 #(
		.INIT('h8)
	) name12 (
		c_pad,
		_w23_,
		_w34_
	);
	LUT2 #(
		.INIT('h1)
	) name13 (
		\c0_pad ,
		_w34_,
		_w35_
	);
	LUT2 #(
		.INIT('h2)
	) name14 (
		m_pad,
		_w29_,
		_w36_
	);
	LUT2 #(
		.INIT('h4)
	) name15 (
		_w35_,
		_w36_,
		_w37_
	);
	LUT2 #(
		.INIT('h4)
	) name16 (
		d_pad,
		_w24_,
		_w38_
	);
	LUT2 #(
		.INIT('h2)
	) name17 (
		\e0_pad ,
		\h0_pad ,
		_w39_
	);
	LUT2 #(
		.INIT('h1)
	) name18 (
		_w24_,
		_w39_,
		_w40_
	);
	LUT2 #(
		.INIT('h2)
	) name19 (
		m_pad,
		_w38_,
		_w41_
	);
	LUT2 #(
		.INIT('h4)
	) name20 (
		_w40_,
		_w41_,
		_w42_
	);
	LUT2 #(
		.INIT('h1)
	) name21 (
		\d0_pad ,
		_w24_,
		_w43_
	);
	LUT2 #(
		.INIT('h4)
	) name22 (
		e_pad,
		_w24_,
		_w44_
	);
	LUT2 #(
		.INIT('h2)
	) name23 (
		m_pad,
		_w43_,
		_w45_
	);
	LUT2 #(
		.INIT('h4)
	) name24 (
		_w44_,
		_w45_,
		_w46_
	);
	LUT2 #(
		.INIT('h1)
	) name25 (
		t_pad,
		_w24_,
		_w47_
	);
	LUT2 #(
		.INIT('h4)
	) name26 (
		f_pad,
		_w24_,
		_w48_
	);
	LUT2 #(
		.INIT('h2)
	) name27 (
		m_pad,
		_w47_,
		_w49_
	);
	LUT2 #(
		.INIT('h4)
	) name28 (
		_w48_,
		_w49_,
		_w50_
	);
	LUT2 #(
		.INIT('h1)
	) name29 (
		\b0_pad ,
		_w24_,
		_w51_
	);
	LUT2 #(
		.INIT('h4)
	) name30 (
		g_pad,
		_w24_,
		_w52_
	);
	LUT2 #(
		.INIT('h2)
	) name31 (
		m_pad,
		_w51_,
		_w53_
	);
	LUT2 #(
		.INIT('h4)
	) name32 (
		_w52_,
		_w53_,
		_w54_
	);
	LUT2 #(
		.INIT('h1)
	) name33 (
		v_pad,
		_w24_,
		_w55_
	);
	LUT2 #(
		.INIT('h4)
	) name34 (
		h_pad,
		_w24_,
		_w56_
	);
	LUT2 #(
		.INIT('h2)
	) name35 (
		m_pad,
		_w55_,
		_w57_
	);
	LUT2 #(
		.INIT('h4)
	) name36 (
		_w56_,
		_w57_,
		_w58_
	);
	LUT2 #(
		.INIT('h8)
	) name37 (
		l_pad,
		v_pad,
		_w59_
	);
	LUT2 #(
		.INIT('h4)
	) name38 (
		\h0_pad ,
		_w29_,
		_w60_
	);
	LUT2 #(
		.INIT('h1)
	) name39 (
		\h0_pad ,
		_w24_,
		_w61_
	);
	LUT2 #(
		.INIT('h4)
	) name40 (
		l_pad,
		m_pad,
		_w62_
	);
	LUT2 #(
		.INIT('h4)
	) name41 (
		_w61_,
		_w62_,
		_w63_
	);
	LUT2 #(
		.INIT('h8)
	) name42 (
		m_pad,
		_w60_,
		_w64_
	);
	assign \a0_pad  = t_pad;
	assign \f0_pad  = _w22_ ;
	assign \g0_pad  = _w22_ ;
	assign \i0_pad  = _w28_ ;
	assign \j0_pad  = _w33_ ;
	assign \k0_pad  = _w37_ ;
	assign \l0_pad  = _w42_ ;
	assign \m0_pad  = _w46_ ;
	assign \n0_pad  = _w50_ ;
	assign \o0_pad  = _w54_ ;
	assign \p0_pad  = _w58_ ;
	assign w_pad = _w59_ ;
	assign x_pad = _w60_ ;
	assign y_pad = _w63_ ;
	assign z_pad = _w64_ ;
endmodule;