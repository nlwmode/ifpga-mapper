module top (\inA0_pad , \inA10_pad , \inA11_pad , \inA12_pad , \inA13_pad , \inA14_pad , \inA15_pad , \inA1_pad , \inA2_pad , \inA3_pad , \inA4_pad , \inA5_pad , \inA6_pad , \inA7_pad , \inA8_pad , \inA9_pad , \inB0_pad , \inB10_pad , \inB11_pad , \inB12_pad , \inB13_pad , \inB14_pad , \inB15_pad , \inB1_pad , \inB2_pad , \inB3_pad , \inB4_pad , \inB5_pad , \inB6_pad , \inB7_pad , \inB8_pad , \inB9_pad , \inC0_pad , \inC10_pad , \inC11_pad , \inC12_pad , \inC13_pad , \inC14_pad , \inC15_pad , \inC1_pad , \inC2_pad , \inC3_pad , \inC4_pad , \inC5_pad , \inC6_pad , \inC7_pad , \inC8_pad , \inC9_pad , \inD0_pad , \inD10_pad , \inD11_pad , \inD12_pad , \inD13_pad , \inD14_pad , \inD15_pad , \inD1_pad , \inD2_pad , \inD3_pad , \inD4_pad , \inD5_pad , \inD6_pad , \inD7_pad , \inD8_pad , \inD9_pad , \musel1_pad , \musel2_pad , \musel3_pad , \musel4_pad , \opsel0_pad , \opsel1_pad , \opsel2_pad , \opsel3_pad , \sh0_pad , \sh1_pad , \sh2_pad , \O0_pad , \O10_pad , \O11_pad , \O12_pad , \O13_pad , \O14_pad , \O15_pad , \O1_pad , \O2_pad , \O3_pad , \O4_pad , \O5_pad , \O6_pad , \O7_pad , \O8_pad , \O9_pad );
	input \inA0_pad  ;
	input \inA10_pad  ;
	input \inA11_pad  ;
	input \inA12_pad  ;
	input \inA13_pad  ;
	input \inA14_pad  ;
	input \inA15_pad  ;
	input \inA1_pad  ;
	input \inA2_pad  ;
	input \inA3_pad  ;
	input \inA4_pad  ;
	input \inA5_pad  ;
	input \inA6_pad  ;
	input \inA7_pad  ;
	input \inA8_pad  ;
	input \inA9_pad  ;
	input \inB0_pad  ;
	input \inB10_pad  ;
	input \inB11_pad  ;
	input \inB12_pad  ;
	input \inB13_pad  ;
	input \inB14_pad  ;
	input \inB15_pad  ;
	input \inB1_pad  ;
	input \inB2_pad  ;
	input \inB3_pad  ;
	input \inB4_pad  ;
	input \inB5_pad  ;
	input \inB6_pad  ;
	input \inB7_pad  ;
	input \inB8_pad  ;
	input \inB9_pad  ;
	input \inC0_pad  ;
	input \inC10_pad  ;
	input \inC11_pad  ;
	input \inC12_pad  ;
	input \inC13_pad  ;
	input \inC14_pad  ;
	input \inC15_pad  ;
	input \inC1_pad  ;
	input \inC2_pad  ;
	input \inC3_pad  ;
	input \inC4_pad  ;
	input \inC5_pad  ;
	input \inC6_pad  ;
	input \inC7_pad  ;
	input \inC8_pad  ;
	input \inC9_pad  ;
	input \inD0_pad  ;
	input \inD10_pad  ;
	input \inD11_pad  ;
	input \inD12_pad  ;
	input \inD13_pad  ;
	input \inD14_pad  ;
	input \inD15_pad  ;
	input \inD1_pad  ;
	input \inD2_pad  ;
	input \inD3_pad  ;
	input \inD4_pad  ;
	input \inD5_pad  ;
	input \inD6_pad  ;
	input \inD7_pad  ;
	input \inD8_pad  ;
	input \inD9_pad  ;
	input \musel1_pad  ;
	input \musel2_pad  ;
	input \musel3_pad  ;
	input \musel4_pad  ;
	input \opsel0_pad  ;
	input \opsel1_pad  ;
	input \opsel2_pad  ;
	input \opsel3_pad  ;
	input \sh0_pad  ;
	input \sh1_pad  ;
	input \sh2_pad  ;
	output \O0_pad  ;
	output \O10_pad  ;
	output \O11_pad  ;
	output \O12_pad  ;
	output \O13_pad  ;
	output \O14_pad  ;
	output \O15_pad  ;
	output \O1_pad  ;
	output \O2_pad  ;
	output \O3_pad  ;
	output \O4_pad  ;
	output \O5_pad  ;
	output \O6_pad  ;
	output \O7_pad  ;
	output \O8_pad  ;
	output \O9_pad  ;
	wire _w1121_ ;
	wire _w1120_ ;
	wire _w1119_ ;
	wire _w1118_ ;
	wire _w1117_ ;
	wire _w1116_ ;
	wire _w1115_ ;
	wire _w1114_ ;
	wire _w1113_ ;
	wire _w1112_ ;
	wire _w1111_ ;
	wire _w1110_ ;
	wire _w1109_ ;
	wire _w1108_ ;
	wire _w1107_ ;
	wire _w1106_ ;
	wire _w1105_ ;
	wire _w1104_ ;
	wire _w1103_ ;
	wire _w1102_ ;
	wire _w1101_ ;
	wire _w1100_ ;
	wire _w1099_ ;
	wire _w1098_ ;
	wire _w1097_ ;
	wire _w1096_ ;
	wire _w1095_ ;
	wire _w1094_ ;
	wire _w1093_ ;
	wire _w1092_ ;
	wire _w1091_ ;
	wire _w1090_ ;
	wire _w1089_ ;
	wire _w1088_ ;
	wire _w1087_ ;
	wire _w1086_ ;
	wire _w1085_ ;
	wire _w1084_ ;
	wire _w1083_ ;
	wire _w1082_ ;
	wire _w1081_ ;
	wire _w1080_ ;
	wire _w1079_ ;
	wire _w1078_ ;
	wire _w1077_ ;
	wire _w1076_ ;
	wire _w1075_ ;
	wire _w1074_ ;
	wire _w1073_ ;
	wire _w1072_ ;
	wire _w1071_ ;
	wire _w1070_ ;
	wire _w1069_ ;
	wire _w1068_ ;
	wire _w1067_ ;
	wire _w1066_ ;
	wire _w1065_ ;
	wire _w1064_ ;
	wire _w1063_ ;
	wire _w1062_ ;
	wire _w1061_ ;
	wire _w1060_ ;
	wire _w1059_ ;
	wire _w1058_ ;
	wire _w1057_ ;
	wire _w1056_ ;
	wire _w1055_ ;
	wire _w1054_ ;
	wire _w1053_ ;
	wire _w1052_ ;
	wire _w1051_ ;
	wire _w1050_ ;
	wire _w1049_ ;
	wire _w1048_ ;
	wire _w1047_ ;
	wire _w1046_ ;
	wire _w1045_ ;
	wire _w1044_ ;
	wire _w1043_ ;
	wire _w1042_ ;
	wire _w1041_ ;
	wire _w1040_ ;
	wire _w1039_ ;
	wire _w1038_ ;
	wire _w1037_ ;
	wire _w1036_ ;
	wire _w1035_ ;
	wire _w1034_ ;
	wire _w1033_ ;
	wire _w1032_ ;
	wire _w1031_ ;
	wire _w1030_ ;
	wire _w1029_ ;
	wire _w1028_ ;
	wire _w1027_ ;
	wire _w1026_ ;
	wire _w1025_ ;
	wire _w1024_ ;
	wire _w1023_ ;
	wire _w1022_ ;
	wire _w1021_ ;
	wire _w1020_ ;
	wire _w1019_ ;
	wire _w1018_ ;
	wire _w1017_ ;
	wire _w1016_ ;
	wire _w1015_ ;
	wire _w1014_ ;
	wire _w1013_ ;
	wire _w1012_ ;
	wire _w1011_ ;
	wire _w1010_ ;
	wire _w1009_ ;
	wire _w1008_ ;
	wire _w1007_ ;
	wire _w1006_ ;
	wire _w1005_ ;
	wire _w1004_ ;
	wire _w1003_ ;
	wire _w1002_ ;
	wire _w1001_ ;
	wire _w1000_ ;
	wire _w999_ ;
	wire _w998_ ;
	wire _w997_ ;
	wire _w996_ ;
	wire _w995_ ;
	wire _w994_ ;
	wire _w993_ ;
	wire _w992_ ;
	wire _w991_ ;
	wire _w990_ ;
	wire _w989_ ;
	wire _w988_ ;
	wire _w987_ ;
	wire _w986_ ;
	wire _w985_ ;
	wire _w984_ ;
	wire _w983_ ;
	wire _w982_ ;
	wire _w981_ ;
	wire _w980_ ;
	wire _w979_ ;
	wire _w978_ ;
	wire _w977_ ;
	wire _w976_ ;
	wire _w975_ ;
	wire _w974_ ;
	wire _w973_ ;
	wire _w972_ ;
	wire _w971_ ;
	wire _w970_ ;
	wire _w969_ ;
	wire _w968_ ;
	wire _w967_ ;
	wire _w966_ ;
	wire _w965_ ;
	wire _w964_ ;
	wire _w963_ ;
	wire _w962_ ;
	wire _w961_ ;
	wire _w960_ ;
	wire _w959_ ;
	wire _w958_ ;
	wire _w957_ ;
	wire _w956_ ;
	wire _w955_ ;
	wire _w954_ ;
	wire _w953_ ;
	wire _w952_ ;
	wire _w951_ ;
	wire _w950_ ;
	wire _w949_ ;
	wire _w948_ ;
	wire _w947_ ;
	wire _w946_ ;
	wire _w945_ ;
	wire _w944_ ;
	wire _w943_ ;
	wire _w942_ ;
	wire _w941_ ;
	wire _w940_ ;
	wire _w939_ ;
	wire _w938_ ;
	wire _w937_ ;
	wire _w936_ ;
	wire _w935_ ;
	wire _w934_ ;
	wire _w933_ ;
	wire _w932_ ;
	wire _w931_ ;
	wire _w930_ ;
	wire _w929_ ;
	wire _w928_ ;
	wire _w927_ ;
	wire _w926_ ;
	wire _w925_ ;
	wire _w924_ ;
	wire _w923_ ;
	wire _w922_ ;
	wire _w921_ ;
	wire _w920_ ;
	wire _w919_ ;
	wire _w918_ ;
	wire _w917_ ;
	wire _w916_ ;
	wire _w915_ ;
	wire _w914_ ;
	wire _w913_ ;
	wire _w912_ ;
	wire _w911_ ;
	wire _w910_ ;
	wire _w909_ ;
	wire _w908_ ;
	wire _w907_ ;
	wire _w906_ ;
	wire _w905_ ;
	wire _w904_ ;
	wire _w903_ ;
	wire _w902_ ;
	wire _w901_ ;
	wire _w900_ ;
	wire _w899_ ;
	wire _w898_ ;
	wire _w897_ ;
	wire _w896_ ;
	wire _w895_ ;
	wire _w894_ ;
	wire _w893_ ;
	wire _w892_ ;
	wire _w891_ ;
	wire _w890_ ;
	wire _w889_ ;
	wire _w888_ ;
	wire _w887_ ;
	wire _w886_ ;
	wire _w885_ ;
	wire _w884_ ;
	wire _w883_ ;
	wire _w882_ ;
	wire _w881_ ;
	wire _w880_ ;
	wire _w879_ ;
	wire _w878_ ;
	wire _w877_ ;
	wire _w876_ ;
	wire _w875_ ;
	wire _w874_ ;
	wire _w873_ ;
	wire _w872_ ;
	wire _w871_ ;
	wire _w870_ ;
	wire _w869_ ;
	wire _w868_ ;
	wire _w867_ ;
	wire _w866_ ;
	wire _w865_ ;
	wire _w864_ ;
	wire _w863_ ;
	wire _w862_ ;
	wire _w861_ ;
	wire _w860_ ;
	wire _w859_ ;
	wire _w858_ ;
	wire _w857_ ;
	wire _w856_ ;
	wire _w855_ ;
	wire _w854_ ;
	wire _w853_ ;
	wire _w852_ ;
	wire _w851_ ;
	wire _w850_ ;
	wire _w849_ ;
	wire _w848_ ;
	wire _w847_ ;
	wire _w846_ ;
	wire _w845_ ;
	wire _w844_ ;
	wire _w843_ ;
	wire _w842_ ;
	wire _w841_ ;
	wire _w840_ ;
	wire _w839_ ;
	wire _w838_ ;
	wire _w837_ ;
	wire _w836_ ;
	wire _w835_ ;
	wire _w834_ ;
	wire _w833_ ;
	wire _w832_ ;
	wire _w831_ ;
	wire _w830_ ;
	wire _w829_ ;
	wire _w828_ ;
	wire _w827_ ;
	wire _w826_ ;
	wire _w825_ ;
	wire _w824_ ;
	wire _w823_ ;
	wire _w822_ ;
	wire _w821_ ;
	wire _w820_ ;
	wire _w819_ ;
	wire _w818_ ;
	wire _w817_ ;
	wire _w816_ ;
	wire _w815_ ;
	wire _w814_ ;
	wire _w813_ ;
	wire _w812_ ;
	wire _w811_ ;
	wire _w810_ ;
	wire _w809_ ;
	wire _w808_ ;
	wire _w807_ ;
	wire _w806_ ;
	wire _w805_ ;
	wire _w804_ ;
	wire _w803_ ;
	wire _w802_ ;
	wire _w801_ ;
	wire _w800_ ;
	wire _w799_ ;
	wire _w798_ ;
	wire _w797_ ;
	wire _w796_ ;
	wire _w795_ ;
	wire _w794_ ;
	wire _w793_ ;
	wire _w792_ ;
	wire _w791_ ;
	wire _w790_ ;
	wire _w789_ ;
	wire _w788_ ;
	wire _w787_ ;
	wire _w786_ ;
	wire _w785_ ;
	wire _w784_ ;
	wire _w783_ ;
	wire _w782_ ;
	wire _w781_ ;
	wire _w780_ ;
	wire _w779_ ;
	wire _w778_ ;
	wire _w777_ ;
	wire _w776_ ;
	wire _w775_ ;
	wire _w774_ ;
	wire _w773_ ;
	wire _w772_ ;
	wire _w771_ ;
	wire _w770_ ;
	wire _w769_ ;
	wire _w768_ ;
	wire _w767_ ;
	wire _w766_ ;
	wire _w765_ ;
	wire _w764_ ;
	wire _w763_ ;
	wire _w762_ ;
	wire _w761_ ;
	wire _w760_ ;
	wire _w759_ ;
	wire _w758_ ;
	wire _w757_ ;
	wire _w756_ ;
	wire _w755_ ;
	wire _w754_ ;
	wire _w753_ ;
	wire _w752_ ;
	wire _w751_ ;
	wire _w750_ ;
	wire _w749_ ;
	wire _w748_ ;
	wire _w747_ ;
	wire _w746_ ;
	wire _w745_ ;
	wire _w744_ ;
	wire _w743_ ;
	wire _w742_ ;
	wire _w741_ ;
	wire _w740_ ;
	wire _w739_ ;
	wire _w738_ ;
	wire _w737_ ;
	wire _w736_ ;
	wire _w735_ ;
	wire _w734_ ;
	wire _w733_ ;
	wire _w732_ ;
	wire _w731_ ;
	wire _w730_ ;
	wire _w729_ ;
	wire _w728_ ;
	wire _w727_ ;
	wire _w726_ ;
	wire _w725_ ;
	wire _w724_ ;
	wire _w723_ ;
	wire _w722_ ;
	wire _w721_ ;
	wire _w720_ ;
	wire _w719_ ;
	wire _w718_ ;
	wire _w717_ ;
	wire _w716_ ;
	wire _w715_ ;
	wire _w714_ ;
	wire _w713_ ;
	wire _w712_ ;
	wire _w711_ ;
	wire _w710_ ;
	wire _w709_ ;
	wire _w708_ ;
	wire _w707_ ;
	wire _w706_ ;
	wire _w705_ ;
	wire _w704_ ;
	wire _w703_ ;
	wire _w702_ ;
	wire _w701_ ;
	wire _w700_ ;
	wire _w699_ ;
	wire _w698_ ;
	wire _w697_ ;
	wire _w696_ ;
	wire _w695_ ;
	wire _w694_ ;
	wire _w693_ ;
	wire _w692_ ;
	wire _w691_ ;
	wire _w690_ ;
	wire _w689_ ;
	wire _w688_ ;
	wire _w687_ ;
	wire _w686_ ;
	wire _w685_ ;
	wire _w684_ ;
	wire _w683_ ;
	wire _w682_ ;
	wire _w681_ ;
	wire _w680_ ;
	wire _w679_ ;
	wire _w678_ ;
	wire _w677_ ;
	wire _w676_ ;
	wire _w675_ ;
	wire _w674_ ;
	wire _w673_ ;
	wire _w672_ ;
	wire _w671_ ;
	wire _w670_ ;
	wire _w669_ ;
	wire _w668_ ;
	wire _w667_ ;
	wire _w666_ ;
	wire _w665_ ;
	wire _w664_ ;
	wire _w663_ ;
	wire _w662_ ;
	wire _w661_ ;
	wire _w660_ ;
	wire _w659_ ;
	wire _w658_ ;
	wire _w657_ ;
	wire _w656_ ;
	wire _w655_ ;
	wire _w654_ ;
	wire _w653_ ;
	wire _w652_ ;
	wire _w651_ ;
	wire _w650_ ;
	wire _w649_ ;
	wire _w648_ ;
	wire _w647_ ;
	wire _w646_ ;
	wire _w645_ ;
	wire _w644_ ;
	wire _w643_ ;
	wire _w642_ ;
	wire _w641_ ;
	wire _w640_ ;
	wire _w639_ ;
	wire _w638_ ;
	wire _w637_ ;
	wire _w636_ ;
	wire _w635_ ;
	wire _w634_ ;
	wire _w633_ ;
	wire _w632_ ;
	wire _w631_ ;
	wire _w630_ ;
	wire _w629_ ;
	wire _w628_ ;
	wire _w627_ ;
	wire _w626_ ;
	wire _w625_ ;
	wire _w624_ ;
	wire _w623_ ;
	wire _w622_ ;
	wire _w621_ ;
	wire _w620_ ;
	wire _w619_ ;
	wire _w618_ ;
	wire _w617_ ;
	wire _w332_ ;
	wire _w331_ ;
	wire _w330_ ;
	wire _w329_ ;
	wire _w328_ ;
	wire _w327_ ;
	wire _w326_ ;
	wire _w325_ ;
	wire _w324_ ;
	wire _w323_ ;
	wire _w322_ ;
	wire _w321_ ;
	wire _w320_ ;
	wire _w319_ ;
	wire _w318_ ;
	wire _w317_ ;
	wire _w316_ ;
	wire _w315_ ;
	wire _w314_ ;
	wire _w313_ ;
	wire _w312_ ;
	wire _w311_ ;
	wire _w310_ ;
	wire _w309_ ;
	wire _w308_ ;
	wire _w307_ ;
	wire _w306_ ;
	wire _w305_ ;
	wire _w304_ ;
	wire _w303_ ;
	wire _w302_ ;
	wire _w301_ ;
	wire _w300_ ;
	wire _w299_ ;
	wire _w298_ ;
	wire _w297_ ;
	wire _w296_ ;
	wire _w295_ ;
	wire _w294_ ;
	wire _w293_ ;
	wire _w292_ ;
	wire _w291_ ;
	wire _w290_ ;
	wire _w289_ ;
	wire _w288_ ;
	wire _w287_ ;
	wire _w286_ ;
	wire _w285_ ;
	wire _w284_ ;
	wire _w283_ ;
	wire _w282_ ;
	wire _w281_ ;
	wire _w280_ ;
	wire _w279_ ;
	wire _w278_ ;
	wire _w277_ ;
	wire _w276_ ;
	wire _w275_ ;
	wire _w274_ ;
	wire _w273_ ;
	wire _w272_ ;
	wire _w271_ ;
	wire _w270_ ;
	wire _w269_ ;
	wire _w268_ ;
	wire _w267_ ;
	wire _w266_ ;
	wire _w265_ ;
	wire _w264_ ;
	wire _w263_ ;
	wire _w262_ ;
	wire _w261_ ;
	wire _w260_ ;
	wire _w259_ ;
	wire _w258_ ;
	wire _w257_ ;
	wire _w256_ ;
	wire _w255_ ;
	wire _w254_ ;
	wire _w253_ ;
	wire _w252_ ;
	wire _w251_ ;
	wire _w250_ ;
	wire _w249_ ;
	wire _w248_ ;
	wire _w247_ ;
	wire _w246_ ;
	wire _w245_ ;
	wire _w244_ ;
	wire _w243_ ;
	wire _w242_ ;
	wire _w241_ ;
	wire _w240_ ;
	wire _w239_ ;
	wire _w238_ ;
	wire _w237_ ;
	wire _w236_ ;
	wire _w235_ ;
	wire _w234_ ;
	wire _w233_ ;
	wire _w232_ ;
	wire _w231_ ;
	wire _w230_ ;
	wire _w229_ ;
	wire _w228_ ;
	wire _w227_ ;
	wire _w226_ ;
	wire _w225_ ;
	wire _w224_ ;
	wire _w223_ ;
	wire _w222_ ;
	wire _w221_ ;
	wire _w220_ ;
	wire _w219_ ;
	wire _w218_ ;
	wire _w217_ ;
	wire _w216_ ;
	wire _w215_ ;
	wire _w214_ ;
	wire _w213_ ;
	wire _w212_ ;
	wire _w211_ ;
	wire _w210_ ;
	wire _w209_ ;
	wire _w208_ ;
	wire _w207_ ;
	wire _w206_ ;
	wire _w205_ ;
	wire _w204_ ;
	wire _w203_ ;
	wire _w134_ ;
	wire _w133_ ;
	wire _w132_ ;
	wire _w131_ ;
	wire _w130_ ;
	wire _w129_ ;
	wire _w128_ ;
	wire _w127_ ;
	wire _w126_ ;
	wire _w125_ ;
	wire _w124_ ;
	wire _w123_ ;
	wire _w122_ ;
	wire _w121_ ;
	wire _w120_ ;
	wire _w119_ ;
	wire _w118_ ;
	wire _w117_ ;
	wire _w116_ ;
	wire _w115_ ;
	wire _w114_ ;
	wire _w113_ ;
	wire _w112_ ;
	wire _w111_ ;
	wire _w110_ ;
	wire _w109_ ;
	wire _w108_ ;
	wire _w107_ ;
	wire _w106_ ;
	wire _w105_ ;
	wire _w88_ ;
	wire _w87_ ;
	wire _w86_ ;
	wire _w85_ ;
	wire _w84_ ;
	wire _w83_ ;
	wire _w82_ ;
	wire _w81_ ;
	wire _w80_ ;
	wire _w79_ ;
	wire _w78_ ;
	wire _w77_ ;
	wire _w76_ ;
	wire _w89_ ;
	wire _w90_ ;
	wire _w91_ ;
	wire _w92_ ;
	wire _w93_ ;
	wire _w94_ ;
	wire _w95_ ;
	wire _w96_ ;
	wire _w97_ ;
	wire _w98_ ;
	wire _w99_ ;
	wire _w100_ ;
	wire _w101_ ;
	wire _w102_ ;
	wire _w103_ ;
	wire _w104_ ;
	wire _w135_ ;
	wire _w136_ ;
	wire _w137_ ;
	wire _w138_ ;
	wire _w139_ ;
	wire _w140_ ;
	wire _w141_ ;
	wire _w142_ ;
	wire _w143_ ;
	wire _w144_ ;
	wire _w145_ ;
	wire _w146_ ;
	wire _w147_ ;
	wire _w148_ ;
	wire _w149_ ;
	wire _w150_ ;
	wire _w151_ ;
	wire _w152_ ;
	wire _w153_ ;
	wire _w154_ ;
	wire _w155_ ;
	wire _w156_ ;
	wire _w157_ ;
	wire _w158_ ;
	wire _w159_ ;
	wire _w160_ ;
	wire _w161_ ;
	wire _w162_ ;
	wire _w163_ ;
	wire _w164_ ;
	wire _w165_ ;
	wire _w166_ ;
	wire _w167_ ;
	wire _w168_ ;
	wire _w169_ ;
	wire _w170_ ;
	wire _w171_ ;
	wire _w172_ ;
	wire _w173_ ;
	wire _w174_ ;
	wire _w175_ ;
	wire _w176_ ;
	wire _w177_ ;
	wire _w178_ ;
	wire _w179_ ;
	wire _w180_ ;
	wire _w181_ ;
	wire _w182_ ;
	wire _w183_ ;
	wire _w184_ ;
	wire _w185_ ;
	wire _w186_ ;
	wire _w187_ ;
	wire _w188_ ;
	wire _w189_ ;
	wire _w190_ ;
	wire _w191_ ;
	wire _w192_ ;
	wire _w193_ ;
	wire _w194_ ;
	wire _w195_ ;
	wire _w196_ ;
	wire _w197_ ;
	wire _w198_ ;
	wire _w199_ ;
	wire _w200_ ;
	wire _w201_ ;
	wire _w202_ ;
	wire _w333_ ;
	wire _w334_ ;
	wire _w335_ ;
	wire _w336_ ;
	wire _w337_ ;
	wire _w338_ ;
	wire _w339_ ;
	wire _w340_ ;
	wire _w341_ ;
	wire _w342_ ;
	wire _w343_ ;
	wire _w344_ ;
	wire _w345_ ;
	wire _w346_ ;
	wire _w347_ ;
	wire _w348_ ;
	wire _w349_ ;
	wire _w350_ ;
	wire _w351_ ;
	wire _w352_ ;
	wire _w353_ ;
	wire _w354_ ;
	wire _w355_ ;
	wire _w356_ ;
	wire _w357_ ;
	wire _w358_ ;
	wire _w359_ ;
	wire _w360_ ;
	wire _w361_ ;
	wire _w362_ ;
	wire _w363_ ;
	wire _w364_ ;
	wire _w365_ ;
	wire _w366_ ;
	wire _w367_ ;
	wire _w368_ ;
	wire _w369_ ;
	wire _w370_ ;
	wire _w371_ ;
	wire _w372_ ;
	wire _w373_ ;
	wire _w374_ ;
	wire _w375_ ;
	wire _w376_ ;
	wire _w377_ ;
	wire _w378_ ;
	wire _w379_ ;
	wire _w380_ ;
	wire _w381_ ;
	wire _w382_ ;
	wire _w383_ ;
	wire _w384_ ;
	wire _w385_ ;
	wire _w386_ ;
	wire _w387_ ;
	wire _w388_ ;
	wire _w389_ ;
	wire _w390_ ;
	wire _w391_ ;
	wire _w392_ ;
	wire _w393_ ;
	wire _w394_ ;
	wire _w395_ ;
	wire _w396_ ;
	wire _w397_ ;
	wire _w398_ ;
	wire _w399_ ;
	wire _w400_ ;
	wire _w401_ ;
	wire _w402_ ;
	wire _w403_ ;
	wire _w404_ ;
	wire _w405_ ;
	wire _w406_ ;
	wire _w407_ ;
	wire _w408_ ;
	wire _w409_ ;
	wire _w410_ ;
	wire _w411_ ;
	wire _w412_ ;
	wire _w413_ ;
	wire _w414_ ;
	wire _w415_ ;
	wire _w416_ ;
	wire _w417_ ;
	wire _w418_ ;
	wire _w419_ ;
	wire _w420_ ;
	wire _w421_ ;
	wire _w422_ ;
	wire _w423_ ;
	wire _w424_ ;
	wire _w425_ ;
	wire _w426_ ;
	wire _w427_ ;
	wire _w428_ ;
	wire _w429_ ;
	wire _w430_ ;
	wire _w431_ ;
	wire _w432_ ;
	wire _w433_ ;
	wire _w434_ ;
	wire _w435_ ;
	wire _w436_ ;
	wire _w437_ ;
	wire _w438_ ;
	wire _w439_ ;
	wire _w440_ ;
	wire _w441_ ;
	wire _w442_ ;
	wire _w443_ ;
	wire _w444_ ;
	wire _w445_ ;
	wire _w446_ ;
	wire _w447_ ;
	wire _w448_ ;
	wire _w449_ ;
	wire _w450_ ;
	wire _w451_ ;
	wire _w452_ ;
	wire _w453_ ;
	wire _w454_ ;
	wire _w455_ ;
	wire _w456_ ;
	wire _w457_ ;
	wire _w458_ ;
	wire _w459_ ;
	wire _w460_ ;
	wire _w461_ ;
	wire _w462_ ;
	wire _w463_ ;
	wire _w464_ ;
	wire _w465_ ;
	wire _w466_ ;
	wire _w467_ ;
	wire _w468_ ;
	wire _w469_ ;
	wire _w470_ ;
	wire _w471_ ;
	wire _w472_ ;
	wire _w473_ ;
	wire _w474_ ;
	wire _w475_ ;
	wire _w476_ ;
	wire _w477_ ;
	wire _w478_ ;
	wire _w479_ ;
	wire _w480_ ;
	wire _w481_ ;
	wire _w482_ ;
	wire _w483_ ;
	wire _w484_ ;
	wire _w485_ ;
	wire _w486_ ;
	wire _w487_ ;
	wire _w488_ ;
	wire _w489_ ;
	wire _w490_ ;
	wire _w491_ ;
	wire _w492_ ;
	wire _w493_ ;
	wire _w494_ ;
	wire _w495_ ;
	wire _w496_ ;
	wire _w497_ ;
	wire _w498_ ;
	wire _w499_ ;
	wire _w500_ ;
	wire _w501_ ;
	wire _w502_ ;
	wire _w503_ ;
	wire _w504_ ;
	wire _w505_ ;
	wire _w506_ ;
	wire _w507_ ;
	wire _w508_ ;
	wire _w509_ ;
	wire _w510_ ;
	wire _w511_ ;
	wire _w512_ ;
	wire _w513_ ;
	wire _w514_ ;
	wire _w515_ ;
	wire _w516_ ;
	wire _w517_ ;
	wire _w518_ ;
	wire _w519_ ;
	wire _w520_ ;
	wire _w521_ ;
	wire _w522_ ;
	wire _w523_ ;
	wire _w524_ ;
	wire _w525_ ;
	wire _w526_ ;
	wire _w527_ ;
	wire _w528_ ;
	wire _w529_ ;
	wire _w530_ ;
	wire _w531_ ;
	wire _w532_ ;
	wire _w533_ ;
	wire _w534_ ;
	wire _w535_ ;
	wire _w536_ ;
	wire _w537_ ;
	wire _w538_ ;
	wire _w539_ ;
	wire _w540_ ;
	wire _w541_ ;
	wire _w542_ ;
	wire _w543_ ;
	wire _w544_ ;
	wire _w545_ ;
	wire _w546_ ;
	wire _w547_ ;
	wire _w548_ ;
	wire _w549_ ;
	wire _w550_ ;
	wire _w551_ ;
	wire _w552_ ;
	wire _w553_ ;
	wire _w554_ ;
	wire _w555_ ;
	wire _w556_ ;
	wire _w557_ ;
	wire _w558_ ;
	wire _w559_ ;
	wire _w560_ ;
	wire _w561_ ;
	wire _w562_ ;
	wire _w563_ ;
	wire _w564_ ;
	wire _w565_ ;
	wire _w566_ ;
	wire _w567_ ;
	wire _w568_ ;
	wire _w569_ ;
	wire _w570_ ;
	wire _w571_ ;
	wire _w572_ ;
	wire _w573_ ;
	wire _w574_ ;
	wire _w575_ ;
	wire _w576_ ;
	wire _w577_ ;
	wire _w578_ ;
	wire _w579_ ;
	wire _w580_ ;
	wire _w581_ ;
	wire _w582_ ;
	wire _w583_ ;
	wire _w584_ ;
	wire _w585_ ;
	wire _w586_ ;
	wire _w587_ ;
	wire _w588_ ;
	wire _w589_ ;
	wire _w590_ ;
	wire _w591_ ;
	wire _w592_ ;
	wire _w593_ ;
	wire _w594_ ;
	wire _w595_ ;
	wire _w596_ ;
	wire _w597_ ;
	wire _w598_ ;
	wire _w599_ ;
	wire _w600_ ;
	wire _w601_ ;
	wire _w602_ ;
	wire _w603_ ;
	wire _w604_ ;
	wire _w605_ ;
	wire _w606_ ;
	wire _w607_ ;
	wire _w608_ ;
	wire _w609_ ;
	wire _w610_ ;
	wire _w611_ ;
	wire _w612_ ;
	wire _w613_ ;
	wire _w614_ ;
	wire _w615_ ;
	wire _w616_ ;
	LUT2 #(
		.INIT('h4)
	) name0 (
		\opsel2_pad ,
		\opsel3_pad ,
		_w76_
	);
	LUT2 #(
		.INIT('h4)
	) name1 (
		\musel3_pad ,
		\musel4_pad ,
		_w77_
	);
	LUT2 #(
		.INIT('h1)
	) name2 (
		\musel1_pad ,
		\musel2_pad ,
		_w78_
	);
	LUT2 #(
		.INIT('h8)
	) name3 (
		_w77_,
		_w78_,
		_w79_
	);
	LUT2 #(
		.INIT('h8)
	) name4 (
		\inD3_pad ,
		_w79_,
		_w80_
	);
	LUT2 #(
		.INIT('h2)
	) name5 (
		\musel3_pad ,
		\musel4_pad ,
		_w81_
	);
	LUT2 #(
		.INIT('h8)
	) name6 (
		\musel1_pad ,
		\musel2_pad ,
		_w82_
	);
	LUT2 #(
		.INIT('h1)
	) name7 (
		_w78_,
		_w82_,
		_w83_
	);
	LUT2 #(
		.INIT('h8)
	) name8 (
		\inB3_pad ,
		_w83_,
		_w84_
	);
	LUT2 #(
		.INIT('h8)
	) name9 (
		\inD3_pad ,
		_w82_,
		_w85_
	);
	LUT2 #(
		.INIT('h1)
	) name10 (
		_w84_,
		_w85_,
		_w86_
	);
	LUT2 #(
		.INIT('h2)
	) name11 (
		_w81_,
		_w86_,
		_w87_
	);
	LUT2 #(
		.INIT('h1)
	) name12 (
		_w80_,
		_w87_,
		_w88_
	);
	LUT2 #(
		.INIT('h1)
	) name13 (
		\sh2_pad ,
		_w88_,
		_w89_
	);
	LUT2 #(
		.INIT('h8)
	) name14 (
		\inD0_pad ,
		_w79_,
		_w90_
	);
	LUT2 #(
		.INIT('h8)
	) name15 (
		\inB0_pad ,
		_w83_,
		_w91_
	);
	LUT2 #(
		.INIT('h8)
	) name16 (
		\inD0_pad ,
		_w82_,
		_w92_
	);
	LUT2 #(
		.INIT('h1)
	) name17 (
		_w91_,
		_w92_,
		_w93_
	);
	LUT2 #(
		.INIT('h2)
	) name18 (
		_w81_,
		_w93_,
		_w94_
	);
	LUT2 #(
		.INIT('h1)
	) name19 (
		_w90_,
		_w94_,
		_w95_
	);
	LUT2 #(
		.INIT('h2)
	) name20 (
		\sh2_pad ,
		_w95_,
		_w96_
	);
	LUT2 #(
		.INIT('h1)
	) name21 (
		_w89_,
		_w96_,
		_w97_
	);
	LUT2 #(
		.INIT('h2)
	) name22 (
		\sh1_pad ,
		_w97_,
		_w98_
	);
	LUT2 #(
		.INIT('h8)
	) name23 (
		\inD5_pad ,
		_w79_,
		_w99_
	);
	LUT2 #(
		.INIT('h8)
	) name24 (
		\inB5_pad ,
		_w83_,
		_w100_
	);
	LUT2 #(
		.INIT('h8)
	) name25 (
		\inD5_pad ,
		_w82_,
		_w101_
	);
	LUT2 #(
		.INIT('h1)
	) name26 (
		_w100_,
		_w101_,
		_w102_
	);
	LUT2 #(
		.INIT('h2)
	) name27 (
		_w81_,
		_w102_,
		_w103_
	);
	LUT2 #(
		.INIT('h1)
	) name28 (
		_w99_,
		_w103_,
		_w104_
	);
	LUT2 #(
		.INIT('h2)
	) name29 (
		\sh2_pad ,
		_w104_,
		_w105_
	);
	LUT2 #(
		.INIT('h8)
	) name30 (
		\inD1_pad ,
		_w79_,
		_w106_
	);
	LUT2 #(
		.INIT('h8)
	) name31 (
		\inB1_pad ,
		_w83_,
		_w107_
	);
	LUT2 #(
		.INIT('h8)
	) name32 (
		\inD1_pad ,
		_w82_,
		_w108_
	);
	LUT2 #(
		.INIT('h1)
	) name33 (
		_w107_,
		_w108_,
		_w109_
	);
	LUT2 #(
		.INIT('h2)
	) name34 (
		_w81_,
		_w109_,
		_w110_
	);
	LUT2 #(
		.INIT('h1)
	) name35 (
		_w106_,
		_w110_,
		_w111_
	);
	LUT2 #(
		.INIT('h1)
	) name36 (
		\sh2_pad ,
		_w111_,
		_w112_
	);
	LUT2 #(
		.INIT('h1)
	) name37 (
		_w105_,
		_w112_,
		_w113_
	);
	LUT2 #(
		.INIT('h1)
	) name38 (
		\sh1_pad ,
		_w113_,
		_w114_
	);
	LUT2 #(
		.INIT('h1)
	) name39 (
		_w98_,
		_w114_,
		_w115_
	);
	LUT2 #(
		.INIT('h2)
	) name40 (
		\sh0_pad ,
		_w115_,
		_w116_
	);
	LUT2 #(
		.INIT('h8)
	) name41 (
		\inD8_pad ,
		_w79_,
		_w117_
	);
	LUT2 #(
		.INIT('h8)
	) name42 (
		\inB8_pad ,
		_w83_,
		_w118_
	);
	LUT2 #(
		.INIT('h8)
	) name43 (
		\inD8_pad ,
		_w82_,
		_w119_
	);
	LUT2 #(
		.INIT('h1)
	) name44 (
		_w118_,
		_w119_,
		_w120_
	);
	LUT2 #(
		.INIT('h2)
	) name45 (
		_w81_,
		_w120_,
		_w121_
	);
	LUT2 #(
		.INIT('h1)
	) name46 (
		_w117_,
		_w121_,
		_w122_
	);
	LUT2 #(
		.INIT('h2)
	) name47 (
		\sh2_pad ,
		_w122_,
		_w123_
	);
	LUT2 #(
		.INIT('h8)
	) name48 (
		\inD2_pad ,
		_w79_,
		_w124_
	);
	LUT2 #(
		.INIT('h8)
	) name49 (
		\inB2_pad ,
		_w83_,
		_w125_
	);
	LUT2 #(
		.INIT('h8)
	) name50 (
		\inD2_pad ,
		_w82_,
		_w126_
	);
	LUT2 #(
		.INIT('h1)
	) name51 (
		_w125_,
		_w126_,
		_w127_
	);
	LUT2 #(
		.INIT('h2)
	) name52 (
		_w81_,
		_w127_,
		_w128_
	);
	LUT2 #(
		.INIT('h1)
	) name53 (
		_w124_,
		_w128_,
		_w129_
	);
	LUT2 #(
		.INIT('h1)
	) name54 (
		\sh2_pad ,
		_w129_,
		_w130_
	);
	LUT2 #(
		.INIT('h2)
	) name55 (
		\sh1_pad ,
		_w123_,
		_w131_
	);
	LUT2 #(
		.INIT('h4)
	) name56 (
		_w130_,
		_w131_,
		_w132_
	);
	LUT2 #(
		.INIT('h1)
	) name57 (
		\sh2_pad ,
		_w95_,
		_w133_
	);
	LUT2 #(
		.INIT('h8)
	) name58 (
		\inD4_pad ,
		_w79_,
		_w134_
	);
	LUT2 #(
		.INIT('h8)
	) name59 (
		\inB4_pad ,
		_w83_,
		_w135_
	);
	LUT2 #(
		.INIT('h8)
	) name60 (
		\inD4_pad ,
		_w82_,
		_w136_
	);
	LUT2 #(
		.INIT('h1)
	) name61 (
		_w135_,
		_w136_,
		_w137_
	);
	LUT2 #(
		.INIT('h2)
	) name62 (
		_w81_,
		_w137_,
		_w138_
	);
	LUT2 #(
		.INIT('h1)
	) name63 (
		_w134_,
		_w138_,
		_w139_
	);
	LUT2 #(
		.INIT('h2)
	) name64 (
		\sh2_pad ,
		_w139_,
		_w140_
	);
	LUT2 #(
		.INIT('h1)
	) name65 (
		\sh1_pad ,
		_w133_,
		_w141_
	);
	LUT2 #(
		.INIT('h4)
	) name66 (
		_w140_,
		_w141_,
		_w142_
	);
	LUT2 #(
		.INIT('h1)
	) name67 (
		\sh0_pad ,
		_w132_,
		_w143_
	);
	LUT2 #(
		.INIT('h4)
	) name68 (
		_w142_,
		_w143_,
		_w144_
	);
	LUT2 #(
		.INIT('h1)
	) name69 (
		_w116_,
		_w144_,
		_w145_
	);
	LUT2 #(
		.INIT('h1)
	) name70 (
		\opsel0_pad ,
		\opsel1_pad ,
		_w146_
	);
	LUT2 #(
		.INIT('h4)
	) name71 (
		_w145_,
		_w146_,
		_w147_
	);
	LUT2 #(
		.INIT('h8)
	) name72 (
		\opsel0_pad ,
		\opsel1_pad ,
		_w148_
	);
	LUT2 #(
		.INIT('h1)
	) name73 (
		_w146_,
		_w148_,
		_w149_
	);
	LUT2 #(
		.INIT('h4)
	) name74 (
		\musel2_pad ,
		\musel3_pad ,
		_w150_
	);
	LUT2 #(
		.INIT('h8)
	) name75 (
		\inD0_pad ,
		_w150_,
		_w151_
	);
	LUT2 #(
		.INIT('h2)
	) name76 (
		\musel2_pad ,
		\musel3_pad ,
		_w152_
	);
	LUT2 #(
		.INIT('h8)
	) name77 (
		\inB0_pad ,
		_w152_,
		_w153_
	);
	LUT2 #(
		.INIT('h1)
	) name78 (
		_w151_,
		_w153_,
		_w154_
	);
	LUT2 #(
		.INIT('h1)
	) name79 (
		\musel1_pad ,
		_w154_,
		_w155_
	);
	LUT2 #(
		.INIT('h2)
	) name80 (
		\musel1_pad ,
		\musel3_pad ,
		_w156_
	);
	LUT2 #(
		.INIT('h2)
	) name81 (
		\inA0_pad ,
		\musel2_pad ,
		_w157_
	);
	LUT2 #(
		.INIT('h8)
	) name82 (
		\inC0_pad ,
		\musel2_pad ,
		_w158_
	);
	LUT2 #(
		.INIT('h1)
	) name83 (
		_w157_,
		_w158_,
		_w159_
	);
	LUT2 #(
		.INIT('h2)
	) name84 (
		_w156_,
		_w159_,
		_w160_
	);
	LUT2 #(
		.INIT('h1)
	) name85 (
		_w155_,
		_w160_,
		_w161_
	);
	LUT2 #(
		.INIT('h1)
	) name86 (
		\musel4_pad ,
		_w161_,
		_w162_
	);
	LUT2 #(
		.INIT('h8)
	) name87 (
		\inC0_pad ,
		_w79_,
		_w163_
	);
	LUT2 #(
		.INIT('h8)
	) name88 (
		\inA0_pad ,
		_w83_,
		_w164_
	);
	LUT2 #(
		.INIT('h8)
	) name89 (
		\musel1_pad ,
		_w158_,
		_w165_
	);
	LUT2 #(
		.INIT('h1)
	) name90 (
		_w164_,
		_w165_,
		_w166_
	);
	LUT2 #(
		.INIT('h2)
	) name91 (
		_w81_,
		_w166_,
		_w167_
	);
	LUT2 #(
		.INIT('h1)
	) name92 (
		_w163_,
		_w167_,
		_w168_
	);
	LUT2 #(
		.INIT('h1)
	) name93 (
		_w162_,
		_w168_,
		_w169_
	);
	LUT2 #(
		.INIT('h8)
	) name94 (
		_w162_,
		_w168_,
		_w170_
	);
	LUT2 #(
		.INIT('h1)
	) name95 (
		_w169_,
		_w170_,
		_w171_
	);
	LUT2 #(
		.INIT('h2)
	) name96 (
		_w149_,
		_w171_,
		_w172_
	);
	LUT2 #(
		.INIT('h1)
	) name97 (
		_w147_,
		_w172_,
		_w173_
	);
	LUT2 #(
		.INIT('h2)
	) name98 (
		_w76_,
		_w173_,
		_w174_
	);
	LUT2 #(
		.INIT('h2)
	) name99 (
		\opsel2_pad ,
		_w146_,
		_w175_
	);
	LUT2 #(
		.INIT('h2)
	) name100 (
		\inC0_pad ,
		\musel1_pad ,
		_w176_
	);
	LUT2 #(
		.INIT('h1)
	) name101 (
		_w157_,
		_w176_,
		_w177_
	);
	LUT2 #(
		.INIT('h2)
	) name102 (
		_w77_,
		_w78_,
		_w178_
	);
	LUT2 #(
		.INIT('h4)
	) name103 (
		_w177_,
		_w178_,
		_w179_
	);
	LUT2 #(
		.INIT('h1)
	) name104 (
		_w175_,
		_w179_,
		_w180_
	);
	LUT2 #(
		.INIT('h8)
	) name105 (
		_w145_,
		_w175_,
		_w181_
	);
	LUT2 #(
		.INIT('h4)
	) name106 (
		\opsel2_pad ,
		_w146_,
		_w182_
	);
	LUT2 #(
		.INIT('h1)
	) name107 (
		\opsel3_pad ,
		_w182_,
		_w183_
	);
	LUT2 #(
		.INIT('h4)
	) name108 (
		_w180_,
		_w183_,
		_w184_
	);
	LUT2 #(
		.INIT('h4)
	) name109 (
		_w181_,
		_w184_,
		_w185_
	);
	LUT2 #(
		.INIT('h1)
	) name110 (
		_w174_,
		_w185_,
		_w186_
	);
	LUT2 #(
		.INIT('h8)
	) name111 (
		\inD14_pad ,
		_w79_,
		_w187_
	);
	LUT2 #(
		.INIT('h8)
	) name112 (
		\inB14_pad ,
		_w83_,
		_w188_
	);
	LUT2 #(
		.INIT('h8)
	) name113 (
		\inD14_pad ,
		_w82_,
		_w189_
	);
	LUT2 #(
		.INIT('h1)
	) name114 (
		_w188_,
		_w189_,
		_w190_
	);
	LUT2 #(
		.INIT('h2)
	) name115 (
		_w81_,
		_w190_,
		_w191_
	);
	LUT2 #(
		.INIT('h1)
	) name116 (
		_w187_,
		_w191_,
		_w192_
	);
	LUT2 #(
		.INIT('h2)
	) name117 (
		\sh2_pad ,
		_w192_,
		_w193_
	);
	LUT2 #(
		.INIT('h8)
	) name118 (
		\inD10_pad ,
		_w79_,
		_w194_
	);
	LUT2 #(
		.INIT('h8)
	) name119 (
		\inB10_pad ,
		_w83_,
		_w195_
	);
	LUT2 #(
		.INIT('h8)
	) name120 (
		\inD10_pad ,
		_w82_,
		_w196_
	);
	LUT2 #(
		.INIT('h1)
	) name121 (
		_w195_,
		_w196_,
		_w197_
	);
	LUT2 #(
		.INIT('h2)
	) name122 (
		_w81_,
		_w197_,
		_w198_
	);
	LUT2 #(
		.INIT('h1)
	) name123 (
		_w194_,
		_w198_,
		_w199_
	);
	LUT2 #(
		.INIT('h1)
	) name124 (
		\sh2_pad ,
		_w199_,
		_w200_
	);
	LUT2 #(
		.INIT('h1)
	) name125 (
		_w193_,
		_w200_,
		_w201_
	);
	LUT2 #(
		.INIT('h1)
	) name126 (
		\sh1_pad ,
		_w201_,
		_w202_
	);
	LUT2 #(
		.INIT('h8)
	) name127 (
		\inD12_pad ,
		_w79_,
		_w203_
	);
	LUT2 #(
		.INIT('h8)
	) name128 (
		\inB12_pad ,
		_w83_,
		_w204_
	);
	LUT2 #(
		.INIT('h8)
	) name129 (
		\inD12_pad ,
		_w82_,
		_w205_
	);
	LUT2 #(
		.INIT('h1)
	) name130 (
		_w204_,
		_w205_,
		_w206_
	);
	LUT2 #(
		.INIT('h2)
	) name131 (
		_w81_,
		_w206_,
		_w207_
	);
	LUT2 #(
		.INIT('h1)
	) name132 (
		_w203_,
		_w207_,
		_w208_
	);
	LUT2 #(
		.INIT('h1)
	) name133 (
		\sh2_pad ,
		_w208_,
		_w209_
	);
	LUT2 #(
		.INIT('h8)
	) name134 (
		\inD15_pad ,
		_w79_,
		_w210_
	);
	LUT2 #(
		.INIT('h8)
	) name135 (
		\inB15_pad ,
		_w83_,
		_w211_
	);
	LUT2 #(
		.INIT('h8)
	) name136 (
		\inD15_pad ,
		_w82_,
		_w212_
	);
	LUT2 #(
		.INIT('h1)
	) name137 (
		_w211_,
		_w212_,
		_w213_
	);
	LUT2 #(
		.INIT('h2)
	) name138 (
		_w81_,
		_w213_,
		_w214_
	);
	LUT2 #(
		.INIT('h1)
	) name139 (
		_w210_,
		_w214_,
		_w215_
	);
	LUT2 #(
		.INIT('h2)
	) name140 (
		\sh2_pad ,
		_w215_,
		_w216_
	);
	LUT2 #(
		.INIT('h1)
	) name141 (
		_w209_,
		_w216_,
		_w217_
	);
	LUT2 #(
		.INIT('h2)
	) name142 (
		\sh1_pad ,
		_w217_,
		_w218_
	);
	LUT2 #(
		.INIT('h1)
	) name143 (
		_w202_,
		_w218_,
		_w219_
	);
	LUT2 #(
		.INIT('h1)
	) name144 (
		\sh0_pad ,
		_w219_,
		_w220_
	);
	LUT2 #(
		.INIT('h2)
	) name145 (
		\sh2_pad ,
		_w199_,
		_w221_
	);
	LUT2 #(
		.INIT('h8)
	) name146 (
		\inD13_pad ,
		_w79_,
		_w222_
	);
	LUT2 #(
		.INIT('h8)
	) name147 (
		\inB13_pad ,
		_w83_,
		_w223_
	);
	LUT2 #(
		.INIT('h8)
	) name148 (
		\inD13_pad ,
		_w82_,
		_w224_
	);
	LUT2 #(
		.INIT('h1)
	) name149 (
		_w223_,
		_w224_,
		_w225_
	);
	LUT2 #(
		.INIT('h2)
	) name150 (
		_w81_,
		_w225_,
		_w226_
	);
	LUT2 #(
		.INIT('h1)
	) name151 (
		_w222_,
		_w226_,
		_w227_
	);
	LUT2 #(
		.INIT('h1)
	) name152 (
		\sh2_pad ,
		_w227_,
		_w228_
	);
	LUT2 #(
		.INIT('h2)
	) name153 (
		\sh1_pad ,
		_w221_,
		_w229_
	);
	LUT2 #(
		.INIT('h4)
	) name154 (
		_w228_,
		_w229_,
		_w230_
	);
	LUT2 #(
		.INIT('h8)
	) name155 (
		\inD11_pad ,
		_w79_,
		_w231_
	);
	LUT2 #(
		.INIT('h8)
	) name156 (
		\inB11_pad ,
		_w83_,
		_w232_
	);
	LUT2 #(
		.INIT('h8)
	) name157 (
		\inD11_pad ,
		_w82_,
		_w233_
	);
	LUT2 #(
		.INIT('h1)
	) name158 (
		_w232_,
		_w233_,
		_w234_
	);
	LUT2 #(
		.INIT('h2)
	) name159 (
		_w81_,
		_w234_,
		_w235_
	);
	LUT2 #(
		.INIT('h1)
	) name160 (
		_w231_,
		_w235_,
		_w236_
	);
	LUT2 #(
		.INIT('h1)
	) name161 (
		\sh2_pad ,
		_w236_,
		_w237_
	);
	LUT2 #(
		.INIT('h1)
	) name162 (
		_w216_,
		_w237_,
		_w238_
	);
	LUT2 #(
		.INIT('h4)
	) name163 (
		\sh1_pad ,
		_w238_,
		_w239_
	);
	LUT2 #(
		.INIT('h2)
	) name164 (
		\sh0_pad ,
		_w230_,
		_w240_
	);
	LUT2 #(
		.INIT('h4)
	) name165 (
		_w239_,
		_w240_,
		_w241_
	);
	LUT2 #(
		.INIT('h1)
	) name166 (
		_w220_,
		_w241_,
		_w242_
	);
	LUT2 #(
		.INIT('h2)
	) name167 (
		_w146_,
		_w242_,
		_w243_
	);
	LUT2 #(
		.INIT('h8)
	) name168 (
		\inC9_pad ,
		_w79_,
		_w244_
	);
	LUT2 #(
		.INIT('h8)
	) name169 (
		\inA9_pad ,
		_w83_,
		_w245_
	);
	LUT2 #(
		.INIT('h8)
	) name170 (
		\inC9_pad ,
		\musel2_pad ,
		_w246_
	);
	LUT2 #(
		.INIT('h8)
	) name171 (
		\musel1_pad ,
		_w246_,
		_w247_
	);
	LUT2 #(
		.INIT('h1)
	) name172 (
		_w245_,
		_w247_,
		_w248_
	);
	LUT2 #(
		.INIT('h2)
	) name173 (
		_w81_,
		_w248_,
		_w249_
	);
	LUT2 #(
		.INIT('h1)
	) name174 (
		_w244_,
		_w249_,
		_w250_
	);
	LUT2 #(
		.INIT('h1)
	) name175 (
		\opsel1_pad ,
		_w76_,
		_w251_
	);
	LUT2 #(
		.INIT('h2)
	) name176 (
		\opsel2_pad ,
		\opsel3_pad ,
		_w252_
	);
	LUT2 #(
		.INIT('h2)
	) name177 (
		\opsel1_pad ,
		_w252_,
		_w253_
	);
	LUT2 #(
		.INIT('h1)
	) name178 (
		\opsel0_pad ,
		_w251_,
		_w254_
	);
	LUT2 #(
		.INIT('h4)
	) name179 (
		_w253_,
		_w254_,
		_w255_
	);
	LUT2 #(
		.INIT('h1)
	) name180 (
		_w250_,
		_w255_,
		_w256_
	);
	LUT2 #(
		.INIT('h8)
	) name181 (
		_w250_,
		_w255_,
		_w257_
	);
	LUT2 #(
		.INIT('h1)
	) name182 (
		_w256_,
		_w257_,
		_w258_
	);
	LUT2 #(
		.INIT('h8)
	) name183 (
		\inD9_pad ,
		_w150_,
		_w259_
	);
	LUT2 #(
		.INIT('h8)
	) name184 (
		\inB9_pad ,
		_w152_,
		_w260_
	);
	LUT2 #(
		.INIT('h1)
	) name185 (
		_w259_,
		_w260_,
		_w261_
	);
	LUT2 #(
		.INIT('h1)
	) name186 (
		\musel1_pad ,
		_w261_,
		_w262_
	);
	LUT2 #(
		.INIT('h2)
	) name187 (
		\inA9_pad ,
		\musel2_pad ,
		_w263_
	);
	LUT2 #(
		.INIT('h1)
	) name188 (
		_w246_,
		_w263_,
		_w264_
	);
	LUT2 #(
		.INIT('h2)
	) name189 (
		_w156_,
		_w264_,
		_w265_
	);
	LUT2 #(
		.INIT('h1)
	) name190 (
		_w262_,
		_w265_,
		_w266_
	);
	LUT2 #(
		.INIT('h1)
	) name191 (
		\musel4_pad ,
		_w266_,
		_w267_
	);
	LUT2 #(
		.INIT('h2)
	) name192 (
		_w258_,
		_w267_,
		_w268_
	);
	LUT2 #(
		.INIT('h4)
	) name193 (
		_w258_,
		_w267_,
		_w269_
	);
	LUT2 #(
		.INIT('h8)
	) name194 (
		\inC8_pad ,
		_w79_,
		_w270_
	);
	LUT2 #(
		.INIT('h8)
	) name195 (
		\inA8_pad ,
		_w83_,
		_w271_
	);
	LUT2 #(
		.INIT('h8)
	) name196 (
		\inC8_pad ,
		\musel2_pad ,
		_w272_
	);
	LUT2 #(
		.INIT('h8)
	) name197 (
		\musel1_pad ,
		_w272_,
		_w273_
	);
	LUT2 #(
		.INIT('h1)
	) name198 (
		_w271_,
		_w273_,
		_w274_
	);
	LUT2 #(
		.INIT('h2)
	) name199 (
		_w81_,
		_w274_,
		_w275_
	);
	LUT2 #(
		.INIT('h1)
	) name200 (
		_w270_,
		_w275_,
		_w276_
	);
	LUT2 #(
		.INIT('h1)
	) name201 (
		_w255_,
		_w276_,
		_w277_
	);
	LUT2 #(
		.INIT('h8)
	) name202 (
		_w255_,
		_w276_,
		_w278_
	);
	LUT2 #(
		.INIT('h1)
	) name203 (
		_w277_,
		_w278_,
		_w279_
	);
	LUT2 #(
		.INIT('h8)
	) name204 (
		\inD8_pad ,
		_w150_,
		_w280_
	);
	LUT2 #(
		.INIT('h8)
	) name205 (
		\inB8_pad ,
		_w152_,
		_w281_
	);
	LUT2 #(
		.INIT('h1)
	) name206 (
		_w280_,
		_w281_,
		_w282_
	);
	LUT2 #(
		.INIT('h1)
	) name207 (
		\musel1_pad ,
		_w282_,
		_w283_
	);
	LUT2 #(
		.INIT('h2)
	) name208 (
		\inA8_pad ,
		\musel2_pad ,
		_w284_
	);
	LUT2 #(
		.INIT('h1)
	) name209 (
		_w272_,
		_w284_,
		_w285_
	);
	LUT2 #(
		.INIT('h2)
	) name210 (
		_w156_,
		_w285_,
		_w286_
	);
	LUT2 #(
		.INIT('h1)
	) name211 (
		_w283_,
		_w286_,
		_w287_
	);
	LUT2 #(
		.INIT('h1)
	) name212 (
		\musel4_pad ,
		_w287_,
		_w288_
	);
	LUT2 #(
		.INIT('h2)
	) name213 (
		_w279_,
		_w288_,
		_w289_
	);
	LUT2 #(
		.INIT('h4)
	) name214 (
		_w279_,
		_w288_,
		_w290_
	);
	LUT2 #(
		.INIT('h8)
	) name215 (
		\inC4_pad ,
		_w79_,
		_w291_
	);
	LUT2 #(
		.INIT('h4)
	) name216 (
		\inA4_pad ,
		_w83_,
		_w292_
	);
	LUT2 #(
		.INIT('h8)
	) name217 (
		\inC4_pad ,
		\musel2_pad ,
		_w293_
	);
	LUT2 #(
		.INIT('h1)
	) name218 (
		_w83_,
		_w293_,
		_w294_
	);
	LUT2 #(
		.INIT('h2)
	) name219 (
		_w81_,
		_w292_,
		_w295_
	);
	LUT2 #(
		.INIT('h4)
	) name220 (
		_w294_,
		_w295_,
		_w296_
	);
	LUT2 #(
		.INIT('h1)
	) name221 (
		_w291_,
		_w296_,
		_w297_
	);
	LUT2 #(
		.INIT('h1)
	) name222 (
		_w255_,
		_w297_,
		_w298_
	);
	LUT2 #(
		.INIT('h8)
	) name223 (
		_w255_,
		_w297_,
		_w299_
	);
	LUT2 #(
		.INIT('h1)
	) name224 (
		_w298_,
		_w299_,
		_w300_
	);
	LUT2 #(
		.INIT('h8)
	) name225 (
		\inD4_pad ,
		_w150_,
		_w301_
	);
	LUT2 #(
		.INIT('h8)
	) name226 (
		\inB4_pad ,
		_w152_,
		_w302_
	);
	LUT2 #(
		.INIT('h1)
	) name227 (
		_w301_,
		_w302_,
		_w303_
	);
	LUT2 #(
		.INIT('h1)
	) name228 (
		\musel1_pad ,
		_w303_,
		_w304_
	);
	LUT2 #(
		.INIT('h2)
	) name229 (
		\inA4_pad ,
		\musel2_pad ,
		_w305_
	);
	LUT2 #(
		.INIT('h1)
	) name230 (
		_w293_,
		_w305_,
		_w306_
	);
	LUT2 #(
		.INIT('h2)
	) name231 (
		_w156_,
		_w306_,
		_w307_
	);
	LUT2 #(
		.INIT('h1)
	) name232 (
		_w304_,
		_w307_,
		_w308_
	);
	LUT2 #(
		.INIT('h1)
	) name233 (
		\musel4_pad ,
		_w308_,
		_w309_
	);
	LUT2 #(
		.INIT('h2)
	) name234 (
		_w300_,
		_w309_,
		_w310_
	);
	LUT2 #(
		.INIT('h8)
	) name235 (
		\inC3_pad ,
		_w79_,
		_w311_
	);
	LUT2 #(
		.INIT('h8)
	) name236 (
		\inA3_pad ,
		_w83_,
		_w312_
	);
	LUT2 #(
		.INIT('h8)
	) name237 (
		\inC3_pad ,
		\musel2_pad ,
		_w313_
	);
	LUT2 #(
		.INIT('h8)
	) name238 (
		\musel1_pad ,
		_w313_,
		_w314_
	);
	LUT2 #(
		.INIT('h1)
	) name239 (
		_w312_,
		_w314_,
		_w315_
	);
	LUT2 #(
		.INIT('h2)
	) name240 (
		_w81_,
		_w315_,
		_w316_
	);
	LUT2 #(
		.INIT('h1)
	) name241 (
		_w311_,
		_w316_,
		_w317_
	);
	LUT2 #(
		.INIT('h1)
	) name242 (
		_w255_,
		_w317_,
		_w318_
	);
	LUT2 #(
		.INIT('h8)
	) name243 (
		_w255_,
		_w317_,
		_w319_
	);
	LUT2 #(
		.INIT('h1)
	) name244 (
		_w318_,
		_w319_,
		_w320_
	);
	LUT2 #(
		.INIT('h8)
	) name245 (
		\inD3_pad ,
		_w150_,
		_w321_
	);
	LUT2 #(
		.INIT('h8)
	) name246 (
		\inB3_pad ,
		_w152_,
		_w322_
	);
	LUT2 #(
		.INIT('h1)
	) name247 (
		_w321_,
		_w322_,
		_w323_
	);
	LUT2 #(
		.INIT('h1)
	) name248 (
		\musel1_pad ,
		_w323_,
		_w324_
	);
	LUT2 #(
		.INIT('h2)
	) name249 (
		\inA3_pad ,
		\musel2_pad ,
		_w325_
	);
	LUT2 #(
		.INIT('h1)
	) name250 (
		_w313_,
		_w325_,
		_w326_
	);
	LUT2 #(
		.INIT('h2)
	) name251 (
		_w156_,
		_w326_,
		_w327_
	);
	LUT2 #(
		.INIT('h1)
	) name252 (
		_w324_,
		_w327_,
		_w328_
	);
	LUT2 #(
		.INIT('h1)
	) name253 (
		\musel4_pad ,
		_w328_,
		_w329_
	);
	LUT2 #(
		.INIT('h4)
	) name254 (
		_w320_,
		_w329_,
		_w330_
	);
	LUT2 #(
		.INIT('h8)
	) name255 (
		\inC2_pad ,
		_w79_,
		_w331_
	);
	LUT2 #(
		.INIT('h8)
	) name256 (
		\inA2_pad ,
		_w83_,
		_w332_
	);
	LUT2 #(
		.INIT('h8)
	) name257 (
		\inC2_pad ,
		\musel2_pad ,
		_w333_
	);
	LUT2 #(
		.INIT('h8)
	) name258 (
		\musel1_pad ,
		_w333_,
		_w334_
	);
	LUT2 #(
		.INIT('h1)
	) name259 (
		_w332_,
		_w334_,
		_w335_
	);
	LUT2 #(
		.INIT('h2)
	) name260 (
		_w81_,
		_w335_,
		_w336_
	);
	LUT2 #(
		.INIT('h1)
	) name261 (
		_w331_,
		_w336_,
		_w337_
	);
	LUT2 #(
		.INIT('h1)
	) name262 (
		_w255_,
		_w337_,
		_w338_
	);
	LUT2 #(
		.INIT('h8)
	) name263 (
		_w255_,
		_w337_,
		_w339_
	);
	LUT2 #(
		.INIT('h1)
	) name264 (
		_w338_,
		_w339_,
		_w340_
	);
	LUT2 #(
		.INIT('h8)
	) name265 (
		\inD2_pad ,
		_w150_,
		_w341_
	);
	LUT2 #(
		.INIT('h8)
	) name266 (
		\inB2_pad ,
		_w152_,
		_w342_
	);
	LUT2 #(
		.INIT('h1)
	) name267 (
		_w341_,
		_w342_,
		_w343_
	);
	LUT2 #(
		.INIT('h1)
	) name268 (
		\musel1_pad ,
		_w343_,
		_w344_
	);
	LUT2 #(
		.INIT('h2)
	) name269 (
		\inA2_pad ,
		\musel2_pad ,
		_w345_
	);
	LUT2 #(
		.INIT('h1)
	) name270 (
		_w333_,
		_w345_,
		_w346_
	);
	LUT2 #(
		.INIT('h2)
	) name271 (
		_w156_,
		_w346_,
		_w347_
	);
	LUT2 #(
		.INIT('h1)
	) name272 (
		_w344_,
		_w347_,
		_w348_
	);
	LUT2 #(
		.INIT('h1)
	) name273 (
		\musel4_pad ,
		_w348_,
		_w349_
	);
	LUT2 #(
		.INIT('h2)
	) name274 (
		_w340_,
		_w349_,
		_w350_
	);
	LUT2 #(
		.INIT('h2)
	) name275 (
		_w320_,
		_w329_,
		_w351_
	);
	LUT2 #(
		.INIT('h1)
	) name276 (
		_w350_,
		_w351_,
		_w352_
	);
	LUT2 #(
		.INIT('h8)
	) name277 (
		\inC1_pad ,
		_w79_,
		_w353_
	);
	LUT2 #(
		.INIT('h8)
	) name278 (
		\inA1_pad ,
		_w83_,
		_w354_
	);
	LUT2 #(
		.INIT('h8)
	) name279 (
		\inC1_pad ,
		\musel2_pad ,
		_w355_
	);
	LUT2 #(
		.INIT('h8)
	) name280 (
		\musel1_pad ,
		_w355_,
		_w356_
	);
	LUT2 #(
		.INIT('h1)
	) name281 (
		_w354_,
		_w356_,
		_w357_
	);
	LUT2 #(
		.INIT('h2)
	) name282 (
		_w81_,
		_w357_,
		_w358_
	);
	LUT2 #(
		.INIT('h1)
	) name283 (
		_w353_,
		_w358_,
		_w359_
	);
	LUT2 #(
		.INIT('h1)
	) name284 (
		_w255_,
		_w359_,
		_w360_
	);
	LUT2 #(
		.INIT('h8)
	) name285 (
		_w255_,
		_w359_,
		_w361_
	);
	LUT2 #(
		.INIT('h1)
	) name286 (
		_w360_,
		_w361_,
		_w362_
	);
	LUT2 #(
		.INIT('h8)
	) name287 (
		\inD1_pad ,
		_w150_,
		_w363_
	);
	LUT2 #(
		.INIT('h8)
	) name288 (
		\inB1_pad ,
		_w152_,
		_w364_
	);
	LUT2 #(
		.INIT('h1)
	) name289 (
		_w363_,
		_w364_,
		_w365_
	);
	LUT2 #(
		.INIT('h1)
	) name290 (
		\musel1_pad ,
		_w365_,
		_w366_
	);
	LUT2 #(
		.INIT('h2)
	) name291 (
		\inA1_pad ,
		\musel2_pad ,
		_w367_
	);
	LUT2 #(
		.INIT('h1)
	) name292 (
		_w355_,
		_w367_,
		_w368_
	);
	LUT2 #(
		.INIT('h2)
	) name293 (
		_w156_,
		_w368_,
		_w369_
	);
	LUT2 #(
		.INIT('h1)
	) name294 (
		_w366_,
		_w369_,
		_w370_
	);
	LUT2 #(
		.INIT('h1)
	) name295 (
		\musel4_pad ,
		_w370_,
		_w371_
	);
	LUT2 #(
		.INIT('h2)
	) name296 (
		_w362_,
		_w371_,
		_w372_
	);
	LUT2 #(
		.INIT('h4)
	) name297 (
		_w169_,
		_w255_,
		_w373_
	);
	LUT2 #(
		.INIT('h4)
	) name298 (
		_w372_,
		_w373_,
		_w374_
	);
	LUT2 #(
		.INIT('h8)
	) name299 (
		_w352_,
		_w374_,
		_w375_
	);
	LUT2 #(
		.INIT('h4)
	) name300 (
		_w340_,
		_w349_,
		_w376_
	);
	LUT2 #(
		.INIT('h4)
	) name301 (
		_w362_,
		_w371_,
		_w377_
	);
	LUT2 #(
		.INIT('h4)
	) name302 (
		_w168_,
		_w255_,
		_w378_
	);
	LUT2 #(
		.INIT('h2)
	) name303 (
		_w168_,
		_w255_,
		_w379_
	);
	LUT2 #(
		.INIT('h2)
	) name304 (
		_w162_,
		_w378_,
		_w380_
	);
	LUT2 #(
		.INIT('h4)
	) name305 (
		_w379_,
		_w380_,
		_w381_
	);
	LUT2 #(
		.INIT('h1)
	) name306 (
		_w376_,
		_w377_,
		_w382_
	);
	LUT2 #(
		.INIT('h4)
	) name307 (
		_w381_,
		_w382_,
		_w383_
	);
	LUT2 #(
		.INIT('h2)
	) name308 (
		_w352_,
		_w383_,
		_w384_
	);
	LUT2 #(
		.INIT('h1)
	) name309 (
		_w330_,
		_w375_,
		_w385_
	);
	LUT2 #(
		.INIT('h4)
	) name310 (
		_w384_,
		_w385_,
		_w386_
	);
	LUT2 #(
		.INIT('h1)
	) name311 (
		_w310_,
		_w386_,
		_w387_
	);
	LUT2 #(
		.INIT('h8)
	) name312 (
		\inC6_pad ,
		_w79_,
		_w388_
	);
	LUT2 #(
		.INIT('h4)
	) name313 (
		\inA6_pad ,
		_w83_,
		_w389_
	);
	LUT2 #(
		.INIT('h8)
	) name314 (
		\inC6_pad ,
		\musel2_pad ,
		_w390_
	);
	LUT2 #(
		.INIT('h1)
	) name315 (
		_w83_,
		_w390_,
		_w391_
	);
	LUT2 #(
		.INIT('h2)
	) name316 (
		_w81_,
		_w389_,
		_w392_
	);
	LUT2 #(
		.INIT('h4)
	) name317 (
		_w391_,
		_w392_,
		_w393_
	);
	LUT2 #(
		.INIT('h1)
	) name318 (
		_w388_,
		_w393_,
		_w394_
	);
	LUT2 #(
		.INIT('h1)
	) name319 (
		_w255_,
		_w394_,
		_w395_
	);
	LUT2 #(
		.INIT('h8)
	) name320 (
		_w255_,
		_w394_,
		_w396_
	);
	LUT2 #(
		.INIT('h1)
	) name321 (
		_w395_,
		_w396_,
		_w397_
	);
	LUT2 #(
		.INIT('h8)
	) name322 (
		\inD6_pad ,
		_w150_,
		_w398_
	);
	LUT2 #(
		.INIT('h8)
	) name323 (
		\inB6_pad ,
		_w152_,
		_w399_
	);
	LUT2 #(
		.INIT('h1)
	) name324 (
		_w398_,
		_w399_,
		_w400_
	);
	LUT2 #(
		.INIT('h1)
	) name325 (
		\musel1_pad ,
		_w400_,
		_w401_
	);
	LUT2 #(
		.INIT('h2)
	) name326 (
		\inA6_pad ,
		\musel2_pad ,
		_w402_
	);
	LUT2 #(
		.INIT('h1)
	) name327 (
		_w390_,
		_w402_,
		_w403_
	);
	LUT2 #(
		.INIT('h2)
	) name328 (
		_w156_,
		_w403_,
		_w404_
	);
	LUT2 #(
		.INIT('h1)
	) name329 (
		_w401_,
		_w404_,
		_w405_
	);
	LUT2 #(
		.INIT('h1)
	) name330 (
		\musel4_pad ,
		_w405_,
		_w406_
	);
	LUT2 #(
		.INIT('h2)
	) name331 (
		_w397_,
		_w406_,
		_w407_
	);
	LUT2 #(
		.INIT('h8)
	) name332 (
		\inC7_pad ,
		_w79_,
		_w408_
	);
	LUT2 #(
		.INIT('h4)
	) name333 (
		\inA7_pad ,
		_w83_,
		_w409_
	);
	LUT2 #(
		.INIT('h8)
	) name334 (
		\inC7_pad ,
		\musel2_pad ,
		_w410_
	);
	LUT2 #(
		.INIT('h1)
	) name335 (
		_w83_,
		_w410_,
		_w411_
	);
	LUT2 #(
		.INIT('h2)
	) name336 (
		_w81_,
		_w409_,
		_w412_
	);
	LUT2 #(
		.INIT('h4)
	) name337 (
		_w411_,
		_w412_,
		_w413_
	);
	LUT2 #(
		.INIT('h1)
	) name338 (
		_w408_,
		_w413_,
		_w414_
	);
	LUT2 #(
		.INIT('h1)
	) name339 (
		_w255_,
		_w414_,
		_w415_
	);
	LUT2 #(
		.INIT('h8)
	) name340 (
		_w255_,
		_w414_,
		_w416_
	);
	LUT2 #(
		.INIT('h1)
	) name341 (
		_w415_,
		_w416_,
		_w417_
	);
	LUT2 #(
		.INIT('h8)
	) name342 (
		\inD7_pad ,
		_w150_,
		_w418_
	);
	LUT2 #(
		.INIT('h8)
	) name343 (
		\inB7_pad ,
		_w152_,
		_w419_
	);
	LUT2 #(
		.INIT('h1)
	) name344 (
		_w418_,
		_w419_,
		_w420_
	);
	LUT2 #(
		.INIT('h1)
	) name345 (
		\musel1_pad ,
		_w420_,
		_w421_
	);
	LUT2 #(
		.INIT('h2)
	) name346 (
		\inA7_pad ,
		\musel2_pad ,
		_w422_
	);
	LUT2 #(
		.INIT('h1)
	) name347 (
		_w410_,
		_w422_,
		_w423_
	);
	LUT2 #(
		.INIT('h2)
	) name348 (
		_w156_,
		_w423_,
		_w424_
	);
	LUT2 #(
		.INIT('h1)
	) name349 (
		_w421_,
		_w424_,
		_w425_
	);
	LUT2 #(
		.INIT('h1)
	) name350 (
		\musel4_pad ,
		_w425_,
		_w426_
	);
	LUT2 #(
		.INIT('h2)
	) name351 (
		_w417_,
		_w426_,
		_w427_
	);
	LUT2 #(
		.INIT('h1)
	) name352 (
		_w407_,
		_w427_,
		_w428_
	);
	LUT2 #(
		.INIT('h8)
	) name353 (
		\inC5_pad ,
		_w79_,
		_w429_
	);
	LUT2 #(
		.INIT('h4)
	) name354 (
		\inA5_pad ,
		_w83_,
		_w430_
	);
	LUT2 #(
		.INIT('h8)
	) name355 (
		\inC5_pad ,
		\musel2_pad ,
		_w431_
	);
	LUT2 #(
		.INIT('h1)
	) name356 (
		_w83_,
		_w431_,
		_w432_
	);
	LUT2 #(
		.INIT('h2)
	) name357 (
		_w81_,
		_w430_,
		_w433_
	);
	LUT2 #(
		.INIT('h4)
	) name358 (
		_w432_,
		_w433_,
		_w434_
	);
	LUT2 #(
		.INIT('h1)
	) name359 (
		_w429_,
		_w434_,
		_w435_
	);
	LUT2 #(
		.INIT('h1)
	) name360 (
		_w255_,
		_w435_,
		_w436_
	);
	LUT2 #(
		.INIT('h8)
	) name361 (
		_w255_,
		_w435_,
		_w437_
	);
	LUT2 #(
		.INIT('h1)
	) name362 (
		_w436_,
		_w437_,
		_w438_
	);
	LUT2 #(
		.INIT('h8)
	) name363 (
		\inD5_pad ,
		_w150_,
		_w439_
	);
	LUT2 #(
		.INIT('h8)
	) name364 (
		\inB5_pad ,
		_w152_,
		_w440_
	);
	LUT2 #(
		.INIT('h1)
	) name365 (
		_w439_,
		_w440_,
		_w441_
	);
	LUT2 #(
		.INIT('h1)
	) name366 (
		\musel1_pad ,
		_w441_,
		_w442_
	);
	LUT2 #(
		.INIT('h2)
	) name367 (
		\inA5_pad ,
		\musel2_pad ,
		_w443_
	);
	LUT2 #(
		.INIT('h1)
	) name368 (
		_w431_,
		_w443_,
		_w444_
	);
	LUT2 #(
		.INIT('h2)
	) name369 (
		_w156_,
		_w444_,
		_w445_
	);
	LUT2 #(
		.INIT('h1)
	) name370 (
		_w442_,
		_w445_,
		_w446_
	);
	LUT2 #(
		.INIT('h1)
	) name371 (
		\musel4_pad ,
		_w446_,
		_w447_
	);
	LUT2 #(
		.INIT('h2)
	) name372 (
		_w438_,
		_w447_,
		_w448_
	);
	LUT2 #(
		.INIT('h2)
	) name373 (
		_w428_,
		_w448_,
		_w449_
	);
	LUT2 #(
		.INIT('h8)
	) name374 (
		_w387_,
		_w449_,
		_w450_
	);
	LUT2 #(
		.INIT('h4)
	) name375 (
		_w417_,
		_w426_,
		_w451_
	);
	LUT2 #(
		.INIT('h4)
	) name376 (
		_w300_,
		_w309_,
		_w452_
	);
	LUT2 #(
		.INIT('h4)
	) name377 (
		_w448_,
		_w452_,
		_w453_
	);
	LUT2 #(
		.INIT('h4)
	) name378 (
		_w438_,
		_w447_,
		_w454_
	);
	LUT2 #(
		.INIT('h4)
	) name379 (
		_w397_,
		_w406_,
		_w455_
	);
	LUT2 #(
		.INIT('h1)
	) name380 (
		_w454_,
		_w455_,
		_w456_
	);
	LUT2 #(
		.INIT('h4)
	) name381 (
		_w453_,
		_w456_,
		_w457_
	);
	LUT2 #(
		.INIT('h2)
	) name382 (
		_w428_,
		_w457_,
		_w458_
	);
	LUT2 #(
		.INIT('h1)
	) name383 (
		_w451_,
		_w458_,
		_w459_
	);
	LUT2 #(
		.INIT('h4)
	) name384 (
		_w450_,
		_w459_,
		_w460_
	);
	LUT2 #(
		.INIT('h4)
	) name385 (
		_w290_,
		_w460_,
		_w461_
	);
	LUT2 #(
		.INIT('h1)
	) name386 (
		_w289_,
		_w461_,
		_w462_
	);
	LUT2 #(
		.INIT('h1)
	) name387 (
		_w269_,
		_w462_,
		_w463_
	);
	LUT2 #(
		.INIT('h1)
	) name388 (
		_w268_,
		_w463_,
		_w464_
	);
	LUT2 #(
		.INIT('h8)
	) name389 (
		\inC10_pad ,
		_w79_,
		_w465_
	);
	LUT2 #(
		.INIT('h8)
	) name390 (
		\inA10_pad ,
		_w83_,
		_w466_
	);
	LUT2 #(
		.INIT('h8)
	) name391 (
		\inC10_pad ,
		\musel2_pad ,
		_w467_
	);
	LUT2 #(
		.INIT('h8)
	) name392 (
		\musel1_pad ,
		_w467_,
		_w468_
	);
	LUT2 #(
		.INIT('h1)
	) name393 (
		_w466_,
		_w468_,
		_w469_
	);
	LUT2 #(
		.INIT('h2)
	) name394 (
		_w81_,
		_w469_,
		_w470_
	);
	LUT2 #(
		.INIT('h1)
	) name395 (
		_w465_,
		_w470_,
		_w471_
	);
	LUT2 #(
		.INIT('h1)
	) name396 (
		_w255_,
		_w471_,
		_w472_
	);
	LUT2 #(
		.INIT('h8)
	) name397 (
		_w255_,
		_w471_,
		_w473_
	);
	LUT2 #(
		.INIT('h1)
	) name398 (
		_w472_,
		_w473_,
		_w474_
	);
	LUT2 #(
		.INIT('h8)
	) name399 (
		\inD10_pad ,
		_w150_,
		_w475_
	);
	LUT2 #(
		.INIT('h8)
	) name400 (
		\inB10_pad ,
		_w152_,
		_w476_
	);
	LUT2 #(
		.INIT('h1)
	) name401 (
		_w475_,
		_w476_,
		_w477_
	);
	LUT2 #(
		.INIT('h1)
	) name402 (
		\musel1_pad ,
		_w477_,
		_w478_
	);
	LUT2 #(
		.INIT('h2)
	) name403 (
		\inA10_pad ,
		\musel2_pad ,
		_w479_
	);
	LUT2 #(
		.INIT('h1)
	) name404 (
		_w467_,
		_w479_,
		_w480_
	);
	LUT2 #(
		.INIT('h2)
	) name405 (
		_w156_,
		_w480_,
		_w481_
	);
	LUT2 #(
		.INIT('h1)
	) name406 (
		_w478_,
		_w481_,
		_w482_
	);
	LUT2 #(
		.INIT('h1)
	) name407 (
		\musel4_pad ,
		_w482_,
		_w483_
	);
	LUT2 #(
		.INIT('h4)
	) name408 (
		_w474_,
		_w483_,
		_w484_
	);
	LUT2 #(
		.INIT('h2)
	) name409 (
		_w474_,
		_w483_,
		_w485_
	);
	LUT2 #(
		.INIT('h1)
	) name410 (
		_w484_,
		_w485_,
		_w486_
	);
	LUT2 #(
		.INIT('h1)
	) name411 (
		_w464_,
		_w486_,
		_w487_
	);
	LUT2 #(
		.INIT('h2)
	) name412 (
		_w464_,
		_w485_,
		_w488_
	);
	LUT2 #(
		.INIT('h4)
	) name413 (
		_w484_,
		_w488_,
		_w489_
	);
	LUT2 #(
		.INIT('h2)
	) name414 (
		_w149_,
		_w487_,
		_w490_
	);
	LUT2 #(
		.INIT('h4)
	) name415 (
		_w489_,
		_w490_,
		_w491_
	);
	LUT2 #(
		.INIT('h1)
	) name416 (
		_w243_,
		_w491_,
		_w492_
	);
	LUT2 #(
		.INIT('h2)
	) name417 (
		_w76_,
		_w492_,
		_w493_
	);
	LUT2 #(
		.INIT('h2)
	) name418 (
		\inA15_pad ,
		\musel2_pad ,
		_w494_
	);
	LUT2 #(
		.INIT('h2)
	) name419 (
		\inC15_pad ,
		\musel1_pad ,
		_w495_
	);
	LUT2 #(
		.INIT('h1)
	) name420 (
		_w494_,
		_w495_,
		_w496_
	);
	LUT2 #(
		.INIT('h4)
	) name421 (
		_w78_,
		_w496_,
		_w497_
	);
	LUT2 #(
		.INIT('h2)
	) name422 (
		\inC10_pad ,
		\musel1_pad ,
		_w498_
	);
	LUT2 #(
		.INIT('h1)
	) name423 (
		_w479_,
		_w498_,
		_w499_
	);
	LUT2 #(
		.INIT('h2)
	) name424 (
		_w497_,
		_w499_,
		_w500_
	);
	LUT2 #(
		.INIT('h1)
	) name425 (
		_w78_,
		_w496_,
		_w501_
	);
	LUT2 #(
		.INIT('h8)
	) name426 (
		_w499_,
		_w501_,
		_w502_
	);
	LUT2 #(
		.INIT('h1)
	) name427 (
		_w500_,
		_w502_,
		_w503_
	);
	LUT2 #(
		.INIT('h2)
	) name428 (
		\inC9_pad ,
		\musel1_pad ,
		_w504_
	);
	LUT2 #(
		.INIT('h1)
	) name429 (
		_w263_,
		_w504_,
		_w505_
	);
	LUT2 #(
		.INIT('h2)
	) name430 (
		_w497_,
		_w505_,
		_w506_
	);
	LUT2 #(
		.INIT('h8)
	) name431 (
		_w501_,
		_w505_,
		_w507_
	);
	LUT2 #(
		.INIT('h1)
	) name432 (
		_w506_,
		_w507_,
		_w508_
	);
	LUT2 #(
		.INIT('h2)
	) name433 (
		\inC8_pad ,
		\musel1_pad ,
		_w509_
	);
	LUT2 #(
		.INIT('h1)
	) name434 (
		_w284_,
		_w509_,
		_w510_
	);
	LUT2 #(
		.INIT('h2)
	) name435 (
		_w497_,
		_w510_,
		_w511_
	);
	LUT2 #(
		.INIT('h8)
	) name436 (
		_w501_,
		_w510_,
		_w512_
	);
	LUT2 #(
		.INIT('h1)
	) name437 (
		_w511_,
		_w512_,
		_w513_
	);
	LUT2 #(
		.INIT('h2)
	) name438 (
		\inC2_pad ,
		\musel1_pad ,
		_w514_
	);
	LUT2 #(
		.INIT('h1)
	) name439 (
		_w345_,
		_w514_,
		_w515_
	);
	LUT2 #(
		.INIT('h1)
	) name440 (
		_w496_,
		_w515_,
		_w516_
	);
	LUT2 #(
		.INIT('h8)
	) name441 (
		_w496_,
		_w515_,
		_w517_
	);
	LUT2 #(
		.INIT('h2)
	) name442 (
		_w178_,
		_w516_,
		_w518_
	);
	LUT2 #(
		.INIT('h4)
	) name443 (
		_w517_,
		_w518_,
		_w519_
	);
	LUT2 #(
		.INIT('h2)
	) name444 (
		\inC3_pad ,
		\musel1_pad ,
		_w520_
	);
	LUT2 #(
		.INIT('h1)
	) name445 (
		_w325_,
		_w520_,
		_w521_
	);
	LUT2 #(
		.INIT('h2)
	) name446 (
		_w497_,
		_w521_,
		_w522_
	);
	LUT2 #(
		.INIT('h8)
	) name447 (
		_w501_,
		_w521_,
		_w523_
	);
	LUT2 #(
		.INIT('h1)
	) name448 (
		_w522_,
		_w523_,
		_w524_
	);
	LUT2 #(
		.INIT('h2)
	) name449 (
		_w178_,
		_w496_,
		_w525_
	);
	LUT2 #(
		.INIT('h8)
	) name450 (
		_w177_,
		_w525_,
		_w526_
	);
	LUT2 #(
		.INIT('h2)
	) name451 (
		_w179_,
		_w521_,
		_w527_
	);
	LUT2 #(
		.INIT('h1)
	) name452 (
		_w526_,
		_w527_,
		_w528_
	);
	LUT2 #(
		.INIT('h2)
	) name453 (
		\inC1_pad ,
		\musel1_pad ,
		_w529_
	);
	LUT2 #(
		.INIT('h1)
	) name454 (
		_w367_,
		_w529_,
		_w530_
	);
	LUT2 #(
		.INIT('h8)
	) name455 (
		_w501_,
		_w530_,
		_w531_
	);
	LUT2 #(
		.INIT('h2)
	) name456 (
		_w497_,
		_w530_,
		_w532_
	);
	LUT2 #(
		.INIT('h1)
	) name457 (
		_w531_,
		_w532_,
		_w533_
	);
	LUT2 #(
		.INIT('h2)
	) name458 (
		_w519_,
		_w524_,
		_w534_
	);
	LUT2 #(
		.INIT('h1)
	) name459 (
		_w528_,
		_w533_,
		_w535_
	);
	LUT2 #(
		.INIT('h8)
	) name460 (
		_w534_,
		_w535_,
		_w536_
	);
	LUT2 #(
		.INIT('h2)
	) name461 (
		\inA11_pad ,
		\musel2_pad ,
		_w537_
	);
	LUT2 #(
		.INIT('h2)
	) name462 (
		\inC11_pad ,
		\musel1_pad ,
		_w538_
	);
	LUT2 #(
		.INIT('h1)
	) name463 (
		_w537_,
		_w538_,
		_w539_
	);
	LUT2 #(
		.INIT('h8)
	) name464 (
		_w496_,
		_w539_,
		_w540_
	);
	LUT2 #(
		.INIT('h2)
	) name465 (
		_w501_,
		_w539_,
		_w541_
	);
	LUT2 #(
		.INIT('h2)
	) name466 (
		_w178_,
		_w540_,
		_w542_
	);
	LUT2 #(
		.INIT('h4)
	) name467 (
		_w541_,
		_w542_,
		_w543_
	);
	LUT2 #(
		.INIT('h1)
	) name468 (
		_w503_,
		_w508_,
		_w544_
	);
	LUT2 #(
		.INIT('h4)
	) name469 (
		_w513_,
		_w543_,
		_w545_
	);
	LUT2 #(
		.INIT('h8)
	) name470 (
		_w544_,
		_w545_,
		_w546_
	);
	LUT2 #(
		.INIT('h8)
	) name471 (
		_w536_,
		_w546_,
		_w547_
	);
	LUT2 #(
		.INIT('h8)
	) name472 (
		_w501_,
		_w547_,
		_w548_
	);
	LUT2 #(
		.INIT('h2)
	) name473 (
		_w77_,
		_w548_,
		_w549_
	);
	LUT2 #(
		.INIT('h4)
	) name474 (
		_w503_,
		_w549_,
		_w550_
	);
	LUT2 #(
		.INIT('h1)
	) name475 (
		_w175_,
		_w550_,
		_w551_
	);
	LUT2 #(
		.INIT('h8)
	) name476 (
		_w175_,
		_w242_,
		_w552_
	);
	LUT2 #(
		.INIT('h2)
	) name477 (
		_w183_,
		_w551_,
		_w553_
	);
	LUT2 #(
		.INIT('h4)
	) name478 (
		_w552_,
		_w553_,
		_w554_
	);
	LUT2 #(
		.INIT('h1)
	) name479 (
		_w493_,
		_w554_,
		_w555_
	);
	LUT2 #(
		.INIT('h8)
	) name480 (
		\sh0_pad ,
		\sh1_pad ,
		_w556_
	);
	LUT2 #(
		.INIT('h2)
	) name481 (
		_w215_,
		_w556_,
		_w557_
	);
	LUT2 #(
		.INIT('h8)
	) name482 (
		_w236_,
		_w556_,
		_w558_
	);
	LUT2 #(
		.INIT('h1)
	) name483 (
		_w557_,
		_w558_,
		_w559_
	);
	LUT2 #(
		.INIT('h2)
	) name484 (
		\sh2_pad ,
		_w559_,
		_w560_
	);
	LUT2 #(
		.INIT('h2)
	) name485 (
		\sh1_pad ,
		_w192_,
		_w561_
	);
	LUT2 #(
		.INIT('h1)
	) name486 (
		\sh1_pad ,
		_w208_,
		_w562_
	);
	LUT2 #(
		.INIT('h1)
	) name487 (
		_w561_,
		_w562_,
		_w563_
	);
	LUT2 #(
		.INIT('h2)
	) name488 (
		\sh0_pad ,
		_w563_,
		_w564_
	);
	LUT2 #(
		.INIT('h1)
	) name489 (
		\sh1_pad ,
		_w236_,
		_w565_
	);
	LUT2 #(
		.INIT('h2)
	) name490 (
		\sh1_pad ,
		_w227_,
		_w566_
	);
	LUT2 #(
		.INIT('h1)
	) name491 (
		_w565_,
		_w566_,
		_w567_
	);
	LUT2 #(
		.INIT('h1)
	) name492 (
		\sh0_pad ,
		_w567_,
		_w568_
	);
	LUT2 #(
		.INIT('h1)
	) name493 (
		\sh2_pad ,
		_w564_,
		_w569_
	);
	LUT2 #(
		.INIT('h4)
	) name494 (
		_w568_,
		_w569_,
		_w570_
	);
	LUT2 #(
		.INIT('h1)
	) name495 (
		_w560_,
		_w570_,
		_w571_
	);
	LUT2 #(
		.INIT('h8)
	) name496 (
		_w146_,
		_w571_,
		_w572_
	);
	LUT2 #(
		.INIT('h8)
	) name497 (
		\inC11_pad ,
		_w79_,
		_w573_
	);
	LUT2 #(
		.INIT('h8)
	) name498 (
		\inA11_pad ,
		_w83_,
		_w574_
	);
	LUT2 #(
		.INIT('h8)
	) name499 (
		\inC11_pad ,
		\musel2_pad ,
		_w575_
	);
	LUT2 #(
		.INIT('h8)
	) name500 (
		\musel1_pad ,
		_w575_,
		_w576_
	);
	LUT2 #(
		.INIT('h1)
	) name501 (
		_w574_,
		_w576_,
		_w577_
	);
	LUT2 #(
		.INIT('h2)
	) name502 (
		_w81_,
		_w577_,
		_w578_
	);
	LUT2 #(
		.INIT('h1)
	) name503 (
		_w573_,
		_w578_,
		_w579_
	);
	LUT2 #(
		.INIT('h1)
	) name504 (
		_w255_,
		_w579_,
		_w580_
	);
	LUT2 #(
		.INIT('h8)
	) name505 (
		_w255_,
		_w579_,
		_w581_
	);
	LUT2 #(
		.INIT('h1)
	) name506 (
		_w580_,
		_w581_,
		_w582_
	);
	LUT2 #(
		.INIT('h8)
	) name507 (
		\inD11_pad ,
		_w150_,
		_w583_
	);
	LUT2 #(
		.INIT('h8)
	) name508 (
		\inB11_pad ,
		_w152_,
		_w584_
	);
	LUT2 #(
		.INIT('h1)
	) name509 (
		_w583_,
		_w584_,
		_w585_
	);
	LUT2 #(
		.INIT('h1)
	) name510 (
		\musel1_pad ,
		_w585_,
		_w586_
	);
	LUT2 #(
		.INIT('h1)
	) name511 (
		_w537_,
		_w575_,
		_w587_
	);
	LUT2 #(
		.INIT('h2)
	) name512 (
		_w156_,
		_w587_,
		_w588_
	);
	LUT2 #(
		.INIT('h1)
	) name513 (
		_w586_,
		_w588_,
		_w589_
	);
	LUT2 #(
		.INIT('h1)
	) name514 (
		\musel4_pad ,
		_w589_,
		_w590_
	);
	LUT2 #(
		.INIT('h2)
	) name515 (
		_w582_,
		_w590_,
		_w591_
	);
	LUT2 #(
		.INIT('h4)
	) name516 (
		_w582_,
		_w590_,
		_w592_
	);
	LUT2 #(
		.INIT('h1)
	) name517 (
		_w591_,
		_w592_,
		_w593_
	);
	LUT2 #(
		.INIT('h8)
	) name518 (
		_w488_,
		_w593_,
		_w594_
	);
	LUT2 #(
		.INIT('h1)
	) name519 (
		_w484_,
		_w593_,
		_w595_
	);
	LUT2 #(
		.INIT('h4)
	) name520 (
		_w488_,
		_w595_,
		_w596_
	);
	LUT2 #(
		.INIT('h2)
	) name521 (
		_w149_,
		_w594_,
		_w597_
	);
	LUT2 #(
		.INIT('h4)
	) name522 (
		_w596_,
		_w597_,
		_w598_
	);
	LUT2 #(
		.INIT('h1)
	) name523 (
		_w572_,
		_w598_,
		_w599_
	);
	LUT2 #(
		.INIT('h2)
	) name524 (
		_w76_,
		_w599_,
		_w600_
	);
	LUT2 #(
		.INIT('h2)
	) name525 (
		_w543_,
		_w548_,
		_w601_
	);
	LUT2 #(
		.INIT('h1)
	) name526 (
		_w175_,
		_w601_,
		_w602_
	);
	LUT2 #(
		.INIT('h2)
	) name527 (
		_w175_,
		_w571_,
		_w603_
	);
	LUT2 #(
		.INIT('h2)
	) name528 (
		_w183_,
		_w602_,
		_w604_
	);
	LUT2 #(
		.INIT('h4)
	) name529 (
		_w603_,
		_w604_,
		_w605_
	);
	LUT2 #(
		.INIT('h1)
	) name530 (
		_w600_,
		_w605_,
		_w606_
	);
	LUT2 #(
		.INIT('h4)
	) name531 (
		_w215_,
		_w556_,
		_w607_
	);
	LUT2 #(
		.INIT('h1)
	) name532 (
		\sh0_pad ,
		_w563_,
		_w608_
	);
	LUT2 #(
		.INIT('h2)
	) name533 (
		\sh0_pad ,
		\sh1_pad ,
		_w609_
	);
	LUT2 #(
		.INIT('h4)
	) name534 (
		_w227_,
		_w609_,
		_w610_
	);
	LUT2 #(
		.INIT('h1)
	) name535 (
		_w607_,
		_w610_,
		_w611_
	);
	LUT2 #(
		.INIT('h4)
	) name536 (
		_w608_,
		_w611_,
		_w612_
	);
	LUT2 #(
		.INIT('h1)
	) name537 (
		\sh2_pad ,
		_w612_,
		_w613_
	);
	LUT2 #(
		.INIT('h8)
	) name538 (
		_w208_,
		_w556_,
		_w614_
	);
	LUT2 #(
		.INIT('h2)
	) name539 (
		\sh2_pad ,
		_w557_,
		_w615_
	);
	LUT2 #(
		.INIT('h4)
	) name540 (
		_w614_,
		_w615_,
		_w616_
	);
	LUT2 #(
		.INIT('h1)
	) name541 (
		_w613_,
		_w616_,
		_w617_
	);
	LUT2 #(
		.INIT('h2)
	) name542 (
		_w146_,
		_w617_,
		_w618_
	);
	LUT2 #(
		.INIT('h8)
	) name543 (
		\inC12_pad ,
		_w79_,
		_w619_
	);
	LUT2 #(
		.INIT('h8)
	) name544 (
		\inA12_pad ,
		_w83_,
		_w620_
	);
	LUT2 #(
		.INIT('h8)
	) name545 (
		\inC12_pad ,
		\musel2_pad ,
		_w621_
	);
	LUT2 #(
		.INIT('h8)
	) name546 (
		\musel1_pad ,
		_w621_,
		_w622_
	);
	LUT2 #(
		.INIT('h1)
	) name547 (
		_w620_,
		_w622_,
		_w623_
	);
	LUT2 #(
		.INIT('h2)
	) name548 (
		_w81_,
		_w623_,
		_w624_
	);
	LUT2 #(
		.INIT('h1)
	) name549 (
		_w619_,
		_w624_,
		_w625_
	);
	LUT2 #(
		.INIT('h1)
	) name550 (
		_w255_,
		_w625_,
		_w626_
	);
	LUT2 #(
		.INIT('h8)
	) name551 (
		_w255_,
		_w625_,
		_w627_
	);
	LUT2 #(
		.INIT('h1)
	) name552 (
		_w626_,
		_w627_,
		_w628_
	);
	LUT2 #(
		.INIT('h8)
	) name553 (
		\inD12_pad ,
		_w150_,
		_w629_
	);
	LUT2 #(
		.INIT('h8)
	) name554 (
		\inB12_pad ,
		_w152_,
		_w630_
	);
	LUT2 #(
		.INIT('h1)
	) name555 (
		_w629_,
		_w630_,
		_w631_
	);
	LUT2 #(
		.INIT('h1)
	) name556 (
		\musel1_pad ,
		_w631_,
		_w632_
	);
	LUT2 #(
		.INIT('h2)
	) name557 (
		\inA12_pad ,
		\musel2_pad ,
		_w633_
	);
	LUT2 #(
		.INIT('h1)
	) name558 (
		_w621_,
		_w633_,
		_w634_
	);
	LUT2 #(
		.INIT('h2)
	) name559 (
		_w156_,
		_w634_,
		_w635_
	);
	LUT2 #(
		.INIT('h1)
	) name560 (
		_w632_,
		_w635_,
		_w636_
	);
	LUT2 #(
		.INIT('h1)
	) name561 (
		\musel4_pad ,
		_w636_,
		_w637_
	);
	LUT2 #(
		.INIT('h2)
	) name562 (
		_w628_,
		_w637_,
		_w638_
	);
	LUT2 #(
		.INIT('h4)
	) name563 (
		_w628_,
		_w637_,
		_w639_
	);
	LUT2 #(
		.INIT('h1)
	) name564 (
		_w638_,
		_w639_,
		_w640_
	);
	LUT2 #(
		.INIT('h1)
	) name565 (
		_w268_,
		_w289_,
		_w641_
	);
	LUT2 #(
		.INIT('h1)
	) name566 (
		_w485_,
		_w591_,
		_w642_
	);
	LUT2 #(
		.INIT('h8)
	) name567 (
		_w641_,
		_w642_,
		_w643_
	);
	LUT2 #(
		.INIT('h4)
	) name568 (
		_w460_,
		_w643_,
		_w644_
	);
	LUT2 #(
		.INIT('h1)
	) name569 (
		_w640_,
		_w644_,
		_w645_
	);
	LUT2 #(
		.INIT('h8)
	) name570 (
		_w640_,
		_w644_,
		_w646_
	);
	LUT2 #(
		.INIT('h2)
	) name571 (
		_w149_,
		_w645_,
		_w647_
	);
	LUT2 #(
		.INIT('h4)
	) name572 (
		_w646_,
		_w647_,
		_w648_
	);
	LUT2 #(
		.INIT('h1)
	) name573 (
		_w618_,
		_w648_,
		_w649_
	);
	LUT2 #(
		.INIT('h2)
	) name574 (
		_w76_,
		_w649_,
		_w650_
	);
	LUT2 #(
		.INIT('h2)
	) name575 (
		\inC4_pad ,
		\musel1_pad ,
		_w651_
	);
	LUT2 #(
		.INIT('h1)
	) name576 (
		_w305_,
		_w651_,
		_w652_
	);
	LUT2 #(
		.INIT('h2)
	) name577 (
		_w497_,
		_w652_,
		_w653_
	);
	LUT2 #(
		.INIT('h8)
	) name578 (
		_w501_,
		_w652_,
		_w654_
	);
	LUT2 #(
		.INIT('h1)
	) name579 (
		_w653_,
		_w654_,
		_w655_
	);
	LUT2 #(
		.INIT('h2)
	) name580 (
		\inC6_pad ,
		\musel1_pad ,
		_w656_
	);
	LUT2 #(
		.INIT('h1)
	) name581 (
		_w402_,
		_w656_,
		_w657_
	);
	LUT2 #(
		.INIT('h1)
	) name582 (
		_w78_,
		_w657_,
		_w658_
	);
	LUT2 #(
		.INIT('h2)
	) name583 (
		\inC5_pad ,
		\musel1_pad ,
		_w659_
	);
	LUT2 #(
		.INIT('h1)
	) name584 (
		_w443_,
		_w659_,
		_w660_
	);
	LUT2 #(
		.INIT('h8)
	) name585 (
		_w496_,
		_w660_,
		_w661_
	);
	LUT2 #(
		.INIT('h2)
	) name586 (
		_w501_,
		_w660_,
		_w662_
	);
	LUT2 #(
		.INIT('h2)
	) name587 (
		_w178_,
		_w661_,
		_w663_
	);
	LUT2 #(
		.INIT('h4)
	) name588 (
		_w662_,
		_w663_,
		_w664_
	);
	LUT2 #(
		.INIT('h2)
	) name589 (
		\inC7_pad ,
		\musel1_pad ,
		_w665_
	);
	LUT2 #(
		.INIT('h1)
	) name590 (
		_w422_,
		_w665_,
		_w666_
	);
	LUT2 #(
		.INIT('h8)
	) name591 (
		_w525_,
		_w666_,
		_w667_
	);
	LUT2 #(
		.INIT('h4)
	) name592 (
		_w658_,
		_w667_,
		_w668_
	);
	LUT2 #(
		.INIT('h4)
	) name593 (
		_w655_,
		_w668_,
		_w669_
	);
	LUT2 #(
		.INIT('h8)
	) name594 (
		_w664_,
		_w669_,
		_w670_
	);
	LUT2 #(
		.INIT('h8)
	) name595 (
		_w547_,
		_w670_,
		_w671_
	);
	LUT2 #(
		.INIT('h2)
	) name596 (
		\inC12_pad ,
		\musel1_pad ,
		_w672_
	);
	LUT2 #(
		.INIT('h1)
	) name597 (
		_w633_,
		_w672_,
		_w673_
	);
	LUT2 #(
		.INIT('h8)
	) name598 (
		_w496_,
		_w673_,
		_w674_
	);
	LUT2 #(
		.INIT('h2)
	) name599 (
		_w501_,
		_w673_,
		_w675_
	);
	LUT2 #(
		.INIT('h2)
	) name600 (
		_w178_,
		_w674_,
		_w676_
	);
	LUT2 #(
		.INIT('h4)
	) name601 (
		_w675_,
		_w676_,
		_w677_
	);
	LUT2 #(
		.INIT('h8)
	) name602 (
		_w671_,
		_w677_,
		_w678_
	);
	LUT2 #(
		.INIT('h1)
	) name603 (
		_w671_,
		_w677_,
		_w679_
	);
	LUT2 #(
		.INIT('h1)
	) name604 (
		_w678_,
		_w679_,
		_w680_
	);
	LUT2 #(
		.INIT('h1)
	) name605 (
		_w175_,
		_w680_,
		_w681_
	);
	LUT2 #(
		.INIT('h8)
	) name606 (
		_w175_,
		_w617_,
		_w682_
	);
	LUT2 #(
		.INIT('h2)
	) name607 (
		_w183_,
		_w681_,
		_w683_
	);
	LUT2 #(
		.INIT('h4)
	) name608 (
		_w682_,
		_w683_,
		_w684_
	);
	LUT2 #(
		.INIT('h1)
	) name609 (
		_w650_,
		_w684_,
		_w685_
	);
	LUT2 #(
		.INIT('h8)
	) name610 (
		\sh2_pad ,
		_w556_,
		_w686_
	);
	LUT2 #(
		.INIT('h4)
	) name611 (
		_w227_,
		_w686_,
		_w687_
	);
	LUT2 #(
		.INIT('h1)
	) name612 (
		\sh1_pad ,
		\sh2_pad ,
		_w688_
	);
	LUT2 #(
		.INIT('h1)
	) name613 (
		_w686_,
		_w688_,
		_w689_
	);
	LUT2 #(
		.INIT('h4)
	) name614 (
		_w215_,
		_w689_,
		_w690_
	);
	LUT2 #(
		.INIT('h4)
	) name615 (
		\sh0_pad ,
		_w227_,
		_w691_
	);
	LUT2 #(
		.INIT('h8)
	) name616 (
		\sh0_pad ,
		_w192_,
		_w692_
	);
	LUT2 #(
		.INIT('h2)
	) name617 (
		_w688_,
		_w691_,
		_w693_
	);
	LUT2 #(
		.INIT('h4)
	) name618 (
		_w692_,
		_w693_,
		_w694_
	);
	LUT2 #(
		.INIT('h1)
	) name619 (
		_w687_,
		_w690_,
		_w695_
	);
	LUT2 #(
		.INIT('h4)
	) name620 (
		_w694_,
		_w695_,
		_w696_
	);
	LUT2 #(
		.INIT('h2)
	) name621 (
		_w146_,
		_w696_,
		_w697_
	);
	LUT2 #(
		.INIT('h8)
	) name622 (
		\inC13_pad ,
		_w79_,
		_w698_
	);
	LUT2 #(
		.INIT('h8)
	) name623 (
		\inA13_pad ,
		_w83_,
		_w699_
	);
	LUT2 #(
		.INIT('h8)
	) name624 (
		\inC13_pad ,
		\musel2_pad ,
		_w700_
	);
	LUT2 #(
		.INIT('h8)
	) name625 (
		\musel1_pad ,
		_w700_,
		_w701_
	);
	LUT2 #(
		.INIT('h1)
	) name626 (
		_w699_,
		_w701_,
		_w702_
	);
	LUT2 #(
		.INIT('h2)
	) name627 (
		_w81_,
		_w702_,
		_w703_
	);
	LUT2 #(
		.INIT('h1)
	) name628 (
		_w698_,
		_w703_,
		_w704_
	);
	LUT2 #(
		.INIT('h1)
	) name629 (
		_w255_,
		_w704_,
		_w705_
	);
	LUT2 #(
		.INIT('h8)
	) name630 (
		_w255_,
		_w704_,
		_w706_
	);
	LUT2 #(
		.INIT('h1)
	) name631 (
		_w705_,
		_w706_,
		_w707_
	);
	LUT2 #(
		.INIT('h8)
	) name632 (
		\inD13_pad ,
		_w150_,
		_w708_
	);
	LUT2 #(
		.INIT('h8)
	) name633 (
		\inB13_pad ,
		_w152_,
		_w709_
	);
	LUT2 #(
		.INIT('h1)
	) name634 (
		_w708_,
		_w709_,
		_w710_
	);
	LUT2 #(
		.INIT('h1)
	) name635 (
		\musel1_pad ,
		_w710_,
		_w711_
	);
	LUT2 #(
		.INIT('h2)
	) name636 (
		\inA13_pad ,
		\musel2_pad ,
		_w712_
	);
	LUT2 #(
		.INIT('h1)
	) name637 (
		_w700_,
		_w712_,
		_w713_
	);
	LUT2 #(
		.INIT('h2)
	) name638 (
		_w156_,
		_w713_,
		_w714_
	);
	LUT2 #(
		.INIT('h1)
	) name639 (
		_w711_,
		_w714_,
		_w715_
	);
	LUT2 #(
		.INIT('h1)
	) name640 (
		\musel4_pad ,
		_w715_,
		_w716_
	);
	LUT2 #(
		.INIT('h2)
	) name641 (
		_w707_,
		_w716_,
		_w717_
	);
	LUT2 #(
		.INIT('h4)
	) name642 (
		_w707_,
		_w716_,
		_w718_
	);
	LUT2 #(
		.INIT('h1)
	) name643 (
		_w717_,
		_w718_,
		_w719_
	);
	LUT2 #(
		.INIT('h4)
	) name644 (
		_w638_,
		_w644_,
		_w720_
	);
	LUT2 #(
		.INIT('h1)
	) name645 (
		_w639_,
		_w720_,
		_w721_
	);
	LUT2 #(
		.INIT('h4)
	) name646 (
		_w719_,
		_w721_,
		_w722_
	);
	LUT2 #(
		.INIT('h8)
	) name647 (
		_w719_,
		_w720_,
		_w723_
	);
	LUT2 #(
		.INIT('h2)
	) name648 (
		_w149_,
		_w723_,
		_w724_
	);
	LUT2 #(
		.INIT('h4)
	) name649 (
		_w722_,
		_w724_,
		_w725_
	);
	LUT2 #(
		.INIT('h1)
	) name650 (
		_w697_,
		_w725_,
		_w726_
	);
	LUT2 #(
		.INIT('h2)
	) name651 (
		_w76_,
		_w726_,
		_w727_
	);
	LUT2 #(
		.INIT('h8)
	) name652 (
		_w175_,
		_w696_,
		_w728_
	);
	LUT2 #(
		.INIT('h2)
	) name653 (
		\inC13_pad ,
		\musel1_pad ,
		_w729_
	);
	LUT2 #(
		.INIT('h1)
	) name654 (
		_w712_,
		_w729_,
		_w730_
	);
	LUT2 #(
		.INIT('h2)
	) name655 (
		_w497_,
		_w730_,
		_w731_
	);
	LUT2 #(
		.INIT('h8)
	) name656 (
		_w501_,
		_w730_,
		_w732_
	);
	LUT2 #(
		.INIT('h1)
	) name657 (
		_w731_,
		_w732_,
		_w733_
	);
	LUT2 #(
		.INIT('h2)
	) name658 (
		_w77_,
		_w733_,
		_w734_
	);
	LUT2 #(
		.INIT('h1)
	) name659 (
		_w678_,
		_w734_,
		_w735_
	);
	LUT2 #(
		.INIT('h2)
	) name660 (
		_w678_,
		_w733_,
		_w736_
	);
	LUT2 #(
		.INIT('h1)
	) name661 (
		_w735_,
		_w736_,
		_w737_
	);
	LUT2 #(
		.INIT('h1)
	) name662 (
		_w175_,
		_w737_,
		_w738_
	);
	LUT2 #(
		.INIT('h2)
	) name663 (
		_w183_,
		_w728_,
		_w739_
	);
	LUT2 #(
		.INIT('h4)
	) name664 (
		_w738_,
		_w739_,
		_w740_
	);
	LUT2 #(
		.INIT('h1)
	) name665 (
		_w727_,
		_w740_,
		_w741_
	);
	LUT2 #(
		.INIT('h4)
	) name666 (
		_w717_,
		_w720_,
		_w742_
	);
	LUT2 #(
		.INIT('h8)
	) name667 (
		\inC14_pad ,
		_w79_,
		_w743_
	);
	LUT2 #(
		.INIT('h8)
	) name668 (
		\inA14_pad ,
		_w83_,
		_w744_
	);
	LUT2 #(
		.INIT('h8)
	) name669 (
		\inC14_pad ,
		\musel2_pad ,
		_w745_
	);
	LUT2 #(
		.INIT('h8)
	) name670 (
		\musel1_pad ,
		_w745_,
		_w746_
	);
	LUT2 #(
		.INIT('h1)
	) name671 (
		_w744_,
		_w746_,
		_w747_
	);
	LUT2 #(
		.INIT('h2)
	) name672 (
		_w81_,
		_w747_,
		_w748_
	);
	LUT2 #(
		.INIT('h1)
	) name673 (
		_w743_,
		_w748_,
		_w749_
	);
	LUT2 #(
		.INIT('h1)
	) name674 (
		_w255_,
		_w749_,
		_w750_
	);
	LUT2 #(
		.INIT('h8)
	) name675 (
		_w255_,
		_w749_,
		_w751_
	);
	LUT2 #(
		.INIT('h1)
	) name676 (
		_w750_,
		_w751_,
		_w752_
	);
	LUT2 #(
		.INIT('h8)
	) name677 (
		\inD14_pad ,
		_w150_,
		_w753_
	);
	LUT2 #(
		.INIT('h8)
	) name678 (
		\inB14_pad ,
		_w152_,
		_w754_
	);
	LUT2 #(
		.INIT('h1)
	) name679 (
		_w753_,
		_w754_,
		_w755_
	);
	LUT2 #(
		.INIT('h1)
	) name680 (
		\musel1_pad ,
		_w755_,
		_w756_
	);
	LUT2 #(
		.INIT('h2)
	) name681 (
		\inA14_pad ,
		\musel2_pad ,
		_w757_
	);
	LUT2 #(
		.INIT('h1)
	) name682 (
		_w745_,
		_w757_,
		_w758_
	);
	LUT2 #(
		.INIT('h2)
	) name683 (
		_w156_,
		_w758_,
		_w759_
	);
	LUT2 #(
		.INIT('h1)
	) name684 (
		_w756_,
		_w759_,
		_w760_
	);
	LUT2 #(
		.INIT('h1)
	) name685 (
		\musel4_pad ,
		_w760_,
		_w761_
	);
	LUT2 #(
		.INIT('h2)
	) name686 (
		_w752_,
		_w761_,
		_w762_
	);
	LUT2 #(
		.INIT('h4)
	) name687 (
		_w752_,
		_w761_,
		_w763_
	);
	LUT2 #(
		.INIT('h1)
	) name688 (
		_w762_,
		_w763_,
		_w764_
	);
	LUT2 #(
		.INIT('h4)
	) name689 (
		_w718_,
		_w764_,
		_w765_
	);
	LUT2 #(
		.INIT('h4)
	) name690 (
		_w742_,
		_w765_,
		_w766_
	);
	LUT2 #(
		.INIT('h4)
	) name691 (
		_w718_,
		_w721_,
		_w767_
	);
	LUT2 #(
		.INIT('h1)
	) name692 (
		_w717_,
		_w764_,
		_w768_
	);
	LUT2 #(
		.INIT('h4)
	) name693 (
		_w767_,
		_w768_,
		_w769_
	);
	LUT2 #(
		.INIT('h1)
	) name694 (
		_w766_,
		_w769_,
		_w770_
	);
	LUT2 #(
		.INIT('h2)
	) name695 (
		_w149_,
		_w770_,
		_w771_
	);
	LUT2 #(
		.INIT('h8)
	) name696 (
		\sh0_pad ,
		\sh2_pad ,
		_w772_
	);
	LUT2 #(
		.INIT('h1)
	) name697 (
		_w688_,
		_w772_,
		_w773_
	);
	LUT2 #(
		.INIT('h1)
	) name698 (
		_w609_,
		_w773_,
		_w774_
	);
	LUT2 #(
		.INIT('h4)
	) name699 (
		_w192_,
		_w774_,
		_w775_
	);
	LUT2 #(
		.INIT('h1)
	) name700 (
		_w215_,
		_w774_,
		_w776_
	);
	LUT2 #(
		.INIT('h1)
	) name701 (
		_w775_,
		_w776_,
		_w777_
	);
	LUT2 #(
		.INIT('h2)
	) name702 (
		_w146_,
		_w777_,
		_w778_
	);
	LUT2 #(
		.INIT('h1)
	) name703 (
		_w771_,
		_w778_,
		_w779_
	);
	LUT2 #(
		.INIT('h2)
	) name704 (
		_w76_,
		_w779_,
		_w780_
	);
	LUT2 #(
		.INIT('h8)
	) name705 (
		_w175_,
		_w777_,
		_w781_
	);
	LUT2 #(
		.INIT('h2)
	) name706 (
		\inC14_pad ,
		\musel1_pad ,
		_w782_
	);
	LUT2 #(
		.INIT('h1)
	) name707 (
		_w757_,
		_w782_,
		_w783_
	);
	LUT2 #(
		.INIT('h8)
	) name708 (
		_w496_,
		_w783_,
		_w784_
	);
	LUT2 #(
		.INIT('h2)
	) name709 (
		_w501_,
		_w783_,
		_w785_
	);
	LUT2 #(
		.INIT('h2)
	) name710 (
		_w178_,
		_w784_,
		_w786_
	);
	LUT2 #(
		.INIT('h4)
	) name711 (
		_w785_,
		_w786_,
		_w787_
	);
	LUT2 #(
		.INIT('h8)
	) name712 (
		_w736_,
		_w787_,
		_w788_
	);
	LUT2 #(
		.INIT('h1)
	) name713 (
		_w736_,
		_w787_,
		_w789_
	);
	LUT2 #(
		.INIT('h1)
	) name714 (
		_w788_,
		_w789_,
		_w790_
	);
	LUT2 #(
		.INIT('h1)
	) name715 (
		_w175_,
		_w790_,
		_w791_
	);
	LUT2 #(
		.INIT('h2)
	) name716 (
		_w183_,
		_w781_,
		_w792_
	);
	LUT2 #(
		.INIT('h4)
	) name717 (
		_w791_,
		_w792_,
		_w793_
	);
	LUT2 #(
		.INIT('h1)
	) name718 (
		_w780_,
		_w793_,
		_w794_
	);
	LUT2 #(
		.INIT('h2)
	) name719 (
		_w146_,
		_w215_,
		_w795_
	);
	LUT2 #(
		.INIT('h1)
	) name720 (
		_w762_,
		_w766_,
		_w796_
	);
	LUT2 #(
		.INIT('h8)
	) name721 (
		\inC15_pad ,
		_w79_,
		_w797_
	);
	LUT2 #(
		.INIT('h8)
	) name722 (
		\inA15_pad ,
		_w83_,
		_w798_
	);
	LUT2 #(
		.INIT('h8)
	) name723 (
		\inC15_pad ,
		\musel2_pad ,
		_w799_
	);
	LUT2 #(
		.INIT('h8)
	) name724 (
		\musel1_pad ,
		_w799_,
		_w800_
	);
	LUT2 #(
		.INIT('h1)
	) name725 (
		_w798_,
		_w800_,
		_w801_
	);
	LUT2 #(
		.INIT('h2)
	) name726 (
		_w81_,
		_w801_,
		_w802_
	);
	LUT2 #(
		.INIT('h1)
	) name727 (
		_w797_,
		_w802_,
		_w803_
	);
	LUT2 #(
		.INIT('h8)
	) name728 (
		\inD15_pad ,
		_w150_,
		_w804_
	);
	LUT2 #(
		.INIT('h8)
	) name729 (
		\inB15_pad ,
		_w152_,
		_w805_
	);
	LUT2 #(
		.INIT('h1)
	) name730 (
		_w804_,
		_w805_,
		_w806_
	);
	LUT2 #(
		.INIT('h1)
	) name731 (
		\musel1_pad ,
		_w806_,
		_w807_
	);
	LUT2 #(
		.INIT('h1)
	) name732 (
		_w494_,
		_w799_,
		_w808_
	);
	LUT2 #(
		.INIT('h2)
	) name733 (
		_w156_,
		_w808_,
		_w809_
	);
	LUT2 #(
		.INIT('h1)
	) name734 (
		_w807_,
		_w809_,
		_w810_
	);
	LUT2 #(
		.INIT('h1)
	) name735 (
		\musel4_pad ,
		_w810_,
		_w811_
	);
	LUT2 #(
		.INIT('h2)
	) name736 (
		_w803_,
		_w811_,
		_w812_
	);
	LUT2 #(
		.INIT('h4)
	) name737 (
		_w803_,
		_w811_,
		_w813_
	);
	LUT2 #(
		.INIT('h1)
	) name738 (
		_w812_,
		_w813_,
		_w814_
	);
	LUT2 #(
		.INIT('h8)
	) name739 (
		_w255_,
		_w814_,
		_w815_
	);
	LUT2 #(
		.INIT('h1)
	) name740 (
		_w255_,
		_w814_,
		_w816_
	);
	LUT2 #(
		.INIT('h1)
	) name741 (
		_w815_,
		_w816_,
		_w817_
	);
	LUT2 #(
		.INIT('h1)
	) name742 (
		_w763_,
		_w817_,
		_w818_
	);
	LUT2 #(
		.INIT('h4)
	) name743 (
		_w796_,
		_w818_,
		_w819_
	);
	LUT2 #(
		.INIT('h8)
	) name744 (
		_w796_,
		_w817_,
		_w820_
	);
	LUT2 #(
		.INIT('h2)
	) name745 (
		_w149_,
		_w819_,
		_w821_
	);
	LUT2 #(
		.INIT('h4)
	) name746 (
		_w820_,
		_w821_,
		_w822_
	);
	LUT2 #(
		.INIT('h1)
	) name747 (
		_w795_,
		_w822_,
		_w823_
	);
	LUT2 #(
		.INIT('h2)
	) name748 (
		_w76_,
		_w823_,
		_w824_
	);
	LUT2 #(
		.INIT('h8)
	) name749 (
		_w175_,
		_w215_,
		_w825_
	);
	LUT2 #(
		.INIT('h1)
	) name750 (
		_w175_,
		_w788_,
		_w826_
	);
	LUT2 #(
		.INIT('h2)
	) name751 (
		_w183_,
		_w825_,
		_w827_
	);
	LUT2 #(
		.INIT('h4)
	) name752 (
		_w826_,
		_w827_,
		_w828_
	);
	LUT2 #(
		.INIT('h1)
	) name753 (
		_w824_,
		_w828_,
		_w829_
	);
	LUT2 #(
		.INIT('h8)
	) name754 (
		\inD9_pad ,
		_w79_,
		_w830_
	);
	LUT2 #(
		.INIT('h8)
	) name755 (
		\inB9_pad ,
		_w83_,
		_w831_
	);
	LUT2 #(
		.INIT('h8)
	) name756 (
		\inD9_pad ,
		_w82_,
		_w832_
	);
	LUT2 #(
		.INIT('h1)
	) name757 (
		_w831_,
		_w832_,
		_w833_
	);
	LUT2 #(
		.INIT('h2)
	) name758 (
		_w81_,
		_w833_,
		_w834_
	);
	LUT2 #(
		.INIT('h1)
	) name759 (
		_w830_,
		_w834_,
		_w835_
	);
	LUT2 #(
		.INIT('h2)
	) name760 (
		\sh2_pad ,
		_w835_,
		_w836_
	);
	LUT2 #(
		.INIT('h1)
	) name761 (
		_w89_,
		_w836_,
		_w837_
	);
	LUT2 #(
		.INIT('h2)
	) name762 (
		\sh1_pad ,
		_w837_,
		_w838_
	);
	LUT2 #(
		.INIT('h1)
	) name763 (
		_w114_,
		_w838_,
		_w839_
	);
	LUT2 #(
		.INIT('h1)
	) name764 (
		\sh0_pad ,
		_w839_,
		_w840_
	);
	LUT2 #(
		.INIT('h8)
	) name765 (
		\inD6_pad ,
		_w79_,
		_w841_
	);
	LUT2 #(
		.INIT('h8)
	) name766 (
		\inB6_pad ,
		_w83_,
		_w842_
	);
	LUT2 #(
		.INIT('h8)
	) name767 (
		\inD6_pad ,
		_w82_,
		_w843_
	);
	LUT2 #(
		.INIT('h1)
	) name768 (
		_w842_,
		_w843_,
		_w844_
	);
	LUT2 #(
		.INIT('h2)
	) name769 (
		_w81_,
		_w844_,
		_w845_
	);
	LUT2 #(
		.INIT('h1)
	) name770 (
		_w841_,
		_w845_,
		_w846_
	);
	LUT2 #(
		.INIT('h2)
	) name771 (
		\sh2_pad ,
		_w846_,
		_w847_
	);
	LUT2 #(
		.INIT('h1)
	) name772 (
		_w130_,
		_w847_,
		_w848_
	);
	LUT2 #(
		.INIT('h1)
	) name773 (
		\sh1_pad ,
		_w848_,
		_w849_
	);
	LUT2 #(
		.INIT('h1)
	) name774 (
		\sh2_pad ,
		_w139_,
		_w850_
	);
	LUT2 #(
		.INIT('h2)
	) name775 (
		\sh2_pad ,
		_w111_,
		_w851_
	);
	LUT2 #(
		.INIT('h1)
	) name776 (
		_w850_,
		_w851_,
		_w852_
	);
	LUT2 #(
		.INIT('h2)
	) name777 (
		\sh1_pad ,
		_w852_,
		_w853_
	);
	LUT2 #(
		.INIT('h1)
	) name778 (
		_w849_,
		_w853_,
		_w854_
	);
	LUT2 #(
		.INIT('h2)
	) name779 (
		\sh0_pad ,
		_w854_,
		_w855_
	);
	LUT2 #(
		.INIT('h1)
	) name780 (
		_w840_,
		_w855_,
		_w856_
	);
	LUT2 #(
		.INIT('h2)
	) name781 (
		_w146_,
		_w856_,
		_w857_
	);
	LUT2 #(
		.INIT('h1)
	) name782 (
		_w372_,
		_w377_,
		_w858_
	);
	LUT2 #(
		.INIT('h1)
	) name783 (
		_w169_,
		_w379_,
		_w859_
	);
	LUT2 #(
		.INIT('h1)
	) name784 (
		_w858_,
		_w859_,
		_w860_
	);
	LUT2 #(
		.INIT('h8)
	) name785 (
		_w858_,
		_w859_,
		_w861_
	);
	LUT2 #(
		.INIT('h2)
	) name786 (
		_w149_,
		_w860_,
		_w862_
	);
	LUT2 #(
		.INIT('h4)
	) name787 (
		_w861_,
		_w862_,
		_w863_
	);
	LUT2 #(
		.INIT('h1)
	) name788 (
		_w857_,
		_w863_,
		_w864_
	);
	LUT2 #(
		.INIT('h2)
	) name789 (
		_w76_,
		_w864_,
		_w865_
	);
	LUT2 #(
		.INIT('h2)
	) name790 (
		_w175_,
		_w856_,
		_w866_
	);
	LUT2 #(
		.INIT('h2)
	) name791 (
		_w77_,
		_w533_,
		_w867_
	);
	LUT2 #(
		.INIT('h1)
	) name792 (
		_w526_,
		_w867_,
		_w868_
	);
	LUT2 #(
		.INIT('h1)
	) name793 (
		_w78_,
		_w530_,
		_w869_
	);
	LUT2 #(
		.INIT('h2)
	) name794 (
		_w526_,
		_w869_,
		_w870_
	);
	LUT2 #(
		.INIT('h1)
	) name795 (
		_w175_,
		_w870_,
		_w871_
	);
	LUT2 #(
		.INIT('h4)
	) name796 (
		_w868_,
		_w871_,
		_w872_
	);
	LUT2 #(
		.INIT('h1)
	) name797 (
		_w866_,
		_w872_,
		_w873_
	);
	LUT2 #(
		.INIT('h2)
	) name798 (
		_w183_,
		_w873_,
		_w874_
	);
	LUT2 #(
		.INIT('h1)
	) name799 (
		_w865_,
		_w874_,
		_w875_
	);
	LUT2 #(
		.INIT('h1)
	) name800 (
		_w221_,
		_w850_,
		_w876_
	);
	LUT2 #(
		.INIT('h2)
	) name801 (
		\sh1_pad ,
		_w876_,
		_w877_
	);
	LUT2 #(
		.INIT('h1)
	) name802 (
		_w849_,
		_w877_,
		_w878_
	);
	LUT2 #(
		.INIT('h1)
	) name803 (
		\sh0_pad ,
		_w878_,
		_w879_
	);
	LUT2 #(
		.INIT('h8)
	) name804 (
		\inD7_pad ,
		_w79_,
		_w880_
	);
	LUT2 #(
		.INIT('h8)
	) name805 (
		\inB7_pad ,
		_w83_,
		_w881_
	);
	LUT2 #(
		.INIT('h8)
	) name806 (
		\inD7_pad ,
		_w82_,
		_w882_
	);
	LUT2 #(
		.INIT('h1)
	) name807 (
		_w881_,
		_w882_,
		_w883_
	);
	LUT2 #(
		.INIT('h2)
	) name808 (
		_w81_,
		_w883_,
		_w884_
	);
	LUT2 #(
		.INIT('h1)
	) name809 (
		_w880_,
		_w884_,
		_w885_
	);
	LUT2 #(
		.INIT('h2)
	) name810 (
		\sh2_pad ,
		_w885_,
		_w886_
	);
	LUT2 #(
		.INIT('h1)
	) name811 (
		_w89_,
		_w886_,
		_w887_
	);
	LUT2 #(
		.INIT('h1)
	) name812 (
		\sh1_pad ,
		_w887_,
		_w888_
	);
	LUT2 #(
		.INIT('h1)
	) name813 (
		\sh2_pad ,
		_w104_,
		_w889_
	);
	LUT2 #(
		.INIT('h2)
	) name814 (
		\sh2_pad ,
		_w129_,
		_w890_
	);
	LUT2 #(
		.INIT('h1)
	) name815 (
		_w889_,
		_w890_,
		_w891_
	);
	LUT2 #(
		.INIT('h2)
	) name816 (
		\sh1_pad ,
		_w891_,
		_w892_
	);
	LUT2 #(
		.INIT('h1)
	) name817 (
		_w888_,
		_w892_,
		_w893_
	);
	LUT2 #(
		.INIT('h2)
	) name818 (
		\sh0_pad ,
		_w893_,
		_w894_
	);
	LUT2 #(
		.INIT('h1)
	) name819 (
		_w879_,
		_w894_,
		_w895_
	);
	LUT2 #(
		.INIT('h2)
	) name820 (
		_w146_,
		_w895_,
		_w896_
	);
	LUT2 #(
		.INIT('h1)
	) name821 (
		_w350_,
		_w376_,
		_w897_
	);
	LUT2 #(
		.INIT('h4)
	) name822 (
		_w372_,
		_w859_,
		_w898_
	);
	LUT2 #(
		.INIT('h8)
	) name823 (
		_w897_,
		_w898_,
		_w899_
	);
	LUT2 #(
		.INIT('h1)
	) name824 (
		_w377_,
		_w898_,
		_w900_
	);
	LUT2 #(
		.INIT('h4)
	) name825 (
		_w897_,
		_w900_,
		_w901_
	);
	LUT2 #(
		.INIT('h2)
	) name826 (
		_w149_,
		_w899_,
		_w902_
	);
	LUT2 #(
		.INIT('h4)
	) name827 (
		_w901_,
		_w902_,
		_w903_
	);
	LUT2 #(
		.INIT('h1)
	) name828 (
		_w896_,
		_w903_,
		_w904_
	);
	LUT2 #(
		.INIT('h2)
	) name829 (
		_w76_,
		_w904_,
		_w905_
	);
	LUT2 #(
		.INIT('h2)
	) name830 (
		_w175_,
		_w895_,
		_w906_
	);
	LUT2 #(
		.INIT('h1)
	) name831 (
		_w519_,
		_w870_,
		_w907_
	);
	LUT2 #(
		.INIT('h8)
	) name832 (
		_w519_,
		_w870_,
		_w908_
	);
	LUT2 #(
		.INIT('h1)
	) name833 (
		_w175_,
		_w907_,
		_w909_
	);
	LUT2 #(
		.INIT('h4)
	) name834 (
		_w908_,
		_w909_,
		_w910_
	);
	LUT2 #(
		.INIT('h1)
	) name835 (
		_w906_,
		_w910_,
		_w911_
	);
	LUT2 #(
		.INIT('h2)
	) name836 (
		_w183_,
		_w911_,
		_w912_
	);
	LUT2 #(
		.INIT('h1)
	) name837 (
		_w905_,
		_w912_,
		_w913_
	);
	LUT2 #(
		.INIT('h2)
	) name838 (
		\sh2_pad ,
		_w236_,
		_w914_
	);
	LUT2 #(
		.INIT('h1)
	) name839 (
		_w889_,
		_w914_,
		_w915_
	);
	LUT2 #(
		.INIT('h2)
	) name840 (
		\sh1_pad ,
		_w915_,
		_w916_
	);
	LUT2 #(
		.INIT('h1)
	) name841 (
		_w888_,
		_w916_,
		_w917_
	);
	LUT2 #(
		.INIT('h1)
	) name842 (
		\sh0_pad ,
		_w917_,
		_w918_
	);
	LUT2 #(
		.INIT('h1)
	) name843 (
		_w123_,
		_w850_,
		_w919_
	);
	LUT2 #(
		.INIT('h1)
	) name844 (
		\sh1_pad ,
		_w919_,
		_w920_
	);
	LUT2 #(
		.INIT('h1)
	) name845 (
		\sh2_pad ,
		_w846_,
		_w921_
	);
	LUT2 #(
		.INIT('h2)
	) name846 (
		\sh2_pad ,
		_w88_,
		_w922_
	);
	LUT2 #(
		.INIT('h1)
	) name847 (
		_w921_,
		_w922_,
		_w923_
	);
	LUT2 #(
		.INIT('h2)
	) name848 (
		\sh1_pad ,
		_w923_,
		_w924_
	);
	LUT2 #(
		.INIT('h1)
	) name849 (
		_w920_,
		_w924_,
		_w925_
	);
	LUT2 #(
		.INIT('h2)
	) name850 (
		\sh0_pad ,
		_w925_,
		_w926_
	);
	LUT2 #(
		.INIT('h1)
	) name851 (
		_w918_,
		_w926_,
		_w927_
	);
	LUT2 #(
		.INIT('h2)
	) name852 (
		_w146_,
		_w927_,
		_w928_
	);
	LUT2 #(
		.INIT('h1)
	) name853 (
		_w350_,
		_w900_,
		_w929_
	);
	LUT2 #(
		.INIT('h1)
	) name854 (
		_w330_,
		_w351_,
		_w930_
	);
	LUT2 #(
		.INIT('h8)
	) name855 (
		_w929_,
		_w930_,
		_w931_
	);
	LUT2 #(
		.INIT('h1)
	) name856 (
		_w376_,
		_w930_,
		_w932_
	);
	LUT2 #(
		.INIT('h4)
	) name857 (
		_w929_,
		_w932_,
		_w933_
	);
	LUT2 #(
		.INIT('h2)
	) name858 (
		_w149_,
		_w931_,
		_w934_
	);
	LUT2 #(
		.INIT('h4)
	) name859 (
		_w933_,
		_w934_,
		_w935_
	);
	LUT2 #(
		.INIT('h1)
	) name860 (
		_w928_,
		_w935_,
		_w936_
	);
	LUT2 #(
		.INIT('h2)
	) name861 (
		_w76_,
		_w936_,
		_w937_
	);
	LUT2 #(
		.INIT('h2)
	) name862 (
		_w77_,
		_w524_,
		_w938_
	);
	LUT2 #(
		.INIT('h4)
	) name863 (
		_w908_,
		_w938_,
		_w939_
	);
	LUT2 #(
		.INIT('h8)
	) name864 (
		_w524_,
		_w908_,
		_w940_
	);
	LUT2 #(
		.INIT('h1)
	) name865 (
		_w175_,
		_w939_,
		_w941_
	);
	LUT2 #(
		.INIT('h4)
	) name866 (
		_w940_,
		_w941_,
		_w942_
	);
	LUT2 #(
		.INIT('h8)
	) name867 (
		_w175_,
		_w927_,
		_w943_
	);
	LUT2 #(
		.INIT('h2)
	) name868 (
		_w183_,
		_w942_,
		_w944_
	);
	LUT2 #(
		.INIT('h4)
	) name869 (
		_w943_,
		_w944_,
		_w945_
	);
	LUT2 #(
		.INIT('h1)
	) name870 (
		_w937_,
		_w945_,
		_w946_
	);
	LUT2 #(
		.INIT('h2)
	) name871 (
		\sh2_pad ,
		_w208_,
		_w947_
	);
	LUT2 #(
		.INIT('h1)
	) name872 (
		_w921_,
		_w947_,
		_w948_
	);
	LUT2 #(
		.INIT('h2)
	) name873 (
		\sh1_pad ,
		_w948_,
		_w949_
	);
	LUT2 #(
		.INIT('h1)
	) name874 (
		_w920_,
		_w949_,
		_w950_
	);
	LUT2 #(
		.INIT('h1)
	) name875 (
		\sh0_pad ,
		_w950_,
		_w951_
	);
	LUT2 #(
		.INIT('h1)
	) name876 (
		_w836_,
		_w889_,
		_w952_
	);
	LUT2 #(
		.INIT('h1)
	) name877 (
		\sh1_pad ,
		_w952_,
		_w953_
	);
	LUT2 #(
		.INIT('h1)
	) name878 (
		\sh2_pad ,
		_w885_,
		_w954_
	);
	LUT2 #(
		.INIT('h1)
	) name879 (
		_w140_,
		_w954_,
		_w955_
	);
	LUT2 #(
		.INIT('h2)
	) name880 (
		\sh1_pad ,
		_w955_,
		_w956_
	);
	LUT2 #(
		.INIT('h1)
	) name881 (
		_w953_,
		_w956_,
		_w957_
	);
	LUT2 #(
		.INIT('h2)
	) name882 (
		\sh0_pad ,
		_w957_,
		_w958_
	);
	LUT2 #(
		.INIT('h1)
	) name883 (
		_w951_,
		_w958_,
		_w959_
	);
	LUT2 #(
		.INIT('h2)
	) name884 (
		_w146_,
		_w959_,
		_w960_
	);
	LUT2 #(
		.INIT('h1)
	) name885 (
		_w310_,
		_w452_,
		_w961_
	);
	LUT2 #(
		.INIT('h4)
	) name886 (
		_w386_,
		_w961_,
		_w962_
	);
	LUT2 #(
		.INIT('h2)
	) name887 (
		_w386_,
		_w961_,
		_w963_
	);
	LUT2 #(
		.INIT('h2)
	) name888 (
		_w149_,
		_w962_,
		_w964_
	);
	LUT2 #(
		.INIT('h4)
	) name889 (
		_w963_,
		_w964_,
		_w965_
	);
	LUT2 #(
		.INIT('h1)
	) name890 (
		_w960_,
		_w965_,
		_w966_
	);
	LUT2 #(
		.INIT('h2)
	) name891 (
		_w76_,
		_w966_,
		_w967_
	);
	LUT2 #(
		.INIT('h8)
	) name892 (
		_w501_,
		_w536_,
		_w968_
	);
	LUT2 #(
		.INIT('h2)
	) name893 (
		_w77_,
		_w655_,
		_w969_
	);
	LUT2 #(
		.INIT('h8)
	) name894 (
		_w968_,
		_w969_,
		_w970_
	);
	LUT2 #(
		.INIT('h1)
	) name895 (
		_w968_,
		_w969_,
		_w971_
	);
	LUT2 #(
		.INIT('h1)
	) name896 (
		_w970_,
		_w971_,
		_w972_
	);
	LUT2 #(
		.INIT('h1)
	) name897 (
		_w175_,
		_w972_,
		_w973_
	);
	LUT2 #(
		.INIT('h8)
	) name898 (
		_w175_,
		_w959_,
		_w974_
	);
	LUT2 #(
		.INIT('h2)
	) name899 (
		_w183_,
		_w973_,
		_w975_
	);
	LUT2 #(
		.INIT('h4)
	) name900 (
		_w974_,
		_w975_,
		_w976_
	);
	LUT2 #(
		.INIT('h1)
	) name901 (
		_w967_,
		_w976_,
		_w977_
	);
	LUT2 #(
		.INIT('h2)
	) name902 (
		\sh2_pad ,
		_w227_,
		_w978_
	);
	LUT2 #(
		.INIT('h1)
	) name903 (
		_w954_,
		_w978_,
		_w979_
	);
	LUT2 #(
		.INIT('h2)
	) name904 (
		\sh1_pad ,
		_w979_,
		_w980_
	);
	LUT2 #(
		.INIT('h1)
	) name905 (
		_w953_,
		_w980_,
		_w981_
	);
	LUT2 #(
		.INIT('h1)
	) name906 (
		\sh0_pad ,
		_w981_,
		_w982_
	);
	LUT2 #(
		.INIT('h1)
	) name907 (
		_w221_,
		_w921_,
		_w983_
	);
	LUT2 #(
		.INIT('h1)
	) name908 (
		\sh1_pad ,
		_w983_,
		_w984_
	);
	LUT2 #(
		.INIT('h1)
	) name909 (
		\sh2_pad ,
		_w122_,
		_w985_
	);
	LUT2 #(
		.INIT('h1)
	) name910 (
		_w105_,
		_w985_,
		_w986_
	);
	LUT2 #(
		.INIT('h2)
	) name911 (
		\sh1_pad ,
		_w986_,
		_w987_
	);
	LUT2 #(
		.INIT('h1)
	) name912 (
		_w984_,
		_w987_,
		_w988_
	);
	LUT2 #(
		.INIT('h2)
	) name913 (
		\sh0_pad ,
		_w988_,
		_w989_
	);
	LUT2 #(
		.INIT('h1)
	) name914 (
		_w982_,
		_w989_,
		_w990_
	);
	LUT2 #(
		.INIT('h2)
	) name915 (
		_w146_,
		_w990_,
		_w991_
	);
	LUT2 #(
		.INIT('h1)
	) name916 (
		_w448_,
		_w454_,
		_w992_
	);
	LUT2 #(
		.INIT('h1)
	) name917 (
		_w452_,
		_w992_,
		_w993_
	);
	LUT2 #(
		.INIT('h4)
	) name918 (
		_w387_,
		_w993_,
		_w994_
	);
	LUT2 #(
		.INIT('h8)
	) name919 (
		_w387_,
		_w992_,
		_w995_
	);
	LUT2 #(
		.INIT('h2)
	) name920 (
		_w149_,
		_w994_,
		_w996_
	);
	LUT2 #(
		.INIT('h4)
	) name921 (
		_w995_,
		_w996_,
		_w997_
	);
	LUT2 #(
		.INIT('h1)
	) name922 (
		_w991_,
		_w997_,
		_w998_
	);
	LUT2 #(
		.INIT('h2)
	) name923 (
		_w76_,
		_w998_,
		_w999_
	);
	LUT2 #(
		.INIT('h1)
	) name924 (
		_w664_,
		_w970_,
		_w1000_
	);
	LUT2 #(
		.INIT('h1)
	) name925 (
		_w78_,
		_w660_,
		_w1001_
	);
	LUT2 #(
		.INIT('h2)
	) name926 (
		_w970_,
		_w1001_,
		_w1002_
	);
	LUT2 #(
		.INIT('h1)
	) name927 (
		_w1000_,
		_w1002_,
		_w1003_
	);
	LUT2 #(
		.INIT('h1)
	) name928 (
		_w175_,
		_w1003_,
		_w1004_
	);
	LUT2 #(
		.INIT('h8)
	) name929 (
		_w175_,
		_w990_,
		_w1005_
	);
	LUT2 #(
		.INIT('h2)
	) name930 (
		_w183_,
		_w1004_,
		_w1006_
	);
	LUT2 #(
		.INIT('h4)
	) name931 (
		_w1005_,
		_w1006_,
		_w1007_
	);
	LUT2 #(
		.INIT('h1)
	) name932 (
		_w999_,
		_w1007_,
		_w1008_
	);
	LUT2 #(
		.INIT('h1)
	) name933 (
		_w193_,
		_w985_,
		_w1009_
	);
	LUT2 #(
		.INIT('h2)
	) name934 (
		\sh1_pad ,
		_w1009_,
		_w1010_
	);
	LUT2 #(
		.INIT('h1)
	) name935 (
		_w984_,
		_w1010_,
		_w1011_
	);
	LUT2 #(
		.INIT('h1)
	) name936 (
		\sh0_pad ,
		_w1011_,
		_w1012_
	);
	LUT2 #(
		.INIT('h1)
	) name937 (
		_w914_,
		_w954_,
		_w1013_
	);
	LUT2 #(
		.INIT('h1)
	) name938 (
		\sh1_pad ,
		_w1013_,
		_w1014_
	);
	LUT2 #(
		.INIT('h1)
	) name939 (
		\sh2_pad ,
		_w835_,
		_w1015_
	);
	LUT2 #(
		.INIT('h1)
	) name940 (
		_w847_,
		_w1015_,
		_w1016_
	);
	LUT2 #(
		.INIT('h2)
	) name941 (
		\sh1_pad ,
		_w1016_,
		_w1017_
	);
	LUT2 #(
		.INIT('h1)
	) name942 (
		_w1014_,
		_w1017_,
		_w1018_
	);
	LUT2 #(
		.INIT('h2)
	) name943 (
		\sh0_pad ,
		_w1018_,
		_w1019_
	);
	LUT2 #(
		.INIT('h1)
	) name944 (
		_w1012_,
		_w1019_,
		_w1020_
	);
	LUT2 #(
		.INIT('h2)
	) name945 (
		_w146_,
		_w1020_,
		_w1021_
	);
	LUT2 #(
		.INIT('h1)
	) name946 (
		_w407_,
		_w455_,
		_w1022_
	);
	LUT2 #(
		.INIT('h1)
	) name947 (
		_w387_,
		_w454_,
		_w1023_
	);
	LUT2 #(
		.INIT('h1)
	) name948 (
		_w448_,
		_w1023_,
		_w1024_
	);
	LUT2 #(
		.INIT('h1)
	) name949 (
		_w453_,
		_w1022_,
		_w1025_
	);
	LUT2 #(
		.INIT('h4)
	) name950 (
		_w1024_,
		_w1025_,
		_w1026_
	);
	LUT2 #(
		.INIT('h4)
	) name951 (
		_w407_,
		_w1024_,
		_w1027_
	);
	LUT2 #(
		.INIT('h4)
	) name952 (
		_w455_,
		_w1027_,
		_w1028_
	);
	LUT2 #(
		.INIT('h2)
	) name953 (
		_w149_,
		_w1026_,
		_w1029_
	);
	LUT2 #(
		.INIT('h4)
	) name954 (
		_w1028_,
		_w1029_,
		_w1030_
	);
	LUT2 #(
		.INIT('h1)
	) name955 (
		_w1021_,
		_w1030_,
		_w1031_
	);
	LUT2 #(
		.INIT('h2)
	) name956 (
		_w76_,
		_w1031_,
		_w1032_
	);
	LUT2 #(
		.INIT('h8)
	) name957 (
		_w175_,
		_w1020_,
		_w1033_
	);
	LUT2 #(
		.INIT('h8)
	) name958 (
		_w496_,
		_w657_,
		_w1034_
	);
	LUT2 #(
		.INIT('h2)
	) name959 (
		_w501_,
		_w657_,
		_w1035_
	);
	LUT2 #(
		.INIT('h2)
	) name960 (
		_w178_,
		_w1034_,
		_w1036_
	);
	LUT2 #(
		.INIT('h4)
	) name961 (
		_w1035_,
		_w1036_,
		_w1037_
	);
	LUT2 #(
		.INIT('h8)
	) name962 (
		_w1002_,
		_w1037_,
		_w1038_
	);
	LUT2 #(
		.INIT('h1)
	) name963 (
		_w1002_,
		_w1037_,
		_w1039_
	);
	LUT2 #(
		.INIT('h1)
	) name964 (
		_w1038_,
		_w1039_,
		_w1040_
	);
	LUT2 #(
		.INIT('h1)
	) name965 (
		_w175_,
		_w1040_,
		_w1041_
	);
	LUT2 #(
		.INIT('h2)
	) name966 (
		_w183_,
		_w1033_,
		_w1042_
	);
	LUT2 #(
		.INIT('h4)
	) name967 (
		_w1041_,
		_w1042_,
		_w1043_
	);
	LUT2 #(
		.INIT('h1)
	) name968 (
		_w1032_,
		_w1043_,
		_w1044_
	);
	LUT2 #(
		.INIT('h1)
	) name969 (
		_w216_,
		_w1015_,
		_w1045_
	);
	LUT2 #(
		.INIT('h2)
	) name970 (
		\sh1_pad ,
		_w1045_,
		_w1046_
	);
	LUT2 #(
		.INIT('h1)
	) name971 (
		_w1014_,
		_w1046_,
		_w1047_
	);
	LUT2 #(
		.INIT('h1)
	) name972 (
		\sh0_pad ,
		_w1047_,
		_w1048_
	);
	LUT2 #(
		.INIT('h1)
	) name973 (
		_w947_,
		_w985_,
		_w1049_
	);
	LUT2 #(
		.INIT('h1)
	) name974 (
		\sh1_pad ,
		_w1049_,
		_w1050_
	);
	LUT2 #(
		.INIT('h1)
	) name975 (
		_w200_,
		_w886_,
		_w1051_
	);
	LUT2 #(
		.INIT('h2)
	) name976 (
		\sh1_pad ,
		_w1051_,
		_w1052_
	);
	LUT2 #(
		.INIT('h1)
	) name977 (
		_w1050_,
		_w1052_,
		_w1053_
	);
	LUT2 #(
		.INIT('h2)
	) name978 (
		\sh0_pad ,
		_w1053_,
		_w1054_
	);
	LUT2 #(
		.INIT('h1)
	) name979 (
		_w1048_,
		_w1054_,
		_w1055_
	);
	LUT2 #(
		.INIT('h2)
	) name980 (
		_w146_,
		_w1055_,
		_w1056_
	);
	LUT2 #(
		.INIT('h1)
	) name981 (
		_w427_,
		_w451_,
		_w1057_
	);
	LUT2 #(
		.INIT('h8)
	) name982 (
		_w1027_,
		_w1057_,
		_w1058_
	);
	LUT2 #(
		.INIT('h1)
	) name983 (
		_w455_,
		_w1057_,
		_w1059_
	);
	LUT2 #(
		.INIT('h4)
	) name984 (
		_w1027_,
		_w1059_,
		_w1060_
	);
	LUT2 #(
		.INIT('h2)
	) name985 (
		_w149_,
		_w1058_,
		_w1061_
	);
	LUT2 #(
		.INIT('h4)
	) name986 (
		_w1060_,
		_w1061_,
		_w1062_
	);
	LUT2 #(
		.INIT('h1)
	) name987 (
		_w1056_,
		_w1062_,
		_w1063_
	);
	LUT2 #(
		.INIT('h2)
	) name988 (
		_w76_,
		_w1063_,
		_w1064_
	);
	LUT2 #(
		.INIT('h2)
	) name989 (
		_w77_,
		_w666_,
		_w1065_
	);
	LUT2 #(
		.INIT('h8)
	) name990 (
		_w497_,
		_w1065_,
		_w1066_
	);
	LUT2 #(
		.INIT('h1)
	) name991 (
		_w667_,
		_w1066_,
		_w1067_
	);
	LUT2 #(
		.INIT('h2)
	) name992 (
		_w1038_,
		_w1067_,
		_w1068_
	);
	LUT2 #(
		.INIT('h4)
	) name993 (
		_w1038_,
		_w1067_,
		_w1069_
	);
	LUT2 #(
		.INIT('h1)
	) name994 (
		_w1068_,
		_w1069_,
		_w1070_
	);
	LUT2 #(
		.INIT('h1)
	) name995 (
		_w175_,
		_w1070_,
		_w1071_
	);
	LUT2 #(
		.INIT('h8)
	) name996 (
		_w175_,
		_w1055_,
		_w1072_
	);
	LUT2 #(
		.INIT('h2)
	) name997 (
		_w183_,
		_w1072_,
		_w1073_
	);
	LUT2 #(
		.INIT('h4)
	) name998 (
		_w1071_,
		_w1073_,
		_w1074_
	);
	LUT2 #(
		.INIT('h1)
	) name999 (
		_w1064_,
		_w1074_,
		_w1075_
	);
	LUT2 #(
		.INIT('h1)
	) name1000 (
		_w200_,
		_w216_,
		_w1076_
	);
	LUT2 #(
		.INIT('h2)
	) name1001 (
		\sh1_pad ,
		_w1076_,
		_w1077_
	);
	LUT2 #(
		.INIT('h1)
	) name1002 (
		_w1050_,
		_w1077_,
		_w1078_
	);
	LUT2 #(
		.INIT('h1)
	) name1003 (
		\sh0_pad ,
		_w1078_,
		_w1079_
	);
	LUT2 #(
		.INIT('h1)
	) name1004 (
		_w978_,
		_w1015_,
		_w1080_
	);
	LUT2 #(
		.INIT('h1)
	) name1005 (
		\sh1_pad ,
		_w1080_,
		_w1081_
	);
	LUT2 #(
		.INIT('h1)
	) name1006 (
		_w123_,
		_w237_,
		_w1082_
	);
	LUT2 #(
		.INIT('h2)
	) name1007 (
		\sh1_pad ,
		_w1082_,
		_w1083_
	);
	LUT2 #(
		.INIT('h1)
	) name1008 (
		_w1081_,
		_w1083_,
		_w1084_
	);
	LUT2 #(
		.INIT('h2)
	) name1009 (
		\sh0_pad ,
		_w1084_,
		_w1085_
	);
	LUT2 #(
		.INIT('h1)
	) name1010 (
		_w1079_,
		_w1085_,
		_w1086_
	);
	LUT2 #(
		.INIT('h2)
	) name1011 (
		_w146_,
		_w1086_,
		_w1087_
	);
	LUT2 #(
		.INIT('h1)
	) name1012 (
		_w289_,
		_w290_,
		_w1088_
	);
	LUT2 #(
		.INIT('h4)
	) name1013 (
		_w460_,
		_w1088_,
		_w1089_
	);
	LUT2 #(
		.INIT('h2)
	) name1014 (
		_w460_,
		_w1088_,
		_w1090_
	);
	LUT2 #(
		.INIT('h2)
	) name1015 (
		_w149_,
		_w1089_,
		_w1091_
	);
	LUT2 #(
		.INIT('h4)
	) name1016 (
		_w1090_,
		_w1091_,
		_w1092_
	);
	LUT2 #(
		.INIT('h1)
	) name1017 (
		_w1087_,
		_w1092_,
		_w1093_
	);
	LUT2 #(
		.INIT('h2)
	) name1018 (
		_w76_,
		_w1093_,
		_w1094_
	);
	LUT2 #(
		.INIT('h2)
	) name1019 (
		_w175_,
		_w1086_,
		_w1095_
	);
	LUT2 #(
		.INIT('h4)
	) name1020 (
		_w175_,
		_w549_,
		_w1096_
	);
	LUT2 #(
		.INIT('h4)
	) name1021 (
		_w513_,
		_w1096_,
		_w1097_
	);
	LUT2 #(
		.INIT('h1)
	) name1022 (
		_w1095_,
		_w1097_,
		_w1098_
	);
	LUT2 #(
		.INIT('h2)
	) name1023 (
		_w183_,
		_w1098_,
		_w1099_
	);
	LUT2 #(
		.INIT('h1)
	) name1024 (
		_w1094_,
		_w1099_,
		_w1100_
	);
	LUT2 #(
		.INIT('h2)
	) name1025 (
		\sh1_pad ,
		_w238_,
		_w1101_
	);
	LUT2 #(
		.INIT('h1)
	) name1026 (
		_w1081_,
		_w1101_,
		_w1102_
	);
	LUT2 #(
		.INIT('h1)
	) name1027 (
		\sh0_pad ,
		_w1102_,
		_w1103_
	);
	LUT2 #(
		.INIT('h1)
	) name1028 (
		_w209_,
		_w836_,
		_w1104_
	);
	LUT2 #(
		.INIT('h2)
	) name1029 (
		\sh1_pad ,
		_w1104_,
		_w1105_
	);
	LUT2 #(
		.INIT('h1)
	) name1030 (
		_w202_,
		_w1105_,
		_w1106_
	);
	LUT2 #(
		.INIT('h2)
	) name1031 (
		\sh0_pad ,
		_w1106_,
		_w1107_
	);
	LUT2 #(
		.INIT('h1)
	) name1032 (
		_w1103_,
		_w1107_,
		_w1108_
	);
	LUT2 #(
		.INIT('h2)
	) name1033 (
		_w146_,
		_w1108_,
		_w1109_
	);
	LUT2 #(
		.INIT('h1)
	) name1034 (
		_w268_,
		_w269_,
		_w1110_
	);
	LUT2 #(
		.INIT('h1)
	) name1035 (
		_w462_,
		_w1110_,
		_w1111_
	);
	LUT2 #(
		.INIT('h8)
	) name1036 (
		_w462_,
		_w1110_,
		_w1112_
	);
	LUT2 #(
		.INIT('h2)
	) name1037 (
		_w149_,
		_w1111_,
		_w1113_
	);
	LUT2 #(
		.INIT('h4)
	) name1038 (
		_w1112_,
		_w1113_,
		_w1114_
	);
	LUT2 #(
		.INIT('h1)
	) name1039 (
		_w1109_,
		_w1114_,
		_w1115_
	);
	LUT2 #(
		.INIT('h2)
	) name1040 (
		_w76_,
		_w1115_,
		_w1116_
	);
	LUT2 #(
		.INIT('h2)
	) name1041 (
		_w175_,
		_w1108_,
		_w1117_
	);
	LUT2 #(
		.INIT('h4)
	) name1042 (
		_w508_,
		_w1096_,
		_w1118_
	);
	LUT2 #(
		.INIT('h1)
	) name1043 (
		_w1117_,
		_w1118_,
		_w1119_
	);
	LUT2 #(
		.INIT('h2)
	) name1044 (
		_w183_,
		_w1119_,
		_w1120_
	);
	LUT2 #(
		.INIT('h1)
	) name1045 (
		_w1116_,
		_w1120_,
		_w1121_
	);
	assign \O0_pad  = _w186_ ;
	assign \O10_pad  = _w555_ ;
	assign \O11_pad  = _w606_ ;
	assign \O12_pad  = _w685_ ;
	assign \O13_pad  = _w741_ ;
	assign \O14_pad  = _w794_ ;
	assign \O15_pad  = _w829_ ;
	assign \O1_pad  = _w875_ ;
	assign \O2_pad  = _w913_ ;
	assign \O3_pad  = _w946_ ;
	assign \O4_pad  = _w977_ ;
	assign \O5_pad  = _w1008_ ;
	assign \O6_pad  = _w1044_ ;
	assign \O7_pad  = _w1075_ ;
	assign \O8_pad  = _w1100_ ;
	assign \O9_pad  = _w1121_ ;
endmodule;