module top (\addroundkey_ready_o_reg/NET0131 , \addroundkey_round_reg[0]/NET0131 , \addroundkey_round_reg[1]/NET0131 , \addroundkey_round_reg[2]/NET0131 , \addroundkey_round_reg[3]/NET0131 , \addroundkey_start_i_reg/NET0131 , \data_i[0]_pad , \data_i[100]_pad , \data_i[101]_pad , \data_i[102]_pad , \data_i[103]_pad , \data_i[104]_pad , \data_i[105]_pad , \data_i[106]_pad , \data_i[107]_pad , \data_i[108]_pad , \data_i[109]_pad , \data_i[10]_pad , \data_i[110]_pad , \data_i[111]_pad , \data_i[112]_pad , \data_i[113]_pad , \data_i[114]_pad , \data_i[115]_pad , \data_i[116]_pad , \data_i[117]_pad , \data_i[118]_pad , \data_i[119]_pad , \data_i[11]_pad , \data_i[120]_pad , \data_i[121]_pad , \data_i[122]_pad , \data_i[123]_pad , \data_i[124]_pad , \data_i[125]_pad , \data_i[126]_pad , \data_i[127]_pad , \data_i[12]_pad , \data_i[13]_pad , \data_i[14]_pad , \data_i[15]_pad , \data_i[16]_pad , \data_i[17]_pad , \data_i[18]_pad , \data_i[19]_pad , \data_i[1]_pad , \data_i[20]_pad , \data_i[21]_pad , \data_i[22]_pad , \data_i[23]_pad , \data_i[24]_pad , \data_i[25]_pad , \data_i[26]_pad , \data_i[27]_pad , \data_i[28]_pad , \data_i[29]_pad , \data_i[2]_pad , \data_i[30]_pad , \data_i[31]_pad , \data_i[32]_pad , \data_i[33]_pad , \data_i[34]_pad , \data_i[35]_pad , \data_i[36]_pad , \data_i[37]_pad , \data_i[38]_pad , \data_i[39]_pad , \data_i[3]_pad , \data_i[40]_pad , \data_i[41]_pad , \data_i[42]_pad , \data_i[43]_pad , \data_i[44]_pad , \data_i[45]_pad , \data_i[46]_pad , \data_i[47]_pad , \data_i[48]_pad , \data_i[49]_pad , \data_i[4]_pad , \data_i[50]_pad , \data_i[51]_pad , \data_i[52]_pad , \data_i[53]_pad , \data_i[54]_pad , \data_i[55]_pad , \data_i[56]_pad , \data_i[57]_pad , \data_i[58]_pad , \data_i[59]_pad , \data_i[5]_pad , \data_i[60]_pad , \data_i[61]_pad , \data_i[62]_pad , \data_i[63]_pad , \data_i[64]_pad , \data_i[65]_pad , \data_i[66]_pad , \data_i[67]_pad , \data_i[68]_pad , \data_i[69]_pad , \data_i[6]_pad , \data_i[70]_pad , \data_i[71]_pad , \data_i[72]_pad , \data_i[73]_pad , \data_i[74]_pad , \data_i[75]_pad , \data_i[76]_pad , \data_i[77]_pad , \data_i[78]_pad , \data_i[79]_pad , \data_i[7]_pad , \data_i[80]_pad , \data_i[81]_pad , \data_i[82]_pad , \data_i[83]_pad , \data_i[84]_pad , \data_i[85]_pad , \data_i[86]_pad , \data_i[87]_pad , \data_i[88]_pad , \data_i[89]_pad , \data_i[8]_pad , \data_i[90]_pad , \data_i[91]_pad , \data_i[92]_pad , \data_i[93]_pad , \data_i[94]_pad , \data_i[95]_pad , \data_i[96]_pad , \data_i[97]_pad , \data_i[98]_pad , \data_i[99]_pad , \data_i[9]_pad , \data_o[0]_pad , \data_o[100]_pad , \data_o[101]_pad , \data_o[102]_pad , \data_o[103]_pad , \data_o[104]_pad , \data_o[105]_pad , \data_o[106]_pad , \data_o[107]_pad , \data_o[108]_pad , \data_o[109]_pad , \data_o[10]_pad , \data_o[110]_pad , \data_o[111]_pad , \data_o[112]_pad , \data_o[113]_pad , \data_o[114]_pad , \data_o[115]_pad , \data_o[116]_pad , \data_o[117]_pad , \data_o[118]_pad , \data_o[119]_pad , \data_o[11]_pad , \data_o[120]_pad , \data_o[121]_pad , \data_o[122]_pad , \data_o[123]_pad , \data_o[124]_pad , \data_o[125]_pad , \data_o[126]_pad , \data_o[127]_pad , \data_o[12]_pad , \data_o[13]_pad , \data_o[14]_pad , \data_o[15]_pad , \data_o[16]_pad , \data_o[17]_pad , \data_o[18]_pad , \data_o[19]_pad , \data_o[1]_pad , \data_o[20]_pad , \data_o[21]_pad , \data_o[22]_pad , \data_o[23]_pad , \data_o[24]_pad , \data_o[25]_pad , \data_o[26]_pad , \data_o[27]_pad , \data_o[28]_pad , \data_o[29]_pad , \data_o[2]_pad , \data_o[30]_pad , \data_o[31]_pad , \data_o[32]_pad , \data_o[33]_pad , \data_o[34]_pad , \data_o[35]_pad , \data_o[36]_pad , \data_o[37]_pad , \data_o[38]_pad , \data_o[39]_pad , \data_o[3]_pad , \data_o[40]_pad , \data_o[41]_pad , \data_o[42]_pad , \data_o[43]_pad , \data_o[44]_pad , \data_o[45]_pad , \data_o[46]_pad , \data_o[47]_pad , \data_o[48]_pad , \data_o[49]_pad , \data_o[4]_pad , \data_o[50]_pad , \data_o[51]_pad , \data_o[52]_pad , \data_o[53]_pad , \data_o[54]_pad , \data_o[55]_pad , \data_o[56]_pad , \data_o[57]_pad , \data_o[58]_pad , \data_o[59]_pad , \data_o[5]_pad , \data_o[60]_pad , \data_o[61]_pad , \data_o[62]_pad , \data_o[63]_pad , \data_o[64]_pad , \data_o[65]_pad , \data_o[66]_pad , \data_o[67]_pad , \data_o[68]_pad , \data_o[69]_pad , \data_o[6]_pad , \data_o[70]_pad , \data_o[71]_pad , \data_o[72]_pad , \data_o[73]_pad , \data_o[74]_pad , \data_o[75]_pad , \data_o[76]_pad , \data_o[77]_pad , \data_o[78]_pad , \data_o[79]_pad , \data_o[7]_pad , \data_o[80]_pad , \data_o[81]_pad , \data_o[82]_pad , \data_o[83]_pad , \data_o[84]_pad , \data_o[85]_pad , \data_o[86]_pad , \data_o[87]_pad , \data_o[88]_pad , \data_o[89]_pad , \data_o[8]_pad , \data_o[90]_pad , \data_o[91]_pad , \data_o[92]_pad , \data_o[93]_pad , \data_o[94]_pad , \data_o[95]_pad , \data_o[96]_pad , \data_o[97]_pad , \data_o[98]_pad , \data_o[99]_pad , \data_o[9]_pad , decrypt_i_pad, \first_round_reg_reg/NET0131 , \key_i[0]_pad , \key_i[100]_pad , \key_i[101]_pad , \key_i[102]_pad , \key_i[103]_pad , \key_i[104]_pad , \key_i[105]_pad , \key_i[106]_pad , \key_i[107]_pad , \key_i[108]_pad , \key_i[109]_pad , \key_i[10]_pad , \key_i[110]_pad , \key_i[111]_pad , \key_i[112]_pad , \key_i[113]_pad , \key_i[114]_pad , \key_i[115]_pad , \key_i[116]_pad , \key_i[117]_pad , \key_i[118]_pad , \key_i[119]_pad , \key_i[11]_pad , \key_i[120]_pad , \key_i[121]_pad , \key_i[122]_pad , \key_i[123]_pad , \key_i[124]_pad , \key_i[125]_pad , \key_i[126]_pad , \key_i[127]_pad , \key_i[12]_pad , \key_i[13]_pad , \key_i[14]_pad , \key_i[15]_pad , \key_i[16]_pad , \key_i[17]_pad , \key_i[18]_pad , \key_i[19]_pad , \key_i[1]_pad , \key_i[20]_pad , \key_i[21]_pad , \key_i[22]_pad , \key_i[23]_pad , \key_i[24]_pad , \key_i[25]_pad , \key_i[26]_pad , \key_i[27]_pad , \key_i[28]_pad , \key_i[29]_pad , \key_i[2]_pad , \key_i[30]_pad , \key_i[31]_pad , \key_i[32]_pad , \key_i[33]_pad , \key_i[34]_pad , \key_i[35]_pad , \key_i[36]_pad , \key_i[37]_pad , \key_i[38]_pad , \key_i[39]_pad , \key_i[3]_pad , \key_i[40]_pad , \key_i[41]_pad , \key_i[42]_pad , \key_i[43]_pad , \key_i[44]_pad , \key_i[45]_pad , \key_i[46]_pad , \key_i[47]_pad , \key_i[48]_pad , \key_i[49]_pad , \key_i[4]_pad , \key_i[50]_pad , \key_i[51]_pad , \key_i[52]_pad , \key_i[53]_pad , \key_i[54]_pad , \key_i[55]_pad , \key_i[56]_pad , \key_i[57]_pad , \key_i[58]_pad , \key_i[59]_pad , \key_i[5]_pad , \key_i[60]_pad , \key_i[61]_pad , \key_i[62]_pad , \key_i[63]_pad , \key_i[64]_pad , \key_i[65]_pad , \key_i[66]_pad , \key_i[67]_pad , \key_i[68]_pad , \key_i[69]_pad , \key_i[6]_pad , \key_i[70]_pad , \key_i[71]_pad , \key_i[72]_pad , \key_i[73]_pad , \key_i[74]_pad , \key_i[75]_pad , \key_i[76]_pad , \key_i[77]_pad , \key_i[78]_pad , \key_i[79]_pad , \key_i[7]_pad , \key_i[80]_pad , \key_i[81]_pad , \key_i[82]_pad , \key_i[83]_pad , \key_i[84]_pad , \key_i[85]_pad , \key_i[86]_pad , \key_i[87]_pad , \key_i[88]_pad , \key_i[89]_pad , \key_i[8]_pad , \key_i[90]_pad , \key_i[91]_pad , \key_i[92]_pad , \key_i[93]_pad , \key_i[94]_pad , \key_i[95]_pad , \key_i[96]_pad , \key_i[97]_pad , \key_i[98]_pad , \key_i[99]_pad , \key_i[9]_pad , \ks1_col_reg[0]/NET0131 , \ks1_col_reg[16]/NET0131 , \ks1_col_reg[17]/NET0131 , \ks1_col_reg[18]/NET0131 , \ks1_col_reg[19]/NET0131 , \ks1_col_reg[1]/NET0131 , \ks1_col_reg[20]/NET0131 , \ks1_col_reg[21]/NET0131 , \ks1_col_reg[22]/NET0131 , \ks1_col_reg[23]/NET0131 , \ks1_col_reg[24]/NET0131 , \ks1_col_reg[25]/NET0131 , \ks1_col_reg[26]/NET0131 , \ks1_col_reg[27]/NET0131 , \ks1_col_reg[28]/NET0131 , \ks1_col_reg[29]/NET0131 , \ks1_col_reg[2]/NET0131 , \ks1_col_reg[30]/NET0131 , \ks1_col_reg[31]/NET0131 , \ks1_col_reg[3]/NET0131 , \ks1_col_reg[4]/NET0131 , \ks1_col_reg[5]/NET0131 , \ks1_col_reg[6]/NET0131 , \ks1_col_reg[7]/NET0131 , \ks1_key_reg_reg[0]/NET0131 , \ks1_key_reg_reg[100]/NET0131 , \ks1_key_reg_reg[101]/NET0131 , \ks1_key_reg_reg[102]/NET0131 , \ks1_key_reg_reg[103]/NET0131 , \ks1_key_reg_reg[104]/NET0131 , \ks1_key_reg_reg[105]/NET0131 , \ks1_key_reg_reg[106]/NET0131 , \ks1_key_reg_reg[107]/NET0131 , \ks1_key_reg_reg[108]/NET0131 , \ks1_key_reg_reg[109]/P0002 , \ks1_key_reg_reg[10]/NET0131 , \ks1_key_reg_reg[110]/P0002 , \ks1_key_reg_reg[111]/NET0131 , \ks1_key_reg_reg[112]/NET0131 , \ks1_key_reg_reg[113]/NET0131 , \ks1_key_reg_reg[114]/NET0131 , \ks1_key_reg_reg[115]/NET0131 , \ks1_key_reg_reg[116]/NET0131 , \ks1_key_reg_reg[117]/NET0131 , \ks1_key_reg_reg[118]/NET0131 , \ks1_key_reg_reg[119]/NET0131 , \ks1_key_reg_reg[11]/NET0131 , \ks1_key_reg_reg[120]/NET0131 , \ks1_key_reg_reg[121]/NET0131 , \ks1_key_reg_reg[122]/NET0131 , \ks1_key_reg_reg[123]/NET0131 , \ks1_key_reg_reg[124]/NET0131 , \ks1_key_reg_reg[125]/NET0131 , \ks1_key_reg_reg[126]/NET0131 , \ks1_key_reg_reg[127]/NET0131 , \ks1_key_reg_reg[12]/NET0131 , \ks1_key_reg_reg[13]/NET0131 , \ks1_key_reg_reg[14]/NET0131 , \ks1_key_reg_reg[15]/NET0131 , \ks1_key_reg_reg[16]/NET0131 , \ks1_key_reg_reg[17]/NET0131 , \ks1_key_reg_reg[18]/NET0131 , \ks1_key_reg_reg[19]/NET0131 , \ks1_key_reg_reg[1]/NET0131 , \ks1_key_reg_reg[20]/NET0131 , \ks1_key_reg_reg[21]/NET0131 , \ks1_key_reg_reg[22]/NET0131 , \ks1_key_reg_reg[23]/NET0131 , \ks1_key_reg_reg[24]/NET0131 , \ks1_key_reg_reg[25]/NET0131 , \ks1_key_reg_reg[26]/NET0131 , \ks1_key_reg_reg[27]/NET0131 , \ks1_key_reg_reg[28]/NET0131 , \ks1_key_reg_reg[29]/NET0131 , \ks1_key_reg_reg[2]/NET0131 , \ks1_key_reg_reg[30]/NET0131 , \ks1_key_reg_reg[31]/NET0131 , \ks1_key_reg_reg[32]/NET0131 , \ks1_key_reg_reg[33]/NET0131 , \ks1_key_reg_reg[34]/NET0131 , \ks1_key_reg_reg[35]/NET0131 , \ks1_key_reg_reg[36]/NET0131 , \ks1_key_reg_reg[37]/NET0131 , \ks1_key_reg_reg[38]/NET0131 , \ks1_key_reg_reg[39]/NET0131 , \ks1_key_reg_reg[3]/NET0131 , \ks1_key_reg_reg[40]/P0002 , \ks1_key_reg_reg[41]/P0002 , \ks1_key_reg_reg[42]/P0002 , \ks1_key_reg_reg[43]/P0002 , \ks1_key_reg_reg[44]/P0002 , \ks1_key_reg_reg[45]/P0002 , \ks1_key_reg_reg[46]/P0002 , \ks1_key_reg_reg[47]/P0002 , \ks1_key_reg_reg[48]/NET0131 , \ks1_key_reg_reg[49]/NET0131 , \ks1_key_reg_reg[4]/NET0131 , \ks1_key_reg_reg[50]/NET0131 , \ks1_key_reg_reg[51]/NET0131 , \ks1_key_reg_reg[52]/NET0131 , \ks1_key_reg_reg[53]/NET0131 , \ks1_key_reg_reg[54]/NET0131 , \ks1_key_reg_reg[55]/NET0131 , \ks1_key_reg_reg[56]/NET0131 , \ks1_key_reg_reg[57]/NET0131 , \ks1_key_reg_reg[58]/NET0131 , \ks1_key_reg_reg[59]/NET0131 , \ks1_key_reg_reg[5]/NET0131 , \ks1_key_reg_reg[60]/NET0131 , \ks1_key_reg_reg[61]/NET0131 , \ks1_key_reg_reg[62]/NET0131 , \ks1_key_reg_reg[63]/NET0131 , \ks1_key_reg_reg[64]/NET0131 , \ks1_key_reg_reg[65]/NET0131 , \ks1_key_reg_reg[66]/NET0131 , \ks1_key_reg_reg[67]/NET0131 , \ks1_key_reg_reg[68]/NET0131 , \ks1_key_reg_reg[69]/NET0131 , \ks1_key_reg_reg[6]/NET0131 , \ks1_key_reg_reg[70]/NET0131 , \ks1_key_reg_reg[71]/NET0131 , \ks1_key_reg_reg[72]/P0002 , \ks1_key_reg_reg[73]/NET0131 , \ks1_key_reg_reg[74]/NET0131 , \ks1_key_reg_reg[75]/P0002 , \ks1_key_reg_reg[76]/P0002 , \ks1_key_reg_reg[77]/P0002 , \ks1_key_reg_reg[78]/P0002 , \ks1_key_reg_reg[79]/P0002 , \ks1_key_reg_reg[7]/NET0131 , \ks1_key_reg_reg[80]/NET0131 , \ks1_key_reg_reg[81]/NET0131 , \ks1_key_reg_reg[82]/NET0131 , \ks1_key_reg_reg[83]/NET0131 , \ks1_key_reg_reg[84]/NET0131 , \ks1_key_reg_reg[85]/NET0131 , \ks1_key_reg_reg[86]/NET0131 , \ks1_key_reg_reg[87]/NET0131 , \ks1_key_reg_reg[88]/NET0131 , \ks1_key_reg_reg[89]/NET0131 , \ks1_key_reg_reg[8]/NET0131 , \ks1_key_reg_reg[90]/NET0131 , \ks1_key_reg_reg[91]/NET0131 , \ks1_key_reg_reg[92]/NET0131 , \ks1_key_reg_reg[93]/NET0131 , \ks1_key_reg_reg[94]/NET0131 , \ks1_key_reg_reg[95]/NET0131 , \ks1_key_reg_reg[96]/NET0131 , \ks1_key_reg_reg[97]/NET0131 , \ks1_key_reg_reg[98]/NET0131 , \ks1_key_reg_reg[99]/NET0131 , \ks1_key_reg_reg[9]/NET0131 , \ks1_ready_o_reg/NET0131 , \ks1_state_reg[0]/NET0131 , \ks1_state_reg[1]/NET0131 , \ks1_state_reg[2]/NET0131 , load_i_pad, \mix1_data_o_reg_reg[0]/NET0131 , \mix1_data_o_reg_reg[100]/NET0131 , \mix1_data_o_reg_reg[101]/NET0131 , \mix1_data_o_reg_reg[102]/NET0131 , \mix1_data_o_reg_reg[103]/NET0131 , \mix1_data_o_reg_reg[104]/NET0131 , \mix1_data_o_reg_reg[105]/NET0131 , \mix1_data_o_reg_reg[106]/NET0131 , \mix1_data_o_reg_reg[107]/NET0131 , \mix1_data_o_reg_reg[108]/NET0131 , \mix1_data_o_reg_reg[109]/NET0131 , \mix1_data_o_reg_reg[10]/NET0131 , \mix1_data_o_reg_reg[110]/NET0131 , \mix1_data_o_reg_reg[111]/NET0131 , \mix1_data_o_reg_reg[112]/NET0131 , \mix1_data_o_reg_reg[113]/NET0131 , \mix1_data_o_reg_reg[114]/NET0131 , \mix1_data_o_reg_reg[115]/NET0131 , \mix1_data_o_reg_reg[116]/NET0131 , \mix1_data_o_reg_reg[117]/NET0131 , \mix1_data_o_reg_reg[118]/NET0131 , \mix1_data_o_reg_reg[119]/NET0131 , \mix1_data_o_reg_reg[11]/NET0131 , \mix1_data_o_reg_reg[120]/NET0131 , \mix1_data_o_reg_reg[121]/NET0131 , \mix1_data_o_reg_reg[122]/NET0131 , \mix1_data_o_reg_reg[123]/NET0131 , \mix1_data_o_reg_reg[124]/NET0131 , \mix1_data_o_reg_reg[125]/NET0131 , \mix1_data_o_reg_reg[126]/NET0131 , \mix1_data_o_reg_reg[127]/NET0131 , \mix1_data_o_reg_reg[12]/NET0131 , \mix1_data_o_reg_reg[13]/NET0131 , \mix1_data_o_reg_reg[14]/NET0131 , \mix1_data_o_reg_reg[15]/NET0131 , \mix1_data_o_reg_reg[16]/NET0131 , \mix1_data_o_reg_reg[17]/NET0131 , \mix1_data_o_reg_reg[18]/NET0131 , \mix1_data_o_reg_reg[19]/NET0131 , \mix1_data_o_reg_reg[1]/NET0131 , \mix1_data_o_reg_reg[20]/NET0131 , \mix1_data_o_reg_reg[21]/NET0131 , \mix1_data_o_reg_reg[22]/NET0131 , \mix1_data_o_reg_reg[23]/NET0131 , \mix1_data_o_reg_reg[24]/NET0131 , \mix1_data_o_reg_reg[25]/NET0131 , \mix1_data_o_reg_reg[26]/NET0131 , \mix1_data_o_reg_reg[27]/NET0131 , \mix1_data_o_reg_reg[28]/NET0131 , \mix1_data_o_reg_reg[29]/NET0131 , \mix1_data_o_reg_reg[2]/NET0131 , \mix1_data_o_reg_reg[30]/NET0131 , \mix1_data_o_reg_reg[31]/NET0131 , \mix1_data_o_reg_reg[32]/NET0131 , \mix1_data_o_reg_reg[33]/NET0131 , \mix1_data_o_reg_reg[34]/NET0131 , \mix1_data_o_reg_reg[35]/NET0131 , \mix1_data_o_reg_reg[36]/NET0131 , \mix1_data_o_reg_reg[37]/NET0131 , \mix1_data_o_reg_reg[38]/NET0131 , \mix1_data_o_reg_reg[39]/NET0131 , \mix1_data_o_reg_reg[3]/NET0131 , \mix1_data_o_reg_reg[40]/NET0131 , \mix1_data_o_reg_reg[41]/NET0131 , \mix1_data_o_reg_reg[42]/NET0131 , \mix1_data_o_reg_reg[43]/NET0131 , \mix1_data_o_reg_reg[44]/NET0131 , \mix1_data_o_reg_reg[45]/NET0131 , \mix1_data_o_reg_reg[46]/NET0131 , \mix1_data_o_reg_reg[47]/NET0131 , \mix1_data_o_reg_reg[48]/NET0131 , \mix1_data_o_reg_reg[49]/NET0131 , \mix1_data_o_reg_reg[4]/NET0131 , \mix1_data_o_reg_reg[50]/NET0131 , \mix1_data_o_reg_reg[51]/NET0131 , \mix1_data_o_reg_reg[52]/NET0131 , \mix1_data_o_reg_reg[53]/NET0131 , \mix1_data_o_reg_reg[54]/NET0131 , \mix1_data_o_reg_reg[55]/NET0131 , \mix1_data_o_reg_reg[56]/NET0131 , \mix1_data_o_reg_reg[57]/NET0131 , \mix1_data_o_reg_reg[58]/NET0131 , \mix1_data_o_reg_reg[59]/NET0131 , \mix1_data_o_reg_reg[5]/NET0131 , \mix1_data_o_reg_reg[60]/NET0131 , \mix1_data_o_reg_reg[61]/NET0131 , \mix1_data_o_reg_reg[62]/NET0131 , \mix1_data_o_reg_reg[63]/NET0131 , \mix1_data_o_reg_reg[64]/NET0131 , \mix1_data_o_reg_reg[65]/NET0131 , \mix1_data_o_reg_reg[66]/NET0131 , \mix1_data_o_reg_reg[67]/NET0131 , \mix1_data_o_reg_reg[68]/NET0131 , \mix1_data_o_reg_reg[69]/NET0131 , \mix1_data_o_reg_reg[6]/NET0131 , \mix1_data_o_reg_reg[70]/NET0131 , \mix1_data_o_reg_reg[71]/NET0131 , \mix1_data_o_reg_reg[72]/NET0131 , \mix1_data_o_reg_reg[73]/NET0131 , \mix1_data_o_reg_reg[74]/NET0131 , \mix1_data_o_reg_reg[75]/NET0131 , \mix1_data_o_reg_reg[76]/NET0131 , \mix1_data_o_reg_reg[77]/NET0131 , \mix1_data_o_reg_reg[78]/NET0131 , \mix1_data_o_reg_reg[79]/NET0131 , \mix1_data_o_reg_reg[7]/NET0131 , \mix1_data_o_reg_reg[80]/NET0131 , \mix1_data_o_reg_reg[81]/NET0131 , \mix1_data_o_reg_reg[82]/NET0131 , \mix1_data_o_reg_reg[83]/NET0131 , \mix1_data_o_reg_reg[84]/NET0131 , \mix1_data_o_reg_reg[85]/NET0131 , \mix1_data_o_reg_reg[86]/NET0131 , \mix1_data_o_reg_reg[87]/NET0131 , \mix1_data_o_reg_reg[88]/NET0131 , \mix1_data_o_reg_reg[89]/NET0131 , \mix1_data_o_reg_reg[8]/NET0131 , \mix1_data_o_reg_reg[90]/NET0131 , \mix1_data_o_reg_reg[91]/NET0131 , \mix1_data_o_reg_reg[92]/NET0131 , \mix1_data_o_reg_reg[93]/NET0131 , \mix1_data_o_reg_reg[94]/NET0131 , \mix1_data_o_reg_reg[95]/NET0131 , \mix1_data_o_reg_reg[96]/NET0131 , \mix1_data_o_reg_reg[97]/NET0131 , \mix1_data_o_reg_reg[98]/NET0131 , \mix1_data_o_reg_reg[99]/NET0131 , \mix1_data_o_reg_reg[9]/NET0131 , \mix1_data_reg_reg[100]/NET0131 , \mix1_data_reg_reg[101]/NET0131 , \mix1_data_reg_reg[102]/NET0131 , \mix1_data_reg_reg[103]/NET0131 , \mix1_data_reg_reg[104]/NET0131 , \mix1_data_reg_reg[105]/NET0131 , \mix1_data_reg_reg[106]/NET0131 , \mix1_data_reg_reg[107]/NET0131 , \mix1_data_reg_reg[108]/NET0131 , \mix1_data_reg_reg[109]/NET0131 , \mix1_data_reg_reg[110]/NET0131 , \mix1_data_reg_reg[111]/NET0131 , \mix1_data_reg_reg[112]/NET0131 , \mix1_data_reg_reg[113]/NET0131 , \mix1_data_reg_reg[114]/NET0131 , \mix1_data_reg_reg[115]/NET0131 , \mix1_data_reg_reg[116]/NET0131 , \mix1_data_reg_reg[117]/NET0131 , \mix1_data_reg_reg[118]/NET0131 , \mix1_data_reg_reg[119]/NET0131 , \mix1_data_reg_reg[120]/NET0131 , \mix1_data_reg_reg[121]/NET0131 , \mix1_data_reg_reg[122]/NET0131 , \mix1_data_reg_reg[123]/NET0131 , \mix1_data_reg_reg[124]/NET0131 , \mix1_data_reg_reg[125]/NET0131 , \mix1_data_reg_reg[126]/NET0131 , \mix1_data_reg_reg[127]/NET0131 , \mix1_data_reg_reg[32]/NET0131 , \mix1_data_reg_reg[33]/NET0131 , \mix1_data_reg_reg[34]/NET0131 , \mix1_data_reg_reg[35]/NET0131 , \mix1_data_reg_reg[36]/NET0131 , \mix1_data_reg_reg[37]/NET0131 , \mix1_data_reg_reg[38]/NET0131 , \mix1_data_reg_reg[39]/NET0131 , \mix1_data_reg_reg[40]/NET0131 , \mix1_data_reg_reg[41]/NET0131 , \mix1_data_reg_reg[42]/NET0131 , \mix1_data_reg_reg[43]/NET0131 , \mix1_data_reg_reg[44]/NET0131 , \mix1_data_reg_reg[45]/NET0131 , \mix1_data_reg_reg[46]/NET0131 , \mix1_data_reg_reg[47]/NET0131 , \mix1_data_reg_reg[48]/NET0131 , \mix1_data_reg_reg[49]/NET0131 , \mix1_data_reg_reg[50]/NET0131 , \mix1_data_reg_reg[51]/NET0131 , \mix1_data_reg_reg[52]/NET0131 , \mix1_data_reg_reg[53]/NET0131 , \mix1_data_reg_reg[54]/NET0131 , \mix1_data_reg_reg[55]/NET0131 , \mix1_data_reg_reg[56]/NET0131 , \mix1_data_reg_reg[57]/NET0131 , \mix1_data_reg_reg[58]/NET0131 , \mix1_data_reg_reg[59]/NET0131 , \mix1_data_reg_reg[60]/NET0131 , \mix1_data_reg_reg[61]/NET0131 , \mix1_data_reg_reg[62]/NET0131 , \mix1_data_reg_reg[63]/NET0131 , \mix1_data_reg_reg[64]/NET0131 , \mix1_data_reg_reg[65]/NET0131 , \mix1_data_reg_reg[66]/NET0131 , \mix1_data_reg_reg[67]/NET0131 , \mix1_data_reg_reg[68]/NET0131 , \mix1_data_reg_reg[69]/NET0131 , \mix1_data_reg_reg[70]/NET0131 , \mix1_data_reg_reg[71]/NET0131 , \mix1_data_reg_reg[72]/NET0131 , \mix1_data_reg_reg[73]/NET0131 , \mix1_data_reg_reg[74]/NET0131 , \mix1_data_reg_reg[75]/NET0131 , \mix1_data_reg_reg[76]/NET0131 , \mix1_data_reg_reg[77]/NET0131 , \mix1_data_reg_reg[78]/NET0131 , \mix1_data_reg_reg[79]/NET0131 , \mix1_data_reg_reg[80]/NET0131 , \mix1_data_reg_reg[81]/NET0131 , \mix1_data_reg_reg[82]/NET0131 , \mix1_data_reg_reg[83]/NET0131 , \mix1_data_reg_reg[84]/NET0131 , \mix1_data_reg_reg[85]/NET0131 , \mix1_data_reg_reg[86]/NET0131 , \mix1_data_reg_reg[87]/NET0131 , \mix1_data_reg_reg[88]/NET0131 , \mix1_data_reg_reg[89]/NET0131 , \mix1_data_reg_reg[90]/NET0131 , \mix1_data_reg_reg[91]/NET0131 , \mix1_data_reg_reg[92]/NET0131 , \mix1_data_reg_reg[93]/NET0131 , \mix1_data_reg_reg[94]/NET0131 , \mix1_data_reg_reg[95]/NET0131 , \mix1_data_reg_reg[96]/NET0131 , \mix1_data_reg_reg[97]/NET0131 , \mix1_data_reg_reg[98]/NET0131 , \mix1_data_reg_reg[99]/NET0131 , \mix1_ready_o_reg/NET0131 , \mix1_state_reg[0]/NET0131 , \mix1_state_reg[1]/NET0131 , \round_reg[0]/NET0131 , \round_reg[1]/NET0131 , \round_reg[2]/NET0131 , \round_reg[3]/NET0131 , \sbox1_ah_reg_reg[0]/NET0131 , \sbox1_ah_reg_reg[1]/NET0131 , \sbox1_ah_reg_reg[2]/NET0131 , \sbox1_ah_reg_reg[3]/NET0131 , \sbox1_alph_reg[0]/NET0131 , \sbox1_alph_reg[1]/NET0131 , \sbox1_alph_reg[2]/NET0131 , \sbox1_alph_reg[3]/NET0131 , \sbox1_to_invert_reg[0]/NET0131 , \sbox1_to_invert_reg[1]/NET0131 , \sbox1_to_invert_reg[2]/NET0131 , \sbox1_to_invert_reg[3]/NET0131 , \state_reg/NET0131 , \sub1_data_reg_reg[0]/NET0131 , \sub1_data_reg_reg[100]/NET0131 , \sub1_data_reg_reg[101]/NET0131 , \sub1_data_reg_reg[102]/NET0131 , \sub1_data_reg_reg[103]/NET0131 , \sub1_data_reg_reg[104]/NET0131 , \sub1_data_reg_reg[105]/NET0131 , \sub1_data_reg_reg[106]/NET0131 , \sub1_data_reg_reg[107]/NET0131 , \sub1_data_reg_reg[108]/NET0131 , \sub1_data_reg_reg[109]/NET0131 , \sub1_data_reg_reg[10]/NET0131 , \sub1_data_reg_reg[110]/NET0131 , \sub1_data_reg_reg[111]/NET0131 , \sub1_data_reg_reg[112]/NET0131 , \sub1_data_reg_reg[113]/NET0131 , \sub1_data_reg_reg[114]/NET0131 , \sub1_data_reg_reg[115]/NET0131 , \sub1_data_reg_reg[116]/NET0131 , \sub1_data_reg_reg[117]/NET0131 , \sub1_data_reg_reg[118]/NET0131 , \sub1_data_reg_reg[119]/NET0131 , \sub1_data_reg_reg[11]/NET0131 , \sub1_data_reg_reg[120]/NET0131 , \sub1_data_reg_reg[121]/NET0131 , \sub1_data_reg_reg[122]/NET0131 , \sub1_data_reg_reg[123]/NET0131 , \sub1_data_reg_reg[124]/NET0131 , \sub1_data_reg_reg[125]/NET0131 , \sub1_data_reg_reg[126]/NET0131 , \sub1_data_reg_reg[127]/NET0131 , \sub1_data_reg_reg[12]/NET0131 , \sub1_data_reg_reg[13]/NET0131 , \sub1_data_reg_reg[14]/NET0131 , \sub1_data_reg_reg[15]/NET0131 , \sub1_data_reg_reg[16]/NET0131 , \sub1_data_reg_reg[17]/NET0131 , \sub1_data_reg_reg[18]/NET0131 , \sub1_data_reg_reg[19]/NET0131 , \sub1_data_reg_reg[1]/NET0131 , \sub1_data_reg_reg[20]/NET0131 , \sub1_data_reg_reg[21]/NET0131 , \sub1_data_reg_reg[22]/NET0131 , \sub1_data_reg_reg[23]/NET0131 , \sub1_data_reg_reg[24]/NET0131 , \sub1_data_reg_reg[25]/NET0131 , \sub1_data_reg_reg[26]/NET0131 , \sub1_data_reg_reg[27]/NET0131 , \sub1_data_reg_reg[28]/NET0131 , \sub1_data_reg_reg[29]/NET0131 , \sub1_data_reg_reg[2]/NET0131 , \sub1_data_reg_reg[30]/NET0131 , \sub1_data_reg_reg[31]/NET0131 , \sub1_data_reg_reg[32]/NET0131 , \sub1_data_reg_reg[33]/NET0131 , \sub1_data_reg_reg[34]/NET0131 , \sub1_data_reg_reg[35]/NET0131 , \sub1_data_reg_reg[36]/NET0131 , \sub1_data_reg_reg[37]/NET0131 , \sub1_data_reg_reg[38]/NET0131 , \sub1_data_reg_reg[39]/NET0131 , \sub1_data_reg_reg[3]/NET0131 , \sub1_data_reg_reg[40]/NET0131 , \sub1_data_reg_reg[41]/NET0131 , \sub1_data_reg_reg[42]/NET0131 , \sub1_data_reg_reg[43]/NET0131 , \sub1_data_reg_reg[44]/NET0131 , \sub1_data_reg_reg[45]/NET0131 , \sub1_data_reg_reg[46]/NET0131 , \sub1_data_reg_reg[47]/NET0131 , \sub1_data_reg_reg[48]/NET0131 , \sub1_data_reg_reg[49]/NET0131 , \sub1_data_reg_reg[4]/NET0131 , \sub1_data_reg_reg[50]/NET0131 , \sub1_data_reg_reg[51]/NET0131 , \sub1_data_reg_reg[52]/NET0131 , \sub1_data_reg_reg[53]/NET0131 , \sub1_data_reg_reg[54]/NET0131 , \sub1_data_reg_reg[55]/NET0131 , \sub1_data_reg_reg[56]/NET0131 , \sub1_data_reg_reg[57]/NET0131 , \sub1_data_reg_reg[58]/NET0131 , \sub1_data_reg_reg[59]/NET0131 , \sub1_data_reg_reg[5]/NET0131 , \sub1_data_reg_reg[60]/NET0131 , \sub1_data_reg_reg[61]/NET0131 , \sub1_data_reg_reg[62]/NET0131 , \sub1_data_reg_reg[63]/NET0131 , \sub1_data_reg_reg[64]/NET0131 , \sub1_data_reg_reg[65]/NET0131 , \sub1_data_reg_reg[66]/NET0131 , \sub1_data_reg_reg[67]/NET0131 , \sub1_data_reg_reg[68]/NET0131 , \sub1_data_reg_reg[69]/NET0131 , \sub1_data_reg_reg[6]/NET0131 , \sub1_data_reg_reg[70]/NET0131 , \sub1_data_reg_reg[71]/NET0131 , \sub1_data_reg_reg[72]/NET0131 , \sub1_data_reg_reg[73]/NET0131 , \sub1_data_reg_reg[74]/NET0131 , \sub1_data_reg_reg[75]/NET0131 , \sub1_data_reg_reg[76]/NET0131 , \sub1_data_reg_reg[77]/NET0131 , \sub1_data_reg_reg[78]/NET0131 , \sub1_data_reg_reg[79]/NET0131 , \sub1_data_reg_reg[7]/NET0131 , \sub1_data_reg_reg[80]/NET0131 , \sub1_data_reg_reg[81]/NET0131 , \sub1_data_reg_reg[82]/NET0131 , \sub1_data_reg_reg[83]/NET0131 , \sub1_data_reg_reg[84]/NET0131 , \sub1_data_reg_reg[85]/NET0131 , \sub1_data_reg_reg[86]/NET0131 , \sub1_data_reg_reg[87]/NET0131 , \sub1_data_reg_reg[88]/NET0131 , \sub1_data_reg_reg[89]/NET0131 , \sub1_data_reg_reg[8]/NET0131 , \sub1_data_reg_reg[90]/NET0131 , \sub1_data_reg_reg[91]/NET0131 , \sub1_data_reg_reg[92]/NET0131 , \sub1_data_reg_reg[93]/NET0131 , \sub1_data_reg_reg[94]/NET0131 , \sub1_data_reg_reg[95]/NET0131 , \sub1_data_reg_reg[96]/NET0131 , \sub1_data_reg_reg[97]/NET0131 , \sub1_data_reg_reg[98]/NET0131 , \sub1_data_reg_reg[99]/NET0131 , \sub1_data_reg_reg[9]/NET0131 , \sub1_ready_o_reg/NET0131 , \sub1_state_reg[0]/NET0131 , \sub1_state_reg[1]/NET0131 , \sub1_state_reg[2]/NET0131 , \sub1_state_reg[3]/NET0131 , \sub1_state_reg[4]/NET0131 , \_al_n0 , \_al_n1 , \g27929/_0_ , \g27942/_3_ , \g27943/_3_ , \g27944/_3_ , \g27945/_0_ , \g27995/_0_ , \g27998/_0_ , \g28019/_0_ , \g28020/_0_ , \g28021/_0_ , \g28022/_0_ , \g28023/_0_ , \g28024/_0_ , \g28025/_0_ , \g28026/_0_ , \g28027/_0_ , \g28028/_0_ , \g28029/_0_ , \g28030/_0_ , \g28031/_0_ , \g28032/_0_ , \g28033/_0_ , \g28034/_0_ , \g28044/_0_ , \g28045/_0_ , \g28046/_0_ , \g28047/_0_ , \g28048/_0_ , \g28049/_0_ , \g28050/_0_ , \g28051/_0_ , \g28151/_0_ , \g28177/_0_ , \g28178/_0_ , \g28179/_0_ , \g28180/_0_ , \g28181/_0_ , \g28182/_0_ , \g28183/_0_ , \g28184/_0_ , \g28185/_0_ , \g28186/_0_ , \g28187/_0_ , \g28188/_0_ , \g28189/_0_ , \g28190/_0_ , \g28191/_0_ , \g28192/_0_ , \g28193/_0_ , \g28194/_0_ , \g28195/_0_ , \g28196/_0_ , \g28197/_0_ , \g28198/_0_ , \g28199/_0_ , \g28200/_0_ , \g28201/_0_ , \g28202/_0_ , \g28203/_0_ , \g28253/_0_ , \g28254/_0_ , \g28255/_0_ , \g28256/_0_ , \g28257/_0_ , \g28258/_0_ , \g28259/_0_ , \g28260/_0_ , \g28261/_0_ , \g28262/_0_ , \g28263/_0_ , \g28264/_0_ , \g28265/_0_ , \g28266/_0_ , \g28267/_0_ , \g28268/_0_ , \g28269/_0_ , \g28270/_0_ , \g28271/_0_ , \g28272/_0_ , \g28273/_0_ , \g28274/_0_ , \g28275/_0_ , \g28276/_0_ , \g28277/_0_ , \g28278/_0_ , \g28279/_0_ , \g28384/_2_ , \g28385/_2_ , \g28388/_2_ , \g28389/_2_ , \g28394/_2_ , \g28395/_2_ , \g28401/_2_ , \g28402/_2_ , \g28403/_0_ , \g28404/_0_ , \g28408/_0_ , \g28410/_0_ , \g28440/_0_ , \g28441/_0_ , \g28442/_0_ , \g28443/_0_ , \g28444/_0_ , \g28445/_0_ , \g28446/_0_ , \g28447/_0_ , \g28448/_0_ , \g28449/_0_ , \g28450/_0_ , \g28451/_0_ , \g28452/_0_ , \g28453/_0_ , \g28538/_0_ , \g28539/_0_ , \g28540/_0_ , \g28541/_0_ , \g28542/_0_ , \g28543/_0_ , \g28544/_0_ , \g28545/_0_ , \g28546/_0_ , \g28547/_0_ , \g28548/_0_ , \g28549/_0_ , \g28550/_0_ , \g28551/_0_ , \g28552/_0_ , \g28557/_0_ , \g28558/_0_ , \g28563/_0_ , \g28564/_0_ , \g28565/_0_ , \g28566/_0_ , \g28567/_0_ , \g28625/_2_ , \g28626/_2_ , \g28633/_2_ , \g28639/_2_ , \g28655/_2_ , \g28656/_2_ , \g28657/_2_ , \g28660/_2_ , \g28661/_2_ , \g28662/_2_ , \g28666/_2_ , \g28667/_2_ , \g28668/_2_ , \g28678/_2_ , \g28679/_2_ , \g28680/_2_ , \g28690/_0_ , \g28710/_0_ , \g28716/_0_ , \g28795/_0_ , \g28796/_0_ , \g28798/_0_ , \g28799/_0_ , \g28800/_0_ , \g28801/_0_ , \g28804/_0_ , \g28825/_2_ , \g28826/_2_ , \g28830/_2_ , \g28834/_2_ , \g28842/_2_ , \g28843/_2_ , \g28845/_2_ , \g28848/_2_ , \g28890/_0_ , \g28936/_0_ , \g28982/_0_ , \g29050/_0_ , \g29051/_0_ , \g29052/_0_ , \g29053/_0_ , \g29054/_0_ , \g29055/_0_ , \g29056/_0_ , \g29057/_0_ , \g29058/_0_ , \g29059/_0_ , \g29060/_0_ , \g29061/_0_ , \g29328/_0_ , \g29329/_0_ , \g29330/_0_ , \g29331/_0_ , \g29332/_0_ , \g29333/_0_ , \g29334/_0_ , \g29335/_0_ , \g29336/_0_ , \g29337/_0_ , \g29338/_0_ , \g29339/_0_ , \g29340/_0_ , \g29341/_0_ , \g29342/_0_ , \g29343/_0_ , \g29344/_0_ , \g29345/_0_ , \g29346/_0_ , \g29347/_0_ , \g29348/_0_ , \g29349/_0_ , \g29350/_0_ , \g29351/_0_ , \g29352/_0_ , \g29353/_0_ , \g29354/_0_ , \g29355/_0_ , \g29356/_0_ , \g29357/_0_ , \g29358/_0_ , \g29359/_0_ , \g29360/_0_ , \g29361/_0_ , \g29362/_0_ , \g29363/_0_ , \g29364/_0_ , \g29365/_0_ , \g29366/_0_ , \g29367/_0_ , \g29395/_0_ , \g29396/_0_ , \g29453/_0_ , \g29454/_0_ , \g29455/_0_ , \g29456/_0_ , \g29457/_0_ , \g29458/_0_ , \g29459/_0_ , \g29460/_0_ , \g29461/_0_ , \g29462/_0_ , \g29463/_0_ , \g29464/_0_ , \g29465/_0_ , \g29466/_0_ , \g29467/_0_ , \g29468/_0_ , \g29469/_0_ , \g29470/_0_ , \g29471/_0_ , \g29472/_0_ , \g29473/_0_ , \g29474/_0_ , \g29475/_0_ , \g29476/_0_ , \g29477/_0_ , \g29478/_0_ , \g29479/_0_ , \g29480/_0_ , \g29481/_0_ , \g29482/_0_ , \g29483/_0_ , \g29484/_0_ , \g29485/_0_ , \g29486/_0_ , \g29487/_0_ , \g29488/_0_ , \g29489/_0_ , \g29490/_0_ , \g29491/_0_ , \g29492/_0_ , \g29493/_0_ , \g29494/_0_ , \g29495/_0_ , \g29496/_0_ , \g29497/_0_ , \g29498/_0_ , \g29499/_0_ , \g29500/_0_ , \g29501/_0_ , \g29502/_0_ , \g29503/_0_ , \g29504/_0_ , \g29505/_0_ , \g29506/_0_ , \g29507/_0_ , \g29508/_0_ , \g29509/_0_ , \g29510/_0_ , \g29511/_0_ , \g29512/_0_ , \g29513/_0_ , \g29514/_0_ , \g29515/_0_ , \g29516/_0_ , \g29517/_0_ , \g29518/_0_ , \g29519/_0_ , \g29520/_0_ , \g29521/_0_ , \g29522/_0_ , \g29523/_0_ , \g29524/_0_ , \g29525/_0_ , \g29526/_0_ , \g29527/_0_ , \g29528/_0_ , \g29529/_0_ , \g29530/_0_ , \g29531/_0_ , \g29532/_0_ , \g29533/_0_ , \g29534/_0_ , \g29535/_0_ , \g29536/_0_ , \g29537/_0_ , \g29538/_0_ , \g29539/_0_ , \g29540/_0_ , \g29541/_0_ , \g29542/_0_ , \g29543/_0_ , \g29544/_0_ , \g29545/_0_ , \g29546/_0_ , \g29547/_0_ , \g29548/_0_ , \g29549/_0_ , \g29550/_0_ , \g29551/_0_ , \g29552/_0_ , \g29553/_0_ , \g29554/_0_ , \g29555/_0_ , \g29556/_0_ , \g29557/_0_ , \g29558/_0_ , \g29559/_0_ , \g29560/_0_ , \g29561/_0_ , \g29562/_0_ , \g29563/_0_ , \g29564/_0_ , \g29565/_0_ , \g29566/_0_ , \g29567/_0_ , \g29568/_0_ , \g29569/_0_ , \g29570/_0_ , \g29571/_0_ , \g29572/_0_ , \g29573/_0_ , \g29574/_0_ , \g29575/_0_ , \g29576/_0_ , \g29577/_0_ , \g29578/_0_ , \g29579/_0_ , \g29580/_0_ , \g29582/_0_ , \g29583/_0_ , \g29584/_0_ , \g29585/_0_ , \g29586/_0_ , \g29587/_0_ , \g29588/_0_ , \g29589/_0_ , \g29590/_0_ , \g29591/_0_ , \g29592/_0_ , \g29593/_0_ , \g29634/_0_ , \g29635/_0_ , \g29636/_0_ , \g29637/_0_ , \g29645/_0_ , \g29646/_0_ , \g29647/_0_ , \g29824/_0_ , \g29828/_0_ , \g29832/_0_ , \g29836/_0_ , \g29837/_0_ , \g29838/_0_ , \g29839/_0_ , \g29840/_0_ , \g29841/_0_ , \g29842/_0_ , \g29843/_0_ , \g29844/_0_ , \g29845/_0_ , \g29846/_0_ , \g29847/_0_ , \g29848/_0_ , \g29849/_0_ , \g29850/_0_ , \g29851/_0_ , \g29852/_0_ , \g29853/_0_ , \g29854/_0_ , \g29855/_0_ , \g29856/_0_ , \g29857/_0_ , \g29858/_0_ , \g29859/_0_ , \g29860/_0_ , \g29861/_0_ , \g29862/_0_ , \g29863/_0_ , \g29864/_0_ , \g29865/_0_ , \g29866/_0_ , \g29867/_0_ , \g29868/_0_ , \g30081/_0_ , \g30082/_0_ , \g30083/_0_ , \g30084/_0_ , \g30085/_0_ , \g30086/_0_ , \g30087/_0_ , \g30088/_0_ , \g30089/_0_ , \g30090/_0_ , \g30091/_0_ , \g30092/_0_ , \g30093/_0_ , \g30094/_0_ , \g30095/_0_ , \g30096/_0_ , \g30135/_0_ , \g30137/_0_ , \g30164/_0_ , \g30165/_0_ , \g30166/_0_ , \g30167/_0_ , \g30168/_0_ , \g30169/_0_ , \g30170/_0_ , \g30231/_0_ , \g30232/_0_ , \g30233/_0_ , \g30234/_0_ , \g30235/_0_ , \g30236/_0_ , \g30237/_0_ , \g30238/_0_ , \g30286/_0_ , \g30287/_0_ , \g30288/_0_ , \g30289/_0_ , \g30290/_0_ , \g30291/_0_ , \g30292/_0_ , \g30293/_0_ , \g30294/_0_ , \g30295/_0_ , \g30296/_0_ , \g30297/_0_ , \g30298/_0_ , \g30299/_0_ , \g30300/_0_ , \g30301/_0_ , \g30303/_0_ , \g30304/_0_ , \g30305/_0_ , \g30306/_0_ , \g30307/_0_ , \g30308/_0_ , \g30309/_0_ , \g30310/_0_ , \g30311/_0_ , \g30312/_0_ , \g30313/_0_ , \g30314/_0_ , \g30315/_0_ , \g30316/_0_ , \g30317/_0_ , \g30318/_0_ , \g30319/_0_ , \g30481/_0_ , \g30482/_0_ , \g30483/_0_ , \g30484/_0_ , \g30493/_0_ , \g30495/_0_ , \g30536/_0_ , \g30537/_0_ , \g30538/_0_ , \g30735/_0_ , \g30927/_0_ , \g30928/_0_ , \g30929/_0_ , \g30971/_0_ , \g30972/_0_ , \g30973/_0_ , \g30974/_0_ , \g31129/_0_ , \g31130/_0_ , \g31131/_0_ , \g31132/_0_ , \g31133/_0_ , \g31134/_0_ , \g31135/_0_ , \g31136/_0_ , \g31137/_0_ , \g31138/_0_ , \g31139/_0_ , \g31140/_0_ , \g31141/_0_ , \g31142/_0_ , \g31143/_0_ , \g31144/_0_ , \g31352/_0_ , \g31353/_0_ , \g31354/_0_ , \g31355/_0_ , \g31356/_0_ , \g31357/_0_ , \g31358/_0_ , \g31359/_0_ , \g31360/_0_ , \g31361/_0_ , \g31362/_0_ , \g31363/_0_ , \g31364/_0_ , \g31365/_0_ , \g31366/_0_ , \g31367/_0_ , \g31706/_0_ , \g32001/_0_ , \g32008/_0_ , \g32009/_0_ , \g32010/_0_ , \g32011/_0_ , \g32118/_0_ , \g33261/_0_ , \g33262/_0_ , \g33263/_0_ , \g33264/_0_ , \g33265/_0_ , \g33266/_0_ , \g33450/_0_ , \g33451/_0_ , \g33453/_0_ , \g33485/_0_ , \g33679/_2_ , \g34838/_2_ , \g34971/_0_ , \g34972/_0_ , \g34973/_0_ , \g34974/_0_ , \g34975/_0_ , \g34976/_0_ , \g34977/_0_ , \g34978/_0_ , \g34979/_0_ , \g34980/_0_ , \g34981/_0_ , \g34982/_0_ , \g34983/_0_ , \g34984/_0_ , \g34985/_0_ , \g34986/_0_ , \g34987/_0_ , \g34988/_0_ , \g34989/_0_ , \g34990/_0_ , \g34991/_0_ , \g34992/_0_ , \g34993/_0_ , \g34994/_0_ , \g34995/_0_ , \g34996/_0_ , \g34997/_0_ , \g34998/_0_ , \g34999/_0_ , \g35000/_0_ , \g35001/_0_ , \g35002/_0_ , \g35003/_0_ , \g35004/_0_ , \g35005/_0_ , \g35006/_0_ , \g35007/_0_ , \g35008/_0_ , \g35009/_0_ , \g35010/_0_ , \g35011/_0_ , \g35012/_0_ , \g35013/_0_ , \g35014/_0_ , \g35015/_0_ , \g35016/_0_ , \g35017/_0_ , \g35018/_0_ , \g35019/_0_ , \g35020/_0_ , \g35021/_0_ , \g35022/_0_ , \g35023/_0_ , \g35024/_0_ , \g35025/_0_ , \g35026/_0_ , \g35027/_0_ , \g35028/_0_ , \g35029/_0_ , \g35030/_0_ , \g35031/_0_ , \g35032/_0_ , \g35033/_0_ , \g35034/_0_ , \g35035/_0_ , \g35036/_0_ , \g35037/_0_ , \g35038/_0_ , \g35039/_0_ , \g35040/_0_ , \g35041/_0_ , \g35042/_0_ , \g35043/_0_ , \g35044/_0_ , \g35045/_0_ , \g35046/_0_ , \g35047/_0_ , \g35048/_0_ , \g35049/_0_ , \g35050/_0_ , \g35051/_0_ , \g35052/_0_ , \g35053/_0_ , \g35054/_0_ , \g35055/_0_ , \g35056/_0_ , \g35057/_0_ , \g35058/_0_ , \g35059/_0_ , \g35060/_0_ , \g35061/_0_ , \g35062/_0_ , \g35063/_0_ , \g35064/_0_ , \g35065/_0_ , \g35066/_0_ , \g35538/_0_ , \g35956/_0_ , \g36298/_1_ , \g36324/_0_ , \g36375/_0_ , \g38269/_0_ , \g38473/_0_ , \g38501/_0_ , \g38569/_0_ , \g38629/_0_ , \g38721_dup/_3_ , \g38735/_0_ , \g38753/_0_ , \g38849/_3_ , \g39071/_0_ , \g39073/_0_ , \g39077/_0_ , \g39080/_0_ , \g39135/_0_ , \g39138/_0_ , \g39182/_0_ , \g39197/_3_ , \g39207/_3_ , \g39241/_0_ , \g39272/_0_ , \g39307/_0_ , \g39308/_0_ , \g39361/_0_ , \g39494/_0_ , \g39558/_0_ , \g39575/_0_ , \g39583/_0_ );
	input \addroundkey_ready_o_reg/NET0131  ;
	input \addroundkey_round_reg[0]/NET0131  ;
	input \addroundkey_round_reg[1]/NET0131  ;
	input \addroundkey_round_reg[2]/NET0131  ;
	input \addroundkey_round_reg[3]/NET0131  ;
	input \addroundkey_start_i_reg/NET0131  ;
	input \data_i[0]_pad  ;
	input \data_i[100]_pad  ;
	input \data_i[101]_pad  ;
	input \data_i[102]_pad  ;
	input \data_i[103]_pad  ;
	input \data_i[104]_pad  ;
	input \data_i[105]_pad  ;
	input \data_i[106]_pad  ;
	input \data_i[107]_pad  ;
	input \data_i[108]_pad  ;
	input \data_i[109]_pad  ;
	input \data_i[10]_pad  ;
	input \data_i[110]_pad  ;
	input \data_i[111]_pad  ;
	input \data_i[112]_pad  ;
	input \data_i[113]_pad  ;
	input \data_i[114]_pad  ;
	input \data_i[115]_pad  ;
	input \data_i[116]_pad  ;
	input \data_i[117]_pad  ;
	input \data_i[118]_pad  ;
	input \data_i[119]_pad  ;
	input \data_i[11]_pad  ;
	input \data_i[120]_pad  ;
	input \data_i[121]_pad  ;
	input \data_i[122]_pad  ;
	input \data_i[123]_pad  ;
	input \data_i[124]_pad  ;
	input \data_i[125]_pad  ;
	input \data_i[126]_pad  ;
	input \data_i[127]_pad  ;
	input \data_i[12]_pad  ;
	input \data_i[13]_pad  ;
	input \data_i[14]_pad  ;
	input \data_i[15]_pad  ;
	input \data_i[16]_pad  ;
	input \data_i[17]_pad  ;
	input \data_i[18]_pad  ;
	input \data_i[19]_pad  ;
	input \data_i[1]_pad  ;
	input \data_i[20]_pad  ;
	input \data_i[21]_pad  ;
	input \data_i[22]_pad  ;
	input \data_i[23]_pad  ;
	input \data_i[24]_pad  ;
	input \data_i[25]_pad  ;
	input \data_i[26]_pad  ;
	input \data_i[27]_pad  ;
	input \data_i[28]_pad  ;
	input \data_i[29]_pad  ;
	input \data_i[2]_pad  ;
	input \data_i[30]_pad  ;
	input \data_i[31]_pad  ;
	input \data_i[32]_pad  ;
	input \data_i[33]_pad  ;
	input \data_i[34]_pad  ;
	input \data_i[35]_pad  ;
	input \data_i[36]_pad  ;
	input \data_i[37]_pad  ;
	input \data_i[38]_pad  ;
	input \data_i[39]_pad  ;
	input \data_i[3]_pad  ;
	input \data_i[40]_pad  ;
	input \data_i[41]_pad  ;
	input \data_i[42]_pad  ;
	input \data_i[43]_pad  ;
	input \data_i[44]_pad  ;
	input \data_i[45]_pad  ;
	input \data_i[46]_pad  ;
	input \data_i[47]_pad  ;
	input \data_i[48]_pad  ;
	input \data_i[49]_pad  ;
	input \data_i[4]_pad  ;
	input \data_i[50]_pad  ;
	input \data_i[51]_pad  ;
	input \data_i[52]_pad  ;
	input \data_i[53]_pad  ;
	input \data_i[54]_pad  ;
	input \data_i[55]_pad  ;
	input \data_i[56]_pad  ;
	input \data_i[57]_pad  ;
	input \data_i[58]_pad  ;
	input \data_i[59]_pad  ;
	input \data_i[5]_pad  ;
	input \data_i[60]_pad  ;
	input \data_i[61]_pad  ;
	input \data_i[62]_pad  ;
	input \data_i[63]_pad  ;
	input \data_i[64]_pad  ;
	input \data_i[65]_pad  ;
	input \data_i[66]_pad  ;
	input \data_i[67]_pad  ;
	input \data_i[68]_pad  ;
	input \data_i[69]_pad  ;
	input \data_i[6]_pad  ;
	input \data_i[70]_pad  ;
	input \data_i[71]_pad  ;
	input \data_i[72]_pad  ;
	input \data_i[73]_pad  ;
	input \data_i[74]_pad  ;
	input \data_i[75]_pad  ;
	input \data_i[76]_pad  ;
	input \data_i[77]_pad  ;
	input \data_i[78]_pad  ;
	input \data_i[79]_pad  ;
	input \data_i[7]_pad  ;
	input \data_i[80]_pad  ;
	input \data_i[81]_pad  ;
	input \data_i[82]_pad  ;
	input \data_i[83]_pad  ;
	input \data_i[84]_pad  ;
	input \data_i[85]_pad  ;
	input \data_i[86]_pad  ;
	input \data_i[87]_pad  ;
	input \data_i[88]_pad  ;
	input \data_i[89]_pad  ;
	input \data_i[8]_pad  ;
	input \data_i[90]_pad  ;
	input \data_i[91]_pad  ;
	input \data_i[92]_pad  ;
	input \data_i[93]_pad  ;
	input \data_i[94]_pad  ;
	input \data_i[95]_pad  ;
	input \data_i[96]_pad  ;
	input \data_i[97]_pad  ;
	input \data_i[98]_pad  ;
	input \data_i[99]_pad  ;
	input \data_i[9]_pad  ;
	input \data_o[0]_pad  ;
	input \data_o[100]_pad  ;
	input \data_o[101]_pad  ;
	input \data_o[102]_pad  ;
	input \data_o[103]_pad  ;
	input \data_o[104]_pad  ;
	input \data_o[105]_pad  ;
	input \data_o[106]_pad  ;
	input \data_o[107]_pad  ;
	input \data_o[108]_pad  ;
	input \data_o[109]_pad  ;
	input \data_o[10]_pad  ;
	input \data_o[110]_pad  ;
	input \data_o[111]_pad  ;
	input \data_o[112]_pad  ;
	input \data_o[113]_pad  ;
	input \data_o[114]_pad  ;
	input \data_o[115]_pad  ;
	input \data_o[116]_pad  ;
	input \data_o[117]_pad  ;
	input \data_o[118]_pad  ;
	input \data_o[119]_pad  ;
	input \data_o[11]_pad  ;
	input \data_o[120]_pad  ;
	input \data_o[121]_pad  ;
	input \data_o[122]_pad  ;
	input \data_o[123]_pad  ;
	input \data_o[124]_pad  ;
	input \data_o[125]_pad  ;
	input \data_o[126]_pad  ;
	input \data_o[127]_pad  ;
	input \data_o[12]_pad  ;
	input \data_o[13]_pad  ;
	input \data_o[14]_pad  ;
	input \data_o[15]_pad  ;
	input \data_o[16]_pad  ;
	input \data_o[17]_pad  ;
	input \data_o[18]_pad  ;
	input \data_o[19]_pad  ;
	input \data_o[1]_pad  ;
	input \data_o[20]_pad  ;
	input \data_o[21]_pad  ;
	input \data_o[22]_pad  ;
	input \data_o[23]_pad  ;
	input \data_o[24]_pad  ;
	input \data_o[25]_pad  ;
	input \data_o[26]_pad  ;
	input \data_o[27]_pad  ;
	input \data_o[28]_pad  ;
	input \data_o[29]_pad  ;
	input \data_o[2]_pad  ;
	input \data_o[30]_pad  ;
	input \data_o[31]_pad  ;
	input \data_o[32]_pad  ;
	input \data_o[33]_pad  ;
	input \data_o[34]_pad  ;
	input \data_o[35]_pad  ;
	input \data_o[36]_pad  ;
	input \data_o[37]_pad  ;
	input \data_o[38]_pad  ;
	input \data_o[39]_pad  ;
	input \data_o[3]_pad  ;
	input \data_o[40]_pad  ;
	input \data_o[41]_pad  ;
	input \data_o[42]_pad  ;
	input \data_o[43]_pad  ;
	input \data_o[44]_pad  ;
	input \data_o[45]_pad  ;
	input \data_o[46]_pad  ;
	input \data_o[47]_pad  ;
	input \data_o[48]_pad  ;
	input \data_o[49]_pad  ;
	input \data_o[4]_pad  ;
	input \data_o[50]_pad  ;
	input \data_o[51]_pad  ;
	input \data_o[52]_pad  ;
	input \data_o[53]_pad  ;
	input \data_o[54]_pad  ;
	input \data_o[55]_pad  ;
	input \data_o[56]_pad  ;
	input \data_o[57]_pad  ;
	input \data_o[58]_pad  ;
	input \data_o[59]_pad  ;
	input \data_o[5]_pad  ;
	input \data_o[60]_pad  ;
	input \data_o[61]_pad  ;
	input \data_o[62]_pad  ;
	input \data_o[63]_pad  ;
	input \data_o[64]_pad  ;
	input \data_o[65]_pad  ;
	input \data_o[66]_pad  ;
	input \data_o[67]_pad  ;
	input \data_o[68]_pad  ;
	input \data_o[69]_pad  ;
	input \data_o[6]_pad  ;
	input \data_o[70]_pad  ;
	input \data_o[71]_pad  ;
	input \data_o[72]_pad  ;
	input \data_o[73]_pad  ;
	input \data_o[74]_pad  ;
	input \data_o[75]_pad  ;
	input \data_o[76]_pad  ;
	input \data_o[77]_pad  ;
	input \data_o[78]_pad  ;
	input \data_o[79]_pad  ;
	input \data_o[7]_pad  ;
	input \data_o[80]_pad  ;
	input \data_o[81]_pad  ;
	input \data_o[82]_pad  ;
	input \data_o[83]_pad  ;
	input \data_o[84]_pad  ;
	input \data_o[85]_pad  ;
	input \data_o[86]_pad  ;
	input \data_o[87]_pad  ;
	input \data_o[88]_pad  ;
	input \data_o[89]_pad  ;
	input \data_o[8]_pad  ;
	input \data_o[90]_pad  ;
	input \data_o[91]_pad  ;
	input \data_o[92]_pad  ;
	input \data_o[93]_pad  ;
	input \data_o[94]_pad  ;
	input \data_o[95]_pad  ;
	input \data_o[96]_pad  ;
	input \data_o[97]_pad  ;
	input \data_o[98]_pad  ;
	input \data_o[99]_pad  ;
	input \data_o[9]_pad  ;
	input decrypt_i_pad ;
	input \first_round_reg_reg/NET0131  ;
	input \key_i[0]_pad  ;
	input \key_i[100]_pad  ;
	input \key_i[101]_pad  ;
	input \key_i[102]_pad  ;
	input \key_i[103]_pad  ;
	input \key_i[104]_pad  ;
	input \key_i[105]_pad  ;
	input \key_i[106]_pad  ;
	input \key_i[107]_pad  ;
	input \key_i[108]_pad  ;
	input \key_i[109]_pad  ;
	input \key_i[10]_pad  ;
	input \key_i[110]_pad  ;
	input \key_i[111]_pad  ;
	input \key_i[112]_pad  ;
	input \key_i[113]_pad  ;
	input \key_i[114]_pad  ;
	input \key_i[115]_pad  ;
	input \key_i[116]_pad  ;
	input \key_i[117]_pad  ;
	input \key_i[118]_pad  ;
	input \key_i[119]_pad  ;
	input \key_i[11]_pad  ;
	input \key_i[120]_pad  ;
	input \key_i[121]_pad  ;
	input \key_i[122]_pad  ;
	input \key_i[123]_pad  ;
	input \key_i[124]_pad  ;
	input \key_i[125]_pad  ;
	input \key_i[126]_pad  ;
	input \key_i[127]_pad  ;
	input \key_i[12]_pad  ;
	input \key_i[13]_pad  ;
	input \key_i[14]_pad  ;
	input \key_i[15]_pad  ;
	input \key_i[16]_pad  ;
	input \key_i[17]_pad  ;
	input \key_i[18]_pad  ;
	input \key_i[19]_pad  ;
	input \key_i[1]_pad  ;
	input \key_i[20]_pad  ;
	input \key_i[21]_pad  ;
	input \key_i[22]_pad  ;
	input \key_i[23]_pad  ;
	input \key_i[24]_pad  ;
	input \key_i[25]_pad  ;
	input \key_i[26]_pad  ;
	input \key_i[27]_pad  ;
	input \key_i[28]_pad  ;
	input \key_i[29]_pad  ;
	input \key_i[2]_pad  ;
	input \key_i[30]_pad  ;
	input \key_i[31]_pad  ;
	input \key_i[32]_pad  ;
	input \key_i[33]_pad  ;
	input \key_i[34]_pad  ;
	input \key_i[35]_pad  ;
	input \key_i[36]_pad  ;
	input \key_i[37]_pad  ;
	input \key_i[38]_pad  ;
	input \key_i[39]_pad  ;
	input \key_i[3]_pad  ;
	input \key_i[40]_pad  ;
	input \key_i[41]_pad  ;
	input \key_i[42]_pad  ;
	input \key_i[43]_pad  ;
	input \key_i[44]_pad  ;
	input \key_i[45]_pad  ;
	input \key_i[46]_pad  ;
	input \key_i[47]_pad  ;
	input \key_i[48]_pad  ;
	input \key_i[49]_pad  ;
	input \key_i[4]_pad  ;
	input \key_i[50]_pad  ;
	input \key_i[51]_pad  ;
	input \key_i[52]_pad  ;
	input \key_i[53]_pad  ;
	input \key_i[54]_pad  ;
	input \key_i[55]_pad  ;
	input \key_i[56]_pad  ;
	input \key_i[57]_pad  ;
	input \key_i[58]_pad  ;
	input \key_i[59]_pad  ;
	input \key_i[5]_pad  ;
	input \key_i[60]_pad  ;
	input \key_i[61]_pad  ;
	input \key_i[62]_pad  ;
	input \key_i[63]_pad  ;
	input \key_i[64]_pad  ;
	input \key_i[65]_pad  ;
	input \key_i[66]_pad  ;
	input \key_i[67]_pad  ;
	input \key_i[68]_pad  ;
	input \key_i[69]_pad  ;
	input \key_i[6]_pad  ;
	input \key_i[70]_pad  ;
	input \key_i[71]_pad  ;
	input \key_i[72]_pad  ;
	input \key_i[73]_pad  ;
	input \key_i[74]_pad  ;
	input \key_i[75]_pad  ;
	input \key_i[76]_pad  ;
	input \key_i[77]_pad  ;
	input \key_i[78]_pad  ;
	input \key_i[79]_pad  ;
	input \key_i[7]_pad  ;
	input \key_i[80]_pad  ;
	input \key_i[81]_pad  ;
	input \key_i[82]_pad  ;
	input \key_i[83]_pad  ;
	input \key_i[84]_pad  ;
	input \key_i[85]_pad  ;
	input \key_i[86]_pad  ;
	input \key_i[87]_pad  ;
	input \key_i[88]_pad  ;
	input \key_i[89]_pad  ;
	input \key_i[8]_pad  ;
	input \key_i[90]_pad  ;
	input \key_i[91]_pad  ;
	input \key_i[92]_pad  ;
	input \key_i[93]_pad  ;
	input \key_i[94]_pad  ;
	input \key_i[95]_pad  ;
	input \key_i[96]_pad  ;
	input \key_i[97]_pad  ;
	input \key_i[98]_pad  ;
	input \key_i[99]_pad  ;
	input \key_i[9]_pad  ;
	input \ks1_col_reg[0]/NET0131  ;
	input \ks1_col_reg[16]/NET0131  ;
	input \ks1_col_reg[17]/NET0131  ;
	input \ks1_col_reg[18]/NET0131  ;
	input \ks1_col_reg[19]/NET0131  ;
	input \ks1_col_reg[1]/NET0131  ;
	input \ks1_col_reg[20]/NET0131  ;
	input \ks1_col_reg[21]/NET0131  ;
	input \ks1_col_reg[22]/NET0131  ;
	input \ks1_col_reg[23]/NET0131  ;
	input \ks1_col_reg[24]/NET0131  ;
	input \ks1_col_reg[25]/NET0131  ;
	input \ks1_col_reg[26]/NET0131  ;
	input \ks1_col_reg[27]/NET0131  ;
	input \ks1_col_reg[28]/NET0131  ;
	input \ks1_col_reg[29]/NET0131  ;
	input \ks1_col_reg[2]/NET0131  ;
	input \ks1_col_reg[30]/NET0131  ;
	input \ks1_col_reg[31]/NET0131  ;
	input \ks1_col_reg[3]/NET0131  ;
	input \ks1_col_reg[4]/NET0131  ;
	input \ks1_col_reg[5]/NET0131  ;
	input \ks1_col_reg[6]/NET0131  ;
	input \ks1_col_reg[7]/NET0131  ;
	input \ks1_key_reg_reg[0]/NET0131  ;
	input \ks1_key_reg_reg[100]/NET0131  ;
	input \ks1_key_reg_reg[101]/NET0131  ;
	input \ks1_key_reg_reg[102]/NET0131  ;
	input \ks1_key_reg_reg[103]/NET0131  ;
	input \ks1_key_reg_reg[104]/NET0131  ;
	input \ks1_key_reg_reg[105]/NET0131  ;
	input \ks1_key_reg_reg[106]/NET0131  ;
	input \ks1_key_reg_reg[107]/NET0131  ;
	input \ks1_key_reg_reg[108]/NET0131  ;
	input \ks1_key_reg_reg[109]/P0002  ;
	input \ks1_key_reg_reg[10]/NET0131  ;
	input \ks1_key_reg_reg[110]/P0002  ;
	input \ks1_key_reg_reg[111]/NET0131  ;
	input \ks1_key_reg_reg[112]/NET0131  ;
	input \ks1_key_reg_reg[113]/NET0131  ;
	input \ks1_key_reg_reg[114]/NET0131  ;
	input \ks1_key_reg_reg[115]/NET0131  ;
	input \ks1_key_reg_reg[116]/NET0131  ;
	input \ks1_key_reg_reg[117]/NET0131  ;
	input \ks1_key_reg_reg[118]/NET0131  ;
	input \ks1_key_reg_reg[119]/NET0131  ;
	input \ks1_key_reg_reg[11]/NET0131  ;
	input \ks1_key_reg_reg[120]/NET0131  ;
	input \ks1_key_reg_reg[121]/NET0131  ;
	input \ks1_key_reg_reg[122]/NET0131  ;
	input \ks1_key_reg_reg[123]/NET0131  ;
	input \ks1_key_reg_reg[124]/NET0131  ;
	input \ks1_key_reg_reg[125]/NET0131  ;
	input \ks1_key_reg_reg[126]/NET0131  ;
	input \ks1_key_reg_reg[127]/NET0131  ;
	input \ks1_key_reg_reg[12]/NET0131  ;
	input \ks1_key_reg_reg[13]/NET0131  ;
	input \ks1_key_reg_reg[14]/NET0131  ;
	input \ks1_key_reg_reg[15]/NET0131  ;
	input \ks1_key_reg_reg[16]/NET0131  ;
	input \ks1_key_reg_reg[17]/NET0131  ;
	input \ks1_key_reg_reg[18]/NET0131  ;
	input \ks1_key_reg_reg[19]/NET0131  ;
	input \ks1_key_reg_reg[1]/NET0131  ;
	input \ks1_key_reg_reg[20]/NET0131  ;
	input \ks1_key_reg_reg[21]/NET0131  ;
	input \ks1_key_reg_reg[22]/NET0131  ;
	input \ks1_key_reg_reg[23]/NET0131  ;
	input \ks1_key_reg_reg[24]/NET0131  ;
	input \ks1_key_reg_reg[25]/NET0131  ;
	input \ks1_key_reg_reg[26]/NET0131  ;
	input \ks1_key_reg_reg[27]/NET0131  ;
	input \ks1_key_reg_reg[28]/NET0131  ;
	input \ks1_key_reg_reg[29]/NET0131  ;
	input \ks1_key_reg_reg[2]/NET0131  ;
	input \ks1_key_reg_reg[30]/NET0131  ;
	input \ks1_key_reg_reg[31]/NET0131  ;
	input \ks1_key_reg_reg[32]/NET0131  ;
	input \ks1_key_reg_reg[33]/NET0131  ;
	input \ks1_key_reg_reg[34]/NET0131  ;
	input \ks1_key_reg_reg[35]/NET0131  ;
	input \ks1_key_reg_reg[36]/NET0131  ;
	input \ks1_key_reg_reg[37]/NET0131  ;
	input \ks1_key_reg_reg[38]/NET0131  ;
	input \ks1_key_reg_reg[39]/NET0131  ;
	input \ks1_key_reg_reg[3]/NET0131  ;
	input \ks1_key_reg_reg[40]/P0002  ;
	input \ks1_key_reg_reg[41]/P0002  ;
	input \ks1_key_reg_reg[42]/P0002  ;
	input \ks1_key_reg_reg[43]/P0002  ;
	input \ks1_key_reg_reg[44]/P0002  ;
	input \ks1_key_reg_reg[45]/P0002  ;
	input \ks1_key_reg_reg[46]/P0002  ;
	input \ks1_key_reg_reg[47]/P0002  ;
	input \ks1_key_reg_reg[48]/NET0131  ;
	input \ks1_key_reg_reg[49]/NET0131  ;
	input \ks1_key_reg_reg[4]/NET0131  ;
	input \ks1_key_reg_reg[50]/NET0131  ;
	input \ks1_key_reg_reg[51]/NET0131  ;
	input \ks1_key_reg_reg[52]/NET0131  ;
	input \ks1_key_reg_reg[53]/NET0131  ;
	input \ks1_key_reg_reg[54]/NET0131  ;
	input \ks1_key_reg_reg[55]/NET0131  ;
	input \ks1_key_reg_reg[56]/NET0131  ;
	input \ks1_key_reg_reg[57]/NET0131  ;
	input \ks1_key_reg_reg[58]/NET0131  ;
	input \ks1_key_reg_reg[59]/NET0131  ;
	input \ks1_key_reg_reg[5]/NET0131  ;
	input \ks1_key_reg_reg[60]/NET0131  ;
	input \ks1_key_reg_reg[61]/NET0131  ;
	input \ks1_key_reg_reg[62]/NET0131  ;
	input \ks1_key_reg_reg[63]/NET0131  ;
	input \ks1_key_reg_reg[64]/NET0131  ;
	input \ks1_key_reg_reg[65]/NET0131  ;
	input \ks1_key_reg_reg[66]/NET0131  ;
	input \ks1_key_reg_reg[67]/NET0131  ;
	input \ks1_key_reg_reg[68]/NET0131  ;
	input \ks1_key_reg_reg[69]/NET0131  ;
	input \ks1_key_reg_reg[6]/NET0131  ;
	input \ks1_key_reg_reg[70]/NET0131  ;
	input \ks1_key_reg_reg[71]/NET0131  ;
	input \ks1_key_reg_reg[72]/P0002  ;
	input \ks1_key_reg_reg[73]/NET0131  ;
	input \ks1_key_reg_reg[74]/NET0131  ;
	input \ks1_key_reg_reg[75]/P0002  ;
	input \ks1_key_reg_reg[76]/P0002  ;
	input \ks1_key_reg_reg[77]/P0002  ;
	input \ks1_key_reg_reg[78]/P0002  ;
	input \ks1_key_reg_reg[79]/P0002  ;
	input \ks1_key_reg_reg[7]/NET0131  ;
	input \ks1_key_reg_reg[80]/NET0131  ;
	input \ks1_key_reg_reg[81]/NET0131  ;
	input \ks1_key_reg_reg[82]/NET0131  ;
	input \ks1_key_reg_reg[83]/NET0131  ;
	input \ks1_key_reg_reg[84]/NET0131  ;
	input \ks1_key_reg_reg[85]/NET0131  ;
	input \ks1_key_reg_reg[86]/NET0131  ;
	input \ks1_key_reg_reg[87]/NET0131  ;
	input \ks1_key_reg_reg[88]/NET0131  ;
	input \ks1_key_reg_reg[89]/NET0131  ;
	input \ks1_key_reg_reg[8]/NET0131  ;
	input \ks1_key_reg_reg[90]/NET0131  ;
	input \ks1_key_reg_reg[91]/NET0131  ;
	input \ks1_key_reg_reg[92]/NET0131  ;
	input \ks1_key_reg_reg[93]/NET0131  ;
	input \ks1_key_reg_reg[94]/NET0131  ;
	input \ks1_key_reg_reg[95]/NET0131  ;
	input \ks1_key_reg_reg[96]/NET0131  ;
	input \ks1_key_reg_reg[97]/NET0131  ;
	input \ks1_key_reg_reg[98]/NET0131  ;
	input \ks1_key_reg_reg[99]/NET0131  ;
	input \ks1_key_reg_reg[9]/NET0131  ;
	input \ks1_ready_o_reg/NET0131  ;
	input \ks1_state_reg[0]/NET0131  ;
	input \ks1_state_reg[1]/NET0131  ;
	input \ks1_state_reg[2]/NET0131  ;
	input load_i_pad ;
	input \mix1_data_o_reg_reg[0]/NET0131  ;
	input \mix1_data_o_reg_reg[100]/NET0131  ;
	input \mix1_data_o_reg_reg[101]/NET0131  ;
	input \mix1_data_o_reg_reg[102]/NET0131  ;
	input \mix1_data_o_reg_reg[103]/NET0131  ;
	input \mix1_data_o_reg_reg[104]/NET0131  ;
	input \mix1_data_o_reg_reg[105]/NET0131  ;
	input \mix1_data_o_reg_reg[106]/NET0131  ;
	input \mix1_data_o_reg_reg[107]/NET0131  ;
	input \mix1_data_o_reg_reg[108]/NET0131  ;
	input \mix1_data_o_reg_reg[109]/NET0131  ;
	input \mix1_data_o_reg_reg[10]/NET0131  ;
	input \mix1_data_o_reg_reg[110]/NET0131  ;
	input \mix1_data_o_reg_reg[111]/NET0131  ;
	input \mix1_data_o_reg_reg[112]/NET0131  ;
	input \mix1_data_o_reg_reg[113]/NET0131  ;
	input \mix1_data_o_reg_reg[114]/NET0131  ;
	input \mix1_data_o_reg_reg[115]/NET0131  ;
	input \mix1_data_o_reg_reg[116]/NET0131  ;
	input \mix1_data_o_reg_reg[117]/NET0131  ;
	input \mix1_data_o_reg_reg[118]/NET0131  ;
	input \mix1_data_o_reg_reg[119]/NET0131  ;
	input \mix1_data_o_reg_reg[11]/NET0131  ;
	input \mix1_data_o_reg_reg[120]/NET0131  ;
	input \mix1_data_o_reg_reg[121]/NET0131  ;
	input \mix1_data_o_reg_reg[122]/NET0131  ;
	input \mix1_data_o_reg_reg[123]/NET0131  ;
	input \mix1_data_o_reg_reg[124]/NET0131  ;
	input \mix1_data_o_reg_reg[125]/NET0131  ;
	input \mix1_data_o_reg_reg[126]/NET0131  ;
	input \mix1_data_o_reg_reg[127]/NET0131  ;
	input \mix1_data_o_reg_reg[12]/NET0131  ;
	input \mix1_data_o_reg_reg[13]/NET0131  ;
	input \mix1_data_o_reg_reg[14]/NET0131  ;
	input \mix1_data_o_reg_reg[15]/NET0131  ;
	input \mix1_data_o_reg_reg[16]/NET0131  ;
	input \mix1_data_o_reg_reg[17]/NET0131  ;
	input \mix1_data_o_reg_reg[18]/NET0131  ;
	input \mix1_data_o_reg_reg[19]/NET0131  ;
	input \mix1_data_o_reg_reg[1]/NET0131  ;
	input \mix1_data_o_reg_reg[20]/NET0131  ;
	input \mix1_data_o_reg_reg[21]/NET0131  ;
	input \mix1_data_o_reg_reg[22]/NET0131  ;
	input \mix1_data_o_reg_reg[23]/NET0131  ;
	input \mix1_data_o_reg_reg[24]/NET0131  ;
	input \mix1_data_o_reg_reg[25]/NET0131  ;
	input \mix1_data_o_reg_reg[26]/NET0131  ;
	input \mix1_data_o_reg_reg[27]/NET0131  ;
	input \mix1_data_o_reg_reg[28]/NET0131  ;
	input \mix1_data_o_reg_reg[29]/NET0131  ;
	input \mix1_data_o_reg_reg[2]/NET0131  ;
	input \mix1_data_o_reg_reg[30]/NET0131  ;
	input \mix1_data_o_reg_reg[31]/NET0131  ;
	input \mix1_data_o_reg_reg[32]/NET0131  ;
	input \mix1_data_o_reg_reg[33]/NET0131  ;
	input \mix1_data_o_reg_reg[34]/NET0131  ;
	input \mix1_data_o_reg_reg[35]/NET0131  ;
	input \mix1_data_o_reg_reg[36]/NET0131  ;
	input \mix1_data_o_reg_reg[37]/NET0131  ;
	input \mix1_data_o_reg_reg[38]/NET0131  ;
	input \mix1_data_o_reg_reg[39]/NET0131  ;
	input \mix1_data_o_reg_reg[3]/NET0131  ;
	input \mix1_data_o_reg_reg[40]/NET0131  ;
	input \mix1_data_o_reg_reg[41]/NET0131  ;
	input \mix1_data_o_reg_reg[42]/NET0131  ;
	input \mix1_data_o_reg_reg[43]/NET0131  ;
	input \mix1_data_o_reg_reg[44]/NET0131  ;
	input \mix1_data_o_reg_reg[45]/NET0131  ;
	input \mix1_data_o_reg_reg[46]/NET0131  ;
	input \mix1_data_o_reg_reg[47]/NET0131  ;
	input \mix1_data_o_reg_reg[48]/NET0131  ;
	input \mix1_data_o_reg_reg[49]/NET0131  ;
	input \mix1_data_o_reg_reg[4]/NET0131  ;
	input \mix1_data_o_reg_reg[50]/NET0131  ;
	input \mix1_data_o_reg_reg[51]/NET0131  ;
	input \mix1_data_o_reg_reg[52]/NET0131  ;
	input \mix1_data_o_reg_reg[53]/NET0131  ;
	input \mix1_data_o_reg_reg[54]/NET0131  ;
	input \mix1_data_o_reg_reg[55]/NET0131  ;
	input \mix1_data_o_reg_reg[56]/NET0131  ;
	input \mix1_data_o_reg_reg[57]/NET0131  ;
	input \mix1_data_o_reg_reg[58]/NET0131  ;
	input \mix1_data_o_reg_reg[59]/NET0131  ;
	input \mix1_data_o_reg_reg[5]/NET0131  ;
	input \mix1_data_o_reg_reg[60]/NET0131  ;
	input \mix1_data_o_reg_reg[61]/NET0131  ;
	input \mix1_data_o_reg_reg[62]/NET0131  ;
	input \mix1_data_o_reg_reg[63]/NET0131  ;
	input \mix1_data_o_reg_reg[64]/NET0131  ;
	input \mix1_data_o_reg_reg[65]/NET0131  ;
	input \mix1_data_o_reg_reg[66]/NET0131  ;
	input \mix1_data_o_reg_reg[67]/NET0131  ;
	input \mix1_data_o_reg_reg[68]/NET0131  ;
	input \mix1_data_o_reg_reg[69]/NET0131  ;
	input \mix1_data_o_reg_reg[6]/NET0131  ;
	input \mix1_data_o_reg_reg[70]/NET0131  ;
	input \mix1_data_o_reg_reg[71]/NET0131  ;
	input \mix1_data_o_reg_reg[72]/NET0131  ;
	input \mix1_data_o_reg_reg[73]/NET0131  ;
	input \mix1_data_o_reg_reg[74]/NET0131  ;
	input \mix1_data_o_reg_reg[75]/NET0131  ;
	input \mix1_data_o_reg_reg[76]/NET0131  ;
	input \mix1_data_o_reg_reg[77]/NET0131  ;
	input \mix1_data_o_reg_reg[78]/NET0131  ;
	input \mix1_data_o_reg_reg[79]/NET0131  ;
	input \mix1_data_o_reg_reg[7]/NET0131  ;
	input \mix1_data_o_reg_reg[80]/NET0131  ;
	input \mix1_data_o_reg_reg[81]/NET0131  ;
	input \mix1_data_o_reg_reg[82]/NET0131  ;
	input \mix1_data_o_reg_reg[83]/NET0131  ;
	input \mix1_data_o_reg_reg[84]/NET0131  ;
	input \mix1_data_o_reg_reg[85]/NET0131  ;
	input \mix1_data_o_reg_reg[86]/NET0131  ;
	input \mix1_data_o_reg_reg[87]/NET0131  ;
	input \mix1_data_o_reg_reg[88]/NET0131  ;
	input \mix1_data_o_reg_reg[89]/NET0131  ;
	input \mix1_data_o_reg_reg[8]/NET0131  ;
	input \mix1_data_o_reg_reg[90]/NET0131  ;
	input \mix1_data_o_reg_reg[91]/NET0131  ;
	input \mix1_data_o_reg_reg[92]/NET0131  ;
	input \mix1_data_o_reg_reg[93]/NET0131  ;
	input \mix1_data_o_reg_reg[94]/NET0131  ;
	input \mix1_data_o_reg_reg[95]/NET0131  ;
	input \mix1_data_o_reg_reg[96]/NET0131  ;
	input \mix1_data_o_reg_reg[97]/NET0131  ;
	input \mix1_data_o_reg_reg[98]/NET0131  ;
	input \mix1_data_o_reg_reg[99]/NET0131  ;
	input \mix1_data_o_reg_reg[9]/NET0131  ;
	input \mix1_data_reg_reg[100]/NET0131  ;
	input \mix1_data_reg_reg[101]/NET0131  ;
	input \mix1_data_reg_reg[102]/NET0131  ;
	input \mix1_data_reg_reg[103]/NET0131  ;
	input \mix1_data_reg_reg[104]/NET0131  ;
	input \mix1_data_reg_reg[105]/NET0131  ;
	input \mix1_data_reg_reg[106]/NET0131  ;
	input \mix1_data_reg_reg[107]/NET0131  ;
	input \mix1_data_reg_reg[108]/NET0131  ;
	input \mix1_data_reg_reg[109]/NET0131  ;
	input \mix1_data_reg_reg[110]/NET0131  ;
	input \mix1_data_reg_reg[111]/NET0131  ;
	input \mix1_data_reg_reg[112]/NET0131  ;
	input \mix1_data_reg_reg[113]/NET0131  ;
	input \mix1_data_reg_reg[114]/NET0131  ;
	input \mix1_data_reg_reg[115]/NET0131  ;
	input \mix1_data_reg_reg[116]/NET0131  ;
	input \mix1_data_reg_reg[117]/NET0131  ;
	input \mix1_data_reg_reg[118]/NET0131  ;
	input \mix1_data_reg_reg[119]/NET0131  ;
	input \mix1_data_reg_reg[120]/NET0131  ;
	input \mix1_data_reg_reg[121]/NET0131  ;
	input \mix1_data_reg_reg[122]/NET0131  ;
	input \mix1_data_reg_reg[123]/NET0131  ;
	input \mix1_data_reg_reg[124]/NET0131  ;
	input \mix1_data_reg_reg[125]/NET0131  ;
	input \mix1_data_reg_reg[126]/NET0131  ;
	input \mix1_data_reg_reg[127]/NET0131  ;
	input \mix1_data_reg_reg[32]/NET0131  ;
	input \mix1_data_reg_reg[33]/NET0131  ;
	input \mix1_data_reg_reg[34]/NET0131  ;
	input \mix1_data_reg_reg[35]/NET0131  ;
	input \mix1_data_reg_reg[36]/NET0131  ;
	input \mix1_data_reg_reg[37]/NET0131  ;
	input \mix1_data_reg_reg[38]/NET0131  ;
	input \mix1_data_reg_reg[39]/NET0131  ;
	input \mix1_data_reg_reg[40]/NET0131  ;
	input \mix1_data_reg_reg[41]/NET0131  ;
	input \mix1_data_reg_reg[42]/NET0131  ;
	input \mix1_data_reg_reg[43]/NET0131  ;
	input \mix1_data_reg_reg[44]/NET0131  ;
	input \mix1_data_reg_reg[45]/NET0131  ;
	input \mix1_data_reg_reg[46]/NET0131  ;
	input \mix1_data_reg_reg[47]/NET0131  ;
	input \mix1_data_reg_reg[48]/NET0131  ;
	input \mix1_data_reg_reg[49]/NET0131  ;
	input \mix1_data_reg_reg[50]/NET0131  ;
	input \mix1_data_reg_reg[51]/NET0131  ;
	input \mix1_data_reg_reg[52]/NET0131  ;
	input \mix1_data_reg_reg[53]/NET0131  ;
	input \mix1_data_reg_reg[54]/NET0131  ;
	input \mix1_data_reg_reg[55]/NET0131  ;
	input \mix1_data_reg_reg[56]/NET0131  ;
	input \mix1_data_reg_reg[57]/NET0131  ;
	input \mix1_data_reg_reg[58]/NET0131  ;
	input \mix1_data_reg_reg[59]/NET0131  ;
	input \mix1_data_reg_reg[60]/NET0131  ;
	input \mix1_data_reg_reg[61]/NET0131  ;
	input \mix1_data_reg_reg[62]/NET0131  ;
	input \mix1_data_reg_reg[63]/NET0131  ;
	input \mix1_data_reg_reg[64]/NET0131  ;
	input \mix1_data_reg_reg[65]/NET0131  ;
	input \mix1_data_reg_reg[66]/NET0131  ;
	input \mix1_data_reg_reg[67]/NET0131  ;
	input \mix1_data_reg_reg[68]/NET0131  ;
	input \mix1_data_reg_reg[69]/NET0131  ;
	input \mix1_data_reg_reg[70]/NET0131  ;
	input \mix1_data_reg_reg[71]/NET0131  ;
	input \mix1_data_reg_reg[72]/NET0131  ;
	input \mix1_data_reg_reg[73]/NET0131  ;
	input \mix1_data_reg_reg[74]/NET0131  ;
	input \mix1_data_reg_reg[75]/NET0131  ;
	input \mix1_data_reg_reg[76]/NET0131  ;
	input \mix1_data_reg_reg[77]/NET0131  ;
	input \mix1_data_reg_reg[78]/NET0131  ;
	input \mix1_data_reg_reg[79]/NET0131  ;
	input \mix1_data_reg_reg[80]/NET0131  ;
	input \mix1_data_reg_reg[81]/NET0131  ;
	input \mix1_data_reg_reg[82]/NET0131  ;
	input \mix1_data_reg_reg[83]/NET0131  ;
	input \mix1_data_reg_reg[84]/NET0131  ;
	input \mix1_data_reg_reg[85]/NET0131  ;
	input \mix1_data_reg_reg[86]/NET0131  ;
	input \mix1_data_reg_reg[87]/NET0131  ;
	input \mix1_data_reg_reg[88]/NET0131  ;
	input \mix1_data_reg_reg[89]/NET0131  ;
	input \mix1_data_reg_reg[90]/NET0131  ;
	input \mix1_data_reg_reg[91]/NET0131  ;
	input \mix1_data_reg_reg[92]/NET0131  ;
	input \mix1_data_reg_reg[93]/NET0131  ;
	input \mix1_data_reg_reg[94]/NET0131  ;
	input \mix1_data_reg_reg[95]/NET0131  ;
	input \mix1_data_reg_reg[96]/NET0131  ;
	input \mix1_data_reg_reg[97]/NET0131  ;
	input \mix1_data_reg_reg[98]/NET0131  ;
	input \mix1_data_reg_reg[99]/NET0131  ;
	input \mix1_ready_o_reg/NET0131  ;
	input \mix1_state_reg[0]/NET0131  ;
	input \mix1_state_reg[1]/NET0131  ;
	input \round_reg[0]/NET0131  ;
	input \round_reg[1]/NET0131  ;
	input \round_reg[2]/NET0131  ;
	input \round_reg[3]/NET0131  ;
	input \sbox1_ah_reg_reg[0]/NET0131  ;
	input \sbox1_ah_reg_reg[1]/NET0131  ;
	input \sbox1_ah_reg_reg[2]/NET0131  ;
	input \sbox1_ah_reg_reg[3]/NET0131  ;
	input \sbox1_alph_reg[0]/NET0131  ;
	input \sbox1_alph_reg[1]/NET0131  ;
	input \sbox1_alph_reg[2]/NET0131  ;
	input \sbox1_alph_reg[3]/NET0131  ;
	input \sbox1_to_invert_reg[0]/NET0131  ;
	input \sbox1_to_invert_reg[1]/NET0131  ;
	input \sbox1_to_invert_reg[2]/NET0131  ;
	input \sbox1_to_invert_reg[3]/NET0131  ;
	input \state_reg/NET0131  ;
	input \sub1_data_reg_reg[0]/NET0131  ;
	input \sub1_data_reg_reg[100]/NET0131  ;
	input \sub1_data_reg_reg[101]/NET0131  ;
	input \sub1_data_reg_reg[102]/NET0131  ;
	input \sub1_data_reg_reg[103]/NET0131  ;
	input \sub1_data_reg_reg[104]/NET0131  ;
	input \sub1_data_reg_reg[105]/NET0131  ;
	input \sub1_data_reg_reg[106]/NET0131  ;
	input \sub1_data_reg_reg[107]/NET0131  ;
	input \sub1_data_reg_reg[108]/NET0131  ;
	input \sub1_data_reg_reg[109]/NET0131  ;
	input \sub1_data_reg_reg[10]/NET0131  ;
	input \sub1_data_reg_reg[110]/NET0131  ;
	input \sub1_data_reg_reg[111]/NET0131  ;
	input \sub1_data_reg_reg[112]/NET0131  ;
	input \sub1_data_reg_reg[113]/NET0131  ;
	input \sub1_data_reg_reg[114]/NET0131  ;
	input \sub1_data_reg_reg[115]/NET0131  ;
	input \sub1_data_reg_reg[116]/NET0131  ;
	input \sub1_data_reg_reg[117]/NET0131  ;
	input \sub1_data_reg_reg[118]/NET0131  ;
	input \sub1_data_reg_reg[119]/NET0131  ;
	input \sub1_data_reg_reg[11]/NET0131  ;
	input \sub1_data_reg_reg[120]/NET0131  ;
	input \sub1_data_reg_reg[121]/NET0131  ;
	input \sub1_data_reg_reg[122]/NET0131  ;
	input \sub1_data_reg_reg[123]/NET0131  ;
	input \sub1_data_reg_reg[124]/NET0131  ;
	input \sub1_data_reg_reg[125]/NET0131  ;
	input \sub1_data_reg_reg[126]/NET0131  ;
	input \sub1_data_reg_reg[127]/NET0131  ;
	input \sub1_data_reg_reg[12]/NET0131  ;
	input \sub1_data_reg_reg[13]/NET0131  ;
	input \sub1_data_reg_reg[14]/NET0131  ;
	input \sub1_data_reg_reg[15]/NET0131  ;
	input \sub1_data_reg_reg[16]/NET0131  ;
	input \sub1_data_reg_reg[17]/NET0131  ;
	input \sub1_data_reg_reg[18]/NET0131  ;
	input \sub1_data_reg_reg[19]/NET0131  ;
	input \sub1_data_reg_reg[1]/NET0131  ;
	input \sub1_data_reg_reg[20]/NET0131  ;
	input \sub1_data_reg_reg[21]/NET0131  ;
	input \sub1_data_reg_reg[22]/NET0131  ;
	input \sub1_data_reg_reg[23]/NET0131  ;
	input \sub1_data_reg_reg[24]/NET0131  ;
	input \sub1_data_reg_reg[25]/NET0131  ;
	input \sub1_data_reg_reg[26]/NET0131  ;
	input \sub1_data_reg_reg[27]/NET0131  ;
	input \sub1_data_reg_reg[28]/NET0131  ;
	input \sub1_data_reg_reg[29]/NET0131  ;
	input \sub1_data_reg_reg[2]/NET0131  ;
	input \sub1_data_reg_reg[30]/NET0131  ;
	input \sub1_data_reg_reg[31]/NET0131  ;
	input \sub1_data_reg_reg[32]/NET0131  ;
	input \sub1_data_reg_reg[33]/NET0131  ;
	input \sub1_data_reg_reg[34]/NET0131  ;
	input \sub1_data_reg_reg[35]/NET0131  ;
	input \sub1_data_reg_reg[36]/NET0131  ;
	input \sub1_data_reg_reg[37]/NET0131  ;
	input \sub1_data_reg_reg[38]/NET0131  ;
	input \sub1_data_reg_reg[39]/NET0131  ;
	input \sub1_data_reg_reg[3]/NET0131  ;
	input \sub1_data_reg_reg[40]/NET0131  ;
	input \sub1_data_reg_reg[41]/NET0131  ;
	input \sub1_data_reg_reg[42]/NET0131  ;
	input \sub1_data_reg_reg[43]/NET0131  ;
	input \sub1_data_reg_reg[44]/NET0131  ;
	input \sub1_data_reg_reg[45]/NET0131  ;
	input \sub1_data_reg_reg[46]/NET0131  ;
	input \sub1_data_reg_reg[47]/NET0131  ;
	input \sub1_data_reg_reg[48]/NET0131  ;
	input \sub1_data_reg_reg[49]/NET0131  ;
	input \sub1_data_reg_reg[4]/NET0131  ;
	input \sub1_data_reg_reg[50]/NET0131  ;
	input \sub1_data_reg_reg[51]/NET0131  ;
	input \sub1_data_reg_reg[52]/NET0131  ;
	input \sub1_data_reg_reg[53]/NET0131  ;
	input \sub1_data_reg_reg[54]/NET0131  ;
	input \sub1_data_reg_reg[55]/NET0131  ;
	input \sub1_data_reg_reg[56]/NET0131  ;
	input \sub1_data_reg_reg[57]/NET0131  ;
	input \sub1_data_reg_reg[58]/NET0131  ;
	input \sub1_data_reg_reg[59]/NET0131  ;
	input \sub1_data_reg_reg[5]/NET0131  ;
	input \sub1_data_reg_reg[60]/NET0131  ;
	input \sub1_data_reg_reg[61]/NET0131  ;
	input \sub1_data_reg_reg[62]/NET0131  ;
	input \sub1_data_reg_reg[63]/NET0131  ;
	input \sub1_data_reg_reg[64]/NET0131  ;
	input \sub1_data_reg_reg[65]/NET0131  ;
	input \sub1_data_reg_reg[66]/NET0131  ;
	input \sub1_data_reg_reg[67]/NET0131  ;
	input \sub1_data_reg_reg[68]/NET0131  ;
	input \sub1_data_reg_reg[69]/NET0131  ;
	input \sub1_data_reg_reg[6]/NET0131  ;
	input \sub1_data_reg_reg[70]/NET0131  ;
	input \sub1_data_reg_reg[71]/NET0131  ;
	input \sub1_data_reg_reg[72]/NET0131  ;
	input \sub1_data_reg_reg[73]/NET0131  ;
	input \sub1_data_reg_reg[74]/NET0131  ;
	input \sub1_data_reg_reg[75]/NET0131  ;
	input \sub1_data_reg_reg[76]/NET0131  ;
	input \sub1_data_reg_reg[77]/NET0131  ;
	input \sub1_data_reg_reg[78]/NET0131  ;
	input \sub1_data_reg_reg[79]/NET0131  ;
	input \sub1_data_reg_reg[7]/NET0131  ;
	input \sub1_data_reg_reg[80]/NET0131  ;
	input \sub1_data_reg_reg[81]/NET0131  ;
	input \sub1_data_reg_reg[82]/NET0131  ;
	input \sub1_data_reg_reg[83]/NET0131  ;
	input \sub1_data_reg_reg[84]/NET0131  ;
	input \sub1_data_reg_reg[85]/NET0131  ;
	input \sub1_data_reg_reg[86]/NET0131  ;
	input \sub1_data_reg_reg[87]/NET0131  ;
	input \sub1_data_reg_reg[88]/NET0131  ;
	input \sub1_data_reg_reg[89]/NET0131  ;
	input \sub1_data_reg_reg[8]/NET0131  ;
	input \sub1_data_reg_reg[90]/NET0131  ;
	input \sub1_data_reg_reg[91]/NET0131  ;
	input \sub1_data_reg_reg[92]/NET0131  ;
	input \sub1_data_reg_reg[93]/NET0131  ;
	input \sub1_data_reg_reg[94]/NET0131  ;
	input \sub1_data_reg_reg[95]/NET0131  ;
	input \sub1_data_reg_reg[96]/NET0131  ;
	input \sub1_data_reg_reg[97]/NET0131  ;
	input \sub1_data_reg_reg[98]/NET0131  ;
	input \sub1_data_reg_reg[99]/NET0131  ;
	input \sub1_data_reg_reg[9]/NET0131  ;
	input \sub1_ready_o_reg/NET0131  ;
	input \sub1_state_reg[0]/NET0131  ;
	input \sub1_state_reg[1]/NET0131  ;
	input \sub1_state_reg[2]/NET0131  ;
	input \sub1_state_reg[3]/NET0131  ;
	input \sub1_state_reg[4]/NET0131  ;
	output \_al_n0  ;
	output \_al_n1  ;
	output \g27929/_0_  ;
	output \g27942/_3_  ;
	output \g27943/_3_  ;
	output \g27944/_3_  ;
	output \g27945/_0_  ;
	output \g27995/_0_  ;
	output \g27998/_0_  ;
	output \g28019/_0_  ;
	output \g28020/_0_  ;
	output \g28021/_0_  ;
	output \g28022/_0_  ;
	output \g28023/_0_  ;
	output \g28024/_0_  ;
	output \g28025/_0_  ;
	output \g28026/_0_  ;
	output \g28027/_0_  ;
	output \g28028/_0_  ;
	output \g28029/_0_  ;
	output \g28030/_0_  ;
	output \g28031/_0_  ;
	output \g28032/_0_  ;
	output \g28033/_0_  ;
	output \g28034/_0_  ;
	output \g28044/_0_  ;
	output \g28045/_0_  ;
	output \g28046/_0_  ;
	output \g28047/_0_  ;
	output \g28048/_0_  ;
	output \g28049/_0_  ;
	output \g28050/_0_  ;
	output \g28051/_0_  ;
	output \g28151/_0_  ;
	output \g28177/_0_  ;
	output \g28178/_0_  ;
	output \g28179/_0_  ;
	output \g28180/_0_  ;
	output \g28181/_0_  ;
	output \g28182/_0_  ;
	output \g28183/_0_  ;
	output \g28184/_0_  ;
	output \g28185/_0_  ;
	output \g28186/_0_  ;
	output \g28187/_0_  ;
	output \g28188/_0_  ;
	output \g28189/_0_  ;
	output \g28190/_0_  ;
	output \g28191/_0_  ;
	output \g28192/_0_  ;
	output \g28193/_0_  ;
	output \g28194/_0_  ;
	output \g28195/_0_  ;
	output \g28196/_0_  ;
	output \g28197/_0_  ;
	output \g28198/_0_  ;
	output \g28199/_0_  ;
	output \g28200/_0_  ;
	output \g28201/_0_  ;
	output \g28202/_0_  ;
	output \g28203/_0_  ;
	output \g28253/_0_  ;
	output \g28254/_0_  ;
	output \g28255/_0_  ;
	output \g28256/_0_  ;
	output \g28257/_0_  ;
	output \g28258/_0_  ;
	output \g28259/_0_  ;
	output \g28260/_0_  ;
	output \g28261/_0_  ;
	output \g28262/_0_  ;
	output \g28263/_0_  ;
	output \g28264/_0_  ;
	output \g28265/_0_  ;
	output \g28266/_0_  ;
	output \g28267/_0_  ;
	output \g28268/_0_  ;
	output \g28269/_0_  ;
	output \g28270/_0_  ;
	output \g28271/_0_  ;
	output \g28272/_0_  ;
	output \g28273/_0_  ;
	output \g28274/_0_  ;
	output \g28275/_0_  ;
	output \g28276/_0_  ;
	output \g28277/_0_  ;
	output \g28278/_0_  ;
	output \g28279/_0_  ;
	output \g28384/_2_  ;
	output \g28385/_2_  ;
	output \g28388/_2_  ;
	output \g28389/_2_  ;
	output \g28394/_2_  ;
	output \g28395/_2_  ;
	output \g28401/_2_  ;
	output \g28402/_2_  ;
	output \g28403/_0_  ;
	output \g28404/_0_  ;
	output \g28408/_0_  ;
	output \g28410/_0_  ;
	output \g28440/_0_  ;
	output \g28441/_0_  ;
	output \g28442/_0_  ;
	output \g28443/_0_  ;
	output \g28444/_0_  ;
	output \g28445/_0_  ;
	output \g28446/_0_  ;
	output \g28447/_0_  ;
	output \g28448/_0_  ;
	output \g28449/_0_  ;
	output \g28450/_0_  ;
	output \g28451/_0_  ;
	output \g28452/_0_  ;
	output \g28453/_0_  ;
	output \g28538/_0_  ;
	output \g28539/_0_  ;
	output \g28540/_0_  ;
	output \g28541/_0_  ;
	output \g28542/_0_  ;
	output \g28543/_0_  ;
	output \g28544/_0_  ;
	output \g28545/_0_  ;
	output \g28546/_0_  ;
	output \g28547/_0_  ;
	output \g28548/_0_  ;
	output \g28549/_0_  ;
	output \g28550/_0_  ;
	output \g28551/_0_  ;
	output \g28552/_0_  ;
	output \g28557/_0_  ;
	output \g28558/_0_  ;
	output \g28563/_0_  ;
	output \g28564/_0_  ;
	output \g28565/_0_  ;
	output \g28566/_0_  ;
	output \g28567/_0_  ;
	output \g28625/_2_  ;
	output \g28626/_2_  ;
	output \g28633/_2_  ;
	output \g28639/_2_  ;
	output \g28655/_2_  ;
	output \g28656/_2_  ;
	output \g28657/_2_  ;
	output \g28660/_2_  ;
	output \g28661/_2_  ;
	output \g28662/_2_  ;
	output \g28666/_2_  ;
	output \g28667/_2_  ;
	output \g28668/_2_  ;
	output \g28678/_2_  ;
	output \g28679/_2_  ;
	output \g28680/_2_  ;
	output \g28690/_0_  ;
	output \g28710/_0_  ;
	output \g28716/_0_  ;
	output \g28795/_0_  ;
	output \g28796/_0_  ;
	output \g28798/_0_  ;
	output \g28799/_0_  ;
	output \g28800/_0_  ;
	output \g28801/_0_  ;
	output \g28804/_0_  ;
	output \g28825/_2_  ;
	output \g28826/_2_  ;
	output \g28830/_2_  ;
	output \g28834/_2_  ;
	output \g28842/_2_  ;
	output \g28843/_2_  ;
	output \g28845/_2_  ;
	output \g28848/_2_  ;
	output \g28890/_0_  ;
	output \g28936/_0_  ;
	output \g28982/_0_  ;
	output \g29050/_0_  ;
	output \g29051/_0_  ;
	output \g29052/_0_  ;
	output \g29053/_0_  ;
	output \g29054/_0_  ;
	output \g29055/_0_  ;
	output \g29056/_0_  ;
	output \g29057/_0_  ;
	output \g29058/_0_  ;
	output \g29059/_0_  ;
	output \g29060/_0_  ;
	output \g29061/_0_  ;
	output \g29328/_0_  ;
	output \g29329/_0_  ;
	output \g29330/_0_  ;
	output \g29331/_0_  ;
	output \g29332/_0_  ;
	output \g29333/_0_  ;
	output \g29334/_0_  ;
	output \g29335/_0_  ;
	output \g29336/_0_  ;
	output \g29337/_0_  ;
	output \g29338/_0_  ;
	output \g29339/_0_  ;
	output \g29340/_0_  ;
	output \g29341/_0_  ;
	output \g29342/_0_  ;
	output \g29343/_0_  ;
	output \g29344/_0_  ;
	output \g29345/_0_  ;
	output \g29346/_0_  ;
	output \g29347/_0_  ;
	output \g29348/_0_  ;
	output \g29349/_0_  ;
	output \g29350/_0_  ;
	output \g29351/_0_  ;
	output \g29352/_0_  ;
	output \g29353/_0_  ;
	output \g29354/_0_  ;
	output \g29355/_0_  ;
	output \g29356/_0_  ;
	output \g29357/_0_  ;
	output \g29358/_0_  ;
	output \g29359/_0_  ;
	output \g29360/_0_  ;
	output \g29361/_0_  ;
	output \g29362/_0_  ;
	output \g29363/_0_  ;
	output \g29364/_0_  ;
	output \g29365/_0_  ;
	output \g29366/_0_  ;
	output \g29367/_0_  ;
	output \g29395/_0_  ;
	output \g29396/_0_  ;
	output \g29453/_0_  ;
	output \g29454/_0_  ;
	output \g29455/_0_  ;
	output \g29456/_0_  ;
	output \g29457/_0_  ;
	output \g29458/_0_  ;
	output \g29459/_0_  ;
	output \g29460/_0_  ;
	output \g29461/_0_  ;
	output \g29462/_0_  ;
	output \g29463/_0_  ;
	output \g29464/_0_  ;
	output \g29465/_0_  ;
	output \g29466/_0_  ;
	output \g29467/_0_  ;
	output \g29468/_0_  ;
	output \g29469/_0_  ;
	output \g29470/_0_  ;
	output \g29471/_0_  ;
	output \g29472/_0_  ;
	output \g29473/_0_  ;
	output \g29474/_0_  ;
	output \g29475/_0_  ;
	output \g29476/_0_  ;
	output \g29477/_0_  ;
	output \g29478/_0_  ;
	output \g29479/_0_  ;
	output \g29480/_0_  ;
	output \g29481/_0_  ;
	output \g29482/_0_  ;
	output \g29483/_0_  ;
	output \g29484/_0_  ;
	output \g29485/_0_  ;
	output \g29486/_0_  ;
	output \g29487/_0_  ;
	output \g29488/_0_  ;
	output \g29489/_0_  ;
	output \g29490/_0_  ;
	output \g29491/_0_  ;
	output \g29492/_0_  ;
	output \g29493/_0_  ;
	output \g29494/_0_  ;
	output \g29495/_0_  ;
	output \g29496/_0_  ;
	output \g29497/_0_  ;
	output \g29498/_0_  ;
	output \g29499/_0_  ;
	output \g29500/_0_  ;
	output \g29501/_0_  ;
	output \g29502/_0_  ;
	output \g29503/_0_  ;
	output \g29504/_0_  ;
	output \g29505/_0_  ;
	output \g29506/_0_  ;
	output \g29507/_0_  ;
	output \g29508/_0_  ;
	output \g29509/_0_  ;
	output \g29510/_0_  ;
	output \g29511/_0_  ;
	output \g29512/_0_  ;
	output \g29513/_0_  ;
	output \g29514/_0_  ;
	output \g29515/_0_  ;
	output \g29516/_0_  ;
	output \g29517/_0_  ;
	output \g29518/_0_  ;
	output \g29519/_0_  ;
	output \g29520/_0_  ;
	output \g29521/_0_  ;
	output \g29522/_0_  ;
	output \g29523/_0_  ;
	output \g29524/_0_  ;
	output \g29525/_0_  ;
	output \g29526/_0_  ;
	output \g29527/_0_  ;
	output \g29528/_0_  ;
	output \g29529/_0_  ;
	output \g29530/_0_  ;
	output \g29531/_0_  ;
	output \g29532/_0_  ;
	output \g29533/_0_  ;
	output \g29534/_0_  ;
	output \g29535/_0_  ;
	output \g29536/_0_  ;
	output \g29537/_0_  ;
	output \g29538/_0_  ;
	output \g29539/_0_  ;
	output \g29540/_0_  ;
	output \g29541/_0_  ;
	output \g29542/_0_  ;
	output \g29543/_0_  ;
	output \g29544/_0_  ;
	output \g29545/_0_  ;
	output \g29546/_0_  ;
	output \g29547/_0_  ;
	output \g29548/_0_  ;
	output \g29549/_0_  ;
	output \g29550/_0_  ;
	output \g29551/_0_  ;
	output \g29552/_0_  ;
	output \g29553/_0_  ;
	output \g29554/_0_  ;
	output \g29555/_0_  ;
	output \g29556/_0_  ;
	output \g29557/_0_  ;
	output \g29558/_0_  ;
	output \g29559/_0_  ;
	output \g29560/_0_  ;
	output \g29561/_0_  ;
	output \g29562/_0_  ;
	output \g29563/_0_  ;
	output \g29564/_0_  ;
	output \g29565/_0_  ;
	output \g29566/_0_  ;
	output \g29567/_0_  ;
	output \g29568/_0_  ;
	output \g29569/_0_  ;
	output \g29570/_0_  ;
	output \g29571/_0_  ;
	output \g29572/_0_  ;
	output \g29573/_0_  ;
	output \g29574/_0_  ;
	output \g29575/_0_  ;
	output \g29576/_0_  ;
	output \g29577/_0_  ;
	output \g29578/_0_  ;
	output \g29579/_0_  ;
	output \g29580/_0_  ;
	output \g29582/_0_  ;
	output \g29583/_0_  ;
	output \g29584/_0_  ;
	output \g29585/_0_  ;
	output \g29586/_0_  ;
	output \g29587/_0_  ;
	output \g29588/_0_  ;
	output \g29589/_0_  ;
	output \g29590/_0_  ;
	output \g29591/_0_  ;
	output \g29592/_0_  ;
	output \g29593/_0_  ;
	output \g29634/_0_  ;
	output \g29635/_0_  ;
	output \g29636/_0_  ;
	output \g29637/_0_  ;
	output \g29645/_0_  ;
	output \g29646/_0_  ;
	output \g29647/_0_  ;
	output \g29824/_0_  ;
	output \g29828/_0_  ;
	output \g29832/_0_  ;
	output \g29836/_0_  ;
	output \g29837/_0_  ;
	output \g29838/_0_  ;
	output \g29839/_0_  ;
	output \g29840/_0_  ;
	output \g29841/_0_  ;
	output \g29842/_0_  ;
	output \g29843/_0_  ;
	output \g29844/_0_  ;
	output \g29845/_0_  ;
	output \g29846/_0_  ;
	output \g29847/_0_  ;
	output \g29848/_0_  ;
	output \g29849/_0_  ;
	output \g29850/_0_  ;
	output \g29851/_0_  ;
	output \g29852/_0_  ;
	output \g29853/_0_  ;
	output \g29854/_0_  ;
	output \g29855/_0_  ;
	output \g29856/_0_  ;
	output \g29857/_0_  ;
	output \g29858/_0_  ;
	output \g29859/_0_  ;
	output \g29860/_0_  ;
	output \g29861/_0_  ;
	output \g29862/_0_  ;
	output \g29863/_0_  ;
	output \g29864/_0_  ;
	output \g29865/_0_  ;
	output \g29866/_0_  ;
	output \g29867/_0_  ;
	output \g29868/_0_  ;
	output \g30081/_0_  ;
	output \g30082/_0_  ;
	output \g30083/_0_  ;
	output \g30084/_0_  ;
	output \g30085/_0_  ;
	output \g30086/_0_  ;
	output \g30087/_0_  ;
	output \g30088/_0_  ;
	output \g30089/_0_  ;
	output \g30090/_0_  ;
	output \g30091/_0_  ;
	output \g30092/_0_  ;
	output \g30093/_0_  ;
	output \g30094/_0_  ;
	output \g30095/_0_  ;
	output \g30096/_0_  ;
	output \g30135/_0_  ;
	output \g30137/_0_  ;
	output \g30164/_0_  ;
	output \g30165/_0_  ;
	output \g30166/_0_  ;
	output \g30167/_0_  ;
	output \g30168/_0_  ;
	output \g30169/_0_  ;
	output \g30170/_0_  ;
	output \g30231/_0_  ;
	output \g30232/_0_  ;
	output \g30233/_0_  ;
	output \g30234/_0_  ;
	output \g30235/_0_  ;
	output \g30236/_0_  ;
	output \g30237/_0_  ;
	output \g30238/_0_  ;
	output \g30286/_0_  ;
	output \g30287/_0_  ;
	output \g30288/_0_  ;
	output \g30289/_0_  ;
	output \g30290/_0_  ;
	output \g30291/_0_  ;
	output \g30292/_0_  ;
	output \g30293/_0_  ;
	output \g30294/_0_  ;
	output \g30295/_0_  ;
	output \g30296/_0_  ;
	output \g30297/_0_  ;
	output \g30298/_0_  ;
	output \g30299/_0_  ;
	output \g30300/_0_  ;
	output \g30301/_0_  ;
	output \g30303/_0_  ;
	output \g30304/_0_  ;
	output \g30305/_0_  ;
	output \g30306/_0_  ;
	output \g30307/_0_  ;
	output \g30308/_0_  ;
	output \g30309/_0_  ;
	output \g30310/_0_  ;
	output \g30311/_0_  ;
	output \g30312/_0_  ;
	output \g30313/_0_  ;
	output \g30314/_0_  ;
	output \g30315/_0_  ;
	output \g30316/_0_  ;
	output \g30317/_0_  ;
	output \g30318/_0_  ;
	output \g30319/_0_  ;
	output \g30481/_0_  ;
	output \g30482/_0_  ;
	output \g30483/_0_  ;
	output \g30484/_0_  ;
	output \g30493/_0_  ;
	output \g30495/_0_  ;
	output \g30536/_0_  ;
	output \g30537/_0_  ;
	output \g30538/_0_  ;
	output \g30735/_0_  ;
	output \g30927/_0_  ;
	output \g30928/_0_  ;
	output \g30929/_0_  ;
	output \g30971/_0_  ;
	output \g30972/_0_  ;
	output \g30973/_0_  ;
	output \g30974/_0_  ;
	output \g31129/_0_  ;
	output \g31130/_0_  ;
	output \g31131/_0_  ;
	output \g31132/_0_  ;
	output \g31133/_0_  ;
	output \g31134/_0_  ;
	output \g31135/_0_  ;
	output \g31136/_0_  ;
	output \g31137/_0_  ;
	output \g31138/_0_  ;
	output \g31139/_0_  ;
	output \g31140/_0_  ;
	output \g31141/_0_  ;
	output \g31142/_0_  ;
	output \g31143/_0_  ;
	output \g31144/_0_  ;
	output \g31352/_0_  ;
	output \g31353/_0_  ;
	output \g31354/_0_  ;
	output \g31355/_0_  ;
	output \g31356/_0_  ;
	output \g31357/_0_  ;
	output \g31358/_0_  ;
	output \g31359/_0_  ;
	output \g31360/_0_  ;
	output \g31361/_0_  ;
	output \g31362/_0_  ;
	output \g31363/_0_  ;
	output \g31364/_0_  ;
	output \g31365/_0_  ;
	output \g31366/_0_  ;
	output \g31367/_0_  ;
	output \g31706/_0_  ;
	output \g32001/_0_  ;
	output \g32008/_0_  ;
	output \g32009/_0_  ;
	output \g32010/_0_  ;
	output \g32011/_0_  ;
	output \g32118/_0_  ;
	output \g33261/_0_  ;
	output \g33262/_0_  ;
	output \g33263/_0_  ;
	output \g33264/_0_  ;
	output \g33265/_0_  ;
	output \g33266/_0_  ;
	output \g33450/_0_  ;
	output \g33451/_0_  ;
	output \g33453/_0_  ;
	output \g33485/_0_  ;
	output \g33679/_2_  ;
	output \g34838/_2_  ;
	output \g34971/_0_  ;
	output \g34972/_0_  ;
	output \g34973/_0_  ;
	output \g34974/_0_  ;
	output \g34975/_0_  ;
	output \g34976/_0_  ;
	output \g34977/_0_  ;
	output \g34978/_0_  ;
	output \g34979/_0_  ;
	output \g34980/_0_  ;
	output \g34981/_0_  ;
	output \g34982/_0_  ;
	output \g34983/_0_  ;
	output \g34984/_0_  ;
	output \g34985/_0_  ;
	output \g34986/_0_  ;
	output \g34987/_0_  ;
	output \g34988/_0_  ;
	output \g34989/_0_  ;
	output \g34990/_0_  ;
	output \g34991/_0_  ;
	output \g34992/_0_  ;
	output \g34993/_0_  ;
	output \g34994/_0_  ;
	output \g34995/_0_  ;
	output \g34996/_0_  ;
	output \g34997/_0_  ;
	output \g34998/_0_  ;
	output \g34999/_0_  ;
	output \g35000/_0_  ;
	output \g35001/_0_  ;
	output \g35002/_0_  ;
	output \g35003/_0_  ;
	output \g35004/_0_  ;
	output \g35005/_0_  ;
	output \g35006/_0_  ;
	output \g35007/_0_  ;
	output \g35008/_0_  ;
	output \g35009/_0_  ;
	output \g35010/_0_  ;
	output \g35011/_0_  ;
	output \g35012/_0_  ;
	output \g35013/_0_  ;
	output \g35014/_0_  ;
	output \g35015/_0_  ;
	output \g35016/_0_  ;
	output \g35017/_0_  ;
	output \g35018/_0_  ;
	output \g35019/_0_  ;
	output \g35020/_0_  ;
	output \g35021/_0_  ;
	output \g35022/_0_  ;
	output \g35023/_0_  ;
	output \g35024/_0_  ;
	output \g35025/_0_  ;
	output \g35026/_0_  ;
	output \g35027/_0_  ;
	output \g35028/_0_  ;
	output \g35029/_0_  ;
	output \g35030/_0_  ;
	output \g35031/_0_  ;
	output \g35032/_0_  ;
	output \g35033/_0_  ;
	output \g35034/_0_  ;
	output \g35035/_0_  ;
	output \g35036/_0_  ;
	output \g35037/_0_  ;
	output \g35038/_0_  ;
	output \g35039/_0_  ;
	output \g35040/_0_  ;
	output \g35041/_0_  ;
	output \g35042/_0_  ;
	output \g35043/_0_  ;
	output \g35044/_0_  ;
	output \g35045/_0_  ;
	output \g35046/_0_  ;
	output \g35047/_0_  ;
	output \g35048/_0_  ;
	output \g35049/_0_  ;
	output \g35050/_0_  ;
	output \g35051/_0_  ;
	output \g35052/_0_  ;
	output \g35053/_0_  ;
	output \g35054/_0_  ;
	output \g35055/_0_  ;
	output \g35056/_0_  ;
	output \g35057/_0_  ;
	output \g35058/_0_  ;
	output \g35059/_0_  ;
	output \g35060/_0_  ;
	output \g35061/_0_  ;
	output \g35062/_0_  ;
	output \g35063/_0_  ;
	output \g35064/_0_  ;
	output \g35065/_0_  ;
	output \g35066/_0_  ;
	output \g35538/_0_  ;
	output \g35956/_0_  ;
	output \g36298/_1_  ;
	output \g36324/_0_  ;
	output \g36375/_0_  ;
	output \g38269/_0_  ;
	output \g38473/_0_  ;
	output \g38501/_0_  ;
	output \g38569/_0_  ;
	output \g38629/_0_  ;
	output \g38721_dup/_3_  ;
	output \g38735/_0_  ;
	output \g38753/_0_  ;
	output \g38849/_3_  ;
	output \g39071/_0_  ;
	output \g39073/_0_  ;
	output \g39077/_0_  ;
	output \g39080/_0_  ;
	output \g39135/_0_  ;
	output \g39138/_0_  ;
	output \g39182/_0_  ;
	output \g39197/_3_  ;
	output \g39207/_3_  ;
	output \g39241/_0_  ;
	output \g39272/_0_  ;
	output \g39307/_0_  ;
	output \g39308/_0_  ;
	output \g39361/_0_  ;
	output \g39494/_0_  ;
	output \g39558/_0_  ;
	output \g39575/_0_  ;
	output \g39583/_0_  ;
	wire _w4661_ ;
	wire _w4660_ ;
	wire _w4659_ ;
	wire _w4658_ ;
	wire _w4657_ ;
	wire _w4656_ ;
	wire _w4655_ ;
	wire _w4654_ ;
	wire _w4653_ ;
	wire _w4652_ ;
	wire _w4651_ ;
	wire _w4650_ ;
	wire _w4649_ ;
	wire _w4648_ ;
	wire _w4647_ ;
	wire _w4646_ ;
	wire _w4645_ ;
	wire _w4644_ ;
	wire _w4643_ ;
	wire _w4642_ ;
	wire _w4641_ ;
	wire _w4640_ ;
	wire _w4639_ ;
	wire _w4638_ ;
	wire _w4637_ ;
	wire _w4636_ ;
	wire _w4635_ ;
	wire _w4634_ ;
	wire _w4633_ ;
	wire _w4632_ ;
	wire _w4631_ ;
	wire _w4630_ ;
	wire _w4629_ ;
	wire _w4628_ ;
	wire _w4627_ ;
	wire _w4626_ ;
	wire _w4625_ ;
	wire _w4624_ ;
	wire _w4623_ ;
	wire _w4622_ ;
	wire _w4621_ ;
	wire _w4620_ ;
	wire _w4619_ ;
	wire _w4618_ ;
	wire _w4617_ ;
	wire _w4616_ ;
	wire _w4615_ ;
	wire _w4614_ ;
	wire _w4613_ ;
	wire _w4612_ ;
	wire _w4611_ ;
	wire _w4610_ ;
	wire _w4609_ ;
	wire _w4608_ ;
	wire _w4607_ ;
	wire _w4606_ ;
	wire _w4605_ ;
	wire _w4604_ ;
	wire _w4603_ ;
	wire _w4602_ ;
	wire _w4601_ ;
	wire _w4600_ ;
	wire _w4599_ ;
	wire _w4598_ ;
	wire _w4597_ ;
	wire _w4596_ ;
	wire _w4595_ ;
	wire _w4594_ ;
	wire _w4593_ ;
	wire _w4592_ ;
	wire _w4591_ ;
	wire _w4590_ ;
	wire _w4589_ ;
	wire _w4588_ ;
	wire _w4587_ ;
	wire _w4586_ ;
	wire _w4585_ ;
	wire _w4584_ ;
	wire _w4583_ ;
	wire _w4582_ ;
	wire _w4581_ ;
	wire _w4580_ ;
	wire _w4579_ ;
	wire _w4578_ ;
	wire _w4577_ ;
	wire _w4576_ ;
	wire _w4575_ ;
	wire _w4574_ ;
	wire _w4573_ ;
	wire _w4572_ ;
	wire _w4571_ ;
	wire _w4570_ ;
	wire _w4569_ ;
	wire _w4568_ ;
	wire _w4567_ ;
	wire _w4566_ ;
	wire _w4565_ ;
	wire _w4564_ ;
	wire _w4563_ ;
	wire _w4562_ ;
	wire _w4561_ ;
	wire _w4560_ ;
	wire _w4559_ ;
	wire _w4558_ ;
	wire _w4557_ ;
	wire _w4556_ ;
	wire _w4555_ ;
	wire _w4554_ ;
	wire _w4553_ ;
	wire _w4552_ ;
	wire _w4551_ ;
	wire _w4550_ ;
	wire _w4549_ ;
	wire _w4548_ ;
	wire _w4547_ ;
	wire _w4546_ ;
	wire _w4545_ ;
	wire _w4544_ ;
	wire _w4543_ ;
	wire _w4542_ ;
	wire _w4541_ ;
	wire _w4540_ ;
	wire _w4539_ ;
	wire _w4538_ ;
	wire _w4537_ ;
	wire _w4536_ ;
	wire _w4535_ ;
	wire _w4534_ ;
	wire _w4533_ ;
	wire _w4532_ ;
	wire _w4531_ ;
	wire _w4530_ ;
	wire _w4529_ ;
	wire _w4528_ ;
	wire _w4527_ ;
	wire _w4526_ ;
	wire _w4525_ ;
	wire _w4524_ ;
	wire _w4523_ ;
	wire _w4522_ ;
	wire _w4521_ ;
	wire _w4520_ ;
	wire _w4519_ ;
	wire _w4518_ ;
	wire _w4517_ ;
	wire _w4516_ ;
	wire _w4515_ ;
	wire _w4514_ ;
	wire _w4513_ ;
	wire _w4512_ ;
	wire _w4511_ ;
	wire _w4510_ ;
	wire _w4509_ ;
	wire _w4508_ ;
	wire _w4507_ ;
	wire _w4506_ ;
	wire _w4505_ ;
	wire _w4504_ ;
	wire _w4503_ ;
	wire _w4502_ ;
	wire _w4501_ ;
	wire _w4500_ ;
	wire _w4499_ ;
	wire _w4498_ ;
	wire _w4497_ ;
	wire _w4496_ ;
	wire _w4495_ ;
	wire _w4494_ ;
	wire _w4493_ ;
	wire _w4492_ ;
	wire _w4491_ ;
	wire _w4490_ ;
	wire _w4489_ ;
	wire _w4488_ ;
	wire _w4487_ ;
	wire _w4486_ ;
	wire _w4485_ ;
	wire _w4484_ ;
	wire _w4483_ ;
	wire _w4482_ ;
	wire _w4481_ ;
	wire _w4480_ ;
	wire _w4479_ ;
	wire _w4478_ ;
	wire _w4477_ ;
	wire _w4476_ ;
	wire _w4475_ ;
	wire _w4474_ ;
	wire _w4473_ ;
	wire _w4472_ ;
	wire _w4471_ ;
	wire _w4470_ ;
	wire _w4469_ ;
	wire _w4468_ ;
	wire _w4467_ ;
	wire _w4466_ ;
	wire _w4465_ ;
	wire _w4464_ ;
	wire _w4463_ ;
	wire _w4462_ ;
	wire _w4461_ ;
	wire _w4460_ ;
	wire _w4459_ ;
	wire _w4458_ ;
	wire _w4457_ ;
	wire _w4456_ ;
	wire _w4455_ ;
	wire _w4454_ ;
	wire _w4453_ ;
	wire _w4452_ ;
	wire _w4451_ ;
	wire _w4450_ ;
	wire _w4449_ ;
	wire _w4448_ ;
	wire _w4447_ ;
	wire _w4446_ ;
	wire _w4445_ ;
	wire _w4444_ ;
	wire _w4443_ ;
	wire _w4442_ ;
	wire _w4441_ ;
	wire _w4440_ ;
	wire _w4439_ ;
	wire _w4438_ ;
	wire _w4437_ ;
	wire _w4436_ ;
	wire _w4435_ ;
	wire _w4434_ ;
	wire _w4433_ ;
	wire _w4432_ ;
	wire _w4431_ ;
	wire _w4430_ ;
	wire _w4429_ ;
	wire _w4428_ ;
	wire _w4427_ ;
	wire _w4426_ ;
	wire _w4425_ ;
	wire _w4424_ ;
	wire _w4423_ ;
	wire _w4422_ ;
	wire _w4421_ ;
	wire _w4420_ ;
	wire _w4419_ ;
	wire _w4418_ ;
	wire _w4417_ ;
	wire _w4416_ ;
	wire _w4415_ ;
	wire _w4414_ ;
	wire _w4413_ ;
	wire _w4412_ ;
	wire _w4411_ ;
	wire _w4410_ ;
	wire _w4409_ ;
	wire _w4408_ ;
	wire _w4407_ ;
	wire _w4406_ ;
	wire _w4405_ ;
	wire _w4404_ ;
	wire _w4403_ ;
	wire _w4402_ ;
	wire _w4401_ ;
	wire _w4400_ ;
	wire _w4399_ ;
	wire _w4398_ ;
	wire _w4397_ ;
	wire _w4396_ ;
	wire _w4395_ ;
	wire _w4394_ ;
	wire _w4393_ ;
	wire _w4392_ ;
	wire _w4391_ ;
	wire _w4390_ ;
	wire _w4389_ ;
	wire _w4388_ ;
	wire _w4387_ ;
	wire _w4386_ ;
	wire _w4385_ ;
	wire _w4384_ ;
	wire _w4383_ ;
	wire _w4382_ ;
	wire _w4381_ ;
	wire _w4380_ ;
	wire _w4379_ ;
	wire _w4378_ ;
	wire _w4377_ ;
	wire _w4376_ ;
	wire _w4375_ ;
	wire _w4374_ ;
	wire _w4373_ ;
	wire _w4372_ ;
	wire _w4371_ ;
	wire _w4370_ ;
	wire _w4369_ ;
	wire _w4368_ ;
	wire _w4367_ ;
	wire _w4366_ ;
	wire _w4365_ ;
	wire _w4364_ ;
	wire _w4363_ ;
	wire _w4362_ ;
	wire _w4361_ ;
	wire _w4360_ ;
	wire _w4359_ ;
	wire _w4358_ ;
	wire _w4357_ ;
	wire _w4356_ ;
	wire _w4355_ ;
	wire _w4354_ ;
	wire _w4353_ ;
	wire _w4352_ ;
	wire _w4351_ ;
	wire _w4350_ ;
	wire _w4349_ ;
	wire _w4348_ ;
	wire _w4347_ ;
	wire _w4346_ ;
	wire _w4345_ ;
	wire _w4344_ ;
	wire _w4343_ ;
	wire _w4342_ ;
	wire _w4341_ ;
	wire _w4340_ ;
	wire _w4339_ ;
	wire _w4338_ ;
	wire _w4337_ ;
	wire _w4336_ ;
	wire _w4335_ ;
	wire _w4334_ ;
	wire _w4333_ ;
	wire _w4332_ ;
	wire _w4331_ ;
	wire _w4330_ ;
	wire _w4329_ ;
	wire _w4328_ ;
	wire _w4327_ ;
	wire _w4326_ ;
	wire _w4325_ ;
	wire _w4324_ ;
	wire _w4323_ ;
	wire _w4322_ ;
	wire _w4321_ ;
	wire _w4320_ ;
	wire _w4319_ ;
	wire _w4318_ ;
	wire _w4317_ ;
	wire _w4316_ ;
	wire _w4315_ ;
	wire _w4314_ ;
	wire _w4313_ ;
	wire _w4312_ ;
	wire _w4311_ ;
	wire _w4310_ ;
	wire _w4309_ ;
	wire _w4308_ ;
	wire _w4307_ ;
	wire _w4306_ ;
	wire _w4305_ ;
	wire _w4304_ ;
	wire _w4303_ ;
	wire _w4302_ ;
	wire _w4301_ ;
	wire _w4300_ ;
	wire _w4299_ ;
	wire _w4298_ ;
	wire _w4297_ ;
	wire _w4296_ ;
	wire _w4295_ ;
	wire _w4294_ ;
	wire _w4293_ ;
	wire _w4292_ ;
	wire _w4291_ ;
	wire _w4290_ ;
	wire _w4289_ ;
	wire _w4288_ ;
	wire _w4287_ ;
	wire _w4286_ ;
	wire _w4285_ ;
	wire _w4284_ ;
	wire _w4283_ ;
	wire _w4282_ ;
	wire _w4281_ ;
	wire _w4280_ ;
	wire _w4279_ ;
	wire _w4278_ ;
	wire _w4277_ ;
	wire _w4276_ ;
	wire _w4275_ ;
	wire _w4274_ ;
	wire _w4273_ ;
	wire _w4272_ ;
	wire _w4271_ ;
	wire _w4270_ ;
	wire _w4269_ ;
	wire _w4268_ ;
	wire _w4267_ ;
	wire _w4266_ ;
	wire _w4265_ ;
	wire _w4264_ ;
	wire _w4263_ ;
	wire _w4262_ ;
	wire _w4261_ ;
	wire _w4260_ ;
	wire _w4259_ ;
	wire _w4258_ ;
	wire _w4257_ ;
	wire _w4256_ ;
	wire _w4255_ ;
	wire _w4254_ ;
	wire _w4253_ ;
	wire _w4252_ ;
	wire _w4251_ ;
	wire _w4250_ ;
	wire _w4249_ ;
	wire _w4248_ ;
	wire _w4247_ ;
	wire _w4246_ ;
	wire _w4245_ ;
	wire _w4244_ ;
	wire _w4243_ ;
	wire _w4242_ ;
	wire _w4241_ ;
	wire _w4240_ ;
	wire _w4239_ ;
	wire _w4238_ ;
	wire _w4237_ ;
	wire _w4236_ ;
	wire _w4235_ ;
	wire _w4234_ ;
	wire _w4233_ ;
	wire _w4232_ ;
	wire _w4231_ ;
	wire _w4230_ ;
	wire _w4229_ ;
	wire _w4228_ ;
	wire _w4227_ ;
	wire _w4226_ ;
	wire _w4225_ ;
	wire _w4224_ ;
	wire _w4223_ ;
	wire _w4222_ ;
	wire _w4221_ ;
	wire _w4220_ ;
	wire _w4219_ ;
	wire _w4218_ ;
	wire _w4217_ ;
	wire _w4216_ ;
	wire _w4215_ ;
	wire _w4214_ ;
	wire _w4213_ ;
	wire _w4212_ ;
	wire _w4211_ ;
	wire _w4210_ ;
	wire _w4209_ ;
	wire _w4208_ ;
	wire _w4207_ ;
	wire _w4206_ ;
	wire _w4205_ ;
	wire _w4204_ ;
	wire _w4203_ ;
	wire _w4202_ ;
	wire _w4201_ ;
	wire _w4200_ ;
	wire _w4199_ ;
	wire _w4198_ ;
	wire _w4197_ ;
	wire _w4196_ ;
	wire _w4195_ ;
	wire _w4194_ ;
	wire _w4193_ ;
	wire _w4192_ ;
	wire _w4191_ ;
	wire _w4190_ ;
	wire _w4189_ ;
	wire _w4188_ ;
	wire _w4187_ ;
	wire _w4186_ ;
	wire _w4185_ ;
	wire _w4184_ ;
	wire _w4183_ ;
	wire _w4182_ ;
	wire _w4181_ ;
	wire _w4180_ ;
	wire _w4179_ ;
	wire _w4178_ ;
	wire _w4177_ ;
	wire _w4176_ ;
	wire _w4175_ ;
	wire _w4174_ ;
	wire _w4173_ ;
	wire _w4172_ ;
	wire _w4171_ ;
	wire _w4170_ ;
	wire _w4169_ ;
	wire _w4168_ ;
	wire _w4167_ ;
	wire _w4166_ ;
	wire _w4165_ ;
	wire _w4164_ ;
	wire _w4163_ ;
	wire _w4162_ ;
	wire _w4161_ ;
	wire _w4160_ ;
	wire _w4159_ ;
	wire _w4158_ ;
	wire _w4157_ ;
	wire _w4156_ ;
	wire _w4155_ ;
	wire _w4154_ ;
	wire _w4153_ ;
	wire _w4152_ ;
	wire _w4151_ ;
	wire _w4150_ ;
	wire _w4149_ ;
	wire _w4148_ ;
	wire _w4147_ ;
	wire _w4146_ ;
	wire _w4145_ ;
	wire _w4144_ ;
	wire _w4143_ ;
	wire _w4142_ ;
	wire _w4141_ ;
	wire _w4140_ ;
	wire _w4139_ ;
	wire _w4138_ ;
	wire _w4137_ ;
	wire _w4136_ ;
	wire _w4135_ ;
	wire _w4134_ ;
	wire _w4133_ ;
	wire _w4132_ ;
	wire _w4131_ ;
	wire _w4130_ ;
	wire _w4129_ ;
	wire _w4128_ ;
	wire _w4127_ ;
	wire _w4126_ ;
	wire _w4125_ ;
	wire _w4124_ ;
	wire _w4123_ ;
	wire _w4122_ ;
	wire _w4121_ ;
	wire _w4120_ ;
	wire _w4119_ ;
	wire _w4118_ ;
	wire _w4117_ ;
	wire _w4116_ ;
	wire _w4115_ ;
	wire _w4114_ ;
	wire _w4113_ ;
	wire _w4112_ ;
	wire _w4111_ ;
	wire _w4110_ ;
	wire _w4109_ ;
	wire _w4108_ ;
	wire _w4107_ ;
	wire _w4106_ ;
	wire _w4105_ ;
	wire _w4104_ ;
	wire _w4103_ ;
	wire _w4102_ ;
	wire _w4101_ ;
	wire _w4100_ ;
	wire _w4099_ ;
	wire _w4098_ ;
	wire _w4097_ ;
	wire _w4096_ ;
	wire _w4095_ ;
	wire _w4094_ ;
	wire _w4093_ ;
	wire _w4092_ ;
	wire _w4091_ ;
	wire _w4090_ ;
	wire _w4089_ ;
	wire _w4088_ ;
	wire _w4087_ ;
	wire _w4086_ ;
	wire _w4085_ ;
	wire _w4084_ ;
	wire _w4083_ ;
	wire _w4082_ ;
	wire _w4081_ ;
	wire _w4080_ ;
	wire _w4079_ ;
	wire _w4078_ ;
	wire _w4077_ ;
	wire _w4076_ ;
	wire _w4075_ ;
	wire _w4074_ ;
	wire _w4073_ ;
	wire _w4072_ ;
	wire _w4071_ ;
	wire _w4070_ ;
	wire _w4069_ ;
	wire _w4068_ ;
	wire _w4067_ ;
	wire _w4066_ ;
	wire _w4065_ ;
	wire _w4064_ ;
	wire _w4063_ ;
	wire _w4062_ ;
	wire _w4061_ ;
	wire _w4060_ ;
	wire _w4059_ ;
	wire _w4058_ ;
	wire _w4057_ ;
	wire _w4056_ ;
	wire _w4055_ ;
	wire _w4054_ ;
	wire _w4053_ ;
	wire _w4052_ ;
	wire _w4051_ ;
	wire _w4050_ ;
	wire _w4049_ ;
	wire _w4048_ ;
	wire _w4047_ ;
	wire _w4046_ ;
	wire _w4045_ ;
	wire _w4044_ ;
	wire _w4043_ ;
	wire _w4042_ ;
	wire _w4041_ ;
	wire _w4040_ ;
	wire _w4039_ ;
	wire _w4038_ ;
	wire _w4037_ ;
	wire _w4036_ ;
	wire _w4035_ ;
	wire _w4034_ ;
	wire _w4033_ ;
	wire _w4032_ ;
	wire _w4031_ ;
	wire _w4030_ ;
	wire _w4029_ ;
	wire _w4028_ ;
	wire _w4027_ ;
	wire _w4026_ ;
	wire _w4025_ ;
	wire _w4024_ ;
	wire _w4023_ ;
	wire _w4022_ ;
	wire _w4021_ ;
	wire _w4020_ ;
	wire _w4019_ ;
	wire _w4018_ ;
	wire _w4017_ ;
	wire _w4016_ ;
	wire _w4015_ ;
	wire _w4014_ ;
	wire _w4013_ ;
	wire _w4012_ ;
	wire _w4011_ ;
	wire _w4010_ ;
	wire _w4009_ ;
	wire _w4008_ ;
	wire _w4007_ ;
	wire _w4006_ ;
	wire _w4005_ ;
	wire _w4004_ ;
	wire _w4003_ ;
	wire _w4002_ ;
	wire _w4001_ ;
	wire _w4000_ ;
	wire _w3999_ ;
	wire _w3998_ ;
	wire _w3997_ ;
	wire _w3996_ ;
	wire _w3995_ ;
	wire _w3994_ ;
	wire _w3993_ ;
	wire _w3992_ ;
	wire _w3991_ ;
	wire _w3990_ ;
	wire _w3989_ ;
	wire _w3988_ ;
	wire _w3987_ ;
	wire _w3986_ ;
	wire _w3985_ ;
	wire _w3984_ ;
	wire _w3983_ ;
	wire _w3982_ ;
	wire _w3981_ ;
	wire _w3980_ ;
	wire _w3979_ ;
	wire _w3978_ ;
	wire _w3977_ ;
	wire _w3976_ ;
	wire _w3975_ ;
	wire _w3974_ ;
	wire _w3973_ ;
	wire _w3972_ ;
	wire _w3971_ ;
	wire _w3970_ ;
	wire _w3969_ ;
	wire _w3968_ ;
	wire _w3967_ ;
	wire _w3966_ ;
	wire _w3965_ ;
	wire _w3964_ ;
	wire _w3963_ ;
	wire _w3962_ ;
	wire _w3961_ ;
	wire _w3960_ ;
	wire _w3959_ ;
	wire _w3958_ ;
	wire _w3957_ ;
	wire _w3956_ ;
	wire _w3955_ ;
	wire _w3954_ ;
	wire _w3953_ ;
	wire _w3952_ ;
	wire _w3951_ ;
	wire _w3950_ ;
	wire _w3949_ ;
	wire _w3948_ ;
	wire _w3947_ ;
	wire _w3946_ ;
	wire _w3945_ ;
	wire _w3944_ ;
	wire _w3943_ ;
	wire _w3942_ ;
	wire _w3941_ ;
	wire _w3940_ ;
	wire _w3939_ ;
	wire _w3938_ ;
	wire _w3937_ ;
	wire _w3936_ ;
	wire _w3935_ ;
	wire _w3934_ ;
	wire _w3933_ ;
	wire _w3932_ ;
	wire _w3931_ ;
	wire _w3930_ ;
	wire _w3929_ ;
	wire _w3928_ ;
	wire _w3927_ ;
	wire _w3926_ ;
	wire _w3925_ ;
	wire _w3924_ ;
	wire _w3923_ ;
	wire _w3922_ ;
	wire _w3921_ ;
	wire _w3920_ ;
	wire _w3919_ ;
	wire _w3918_ ;
	wire _w3917_ ;
	wire _w3916_ ;
	wire _w3915_ ;
	wire _w3914_ ;
	wire _w3913_ ;
	wire _w3912_ ;
	wire _w3911_ ;
	wire _w3910_ ;
	wire _w3909_ ;
	wire _w3908_ ;
	wire _w3907_ ;
	wire _w3906_ ;
	wire _w3905_ ;
	wire _w3904_ ;
	wire _w3903_ ;
	wire _w3902_ ;
	wire _w3901_ ;
	wire _w3900_ ;
	wire _w3899_ ;
	wire _w3898_ ;
	wire _w3897_ ;
	wire _w3896_ ;
	wire _w3895_ ;
	wire _w3894_ ;
	wire _w3893_ ;
	wire _w3892_ ;
	wire _w3891_ ;
	wire _w3890_ ;
	wire _w3889_ ;
	wire _w3888_ ;
	wire _w3887_ ;
	wire _w3886_ ;
	wire _w3885_ ;
	wire _w3884_ ;
	wire _w3883_ ;
	wire _w3882_ ;
	wire _w3881_ ;
	wire _w3880_ ;
	wire _w3879_ ;
	wire _w3878_ ;
	wire _w3877_ ;
	wire _w3876_ ;
	wire _w3875_ ;
	wire _w3874_ ;
	wire _w3873_ ;
	wire _w3872_ ;
	wire _w3871_ ;
	wire _w3870_ ;
	wire _w3869_ ;
	wire _w3868_ ;
	wire _w3867_ ;
	wire _w3866_ ;
	wire _w3865_ ;
	wire _w3864_ ;
	wire _w3863_ ;
	wire _w3862_ ;
	wire _w3861_ ;
	wire _w3860_ ;
	wire _w3859_ ;
	wire _w3858_ ;
	wire _w3857_ ;
	wire _w3856_ ;
	wire _w3855_ ;
	wire _w3854_ ;
	wire _w3853_ ;
	wire _w3852_ ;
	wire _w3851_ ;
	wire _w3850_ ;
	wire _w3849_ ;
	wire _w3848_ ;
	wire _w3847_ ;
	wire _w3846_ ;
	wire _w3845_ ;
	wire _w3844_ ;
	wire _w3843_ ;
	wire _w3842_ ;
	wire _w3841_ ;
	wire _w3840_ ;
	wire _w3839_ ;
	wire _w3838_ ;
	wire _w3837_ ;
	wire _w3836_ ;
	wire _w3835_ ;
	wire _w3834_ ;
	wire _w3833_ ;
	wire _w3832_ ;
	wire _w3831_ ;
	wire _w3830_ ;
	wire _w3829_ ;
	wire _w3828_ ;
	wire _w3827_ ;
	wire _w3826_ ;
	wire _w3825_ ;
	wire _w3824_ ;
	wire _w3823_ ;
	wire _w3822_ ;
	wire _w3821_ ;
	wire _w3820_ ;
	wire _w3819_ ;
	wire _w3818_ ;
	wire _w3817_ ;
	wire _w3816_ ;
	wire _w3815_ ;
	wire _w3814_ ;
	wire _w3813_ ;
	wire _w3812_ ;
	wire _w3811_ ;
	wire _w3810_ ;
	wire _w3809_ ;
	wire _w3808_ ;
	wire _w3807_ ;
	wire _w3806_ ;
	wire _w3805_ ;
	wire _w3804_ ;
	wire _w3803_ ;
	wire _w3802_ ;
	wire _w3801_ ;
	wire _w3800_ ;
	wire _w3799_ ;
	wire _w3798_ ;
	wire _w3797_ ;
	wire _w3796_ ;
	wire _w3795_ ;
	wire _w3794_ ;
	wire _w3793_ ;
	wire _w3792_ ;
	wire _w3791_ ;
	wire _w3790_ ;
	wire _w3789_ ;
	wire _w3788_ ;
	wire _w3787_ ;
	wire _w3786_ ;
	wire _w3785_ ;
	wire _w3784_ ;
	wire _w3783_ ;
	wire _w3782_ ;
	wire _w3781_ ;
	wire _w3780_ ;
	wire _w3779_ ;
	wire _w3778_ ;
	wire _w3777_ ;
	wire _w3776_ ;
	wire _w3775_ ;
	wire _w3774_ ;
	wire _w3773_ ;
	wire _w3772_ ;
	wire _w3771_ ;
	wire _w3770_ ;
	wire _w3769_ ;
	wire _w3768_ ;
	wire _w3767_ ;
	wire _w3766_ ;
	wire _w3765_ ;
	wire _w3764_ ;
	wire _w3763_ ;
	wire _w3762_ ;
	wire _w3761_ ;
	wire _w3760_ ;
	wire _w3759_ ;
	wire _w3758_ ;
	wire _w3757_ ;
	wire _w3756_ ;
	wire _w3755_ ;
	wire _w3754_ ;
	wire _w3753_ ;
	wire _w3752_ ;
	wire _w3751_ ;
	wire _w3750_ ;
	wire _w3749_ ;
	wire _w3748_ ;
	wire _w3747_ ;
	wire _w3746_ ;
	wire _w3745_ ;
	wire _w3744_ ;
	wire _w3743_ ;
	wire _w3742_ ;
	wire _w3741_ ;
	wire _w3740_ ;
	wire _w3739_ ;
	wire _w3738_ ;
	wire _w3737_ ;
	wire _w3736_ ;
	wire _w3735_ ;
	wire _w3734_ ;
	wire _w3733_ ;
	wire _w3732_ ;
	wire _w3731_ ;
	wire _w3730_ ;
	wire _w3729_ ;
	wire _w3728_ ;
	wire _w3727_ ;
	wire _w3726_ ;
	wire _w3725_ ;
	wire _w3724_ ;
	wire _w3723_ ;
	wire _w3722_ ;
	wire _w3721_ ;
	wire _w3720_ ;
	wire _w3719_ ;
	wire _w3718_ ;
	wire _w3717_ ;
	wire _w3716_ ;
	wire _w3715_ ;
	wire _w3714_ ;
	wire _w3713_ ;
	wire _w3712_ ;
	wire _w3711_ ;
	wire _w3710_ ;
	wire _w3709_ ;
	wire _w3708_ ;
	wire _w3707_ ;
	wire _w3706_ ;
	wire _w3705_ ;
	wire _w3704_ ;
	wire _w3703_ ;
	wire _w3702_ ;
	wire _w3701_ ;
	wire _w3700_ ;
	wire _w3699_ ;
	wire _w3698_ ;
	wire _w3697_ ;
	wire _w3696_ ;
	wire _w3695_ ;
	wire _w3694_ ;
	wire _w3693_ ;
	wire _w3692_ ;
	wire _w3691_ ;
	wire _w3690_ ;
	wire _w3689_ ;
	wire _w3688_ ;
	wire _w3687_ ;
	wire _w3686_ ;
	wire _w3685_ ;
	wire _w3684_ ;
	wire _w3683_ ;
	wire _w3682_ ;
	wire _w3681_ ;
	wire _w3680_ ;
	wire _w3679_ ;
	wire _w3678_ ;
	wire _w3677_ ;
	wire _w3676_ ;
	wire _w3675_ ;
	wire _w3674_ ;
	wire _w3673_ ;
	wire _w3672_ ;
	wire _w3671_ ;
	wire _w3670_ ;
	wire _w3669_ ;
	wire _w3668_ ;
	wire _w3667_ ;
	wire _w3666_ ;
	wire _w3665_ ;
	wire _w3664_ ;
	wire _w3663_ ;
	wire _w3662_ ;
	wire _w3661_ ;
	wire _w3660_ ;
	wire _w3659_ ;
	wire _w3658_ ;
	wire _w3657_ ;
	wire _w3656_ ;
	wire _w3655_ ;
	wire _w3654_ ;
	wire _w3653_ ;
	wire _w3652_ ;
	wire _w3651_ ;
	wire _w3650_ ;
	wire _w3649_ ;
	wire _w3648_ ;
	wire _w3647_ ;
	wire _w3646_ ;
	wire _w3645_ ;
	wire _w3644_ ;
	wire _w3643_ ;
	wire _w3642_ ;
	wire _w3641_ ;
	wire _w3640_ ;
	wire _w3639_ ;
	wire _w3638_ ;
	wire _w3637_ ;
	wire _w3636_ ;
	wire _w3635_ ;
	wire _w3634_ ;
	wire _w3633_ ;
	wire _w3632_ ;
	wire _w3631_ ;
	wire _w3630_ ;
	wire _w3629_ ;
	wire _w3628_ ;
	wire _w3627_ ;
	wire _w3626_ ;
	wire _w3625_ ;
	wire _w3624_ ;
	wire _w3623_ ;
	wire _w3622_ ;
	wire _w3621_ ;
	wire _w3620_ ;
	wire _w3619_ ;
	wire _w3618_ ;
	wire _w3617_ ;
	wire _w3616_ ;
	wire _w3615_ ;
	wire _w3614_ ;
	wire _w3613_ ;
	wire _w3612_ ;
	wire _w3611_ ;
	wire _w3610_ ;
	wire _w3609_ ;
	wire _w3608_ ;
	wire _w3607_ ;
	wire _w3606_ ;
	wire _w3605_ ;
	wire _w3604_ ;
	wire _w3603_ ;
	wire _w3602_ ;
	wire _w3601_ ;
	wire _w3600_ ;
	wire _w3599_ ;
	wire _w3598_ ;
	wire _w3597_ ;
	wire _w3596_ ;
	wire _w3595_ ;
	wire _w3594_ ;
	wire _w3593_ ;
	wire _w3592_ ;
	wire _w3591_ ;
	wire _w3590_ ;
	wire _w3589_ ;
	wire _w3588_ ;
	wire _w3587_ ;
	wire _w3586_ ;
	wire _w3585_ ;
	wire _w3584_ ;
	wire _w3583_ ;
	wire _w3582_ ;
	wire _w3581_ ;
	wire _w3580_ ;
	wire _w3579_ ;
	wire _w3578_ ;
	wire _w3577_ ;
	wire _w3576_ ;
	wire _w3575_ ;
	wire _w3574_ ;
	wire _w3573_ ;
	wire _w3572_ ;
	wire _w3571_ ;
	wire _w3570_ ;
	wire _w3569_ ;
	wire _w3568_ ;
	wire _w3567_ ;
	wire _w3566_ ;
	wire _w3565_ ;
	wire _w3564_ ;
	wire _w3563_ ;
	wire _w3562_ ;
	wire _w3561_ ;
	wire _w3560_ ;
	wire _w3559_ ;
	wire _w3558_ ;
	wire _w3557_ ;
	wire _w3556_ ;
	wire _w3555_ ;
	wire _w3554_ ;
	wire _w3553_ ;
	wire _w3552_ ;
	wire _w3551_ ;
	wire _w3550_ ;
	wire _w3549_ ;
	wire _w3548_ ;
	wire _w3547_ ;
	wire _w3546_ ;
	wire _w3545_ ;
	wire _w3544_ ;
	wire _w3543_ ;
	wire _w3542_ ;
	wire _w3541_ ;
	wire _w3540_ ;
	wire _w3539_ ;
	wire _w3538_ ;
	wire _w3537_ ;
	wire _w3536_ ;
	wire _w3535_ ;
	wire _w3534_ ;
	wire _w3533_ ;
	wire _w3532_ ;
	wire _w3531_ ;
	wire _w3530_ ;
	wire _w3529_ ;
	wire _w3528_ ;
	wire _w3527_ ;
	wire _w3526_ ;
	wire _w3525_ ;
	wire _w3524_ ;
	wire _w3523_ ;
	wire _w3522_ ;
	wire _w3521_ ;
	wire _w3520_ ;
	wire _w3519_ ;
	wire _w3518_ ;
	wire _w3517_ ;
	wire _w3516_ ;
	wire _w3515_ ;
	wire _w3514_ ;
	wire _w3513_ ;
	wire _w3512_ ;
	wire _w3511_ ;
	wire _w3510_ ;
	wire _w3509_ ;
	wire _w3508_ ;
	wire _w3507_ ;
	wire _w3506_ ;
	wire _w3505_ ;
	wire _w3504_ ;
	wire _w3503_ ;
	wire _w3502_ ;
	wire _w3501_ ;
	wire _w3500_ ;
	wire _w3499_ ;
	wire _w3498_ ;
	wire _w3497_ ;
	wire _w3496_ ;
	wire _w3495_ ;
	wire _w3494_ ;
	wire _w3493_ ;
	wire _w3492_ ;
	wire _w3491_ ;
	wire _w3490_ ;
	wire _w3489_ ;
	wire _w3488_ ;
	wire _w3487_ ;
	wire _w3486_ ;
	wire _w3485_ ;
	wire _w3484_ ;
	wire _w3483_ ;
	wire _w3482_ ;
	wire _w3481_ ;
	wire _w3480_ ;
	wire _w3479_ ;
	wire _w3478_ ;
	wire _w3477_ ;
	wire _w3476_ ;
	wire _w3475_ ;
	wire _w3474_ ;
	wire _w3473_ ;
	wire _w3472_ ;
	wire _w3471_ ;
	wire _w3470_ ;
	wire _w3469_ ;
	wire _w3468_ ;
	wire _w3467_ ;
	wire _w3466_ ;
	wire _w3465_ ;
	wire _w3464_ ;
	wire _w3463_ ;
	wire _w3462_ ;
	wire _w3461_ ;
	wire _w3460_ ;
	wire _w3459_ ;
	wire _w3458_ ;
	wire _w3457_ ;
	wire _w3456_ ;
	wire _w3455_ ;
	wire _w3454_ ;
	wire _w3453_ ;
	wire _w3452_ ;
	wire _w3451_ ;
	wire _w3450_ ;
	wire _w3449_ ;
	wire _w3448_ ;
	wire _w3447_ ;
	wire _w3446_ ;
	wire _w3445_ ;
	wire _w3444_ ;
	wire _w3443_ ;
	wire _w3442_ ;
	wire _w3441_ ;
	wire _w3440_ ;
	wire _w3439_ ;
	wire _w3438_ ;
	wire _w3437_ ;
	wire _w3436_ ;
	wire _w3435_ ;
	wire _w3434_ ;
	wire _w3433_ ;
	wire _w3432_ ;
	wire _w3431_ ;
	wire _w3430_ ;
	wire _w3429_ ;
	wire _w3428_ ;
	wire _w3427_ ;
	wire _w3426_ ;
	wire _w3425_ ;
	wire _w3424_ ;
	wire _w3423_ ;
	wire _w3422_ ;
	wire _w3421_ ;
	wire _w3420_ ;
	wire _w3419_ ;
	wire _w3418_ ;
	wire _w3417_ ;
	wire _w3416_ ;
	wire _w3415_ ;
	wire _w3414_ ;
	wire _w3413_ ;
	wire _w3412_ ;
	wire _w3411_ ;
	wire _w3410_ ;
	wire _w3409_ ;
	wire _w3408_ ;
	wire _w3407_ ;
	wire _w3406_ ;
	wire _w3405_ ;
	wire _w3404_ ;
	wire _w3403_ ;
	wire _w3402_ ;
	wire _w3401_ ;
	wire _w3400_ ;
	wire _w3399_ ;
	wire _w3398_ ;
	wire _w3397_ ;
	wire _w3396_ ;
	wire _w3395_ ;
	wire _w3394_ ;
	wire _w3393_ ;
	wire _w3392_ ;
	wire _w3391_ ;
	wire _w3390_ ;
	wire _w3389_ ;
	wire _w3388_ ;
	wire _w3387_ ;
	wire _w3386_ ;
	wire _w3385_ ;
	wire _w3384_ ;
	wire _w3383_ ;
	wire _w3382_ ;
	wire _w3381_ ;
	wire _w3380_ ;
	wire _w3379_ ;
	wire _w3378_ ;
	wire _w3377_ ;
	wire _w3376_ ;
	wire _w3375_ ;
	wire _w3374_ ;
	wire _w3373_ ;
	wire _w3372_ ;
	wire _w3371_ ;
	wire _w3370_ ;
	wire _w3369_ ;
	wire _w3368_ ;
	wire _w3367_ ;
	wire _w3366_ ;
	wire _w3365_ ;
	wire _w3364_ ;
	wire _w3363_ ;
	wire _w3362_ ;
	wire _w3361_ ;
	wire _w3360_ ;
	wire _w3359_ ;
	wire _w3358_ ;
	wire _w3357_ ;
	wire _w3356_ ;
	wire _w3355_ ;
	wire _w3354_ ;
	wire _w3353_ ;
	wire _w3352_ ;
	wire _w3351_ ;
	wire _w3350_ ;
	wire _w3349_ ;
	wire _w3348_ ;
	wire _w3347_ ;
	wire _w3346_ ;
	wire _w3345_ ;
	wire _w3344_ ;
	wire _w3343_ ;
	wire _w3342_ ;
	wire _w3341_ ;
	wire _w3340_ ;
	wire _w3339_ ;
	wire _w3338_ ;
	wire _w3337_ ;
	wire _w3336_ ;
	wire _w3335_ ;
	wire _w3334_ ;
	wire _w3333_ ;
	wire _w3332_ ;
	wire _w3331_ ;
	wire _w3330_ ;
	wire _w3329_ ;
	wire _w3328_ ;
	wire _w3327_ ;
	wire _w3326_ ;
	wire _w3325_ ;
	wire _w3324_ ;
	wire _w3323_ ;
	wire _w3322_ ;
	wire _w3321_ ;
	wire _w3320_ ;
	wire _w3319_ ;
	wire _w3318_ ;
	wire _w3317_ ;
	wire _w3316_ ;
	wire _w3315_ ;
	wire _w3314_ ;
	wire _w3313_ ;
	wire _w3312_ ;
	wire _w3311_ ;
	wire _w3310_ ;
	wire _w3309_ ;
	wire _w3308_ ;
	wire _w3307_ ;
	wire _w3306_ ;
	wire _w3305_ ;
	wire _w3304_ ;
	wire _w3303_ ;
	wire _w3302_ ;
	wire _w3301_ ;
	wire _w3300_ ;
	wire _w3299_ ;
	wire _w3298_ ;
	wire _w3297_ ;
	wire _w3296_ ;
	wire _w3295_ ;
	wire _w3294_ ;
	wire _w3293_ ;
	wire _w3292_ ;
	wire _w3291_ ;
	wire _w3290_ ;
	wire _w3289_ ;
	wire _w3288_ ;
	wire _w3287_ ;
	wire _w3286_ ;
	wire _w2037_ ;
	wire _w2036_ ;
	wire _w2035_ ;
	wire _w2034_ ;
	wire _w2033_ ;
	wire _w2032_ ;
	wire _w2031_ ;
	wire _w2030_ ;
	wire _w2029_ ;
	wire _w2028_ ;
	wire _w2027_ ;
	wire _w2026_ ;
	wire _w2025_ ;
	wire _w2024_ ;
	wire _w2023_ ;
	wire _w2022_ ;
	wire _w2021_ ;
	wire _w2020_ ;
	wire _w2019_ ;
	wire _w2018_ ;
	wire _w2017_ ;
	wire _w2016_ ;
	wire _w2015_ ;
	wire _w2014_ ;
	wire _w2013_ ;
	wire _w2012_ ;
	wire _w2011_ ;
	wire _w2010_ ;
	wire _w2009_ ;
	wire _w2008_ ;
	wire _w2007_ ;
	wire _w2006_ ;
	wire _w2005_ ;
	wire _w2004_ ;
	wire _w2003_ ;
	wire _w2002_ ;
	wire _w2001_ ;
	wire _w2000_ ;
	wire _w1999_ ;
	wire _w1998_ ;
	wire _w1997_ ;
	wire _w1996_ ;
	wire _w1995_ ;
	wire _w1994_ ;
	wire _w1993_ ;
	wire _w1992_ ;
	wire _w1991_ ;
	wire _w1990_ ;
	wire _w1989_ ;
	wire _w1988_ ;
	wire _w1987_ ;
	wire _w1986_ ;
	wire _w1985_ ;
	wire _w1984_ ;
	wire _w1983_ ;
	wire _w1982_ ;
	wire _w1981_ ;
	wire _w1980_ ;
	wire _w1979_ ;
	wire _w1978_ ;
	wire _w1977_ ;
	wire _w1976_ ;
	wire _w1975_ ;
	wire _w1974_ ;
	wire _w1973_ ;
	wire _w1972_ ;
	wire _w1971_ ;
	wire _w1970_ ;
	wire _w1969_ ;
	wire _w1968_ ;
	wire _w1967_ ;
	wire _w1966_ ;
	wire _w1965_ ;
	wire _w1964_ ;
	wire _w1963_ ;
	wire _w1962_ ;
	wire _w1961_ ;
	wire _w1960_ ;
	wire _w1959_ ;
	wire _w1958_ ;
	wire _w1957_ ;
	wire _w1956_ ;
	wire _w1955_ ;
	wire _w1954_ ;
	wire _w1953_ ;
	wire _w1952_ ;
	wire _w1951_ ;
	wire _w1950_ ;
	wire _w1949_ ;
	wire _w1948_ ;
	wire _w1947_ ;
	wire _w1946_ ;
	wire _w1945_ ;
	wire _w1944_ ;
	wire _w1943_ ;
	wire _w1942_ ;
	wire _w1941_ ;
	wire _w1940_ ;
	wire _w1939_ ;
	wire _w1938_ ;
	wire _w1937_ ;
	wire _w1936_ ;
	wire _w1935_ ;
	wire _w1934_ ;
	wire _w1933_ ;
	wire _w1932_ ;
	wire _w1931_ ;
	wire _w1930_ ;
	wire _w1929_ ;
	wire _w1928_ ;
	wire _w1927_ ;
	wire _w1926_ ;
	wire _w1925_ ;
	wire _w1924_ ;
	wire _w1923_ ;
	wire _w1922_ ;
	wire _w1921_ ;
	wire _w1920_ ;
	wire _w1919_ ;
	wire _w1918_ ;
	wire _w1917_ ;
	wire _w1916_ ;
	wire _w1915_ ;
	wire _w1914_ ;
	wire _w1913_ ;
	wire _w1912_ ;
	wire _w1911_ ;
	wire _w1910_ ;
	wire _w1909_ ;
	wire _w1908_ ;
	wire _w1907_ ;
	wire _w1906_ ;
	wire _w1905_ ;
	wire _w1904_ ;
	wire _w1903_ ;
	wire _w1902_ ;
	wire _w1901_ ;
	wire _w1900_ ;
	wire _w1899_ ;
	wire _w1898_ ;
	wire _w1897_ ;
	wire _w1896_ ;
	wire _w1895_ ;
	wire _w1894_ ;
	wire _w1893_ ;
	wire _w1892_ ;
	wire _w1891_ ;
	wire _w1890_ ;
	wire _w1889_ ;
	wire _w1888_ ;
	wire _w1887_ ;
	wire _w1886_ ;
	wire _w1885_ ;
	wire _w1884_ ;
	wire _w1883_ ;
	wire _w1882_ ;
	wire _w1881_ ;
	wire _w1880_ ;
	wire _w1879_ ;
	wire _w1878_ ;
	wire _w1877_ ;
	wire _w1876_ ;
	wire _w1875_ ;
	wire _w1874_ ;
	wire _w1873_ ;
	wire _w1872_ ;
	wire _w1871_ ;
	wire _w1870_ ;
	wire _w1869_ ;
	wire _w1868_ ;
	wire _w1867_ ;
	wire _w1866_ ;
	wire _w1865_ ;
	wire _w1864_ ;
	wire _w1863_ ;
	wire _w1862_ ;
	wire _w1861_ ;
	wire _w1860_ ;
	wire _w1859_ ;
	wire _w1858_ ;
	wire _w1857_ ;
	wire _w1856_ ;
	wire _w1855_ ;
	wire _w1854_ ;
	wire _w1853_ ;
	wire _w1852_ ;
	wire _w1851_ ;
	wire _w1850_ ;
	wire _w1849_ ;
	wire _w1848_ ;
	wire _w1847_ ;
	wire _w1846_ ;
	wire _w1845_ ;
	wire _w1844_ ;
	wire _w1843_ ;
	wire _w1842_ ;
	wire _w1841_ ;
	wire _w1840_ ;
	wire _w1839_ ;
	wire _w1838_ ;
	wire _w1837_ ;
	wire _w1836_ ;
	wire _w1835_ ;
	wire _w1834_ ;
	wire _w1833_ ;
	wire _w1832_ ;
	wire _w1831_ ;
	wire _w1830_ ;
	wire _w1829_ ;
	wire _w1828_ ;
	wire _w1827_ ;
	wire _w1826_ ;
	wire _w1825_ ;
	wire _w1824_ ;
	wire _w1823_ ;
	wire _w1822_ ;
	wire _w1821_ ;
	wire _w1820_ ;
	wire _w1819_ ;
	wire _w1818_ ;
	wire _w1817_ ;
	wire _w1816_ ;
	wire _w1815_ ;
	wire _w1814_ ;
	wire _w1813_ ;
	wire _w1812_ ;
	wire _w1811_ ;
	wire _w1810_ ;
	wire _w1809_ ;
	wire _w1808_ ;
	wire _w1807_ ;
	wire _w1806_ ;
	wire _w1805_ ;
	wire _w1804_ ;
	wire _w1803_ ;
	wire _w1802_ ;
	wire _w1801_ ;
	wire _w1800_ ;
	wire _w1799_ ;
	wire _w1798_ ;
	wire _w1797_ ;
	wire _w1796_ ;
	wire _w1795_ ;
	wire _w1794_ ;
	wire _w1793_ ;
	wire _w1792_ ;
	wire _w1791_ ;
	wire _w1790_ ;
	wire _w1789_ ;
	wire _w1788_ ;
	wire _w1787_ ;
	wire _w1786_ ;
	wire _w1785_ ;
	wire _w1784_ ;
	wire _w1783_ ;
	wire _w1782_ ;
	wire _w1781_ ;
	wire _w1780_ ;
	wire _w1779_ ;
	wire _w1778_ ;
	wire _w1777_ ;
	wire _w1776_ ;
	wire _w1775_ ;
	wire _w1774_ ;
	wire _w1773_ ;
	wire _w1772_ ;
	wire _w1771_ ;
	wire _w1770_ ;
	wire _w1769_ ;
	wire _w1768_ ;
	wire _w1767_ ;
	wire _w1766_ ;
	wire _w1765_ ;
	wire _w1764_ ;
	wire _w1763_ ;
	wire _w1762_ ;
	wire _w1761_ ;
	wire _w1760_ ;
	wire _w1759_ ;
	wire _w1758_ ;
	wire _w1757_ ;
	wire _w1756_ ;
	wire _w1755_ ;
	wire _w1754_ ;
	wire _w1753_ ;
	wire _w1752_ ;
	wire _w1751_ ;
	wire _w1750_ ;
	wire _w1749_ ;
	wire _w1748_ ;
	wire _w1747_ ;
	wire _w1746_ ;
	wire _w1745_ ;
	wire _w1744_ ;
	wire _w1743_ ;
	wire _w1742_ ;
	wire _w1741_ ;
	wire _w1740_ ;
	wire _w1739_ ;
	wire _w1738_ ;
	wire _w1737_ ;
	wire _w1736_ ;
	wire _w1735_ ;
	wire _w1734_ ;
	wire _w1733_ ;
	wire _w1732_ ;
	wire _w1731_ ;
	wire _w1730_ ;
	wire _w1729_ ;
	wire _w1728_ ;
	wire _w1727_ ;
	wire _w1726_ ;
	wire _w1725_ ;
	wire _w1724_ ;
	wire _w1723_ ;
	wire _w1722_ ;
	wire _w1721_ ;
	wire _w1720_ ;
	wire _w1719_ ;
	wire _w1718_ ;
	wire _w1717_ ;
	wire _w1716_ ;
	wire _w1715_ ;
	wire _w1714_ ;
	wire _w1713_ ;
	wire _w1712_ ;
	wire _w1711_ ;
	wire _w1710_ ;
	wire _w1709_ ;
	wire _w1708_ ;
	wire _w1707_ ;
	wire _w1706_ ;
	wire _w1705_ ;
	wire _w1704_ ;
	wire _w1703_ ;
	wire _w1702_ ;
	wire _w1701_ ;
	wire _w1700_ ;
	wire _w1699_ ;
	wire _w1698_ ;
	wire _w1697_ ;
	wire _w1696_ ;
	wire _w1695_ ;
	wire _w1694_ ;
	wire _w1693_ ;
	wire _w1692_ ;
	wire _w1691_ ;
	wire _w1690_ ;
	wire _w1689_ ;
	wire _w1688_ ;
	wire _w1687_ ;
	wire _w1686_ ;
	wire _w1685_ ;
	wire _w1684_ ;
	wire _w1683_ ;
	wire _w1682_ ;
	wire _w1681_ ;
	wire _w1680_ ;
	wire _w1679_ ;
	wire _w1678_ ;
	wire _w1677_ ;
	wire _w1676_ ;
	wire _w1675_ ;
	wire _w1674_ ;
	wire _w1673_ ;
	wire _w1672_ ;
	wire _w1671_ ;
	wire _w1670_ ;
	wire _w1669_ ;
	wire _w1668_ ;
	wire _w1667_ ;
	wire _w1666_ ;
	wire _w1665_ ;
	wire _w1664_ ;
	wire _w1663_ ;
	wire _w1662_ ;
	wire _w1661_ ;
	wire _w1660_ ;
	wire _w1659_ ;
	wire _w1658_ ;
	wire _w1657_ ;
	wire _w1656_ ;
	wire _w1655_ ;
	wire _w1654_ ;
	wire _w1653_ ;
	wire _w1652_ ;
	wire _w1651_ ;
	wire _w1650_ ;
	wire _w1649_ ;
	wire _w1648_ ;
	wire _w1647_ ;
	wire _w1646_ ;
	wire _w1645_ ;
	wire _w1644_ ;
	wire _w1643_ ;
	wire _w1642_ ;
	wire _w1641_ ;
	wire _w1640_ ;
	wire _w1639_ ;
	wire _w1638_ ;
	wire _w1637_ ;
	wire _w1636_ ;
	wire _w1635_ ;
	wire _w1634_ ;
	wire _w1633_ ;
	wire _w1632_ ;
	wire _w1631_ ;
	wire _w1630_ ;
	wire _w1629_ ;
	wire _w1628_ ;
	wire _w1627_ ;
	wire _w1626_ ;
	wire _w1625_ ;
	wire _w1624_ ;
	wire _w1623_ ;
	wire _w1622_ ;
	wire _w1621_ ;
	wire _w1620_ ;
	wire _w1619_ ;
	wire _w1618_ ;
	wire _w1617_ ;
	wire _w1616_ ;
	wire _w1615_ ;
	wire _w1614_ ;
	wire _w1613_ ;
	wire _w1612_ ;
	wire _w1611_ ;
	wire _w1610_ ;
	wire _w1609_ ;
	wire _w1608_ ;
	wire _w1607_ ;
	wire _w1606_ ;
	wire _w1605_ ;
	wire _w1604_ ;
	wire _w1603_ ;
	wire _w1602_ ;
	wire _w1601_ ;
	wire _w1600_ ;
	wire _w1599_ ;
	wire _w1598_ ;
	wire _w1597_ ;
	wire _w1596_ ;
	wire _w1595_ ;
	wire _w1594_ ;
	wire _w1593_ ;
	wire _w1592_ ;
	wire _w1591_ ;
	wire _w1590_ ;
	wire _w1589_ ;
	wire _w1588_ ;
	wire _w1587_ ;
	wire _w1586_ ;
	wire _w1585_ ;
	wire _w1584_ ;
	wire _w1583_ ;
	wire _w1582_ ;
	wire _w1581_ ;
	wire _w1580_ ;
	wire _w1579_ ;
	wire _w1578_ ;
	wire _w1577_ ;
	wire _w1576_ ;
	wire _w1575_ ;
	wire _w1574_ ;
	wire _w1573_ ;
	wire _w1572_ ;
	wire _w1571_ ;
	wire _w1570_ ;
	wire _w1569_ ;
	wire _w1568_ ;
	wire _w1567_ ;
	wire _w1566_ ;
	wire _w1565_ ;
	wire _w1564_ ;
	wire _w1563_ ;
	wire _w1562_ ;
	wire _w1561_ ;
	wire _w1560_ ;
	wire _w1559_ ;
	wire _w1558_ ;
	wire _w1557_ ;
	wire _w1556_ ;
	wire _w1555_ ;
	wire _w1554_ ;
	wire _w1553_ ;
	wire _w1552_ ;
	wire _w1551_ ;
	wire _w1550_ ;
	wire _w1549_ ;
	wire _w1548_ ;
	wire _w1547_ ;
	wire _w1546_ ;
	wire _w1545_ ;
	wire _w1544_ ;
	wire _w1543_ ;
	wire _w1542_ ;
	wire _w1541_ ;
	wire _w1540_ ;
	wire _w1539_ ;
	wire _w1538_ ;
	wire _w1537_ ;
	wire _w1536_ ;
	wire _w1535_ ;
	wire _w1534_ ;
	wire _w1533_ ;
	wire _w1532_ ;
	wire _w1531_ ;
	wire _w1530_ ;
	wire _w1529_ ;
	wire _w1528_ ;
	wire _w1527_ ;
	wire _w1526_ ;
	wire _w1525_ ;
	wire _w1524_ ;
	wire _w1523_ ;
	wire _w1522_ ;
	wire _w1521_ ;
	wire _w1520_ ;
	wire _w1519_ ;
	wire _w1518_ ;
	wire _w1517_ ;
	wire _w1516_ ;
	wire _w1515_ ;
	wire _w1514_ ;
	wire _w1513_ ;
	wire _w1512_ ;
	wire _w1511_ ;
	wire _w1510_ ;
	wire _w1509_ ;
	wire _w1508_ ;
	wire _w1507_ ;
	wire _w1506_ ;
	wire _w1505_ ;
	wire _w1504_ ;
	wire _w1503_ ;
	wire _w1502_ ;
	wire _w1501_ ;
	wire _w1500_ ;
	wire _w1499_ ;
	wire _w1498_ ;
	wire _w1497_ ;
	wire _w1496_ ;
	wire _w1495_ ;
	wire _w1494_ ;
	wire _w1493_ ;
	wire _w1492_ ;
	wire _w1491_ ;
	wire _w1490_ ;
	wire _w1489_ ;
	wire _w1488_ ;
	wire _w1487_ ;
	wire _w1486_ ;
	wire _w1485_ ;
	wire _w1484_ ;
	wire _w1483_ ;
	wire _w1482_ ;
	wire _w1481_ ;
	wire _w1480_ ;
	wire _w1479_ ;
	wire _w1478_ ;
	wire _w1477_ ;
	wire _w1476_ ;
	wire _w1475_ ;
	wire _w1474_ ;
	wire _w1473_ ;
	wire _w1472_ ;
	wire _w1471_ ;
	wire _w1470_ ;
	wire _w1185_ ;
	wire _w1184_ ;
	wire _w1183_ ;
	wire _w1182_ ;
	wire _w1181_ ;
	wire _w1180_ ;
	wire _w1179_ ;
	wire _w1178_ ;
	wire _w1177_ ;
	wire _w1176_ ;
	wire _w1175_ ;
	wire _w1174_ ;
	wire _w1173_ ;
	wire _w1172_ ;
	wire _w1171_ ;
	wire _w1170_ ;
	wire _w1169_ ;
	wire _w1168_ ;
	wire _w1167_ ;
	wire _w1166_ ;
	wire _w1165_ ;
	wire _w1164_ ;
	wire _w1163_ ;
	wire _w1162_ ;
	wire _w1161_ ;
	wire _w1160_ ;
	wire _w1159_ ;
	wire _w1158_ ;
	wire _w1157_ ;
	wire _w1156_ ;
	wire _w1155_ ;
	wire _w1154_ ;
	wire _w1153_ ;
	wire _w1152_ ;
	wire _w1151_ ;
	wire _w1150_ ;
	wire _w1149_ ;
	wire _w1148_ ;
	wire _w1147_ ;
	wire _w1146_ ;
	wire _w1145_ ;
	wire _w1144_ ;
	wire _w1143_ ;
	wire _w1142_ ;
	wire _w1141_ ;
	wire _w1140_ ;
	wire _w1139_ ;
	wire _w1138_ ;
	wire _w1137_ ;
	wire _w1136_ ;
	wire _w1135_ ;
	wire _w1134_ ;
	wire _w1133_ ;
	wire _w1132_ ;
	wire _w1131_ ;
	wire _w1130_ ;
	wire _w1129_ ;
	wire _w1128_ ;
	wire _w1127_ ;
	wire _w1126_ ;
	wire _w1125_ ;
	wire _w1124_ ;
	wire _w1123_ ;
	wire _w1122_ ;
	wire _w1121_ ;
	wire _w1120_ ;
	wire _w1119_ ;
	wire _w1118_ ;
	wire _w1117_ ;
	wire _w1116_ ;
	wire _w1115_ ;
	wire _w1114_ ;
	wire _w1113_ ;
	wire _w1112_ ;
	wire _w1111_ ;
	wire _w1110_ ;
	wire _w1109_ ;
	wire _w1108_ ;
	wire _w1107_ ;
	wire _w1106_ ;
	wire _w1105_ ;
	wire _w1104_ ;
	wire _w1103_ ;
	wire _w1102_ ;
	wire _w1101_ ;
	wire _w1100_ ;
	wire _w1099_ ;
	wire _w1098_ ;
	wire _w1097_ ;
	wire _w1096_ ;
	wire _w1095_ ;
	wire _w1094_ ;
	wire _w1093_ ;
	wire _w1092_ ;
	wire _w1091_ ;
	wire _w1090_ ;
	wire _w1089_ ;
	wire _w1088_ ;
	wire _w1087_ ;
	wire _w1086_ ;
	wire _w1085_ ;
	wire _w1084_ ;
	wire _w1083_ ;
	wire _w1082_ ;
	wire _w1081_ ;
	wire _w1080_ ;
	wire _w1079_ ;
	wire _w1078_ ;
	wire _w1077_ ;
	wire _w1076_ ;
	wire _w1075_ ;
	wire _w1074_ ;
	wire _w1073_ ;
	wire _w1072_ ;
	wire _w1071_ ;
	wire _w1070_ ;
	wire _w1069_ ;
	wire _w1068_ ;
	wire _w1067_ ;
	wire _w1066_ ;
	wire _w1065_ ;
	wire _w1064_ ;
	wire _w1063_ ;
	wire _w1062_ ;
	wire _w1061_ ;
	wire _w1060_ ;
	wire _w1059_ ;
	wire _w1058_ ;
	wire _w1057_ ;
	wire _w1056_ ;
	wire _w987_ ;
	wire _w986_ ;
	wire _w985_ ;
	wire _w984_ ;
	wire _w983_ ;
	wire _w982_ ;
	wire _w981_ ;
	wire _w980_ ;
	wire _w979_ ;
	wire _w978_ ;
	wire _w977_ ;
	wire _w976_ ;
	wire _w975_ ;
	wire _w974_ ;
	wire _w973_ ;
	wire _w972_ ;
	wire _w971_ ;
	wire _w970_ ;
	wire _w969_ ;
	wire _w968_ ;
	wire _w967_ ;
	wire _w966_ ;
	wire _w965_ ;
	wire _w964_ ;
	wire _w963_ ;
	wire _w962_ ;
	wire _w961_ ;
	wire _w960_ ;
	wire _w959_ ;
	wire _w958_ ;
	wire _w941_ ;
	wire _w940_ ;
	wire _w939_ ;
	wire _w938_ ;
	wire _w937_ ;
	wire _w936_ ;
	wire _w935_ ;
	wire _w934_ ;
	wire _w933_ ;
	wire _w932_ ;
	wire _w931_ ;
	wire _w930_ ;
	wire _w929_ ;
	wire _w942_ ;
	wire _w943_ ;
	wire _w944_ ;
	wire _w945_ ;
	wire _w946_ ;
	wire _w947_ ;
	wire _w948_ ;
	wire _w949_ ;
	wire _w950_ ;
	wire _w951_ ;
	wire _w952_ ;
	wire _w953_ ;
	wire _w954_ ;
	wire _w955_ ;
	wire _w956_ ;
	wire _w957_ ;
	wire _w988_ ;
	wire _w989_ ;
	wire _w990_ ;
	wire _w991_ ;
	wire _w992_ ;
	wire _w993_ ;
	wire _w994_ ;
	wire _w995_ ;
	wire _w996_ ;
	wire _w997_ ;
	wire _w998_ ;
	wire _w999_ ;
	wire _w1000_ ;
	wire _w1001_ ;
	wire _w1002_ ;
	wire _w1003_ ;
	wire _w1004_ ;
	wire _w1005_ ;
	wire _w1006_ ;
	wire _w1007_ ;
	wire _w1008_ ;
	wire _w1009_ ;
	wire _w1010_ ;
	wire _w1011_ ;
	wire _w1012_ ;
	wire _w1013_ ;
	wire _w1014_ ;
	wire _w1015_ ;
	wire _w1016_ ;
	wire _w1017_ ;
	wire _w1018_ ;
	wire _w1019_ ;
	wire _w1020_ ;
	wire _w1021_ ;
	wire _w1022_ ;
	wire _w1023_ ;
	wire _w1024_ ;
	wire _w1025_ ;
	wire _w1026_ ;
	wire _w1027_ ;
	wire _w1028_ ;
	wire _w1029_ ;
	wire _w1030_ ;
	wire _w1031_ ;
	wire _w1032_ ;
	wire _w1033_ ;
	wire _w1034_ ;
	wire _w1035_ ;
	wire _w1036_ ;
	wire _w1037_ ;
	wire _w1038_ ;
	wire _w1039_ ;
	wire _w1040_ ;
	wire _w1041_ ;
	wire _w1042_ ;
	wire _w1043_ ;
	wire _w1044_ ;
	wire _w1045_ ;
	wire _w1046_ ;
	wire _w1047_ ;
	wire _w1048_ ;
	wire _w1049_ ;
	wire _w1050_ ;
	wire _w1051_ ;
	wire _w1052_ ;
	wire _w1053_ ;
	wire _w1054_ ;
	wire _w1055_ ;
	wire _w1186_ ;
	wire _w1187_ ;
	wire _w1188_ ;
	wire _w1189_ ;
	wire _w1190_ ;
	wire _w1191_ ;
	wire _w1192_ ;
	wire _w1193_ ;
	wire _w1194_ ;
	wire _w1195_ ;
	wire _w1196_ ;
	wire _w1197_ ;
	wire _w1198_ ;
	wire _w1199_ ;
	wire _w1200_ ;
	wire _w1201_ ;
	wire _w1202_ ;
	wire _w1203_ ;
	wire _w1204_ ;
	wire _w1205_ ;
	wire _w1206_ ;
	wire _w1207_ ;
	wire _w1208_ ;
	wire _w1209_ ;
	wire _w1210_ ;
	wire _w1211_ ;
	wire _w1212_ ;
	wire _w1213_ ;
	wire _w1214_ ;
	wire _w1215_ ;
	wire _w1216_ ;
	wire _w1217_ ;
	wire _w1218_ ;
	wire _w1219_ ;
	wire _w1220_ ;
	wire _w1221_ ;
	wire _w1222_ ;
	wire _w1223_ ;
	wire _w1224_ ;
	wire _w1225_ ;
	wire _w1226_ ;
	wire _w1227_ ;
	wire _w1228_ ;
	wire _w1229_ ;
	wire _w1230_ ;
	wire _w1231_ ;
	wire _w1232_ ;
	wire _w1233_ ;
	wire _w1234_ ;
	wire _w1235_ ;
	wire _w1236_ ;
	wire _w1237_ ;
	wire _w1238_ ;
	wire _w1239_ ;
	wire _w1240_ ;
	wire _w1241_ ;
	wire _w1242_ ;
	wire _w1243_ ;
	wire _w1244_ ;
	wire _w1245_ ;
	wire _w1246_ ;
	wire _w1247_ ;
	wire _w1248_ ;
	wire _w1249_ ;
	wire _w1250_ ;
	wire _w1251_ ;
	wire _w1252_ ;
	wire _w1253_ ;
	wire _w1254_ ;
	wire _w1255_ ;
	wire _w1256_ ;
	wire _w1257_ ;
	wire _w1258_ ;
	wire _w1259_ ;
	wire _w1260_ ;
	wire _w1261_ ;
	wire _w1262_ ;
	wire _w1263_ ;
	wire _w1264_ ;
	wire _w1265_ ;
	wire _w1266_ ;
	wire _w1267_ ;
	wire _w1268_ ;
	wire _w1269_ ;
	wire _w1270_ ;
	wire _w1271_ ;
	wire _w1272_ ;
	wire _w1273_ ;
	wire _w1274_ ;
	wire _w1275_ ;
	wire _w1276_ ;
	wire _w1277_ ;
	wire _w1278_ ;
	wire _w1279_ ;
	wire _w1280_ ;
	wire _w1281_ ;
	wire _w1282_ ;
	wire _w1283_ ;
	wire _w1284_ ;
	wire _w1285_ ;
	wire _w1286_ ;
	wire _w1287_ ;
	wire _w1288_ ;
	wire _w1289_ ;
	wire _w1290_ ;
	wire _w1291_ ;
	wire _w1292_ ;
	wire _w1293_ ;
	wire _w1294_ ;
	wire _w1295_ ;
	wire _w1296_ ;
	wire _w1297_ ;
	wire _w1298_ ;
	wire _w1299_ ;
	wire _w1300_ ;
	wire _w1301_ ;
	wire _w1302_ ;
	wire _w1303_ ;
	wire _w1304_ ;
	wire _w1305_ ;
	wire _w1306_ ;
	wire _w1307_ ;
	wire _w1308_ ;
	wire _w1309_ ;
	wire _w1310_ ;
	wire _w1311_ ;
	wire _w1312_ ;
	wire _w1313_ ;
	wire _w1314_ ;
	wire _w1315_ ;
	wire _w1316_ ;
	wire _w1317_ ;
	wire _w1318_ ;
	wire _w1319_ ;
	wire _w1320_ ;
	wire _w1321_ ;
	wire _w1322_ ;
	wire _w1323_ ;
	wire _w1324_ ;
	wire _w1325_ ;
	wire _w1326_ ;
	wire _w1327_ ;
	wire _w1328_ ;
	wire _w1329_ ;
	wire _w1330_ ;
	wire _w1331_ ;
	wire _w1332_ ;
	wire _w1333_ ;
	wire _w1334_ ;
	wire _w1335_ ;
	wire _w1336_ ;
	wire _w1337_ ;
	wire _w1338_ ;
	wire _w1339_ ;
	wire _w1340_ ;
	wire _w1341_ ;
	wire _w1342_ ;
	wire _w1343_ ;
	wire _w1344_ ;
	wire _w1345_ ;
	wire _w1346_ ;
	wire _w1347_ ;
	wire _w1348_ ;
	wire _w1349_ ;
	wire _w1350_ ;
	wire _w1351_ ;
	wire _w1352_ ;
	wire _w1353_ ;
	wire _w1354_ ;
	wire _w1355_ ;
	wire _w1356_ ;
	wire _w1357_ ;
	wire _w1358_ ;
	wire _w1359_ ;
	wire _w1360_ ;
	wire _w1361_ ;
	wire _w1362_ ;
	wire _w1363_ ;
	wire _w1364_ ;
	wire _w1365_ ;
	wire _w1366_ ;
	wire _w1367_ ;
	wire _w1368_ ;
	wire _w1369_ ;
	wire _w1370_ ;
	wire _w1371_ ;
	wire _w1372_ ;
	wire _w1373_ ;
	wire _w1374_ ;
	wire _w1375_ ;
	wire _w1376_ ;
	wire _w1377_ ;
	wire _w1378_ ;
	wire _w1379_ ;
	wire _w1380_ ;
	wire _w1381_ ;
	wire _w1382_ ;
	wire _w1383_ ;
	wire _w1384_ ;
	wire _w1385_ ;
	wire _w1386_ ;
	wire _w1387_ ;
	wire _w1388_ ;
	wire _w1389_ ;
	wire _w1390_ ;
	wire _w1391_ ;
	wire _w1392_ ;
	wire _w1393_ ;
	wire _w1394_ ;
	wire _w1395_ ;
	wire _w1396_ ;
	wire _w1397_ ;
	wire _w1398_ ;
	wire _w1399_ ;
	wire _w1400_ ;
	wire _w1401_ ;
	wire _w1402_ ;
	wire _w1403_ ;
	wire _w1404_ ;
	wire _w1405_ ;
	wire _w1406_ ;
	wire _w1407_ ;
	wire _w1408_ ;
	wire _w1409_ ;
	wire _w1410_ ;
	wire _w1411_ ;
	wire _w1412_ ;
	wire _w1413_ ;
	wire _w1414_ ;
	wire _w1415_ ;
	wire _w1416_ ;
	wire _w1417_ ;
	wire _w1418_ ;
	wire _w1419_ ;
	wire _w1420_ ;
	wire _w1421_ ;
	wire _w1422_ ;
	wire _w1423_ ;
	wire _w1424_ ;
	wire _w1425_ ;
	wire _w1426_ ;
	wire _w1427_ ;
	wire _w1428_ ;
	wire _w1429_ ;
	wire _w1430_ ;
	wire _w1431_ ;
	wire _w1432_ ;
	wire _w1433_ ;
	wire _w1434_ ;
	wire _w1435_ ;
	wire _w1436_ ;
	wire _w1437_ ;
	wire _w1438_ ;
	wire _w1439_ ;
	wire _w1440_ ;
	wire _w1441_ ;
	wire _w1442_ ;
	wire _w1443_ ;
	wire _w1444_ ;
	wire _w1445_ ;
	wire _w1446_ ;
	wire _w1447_ ;
	wire _w1448_ ;
	wire _w1449_ ;
	wire _w1450_ ;
	wire _w1451_ ;
	wire _w1452_ ;
	wire _w1453_ ;
	wire _w1454_ ;
	wire _w1455_ ;
	wire _w1456_ ;
	wire _w1457_ ;
	wire _w1458_ ;
	wire _w1459_ ;
	wire _w1460_ ;
	wire _w1461_ ;
	wire _w1462_ ;
	wire _w1463_ ;
	wire _w1464_ ;
	wire _w1465_ ;
	wire _w1466_ ;
	wire _w1467_ ;
	wire _w1468_ ;
	wire _w1469_ ;
	wire _w2038_ ;
	wire _w2039_ ;
	wire _w2040_ ;
	wire _w2041_ ;
	wire _w2042_ ;
	wire _w2043_ ;
	wire _w2044_ ;
	wire _w2045_ ;
	wire _w2046_ ;
	wire _w2047_ ;
	wire _w2048_ ;
	wire _w2049_ ;
	wire _w2050_ ;
	wire _w2051_ ;
	wire _w2052_ ;
	wire _w2053_ ;
	wire _w2054_ ;
	wire _w2055_ ;
	wire _w2056_ ;
	wire _w2057_ ;
	wire _w2058_ ;
	wire _w2059_ ;
	wire _w2060_ ;
	wire _w2061_ ;
	wire _w2062_ ;
	wire _w2063_ ;
	wire _w2064_ ;
	wire _w2065_ ;
	wire _w2066_ ;
	wire _w2067_ ;
	wire _w2068_ ;
	wire _w2069_ ;
	wire _w2070_ ;
	wire _w2071_ ;
	wire _w2072_ ;
	wire _w2073_ ;
	wire _w2074_ ;
	wire _w2075_ ;
	wire _w2076_ ;
	wire _w2077_ ;
	wire _w2078_ ;
	wire _w2079_ ;
	wire _w2080_ ;
	wire _w2081_ ;
	wire _w2082_ ;
	wire _w2083_ ;
	wire _w2084_ ;
	wire _w2085_ ;
	wire _w2086_ ;
	wire _w2087_ ;
	wire _w2088_ ;
	wire _w2089_ ;
	wire _w2090_ ;
	wire _w2091_ ;
	wire _w2092_ ;
	wire _w2093_ ;
	wire _w2094_ ;
	wire _w2095_ ;
	wire _w2096_ ;
	wire _w2097_ ;
	wire _w2098_ ;
	wire _w2099_ ;
	wire _w2100_ ;
	wire _w2101_ ;
	wire _w2102_ ;
	wire _w2103_ ;
	wire _w2104_ ;
	wire _w2105_ ;
	wire _w2106_ ;
	wire _w2107_ ;
	wire _w2108_ ;
	wire _w2109_ ;
	wire _w2110_ ;
	wire _w2111_ ;
	wire _w2112_ ;
	wire _w2113_ ;
	wire _w2114_ ;
	wire _w2115_ ;
	wire _w2116_ ;
	wire _w2117_ ;
	wire _w2118_ ;
	wire _w2119_ ;
	wire _w2120_ ;
	wire _w2121_ ;
	wire _w2122_ ;
	wire _w2123_ ;
	wire _w2124_ ;
	wire _w2125_ ;
	wire _w2126_ ;
	wire _w2127_ ;
	wire _w2128_ ;
	wire _w2129_ ;
	wire _w2130_ ;
	wire _w2131_ ;
	wire _w2132_ ;
	wire _w2133_ ;
	wire _w2134_ ;
	wire _w2135_ ;
	wire _w2136_ ;
	wire _w2137_ ;
	wire _w2138_ ;
	wire _w2139_ ;
	wire _w2140_ ;
	wire _w2141_ ;
	wire _w2142_ ;
	wire _w2143_ ;
	wire _w2144_ ;
	wire _w2145_ ;
	wire _w2146_ ;
	wire _w2147_ ;
	wire _w2148_ ;
	wire _w2149_ ;
	wire _w2150_ ;
	wire _w2151_ ;
	wire _w2152_ ;
	wire _w2153_ ;
	wire _w2154_ ;
	wire _w2155_ ;
	wire _w2156_ ;
	wire _w2157_ ;
	wire _w2158_ ;
	wire _w2159_ ;
	wire _w2160_ ;
	wire _w2161_ ;
	wire _w2162_ ;
	wire _w2163_ ;
	wire _w2164_ ;
	wire _w2165_ ;
	wire _w2166_ ;
	wire _w2167_ ;
	wire _w2168_ ;
	wire _w2169_ ;
	wire _w2170_ ;
	wire _w2171_ ;
	wire _w2172_ ;
	wire _w2173_ ;
	wire _w2174_ ;
	wire _w2175_ ;
	wire _w2176_ ;
	wire _w2177_ ;
	wire _w2178_ ;
	wire _w2179_ ;
	wire _w2180_ ;
	wire _w2181_ ;
	wire _w2182_ ;
	wire _w2183_ ;
	wire _w2184_ ;
	wire _w2185_ ;
	wire _w2186_ ;
	wire _w2187_ ;
	wire _w2188_ ;
	wire _w2189_ ;
	wire _w2190_ ;
	wire _w2191_ ;
	wire _w2192_ ;
	wire _w2193_ ;
	wire _w2194_ ;
	wire _w2195_ ;
	wire _w2196_ ;
	wire _w2197_ ;
	wire _w2198_ ;
	wire _w2199_ ;
	wire _w2200_ ;
	wire _w2201_ ;
	wire _w2202_ ;
	wire _w2203_ ;
	wire _w2204_ ;
	wire _w2205_ ;
	wire _w2206_ ;
	wire _w2207_ ;
	wire _w2208_ ;
	wire _w2209_ ;
	wire _w2210_ ;
	wire _w2211_ ;
	wire _w2212_ ;
	wire _w2213_ ;
	wire _w2214_ ;
	wire _w2215_ ;
	wire _w2216_ ;
	wire _w2217_ ;
	wire _w2218_ ;
	wire _w2219_ ;
	wire _w2220_ ;
	wire _w2221_ ;
	wire _w2222_ ;
	wire _w2223_ ;
	wire _w2224_ ;
	wire _w2225_ ;
	wire _w2226_ ;
	wire _w2227_ ;
	wire _w2228_ ;
	wire _w2229_ ;
	wire _w2230_ ;
	wire _w2231_ ;
	wire _w2232_ ;
	wire _w2233_ ;
	wire _w2234_ ;
	wire _w2235_ ;
	wire _w2236_ ;
	wire _w2237_ ;
	wire _w2238_ ;
	wire _w2239_ ;
	wire _w2240_ ;
	wire _w2241_ ;
	wire _w2242_ ;
	wire _w2243_ ;
	wire _w2244_ ;
	wire _w2245_ ;
	wire _w2246_ ;
	wire _w2247_ ;
	wire _w2248_ ;
	wire _w2249_ ;
	wire _w2250_ ;
	wire _w2251_ ;
	wire _w2252_ ;
	wire _w2253_ ;
	wire _w2254_ ;
	wire _w2255_ ;
	wire _w2256_ ;
	wire _w2257_ ;
	wire _w2258_ ;
	wire _w2259_ ;
	wire _w2260_ ;
	wire _w2261_ ;
	wire _w2262_ ;
	wire _w2263_ ;
	wire _w2264_ ;
	wire _w2265_ ;
	wire _w2266_ ;
	wire _w2267_ ;
	wire _w2268_ ;
	wire _w2269_ ;
	wire _w2270_ ;
	wire _w2271_ ;
	wire _w2272_ ;
	wire _w2273_ ;
	wire _w2274_ ;
	wire _w2275_ ;
	wire _w2276_ ;
	wire _w2277_ ;
	wire _w2278_ ;
	wire _w2279_ ;
	wire _w2280_ ;
	wire _w2281_ ;
	wire _w2282_ ;
	wire _w2283_ ;
	wire _w2284_ ;
	wire _w2285_ ;
	wire _w2286_ ;
	wire _w2287_ ;
	wire _w2288_ ;
	wire _w2289_ ;
	wire _w2290_ ;
	wire _w2291_ ;
	wire _w2292_ ;
	wire _w2293_ ;
	wire _w2294_ ;
	wire _w2295_ ;
	wire _w2296_ ;
	wire _w2297_ ;
	wire _w2298_ ;
	wire _w2299_ ;
	wire _w2300_ ;
	wire _w2301_ ;
	wire _w2302_ ;
	wire _w2303_ ;
	wire _w2304_ ;
	wire _w2305_ ;
	wire _w2306_ ;
	wire _w2307_ ;
	wire _w2308_ ;
	wire _w2309_ ;
	wire _w2310_ ;
	wire _w2311_ ;
	wire _w2312_ ;
	wire _w2313_ ;
	wire _w2314_ ;
	wire _w2315_ ;
	wire _w2316_ ;
	wire _w2317_ ;
	wire _w2318_ ;
	wire _w2319_ ;
	wire _w2320_ ;
	wire _w2321_ ;
	wire _w2322_ ;
	wire _w2323_ ;
	wire _w2324_ ;
	wire _w2325_ ;
	wire _w2326_ ;
	wire _w2327_ ;
	wire _w2328_ ;
	wire _w2329_ ;
	wire _w2330_ ;
	wire _w2331_ ;
	wire _w2332_ ;
	wire _w2333_ ;
	wire _w2334_ ;
	wire _w2335_ ;
	wire _w2336_ ;
	wire _w2337_ ;
	wire _w2338_ ;
	wire _w2339_ ;
	wire _w2340_ ;
	wire _w2341_ ;
	wire _w2342_ ;
	wire _w2343_ ;
	wire _w2344_ ;
	wire _w2345_ ;
	wire _w2346_ ;
	wire _w2347_ ;
	wire _w2348_ ;
	wire _w2349_ ;
	wire _w2350_ ;
	wire _w2351_ ;
	wire _w2352_ ;
	wire _w2353_ ;
	wire _w2354_ ;
	wire _w2355_ ;
	wire _w2356_ ;
	wire _w2357_ ;
	wire _w2358_ ;
	wire _w2359_ ;
	wire _w2360_ ;
	wire _w2361_ ;
	wire _w2362_ ;
	wire _w2363_ ;
	wire _w2364_ ;
	wire _w2365_ ;
	wire _w2366_ ;
	wire _w2367_ ;
	wire _w2368_ ;
	wire _w2369_ ;
	wire _w2370_ ;
	wire _w2371_ ;
	wire _w2372_ ;
	wire _w2373_ ;
	wire _w2374_ ;
	wire _w2375_ ;
	wire _w2376_ ;
	wire _w2377_ ;
	wire _w2378_ ;
	wire _w2379_ ;
	wire _w2380_ ;
	wire _w2381_ ;
	wire _w2382_ ;
	wire _w2383_ ;
	wire _w2384_ ;
	wire _w2385_ ;
	wire _w2386_ ;
	wire _w2387_ ;
	wire _w2388_ ;
	wire _w2389_ ;
	wire _w2390_ ;
	wire _w2391_ ;
	wire _w2392_ ;
	wire _w2393_ ;
	wire _w2394_ ;
	wire _w2395_ ;
	wire _w2396_ ;
	wire _w2397_ ;
	wire _w2398_ ;
	wire _w2399_ ;
	wire _w2400_ ;
	wire _w2401_ ;
	wire _w2402_ ;
	wire _w2403_ ;
	wire _w2404_ ;
	wire _w2405_ ;
	wire _w2406_ ;
	wire _w2407_ ;
	wire _w2408_ ;
	wire _w2409_ ;
	wire _w2410_ ;
	wire _w2411_ ;
	wire _w2412_ ;
	wire _w2413_ ;
	wire _w2414_ ;
	wire _w2415_ ;
	wire _w2416_ ;
	wire _w2417_ ;
	wire _w2418_ ;
	wire _w2419_ ;
	wire _w2420_ ;
	wire _w2421_ ;
	wire _w2422_ ;
	wire _w2423_ ;
	wire _w2424_ ;
	wire _w2425_ ;
	wire _w2426_ ;
	wire _w2427_ ;
	wire _w2428_ ;
	wire _w2429_ ;
	wire _w2430_ ;
	wire _w2431_ ;
	wire _w2432_ ;
	wire _w2433_ ;
	wire _w2434_ ;
	wire _w2435_ ;
	wire _w2436_ ;
	wire _w2437_ ;
	wire _w2438_ ;
	wire _w2439_ ;
	wire _w2440_ ;
	wire _w2441_ ;
	wire _w2442_ ;
	wire _w2443_ ;
	wire _w2444_ ;
	wire _w2445_ ;
	wire _w2446_ ;
	wire _w2447_ ;
	wire _w2448_ ;
	wire _w2449_ ;
	wire _w2450_ ;
	wire _w2451_ ;
	wire _w2452_ ;
	wire _w2453_ ;
	wire _w2454_ ;
	wire _w2455_ ;
	wire _w2456_ ;
	wire _w2457_ ;
	wire _w2458_ ;
	wire _w2459_ ;
	wire _w2460_ ;
	wire _w2461_ ;
	wire _w2462_ ;
	wire _w2463_ ;
	wire _w2464_ ;
	wire _w2465_ ;
	wire _w2466_ ;
	wire _w2467_ ;
	wire _w2468_ ;
	wire _w2469_ ;
	wire _w2470_ ;
	wire _w2471_ ;
	wire _w2472_ ;
	wire _w2473_ ;
	wire _w2474_ ;
	wire _w2475_ ;
	wire _w2476_ ;
	wire _w2477_ ;
	wire _w2478_ ;
	wire _w2479_ ;
	wire _w2480_ ;
	wire _w2481_ ;
	wire _w2482_ ;
	wire _w2483_ ;
	wire _w2484_ ;
	wire _w2485_ ;
	wire _w2486_ ;
	wire _w2487_ ;
	wire _w2488_ ;
	wire _w2489_ ;
	wire _w2490_ ;
	wire _w2491_ ;
	wire _w2492_ ;
	wire _w2493_ ;
	wire _w2494_ ;
	wire _w2495_ ;
	wire _w2496_ ;
	wire _w2497_ ;
	wire _w2498_ ;
	wire _w2499_ ;
	wire _w2500_ ;
	wire _w2501_ ;
	wire _w2502_ ;
	wire _w2503_ ;
	wire _w2504_ ;
	wire _w2505_ ;
	wire _w2506_ ;
	wire _w2507_ ;
	wire _w2508_ ;
	wire _w2509_ ;
	wire _w2510_ ;
	wire _w2511_ ;
	wire _w2512_ ;
	wire _w2513_ ;
	wire _w2514_ ;
	wire _w2515_ ;
	wire _w2516_ ;
	wire _w2517_ ;
	wire _w2518_ ;
	wire _w2519_ ;
	wire _w2520_ ;
	wire _w2521_ ;
	wire _w2522_ ;
	wire _w2523_ ;
	wire _w2524_ ;
	wire _w2525_ ;
	wire _w2526_ ;
	wire _w2527_ ;
	wire _w2528_ ;
	wire _w2529_ ;
	wire _w2530_ ;
	wire _w2531_ ;
	wire _w2532_ ;
	wire _w2533_ ;
	wire _w2534_ ;
	wire _w2535_ ;
	wire _w2536_ ;
	wire _w2537_ ;
	wire _w2538_ ;
	wire _w2539_ ;
	wire _w2540_ ;
	wire _w2541_ ;
	wire _w2542_ ;
	wire _w2543_ ;
	wire _w2544_ ;
	wire _w2545_ ;
	wire _w2546_ ;
	wire _w2547_ ;
	wire _w2548_ ;
	wire _w2549_ ;
	wire _w2550_ ;
	wire _w2551_ ;
	wire _w2552_ ;
	wire _w2553_ ;
	wire _w2554_ ;
	wire _w2555_ ;
	wire _w2556_ ;
	wire _w2557_ ;
	wire _w2558_ ;
	wire _w2559_ ;
	wire _w2560_ ;
	wire _w2561_ ;
	wire _w2562_ ;
	wire _w2563_ ;
	wire _w2564_ ;
	wire _w2565_ ;
	wire _w2566_ ;
	wire _w2567_ ;
	wire _w2568_ ;
	wire _w2569_ ;
	wire _w2570_ ;
	wire _w2571_ ;
	wire _w2572_ ;
	wire _w2573_ ;
	wire _w2574_ ;
	wire _w2575_ ;
	wire _w2576_ ;
	wire _w2577_ ;
	wire _w2578_ ;
	wire _w2579_ ;
	wire _w2580_ ;
	wire _w2581_ ;
	wire _w2582_ ;
	wire _w2583_ ;
	wire _w2584_ ;
	wire _w2585_ ;
	wire _w2586_ ;
	wire _w2587_ ;
	wire _w2588_ ;
	wire _w2589_ ;
	wire _w2590_ ;
	wire _w2591_ ;
	wire _w2592_ ;
	wire _w2593_ ;
	wire _w2594_ ;
	wire _w2595_ ;
	wire _w2596_ ;
	wire _w2597_ ;
	wire _w2598_ ;
	wire _w2599_ ;
	wire _w2600_ ;
	wire _w2601_ ;
	wire _w2602_ ;
	wire _w2603_ ;
	wire _w2604_ ;
	wire _w2605_ ;
	wire _w2606_ ;
	wire _w2607_ ;
	wire _w2608_ ;
	wire _w2609_ ;
	wire _w2610_ ;
	wire _w2611_ ;
	wire _w2612_ ;
	wire _w2613_ ;
	wire _w2614_ ;
	wire _w2615_ ;
	wire _w2616_ ;
	wire _w2617_ ;
	wire _w2618_ ;
	wire _w2619_ ;
	wire _w2620_ ;
	wire _w2621_ ;
	wire _w2622_ ;
	wire _w2623_ ;
	wire _w2624_ ;
	wire _w2625_ ;
	wire _w2626_ ;
	wire _w2627_ ;
	wire _w2628_ ;
	wire _w2629_ ;
	wire _w2630_ ;
	wire _w2631_ ;
	wire _w2632_ ;
	wire _w2633_ ;
	wire _w2634_ ;
	wire _w2635_ ;
	wire _w2636_ ;
	wire _w2637_ ;
	wire _w2638_ ;
	wire _w2639_ ;
	wire _w2640_ ;
	wire _w2641_ ;
	wire _w2642_ ;
	wire _w2643_ ;
	wire _w2644_ ;
	wire _w2645_ ;
	wire _w2646_ ;
	wire _w2647_ ;
	wire _w2648_ ;
	wire _w2649_ ;
	wire _w2650_ ;
	wire _w2651_ ;
	wire _w2652_ ;
	wire _w2653_ ;
	wire _w2654_ ;
	wire _w2655_ ;
	wire _w2656_ ;
	wire _w2657_ ;
	wire _w2658_ ;
	wire _w2659_ ;
	wire _w2660_ ;
	wire _w2661_ ;
	wire _w2662_ ;
	wire _w2663_ ;
	wire _w2664_ ;
	wire _w2665_ ;
	wire _w2666_ ;
	wire _w2667_ ;
	wire _w2668_ ;
	wire _w2669_ ;
	wire _w2670_ ;
	wire _w2671_ ;
	wire _w2672_ ;
	wire _w2673_ ;
	wire _w2674_ ;
	wire _w2675_ ;
	wire _w2676_ ;
	wire _w2677_ ;
	wire _w2678_ ;
	wire _w2679_ ;
	wire _w2680_ ;
	wire _w2681_ ;
	wire _w2682_ ;
	wire _w2683_ ;
	wire _w2684_ ;
	wire _w2685_ ;
	wire _w2686_ ;
	wire _w2687_ ;
	wire _w2688_ ;
	wire _w2689_ ;
	wire _w2690_ ;
	wire _w2691_ ;
	wire _w2692_ ;
	wire _w2693_ ;
	wire _w2694_ ;
	wire _w2695_ ;
	wire _w2696_ ;
	wire _w2697_ ;
	wire _w2698_ ;
	wire _w2699_ ;
	wire _w2700_ ;
	wire _w2701_ ;
	wire _w2702_ ;
	wire _w2703_ ;
	wire _w2704_ ;
	wire _w2705_ ;
	wire _w2706_ ;
	wire _w2707_ ;
	wire _w2708_ ;
	wire _w2709_ ;
	wire _w2710_ ;
	wire _w2711_ ;
	wire _w2712_ ;
	wire _w2713_ ;
	wire _w2714_ ;
	wire _w2715_ ;
	wire _w2716_ ;
	wire _w2717_ ;
	wire _w2718_ ;
	wire _w2719_ ;
	wire _w2720_ ;
	wire _w2721_ ;
	wire _w2722_ ;
	wire _w2723_ ;
	wire _w2724_ ;
	wire _w2725_ ;
	wire _w2726_ ;
	wire _w2727_ ;
	wire _w2728_ ;
	wire _w2729_ ;
	wire _w2730_ ;
	wire _w2731_ ;
	wire _w2732_ ;
	wire _w2733_ ;
	wire _w2734_ ;
	wire _w2735_ ;
	wire _w2736_ ;
	wire _w2737_ ;
	wire _w2738_ ;
	wire _w2739_ ;
	wire _w2740_ ;
	wire _w2741_ ;
	wire _w2742_ ;
	wire _w2743_ ;
	wire _w2744_ ;
	wire _w2745_ ;
	wire _w2746_ ;
	wire _w2747_ ;
	wire _w2748_ ;
	wire _w2749_ ;
	wire _w2750_ ;
	wire _w2751_ ;
	wire _w2752_ ;
	wire _w2753_ ;
	wire _w2754_ ;
	wire _w2755_ ;
	wire _w2756_ ;
	wire _w2757_ ;
	wire _w2758_ ;
	wire _w2759_ ;
	wire _w2760_ ;
	wire _w2761_ ;
	wire _w2762_ ;
	wire _w2763_ ;
	wire _w2764_ ;
	wire _w2765_ ;
	wire _w2766_ ;
	wire _w2767_ ;
	wire _w2768_ ;
	wire _w2769_ ;
	wire _w2770_ ;
	wire _w2771_ ;
	wire _w2772_ ;
	wire _w2773_ ;
	wire _w2774_ ;
	wire _w2775_ ;
	wire _w2776_ ;
	wire _w2777_ ;
	wire _w2778_ ;
	wire _w2779_ ;
	wire _w2780_ ;
	wire _w2781_ ;
	wire _w2782_ ;
	wire _w2783_ ;
	wire _w2784_ ;
	wire _w2785_ ;
	wire _w2786_ ;
	wire _w2787_ ;
	wire _w2788_ ;
	wire _w2789_ ;
	wire _w2790_ ;
	wire _w2791_ ;
	wire _w2792_ ;
	wire _w2793_ ;
	wire _w2794_ ;
	wire _w2795_ ;
	wire _w2796_ ;
	wire _w2797_ ;
	wire _w2798_ ;
	wire _w2799_ ;
	wire _w2800_ ;
	wire _w2801_ ;
	wire _w2802_ ;
	wire _w2803_ ;
	wire _w2804_ ;
	wire _w2805_ ;
	wire _w2806_ ;
	wire _w2807_ ;
	wire _w2808_ ;
	wire _w2809_ ;
	wire _w2810_ ;
	wire _w2811_ ;
	wire _w2812_ ;
	wire _w2813_ ;
	wire _w2814_ ;
	wire _w2815_ ;
	wire _w2816_ ;
	wire _w2817_ ;
	wire _w2818_ ;
	wire _w2819_ ;
	wire _w2820_ ;
	wire _w2821_ ;
	wire _w2822_ ;
	wire _w2823_ ;
	wire _w2824_ ;
	wire _w2825_ ;
	wire _w2826_ ;
	wire _w2827_ ;
	wire _w2828_ ;
	wire _w2829_ ;
	wire _w2830_ ;
	wire _w2831_ ;
	wire _w2832_ ;
	wire _w2833_ ;
	wire _w2834_ ;
	wire _w2835_ ;
	wire _w2836_ ;
	wire _w2837_ ;
	wire _w2838_ ;
	wire _w2839_ ;
	wire _w2840_ ;
	wire _w2841_ ;
	wire _w2842_ ;
	wire _w2843_ ;
	wire _w2844_ ;
	wire _w2845_ ;
	wire _w2846_ ;
	wire _w2847_ ;
	wire _w2848_ ;
	wire _w2849_ ;
	wire _w2850_ ;
	wire _w2851_ ;
	wire _w2852_ ;
	wire _w2853_ ;
	wire _w2854_ ;
	wire _w2855_ ;
	wire _w2856_ ;
	wire _w2857_ ;
	wire _w2858_ ;
	wire _w2859_ ;
	wire _w2860_ ;
	wire _w2861_ ;
	wire _w2862_ ;
	wire _w2863_ ;
	wire _w2864_ ;
	wire _w2865_ ;
	wire _w2866_ ;
	wire _w2867_ ;
	wire _w2868_ ;
	wire _w2869_ ;
	wire _w2870_ ;
	wire _w2871_ ;
	wire _w2872_ ;
	wire _w2873_ ;
	wire _w2874_ ;
	wire _w2875_ ;
	wire _w2876_ ;
	wire _w2877_ ;
	wire _w2878_ ;
	wire _w2879_ ;
	wire _w2880_ ;
	wire _w2881_ ;
	wire _w2882_ ;
	wire _w2883_ ;
	wire _w2884_ ;
	wire _w2885_ ;
	wire _w2886_ ;
	wire _w2887_ ;
	wire _w2888_ ;
	wire _w2889_ ;
	wire _w2890_ ;
	wire _w2891_ ;
	wire _w2892_ ;
	wire _w2893_ ;
	wire _w2894_ ;
	wire _w2895_ ;
	wire _w2896_ ;
	wire _w2897_ ;
	wire _w2898_ ;
	wire _w2899_ ;
	wire _w2900_ ;
	wire _w2901_ ;
	wire _w2902_ ;
	wire _w2903_ ;
	wire _w2904_ ;
	wire _w2905_ ;
	wire _w2906_ ;
	wire _w2907_ ;
	wire _w2908_ ;
	wire _w2909_ ;
	wire _w2910_ ;
	wire _w2911_ ;
	wire _w2912_ ;
	wire _w2913_ ;
	wire _w2914_ ;
	wire _w2915_ ;
	wire _w2916_ ;
	wire _w2917_ ;
	wire _w2918_ ;
	wire _w2919_ ;
	wire _w2920_ ;
	wire _w2921_ ;
	wire _w2922_ ;
	wire _w2923_ ;
	wire _w2924_ ;
	wire _w2925_ ;
	wire _w2926_ ;
	wire _w2927_ ;
	wire _w2928_ ;
	wire _w2929_ ;
	wire _w2930_ ;
	wire _w2931_ ;
	wire _w2932_ ;
	wire _w2933_ ;
	wire _w2934_ ;
	wire _w2935_ ;
	wire _w2936_ ;
	wire _w2937_ ;
	wire _w2938_ ;
	wire _w2939_ ;
	wire _w2940_ ;
	wire _w2941_ ;
	wire _w2942_ ;
	wire _w2943_ ;
	wire _w2944_ ;
	wire _w2945_ ;
	wire _w2946_ ;
	wire _w2947_ ;
	wire _w2948_ ;
	wire _w2949_ ;
	wire _w2950_ ;
	wire _w2951_ ;
	wire _w2952_ ;
	wire _w2953_ ;
	wire _w2954_ ;
	wire _w2955_ ;
	wire _w2956_ ;
	wire _w2957_ ;
	wire _w2958_ ;
	wire _w2959_ ;
	wire _w2960_ ;
	wire _w2961_ ;
	wire _w2962_ ;
	wire _w2963_ ;
	wire _w2964_ ;
	wire _w2965_ ;
	wire _w2966_ ;
	wire _w2967_ ;
	wire _w2968_ ;
	wire _w2969_ ;
	wire _w2970_ ;
	wire _w2971_ ;
	wire _w2972_ ;
	wire _w2973_ ;
	wire _w2974_ ;
	wire _w2975_ ;
	wire _w2976_ ;
	wire _w2977_ ;
	wire _w2978_ ;
	wire _w2979_ ;
	wire _w2980_ ;
	wire _w2981_ ;
	wire _w2982_ ;
	wire _w2983_ ;
	wire _w2984_ ;
	wire _w2985_ ;
	wire _w2986_ ;
	wire _w2987_ ;
	wire _w2988_ ;
	wire _w2989_ ;
	wire _w2990_ ;
	wire _w2991_ ;
	wire _w2992_ ;
	wire _w2993_ ;
	wire _w2994_ ;
	wire _w2995_ ;
	wire _w2996_ ;
	wire _w2997_ ;
	wire _w2998_ ;
	wire _w2999_ ;
	wire _w3000_ ;
	wire _w3001_ ;
	wire _w3002_ ;
	wire _w3003_ ;
	wire _w3004_ ;
	wire _w3005_ ;
	wire _w3006_ ;
	wire _w3007_ ;
	wire _w3008_ ;
	wire _w3009_ ;
	wire _w3010_ ;
	wire _w3011_ ;
	wire _w3012_ ;
	wire _w3013_ ;
	wire _w3014_ ;
	wire _w3015_ ;
	wire _w3016_ ;
	wire _w3017_ ;
	wire _w3018_ ;
	wire _w3019_ ;
	wire _w3020_ ;
	wire _w3021_ ;
	wire _w3022_ ;
	wire _w3023_ ;
	wire _w3024_ ;
	wire _w3025_ ;
	wire _w3026_ ;
	wire _w3027_ ;
	wire _w3028_ ;
	wire _w3029_ ;
	wire _w3030_ ;
	wire _w3031_ ;
	wire _w3032_ ;
	wire _w3033_ ;
	wire _w3034_ ;
	wire _w3035_ ;
	wire _w3036_ ;
	wire _w3037_ ;
	wire _w3038_ ;
	wire _w3039_ ;
	wire _w3040_ ;
	wire _w3041_ ;
	wire _w3042_ ;
	wire _w3043_ ;
	wire _w3044_ ;
	wire _w3045_ ;
	wire _w3046_ ;
	wire _w3047_ ;
	wire _w3048_ ;
	wire _w3049_ ;
	wire _w3050_ ;
	wire _w3051_ ;
	wire _w3052_ ;
	wire _w3053_ ;
	wire _w3054_ ;
	wire _w3055_ ;
	wire _w3056_ ;
	wire _w3057_ ;
	wire _w3058_ ;
	wire _w3059_ ;
	wire _w3060_ ;
	wire _w3061_ ;
	wire _w3062_ ;
	wire _w3063_ ;
	wire _w3064_ ;
	wire _w3065_ ;
	wire _w3066_ ;
	wire _w3067_ ;
	wire _w3068_ ;
	wire _w3069_ ;
	wire _w3070_ ;
	wire _w3071_ ;
	wire _w3072_ ;
	wire _w3073_ ;
	wire _w3074_ ;
	wire _w3075_ ;
	wire _w3076_ ;
	wire _w3077_ ;
	wire _w3078_ ;
	wire _w3079_ ;
	wire _w3080_ ;
	wire _w3081_ ;
	wire _w3082_ ;
	wire _w3083_ ;
	wire _w3084_ ;
	wire _w3085_ ;
	wire _w3086_ ;
	wire _w3087_ ;
	wire _w3088_ ;
	wire _w3089_ ;
	wire _w3090_ ;
	wire _w3091_ ;
	wire _w3092_ ;
	wire _w3093_ ;
	wire _w3094_ ;
	wire _w3095_ ;
	wire _w3096_ ;
	wire _w3097_ ;
	wire _w3098_ ;
	wire _w3099_ ;
	wire _w3100_ ;
	wire _w3101_ ;
	wire _w3102_ ;
	wire _w3103_ ;
	wire _w3104_ ;
	wire _w3105_ ;
	wire _w3106_ ;
	wire _w3107_ ;
	wire _w3108_ ;
	wire _w3109_ ;
	wire _w3110_ ;
	wire _w3111_ ;
	wire _w3112_ ;
	wire _w3113_ ;
	wire _w3114_ ;
	wire _w3115_ ;
	wire _w3116_ ;
	wire _w3117_ ;
	wire _w3118_ ;
	wire _w3119_ ;
	wire _w3120_ ;
	wire _w3121_ ;
	wire _w3122_ ;
	wire _w3123_ ;
	wire _w3124_ ;
	wire _w3125_ ;
	wire _w3126_ ;
	wire _w3127_ ;
	wire _w3128_ ;
	wire _w3129_ ;
	wire _w3130_ ;
	wire _w3131_ ;
	wire _w3132_ ;
	wire _w3133_ ;
	wire _w3134_ ;
	wire _w3135_ ;
	wire _w3136_ ;
	wire _w3137_ ;
	wire _w3138_ ;
	wire _w3139_ ;
	wire _w3140_ ;
	wire _w3141_ ;
	wire _w3142_ ;
	wire _w3143_ ;
	wire _w3144_ ;
	wire _w3145_ ;
	wire _w3146_ ;
	wire _w3147_ ;
	wire _w3148_ ;
	wire _w3149_ ;
	wire _w3150_ ;
	wire _w3151_ ;
	wire _w3152_ ;
	wire _w3153_ ;
	wire _w3154_ ;
	wire _w3155_ ;
	wire _w3156_ ;
	wire _w3157_ ;
	wire _w3158_ ;
	wire _w3159_ ;
	wire _w3160_ ;
	wire _w3161_ ;
	wire _w3162_ ;
	wire _w3163_ ;
	wire _w3164_ ;
	wire _w3165_ ;
	wire _w3166_ ;
	wire _w3167_ ;
	wire _w3168_ ;
	wire _w3169_ ;
	wire _w3170_ ;
	wire _w3171_ ;
	wire _w3172_ ;
	wire _w3173_ ;
	wire _w3174_ ;
	wire _w3175_ ;
	wire _w3176_ ;
	wire _w3177_ ;
	wire _w3178_ ;
	wire _w3179_ ;
	wire _w3180_ ;
	wire _w3181_ ;
	wire _w3182_ ;
	wire _w3183_ ;
	wire _w3184_ ;
	wire _w3185_ ;
	wire _w3186_ ;
	wire _w3187_ ;
	wire _w3188_ ;
	wire _w3189_ ;
	wire _w3190_ ;
	wire _w3191_ ;
	wire _w3192_ ;
	wire _w3193_ ;
	wire _w3194_ ;
	wire _w3195_ ;
	wire _w3196_ ;
	wire _w3197_ ;
	wire _w3198_ ;
	wire _w3199_ ;
	wire _w3200_ ;
	wire _w3201_ ;
	wire _w3202_ ;
	wire _w3203_ ;
	wire _w3204_ ;
	wire _w3205_ ;
	wire _w3206_ ;
	wire _w3207_ ;
	wire _w3208_ ;
	wire _w3209_ ;
	wire _w3210_ ;
	wire _w3211_ ;
	wire _w3212_ ;
	wire _w3213_ ;
	wire _w3214_ ;
	wire _w3215_ ;
	wire _w3216_ ;
	wire _w3217_ ;
	wire _w3218_ ;
	wire _w3219_ ;
	wire _w3220_ ;
	wire _w3221_ ;
	wire _w3222_ ;
	wire _w3223_ ;
	wire _w3224_ ;
	wire _w3225_ ;
	wire _w3226_ ;
	wire _w3227_ ;
	wire _w3228_ ;
	wire _w3229_ ;
	wire _w3230_ ;
	wire _w3231_ ;
	wire _w3232_ ;
	wire _w3233_ ;
	wire _w3234_ ;
	wire _w3235_ ;
	wire _w3236_ ;
	wire _w3237_ ;
	wire _w3238_ ;
	wire _w3239_ ;
	wire _w3240_ ;
	wire _w3241_ ;
	wire _w3242_ ;
	wire _w3243_ ;
	wire _w3244_ ;
	wire _w3245_ ;
	wire _w3246_ ;
	wire _w3247_ ;
	wire _w3248_ ;
	wire _w3249_ ;
	wire _w3250_ ;
	wire _w3251_ ;
	wire _w3252_ ;
	wire _w3253_ ;
	wire _w3254_ ;
	wire _w3255_ ;
	wire _w3256_ ;
	wire _w3257_ ;
	wire _w3258_ ;
	wire _w3259_ ;
	wire _w3260_ ;
	wire _w3261_ ;
	wire _w3262_ ;
	wire _w3263_ ;
	wire _w3264_ ;
	wire _w3265_ ;
	wire _w3266_ ;
	wire _w3267_ ;
	wire _w3268_ ;
	wire _w3269_ ;
	wire _w3270_ ;
	wire _w3271_ ;
	wire _w3272_ ;
	wire _w3273_ ;
	wire _w3274_ ;
	wire _w3275_ ;
	wire _w3276_ ;
	wire _w3277_ ;
	wire _w3278_ ;
	wire _w3279_ ;
	wire _w3280_ ;
	wire _w3281_ ;
	wire _w3282_ ;
	wire _w3283_ ;
	wire _w3284_ ;
	wire _w3285_ ;
	LUT3 #(
		.INIT('h10)
	) name0 (
		\ks1_state_reg[0]/NET0131 ,
		\ks1_state_reg[1]/NET0131 ,
		\ks1_state_reg[2]/NET0131 ,
		_w929_
	);
	LUT4 #(
		.INIT('h0001)
	) name1 (
		\round_reg[0]/NET0131 ,
		\round_reg[1]/NET0131 ,
		\round_reg[2]/NET0131 ,
		\round_reg[3]/NET0131 ,
		_w930_
	);
	LUT2 #(
		.INIT('h8)
	) name2 (
		\addroundkey_start_i_reg/NET0131 ,
		_w930_,
		_w931_
	);
	LUT4 #(
		.INIT('h8421)
	) name3 (
		\addroundkey_round_reg[0]/NET0131 ,
		\addroundkey_round_reg[2]/NET0131 ,
		\round_reg[0]/NET0131 ,
		\round_reg[2]/NET0131 ,
		_w932_
	);
	LUT4 #(
		.INIT('h8421)
	) name4 (
		\addroundkey_round_reg[1]/NET0131 ,
		\addroundkey_round_reg[3]/NET0131 ,
		\round_reg[1]/NET0131 ,
		\round_reg[3]/NET0131 ,
		_w933_
	);
	LUT2 #(
		.INIT('h8)
	) name5 (
		_w932_,
		_w933_,
		_w934_
	);
	LUT3 #(
		.INIT('h01)
	) name6 (
		\addroundkey_round_reg[1]/NET0131 ,
		\addroundkey_round_reg[2]/NET0131 ,
		\addroundkey_round_reg[3]/NET0131 ,
		_w935_
	);
	LUT4 #(
		.INIT('hd500)
	) name7 (
		\ks1_ready_o_reg/NET0131 ,
		_w932_,
		_w933_,
		_w935_,
		_w936_
	);
	LUT3 #(
		.INIT('hc8)
	) name8 (
		\addroundkey_start_i_reg/NET0131 ,
		\key_i[14]_pad ,
		_w936_,
		_w937_
	);
	LUT2 #(
		.INIT('h2)
	) name9 (
		\addroundkey_start_i_reg/NET0131 ,
		_w930_,
		_w938_
	);
	LUT3 #(
		.INIT('h02)
	) name10 (
		\ks1_key_reg_reg[14]/NET0131 ,
		_w936_,
		_w938_,
		_w939_
	);
	LUT4 #(
		.INIT('h0001)
	) name11 (
		\addroundkey_round_reg[1]/NET0131 ,
		\addroundkey_round_reg[2]/NET0131 ,
		\addroundkey_round_reg[3]/NET0131 ,
		\key_i[14]_pad ,
		_w940_
	);
	LUT4 #(
		.INIT('h00fe)
	) name12 (
		\addroundkey_round_reg[1]/NET0131 ,
		\addroundkey_round_reg[2]/NET0131 ,
		\addroundkey_round_reg[3]/NET0131 ,
		\ks1_key_reg_reg[14]/NET0131 ,
		_w941_
	);
	LUT4 #(
		.INIT('h0008)
	) name13 (
		\addroundkey_start_i_reg/NET0131 ,
		_w930_,
		_w941_,
		_w940_,
		_w942_
	);
	LUT4 #(
		.INIT('h00ab)
	) name14 (
		_w931_,
		_w937_,
		_w939_,
		_w942_,
		_w943_
	);
	LUT2 #(
		.INIT('h4)
	) name15 (
		\addroundkey_start_i_reg/NET0131 ,
		\ks1_ready_o_reg/NET0131 ,
		_w944_
	);
	LUT3 #(
		.INIT('h70)
	) name16 (
		_w932_,
		_w933_,
		_w944_,
		_w945_
	);
	LUT2 #(
		.INIT('h1)
	) name17 (
		\ks1_state_reg[0]/NET0131 ,
		\ks1_state_reg[2]/NET0131 ,
		_w946_
	);
	LUT3 #(
		.INIT('h01)
	) name18 (
		\ks1_state_reg[0]/NET0131 ,
		\ks1_state_reg[1]/NET0131 ,
		\ks1_state_reg[2]/NET0131 ,
		_w947_
	);
	LUT3 #(
		.INIT('he0)
	) name19 (
		_w938_,
		_w945_,
		_w947_,
		_w948_
	);
	LUT3 #(
		.INIT('he1)
	) name20 (
		\ks1_state_reg[0]/NET0131 ,
		\ks1_state_reg[1]/NET0131 ,
		\ks1_state_reg[2]/NET0131 ,
		_w949_
	);
	LUT4 #(
		.INIT('h1f00)
	) name21 (
		_w938_,
		_w945_,
		_w947_,
		_w949_,
		_w950_
	);
	LUT2 #(
		.INIT('h8)
	) name22 (
		decrypt_i_pad,
		_w950_,
		_w951_
	);
	LUT4 #(
		.INIT('h953c)
	) name23 (
		\sbox1_to_invert_reg[0]/NET0131 ,
		\sbox1_to_invert_reg[1]/NET0131 ,
		\sbox1_to_invert_reg[2]/NET0131 ,
		\sbox1_to_invert_reg[3]/NET0131 ,
		_w952_
	);
	LUT2 #(
		.INIT('h8)
	) name24 (
		\sbox1_ah_reg_reg[1]/NET0131 ,
		_w952_,
		_w953_
	);
	LUT4 #(
		.INIT('hb689)
	) name25 (
		\sbox1_to_invert_reg[0]/NET0131 ,
		\sbox1_to_invert_reg[1]/NET0131 ,
		\sbox1_to_invert_reg[2]/NET0131 ,
		\sbox1_to_invert_reg[3]/NET0131 ,
		_w954_
	);
	LUT2 #(
		.INIT('h2)
	) name26 (
		\sbox1_ah_reg_reg[0]/NET0131 ,
		_w954_,
		_w955_
	);
	LUT4 #(
		.INIT('h53e8)
	) name27 (
		\sbox1_to_invert_reg[0]/NET0131 ,
		\sbox1_to_invert_reg[1]/NET0131 ,
		\sbox1_to_invert_reg[2]/NET0131 ,
		\sbox1_to_invert_reg[3]/NET0131 ,
		_w956_
	);
	LUT4 #(
		.INIT('hd227)
	) name28 (
		\sbox1_to_invert_reg[0]/NET0131 ,
		\sbox1_to_invert_reg[1]/NET0131 ,
		\sbox1_to_invert_reg[2]/NET0131 ,
		\sbox1_to_invert_reg[3]/NET0131 ,
		_w957_
	);
	LUT4 #(
		.INIT('h3f95)
	) name29 (
		\sbox1_ah_reg_reg[2]/NET0131 ,
		\sbox1_ah_reg_reg[3]/NET0131 ,
		_w956_,
		_w957_,
		_w958_
	);
	LUT3 #(
		.INIT('h69)
	) name30 (
		_w953_,
		_w955_,
		_w958_,
		_w959_
	);
	LUT2 #(
		.INIT('h8)
	) name31 (
		\sbox1_ah_reg_reg[2]/NET0131 ,
		_w956_,
		_w960_
	);
	LUT4 #(
		.INIT('hf359)
	) name32 (
		\sbox1_ah_reg_reg[1]/NET0131 ,
		\sbox1_ah_reg_reg[3]/NET0131 ,
		_w954_,
		_w957_,
		_w961_
	);
	LUT2 #(
		.INIT('h9)
	) name33 (
		\sbox1_ah_reg_reg[0]/NET0131 ,
		\sbox1_ah_reg_reg[3]/NET0131 ,
		_w962_
	);
	LUT2 #(
		.INIT('h2)
	) name34 (
		_w952_,
		_w962_,
		_w963_
	);
	LUT3 #(
		.INIT('h69)
	) name35 (
		_w960_,
		_w961_,
		_w963_,
		_w964_
	);
	LUT4 #(
		.INIT('hb8e4)
	) name36 (
		\sbox1_to_invert_reg[0]/NET0131 ,
		\sbox1_to_invert_reg[1]/NET0131 ,
		\sbox1_to_invert_reg[2]/NET0131 ,
		\sbox1_to_invert_reg[3]/NET0131 ,
		_w965_
	);
	LUT2 #(
		.INIT('h8)
	) name37 (
		\sbox1_ah_reg_reg[3]/NET0131 ,
		_w965_,
		_w966_
	);
	LUT4 #(
		.INIT('hdc4a)
	) name38 (
		\sbox1_to_invert_reg[0]/NET0131 ,
		\sbox1_to_invert_reg[1]/NET0131 ,
		\sbox1_to_invert_reg[2]/NET0131 ,
		\sbox1_to_invert_reg[3]/NET0131 ,
		_w967_
	);
	LUT2 #(
		.INIT('h8)
	) name39 (
		\sbox1_ah_reg_reg[2]/NET0131 ,
		_w967_,
		_w968_
	);
	LUT4 #(
		.INIT('h3f95)
	) name40 (
		\sbox1_ah_reg_reg[0]/NET0131 ,
		\sbox1_ah_reg_reg[1]/NET0131 ,
		_w956_,
		_w957_,
		_w969_
	);
	LUT3 #(
		.INIT('h69)
	) name41 (
		_w966_,
		_w968_,
		_w969_,
		_w970_
	);
	LUT3 #(
		.INIT('h69)
	) name42 (
		_w959_,
		_w964_,
		_w970_,
		_w971_
	);
	LUT2 #(
		.INIT('h8)
	) name43 (
		\sbox1_alph_reg[2]/NET0131 ,
		_w967_,
		_w972_
	);
	LUT2 #(
		.INIT('h8)
	) name44 (
		\sbox1_alph_reg[1]/NET0131 ,
		_w956_,
		_w973_
	);
	LUT4 #(
		.INIT('h39f5)
	) name45 (
		\sbox1_alph_reg[0]/NET0131 ,
		\sbox1_alph_reg[3]/NET0131 ,
		_w957_,
		_w965_,
		_w974_
	);
	LUT3 #(
		.INIT('h69)
	) name46 (
		_w972_,
		_w973_,
		_w974_,
		_w975_
	);
	LUT4 #(
		.INIT('h953f)
	) name47 (
		\sbox1_alph_reg[1]/NET0131 ,
		\sbox1_alph_reg[2]/NET0131 ,
		_w965_,
		_w967_,
		_w976_
	);
	LUT4 #(
		.INIT('h60ac)
	) name48 (
		\sbox1_alph_reg[0]/NET0131 ,
		\sbox1_alph_reg[3]/NET0131 ,
		_w956_,
		_w957_,
		_w977_
	);
	LUT2 #(
		.INIT('h9)
	) name49 (
		_w976_,
		_w977_,
		_w978_
	);
	LUT2 #(
		.INIT('h8)
	) name50 (
		\sbox1_alph_reg[0]/NET0131 ,
		_w952_,
		_w979_
	);
	LUT2 #(
		.INIT('h8)
	) name51 (
		\sbox1_alph_reg[3]/NET0131 ,
		_w967_,
		_w980_
	);
	LUT4 #(
		.INIT('h3f95)
	) name52 (
		\sbox1_alph_reg[1]/NET0131 ,
		\sbox1_alph_reg[2]/NET0131 ,
		_w956_,
		_w957_,
		_w981_
	);
	LUT3 #(
		.INIT('h96)
	) name53 (
		_w979_,
		_w980_,
		_w981_,
		_w982_
	);
	LUT2 #(
		.INIT('h6)
	) name54 (
		_w978_,
		_w982_,
		_w983_
	);
	LUT4 #(
		.INIT('h6996)
	) name55 (
		_w964_,
		_w975_,
		_w978_,
		_w982_,
		_w984_
	);
	LUT4 #(
		.INIT('h278d)
	) name56 (
		_w951_,
		_w959_,
		_w971_,
		_w984_,
		_w985_
	);
	LUT4 #(
		.INIT('h80f0)
	) name57 (
		_w932_,
		_w933_,
		_w935_,
		_w944_,
		_w986_
	);
	LUT4 #(
		.INIT('haaac)
	) name58 (
		\key_i[110]_pad ,
		\ks1_key_reg_reg[110]/P0002 ,
		_w938_,
		_w986_,
		_w987_
	);
	LUT2 #(
		.INIT('h9)
	) name59 (
		_w985_,
		_w987_,
		_w988_
	);
	LUT4 #(
		.INIT('haaac)
	) name60 (
		\key_i[78]_pad ,
		\ks1_key_reg_reg[78]/P0002 ,
		_w938_,
		_w986_,
		_w989_
	);
	LUT3 #(
		.INIT('h69)
	) name61 (
		_w985_,
		_w987_,
		_w989_,
		_w990_
	);
	LUT4 #(
		.INIT('haaac)
	) name62 (
		\key_i[46]_pad ,
		\ks1_key_reg_reg[46]/P0002 ,
		_w938_,
		_w986_,
		_w991_
	);
	LUT4 #(
		.INIT('h9669)
	) name63 (
		_w985_,
		_w987_,
		_w989_,
		_w991_,
		_w992_
	);
	LUT4 #(
		.INIT('he22e)
	) name64 (
		\ks1_key_reg_reg[14]/NET0131 ,
		_w929_,
		_w943_,
		_w992_,
		_w993_
	);
	LUT2 #(
		.INIT('h4)
	) name65 (
		\round_reg[2]/NET0131 ,
		\round_reg[3]/NET0131 ,
		_w994_
	);
	LUT4 #(
		.INIT('h0400)
	) name66 (
		\round_reg[0]/NET0131 ,
		\round_reg[1]/NET0131 ,
		\round_reg[2]/NET0131 ,
		\round_reg[3]/NET0131 ,
		_w995_
	);
	LUT2 #(
		.INIT('h2)
	) name67 (
		decrypt_i_pad,
		_w995_,
		_w996_
	);
	LUT3 #(
		.INIT('h02)
	) name68 (
		decrypt_i_pad,
		\mix1_data_o_reg_reg[60]/NET0131 ,
		_w995_,
		_w997_
	);
	LUT3 #(
		.INIT('h01)
	) name69 (
		\sub1_state_reg[0]/NET0131 ,
		\sub1_state_reg[1]/NET0131 ,
		\sub1_state_reg[2]/NET0131 ,
		_w998_
	);
	LUT4 #(
		.INIT('h0100)
	) name70 (
		\sub1_state_reg[0]/NET0131 ,
		\sub1_state_reg[1]/NET0131 ,
		\sub1_state_reg[2]/NET0131 ,
		\sub1_state_reg[3]/NET0131 ,
		_w999_
	);
	LUT4 #(
		.INIT('hae00)
	) name71 (
		\data_o[60]_pad ,
		decrypt_i_pad,
		_w995_,
		_w999_,
		_w1000_
	);
	LUT3 #(
		.INIT('h02)
	) name72 (
		decrypt_i_pad,
		\mix1_data_o_reg_reg[116]/NET0131 ,
		_w995_,
		_w1001_
	);
	LUT4 #(
		.INIT('h0002)
	) name73 (
		\sub1_state_reg[0]/NET0131 ,
		\sub1_state_reg[1]/NET0131 ,
		\sub1_state_reg[2]/NET0131 ,
		\sub1_state_reg[3]/NET0131 ,
		_w1002_
	);
	LUT4 #(
		.INIT('hae00)
	) name74 (
		\data_o[116]_pad ,
		decrypt_i_pad,
		_w995_,
		_w1002_,
		_w1003_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name75 (
		_w997_,
		_w1000_,
		_w1001_,
		_w1003_,
		_w1004_
	);
	LUT3 #(
		.INIT('h02)
	) name76 (
		decrypt_i_pad,
		\mix1_data_o_reg_reg[44]/NET0131 ,
		_w995_,
		_w1005_
	);
	LUT4 #(
		.INIT('h0400)
	) name77 (
		\sub1_state_reg[0]/NET0131 ,
		\sub1_state_reg[1]/NET0131 ,
		\sub1_state_reg[2]/NET0131 ,
		\sub1_state_reg[3]/NET0131 ,
		_w1006_
	);
	LUT4 #(
		.INIT('hae00)
	) name78 (
		\data_o[44]_pad ,
		decrypt_i_pad,
		_w995_,
		_w1006_,
		_w1007_
	);
	LUT3 #(
		.INIT('h02)
	) name79 (
		decrypt_i_pad,
		\mix1_data_o_reg_reg[4]/NET0131 ,
		_w995_,
		_w1008_
	);
	LUT4 #(
		.INIT('h8000)
	) name80 (
		\sub1_state_reg[0]/NET0131 ,
		\sub1_state_reg[1]/NET0131 ,
		\sub1_state_reg[2]/NET0131 ,
		\sub1_state_reg[3]/NET0131 ,
		_w1009_
	);
	LUT4 #(
		.INIT('hae00)
	) name81 (
		\data_o[4]_pad ,
		decrypt_i_pad,
		_w995_,
		_w1009_,
		_w1010_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name82 (
		_w1005_,
		_w1007_,
		_w1008_,
		_w1010_,
		_w1011_
	);
	LUT3 #(
		.INIT('h02)
	) name83 (
		decrypt_i_pad,
		\mix1_data_o_reg_reg[12]/NET0131 ,
		_w995_,
		_w1012_
	);
	LUT4 #(
		.INIT('h4000)
	) name84 (
		\sub1_state_reg[0]/NET0131 ,
		\sub1_state_reg[1]/NET0131 ,
		\sub1_state_reg[2]/NET0131 ,
		\sub1_state_reg[3]/NET0131 ,
		_w1013_
	);
	LUT4 #(
		.INIT('ha0e0)
	) name85 (
		\data_o[12]_pad ,
		decrypt_i_pad,
		_w1013_,
		_w995_,
		_w1014_
	);
	LUT3 #(
		.INIT('h02)
	) name86 (
		decrypt_i_pad,
		\mix1_data_o_reg_reg[100]/NET0131 ,
		_w995_,
		_w1015_
	);
	LUT4 #(
		.INIT('h0008)
	) name87 (
		\sub1_state_reg[0]/NET0131 ,
		\sub1_state_reg[1]/NET0131 ,
		\sub1_state_reg[2]/NET0131 ,
		\sub1_state_reg[3]/NET0131 ,
		_w1016_
	);
	LUT4 #(
		.INIT('hae00)
	) name88 (
		\data_o[100]_pad ,
		decrypt_i_pad,
		_w995_,
		_w1016_,
		_w1017_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name89 (
		_w1012_,
		_w1014_,
		_w1015_,
		_w1017_,
		_w1018_
	);
	LUT3 #(
		.INIT('h02)
	) name90 (
		decrypt_i_pad,
		\mix1_data_o_reg_reg[28]/NET0131 ,
		_w995_,
		_w1019_
	);
	LUT4 #(
		.INIT('h1000)
	) name91 (
		\sub1_state_reg[0]/NET0131 ,
		\sub1_state_reg[1]/NET0131 ,
		\sub1_state_reg[2]/NET0131 ,
		\sub1_state_reg[3]/NET0131 ,
		_w1020_
	);
	LUT4 #(
		.INIT('hae00)
	) name92 (
		\data_o[28]_pad ,
		decrypt_i_pad,
		_w995_,
		_w1020_,
		_w1021_
	);
	LUT3 #(
		.INIT('h02)
	) name93 (
		decrypt_i_pad,
		\mix1_data_o_reg_reg[20]/NET0131 ,
		_w995_,
		_w1022_
	);
	LUT4 #(
		.INIT('h2000)
	) name94 (
		\sub1_state_reg[0]/NET0131 ,
		\sub1_state_reg[1]/NET0131 ,
		\sub1_state_reg[2]/NET0131 ,
		\sub1_state_reg[3]/NET0131 ,
		_w1023_
	);
	LUT4 #(
		.INIT('hae00)
	) name95 (
		\data_o[20]_pad ,
		decrypt_i_pad,
		_w995_,
		_w1023_,
		_w1024_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name96 (
		_w1019_,
		_w1021_,
		_w1022_,
		_w1024_,
		_w1025_
	);
	LUT4 #(
		.INIT('h8000)
	) name97 (
		_w1018_,
		_w1025_,
		_w1004_,
		_w1011_,
		_w1026_
	);
	LUT3 #(
		.INIT('h02)
	) name98 (
		decrypt_i_pad,
		\mix1_data_o_reg_reg[108]/NET0131 ,
		_w995_,
		_w1027_
	);
	LUT4 #(
		.INIT('h0004)
	) name99 (
		\sub1_state_reg[0]/NET0131 ,
		\sub1_state_reg[1]/NET0131 ,
		\sub1_state_reg[2]/NET0131 ,
		\sub1_state_reg[3]/NET0131 ,
		_w1028_
	);
	LUT4 #(
		.INIT('hae00)
	) name100 (
		\data_o[108]_pad ,
		decrypt_i_pad,
		_w995_,
		_w1028_,
		_w1029_
	);
	LUT2 #(
		.INIT('h4)
	) name101 (
		_w1027_,
		_w1029_,
		_w1030_
	);
	LUT3 #(
		.INIT('h02)
	) name102 (
		decrypt_i_pad,
		\mix1_data_o_reg_reg[92]/NET0131 ,
		_w995_,
		_w1031_
	);
	LUT4 #(
		.INIT('h0010)
	) name103 (
		\sub1_state_reg[0]/NET0131 ,
		\sub1_state_reg[1]/NET0131 ,
		\sub1_state_reg[2]/NET0131 ,
		\sub1_state_reg[3]/NET0131 ,
		_w1032_
	);
	LUT4 #(
		.INIT('hae00)
	) name104 (
		\data_o[92]_pad ,
		decrypt_i_pad,
		_w995_,
		_w1032_,
		_w1033_
	);
	LUT3 #(
		.INIT('h02)
	) name105 (
		decrypt_i_pad,
		\mix1_data_o_reg_reg[76]/NET0131 ,
		_w995_,
		_w1034_
	);
	LUT4 #(
		.INIT('h0040)
	) name106 (
		\sub1_state_reg[0]/NET0131 ,
		\sub1_state_reg[1]/NET0131 ,
		\sub1_state_reg[2]/NET0131 ,
		\sub1_state_reg[3]/NET0131 ,
		_w1035_
	);
	LUT4 #(
		.INIT('hae00)
	) name107 (
		\data_o[76]_pad ,
		decrypt_i_pad,
		_w995_,
		_w1035_,
		_w1036_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name108 (
		_w1031_,
		_w1033_,
		_w1034_,
		_w1036_,
		_w1037_
	);
	LUT3 #(
		.INIT('h02)
	) name109 (
		decrypt_i_pad,
		\mix1_data_o_reg_reg[68]/NET0131 ,
		_w995_,
		_w1038_
	);
	LUT4 #(
		.INIT('h0080)
	) name110 (
		\sub1_state_reg[0]/NET0131 ,
		\sub1_state_reg[1]/NET0131 ,
		\sub1_state_reg[2]/NET0131 ,
		\sub1_state_reg[3]/NET0131 ,
		_w1039_
	);
	LUT4 #(
		.INIT('hae00)
	) name111 (
		\data_o[68]_pad ,
		decrypt_i_pad,
		_w995_,
		_w1039_,
		_w1040_
	);
	LUT3 #(
		.INIT('h02)
	) name112 (
		decrypt_i_pad,
		\mix1_data_o_reg_reg[36]/NET0131 ,
		_w995_,
		_w1041_
	);
	LUT4 #(
		.INIT('h0800)
	) name113 (
		\sub1_state_reg[0]/NET0131 ,
		\sub1_state_reg[1]/NET0131 ,
		\sub1_state_reg[2]/NET0131 ,
		\sub1_state_reg[3]/NET0131 ,
		_w1042_
	);
	LUT4 #(
		.INIT('hae00)
	) name114 (
		\data_o[36]_pad ,
		decrypt_i_pad,
		_w995_,
		_w1042_,
		_w1043_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name115 (
		_w1038_,
		_w1040_,
		_w1041_,
		_w1043_,
		_w1044_
	);
	LUT3 #(
		.INIT('h02)
	) name116 (
		decrypt_i_pad,
		\mix1_data_o_reg_reg[52]/NET0131 ,
		_w995_,
		_w1045_
	);
	LUT4 #(
		.INIT('h0200)
	) name117 (
		\sub1_state_reg[0]/NET0131 ,
		\sub1_state_reg[1]/NET0131 ,
		\sub1_state_reg[2]/NET0131 ,
		\sub1_state_reg[3]/NET0131 ,
		_w1046_
	);
	LUT4 #(
		.INIT('hae00)
	) name118 (
		\data_o[52]_pad ,
		decrypt_i_pad,
		_w995_,
		_w1046_,
		_w1047_
	);
	LUT3 #(
		.INIT('h02)
	) name119 (
		decrypt_i_pad,
		\mix1_data_o_reg_reg[84]/NET0131 ,
		_w995_,
		_w1048_
	);
	LUT4 #(
		.INIT('h0020)
	) name120 (
		\sub1_state_reg[0]/NET0131 ,
		\sub1_state_reg[1]/NET0131 ,
		\sub1_state_reg[2]/NET0131 ,
		\sub1_state_reg[3]/NET0131 ,
		_w1049_
	);
	LUT4 #(
		.INIT('hae00)
	) name121 (
		\data_o[84]_pad ,
		decrypt_i_pad,
		_w995_,
		_w1049_,
		_w1050_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name122 (
		_w1045_,
		_w1047_,
		_w1048_,
		_w1050_,
		_w1051_
	);
	LUT4 #(
		.INIT('h4000)
	) name123 (
		_w1030_,
		_w1044_,
		_w1051_,
		_w1037_,
		_w1052_
	);
	LUT4 #(
		.INIT('h0001)
	) name124 (
		\sub1_state_reg[0]/NET0131 ,
		\sub1_state_reg[1]/NET0131 ,
		\sub1_state_reg[2]/NET0131 ,
		\sub1_state_reg[3]/NET0131 ,
		_w1053_
	);
	LUT3 #(
		.INIT('h27)
	) name125 (
		decrypt_i_pad,
		_w930_,
		_w995_,
		_w1054_
	);
	LUT4 #(
		.INIT('hc480)
	) name126 (
		decrypt_i_pad,
		\state_reg/NET0131 ,
		_w930_,
		_w995_,
		_w1055_
	);
	LUT4 #(
		.INIT('h151d)
	) name127 (
		\addroundkey_ready_o_reg/NET0131 ,
		decrypt_i_pad,
		\mix1_ready_o_reg/NET0131 ,
		_w995_,
		_w1056_
	);
	LUT2 #(
		.INIT('h1)
	) name128 (
		_w1055_,
		_w1056_,
		_w1057_
	);
	LUT3 #(
		.INIT('h51)
	) name129 (
		\data_o[124]_pad ,
		decrypt_i_pad,
		_w995_,
		_w1058_
	);
	LUT3 #(
		.INIT('h02)
	) name130 (
		decrypt_i_pad,
		\mix1_data_o_reg_reg[124]/NET0131 ,
		_w995_,
		_w1059_
	);
	LUT2 #(
		.INIT('h4)
	) name131 (
		\sub1_state_reg[4]/NET0131 ,
		_w1053_,
		_w1060_
	);
	LUT3 #(
		.INIT('h04)
	) name132 (
		_w1059_,
		_w1060_,
		_w1058_,
		_w1061_
	);
	LUT2 #(
		.INIT('h8)
	) name133 (
		_w1057_,
		_w1061_,
		_w1062_
	);
	LUT4 #(
		.INIT('h00f8)
	) name134 (
		_w1026_,
		_w1052_,
		_w1053_,
		_w1062_,
		_w1063_
	);
	LUT3 #(
		.INIT('h08)
	) name135 (
		\ks1_state_reg[0]/NET0131 ,
		\ks1_state_reg[1]/NET0131 ,
		\ks1_state_reg[2]/NET0131 ,
		_w1064_
	);
	LUT3 #(
		.INIT('hc8)
	) name136 (
		\addroundkey_start_i_reg/NET0131 ,
		\key_i[4]_pad ,
		_w936_,
		_w1065_
	);
	LUT3 #(
		.INIT('h02)
	) name137 (
		\ks1_key_reg_reg[4]/NET0131 ,
		_w936_,
		_w938_,
		_w1066_
	);
	LUT4 #(
		.INIT('h0001)
	) name138 (
		\addroundkey_round_reg[1]/NET0131 ,
		\addroundkey_round_reg[2]/NET0131 ,
		\addroundkey_round_reg[3]/NET0131 ,
		\key_i[4]_pad ,
		_w1067_
	);
	LUT4 #(
		.INIT('h00fe)
	) name139 (
		\addroundkey_round_reg[1]/NET0131 ,
		\addroundkey_round_reg[2]/NET0131 ,
		\addroundkey_round_reg[3]/NET0131 ,
		\ks1_key_reg_reg[4]/NET0131 ,
		_w1068_
	);
	LUT4 #(
		.INIT('h0008)
	) name140 (
		\addroundkey_start_i_reg/NET0131 ,
		_w930_,
		_w1068_,
		_w1067_,
		_w1069_
	);
	LUT4 #(
		.INIT('h00ab)
	) name141 (
		_w931_,
		_w1065_,
		_w1066_,
		_w1069_,
		_w1070_
	);
	LUT3 #(
		.INIT('h04)
	) name142 (
		\ks1_state_reg[0]/NET0131 ,
		\ks1_state_reg[1]/NET0131 ,
		\ks1_state_reg[2]/NET0131 ,
		_w1071_
	);
	LUT3 #(
		.INIT('hc8)
	) name143 (
		\addroundkey_start_i_reg/NET0131 ,
		\key_i[12]_pad ,
		_w936_,
		_w1072_
	);
	LUT3 #(
		.INIT('h02)
	) name144 (
		\ks1_key_reg_reg[12]/NET0131 ,
		_w936_,
		_w938_,
		_w1073_
	);
	LUT4 #(
		.INIT('h0001)
	) name145 (
		\addroundkey_round_reg[1]/NET0131 ,
		\addroundkey_round_reg[2]/NET0131 ,
		\addroundkey_round_reg[3]/NET0131 ,
		\key_i[12]_pad ,
		_w1074_
	);
	LUT4 #(
		.INIT('h00fe)
	) name146 (
		\addroundkey_round_reg[1]/NET0131 ,
		\addroundkey_round_reg[2]/NET0131 ,
		\addroundkey_round_reg[3]/NET0131 ,
		\ks1_key_reg_reg[12]/NET0131 ,
		_w1075_
	);
	LUT4 #(
		.INIT('h0008)
	) name147 (
		\addroundkey_start_i_reg/NET0131 ,
		_w930_,
		_w1075_,
		_w1074_,
		_w1076_
	);
	LUT4 #(
		.INIT('h00ab)
	) name148 (
		_w931_,
		_w1072_,
		_w1073_,
		_w1076_,
		_w1077_
	);
	LUT4 #(
		.INIT('hdd0d)
	) name149 (
		_w1064_,
		_w1070_,
		_w1071_,
		_w1077_,
		_w1078_
	);
	LUT3 #(
		.INIT('h02)
	) name150 (
		\ks1_state_reg[0]/NET0131 ,
		\ks1_state_reg[1]/NET0131 ,
		\ks1_state_reg[2]/NET0131 ,
		_w1079_
	);
	LUT3 #(
		.INIT('hc8)
	) name151 (
		\addroundkey_start_i_reg/NET0131 ,
		\key_i[20]_pad ,
		_w936_,
		_w1080_
	);
	LUT3 #(
		.INIT('h02)
	) name152 (
		\ks1_key_reg_reg[20]/NET0131 ,
		_w936_,
		_w938_,
		_w1081_
	);
	LUT4 #(
		.INIT('h0001)
	) name153 (
		\addroundkey_round_reg[1]/NET0131 ,
		\addroundkey_round_reg[2]/NET0131 ,
		\addroundkey_round_reg[3]/NET0131 ,
		\key_i[20]_pad ,
		_w1082_
	);
	LUT4 #(
		.INIT('h00fe)
	) name154 (
		\addroundkey_round_reg[1]/NET0131 ,
		\addroundkey_round_reg[2]/NET0131 ,
		\addroundkey_round_reg[3]/NET0131 ,
		\ks1_key_reg_reg[20]/NET0131 ,
		_w1083_
	);
	LUT4 #(
		.INIT('h0008)
	) name155 (
		\addroundkey_start_i_reg/NET0131 ,
		_w930_,
		_w1083_,
		_w1082_,
		_w1084_
	);
	LUT4 #(
		.INIT('h00ab)
	) name156 (
		_w931_,
		_w1080_,
		_w1081_,
		_w1084_,
		_w1085_
	);
	LUT3 #(
		.INIT('hc8)
	) name157 (
		\addroundkey_start_i_reg/NET0131 ,
		\key_i[28]_pad ,
		_w936_,
		_w1086_
	);
	LUT3 #(
		.INIT('h02)
	) name158 (
		\ks1_key_reg_reg[28]/NET0131 ,
		_w936_,
		_w938_,
		_w1087_
	);
	LUT4 #(
		.INIT('h0001)
	) name159 (
		\addroundkey_round_reg[1]/NET0131 ,
		\addroundkey_round_reg[2]/NET0131 ,
		\addroundkey_round_reg[3]/NET0131 ,
		\key_i[28]_pad ,
		_w1088_
	);
	LUT4 #(
		.INIT('h00fe)
	) name160 (
		\addroundkey_round_reg[1]/NET0131 ,
		\addroundkey_round_reg[2]/NET0131 ,
		\addroundkey_round_reg[3]/NET0131 ,
		\ks1_key_reg_reg[28]/NET0131 ,
		_w1089_
	);
	LUT4 #(
		.INIT('h0008)
	) name161 (
		\addroundkey_start_i_reg/NET0131 ,
		_w930_,
		_w1089_,
		_w1088_,
		_w1090_
	);
	LUT4 #(
		.INIT('h00ab)
	) name162 (
		_w931_,
		_w1086_,
		_w1087_,
		_w1090_,
		_w1091_
	);
	LUT4 #(
		.INIT('hf351)
	) name163 (
		_w948_,
		_w1079_,
		_w1085_,
		_w1091_,
		_w1092_
	);
	LUT4 #(
		.INIT('hd000)
	) name164 (
		_w950_,
		_w1063_,
		_w1078_,
		_w1092_,
		_w1093_
	);
	LUT2 #(
		.INIT('h1)
	) name165 (
		_w951_,
		_w1093_,
		_w1094_
	);
	LUT3 #(
		.INIT('h02)
	) name166 (
		decrypt_i_pad,
		\mix1_data_o_reg_reg[70]/NET0131 ,
		_w995_,
		_w1095_
	);
	LUT4 #(
		.INIT('hae00)
	) name167 (
		\data_o[70]_pad ,
		decrypt_i_pad,
		_w995_,
		_w1039_,
		_w1096_
	);
	LUT3 #(
		.INIT('h02)
	) name168 (
		decrypt_i_pad,
		\mix1_data_o_reg_reg[30]/NET0131 ,
		_w995_,
		_w1097_
	);
	LUT4 #(
		.INIT('hae00)
	) name169 (
		\data_o[30]_pad ,
		decrypt_i_pad,
		_w995_,
		_w1020_,
		_w1098_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name170 (
		_w1095_,
		_w1096_,
		_w1097_,
		_w1098_,
		_w1099_
	);
	LUT3 #(
		.INIT('h02)
	) name171 (
		decrypt_i_pad,
		\mix1_data_o_reg_reg[54]/NET0131 ,
		_w995_,
		_w1100_
	);
	LUT4 #(
		.INIT('hae00)
	) name172 (
		\data_o[54]_pad ,
		decrypt_i_pad,
		_w995_,
		_w1046_,
		_w1101_
	);
	LUT3 #(
		.INIT('h02)
	) name173 (
		decrypt_i_pad,
		\mix1_data_o_reg_reg[22]/NET0131 ,
		_w995_,
		_w1102_
	);
	LUT4 #(
		.INIT('hae00)
	) name174 (
		\data_o[22]_pad ,
		decrypt_i_pad,
		_w995_,
		_w1023_,
		_w1103_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name175 (
		_w1100_,
		_w1101_,
		_w1102_,
		_w1103_,
		_w1104_
	);
	LUT3 #(
		.INIT('h02)
	) name176 (
		decrypt_i_pad,
		\mix1_data_o_reg_reg[118]/NET0131 ,
		_w995_,
		_w1105_
	);
	LUT4 #(
		.INIT('hae00)
	) name177 (
		\data_o[118]_pad ,
		decrypt_i_pad,
		_w995_,
		_w1002_,
		_w1106_
	);
	LUT3 #(
		.INIT('h02)
	) name178 (
		decrypt_i_pad,
		\mix1_data_o_reg_reg[110]/NET0131 ,
		_w995_,
		_w1107_
	);
	LUT4 #(
		.INIT('hae00)
	) name179 (
		\data_o[110]_pad ,
		decrypt_i_pad,
		_w995_,
		_w1028_,
		_w1108_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name180 (
		_w1105_,
		_w1106_,
		_w1107_,
		_w1108_,
		_w1109_
	);
	LUT3 #(
		.INIT('h02)
	) name181 (
		decrypt_i_pad,
		\mix1_data_o_reg_reg[102]/NET0131 ,
		_w995_,
		_w1110_
	);
	LUT4 #(
		.INIT('hae00)
	) name182 (
		\data_o[102]_pad ,
		decrypt_i_pad,
		_w995_,
		_w1016_,
		_w1111_
	);
	LUT3 #(
		.INIT('h02)
	) name183 (
		decrypt_i_pad,
		\mix1_data_o_reg_reg[46]/NET0131 ,
		_w995_,
		_w1112_
	);
	LUT4 #(
		.INIT('hae00)
	) name184 (
		\data_o[46]_pad ,
		decrypt_i_pad,
		_w995_,
		_w1006_,
		_w1113_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name185 (
		_w1110_,
		_w1111_,
		_w1112_,
		_w1113_,
		_w1114_
	);
	LUT4 #(
		.INIT('h8000)
	) name186 (
		_w1109_,
		_w1114_,
		_w1099_,
		_w1104_,
		_w1115_
	);
	LUT3 #(
		.INIT('h02)
	) name187 (
		decrypt_i_pad,
		\mix1_data_o_reg_reg[14]/NET0131 ,
		_w995_,
		_w1116_
	);
	LUT4 #(
		.INIT('ha0e0)
	) name188 (
		\data_o[14]_pad ,
		decrypt_i_pad,
		_w1013_,
		_w995_,
		_w1117_
	);
	LUT2 #(
		.INIT('h4)
	) name189 (
		_w1116_,
		_w1117_,
		_w1118_
	);
	LUT3 #(
		.INIT('h02)
	) name190 (
		decrypt_i_pad,
		\mix1_data_o_reg_reg[62]/NET0131 ,
		_w995_,
		_w1119_
	);
	LUT4 #(
		.INIT('hae00)
	) name191 (
		\data_o[62]_pad ,
		decrypt_i_pad,
		_w995_,
		_w999_,
		_w1120_
	);
	LUT3 #(
		.INIT('h02)
	) name192 (
		decrypt_i_pad,
		\mix1_data_o_reg_reg[86]/NET0131 ,
		_w995_,
		_w1121_
	);
	LUT4 #(
		.INIT('hae00)
	) name193 (
		\data_o[86]_pad ,
		decrypt_i_pad,
		_w995_,
		_w1049_,
		_w1122_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name194 (
		_w1119_,
		_w1120_,
		_w1121_,
		_w1122_,
		_w1123_
	);
	LUT3 #(
		.INIT('h02)
	) name195 (
		decrypt_i_pad,
		\mix1_data_o_reg_reg[6]/NET0131 ,
		_w995_,
		_w1124_
	);
	LUT4 #(
		.INIT('hae00)
	) name196 (
		\data_o[6]_pad ,
		decrypt_i_pad,
		_w995_,
		_w1009_,
		_w1125_
	);
	LUT3 #(
		.INIT('h02)
	) name197 (
		decrypt_i_pad,
		\mix1_data_o_reg_reg[94]/NET0131 ,
		_w995_,
		_w1126_
	);
	LUT4 #(
		.INIT('hae00)
	) name198 (
		\data_o[94]_pad ,
		decrypt_i_pad,
		_w995_,
		_w1032_,
		_w1127_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name199 (
		_w1124_,
		_w1125_,
		_w1126_,
		_w1127_,
		_w1128_
	);
	LUT3 #(
		.INIT('h02)
	) name200 (
		decrypt_i_pad,
		\mix1_data_o_reg_reg[78]/NET0131 ,
		_w995_,
		_w1129_
	);
	LUT4 #(
		.INIT('hae00)
	) name201 (
		\data_o[78]_pad ,
		decrypt_i_pad,
		_w995_,
		_w1035_,
		_w1130_
	);
	LUT3 #(
		.INIT('h02)
	) name202 (
		decrypt_i_pad,
		\mix1_data_o_reg_reg[38]/NET0131 ,
		_w995_,
		_w1131_
	);
	LUT4 #(
		.INIT('hae00)
	) name203 (
		\data_o[38]_pad ,
		decrypt_i_pad,
		_w995_,
		_w1042_,
		_w1132_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name204 (
		_w1129_,
		_w1130_,
		_w1131_,
		_w1132_,
		_w1133_
	);
	LUT4 #(
		.INIT('h4000)
	) name205 (
		_w1118_,
		_w1128_,
		_w1133_,
		_w1123_,
		_w1134_
	);
	LUT3 #(
		.INIT('h51)
	) name206 (
		\data_o[126]_pad ,
		decrypt_i_pad,
		_w995_,
		_w1135_
	);
	LUT3 #(
		.INIT('h02)
	) name207 (
		decrypt_i_pad,
		\mix1_data_o_reg_reg[126]/NET0131 ,
		_w995_,
		_w1136_
	);
	LUT3 #(
		.INIT('h02)
	) name208 (
		_w1060_,
		_w1136_,
		_w1135_,
		_w1137_
	);
	LUT2 #(
		.INIT('h8)
	) name209 (
		_w1057_,
		_w1137_,
		_w1138_
	);
	LUT4 #(
		.INIT('h00ea)
	) name210 (
		_w1053_,
		_w1115_,
		_w1134_,
		_w1138_,
		_w1139_
	);
	LUT2 #(
		.INIT('h4)
	) name211 (
		_w943_,
		_w1071_,
		_w1140_
	);
	LUT3 #(
		.INIT('hc8)
	) name212 (
		\addroundkey_start_i_reg/NET0131 ,
		\key_i[30]_pad ,
		_w936_,
		_w1141_
	);
	LUT3 #(
		.INIT('h02)
	) name213 (
		\ks1_key_reg_reg[30]/NET0131 ,
		_w936_,
		_w938_,
		_w1142_
	);
	LUT4 #(
		.INIT('h0001)
	) name214 (
		\addroundkey_round_reg[1]/NET0131 ,
		\addroundkey_round_reg[2]/NET0131 ,
		\addroundkey_round_reg[3]/NET0131 ,
		\key_i[30]_pad ,
		_w1143_
	);
	LUT4 #(
		.INIT('h00fe)
	) name215 (
		\addroundkey_round_reg[1]/NET0131 ,
		\addroundkey_round_reg[2]/NET0131 ,
		\addroundkey_round_reg[3]/NET0131 ,
		\ks1_key_reg_reg[30]/NET0131 ,
		_w1144_
	);
	LUT4 #(
		.INIT('h0008)
	) name216 (
		\addroundkey_start_i_reg/NET0131 ,
		_w930_,
		_w1144_,
		_w1143_,
		_w1145_
	);
	LUT4 #(
		.INIT('h00ab)
	) name217 (
		_w931_,
		_w1141_,
		_w1142_,
		_w1145_,
		_w1146_
	);
	LUT4 #(
		.INIT('h5553)
	) name218 (
		\key_i[6]_pad ,
		\ks1_key_reg_reg[6]/NET0131 ,
		_w938_,
		_w986_,
		_w1147_
	);
	LUT4 #(
		.INIT('h5553)
	) name219 (
		\key_i[22]_pad ,
		\ks1_key_reg_reg[22]/NET0131 ,
		_w938_,
		_w986_,
		_w1148_
	);
	LUT4 #(
		.INIT('hf531)
	) name220 (
		_w1064_,
		_w1079_,
		_w1147_,
		_w1148_,
		_w1149_
	);
	LUT3 #(
		.INIT('hd0)
	) name221 (
		_w948_,
		_w1146_,
		_w1149_,
		_w1150_
	);
	LUT4 #(
		.INIT('h0d00)
	) name222 (
		_w950_,
		_w1139_,
		_w1140_,
		_w1150_,
		_w1151_
	);
	LUT3 #(
		.INIT('h02)
	) name223 (
		decrypt_i_pad,
		\mix1_data_o_reg_reg[67]/NET0131 ,
		_w995_,
		_w1152_
	);
	LUT4 #(
		.INIT('hae00)
	) name224 (
		\data_o[67]_pad ,
		decrypt_i_pad,
		_w995_,
		_w1039_,
		_w1153_
	);
	LUT3 #(
		.INIT('h02)
	) name225 (
		decrypt_i_pad,
		\mix1_data_o_reg_reg[115]/NET0131 ,
		_w995_,
		_w1154_
	);
	LUT4 #(
		.INIT('hae00)
	) name226 (
		\data_o[115]_pad ,
		decrypt_i_pad,
		_w995_,
		_w1002_,
		_w1155_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name227 (
		_w1152_,
		_w1153_,
		_w1154_,
		_w1155_,
		_w1156_
	);
	LUT3 #(
		.INIT('h02)
	) name228 (
		decrypt_i_pad,
		\mix1_data_o_reg_reg[43]/NET0131 ,
		_w995_,
		_w1157_
	);
	LUT4 #(
		.INIT('hae00)
	) name229 (
		\data_o[43]_pad ,
		decrypt_i_pad,
		_w995_,
		_w1006_,
		_w1158_
	);
	LUT3 #(
		.INIT('h02)
	) name230 (
		decrypt_i_pad,
		\mix1_data_o_reg_reg[51]/NET0131 ,
		_w995_,
		_w1159_
	);
	LUT4 #(
		.INIT('hae00)
	) name231 (
		\data_o[51]_pad ,
		decrypt_i_pad,
		_w995_,
		_w1046_,
		_w1160_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name232 (
		_w1157_,
		_w1158_,
		_w1159_,
		_w1160_,
		_w1161_
	);
	LUT3 #(
		.INIT('h02)
	) name233 (
		decrypt_i_pad,
		\mix1_data_o_reg_reg[99]/NET0131 ,
		_w995_,
		_w1162_
	);
	LUT4 #(
		.INIT('hae00)
	) name234 (
		\data_o[99]_pad ,
		decrypt_i_pad,
		_w995_,
		_w1016_,
		_w1163_
	);
	LUT3 #(
		.INIT('h02)
	) name235 (
		decrypt_i_pad,
		\mix1_data_o_reg_reg[83]/NET0131 ,
		_w995_,
		_w1164_
	);
	LUT4 #(
		.INIT('hae00)
	) name236 (
		\data_o[83]_pad ,
		decrypt_i_pad,
		_w995_,
		_w1049_,
		_w1165_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name237 (
		_w1162_,
		_w1163_,
		_w1164_,
		_w1165_,
		_w1166_
	);
	LUT3 #(
		.INIT('h02)
	) name238 (
		decrypt_i_pad,
		\mix1_data_o_reg_reg[35]/NET0131 ,
		_w995_,
		_w1167_
	);
	LUT4 #(
		.INIT('hae00)
	) name239 (
		\data_o[35]_pad ,
		decrypt_i_pad,
		_w995_,
		_w1042_,
		_w1168_
	);
	LUT3 #(
		.INIT('h02)
	) name240 (
		decrypt_i_pad,
		\mix1_data_o_reg_reg[91]/NET0131 ,
		_w995_,
		_w1169_
	);
	LUT4 #(
		.INIT('hae00)
	) name241 (
		\data_o[91]_pad ,
		decrypt_i_pad,
		_w995_,
		_w1032_,
		_w1170_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name242 (
		_w1167_,
		_w1168_,
		_w1169_,
		_w1170_,
		_w1171_
	);
	LUT4 #(
		.INIT('h8000)
	) name243 (
		_w1166_,
		_w1171_,
		_w1156_,
		_w1161_,
		_w1172_
	);
	LUT3 #(
		.INIT('h02)
	) name244 (
		decrypt_i_pad,
		\mix1_data_o_reg_reg[27]/NET0131 ,
		_w995_,
		_w1173_
	);
	LUT4 #(
		.INIT('hae00)
	) name245 (
		\data_o[27]_pad ,
		decrypt_i_pad,
		_w995_,
		_w1020_,
		_w1174_
	);
	LUT2 #(
		.INIT('h4)
	) name246 (
		_w1173_,
		_w1174_,
		_w1175_
	);
	LUT3 #(
		.INIT('h02)
	) name247 (
		decrypt_i_pad,
		\mix1_data_o_reg_reg[59]/NET0131 ,
		_w995_,
		_w1176_
	);
	LUT4 #(
		.INIT('hae00)
	) name248 (
		\data_o[59]_pad ,
		decrypt_i_pad,
		_w995_,
		_w999_,
		_w1177_
	);
	LUT3 #(
		.INIT('h02)
	) name249 (
		decrypt_i_pad,
		\mix1_data_o_reg_reg[107]/NET0131 ,
		_w995_,
		_w1178_
	);
	LUT4 #(
		.INIT('hae00)
	) name250 (
		\data_o[107]_pad ,
		decrypt_i_pad,
		_w995_,
		_w1028_,
		_w1179_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name251 (
		_w1176_,
		_w1177_,
		_w1178_,
		_w1179_,
		_w1180_
	);
	LUT3 #(
		.INIT('h02)
	) name252 (
		decrypt_i_pad,
		\mix1_data_o_reg_reg[3]/NET0131 ,
		_w995_,
		_w1181_
	);
	LUT4 #(
		.INIT('hae00)
	) name253 (
		\data_o[3]_pad ,
		decrypt_i_pad,
		_w995_,
		_w1009_,
		_w1182_
	);
	LUT3 #(
		.INIT('h02)
	) name254 (
		decrypt_i_pad,
		\mix1_data_o_reg_reg[75]/NET0131 ,
		_w995_,
		_w1183_
	);
	LUT4 #(
		.INIT('hae00)
	) name255 (
		\data_o[75]_pad ,
		decrypt_i_pad,
		_w995_,
		_w1035_,
		_w1184_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name256 (
		_w1181_,
		_w1182_,
		_w1183_,
		_w1184_,
		_w1185_
	);
	LUT3 #(
		.INIT('h02)
	) name257 (
		decrypt_i_pad,
		\mix1_data_o_reg_reg[19]/NET0131 ,
		_w995_,
		_w1186_
	);
	LUT4 #(
		.INIT('hae00)
	) name258 (
		\data_o[19]_pad ,
		decrypt_i_pad,
		_w995_,
		_w1023_,
		_w1187_
	);
	LUT3 #(
		.INIT('h02)
	) name259 (
		decrypt_i_pad,
		\mix1_data_o_reg_reg[11]/NET0131 ,
		_w995_,
		_w1188_
	);
	LUT4 #(
		.INIT('ha0e0)
	) name260 (
		\data_o[11]_pad ,
		decrypt_i_pad,
		_w1013_,
		_w995_,
		_w1189_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name261 (
		_w1186_,
		_w1187_,
		_w1188_,
		_w1189_,
		_w1190_
	);
	LUT4 #(
		.INIT('h4000)
	) name262 (
		_w1175_,
		_w1185_,
		_w1190_,
		_w1180_,
		_w1191_
	);
	LUT3 #(
		.INIT('h51)
	) name263 (
		\data_o[123]_pad ,
		decrypt_i_pad,
		_w995_,
		_w1192_
	);
	LUT3 #(
		.INIT('h02)
	) name264 (
		decrypt_i_pad,
		\mix1_data_o_reg_reg[123]/NET0131 ,
		_w995_,
		_w1193_
	);
	LUT3 #(
		.INIT('h02)
	) name265 (
		_w1060_,
		_w1193_,
		_w1192_,
		_w1194_
	);
	LUT2 #(
		.INIT('h8)
	) name266 (
		_w1057_,
		_w1194_,
		_w1195_
	);
	LUT4 #(
		.INIT('h00ea)
	) name267 (
		_w1053_,
		_w1172_,
		_w1191_,
		_w1195_,
		_w1196_
	);
	LUT3 #(
		.INIT('hc8)
	) name268 (
		\addroundkey_start_i_reg/NET0131 ,
		\key_i[3]_pad ,
		_w936_,
		_w1197_
	);
	LUT3 #(
		.INIT('h02)
	) name269 (
		\ks1_key_reg_reg[3]/NET0131 ,
		_w936_,
		_w938_,
		_w1198_
	);
	LUT4 #(
		.INIT('h0001)
	) name270 (
		\addroundkey_round_reg[1]/NET0131 ,
		\addroundkey_round_reg[2]/NET0131 ,
		\addroundkey_round_reg[3]/NET0131 ,
		\key_i[3]_pad ,
		_w1199_
	);
	LUT4 #(
		.INIT('h00fe)
	) name271 (
		\addroundkey_round_reg[1]/NET0131 ,
		\addroundkey_round_reg[2]/NET0131 ,
		\addroundkey_round_reg[3]/NET0131 ,
		\ks1_key_reg_reg[3]/NET0131 ,
		_w1200_
	);
	LUT4 #(
		.INIT('h0008)
	) name272 (
		\addroundkey_start_i_reg/NET0131 ,
		_w930_,
		_w1200_,
		_w1199_,
		_w1201_
	);
	LUT4 #(
		.INIT('h00ab)
	) name273 (
		_w931_,
		_w1197_,
		_w1198_,
		_w1201_,
		_w1202_
	);
	LUT3 #(
		.INIT('hc8)
	) name274 (
		\addroundkey_start_i_reg/NET0131 ,
		\key_i[19]_pad ,
		_w936_,
		_w1203_
	);
	LUT3 #(
		.INIT('h02)
	) name275 (
		\ks1_key_reg_reg[19]/NET0131 ,
		_w936_,
		_w938_,
		_w1204_
	);
	LUT4 #(
		.INIT('h0001)
	) name276 (
		\addroundkey_round_reg[1]/NET0131 ,
		\addroundkey_round_reg[2]/NET0131 ,
		\addroundkey_round_reg[3]/NET0131 ,
		\key_i[19]_pad ,
		_w1205_
	);
	LUT4 #(
		.INIT('h00fe)
	) name277 (
		\addroundkey_round_reg[1]/NET0131 ,
		\addroundkey_round_reg[2]/NET0131 ,
		\addroundkey_round_reg[3]/NET0131 ,
		\ks1_key_reg_reg[19]/NET0131 ,
		_w1206_
	);
	LUT4 #(
		.INIT('h0008)
	) name278 (
		\addroundkey_start_i_reg/NET0131 ,
		_w930_,
		_w1206_,
		_w1205_,
		_w1207_
	);
	LUT4 #(
		.INIT('h00ab)
	) name279 (
		_w931_,
		_w1203_,
		_w1204_,
		_w1207_,
		_w1208_
	);
	LUT4 #(
		.INIT('hf531)
	) name280 (
		_w1064_,
		_w1079_,
		_w1202_,
		_w1208_,
		_w1209_
	);
	LUT3 #(
		.INIT('hc8)
	) name281 (
		\addroundkey_start_i_reg/NET0131 ,
		\key_i[11]_pad ,
		_w936_,
		_w1210_
	);
	LUT3 #(
		.INIT('h02)
	) name282 (
		\ks1_key_reg_reg[11]/NET0131 ,
		_w936_,
		_w938_,
		_w1211_
	);
	LUT4 #(
		.INIT('h0001)
	) name283 (
		\addroundkey_round_reg[1]/NET0131 ,
		\addroundkey_round_reg[2]/NET0131 ,
		\addroundkey_round_reg[3]/NET0131 ,
		\key_i[11]_pad ,
		_w1212_
	);
	LUT4 #(
		.INIT('h00fe)
	) name284 (
		\addroundkey_round_reg[1]/NET0131 ,
		\addroundkey_round_reg[2]/NET0131 ,
		\addroundkey_round_reg[3]/NET0131 ,
		\ks1_key_reg_reg[11]/NET0131 ,
		_w1213_
	);
	LUT4 #(
		.INIT('h0008)
	) name285 (
		\addroundkey_start_i_reg/NET0131 ,
		_w930_,
		_w1213_,
		_w1212_,
		_w1214_
	);
	LUT4 #(
		.INIT('h00ab)
	) name286 (
		_w931_,
		_w1210_,
		_w1211_,
		_w1214_,
		_w1215_
	);
	LUT3 #(
		.INIT('hc8)
	) name287 (
		\addroundkey_start_i_reg/NET0131 ,
		\key_i[27]_pad ,
		_w936_,
		_w1216_
	);
	LUT3 #(
		.INIT('h02)
	) name288 (
		\ks1_key_reg_reg[27]/NET0131 ,
		_w936_,
		_w938_,
		_w1217_
	);
	LUT4 #(
		.INIT('h0001)
	) name289 (
		\addroundkey_round_reg[1]/NET0131 ,
		\addroundkey_round_reg[2]/NET0131 ,
		\addroundkey_round_reg[3]/NET0131 ,
		\key_i[27]_pad ,
		_w1218_
	);
	LUT4 #(
		.INIT('h00fe)
	) name290 (
		\addroundkey_round_reg[1]/NET0131 ,
		\addroundkey_round_reg[2]/NET0131 ,
		\addroundkey_round_reg[3]/NET0131 ,
		\ks1_key_reg_reg[27]/NET0131 ,
		_w1219_
	);
	LUT4 #(
		.INIT('h0008)
	) name291 (
		\addroundkey_start_i_reg/NET0131 ,
		_w930_,
		_w1219_,
		_w1218_,
		_w1220_
	);
	LUT4 #(
		.INIT('h00ab)
	) name292 (
		_w931_,
		_w1216_,
		_w1217_,
		_w1220_,
		_w1221_
	);
	LUT4 #(
		.INIT('hf351)
	) name293 (
		_w948_,
		_w1071_,
		_w1215_,
		_w1221_,
		_w1222_
	);
	LUT4 #(
		.INIT('hd000)
	) name294 (
		_w950_,
		_w1196_,
		_w1209_,
		_w1222_,
		_w1223_
	);
	LUT3 #(
		.INIT('h02)
	) name295 (
		decrypt_i_pad,
		\mix1_data_o_reg_reg[9]/NET0131 ,
		_w995_,
		_w1224_
	);
	LUT4 #(
		.INIT('ha0e0)
	) name296 (
		\data_o[9]_pad ,
		decrypt_i_pad,
		_w1013_,
		_w995_,
		_w1225_
	);
	LUT3 #(
		.INIT('h02)
	) name297 (
		decrypt_i_pad,
		\mix1_data_o_reg_reg[57]/NET0131 ,
		_w995_,
		_w1226_
	);
	LUT4 #(
		.INIT('hae00)
	) name298 (
		\data_o[57]_pad ,
		decrypt_i_pad,
		_w995_,
		_w999_,
		_w1227_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name299 (
		_w1224_,
		_w1225_,
		_w1226_,
		_w1227_,
		_w1228_
	);
	LUT3 #(
		.INIT('h02)
	) name300 (
		decrypt_i_pad,
		\mix1_data_o_reg_reg[49]/NET0131 ,
		_w995_,
		_w1229_
	);
	LUT4 #(
		.INIT('hae00)
	) name301 (
		\data_o[49]_pad ,
		decrypt_i_pad,
		_w995_,
		_w1046_,
		_w1230_
	);
	LUT3 #(
		.INIT('h02)
	) name302 (
		decrypt_i_pad,
		\mix1_data_o_reg_reg[89]/NET0131 ,
		_w995_,
		_w1231_
	);
	LUT4 #(
		.INIT('hae00)
	) name303 (
		\data_o[89]_pad ,
		decrypt_i_pad,
		_w995_,
		_w1032_,
		_w1232_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name304 (
		_w1229_,
		_w1230_,
		_w1231_,
		_w1232_,
		_w1233_
	);
	LUT3 #(
		.INIT('h02)
	) name305 (
		decrypt_i_pad,
		\mix1_data_o_reg_reg[105]/NET0131 ,
		_w995_,
		_w1234_
	);
	LUT4 #(
		.INIT('hae00)
	) name306 (
		\data_o[105]_pad ,
		decrypt_i_pad,
		_w995_,
		_w1028_,
		_w1235_
	);
	LUT3 #(
		.INIT('h02)
	) name307 (
		decrypt_i_pad,
		\mix1_data_o_reg_reg[81]/NET0131 ,
		_w995_,
		_w1236_
	);
	LUT4 #(
		.INIT('hae00)
	) name308 (
		\data_o[81]_pad ,
		decrypt_i_pad,
		_w995_,
		_w1049_,
		_w1237_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name309 (
		_w1234_,
		_w1235_,
		_w1236_,
		_w1237_,
		_w1238_
	);
	LUT3 #(
		.INIT('h02)
	) name310 (
		decrypt_i_pad,
		\mix1_data_o_reg_reg[113]/NET0131 ,
		_w995_,
		_w1239_
	);
	LUT4 #(
		.INIT('hae00)
	) name311 (
		\data_o[113]_pad ,
		decrypt_i_pad,
		_w995_,
		_w1002_,
		_w1240_
	);
	LUT3 #(
		.INIT('h02)
	) name312 (
		decrypt_i_pad,
		\mix1_data_o_reg_reg[17]/NET0131 ,
		_w995_,
		_w1241_
	);
	LUT4 #(
		.INIT('hae00)
	) name313 (
		\data_o[17]_pad ,
		decrypt_i_pad,
		_w995_,
		_w1023_,
		_w1242_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name314 (
		_w1239_,
		_w1240_,
		_w1241_,
		_w1242_,
		_w1243_
	);
	LUT4 #(
		.INIT('h8000)
	) name315 (
		_w1238_,
		_w1243_,
		_w1228_,
		_w1233_,
		_w1244_
	);
	LUT3 #(
		.INIT('h02)
	) name316 (
		decrypt_i_pad,
		\mix1_data_o_reg_reg[97]/NET0131 ,
		_w995_,
		_w1245_
	);
	LUT4 #(
		.INIT('hae00)
	) name317 (
		\data_o[97]_pad ,
		decrypt_i_pad,
		_w995_,
		_w1016_,
		_w1246_
	);
	LUT2 #(
		.INIT('h4)
	) name318 (
		_w1245_,
		_w1246_,
		_w1247_
	);
	LUT3 #(
		.INIT('h02)
	) name319 (
		decrypt_i_pad,
		\mix1_data_o_reg_reg[73]/NET0131 ,
		_w995_,
		_w1248_
	);
	LUT4 #(
		.INIT('hae00)
	) name320 (
		\data_o[73]_pad ,
		decrypt_i_pad,
		_w995_,
		_w1035_,
		_w1249_
	);
	LUT3 #(
		.INIT('h02)
	) name321 (
		decrypt_i_pad,
		\mix1_data_o_reg_reg[1]/NET0131 ,
		_w995_,
		_w1250_
	);
	LUT4 #(
		.INIT('hae00)
	) name322 (
		\data_o[1]_pad ,
		decrypt_i_pad,
		_w995_,
		_w1009_,
		_w1251_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name323 (
		_w1248_,
		_w1249_,
		_w1250_,
		_w1251_,
		_w1252_
	);
	LUT3 #(
		.INIT('h02)
	) name324 (
		decrypt_i_pad,
		\mix1_data_o_reg_reg[41]/NET0131 ,
		_w995_,
		_w1253_
	);
	LUT4 #(
		.INIT('hae00)
	) name325 (
		\data_o[41]_pad ,
		decrypt_i_pad,
		_w995_,
		_w1006_,
		_w1254_
	);
	LUT3 #(
		.INIT('h02)
	) name326 (
		decrypt_i_pad,
		\mix1_data_o_reg_reg[25]/NET0131 ,
		_w995_,
		_w1255_
	);
	LUT4 #(
		.INIT('hae00)
	) name327 (
		\data_o[25]_pad ,
		decrypt_i_pad,
		_w995_,
		_w1020_,
		_w1256_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name328 (
		_w1253_,
		_w1254_,
		_w1255_,
		_w1256_,
		_w1257_
	);
	LUT3 #(
		.INIT('h02)
	) name329 (
		decrypt_i_pad,
		\mix1_data_o_reg_reg[65]/NET0131 ,
		_w995_,
		_w1258_
	);
	LUT4 #(
		.INIT('hae00)
	) name330 (
		\data_o[65]_pad ,
		decrypt_i_pad,
		_w995_,
		_w1039_,
		_w1259_
	);
	LUT3 #(
		.INIT('h02)
	) name331 (
		decrypt_i_pad,
		\mix1_data_o_reg_reg[33]/NET0131 ,
		_w995_,
		_w1260_
	);
	LUT4 #(
		.INIT('hae00)
	) name332 (
		\data_o[33]_pad ,
		decrypt_i_pad,
		_w995_,
		_w1042_,
		_w1261_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name333 (
		_w1258_,
		_w1259_,
		_w1260_,
		_w1261_,
		_w1262_
	);
	LUT4 #(
		.INIT('h4000)
	) name334 (
		_w1247_,
		_w1257_,
		_w1262_,
		_w1252_,
		_w1263_
	);
	LUT3 #(
		.INIT('h51)
	) name335 (
		\data_o[121]_pad ,
		decrypt_i_pad,
		_w995_,
		_w1264_
	);
	LUT3 #(
		.INIT('h02)
	) name336 (
		decrypt_i_pad,
		\mix1_data_o_reg_reg[121]/NET0131 ,
		_w995_,
		_w1265_
	);
	LUT3 #(
		.INIT('h02)
	) name337 (
		_w1060_,
		_w1265_,
		_w1264_,
		_w1266_
	);
	LUT2 #(
		.INIT('h8)
	) name338 (
		_w1057_,
		_w1266_,
		_w1267_
	);
	LUT4 #(
		.INIT('h00ea)
	) name339 (
		_w1053_,
		_w1244_,
		_w1263_,
		_w1267_,
		_w1268_
	);
	LUT3 #(
		.INIT('hc8)
	) name340 (
		\addroundkey_start_i_reg/NET0131 ,
		\key_i[9]_pad ,
		_w936_,
		_w1269_
	);
	LUT3 #(
		.INIT('h02)
	) name341 (
		\ks1_key_reg_reg[9]/NET0131 ,
		_w936_,
		_w938_,
		_w1270_
	);
	LUT4 #(
		.INIT('h0001)
	) name342 (
		\addroundkey_round_reg[1]/NET0131 ,
		\addroundkey_round_reg[2]/NET0131 ,
		\addroundkey_round_reg[3]/NET0131 ,
		\key_i[9]_pad ,
		_w1271_
	);
	LUT4 #(
		.INIT('h00fe)
	) name343 (
		\addroundkey_round_reg[1]/NET0131 ,
		\addroundkey_round_reg[2]/NET0131 ,
		\addroundkey_round_reg[3]/NET0131 ,
		\ks1_key_reg_reg[9]/NET0131 ,
		_w1272_
	);
	LUT4 #(
		.INIT('h0008)
	) name344 (
		\addroundkey_start_i_reg/NET0131 ,
		_w930_,
		_w1272_,
		_w1271_,
		_w1273_
	);
	LUT4 #(
		.INIT('h00ab)
	) name345 (
		_w931_,
		_w1269_,
		_w1270_,
		_w1273_,
		_w1274_
	);
	LUT3 #(
		.INIT('hc8)
	) name346 (
		\addroundkey_start_i_reg/NET0131 ,
		\key_i[17]_pad ,
		_w936_,
		_w1275_
	);
	LUT3 #(
		.INIT('h02)
	) name347 (
		\ks1_key_reg_reg[17]/NET0131 ,
		_w936_,
		_w938_,
		_w1276_
	);
	LUT4 #(
		.INIT('h0001)
	) name348 (
		\addroundkey_round_reg[1]/NET0131 ,
		\addroundkey_round_reg[2]/NET0131 ,
		\addroundkey_round_reg[3]/NET0131 ,
		\key_i[17]_pad ,
		_w1277_
	);
	LUT4 #(
		.INIT('h00fe)
	) name349 (
		\addroundkey_round_reg[1]/NET0131 ,
		\addroundkey_round_reg[2]/NET0131 ,
		\addroundkey_round_reg[3]/NET0131 ,
		\ks1_key_reg_reg[17]/NET0131 ,
		_w1278_
	);
	LUT4 #(
		.INIT('h0008)
	) name350 (
		\addroundkey_start_i_reg/NET0131 ,
		_w930_,
		_w1278_,
		_w1277_,
		_w1279_
	);
	LUT4 #(
		.INIT('h00ab)
	) name351 (
		_w931_,
		_w1275_,
		_w1276_,
		_w1279_,
		_w1280_
	);
	LUT4 #(
		.INIT('hf531)
	) name352 (
		_w1071_,
		_w1079_,
		_w1274_,
		_w1280_,
		_w1281_
	);
	LUT3 #(
		.INIT('hc8)
	) name353 (
		\addroundkey_start_i_reg/NET0131 ,
		\key_i[25]_pad ,
		_w936_,
		_w1282_
	);
	LUT3 #(
		.INIT('h02)
	) name354 (
		\ks1_key_reg_reg[25]/NET0131 ,
		_w936_,
		_w938_,
		_w1283_
	);
	LUT4 #(
		.INIT('h0001)
	) name355 (
		\addroundkey_round_reg[1]/NET0131 ,
		\addroundkey_round_reg[2]/NET0131 ,
		\addroundkey_round_reg[3]/NET0131 ,
		\key_i[25]_pad ,
		_w1284_
	);
	LUT4 #(
		.INIT('h00fe)
	) name356 (
		\addroundkey_round_reg[1]/NET0131 ,
		\addroundkey_round_reg[2]/NET0131 ,
		\addroundkey_round_reg[3]/NET0131 ,
		\ks1_key_reg_reg[25]/NET0131 ,
		_w1285_
	);
	LUT4 #(
		.INIT('h0008)
	) name357 (
		\addroundkey_start_i_reg/NET0131 ,
		_w930_,
		_w1285_,
		_w1284_,
		_w1286_
	);
	LUT4 #(
		.INIT('h00ab)
	) name358 (
		_w931_,
		_w1282_,
		_w1283_,
		_w1286_,
		_w1287_
	);
	LUT3 #(
		.INIT('hc8)
	) name359 (
		\addroundkey_start_i_reg/NET0131 ,
		\key_i[1]_pad ,
		_w936_,
		_w1288_
	);
	LUT3 #(
		.INIT('h02)
	) name360 (
		\ks1_key_reg_reg[1]/NET0131 ,
		_w936_,
		_w938_,
		_w1289_
	);
	LUT4 #(
		.INIT('h0001)
	) name361 (
		\addroundkey_round_reg[1]/NET0131 ,
		\addroundkey_round_reg[2]/NET0131 ,
		\addroundkey_round_reg[3]/NET0131 ,
		\key_i[1]_pad ,
		_w1290_
	);
	LUT4 #(
		.INIT('h00fe)
	) name362 (
		\addroundkey_round_reg[1]/NET0131 ,
		\addroundkey_round_reg[2]/NET0131 ,
		\addroundkey_round_reg[3]/NET0131 ,
		\ks1_key_reg_reg[1]/NET0131 ,
		_w1291_
	);
	LUT4 #(
		.INIT('h0008)
	) name363 (
		\addroundkey_start_i_reg/NET0131 ,
		_w930_,
		_w1291_,
		_w1290_,
		_w1292_
	);
	LUT4 #(
		.INIT('h00ab)
	) name364 (
		_w931_,
		_w1288_,
		_w1289_,
		_w1292_,
		_w1293_
	);
	LUT4 #(
		.INIT('hf531)
	) name365 (
		_w948_,
		_w1064_,
		_w1287_,
		_w1293_,
		_w1294_
	);
	LUT4 #(
		.INIT('hd000)
	) name366 (
		_w950_,
		_w1268_,
		_w1281_,
		_w1294_,
		_w1295_
	);
	LUT4 #(
		.INIT('h2882)
	) name367 (
		_w951_,
		_w1151_,
		_w1223_,
		_w1295_,
		_w1296_
	);
	LUT2 #(
		.INIT('h1)
	) name368 (
		_w1094_,
		_w1296_,
		_w1297_
	);
	LUT3 #(
		.INIT('h02)
	) name369 (
		decrypt_i_pad,
		\mix1_data_o_reg_reg[72]/NET0131 ,
		_w995_,
		_w1298_
	);
	LUT4 #(
		.INIT('hae00)
	) name370 (
		\data_o[72]_pad ,
		decrypt_i_pad,
		_w995_,
		_w1035_,
		_w1299_
	);
	LUT3 #(
		.INIT('h02)
	) name371 (
		decrypt_i_pad,
		\mix1_data_o_reg_reg[56]/NET0131 ,
		_w995_,
		_w1300_
	);
	LUT4 #(
		.INIT('hae00)
	) name372 (
		\data_o[56]_pad ,
		decrypt_i_pad,
		_w995_,
		_w999_,
		_w1301_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name373 (
		_w1298_,
		_w1299_,
		_w1300_,
		_w1301_,
		_w1302_
	);
	LUT3 #(
		.INIT('h02)
	) name374 (
		decrypt_i_pad,
		\mix1_data_o_reg_reg[88]/NET0131 ,
		_w995_,
		_w1303_
	);
	LUT4 #(
		.INIT('hae00)
	) name375 (
		\data_o[88]_pad ,
		decrypt_i_pad,
		_w995_,
		_w1032_,
		_w1304_
	);
	LUT3 #(
		.INIT('h02)
	) name376 (
		decrypt_i_pad,
		\mix1_data_o_reg_reg[40]/NET0131 ,
		_w995_,
		_w1305_
	);
	LUT4 #(
		.INIT('hae00)
	) name377 (
		\data_o[40]_pad ,
		decrypt_i_pad,
		_w995_,
		_w1006_,
		_w1306_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name378 (
		_w1303_,
		_w1304_,
		_w1305_,
		_w1306_,
		_w1307_
	);
	LUT3 #(
		.INIT('h02)
	) name379 (
		decrypt_i_pad,
		\mix1_data_o_reg_reg[112]/NET0131 ,
		_w995_,
		_w1308_
	);
	LUT4 #(
		.INIT('hae00)
	) name380 (
		\data_o[112]_pad ,
		decrypt_i_pad,
		_w995_,
		_w1002_,
		_w1309_
	);
	LUT3 #(
		.INIT('h02)
	) name381 (
		decrypt_i_pad,
		\mix1_data_o_reg_reg[96]/NET0131 ,
		_w995_,
		_w1310_
	);
	LUT4 #(
		.INIT('hae00)
	) name382 (
		\data_o[96]_pad ,
		decrypt_i_pad,
		_w995_,
		_w1016_,
		_w1311_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name383 (
		_w1308_,
		_w1309_,
		_w1310_,
		_w1311_,
		_w1312_
	);
	LUT3 #(
		.INIT('h02)
	) name384 (
		decrypt_i_pad,
		\mix1_data_o_reg_reg[104]/NET0131 ,
		_w995_,
		_w1313_
	);
	LUT4 #(
		.INIT('hae00)
	) name385 (
		\data_o[104]_pad ,
		decrypt_i_pad,
		_w995_,
		_w1028_,
		_w1314_
	);
	LUT3 #(
		.INIT('h02)
	) name386 (
		decrypt_i_pad,
		\mix1_data_o_reg_reg[64]/NET0131 ,
		_w995_,
		_w1315_
	);
	LUT4 #(
		.INIT('hae00)
	) name387 (
		\data_o[64]_pad ,
		decrypt_i_pad,
		_w995_,
		_w1039_,
		_w1316_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name388 (
		_w1313_,
		_w1314_,
		_w1315_,
		_w1316_,
		_w1317_
	);
	LUT4 #(
		.INIT('h8000)
	) name389 (
		_w1312_,
		_w1317_,
		_w1302_,
		_w1307_,
		_w1318_
	);
	LUT3 #(
		.INIT('h02)
	) name390 (
		decrypt_i_pad,
		\mix1_data_o_reg_reg[80]/NET0131 ,
		_w995_,
		_w1319_
	);
	LUT4 #(
		.INIT('hae00)
	) name391 (
		\data_o[80]_pad ,
		decrypt_i_pad,
		_w995_,
		_w1049_,
		_w1320_
	);
	LUT2 #(
		.INIT('h4)
	) name392 (
		_w1319_,
		_w1320_,
		_w1321_
	);
	LUT3 #(
		.INIT('h02)
	) name393 (
		decrypt_i_pad,
		\mix1_data_o_reg_reg[8]/NET0131 ,
		_w995_,
		_w1322_
	);
	LUT4 #(
		.INIT('ha0e0)
	) name394 (
		\data_o[8]_pad ,
		decrypt_i_pad,
		_w1013_,
		_w995_,
		_w1323_
	);
	LUT3 #(
		.INIT('h02)
	) name395 (
		decrypt_i_pad,
		\mix1_data_o_reg_reg[32]/NET0131 ,
		_w995_,
		_w1324_
	);
	LUT4 #(
		.INIT('hae00)
	) name396 (
		\data_o[32]_pad ,
		decrypt_i_pad,
		_w995_,
		_w1042_,
		_w1325_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name397 (
		_w1322_,
		_w1323_,
		_w1324_,
		_w1325_,
		_w1326_
	);
	LUT3 #(
		.INIT('h02)
	) name398 (
		decrypt_i_pad,
		\mix1_data_o_reg_reg[48]/NET0131 ,
		_w995_,
		_w1327_
	);
	LUT4 #(
		.INIT('hae00)
	) name399 (
		\data_o[48]_pad ,
		decrypt_i_pad,
		_w995_,
		_w1046_,
		_w1328_
	);
	LUT3 #(
		.INIT('h02)
	) name400 (
		decrypt_i_pad,
		\mix1_data_o_reg_reg[0]/NET0131 ,
		_w995_,
		_w1329_
	);
	LUT4 #(
		.INIT('hae00)
	) name401 (
		\data_o[0]_pad ,
		decrypt_i_pad,
		_w995_,
		_w1009_,
		_w1330_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name402 (
		_w1327_,
		_w1328_,
		_w1329_,
		_w1330_,
		_w1331_
	);
	LUT3 #(
		.INIT('h02)
	) name403 (
		decrypt_i_pad,
		\mix1_data_o_reg_reg[16]/NET0131 ,
		_w995_,
		_w1332_
	);
	LUT4 #(
		.INIT('hae00)
	) name404 (
		\data_o[16]_pad ,
		decrypt_i_pad,
		_w995_,
		_w1023_,
		_w1333_
	);
	LUT3 #(
		.INIT('h02)
	) name405 (
		decrypt_i_pad,
		\mix1_data_o_reg_reg[24]/NET0131 ,
		_w995_,
		_w1334_
	);
	LUT4 #(
		.INIT('hae00)
	) name406 (
		\data_o[24]_pad ,
		decrypt_i_pad,
		_w995_,
		_w1020_,
		_w1335_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name407 (
		_w1332_,
		_w1333_,
		_w1334_,
		_w1335_,
		_w1336_
	);
	LUT4 #(
		.INIT('h4000)
	) name408 (
		_w1321_,
		_w1331_,
		_w1336_,
		_w1326_,
		_w1337_
	);
	LUT3 #(
		.INIT('h51)
	) name409 (
		\data_o[120]_pad ,
		decrypt_i_pad,
		_w995_,
		_w1338_
	);
	LUT3 #(
		.INIT('h02)
	) name410 (
		decrypt_i_pad,
		\mix1_data_o_reg_reg[120]/NET0131 ,
		_w995_,
		_w1339_
	);
	LUT3 #(
		.INIT('h02)
	) name411 (
		_w1060_,
		_w1339_,
		_w1338_,
		_w1340_
	);
	LUT2 #(
		.INIT('h8)
	) name412 (
		_w1057_,
		_w1340_,
		_w1341_
	);
	LUT4 #(
		.INIT('h00ea)
	) name413 (
		_w1053_,
		_w1318_,
		_w1337_,
		_w1341_,
		_w1342_
	);
	LUT4 #(
		.INIT('h5553)
	) name414 (
		\key_i[16]_pad ,
		\ks1_key_reg_reg[16]/NET0131 ,
		_w938_,
		_w986_,
		_w1343_
	);
	LUT2 #(
		.INIT('h2)
	) name415 (
		_w1079_,
		_w1343_,
		_w1344_
	);
	LUT3 #(
		.INIT('hc8)
	) name416 (
		\addroundkey_start_i_reg/NET0131 ,
		\key_i[8]_pad ,
		_w936_,
		_w1345_
	);
	LUT3 #(
		.INIT('h02)
	) name417 (
		\ks1_key_reg_reg[8]/NET0131 ,
		_w936_,
		_w938_,
		_w1346_
	);
	LUT4 #(
		.INIT('h0001)
	) name418 (
		\addroundkey_round_reg[1]/NET0131 ,
		\addroundkey_round_reg[2]/NET0131 ,
		\addroundkey_round_reg[3]/NET0131 ,
		\key_i[8]_pad ,
		_w1347_
	);
	LUT4 #(
		.INIT('h00fe)
	) name419 (
		\addroundkey_round_reg[1]/NET0131 ,
		\addroundkey_round_reg[2]/NET0131 ,
		\addroundkey_round_reg[3]/NET0131 ,
		\ks1_key_reg_reg[8]/NET0131 ,
		_w1348_
	);
	LUT4 #(
		.INIT('h0008)
	) name420 (
		\addroundkey_start_i_reg/NET0131 ,
		_w930_,
		_w1348_,
		_w1347_,
		_w1349_
	);
	LUT4 #(
		.INIT('h00ab)
	) name421 (
		_w931_,
		_w1345_,
		_w1346_,
		_w1349_,
		_w1350_
	);
	LUT3 #(
		.INIT('h31)
	) name422 (
		_w1071_,
		_w1344_,
		_w1350_,
		_w1351_
	);
	LUT3 #(
		.INIT('hc8)
	) name423 (
		\addroundkey_start_i_reg/NET0131 ,
		\key_i[24]_pad ,
		_w936_,
		_w1352_
	);
	LUT3 #(
		.INIT('h02)
	) name424 (
		\ks1_key_reg_reg[24]/NET0131 ,
		_w936_,
		_w938_,
		_w1353_
	);
	LUT4 #(
		.INIT('h0001)
	) name425 (
		\addroundkey_round_reg[1]/NET0131 ,
		\addroundkey_round_reg[2]/NET0131 ,
		\addroundkey_round_reg[3]/NET0131 ,
		\key_i[24]_pad ,
		_w1354_
	);
	LUT4 #(
		.INIT('h00fe)
	) name426 (
		\addroundkey_round_reg[1]/NET0131 ,
		\addroundkey_round_reg[2]/NET0131 ,
		\addroundkey_round_reg[3]/NET0131 ,
		\ks1_key_reg_reg[24]/NET0131 ,
		_w1355_
	);
	LUT4 #(
		.INIT('h0008)
	) name427 (
		\addroundkey_start_i_reg/NET0131 ,
		_w930_,
		_w1355_,
		_w1354_,
		_w1356_
	);
	LUT4 #(
		.INIT('h00ab)
	) name428 (
		_w931_,
		_w1352_,
		_w1353_,
		_w1356_,
		_w1357_
	);
	LUT3 #(
		.INIT('hc8)
	) name429 (
		\addroundkey_start_i_reg/NET0131 ,
		\key_i[0]_pad ,
		_w936_,
		_w1358_
	);
	LUT3 #(
		.INIT('h02)
	) name430 (
		\ks1_key_reg_reg[0]/NET0131 ,
		_w936_,
		_w938_,
		_w1359_
	);
	LUT4 #(
		.INIT('h0001)
	) name431 (
		\addroundkey_round_reg[1]/NET0131 ,
		\addroundkey_round_reg[2]/NET0131 ,
		\addroundkey_round_reg[3]/NET0131 ,
		\key_i[0]_pad ,
		_w1360_
	);
	LUT4 #(
		.INIT('h00fe)
	) name432 (
		\addroundkey_round_reg[1]/NET0131 ,
		\addroundkey_round_reg[2]/NET0131 ,
		\addroundkey_round_reg[3]/NET0131 ,
		\ks1_key_reg_reg[0]/NET0131 ,
		_w1361_
	);
	LUT4 #(
		.INIT('h0008)
	) name433 (
		\addroundkey_start_i_reg/NET0131 ,
		_w930_,
		_w1361_,
		_w1360_,
		_w1362_
	);
	LUT4 #(
		.INIT('h00ab)
	) name434 (
		_w931_,
		_w1358_,
		_w1359_,
		_w1362_,
		_w1363_
	);
	LUT4 #(
		.INIT('hf531)
	) name435 (
		_w948_,
		_w1064_,
		_w1357_,
		_w1363_,
		_w1364_
	);
	LUT4 #(
		.INIT('hd000)
	) name436 (
		_w950_,
		_w1342_,
		_w1351_,
		_w1364_,
		_w1365_
	);
	LUT3 #(
		.INIT('h02)
	) name437 (
		decrypt_i_pad,
		\mix1_data_o_reg_reg[21]/NET0131 ,
		_w995_,
		_w1366_
	);
	LUT4 #(
		.INIT('hae00)
	) name438 (
		\data_o[21]_pad ,
		decrypt_i_pad,
		_w995_,
		_w1023_,
		_w1367_
	);
	LUT3 #(
		.INIT('h02)
	) name439 (
		decrypt_i_pad,
		\mix1_data_o_reg_reg[13]/NET0131 ,
		_w995_,
		_w1368_
	);
	LUT4 #(
		.INIT('ha0e0)
	) name440 (
		\data_o[13]_pad ,
		decrypt_i_pad,
		_w1013_,
		_w995_,
		_w1369_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name441 (
		_w1366_,
		_w1367_,
		_w1368_,
		_w1369_,
		_w1370_
	);
	LUT3 #(
		.INIT('h02)
	) name442 (
		decrypt_i_pad,
		\mix1_data_o_reg_reg[5]/NET0131 ,
		_w995_,
		_w1371_
	);
	LUT4 #(
		.INIT('hae00)
	) name443 (
		\data_o[5]_pad ,
		decrypt_i_pad,
		_w995_,
		_w1009_,
		_w1372_
	);
	LUT3 #(
		.INIT('h02)
	) name444 (
		decrypt_i_pad,
		\mix1_data_o_reg_reg[53]/NET0131 ,
		_w995_,
		_w1373_
	);
	LUT4 #(
		.INIT('hae00)
	) name445 (
		\data_o[53]_pad ,
		decrypt_i_pad,
		_w995_,
		_w1046_,
		_w1374_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name446 (
		_w1371_,
		_w1372_,
		_w1373_,
		_w1374_,
		_w1375_
	);
	LUT3 #(
		.INIT('h02)
	) name447 (
		decrypt_i_pad,
		\mix1_data_o_reg_reg[61]/NET0131 ,
		_w995_,
		_w1376_
	);
	LUT4 #(
		.INIT('hae00)
	) name448 (
		\data_o[61]_pad ,
		decrypt_i_pad,
		_w995_,
		_w999_,
		_w1377_
	);
	LUT3 #(
		.INIT('h02)
	) name449 (
		decrypt_i_pad,
		\mix1_data_o_reg_reg[29]/NET0131 ,
		_w995_,
		_w1378_
	);
	LUT4 #(
		.INIT('hae00)
	) name450 (
		\data_o[29]_pad ,
		decrypt_i_pad,
		_w995_,
		_w1020_,
		_w1379_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name451 (
		_w1376_,
		_w1377_,
		_w1378_,
		_w1379_,
		_w1380_
	);
	LUT3 #(
		.INIT('h02)
	) name452 (
		decrypt_i_pad,
		\mix1_data_o_reg_reg[85]/NET0131 ,
		_w995_,
		_w1381_
	);
	LUT4 #(
		.INIT('hae00)
	) name453 (
		\data_o[85]_pad ,
		decrypt_i_pad,
		_w995_,
		_w1049_,
		_w1382_
	);
	LUT3 #(
		.INIT('h02)
	) name454 (
		decrypt_i_pad,
		\mix1_data_o_reg_reg[69]/NET0131 ,
		_w995_,
		_w1383_
	);
	LUT4 #(
		.INIT('hae00)
	) name455 (
		\data_o[69]_pad ,
		decrypt_i_pad,
		_w995_,
		_w1039_,
		_w1384_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name456 (
		_w1381_,
		_w1382_,
		_w1383_,
		_w1384_,
		_w1385_
	);
	LUT4 #(
		.INIT('h8000)
	) name457 (
		_w1380_,
		_w1385_,
		_w1370_,
		_w1375_,
		_w1386_
	);
	LUT3 #(
		.INIT('h02)
	) name458 (
		decrypt_i_pad,
		\mix1_data_o_reg_reg[109]/NET0131 ,
		_w995_,
		_w1387_
	);
	LUT4 #(
		.INIT('hae00)
	) name459 (
		\data_o[109]_pad ,
		decrypt_i_pad,
		_w995_,
		_w1028_,
		_w1388_
	);
	LUT2 #(
		.INIT('h4)
	) name460 (
		_w1387_,
		_w1388_,
		_w1389_
	);
	LUT3 #(
		.INIT('h02)
	) name461 (
		decrypt_i_pad,
		\mix1_data_o_reg_reg[117]/NET0131 ,
		_w995_,
		_w1390_
	);
	LUT4 #(
		.INIT('hae00)
	) name462 (
		\data_o[117]_pad ,
		decrypt_i_pad,
		_w995_,
		_w1002_,
		_w1391_
	);
	LUT3 #(
		.INIT('h02)
	) name463 (
		decrypt_i_pad,
		\mix1_data_o_reg_reg[37]/NET0131 ,
		_w995_,
		_w1392_
	);
	LUT4 #(
		.INIT('hae00)
	) name464 (
		\data_o[37]_pad ,
		decrypt_i_pad,
		_w995_,
		_w1042_,
		_w1393_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name465 (
		_w1390_,
		_w1391_,
		_w1392_,
		_w1393_,
		_w1394_
	);
	LUT3 #(
		.INIT('h02)
	) name466 (
		decrypt_i_pad,
		\mix1_data_o_reg_reg[45]/NET0131 ,
		_w995_,
		_w1395_
	);
	LUT4 #(
		.INIT('hae00)
	) name467 (
		\data_o[45]_pad ,
		decrypt_i_pad,
		_w995_,
		_w1006_,
		_w1396_
	);
	LUT3 #(
		.INIT('h02)
	) name468 (
		decrypt_i_pad,
		\mix1_data_o_reg_reg[93]/NET0131 ,
		_w995_,
		_w1397_
	);
	LUT4 #(
		.INIT('hae00)
	) name469 (
		\data_o[93]_pad ,
		decrypt_i_pad,
		_w995_,
		_w1032_,
		_w1398_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name470 (
		_w1395_,
		_w1396_,
		_w1397_,
		_w1398_,
		_w1399_
	);
	LUT3 #(
		.INIT('h02)
	) name471 (
		decrypt_i_pad,
		\mix1_data_o_reg_reg[77]/NET0131 ,
		_w995_,
		_w1400_
	);
	LUT4 #(
		.INIT('hae00)
	) name472 (
		\data_o[77]_pad ,
		decrypt_i_pad,
		_w995_,
		_w1035_,
		_w1401_
	);
	LUT3 #(
		.INIT('h02)
	) name473 (
		decrypt_i_pad,
		\mix1_data_o_reg_reg[101]/NET0131 ,
		_w995_,
		_w1402_
	);
	LUT4 #(
		.INIT('hae00)
	) name474 (
		\data_o[101]_pad ,
		decrypt_i_pad,
		_w995_,
		_w1016_,
		_w1403_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name475 (
		_w1400_,
		_w1401_,
		_w1402_,
		_w1403_,
		_w1404_
	);
	LUT4 #(
		.INIT('h4000)
	) name476 (
		_w1389_,
		_w1399_,
		_w1404_,
		_w1394_,
		_w1405_
	);
	LUT3 #(
		.INIT('h51)
	) name477 (
		\data_o[125]_pad ,
		decrypt_i_pad,
		_w995_,
		_w1406_
	);
	LUT3 #(
		.INIT('h02)
	) name478 (
		decrypt_i_pad,
		\mix1_data_o_reg_reg[125]/NET0131 ,
		_w995_,
		_w1407_
	);
	LUT3 #(
		.INIT('h02)
	) name479 (
		_w1060_,
		_w1407_,
		_w1406_,
		_w1408_
	);
	LUT2 #(
		.INIT('h8)
	) name480 (
		_w1057_,
		_w1408_,
		_w1409_
	);
	LUT4 #(
		.INIT('h00ea)
	) name481 (
		_w1053_,
		_w1386_,
		_w1405_,
		_w1409_,
		_w1410_
	);
	LUT4 #(
		.INIT('h5553)
	) name482 (
		\key_i[5]_pad ,
		\ks1_key_reg_reg[5]/NET0131 ,
		_w938_,
		_w986_,
		_w1411_
	);
	LUT2 #(
		.INIT('h2)
	) name483 (
		_w1064_,
		_w1411_,
		_w1412_
	);
	LUT3 #(
		.INIT('hc8)
	) name484 (
		\addroundkey_start_i_reg/NET0131 ,
		\key_i[21]_pad ,
		_w936_,
		_w1413_
	);
	LUT3 #(
		.INIT('h02)
	) name485 (
		\ks1_key_reg_reg[21]/NET0131 ,
		_w936_,
		_w938_,
		_w1414_
	);
	LUT4 #(
		.INIT('h0001)
	) name486 (
		\addroundkey_round_reg[1]/NET0131 ,
		\addroundkey_round_reg[2]/NET0131 ,
		\addroundkey_round_reg[3]/NET0131 ,
		\key_i[21]_pad ,
		_w1415_
	);
	LUT4 #(
		.INIT('h00fe)
	) name487 (
		\addroundkey_round_reg[1]/NET0131 ,
		\addroundkey_round_reg[2]/NET0131 ,
		\addroundkey_round_reg[3]/NET0131 ,
		\ks1_key_reg_reg[21]/NET0131 ,
		_w1416_
	);
	LUT4 #(
		.INIT('h0008)
	) name488 (
		\addroundkey_start_i_reg/NET0131 ,
		_w930_,
		_w1416_,
		_w1415_,
		_w1417_
	);
	LUT4 #(
		.INIT('h00ab)
	) name489 (
		_w931_,
		_w1413_,
		_w1414_,
		_w1417_,
		_w1418_
	);
	LUT3 #(
		.INIT('h31)
	) name490 (
		_w1079_,
		_w1412_,
		_w1418_,
		_w1419_
	);
	LUT3 #(
		.INIT('hc8)
	) name491 (
		\addroundkey_start_i_reg/NET0131 ,
		\key_i[29]_pad ,
		_w936_,
		_w1420_
	);
	LUT3 #(
		.INIT('h02)
	) name492 (
		\ks1_key_reg_reg[29]/NET0131 ,
		_w936_,
		_w938_,
		_w1421_
	);
	LUT4 #(
		.INIT('h0001)
	) name493 (
		\addroundkey_round_reg[1]/NET0131 ,
		\addroundkey_round_reg[2]/NET0131 ,
		\addroundkey_round_reg[3]/NET0131 ,
		\key_i[29]_pad ,
		_w1422_
	);
	LUT4 #(
		.INIT('h00fe)
	) name494 (
		\addroundkey_round_reg[1]/NET0131 ,
		\addroundkey_round_reg[2]/NET0131 ,
		\addroundkey_round_reg[3]/NET0131 ,
		\ks1_key_reg_reg[29]/NET0131 ,
		_w1423_
	);
	LUT4 #(
		.INIT('h0008)
	) name495 (
		\addroundkey_start_i_reg/NET0131 ,
		_w930_,
		_w1423_,
		_w1422_,
		_w1424_
	);
	LUT4 #(
		.INIT('h00ab)
	) name496 (
		_w931_,
		_w1420_,
		_w1421_,
		_w1424_,
		_w1425_
	);
	LUT3 #(
		.INIT('hc8)
	) name497 (
		\addroundkey_start_i_reg/NET0131 ,
		\key_i[13]_pad ,
		_w936_,
		_w1426_
	);
	LUT3 #(
		.INIT('h02)
	) name498 (
		\ks1_key_reg_reg[13]/NET0131 ,
		_w936_,
		_w938_,
		_w1427_
	);
	LUT4 #(
		.INIT('h0001)
	) name499 (
		\addroundkey_round_reg[1]/NET0131 ,
		\addroundkey_round_reg[2]/NET0131 ,
		\addroundkey_round_reg[3]/NET0131 ,
		\key_i[13]_pad ,
		_w1428_
	);
	LUT4 #(
		.INIT('h00fe)
	) name500 (
		\addroundkey_round_reg[1]/NET0131 ,
		\addroundkey_round_reg[2]/NET0131 ,
		\addroundkey_round_reg[3]/NET0131 ,
		\ks1_key_reg_reg[13]/NET0131 ,
		_w1429_
	);
	LUT4 #(
		.INIT('h0008)
	) name501 (
		\addroundkey_start_i_reg/NET0131 ,
		_w930_,
		_w1429_,
		_w1428_,
		_w1430_
	);
	LUT4 #(
		.INIT('h00ab)
	) name502 (
		_w931_,
		_w1426_,
		_w1427_,
		_w1430_,
		_w1431_
	);
	LUT4 #(
		.INIT('hf531)
	) name503 (
		_w948_,
		_w1071_,
		_w1425_,
		_w1431_,
		_w1432_
	);
	LUT4 #(
		.INIT('hd000)
	) name504 (
		_w950_,
		_w1410_,
		_w1419_,
		_w1432_,
		_w1433_
	);
	LUT4 #(
		.INIT('h2882)
	) name505 (
		_w951_,
		_w1223_,
		_w1365_,
		_w1433_,
		_w1434_
	);
	LUT2 #(
		.INIT('h1)
	) name506 (
		_w951_,
		_w1151_,
		_w1435_
	);
	LUT4 #(
		.INIT('heee1)
	) name507 (
		_w1094_,
		_w1296_,
		_w1434_,
		_w1435_,
		_w1436_
	);
	LUT3 #(
		.INIT('h02)
	) name508 (
		decrypt_i_pad,
		\mix1_data_o_reg_reg[58]/NET0131 ,
		_w995_,
		_w1437_
	);
	LUT4 #(
		.INIT('hae00)
	) name509 (
		\data_o[58]_pad ,
		decrypt_i_pad,
		_w995_,
		_w999_,
		_w1438_
	);
	LUT3 #(
		.INIT('h02)
	) name510 (
		decrypt_i_pad,
		\mix1_data_o_reg_reg[98]/NET0131 ,
		_w995_,
		_w1439_
	);
	LUT4 #(
		.INIT('hae00)
	) name511 (
		\data_o[98]_pad ,
		decrypt_i_pad,
		_w995_,
		_w1016_,
		_w1440_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name512 (
		_w1437_,
		_w1438_,
		_w1439_,
		_w1440_,
		_w1441_
	);
	LUT3 #(
		.INIT('h02)
	) name513 (
		decrypt_i_pad,
		\mix1_data_o_reg_reg[50]/NET0131 ,
		_w995_,
		_w1442_
	);
	LUT4 #(
		.INIT('hae00)
	) name514 (
		\data_o[50]_pad ,
		decrypt_i_pad,
		_w995_,
		_w1046_,
		_w1443_
	);
	LUT3 #(
		.INIT('h02)
	) name515 (
		decrypt_i_pad,
		\mix1_data_o_reg_reg[90]/NET0131 ,
		_w995_,
		_w1444_
	);
	LUT4 #(
		.INIT('hae00)
	) name516 (
		\data_o[90]_pad ,
		decrypt_i_pad,
		_w995_,
		_w1032_,
		_w1445_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name517 (
		_w1442_,
		_w1443_,
		_w1444_,
		_w1445_,
		_w1446_
	);
	LUT3 #(
		.INIT('h02)
	) name518 (
		decrypt_i_pad,
		\mix1_data_o_reg_reg[106]/NET0131 ,
		_w995_,
		_w1447_
	);
	LUT4 #(
		.INIT('hae00)
	) name519 (
		\data_o[106]_pad ,
		decrypt_i_pad,
		_w995_,
		_w1028_,
		_w1448_
	);
	LUT3 #(
		.INIT('h02)
	) name520 (
		decrypt_i_pad,
		\mix1_data_o_reg_reg[82]/NET0131 ,
		_w995_,
		_w1449_
	);
	LUT4 #(
		.INIT('hae00)
	) name521 (
		\data_o[82]_pad ,
		decrypt_i_pad,
		_w995_,
		_w1049_,
		_w1450_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name522 (
		_w1447_,
		_w1448_,
		_w1449_,
		_w1450_,
		_w1451_
	);
	LUT3 #(
		.INIT('h02)
	) name523 (
		decrypt_i_pad,
		\mix1_data_o_reg_reg[114]/NET0131 ,
		_w995_,
		_w1452_
	);
	LUT4 #(
		.INIT('hae00)
	) name524 (
		\data_o[114]_pad ,
		decrypt_i_pad,
		_w995_,
		_w1002_,
		_w1453_
	);
	LUT3 #(
		.INIT('h02)
	) name525 (
		decrypt_i_pad,
		\mix1_data_o_reg_reg[18]/NET0131 ,
		_w995_,
		_w1454_
	);
	LUT4 #(
		.INIT('hae00)
	) name526 (
		\data_o[18]_pad ,
		decrypt_i_pad,
		_w995_,
		_w1023_,
		_w1455_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name527 (
		_w1452_,
		_w1453_,
		_w1454_,
		_w1455_,
		_w1456_
	);
	LUT4 #(
		.INIT('h8000)
	) name528 (
		_w1451_,
		_w1456_,
		_w1441_,
		_w1446_,
		_w1457_
	);
	LUT3 #(
		.INIT('h02)
	) name529 (
		decrypt_i_pad,
		\mix1_data_o_reg_reg[34]/NET0131 ,
		_w995_,
		_w1458_
	);
	LUT4 #(
		.INIT('hae00)
	) name530 (
		\data_o[34]_pad ,
		decrypt_i_pad,
		_w995_,
		_w1042_,
		_w1459_
	);
	LUT2 #(
		.INIT('h4)
	) name531 (
		_w1458_,
		_w1459_,
		_w1460_
	);
	LUT3 #(
		.INIT('h02)
	) name532 (
		decrypt_i_pad,
		\mix1_data_o_reg_reg[74]/NET0131 ,
		_w995_,
		_w1461_
	);
	LUT4 #(
		.INIT('hae00)
	) name533 (
		\data_o[74]_pad ,
		decrypt_i_pad,
		_w995_,
		_w1035_,
		_w1462_
	);
	LUT3 #(
		.INIT('h02)
	) name534 (
		decrypt_i_pad,
		\mix1_data_o_reg_reg[2]/NET0131 ,
		_w995_,
		_w1463_
	);
	LUT4 #(
		.INIT('hae00)
	) name535 (
		\data_o[2]_pad ,
		decrypt_i_pad,
		_w995_,
		_w1009_,
		_w1464_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name536 (
		_w1461_,
		_w1462_,
		_w1463_,
		_w1464_,
		_w1465_
	);
	LUT3 #(
		.INIT('h02)
	) name537 (
		decrypt_i_pad,
		\mix1_data_o_reg_reg[42]/NET0131 ,
		_w995_,
		_w1466_
	);
	LUT4 #(
		.INIT('hae00)
	) name538 (
		\data_o[42]_pad ,
		decrypt_i_pad,
		_w995_,
		_w1006_,
		_w1467_
	);
	LUT3 #(
		.INIT('h02)
	) name539 (
		decrypt_i_pad,
		\mix1_data_o_reg_reg[26]/NET0131 ,
		_w995_,
		_w1468_
	);
	LUT4 #(
		.INIT('hae00)
	) name540 (
		\data_o[26]_pad ,
		decrypt_i_pad,
		_w995_,
		_w1020_,
		_w1469_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name541 (
		_w1466_,
		_w1467_,
		_w1468_,
		_w1469_,
		_w1470_
	);
	LUT3 #(
		.INIT('h02)
	) name542 (
		decrypt_i_pad,
		\mix1_data_o_reg_reg[66]/NET0131 ,
		_w995_,
		_w1471_
	);
	LUT4 #(
		.INIT('hae00)
	) name543 (
		\data_o[66]_pad ,
		decrypt_i_pad,
		_w995_,
		_w1039_,
		_w1472_
	);
	LUT3 #(
		.INIT('h02)
	) name544 (
		decrypt_i_pad,
		\mix1_data_o_reg_reg[10]/NET0131 ,
		_w995_,
		_w1473_
	);
	LUT4 #(
		.INIT('ha0e0)
	) name545 (
		\data_o[10]_pad ,
		decrypt_i_pad,
		_w1013_,
		_w995_,
		_w1474_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name546 (
		_w1471_,
		_w1472_,
		_w1473_,
		_w1474_,
		_w1475_
	);
	LUT4 #(
		.INIT('h4000)
	) name547 (
		_w1460_,
		_w1470_,
		_w1475_,
		_w1465_,
		_w1476_
	);
	LUT3 #(
		.INIT('h51)
	) name548 (
		\data_o[122]_pad ,
		decrypt_i_pad,
		_w995_,
		_w1477_
	);
	LUT3 #(
		.INIT('h02)
	) name549 (
		decrypt_i_pad,
		\mix1_data_o_reg_reg[122]/NET0131 ,
		_w995_,
		_w1478_
	);
	LUT3 #(
		.INIT('h02)
	) name550 (
		_w1060_,
		_w1478_,
		_w1477_,
		_w1479_
	);
	LUT2 #(
		.INIT('h8)
	) name551 (
		_w1057_,
		_w1479_,
		_w1480_
	);
	LUT4 #(
		.INIT('h00ea)
	) name552 (
		_w1053_,
		_w1457_,
		_w1476_,
		_w1480_,
		_w1481_
	);
	LUT3 #(
		.INIT('hc8)
	) name553 (
		\addroundkey_start_i_reg/NET0131 ,
		\key_i[26]_pad ,
		_w936_,
		_w1482_
	);
	LUT3 #(
		.INIT('h02)
	) name554 (
		\ks1_key_reg_reg[26]/NET0131 ,
		_w936_,
		_w938_,
		_w1483_
	);
	LUT4 #(
		.INIT('h0001)
	) name555 (
		\addroundkey_round_reg[1]/NET0131 ,
		\addroundkey_round_reg[2]/NET0131 ,
		\addroundkey_round_reg[3]/NET0131 ,
		\key_i[26]_pad ,
		_w1484_
	);
	LUT4 #(
		.INIT('h00fe)
	) name556 (
		\addroundkey_round_reg[1]/NET0131 ,
		\addroundkey_round_reg[2]/NET0131 ,
		\addroundkey_round_reg[3]/NET0131 ,
		\ks1_key_reg_reg[26]/NET0131 ,
		_w1485_
	);
	LUT4 #(
		.INIT('h0008)
	) name557 (
		\addroundkey_start_i_reg/NET0131 ,
		_w930_,
		_w1485_,
		_w1484_,
		_w1486_
	);
	LUT4 #(
		.INIT('h00ab)
	) name558 (
		_w931_,
		_w1482_,
		_w1483_,
		_w1486_,
		_w1487_
	);
	LUT3 #(
		.INIT('hc8)
	) name559 (
		\addroundkey_start_i_reg/NET0131 ,
		\key_i[18]_pad ,
		_w936_,
		_w1488_
	);
	LUT3 #(
		.INIT('h02)
	) name560 (
		\ks1_key_reg_reg[18]/NET0131 ,
		_w936_,
		_w938_,
		_w1489_
	);
	LUT4 #(
		.INIT('h0001)
	) name561 (
		\addroundkey_round_reg[1]/NET0131 ,
		\addroundkey_round_reg[2]/NET0131 ,
		\addroundkey_round_reg[3]/NET0131 ,
		\key_i[18]_pad ,
		_w1490_
	);
	LUT4 #(
		.INIT('h00fe)
	) name562 (
		\addroundkey_round_reg[1]/NET0131 ,
		\addroundkey_round_reg[2]/NET0131 ,
		\addroundkey_round_reg[3]/NET0131 ,
		\ks1_key_reg_reg[18]/NET0131 ,
		_w1491_
	);
	LUT4 #(
		.INIT('h0008)
	) name563 (
		\addroundkey_start_i_reg/NET0131 ,
		_w930_,
		_w1491_,
		_w1490_,
		_w1492_
	);
	LUT4 #(
		.INIT('h00ab)
	) name564 (
		_w931_,
		_w1488_,
		_w1489_,
		_w1492_,
		_w1493_
	);
	LUT4 #(
		.INIT('hf531)
	) name565 (
		_w948_,
		_w1079_,
		_w1487_,
		_w1493_,
		_w1494_
	);
	LUT3 #(
		.INIT('hc8)
	) name566 (
		\addroundkey_start_i_reg/NET0131 ,
		\key_i[10]_pad ,
		_w936_,
		_w1495_
	);
	LUT3 #(
		.INIT('h02)
	) name567 (
		\ks1_key_reg_reg[10]/NET0131 ,
		_w936_,
		_w938_,
		_w1496_
	);
	LUT4 #(
		.INIT('h0001)
	) name568 (
		\addroundkey_round_reg[1]/NET0131 ,
		\addroundkey_round_reg[2]/NET0131 ,
		\addroundkey_round_reg[3]/NET0131 ,
		\key_i[10]_pad ,
		_w1497_
	);
	LUT4 #(
		.INIT('h00fe)
	) name569 (
		\addroundkey_round_reg[1]/NET0131 ,
		\addroundkey_round_reg[2]/NET0131 ,
		\addroundkey_round_reg[3]/NET0131 ,
		\ks1_key_reg_reg[10]/NET0131 ,
		_w1498_
	);
	LUT4 #(
		.INIT('h0008)
	) name570 (
		\addroundkey_start_i_reg/NET0131 ,
		_w930_,
		_w1498_,
		_w1497_,
		_w1499_
	);
	LUT4 #(
		.INIT('h00ab)
	) name571 (
		_w931_,
		_w1495_,
		_w1496_,
		_w1499_,
		_w1500_
	);
	LUT3 #(
		.INIT('hc8)
	) name572 (
		\addroundkey_start_i_reg/NET0131 ,
		\key_i[2]_pad ,
		_w936_,
		_w1501_
	);
	LUT3 #(
		.INIT('h02)
	) name573 (
		\ks1_key_reg_reg[2]/NET0131 ,
		_w936_,
		_w938_,
		_w1502_
	);
	LUT4 #(
		.INIT('h0001)
	) name574 (
		\addroundkey_round_reg[1]/NET0131 ,
		\addroundkey_round_reg[2]/NET0131 ,
		\addroundkey_round_reg[3]/NET0131 ,
		\key_i[2]_pad ,
		_w1503_
	);
	LUT4 #(
		.INIT('h00fe)
	) name575 (
		\addroundkey_round_reg[1]/NET0131 ,
		\addroundkey_round_reg[2]/NET0131 ,
		\addroundkey_round_reg[3]/NET0131 ,
		\ks1_key_reg_reg[2]/NET0131 ,
		_w1504_
	);
	LUT4 #(
		.INIT('h0008)
	) name576 (
		\addroundkey_start_i_reg/NET0131 ,
		_w930_,
		_w1504_,
		_w1503_,
		_w1505_
	);
	LUT4 #(
		.INIT('h00ab)
	) name577 (
		_w931_,
		_w1501_,
		_w1502_,
		_w1505_,
		_w1506_
	);
	LUT4 #(
		.INIT('hf351)
	) name578 (
		_w1064_,
		_w1071_,
		_w1500_,
		_w1506_,
		_w1507_
	);
	LUT4 #(
		.INIT('hd000)
	) name579 (
		_w950_,
		_w1481_,
		_w1494_,
		_w1507_,
		_w1508_
	);
	LUT2 #(
		.INIT('h1)
	) name580 (
		_w951_,
		_w1508_,
		_w1509_
	);
	LUT3 #(
		.INIT('hc8)
	) name581 (
		\addroundkey_start_i_reg/NET0131 ,
		\key_i[23]_pad ,
		_w936_,
		_w1510_
	);
	LUT3 #(
		.INIT('h02)
	) name582 (
		\ks1_key_reg_reg[23]/NET0131 ,
		_w936_,
		_w938_,
		_w1511_
	);
	LUT4 #(
		.INIT('h0001)
	) name583 (
		\addroundkey_round_reg[1]/NET0131 ,
		\addroundkey_round_reg[2]/NET0131 ,
		\addroundkey_round_reg[3]/NET0131 ,
		\key_i[23]_pad ,
		_w1512_
	);
	LUT4 #(
		.INIT('h00fe)
	) name584 (
		\addroundkey_round_reg[1]/NET0131 ,
		\addroundkey_round_reg[2]/NET0131 ,
		\addroundkey_round_reg[3]/NET0131 ,
		\ks1_key_reg_reg[23]/NET0131 ,
		_w1513_
	);
	LUT4 #(
		.INIT('h0008)
	) name585 (
		\addroundkey_start_i_reg/NET0131 ,
		_w930_,
		_w1513_,
		_w1512_,
		_w1514_
	);
	LUT4 #(
		.INIT('h00ab)
	) name586 (
		_w931_,
		_w1510_,
		_w1511_,
		_w1514_,
		_w1515_
	);
	LUT3 #(
		.INIT('hc8)
	) name587 (
		\addroundkey_start_i_reg/NET0131 ,
		\key_i[7]_pad ,
		_w936_,
		_w1516_
	);
	LUT3 #(
		.INIT('h02)
	) name588 (
		\ks1_key_reg_reg[7]/NET0131 ,
		_w936_,
		_w938_,
		_w1517_
	);
	LUT4 #(
		.INIT('h0001)
	) name589 (
		\addroundkey_round_reg[1]/NET0131 ,
		\addroundkey_round_reg[2]/NET0131 ,
		\addroundkey_round_reg[3]/NET0131 ,
		\key_i[7]_pad ,
		_w1518_
	);
	LUT4 #(
		.INIT('h00fe)
	) name590 (
		\addroundkey_round_reg[1]/NET0131 ,
		\addroundkey_round_reg[2]/NET0131 ,
		\addroundkey_round_reg[3]/NET0131 ,
		\ks1_key_reg_reg[7]/NET0131 ,
		_w1519_
	);
	LUT4 #(
		.INIT('h0008)
	) name591 (
		\addroundkey_start_i_reg/NET0131 ,
		_w930_,
		_w1519_,
		_w1518_,
		_w1520_
	);
	LUT4 #(
		.INIT('h00ab)
	) name592 (
		_w931_,
		_w1516_,
		_w1517_,
		_w1520_,
		_w1521_
	);
	LUT4 #(
		.INIT('hf351)
	) name593 (
		_w1064_,
		_w1079_,
		_w1515_,
		_w1521_,
		_w1522_
	);
	LUT3 #(
		.INIT('hc8)
	) name594 (
		\addroundkey_start_i_reg/NET0131 ,
		\key_i[15]_pad ,
		_w936_,
		_w1523_
	);
	LUT3 #(
		.INIT('h02)
	) name595 (
		\ks1_key_reg_reg[15]/NET0131 ,
		_w936_,
		_w938_,
		_w1524_
	);
	LUT4 #(
		.INIT('h0001)
	) name596 (
		\addroundkey_round_reg[1]/NET0131 ,
		\addroundkey_round_reg[2]/NET0131 ,
		\addroundkey_round_reg[3]/NET0131 ,
		\key_i[15]_pad ,
		_w1525_
	);
	LUT4 #(
		.INIT('h00fe)
	) name597 (
		\addroundkey_round_reg[1]/NET0131 ,
		\addroundkey_round_reg[2]/NET0131 ,
		\addroundkey_round_reg[3]/NET0131 ,
		\ks1_key_reg_reg[15]/NET0131 ,
		_w1526_
	);
	LUT4 #(
		.INIT('h0008)
	) name598 (
		\addroundkey_start_i_reg/NET0131 ,
		_w930_,
		_w1526_,
		_w1525_,
		_w1527_
	);
	LUT4 #(
		.INIT('h00ab)
	) name599 (
		_w931_,
		_w1523_,
		_w1524_,
		_w1527_,
		_w1528_
	);
	LUT3 #(
		.INIT('hc8)
	) name600 (
		\addroundkey_start_i_reg/NET0131 ,
		\key_i[31]_pad ,
		_w936_,
		_w1529_
	);
	LUT3 #(
		.INIT('h02)
	) name601 (
		\ks1_key_reg_reg[31]/NET0131 ,
		_w936_,
		_w938_,
		_w1530_
	);
	LUT4 #(
		.INIT('h0001)
	) name602 (
		\addroundkey_round_reg[1]/NET0131 ,
		\addroundkey_round_reg[2]/NET0131 ,
		\addroundkey_round_reg[3]/NET0131 ,
		\key_i[31]_pad ,
		_w1531_
	);
	LUT4 #(
		.INIT('h00fe)
	) name603 (
		\addroundkey_round_reg[1]/NET0131 ,
		\addroundkey_round_reg[2]/NET0131 ,
		\addroundkey_round_reg[3]/NET0131 ,
		\ks1_key_reg_reg[31]/NET0131 ,
		_w1532_
	);
	LUT4 #(
		.INIT('h0008)
	) name604 (
		\addroundkey_start_i_reg/NET0131 ,
		_w930_,
		_w1532_,
		_w1531_,
		_w1533_
	);
	LUT4 #(
		.INIT('h00ab)
	) name605 (
		_w931_,
		_w1529_,
		_w1530_,
		_w1533_,
		_w1534_
	);
	LUT4 #(
		.INIT('hf351)
	) name606 (
		_w948_,
		_w1071_,
		_w1528_,
		_w1534_,
		_w1535_
	);
	LUT3 #(
		.INIT('h02)
	) name607 (
		decrypt_i_pad,
		\mix1_data_o_reg_reg[87]/NET0131 ,
		_w995_,
		_w1536_
	);
	LUT4 #(
		.INIT('hae00)
	) name608 (
		\data_o[87]_pad ,
		decrypt_i_pad,
		_w995_,
		_w1049_,
		_w1537_
	);
	LUT3 #(
		.INIT('h02)
	) name609 (
		decrypt_i_pad,
		\mix1_data_o_reg_reg[63]/NET0131 ,
		_w995_,
		_w1538_
	);
	LUT4 #(
		.INIT('hae00)
	) name610 (
		\data_o[63]_pad ,
		decrypt_i_pad,
		_w995_,
		_w999_,
		_w1539_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name611 (
		_w1536_,
		_w1537_,
		_w1538_,
		_w1539_,
		_w1540_
	);
	LUT3 #(
		.INIT('h02)
	) name612 (
		decrypt_i_pad,
		\mix1_data_o_reg_reg[55]/NET0131 ,
		_w995_,
		_w1541_
	);
	LUT4 #(
		.INIT('hae00)
	) name613 (
		\data_o[55]_pad ,
		decrypt_i_pad,
		_w995_,
		_w1046_,
		_w1542_
	);
	LUT3 #(
		.INIT('h02)
	) name614 (
		decrypt_i_pad,
		\mix1_data_o_reg_reg[95]/NET0131 ,
		_w995_,
		_w1543_
	);
	LUT4 #(
		.INIT('hae00)
	) name615 (
		\data_o[95]_pad ,
		decrypt_i_pad,
		_w995_,
		_w1032_,
		_w1544_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name616 (
		_w1541_,
		_w1542_,
		_w1543_,
		_w1544_,
		_w1545_
	);
	LUT3 #(
		.INIT('h02)
	) name617 (
		decrypt_i_pad,
		\mix1_data_o_reg_reg[15]/NET0131 ,
		_w995_,
		_w1546_
	);
	LUT4 #(
		.INIT('ha0e0)
	) name618 (
		\data_o[15]_pad ,
		decrypt_i_pad,
		_w1013_,
		_w995_,
		_w1547_
	);
	LUT3 #(
		.INIT('h02)
	) name619 (
		decrypt_i_pad,
		\mix1_data_o_reg_reg[39]/NET0131 ,
		_w995_,
		_w1548_
	);
	LUT4 #(
		.INIT('hae00)
	) name620 (
		\data_o[39]_pad ,
		decrypt_i_pad,
		_w995_,
		_w1042_,
		_w1549_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name621 (
		_w1546_,
		_w1547_,
		_w1548_,
		_w1549_,
		_w1550_
	);
	LUT3 #(
		.INIT('h02)
	) name622 (
		decrypt_i_pad,
		\mix1_data_o_reg_reg[31]/NET0131 ,
		_w995_,
		_w1551_
	);
	LUT4 #(
		.INIT('hae00)
	) name623 (
		\data_o[31]_pad ,
		decrypt_i_pad,
		_w995_,
		_w1020_,
		_w1552_
	);
	LUT3 #(
		.INIT('h02)
	) name624 (
		decrypt_i_pad,
		\mix1_data_o_reg_reg[23]/NET0131 ,
		_w995_,
		_w1553_
	);
	LUT4 #(
		.INIT('hae00)
	) name625 (
		\data_o[23]_pad ,
		decrypt_i_pad,
		_w995_,
		_w1023_,
		_w1554_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name626 (
		_w1551_,
		_w1552_,
		_w1553_,
		_w1554_,
		_w1555_
	);
	LUT4 #(
		.INIT('h8000)
	) name627 (
		_w1550_,
		_w1555_,
		_w1540_,
		_w1545_,
		_w1556_
	);
	LUT3 #(
		.INIT('h02)
	) name628 (
		decrypt_i_pad,
		\mix1_data_o_reg_reg[119]/NET0131 ,
		_w995_,
		_w1557_
	);
	LUT4 #(
		.INIT('hae00)
	) name629 (
		\data_o[119]_pad ,
		decrypt_i_pad,
		_w995_,
		_w1002_,
		_w1558_
	);
	LUT2 #(
		.INIT('h4)
	) name630 (
		_w1557_,
		_w1558_,
		_w1559_
	);
	LUT3 #(
		.INIT('h02)
	) name631 (
		decrypt_i_pad,
		\mix1_data_o_reg_reg[79]/NET0131 ,
		_w995_,
		_w1560_
	);
	LUT4 #(
		.INIT('hae00)
	) name632 (
		\data_o[79]_pad ,
		decrypt_i_pad,
		_w995_,
		_w1035_,
		_w1561_
	);
	LUT3 #(
		.INIT('h02)
	) name633 (
		decrypt_i_pad,
		\mix1_data_o_reg_reg[7]/NET0131 ,
		_w995_,
		_w1562_
	);
	LUT4 #(
		.INIT('hae00)
	) name634 (
		\data_o[7]_pad ,
		decrypt_i_pad,
		_w995_,
		_w1009_,
		_w1563_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name635 (
		_w1560_,
		_w1561_,
		_w1562_,
		_w1563_,
		_w1564_
	);
	LUT3 #(
		.INIT('h02)
	) name636 (
		decrypt_i_pad,
		\mix1_data_o_reg_reg[47]/NET0131 ,
		_w995_,
		_w1565_
	);
	LUT4 #(
		.INIT('hae00)
	) name637 (
		\data_o[47]_pad ,
		decrypt_i_pad,
		_w995_,
		_w1006_,
		_w1566_
	);
	LUT3 #(
		.INIT('h02)
	) name638 (
		decrypt_i_pad,
		\mix1_data_o_reg_reg[103]/NET0131 ,
		_w995_,
		_w1567_
	);
	LUT4 #(
		.INIT('hae00)
	) name639 (
		\data_o[103]_pad ,
		decrypt_i_pad,
		_w995_,
		_w1016_,
		_w1568_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name640 (
		_w1565_,
		_w1566_,
		_w1567_,
		_w1568_,
		_w1569_
	);
	LUT3 #(
		.INIT('h02)
	) name641 (
		decrypt_i_pad,
		\mix1_data_o_reg_reg[71]/NET0131 ,
		_w995_,
		_w1570_
	);
	LUT4 #(
		.INIT('hae00)
	) name642 (
		\data_o[71]_pad ,
		decrypt_i_pad,
		_w995_,
		_w1039_,
		_w1571_
	);
	LUT3 #(
		.INIT('h02)
	) name643 (
		decrypt_i_pad,
		\mix1_data_o_reg_reg[111]/NET0131 ,
		_w995_,
		_w1572_
	);
	LUT4 #(
		.INIT('hae00)
	) name644 (
		\data_o[111]_pad ,
		decrypt_i_pad,
		_w995_,
		_w1028_,
		_w1573_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name645 (
		_w1570_,
		_w1571_,
		_w1572_,
		_w1573_,
		_w1574_
	);
	LUT4 #(
		.INIT('h4000)
	) name646 (
		_w1559_,
		_w1569_,
		_w1574_,
		_w1564_,
		_w1575_
	);
	LUT3 #(
		.INIT('h51)
	) name647 (
		\data_o[127]_pad ,
		decrypt_i_pad,
		_w995_,
		_w1576_
	);
	LUT3 #(
		.INIT('h02)
	) name648 (
		decrypt_i_pad,
		\mix1_data_o_reg_reg[127]/NET0131 ,
		_w995_,
		_w1577_
	);
	LUT3 #(
		.INIT('h02)
	) name649 (
		_w1060_,
		_w1577_,
		_w1576_,
		_w1578_
	);
	LUT2 #(
		.INIT('h8)
	) name650 (
		_w1057_,
		_w1578_,
		_w1579_
	);
	LUT4 #(
		.INIT('h00ea)
	) name651 (
		_w1053_,
		_w1556_,
		_w1575_,
		_w1579_,
		_w1580_
	);
	LUT4 #(
		.INIT('hea40)
	) name652 (
		_w950_,
		_w1522_,
		_w1535_,
		_w1580_,
		_w1581_
	);
	LUT4 #(
		.INIT('h8228)
	) name653 (
		_w951_,
		_w1093_,
		_w1295_,
		_w1581_,
		_w1582_
	);
	LUT2 #(
		.INIT('h1)
	) name654 (
		_w1509_,
		_w1582_,
		_w1583_
	);
	LUT4 #(
		.INIT('h111e)
	) name655 (
		_w1094_,
		_w1296_,
		_w1509_,
		_w1582_,
		_w1584_
	);
	LUT4 #(
		.INIT('h2882)
	) name656 (
		_w951_,
		_w1093_,
		_w1508_,
		_w1581_,
		_w1585_
	);
	LUT2 #(
		.INIT('h1)
	) name657 (
		_w951_,
		_w1433_,
		_w1586_
	);
	LUT2 #(
		.INIT('h1)
	) name658 (
		_w1585_,
		_w1586_,
		_w1587_
	);
	LUT2 #(
		.INIT('h6)
	) name659 (
		_w1436_,
		_w1587_,
		_w1588_
	);
	LUT3 #(
		.INIT('h21)
	) name660 (
		_w1436_,
		_w1584_,
		_w1587_,
		_w1589_
	);
	LUT4 #(
		.INIT('h2882)
	) name661 (
		_w951_,
		_w1433_,
		_w1508_,
		_w1581_,
		_w1590_
	);
	LUT2 #(
		.INIT('h4)
	) name662 (
		_w951_,
		_w1365_,
		_w1591_
	);
	LUT2 #(
		.INIT('h1)
	) name663 (
		_w1590_,
		_w1591_,
		_w1592_
	);
	LUT4 #(
		.INIT('h9669)
	) name664 (
		_w1436_,
		_w1584_,
		_w1587_,
		_w1592_,
		_w1593_
	);
	LUT4 #(
		.INIT('h2882)
	) name665 (
		_w1436_,
		_w1584_,
		_w1587_,
		_w1592_,
		_w1594_
	);
	LUT2 #(
		.INIT('h1)
	) name666 (
		_w951_,
		_w1295_,
		_w1595_
	);
	LUT4 #(
		.INIT('h2882)
	) name667 (
		_w951_,
		_w1151_,
		_w1223_,
		_w1365_,
		_w1596_
	);
	LUT2 #(
		.INIT('h1)
	) name668 (
		_w951_,
		_w1581_,
		_w1597_
	);
	LUT4 #(
		.INIT('h2882)
	) name669 (
		_w951_,
		_w1093_,
		_w1151_,
		_w1295_,
		_w1598_
	);
	LUT2 #(
		.INIT('h1)
	) name670 (
		_w1597_,
		_w1598_,
		_w1599_
	);
	LUT4 #(
		.INIT('h111e)
	) name671 (
		_w1595_,
		_w1596_,
		_w1597_,
		_w1598_,
		_w1600_
	);
	LUT3 #(
		.INIT('h31)
	) name672 (
		_w1593_,
		_w1594_,
		_w1600_,
		_w1601_
	);
	LUT4 #(
		.INIT('h111e)
	) name673 (
		_w1509_,
		_w1582_,
		_w1595_,
		_w1596_,
		_w1602_
	);
	LUT3 #(
		.INIT('h06)
	) name674 (
		_w1436_,
		_w1587_,
		_w1602_,
		_w1603_
	);
	LUT4 #(
		.INIT('heee1)
	) name675 (
		_w1585_,
		_w1586_,
		_w1597_,
		_w1598_,
		_w1604_
	);
	LUT4 #(
		.INIT('h111e)
	) name676 (
		_w1585_,
		_w1586_,
		_w1597_,
		_w1598_,
		_w1605_
	);
	LUT4 #(
		.INIT('h2882)
	) name677 (
		_w951_,
		_w1365_,
		_w1433_,
		_w1508_,
		_w1606_
	);
	LUT2 #(
		.INIT('h1)
	) name678 (
		_w951_,
		_w1223_,
		_w1607_
	);
	LUT4 #(
		.INIT('heee1)
	) name679 (
		_w1509_,
		_w1582_,
		_w1606_,
		_w1607_,
		_w1608_
	);
	LUT2 #(
		.INIT('h6)
	) name680 (
		_w1604_,
		_w1608_,
		_w1609_
	);
	LUT4 #(
		.INIT('h0660)
	) name681 (
		_w1584_,
		_w1600_,
		_w1604_,
		_w1608_,
		_w1610_
	);
	LUT3 #(
		.INIT('h18)
	) name682 (
		_w1583_,
		_w1587_,
		_w1599_,
		_w1611_
	);
	LUT3 #(
		.INIT('h96)
	) name683 (
		_w1603_,
		_w1610_,
		_w1611_,
		_w1612_
	);
	LUT2 #(
		.INIT('h6)
	) name684 (
		_w1601_,
		_w1612_,
		_w1613_
	);
	LUT3 #(
		.INIT('h28)
	) name685 (
		_w1602_,
		_w1604_,
		_w1608_,
		_w1614_
	);
	LUT2 #(
		.INIT('h9)
	) name686 (
		_w1589_,
		_w1614_,
		_w1615_
	);
	LUT2 #(
		.INIT('h1)
	) name687 (
		_w1436_,
		_w1600_,
		_w1616_
	);
	LUT3 #(
		.INIT('h1e)
	) name688 (
		_w1593_,
		_w1604_,
		_w1616_,
		_w1617_
	);
	LUT2 #(
		.INIT('h9)
	) name689 (
		_w1615_,
		_w1617_,
		_w1618_
	);
	LUT2 #(
		.INIT('h4)
	) name690 (
		_w1593_,
		_w1609_,
		_w1619_
	);
	LUT3 #(
		.INIT('h60)
	) name691 (
		_w1436_,
		_w1587_,
		_w1600_,
		_w1620_
	);
	LUT2 #(
		.INIT('h1)
	) name692 (
		_w1584_,
		_w1604_,
		_w1621_
	);
	LUT3 #(
		.INIT('h06)
	) name693 (
		_w1584_,
		_w1600_,
		_w1604_,
		_w1622_
	);
	LUT3 #(
		.INIT('h8d)
	) name694 (
		_w1620_,
		_w1621_,
		_w1622_,
		_w1623_
	);
	LUT2 #(
		.INIT('h9)
	) name695 (
		_w1436_,
		_w1600_,
		_w1624_
	);
	LUT4 #(
		.INIT('h9655)
	) name696 (
		_w1297_,
		_w1436_,
		_w1600_,
		_w1602_,
		_w1625_
	);
	LUT3 #(
		.INIT('h69)
	) name697 (
		_w1619_,
		_w1623_,
		_w1625_,
		_w1626_
	);
	LUT2 #(
		.INIT('h8)
	) name698 (
		\sbox1_alph_reg[1]/NET0131 ,
		_w952_,
		_w1627_
	);
	LUT2 #(
		.INIT('h8)
	) name699 (
		\sbox1_alph_reg[3]/NET0131 ,
		_w956_,
		_w1628_
	);
	LUT4 #(
		.INIT('hf539)
	) name700 (
		\sbox1_alph_reg[0]/NET0131 ,
		\sbox1_alph_reg[2]/NET0131 ,
		_w954_,
		_w957_,
		_w1629_
	);
	LUT3 #(
		.INIT('h69)
	) name701 (
		_w1627_,
		_w1628_,
		_w1629_,
		_w1630_
	);
	LUT2 #(
		.INIT('h6)
	) name702 (
		_w959_,
		_w1630_,
		_w1631_
	);
	LUT3 #(
		.INIT('h96)
	) name703 (
		_w959_,
		_w978_,
		_w982_,
		_w1632_
	);
	LUT4 #(
		.INIT('hdd2d)
	) name704 (
		\sbox1_ah_reg_reg[2]/NET0131 ,
		_w952_,
		_w956_,
		_w962_,
		_w1633_
	);
	LUT2 #(
		.INIT('h2)
	) name705 (
		\sbox1_ah_reg_reg[1]/NET0131 ,
		_w954_,
		_w1634_
	);
	LUT2 #(
		.INIT('h9)
	) name706 (
		_w1633_,
		_w1634_,
		_w1635_
	);
	LUT3 #(
		.INIT('h53)
	) name707 (
		\sbox1_ah_reg_reg[2]/NET0131 ,
		\sbox1_ah_reg_reg[3]/NET0131 ,
		_w957_,
		_w1636_
	);
	LUT3 #(
		.INIT('h69)
	) name708 (
		_w955_,
		_w958_,
		_w1636_,
		_w1637_
	);
	LUT2 #(
		.INIT('h6)
	) name709 (
		_w1635_,
		_w1637_,
		_w1638_
	);
	LUT2 #(
		.INIT('h6)
	) name710 (
		_w1632_,
		_w1638_,
		_w1639_
	);
	LUT4 #(
		.INIT('h4114)
	) name711 (
		_w951_,
		_w984_,
		_w1632_,
		_w1638_,
		_w1640_
	);
	LUT4 #(
		.INIT('haaac)
	) name712 (
		\key_i[104]_pad ,
		\ks1_key_reg_reg[104]/NET0131 ,
		_w938_,
		_w986_,
		_w1641_
	);
	LUT3 #(
		.INIT('h96)
	) name713 (
		_w1631_,
		_w1640_,
		_w1641_,
		_w1642_
	);
	LUT4 #(
		.INIT('haaac)
	) name714 (
		\key_i[72]_pad ,
		\ks1_key_reg_reg[72]/P0002 ,
		_w938_,
		_w986_,
		_w1643_
	);
	LUT4 #(
		.INIT('h6996)
	) name715 (
		_w1631_,
		_w1640_,
		_w1641_,
		_w1643_,
		_w1644_
	);
	LUT4 #(
		.INIT('haaac)
	) name716 (
		\key_i[40]_pad ,
		\ks1_key_reg_reg[40]/P0002 ,
		_w938_,
		_w986_,
		_w1645_
	);
	LUT2 #(
		.INIT('h6)
	) name717 (
		_w1644_,
		_w1645_,
		_w1646_
	);
	LUT4 #(
		.INIT('h2882)
	) name718 (
		_w929_,
		_w1350_,
		_w1644_,
		_w1645_,
		_w1647_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name719 (
		\ks1_key_reg_reg[8]/NET0131 ,
		\ks1_state_reg[0]/NET0131 ,
		\ks1_state_reg[1]/NET0131 ,
		\ks1_state_reg[2]/NET0131 ,
		_w1648_
	);
	LUT2 #(
		.INIT('he)
	) name720 (
		_w1647_,
		_w1648_,
		_w1649_
	);
	LUT4 #(
		.INIT('h5553)
	) name721 (
		\key_i[74]_pad ,
		\ks1_key_reg_reg[74]/NET0131 ,
		_w938_,
		_w986_,
		_w1650_
	);
	LUT3 #(
		.INIT('hc8)
	) name722 (
		\addroundkey_start_i_reg/NET0131 ,
		\key_i[106]_pad ,
		_w936_,
		_w1651_
	);
	LUT3 #(
		.INIT('h02)
	) name723 (
		\ks1_key_reg_reg[106]/NET0131 ,
		_w936_,
		_w938_,
		_w1652_
	);
	LUT4 #(
		.INIT('h0001)
	) name724 (
		\addroundkey_round_reg[1]/NET0131 ,
		\addroundkey_round_reg[2]/NET0131 ,
		\addroundkey_round_reg[3]/NET0131 ,
		\key_i[106]_pad ,
		_w1653_
	);
	LUT4 #(
		.INIT('h00fe)
	) name725 (
		\addroundkey_round_reg[1]/NET0131 ,
		\addroundkey_round_reg[2]/NET0131 ,
		\addroundkey_round_reg[3]/NET0131 ,
		\ks1_key_reg_reg[106]/NET0131 ,
		_w1654_
	);
	LUT4 #(
		.INIT('h0008)
	) name726 (
		\addroundkey_start_i_reg/NET0131 ,
		_w930_,
		_w1654_,
		_w1653_,
		_w1655_
	);
	LUT4 #(
		.INIT('h00ab)
	) name727 (
		_w931_,
		_w1651_,
		_w1652_,
		_w1655_,
		_w1656_
	);
	LUT3 #(
		.INIT('h96)
	) name728 (
		_w959_,
		_w978_,
		_w1630_,
		_w1657_
	);
	LUT3 #(
		.INIT('h96)
	) name729 (
		_w964_,
		_w1635_,
		_w1637_,
		_w1658_
	);
	LUT3 #(
		.INIT('h82)
	) name730 (
		_w951_,
		_w1631_,
		_w1658_,
		_w1659_
	);
	LUT3 #(
		.INIT('h14)
	) name731 (
		_w951_,
		_w1632_,
		_w1638_,
		_w1660_
	);
	LUT3 #(
		.INIT('h56)
	) name732 (
		_w1657_,
		_w1659_,
		_w1660_,
		_w1661_
	);
	LUT4 #(
		.INIT('h9996)
	) name733 (
		_w1656_,
		_w1657_,
		_w1659_,
		_w1660_,
		_w1662_
	);
	LUT4 #(
		.INIT('h6669)
	) name734 (
		_w1656_,
		_w1657_,
		_w1659_,
		_w1660_,
		_w1663_
	);
	LUT4 #(
		.INIT('haaac)
	) name735 (
		\key_i[42]_pad ,
		\ks1_key_reg_reg[42]/P0002 ,
		_w938_,
		_w986_,
		_w1664_
	);
	LUT3 #(
		.INIT('h69)
	) name736 (
		_w1650_,
		_w1662_,
		_w1664_,
		_w1665_
	);
	LUT3 #(
		.INIT('h96)
	) name737 (
		_w1650_,
		_w1662_,
		_w1664_,
		_w1666_
	);
	LUT4 #(
		.INIT('h2ee2)
	) name738 (
		\ks1_key_reg_reg[10]/NET0131 ,
		_w929_,
		_w1500_,
		_w1665_,
		_w1667_
	);
	LUT3 #(
		.INIT('h1e)
	) name739 (
		\sub1_state_reg[0]/NET0131 ,
		\sub1_state_reg[1]/NET0131 ,
		\sub1_state_reg[2]/NET0131 ,
		_w1668_
	);
	LUT2 #(
		.INIT('h6)
	) name740 (
		\sub1_state_reg[0]/NET0131 ,
		\sub1_state_reg[1]/NET0131 ,
		_w1669_
	);
	LUT4 #(
		.INIT('h0018)
	) name741 (
		\sub1_state_reg[0]/NET0131 ,
		\sub1_state_reg[1]/NET0131 ,
		\sub1_state_reg[2]/NET0131 ,
		\sub1_state_reg[4]/NET0131 ,
		_w1670_
	);
	LUT4 #(
		.INIT('h0154)
	) name742 (
		\sub1_state_reg[0]/NET0131 ,
		\sub1_state_reg[1]/NET0131 ,
		\sub1_state_reg[2]/NET0131 ,
		\sub1_state_reg[3]/NET0131 ,
		_w1671_
	);
	LUT2 #(
		.INIT('h8)
	) name743 (
		_w1670_,
		_w1671_,
		_w1672_
	);
	LUT4 #(
		.INIT('h3222)
	) name744 (
		\sub1_data_reg_reg[102]/NET0131 ,
		_w1053_,
		_w1670_,
		_w1671_,
		_w1673_
	);
	LUT3 #(
		.INIT('h20)
	) name745 (
		\sub1_data_reg_reg[102]/NET0131 ,
		\sub1_state_reg[4]/NET0131 ,
		_w1053_,
		_w1674_
	);
	LUT4 #(
		.INIT('h4114)
	) name746 (
		decrypt_i_pad,
		_w959_,
		_w964_,
		_w970_,
		_w1675_
	);
	LUT2 #(
		.INIT('h2)
	) name747 (
		decrypt_i_pad,
		\sub1_data_reg_reg[70]/NET0131 ,
		_w1676_
	);
	LUT2 #(
		.INIT('h8)
	) name748 (
		\sub1_state_reg[4]/NET0131 ,
		_w1053_,
		_w1677_
	);
	LUT3 #(
		.INIT('h08)
	) name749 (
		\sub1_state_reg[4]/NET0131 ,
		_w1053_,
		_w1676_,
		_w1678_
	);
	LUT3 #(
		.INIT('h45)
	) name750 (
		_w1674_,
		_w1675_,
		_w1678_,
		_w1679_
	);
	LUT4 #(
		.INIT('h70ff)
	) name751 (
		_w985_,
		_w1672_,
		_w1673_,
		_w1679_,
		_w1680_
	);
	LUT3 #(
		.INIT('h69)
	) name752 (
		_w975_,
		_w1635_,
		_w1637_,
		_w1681_
	);
	LUT3 #(
		.INIT('h96)
	) name753 (
		_w970_,
		_w1635_,
		_w1637_,
		_w1682_
	);
	LUT4 #(
		.INIT('heb41)
	) name754 (
		_w951_,
		_w984_,
		_w1682_,
		_w1681_,
		_w1683_
	);
	LUT4 #(
		.INIT('h3222)
	) name755 (
		\sub1_data_reg_reg[101]/NET0131 ,
		_w1053_,
		_w1670_,
		_w1671_,
		_w1684_
	);
	LUT3 #(
		.INIT('hd0)
	) name756 (
		_w1672_,
		_w1683_,
		_w1684_,
		_w1685_
	);
	LUT3 #(
		.INIT('h20)
	) name757 (
		\sub1_data_reg_reg[101]/NET0131 ,
		\sub1_state_reg[4]/NET0131 ,
		_w1053_,
		_w1686_
	);
	LUT2 #(
		.INIT('h2)
	) name758 (
		decrypt_i_pad,
		\sub1_data_reg_reg[69]/NET0131 ,
		_w1687_
	);
	LUT3 #(
		.INIT('h08)
	) name759 (
		\sub1_state_reg[4]/NET0131 ,
		_w1053_,
		_w1687_,
		_w1688_
	);
	LUT4 #(
		.INIT('heb00)
	) name760 (
		decrypt_i_pad,
		_w984_,
		_w1682_,
		_w1688_,
		_w1689_
	);
	LUT2 #(
		.INIT('h1)
	) name761 (
		_w1686_,
		_w1689_,
		_w1690_
	);
	LUT2 #(
		.INIT('hb)
	) name762 (
		_w1685_,
		_w1690_,
		_w1691_
	);
	LUT4 #(
		.INIT('h0006)
	) name763 (
		\sub1_state_reg[0]/NET0131 ,
		\sub1_state_reg[1]/NET0131 ,
		\sub1_state_reg[2]/NET0131 ,
		\sub1_state_reg[4]/NET0131 ,
		_w1692_
	);
	LUT2 #(
		.INIT('h8)
	) name764 (
		_w1671_,
		_w1692_,
		_w1693_
	);
	LUT4 #(
		.INIT('h3222)
	) name765 (
		\sub1_data_reg_reg[117]/NET0131 ,
		_w1053_,
		_w1671_,
		_w1692_,
		_w1694_
	);
	LUT3 #(
		.INIT('hd8)
	) name766 (
		decrypt_i_pad,
		\sub1_data_reg_reg[21]/NET0131 ,
		\sub1_data_reg_reg[85]/NET0131 ,
		_w1695_
	);
	LUT4 #(
		.INIT('h1fdf)
	) name767 (
		\sub1_data_reg_reg[117]/NET0131 ,
		\sub1_state_reg[4]/NET0131 ,
		_w1053_,
		_w1695_,
		_w1696_
	);
	LUT4 #(
		.INIT('hb0ff)
	) name768 (
		_w1683_,
		_w1693_,
		_w1694_,
		_w1696_,
		_w1697_
	);
	LUT4 #(
		.INIT('h3222)
	) name769 (
		\sub1_data_reg_reg[118]/NET0131 ,
		_w1053_,
		_w1671_,
		_w1692_,
		_w1698_
	);
	LUT3 #(
		.INIT('hd8)
	) name770 (
		decrypt_i_pad,
		\sub1_data_reg_reg[22]/NET0131 ,
		\sub1_data_reg_reg[86]/NET0131 ,
		_w1699_
	);
	LUT4 #(
		.INIT('h1fdf)
	) name771 (
		\sub1_data_reg_reg[118]/NET0131 ,
		\sub1_state_reg[4]/NET0131 ,
		_w1053_,
		_w1699_,
		_w1700_
	);
	LUT4 #(
		.INIT('h70ff)
	) name772 (
		_w985_,
		_w1693_,
		_w1698_,
		_w1700_,
		_w1701_
	);
	LUT4 #(
		.INIT('h0900)
	) name773 (
		\sub1_state_reg[4]/NET0131 ,
		_w1053_,
		_w1668_,
		_w1669_,
		_w1702_
	);
	LUT4 #(
		.INIT('h1044)
	) name774 (
		\sub1_state_reg[0]/NET0131 ,
		\sub1_state_reg[3]/NET0131 ,
		\sub1_state_reg[4]/NET0131 ,
		_w998_,
		_w1703_
	);
	LUT2 #(
		.INIT('h8)
	) name775 (
		_w1702_,
		_w1703_,
		_w1704_
	);
	LUT4 #(
		.INIT('h3222)
	) name776 (
		\sub1_data_reg_reg[21]/NET0131 ,
		_w1053_,
		_w1702_,
		_w1703_,
		_w1705_
	);
	LUT3 #(
		.INIT('he4)
	) name777 (
		decrypt_i_pad,
		\sub1_data_reg_reg[117]/NET0131 ,
		\sub1_data_reg_reg[53]/NET0131 ,
		_w1706_
	);
	LUT4 #(
		.INIT('h1fdf)
	) name778 (
		\sub1_data_reg_reg[21]/NET0131 ,
		\sub1_state_reg[4]/NET0131 ,
		_w1053_,
		_w1706_,
		_w1707_
	);
	LUT4 #(
		.INIT('hb0ff)
	) name779 (
		_w1683_,
		_w1704_,
		_w1705_,
		_w1707_,
		_w1708_
	);
	LUT4 #(
		.INIT('h3222)
	) name780 (
		\sub1_data_reg_reg[22]/NET0131 ,
		_w1053_,
		_w1702_,
		_w1703_,
		_w1709_
	);
	LUT3 #(
		.INIT('he4)
	) name781 (
		decrypt_i_pad,
		\sub1_data_reg_reg[118]/NET0131 ,
		\sub1_data_reg_reg[54]/NET0131 ,
		_w1710_
	);
	LUT4 #(
		.INIT('h1fdf)
	) name782 (
		\sub1_data_reg_reg[22]/NET0131 ,
		\sub1_state_reg[4]/NET0131 ,
		_w1053_,
		_w1710_,
		_w1711_
	);
	LUT4 #(
		.INIT('h70ff)
	) name783 (
		_w985_,
		_w1704_,
		_w1709_,
		_w1711_,
		_w1712_
	);
	LUT2 #(
		.INIT('h8)
	) name784 (
		_w1670_,
		_w1703_,
		_w1713_
	);
	LUT4 #(
		.INIT('h8b88)
	) name785 (
		\sub1_state_reg[4]/NET0131 ,
		_w1053_,
		_w1683_,
		_w1713_,
		_w1714_
	);
	LUT3 #(
		.INIT('h40)
	) name786 (
		_w1053_,
		_w1683_,
		_w1713_,
		_w1715_
	);
	LUT2 #(
		.INIT('h1)
	) name787 (
		decrypt_i_pad,
		\sub1_data_reg_reg[69]/NET0131 ,
		_w1716_
	);
	LUT3 #(
		.INIT('h08)
	) name788 (
		\sub1_state_reg[4]/NET0131 ,
		_w1053_,
		_w1716_,
		_w1717_
	);
	LUT3 #(
		.INIT('hd0)
	) name789 (
		decrypt_i_pad,
		_w1683_,
		_w1717_,
		_w1718_
	);
	LUT4 #(
		.INIT('hffce)
	) name790 (
		\sub1_data_reg_reg[37]/NET0131 ,
		_w1715_,
		_w1714_,
		_w1718_,
		_w1719_
	);
	LUT2 #(
		.INIT('h1)
	) name791 (
		decrypt_i_pad,
		\sub1_data_reg_reg[70]/NET0131 ,
		_w1720_
	);
	LUT3 #(
		.INIT('h08)
	) name792 (
		\sub1_state_reg[4]/NET0131 ,
		_w1053_,
		_w1720_,
		_w1721_
	);
	LUT3 #(
		.INIT('h70)
	) name793 (
		decrypt_i_pad,
		_w985_,
		_w1721_,
		_w1722_
	);
	LUT3 #(
		.INIT('h20)
	) name794 (
		\sub1_data_reg_reg[38]/NET0131 ,
		\sub1_state_reg[4]/NET0131 ,
		_w1053_,
		_w1723_
	);
	LUT4 #(
		.INIT('h3222)
	) name795 (
		\sub1_data_reg_reg[38]/NET0131 ,
		_w1053_,
		_w1670_,
		_w1703_,
		_w1724_
	);
	LUT4 #(
		.INIT('h080f)
	) name796 (
		_w985_,
		_w1713_,
		_w1723_,
		_w1724_,
		_w1725_
	);
	LUT2 #(
		.INIT('hb)
	) name797 (
		_w1722_,
		_w1725_,
		_w1726_
	);
	LUT2 #(
		.INIT('h8)
	) name798 (
		_w1692_,
		_w1703_,
		_w1727_
	);
	LUT4 #(
		.INIT('h3222)
	) name799 (
		\sub1_data_reg_reg[53]/NET0131 ,
		_w1053_,
		_w1692_,
		_w1703_,
		_w1728_
	);
	LUT3 #(
		.INIT('he4)
	) name800 (
		decrypt_i_pad,
		\sub1_data_reg_reg[21]/NET0131 ,
		\sub1_data_reg_reg[85]/NET0131 ,
		_w1729_
	);
	LUT4 #(
		.INIT('h1fdf)
	) name801 (
		\sub1_data_reg_reg[53]/NET0131 ,
		\sub1_state_reg[4]/NET0131 ,
		_w1053_,
		_w1729_,
		_w1730_
	);
	LUT4 #(
		.INIT('hb0ff)
	) name802 (
		_w1683_,
		_w1727_,
		_w1728_,
		_w1730_,
		_w1731_
	);
	LUT4 #(
		.INIT('h3222)
	) name803 (
		\sub1_data_reg_reg[54]/NET0131 ,
		_w1053_,
		_w1692_,
		_w1703_,
		_w1732_
	);
	LUT3 #(
		.INIT('he4)
	) name804 (
		decrypt_i_pad,
		\sub1_data_reg_reg[22]/NET0131 ,
		\sub1_data_reg_reg[86]/NET0131 ,
		_w1733_
	);
	LUT4 #(
		.INIT('h1fdf)
	) name805 (
		\sub1_data_reg_reg[54]/NET0131 ,
		\sub1_state_reg[4]/NET0131 ,
		_w1053_,
		_w1733_,
		_w1734_
	);
	LUT4 #(
		.INIT('h70ff)
	) name806 (
		_w985_,
		_w1727_,
		_w1732_,
		_w1734_,
		_w1735_
	);
	LUT4 #(
		.INIT('h0009)
	) name807 (
		\sub1_state_reg[4]/NET0131 ,
		_w1053_,
		_w1668_,
		_w1669_,
		_w1736_
	);
	LUT3 #(
		.INIT('hd8)
	) name808 (
		decrypt_i_pad,
		\sub1_data_reg_reg[101]/NET0131 ,
		\sub1_data_reg_reg[37]/NET0131 ,
		_w1737_
	);
	LUT3 #(
		.INIT('h80)
	) name809 (
		\sub1_state_reg[4]/NET0131 ,
		_w1053_,
		_w1737_,
		_w1738_
	);
	LUT4 #(
		.INIT('hff2a)
	) name810 (
		\sub1_data_reg_reg[5]/NET0131 ,
		_w1703_,
		_w1736_,
		_w1738_,
		_w1739_
	);
	LUT3 #(
		.INIT('hd8)
	) name811 (
		decrypt_i_pad,
		\sub1_data_reg_reg[102]/NET0131 ,
		\sub1_data_reg_reg[38]/NET0131 ,
		_w1740_
	);
	LUT3 #(
		.INIT('h80)
	) name812 (
		\sub1_state_reg[4]/NET0131 ,
		_w1053_,
		_w1740_,
		_w1741_
	);
	LUT4 #(
		.INIT('hff2a)
	) name813 (
		\sub1_data_reg_reg[6]/NET0131 ,
		_w1703_,
		_w1736_,
		_w1741_,
		_w1742_
	);
	LUT2 #(
		.INIT('h8)
	) name814 (
		_w1671_,
		_w1736_,
		_w1743_
	);
	LUT4 #(
		.INIT('h3222)
	) name815 (
		\sub1_data_reg_reg[69]/NET0131 ,
		_w1053_,
		_w1671_,
		_w1736_,
		_w1744_
	);
	LUT3 #(
		.INIT('he4)
	) name816 (
		decrypt_i_pad,
		\sub1_data_reg_reg[101]/NET0131 ,
		\sub1_data_reg_reg[37]/NET0131 ,
		_w1745_
	);
	LUT4 #(
		.INIT('h1fdf)
	) name817 (
		\sub1_data_reg_reg[69]/NET0131 ,
		\sub1_state_reg[4]/NET0131 ,
		_w1053_,
		_w1745_,
		_w1746_
	);
	LUT4 #(
		.INIT('hb0ff)
	) name818 (
		_w1683_,
		_w1743_,
		_w1744_,
		_w1746_,
		_w1747_
	);
	LUT4 #(
		.INIT('h3222)
	) name819 (
		\sub1_data_reg_reg[70]/NET0131 ,
		_w1053_,
		_w1671_,
		_w1736_,
		_w1748_
	);
	LUT3 #(
		.INIT('he4)
	) name820 (
		decrypt_i_pad,
		\sub1_data_reg_reg[102]/NET0131 ,
		\sub1_data_reg_reg[38]/NET0131 ,
		_w1749_
	);
	LUT4 #(
		.INIT('h1fdf)
	) name821 (
		\sub1_data_reg_reg[70]/NET0131 ,
		\sub1_state_reg[4]/NET0131 ,
		_w1053_,
		_w1749_,
		_w1750_
	);
	LUT4 #(
		.INIT('h70ff)
	) name822 (
		_w985_,
		_w1743_,
		_w1748_,
		_w1750_,
		_w1751_
	);
	LUT2 #(
		.INIT('h8)
	) name823 (
		_w1671_,
		_w1702_,
		_w1752_
	);
	LUT4 #(
		.INIT('h3222)
	) name824 (
		\sub1_data_reg_reg[85]/NET0131 ,
		_w1053_,
		_w1671_,
		_w1702_,
		_w1753_
	);
	LUT3 #(
		.INIT('hd8)
	) name825 (
		decrypt_i_pad,
		\sub1_data_reg_reg[117]/NET0131 ,
		\sub1_data_reg_reg[53]/NET0131 ,
		_w1754_
	);
	LUT4 #(
		.INIT('h1fdf)
	) name826 (
		\sub1_data_reg_reg[85]/NET0131 ,
		\sub1_state_reg[4]/NET0131 ,
		_w1053_,
		_w1754_,
		_w1755_
	);
	LUT4 #(
		.INIT('hb0ff)
	) name827 (
		_w1683_,
		_w1752_,
		_w1753_,
		_w1755_,
		_w1756_
	);
	LUT4 #(
		.INIT('h3222)
	) name828 (
		\sub1_data_reg_reg[86]/NET0131 ,
		_w1053_,
		_w1671_,
		_w1702_,
		_w1757_
	);
	LUT3 #(
		.INIT('hd8)
	) name829 (
		decrypt_i_pad,
		\sub1_data_reg_reg[118]/NET0131 ,
		\sub1_data_reg_reg[54]/NET0131 ,
		_w1758_
	);
	LUT4 #(
		.INIT('h1fdf)
	) name830 (
		\sub1_data_reg_reg[86]/NET0131 ,
		\sub1_state_reg[4]/NET0131 ,
		_w1053_,
		_w1758_,
		_w1759_
	);
	LUT4 #(
		.INIT('h70ff)
	) name831 (
		_w985_,
		_w1752_,
		_w1757_,
		_w1759_,
		_w1760_
	);
	LUT2 #(
		.INIT('h2)
	) name832 (
		\sub1_state_reg[0]/NET0131 ,
		\sub1_state_reg[3]/NET0131 ,
		_w1761_
	);
	LUT2 #(
		.INIT('h8)
	) name833 (
		_w1670_,
		_w1761_,
		_w1762_
	);
	LUT4 #(
		.INIT('h3222)
	) name834 (
		\sub1_data_reg_reg[109]/NET0131 ,
		_w1053_,
		_w1670_,
		_w1761_,
		_w1763_
	);
	LUT4 #(
		.INIT('h35ff)
	) name835 (
		\sub1_data_reg_reg[109]/NET0131 ,
		\sub1_data_reg_reg[45]/NET0131 ,
		\sub1_state_reg[4]/NET0131 ,
		_w1053_,
		_w1764_
	);
	LUT4 #(
		.INIT('hb0ff)
	) name836 (
		_w1683_,
		_w1762_,
		_w1763_,
		_w1764_,
		_w1765_
	);
	LUT4 #(
		.INIT('h3222)
	) name837 (
		\sub1_data_reg_reg[110]/NET0131 ,
		_w1053_,
		_w1670_,
		_w1761_,
		_w1766_
	);
	LUT4 #(
		.INIT('h35ff)
	) name838 (
		\sub1_data_reg_reg[110]/NET0131 ,
		\sub1_data_reg_reg[46]/NET0131 ,
		\sub1_state_reg[4]/NET0131 ,
		_w1053_,
		_w1767_
	);
	LUT4 #(
		.INIT('h70ff)
	) name839 (
		_w985_,
		_w1762_,
		_w1766_,
		_w1767_,
		_w1768_
	);
	LUT2 #(
		.INIT('h8)
	) name840 (
		\sub1_state_reg[0]/NET0131 ,
		\sub1_state_reg[3]/NET0131 ,
		_w1769_
	);
	LUT2 #(
		.INIT('h8)
	) name841 (
		_w1736_,
		_w1769_,
		_w1770_
	);
	LUT4 #(
		.INIT('h3222)
	) name842 (
		\sub1_data_reg_reg[13]/NET0131 ,
		_w1053_,
		_w1736_,
		_w1769_,
		_w1771_
	);
	LUT4 #(
		.INIT('h35ff)
	) name843 (
		\sub1_data_reg_reg[13]/NET0131 ,
		\sub1_data_reg_reg[77]/NET0131 ,
		\sub1_state_reg[4]/NET0131 ,
		_w1053_,
		_w1772_
	);
	LUT4 #(
		.INIT('hb0ff)
	) name844 (
		_w1683_,
		_w1770_,
		_w1771_,
		_w1772_,
		_w1773_
	);
	LUT4 #(
		.INIT('h3222)
	) name845 (
		\sub1_data_reg_reg[14]/NET0131 ,
		_w1053_,
		_w1736_,
		_w1769_,
		_w1774_
	);
	LUT4 #(
		.INIT('h35ff)
	) name846 (
		\sub1_data_reg_reg[14]/NET0131 ,
		\sub1_data_reg_reg[78]/NET0131 ,
		\sub1_state_reg[4]/NET0131 ,
		_w1053_,
		_w1775_
	);
	LUT4 #(
		.INIT('h70ff)
	) name847 (
		_w985_,
		_w1770_,
		_w1774_,
		_w1775_,
		_w1776_
	);
	LUT2 #(
		.INIT('h8)
	) name848 (
		_w1670_,
		_w1769_,
		_w1777_
	);
	LUT4 #(
		.INIT('h3222)
	) name849 (
		\sub1_data_reg_reg[45]/NET0131 ,
		_w1053_,
		_w1670_,
		_w1769_,
		_w1778_
	);
	LUT4 #(
		.INIT('h53ff)
	) name850 (
		\sub1_data_reg_reg[109]/NET0131 ,
		\sub1_data_reg_reg[45]/NET0131 ,
		\sub1_state_reg[4]/NET0131 ,
		_w1053_,
		_w1779_
	);
	LUT4 #(
		.INIT('hb0ff)
	) name851 (
		_w1683_,
		_w1777_,
		_w1778_,
		_w1779_,
		_w1780_
	);
	LUT4 #(
		.INIT('h3222)
	) name852 (
		\sub1_data_reg_reg[46]/NET0131 ,
		_w1053_,
		_w1670_,
		_w1769_,
		_w1781_
	);
	LUT4 #(
		.INIT('h53ff)
	) name853 (
		\sub1_data_reg_reg[110]/NET0131 ,
		\sub1_data_reg_reg[46]/NET0131 ,
		\sub1_state_reg[4]/NET0131 ,
		_w1053_,
		_w1782_
	);
	LUT4 #(
		.INIT('h70ff)
	) name854 (
		_w985_,
		_w1777_,
		_w1781_,
		_w1782_,
		_w1783_
	);
	LUT2 #(
		.INIT('h8)
	) name855 (
		_w1736_,
		_w1761_,
		_w1784_
	);
	LUT4 #(
		.INIT('h3222)
	) name856 (
		\sub1_data_reg_reg[77]/NET0131 ,
		_w1053_,
		_w1736_,
		_w1761_,
		_w1785_
	);
	LUT4 #(
		.INIT('h53ff)
	) name857 (
		\sub1_data_reg_reg[13]/NET0131 ,
		\sub1_data_reg_reg[77]/NET0131 ,
		\sub1_state_reg[4]/NET0131 ,
		_w1053_,
		_w1786_
	);
	LUT4 #(
		.INIT('hb0ff)
	) name858 (
		_w1683_,
		_w1784_,
		_w1785_,
		_w1786_,
		_w1787_
	);
	LUT4 #(
		.INIT('h3222)
	) name859 (
		\sub1_data_reg_reg[78]/NET0131 ,
		_w1053_,
		_w1736_,
		_w1761_,
		_w1788_
	);
	LUT4 #(
		.INIT('h53ff)
	) name860 (
		\sub1_data_reg_reg[14]/NET0131 ,
		\sub1_data_reg_reg[78]/NET0131 ,
		\sub1_state_reg[4]/NET0131 ,
		_w1053_,
		_w1789_
	);
	LUT4 #(
		.INIT('h70ff)
	) name861 (
		_w985_,
		_w1784_,
		_w1788_,
		_w1789_,
		_w1790_
	);
	LUT3 #(
		.INIT('h1b)
	) name862 (
		decrypt_i_pad,
		\sub1_data_reg_reg[32]/NET0131 ,
		\sub1_data_reg_reg[96]/NET0131 ,
		_w1791_
	);
	LUT4 #(
		.INIT('h2aea)
	) name863 (
		\sub1_data_reg_reg[0]/NET0131 ,
		\sub1_state_reg[4]/NET0131 ,
		_w1053_,
		_w1791_,
		_w1792_
	);
	LUT4 #(
		.INIT('h6996)
	) name864 (
		_w970_,
		_w978_,
		_w1635_,
		_w1637_,
		_w1793_
	);
	LUT4 #(
		.INIT('h782d)
	) name865 (
		_w951_,
		_w959_,
		_w984_,
		_w1793_,
		_w1794_
	);
	LUT4 #(
		.INIT('h4515)
	) name866 (
		_w1053_,
		_w1639_,
		_w1672_,
		_w1794_,
		_w1795_
	);
	LUT3 #(
		.INIT('ha8)
	) name867 (
		\sub1_data_reg_reg[103]/NET0131 ,
		_w1060_,
		_w1795_,
		_w1796_
	);
	LUT4 #(
		.INIT('h4010)
	) name868 (
		_w1053_,
		_w1639_,
		_w1672_,
		_w1794_,
		_w1797_
	);
	LUT2 #(
		.INIT('h2)
	) name869 (
		decrypt_i_pad,
		\sub1_data_reg_reg[71]/NET0131 ,
		_w1798_
	);
	LUT3 #(
		.INIT('h08)
	) name870 (
		\sub1_state_reg[4]/NET0131 ,
		_w1053_,
		_w1798_,
		_w1799_
	);
	LUT4 #(
		.INIT('heb00)
	) name871 (
		decrypt_i_pad,
		_w1639_,
		_w1794_,
		_w1799_,
		_w1800_
	);
	LUT2 #(
		.INIT('h1)
	) name872 (
		_w1797_,
		_w1800_,
		_w1801_
	);
	LUT2 #(
		.INIT('hb)
	) name873 (
		_w1796_,
		_w1801_,
		_w1802_
	);
	LUT4 #(
		.INIT('h3222)
	) name874 (
		\sub1_data_reg_reg[112]/NET0131 ,
		_w1053_,
		_w1671_,
		_w1692_,
		_w1803_
	);
	LUT4 #(
		.INIT('h6f00)
	) name875 (
		_w1631_,
		_w1640_,
		_w1693_,
		_w1803_,
		_w1804_
	);
	LUT3 #(
		.INIT('hd8)
	) name876 (
		decrypt_i_pad,
		\sub1_data_reg_reg[16]/NET0131 ,
		\sub1_data_reg_reg[80]/NET0131 ,
		_w1805_
	);
	LUT4 #(
		.INIT('h1fdf)
	) name877 (
		\sub1_data_reg_reg[112]/NET0131 ,
		\sub1_state_reg[4]/NET0131 ,
		_w1053_,
		_w1805_,
		_w1806_
	);
	LUT2 #(
		.INIT('hb)
	) name878 (
		_w1804_,
		_w1806_,
		_w1807_
	);
	LUT4 #(
		.INIT('h6996)
	) name879 (
		_w959_,
		_w964_,
		_w975_,
		_w1630_,
		_w1808_
	);
	LUT4 #(
		.INIT('h1b4e)
	) name880 (
		_w951_,
		_w970_,
		_w1793_,
		_w1808_,
		_w1809_
	);
	LUT4 #(
		.INIT('h3222)
	) name881 (
		\sub1_data_reg_reg[115]/NET0131 ,
		_w1053_,
		_w1671_,
		_w1692_,
		_w1810_
	);
	LUT3 #(
		.INIT('hd8)
	) name882 (
		decrypt_i_pad,
		\sub1_data_reg_reg[19]/NET0131 ,
		\sub1_data_reg_reg[83]/NET0131 ,
		_w1811_
	);
	LUT4 #(
		.INIT('h1fdf)
	) name883 (
		\sub1_data_reg_reg[115]/NET0131 ,
		\sub1_state_reg[4]/NET0131 ,
		_w1053_,
		_w1811_,
		_w1812_
	);
	LUT4 #(
		.INIT('hd0ff)
	) name884 (
		_w1693_,
		_w1809_,
		_w1810_,
		_w1812_,
		_w1813_
	);
	LUT3 #(
		.INIT('h96)
	) name885 (
		_w983_,
		_w1631_,
		_w1658_,
		_w1814_
	);
	LUT4 #(
		.INIT('h8008)
	) name886 (
		decrypt_i_pad,
		_w950_,
		_w959_,
		_w1630_,
		_w1815_
	);
	LUT3 #(
		.INIT('h0b)
	) name887 (
		_w951_,
		_w1682_,
		_w1815_,
		_w1816_
	);
	LUT4 #(
		.INIT('h3222)
	) name888 (
		\sub1_data_reg_reg[116]/NET0131 ,
		_w1053_,
		_w1671_,
		_w1692_,
		_w1817_
	);
	LUT4 #(
		.INIT('h7d00)
	) name889 (
		_w1693_,
		_w1814_,
		_w1816_,
		_w1817_,
		_w1818_
	);
	LUT3 #(
		.INIT('hd8)
	) name890 (
		decrypt_i_pad,
		\sub1_data_reg_reg[20]/NET0131 ,
		\sub1_data_reg_reg[84]/NET0131 ,
		_w1819_
	);
	LUT4 #(
		.INIT('h1fdf)
	) name891 (
		\sub1_data_reg_reg[116]/NET0131 ,
		\sub1_state_reg[4]/NET0131 ,
		_w1053_,
		_w1819_,
		_w1820_
	);
	LUT2 #(
		.INIT('hb)
	) name892 (
		_w1818_,
		_w1820_,
		_w1821_
	);
	LUT4 #(
		.INIT('h3222)
	) name893 (
		\sub1_data_reg_reg[119]/NET0131 ,
		_w1053_,
		_w1671_,
		_w1692_,
		_w1822_
	);
	LUT4 #(
		.INIT('hb700)
	) name894 (
		_w1639_,
		_w1693_,
		_w1794_,
		_w1822_,
		_w1823_
	);
	LUT3 #(
		.INIT('hd8)
	) name895 (
		decrypt_i_pad,
		\sub1_data_reg_reg[23]/NET0131 ,
		\sub1_data_reg_reg[87]/NET0131 ,
		_w1824_
	);
	LUT4 #(
		.INIT('h1fdf)
	) name896 (
		\sub1_data_reg_reg[119]/NET0131 ,
		\sub1_state_reg[4]/NET0131 ,
		_w1053_,
		_w1824_,
		_w1825_
	);
	LUT2 #(
		.INIT('hb)
	) name897 (
		_w1823_,
		_w1825_,
		_w1826_
	);
	LUT4 #(
		.INIT('h3222)
	) name898 (
		\sub1_data_reg_reg[16]/NET0131 ,
		_w1053_,
		_w1702_,
		_w1703_,
		_w1827_
	);
	LUT4 #(
		.INIT('h6f00)
	) name899 (
		_w1631_,
		_w1640_,
		_w1704_,
		_w1827_,
		_w1828_
	);
	LUT3 #(
		.INIT('he4)
	) name900 (
		decrypt_i_pad,
		\sub1_data_reg_reg[112]/NET0131 ,
		\sub1_data_reg_reg[48]/NET0131 ,
		_w1829_
	);
	LUT4 #(
		.INIT('h1fdf)
	) name901 (
		\sub1_data_reg_reg[16]/NET0131 ,
		\sub1_state_reg[4]/NET0131 ,
		_w1053_,
		_w1829_,
		_w1830_
	);
	LUT2 #(
		.INIT('hb)
	) name902 (
		_w1828_,
		_w1830_,
		_w1831_
	);
	LUT4 #(
		.INIT('h3222)
	) name903 (
		\sub1_data_reg_reg[19]/NET0131 ,
		_w1053_,
		_w1702_,
		_w1703_,
		_w1832_
	);
	LUT3 #(
		.INIT('he4)
	) name904 (
		decrypt_i_pad,
		\sub1_data_reg_reg[115]/NET0131 ,
		\sub1_data_reg_reg[51]/NET0131 ,
		_w1833_
	);
	LUT4 #(
		.INIT('h1fdf)
	) name905 (
		\sub1_data_reg_reg[19]/NET0131 ,
		\sub1_state_reg[4]/NET0131 ,
		_w1053_,
		_w1833_,
		_w1834_
	);
	LUT4 #(
		.INIT('hd0ff)
	) name906 (
		_w1704_,
		_w1809_,
		_w1832_,
		_w1834_,
		_w1835_
	);
	LUT4 #(
		.INIT('h3222)
	) name907 (
		\sub1_data_reg_reg[20]/NET0131 ,
		_w1053_,
		_w1702_,
		_w1703_,
		_w1836_
	);
	LUT4 #(
		.INIT('h7d00)
	) name908 (
		_w1704_,
		_w1814_,
		_w1816_,
		_w1836_,
		_w1837_
	);
	LUT3 #(
		.INIT('he4)
	) name909 (
		decrypt_i_pad,
		\sub1_data_reg_reg[116]/NET0131 ,
		\sub1_data_reg_reg[52]/NET0131 ,
		_w1838_
	);
	LUT4 #(
		.INIT('h1fdf)
	) name910 (
		\sub1_data_reg_reg[20]/NET0131 ,
		\sub1_state_reg[4]/NET0131 ,
		_w1053_,
		_w1838_,
		_w1839_
	);
	LUT2 #(
		.INIT('hb)
	) name911 (
		_w1837_,
		_w1839_,
		_w1840_
	);
	LUT4 #(
		.INIT('h3222)
	) name912 (
		\sub1_data_reg_reg[23]/NET0131 ,
		_w1053_,
		_w1702_,
		_w1703_,
		_w1841_
	);
	LUT4 #(
		.INIT('hb700)
	) name913 (
		_w1639_,
		_w1704_,
		_w1794_,
		_w1841_,
		_w1842_
	);
	LUT3 #(
		.INIT('he4)
	) name914 (
		decrypt_i_pad,
		\sub1_data_reg_reg[119]/NET0131 ,
		\sub1_data_reg_reg[55]/NET0131 ,
		_w1843_
	);
	LUT4 #(
		.INIT('h1fdf)
	) name915 (
		\sub1_data_reg_reg[23]/NET0131 ,
		\sub1_state_reg[4]/NET0131 ,
		_w1053_,
		_w1843_,
		_w1844_
	);
	LUT2 #(
		.INIT('hb)
	) name916 (
		_w1842_,
		_w1844_,
		_w1845_
	);
	LUT4 #(
		.INIT('h1551)
	) name917 (
		_w1053_,
		_w1713_,
		_w1814_,
		_w1816_,
		_w1846_
	);
	LUT3 #(
		.INIT('ha8)
	) name918 (
		\sub1_data_reg_reg[36]/NET0131 ,
		_w1060_,
		_w1846_,
		_w1847_
	);
	LUT4 #(
		.INIT('h0440)
	) name919 (
		_w1053_,
		_w1713_,
		_w1814_,
		_w1816_,
		_w1848_
	);
	LUT2 #(
		.INIT('h1)
	) name920 (
		decrypt_i_pad,
		\sub1_data_reg_reg[68]/NET0131 ,
		_w1849_
	);
	LUT3 #(
		.INIT('h08)
	) name921 (
		\sub1_state_reg[4]/NET0131 ,
		_w1053_,
		_w1849_,
		_w1850_
	);
	LUT4 #(
		.INIT('h7d00)
	) name922 (
		decrypt_i_pad,
		_w1814_,
		_w1816_,
		_w1850_,
		_w1851_
	);
	LUT2 #(
		.INIT('h1)
	) name923 (
		_w1848_,
		_w1851_,
		_w1852_
	);
	LUT2 #(
		.INIT('hb)
	) name924 (
		_w1847_,
		_w1852_,
		_w1853_
	);
	LUT3 #(
		.INIT('he4)
	) name925 (
		decrypt_i_pad,
		\sub1_data_reg_reg[35]/NET0131 ,
		\sub1_data_reg_reg[99]/NET0131 ,
		_w1854_
	);
	LUT3 #(
		.INIT('h80)
	) name926 (
		\sub1_state_reg[4]/NET0131 ,
		_w1053_,
		_w1854_,
		_w1855_
	);
	LUT4 #(
		.INIT('hff2a)
	) name927 (
		\sub1_data_reg_reg[3]/NET0131 ,
		_w1703_,
		_w1736_,
		_w1855_,
		_w1856_
	);
	LUT4 #(
		.INIT('h3222)
	) name928 (
		\sub1_data_reg_reg[48]/NET0131 ,
		_w1053_,
		_w1692_,
		_w1703_,
		_w1857_
	);
	LUT4 #(
		.INIT('h6f00)
	) name929 (
		_w1631_,
		_w1640_,
		_w1727_,
		_w1857_,
		_w1858_
	);
	LUT3 #(
		.INIT('he4)
	) name930 (
		decrypt_i_pad,
		\sub1_data_reg_reg[16]/NET0131 ,
		\sub1_data_reg_reg[80]/NET0131 ,
		_w1859_
	);
	LUT4 #(
		.INIT('h1fdf)
	) name931 (
		\sub1_data_reg_reg[48]/NET0131 ,
		\sub1_state_reg[4]/NET0131 ,
		_w1053_,
		_w1859_,
		_w1860_
	);
	LUT2 #(
		.INIT('hb)
	) name932 (
		_w1858_,
		_w1860_,
		_w1861_
	);
	LUT3 #(
		.INIT('hd8)
	) name933 (
		decrypt_i_pad,
		\sub1_data_reg_reg[100]/NET0131 ,
		\sub1_data_reg_reg[36]/NET0131 ,
		_w1862_
	);
	LUT3 #(
		.INIT('h80)
	) name934 (
		\sub1_state_reg[4]/NET0131 ,
		_w1053_,
		_w1862_,
		_w1863_
	);
	LUT4 #(
		.INIT('hff2a)
	) name935 (
		\sub1_data_reg_reg[4]/NET0131 ,
		_w1703_,
		_w1736_,
		_w1863_,
		_w1864_
	);
	LUT4 #(
		.INIT('h3222)
	) name936 (
		\sub1_data_reg_reg[51]/NET0131 ,
		_w1053_,
		_w1692_,
		_w1703_,
		_w1865_
	);
	LUT3 #(
		.INIT('he4)
	) name937 (
		decrypt_i_pad,
		\sub1_data_reg_reg[19]/NET0131 ,
		\sub1_data_reg_reg[83]/NET0131 ,
		_w1866_
	);
	LUT4 #(
		.INIT('h1fdf)
	) name938 (
		\sub1_data_reg_reg[51]/NET0131 ,
		\sub1_state_reg[4]/NET0131 ,
		_w1053_,
		_w1866_,
		_w1867_
	);
	LUT4 #(
		.INIT('hd0ff)
	) name939 (
		_w1727_,
		_w1809_,
		_w1865_,
		_w1867_,
		_w1868_
	);
	LUT4 #(
		.INIT('h3222)
	) name940 (
		\sub1_data_reg_reg[52]/NET0131 ,
		_w1053_,
		_w1692_,
		_w1703_,
		_w1869_
	);
	LUT4 #(
		.INIT('h7d00)
	) name941 (
		_w1727_,
		_w1814_,
		_w1816_,
		_w1869_,
		_w1870_
	);
	LUT3 #(
		.INIT('he4)
	) name942 (
		decrypt_i_pad,
		\sub1_data_reg_reg[20]/NET0131 ,
		\sub1_data_reg_reg[84]/NET0131 ,
		_w1871_
	);
	LUT4 #(
		.INIT('h1fdf)
	) name943 (
		\sub1_data_reg_reg[52]/NET0131 ,
		\sub1_state_reg[4]/NET0131 ,
		_w1053_,
		_w1871_,
		_w1872_
	);
	LUT2 #(
		.INIT('hb)
	) name944 (
		_w1870_,
		_w1872_,
		_w1873_
	);
	LUT4 #(
		.INIT('h3222)
	) name945 (
		\sub1_data_reg_reg[55]/NET0131 ,
		_w1053_,
		_w1692_,
		_w1703_,
		_w1874_
	);
	LUT4 #(
		.INIT('hb700)
	) name946 (
		_w1639_,
		_w1727_,
		_w1794_,
		_w1874_,
		_w1875_
	);
	LUT3 #(
		.INIT('he4)
	) name947 (
		decrypt_i_pad,
		\sub1_data_reg_reg[23]/NET0131 ,
		\sub1_data_reg_reg[87]/NET0131 ,
		_w1876_
	);
	LUT4 #(
		.INIT('h1fdf)
	) name948 (
		\sub1_data_reg_reg[55]/NET0131 ,
		\sub1_state_reg[4]/NET0131 ,
		_w1053_,
		_w1876_,
		_w1877_
	);
	LUT2 #(
		.INIT('hb)
	) name949 (
		_w1875_,
		_w1877_,
		_w1878_
	);
	LUT4 #(
		.INIT('h3222)
	) name950 (
		\sub1_data_reg_reg[64]/NET0131 ,
		_w1053_,
		_w1671_,
		_w1736_,
		_w1879_
	);
	LUT4 #(
		.INIT('h6f00)
	) name951 (
		_w1631_,
		_w1640_,
		_w1743_,
		_w1879_,
		_w1880_
	);
	LUT3 #(
		.INIT('hd8)
	) name952 (
		decrypt_i_pad,
		\sub1_data_reg_reg[32]/NET0131 ,
		\sub1_data_reg_reg[96]/NET0131 ,
		_w1881_
	);
	LUT4 #(
		.INIT('h1fdf)
	) name953 (
		\sub1_data_reg_reg[64]/NET0131 ,
		\sub1_state_reg[4]/NET0131 ,
		_w1053_,
		_w1881_,
		_w1882_
	);
	LUT2 #(
		.INIT('hb)
	) name954 (
		_w1880_,
		_w1882_,
		_w1883_
	);
	LUT4 #(
		.INIT('h3222)
	) name955 (
		\sub1_data_reg_reg[67]/NET0131 ,
		_w1053_,
		_w1671_,
		_w1736_,
		_w1884_
	);
	LUT3 #(
		.INIT('hd8)
	) name956 (
		decrypt_i_pad,
		\sub1_data_reg_reg[35]/NET0131 ,
		\sub1_data_reg_reg[99]/NET0131 ,
		_w1885_
	);
	LUT4 #(
		.INIT('h1fdf)
	) name957 (
		\sub1_data_reg_reg[67]/NET0131 ,
		\sub1_state_reg[4]/NET0131 ,
		_w1053_,
		_w1885_,
		_w1886_
	);
	LUT4 #(
		.INIT('hd0ff)
	) name958 (
		_w1743_,
		_w1809_,
		_w1884_,
		_w1886_,
		_w1887_
	);
	LUT4 #(
		.INIT('h3222)
	) name959 (
		\sub1_data_reg_reg[68]/NET0131 ,
		_w1053_,
		_w1671_,
		_w1736_,
		_w1888_
	);
	LUT4 #(
		.INIT('h7d00)
	) name960 (
		_w1743_,
		_w1814_,
		_w1816_,
		_w1888_,
		_w1889_
	);
	LUT3 #(
		.INIT('he4)
	) name961 (
		decrypt_i_pad,
		\sub1_data_reg_reg[100]/NET0131 ,
		\sub1_data_reg_reg[36]/NET0131 ,
		_w1890_
	);
	LUT4 #(
		.INIT('h1fdf)
	) name962 (
		\sub1_data_reg_reg[68]/NET0131 ,
		\sub1_state_reg[4]/NET0131 ,
		_w1053_,
		_w1890_,
		_w1891_
	);
	LUT2 #(
		.INIT('hb)
	) name963 (
		_w1889_,
		_w1891_,
		_w1892_
	);
	LUT4 #(
		.INIT('h3222)
	) name964 (
		\sub1_data_reg_reg[71]/NET0131 ,
		_w1053_,
		_w1671_,
		_w1736_,
		_w1893_
	);
	LUT4 #(
		.INIT('hb700)
	) name965 (
		_w1639_,
		_w1743_,
		_w1794_,
		_w1893_,
		_w1894_
	);
	LUT3 #(
		.INIT('he4)
	) name966 (
		decrypt_i_pad,
		\sub1_data_reg_reg[103]/NET0131 ,
		\sub1_data_reg_reg[39]/NET0131 ,
		_w1895_
	);
	LUT4 #(
		.INIT('h1fdf)
	) name967 (
		\sub1_data_reg_reg[71]/NET0131 ,
		\sub1_state_reg[4]/NET0131 ,
		_w1053_,
		_w1895_,
		_w1896_
	);
	LUT2 #(
		.INIT('hb)
	) name968 (
		_w1894_,
		_w1896_,
		_w1897_
	);
	LUT3 #(
		.INIT('hd8)
	) name969 (
		decrypt_i_pad,
		\sub1_data_reg_reg[103]/NET0131 ,
		\sub1_data_reg_reg[39]/NET0131 ,
		_w1898_
	);
	LUT3 #(
		.INIT('h80)
	) name970 (
		\sub1_state_reg[4]/NET0131 ,
		_w1053_,
		_w1898_,
		_w1899_
	);
	LUT4 #(
		.INIT('hff2a)
	) name971 (
		\sub1_data_reg_reg[7]/NET0131 ,
		_w1703_,
		_w1736_,
		_w1899_,
		_w1900_
	);
	LUT4 #(
		.INIT('h3222)
	) name972 (
		\sub1_data_reg_reg[80]/NET0131 ,
		_w1053_,
		_w1671_,
		_w1702_,
		_w1901_
	);
	LUT4 #(
		.INIT('h6f00)
	) name973 (
		_w1631_,
		_w1640_,
		_w1752_,
		_w1901_,
		_w1902_
	);
	LUT3 #(
		.INIT('hd8)
	) name974 (
		decrypt_i_pad,
		\sub1_data_reg_reg[112]/NET0131 ,
		\sub1_data_reg_reg[48]/NET0131 ,
		_w1903_
	);
	LUT4 #(
		.INIT('h1fdf)
	) name975 (
		\sub1_data_reg_reg[80]/NET0131 ,
		\sub1_state_reg[4]/NET0131 ,
		_w1053_,
		_w1903_,
		_w1904_
	);
	LUT2 #(
		.INIT('hb)
	) name976 (
		_w1902_,
		_w1904_,
		_w1905_
	);
	LUT4 #(
		.INIT('h3222)
	) name977 (
		\sub1_data_reg_reg[83]/NET0131 ,
		_w1053_,
		_w1671_,
		_w1702_,
		_w1906_
	);
	LUT3 #(
		.INIT('hd8)
	) name978 (
		decrypt_i_pad,
		\sub1_data_reg_reg[115]/NET0131 ,
		\sub1_data_reg_reg[51]/NET0131 ,
		_w1907_
	);
	LUT4 #(
		.INIT('h1fdf)
	) name979 (
		\sub1_data_reg_reg[83]/NET0131 ,
		\sub1_state_reg[4]/NET0131 ,
		_w1053_,
		_w1907_,
		_w1908_
	);
	LUT4 #(
		.INIT('hd0ff)
	) name980 (
		_w1752_,
		_w1809_,
		_w1906_,
		_w1908_,
		_w1909_
	);
	LUT4 #(
		.INIT('h3222)
	) name981 (
		\sub1_data_reg_reg[84]/NET0131 ,
		_w1053_,
		_w1671_,
		_w1702_,
		_w1910_
	);
	LUT4 #(
		.INIT('h7d00)
	) name982 (
		_w1752_,
		_w1814_,
		_w1816_,
		_w1910_,
		_w1911_
	);
	LUT3 #(
		.INIT('hd8)
	) name983 (
		decrypt_i_pad,
		\sub1_data_reg_reg[116]/NET0131 ,
		\sub1_data_reg_reg[52]/NET0131 ,
		_w1912_
	);
	LUT4 #(
		.INIT('h1fdf)
	) name984 (
		\sub1_data_reg_reg[84]/NET0131 ,
		\sub1_state_reg[4]/NET0131 ,
		_w1053_,
		_w1912_,
		_w1913_
	);
	LUT2 #(
		.INIT('hb)
	) name985 (
		_w1911_,
		_w1913_,
		_w1914_
	);
	LUT4 #(
		.INIT('h3222)
	) name986 (
		\sub1_data_reg_reg[87]/NET0131 ,
		_w1053_,
		_w1671_,
		_w1702_,
		_w1915_
	);
	LUT4 #(
		.INIT('hb700)
	) name987 (
		_w1639_,
		_w1752_,
		_w1794_,
		_w1915_,
		_w1916_
	);
	LUT3 #(
		.INIT('hd8)
	) name988 (
		decrypt_i_pad,
		\sub1_data_reg_reg[119]/NET0131 ,
		\sub1_data_reg_reg[55]/NET0131 ,
		_w1917_
	);
	LUT4 #(
		.INIT('h1fdf)
	) name989 (
		\sub1_data_reg_reg[87]/NET0131 ,
		\sub1_state_reg[4]/NET0131 ,
		_w1053_,
		_w1917_,
		_w1918_
	);
	LUT2 #(
		.INIT('hb)
	) name990 (
		_w1916_,
		_w1918_,
		_w1919_
	);
	LUT4 #(
		.INIT('h3222)
	) name991 (
		\sub1_data_reg_reg[96]/NET0131 ,
		_w1053_,
		_w1670_,
		_w1671_,
		_w1920_
	);
	LUT4 #(
		.INIT('h6f00)
	) name992 (
		_w1631_,
		_w1640_,
		_w1672_,
		_w1920_,
		_w1921_
	);
	LUT3 #(
		.INIT('h20)
	) name993 (
		\sub1_data_reg_reg[96]/NET0131 ,
		\sub1_state_reg[4]/NET0131 ,
		_w1053_,
		_w1922_
	);
	LUT2 #(
		.INIT('h2)
	) name994 (
		decrypt_i_pad,
		\sub1_data_reg_reg[64]/NET0131 ,
		_w1923_
	);
	LUT3 #(
		.INIT('h08)
	) name995 (
		\sub1_state_reg[4]/NET0131 ,
		_w1053_,
		_w1923_,
		_w1924_
	);
	LUT4 #(
		.INIT('hbe00)
	) name996 (
		decrypt_i_pad,
		_w1631_,
		_w1640_,
		_w1924_,
		_w1925_
	);
	LUT3 #(
		.INIT('hfe)
	) name997 (
		_w1922_,
		_w1925_,
		_w1921_,
		_w1926_
	);
	LUT4 #(
		.INIT('h3222)
	) name998 (
		\sub1_data_reg_reg[104]/NET0131 ,
		_w1053_,
		_w1670_,
		_w1761_,
		_w1927_
	);
	LUT4 #(
		.INIT('h6f00)
	) name999 (
		_w1631_,
		_w1640_,
		_w1762_,
		_w1927_,
		_w1928_
	);
	LUT4 #(
		.INIT('h35ff)
	) name1000 (
		\sub1_data_reg_reg[104]/NET0131 ,
		\sub1_data_reg_reg[40]/NET0131 ,
		\sub1_state_reg[4]/NET0131 ,
		_w1053_,
		_w1929_
	);
	LUT2 #(
		.INIT('hb)
	) name1001 (
		_w1928_,
		_w1929_,
		_w1930_
	);
	LUT4 #(
		.INIT('h3222)
	) name1002 (
		\sub1_data_reg_reg[107]/NET0131 ,
		_w1053_,
		_w1670_,
		_w1761_,
		_w1931_
	);
	LUT4 #(
		.INIT('h35ff)
	) name1003 (
		\sub1_data_reg_reg[107]/NET0131 ,
		\sub1_data_reg_reg[43]/NET0131 ,
		\sub1_state_reg[4]/NET0131 ,
		_w1053_,
		_w1932_
	);
	LUT4 #(
		.INIT('hd0ff)
	) name1004 (
		_w1762_,
		_w1809_,
		_w1931_,
		_w1932_,
		_w1933_
	);
	LUT4 #(
		.INIT('h3222)
	) name1005 (
		\sub1_data_reg_reg[108]/NET0131 ,
		_w1053_,
		_w1670_,
		_w1761_,
		_w1934_
	);
	LUT4 #(
		.INIT('h7d00)
	) name1006 (
		_w1762_,
		_w1814_,
		_w1816_,
		_w1934_,
		_w1935_
	);
	LUT4 #(
		.INIT('h35ff)
	) name1007 (
		\sub1_data_reg_reg[108]/NET0131 ,
		\sub1_data_reg_reg[44]/NET0131 ,
		\sub1_state_reg[4]/NET0131 ,
		_w1053_,
		_w1936_
	);
	LUT2 #(
		.INIT('hb)
	) name1008 (
		_w1935_,
		_w1936_,
		_w1937_
	);
	LUT4 #(
		.INIT('h3222)
	) name1009 (
		\sub1_data_reg_reg[111]/NET0131 ,
		_w1053_,
		_w1670_,
		_w1761_,
		_w1938_
	);
	LUT4 #(
		.INIT('hb700)
	) name1010 (
		_w1639_,
		_w1762_,
		_w1794_,
		_w1938_,
		_w1939_
	);
	LUT4 #(
		.INIT('h35ff)
	) name1011 (
		\sub1_data_reg_reg[111]/NET0131 ,
		\sub1_data_reg_reg[47]/NET0131 ,
		\sub1_state_reg[4]/NET0131 ,
		_w1053_,
		_w1940_
	);
	LUT2 #(
		.INIT('hb)
	) name1012 (
		_w1939_,
		_w1940_,
		_w1941_
	);
	LUT4 #(
		.INIT('h3222)
	) name1013 (
		\sub1_data_reg_reg[11]/NET0131 ,
		_w1053_,
		_w1736_,
		_w1769_,
		_w1942_
	);
	LUT4 #(
		.INIT('h35ff)
	) name1014 (
		\sub1_data_reg_reg[11]/NET0131 ,
		\sub1_data_reg_reg[75]/NET0131 ,
		\sub1_state_reg[4]/NET0131 ,
		_w1053_,
		_w1943_
	);
	LUT4 #(
		.INIT('hd0ff)
	) name1015 (
		_w1770_,
		_w1809_,
		_w1942_,
		_w1943_,
		_w1944_
	);
	LUT3 #(
		.INIT('h3a)
	) name1016 (
		\ks1_col_reg[30]/NET0131 ,
		_w985_,
		_w1071_,
		_w1945_
	);
	LUT3 #(
		.INIT('he2)
	) name1017 (
		\ks1_col_reg[21]/NET0131 ,
		_w1064_,
		_w1683_,
		_w1946_
	);
	LUT4 #(
		.INIT('h3222)
	) name1018 (
		\sub1_data_reg_reg[12]/NET0131 ,
		_w1053_,
		_w1736_,
		_w1769_,
		_w1947_
	);
	LUT4 #(
		.INIT('h7d00)
	) name1019 (
		_w1770_,
		_w1814_,
		_w1816_,
		_w1947_,
		_w1948_
	);
	LUT4 #(
		.INIT('h35ff)
	) name1020 (
		\sub1_data_reg_reg[12]/NET0131 ,
		\sub1_data_reg_reg[76]/NET0131 ,
		\sub1_state_reg[4]/NET0131 ,
		_w1053_,
		_w1949_
	);
	LUT2 #(
		.INIT('hb)
	) name1021 (
		_w1948_,
		_w1949_,
		_w1950_
	);
	LUT3 #(
		.INIT('h3a)
	) name1022 (
		\ks1_col_reg[22]/NET0131 ,
		_w985_,
		_w1064_,
		_w1951_
	);
	LUT4 #(
		.INIT('h3222)
	) name1023 (
		\sub1_data_reg_reg[15]/NET0131 ,
		_w1053_,
		_w1736_,
		_w1769_,
		_w1952_
	);
	LUT4 #(
		.INIT('hb700)
	) name1024 (
		_w1639_,
		_w1770_,
		_w1794_,
		_w1952_,
		_w1953_
	);
	LUT4 #(
		.INIT('h35ff)
	) name1025 (
		\sub1_data_reg_reg[15]/NET0131 ,
		\sub1_data_reg_reg[79]/NET0131 ,
		\sub1_state_reg[4]/NET0131 ,
		_w1053_,
		_w1954_
	);
	LUT2 #(
		.INIT('hb)
	) name1026 (
		_w1953_,
		_w1954_,
		_w1955_
	);
	LUT3 #(
		.INIT('h3a)
	) name1027 (
		\ks1_col_reg[6]/NET0131 ,
		_w985_,
		_w1079_,
		_w1956_
	);
	LUT3 #(
		.INIT('he2)
	) name1028 (
		\ks1_col_reg[29]/NET0131 ,
		_w1071_,
		_w1683_,
		_w1957_
	);
	LUT3 #(
		.INIT('he2)
	) name1029 (
		\ks1_col_reg[5]/NET0131 ,
		_w1079_,
		_w1683_,
		_w1958_
	);
	LUT4 #(
		.INIT('h3222)
	) name1030 (
		\sub1_data_reg_reg[40]/NET0131 ,
		_w1053_,
		_w1670_,
		_w1769_,
		_w1959_
	);
	LUT4 #(
		.INIT('h6f00)
	) name1031 (
		_w1631_,
		_w1640_,
		_w1777_,
		_w1959_,
		_w1960_
	);
	LUT4 #(
		.INIT('h53ff)
	) name1032 (
		\sub1_data_reg_reg[104]/NET0131 ,
		\sub1_data_reg_reg[40]/NET0131 ,
		\sub1_state_reg[4]/NET0131 ,
		_w1053_,
		_w1961_
	);
	LUT2 #(
		.INIT('hb)
	) name1033 (
		_w1960_,
		_w1961_,
		_w1962_
	);
	LUT4 #(
		.INIT('h3222)
	) name1034 (
		\sub1_data_reg_reg[43]/NET0131 ,
		_w1053_,
		_w1670_,
		_w1769_,
		_w1963_
	);
	LUT4 #(
		.INIT('h53ff)
	) name1035 (
		\sub1_data_reg_reg[107]/NET0131 ,
		\sub1_data_reg_reg[43]/NET0131 ,
		\sub1_state_reg[4]/NET0131 ,
		_w1053_,
		_w1964_
	);
	LUT4 #(
		.INIT('hd0ff)
	) name1036 (
		_w1777_,
		_w1809_,
		_w1963_,
		_w1964_,
		_w1965_
	);
	LUT4 #(
		.INIT('h3222)
	) name1037 (
		\sub1_data_reg_reg[44]/NET0131 ,
		_w1053_,
		_w1670_,
		_w1769_,
		_w1966_
	);
	LUT4 #(
		.INIT('h7d00)
	) name1038 (
		_w1777_,
		_w1814_,
		_w1816_,
		_w1966_,
		_w1967_
	);
	LUT4 #(
		.INIT('h53ff)
	) name1039 (
		\sub1_data_reg_reg[108]/NET0131 ,
		\sub1_data_reg_reg[44]/NET0131 ,
		\sub1_state_reg[4]/NET0131 ,
		_w1053_,
		_w1968_
	);
	LUT2 #(
		.INIT('hb)
	) name1040 (
		_w1967_,
		_w1968_,
		_w1969_
	);
	LUT4 #(
		.INIT('h3222)
	) name1041 (
		\sub1_data_reg_reg[47]/NET0131 ,
		_w1053_,
		_w1670_,
		_w1769_,
		_w1970_
	);
	LUT4 #(
		.INIT('hb700)
	) name1042 (
		_w1639_,
		_w1777_,
		_w1794_,
		_w1970_,
		_w1971_
	);
	LUT4 #(
		.INIT('h53ff)
	) name1043 (
		\sub1_data_reg_reg[111]/NET0131 ,
		\sub1_data_reg_reg[47]/NET0131 ,
		\sub1_state_reg[4]/NET0131 ,
		_w1053_,
		_w1972_
	);
	LUT2 #(
		.INIT('hb)
	) name1044 (
		_w1971_,
		_w1972_,
		_w1973_
	);
	LUT4 #(
		.INIT('h3222)
	) name1045 (
		\sub1_data_reg_reg[72]/NET0131 ,
		_w1053_,
		_w1736_,
		_w1761_,
		_w1974_
	);
	LUT4 #(
		.INIT('h6f00)
	) name1046 (
		_w1631_,
		_w1640_,
		_w1784_,
		_w1974_,
		_w1975_
	);
	LUT4 #(
		.INIT('h35ff)
	) name1047 (
		\sub1_data_reg_reg[72]/NET0131 ,
		\sub1_data_reg_reg[8]/NET0131 ,
		\sub1_state_reg[4]/NET0131 ,
		_w1053_,
		_w1976_
	);
	LUT2 #(
		.INIT('hb)
	) name1048 (
		_w1975_,
		_w1976_,
		_w1977_
	);
	LUT4 #(
		.INIT('h3222)
	) name1049 (
		\sub1_data_reg_reg[75]/NET0131 ,
		_w1053_,
		_w1736_,
		_w1761_,
		_w1978_
	);
	LUT4 #(
		.INIT('h53ff)
	) name1050 (
		\sub1_data_reg_reg[11]/NET0131 ,
		\sub1_data_reg_reg[75]/NET0131 ,
		\sub1_state_reg[4]/NET0131 ,
		_w1053_,
		_w1979_
	);
	LUT4 #(
		.INIT('hd0ff)
	) name1051 (
		_w1784_,
		_w1809_,
		_w1978_,
		_w1979_,
		_w1980_
	);
	LUT4 #(
		.INIT('h3222)
	) name1052 (
		\sub1_data_reg_reg[76]/NET0131 ,
		_w1053_,
		_w1736_,
		_w1761_,
		_w1981_
	);
	LUT4 #(
		.INIT('h7d00)
	) name1053 (
		_w1784_,
		_w1814_,
		_w1816_,
		_w1981_,
		_w1982_
	);
	LUT4 #(
		.INIT('h53ff)
	) name1054 (
		\sub1_data_reg_reg[12]/NET0131 ,
		\sub1_data_reg_reg[76]/NET0131 ,
		\sub1_state_reg[4]/NET0131 ,
		_w1053_,
		_w1983_
	);
	LUT2 #(
		.INIT('hb)
	) name1055 (
		_w1982_,
		_w1983_,
		_w1984_
	);
	LUT4 #(
		.INIT('h3222)
	) name1056 (
		\sub1_data_reg_reg[79]/NET0131 ,
		_w1053_,
		_w1736_,
		_w1761_,
		_w1985_
	);
	LUT4 #(
		.INIT('hb700)
	) name1057 (
		_w1639_,
		_w1784_,
		_w1794_,
		_w1985_,
		_w1986_
	);
	LUT4 #(
		.INIT('h53ff)
	) name1058 (
		\sub1_data_reg_reg[15]/NET0131 ,
		\sub1_data_reg_reg[79]/NET0131 ,
		\sub1_state_reg[4]/NET0131 ,
		_w1053_,
		_w1987_
	);
	LUT2 #(
		.INIT('hb)
	) name1059 (
		_w1986_,
		_w1987_,
		_w1988_
	);
	LUT4 #(
		.INIT('h3222)
	) name1060 (
		\sub1_data_reg_reg[8]/NET0131 ,
		_w1053_,
		_w1736_,
		_w1769_,
		_w1989_
	);
	LUT4 #(
		.INIT('h6f00)
	) name1061 (
		_w1631_,
		_w1640_,
		_w1770_,
		_w1989_,
		_w1990_
	);
	LUT4 #(
		.INIT('h53ff)
	) name1062 (
		\sub1_data_reg_reg[72]/NET0131 ,
		\sub1_data_reg_reg[8]/NET0131 ,
		\sub1_state_reg[4]/NET0131 ,
		_w1053_,
		_w1991_
	);
	LUT2 #(
		.INIT('hb)
	) name1063 (
		_w1990_,
		_w1991_,
		_w1992_
	);
	LUT4 #(
		.INIT('h1455)
	) name1064 (
		_w1053_,
		_w1631_,
		_w1640_,
		_w1713_,
		_w1993_
	);
	LUT3 #(
		.INIT('ha8)
	) name1065 (
		\sub1_data_reg_reg[32]/NET0131 ,
		_w1060_,
		_w1993_,
		_w1994_
	);
	LUT4 #(
		.INIT('h1400)
	) name1066 (
		_w1053_,
		_w1631_,
		_w1640_,
		_w1713_,
		_w1995_
	);
	LUT2 #(
		.INIT('h1)
	) name1067 (
		decrypt_i_pad,
		\sub1_data_reg_reg[64]/NET0131 ,
		_w1996_
	);
	LUT3 #(
		.INIT('h08)
	) name1068 (
		\sub1_state_reg[4]/NET0131 ,
		_w1053_,
		_w1996_,
		_w1997_
	);
	LUT4 #(
		.INIT('h7d00)
	) name1069 (
		decrypt_i_pad,
		_w1631_,
		_w1640_,
		_w1997_,
		_w1998_
	);
	LUT2 #(
		.INIT('h1)
	) name1070 (
		_w1995_,
		_w1998_,
		_w1999_
	);
	LUT2 #(
		.INIT('hb)
	) name1071 (
		_w1994_,
		_w1999_,
		_w2000_
	);
	LUT4 #(
		.INIT('h88b8)
	) name1072 (
		\sub1_state_reg[4]/NET0131 ,
		_w1053_,
		_w1713_,
		_w1809_,
		_w2001_
	);
	LUT3 #(
		.INIT('h40)
	) name1073 (
		_w1053_,
		_w1713_,
		_w1809_,
		_w2002_
	);
	LUT2 #(
		.INIT('h1)
	) name1074 (
		decrypt_i_pad,
		\sub1_data_reg_reg[67]/NET0131 ,
		_w2003_
	);
	LUT3 #(
		.INIT('h08)
	) name1075 (
		\sub1_state_reg[4]/NET0131 ,
		_w1053_,
		_w2003_,
		_w2004_
	);
	LUT3 #(
		.INIT('hd0)
	) name1076 (
		decrypt_i_pad,
		_w1809_,
		_w2004_,
		_w2005_
	);
	LUT4 #(
		.INIT('hffce)
	) name1077 (
		\sub1_data_reg_reg[35]/NET0131 ,
		_w2002_,
		_w2001_,
		_w2005_,
		_w2006_
	);
	LUT4 #(
		.INIT('h4515)
	) name1078 (
		_w1053_,
		_w1639_,
		_w1713_,
		_w1794_,
		_w2007_
	);
	LUT3 #(
		.INIT('ha8)
	) name1079 (
		\sub1_data_reg_reg[39]/NET0131 ,
		_w1060_,
		_w2007_,
		_w2008_
	);
	LUT4 #(
		.INIT('h4010)
	) name1080 (
		_w1053_,
		_w1639_,
		_w1713_,
		_w1794_,
		_w2009_
	);
	LUT2 #(
		.INIT('h1)
	) name1081 (
		decrypt_i_pad,
		\sub1_data_reg_reg[71]/NET0131 ,
		_w2010_
	);
	LUT3 #(
		.INIT('h08)
	) name1082 (
		\sub1_state_reg[4]/NET0131 ,
		_w1053_,
		_w2010_,
		_w2011_
	);
	LUT4 #(
		.INIT('hd700)
	) name1083 (
		decrypt_i_pad,
		_w1639_,
		_w1794_,
		_w2011_,
		_w2012_
	);
	LUT2 #(
		.INIT('h1)
	) name1084 (
		_w2009_,
		_w2012_,
		_w2013_
	);
	LUT2 #(
		.INIT('hb)
	) name1085 (
		_w2008_,
		_w2013_,
		_w2014_
	);
	LUT4 #(
		.INIT('h1551)
	) name1086 (
		_w1053_,
		_w1672_,
		_w1814_,
		_w1816_,
		_w2015_
	);
	LUT3 #(
		.INIT('ha8)
	) name1087 (
		\sub1_data_reg_reg[100]/NET0131 ,
		_w1060_,
		_w2015_,
		_w2016_
	);
	LUT4 #(
		.INIT('h0440)
	) name1088 (
		_w1053_,
		_w1672_,
		_w1814_,
		_w1816_,
		_w2017_
	);
	LUT2 #(
		.INIT('h2)
	) name1089 (
		decrypt_i_pad,
		\sub1_data_reg_reg[68]/NET0131 ,
		_w2018_
	);
	LUT3 #(
		.INIT('h08)
	) name1090 (
		\sub1_state_reg[4]/NET0131 ,
		_w1053_,
		_w2018_,
		_w2019_
	);
	LUT4 #(
		.INIT('hbe00)
	) name1091 (
		decrypt_i_pad,
		_w1814_,
		_w1816_,
		_w2019_,
		_w2020_
	);
	LUT2 #(
		.INIT('h1)
	) name1092 (
		_w2017_,
		_w2020_,
		_w2021_
	);
	LUT2 #(
		.INIT('hb)
	) name1093 (
		_w2016_,
		_w2021_,
		_w2022_
	);
	LUT4 #(
		.INIT('h88b8)
	) name1094 (
		\sub1_state_reg[4]/NET0131 ,
		_w1053_,
		_w1672_,
		_w1809_,
		_w2023_
	);
	LUT2 #(
		.INIT('h2)
	) name1095 (
		decrypt_i_pad,
		\sub1_data_reg_reg[67]/NET0131 ,
		_w2024_
	);
	LUT3 #(
		.INIT('h08)
	) name1096 (
		\sub1_state_reg[4]/NET0131 ,
		_w1053_,
		_w2024_,
		_w2025_
	);
	LUT4 #(
		.INIT('hbe00)
	) name1097 (
		decrypt_i_pad,
		_w970_,
		_w1808_,
		_w2025_,
		_w2026_
	);
	LUT4 #(
		.INIT('h00bf)
	) name1098 (
		_w1053_,
		_w1672_,
		_w1809_,
		_w2026_,
		_w2027_
	);
	LUT3 #(
		.INIT('h2f)
	) name1099 (
		\sub1_data_reg_reg[99]/NET0131 ,
		_w2023_,
		_w2027_,
		_w2028_
	);
	LUT2 #(
		.INIT('h8)
	) name1100 (
		_w1692_,
		_w1761_,
		_w2029_
	);
	LUT3 #(
		.INIT('hca)
	) name1101 (
		\sub1_data_reg_reg[125]/NET0131 ,
		_w1683_,
		_w2029_,
		_w2030_
	);
	LUT3 #(
		.INIT('h3a)
	) name1102 (
		\sub1_data_reg_reg[126]/NET0131 ,
		_w985_,
		_w2029_,
		_w2031_
	);
	LUT2 #(
		.INIT('h8)
	) name1103 (
		_w1702_,
		_w1769_,
		_w2032_
	);
	LUT3 #(
		.INIT('hca)
	) name1104 (
		\sub1_data_reg_reg[29]/NET0131 ,
		_w1683_,
		_w2032_,
		_w2033_
	);
	LUT3 #(
		.INIT('h3a)
	) name1105 (
		\sub1_data_reg_reg[30]/NET0131 ,
		_w985_,
		_w2032_,
		_w2034_
	);
	LUT2 #(
		.INIT('h8)
	) name1106 (
		_w1692_,
		_w1769_,
		_w2035_
	);
	LUT3 #(
		.INIT('hca)
	) name1107 (
		\sub1_data_reg_reg[61]/NET0131 ,
		_w1683_,
		_w2035_,
		_w2036_
	);
	LUT3 #(
		.INIT('h3a)
	) name1108 (
		\sub1_data_reg_reg[62]/NET0131 ,
		_w985_,
		_w2035_,
		_w2037_
	);
	LUT2 #(
		.INIT('h8)
	) name1109 (
		_w1702_,
		_w1761_,
		_w2038_
	);
	LUT3 #(
		.INIT('hca)
	) name1110 (
		\sub1_data_reg_reg[93]/NET0131 ,
		_w1683_,
		_w2038_,
		_w2039_
	);
	LUT3 #(
		.INIT('h3a)
	) name1111 (
		\sub1_data_reg_reg[94]/NET0131 ,
		_w985_,
		_w2038_,
		_w2040_
	);
	LUT4 #(
		.INIT('h5553)
	) name1112 (
		\key_i[73]_pad ,
		\ks1_key_reg_reg[73]/NET0131 ,
		_w938_,
		_w986_,
		_w2041_
	);
	LUT2 #(
		.INIT('h2)
	) name1113 (
		_w951_,
		_w1658_,
		_w2042_
	);
	LUT4 #(
		.INIT('h1441)
	) name1114 (
		_w951_,
		_w1632_,
		_w1638_,
		_w1808_,
		_w2043_
	);
	LUT4 #(
		.INIT('haaac)
	) name1115 (
		\key_i[105]_pad ,
		\ks1_key_reg_reg[105]/NET0131 ,
		_w938_,
		_w986_,
		_w2044_
	);
	LUT3 #(
		.INIT('h1e)
	) name1116 (
		_w2042_,
		_w2043_,
		_w2044_,
		_w2045_
	);
	LUT4 #(
		.INIT('ha956)
	) name1117 (
		_w2041_,
		_w2042_,
		_w2043_,
		_w2044_,
		_w2046_
	);
	LUT3 #(
		.INIT('h2e)
	) name1118 (
		\ks1_key_reg_reg[73]/NET0131 ,
		_w929_,
		_w2046_,
		_w2047_
	);
	LUT4 #(
		.INIT('h2ee2)
	) name1119 (
		\ks1_key_reg_reg[74]/NET0131 ,
		_w929_,
		_w1650_,
		_w1662_,
		_w2048_
	);
	LUT4 #(
		.INIT('h3222)
	) name1120 (
		\sub1_data_reg_reg[113]/NET0131 ,
		_w1053_,
		_w1671_,
		_w1692_,
		_w2049_
	);
	LUT4 #(
		.INIT('hfd00)
	) name1121 (
		_w1693_,
		_w2042_,
		_w2043_,
		_w2049_,
		_w2050_
	);
	LUT3 #(
		.INIT('hd8)
	) name1122 (
		decrypt_i_pad,
		\sub1_data_reg_reg[17]/NET0131 ,
		\sub1_data_reg_reg[81]/NET0131 ,
		_w2051_
	);
	LUT4 #(
		.INIT('h1fdf)
	) name1123 (
		\sub1_data_reg_reg[113]/NET0131 ,
		\sub1_state_reg[4]/NET0131 ,
		_w1053_,
		_w2051_,
		_w2052_
	);
	LUT2 #(
		.INIT('hb)
	) name1124 (
		_w2050_,
		_w2052_,
		_w2053_
	);
	LUT4 #(
		.INIT('ha900)
	) name1125 (
		_w1657_,
		_w1659_,
		_w1660_,
		_w1693_,
		_w2054_
	);
	LUT4 #(
		.INIT('h3222)
	) name1126 (
		\sub1_data_reg_reg[114]/NET0131 ,
		_w1053_,
		_w1671_,
		_w1692_,
		_w2055_
	);
	LUT3 #(
		.INIT('hd8)
	) name1127 (
		decrypt_i_pad,
		\sub1_data_reg_reg[18]/NET0131 ,
		\sub1_data_reg_reg[82]/NET0131 ,
		_w2056_
	);
	LUT4 #(
		.INIT('h1fdf)
	) name1128 (
		\sub1_data_reg_reg[114]/NET0131 ,
		\sub1_state_reg[4]/NET0131 ,
		_w1053_,
		_w2056_,
		_w2057_
	);
	LUT3 #(
		.INIT('h4f)
	) name1129 (
		_w2054_,
		_w2055_,
		_w2057_,
		_w2058_
	);
	LUT4 #(
		.INIT('h3222)
	) name1130 (
		\sub1_data_reg_reg[17]/NET0131 ,
		_w1053_,
		_w1702_,
		_w1703_,
		_w2059_
	);
	LUT4 #(
		.INIT('hfd00)
	) name1131 (
		_w1704_,
		_w2042_,
		_w2043_,
		_w2059_,
		_w2060_
	);
	LUT3 #(
		.INIT('he4)
	) name1132 (
		decrypt_i_pad,
		\sub1_data_reg_reg[113]/NET0131 ,
		\sub1_data_reg_reg[49]/NET0131 ,
		_w2061_
	);
	LUT4 #(
		.INIT('h1fdf)
	) name1133 (
		\sub1_data_reg_reg[17]/NET0131 ,
		\sub1_state_reg[4]/NET0131 ,
		_w1053_,
		_w2061_,
		_w2062_
	);
	LUT2 #(
		.INIT('hb)
	) name1134 (
		_w2060_,
		_w2062_,
		_w2063_
	);
	LUT4 #(
		.INIT('ha900)
	) name1135 (
		_w1657_,
		_w1659_,
		_w1660_,
		_w1704_,
		_w2064_
	);
	LUT4 #(
		.INIT('h3222)
	) name1136 (
		\sub1_data_reg_reg[18]/NET0131 ,
		_w1053_,
		_w1702_,
		_w1703_,
		_w2065_
	);
	LUT3 #(
		.INIT('he4)
	) name1137 (
		decrypt_i_pad,
		\sub1_data_reg_reg[114]/NET0131 ,
		\sub1_data_reg_reg[50]/NET0131 ,
		_w2066_
	);
	LUT4 #(
		.INIT('h1fdf)
	) name1138 (
		\sub1_data_reg_reg[18]/NET0131 ,
		\sub1_state_reg[4]/NET0131 ,
		_w1053_,
		_w2066_,
		_w2067_
	);
	LUT3 #(
		.INIT('h4f)
	) name1139 (
		_w2064_,
		_w2065_,
		_w2067_,
		_w2068_
	);
	LUT3 #(
		.INIT('h1b)
	) name1140 (
		decrypt_i_pad,
		\sub1_data_reg_reg[33]/NET0131 ,
		\sub1_data_reg_reg[97]/NET0131 ,
		_w2069_
	);
	LUT4 #(
		.INIT('h2aea)
	) name1141 (
		\sub1_data_reg_reg[1]/NET0131 ,
		\sub1_state_reg[4]/NET0131 ,
		_w1053_,
		_w2069_,
		_w2070_
	);
	LUT3 #(
		.INIT('he4)
	) name1142 (
		decrypt_i_pad,
		\sub1_data_reg_reg[34]/NET0131 ,
		\sub1_data_reg_reg[98]/NET0131 ,
		_w2071_
	);
	LUT3 #(
		.INIT('h80)
	) name1143 (
		\sub1_state_reg[4]/NET0131 ,
		_w1053_,
		_w2071_,
		_w2072_
	);
	LUT4 #(
		.INIT('hff2a)
	) name1144 (
		\sub1_data_reg_reg[2]/NET0131 ,
		_w1703_,
		_w1736_,
		_w2072_,
		_w2073_
	);
	LUT4 #(
		.INIT('h3222)
	) name1145 (
		\sub1_data_reg_reg[49]/NET0131 ,
		_w1053_,
		_w1692_,
		_w1703_,
		_w2074_
	);
	LUT4 #(
		.INIT('hfd00)
	) name1146 (
		_w1727_,
		_w2042_,
		_w2043_,
		_w2074_,
		_w2075_
	);
	LUT3 #(
		.INIT('he4)
	) name1147 (
		decrypt_i_pad,
		\sub1_data_reg_reg[17]/NET0131 ,
		\sub1_data_reg_reg[81]/NET0131 ,
		_w2076_
	);
	LUT4 #(
		.INIT('h1fdf)
	) name1148 (
		\sub1_data_reg_reg[49]/NET0131 ,
		\sub1_state_reg[4]/NET0131 ,
		_w1053_,
		_w2076_,
		_w2077_
	);
	LUT2 #(
		.INIT('hb)
	) name1149 (
		_w2075_,
		_w2077_,
		_w2078_
	);
	LUT4 #(
		.INIT('ha900)
	) name1150 (
		_w1657_,
		_w1659_,
		_w1660_,
		_w1727_,
		_w2079_
	);
	LUT4 #(
		.INIT('h3222)
	) name1151 (
		\sub1_data_reg_reg[50]/NET0131 ,
		_w1053_,
		_w1692_,
		_w1703_,
		_w2080_
	);
	LUT3 #(
		.INIT('he4)
	) name1152 (
		decrypt_i_pad,
		\sub1_data_reg_reg[18]/NET0131 ,
		\sub1_data_reg_reg[82]/NET0131 ,
		_w2081_
	);
	LUT4 #(
		.INIT('h1fdf)
	) name1153 (
		\sub1_data_reg_reg[50]/NET0131 ,
		\sub1_state_reg[4]/NET0131 ,
		_w1053_,
		_w2081_,
		_w2082_
	);
	LUT3 #(
		.INIT('h4f)
	) name1154 (
		_w2079_,
		_w2080_,
		_w2082_,
		_w2083_
	);
	LUT4 #(
		.INIT('h3222)
	) name1155 (
		\sub1_data_reg_reg[65]/NET0131 ,
		_w1053_,
		_w1671_,
		_w1736_,
		_w2084_
	);
	LUT4 #(
		.INIT('hfd00)
	) name1156 (
		_w1743_,
		_w2042_,
		_w2043_,
		_w2084_,
		_w2085_
	);
	LUT3 #(
		.INIT('hd8)
	) name1157 (
		decrypt_i_pad,
		\sub1_data_reg_reg[33]/NET0131 ,
		\sub1_data_reg_reg[97]/NET0131 ,
		_w2086_
	);
	LUT4 #(
		.INIT('h1fdf)
	) name1158 (
		\sub1_data_reg_reg[65]/NET0131 ,
		\sub1_state_reg[4]/NET0131 ,
		_w1053_,
		_w2086_,
		_w2087_
	);
	LUT2 #(
		.INIT('hb)
	) name1159 (
		_w2085_,
		_w2087_,
		_w2088_
	);
	LUT4 #(
		.INIT('ha900)
	) name1160 (
		_w1657_,
		_w1659_,
		_w1660_,
		_w1743_,
		_w2089_
	);
	LUT4 #(
		.INIT('h3222)
	) name1161 (
		\sub1_data_reg_reg[66]/NET0131 ,
		_w1053_,
		_w1671_,
		_w1736_,
		_w2090_
	);
	LUT3 #(
		.INIT('hd8)
	) name1162 (
		decrypt_i_pad,
		\sub1_data_reg_reg[34]/NET0131 ,
		\sub1_data_reg_reg[98]/NET0131 ,
		_w2091_
	);
	LUT4 #(
		.INIT('h1fdf)
	) name1163 (
		\sub1_data_reg_reg[66]/NET0131 ,
		\sub1_state_reg[4]/NET0131 ,
		_w1053_,
		_w2091_,
		_w2092_
	);
	LUT3 #(
		.INIT('h4f)
	) name1164 (
		_w2089_,
		_w2090_,
		_w2092_,
		_w2093_
	);
	LUT4 #(
		.INIT('h3222)
	) name1165 (
		\sub1_data_reg_reg[81]/NET0131 ,
		_w1053_,
		_w1671_,
		_w1702_,
		_w2094_
	);
	LUT4 #(
		.INIT('hfd00)
	) name1166 (
		_w1752_,
		_w2042_,
		_w2043_,
		_w2094_,
		_w2095_
	);
	LUT3 #(
		.INIT('hd8)
	) name1167 (
		decrypt_i_pad,
		\sub1_data_reg_reg[113]/NET0131 ,
		\sub1_data_reg_reg[49]/NET0131 ,
		_w2096_
	);
	LUT4 #(
		.INIT('h1fdf)
	) name1168 (
		\sub1_data_reg_reg[81]/NET0131 ,
		\sub1_state_reg[4]/NET0131 ,
		_w1053_,
		_w2096_,
		_w2097_
	);
	LUT2 #(
		.INIT('hb)
	) name1169 (
		_w2095_,
		_w2097_,
		_w2098_
	);
	LUT4 #(
		.INIT('ha900)
	) name1170 (
		_w1657_,
		_w1659_,
		_w1660_,
		_w1752_,
		_w2099_
	);
	LUT4 #(
		.INIT('h3222)
	) name1171 (
		\sub1_data_reg_reg[82]/NET0131 ,
		_w1053_,
		_w1671_,
		_w1702_,
		_w2100_
	);
	LUT3 #(
		.INIT('hd8)
	) name1172 (
		decrypt_i_pad,
		\sub1_data_reg_reg[114]/NET0131 ,
		\sub1_data_reg_reg[50]/NET0131 ,
		_w2101_
	);
	LUT4 #(
		.INIT('h1fdf)
	) name1173 (
		\sub1_data_reg_reg[82]/NET0131 ,
		\sub1_state_reg[4]/NET0131 ,
		_w1053_,
		_w2101_,
		_w2102_
	);
	LUT3 #(
		.INIT('h4f)
	) name1174 (
		_w2099_,
		_w2100_,
		_w2102_,
		_w2103_
	);
	LUT4 #(
		.INIT('h3222)
	) name1175 (
		\sub1_data_reg_reg[97]/NET0131 ,
		_w1053_,
		_w1670_,
		_w1671_,
		_w2104_
	);
	LUT4 #(
		.INIT('hfd00)
	) name1176 (
		_w1672_,
		_w2042_,
		_w2043_,
		_w2104_,
		_w2105_
	);
	LUT3 #(
		.INIT('h20)
	) name1177 (
		\sub1_data_reg_reg[97]/NET0131 ,
		\sub1_state_reg[4]/NET0131 ,
		_w1053_,
		_w2106_
	);
	LUT4 #(
		.INIT('h4114)
	) name1178 (
		decrypt_i_pad,
		_w1632_,
		_w1638_,
		_w1808_,
		_w2107_
	);
	LUT2 #(
		.INIT('h2)
	) name1179 (
		decrypt_i_pad,
		\sub1_data_reg_reg[65]/NET0131 ,
		_w2108_
	);
	LUT3 #(
		.INIT('h08)
	) name1180 (
		\sub1_state_reg[4]/NET0131 ,
		_w1053_,
		_w2108_,
		_w2109_
	);
	LUT3 #(
		.INIT('h45)
	) name1181 (
		_w2106_,
		_w2107_,
		_w2109_,
		_w2110_
	);
	LUT2 #(
		.INIT('hb)
	) name1182 (
		_w2105_,
		_w2110_,
		_w2111_
	);
	LUT4 #(
		.INIT('ha900)
	) name1183 (
		_w1657_,
		_w1659_,
		_w1660_,
		_w1672_,
		_w2112_
	);
	LUT4 #(
		.INIT('h202a)
	) name1184 (
		\sub1_data_reg_reg[98]/NET0131 ,
		\sub1_state_reg[4]/NET0131 ,
		_w1053_,
		_w2112_,
		_w2113_
	);
	LUT3 #(
		.INIT('h40)
	) name1185 (
		_w1053_,
		_w1661_,
		_w1672_,
		_w2114_
	);
	LUT4 #(
		.INIT('h4441)
	) name1186 (
		decrypt_i_pad,
		_w1657_,
		_w1659_,
		_w1660_,
		_w2115_
	);
	LUT2 #(
		.INIT('h2)
	) name1187 (
		decrypt_i_pad,
		\sub1_data_reg_reg[66]/NET0131 ,
		_w2116_
	);
	LUT3 #(
		.INIT('h08)
	) name1188 (
		\sub1_state_reg[4]/NET0131 ,
		_w1053_,
		_w2116_,
		_w2117_
	);
	LUT2 #(
		.INIT('h4)
	) name1189 (
		_w2115_,
		_w2117_,
		_w2118_
	);
	LUT3 #(
		.INIT('hfe)
	) name1190 (
		_w2114_,
		_w2113_,
		_w2118_,
		_w2119_
	);
	LUT4 #(
		.INIT('h3222)
	) name1191 (
		\sub1_data_reg_reg[105]/NET0131 ,
		_w1053_,
		_w1670_,
		_w1761_,
		_w2120_
	);
	LUT4 #(
		.INIT('hfd00)
	) name1192 (
		_w1762_,
		_w2042_,
		_w2043_,
		_w2120_,
		_w2121_
	);
	LUT4 #(
		.INIT('h35ff)
	) name1193 (
		\sub1_data_reg_reg[105]/NET0131 ,
		\sub1_data_reg_reg[41]/NET0131 ,
		\sub1_state_reg[4]/NET0131 ,
		_w1053_,
		_w2122_
	);
	LUT2 #(
		.INIT('hb)
	) name1194 (
		_w2121_,
		_w2122_,
		_w2123_
	);
	LUT4 #(
		.INIT('ha900)
	) name1195 (
		_w1657_,
		_w1659_,
		_w1660_,
		_w1762_,
		_w2124_
	);
	LUT4 #(
		.INIT('h3222)
	) name1196 (
		\sub1_data_reg_reg[106]/NET0131 ,
		_w1053_,
		_w1670_,
		_w1761_,
		_w2125_
	);
	LUT4 #(
		.INIT('h35ff)
	) name1197 (
		\sub1_data_reg_reg[106]/NET0131 ,
		\sub1_data_reg_reg[42]/NET0131 ,
		\sub1_state_reg[4]/NET0131 ,
		_w1053_,
		_w2126_
	);
	LUT3 #(
		.INIT('h4f)
	) name1198 (
		_w2124_,
		_w2125_,
		_w2126_,
		_w2127_
	);
	LUT4 #(
		.INIT('h2ee2)
	) name1199 (
		\ks1_col_reg[0]/NET0131 ,
		_w1079_,
		_w1631_,
		_w1640_,
		_w2128_
	);
	LUT3 #(
		.INIT('he2)
	) name1200 (
		\ks1_col_reg[19]/NET0131 ,
		_w1064_,
		_w1809_,
		_w2129_
	);
	LUT4 #(
		.INIT('h2ee2)
	) name1201 (
		\ks1_col_reg[16]/NET0131 ,
		_w1064_,
		_w1631_,
		_w1640_,
		_w2130_
	);
	LUT4 #(
		.INIT('h2ee2)
	) name1202 (
		\ks1_col_reg[20]/NET0131 ,
		_w1064_,
		_w1814_,
		_w1816_,
		_w2131_
	);
	LUT4 #(
		.INIT('ha900)
	) name1203 (
		_w1657_,
		_w1659_,
		_w1660_,
		_w1770_,
		_w2132_
	);
	LUT4 #(
		.INIT('h3222)
	) name1204 (
		\sub1_data_reg_reg[10]/NET0131 ,
		_w1053_,
		_w1736_,
		_w1769_,
		_w2133_
	);
	LUT4 #(
		.INIT('h35ff)
	) name1205 (
		\sub1_data_reg_reg[10]/NET0131 ,
		\sub1_data_reg_reg[74]/NET0131 ,
		\sub1_state_reg[4]/NET0131 ,
		_w1053_,
		_w2134_
	);
	LUT3 #(
		.INIT('h4f)
	) name1206 (
		_w2132_,
		_w2133_,
		_w2134_,
		_w2135_
	);
	LUT4 #(
		.INIT('he22e)
	) name1207 (
		\ks1_col_reg[23]/NET0131 ,
		_w1064_,
		_w1639_,
		_w1794_,
		_w2136_
	);
	LUT4 #(
		.INIT('h2ee2)
	) name1208 (
		\ks1_col_reg[24]/NET0131 ,
		_w1071_,
		_w1631_,
		_w1640_,
		_w2137_
	);
	LUT3 #(
		.INIT('he2)
	) name1209 (
		\ks1_col_reg[27]/NET0131 ,
		_w1071_,
		_w1809_,
		_w2138_
	);
	LUT4 #(
		.INIT('h2ee2)
	) name1210 (
		\ks1_col_reg[28]/NET0131 ,
		_w1071_,
		_w1814_,
		_w1816_,
		_w2139_
	);
	LUT4 #(
		.INIT('he22e)
	) name1211 (
		\ks1_col_reg[31]/NET0131 ,
		_w1071_,
		_w1639_,
		_w1794_,
		_w2140_
	);
	LUT3 #(
		.INIT('he2)
	) name1212 (
		\ks1_col_reg[3]/NET0131 ,
		_w1079_,
		_w1809_,
		_w2141_
	);
	LUT4 #(
		.INIT('h2ee2)
	) name1213 (
		\ks1_col_reg[4]/NET0131 ,
		_w1079_,
		_w1814_,
		_w1816_,
		_w2142_
	);
	LUT4 #(
		.INIT('he22e)
	) name1214 (
		\ks1_col_reg[7]/NET0131 ,
		_w1079_,
		_w1639_,
		_w1794_,
		_w2143_
	);
	LUT4 #(
		.INIT('h3222)
	) name1215 (
		\sub1_data_reg_reg[41]/NET0131 ,
		_w1053_,
		_w1670_,
		_w1769_,
		_w2144_
	);
	LUT4 #(
		.INIT('hfd00)
	) name1216 (
		_w1777_,
		_w2042_,
		_w2043_,
		_w2144_,
		_w2145_
	);
	LUT4 #(
		.INIT('h53ff)
	) name1217 (
		\sub1_data_reg_reg[105]/NET0131 ,
		\sub1_data_reg_reg[41]/NET0131 ,
		\sub1_state_reg[4]/NET0131 ,
		_w1053_,
		_w2146_
	);
	LUT2 #(
		.INIT('hb)
	) name1218 (
		_w2145_,
		_w2146_,
		_w2147_
	);
	LUT4 #(
		.INIT('ha900)
	) name1219 (
		_w1657_,
		_w1659_,
		_w1660_,
		_w1777_,
		_w2148_
	);
	LUT4 #(
		.INIT('h3222)
	) name1220 (
		\sub1_data_reg_reg[42]/NET0131 ,
		_w1053_,
		_w1670_,
		_w1769_,
		_w2149_
	);
	LUT4 #(
		.INIT('h53ff)
	) name1221 (
		\sub1_data_reg_reg[106]/NET0131 ,
		\sub1_data_reg_reg[42]/NET0131 ,
		\sub1_state_reg[4]/NET0131 ,
		_w1053_,
		_w2150_
	);
	LUT3 #(
		.INIT('h4f)
	) name1222 (
		_w2148_,
		_w2149_,
		_w2150_,
		_w2151_
	);
	LUT4 #(
		.INIT('h3222)
	) name1223 (
		\sub1_data_reg_reg[73]/NET0131 ,
		_w1053_,
		_w1736_,
		_w1761_,
		_w2152_
	);
	LUT4 #(
		.INIT('hfd00)
	) name1224 (
		_w1784_,
		_w2042_,
		_w2043_,
		_w2152_,
		_w2153_
	);
	LUT4 #(
		.INIT('h35ff)
	) name1225 (
		\sub1_data_reg_reg[73]/NET0131 ,
		\sub1_data_reg_reg[9]/NET0131 ,
		\sub1_state_reg[4]/NET0131 ,
		_w1053_,
		_w2154_
	);
	LUT2 #(
		.INIT('hb)
	) name1226 (
		_w2153_,
		_w2154_,
		_w2155_
	);
	LUT4 #(
		.INIT('ha900)
	) name1227 (
		_w1657_,
		_w1659_,
		_w1660_,
		_w1784_,
		_w2156_
	);
	LUT4 #(
		.INIT('h3222)
	) name1228 (
		\sub1_data_reg_reg[74]/NET0131 ,
		_w1053_,
		_w1736_,
		_w1761_,
		_w2157_
	);
	LUT4 #(
		.INIT('h53ff)
	) name1229 (
		\sub1_data_reg_reg[10]/NET0131 ,
		\sub1_data_reg_reg[74]/NET0131 ,
		\sub1_state_reg[4]/NET0131 ,
		_w1053_,
		_w2158_
	);
	LUT3 #(
		.INIT('h4f)
	) name1230 (
		_w2156_,
		_w2157_,
		_w2158_,
		_w2159_
	);
	LUT4 #(
		.INIT('h3222)
	) name1231 (
		\sub1_data_reg_reg[9]/NET0131 ,
		_w1053_,
		_w1736_,
		_w1769_,
		_w2160_
	);
	LUT4 #(
		.INIT('hfd00)
	) name1232 (
		_w1770_,
		_w2042_,
		_w2043_,
		_w2160_,
		_w2161_
	);
	LUT4 #(
		.INIT('h53ff)
	) name1233 (
		\sub1_data_reg_reg[73]/NET0131 ,
		\sub1_data_reg_reg[9]/NET0131 ,
		\sub1_state_reg[4]/NET0131 ,
		_w1053_,
		_w2162_
	);
	LUT2 #(
		.INIT('hb)
	) name1234 (
		_w2161_,
		_w2162_,
		_w2163_
	);
	LUT4 #(
		.INIT('h5551)
	) name1235 (
		_w1053_,
		_w1713_,
		_w2042_,
		_w2043_,
		_w2164_
	);
	LUT3 #(
		.INIT('ha8)
	) name1236 (
		\sub1_data_reg_reg[33]/NET0131 ,
		_w1060_,
		_w2164_,
		_w2165_
	);
	LUT4 #(
		.INIT('h4440)
	) name1237 (
		_w1053_,
		_w1713_,
		_w2042_,
		_w2043_,
		_w2166_
	);
	LUT2 #(
		.INIT('h1)
	) name1238 (
		decrypt_i_pad,
		\sub1_data_reg_reg[65]/NET0131 ,
		_w2167_
	);
	LUT3 #(
		.INIT('h08)
	) name1239 (
		\sub1_state_reg[4]/NET0131 ,
		_w1053_,
		_w2167_,
		_w2168_
	);
	LUT4 #(
		.INIT('hfd00)
	) name1240 (
		decrypt_i_pad,
		_w2042_,
		_w2043_,
		_w2168_,
		_w2169_
	);
	LUT2 #(
		.INIT('h1)
	) name1241 (
		_w2166_,
		_w2169_,
		_w2170_
	);
	LUT2 #(
		.INIT('hb)
	) name1242 (
		_w2165_,
		_w2170_,
		_w2171_
	);
	LUT4 #(
		.INIT('ha900)
	) name1243 (
		_w1657_,
		_w1659_,
		_w1660_,
		_w1713_,
		_w2172_
	);
	LUT4 #(
		.INIT('h202a)
	) name1244 (
		\sub1_data_reg_reg[34]/NET0131 ,
		\sub1_state_reg[4]/NET0131 ,
		_w1053_,
		_w2172_,
		_w2173_
	);
	LUT3 #(
		.INIT('h40)
	) name1245 (
		_w1053_,
		_w1661_,
		_w1713_,
		_w2174_
	);
	LUT4 #(
		.INIT('h8882)
	) name1246 (
		decrypt_i_pad,
		_w1657_,
		_w1659_,
		_w1660_,
		_w2175_
	);
	LUT2 #(
		.INIT('h1)
	) name1247 (
		decrypt_i_pad,
		\sub1_data_reg_reg[66]/NET0131 ,
		_w2176_
	);
	LUT3 #(
		.INIT('h08)
	) name1248 (
		\sub1_state_reg[4]/NET0131 ,
		_w1053_,
		_w2176_,
		_w2177_
	);
	LUT2 #(
		.INIT('h4)
	) name1249 (
		_w2175_,
		_w2177_,
		_w2178_
	);
	LUT3 #(
		.INIT('hfe)
	) name1250 (
		_w2174_,
		_w2173_,
		_w2178_,
		_w2179_
	);
	LUT4 #(
		.INIT('h3caa)
	) name1251 (
		\sub1_data_reg_reg[120]/NET0131 ,
		_w1631_,
		_w1640_,
		_w2029_,
		_w2180_
	);
	LUT4 #(
		.INIT('h3caa)
	) name1252 (
		\sub1_data_reg_reg[24]/NET0131 ,
		_w1631_,
		_w1640_,
		_w2032_,
		_w2181_
	);
	LUT4 #(
		.INIT('h3caa)
	) name1253 (
		\sub1_data_reg_reg[56]/NET0131 ,
		_w1631_,
		_w1640_,
		_w2035_,
		_w2182_
	);
	LUT4 #(
		.INIT('h3caa)
	) name1254 (
		\sub1_data_reg_reg[88]/NET0131 ,
		_w1631_,
		_w1640_,
		_w2038_,
		_w2183_
	);
	LUT3 #(
		.INIT('hca)
	) name1255 (
		\sub1_data_reg_reg[123]/NET0131 ,
		_w1809_,
		_w2029_,
		_w2184_
	);
	LUT4 #(
		.INIT('h3caa)
	) name1256 (
		\sub1_data_reg_reg[124]/NET0131 ,
		_w1814_,
		_w1816_,
		_w2029_,
		_w2185_
	);
	LUT4 #(
		.INIT('hc3aa)
	) name1257 (
		\sub1_data_reg_reg[127]/NET0131 ,
		_w1639_,
		_w1794_,
		_w2029_,
		_w2186_
	);
	LUT3 #(
		.INIT('hca)
	) name1258 (
		\sub1_data_reg_reg[27]/NET0131 ,
		_w1809_,
		_w2032_,
		_w2187_
	);
	LUT4 #(
		.INIT('h3caa)
	) name1259 (
		\sub1_data_reg_reg[28]/NET0131 ,
		_w1814_,
		_w1816_,
		_w2032_,
		_w2188_
	);
	LUT4 #(
		.INIT('hc3aa)
	) name1260 (
		\sub1_data_reg_reg[31]/NET0131 ,
		_w1639_,
		_w1794_,
		_w2032_,
		_w2189_
	);
	LUT3 #(
		.INIT('hca)
	) name1261 (
		\sub1_data_reg_reg[59]/NET0131 ,
		_w1809_,
		_w2035_,
		_w2190_
	);
	LUT4 #(
		.INIT('h3caa)
	) name1262 (
		\sub1_data_reg_reg[60]/NET0131 ,
		_w1814_,
		_w1816_,
		_w2035_,
		_w2191_
	);
	LUT4 #(
		.INIT('hc3aa)
	) name1263 (
		\sub1_data_reg_reg[63]/NET0131 ,
		_w1639_,
		_w1794_,
		_w2035_,
		_w2192_
	);
	LUT3 #(
		.INIT('hca)
	) name1264 (
		\sub1_data_reg_reg[91]/NET0131 ,
		_w1809_,
		_w2038_,
		_w2193_
	);
	LUT4 #(
		.INIT('h3caa)
	) name1265 (
		\sub1_data_reg_reg[92]/NET0131 ,
		_w1814_,
		_w1816_,
		_w2038_,
		_w2194_
	);
	LUT4 #(
		.INIT('hc3aa)
	) name1266 (
		\sub1_data_reg_reg[95]/NET0131 ,
		_w1639_,
		_w1794_,
		_w2038_,
		_w2195_
	);
	LUT4 #(
		.INIT('haaac)
	) name1267 (
		\key_i[111]_pad ,
		\ks1_key_reg_reg[111]/NET0131 ,
		_w938_,
		_w986_,
		_w2196_
	);
	LUT3 #(
		.INIT('h69)
	) name1268 (
		_w1639_,
		_w1794_,
		_w2196_,
		_w2197_
	);
	LUT3 #(
		.INIT('h96)
	) name1269 (
		_w1600_,
		_w1604_,
		_w1608_,
		_w2198_
	);
	LUT4 #(
		.INIT('h2228)
	) name1270 (
		_w1064_,
		_w1657_,
		_w1659_,
		_w1660_,
		_w2199_
	);
	LUT4 #(
		.INIT('haa2a)
	) name1271 (
		\ks1_col_reg[18]/NET0131 ,
		\ks1_state_reg[0]/NET0131 ,
		\ks1_state_reg[1]/NET0131 ,
		\ks1_state_reg[2]/NET0131 ,
		_w2200_
	);
	LUT2 #(
		.INIT('he)
	) name1272 (
		_w2199_,
		_w2200_,
		_w2201_
	);
	LUT4 #(
		.INIT('heee2)
	) name1273 (
		\ks1_col_reg[17]/NET0131 ,
		_w1064_,
		_w2042_,
		_w2043_,
		_w2202_
	);
	LUT4 #(
		.INIT('heee2)
	) name1274 (
		\ks1_col_reg[1]/NET0131 ,
		_w1079_,
		_w2042_,
		_w2043_,
		_w2203_
	);
	LUT4 #(
		.INIT('heee2)
	) name1275 (
		\ks1_col_reg[25]/NET0131 ,
		_w1071_,
		_w2042_,
		_w2043_,
		_w2204_
	);
	LUT4 #(
		.INIT('h2228)
	) name1276 (
		_w1071_,
		_w1657_,
		_w1659_,
		_w1660_,
		_w2205_
	);
	LUT4 #(
		.INIT('haa8a)
	) name1277 (
		\ks1_col_reg[26]/NET0131 ,
		\ks1_state_reg[0]/NET0131 ,
		\ks1_state_reg[1]/NET0131 ,
		\ks1_state_reg[2]/NET0131 ,
		_w2206_
	);
	LUT2 #(
		.INIT('he)
	) name1278 (
		_w2205_,
		_w2206_,
		_w2207_
	);
	LUT4 #(
		.INIT('h2228)
	) name1279 (
		_w1079_,
		_w1657_,
		_w1659_,
		_w1660_,
		_w2208_
	);
	LUT4 #(
		.INIT('haaa2)
	) name1280 (
		\ks1_col_reg[2]/NET0131 ,
		\ks1_state_reg[0]/NET0131 ,
		\ks1_state_reg[1]/NET0131 ,
		\ks1_state_reg[2]/NET0131 ,
		_w2209_
	);
	LUT2 #(
		.INIT('he)
	) name1281 (
		_w2208_,
		_w2209_,
		_w2210_
	);
	LUT4 #(
		.INIT('heee2)
	) name1282 (
		\sub1_data_reg_reg[121]/NET0131 ,
		_w2029_,
		_w2042_,
		_w2043_,
		_w2211_
	);
	LUT4 #(
		.INIT('heee2)
	) name1283 (
		\sub1_data_reg_reg[25]/NET0131 ,
		_w2032_,
		_w2042_,
		_w2043_,
		_w2212_
	);
	LUT4 #(
		.INIT('heee2)
	) name1284 (
		\sub1_data_reg_reg[57]/NET0131 ,
		_w2035_,
		_w2042_,
		_w2043_,
		_w2213_
	);
	LUT4 #(
		.INIT('heee2)
	) name1285 (
		\sub1_data_reg_reg[89]/NET0131 ,
		_w2038_,
		_w2042_,
		_w2043_,
		_w2214_
	);
	LUT4 #(
		.INIT('h5600)
	) name1286 (
		_w1657_,
		_w1659_,
		_w1660_,
		_w2029_,
		_w2215_
	);
	LUT3 #(
		.INIT('h2a)
	) name1287 (
		\sub1_data_reg_reg[122]/NET0131 ,
		_w1692_,
		_w1761_,
		_w2216_
	);
	LUT2 #(
		.INIT('he)
	) name1288 (
		_w2215_,
		_w2216_,
		_w2217_
	);
	LUT4 #(
		.INIT('h5600)
	) name1289 (
		_w1657_,
		_w1659_,
		_w1660_,
		_w2032_,
		_w2218_
	);
	LUT3 #(
		.INIT('h2a)
	) name1290 (
		\sub1_data_reg_reg[26]/NET0131 ,
		_w1702_,
		_w1769_,
		_w2219_
	);
	LUT2 #(
		.INIT('he)
	) name1291 (
		_w2218_,
		_w2219_,
		_w2220_
	);
	LUT4 #(
		.INIT('h5600)
	) name1292 (
		_w1657_,
		_w1659_,
		_w1660_,
		_w2035_,
		_w2221_
	);
	LUT3 #(
		.INIT('h2a)
	) name1293 (
		\sub1_data_reg_reg[58]/NET0131 ,
		_w1692_,
		_w1769_,
		_w2222_
	);
	LUT2 #(
		.INIT('he)
	) name1294 (
		_w2221_,
		_w2222_,
		_w2223_
	);
	LUT4 #(
		.INIT('h5600)
	) name1295 (
		_w1657_,
		_w1659_,
		_w1660_,
		_w2038_,
		_w2224_
	);
	LUT3 #(
		.INIT('h2a)
	) name1296 (
		\sub1_data_reg_reg[90]/NET0131 ,
		_w1702_,
		_w1761_,
		_w2225_
	);
	LUT2 #(
		.INIT('he)
	) name1297 (
		_w2224_,
		_w2225_,
		_w2226_
	);
	LUT3 #(
		.INIT('h69)
	) name1298 (
		_w1436_,
		_w1600_,
		_w1602_,
		_w2227_
	);
	LUT2 #(
		.INIT('h9)
	) name1299 (
		_w1584_,
		_w1604_,
		_w2228_
	);
	LUT3 #(
		.INIT('h04)
	) name1300 (
		decrypt_i_pad,
		\round_reg[0]/NET0131 ,
		\round_reg[1]/NET0131 ,
		_w2229_
	);
	LUT4 #(
		.INIT('h0777)
	) name1301 (
		decrypt_i_pad,
		_w930_,
		_w994_,
		_w2229_,
		_w2230_
	);
	LUT4 #(
		.INIT('hcf47)
	) name1302 (
		\addroundkey_ready_o_reg/NET0131 ,
		decrypt_i_pad,
		\sub1_ready_o_reg/NET0131 ,
		_w995_,
		_w2231_
	);
	LUT2 #(
		.INIT('h1)
	) name1303 (
		\mix1_state_reg[0]/NET0131 ,
		\mix1_state_reg[1]/NET0131 ,
		_w2232_
	);
	LUT4 #(
		.INIT('h3100)
	) name1304 (
		\state_reg/NET0131 ,
		_w2231_,
		_w2230_,
		_w2232_,
		_w2233_
	);
	LUT4 #(
		.INIT('hf0b8)
	) name1305 (
		\data_o[114]_pad ,
		decrypt_i_pad,
		\sub1_data_reg_reg[114]/NET0131 ,
		_w995_,
		_w2234_
	);
	LUT3 #(
		.INIT('h04)
	) name1306 (
		\data_o[18]_pad ,
		decrypt_i_pad,
		_w995_,
		_w2235_
	);
	LUT2 #(
		.INIT('h8)
	) name1307 (
		\mix1_state_reg[0]/NET0131 ,
		\mix1_state_reg[1]/NET0131 ,
		_w2236_
	);
	LUT4 #(
		.INIT('hce00)
	) name1308 (
		decrypt_i_pad,
		\sub1_data_reg_reg[18]/NET0131 ,
		_w995_,
		_w2236_,
		_w2237_
	);
	LUT2 #(
		.INIT('h4)
	) name1309 (
		_w2235_,
		_w2237_,
		_w2238_
	);
	LUT3 #(
		.INIT('h04)
	) name1310 (
		\data_o[82]_pad ,
		decrypt_i_pad,
		_w995_,
		_w2239_
	);
	LUT2 #(
		.INIT('h2)
	) name1311 (
		\mix1_state_reg[0]/NET0131 ,
		\mix1_state_reg[1]/NET0131 ,
		_w2240_
	);
	LUT4 #(
		.INIT('hce00)
	) name1312 (
		decrypt_i_pad,
		\sub1_data_reg_reg[82]/NET0131 ,
		_w995_,
		_w2240_,
		_w2241_
	);
	LUT3 #(
		.INIT('h04)
	) name1313 (
		\data_o[50]_pad ,
		decrypt_i_pad,
		_w995_,
		_w2242_
	);
	LUT2 #(
		.INIT('h4)
	) name1314 (
		\mix1_state_reg[0]/NET0131 ,
		\mix1_state_reg[1]/NET0131 ,
		_w2243_
	);
	LUT4 #(
		.INIT('hce00)
	) name1315 (
		decrypt_i_pad,
		\sub1_data_reg_reg[50]/NET0131 ,
		_w995_,
		_w2243_,
		_w2244_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name1316 (
		_w2239_,
		_w2241_,
		_w2242_,
		_w2244_,
		_w2245_
	);
	LUT4 #(
		.INIT('h1300)
	) name1317 (
		_w2233_,
		_w2238_,
		_w2234_,
		_w2245_,
		_w2246_
	);
	LUT4 #(
		.INIT('hf0b8)
	) name1318 (
		\data_o[103]_pad ,
		decrypt_i_pad,
		\sub1_data_reg_reg[103]/NET0131 ,
		_w995_,
		_w2247_
	);
	LUT3 #(
		.INIT('h04)
	) name1319 (
		\data_o[7]_pad ,
		decrypt_i_pad,
		_w995_,
		_w2248_
	);
	LUT4 #(
		.INIT('hce00)
	) name1320 (
		decrypt_i_pad,
		\sub1_data_reg_reg[7]/NET0131 ,
		_w995_,
		_w2236_,
		_w2249_
	);
	LUT2 #(
		.INIT('h4)
	) name1321 (
		_w2248_,
		_w2249_,
		_w2250_
	);
	LUT3 #(
		.INIT('h04)
	) name1322 (
		\data_o[71]_pad ,
		decrypt_i_pad,
		_w995_,
		_w2251_
	);
	LUT4 #(
		.INIT('hce00)
	) name1323 (
		decrypt_i_pad,
		\sub1_data_reg_reg[71]/NET0131 ,
		_w995_,
		_w2240_,
		_w2252_
	);
	LUT3 #(
		.INIT('h04)
	) name1324 (
		\data_o[39]_pad ,
		decrypt_i_pad,
		_w995_,
		_w2253_
	);
	LUT4 #(
		.INIT('hce00)
	) name1325 (
		decrypt_i_pad,
		\sub1_data_reg_reg[39]/NET0131 ,
		_w995_,
		_w2243_,
		_w2254_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name1326 (
		_w2251_,
		_w2252_,
		_w2253_,
		_w2254_,
		_w2255_
	);
	LUT4 #(
		.INIT('h1300)
	) name1327 (
		_w2233_,
		_w2250_,
		_w2247_,
		_w2255_,
		_w2256_
	);
	LUT4 #(
		.INIT('hf0b8)
	) name1328 (
		\data_o[119]_pad ,
		decrypt_i_pad,
		\sub1_data_reg_reg[119]/NET0131 ,
		_w995_,
		_w2257_
	);
	LUT3 #(
		.INIT('h04)
	) name1329 (
		\data_o[23]_pad ,
		decrypt_i_pad,
		_w995_,
		_w2258_
	);
	LUT4 #(
		.INIT('hce00)
	) name1330 (
		decrypt_i_pad,
		\sub1_data_reg_reg[23]/NET0131 ,
		_w995_,
		_w2236_,
		_w2259_
	);
	LUT2 #(
		.INIT('h4)
	) name1331 (
		_w2258_,
		_w2259_,
		_w2260_
	);
	LUT3 #(
		.INIT('h04)
	) name1332 (
		\data_o[55]_pad ,
		decrypt_i_pad,
		_w995_,
		_w2261_
	);
	LUT4 #(
		.INIT('hce00)
	) name1333 (
		decrypt_i_pad,
		\sub1_data_reg_reg[55]/NET0131 ,
		_w995_,
		_w2243_,
		_w2262_
	);
	LUT3 #(
		.INIT('h04)
	) name1334 (
		\data_o[87]_pad ,
		decrypt_i_pad,
		_w995_,
		_w2263_
	);
	LUT4 #(
		.INIT('hce00)
	) name1335 (
		decrypt_i_pad,
		\sub1_data_reg_reg[87]/NET0131 ,
		_w995_,
		_w2240_,
		_w2264_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name1336 (
		_w2261_,
		_w2262_,
		_w2263_,
		_w2264_,
		_w2265_
	);
	LUT4 #(
		.INIT('h1300)
	) name1337 (
		_w2233_,
		_w2260_,
		_w2257_,
		_w2265_,
		_w2266_
	);
	LUT2 #(
		.INIT('h9)
	) name1338 (
		_w2256_,
		_w2266_,
		_w2267_
	);
	LUT4 #(
		.INIT('hf0b8)
	) name1339 (
		\data_o[117]_pad ,
		decrypt_i_pad,
		\sub1_data_reg_reg[117]/NET0131 ,
		_w995_,
		_w2268_
	);
	LUT3 #(
		.INIT('h04)
	) name1340 (
		\data_o[85]_pad ,
		decrypt_i_pad,
		_w995_,
		_w2269_
	);
	LUT4 #(
		.INIT('hce00)
	) name1341 (
		decrypt_i_pad,
		\sub1_data_reg_reg[85]/NET0131 ,
		_w995_,
		_w2240_,
		_w2270_
	);
	LUT2 #(
		.INIT('h4)
	) name1342 (
		_w2269_,
		_w2270_,
		_w2271_
	);
	LUT3 #(
		.INIT('h04)
	) name1343 (
		\data_o[21]_pad ,
		decrypt_i_pad,
		_w995_,
		_w2272_
	);
	LUT4 #(
		.INIT('hce00)
	) name1344 (
		decrypt_i_pad,
		\sub1_data_reg_reg[21]/NET0131 ,
		_w995_,
		_w2236_,
		_w2273_
	);
	LUT3 #(
		.INIT('h04)
	) name1345 (
		\data_o[53]_pad ,
		decrypt_i_pad,
		_w995_,
		_w2274_
	);
	LUT4 #(
		.INIT('hce00)
	) name1346 (
		decrypt_i_pad,
		\sub1_data_reg_reg[53]/NET0131 ,
		_w995_,
		_w2243_,
		_w2275_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name1347 (
		_w2272_,
		_w2273_,
		_w2274_,
		_w2275_,
		_w2276_
	);
	LUT4 #(
		.INIT('h1300)
	) name1348 (
		_w2233_,
		_w2271_,
		_w2268_,
		_w2276_,
		_w2277_
	);
	LUT4 #(
		.INIT('hf0b8)
	) name1349 (
		\data_o[125]_pad ,
		decrypt_i_pad,
		\sub1_data_reg_reg[125]/NET0131 ,
		_w995_,
		_w2278_
	);
	LUT3 #(
		.INIT('h04)
	) name1350 (
		\data_o[93]_pad ,
		decrypt_i_pad,
		_w995_,
		_w2279_
	);
	LUT4 #(
		.INIT('hce00)
	) name1351 (
		decrypt_i_pad,
		\sub1_data_reg_reg[93]/NET0131 ,
		_w995_,
		_w2240_,
		_w2280_
	);
	LUT2 #(
		.INIT('h4)
	) name1352 (
		_w2279_,
		_w2280_,
		_w2281_
	);
	LUT3 #(
		.INIT('h04)
	) name1353 (
		\data_o[29]_pad ,
		decrypt_i_pad,
		_w995_,
		_w2282_
	);
	LUT4 #(
		.INIT('hce00)
	) name1354 (
		decrypt_i_pad,
		\sub1_data_reg_reg[29]/NET0131 ,
		_w995_,
		_w2236_,
		_w2283_
	);
	LUT3 #(
		.INIT('h04)
	) name1355 (
		\data_o[61]_pad ,
		decrypt_i_pad,
		_w995_,
		_w2284_
	);
	LUT4 #(
		.INIT('hce00)
	) name1356 (
		decrypt_i_pad,
		\sub1_data_reg_reg[61]/NET0131 ,
		_w995_,
		_w2243_,
		_w2285_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name1357 (
		_w2282_,
		_w2283_,
		_w2284_,
		_w2285_,
		_w2286_
	);
	LUT4 #(
		.INIT('h1300)
	) name1358 (
		_w2233_,
		_w2281_,
		_w2278_,
		_w2286_,
		_w2287_
	);
	LUT4 #(
		.INIT('hf0b8)
	) name1359 (
		\data_o[101]_pad ,
		decrypt_i_pad,
		\sub1_data_reg_reg[101]/NET0131 ,
		_w995_,
		_w2288_
	);
	LUT3 #(
		.INIT('h04)
	) name1360 (
		\data_o[37]_pad ,
		decrypt_i_pad,
		_w995_,
		_w2289_
	);
	LUT4 #(
		.INIT('hce00)
	) name1361 (
		decrypt_i_pad,
		\sub1_data_reg_reg[37]/NET0131 ,
		_w995_,
		_w2243_,
		_w2290_
	);
	LUT2 #(
		.INIT('h4)
	) name1362 (
		_w2289_,
		_w2290_,
		_w2291_
	);
	LUT3 #(
		.INIT('h04)
	) name1363 (
		\data_o[69]_pad ,
		decrypt_i_pad,
		_w995_,
		_w2292_
	);
	LUT4 #(
		.INIT('hce00)
	) name1364 (
		decrypt_i_pad,
		\sub1_data_reg_reg[69]/NET0131 ,
		_w995_,
		_w2240_,
		_w2293_
	);
	LUT3 #(
		.INIT('h04)
	) name1365 (
		\data_o[5]_pad ,
		decrypt_i_pad,
		_w995_,
		_w2294_
	);
	LUT4 #(
		.INIT('hce00)
	) name1366 (
		decrypt_i_pad,
		\sub1_data_reg_reg[5]/NET0131 ,
		_w995_,
		_w2236_,
		_w2295_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name1367 (
		_w2292_,
		_w2293_,
		_w2294_,
		_w2295_,
		_w2296_
	);
	LUT4 #(
		.INIT('h1300)
	) name1368 (
		_w2233_,
		_w2291_,
		_w2288_,
		_w2296_,
		_w2297_
	);
	LUT4 #(
		.INIT('hf0b8)
	) name1369 (
		\data_o[109]_pad ,
		decrypt_i_pad,
		\sub1_data_reg_reg[109]/NET0131 ,
		_w995_,
		_w2298_
	);
	LUT3 #(
		.INIT('h04)
	) name1370 (
		\data_o[13]_pad ,
		decrypt_i_pad,
		_w995_,
		_w2299_
	);
	LUT4 #(
		.INIT('hce00)
	) name1371 (
		decrypt_i_pad,
		\sub1_data_reg_reg[13]/NET0131 ,
		_w995_,
		_w2236_,
		_w2300_
	);
	LUT2 #(
		.INIT('h4)
	) name1372 (
		_w2299_,
		_w2300_,
		_w2301_
	);
	LUT3 #(
		.INIT('h04)
	) name1373 (
		\data_o[45]_pad ,
		decrypt_i_pad,
		_w995_,
		_w2302_
	);
	LUT4 #(
		.INIT('hce00)
	) name1374 (
		decrypt_i_pad,
		\sub1_data_reg_reg[45]/NET0131 ,
		_w995_,
		_w2243_,
		_w2303_
	);
	LUT3 #(
		.INIT('h04)
	) name1375 (
		\data_o[77]_pad ,
		decrypt_i_pad,
		_w995_,
		_w2304_
	);
	LUT4 #(
		.INIT('hce00)
	) name1376 (
		decrypt_i_pad,
		\sub1_data_reg_reg[77]/NET0131 ,
		_w995_,
		_w2240_,
		_w2305_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name1377 (
		_w2302_,
		_w2303_,
		_w2304_,
		_w2305_,
		_w2306_
	);
	LUT4 #(
		.INIT('h1300)
	) name1378 (
		_w2233_,
		_w2301_,
		_w2298_,
		_w2306_,
		_w2307_
	);
	LUT2 #(
		.INIT('h9)
	) name1379 (
		_w2297_,
		_w2307_,
		_w2308_
	);
	LUT4 #(
		.INIT('h6996)
	) name1380 (
		_w2277_,
		_w2287_,
		_w2297_,
		_w2307_,
		_w2309_
	);
	LUT4 #(
		.INIT('hf0b8)
	) name1381 (
		\data_o[110]_pad ,
		decrypt_i_pad,
		\sub1_data_reg_reg[110]/NET0131 ,
		_w995_,
		_w2310_
	);
	LUT3 #(
		.INIT('h04)
	) name1382 (
		\data_o[14]_pad ,
		decrypt_i_pad,
		_w995_,
		_w2311_
	);
	LUT4 #(
		.INIT('hce00)
	) name1383 (
		decrypt_i_pad,
		\sub1_data_reg_reg[14]/NET0131 ,
		_w995_,
		_w2236_,
		_w2312_
	);
	LUT2 #(
		.INIT('h4)
	) name1384 (
		_w2311_,
		_w2312_,
		_w2313_
	);
	LUT3 #(
		.INIT('h04)
	) name1385 (
		\data_o[46]_pad ,
		decrypt_i_pad,
		_w995_,
		_w2314_
	);
	LUT4 #(
		.INIT('hce00)
	) name1386 (
		decrypt_i_pad,
		\sub1_data_reg_reg[46]/NET0131 ,
		_w995_,
		_w2243_,
		_w2315_
	);
	LUT3 #(
		.INIT('h04)
	) name1387 (
		\data_o[78]_pad ,
		decrypt_i_pad,
		_w995_,
		_w2316_
	);
	LUT4 #(
		.INIT('hce00)
	) name1388 (
		decrypt_i_pad,
		\sub1_data_reg_reg[78]/NET0131 ,
		_w995_,
		_w2240_,
		_w2317_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name1389 (
		_w2314_,
		_w2315_,
		_w2316_,
		_w2317_,
		_w2318_
	);
	LUT4 #(
		.INIT('h1300)
	) name1390 (
		_w2233_,
		_w2313_,
		_w2310_,
		_w2318_,
		_w2319_
	);
	LUT4 #(
		.INIT('hf0b8)
	) name1391 (
		\data_o[126]_pad ,
		decrypt_i_pad,
		\sub1_data_reg_reg[126]/NET0131 ,
		_w995_,
		_w2320_
	);
	LUT3 #(
		.INIT('h04)
	) name1392 (
		\data_o[94]_pad ,
		decrypt_i_pad,
		_w995_,
		_w2321_
	);
	LUT4 #(
		.INIT('hce00)
	) name1393 (
		decrypt_i_pad,
		\sub1_data_reg_reg[94]/NET0131 ,
		_w995_,
		_w2240_,
		_w2322_
	);
	LUT2 #(
		.INIT('h4)
	) name1394 (
		_w2321_,
		_w2322_,
		_w2323_
	);
	LUT3 #(
		.INIT('h04)
	) name1395 (
		\data_o[62]_pad ,
		decrypt_i_pad,
		_w995_,
		_w2324_
	);
	LUT4 #(
		.INIT('hce00)
	) name1396 (
		decrypt_i_pad,
		\sub1_data_reg_reg[62]/NET0131 ,
		_w995_,
		_w2243_,
		_w2325_
	);
	LUT3 #(
		.INIT('h04)
	) name1397 (
		\data_o[30]_pad ,
		decrypt_i_pad,
		_w995_,
		_w2326_
	);
	LUT4 #(
		.INIT('hce00)
	) name1398 (
		decrypt_i_pad,
		\sub1_data_reg_reg[30]/NET0131 ,
		_w995_,
		_w2236_,
		_w2327_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name1399 (
		_w2324_,
		_w2325_,
		_w2326_,
		_w2327_,
		_w2328_
	);
	LUT4 #(
		.INIT('h1300)
	) name1400 (
		_w2233_,
		_w2323_,
		_w2320_,
		_w2328_,
		_w2329_
	);
	LUT2 #(
		.INIT('h9)
	) name1401 (
		_w2319_,
		_w2329_,
		_w2330_
	);
	LUT4 #(
		.INIT('hf0b8)
	) name1402 (
		\data_o[98]_pad ,
		decrypt_i_pad,
		\sub1_data_reg_reg[98]/NET0131 ,
		_w995_,
		_w2331_
	);
	LUT3 #(
		.INIT('h04)
	) name1403 (
		\data_o[2]_pad ,
		decrypt_i_pad,
		_w995_,
		_w2332_
	);
	LUT4 #(
		.INIT('hce00)
	) name1404 (
		decrypt_i_pad,
		\sub1_data_reg_reg[2]/NET0131 ,
		_w995_,
		_w2236_,
		_w2333_
	);
	LUT2 #(
		.INIT('h4)
	) name1405 (
		_w2332_,
		_w2333_,
		_w2334_
	);
	LUT3 #(
		.INIT('h04)
	) name1406 (
		\data_o[66]_pad ,
		decrypt_i_pad,
		_w995_,
		_w2335_
	);
	LUT4 #(
		.INIT('hce00)
	) name1407 (
		decrypt_i_pad,
		\sub1_data_reg_reg[66]/NET0131 ,
		_w995_,
		_w2240_,
		_w2336_
	);
	LUT3 #(
		.INIT('h04)
	) name1408 (
		\data_o[34]_pad ,
		decrypt_i_pad,
		_w995_,
		_w2337_
	);
	LUT4 #(
		.INIT('hce00)
	) name1409 (
		decrypt_i_pad,
		\sub1_data_reg_reg[34]/NET0131 ,
		_w995_,
		_w2243_,
		_w2338_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name1410 (
		_w2335_,
		_w2336_,
		_w2337_,
		_w2338_,
		_w2339_
	);
	LUT4 #(
		.INIT('h1300)
	) name1411 (
		_w2233_,
		_w2334_,
		_w2331_,
		_w2339_,
		_w2340_
	);
	LUT4 #(
		.INIT('h9669)
	) name1412 (
		_w2267_,
		_w2309_,
		_w2330_,
		_w2340_,
		_w2341_
	);
	LUT4 #(
		.INIT('hf0b8)
	) name1413 (
		\data_o[97]_pad ,
		decrypt_i_pad,
		\sub1_data_reg_reg[97]/NET0131 ,
		_w995_,
		_w2342_
	);
	LUT3 #(
		.INIT('h04)
	) name1414 (
		\data_o[33]_pad ,
		decrypt_i_pad,
		_w995_,
		_w2343_
	);
	LUT4 #(
		.INIT('hce00)
	) name1415 (
		decrypt_i_pad,
		\sub1_data_reg_reg[33]/NET0131 ,
		_w995_,
		_w2243_,
		_w2344_
	);
	LUT2 #(
		.INIT('h4)
	) name1416 (
		_w2343_,
		_w2344_,
		_w2345_
	);
	LUT3 #(
		.INIT('h04)
	) name1417 (
		\data_o[1]_pad ,
		decrypt_i_pad,
		_w995_,
		_w2346_
	);
	LUT4 #(
		.INIT('hce00)
	) name1418 (
		decrypt_i_pad,
		\sub1_data_reg_reg[1]/NET0131 ,
		_w995_,
		_w2236_,
		_w2347_
	);
	LUT3 #(
		.INIT('h04)
	) name1419 (
		\data_o[65]_pad ,
		decrypt_i_pad,
		_w995_,
		_w2348_
	);
	LUT4 #(
		.INIT('hce00)
	) name1420 (
		decrypt_i_pad,
		\sub1_data_reg_reg[65]/NET0131 ,
		_w995_,
		_w2240_,
		_w2349_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name1421 (
		_w2346_,
		_w2347_,
		_w2348_,
		_w2349_,
		_w2350_
	);
	LUT4 #(
		.INIT('h1300)
	) name1422 (
		_w2233_,
		_w2345_,
		_w2342_,
		_w2350_,
		_w2351_
	);
	LUT4 #(
		.INIT('hf0b8)
	) name1423 (
		\data_o[113]_pad ,
		decrypt_i_pad,
		\sub1_data_reg_reg[113]/NET0131 ,
		_w995_,
		_w2352_
	);
	LUT3 #(
		.INIT('h04)
	) name1424 (
		\data_o[49]_pad ,
		decrypt_i_pad,
		_w995_,
		_w2353_
	);
	LUT4 #(
		.INIT('hce00)
	) name1425 (
		decrypt_i_pad,
		\sub1_data_reg_reg[49]/NET0131 ,
		_w995_,
		_w2243_,
		_w2354_
	);
	LUT2 #(
		.INIT('h4)
	) name1426 (
		_w2353_,
		_w2354_,
		_w2355_
	);
	LUT3 #(
		.INIT('h04)
	) name1427 (
		\data_o[17]_pad ,
		decrypt_i_pad,
		_w995_,
		_w2356_
	);
	LUT4 #(
		.INIT('hce00)
	) name1428 (
		decrypt_i_pad,
		\sub1_data_reg_reg[17]/NET0131 ,
		_w995_,
		_w2236_,
		_w2357_
	);
	LUT3 #(
		.INIT('h04)
	) name1429 (
		\data_o[81]_pad ,
		decrypt_i_pad,
		_w995_,
		_w2358_
	);
	LUT4 #(
		.INIT('hce00)
	) name1430 (
		decrypt_i_pad,
		\sub1_data_reg_reg[81]/NET0131 ,
		_w995_,
		_w2240_,
		_w2359_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name1431 (
		_w2356_,
		_w2357_,
		_w2358_,
		_w2359_,
		_w2360_
	);
	LUT4 #(
		.INIT('h1300)
	) name1432 (
		_w2233_,
		_w2355_,
		_w2352_,
		_w2360_,
		_w2361_
	);
	LUT2 #(
		.INIT('h9)
	) name1433 (
		_w2351_,
		_w2361_,
		_w2362_
	);
	LUT4 #(
		.INIT('hf0b8)
	) name1434 (
		\data_o[121]_pad ,
		decrypt_i_pad,
		\sub1_data_reg_reg[121]/NET0131 ,
		_w995_,
		_w2363_
	);
	LUT3 #(
		.INIT('h04)
	) name1435 (
		\data_o[89]_pad ,
		decrypt_i_pad,
		_w995_,
		_w2364_
	);
	LUT4 #(
		.INIT('hce00)
	) name1436 (
		decrypt_i_pad,
		\sub1_data_reg_reg[89]/NET0131 ,
		_w995_,
		_w2240_,
		_w2365_
	);
	LUT2 #(
		.INIT('h4)
	) name1437 (
		_w2364_,
		_w2365_,
		_w2366_
	);
	LUT3 #(
		.INIT('h04)
	) name1438 (
		\data_o[25]_pad ,
		decrypt_i_pad,
		_w995_,
		_w2367_
	);
	LUT4 #(
		.INIT('hce00)
	) name1439 (
		decrypt_i_pad,
		\sub1_data_reg_reg[25]/NET0131 ,
		_w995_,
		_w2236_,
		_w2368_
	);
	LUT3 #(
		.INIT('h04)
	) name1440 (
		\data_o[57]_pad ,
		decrypt_i_pad,
		_w995_,
		_w2369_
	);
	LUT4 #(
		.INIT('hce00)
	) name1441 (
		decrypt_i_pad,
		\sub1_data_reg_reg[57]/NET0131 ,
		_w995_,
		_w2243_,
		_w2370_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name1442 (
		_w2367_,
		_w2368_,
		_w2369_,
		_w2370_,
		_w2371_
	);
	LUT4 #(
		.INIT('h1300)
	) name1443 (
		_w2233_,
		_w2366_,
		_w2363_,
		_w2371_,
		_w2372_
	);
	LUT4 #(
		.INIT('hf0b8)
	) name1444 (
		\data_o[105]_pad ,
		decrypt_i_pad,
		\sub1_data_reg_reg[105]/NET0131 ,
		_w995_,
		_w2373_
	);
	LUT3 #(
		.INIT('h04)
	) name1445 (
		\data_o[41]_pad ,
		decrypt_i_pad,
		_w995_,
		_w2374_
	);
	LUT4 #(
		.INIT('hce00)
	) name1446 (
		decrypt_i_pad,
		\sub1_data_reg_reg[41]/NET0131 ,
		_w995_,
		_w2243_,
		_w2375_
	);
	LUT2 #(
		.INIT('h4)
	) name1447 (
		_w2374_,
		_w2375_,
		_w2376_
	);
	LUT3 #(
		.INIT('h04)
	) name1448 (
		\data_o[9]_pad ,
		decrypt_i_pad,
		_w995_,
		_w2377_
	);
	LUT4 #(
		.INIT('hce00)
	) name1449 (
		decrypt_i_pad,
		\sub1_data_reg_reg[9]/NET0131 ,
		_w995_,
		_w2236_,
		_w2378_
	);
	LUT3 #(
		.INIT('h04)
	) name1450 (
		\data_o[73]_pad ,
		decrypt_i_pad,
		_w995_,
		_w2379_
	);
	LUT4 #(
		.INIT('hce00)
	) name1451 (
		decrypt_i_pad,
		\sub1_data_reg_reg[73]/NET0131 ,
		_w995_,
		_w2240_,
		_w2380_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name1452 (
		_w2377_,
		_w2378_,
		_w2379_,
		_w2380_,
		_w2381_
	);
	LUT4 #(
		.INIT('h1300)
	) name1453 (
		_w2233_,
		_w2376_,
		_w2373_,
		_w2381_,
		_w2382_
	);
	LUT4 #(
		.INIT('h6996)
	) name1454 (
		_w2351_,
		_w2361_,
		_w2372_,
		_w2382_,
		_w2383_
	);
	LUT4 #(
		.INIT('h2882)
	) name1455 (
		decrypt_i_pad,
		_w2246_,
		_w2341_,
		_w2383_,
		_w2384_
	);
	LUT4 #(
		.INIT('hf0b8)
	) name1456 (
		\data_o[116]_pad ,
		decrypt_i_pad,
		\sub1_data_reg_reg[116]/NET0131 ,
		_w995_,
		_w2385_
	);
	LUT3 #(
		.INIT('h04)
	) name1457 (
		\data_o[52]_pad ,
		decrypt_i_pad,
		_w995_,
		_w2386_
	);
	LUT4 #(
		.INIT('hce00)
	) name1458 (
		decrypt_i_pad,
		\sub1_data_reg_reg[52]/NET0131 ,
		_w995_,
		_w2243_,
		_w2387_
	);
	LUT2 #(
		.INIT('h4)
	) name1459 (
		_w2386_,
		_w2387_,
		_w2388_
	);
	LUT3 #(
		.INIT('h04)
	) name1460 (
		\data_o[84]_pad ,
		decrypt_i_pad,
		_w995_,
		_w2389_
	);
	LUT4 #(
		.INIT('hce00)
	) name1461 (
		decrypt_i_pad,
		\sub1_data_reg_reg[84]/NET0131 ,
		_w995_,
		_w2240_,
		_w2390_
	);
	LUT3 #(
		.INIT('h04)
	) name1462 (
		\data_o[20]_pad ,
		decrypt_i_pad,
		_w995_,
		_w2391_
	);
	LUT4 #(
		.INIT('hce00)
	) name1463 (
		decrypt_i_pad,
		\sub1_data_reg_reg[20]/NET0131 ,
		_w995_,
		_w2236_,
		_w2392_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name1464 (
		_w2389_,
		_w2390_,
		_w2391_,
		_w2392_,
		_w2393_
	);
	LUT4 #(
		.INIT('h1300)
	) name1465 (
		_w2233_,
		_w2388_,
		_w2385_,
		_w2393_,
		_w2394_
	);
	LUT4 #(
		.INIT('hf0b8)
	) name1466 (
		\data_o[124]_pad ,
		decrypt_i_pad,
		\sub1_data_reg_reg[124]/NET0131 ,
		_w995_,
		_w2395_
	);
	LUT3 #(
		.INIT('h04)
	) name1467 (
		\data_o[60]_pad ,
		decrypt_i_pad,
		_w995_,
		_w2396_
	);
	LUT4 #(
		.INIT('hce00)
	) name1468 (
		decrypt_i_pad,
		\sub1_data_reg_reg[60]/NET0131 ,
		_w995_,
		_w2243_,
		_w2397_
	);
	LUT2 #(
		.INIT('h4)
	) name1469 (
		_w2396_,
		_w2397_,
		_w2398_
	);
	LUT3 #(
		.INIT('h04)
	) name1470 (
		\data_o[28]_pad ,
		decrypt_i_pad,
		_w995_,
		_w2399_
	);
	LUT4 #(
		.INIT('hce00)
	) name1471 (
		decrypt_i_pad,
		\sub1_data_reg_reg[28]/NET0131 ,
		_w995_,
		_w2236_,
		_w2400_
	);
	LUT3 #(
		.INIT('h04)
	) name1472 (
		\data_o[92]_pad ,
		decrypt_i_pad,
		_w995_,
		_w2401_
	);
	LUT4 #(
		.INIT('hce00)
	) name1473 (
		decrypt_i_pad,
		\sub1_data_reg_reg[92]/NET0131 ,
		_w995_,
		_w2240_,
		_w2402_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name1474 (
		_w2399_,
		_w2400_,
		_w2401_,
		_w2402_,
		_w2403_
	);
	LUT4 #(
		.INIT('h1300)
	) name1475 (
		_w2233_,
		_w2398_,
		_w2395_,
		_w2403_,
		_w2404_
	);
	LUT4 #(
		.INIT('hf0b8)
	) name1476 (
		\data_o[108]_pad ,
		decrypt_i_pad,
		\sub1_data_reg_reg[108]/NET0131 ,
		_w995_,
		_w2405_
	);
	LUT3 #(
		.INIT('h04)
	) name1477 (
		\data_o[44]_pad ,
		decrypt_i_pad,
		_w995_,
		_w2406_
	);
	LUT4 #(
		.INIT('hce00)
	) name1478 (
		decrypt_i_pad,
		\sub1_data_reg_reg[44]/NET0131 ,
		_w995_,
		_w2243_,
		_w2407_
	);
	LUT2 #(
		.INIT('h4)
	) name1479 (
		_w2406_,
		_w2407_,
		_w2408_
	);
	LUT3 #(
		.INIT('h04)
	) name1480 (
		\data_o[12]_pad ,
		decrypt_i_pad,
		_w995_,
		_w2409_
	);
	LUT4 #(
		.INIT('hce00)
	) name1481 (
		decrypt_i_pad,
		\sub1_data_reg_reg[12]/NET0131 ,
		_w995_,
		_w2236_,
		_w2410_
	);
	LUT3 #(
		.INIT('h04)
	) name1482 (
		\data_o[76]_pad ,
		decrypt_i_pad,
		_w995_,
		_w2411_
	);
	LUT4 #(
		.INIT('hce00)
	) name1483 (
		decrypt_i_pad,
		\sub1_data_reg_reg[76]/NET0131 ,
		_w995_,
		_w2240_,
		_w2412_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name1484 (
		_w2409_,
		_w2410_,
		_w2411_,
		_w2412_,
		_w2413_
	);
	LUT4 #(
		.INIT('h1300)
	) name1485 (
		_w2233_,
		_w2408_,
		_w2405_,
		_w2413_,
		_w2414_
	);
	LUT2 #(
		.INIT('h9)
	) name1486 (
		_w2404_,
		_w2414_,
		_w2415_
	);
	LUT3 #(
		.INIT('h69)
	) name1487 (
		_w2394_,
		_w2404_,
		_w2414_,
		_w2416_
	);
	LUT4 #(
		.INIT('hf0b8)
	) name1488 (
		\data_o[123]_pad ,
		decrypt_i_pad,
		\sub1_data_reg_reg[123]/NET0131 ,
		_w995_,
		_w2417_
	);
	LUT3 #(
		.INIT('h04)
	) name1489 (
		\data_o[27]_pad ,
		decrypt_i_pad,
		_w995_,
		_w2418_
	);
	LUT4 #(
		.INIT('hce00)
	) name1490 (
		decrypt_i_pad,
		\sub1_data_reg_reg[27]/NET0131 ,
		_w995_,
		_w2236_,
		_w2419_
	);
	LUT2 #(
		.INIT('h4)
	) name1491 (
		_w2418_,
		_w2419_,
		_w2420_
	);
	LUT3 #(
		.INIT('h04)
	) name1492 (
		\data_o[91]_pad ,
		decrypt_i_pad,
		_w995_,
		_w2421_
	);
	LUT4 #(
		.INIT('hce00)
	) name1493 (
		decrypt_i_pad,
		\sub1_data_reg_reg[91]/NET0131 ,
		_w995_,
		_w2240_,
		_w2422_
	);
	LUT3 #(
		.INIT('h04)
	) name1494 (
		\data_o[59]_pad ,
		decrypt_i_pad,
		_w995_,
		_w2423_
	);
	LUT4 #(
		.INIT('hce00)
	) name1495 (
		decrypt_i_pad,
		\sub1_data_reg_reg[59]/NET0131 ,
		_w995_,
		_w2243_,
		_w2424_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name1496 (
		_w2421_,
		_w2422_,
		_w2423_,
		_w2424_,
		_w2425_
	);
	LUT4 #(
		.INIT('h1300)
	) name1497 (
		_w2233_,
		_w2420_,
		_w2417_,
		_w2425_,
		_w2426_
	);
	LUT4 #(
		.INIT('hf0b8)
	) name1498 (
		\data_o[99]_pad ,
		decrypt_i_pad,
		\sub1_data_reg_reg[99]/NET0131 ,
		_w995_,
		_w2427_
	);
	LUT3 #(
		.INIT('h04)
	) name1499 (
		\data_o[3]_pad ,
		decrypt_i_pad,
		_w995_,
		_w2428_
	);
	LUT4 #(
		.INIT('hce00)
	) name1500 (
		decrypt_i_pad,
		\sub1_data_reg_reg[3]/NET0131 ,
		_w995_,
		_w2236_,
		_w2429_
	);
	LUT2 #(
		.INIT('h4)
	) name1501 (
		_w2428_,
		_w2429_,
		_w2430_
	);
	LUT3 #(
		.INIT('h04)
	) name1502 (
		\data_o[35]_pad ,
		decrypt_i_pad,
		_w995_,
		_w2431_
	);
	LUT4 #(
		.INIT('hce00)
	) name1503 (
		decrypt_i_pad,
		\sub1_data_reg_reg[35]/NET0131 ,
		_w995_,
		_w2243_,
		_w2432_
	);
	LUT3 #(
		.INIT('h04)
	) name1504 (
		\data_o[67]_pad ,
		decrypt_i_pad,
		_w995_,
		_w2433_
	);
	LUT4 #(
		.INIT('hce00)
	) name1505 (
		decrypt_i_pad,
		\sub1_data_reg_reg[67]/NET0131 ,
		_w995_,
		_w2240_,
		_w2434_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name1506 (
		_w2431_,
		_w2432_,
		_w2433_,
		_w2434_,
		_w2435_
	);
	LUT4 #(
		.INIT('h1300)
	) name1507 (
		_w2233_,
		_w2430_,
		_w2427_,
		_w2435_,
		_w2436_
	);
	LUT2 #(
		.INIT('h9)
	) name1508 (
		_w2426_,
		_w2436_,
		_w2437_
	);
	LUT4 #(
		.INIT('hf0b8)
	) name1509 (
		\data_o[127]_pad ,
		decrypt_i_pad,
		\sub1_data_reg_reg[127]/NET0131 ,
		_w995_,
		_w2438_
	);
	LUT3 #(
		.INIT('h04)
	) name1510 (
		\data_o[63]_pad ,
		decrypt_i_pad,
		_w995_,
		_w2439_
	);
	LUT4 #(
		.INIT('hce00)
	) name1511 (
		decrypt_i_pad,
		\sub1_data_reg_reg[63]/NET0131 ,
		_w995_,
		_w2243_,
		_w2440_
	);
	LUT2 #(
		.INIT('h4)
	) name1512 (
		_w2439_,
		_w2440_,
		_w2441_
	);
	LUT3 #(
		.INIT('h04)
	) name1513 (
		\data_o[95]_pad ,
		decrypt_i_pad,
		_w995_,
		_w2442_
	);
	LUT4 #(
		.INIT('hce00)
	) name1514 (
		decrypt_i_pad,
		\sub1_data_reg_reg[95]/NET0131 ,
		_w995_,
		_w2240_,
		_w2443_
	);
	LUT3 #(
		.INIT('h04)
	) name1515 (
		\data_o[31]_pad ,
		decrypt_i_pad,
		_w995_,
		_w2444_
	);
	LUT4 #(
		.INIT('hce00)
	) name1516 (
		decrypt_i_pad,
		\sub1_data_reg_reg[31]/NET0131 ,
		_w995_,
		_w2236_,
		_w2445_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name1517 (
		_w2442_,
		_w2443_,
		_w2444_,
		_w2445_,
		_w2446_
	);
	LUT4 #(
		.INIT('h1300)
	) name1518 (
		_w2233_,
		_w2441_,
		_w2438_,
		_w2446_,
		_w2447_
	);
	LUT2 #(
		.INIT('h9)
	) name1519 (
		_w2256_,
		_w2447_,
		_w2448_
	);
	LUT4 #(
		.INIT('h6996)
	) name1520 (
		_w2256_,
		_w2426_,
		_w2436_,
		_w2447_,
		_w2449_
	);
	LUT2 #(
		.INIT('h9)
	) name1521 (
		_w2416_,
		_w2449_,
		_w2450_
	);
	LUT4 #(
		.INIT('he22e)
	) name1522 (
		\mix1_data_reg_reg[100]/NET0131 ,
		_w2233_,
		_w2384_,
		_w2450_,
		_w2451_
	);
	LUT4 #(
		.INIT('h9669)
	) name1523 (
		_w2277_,
		_w2287_,
		_w2307_,
		_w2404_,
		_w2452_
	);
	LUT4 #(
		.INIT('hf0b8)
	) name1524 (
		\data_o[100]_pad ,
		decrypt_i_pad,
		\sub1_data_reg_reg[100]/NET0131 ,
		_w995_,
		_w2453_
	);
	LUT3 #(
		.INIT('h04)
	) name1525 (
		\data_o[4]_pad ,
		decrypt_i_pad,
		_w995_,
		_w2454_
	);
	LUT4 #(
		.INIT('hce00)
	) name1526 (
		decrypt_i_pad,
		\sub1_data_reg_reg[4]/NET0131 ,
		_w995_,
		_w2236_,
		_w2455_
	);
	LUT2 #(
		.INIT('h4)
	) name1527 (
		_w2454_,
		_w2455_,
		_w2456_
	);
	LUT3 #(
		.INIT('h04)
	) name1528 (
		\data_o[36]_pad ,
		decrypt_i_pad,
		_w995_,
		_w2457_
	);
	LUT4 #(
		.INIT('hce00)
	) name1529 (
		decrypt_i_pad,
		\sub1_data_reg_reg[36]/NET0131 ,
		_w995_,
		_w2243_,
		_w2458_
	);
	LUT3 #(
		.INIT('h04)
	) name1530 (
		\data_o[68]_pad ,
		decrypt_i_pad,
		_w995_,
		_w2459_
	);
	LUT4 #(
		.INIT('hce00)
	) name1531 (
		decrypt_i_pad,
		\sub1_data_reg_reg[68]/NET0131 ,
		_w995_,
		_w2240_,
		_w2460_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name1532 (
		_w2457_,
		_w2458_,
		_w2459_,
		_w2460_,
		_w2461_
	);
	LUT4 #(
		.INIT('h1300)
	) name1533 (
		_w2233_,
		_w2456_,
		_w2453_,
		_w2461_,
		_w2462_
	);
	LUT4 #(
		.INIT('hf0b8)
	) name1534 (
		\data_o[102]_pad ,
		decrypt_i_pad,
		\sub1_data_reg_reg[102]/NET0131 ,
		_w995_,
		_w2463_
	);
	LUT3 #(
		.INIT('h04)
	) name1535 (
		\data_o[6]_pad ,
		decrypt_i_pad,
		_w995_,
		_w2464_
	);
	LUT4 #(
		.INIT('hce00)
	) name1536 (
		decrypt_i_pad,
		\sub1_data_reg_reg[6]/NET0131 ,
		_w995_,
		_w2236_,
		_w2465_
	);
	LUT2 #(
		.INIT('h4)
	) name1537 (
		_w2464_,
		_w2465_,
		_w2466_
	);
	LUT3 #(
		.INIT('h04)
	) name1538 (
		\data_o[38]_pad ,
		decrypt_i_pad,
		_w995_,
		_w2467_
	);
	LUT4 #(
		.INIT('hce00)
	) name1539 (
		decrypt_i_pad,
		\sub1_data_reg_reg[38]/NET0131 ,
		_w995_,
		_w2243_,
		_w2468_
	);
	LUT3 #(
		.INIT('h04)
	) name1540 (
		\data_o[70]_pad ,
		decrypt_i_pad,
		_w995_,
		_w2469_
	);
	LUT4 #(
		.INIT('hce00)
	) name1541 (
		decrypt_i_pad,
		\sub1_data_reg_reg[70]/NET0131 ,
		_w995_,
		_w2240_,
		_w2470_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name1542 (
		_w2467_,
		_w2468_,
		_w2469_,
		_w2470_,
		_w2471_
	);
	LUT4 #(
		.INIT('h1300)
	) name1543 (
		_w2233_,
		_w2466_,
		_w2463_,
		_w2471_,
		_w2472_
	);
	LUT2 #(
		.INIT('h9)
	) name1544 (
		_w2329_,
		_w2472_,
		_w2473_
	);
	LUT4 #(
		.INIT('hf0b8)
	) name1545 (
		\data_o[118]_pad ,
		decrypt_i_pad,
		\sub1_data_reg_reg[118]/NET0131 ,
		_w995_,
		_w2474_
	);
	LUT3 #(
		.INIT('h04)
	) name1546 (
		\data_o[86]_pad ,
		decrypt_i_pad,
		_w995_,
		_w2475_
	);
	LUT4 #(
		.INIT('hce00)
	) name1547 (
		decrypt_i_pad,
		\sub1_data_reg_reg[86]/NET0131 ,
		_w995_,
		_w2240_,
		_w2476_
	);
	LUT2 #(
		.INIT('h4)
	) name1548 (
		_w2475_,
		_w2476_,
		_w2477_
	);
	LUT3 #(
		.INIT('h04)
	) name1549 (
		\data_o[54]_pad ,
		decrypt_i_pad,
		_w995_,
		_w2478_
	);
	LUT4 #(
		.INIT('hce00)
	) name1550 (
		decrypt_i_pad,
		\sub1_data_reg_reg[54]/NET0131 ,
		_w995_,
		_w2243_,
		_w2479_
	);
	LUT3 #(
		.INIT('h04)
	) name1551 (
		\data_o[22]_pad ,
		decrypt_i_pad,
		_w995_,
		_w2480_
	);
	LUT4 #(
		.INIT('hce00)
	) name1552 (
		decrypt_i_pad,
		\sub1_data_reg_reg[22]/NET0131 ,
		_w995_,
		_w2236_,
		_w2481_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name1553 (
		_w2478_,
		_w2479_,
		_w2480_,
		_w2481_,
		_w2482_
	);
	LUT4 #(
		.INIT('h1300)
	) name1554 (
		_w2233_,
		_w2477_,
		_w2474_,
		_w2482_,
		_w2483_
	);
	LUT4 #(
		.INIT('h6996)
	) name1555 (
		_w2256_,
		_w2266_,
		_w2319_,
		_w2483_,
		_w2484_
	);
	LUT3 #(
		.INIT('h96)
	) name1556 (
		_w2436_,
		_w2473_,
		_w2484_,
		_w2485_
	);
	LUT4 #(
		.INIT('hf0b8)
	) name1557 (
		\data_o[115]_pad ,
		decrypt_i_pad,
		\sub1_data_reg_reg[115]/NET0131 ,
		_w995_,
		_w2486_
	);
	LUT3 #(
		.INIT('h04)
	) name1558 (
		\data_o[19]_pad ,
		decrypt_i_pad,
		_w995_,
		_w2487_
	);
	LUT4 #(
		.INIT('hce00)
	) name1559 (
		decrypt_i_pad,
		\sub1_data_reg_reg[19]/NET0131 ,
		_w995_,
		_w2236_,
		_w2488_
	);
	LUT2 #(
		.INIT('h4)
	) name1560 (
		_w2487_,
		_w2488_,
		_w2489_
	);
	LUT3 #(
		.INIT('h04)
	) name1561 (
		\data_o[51]_pad ,
		decrypt_i_pad,
		_w995_,
		_w2490_
	);
	LUT4 #(
		.INIT('hce00)
	) name1562 (
		decrypt_i_pad,
		\sub1_data_reg_reg[51]/NET0131 ,
		_w995_,
		_w2243_,
		_w2491_
	);
	LUT3 #(
		.INIT('h04)
	) name1563 (
		\data_o[83]_pad ,
		decrypt_i_pad,
		_w995_,
		_w2492_
	);
	LUT4 #(
		.INIT('hce00)
	) name1564 (
		decrypt_i_pad,
		\sub1_data_reg_reg[83]/NET0131 ,
		_w995_,
		_w2240_,
		_w2493_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name1565 (
		_w2490_,
		_w2491_,
		_w2492_,
		_w2493_,
		_w2494_
	);
	LUT4 #(
		.INIT('h1300)
	) name1566 (
		_w2233_,
		_w2489_,
		_w2486_,
		_w2494_,
		_w2495_
	);
	LUT4 #(
		.INIT('hf0b8)
	) name1567 (
		\data_o[122]_pad ,
		decrypt_i_pad,
		\sub1_data_reg_reg[122]/NET0131 ,
		_w995_,
		_w2496_
	);
	LUT3 #(
		.INIT('h04)
	) name1568 (
		\data_o[90]_pad ,
		decrypt_i_pad,
		_w995_,
		_w2497_
	);
	LUT4 #(
		.INIT('hce00)
	) name1569 (
		decrypt_i_pad,
		\sub1_data_reg_reg[90]/NET0131 ,
		_w995_,
		_w2240_,
		_w2498_
	);
	LUT2 #(
		.INIT('h4)
	) name1570 (
		_w2497_,
		_w2498_,
		_w2499_
	);
	LUT3 #(
		.INIT('h04)
	) name1571 (
		\data_o[58]_pad ,
		decrypt_i_pad,
		_w995_,
		_w2500_
	);
	LUT4 #(
		.INIT('hce00)
	) name1572 (
		decrypt_i_pad,
		\sub1_data_reg_reg[58]/NET0131 ,
		_w995_,
		_w2243_,
		_w2501_
	);
	LUT3 #(
		.INIT('h04)
	) name1573 (
		\data_o[26]_pad ,
		decrypt_i_pad,
		_w995_,
		_w2502_
	);
	LUT4 #(
		.INIT('hce00)
	) name1574 (
		decrypt_i_pad,
		\sub1_data_reg_reg[26]/NET0131 ,
		_w995_,
		_w2236_,
		_w2503_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name1575 (
		_w2500_,
		_w2501_,
		_w2502_,
		_w2503_,
		_w2504_
	);
	LUT4 #(
		.INIT('h1300)
	) name1576 (
		_w2233_,
		_w2499_,
		_w2496_,
		_w2504_,
		_w2505_
	);
	LUT4 #(
		.INIT('h6996)
	) name1577 (
		_w2256_,
		_w2340_,
		_w2447_,
		_w2505_,
		_w2506_
	);
	LUT2 #(
		.INIT('h6)
	) name1578 (
		_w2495_,
		_w2506_,
		_w2507_
	);
	LUT4 #(
		.INIT('hf0b8)
	) name1579 (
		\data_o[111]_pad ,
		decrypt_i_pad,
		\sub1_data_reg_reg[111]/NET0131 ,
		_w995_,
		_w2508_
	);
	LUT3 #(
		.INIT('h04)
	) name1580 (
		\data_o[15]_pad ,
		decrypt_i_pad,
		_w995_,
		_w2509_
	);
	LUT4 #(
		.INIT('hce00)
	) name1581 (
		decrypt_i_pad,
		\sub1_data_reg_reg[15]/NET0131 ,
		_w995_,
		_w2236_,
		_w2510_
	);
	LUT2 #(
		.INIT('h4)
	) name1582 (
		_w2509_,
		_w2510_,
		_w2511_
	);
	LUT3 #(
		.INIT('h04)
	) name1583 (
		\data_o[79]_pad ,
		decrypt_i_pad,
		_w995_,
		_w2512_
	);
	LUT4 #(
		.INIT('hce00)
	) name1584 (
		decrypt_i_pad,
		\sub1_data_reg_reg[79]/NET0131 ,
		_w995_,
		_w2240_,
		_w2513_
	);
	LUT3 #(
		.INIT('h04)
	) name1585 (
		\data_o[47]_pad ,
		decrypt_i_pad,
		_w995_,
		_w2514_
	);
	LUT4 #(
		.INIT('hce00)
	) name1586 (
		decrypt_i_pad,
		\sub1_data_reg_reg[47]/NET0131 ,
		_w995_,
		_w2243_,
		_w2515_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name1587 (
		_w2512_,
		_w2513_,
		_w2514_,
		_w2515_,
		_w2516_
	);
	LUT4 #(
		.INIT('h1300)
	) name1588 (
		_w2233_,
		_w2511_,
		_w2508_,
		_w2516_,
		_w2517_
	);
	LUT2 #(
		.INIT('h9)
	) name1589 (
		_w2266_,
		_w2517_,
		_w2518_
	);
	LUT4 #(
		.INIT('hf0b8)
	) name1590 (
		\data_o[106]_pad ,
		decrypt_i_pad,
		\sub1_data_reg_reg[106]/NET0131 ,
		_w995_,
		_w2519_
	);
	LUT3 #(
		.INIT('h04)
	) name1591 (
		\data_o[74]_pad ,
		decrypt_i_pad,
		_w995_,
		_w2520_
	);
	LUT4 #(
		.INIT('hce00)
	) name1592 (
		decrypt_i_pad,
		\sub1_data_reg_reg[74]/NET0131 ,
		_w995_,
		_w2240_,
		_w2521_
	);
	LUT2 #(
		.INIT('h4)
	) name1593 (
		_w2520_,
		_w2521_,
		_w2522_
	);
	LUT3 #(
		.INIT('h04)
	) name1594 (
		\data_o[10]_pad ,
		decrypt_i_pad,
		_w995_,
		_w2523_
	);
	LUT4 #(
		.INIT('hce00)
	) name1595 (
		decrypt_i_pad,
		\sub1_data_reg_reg[10]/NET0131 ,
		_w995_,
		_w2236_,
		_w2524_
	);
	LUT3 #(
		.INIT('h04)
	) name1596 (
		\data_o[42]_pad ,
		decrypt_i_pad,
		_w995_,
		_w2525_
	);
	LUT4 #(
		.INIT('hce00)
	) name1597 (
		decrypt_i_pad,
		\sub1_data_reg_reg[42]/NET0131 ,
		_w995_,
		_w2243_,
		_w2526_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name1598 (
		_w2523_,
		_w2524_,
		_w2525_,
		_w2526_,
		_w2527_
	);
	LUT4 #(
		.INIT('h1300)
	) name1599 (
		_w2233_,
		_w2522_,
		_w2519_,
		_w2527_,
		_w2528_
	);
	LUT2 #(
		.INIT('h6)
	) name1600 (
		_w2246_,
		_w2528_,
		_w2529_
	);
	LUT4 #(
		.INIT('h9669)
	) name1601 (
		_w2246_,
		_w2266_,
		_w2517_,
		_w2528_,
		_w2530_
	);
	LUT3 #(
		.INIT('h96)
	) name1602 (
		_w2495_,
		_w2506_,
		_w2530_,
		_w2531_
	);
	LUT4 #(
		.INIT('h3993)
	) name1603 (
		decrypt_i_pad,
		_w2462_,
		_w2485_,
		_w2531_,
		_w2532_
	);
	LUT4 #(
		.INIT('he22e)
	) name1604 (
		\mix1_data_reg_reg[101]/NET0131 ,
		_w2233_,
		_w2452_,
		_w2532_,
		_w2533_
	);
	LUT2 #(
		.INIT('h9)
	) name1605 (
		_w2256_,
		_w2517_,
		_w2534_
	);
	LUT2 #(
		.INIT('h6)
	) name1606 (
		_w2340_,
		_w2528_,
		_w2535_
	);
	LUT4 #(
		.INIT('h9669)
	) name1607 (
		_w2256_,
		_w2340_,
		_w2517_,
		_w2528_,
		_w2536_
	);
	LUT4 #(
		.INIT('hf0b8)
	) name1608 (
		\data_o[104]_pad ,
		decrypt_i_pad,
		\sub1_data_reg_reg[104]/NET0131 ,
		_w995_,
		_w2537_
	);
	LUT3 #(
		.INIT('h04)
	) name1609 (
		\data_o[72]_pad ,
		decrypt_i_pad,
		_w995_,
		_w2538_
	);
	LUT4 #(
		.INIT('hce00)
	) name1610 (
		decrypt_i_pad,
		\sub1_data_reg_reg[72]/NET0131 ,
		_w995_,
		_w2240_,
		_w2539_
	);
	LUT2 #(
		.INIT('h4)
	) name1611 (
		_w2538_,
		_w2539_,
		_w2540_
	);
	LUT3 #(
		.INIT('h04)
	) name1612 (
		\data_o[8]_pad ,
		decrypt_i_pad,
		_w995_,
		_w2541_
	);
	LUT4 #(
		.INIT('hce00)
	) name1613 (
		decrypt_i_pad,
		\sub1_data_reg_reg[8]/NET0131 ,
		_w995_,
		_w2236_,
		_w2542_
	);
	LUT3 #(
		.INIT('h04)
	) name1614 (
		\data_o[40]_pad ,
		decrypt_i_pad,
		_w995_,
		_w2543_
	);
	LUT4 #(
		.INIT('hce00)
	) name1615 (
		decrypt_i_pad,
		\sub1_data_reg_reg[40]/NET0131 ,
		_w995_,
		_w2243_,
		_w2544_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name1616 (
		_w2541_,
		_w2542_,
		_w2543_,
		_w2544_,
		_w2545_
	);
	LUT4 #(
		.INIT('h1300)
	) name1617 (
		_w2233_,
		_w2540_,
		_w2537_,
		_w2545_,
		_w2546_
	);
	LUT4 #(
		.INIT('hf0b8)
	) name1618 (
		\data_o[96]_pad ,
		decrypt_i_pad,
		\sub1_data_reg_reg[96]/NET0131 ,
		_w995_,
		_w2547_
	);
	LUT3 #(
		.INIT('h04)
	) name1619 (
		\data_o[0]_pad ,
		decrypt_i_pad,
		_w995_,
		_w2548_
	);
	LUT4 #(
		.INIT('hce00)
	) name1620 (
		decrypt_i_pad,
		\sub1_data_reg_reg[0]/NET0131 ,
		_w995_,
		_w2236_,
		_w2549_
	);
	LUT2 #(
		.INIT('h4)
	) name1621 (
		_w2548_,
		_w2549_,
		_w2550_
	);
	LUT3 #(
		.INIT('h04)
	) name1622 (
		\data_o[32]_pad ,
		decrypt_i_pad,
		_w995_,
		_w2551_
	);
	LUT4 #(
		.INIT('hce00)
	) name1623 (
		decrypt_i_pad,
		\sub1_data_reg_reg[32]/NET0131 ,
		_w995_,
		_w2243_,
		_w2552_
	);
	LUT3 #(
		.INIT('h04)
	) name1624 (
		\data_o[64]_pad ,
		decrypt_i_pad,
		_w995_,
		_w2553_
	);
	LUT4 #(
		.INIT('hce00)
	) name1625 (
		decrypt_i_pad,
		\sub1_data_reg_reg[64]/NET0131 ,
		_w995_,
		_w2240_,
		_w2554_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name1626 (
		_w2551_,
		_w2552_,
		_w2553_,
		_w2554_,
		_w2555_
	);
	LUT4 #(
		.INIT('h1300)
	) name1627 (
		_w2233_,
		_w2550_,
		_w2547_,
		_w2555_,
		_w2556_
	);
	LUT3 #(
		.INIT('h69)
	) name1628 (
		_w2256_,
		_w2517_,
		_w2556_,
		_w2557_
	);
	LUT4 #(
		.INIT('h9669)
	) name1629 (
		_w2256_,
		_w2517_,
		_w2546_,
		_w2556_,
		_w2558_
	);
	LUT3 #(
		.INIT('h96)
	) name1630 (
		_w2309_,
		_w2330_,
		_w2372_,
		_w2559_
	);
	LUT2 #(
		.INIT('h6)
	) name1631 (
		_w2266_,
		_w2447_,
		_w2560_
	);
	LUT4 #(
		.INIT('hf0b8)
	) name1632 (
		\data_o[112]_pad ,
		decrypt_i_pad,
		\sub1_data_reg_reg[112]/NET0131 ,
		_w995_,
		_w2561_
	);
	LUT3 #(
		.INIT('h04)
	) name1633 (
		\data_o[16]_pad ,
		decrypt_i_pad,
		_w995_,
		_w2562_
	);
	LUT4 #(
		.INIT('hce00)
	) name1634 (
		decrypt_i_pad,
		\sub1_data_reg_reg[16]/NET0131 ,
		_w995_,
		_w2236_,
		_w2563_
	);
	LUT2 #(
		.INIT('h4)
	) name1635 (
		_w2562_,
		_w2563_,
		_w2564_
	);
	LUT3 #(
		.INIT('h04)
	) name1636 (
		\data_o[80]_pad ,
		decrypt_i_pad,
		_w995_,
		_w2565_
	);
	LUT4 #(
		.INIT('hce00)
	) name1637 (
		decrypt_i_pad,
		\sub1_data_reg_reg[80]/NET0131 ,
		_w995_,
		_w2240_,
		_w2566_
	);
	LUT3 #(
		.INIT('h04)
	) name1638 (
		\data_o[48]_pad ,
		decrypt_i_pad,
		_w995_,
		_w2567_
	);
	LUT4 #(
		.INIT('hce00)
	) name1639 (
		decrypt_i_pad,
		\sub1_data_reg_reg[48]/NET0131 ,
		_w995_,
		_w2243_,
		_w2568_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name1640 (
		_w2565_,
		_w2566_,
		_w2567_,
		_w2568_,
		_w2569_
	);
	LUT4 #(
		.INIT('h1300)
	) name1641 (
		_w2233_,
		_w2564_,
		_w2561_,
		_w2569_,
		_w2570_
	);
	LUT4 #(
		.INIT('hf0b8)
	) name1642 (
		\data_o[120]_pad ,
		decrypt_i_pad,
		\sub1_data_reg_reg[120]/NET0131 ,
		_w995_,
		_w2571_
	);
	LUT3 #(
		.INIT('h04)
	) name1643 (
		\data_o[56]_pad ,
		decrypt_i_pad,
		_w995_,
		_w2572_
	);
	LUT4 #(
		.INIT('hce00)
	) name1644 (
		decrypt_i_pad,
		\sub1_data_reg_reg[56]/NET0131 ,
		_w995_,
		_w2243_,
		_w2573_
	);
	LUT2 #(
		.INIT('h4)
	) name1645 (
		_w2572_,
		_w2573_,
		_w2574_
	);
	LUT3 #(
		.INIT('h04)
	) name1646 (
		\data_o[24]_pad ,
		decrypt_i_pad,
		_w995_,
		_w2575_
	);
	LUT4 #(
		.INIT('hce00)
	) name1647 (
		decrypt_i_pad,
		\sub1_data_reg_reg[24]/NET0131 ,
		_w995_,
		_w2236_,
		_w2576_
	);
	LUT3 #(
		.INIT('h04)
	) name1648 (
		\data_o[88]_pad ,
		decrypt_i_pad,
		_w995_,
		_w2577_
	);
	LUT4 #(
		.INIT('hce00)
	) name1649 (
		decrypt_i_pad,
		\sub1_data_reg_reg[88]/NET0131 ,
		_w995_,
		_w2240_,
		_w2578_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name1650 (
		_w2575_,
		_w2576_,
		_w2577_,
		_w2578_,
		_w2579_
	);
	LUT4 #(
		.INIT('h1300)
	) name1651 (
		_w2233_,
		_w2574_,
		_w2571_,
		_w2579_,
		_w2580_
	);
	LUT2 #(
		.INIT('h6)
	) name1652 (
		_w2570_,
		_w2580_,
		_w2581_
	);
	LUT3 #(
		.INIT('h69)
	) name1653 (
		_w2382_,
		_w2570_,
		_w2580_,
		_w2582_
	);
	LUT2 #(
		.INIT('h6)
	) name1654 (
		_w2560_,
		_w2582_,
		_w2583_
	);
	LUT4 #(
		.INIT('h2882)
	) name1655 (
		decrypt_i_pad,
		_w2558_,
		_w2559_,
		_w2583_,
		_w2584_
	);
	LUT4 #(
		.INIT('h6996)
	) name1656 (
		_w2437_,
		_w2495_,
		_w2536_,
		_w2584_,
		_w2585_
	);
	LUT3 #(
		.INIT('h2e)
	) name1657 (
		\mix1_data_reg_reg[107]/NET0131 ,
		_w2233_,
		_w2585_,
		_w2586_
	);
	LUT2 #(
		.INIT('h6)
	) name1658 (
		_w2505_,
		_w2528_,
		_w2587_
	);
	LUT3 #(
		.INIT('h96)
	) name1659 (
		_w2319_,
		_w2483_,
		_w2517_,
		_w2588_
	);
	LUT3 #(
		.INIT('h69)
	) name1660 (
		_w2329_,
		_w2447_,
		_w2472_,
		_w2589_
	);
	LUT4 #(
		.INIT('h6996)
	) name1661 (
		_w2309_,
		_w2330_,
		_w2588_,
		_w2589_,
		_w2590_
	);
	LUT4 #(
		.INIT('h8228)
	) name1662 (
		decrypt_i_pad,
		_w2383_,
		_w2587_,
		_w2590_,
		_w2591_
	);
	LUT4 #(
		.INIT('hf0b8)
	) name1663 (
		\data_o[107]_pad ,
		decrypt_i_pad,
		\sub1_data_reg_reg[107]/NET0131 ,
		_w995_,
		_w2592_
	);
	LUT3 #(
		.INIT('h04)
	) name1664 (
		\data_o[75]_pad ,
		decrypt_i_pad,
		_w995_,
		_w2593_
	);
	LUT4 #(
		.INIT('hce00)
	) name1665 (
		decrypt_i_pad,
		\sub1_data_reg_reg[75]/NET0131 ,
		_w995_,
		_w2240_,
		_w2594_
	);
	LUT2 #(
		.INIT('h4)
	) name1666 (
		_w2593_,
		_w2594_,
		_w2595_
	);
	LUT3 #(
		.INIT('h04)
	) name1667 (
		\data_o[11]_pad ,
		decrypt_i_pad,
		_w995_,
		_w2596_
	);
	LUT4 #(
		.INIT('hce00)
	) name1668 (
		decrypt_i_pad,
		\sub1_data_reg_reg[11]/NET0131 ,
		_w995_,
		_w2236_,
		_w2597_
	);
	LUT3 #(
		.INIT('h04)
	) name1669 (
		\data_o[43]_pad ,
		decrypt_i_pad,
		_w995_,
		_w2598_
	);
	LUT4 #(
		.INIT('hce00)
	) name1670 (
		decrypt_i_pad,
		\sub1_data_reg_reg[43]/NET0131 ,
		_w995_,
		_w2243_,
		_w2599_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name1671 (
		_w2596_,
		_w2597_,
		_w2598_,
		_w2599_,
		_w2600_
	);
	LUT4 #(
		.INIT('h1300)
	) name1672 (
		_w2233_,
		_w2595_,
		_w2592_,
		_w2600_,
		_w2601_
	);
	LUT2 #(
		.INIT('h9)
	) name1673 (
		_w2436_,
		_w2601_,
		_w2602_
	);
	LUT4 #(
		.INIT('h9669)
	) name1674 (
		_w2394_,
		_w2404_,
		_w2436_,
		_w2601_,
		_w2603_
	);
	LUT4 #(
		.INIT('h6996)
	) name1675 (
		_w2462_,
		_w2534_,
		_w2591_,
		_w2603_,
		_w2604_
	);
	LUT3 #(
		.INIT('h2e)
	) name1676 (
		\mix1_data_reg_reg[108]/NET0131 ,
		_w2233_,
		_w2604_,
		_w2605_
	);
	LUT2 #(
		.INIT('h9)
	) name1677 (
		_w2277_,
		_w2297_,
		_w2606_
	);
	LUT3 #(
		.INIT('h69)
	) name1678 (
		_w2277_,
		_w2297_,
		_w2462_,
		_w2607_
	);
	LUT3 #(
		.INIT('h69)
	) name1679 (
		_w2588_,
		_w2589_,
		_w2601_,
		_w2608_
	);
	LUT2 #(
		.INIT('h9)
	) name1680 (
		_w2246_,
		_w2505_,
		_w2609_
	);
	LUT4 #(
		.INIT('h9669)
	) name1681 (
		_w2246_,
		_w2266_,
		_w2447_,
		_w2505_,
		_w2610_
	);
	LUT3 #(
		.INIT('h96)
	) name1682 (
		_w2426_,
		_w2536_,
		_w2610_,
		_w2611_
	);
	LUT4 #(
		.INIT('hc66c)
	) name1683 (
		decrypt_i_pad,
		_w2607_,
		_w2608_,
		_w2611_,
		_w2612_
	);
	LUT2 #(
		.INIT('h9)
	) name1684 (
		_w2287_,
		_w2414_,
		_w2613_
	);
	LUT4 #(
		.INIT('he22e)
	) name1685 (
		\mix1_data_reg_reg[109]/NET0131 ,
		_w2233_,
		_w2612_,
		_w2613_,
		_w2614_
	);
	LUT2 #(
		.INIT('h9)
	) name1686 (
		_w2472_,
		_w2483_,
		_w2615_
	);
	LUT4 #(
		.INIT('h6996)
	) name1687 (
		_w2256_,
		_w2266_,
		_w2447_,
		_w2517_,
		_w2616_
	);
	LUT4 #(
		.INIT('h9669)
	) name1688 (
		_w2309_,
		_w2362_,
		_w2615_,
		_w2616_,
		_w2617_
	);
	LUT2 #(
		.INIT('h9)
	) name1689 (
		_w2546_,
		_w2570_,
		_w2618_
	);
	LUT2 #(
		.INIT('h9)
	) name1690 (
		_w2556_,
		_w2580_,
		_w2619_
	);
	LUT4 #(
		.INIT('h6996)
	) name1691 (
		_w2546_,
		_w2556_,
		_w2570_,
		_w2580_,
		_w2620_
	);
	LUT2 #(
		.INIT('h9)
	) name1692 (
		_w2426_,
		_w2601_,
		_w2621_
	);
	LUT4 #(
		.INIT('h7d82)
	) name1693 (
		decrypt_i_pad,
		_w2617_,
		_w2620_,
		_w2621_,
		_w2622_
	);
	LUT2 #(
		.INIT('h6)
	) name1694 (
		_w2436_,
		_w2530_,
		_w2623_
	);
	LUT4 #(
		.INIT('he22e)
	) name1695 (
		\mix1_data_reg_reg[115]/NET0131 ,
		_w2233_,
		_w2622_,
		_w2623_,
		_w2624_
	);
	LUT4 #(
		.INIT('h9669)
	) name1696 (
		_w2266_,
		_w2404_,
		_w2414_,
		_w2517_,
		_w2625_
	);
	LUT3 #(
		.INIT('h69)
	) name1697 (
		_w2462_,
		_w2495_,
		_w2601_,
		_w2626_
	);
	LUT4 #(
		.INIT('h8228)
	) name1698 (
		_w2233_,
		_w2384_,
		_w2625_,
		_w2626_,
		_w2627_
	);
	LUT2 #(
		.INIT('h1)
	) name1699 (
		\mix1_data_reg_reg[116]/NET0131 ,
		_w2233_,
		_w2628_
	);
	LUT2 #(
		.INIT('h1)
	) name1700 (
		_w2627_,
		_w2628_,
		_w2629_
	);
	LUT2 #(
		.INIT('h6)
	) name1701 (
		_w2394_,
		_w2414_,
		_w2630_
	);
	LUT3 #(
		.INIT('h96)
	) name1702 (
		_w2473_,
		_w2484_,
		_w2495_,
		_w2631_
	);
	LUT3 #(
		.INIT('h96)
	) name1703 (
		_w2436_,
		_w2506_,
		_w2530_,
		_w2632_
	);
	LUT4 #(
		.INIT('hc66c)
	) name1704 (
		decrypt_i_pad,
		_w2630_,
		_w2631_,
		_w2632_,
		_w2633_
	);
	LUT4 #(
		.INIT('h8228)
	) name1705 (
		_w2233_,
		_w2287_,
		_w2308_,
		_w2633_,
		_w2634_
	);
	LUT2 #(
		.INIT('h2)
	) name1706 (
		\mix1_data_reg_reg[117]/NET0131 ,
		_w2233_,
		_w2635_
	);
	LUT2 #(
		.INIT('he)
	) name1707 (
		_w2634_,
		_w2635_,
		_w2636_
	);
	LUT4 #(
		.INIT('h6996)
	) name1708 (
		_w2495_,
		_w2584_,
		_w2602_,
		_w2610_,
		_w2637_
	);
	LUT3 #(
		.INIT('h2e)
	) name1709 (
		\mix1_data_reg_reg[123]/NET0131 ,
		_w2233_,
		_w2637_,
		_w2638_
	);
	LUT3 #(
		.INIT('h96)
	) name1710 (
		_w2307_,
		_w2394_,
		_w2404_,
		_w2639_
	);
	LUT3 #(
		.INIT('h69)
	) name1711 (
		_w2426_,
		_w2588_,
		_w2589_,
		_w2640_
	);
	LUT3 #(
		.INIT('h96)
	) name1712 (
		_w2536_,
		_w2601_,
		_w2610_,
		_w2641_
	);
	LUT4 #(
		.INIT('h3993)
	) name1713 (
		decrypt_i_pad,
		_w2606_,
		_w2640_,
		_w2641_,
		_w2642_
	);
	LUT4 #(
		.INIT('he22e)
	) name1714 (
		\mix1_data_reg_reg[125]/NET0131 ,
		_w2233_,
		_w2639_,
		_w2642_,
		_w2643_
	);
	LUT2 #(
		.INIT('h9)
	) name1715 (
		_w2426_,
		_w2495_,
		_w2644_
	);
	LUT4 #(
		.INIT('h9669)
	) name1716 (
		_w2266_,
		_w2426_,
		_w2447_,
		_w2495_,
		_w2645_
	);
	LUT2 #(
		.INIT('h9)
	) name1717 (
		_w2630_,
		_w2645_,
		_w2646_
	);
	LUT4 #(
		.INIT('h8228)
	) name1718 (
		_w2233_,
		_w2462_,
		_w2591_,
		_w2646_,
		_w2647_
	);
	LUT2 #(
		.INIT('h1)
	) name1719 (
		\mix1_data_reg_reg[124]/NET0131 ,
		_w2233_,
		_w2648_
	);
	LUT2 #(
		.INIT('h1)
	) name1720 (
		_w2647_,
		_w2648_,
		_w2649_
	);
	LUT4 #(
		.INIT('h2ee2)
	) name1721 (
		\mix1_data_reg_reg[99]/NET0131 ,
		_w2233_,
		_w2507_,
		_w2622_,
		_w2650_
	);
	LUT3 #(
		.INIT('h69)
	) name1722 (
		_w2287_,
		_w2297_,
		_w2483_,
		_w2651_
	);
	LUT4 #(
		.INIT('h9669)
	) name1723 (
		_w2394_,
		_w2462_,
		_w2495_,
		_w2601_,
		_w2652_
	);
	LUT4 #(
		.INIT('h8228)
	) name1724 (
		decrypt_i_pad,
		_w2449_,
		_w2518_,
		_w2652_,
		_w2653_
	);
	LUT4 #(
		.INIT('h8228)
	) name1725 (
		_w2233_,
		_w2330_,
		_w2651_,
		_w2653_,
		_w2654_
	);
	LUT2 #(
		.INIT('h1)
	) name1726 (
		\mix1_data_reg_reg[102]/NET0131 ,
		_w2233_,
		_w2655_
	);
	LUT2 #(
		.INIT('h1)
	) name1727 (
		_w2654_,
		_w2655_,
		_w2656_
	);
	LUT3 #(
		.INIT('h28)
	) name1728 (
		decrypt_i_pad,
		_w2416_,
		_w2607_,
		_w2657_
	);
	LUT2 #(
		.INIT('h9)
	) name1729 (
		_w2518_,
		_w2589_,
		_w2658_
	);
	LUT4 #(
		.INIT('h2ee2)
	) name1730 (
		\mix1_data_reg_reg[103]/NET0131 ,
		_w2233_,
		_w2657_,
		_w2658_,
		_w2659_
	);
	LUT4 #(
		.INIT('h963c)
	) name1731 (
		decrypt_i_pad,
		_w2362_,
		_w2372_,
		_w2590_,
		_w2660_
	);
	LUT4 #(
		.INIT('he22e)
	) name1732 (
		\mix1_data_reg_reg[105]/NET0131 ,
		_w2233_,
		_w2558_,
		_w2660_,
		_w2661_
	);
	LUT3 #(
		.INIT('h69)
	) name1733 (
		_w2340_,
		_w2351_,
		_w2382_,
		_w2662_
	);
	LUT3 #(
		.INIT('h69)
	) name1734 (
		_w2266_,
		_w2517_,
		_w2546_,
		_w2663_
	);
	LUT3 #(
		.INIT('h69)
	) name1735 (
		_w2256_,
		_w2447_,
		_w2580_,
		_w2664_
	);
	LUT4 #(
		.INIT('h6006)
	) name1736 (
		_w2588_,
		_w2589_,
		_w2663_,
		_w2664_,
		_w2665_
	);
	LUT4 #(
		.INIT('h0990)
	) name1737 (
		_w2588_,
		_w2589_,
		_w2663_,
		_w2664_,
		_w2666_
	);
	LUT4 #(
		.INIT('h3339)
	) name1738 (
		decrypt_i_pad,
		_w2609_,
		_w2666_,
		_w2665_,
		_w2667_
	);
	LUT4 #(
		.INIT('h2ee2)
	) name1739 (
		\mix1_data_reg_reg[106]/NET0131 ,
		_w2233_,
		_w2662_,
		_w2667_,
		_w2668_
	);
	LUT2 #(
		.INIT('h6)
	) name1740 (
		_w2329_,
		_w2483_,
		_w2669_
	);
	LUT4 #(
		.INIT('h6900)
	) name1741 (
		_w2415_,
		_w2602_,
		_w2616_,
		_w2644_,
		_w2670_
	);
	LUT4 #(
		.INIT('h0096)
	) name1742 (
		_w2415_,
		_w2602_,
		_w2616_,
		_w2644_,
		_w2671_
	);
	LUT4 #(
		.INIT('h3339)
	) name1743 (
		decrypt_i_pad,
		_w2472_,
		_w2671_,
		_w2670_,
		_w2672_
	);
	LUT4 #(
		.INIT('h2882)
	) name1744 (
		_w2233_,
		_w2308_,
		_w2669_,
		_w2672_,
		_w2673_
	);
	LUT2 #(
		.INIT('h2)
	) name1745 (
		\mix1_data_reg_reg[110]/NET0131 ,
		_w2233_,
		_w2674_
	);
	LUT2 #(
		.INIT('he)
	) name1746 (
		_w2673_,
		_w2674_,
		_w2675_
	);
	LUT4 #(
		.INIT('h2882)
	) name1747 (
		decrypt_i_pad,
		_w2462_,
		_w2613_,
		_w2639_,
		_w2676_
	);
	LUT4 #(
		.INIT('h6996)
	) name1748 (
		_w2266_,
		_w2319_,
		_w2472_,
		_w2676_,
		_w2677_
	);
	LUT4 #(
		.INIT('h2ee2)
	) name1749 (
		\mix1_data_reg_reg[111]/NET0131 ,
		_w2233_,
		_w2448_,
		_w2677_,
		_w2678_
	);
	LUT4 #(
		.INIT('h8228)
	) name1750 (
		decrypt_i_pad,
		_w2267_,
		_w2309_,
		_w2330_,
		_w2679_
	);
	LUT2 #(
		.INIT('h9)
	) name1751 (
		_w2351_,
		_w2372_,
		_w2680_
	);
	LUT4 #(
		.INIT('h9669)
	) name1752 (
		_w2266_,
		_w2351_,
		_w2372_,
		_w2517_,
		_w2681_
	);
	LUT4 #(
		.INIT('h6996)
	) name1753 (
		_w2382_,
		_w2618_,
		_w2679_,
		_w2681_,
		_w2682_
	);
	LUT3 #(
		.INIT('h2e)
	) name1754 (
		\mix1_data_reg_reg[113]/NET0131 ,
		_w2233_,
		_w2682_,
		_w2683_
	);
	LUT3 #(
		.INIT('h69)
	) name1755 (
		_w2340_,
		_w2361_,
		_w2382_,
		_w2684_
	);
	LUT2 #(
		.INIT('h9)
	) name1756 (
		_w2556_,
		_w2570_,
		_w2685_
	);
	LUT4 #(
		.INIT('h0660)
	) name1757 (
		_w2473_,
		_w2484_,
		_w2616_,
		_w2685_,
		_w2686_
	);
	LUT4 #(
		.INIT('h9009)
	) name1758 (
		_w2473_,
		_w2484_,
		_w2616_,
		_w2685_,
		_w2687_
	);
	LUT4 #(
		.INIT('h3339)
	) name1759 (
		decrypt_i_pad,
		_w2587_,
		_w2687_,
		_w2686_,
		_w2688_
	);
	LUT4 #(
		.INIT('he22e)
	) name1760 (
		\mix1_data_reg_reg[114]/NET0131 ,
		_w2233_,
		_w2684_,
		_w2688_,
		_w2689_
	);
	LUT3 #(
		.INIT('h69)
	) name1761 (
		_w2277_,
		_w2307_,
		_w2319_,
		_w2690_
	);
	LUT4 #(
		.INIT('h8228)
	) name1762 (
		_w2233_,
		_w2473_,
		_w2653_,
		_w2690_,
		_w2691_
	);
	LUT2 #(
		.INIT('h1)
	) name1763 (
		\mix1_data_reg_reg[118]/NET0131 ,
		_w2233_,
		_w2692_
	);
	LUT2 #(
		.INIT('h1)
	) name1764 (
		_w2691_,
		_w2692_,
		_w2693_
	);
	LUT2 #(
		.INIT('h9)
	) name1765 (
		_w2448_,
		_w2588_,
		_w2694_
	);
	LUT4 #(
		.INIT('he22e)
	) name1766 (
		\mix1_data_reg_reg[119]/NET0131 ,
		_w2233_,
		_w2657_,
		_w2694_,
		_w2695_
	);
	LUT4 #(
		.INIT('h69c3)
	) name1767 (
		decrypt_i_pad,
		_w2362_,
		_w2583_,
		_w2590_,
		_w2696_
	);
	LUT3 #(
		.INIT('he2)
	) name1768 (
		\mix1_data_reg_reg[121]/NET0131 ,
		_w2233_,
		_w2696_,
		_w2697_
	);
	LUT2 #(
		.INIT('h9)
	) name1769 (
		_w2361_,
		_w2372_,
		_w2698_
	);
	LUT4 #(
		.INIT('h3339)
	) name1770 (
		decrypt_i_pad,
		_w2535_,
		_w2666_,
		_w2665_,
		_w2699_
	);
	LUT4 #(
		.INIT('h2882)
	) name1771 (
		_w2233_,
		_w2246_,
		_w2698_,
		_w2699_,
		_w2700_
	);
	LUT2 #(
		.INIT('h2)
	) name1772 (
		\mix1_data_reg_reg[122]/NET0131 ,
		_w2233_,
		_w2701_
	);
	LUT2 #(
		.INIT('he)
	) name1773 (
		_w2700_,
		_w2701_,
		_w2702_
	);
	LUT4 #(
		.INIT('h6996)
	) name1774 (
		_w2277_,
		_w2287_,
		_w2319_,
		_w2483_,
		_w2703_
	);
	LUT4 #(
		.INIT('h2ee2)
	) name1775 (
		\mix1_data_reg_reg[126]/NET0131 ,
		_w2233_,
		_w2672_,
		_w2703_,
		_w2704_
	);
	LUT4 #(
		.INIT('h6996)
	) name1776 (
		_w2266_,
		_w2534_,
		_w2669_,
		_w2676_,
		_w2705_
	);
	LUT3 #(
		.INIT('he2)
	) name1777 (
		\mix1_data_reg_reg[127]/NET0131 ,
		_w2233_,
		_w2705_,
		_w2706_
	);
	LUT4 #(
		.INIT('h2ee2)
	) name1778 (
		\mix1_data_reg_reg[35]/NET0131 ,
		_w2243_,
		_w2507_,
		_w2622_,
		_w2707_
	);
	LUT4 #(
		.INIT('he22e)
	) name1779 (
		\mix1_data_reg_reg[36]/NET0131 ,
		_w2243_,
		_w2384_,
		_w2450_,
		_w2708_
	);
	LUT4 #(
		.INIT('he22e)
	) name1780 (
		\mix1_data_reg_reg[37]/NET0131 ,
		_w2243_,
		_w2452_,
		_w2532_,
		_w2709_
	);
	LUT3 #(
		.INIT('h2e)
	) name1781 (
		\mix1_data_reg_reg[43]/NET0131 ,
		_w2243_,
		_w2585_,
		_w2710_
	);
	LUT3 #(
		.INIT('h2e)
	) name1782 (
		\mix1_data_reg_reg[44]/NET0131 ,
		_w2243_,
		_w2604_,
		_w2711_
	);
	LUT4 #(
		.INIT('he22e)
	) name1783 (
		\mix1_data_reg_reg[45]/NET0131 ,
		_w2243_,
		_w2612_,
		_w2613_,
		_w2712_
	);
	LUT4 #(
		.INIT('he22e)
	) name1784 (
		\mix1_data_reg_reg[51]/NET0131 ,
		_w2243_,
		_w2622_,
		_w2623_,
		_w2713_
	);
	LUT4 #(
		.INIT('h8228)
	) name1785 (
		_w2243_,
		_w2287_,
		_w2308_,
		_w2633_,
		_w2714_
	);
	LUT3 #(
		.INIT('h8a)
	) name1786 (
		\mix1_data_reg_reg[53]/NET0131 ,
		\mix1_state_reg[0]/NET0131 ,
		\mix1_state_reg[1]/NET0131 ,
		_w2715_
	);
	LUT2 #(
		.INIT('he)
	) name1787 (
		_w2714_,
		_w2715_,
		_w2716_
	);
	LUT4 #(
		.INIT('h8228)
	) name1788 (
		_w2243_,
		_w2384_,
		_w2625_,
		_w2626_,
		_w2717_
	);
	LUT3 #(
		.INIT('h45)
	) name1789 (
		\mix1_data_reg_reg[52]/NET0131 ,
		\mix1_state_reg[0]/NET0131 ,
		\mix1_state_reg[1]/NET0131 ,
		_w2718_
	);
	LUT2 #(
		.INIT('h1)
	) name1790 (
		_w2717_,
		_w2718_,
		_w2719_
	);
	LUT3 #(
		.INIT('h2e)
	) name1791 (
		\mix1_data_reg_reg[59]/NET0131 ,
		_w2243_,
		_w2637_,
		_w2720_
	);
	LUT4 #(
		.INIT('h8228)
	) name1792 (
		_w2243_,
		_w2462_,
		_w2591_,
		_w2646_,
		_w2721_
	);
	LUT3 #(
		.INIT('h45)
	) name1793 (
		\mix1_data_reg_reg[60]/NET0131 ,
		\mix1_state_reg[0]/NET0131 ,
		\mix1_state_reg[1]/NET0131 ,
		_w2722_
	);
	LUT2 #(
		.INIT('h1)
	) name1794 (
		_w2721_,
		_w2722_,
		_w2723_
	);
	LUT4 #(
		.INIT('he22e)
	) name1795 (
		\mix1_data_reg_reg[61]/NET0131 ,
		_w2243_,
		_w2639_,
		_w2642_,
		_w2724_
	);
	LUT4 #(
		.INIT('he22e)
	) name1796 (
		\mix1_data_reg_reg[68]/NET0131 ,
		_w2240_,
		_w2384_,
		_w2450_,
		_w2725_
	);
	LUT4 #(
		.INIT('he22e)
	) name1797 (
		\mix1_data_reg_reg[69]/NET0131 ,
		_w2240_,
		_w2452_,
		_w2532_,
		_w2726_
	);
	LUT4 #(
		.INIT('h2ee2)
	) name1798 (
		\mix1_data_reg_reg[67]/NET0131 ,
		_w2240_,
		_w2507_,
		_w2622_,
		_w2727_
	);
	LUT3 #(
		.INIT('h2e)
	) name1799 (
		\mix1_data_reg_reg[75]/NET0131 ,
		_w2240_,
		_w2585_,
		_w2728_
	);
	LUT3 #(
		.INIT('h2e)
	) name1800 (
		\mix1_data_reg_reg[76]/NET0131 ,
		_w2240_,
		_w2604_,
		_w2729_
	);
	LUT4 #(
		.INIT('he22e)
	) name1801 (
		\mix1_data_reg_reg[77]/NET0131 ,
		_w2240_,
		_w2612_,
		_w2613_,
		_w2730_
	);
	LUT4 #(
		.INIT('h8228)
	) name1802 (
		_w2240_,
		_w2384_,
		_w2625_,
		_w2626_,
		_w2731_
	);
	LUT3 #(
		.INIT('h51)
	) name1803 (
		\mix1_data_reg_reg[84]/NET0131 ,
		\mix1_state_reg[0]/NET0131 ,
		\mix1_state_reg[1]/NET0131 ,
		_w2732_
	);
	LUT2 #(
		.INIT('h1)
	) name1804 (
		_w2731_,
		_w2732_,
		_w2733_
	);
	LUT4 #(
		.INIT('h8228)
	) name1805 (
		_w2240_,
		_w2287_,
		_w2308_,
		_w2633_,
		_w2734_
	);
	LUT3 #(
		.INIT('ha2)
	) name1806 (
		\mix1_data_reg_reg[85]/NET0131 ,
		\mix1_state_reg[0]/NET0131 ,
		\mix1_state_reg[1]/NET0131 ,
		_w2735_
	);
	LUT2 #(
		.INIT('he)
	) name1807 (
		_w2734_,
		_w2735_,
		_w2736_
	);
	LUT4 #(
		.INIT('he22e)
	) name1808 (
		\mix1_data_reg_reg[83]/NET0131 ,
		_w2240_,
		_w2622_,
		_w2623_,
		_w2737_
	);
	LUT4 #(
		.INIT('h8228)
	) name1809 (
		_w2240_,
		_w2462_,
		_w2591_,
		_w2646_,
		_w2738_
	);
	LUT3 #(
		.INIT('h51)
	) name1810 (
		\mix1_data_reg_reg[92]/NET0131 ,
		\mix1_state_reg[0]/NET0131 ,
		\mix1_state_reg[1]/NET0131 ,
		_w2739_
	);
	LUT2 #(
		.INIT('h1)
	) name1811 (
		_w2738_,
		_w2739_,
		_w2740_
	);
	LUT3 #(
		.INIT('h2e)
	) name1812 (
		\mix1_data_reg_reg[91]/NET0131 ,
		_w2240_,
		_w2637_,
		_w2741_
	);
	LUT4 #(
		.INIT('he22e)
	) name1813 (
		\mix1_data_reg_reg[93]/NET0131 ,
		_w2240_,
		_w2639_,
		_w2642_,
		_w2742_
	);
	LUT4 #(
		.INIT('h3339)
	) name1814 (
		decrypt_i_pad,
		_w2529_,
		_w2687_,
		_w2686_,
		_w2743_
	);
	LUT4 #(
		.INIT('h2882)
	) name1815 (
		_w2233_,
		_w2505_,
		_w2680_,
		_w2743_,
		_w2744_
	);
	LUT2 #(
		.INIT('h2)
	) name1816 (
		\mix1_data_reg_reg[98]/NET0131 ,
		_w2233_,
		_w2745_
	);
	LUT2 #(
		.INIT('he)
	) name1817 (
		_w2744_,
		_w2745_,
		_w2746_
	);
	LUT4 #(
		.INIT('h9669)
	) name1818 (
		_w2256_,
		_w2361_,
		_w2372_,
		_w2447_,
		_w2747_
	);
	LUT4 #(
		.INIT('h6996)
	) name1819 (
		_w2382_,
		_w2619_,
		_w2679_,
		_w2747_,
		_w2748_
	);
	LUT3 #(
		.INIT('h2e)
	) name1820 (
		\mix1_data_reg_reg[97]/NET0131 ,
		_w2233_,
		_w2748_,
		_w2749_
	);
	LUT4 #(
		.INIT('ha222)
	) name1821 (
		\addroundkey_round_reg[3]/NET0131 ,
		\ks1_ready_o_reg/NET0131 ,
		_w932_,
		_w933_,
		_w2750_
	);
	LUT4 #(
		.INIT('h7f80)
	) name1822 (
		\addroundkey_round_reg[0]/NET0131 ,
		\addroundkey_round_reg[1]/NET0131 ,
		\addroundkey_round_reg[2]/NET0131 ,
		\addroundkey_round_reg[3]/NET0131 ,
		_w2751_
	);
	LUT4 #(
		.INIT('h2a00)
	) name1823 (
		\ks1_ready_o_reg/NET0131 ,
		_w932_,
		_w933_,
		_w2751_,
		_w2752_
	);
	LUT3 #(
		.INIT('h80)
	) name1824 (
		\addroundkey_round_reg[3]/NET0131 ,
		\addroundkey_start_i_reg/NET0131 ,
		_w930_,
		_w2753_
	);
	LUT4 #(
		.INIT('h00ab)
	) name1825 (
		\addroundkey_start_i_reg/NET0131 ,
		_w2750_,
		_w2752_,
		_w2753_,
		_w2754_
	);
	LUT4 #(
		.INIT('ha222)
	) name1826 (
		\addroundkey_round_reg[1]/NET0131 ,
		\ks1_ready_o_reg/NET0131 ,
		_w932_,
		_w933_,
		_w2755_
	);
	LUT2 #(
		.INIT('h6)
	) name1827 (
		\addroundkey_round_reg[0]/NET0131 ,
		\addroundkey_round_reg[1]/NET0131 ,
		_w2756_
	);
	LUT4 #(
		.INIT('h2a00)
	) name1828 (
		\ks1_ready_o_reg/NET0131 ,
		_w932_,
		_w933_,
		_w2756_,
		_w2757_
	);
	LUT3 #(
		.INIT('h80)
	) name1829 (
		\addroundkey_round_reg[1]/NET0131 ,
		\addroundkey_start_i_reg/NET0131 ,
		_w930_,
		_w2758_
	);
	LUT4 #(
		.INIT('h00ab)
	) name1830 (
		\addroundkey_start_i_reg/NET0131 ,
		_w2755_,
		_w2757_,
		_w2758_,
		_w2759_
	);
	LUT3 #(
		.INIT('h21)
	) name1831 (
		\addroundkey_round_reg[0]/NET0131 ,
		_w938_,
		_w945_,
		_w2760_
	);
	LUT4 #(
		.INIT('ha222)
	) name1832 (
		\addroundkey_round_reg[2]/NET0131 ,
		\ks1_ready_o_reg/NET0131 ,
		_w932_,
		_w933_,
		_w2761_
	);
	LUT3 #(
		.INIT('h78)
	) name1833 (
		\addroundkey_round_reg[0]/NET0131 ,
		\addroundkey_round_reg[1]/NET0131 ,
		\addroundkey_round_reg[2]/NET0131 ,
		_w2762_
	);
	LUT4 #(
		.INIT('h2a00)
	) name1834 (
		\ks1_ready_o_reg/NET0131 ,
		_w932_,
		_w933_,
		_w2762_,
		_w2763_
	);
	LUT3 #(
		.INIT('h80)
	) name1835 (
		\addroundkey_round_reg[2]/NET0131 ,
		\addroundkey_start_i_reg/NET0131 ,
		_w930_,
		_w2764_
	);
	LUT4 #(
		.INIT('h00ab)
	) name1836 (
		\addroundkey_start_i_reg/NET0131 ,
		_w2761_,
		_w2763_,
		_w2764_,
		_w2765_
	);
	LUT4 #(
		.INIT('hebf7)
	) name1837 (
		_w2754_,
		_w2759_,
		_w2760_,
		_w2765_,
		_w2766_
	);
	LUT4 #(
		.INIT('haaac)
	) name1838 (
		\key_i[124]_pad ,
		\ks1_key_reg_reg[124]/NET0131 ,
		_w938_,
		_w986_,
		_w2767_
	);
	LUT3 #(
		.INIT('h69)
	) name1839 (
		\ks1_col_reg[28]/NET0131 ,
		_w2766_,
		_w2767_,
		_w2768_
	);
	LUT4 #(
		.INIT('haaac)
	) name1840 (
		\key_i[92]_pad ,
		\ks1_key_reg_reg[92]/NET0131 ,
		_w938_,
		_w986_,
		_w2769_
	);
	LUT4 #(
		.INIT('h9669)
	) name1841 (
		\ks1_col_reg[28]/NET0131 ,
		_w2766_,
		_w2767_,
		_w2769_,
		_w2770_
	);
	LUT4 #(
		.INIT('haaac)
	) name1842 (
		\key_i[60]_pad ,
		\ks1_key_reg_reg[60]/NET0131 ,
		_w938_,
		_w986_,
		_w2771_
	);
	LUT4 #(
		.INIT('h2ee2)
	) name1843 (
		\ks1_key_reg_reg[60]/NET0131 ,
		_w929_,
		_w2770_,
		_w2771_,
		_w2772_
	);
	LUT3 #(
		.INIT('h69)
	) name1844 (
		_w1091_,
		_w2770_,
		_w2771_,
		_w2773_
	);
	LUT3 #(
		.INIT('hc4)
	) name1845 (
		\sub1_ready_o_reg/NET0131 ,
		_w1054_,
		_w2230_,
		_w2774_
	);
	LUT2 #(
		.INIT('h4)
	) name1846 (
		decrypt_i_pad,
		\mix1_ready_o_reg/NET0131 ,
		_w2775_
	);
	LUT2 #(
		.INIT('h8)
	) name1847 (
		decrypt_i_pad,
		\sub1_ready_o_reg/NET0131 ,
		_w2776_
	);
	LUT4 #(
		.INIT('haab8)
	) name1848 (
		\data_i[112]_pad ,
		decrypt_i_pad,
		\mix1_data_o_reg_reg[112]/NET0131 ,
		_w930_,
		_w2777_
	);
	LUT4 #(
		.INIT('haba8)
	) name1849 (
		\sub1_data_reg_reg[112]/NET0131 ,
		_w996_,
		_w2776_,
		_w2777_,
		_w2778_
	);
	LUT4 #(
		.INIT('h404c)
	) name1850 (
		\mix1_data_o_reg_reg[112]/NET0131 ,
		_w2774_,
		_w2775_,
		_w2778_,
		_w2779_
	);
	LUT4 #(
		.INIT('h0545)
	) name1851 (
		\sub1_data_reg_reg[112]/NET0131 ,
		\sub1_ready_o_reg/NET0131 ,
		_w1054_,
		_w2230_,
		_w2780_
	);
	LUT4 #(
		.INIT('h1015)
	) name1852 (
		\state_reg/NET0131 ,
		\sub1_data_reg_reg[112]/NET0131 ,
		_w996_,
		_w2777_,
		_w2781_
	);
	LUT4 #(
		.INIT('h0057)
	) name1853 (
		\state_reg/NET0131 ,
		_w2779_,
		_w2780_,
		_w2781_,
		_w2782_
	);
	LUT3 #(
		.INIT('h48)
	) name1854 (
		\key_i[112]_pad ,
		_w931_,
		_w2782_,
		_w2783_
	);
	LUT3 #(
		.INIT('hc4)
	) name1855 (
		\addroundkey_start_i_reg/NET0131 ,
		\ks1_ready_o_reg/NET0131 ,
		_w930_,
		_w2784_
	);
	LUT2 #(
		.INIT('h8)
	) name1856 (
		_w934_,
		_w2784_,
		_w2785_
	);
	LUT4 #(
		.INIT('h3222)
	) name1857 (
		\data_o[112]_pad ,
		_w931_,
		_w934_,
		_w2784_,
		_w2786_
	);
	LUT4 #(
		.INIT('h6f00)
	) name1858 (
		\ks1_key_reg_reg[112]/NET0131 ,
		_w2782_,
		_w2785_,
		_w2786_,
		_w2787_
	);
	LUT2 #(
		.INIT('he)
	) name1859 (
		_w2783_,
		_w2787_,
		_w2788_
	);
	LUT4 #(
		.INIT('h5547)
	) name1860 (
		\data_i[61]_pad ,
		decrypt_i_pad,
		\mix1_data_o_reg_reg[61]/NET0131 ,
		_w930_,
		_w2789_
	);
	LUT4 #(
		.INIT('ha8ab)
	) name1861 (
		\sub1_data_reg_reg[61]/NET0131 ,
		_w996_,
		_w2776_,
		_w2789_,
		_w2790_
	);
	LUT4 #(
		.INIT('h404c)
	) name1862 (
		\mix1_data_o_reg_reg[61]/NET0131 ,
		_w2774_,
		_w2775_,
		_w2790_,
		_w2791_
	);
	LUT4 #(
		.INIT('h0545)
	) name1863 (
		\sub1_data_reg_reg[61]/NET0131 ,
		\sub1_ready_o_reg/NET0131 ,
		_w1054_,
		_w2230_,
		_w2792_
	);
	LUT4 #(
		.INIT('h1510)
	) name1864 (
		\state_reg/NET0131 ,
		\sub1_data_reg_reg[61]/NET0131 ,
		_w996_,
		_w2789_,
		_w2793_
	);
	LUT4 #(
		.INIT('h0057)
	) name1865 (
		\state_reg/NET0131 ,
		_w2791_,
		_w2792_,
		_w2793_,
		_w2794_
	);
	LUT3 #(
		.INIT('h48)
	) name1866 (
		\key_i[61]_pad ,
		_w931_,
		_w2794_,
		_w2795_
	);
	LUT4 #(
		.INIT('h3222)
	) name1867 (
		\data_o[61]_pad ,
		_w931_,
		_w934_,
		_w2784_,
		_w2796_
	);
	LUT4 #(
		.INIT('h7b00)
	) name1868 (
		\ks1_key_reg_reg[61]/NET0131 ,
		_w2785_,
		_w2794_,
		_w2796_,
		_w2797_
	);
	LUT2 #(
		.INIT('he)
	) name1869 (
		_w2795_,
		_w2797_,
		_w2798_
	);
	LUT4 #(
		.INIT('haab8)
	) name1870 (
		\data_i[19]_pad ,
		decrypt_i_pad,
		\mix1_data_o_reg_reg[19]/NET0131 ,
		_w930_,
		_w2799_
	);
	LUT4 #(
		.INIT('haba8)
	) name1871 (
		\sub1_data_reg_reg[19]/NET0131 ,
		_w996_,
		_w2776_,
		_w2799_,
		_w2800_
	);
	LUT4 #(
		.INIT('h404c)
	) name1872 (
		\mix1_data_o_reg_reg[19]/NET0131 ,
		_w2774_,
		_w2775_,
		_w2800_,
		_w2801_
	);
	LUT4 #(
		.INIT('h0545)
	) name1873 (
		\sub1_data_reg_reg[19]/NET0131 ,
		\sub1_ready_o_reg/NET0131 ,
		_w1054_,
		_w2230_,
		_w2802_
	);
	LUT4 #(
		.INIT('h1015)
	) name1874 (
		\state_reg/NET0131 ,
		\sub1_data_reg_reg[19]/NET0131 ,
		_w996_,
		_w2799_,
		_w2803_
	);
	LUT4 #(
		.INIT('h0057)
	) name1875 (
		\state_reg/NET0131 ,
		_w2801_,
		_w2802_,
		_w2803_,
		_w2804_
	);
	LUT3 #(
		.INIT('h48)
	) name1876 (
		\key_i[19]_pad ,
		_w931_,
		_w2804_,
		_w2805_
	);
	LUT4 #(
		.INIT('h3222)
	) name1877 (
		\data_o[19]_pad ,
		_w931_,
		_w934_,
		_w2784_,
		_w2806_
	);
	LUT4 #(
		.INIT('h7b00)
	) name1878 (
		\ks1_key_reg_reg[19]/NET0131 ,
		_w2785_,
		_w2804_,
		_w2806_,
		_w2807_
	);
	LUT2 #(
		.INIT('he)
	) name1879 (
		_w2805_,
		_w2807_,
		_w2808_
	);
	LUT4 #(
		.INIT('h5547)
	) name1880 (
		\data_i[62]_pad ,
		decrypt_i_pad,
		\mix1_data_o_reg_reg[62]/NET0131 ,
		_w930_,
		_w2809_
	);
	LUT4 #(
		.INIT('ha8ab)
	) name1881 (
		\sub1_data_reg_reg[62]/NET0131 ,
		_w996_,
		_w2776_,
		_w2809_,
		_w2810_
	);
	LUT4 #(
		.INIT('h404c)
	) name1882 (
		\mix1_data_o_reg_reg[62]/NET0131 ,
		_w2774_,
		_w2775_,
		_w2810_,
		_w2811_
	);
	LUT4 #(
		.INIT('h0545)
	) name1883 (
		\sub1_data_reg_reg[62]/NET0131 ,
		\sub1_ready_o_reg/NET0131 ,
		_w1054_,
		_w2230_,
		_w2812_
	);
	LUT4 #(
		.INIT('h1510)
	) name1884 (
		\state_reg/NET0131 ,
		\sub1_data_reg_reg[62]/NET0131 ,
		_w996_,
		_w2809_,
		_w2813_
	);
	LUT4 #(
		.INIT('h0057)
	) name1885 (
		\state_reg/NET0131 ,
		_w2811_,
		_w2812_,
		_w2813_,
		_w2814_
	);
	LUT3 #(
		.INIT('h48)
	) name1886 (
		\key_i[62]_pad ,
		_w931_,
		_w2814_,
		_w2815_
	);
	LUT4 #(
		.INIT('h3222)
	) name1887 (
		\data_o[62]_pad ,
		_w931_,
		_w934_,
		_w2784_,
		_w2816_
	);
	LUT4 #(
		.INIT('h7b00)
	) name1888 (
		\ks1_key_reg_reg[62]/NET0131 ,
		_w2785_,
		_w2814_,
		_w2816_,
		_w2817_
	);
	LUT2 #(
		.INIT('he)
	) name1889 (
		_w2815_,
		_w2817_,
		_w2818_
	);
	LUT4 #(
		.INIT('h5547)
	) name1890 (
		\data_i[63]_pad ,
		decrypt_i_pad,
		\mix1_data_o_reg_reg[63]/NET0131 ,
		_w930_,
		_w2819_
	);
	LUT4 #(
		.INIT('ha8ab)
	) name1891 (
		\sub1_data_reg_reg[63]/NET0131 ,
		_w996_,
		_w2776_,
		_w2819_,
		_w2820_
	);
	LUT4 #(
		.INIT('h404c)
	) name1892 (
		\mix1_data_o_reg_reg[63]/NET0131 ,
		_w2774_,
		_w2775_,
		_w2820_,
		_w2821_
	);
	LUT4 #(
		.INIT('h0545)
	) name1893 (
		\sub1_data_reg_reg[63]/NET0131 ,
		\sub1_ready_o_reg/NET0131 ,
		_w1054_,
		_w2230_,
		_w2822_
	);
	LUT4 #(
		.INIT('h1510)
	) name1894 (
		\state_reg/NET0131 ,
		\sub1_data_reg_reg[63]/NET0131 ,
		_w996_,
		_w2819_,
		_w2823_
	);
	LUT4 #(
		.INIT('h0057)
	) name1895 (
		\state_reg/NET0131 ,
		_w2821_,
		_w2822_,
		_w2823_,
		_w2824_
	);
	LUT3 #(
		.INIT('h48)
	) name1896 (
		\key_i[63]_pad ,
		_w931_,
		_w2824_,
		_w2825_
	);
	LUT4 #(
		.INIT('h3222)
	) name1897 (
		\data_o[63]_pad ,
		_w931_,
		_w934_,
		_w2784_,
		_w2826_
	);
	LUT4 #(
		.INIT('h7b00)
	) name1898 (
		\ks1_key_reg_reg[63]/NET0131 ,
		_w2785_,
		_w2824_,
		_w2826_,
		_w2827_
	);
	LUT2 #(
		.INIT('he)
	) name1899 (
		_w2825_,
		_w2827_,
		_w2828_
	);
	LUT4 #(
		.INIT('h5547)
	) name1900 (
		\data_i[1]_pad ,
		decrypt_i_pad,
		\mix1_data_o_reg_reg[1]/NET0131 ,
		_w930_,
		_w2829_
	);
	LUT4 #(
		.INIT('ha8ab)
	) name1901 (
		\sub1_data_reg_reg[1]/NET0131 ,
		_w996_,
		_w2776_,
		_w2829_,
		_w2830_
	);
	LUT4 #(
		.INIT('h404c)
	) name1902 (
		\mix1_data_o_reg_reg[1]/NET0131 ,
		_w2774_,
		_w2775_,
		_w2830_,
		_w2831_
	);
	LUT4 #(
		.INIT('h0545)
	) name1903 (
		\sub1_data_reg_reg[1]/NET0131 ,
		\sub1_ready_o_reg/NET0131 ,
		_w1054_,
		_w2230_,
		_w2832_
	);
	LUT4 #(
		.INIT('h1510)
	) name1904 (
		\state_reg/NET0131 ,
		\sub1_data_reg_reg[1]/NET0131 ,
		_w996_,
		_w2829_,
		_w2833_
	);
	LUT4 #(
		.INIT('h0057)
	) name1905 (
		\state_reg/NET0131 ,
		_w2831_,
		_w2832_,
		_w2833_,
		_w2834_
	);
	LUT3 #(
		.INIT('h48)
	) name1906 (
		\key_i[1]_pad ,
		_w931_,
		_w2834_,
		_w2835_
	);
	LUT4 #(
		.INIT('h3222)
	) name1907 (
		\data_o[1]_pad ,
		_w931_,
		_w934_,
		_w2784_,
		_w2836_
	);
	LUT4 #(
		.INIT('h7b00)
	) name1908 (
		\ks1_key_reg_reg[1]/NET0131 ,
		_w2785_,
		_w2834_,
		_w2836_,
		_w2837_
	);
	LUT2 #(
		.INIT('he)
	) name1909 (
		_w2835_,
		_w2837_,
		_w2838_
	);
	LUT4 #(
		.INIT('haab8)
	) name1910 (
		\data_i[64]_pad ,
		decrypt_i_pad,
		\mix1_data_o_reg_reg[64]/NET0131 ,
		_w930_,
		_w2839_
	);
	LUT4 #(
		.INIT('haba8)
	) name1911 (
		\sub1_data_reg_reg[64]/NET0131 ,
		_w996_,
		_w2776_,
		_w2839_,
		_w2840_
	);
	LUT4 #(
		.INIT('h404c)
	) name1912 (
		\mix1_data_o_reg_reg[64]/NET0131 ,
		_w2774_,
		_w2775_,
		_w2840_,
		_w2841_
	);
	LUT4 #(
		.INIT('h0545)
	) name1913 (
		\sub1_data_reg_reg[64]/NET0131 ,
		\sub1_ready_o_reg/NET0131 ,
		_w1054_,
		_w2230_,
		_w2842_
	);
	LUT4 #(
		.INIT('h1015)
	) name1914 (
		\state_reg/NET0131 ,
		\sub1_data_reg_reg[64]/NET0131 ,
		_w996_,
		_w2839_,
		_w2843_
	);
	LUT4 #(
		.INIT('h0057)
	) name1915 (
		\state_reg/NET0131 ,
		_w2841_,
		_w2842_,
		_w2843_,
		_w2844_
	);
	LUT3 #(
		.INIT('h48)
	) name1916 (
		\key_i[64]_pad ,
		_w931_,
		_w2844_,
		_w2845_
	);
	LUT4 #(
		.INIT('h3222)
	) name1917 (
		\data_o[64]_pad ,
		_w931_,
		_w934_,
		_w2784_,
		_w2846_
	);
	LUT4 #(
		.INIT('h7b00)
	) name1918 (
		\ks1_key_reg_reg[64]/NET0131 ,
		_w2785_,
		_w2844_,
		_w2846_,
		_w2847_
	);
	LUT2 #(
		.INIT('he)
	) name1919 (
		_w2845_,
		_w2847_,
		_w2848_
	);
	LUT4 #(
		.INIT('haab8)
	) name1920 (
		\data_i[101]_pad ,
		decrypt_i_pad,
		\mix1_data_o_reg_reg[101]/NET0131 ,
		_w930_,
		_w2849_
	);
	LUT4 #(
		.INIT('haba8)
	) name1921 (
		\sub1_data_reg_reg[101]/NET0131 ,
		_w996_,
		_w2776_,
		_w2849_,
		_w2850_
	);
	LUT4 #(
		.INIT('h404c)
	) name1922 (
		\mix1_data_o_reg_reg[101]/NET0131 ,
		_w2774_,
		_w2775_,
		_w2850_,
		_w2851_
	);
	LUT4 #(
		.INIT('h0545)
	) name1923 (
		\sub1_data_reg_reg[101]/NET0131 ,
		\sub1_ready_o_reg/NET0131 ,
		_w1054_,
		_w2230_,
		_w2852_
	);
	LUT4 #(
		.INIT('h1015)
	) name1924 (
		\state_reg/NET0131 ,
		\sub1_data_reg_reg[101]/NET0131 ,
		_w996_,
		_w2849_,
		_w2853_
	);
	LUT4 #(
		.INIT('h0057)
	) name1925 (
		\state_reg/NET0131 ,
		_w2851_,
		_w2852_,
		_w2853_,
		_w2854_
	);
	LUT3 #(
		.INIT('h48)
	) name1926 (
		\key_i[101]_pad ,
		_w931_,
		_w2854_,
		_w2855_
	);
	LUT4 #(
		.INIT('h3222)
	) name1927 (
		\data_o[101]_pad ,
		_w931_,
		_w934_,
		_w2784_,
		_w2856_
	);
	LUT4 #(
		.INIT('h7b00)
	) name1928 (
		\ks1_key_reg_reg[101]/NET0131 ,
		_w2785_,
		_w2854_,
		_w2856_,
		_w2857_
	);
	LUT2 #(
		.INIT('he)
	) name1929 (
		_w2855_,
		_w2857_,
		_w2858_
	);
	LUT4 #(
		.INIT('haab8)
	) name1930 (
		\data_i[65]_pad ,
		decrypt_i_pad,
		\mix1_data_o_reg_reg[65]/NET0131 ,
		_w930_,
		_w2859_
	);
	LUT4 #(
		.INIT('haba8)
	) name1931 (
		\sub1_data_reg_reg[65]/NET0131 ,
		_w996_,
		_w2776_,
		_w2859_,
		_w2860_
	);
	LUT4 #(
		.INIT('h404c)
	) name1932 (
		\mix1_data_o_reg_reg[65]/NET0131 ,
		_w2774_,
		_w2775_,
		_w2860_,
		_w2861_
	);
	LUT4 #(
		.INIT('h0545)
	) name1933 (
		\sub1_data_reg_reg[65]/NET0131 ,
		\sub1_ready_o_reg/NET0131 ,
		_w1054_,
		_w2230_,
		_w2862_
	);
	LUT4 #(
		.INIT('h1015)
	) name1934 (
		\state_reg/NET0131 ,
		\sub1_data_reg_reg[65]/NET0131 ,
		_w996_,
		_w2859_,
		_w2863_
	);
	LUT4 #(
		.INIT('h0057)
	) name1935 (
		\state_reg/NET0131 ,
		_w2861_,
		_w2862_,
		_w2863_,
		_w2864_
	);
	LUT3 #(
		.INIT('h48)
	) name1936 (
		\key_i[65]_pad ,
		_w931_,
		_w2864_,
		_w2865_
	);
	LUT4 #(
		.INIT('h3222)
	) name1937 (
		\data_o[65]_pad ,
		_w931_,
		_w934_,
		_w2784_,
		_w2866_
	);
	LUT4 #(
		.INIT('h7b00)
	) name1938 (
		\ks1_key_reg_reg[65]/NET0131 ,
		_w2785_,
		_w2864_,
		_w2866_,
		_w2867_
	);
	LUT2 #(
		.INIT('he)
	) name1939 (
		_w2865_,
		_w2867_,
		_w2868_
	);
	LUT4 #(
		.INIT('haab8)
	) name1940 (
		\data_i[66]_pad ,
		decrypt_i_pad,
		\mix1_data_o_reg_reg[66]/NET0131 ,
		_w930_,
		_w2869_
	);
	LUT4 #(
		.INIT('haba8)
	) name1941 (
		\sub1_data_reg_reg[66]/NET0131 ,
		_w996_,
		_w2776_,
		_w2869_,
		_w2870_
	);
	LUT4 #(
		.INIT('h404c)
	) name1942 (
		\mix1_data_o_reg_reg[66]/NET0131 ,
		_w2774_,
		_w2775_,
		_w2870_,
		_w2871_
	);
	LUT4 #(
		.INIT('h0545)
	) name1943 (
		\sub1_data_reg_reg[66]/NET0131 ,
		\sub1_ready_o_reg/NET0131 ,
		_w1054_,
		_w2230_,
		_w2872_
	);
	LUT4 #(
		.INIT('h1015)
	) name1944 (
		\state_reg/NET0131 ,
		\sub1_data_reg_reg[66]/NET0131 ,
		_w996_,
		_w2869_,
		_w2873_
	);
	LUT4 #(
		.INIT('h0057)
	) name1945 (
		\state_reg/NET0131 ,
		_w2871_,
		_w2872_,
		_w2873_,
		_w2874_
	);
	LUT3 #(
		.INIT('h48)
	) name1946 (
		\key_i[66]_pad ,
		_w931_,
		_w2874_,
		_w2875_
	);
	LUT4 #(
		.INIT('h3222)
	) name1947 (
		\data_o[66]_pad ,
		_w931_,
		_w934_,
		_w2784_,
		_w2876_
	);
	LUT4 #(
		.INIT('h7b00)
	) name1948 (
		\ks1_key_reg_reg[66]/NET0131 ,
		_w2785_,
		_w2874_,
		_w2876_,
		_w2877_
	);
	LUT2 #(
		.INIT('he)
	) name1949 (
		_w2875_,
		_w2877_,
		_w2878_
	);
	LUT4 #(
		.INIT('haab8)
	) name1950 (
		\data_i[20]_pad ,
		decrypt_i_pad,
		\mix1_data_o_reg_reg[20]/NET0131 ,
		_w930_,
		_w2879_
	);
	LUT4 #(
		.INIT('haba8)
	) name1951 (
		\sub1_data_reg_reg[20]/NET0131 ,
		_w996_,
		_w2776_,
		_w2879_,
		_w2880_
	);
	LUT4 #(
		.INIT('h404c)
	) name1952 (
		\mix1_data_o_reg_reg[20]/NET0131 ,
		_w2774_,
		_w2775_,
		_w2880_,
		_w2881_
	);
	LUT4 #(
		.INIT('h0545)
	) name1953 (
		\sub1_data_reg_reg[20]/NET0131 ,
		\sub1_ready_o_reg/NET0131 ,
		_w1054_,
		_w2230_,
		_w2882_
	);
	LUT4 #(
		.INIT('h1015)
	) name1954 (
		\state_reg/NET0131 ,
		\sub1_data_reg_reg[20]/NET0131 ,
		_w996_,
		_w2879_,
		_w2883_
	);
	LUT4 #(
		.INIT('h0057)
	) name1955 (
		\state_reg/NET0131 ,
		_w2881_,
		_w2882_,
		_w2883_,
		_w2884_
	);
	LUT3 #(
		.INIT('h48)
	) name1956 (
		\key_i[20]_pad ,
		_w931_,
		_w2884_,
		_w2885_
	);
	LUT4 #(
		.INIT('h3222)
	) name1957 (
		\data_o[20]_pad ,
		_w931_,
		_w934_,
		_w2784_,
		_w2886_
	);
	LUT4 #(
		.INIT('h7b00)
	) name1958 (
		\ks1_key_reg_reg[20]/NET0131 ,
		_w2785_,
		_w2884_,
		_w2886_,
		_w2887_
	);
	LUT2 #(
		.INIT('he)
	) name1959 (
		_w2885_,
		_w2887_,
		_w2888_
	);
	LUT4 #(
		.INIT('haab8)
	) name1960 (
		\data_i[67]_pad ,
		decrypt_i_pad,
		\mix1_data_o_reg_reg[67]/NET0131 ,
		_w930_,
		_w2889_
	);
	LUT4 #(
		.INIT('haba8)
	) name1961 (
		\sub1_data_reg_reg[67]/NET0131 ,
		_w996_,
		_w2776_,
		_w2889_,
		_w2890_
	);
	LUT4 #(
		.INIT('h404c)
	) name1962 (
		\mix1_data_o_reg_reg[67]/NET0131 ,
		_w2774_,
		_w2775_,
		_w2890_,
		_w2891_
	);
	LUT4 #(
		.INIT('h0545)
	) name1963 (
		\sub1_data_reg_reg[67]/NET0131 ,
		\sub1_ready_o_reg/NET0131 ,
		_w1054_,
		_w2230_,
		_w2892_
	);
	LUT4 #(
		.INIT('h1015)
	) name1964 (
		\state_reg/NET0131 ,
		\sub1_data_reg_reg[67]/NET0131 ,
		_w996_,
		_w2889_,
		_w2893_
	);
	LUT4 #(
		.INIT('h0057)
	) name1965 (
		\state_reg/NET0131 ,
		_w2891_,
		_w2892_,
		_w2893_,
		_w2894_
	);
	LUT3 #(
		.INIT('h48)
	) name1966 (
		\key_i[67]_pad ,
		_w931_,
		_w2894_,
		_w2895_
	);
	LUT4 #(
		.INIT('h3222)
	) name1967 (
		\data_o[67]_pad ,
		_w931_,
		_w934_,
		_w2784_,
		_w2896_
	);
	LUT4 #(
		.INIT('h7b00)
	) name1968 (
		\ks1_key_reg_reg[67]/NET0131 ,
		_w2785_,
		_w2894_,
		_w2896_,
		_w2897_
	);
	LUT2 #(
		.INIT('he)
	) name1969 (
		_w2895_,
		_w2897_,
		_w2898_
	);
	LUT4 #(
		.INIT('haab8)
	) name1970 (
		\data_i[113]_pad ,
		decrypt_i_pad,
		\mix1_data_o_reg_reg[113]/NET0131 ,
		_w930_,
		_w2899_
	);
	LUT4 #(
		.INIT('haba8)
	) name1971 (
		\sub1_data_reg_reg[113]/NET0131 ,
		_w996_,
		_w2776_,
		_w2899_,
		_w2900_
	);
	LUT4 #(
		.INIT('h404c)
	) name1972 (
		\mix1_data_o_reg_reg[113]/NET0131 ,
		_w2774_,
		_w2775_,
		_w2900_,
		_w2901_
	);
	LUT4 #(
		.INIT('h0545)
	) name1973 (
		\sub1_data_reg_reg[113]/NET0131 ,
		\sub1_ready_o_reg/NET0131 ,
		_w1054_,
		_w2230_,
		_w2902_
	);
	LUT4 #(
		.INIT('h1015)
	) name1974 (
		\state_reg/NET0131 ,
		\sub1_data_reg_reg[113]/NET0131 ,
		_w996_,
		_w2899_,
		_w2903_
	);
	LUT4 #(
		.INIT('h0057)
	) name1975 (
		\state_reg/NET0131 ,
		_w2901_,
		_w2902_,
		_w2903_,
		_w2904_
	);
	LUT3 #(
		.INIT('h48)
	) name1976 (
		\key_i[113]_pad ,
		_w931_,
		_w2904_,
		_w2905_
	);
	LUT4 #(
		.INIT('h3222)
	) name1977 (
		\data_o[113]_pad ,
		_w931_,
		_w934_,
		_w2784_,
		_w2906_
	);
	LUT4 #(
		.INIT('h7b00)
	) name1978 (
		\ks1_key_reg_reg[113]/NET0131 ,
		_w2785_,
		_w2904_,
		_w2906_,
		_w2907_
	);
	LUT2 #(
		.INIT('he)
	) name1979 (
		_w2905_,
		_w2907_,
		_w2908_
	);
	LUT4 #(
		.INIT('haab8)
	) name1980 (
		\data_i[21]_pad ,
		decrypt_i_pad,
		\mix1_data_o_reg_reg[21]/NET0131 ,
		_w930_,
		_w2909_
	);
	LUT4 #(
		.INIT('haba8)
	) name1981 (
		\sub1_data_reg_reg[21]/NET0131 ,
		_w996_,
		_w2776_,
		_w2909_,
		_w2910_
	);
	LUT4 #(
		.INIT('h404c)
	) name1982 (
		\mix1_data_o_reg_reg[21]/NET0131 ,
		_w2774_,
		_w2775_,
		_w2910_,
		_w2911_
	);
	LUT4 #(
		.INIT('h0545)
	) name1983 (
		\sub1_data_reg_reg[21]/NET0131 ,
		\sub1_ready_o_reg/NET0131 ,
		_w1054_,
		_w2230_,
		_w2912_
	);
	LUT4 #(
		.INIT('h1015)
	) name1984 (
		\state_reg/NET0131 ,
		\sub1_data_reg_reg[21]/NET0131 ,
		_w996_,
		_w2909_,
		_w2913_
	);
	LUT4 #(
		.INIT('h0057)
	) name1985 (
		\state_reg/NET0131 ,
		_w2911_,
		_w2912_,
		_w2913_,
		_w2914_
	);
	LUT3 #(
		.INIT('h48)
	) name1986 (
		\key_i[21]_pad ,
		_w931_,
		_w2914_,
		_w2915_
	);
	LUT4 #(
		.INIT('h3222)
	) name1987 (
		\data_o[21]_pad ,
		_w931_,
		_w934_,
		_w2784_,
		_w2916_
	);
	LUT4 #(
		.INIT('h7b00)
	) name1988 (
		\ks1_key_reg_reg[21]/NET0131 ,
		_w2785_,
		_w2914_,
		_w2916_,
		_w2917_
	);
	LUT2 #(
		.INIT('he)
	) name1989 (
		_w2915_,
		_w2917_,
		_w2918_
	);
	LUT4 #(
		.INIT('haab8)
	) name1990 (
		\data_i[68]_pad ,
		decrypt_i_pad,
		\mix1_data_o_reg_reg[68]/NET0131 ,
		_w930_,
		_w2919_
	);
	LUT4 #(
		.INIT('haba8)
	) name1991 (
		\sub1_data_reg_reg[68]/NET0131 ,
		_w996_,
		_w2776_,
		_w2919_,
		_w2920_
	);
	LUT4 #(
		.INIT('h404c)
	) name1992 (
		\mix1_data_o_reg_reg[68]/NET0131 ,
		_w2774_,
		_w2775_,
		_w2920_,
		_w2921_
	);
	LUT4 #(
		.INIT('h0545)
	) name1993 (
		\sub1_data_reg_reg[68]/NET0131 ,
		\sub1_ready_o_reg/NET0131 ,
		_w1054_,
		_w2230_,
		_w2922_
	);
	LUT4 #(
		.INIT('h1015)
	) name1994 (
		\state_reg/NET0131 ,
		\sub1_data_reg_reg[68]/NET0131 ,
		_w996_,
		_w2919_,
		_w2923_
	);
	LUT4 #(
		.INIT('h0057)
	) name1995 (
		\state_reg/NET0131 ,
		_w2921_,
		_w2922_,
		_w2923_,
		_w2924_
	);
	LUT3 #(
		.INIT('h48)
	) name1996 (
		\key_i[68]_pad ,
		_w931_,
		_w2924_,
		_w2925_
	);
	LUT4 #(
		.INIT('h3222)
	) name1997 (
		\data_o[68]_pad ,
		_w931_,
		_w934_,
		_w2784_,
		_w2926_
	);
	LUT4 #(
		.INIT('h7b00)
	) name1998 (
		\ks1_key_reg_reg[68]/NET0131 ,
		_w2785_,
		_w2924_,
		_w2926_,
		_w2927_
	);
	LUT2 #(
		.INIT('he)
	) name1999 (
		_w2925_,
		_w2927_,
		_w2928_
	);
	LUT4 #(
		.INIT('haab8)
	) name2000 (
		\data_i[69]_pad ,
		decrypt_i_pad,
		\mix1_data_o_reg_reg[69]/NET0131 ,
		_w930_,
		_w2929_
	);
	LUT4 #(
		.INIT('haba8)
	) name2001 (
		\sub1_data_reg_reg[69]/NET0131 ,
		_w996_,
		_w2776_,
		_w2929_,
		_w2930_
	);
	LUT4 #(
		.INIT('h404c)
	) name2002 (
		\mix1_data_o_reg_reg[69]/NET0131 ,
		_w2774_,
		_w2775_,
		_w2930_,
		_w2931_
	);
	LUT4 #(
		.INIT('h0545)
	) name2003 (
		\sub1_data_reg_reg[69]/NET0131 ,
		\sub1_ready_o_reg/NET0131 ,
		_w1054_,
		_w2230_,
		_w2932_
	);
	LUT4 #(
		.INIT('h1015)
	) name2004 (
		\state_reg/NET0131 ,
		\sub1_data_reg_reg[69]/NET0131 ,
		_w996_,
		_w2929_,
		_w2933_
	);
	LUT4 #(
		.INIT('h0057)
	) name2005 (
		\state_reg/NET0131 ,
		_w2931_,
		_w2932_,
		_w2933_,
		_w2934_
	);
	LUT3 #(
		.INIT('h48)
	) name2006 (
		\key_i[69]_pad ,
		_w931_,
		_w2934_,
		_w2935_
	);
	LUT4 #(
		.INIT('h3222)
	) name2007 (
		\data_o[69]_pad ,
		_w931_,
		_w934_,
		_w2784_,
		_w2936_
	);
	LUT4 #(
		.INIT('h7b00)
	) name2008 (
		\ks1_key_reg_reg[69]/NET0131 ,
		_w2785_,
		_w2934_,
		_w2936_,
		_w2937_
	);
	LUT2 #(
		.INIT('he)
	) name2009 (
		_w2935_,
		_w2937_,
		_w2938_
	);
	LUT4 #(
		.INIT('haab8)
	) name2010 (
		\data_i[102]_pad ,
		decrypt_i_pad,
		\mix1_data_o_reg_reg[102]/NET0131 ,
		_w930_,
		_w2939_
	);
	LUT4 #(
		.INIT('haba8)
	) name2011 (
		\sub1_data_reg_reg[102]/NET0131 ,
		_w996_,
		_w2776_,
		_w2939_,
		_w2940_
	);
	LUT4 #(
		.INIT('h404c)
	) name2012 (
		\mix1_data_o_reg_reg[102]/NET0131 ,
		_w2774_,
		_w2775_,
		_w2940_,
		_w2941_
	);
	LUT4 #(
		.INIT('h0545)
	) name2013 (
		\sub1_data_reg_reg[102]/NET0131 ,
		\sub1_ready_o_reg/NET0131 ,
		_w1054_,
		_w2230_,
		_w2942_
	);
	LUT4 #(
		.INIT('h1015)
	) name2014 (
		\state_reg/NET0131 ,
		\sub1_data_reg_reg[102]/NET0131 ,
		_w996_,
		_w2939_,
		_w2943_
	);
	LUT4 #(
		.INIT('h0057)
	) name2015 (
		\state_reg/NET0131 ,
		_w2941_,
		_w2942_,
		_w2943_,
		_w2944_
	);
	LUT3 #(
		.INIT('h48)
	) name2016 (
		\key_i[102]_pad ,
		_w931_,
		_w2944_,
		_w2945_
	);
	LUT4 #(
		.INIT('h3222)
	) name2017 (
		\data_o[102]_pad ,
		_w931_,
		_w934_,
		_w2784_,
		_w2946_
	);
	LUT4 #(
		.INIT('h7b00)
	) name2018 (
		\ks1_key_reg_reg[102]/NET0131 ,
		_w2785_,
		_w2944_,
		_w2946_,
		_w2947_
	);
	LUT2 #(
		.INIT('he)
	) name2019 (
		_w2945_,
		_w2947_,
		_w2948_
	);
	LUT4 #(
		.INIT('haab8)
	) name2020 (
		\data_i[114]_pad ,
		decrypt_i_pad,
		\mix1_data_o_reg_reg[114]/NET0131 ,
		_w930_,
		_w2949_
	);
	LUT4 #(
		.INIT('haba8)
	) name2021 (
		\sub1_data_reg_reg[114]/NET0131 ,
		_w996_,
		_w2776_,
		_w2949_,
		_w2950_
	);
	LUT4 #(
		.INIT('h404c)
	) name2022 (
		\mix1_data_o_reg_reg[114]/NET0131 ,
		_w2774_,
		_w2775_,
		_w2950_,
		_w2951_
	);
	LUT4 #(
		.INIT('h0545)
	) name2023 (
		\sub1_data_reg_reg[114]/NET0131 ,
		\sub1_ready_o_reg/NET0131 ,
		_w1054_,
		_w2230_,
		_w2952_
	);
	LUT4 #(
		.INIT('h1015)
	) name2024 (
		\state_reg/NET0131 ,
		\sub1_data_reg_reg[114]/NET0131 ,
		_w996_,
		_w2949_,
		_w2953_
	);
	LUT4 #(
		.INIT('h0057)
	) name2025 (
		\state_reg/NET0131 ,
		_w2951_,
		_w2952_,
		_w2953_,
		_w2954_
	);
	LUT3 #(
		.INIT('h48)
	) name2026 (
		\key_i[114]_pad ,
		_w931_,
		_w2954_,
		_w2955_
	);
	LUT4 #(
		.INIT('h3222)
	) name2027 (
		\data_o[114]_pad ,
		_w931_,
		_w934_,
		_w2784_,
		_w2956_
	);
	LUT4 #(
		.INIT('h7b00)
	) name2028 (
		\ks1_key_reg_reg[114]/NET0131 ,
		_w2785_,
		_w2954_,
		_w2956_,
		_w2957_
	);
	LUT2 #(
		.INIT('he)
	) name2029 (
		_w2955_,
		_w2957_,
		_w2958_
	);
	LUT4 #(
		.INIT('h5547)
	) name2030 (
		\data_i[6]_pad ,
		decrypt_i_pad,
		\mix1_data_o_reg_reg[6]/NET0131 ,
		_w930_,
		_w2959_
	);
	LUT4 #(
		.INIT('ha8ab)
	) name2031 (
		\sub1_data_reg_reg[6]/NET0131 ,
		_w996_,
		_w2776_,
		_w2959_,
		_w2960_
	);
	LUT4 #(
		.INIT('h404c)
	) name2032 (
		\mix1_data_o_reg_reg[6]/NET0131 ,
		_w2774_,
		_w2775_,
		_w2960_,
		_w2961_
	);
	LUT4 #(
		.INIT('h0545)
	) name2033 (
		\sub1_data_reg_reg[6]/NET0131 ,
		\sub1_ready_o_reg/NET0131 ,
		_w1054_,
		_w2230_,
		_w2962_
	);
	LUT4 #(
		.INIT('h1510)
	) name2034 (
		\state_reg/NET0131 ,
		\sub1_data_reg_reg[6]/NET0131 ,
		_w996_,
		_w2959_,
		_w2963_
	);
	LUT4 #(
		.INIT('h0057)
	) name2035 (
		\state_reg/NET0131 ,
		_w2961_,
		_w2962_,
		_w2963_,
		_w2964_
	);
	LUT3 #(
		.INIT('h48)
	) name2036 (
		\key_i[6]_pad ,
		_w931_,
		_w2964_,
		_w2965_
	);
	LUT4 #(
		.INIT('h3222)
	) name2037 (
		\data_o[6]_pad ,
		_w931_,
		_w934_,
		_w2784_,
		_w2966_
	);
	LUT4 #(
		.INIT('h7b00)
	) name2038 (
		\ks1_key_reg_reg[6]/NET0131 ,
		_w2785_,
		_w2964_,
		_w2966_,
		_w2967_
	);
	LUT2 #(
		.INIT('he)
	) name2039 (
		_w2965_,
		_w2967_,
		_w2968_
	);
	LUT4 #(
		.INIT('haab8)
	) name2040 (
		\data_i[22]_pad ,
		decrypt_i_pad,
		\mix1_data_o_reg_reg[22]/NET0131 ,
		_w930_,
		_w2969_
	);
	LUT4 #(
		.INIT('haba8)
	) name2041 (
		\sub1_data_reg_reg[22]/NET0131 ,
		_w996_,
		_w2776_,
		_w2969_,
		_w2970_
	);
	LUT4 #(
		.INIT('h404c)
	) name2042 (
		\mix1_data_o_reg_reg[22]/NET0131 ,
		_w2774_,
		_w2775_,
		_w2970_,
		_w2971_
	);
	LUT4 #(
		.INIT('h0545)
	) name2043 (
		\sub1_data_reg_reg[22]/NET0131 ,
		\sub1_ready_o_reg/NET0131 ,
		_w1054_,
		_w2230_,
		_w2972_
	);
	LUT4 #(
		.INIT('h1015)
	) name2044 (
		\state_reg/NET0131 ,
		\sub1_data_reg_reg[22]/NET0131 ,
		_w996_,
		_w2969_,
		_w2973_
	);
	LUT4 #(
		.INIT('h0057)
	) name2045 (
		\state_reg/NET0131 ,
		_w2971_,
		_w2972_,
		_w2973_,
		_w2974_
	);
	LUT3 #(
		.INIT('h48)
	) name2046 (
		\key_i[22]_pad ,
		_w931_,
		_w2974_,
		_w2975_
	);
	LUT4 #(
		.INIT('h3222)
	) name2047 (
		\data_o[22]_pad ,
		_w931_,
		_w934_,
		_w2784_,
		_w2976_
	);
	LUT4 #(
		.INIT('h7b00)
	) name2048 (
		\ks1_key_reg_reg[22]/NET0131 ,
		_w2785_,
		_w2974_,
		_w2976_,
		_w2977_
	);
	LUT2 #(
		.INIT('he)
	) name2049 (
		_w2975_,
		_w2977_,
		_w2978_
	);
	LUT4 #(
		.INIT('haab8)
	) name2050 (
		\data_i[70]_pad ,
		decrypt_i_pad,
		\mix1_data_o_reg_reg[70]/NET0131 ,
		_w930_,
		_w2979_
	);
	LUT4 #(
		.INIT('haba8)
	) name2051 (
		\sub1_data_reg_reg[70]/NET0131 ,
		_w996_,
		_w2776_,
		_w2979_,
		_w2980_
	);
	LUT4 #(
		.INIT('h404c)
	) name2052 (
		\mix1_data_o_reg_reg[70]/NET0131 ,
		_w2774_,
		_w2775_,
		_w2980_,
		_w2981_
	);
	LUT4 #(
		.INIT('h0545)
	) name2053 (
		\sub1_data_reg_reg[70]/NET0131 ,
		\sub1_ready_o_reg/NET0131 ,
		_w1054_,
		_w2230_,
		_w2982_
	);
	LUT4 #(
		.INIT('h1015)
	) name2054 (
		\state_reg/NET0131 ,
		\sub1_data_reg_reg[70]/NET0131 ,
		_w996_,
		_w2979_,
		_w2983_
	);
	LUT4 #(
		.INIT('h0057)
	) name2055 (
		\state_reg/NET0131 ,
		_w2981_,
		_w2982_,
		_w2983_,
		_w2984_
	);
	LUT3 #(
		.INIT('h48)
	) name2056 (
		\key_i[70]_pad ,
		_w931_,
		_w2984_,
		_w2985_
	);
	LUT4 #(
		.INIT('h3222)
	) name2057 (
		\data_o[70]_pad ,
		_w931_,
		_w934_,
		_w2784_,
		_w2986_
	);
	LUT4 #(
		.INIT('h7b00)
	) name2058 (
		\ks1_key_reg_reg[70]/NET0131 ,
		_w2785_,
		_w2984_,
		_w2986_,
		_w2987_
	);
	LUT2 #(
		.INIT('he)
	) name2059 (
		_w2985_,
		_w2987_,
		_w2988_
	);
	LUT4 #(
		.INIT('haab8)
	) name2060 (
		\data_i[71]_pad ,
		decrypt_i_pad,
		\mix1_data_o_reg_reg[71]/NET0131 ,
		_w930_,
		_w2989_
	);
	LUT4 #(
		.INIT('haba8)
	) name2061 (
		\sub1_data_reg_reg[71]/NET0131 ,
		_w996_,
		_w2776_,
		_w2989_,
		_w2990_
	);
	LUT4 #(
		.INIT('h404c)
	) name2062 (
		\mix1_data_o_reg_reg[71]/NET0131 ,
		_w2774_,
		_w2775_,
		_w2990_,
		_w2991_
	);
	LUT4 #(
		.INIT('h0545)
	) name2063 (
		\sub1_data_reg_reg[71]/NET0131 ,
		\sub1_ready_o_reg/NET0131 ,
		_w1054_,
		_w2230_,
		_w2992_
	);
	LUT4 #(
		.INIT('h1015)
	) name2064 (
		\state_reg/NET0131 ,
		\sub1_data_reg_reg[71]/NET0131 ,
		_w996_,
		_w2989_,
		_w2993_
	);
	LUT4 #(
		.INIT('h0057)
	) name2065 (
		\state_reg/NET0131 ,
		_w2991_,
		_w2992_,
		_w2993_,
		_w2994_
	);
	LUT3 #(
		.INIT('h48)
	) name2066 (
		\key_i[71]_pad ,
		_w931_,
		_w2994_,
		_w2995_
	);
	LUT4 #(
		.INIT('h3222)
	) name2067 (
		\data_o[71]_pad ,
		_w931_,
		_w934_,
		_w2784_,
		_w2996_
	);
	LUT4 #(
		.INIT('h7b00)
	) name2068 (
		\ks1_key_reg_reg[71]/NET0131 ,
		_w2785_,
		_w2994_,
		_w2996_,
		_w2997_
	);
	LUT2 #(
		.INIT('he)
	) name2069 (
		_w2995_,
		_w2997_,
		_w2998_
	);
	LUT4 #(
		.INIT('haab8)
	) name2070 (
		\data_i[23]_pad ,
		decrypt_i_pad,
		\mix1_data_o_reg_reg[23]/NET0131 ,
		_w930_,
		_w2999_
	);
	LUT4 #(
		.INIT('haba8)
	) name2071 (
		\sub1_data_reg_reg[23]/NET0131 ,
		_w996_,
		_w2776_,
		_w2999_,
		_w3000_
	);
	LUT4 #(
		.INIT('h404c)
	) name2072 (
		\mix1_data_o_reg_reg[23]/NET0131 ,
		_w2774_,
		_w2775_,
		_w3000_,
		_w3001_
	);
	LUT4 #(
		.INIT('h0545)
	) name2073 (
		\sub1_data_reg_reg[23]/NET0131 ,
		\sub1_ready_o_reg/NET0131 ,
		_w1054_,
		_w2230_,
		_w3002_
	);
	LUT4 #(
		.INIT('h1015)
	) name2074 (
		\state_reg/NET0131 ,
		\sub1_data_reg_reg[23]/NET0131 ,
		_w996_,
		_w2999_,
		_w3003_
	);
	LUT4 #(
		.INIT('h0057)
	) name2075 (
		\state_reg/NET0131 ,
		_w3001_,
		_w3002_,
		_w3003_,
		_w3004_
	);
	LUT3 #(
		.INIT('h48)
	) name2076 (
		\key_i[23]_pad ,
		_w931_,
		_w3004_,
		_w3005_
	);
	LUT4 #(
		.INIT('h3222)
	) name2077 (
		\data_o[23]_pad ,
		_w931_,
		_w934_,
		_w2784_,
		_w3006_
	);
	LUT4 #(
		.INIT('h7b00)
	) name2078 (
		\ks1_key_reg_reg[23]/NET0131 ,
		_w2785_,
		_w3004_,
		_w3006_,
		_w3007_
	);
	LUT2 #(
		.INIT('he)
	) name2079 (
		_w3005_,
		_w3007_,
		_w3008_
	);
	LUT4 #(
		.INIT('haab8)
	) name2080 (
		\data_i[115]_pad ,
		decrypt_i_pad,
		\mix1_data_o_reg_reg[115]/NET0131 ,
		_w930_,
		_w3009_
	);
	LUT4 #(
		.INIT('haba8)
	) name2081 (
		\sub1_data_reg_reg[115]/NET0131 ,
		_w996_,
		_w2776_,
		_w3009_,
		_w3010_
	);
	LUT4 #(
		.INIT('h404c)
	) name2082 (
		\mix1_data_o_reg_reg[115]/NET0131 ,
		_w2774_,
		_w2775_,
		_w3010_,
		_w3011_
	);
	LUT4 #(
		.INIT('h0545)
	) name2083 (
		\sub1_data_reg_reg[115]/NET0131 ,
		\sub1_ready_o_reg/NET0131 ,
		_w1054_,
		_w2230_,
		_w3012_
	);
	LUT4 #(
		.INIT('h1015)
	) name2084 (
		\state_reg/NET0131 ,
		\sub1_data_reg_reg[115]/NET0131 ,
		_w996_,
		_w3009_,
		_w3013_
	);
	LUT4 #(
		.INIT('h0057)
	) name2085 (
		\state_reg/NET0131 ,
		_w3011_,
		_w3012_,
		_w3013_,
		_w3014_
	);
	LUT3 #(
		.INIT('h48)
	) name2086 (
		\key_i[115]_pad ,
		_w931_,
		_w3014_,
		_w3015_
	);
	LUT4 #(
		.INIT('h3222)
	) name2087 (
		\data_o[115]_pad ,
		_w931_,
		_w934_,
		_w2784_,
		_w3016_
	);
	LUT4 #(
		.INIT('h7b00)
	) name2088 (
		\ks1_key_reg_reg[115]/NET0131 ,
		_w2785_,
		_w3014_,
		_w3016_,
		_w3017_
	);
	LUT2 #(
		.INIT('he)
	) name2089 (
		_w3015_,
		_w3017_,
		_w3018_
	);
	LUT4 #(
		.INIT('h5547)
	) name2090 (
		\data_i[72]_pad ,
		decrypt_i_pad,
		\mix1_data_o_reg_reg[72]/NET0131 ,
		_w930_,
		_w3019_
	);
	LUT4 #(
		.INIT('ha8ab)
	) name2091 (
		\sub1_data_reg_reg[72]/NET0131 ,
		_w996_,
		_w2776_,
		_w3019_,
		_w3020_
	);
	LUT4 #(
		.INIT('h404c)
	) name2092 (
		\mix1_data_o_reg_reg[72]/NET0131 ,
		_w2774_,
		_w2775_,
		_w3020_,
		_w3021_
	);
	LUT4 #(
		.INIT('h0545)
	) name2093 (
		\sub1_data_reg_reg[72]/NET0131 ,
		\sub1_ready_o_reg/NET0131 ,
		_w1054_,
		_w2230_,
		_w3022_
	);
	LUT4 #(
		.INIT('h1510)
	) name2094 (
		\state_reg/NET0131 ,
		\sub1_data_reg_reg[72]/NET0131 ,
		_w996_,
		_w3019_,
		_w3023_
	);
	LUT4 #(
		.INIT('h0057)
	) name2095 (
		\state_reg/NET0131 ,
		_w3021_,
		_w3022_,
		_w3023_,
		_w3024_
	);
	LUT3 #(
		.INIT('h48)
	) name2096 (
		\key_i[72]_pad ,
		_w931_,
		_w3024_,
		_w3025_
	);
	LUT4 #(
		.INIT('h3222)
	) name2097 (
		\data_o[72]_pad ,
		_w931_,
		_w934_,
		_w2784_,
		_w3026_
	);
	LUT4 #(
		.INIT('h7b00)
	) name2098 (
		\ks1_key_reg_reg[72]/P0002 ,
		_w2785_,
		_w3024_,
		_w3026_,
		_w3027_
	);
	LUT2 #(
		.INIT('he)
	) name2099 (
		_w3025_,
		_w3027_,
		_w3028_
	);
	LUT4 #(
		.INIT('h5547)
	) name2100 (
		\data_i[24]_pad ,
		decrypt_i_pad,
		\mix1_data_o_reg_reg[24]/NET0131 ,
		_w930_,
		_w3029_
	);
	LUT4 #(
		.INIT('ha8ab)
	) name2101 (
		\sub1_data_reg_reg[24]/NET0131 ,
		_w996_,
		_w2776_,
		_w3029_,
		_w3030_
	);
	LUT4 #(
		.INIT('h404c)
	) name2102 (
		\mix1_data_o_reg_reg[24]/NET0131 ,
		_w2774_,
		_w2775_,
		_w3030_,
		_w3031_
	);
	LUT4 #(
		.INIT('h0545)
	) name2103 (
		\sub1_data_reg_reg[24]/NET0131 ,
		\sub1_ready_o_reg/NET0131 ,
		_w1054_,
		_w2230_,
		_w3032_
	);
	LUT4 #(
		.INIT('h1510)
	) name2104 (
		\state_reg/NET0131 ,
		\sub1_data_reg_reg[24]/NET0131 ,
		_w996_,
		_w3029_,
		_w3033_
	);
	LUT4 #(
		.INIT('h0057)
	) name2105 (
		\state_reg/NET0131 ,
		_w3031_,
		_w3032_,
		_w3033_,
		_w3034_
	);
	LUT3 #(
		.INIT('h48)
	) name2106 (
		\key_i[24]_pad ,
		_w931_,
		_w3034_,
		_w3035_
	);
	LUT4 #(
		.INIT('h3222)
	) name2107 (
		\data_o[24]_pad ,
		_w931_,
		_w934_,
		_w2784_,
		_w3036_
	);
	LUT4 #(
		.INIT('h7b00)
	) name2108 (
		\ks1_key_reg_reg[24]/NET0131 ,
		_w2785_,
		_w3034_,
		_w3036_,
		_w3037_
	);
	LUT2 #(
		.INIT('he)
	) name2109 (
		_w3035_,
		_w3037_,
		_w3038_
	);
	LUT4 #(
		.INIT('h5547)
	) name2110 (
		\data_i[73]_pad ,
		decrypt_i_pad,
		\mix1_data_o_reg_reg[73]/NET0131 ,
		_w930_,
		_w3039_
	);
	LUT4 #(
		.INIT('ha8ab)
	) name2111 (
		\sub1_data_reg_reg[73]/NET0131 ,
		_w996_,
		_w2776_,
		_w3039_,
		_w3040_
	);
	LUT4 #(
		.INIT('h404c)
	) name2112 (
		\mix1_data_o_reg_reg[73]/NET0131 ,
		_w2774_,
		_w2775_,
		_w3040_,
		_w3041_
	);
	LUT4 #(
		.INIT('h0545)
	) name2113 (
		\sub1_data_reg_reg[73]/NET0131 ,
		\sub1_ready_o_reg/NET0131 ,
		_w1054_,
		_w2230_,
		_w3042_
	);
	LUT4 #(
		.INIT('h1510)
	) name2114 (
		\state_reg/NET0131 ,
		\sub1_data_reg_reg[73]/NET0131 ,
		_w996_,
		_w3039_,
		_w3043_
	);
	LUT4 #(
		.INIT('h0057)
	) name2115 (
		\state_reg/NET0131 ,
		_w3041_,
		_w3042_,
		_w3043_,
		_w3044_
	);
	LUT3 #(
		.INIT('h48)
	) name2116 (
		\key_i[73]_pad ,
		_w931_,
		_w3044_,
		_w3045_
	);
	LUT4 #(
		.INIT('h3222)
	) name2117 (
		\data_o[73]_pad ,
		_w931_,
		_w934_,
		_w2784_,
		_w3046_
	);
	LUT4 #(
		.INIT('h7b00)
	) name2118 (
		\ks1_key_reg_reg[73]/NET0131 ,
		_w2785_,
		_w3044_,
		_w3046_,
		_w3047_
	);
	LUT2 #(
		.INIT('he)
	) name2119 (
		_w3045_,
		_w3047_,
		_w3048_
	);
	LUT4 #(
		.INIT('h5547)
	) name2120 (
		\data_i[74]_pad ,
		decrypt_i_pad,
		\mix1_data_o_reg_reg[74]/NET0131 ,
		_w930_,
		_w3049_
	);
	LUT4 #(
		.INIT('ha8ab)
	) name2121 (
		\sub1_data_reg_reg[74]/NET0131 ,
		_w996_,
		_w2776_,
		_w3049_,
		_w3050_
	);
	LUT4 #(
		.INIT('h404c)
	) name2122 (
		\mix1_data_o_reg_reg[74]/NET0131 ,
		_w2774_,
		_w2775_,
		_w3050_,
		_w3051_
	);
	LUT4 #(
		.INIT('h0545)
	) name2123 (
		\sub1_data_reg_reg[74]/NET0131 ,
		\sub1_ready_o_reg/NET0131 ,
		_w1054_,
		_w2230_,
		_w3052_
	);
	LUT4 #(
		.INIT('h1510)
	) name2124 (
		\state_reg/NET0131 ,
		\sub1_data_reg_reg[74]/NET0131 ,
		_w996_,
		_w3049_,
		_w3053_
	);
	LUT4 #(
		.INIT('h0057)
	) name2125 (
		\state_reg/NET0131 ,
		_w3051_,
		_w3052_,
		_w3053_,
		_w3054_
	);
	LUT3 #(
		.INIT('h48)
	) name2126 (
		\key_i[74]_pad ,
		_w931_,
		_w3054_,
		_w3055_
	);
	LUT4 #(
		.INIT('h3222)
	) name2127 (
		\data_o[74]_pad ,
		_w931_,
		_w934_,
		_w2784_,
		_w3056_
	);
	LUT4 #(
		.INIT('h7b00)
	) name2128 (
		\ks1_key_reg_reg[74]/NET0131 ,
		_w2785_,
		_w3054_,
		_w3056_,
		_w3057_
	);
	LUT2 #(
		.INIT('he)
	) name2129 (
		_w3055_,
		_w3057_,
		_w3058_
	);
	LUT4 #(
		.INIT('h5547)
	) name2130 (
		\data_i[25]_pad ,
		decrypt_i_pad,
		\mix1_data_o_reg_reg[25]/NET0131 ,
		_w930_,
		_w3059_
	);
	LUT4 #(
		.INIT('ha8ab)
	) name2131 (
		\sub1_data_reg_reg[25]/NET0131 ,
		_w996_,
		_w2776_,
		_w3059_,
		_w3060_
	);
	LUT4 #(
		.INIT('h404c)
	) name2132 (
		\mix1_data_o_reg_reg[25]/NET0131 ,
		_w2774_,
		_w2775_,
		_w3060_,
		_w3061_
	);
	LUT4 #(
		.INIT('h0545)
	) name2133 (
		\sub1_data_reg_reg[25]/NET0131 ,
		\sub1_ready_o_reg/NET0131 ,
		_w1054_,
		_w2230_,
		_w3062_
	);
	LUT4 #(
		.INIT('h1510)
	) name2134 (
		\state_reg/NET0131 ,
		\sub1_data_reg_reg[25]/NET0131 ,
		_w996_,
		_w3059_,
		_w3063_
	);
	LUT4 #(
		.INIT('h0057)
	) name2135 (
		\state_reg/NET0131 ,
		_w3061_,
		_w3062_,
		_w3063_,
		_w3064_
	);
	LUT3 #(
		.INIT('h48)
	) name2136 (
		\key_i[25]_pad ,
		_w931_,
		_w3064_,
		_w3065_
	);
	LUT4 #(
		.INIT('h3222)
	) name2137 (
		\data_o[25]_pad ,
		_w931_,
		_w934_,
		_w2784_,
		_w3066_
	);
	LUT4 #(
		.INIT('h7b00)
	) name2138 (
		\ks1_key_reg_reg[25]/NET0131 ,
		_w2785_,
		_w3064_,
		_w3066_,
		_w3067_
	);
	LUT2 #(
		.INIT('he)
	) name2139 (
		_w3065_,
		_w3067_,
		_w3068_
	);
	LUT4 #(
		.INIT('h5547)
	) name2140 (
		\data_i[75]_pad ,
		decrypt_i_pad,
		\mix1_data_o_reg_reg[75]/NET0131 ,
		_w930_,
		_w3069_
	);
	LUT4 #(
		.INIT('ha8ab)
	) name2141 (
		\sub1_data_reg_reg[75]/NET0131 ,
		_w996_,
		_w2776_,
		_w3069_,
		_w3070_
	);
	LUT4 #(
		.INIT('h404c)
	) name2142 (
		\mix1_data_o_reg_reg[75]/NET0131 ,
		_w2774_,
		_w2775_,
		_w3070_,
		_w3071_
	);
	LUT4 #(
		.INIT('h0545)
	) name2143 (
		\sub1_data_reg_reg[75]/NET0131 ,
		\sub1_ready_o_reg/NET0131 ,
		_w1054_,
		_w2230_,
		_w3072_
	);
	LUT4 #(
		.INIT('h1510)
	) name2144 (
		\state_reg/NET0131 ,
		\sub1_data_reg_reg[75]/NET0131 ,
		_w996_,
		_w3069_,
		_w3073_
	);
	LUT4 #(
		.INIT('h0057)
	) name2145 (
		\state_reg/NET0131 ,
		_w3071_,
		_w3072_,
		_w3073_,
		_w3074_
	);
	LUT3 #(
		.INIT('h48)
	) name2146 (
		\key_i[75]_pad ,
		_w931_,
		_w3074_,
		_w3075_
	);
	LUT4 #(
		.INIT('h3222)
	) name2147 (
		\data_o[75]_pad ,
		_w931_,
		_w934_,
		_w2784_,
		_w3076_
	);
	LUT4 #(
		.INIT('h7b00)
	) name2148 (
		\ks1_key_reg_reg[75]/P0002 ,
		_w2785_,
		_w3074_,
		_w3076_,
		_w3077_
	);
	LUT2 #(
		.INIT('he)
	) name2149 (
		_w3075_,
		_w3077_,
		_w3078_
	);
	LUT4 #(
		.INIT('h5547)
	) name2150 (
		\data_i[76]_pad ,
		decrypt_i_pad,
		\mix1_data_o_reg_reg[76]/NET0131 ,
		_w930_,
		_w3079_
	);
	LUT4 #(
		.INIT('ha8ab)
	) name2151 (
		\sub1_data_reg_reg[76]/NET0131 ,
		_w996_,
		_w2776_,
		_w3079_,
		_w3080_
	);
	LUT4 #(
		.INIT('h404c)
	) name2152 (
		\mix1_data_o_reg_reg[76]/NET0131 ,
		_w2774_,
		_w2775_,
		_w3080_,
		_w3081_
	);
	LUT4 #(
		.INIT('h0545)
	) name2153 (
		\sub1_data_reg_reg[76]/NET0131 ,
		\sub1_ready_o_reg/NET0131 ,
		_w1054_,
		_w2230_,
		_w3082_
	);
	LUT4 #(
		.INIT('h1510)
	) name2154 (
		\state_reg/NET0131 ,
		\sub1_data_reg_reg[76]/NET0131 ,
		_w996_,
		_w3079_,
		_w3083_
	);
	LUT4 #(
		.INIT('h0057)
	) name2155 (
		\state_reg/NET0131 ,
		_w3081_,
		_w3082_,
		_w3083_,
		_w3084_
	);
	LUT3 #(
		.INIT('h48)
	) name2156 (
		\key_i[76]_pad ,
		_w931_,
		_w3084_,
		_w3085_
	);
	LUT4 #(
		.INIT('h3222)
	) name2157 (
		\data_o[76]_pad ,
		_w931_,
		_w934_,
		_w2784_,
		_w3086_
	);
	LUT4 #(
		.INIT('h7b00)
	) name2158 (
		\ks1_key_reg_reg[76]/P0002 ,
		_w2785_,
		_w3084_,
		_w3086_,
		_w3087_
	);
	LUT2 #(
		.INIT('he)
	) name2159 (
		_w3085_,
		_w3087_,
		_w3088_
	);
	LUT4 #(
		.INIT('h5547)
	) name2160 (
		\data_i[77]_pad ,
		decrypt_i_pad,
		\mix1_data_o_reg_reg[77]/NET0131 ,
		_w930_,
		_w3089_
	);
	LUT4 #(
		.INIT('ha8ab)
	) name2161 (
		\sub1_data_reg_reg[77]/NET0131 ,
		_w996_,
		_w2776_,
		_w3089_,
		_w3090_
	);
	LUT4 #(
		.INIT('h404c)
	) name2162 (
		\mix1_data_o_reg_reg[77]/NET0131 ,
		_w2774_,
		_w2775_,
		_w3090_,
		_w3091_
	);
	LUT4 #(
		.INIT('h0545)
	) name2163 (
		\sub1_data_reg_reg[77]/NET0131 ,
		\sub1_ready_o_reg/NET0131 ,
		_w1054_,
		_w2230_,
		_w3092_
	);
	LUT4 #(
		.INIT('h1510)
	) name2164 (
		\state_reg/NET0131 ,
		\sub1_data_reg_reg[77]/NET0131 ,
		_w996_,
		_w3089_,
		_w3093_
	);
	LUT4 #(
		.INIT('h0057)
	) name2165 (
		\state_reg/NET0131 ,
		_w3091_,
		_w3092_,
		_w3093_,
		_w3094_
	);
	LUT3 #(
		.INIT('h48)
	) name2166 (
		\key_i[77]_pad ,
		_w931_,
		_w3094_,
		_w3095_
	);
	LUT4 #(
		.INIT('h3222)
	) name2167 (
		\data_o[77]_pad ,
		_w931_,
		_w934_,
		_w2784_,
		_w3096_
	);
	LUT4 #(
		.INIT('h7b00)
	) name2168 (
		\ks1_key_reg_reg[77]/P0002 ,
		_w2785_,
		_w3094_,
		_w3096_,
		_w3097_
	);
	LUT2 #(
		.INIT('he)
	) name2169 (
		_w3095_,
		_w3097_,
		_w3098_
	);
	LUT4 #(
		.INIT('h5547)
	) name2170 (
		\data_i[26]_pad ,
		decrypt_i_pad,
		\mix1_data_o_reg_reg[26]/NET0131 ,
		_w930_,
		_w3099_
	);
	LUT4 #(
		.INIT('ha8ab)
	) name2171 (
		\sub1_data_reg_reg[26]/NET0131 ,
		_w996_,
		_w2776_,
		_w3099_,
		_w3100_
	);
	LUT4 #(
		.INIT('h404c)
	) name2172 (
		\mix1_data_o_reg_reg[26]/NET0131 ,
		_w2774_,
		_w2775_,
		_w3100_,
		_w3101_
	);
	LUT4 #(
		.INIT('h0545)
	) name2173 (
		\sub1_data_reg_reg[26]/NET0131 ,
		\sub1_ready_o_reg/NET0131 ,
		_w1054_,
		_w2230_,
		_w3102_
	);
	LUT4 #(
		.INIT('h1510)
	) name2174 (
		\state_reg/NET0131 ,
		\sub1_data_reg_reg[26]/NET0131 ,
		_w996_,
		_w3099_,
		_w3103_
	);
	LUT4 #(
		.INIT('h0057)
	) name2175 (
		\state_reg/NET0131 ,
		_w3101_,
		_w3102_,
		_w3103_,
		_w3104_
	);
	LUT3 #(
		.INIT('h48)
	) name2176 (
		\key_i[26]_pad ,
		_w931_,
		_w3104_,
		_w3105_
	);
	LUT4 #(
		.INIT('h3222)
	) name2177 (
		\data_o[26]_pad ,
		_w931_,
		_w934_,
		_w2784_,
		_w3106_
	);
	LUT4 #(
		.INIT('h7b00)
	) name2178 (
		\ks1_key_reg_reg[26]/NET0131 ,
		_w2785_,
		_w3104_,
		_w3106_,
		_w3107_
	);
	LUT2 #(
		.INIT('he)
	) name2179 (
		_w3105_,
		_w3107_,
		_w3108_
	);
	LUT4 #(
		.INIT('haab8)
	) name2180 (
		\data_i[103]_pad ,
		decrypt_i_pad,
		\mix1_data_o_reg_reg[103]/NET0131 ,
		_w930_,
		_w3109_
	);
	LUT4 #(
		.INIT('haba8)
	) name2181 (
		\sub1_data_reg_reg[103]/NET0131 ,
		_w996_,
		_w2776_,
		_w3109_,
		_w3110_
	);
	LUT4 #(
		.INIT('h404c)
	) name2182 (
		\mix1_data_o_reg_reg[103]/NET0131 ,
		_w2774_,
		_w2775_,
		_w3110_,
		_w3111_
	);
	LUT4 #(
		.INIT('h0545)
	) name2183 (
		\sub1_data_reg_reg[103]/NET0131 ,
		\sub1_ready_o_reg/NET0131 ,
		_w1054_,
		_w2230_,
		_w3112_
	);
	LUT4 #(
		.INIT('h1015)
	) name2184 (
		\state_reg/NET0131 ,
		\sub1_data_reg_reg[103]/NET0131 ,
		_w996_,
		_w3109_,
		_w3113_
	);
	LUT4 #(
		.INIT('h0057)
	) name2185 (
		\state_reg/NET0131 ,
		_w3111_,
		_w3112_,
		_w3113_,
		_w3114_
	);
	LUT3 #(
		.INIT('h48)
	) name2186 (
		\key_i[103]_pad ,
		_w931_,
		_w3114_,
		_w3115_
	);
	LUT4 #(
		.INIT('h3222)
	) name2187 (
		\data_o[103]_pad ,
		_w931_,
		_w934_,
		_w2784_,
		_w3116_
	);
	LUT4 #(
		.INIT('h7b00)
	) name2188 (
		\ks1_key_reg_reg[103]/NET0131 ,
		_w2785_,
		_w3114_,
		_w3116_,
		_w3117_
	);
	LUT2 #(
		.INIT('he)
	) name2189 (
		_w3115_,
		_w3117_,
		_w3118_
	);
	LUT4 #(
		.INIT('h5547)
	) name2190 (
		\data_i[78]_pad ,
		decrypt_i_pad,
		\mix1_data_o_reg_reg[78]/NET0131 ,
		_w930_,
		_w3119_
	);
	LUT4 #(
		.INIT('ha8ab)
	) name2191 (
		\sub1_data_reg_reg[78]/NET0131 ,
		_w996_,
		_w2776_,
		_w3119_,
		_w3120_
	);
	LUT4 #(
		.INIT('h404c)
	) name2192 (
		\mix1_data_o_reg_reg[78]/NET0131 ,
		_w2774_,
		_w2775_,
		_w3120_,
		_w3121_
	);
	LUT4 #(
		.INIT('h0545)
	) name2193 (
		\sub1_data_reg_reg[78]/NET0131 ,
		\sub1_ready_o_reg/NET0131 ,
		_w1054_,
		_w2230_,
		_w3122_
	);
	LUT4 #(
		.INIT('h1510)
	) name2194 (
		\state_reg/NET0131 ,
		\sub1_data_reg_reg[78]/NET0131 ,
		_w996_,
		_w3119_,
		_w3123_
	);
	LUT4 #(
		.INIT('h0057)
	) name2195 (
		\state_reg/NET0131 ,
		_w3121_,
		_w3122_,
		_w3123_,
		_w3124_
	);
	LUT3 #(
		.INIT('h48)
	) name2196 (
		\key_i[78]_pad ,
		_w931_,
		_w3124_,
		_w3125_
	);
	LUT4 #(
		.INIT('h3222)
	) name2197 (
		\data_o[78]_pad ,
		_w931_,
		_w934_,
		_w2784_,
		_w3126_
	);
	LUT4 #(
		.INIT('h7b00)
	) name2198 (
		\ks1_key_reg_reg[78]/P0002 ,
		_w2785_,
		_w3124_,
		_w3126_,
		_w3127_
	);
	LUT2 #(
		.INIT('he)
	) name2199 (
		_w3125_,
		_w3127_,
		_w3128_
	);
	LUT4 #(
		.INIT('haab8)
	) name2200 (
		\data_i[116]_pad ,
		decrypt_i_pad,
		\mix1_data_o_reg_reg[116]/NET0131 ,
		_w930_,
		_w3129_
	);
	LUT4 #(
		.INIT('haba8)
	) name2201 (
		\sub1_data_reg_reg[116]/NET0131 ,
		_w996_,
		_w2776_,
		_w3129_,
		_w3130_
	);
	LUT4 #(
		.INIT('h404c)
	) name2202 (
		\mix1_data_o_reg_reg[116]/NET0131 ,
		_w2774_,
		_w2775_,
		_w3130_,
		_w3131_
	);
	LUT4 #(
		.INIT('h0545)
	) name2203 (
		\sub1_data_reg_reg[116]/NET0131 ,
		\sub1_ready_o_reg/NET0131 ,
		_w1054_,
		_w2230_,
		_w3132_
	);
	LUT4 #(
		.INIT('h1015)
	) name2204 (
		\state_reg/NET0131 ,
		\sub1_data_reg_reg[116]/NET0131 ,
		_w996_,
		_w3129_,
		_w3133_
	);
	LUT4 #(
		.INIT('h0057)
	) name2205 (
		\state_reg/NET0131 ,
		_w3131_,
		_w3132_,
		_w3133_,
		_w3134_
	);
	LUT3 #(
		.INIT('h48)
	) name2206 (
		\key_i[116]_pad ,
		_w931_,
		_w3134_,
		_w3135_
	);
	LUT4 #(
		.INIT('h3222)
	) name2207 (
		\data_o[116]_pad ,
		_w931_,
		_w934_,
		_w2784_,
		_w3136_
	);
	LUT4 #(
		.INIT('h7b00)
	) name2208 (
		\ks1_key_reg_reg[116]/NET0131 ,
		_w2785_,
		_w3134_,
		_w3136_,
		_w3137_
	);
	LUT2 #(
		.INIT('he)
	) name2209 (
		_w3135_,
		_w3137_,
		_w3138_
	);
	LUT4 #(
		.INIT('h5547)
	) name2210 (
		\data_i[79]_pad ,
		decrypt_i_pad,
		\mix1_data_o_reg_reg[79]/NET0131 ,
		_w930_,
		_w3139_
	);
	LUT4 #(
		.INIT('ha8ab)
	) name2211 (
		\sub1_data_reg_reg[79]/NET0131 ,
		_w996_,
		_w2776_,
		_w3139_,
		_w3140_
	);
	LUT4 #(
		.INIT('h404c)
	) name2212 (
		\mix1_data_o_reg_reg[79]/NET0131 ,
		_w2774_,
		_w2775_,
		_w3140_,
		_w3141_
	);
	LUT4 #(
		.INIT('h0545)
	) name2213 (
		\sub1_data_reg_reg[79]/NET0131 ,
		\sub1_ready_o_reg/NET0131 ,
		_w1054_,
		_w2230_,
		_w3142_
	);
	LUT4 #(
		.INIT('h1510)
	) name2214 (
		\state_reg/NET0131 ,
		\sub1_data_reg_reg[79]/NET0131 ,
		_w996_,
		_w3139_,
		_w3143_
	);
	LUT4 #(
		.INIT('h0057)
	) name2215 (
		\state_reg/NET0131 ,
		_w3141_,
		_w3142_,
		_w3143_,
		_w3144_
	);
	LUT3 #(
		.INIT('h48)
	) name2216 (
		\key_i[79]_pad ,
		_w931_,
		_w3144_,
		_w3145_
	);
	LUT4 #(
		.INIT('h3222)
	) name2217 (
		\data_o[79]_pad ,
		_w931_,
		_w934_,
		_w2784_,
		_w3146_
	);
	LUT4 #(
		.INIT('h7b00)
	) name2218 (
		\ks1_key_reg_reg[79]/P0002 ,
		_w2785_,
		_w3144_,
		_w3146_,
		_w3147_
	);
	LUT2 #(
		.INIT('he)
	) name2219 (
		_w3145_,
		_w3147_,
		_w3148_
	);
	LUT4 #(
		.INIT('h5547)
	) name2220 (
		\data_i[27]_pad ,
		decrypt_i_pad,
		\mix1_data_o_reg_reg[27]/NET0131 ,
		_w930_,
		_w3149_
	);
	LUT4 #(
		.INIT('ha8ab)
	) name2221 (
		\sub1_data_reg_reg[27]/NET0131 ,
		_w996_,
		_w2776_,
		_w3149_,
		_w3150_
	);
	LUT4 #(
		.INIT('h404c)
	) name2222 (
		\mix1_data_o_reg_reg[27]/NET0131 ,
		_w2774_,
		_w2775_,
		_w3150_,
		_w3151_
	);
	LUT4 #(
		.INIT('h0545)
	) name2223 (
		\sub1_data_reg_reg[27]/NET0131 ,
		\sub1_ready_o_reg/NET0131 ,
		_w1054_,
		_w2230_,
		_w3152_
	);
	LUT4 #(
		.INIT('h1510)
	) name2224 (
		\state_reg/NET0131 ,
		\sub1_data_reg_reg[27]/NET0131 ,
		_w996_,
		_w3149_,
		_w3153_
	);
	LUT4 #(
		.INIT('h0057)
	) name2225 (
		\state_reg/NET0131 ,
		_w3151_,
		_w3152_,
		_w3153_,
		_w3154_
	);
	LUT3 #(
		.INIT('h48)
	) name2226 (
		\key_i[27]_pad ,
		_w931_,
		_w3154_,
		_w3155_
	);
	LUT4 #(
		.INIT('h3222)
	) name2227 (
		\data_o[27]_pad ,
		_w931_,
		_w934_,
		_w2784_,
		_w3156_
	);
	LUT4 #(
		.INIT('h7b00)
	) name2228 (
		\ks1_key_reg_reg[27]/NET0131 ,
		_w2785_,
		_w3154_,
		_w3156_,
		_w3157_
	);
	LUT2 #(
		.INIT('he)
	) name2229 (
		_w3155_,
		_w3157_,
		_w3158_
	);
	LUT4 #(
		.INIT('h5547)
	) name2230 (
		\data_i[7]_pad ,
		decrypt_i_pad,
		\mix1_data_o_reg_reg[7]/NET0131 ,
		_w930_,
		_w3159_
	);
	LUT4 #(
		.INIT('ha8ab)
	) name2231 (
		\sub1_data_reg_reg[7]/NET0131 ,
		_w996_,
		_w2776_,
		_w3159_,
		_w3160_
	);
	LUT4 #(
		.INIT('h404c)
	) name2232 (
		\mix1_data_o_reg_reg[7]/NET0131 ,
		_w2774_,
		_w2775_,
		_w3160_,
		_w3161_
	);
	LUT4 #(
		.INIT('h0545)
	) name2233 (
		\sub1_data_reg_reg[7]/NET0131 ,
		\sub1_ready_o_reg/NET0131 ,
		_w1054_,
		_w2230_,
		_w3162_
	);
	LUT4 #(
		.INIT('h1510)
	) name2234 (
		\state_reg/NET0131 ,
		\sub1_data_reg_reg[7]/NET0131 ,
		_w996_,
		_w3159_,
		_w3163_
	);
	LUT4 #(
		.INIT('h0057)
	) name2235 (
		\state_reg/NET0131 ,
		_w3161_,
		_w3162_,
		_w3163_,
		_w3164_
	);
	LUT3 #(
		.INIT('h48)
	) name2236 (
		\key_i[7]_pad ,
		_w931_,
		_w3164_,
		_w3165_
	);
	LUT4 #(
		.INIT('h3222)
	) name2237 (
		\data_o[7]_pad ,
		_w931_,
		_w934_,
		_w2784_,
		_w3166_
	);
	LUT4 #(
		.INIT('h7b00)
	) name2238 (
		\ks1_key_reg_reg[7]/NET0131 ,
		_w2785_,
		_w3164_,
		_w3166_,
		_w3167_
	);
	LUT2 #(
		.INIT('he)
	) name2239 (
		_w3165_,
		_w3167_,
		_w3168_
	);
	LUT4 #(
		.INIT('haab8)
	) name2240 (
		\data_i[117]_pad ,
		decrypt_i_pad,
		\mix1_data_o_reg_reg[117]/NET0131 ,
		_w930_,
		_w3169_
	);
	LUT4 #(
		.INIT('haba8)
	) name2241 (
		\sub1_data_reg_reg[117]/NET0131 ,
		_w996_,
		_w2776_,
		_w3169_,
		_w3170_
	);
	LUT4 #(
		.INIT('h404c)
	) name2242 (
		\mix1_data_o_reg_reg[117]/NET0131 ,
		_w2774_,
		_w2775_,
		_w3170_,
		_w3171_
	);
	LUT4 #(
		.INIT('h0545)
	) name2243 (
		\sub1_data_reg_reg[117]/NET0131 ,
		\sub1_ready_o_reg/NET0131 ,
		_w1054_,
		_w2230_,
		_w3172_
	);
	LUT4 #(
		.INIT('h1015)
	) name2244 (
		\state_reg/NET0131 ,
		\sub1_data_reg_reg[117]/NET0131 ,
		_w996_,
		_w3169_,
		_w3173_
	);
	LUT4 #(
		.INIT('h0057)
	) name2245 (
		\state_reg/NET0131 ,
		_w3171_,
		_w3172_,
		_w3173_,
		_w3174_
	);
	LUT3 #(
		.INIT('h48)
	) name2246 (
		\key_i[117]_pad ,
		_w931_,
		_w3174_,
		_w3175_
	);
	LUT4 #(
		.INIT('h3222)
	) name2247 (
		\data_o[117]_pad ,
		_w931_,
		_w934_,
		_w2784_,
		_w3176_
	);
	LUT4 #(
		.INIT('h7b00)
	) name2248 (
		\ks1_key_reg_reg[117]/NET0131 ,
		_w2785_,
		_w3174_,
		_w3176_,
		_w3177_
	);
	LUT2 #(
		.INIT('he)
	) name2249 (
		_w3175_,
		_w3177_,
		_w3178_
	);
	LUT4 #(
		.INIT('haab8)
	) name2250 (
		\data_i[80]_pad ,
		decrypt_i_pad,
		\mix1_data_o_reg_reg[80]/NET0131 ,
		_w930_,
		_w3179_
	);
	LUT4 #(
		.INIT('haba8)
	) name2251 (
		\sub1_data_reg_reg[80]/NET0131 ,
		_w996_,
		_w2776_,
		_w3179_,
		_w3180_
	);
	LUT4 #(
		.INIT('h404c)
	) name2252 (
		\mix1_data_o_reg_reg[80]/NET0131 ,
		_w2774_,
		_w2775_,
		_w3180_,
		_w3181_
	);
	LUT4 #(
		.INIT('h0545)
	) name2253 (
		\sub1_data_reg_reg[80]/NET0131 ,
		\sub1_ready_o_reg/NET0131 ,
		_w1054_,
		_w2230_,
		_w3182_
	);
	LUT4 #(
		.INIT('h1015)
	) name2254 (
		\state_reg/NET0131 ,
		\sub1_data_reg_reg[80]/NET0131 ,
		_w996_,
		_w3179_,
		_w3183_
	);
	LUT4 #(
		.INIT('h0057)
	) name2255 (
		\state_reg/NET0131 ,
		_w3181_,
		_w3182_,
		_w3183_,
		_w3184_
	);
	LUT3 #(
		.INIT('h48)
	) name2256 (
		\key_i[80]_pad ,
		_w931_,
		_w3184_,
		_w3185_
	);
	LUT4 #(
		.INIT('h3222)
	) name2257 (
		\data_o[80]_pad ,
		_w931_,
		_w934_,
		_w2784_,
		_w3186_
	);
	LUT4 #(
		.INIT('h7b00)
	) name2258 (
		\ks1_key_reg_reg[80]/NET0131 ,
		_w2785_,
		_w3184_,
		_w3186_,
		_w3187_
	);
	LUT2 #(
		.INIT('he)
	) name2259 (
		_w3185_,
		_w3187_,
		_w3188_
	);
	LUT4 #(
		.INIT('h5547)
	) name2260 (
		\data_i[28]_pad ,
		decrypt_i_pad,
		\mix1_data_o_reg_reg[28]/NET0131 ,
		_w930_,
		_w3189_
	);
	LUT4 #(
		.INIT('ha8ab)
	) name2261 (
		\sub1_data_reg_reg[28]/NET0131 ,
		_w996_,
		_w2776_,
		_w3189_,
		_w3190_
	);
	LUT4 #(
		.INIT('h404c)
	) name2262 (
		\mix1_data_o_reg_reg[28]/NET0131 ,
		_w2774_,
		_w2775_,
		_w3190_,
		_w3191_
	);
	LUT4 #(
		.INIT('h0545)
	) name2263 (
		\sub1_data_reg_reg[28]/NET0131 ,
		\sub1_ready_o_reg/NET0131 ,
		_w1054_,
		_w2230_,
		_w3192_
	);
	LUT4 #(
		.INIT('h1510)
	) name2264 (
		\state_reg/NET0131 ,
		\sub1_data_reg_reg[28]/NET0131 ,
		_w996_,
		_w3189_,
		_w3193_
	);
	LUT4 #(
		.INIT('h0057)
	) name2265 (
		\state_reg/NET0131 ,
		_w3191_,
		_w3192_,
		_w3193_,
		_w3194_
	);
	LUT3 #(
		.INIT('h48)
	) name2266 (
		\key_i[28]_pad ,
		_w931_,
		_w3194_,
		_w3195_
	);
	LUT4 #(
		.INIT('h3222)
	) name2267 (
		\data_o[28]_pad ,
		_w931_,
		_w934_,
		_w2784_,
		_w3196_
	);
	LUT4 #(
		.INIT('h7b00)
	) name2268 (
		\ks1_key_reg_reg[28]/NET0131 ,
		_w2785_,
		_w3194_,
		_w3196_,
		_w3197_
	);
	LUT2 #(
		.INIT('he)
	) name2269 (
		_w3195_,
		_w3197_,
		_w3198_
	);
	LUT4 #(
		.INIT('haab8)
	) name2270 (
		\data_i[81]_pad ,
		decrypt_i_pad,
		\mix1_data_o_reg_reg[81]/NET0131 ,
		_w930_,
		_w3199_
	);
	LUT4 #(
		.INIT('haba8)
	) name2271 (
		\sub1_data_reg_reg[81]/NET0131 ,
		_w996_,
		_w2776_,
		_w3199_,
		_w3200_
	);
	LUT4 #(
		.INIT('h404c)
	) name2272 (
		\mix1_data_o_reg_reg[81]/NET0131 ,
		_w2774_,
		_w2775_,
		_w3200_,
		_w3201_
	);
	LUT4 #(
		.INIT('h0545)
	) name2273 (
		\sub1_data_reg_reg[81]/NET0131 ,
		\sub1_ready_o_reg/NET0131 ,
		_w1054_,
		_w2230_,
		_w3202_
	);
	LUT4 #(
		.INIT('h1015)
	) name2274 (
		\state_reg/NET0131 ,
		\sub1_data_reg_reg[81]/NET0131 ,
		_w996_,
		_w3199_,
		_w3203_
	);
	LUT4 #(
		.INIT('h0057)
	) name2275 (
		\state_reg/NET0131 ,
		_w3201_,
		_w3202_,
		_w3203_,
		_w3204_
	);
	LUT3 #(
		.INIT('h48)
	) name2276 (
		\key_i[81]_pad ,
		_w931_,
		_w3204_,
		_w3205_
	);
	LUT4 #(
		.INIT('h3222)
	) name2277 (
		\data_o[81]_pad ,
		_w931_,
		_w934_,
		_w2784_,
		_w3206_
	);
	LUT4 #(
		.INIT('h7b00)
	) name2278 (
		\ks1_key_reg_reg[81]/NET0131 ,
		_w2785_,
		_w3204_,
		_w3206_,
		_w3207_
	);
	LUT2 #(
		.INIT('he)
	) name2279 (
		_w3205_,
		_w3207_,
		_w3208_
	);
	LUT4 #(
		.INIT('haab8)
	) name2280 (
		\data_i[82]_pad ,
		decrypt_i_pad,
		\mix1_data_o_reg_reg[82]/NET0131 ,
		_w930_,
		_w3209_
	);
	LUT4 #(
		.INIT('haba8)
	) name2281 (
		\sub1_data_reg_reg[82]/NET0131 ,
		_w996_,
		_w2776_,
		_w3209_,
		_w3210_
	);
	LUT4 #(
		.INIT('h404c)
	) name2282 (
		\mix1_data_o_reg_reg[82]/NET0131 ,
		_w2774_,
		_w2775_,
		_w3210_,
		_w3211_
	);
	LUT4 #(
		.INIT('h0545)
	) name2283 (
		\sub1_data_reg_reg[82]/NET0131 ,
		\sub1_ready_o_reg/NET0131 ,
		_w1054_,
		_w2230_,
		_w3212_
	);
	LUT4 #(
		.INIT('h1015)
	) name2284 (
		\state_reg/NET0131 ,
		\sub1_data_reg_reg[82]/NET0131 ,
		_w996_,
		_w3209_,
		_w3213_
	);
	LUT4 #(
		.INIT('h0057)
	) name2285 (
		\state_reg/NET0131 ,
		_w3211_,
		_w3212_,
		_w3213_,
		_w3214_
	);
	LUT3 #(
		.INIT('h48)
	) name2286 (
		\key_i[82]_pad ,
		_w931_,
		_w3214_,
		_w3215_
	);
	LUT4 #(
		.INIT('h3222)
	) name2287 (
		\data_o[82]_pad ,
		_w931_,
		_w934_,
		_w2784_,
		_w3216_
	);
	LUT4 #(
		.INIT('h7b00)
	) name2288 (
		\ks1_key_reg_reg[82]/NET0131 ,
		_w2785_,
		_w3214_,
		_w3216_,
		_w3217_
	);
	LUT2 #(
		.INIT('he)
	) name2289 (
		_w3215_,
		_w3217_,
		_w3218_
	);
	LUT4 #(
		.INIT('h5547)
	) name2290 (
		\data_i[29]_pad ,
		decrypt_i_pad,
		\mix1_data_o_reg_reg[29]/NET0131 ,
		_w930_,
		_w3219_
	);
	LUT4 #(
		.INIT('ha8ab)
	) name2291 (
		\sub1_data_reg_reg[29]/NET0131 ,
		_w996_,
		_w2776_,
		_w3219_,
		_w3220_
	);
	LUT4 #(
		.INIT('h404c)
	) name2292 (
		\mix1_data_o_reg_reg[29]/NET0131 ,
		_w2774_,
		_w2775_,
		_w3220_,
		_w3221_
	);
	LUT4 #(
		.INIT('h0545)
	) name2293 (
		\sub1_data_reg_reg[29]/NET0131 ,
		\sub1_ready_o_reg/NET0131 ,
		_w1054_,
		_w2230_,
		_w3222_
	);
	LUT4 #(
		.INIT('h1510)
	) name2294 (
		\state_reg/NET0131 ,
		\sub1_data_reg_reg[29]/NET0131 ,
		_w996_,
		_w3219_,
		_w3223_
	);
	LUT4 #(
		.INIT('h0057)
	) name2295 (
		\state_reg/NET0131 ,
		_w3221_,
		_w3222_,
		_w3223_,
		_w3224_
	);
	LUT3 #(
		.INIT('h48)
	) name2296 (
		\key_i[29]_pad ,
		_w931_,
		_w3224_,
		_w3225_
	);
	LUT4 #(
		.INIT('h3222)
	) name2297 (
		\data_o[29]_pad ,
		_w931_,
		_w934_,
		_w2784_,
		_w3226_
	);
	LUT4 #(
		.INIT('h7b00)
	) name2298 (
		\ks1_key_reg_reg[29]/NET0131 ,
		_w2785_,
		_w3224_,
		_w3226_,
		_w3227_
	);
	LUT2 #(
		.INIT('he)
	) name2299 (
		_w3225_,
		_w3227_,
		_w3228_
	);
	LUT4 #(
		.INIT('haab8)
	) name2300 (
		\data_i[83]_pad ,
		decrypt_i_pad,
		\mix1_data_o_reg_reg[83]/NET0131 ,
		_w930_,
		_w3229_
	);
	LUT4 #(
		.INIT('haba8)
	) name2301 (
		\sub1_data_reg_reg[83]/NET0131 ,
		_w996_,
		_w2776_,
		_w3229_,
		_w3230_
	);
	LUT4 #(
		.INIT('h404c)
	) name2302 (
		\mix1_data_o_reg_reg[83]/NET0131 ,
		_w2774_,
		_w2775_,
		_w3230_,
		_w3231_
	);
	LUT4 #(
		.INIT('h0545)
	) name2303 (
		\sub1_data_reg_reg[83]/NET0131 ,
		\sub1_ready_o_reg/NET0131 ,
		_w1054_,
		_w2230_,
		_w3232_
	);
	LUT4 #(
		.INIT('h1015)
	) name2304 (
		\state_reg/NET0131 ,
		\sub1_data_reg_reg[83]/NET0131 ,
		_w996_,
		_w3229_,
		_w3233_
	);
	LUT4 #(
		.INIT('h0057)
	) name2305 (
		\state_reg/NET0131 ,
		_w3231_,
		_w3232_,
		_w3233_,
		_w3234_
	);
	LUT3 #(
		.INIT('h48)
	) name2306 (
		\key_i[83]_pad ,
		_w931_,
		_w3234_,
		_w3235_
	);
	LUT4 #(
		.INIT('h3222)
	) name2307 (
		\data_o[83]_pad ,
		_w931_,
		_w934_,
		_w2784_,
		_w3236_
	);
	LUT4 #(
		.INIT('h7b00)
	) name2308 (
		\ks1_key_reg_reg[83]/NET0131 ,
		_w2785_,
		_w3234_,
		_w3236_,
		_w3237_
	);
	LUT2 #(
		.INIT('he)
	) name2309 (
		_w3235_,
		_w3237_,
		_w3238_
	);
	LUT4 #(
		.INIT('haab8)
	) name2310 (
		\data_i[84]_pad ,
		decrypt_i_pad,
		\mix1_data_o_reg_reg[84]/NET0131 ,
		_w930_,
		_w3239_
	);
	LUT4 #(
		.INIT('haba8)
	) name2311 (
		\sub1_data_reg_reg[84]/NET0131 ,
		_w996_,
		_w2776_,
		_w3239_,
		_w3240_
	);
	LUT4 #(
		.INIT('h404c)
	) name2312 (
		\mix1_data_o_reg_reg[84]/NET0131 ,
		_w2774_,
		_w2775_,
		_w3240_,
		_w3241_
	);
	LUT4 #(
		.INIT('h0545)
	) name2313 (
		\sub1_data_reg_reg[84]/NET0131 ,
		\sub1_ready_o_reg/NET0131 ,
		_w1054_,
		_w2230_,
		_w3242_
	);
	LUT4 #(
		.INIT('h1015)
	) name2314 (
		\state_reg/NET0131 ,
		\sub1_data_reg_reg[84]/NET0131 ,
		_w996_,
		_w3239_,
		_w3243_
	);
	LUT4 #(
		.INIT('h0057)
	) name2315 (
		\state_reg/NET0131 ,
		_w3241_,
		_w3242_,
		_w3243_,
		_w3244_
	);
	LUT3 #(
		.INIT('h48)
	) name2316 (
		\key_i[84]_pad ,
		_w931_,
		_w3244_,
		_w3245_
	);
	LUT4 #(
		.INIT('h3222)
	) name2317 (
		\data_o[84]_pad ,
		_w931_,
		_w934_,
		_w2784_,
		_w3246_
	);
	LUT4 #(
		.INIT('h7b00)
	) name2318 (
		\ks1_key_reg_reg[84]/NET0131 ,
		_w2785_,
		_w3244_,
		_w3246_,
		_w3247_
	);
	LUT2 #(
		.INIT('he)
	) name2319 (
		_w3245_,
		_w3247_,
		_w3248_
	);
	LUT4 #(
		.INIT('haab8)
	) name2320 (
		\data_i[118]_pad ,
		decrypt_i_pad,
		\mix1_data_o_reg_reg[118]/NET0131 ,
		_w930_,
		_w3249_
	);
	LUT4 #(
		.INIT('haba8)
	) name2321 (
		\sub1_data_reg_reg[118]/NET0131 ,
		_w996_,
		_w2776_,
		_w3249_,
		_w3250_
	);
	LUT4 #(
		.INIT('h404c)
	) name2322 (
		\mix1_data_o_reg_reg[118]/NET0131 ,
		_w2774_,
		_w2775_,
		_w3250_,
		_w3251_
	);
	LUT4 #(
		.INIT('h0545)
	) name2323 (
		\sub1_data_reg_reg[118]/NET0131 ,
		\sub1_ready_o_reg/NET0131 ,
		_w1054_,
		_w2230_,
		_w3252_
	);
	LUT4 #(
		.INIT('h1015)
	) name2324 (
		\state_reg/NET0131 ,
		\sub1_data_reg_reg[118]/NET0131 ,
		_w996_,
		_w3249_,
		_w3253_
	);
	LUT4 #(
		.INIT('h0057)
	) name2325 (
		\state_reg/NET0131 ,
		_w3251_,
		_w3252_,
		_w3253_,
		_w3254_
	);
	LUT3 #(
		.INIT('h48)
	) name2326 (
		\key_i[118]_pad ,
		_w931_,
		_w3254_,
		_w3255_
	);
	LUT4 #(
		.INIT('h3222)
	) name2327 (
		\data_o[118]_pad ,
		_w931_,
		_w934_,
		_w2784_,
		_w3256_
	);
	LUT4 #(
		.INIT('h7b00)
	) name2328 (
		\ks1_key_reg_reg[118]/NET0131 ,
		_w2785_,
		_w3254_,
		_w3256_,
		_w3257_
	);
	LUT2 #(
		.INIT('he)
	) name2329 (
		_w3255_,
		_w3257_,
		_w3258_
	);
	LUT4 #(
		.INIT('h5547)
	) name2330 (
		\data_i[2]_pad ,
		decrypt_i_pad,
		\mix1_data_o_reg_reg[2]/NET0131 ,
		_w930_,
		_w3259_
	);
	LUT4 #(
		.INIT('ha8ab)
	) name2331 (
		\sub1_data_reg_reg[2]/NET0131 ,
		_w996_,
		_w2776_,
		_w3259_,
		_w3260_
	);
	LUT4 #(
		.INIT('h404c)
	) name2332 (
		\mix1_data_o_reg_reg[2]/NET0131 ,
		_w2774_,
		_w2775_,
		_w3260_,
		_w3261_
	);
	LUT4 #(
		.INIT('h0545)
	) name2333 (
		\sub1_data_reg_reg[2]/NET0131 ,
		\sub1_ready_o_reg/NET0131 ,
		_w1054_,
		_w2230_,
		_w3262_
	);
	LUT4 #(
		.INIT('h1510)
	) name2334 (
		\state_reg/NET0131 ,
		\sub1_data_reg_reg[2]/NET0131 ,
		_w996_,
		_w3259_,
		_w3263_
	);
	LUT4 #(
		.INIT('h0057)
	) name2335 (
		\state_reg/NET0131 ,
		_w3261_,
		_w3262_,
		_w3263_,
		_w3264_
	);
	LUT3 #(
		.INIT('h48)
	) name2336 (
		\key_i[2]_pad ,
		_w931_,
		_w3264_,
		_w3265_
	);
	LUT4 #(
		.INIT('h3222)
	) name2337 (
		\data_o[2]_pad ,
		_w931_,
		_w934_,
		_w2784_,
		_w3266_
	);
	LUT4 #(
		.INIT('h7b00)
	) name2338 (
		\ks1_key_reg_reg[2]/NET0131 ,
		_w2785_,
		_w3264_,
		_w3266_,
		_w3267_
	);
	LUT2 #(
		.INIT('he)
	) name2339 (
		_w3265_,
		_w3267_,
		_w3268_
	);
	LUT4 #(
		.INIT('haab8)
	) name2340 (
		\data_i[85]_pad ,
		decrypt_i_pad,
		\mix1_data_o_reg_reg[85]/NET0131 ,
		_w930_,
		_w3269_
	);
	LUT4 #(
		.INIT('haba8)
	) name2341 (
		\sub1_data_reg_reg[85]/NET0131 ,
		_w996_,
		_w2776_,
		_w3269_,
		_w3270_
	);
	LUT4 #(
		.INIT('h404c)
	) name2342 (
		\mix1_data_o_reg_reg[85]/NET0131 ,
		_w2774_,
		_w2775_,
		_w3270_,
		_w3271_
	);
	LUT4 #(
		.INIT('h0545)
	) name2343 (
		\sub1_data_reg_reg[85]/NET0131 ,
		\sub1_ready_o_reg/NET0131 ,
		_w1054_,
		_w2230_,
		_w3272_
	);
	LUT4 #(
		.INIT('h1015)
	) name2344 (
		\state_reg/NET0131 ,
		\sub1_data_reg_reg[85]/NET0131 ,
		_w996_,
		_w3269_,
		_w3273_
	);
	LUT4 #(
		.INIT('h0057)
	) name2345 (
		\state_reg/NET0131 ,
		_w3271_,
		_w3272_,
		_w3273_,
		_w3274_
	);
	LUT3 #(
		.INIT('h48)
	) name2346 (
		\key_i[85]_pad ,
		_w931_,
		_w3274_,
		_w3275_
	);
	LUT4 #(
		.INIT('h3222)
	) name2347 (
		\data_o[85]_pad ,
		_w931_,
		_w934_,
		_w2784_,
		_w3276_
	);
	LUT4 #(
		.INIT('h7b00)
	) name2348 (
		\ks1_key_reg_reg[85]/NET0131 ,
		_w2785_,
		_w3274_,
		_w3276_,
		_w3277_
	);
	LUT2 #(
		.INIT('he)
	) name2349 (
		_w3275_,
		_w3277_,
		_w3278_
	);
	LUT4 #(
		.INIT('h5547)
	) name2350 (
		\data_i[30]_pad ,
		decrypt_i_pad,
		\mix1_data_o_reg_reg[30]/NET0131 ,
		_w930_,
		_w3279_
	);
	LUT4 #(
		.INIT('ha8ab)
	) name2351 (
		\sub1_data_reg_reg[30]/NET0131 ,
		_w996_,
		_w2776_,
		_w3279_,
		_w3280_
	);
	LUT4 #(
		.INIT('h404c)
	) name2352 (
		\mix1_data_o_reg_reg[30]/NET0131 ,
		_w2774_,
		_w2775_,
		_w3280_,
		_w3281_
	);
	LUT4 #(
		.INIT('h0545)
	) name2353 (
		\sub1_data_reg_reg[30]/NET0131 ,
		\sub1_ready_o_reg/NET0131 ,
		_w1054_,
		_w2230_,
		_w3282_
	);
	LUT4 #(
		.INIT('h1510)
	) name2354 (
		\state_reg/NET0131 ,
		\sub1_data_reg_reg[30]/NET0131 ,
		_w996_,
		_w3279_,
		_w3283_
	);
	LUT4 #(
		.INIT('h0057)
	) name2355 (
		\state_reg/NET0131 ,
		_w3281_,
		_w3282_,
		_w3283_,
		_w3284_
	);
	LUT3 #(
		.INIT('h48)
	) name2356 (
		\key_i[30]_pad ,
		_w931_,
		_w3284_,
		_w3285_
	);
	LUT4 #(
		.INIT('h3222)
	) name2357 (
		\data_o[30]_pad ,
		_w931_,
		_w934_,
		_w2784_,
		_w3286_
	);
	LUT4 #(
		.INIT('h7b00)
	) name2358 (
		\ks1_key_reg_reg[30]/NET0131 ,
		_w2785_,
		_w3284_,
		_w3286_,
		_w3287_
	);
	LUT2 #(
		.INIT('he)
	) name2359 (
		_w3285_,
		_w3287_,
		_w3288_
	);
	LUT4 #(
		.INIT('haab8)
	) name2360 (
		\data_i[86]_pad ,
		decrypt_i_pad,
		\mix1_data_o_reg_reg[86]/NET0131 ,
		_w930_,
		_w3289_
	);
	LUT4 #(
		.INIT('haba8)
	) name2361 (
		\sub1_data_reg_reg[86]/NET0131 ,
		_w996_,
		_w2776_,
		_w3289_,
		_w3290_
	);
	LUT4 #(
		.INIT('h404c)
	) name2362 (
		\mix1_data_o_reg_reg[86]/NET0131 ,
		_w2774_,
		_w2775_,
		_w3290_,
		_w3291_
	);
	LUT4 #(
		.INIT('h0545)
	) name2363 (
		\sub1_data_reg_reg[86]/NET0131 ,
		\sub1_ready_o_reg/NET0131 ,
		_w1054_,
		_w2230_,
		_w3292_
	);
	LUT4 #(
		.INIT('h1015)
	) name2364 (
		\state_reg/NET0131 ,
		\sub1_data_reg_reg[86]/NET0131 ,
		_w996_,
		_w3289_,
		_w3293_
	);
	LUT4 #(
		.INIT('h0057)
	) name2365 (
		\state_reg/NET0131 ,
		_w3291_,
		_w3292_,
		_w3293_,
		_w3294_
	);
	LUT3 #(
		.INIT('h48)
	) name2366 (
		\key_i[86]_pad ,
		_w931_,
		_w3294_,
		_w3295_
	);
	LUT4 #(
		.INIT('h3222)
	) name2367 (
		\data_o[86]_pad ,
		_w931_,
		_w934_,
		_w2784_,
		_w3296_
	);
	LUT4 #(
		.INIT('h7b00)
	) name2368 (
		\ks1_key_reg_reg[86]/NET0131 ,
		_w2785_,
		_w3294_,
		_w3296_,
		_w3297_
	);
	LUT2 #(
		.INIT('he)
	) name2369 (
		_w3295_,
		_w3297_,
		_w3298_
	);
	LUT4 #(
		.INIT('haab8)
	) name2370 (
		\data_i[87]_pad ,
		decrypt_i_pad,
		\mix1_data_o_reg_reg[87]/NET0131 ,
		_w930_,
		_w3299_
	);
	LUT4 #(
		.INIT('haba8)
	) name2371 (
		\sub1_data_reg_reg[87]/NET0131 ,
		_w996_,
		_w2776_,
		_w3299_,
		_w3300_
	);
	LUT4 #(
		.INIT('h404c)
	) name2372 (
		\mix1_data_o_reg_reg[87]/NET0131 ,
		_w2774_,
		_w2775_,
		_w3300_,
		_w3301_
	);
	LUT4 #(
		.INIT('h0545)
	) name2373 (
		\sub1_data_reg_reg[87]/NET0131 ,
		\sub1_ready_o_reg/NET0131 ,
		_w1054_,
		_w2230_,
		_w3302_
	);
	LUT4 #(
		.INIT('h1015)
	) name2374 (
		\state_reg/NET0131 ,
		\sub1_data_reg_reg[87]/NET0131 ,
		_w996_,
		_w3299_,
		_w3303_
	);
	LUT4 #(
		.INIT('h0057)
	) name2375 (
		\state_reg/NET0131 ,
		_w3301_,
		_w3302_,
		_w3303_,
		_w3304_
	);
	LUT3 #(
		.INIT('h48)
	) name2376 (
		\key_i[87]_pad ,
		_w931_,
		_w3304_,
		_w3305_
	);
	LUT4 #(
		.INIT('h3222)
	) name2377 (
		\data_o[87]_pad ,
		_w931_,
		_w934_,
		_w2784_,
		_w3306_
	);
	LUT4 #(
		.INIT('h7b00)
	) name2378 (
		\ks1_key_reg_reg[87]/NET0131 ,
		_w2785_,
		_w3304_,
		_w3306_,
		_w3307_
	);
	LUT2 #(
		.INIT('he)
	) name2379 (
		_w3305_,
		_w3307_,
		_w3308_
	);
	LUT4 #(
		.INIT('h5547)
	) name2380 (
		\data_i[31]_pad ,
		decrypt_i_pad,
		\mix1_data_o_reg_reg[31]/NET0131 ,
		_w930_,
		_w3309_
	);
	LUT4 #(
		.INIT('ha8ab)
	) name2381 (
		\sub1_data_reg_reg[31]/NET0131 ,
		_w996_,
		_w2776_,
		_w3309_,
		_w3310_
	);
	LUT4 #(
		.INIT('h404c)
	) name2382 (
		\mix1_data_o_reg_reg[31]/NET0131 ,
		_w2774_,
		_w2775_,
		_w3310_,
		_w3311_
	);
	LUT4 #(
		.INIT('h0545)
	) name2383 (
		\sub1_data_reg_reg[31]/NET0131 ,
		\sub1_ready_o_reg/NET0131 ,
		_w1054_,
		_w2230_,
		_w3312_
	);
	LUT4 #(
		.INIT('h1510)
	) name2384 (
		\state_reg/NET0131 ,
		\sub1_data_reg_reg[31]/NET0131 ,
		_w996_,
		_w3309_,
		_w3313_
	);
	LUT4 #(
		.INIT('h0057)
	) name2385 (
		\state_reg/NET0131 ,
		_w3311_,
		_w3312_,
		_w3313_,
		_w3314_
	);
	LUT3 #(
		.INIT('h48)
	) name2386 (
		\key_i[31]_pad ,
		_w931_,
		_w3314_,
		_w3315_
	);
	LUT4 #(
		.INIT('h3222)
	) name2387 (
		\data_o[31]_pad ,
		_w931_,
		_w934_,
		_w2784_,
		_w3316_
	);
	LUT4 #(
		.INIT('h7b00)
	) name2388 (
		\ks1_key_reg_reg[31]/NET0131 ,
		_w2785_,
		_w3314_,
		_w3316_,
		_w3317_
	);
	LUT2 #(
		.INIT('he)
	) name2389 (
		_w3315_,
		_w3317_,
		_w3318_
	);
	LUT4 #(
		.INIT('h5547)
	) name2390 (
		\data_i[88]_pad ,
		decrypt_i_pad,
		\mix1_data_o_reg_reg[88]/NET0131 ,
		_w930_,
		_w3319_
	);
	LUT4 #(
		.INIT('ha8ab)
	) name2391 (
		\sub1_data_reg_reg[88]/NET0131 ,
		_w996_,
		_w2776_,
		_w3319_,
		_w3320_
	);
	LUT4 #(
		.INIT('h404c)
	) name2392 (
		\mix1_data_o_reg_reg[88]/NET0131 ,
		_w2774_,
		_w2775_,
		_w3320_,
		_w3321_
	);
	LUT4 #(
		.INIT('h0545)
	) name2393 (
		\sub1_data_reg_reg[88]/NET0131 ,
		\sub1_ready_o_reg/NET0131 ,
		_w1054_,
		_w2230_,
		_w3322_
	);
	LUT4 #(
		.INIT('h1510)
	) name2394 (
		\state_reg/NET0131 ,
		\sub1_data_reg_reg[88]/NET0131 ,
		_w996_,
		_w3319_,
		_w3323_
	);
	LUT4 #(
		.INIT('h0057)
	) name2395 (
		\state_reg/NET0131 ,
		_w3321_,
		_w3322_,
		_w3323_,
		_w3324_
	);
	LUT3 #(
		.INIT('h48)
	) name2396 (
		\key_i[88]_pad ,
		_w931_,
		_w3324_,
		_w3325_
	);
	LUT4 #(
		.INIT('h3222)
	) name2397 (
		\data_o[88]_pad ,
		_w931_,
		_w934_,
		_w2784_,
		_w3326_
	);
	LUT4 #(
		.INIT('h7b00)
	) name2398 (
		\ks1_key_reg_reg[88]/NET0131 ,
		_w2785_,
		_w3324_,
		_w3326_,
		_w3327_
	);
	LUT2 #(
		.INIT('he)
	) name2399 (
		_w3325_,
		_w3327_,
		_w3328_
	);
	LUT4 #(
		.INIT('haab8)
	) name2400 (
		\data_i[119]_pad ,
		decrypt_i_pad,
		\mix1_data_o_reg_reg[119]/NET0131 ,
		_w930_,
		_w3329_
	);
	LUT4 #(
		.INIT('haba8)
	) name2401 (
		\sub1_data_reg_reg[119]/NET0131 ,
		_w996_,
		_w2776_,
		_w3329_,
		_w3330_
	);
	LUT4 #(
		.INIT('h404c)
	) name2402 (
		\mix1_data_o_reg_reg[119]/NET0131 ,
		_w2774_,
		_w2775_,
		_w3330_,
		_w3331_
	);
	LUT4 #(
		.INIT('h0545)
	) name2403 (
		\sub1_data_reg_reg[119]/NET0131 ,
		\sub1_ready_o_reg/NET0131 ,
		_w1054_,
		_w2230_,
		_w3332_
	);
	LUT4 #(
		.INIT('h1015)
	) name2404 (
		\state_reg/NET0131 ,
		\sub1_data_reg_reg[119]/NET0131 ,
		_w996_,
		_w3329_,
		_w3333_
	);
	LUT4 #(
		.INIT('h0057)
	) name2405 (
		\state_reg/NET0131 ,
		_w3331_,
		_w3332_,
		_w3333_,
		_w3334_
	);
	LUT3 #(
		.INIT('h48)
	) name2406 (
		\key_i[119]_pad ,
		_w931_,
		_w3334_,
		_w3335_
	);
	LUT4 #(
		.INIT('h3222)
	) name2407 (
		\data_o[119]_pad ,
		_w931_,
		_w934_,
		_w2784_,
		_w3336_
	);
	LUT4 #(
		.INIT('h7b00)
	) name2408 (
		\ks1_key_reg_reg[119]/NET0131 ,
		_w2785_,
		_w3334_,
		_w3336_,
		_w3337_
	);
	LUT2 #(
		.INIT('he)
	) name2409 (
		_w3335_,
		_w3337_,
		_w3338_
	);
	LUT4 #(
		.INIT('h5547)
	) name2410 (
		\data_i[89]_pad ,
		decrypt_i_pad,
		\mix1_data_o_reg_reg[89]/NET0131 ,
		_w930_,
		_w3339_
	);
	LUT4 #(
		.INIT('ha8ab)
	) name2411 (
		\sub1_data_reg_reg[89]/NET0131 ,
		_w996_,
		_w2776_,
		_w3339_,
		_w3340_
	);
	LUT4 #(
		.INIT('h404c)
	) name2412 (
		\mix1_data_o_reg_reg[89]/NET0131 ,
		_w2774_,
		_w2775_,
		_w3340_,
		_w3341_
	);
	LUT4 #(
		.INIT('h0545)
	) name2413 (
		\sub1_data_reg_reg[89]/NET0131 ,
		\sub1_ready_o_reg/NET0131 ,
		_w1054_,
		_w2230_,
		_w3342_
	);
	LUT4 #(
		.INIT('h1510)
	) name2414 (
		\state_reg/NET0131 ,
		\sub1_data_reg_reg[89]/NET0131 ,
		_w996_,
		_w3339_,
		_w3343_
	);
	LUT4 #(
		.INIT('h0057)
	) name2415 (
		\state_reg/NET0131 ,
		_w3341_,
		_w3342_,
		_w3343_,
		_w3344_
	);
	LUT3 #(
		.INIT('h48)
	) name2416 (
		\key_i[89]_pad ,
		_w931_,
		_w3344_,
		_w3345_
	);
	LUT4 #(
		.INIT('h3222)
	) name2417 (
		\data_o[89]_pad ,
		_w931_,
		_w934_,
		_w2784_,
		_w3346_
	);
	LUT4 #(
		.INIT('h7b00)
	) name2418 (
		\ks1_key_reg_reg[89]/NET0131 ,
		_w2785_,
		_w3344_,
		_w3346_,
		_w3347_
	);
	LUT2 #(
		.INIT('he)
	) name2419 (
		_w3345_,
		_w3347_,
		_w3348_
	);
	LUT4 #(
		.INIT('h5547)
	) name2420 (
		\data_i[8]_pad ,
		decrypt_i_pad,
		\mix1_data_o_reg_reg[8]/NET0131 ,
		_w930_,
		_w3349_
	);
	LUT4 #(
		.INIT('ha8ab)
	) name2421 (
		\sub1_data_reg_reg[8]/NET0131 ,
		_w996_,
		_w2776_,
		_w3349_,
		_w3350_
	);
	LUT4 #(
		.INIT('h404c)
	) name2422 (
		\mix1_data_o_reg_reg[8]/NET0131 ,
		_w2774_,
		_w2775_,
		_w3350_,
		_w3351_
	);
	LUT4 #(
		.INIT('h0545)
	) name2423 (
		\sub1_data_reg_reg[8]/NET0131 ,
		\sub1_ready_o_reg/NET0131 ,
		_w1054_,
		_w2230_,
		_w3352_
	);
	LUT4 #(
		.INIT('h1510)
	) name2424 (
		\state_reg/NET0131 ,
		\sub1_data_reg_reg[8]/NET0131 ,
		_w996_,
		_w3349_,
		_w3353_
	);
	LUT4 #(
		.INIT('h0057)
	) name2425 (
		\state_reg/NET0131 ,
		_w3351_,
		_w3352_,
		_w3353_,
		_w3354_
	);
	LUT3 #(
		.INIT('h48)
	) name2426 (
		\key_i[8]_pad ,
		_w931_,
		_w3354_,
		_w3355_
	);
	LUT4 #(
		.INIT('h3222)
	) name2427 (
		\data_o[8]_pad ,
		_w931_,
		_w934_,
		_w2784_,
		_w3356_
	);
	LUT4 #(
		.INIT('h7b00)
	) name2428 (
		\ks1_key_reg_reg[8]/NET0131 ,
		_w2785_,
		_w3354_,
		_w3356_,
		_w3357_
	);
	LUT2 #(
		.INIT('he)
	) name2429 (
		_w3355_,
		_w3357_,
		_w3358_
	);
	LUT4 #(
		.INIT('haab8)
	) name2430 (
		\data_i[32]_pad ,
		decrypt_i_pad,
		\mix1_data_o_reg_reg[32]/NET0131 ,
		_w930_,
		_w3359_
	);
	LUT4 #(
		.INIT('haba8)
	) name2431 (
		\sub1_data_reg_reg[32]/NET0131 ,
		_w996_,
		_w2776_,
		_w3359_,
		_w3360_
	);
	LUT4 #(
		.INIT('h404c)
	) name2432 (
		\mix1_data_o_reg_reg[32]/NET0131 ,
		_w2774_,
		_w2775_,
		_w3360_,
		_w3361_
	);
	LUT4 #(
		.INIT('h0545)
	) name2433 (
		\sub1_data_reg_reg[32]/NET0131 ,
		\sub1_ready_o_reg/NET0131 ,
		_w1054_,
		_w2230_,
		_w3362_
	);
	LUT4 #(
		.INIT('h1015)
	) name2434 (
		\state_reg/NET0131 ,
		\sub1_data_reg_reg[32]/NET0131 ,
		_w996_,
		_w3359_,
		_w3363_
	);
	LUT4 #(
		.INIT('h0057)
	) name2435 (
		\state_reg/NET0131 ,
		_w3361_,
		_w3362_,
		_w3363_,
		_w3364_
	);
	LUT3 #(
		.INIT('h48)
	) name2436 (
		\key_i[32]_pad ,
		_w931_,
		_w3364_,
		_w3365_
	);
	LUT4 #(
		.INIT('h3222)
	) name2437 (
		\data_o[32]_pad ,
		_w931_,
		_w934_,
		_w2784_,
		_w3366_
	);
	LUT4 #(
		.INIT('h7b00)
	) name2438 (
		\ks1_key_reg_reg[32]/NET0131 ,
		_w2785_,
		_w3364_,
		_w3366_,
		_w3367_
	);
	LUT2 #(
		.INIT('he)
	) name2439 (
		_w3365_,
		_w3367_,
		_w3368_
	);
	LUT4 #(
		.INIT('h5547)
	) name2440 (
		\data_i[104]_pad ,
		decrypt_i_pad,
		\mix1_data_o_reg_reg[104]/NET0131 ,
		_w930_,
		_w3369_
	);
	LUT4 #(
		.INIT('ha8ab)
	) name2441 (
		\sub1_data_reg_reg[104]/NET0131 ,
		_w996_,
		_w2776_,
		_w3369_,
		_w3370_
	);
	LUT4 #(
		.INIT('h404c)
	) name2442 (
		\mix1_data_o_reg_reg[104]/NET0131 ,
		_w2774_,
		_w2775_,
		_w3370_,
		_w3371_
	);
	LUT4 #(
		.INIT('h0545)
	) name2443 (
		\sub1_data_reg_reg[104]/NET0131 ,
		\sub1_ready_o_reg/NET0131 ,
		_w1054_,
		_w2230_,
		_w3372_
	);
	LUT4 #(
		.INIT('h1510)
	) name2444 (
		\state_reg/NET0131 ,
		\sub1_data_reg_reg[104]/NET0131 ,
		_w996_,
		_w3369_,
		_w3373_
	);
	LUT4 #(
		.INIT('h0057)
	) name2445 (
		\state_reg/NET0131 ,
		_w3371_,
		_w3372_,
		_w3373_,
		_w3374_
	);
	LUT3 #(
		.INIT('h48)
	) name2446 (
		\key_i[104]_pad ,
		_w931_,
		_w3374_,
		_w3375_
	);
	LUT4 #(
		.INIT('h3222)
	) name2447 (
		\data_o[104]_pad ,
		_w931_,
		_w934_,
		_w2784_,
		_w3376_
	);
	LUT4 #(
		.INIT('h7b00)
	) name2448 (
		\ks1_key_reg_reg[104]/NET0131 ,
		_w2785_,
		_w3374_,
		_w3376_,
		_w3377_
	);
	LUT2 #(
		.INIT('he)
	) name2449 (
		_w3375_,
		_w3377_,
		_w3378_
	);
	LUT4 #(
		.INIT('h5547)
	) name2450 (
		\data_i[90]_pad ,
		decrypt_i_pad,
		\mix1_data_o_reg_reg[90]/NET0131 ,
		_w930_,
		_w3379_
	);
	LUT4 #(
		.INIT('ha8ab)
	) name2451 (
		\sub1_data_reg_reg[90]/NET0131 ,
		_w996_,
		_w2776_,
		_w3379_,
		_w3380_
	);
	LUT4 #(
		.INIT('h404c)
	) name2452 (
		\mix1_data_o_reg_reg[90]/NET0131 ,
		_w2774_,
		_w2775_,
		_w3380_,
		_w3381_
	);
	LUT4 #(
		.INIT('h0545)
	) name2453 (
		\sub1_data_reg_reg[90]/NET0131 ,
		\sub1_ready_o_reg/NET0131 ,
		_w1054_,
		_w2230_,
		_w3382_
	);
	LUT4 #(
		.INIT('h1510)
	) name2454 (
		\state_reg/NET0131 ,
		\sub1_data_reg_reg[90]/NET0131 ,
		_w996_,
		_w3379_,
		_w3383_
	);
	LUT4 #(
		.INIT('h0057)
	) name2455 (
		\state_reg/NET0131 ,
		_w3381_,
		_w3382_,
		_w3383_,
		_w3384_
	);
	LUT3 #(
		.INIT('h48)
	) name2456 (
		\key_i[90]_pad ,
		_w931_,
		_w3384_,
		_w3385_
	);
	LUT4 #(
		.INIT('h3222)
	) name2457 (
		\data_o[90]_pad ,
		_w931_,
		_w934_,
		_w2784_,
		_w3386_
	);
	LUT4 #(
		.INIT('h7b00)
	) name2458 (
		\ks1_key_reg_reg[90]/NET0131 ,
		_w2785_,
		_w3384_,
		_w3386_,
		_w3387_
	);
	LUT2 #(
		.INIT('he)
	) name2459 (
		_w3385_,
		_w3387_,
		_w3388_
	);
	LUT4 #(
		.INIT('h5547)
	) name2460 (
		\data_i[105]_pad ,
		decrypt_i_pad,
		\mix1_data_o_reg_reg[105]/NET0131 ,
		_w930_,
		_w3389_
	);
	LUT4 #(
		.INIT('ha8ab)
	) name2461 (
		\sub1_data_reg_reg[105]/NET0131 ,
		_w996_,
		_w2776_,
		_w3389_,
		_w3390_
	);
	LUT4 #(
		.INIT('h404c)
	) name2462 (
		\mix1_data_o_reg_reg[105]/NET0131 ,
		_w2774_,
		_w2775_,
		_w3390_,
		_w3391_
	);
	LUT4 #(
		.INIT('h0545)
	) name2463 (
		\sub1_data_reg_reg[105]/NET0131 ,
		\sub1_ready_o_reg/NET0131 ,
		_w1054_,
		_w2230_,
		_w3392_
	);
	LUT4 #(
		.INIT('h1510)
	) name2464 (
		\state_reg/NET0131 ,
		\sub1_data_reg_reg[105]/NET0131 ,
		_w996_,
		_w3389_,
		_w3393_
	);
	LUT4 #(
		.INIT('h0057)
	) name2465 (
		\state_reg/NET0131 ,
		_w3391_,
		_w3392_,
		_w3393_,
		_w3394_
	);
	LUT3 #(
		.INIT('h48)
	) name2466 (
		\key_i[105]_pad ,
		_w931_,
		_w3394_,
		_w3395_
	);
	LUT4 #(
		.INIT('h3222)
	) name2467 (
		\data_o[105]_pad ,
		_w931_,
		_w934_,
		_w2784_,
		_w3396_
	);
	LUT4 #(
		.INIT('h7b00)
	) name2468 (
		\ks1_key_reg_reg[105]/NET0131 ,
		_w2785_,
		_w3394_,
		_w3396_,
		_w3397_
	);
	LUT2 #(
		.INIT('he)
	) name2469 (
		_w3395_,
		_w3397_,
		_w3398_
	);
	LUT4 #(
		.INIT('h5547)
	) name2470 (
		\data_i[91]_pad ,
		decrypt_i_pad,
		\mix1_data_o_reg_reg[91]/NET0131 ,
		_w930_,
		_w3399_
	);
	LUT4 #(
		.INIT('ha8ab)
	) name2471 (
		\sub1_data_reg_reg[91]/NET0131 ,
		_w996_,
		_w2776_,
		_w3399_,
		_w3400_
	);
	LUT4 #(
		.INIT('h404c)
	) name2472 (
		\mix1_data_o_reg_reg[91]/NET0131 ,
		_w2774_,
		_w2775_,
		_w3400_,
		_w3401_
	);
	LUT4 #(
		.INIT('h0545)
	) name2473 (
		\sub1_data_reg_reg[91]/NET0131 ,
		\sub1_ready_o_reg/NET0131 ,
		_w1054_,
		_w2230_,
		_w3402_
	);
	LUT4 #(
		.INIT('h1510)
	) name2474 (
		\state_reg/NET0131 ,
		\sub1_data_reg_reg[91]/NET0131 ,
		_w996_,
		_w3399_,
		_w3403_
	);
	LUT4 #(
		.INIT('h0057)
	) name2475 (
		\state_reg/NET0131 ,
		_w3401_,
		_w3402_,
		_w3403_,
		_w3404_
	);
	LUT3 #(
		.INIT('h48)
	) name2476 (
		\key_i[91]_pad ,
		_w931_,
		_w3404_,
		_w3405_
	);
	LUT4 #(
		.INIT('h3222)
	) name2477 (
		\data_o[91]_pad ,
		_w931_,
		_w934_,
		_w2784_,
		_w3406_
	);
	LUT4 #(
		.INIT('h7b00)
	) name2478 (
		\ks1_key_reg_reg[91]/NET0131 ,
		_w2785_,
		_w3404_,
		_w3406_,
		_w3407_
	);
	LUT2 #(
		.INIT('he)
	) name2479 (
		_w3405_,
		_w3407_,
		_w3408_
	);
	LUT4 #(
		.INIT('haab8)
	) name2480 (
		\data_i[33]_pad ,
		decrypt_i_pad,
		\mix1_data_o_reg_reg[33]/NET0131 ,
		_w930_,
		_w3409_
	);
	LUT4 #(
		.INIT('haba8)
	) name2481 (
		\sub1_data_reg_reg[33]/NET0131 ,
		_w996_,
		_w2776_,
		_w3409_,
		_w3410_
	);
	LUT4 #(
		.INIT('h404c)
	) name2482 (
		\mix1_data_o_reg_reg[33]/NET0131 ,
		_w2774_,
		_w2775_,
		_w3410_,
		_w3411_
	);
	LUT4 #(
		.INIT('h0545)
	) name2483 (
		\sub1_data_reg_reg[33]/NET0131 ,
		\sub1_ready_o_reg/NET0131 ,
		_w1054_,
		_w2230_,
		_w3412_
	);
	LUT4 #(
		.INIT('h1015)
	) name2484 (
		\state_reg/NET0131 ,
		\sub1_data_reg_reg[33]/NET0131 ,
		_w996_,
		_w3409_,
		_w3413_
	);
	LUT4 #(
		.INIT('h0057)
	) name2485 (
		\state_reg/NET0131 ,
		_w3411_,
		_w3412_,
		_w3413_,
		_w3414_
	);
	LUT3 #(
		.INIT('h48)
	) name2486 (
		\key_i[33]_pad ,
		_w931_,
		_w3414_,
		_w3415_
	);
	LUT4 #(
		.INIT('h3222)
	) name2487 (
		\data_o[33]_pad ,
		_w931_,
		_w934_,
		_w2784_,
		_w3416_
	);
	LUT4 #(
		.INIT('h7b00)
	) name2488 (
		\ks1_key_reg_reg[33]/NET0131 ,
		_w2785_,
		_w3414_,
		_w3416_,
		_w3417_
	);
	LUT2 #(
		.INIT('he)
	) name2489 (
		_w3415_,
		_w3417_,
		_w3418_
	);
	LUT4 #(
		.INIT('h5547)
	) name2490 (
		\data_i[11]_pad ,
		decrypt_i_pad,
		\mix1_data_o_reg_reg[11]/NET0131 ,
		_w930_,
		_w3419_
	);
	LUT4 #(
		.INIT('ha8ab)
	) name2491 (
		\sub1_data_reg_reg[11]/NET0131 ,
		_w996_,
		_w2776_,
		_w3419_,
		_w3420_
	);
	LUT4 #(
		.INIT('h404c)
	) name2492 (
		\mix1_data_o_reg_reg[11]/NET0131 ,
		_w2774_,
		_w2775_,
		_w3420_,
		_w3421_
	);
	LUT4 #(
		.INIT('h0545)
	) name2493 (
		\sub1_data_reg_reg[11]/NET0131 ,
		\sub1_ready_o_reg/NET0131 ,
		_w1054_,
		_w2230_,
		_w3422_
	);
	LUT4 #(
		.INIT('h1510)
	) name2494 (
		\state_reg/NET0131 ,
		\sub1_data_reg_reg[11]/NET0131 ,
		_w996_,
		_w3419_,
		_w3423_
	);
	LUT4 #(
		.INIT('h0057)
	) name2495 (
		\state_reg/NET0131 ,
		_w3421_,
		_w3422_,
		_w3423_,
		_w3424_
	);
	LUT3 #(
		.INIT('h48)
	) name2496 (
		\key_i[11]_pad ,
		_w931_,
		_w3424_,
		_w3425_
	);
	LUT4 #(
		.INIT('h3222)
	) name2497 (
		\data_o[11]_pad ,
		_w931_,
		_w934_,
		_w2784_,
		_w3426_
	);
	LUT4 #(
		.INIT('h7b00)
	) name2498 (
		\ks1_key_reg_reg[11]/NET0131 ,
		_w2785_,
		_w3424_,
		_w3426_,
		_w3427_
	);
	LUT2 #(
		.INIT('he)
	) name2499 (
		_w3425_,
		_w3427_,
		_w3428_
	);
	LUT4 #(
		.INIT('h5547)
	) name2500 (
		\data_i[92]_pad ,
		decrypt_i_pad,
		\mix1_data_o_reg_reg[92]/NET0131 ,
		_w930_,
		_w3429_
	);
	LUT4 #(
		.INIT('ha8ab)
	) name2501 (
		\sub1_data_reg_reg[92]/NET0131 ,
		_w996_,
		_w2776_,
		_w3429_,
		_w3430_
	);
	LUT4 #(
		.INIT('h404c)
	) name2502 (
		\mix1_data_o_reg_reg[92]/NET0131 ,
		_w2774_,
		_w2775_,
		_w3430_,
		_w3431_
	);
	LUT4 #(
		.INIT('h0545)
	) name2503 (
		\sub1_data_reg_reg[92]/NET0131 ,
		\sub1_ready_o_reg/NET0131 ,
		_w1054_,
		_w2230_,
		_w3432_
	);
	LUT4 #(
		.INIT('h1510)
	) name2504 (
		\state_reg/NET0131 ,
		\sub1_data_reg_reg[92]/NET0131 ,
		_w996_,
		_w3429_,
		_w3433_
	);
	LUT4 #(
		.INIT('h0057)
	) name2505 (
		\state_reg/NET0131 ,
		_w3431_,
		_w3432_,
		_w3433_,
		_w3434_
	);
	LUT3 #(
		.INIT('h48)
	) name2506 (
		\key_i[92]_pad ,
		_w931_,
		_w3434_,
		_w3435_
	);
	LUT4 #(
		.INIT('h3222)
	) name2507 (
		\data_o[92]_pad ,
		_w931_,
		_w934_,
		_w2784_,
		_w3436_
	);
	LUT4 #(
		.INIT('h7b00)
	) name2508 (
		\ks1_key_reg_reg[92]/NET0131 ,
		_w2785_,
		_w3434_,
		_w3436_,
		_w3437_
	);
	LUT2 #(
		.INIT('he)
	) name2509 (
		_w3435_,
		_w3437_,
		_w3438_
	);
	LUT4 #(
		.INIT('h5547)
	) name2510 (
		\data_i[93]_pad ,
		decrypt_i_pad,
		\mix1_data_o_reg_reg[93]/NET0131 ,
		_w930_,
		_w3439_
	);
	LUT4 #(
		.INIT('ha8ab)
	) name2511 (
		\sub1_data_reg_reg[93]/NET0131 ,
		_w996_,
		_w2776_,
		_w3439_,
		_w3440_
	);
	LUT4 #(
		.INIT('h404c)
	) name2512 (
		\mix1_data_o_reg_reg[93]/NET0131 ,
		_w2774_,
		_w2775_,
		_w3440_,
		_w3441_
	);
	LUT4 #(
		.INIT('h0545)
	) name2513 (
		\sub1_data_reg_reg[93]/NET0131 ,
		\sub1_ready_o_reg/NET0131 ,
		_w1054_,
		_w2230_,
		_w3442_
	);
	LUT4 #(
		.INIT('h1510)
	) name2514 (
		\state_reg/NET0131 ,
		\sub1_data_reg_reg[93]/NET0131 ,
		_w996_,
		_w3439_,
		_w3443_
	);
	LUT4 #(
		.INIT('h0057)
	) name2515 (
		\state_reg/NET0131 ,
		_w3441_,
		_w3442_,
		_w3443_,
		_w3444_
	);
	LUT3 #(
		.INIT('h48)
	) name2516 (
		\key_i[93]_pad ,
		_w931_,
		_w3444_,
		_w3445_
	);
	LUT4 #(
		.INIT('h3222)
	) name2517 (
		\data_o[93]_pad ,
		_w931_,
		_w934_,
		_w2784_,
		_w3446_
	);
	LUT4 #(
		.INIT('h7b00)
	) name2518 (
		\ks1_key_reg_reg[93]/NET0131 ,
		_w2785_,
		_w3444_,
		_w3446_,
		_w3447_
	);
	LUT2 #(
		.INIT('he)
	) name2519 (
		_w3445_,
		_w3447_,
		_w3448_
	);
	LUT4 #(
		.INIT('haab8)
	) name2520 (
		\data_i[34]_pad ,
		decrypt_i_pad,
		\mix1_data_o_reg_reg[34]/NET0131 ,
		_w930_,
		_w3449_
	);
	LUT4 #(
		.INIT('haba8)
	) name2521 (
		\sub1_data_reg_reg[34]/NET0131 ,
		_w996_,
		_w2776_,
		_w3449_,
		_w3450_
	);
	LUT4 #(
		.INIT('h404c)
	) name2522 (
		\mix1_data_o_reg_reg[34]/NET0131 ,
		_w2774_,
		_w2775_,
		_w3450_,
		_w3451_
	);
	LUT4 #(
		.INIT('h0545)
	) name2523 (
		\sub1_data_reg_reg[34]/NET0131 ,
		\sub1_ready_o_reg/NET0131 ,
		_w1054_,
		_w2230_,
		_w3452_
	);
	LUT4 #(
		.INIT('h1015)
	) name2524 (
		\state_reg/NET0131 ,
		\sub1_data_reg_reg[34]/NET0131 ,
		_w996_,
		_w3449_,
		_w3453_
	);
	LUT4 #(
		.INIT('h0057)
	) name2525 (
		\state_reg/NET0131 ,
		_w3451_,
		_w3452_,
		_w3453_,
		_w3454_
	);
	LUT3 #(
		.INIT('h48)
	) name2526 (
		\key_i[34]_pad ,
		_w931_,
		_w3454_,
		_w3455_
	);
	LUT4 #(
		.INIT('h3222)
	) name2527 (
		\data_o[34]_pad ,
		_w931_,
		_w934_,
		_w2784_,
		_w3456_
	);
	LUT4 #(
		.INIT('h7b00)
	) name2528 (
		\ks1_key_reg_reg[34]/NET0131 ,
		_w2785_,
		_w3454_,
		_w3456_,
		_w3457_
	);
	LUT2 #(
		.INIT('he)
	) name2529 (
		_w3455_,
		_w3457_,
		_w3458_
	);
	LUT4 #(
		.INIT('h5547)
	) name2530 (
		\data_i[94]_pad ,
		decrypt_i_pad,
		\mix1_data_o_reg_reg[94]/NET0131 ,
		_w930_,
		_w3459_
	);
	LUT4 #(
		.INIT('ha8ab)
	) name2531 (
		\sub1_data_reg_reg[94]/NET0131 ,
		_w996_,
		_w2776_,
		_w3459_,
		_w3460_
	);
	LUT4 #(
		.INIT('h404c)
	) name2532 (
		\mix1_data_o_reg_reg[94]/NET0131 ,
		_w2774_,
		_w2775_,
		_w3460_,
		_w3461_
	);
	LUT4 #(
		.INIT('h0545)
	) name2533 (
		\sub1_data_reg_reg[94]/NET0131 ,
		\sub1_ready_o_reg/NET0131 ,
		_w1054_,
		_w2230_,
		_w3462_
	);
	LUT4 #(
		.INIT('h1510)
	) name2534 (
		\state_reg/NET0131 ,
		\sub1_data_reg_reg[94]/NET0131 ,
		_w996_,
		_w3459_,
		_w3463_
	);
	LUT4 #(
		.INIT('h0057)
	) name2535 (
		\state_reg/NET0131 ,
		_w3461_,
		_w3462_,
		_w3463_,
		_w3464_
	);
	LUT3 #(
		.INIT('h48)
	) name2536 (
		\key_i[94]_pad ,
		_w931_,
		_w3464_,
		_w3465_
	);
	LUT4 #(
		.INIT('h3222)
	) name2537 (
		\data_o[94]_pad ,
		_w931_,
		_w934_,
		_w2784_,
		_w3466_
	);
	LUT4 #(
		.INIT('h7b00)
	) name2538 (
		\ks1_key_reg_reg[94]/NET0131 ,
		_w2785_,
		_w3464_,
		_w3466_,
		_w3467_
	);
	LUT2 #(
		.INIT('he)
	) name2539 (
		_w3465_,
		_w3467_,
		_w3468_
	);
	LUT4 #(
		.INIT('h5547)
	) name2540 (
		\data_i[95]_pad ,
		decrypt_i_pad,
		\mix1_data_o_reg_reg[95]/NET0131 ,
		_w930_,
		_w3469_
	);
	LUT4 #(
		.INIT('ha8ab)
	) name2541 (
		\sub1_data_reg_reg[95]/NET0131 ,
		_w996_,
		_w2776_,
		_w3469_,
		_w3470_
	);
	LUT4 #(
		.INIT('h404c)
	) name2542 (
		\mix1_data_o_reg_reg[95]/NET0131 ,
		_w2774_,
		_w2775_,
		_w3470_,
		_w3471_
	);
	LUT4 #(
		.INIT('h0545)
	) name2543 (
		\sub1_data_reg_reg[95]/NET0131 ,
		\sub1_ready_o_reg/NET0131 ,
		_w1054_,
		_w2230_,
		_w3472_
	);
	LUT4 #(
		.INIT('h1510)
	) name2544 (
		\state_reg/NET0131 ,
		\sub1_data_reg_reg[95]/NET0131 ,
		_w996_,
		_w3469_,
		_w3473_
	);
	LUT4 #(
		.INIT('h0057)
	) name2545 (
		\state_reg/NET0131 ,
		_w3471_,
		_w3472_,
		_w3473_,
		_w3474_
	);
	LUT3 #(
		.INIT('h48)
	) name2546 (
		\key_i[95]_pad ,
		_w931_,
		_w3474_,
		_w3475_
	);
	LUT4 #(
		.INIT('h3222)
	) name2547 (
		\data_o[95]_pad ,
		_w931_,
		_w934_,
		_w2784_,
		_w3476_
	);
	LUT4 #(
		.INIT('h7b00)
	) name2548 (
		\ks1_key_reg_reg[95]/NET0131 ,
		_w2785_,
		_w3474_,
		_w3476_,
		_w3477_
	);
	LUT2 #(
		.INIT('he)
	) name2549 (
		_w3475_,
		_w3477_,
		_w3478_
	);
	LUT4 #(
		.INIT('haab8)
	) name2550 (
		\data_i[35]_pad ,
		decrypt_i_pad,
		\mix1_data_o_reg_reg[35]/NET0131 ,
		_w930_,
		_w3479_
	);
	LUT4 #(
		.INIT('haba8)
	) name2551 (
		\sub1_data_reg_reg[35]/NET0131 ,
		_w996_,
		_w2776_,
		_w3479_,
		_w3480_
	);
	LUT4 #(
		.INIT('h404c)
	) name2552 (
		\mix1_data_o_reg_reg[35]/NET0131 ,
		_w2774_,
		_w2775_,
		_w3480_,
		_w3481_
	);
	LUT4 #(
		.INIT('h0545)
	) name2553 (
		\sub1_data_reg_reg[35]/NET0131 ,
		\sub1_ready_o_reg/NET0131 ,
		_w1054_,
		_w2230_,
		_w3482_
	);
	LUT4 #(
		.INIT('h1015)
	) name2554 (
		\state_reg/NET0131 ,
		\sub1_data_reg_reg[35]/NET0131 ,
		_w996_,
		_w3479_,
		_w3483_
	);
	LUT4 #(
		.INIT('h0057)
	) name2555 (
		\state_reg/NET0131 ,
		_w3481_,
		_w3482_,
		_w3483_,
		_w3484_
	);
	LUT3 #(
		.INIT('h48)
	) name2556 (
		\key_i[35]_pad ,
		_w931_,
		_w3484_,
		_w3485_
	);
	LUT4 #(
		.INIT('h3222)
	) name2557 (
		\data_o[35]_pad ,
		_w931_,
		_w934_,
		_w2784_,
		_w3486_
	);
	LUT4 #(
		.INIT('h7b00)
	) name2558 (
		\ks1_key_reg_reg[35]/NET0131 ,
		_w2785_,
		_w3484_,
		_w3486_,
		_w3487_
	);
	LUT2 #(
		.INIT('he)
	) name2559 (
		_w3485_,
		_w3487_,
		_w3488_
	);
	LUT4 #(
		.INIT('ha820)
	) name2560 (
		\data_i[96]_pad ,
		decrypt_i_pad,
		_w930_,
		_w995_,
		_w3489_
	);
	LUT3 #(
		.INIT('h04)
	) name2561 (
		decrypt_i_pad,
		\mix1_data_o_reg_reg[96]/NET0131 ,
		_w930_,
		_w3490_
	);
	LUT3 #(
		.INIT('h08)
	) name2562 (
		decrypt_i_pad,
		\sub1_data_reg_reg[96]/NET0131 ,
		_w995_,
		_w3491_
	);
	LUT4 #(
		.INIT('h5554)
	) name2563 (
		_w2776_,
		_w3489_,
		_w3490_,
		_w3491_,
		_w3492_
	);
	LUT4 #(
		.INIT('h1bbb)
	) name2564 (
		decrypt_i_pad,
		\mix1_ready_o_reg/NET0131 ,
		\sub1_data_reg_reg[96]/NET0131 ,
		\sub1_ready_o_reg/NET0131 ,
		_w3493_
	);
	LUT3 #(
		.INIT('h10)
	) name2565 (
		decrypt_i_pad,
		\mix1_data_o_reg_reg[96]/NET0131 ,
		\mix1_ready_o_reg/NET0131 ,
		_w3494_
	);
	LUT4 #(
		.INIT('haa20)
	) name2566 (
		_w2774_,
		_w3492_,
		_w3493_,
		_w3494_,
		_w3495_
	);
	LUT4 #(
		.INIT('h0545)
	) name2567 (
		\sub1_data_reg_reg[96]/NET0131 ,
		\sub1_ready_o_reg/NET0131 ,
		_w1054_,
		_w2230_,
		_w3496_
	);
	LUT4 #(
		.INIT('h0001)
	) name2568 (
		\state_reg/NET0131 ,
		_w3489_,
		_w3490_,
		_w3491_,
		_w3497_
	);
	LUT4 #(
		.INIT('h0057)
	) name2569 (
		\state_reg/NET0131 ,
		_w3495_,
		_w3496_,
		_w3497_,
		_w3498_
	);
	LUT3 #(
		.INIT('h48)
	) name2570 (
		\key_i[96]_pad ,
		_w931_,
		_w3498_,
		_w3499_
	);
	LUT4 #(
		.INIT('h3222)
	) name2571 (
		\data_o[96]_pad ,
		_w931_,
		_w934_,
		_w2784_,
		_w3500_
	);
	LUT4 #(
		.INIT('h7b00)
	) name2572 (
		\ks1_key_reg_reg[96]/NET0131 ,
		_w2785_,
		_w3498_,
		_w3500_,
		_w3501_
	);
	LUT2 #(
		.INIT('he)
	) name2573 (
		_w3499_,
		_w3501_,
		_w3502_
	);
	LUT4 #(
		.INIT('h5547)
	) name2574 (
		\data_i[120]_pad ,
		decrypt_i_pad,
		\mix1_data_o_reg_reg[120]/NET0131 ,
		_w930_,
		_w3503_
	);
	LUT4 #(
		.INIT('ha8ab)
	) name2575 (
		\sub1_data_reg_reg[120]/NET0131 ,
		_w996_,
		_w2776_,
		_w3503_,
		_w3504_
	);
	LUT4 #(
		.INIT('h404c)
	) name2576 (
		\mix1_data_o_reg_reg[120]/NET0131 ,
		_w2774_,
		_w2775_,
		_w3504_,
		_w3505_
	);
	LUT4 #(
		.INIT('h0545)
	) name2577 (
		\sub1_data_reg_reg[120]/NET0131 ,
		\sub1_ready_o_reg/NET0131 ,
		_w1054_,
		_w2230_,
		_w3506_
	);
	LUT4 #(
		.INIT('h1510)
	) name2578 (
		\state_reg/NET0131 ,
		\sub1_data_reg_reg[120]/NET0131 ,
		_w996_,
		_w3503_,
		_w3507_
	);
	LUT4 #(
		.INIT('h0057)
	) name2579 (
		\state_reg/NET0131 ,
		_w3505_,
		_w3506_,
		_w3507_,
		_w3508_
	);
	LUT3 #(
		.INIT('h48)
	) name2580 (
		\key_i[120]_pad ,
		_w931_,
		_w3508_,
		_w3509_
	);
	LUT4 #(
		.INIT('h3222)
	) name2581 (
		\data_o[120]_pad ,
		_w931_,
		_w934_,
		_w2784_,
		_w3510_
	);
	LUT4 #(
		.INIT('h7b00)
	) name2582 (
		\ks1_key_reg_reg[120]/NET0131 ,
		_w2785_,
		_w3508_,
		_w3510_,
		_w3511_
	);
	LUT2 #(
		.INIT('he)
	) name2583 (
		_w3509_,
		_w3511_,
		_w3512_
	);
	LUT4 #(
		.INIT('haab8)
	) name2584 (
		\data_i[36]_pad ,
		decrypt_i_pad,
		\mix1_data_o_reg_reg[36]/NET0131 ,
		_w930_,
		_w3513_
	);
	LUT4 #(
		.INIT('haba8)
	) name2585 (
		\sub1_data_reg_reg[36]/NET0131 ,
		_w996_,
		_w2776_,
		_w3513_,
		_w3514_
	);
	LUT4 #(
		.INIT('h404c)
	) name2586 (
		\mix1_data_o_reg_reg[36]/NET0131 ,
		_w2774_,
		_w2775_,
		_w3514_,
		_w3515_
	);
	LUT4 #(
		.INIT('h0545)
	) name2587 (
		\sub1_data_reg_reg[36]/NET0131 ,
		\sub1_ready_o_reg/NET0131 ,
		_w1054_,
		_w2230_,
		_w3516_
	);
	LUT4 #(
		.INIT('h1015)
	) name2588 (
		\state_reg/NET0131 ,
		\sub1_data_reg_reg[36]/NET0131 ,
		_w996_,
		_w3513_,
		_w3517_
	);
	LUT4 #(
		.INIT('h0057)
	) name2589 (
		\state_reg/NET0131 ,
		_w3515_,
		_w3516_,
		_w3517_,
		_w3518_
	);
	LUT3 #(
		.INIT('h48)
	) name2590 (
		\key_i[36]_pad ,
		_w931_,
		_w3518_,
		_w3519_
	);
	LUT4 #(
		.INIT('h3222)
	) name2591 (
		\data_o[36]_pad ,
		_w931_,
		_w934_,
		_w2784_,
		_w3520_
	);
	LUT4 #(
		.INIT('h7b00)
	) name2592 (
		\ks1_key_reg_reg[36]/NET0131 ,
		_w2785_,
		_w3518_,
		_w3520_,
		_w3521_
	);
	LUT2 #(
		.INIT('he)
	) name2593 (
		_w3519_,
		_w3521_,
		_w3522_
	);
	LUT4 #(
		.INIT('ha820)
	) name2594 (
		\data_i[97]_pad ,
		decrypt_i_pad,
		_w930_,
		_w995_,
		_w3523_
	);
	LUT3 #(
		.INIT('h04)
	) name2595 (
		decrypt_i_pad,
		\mix1_data_o_reg_reg[97]/NET0131 ,
		_w930_,
		_w3524_
	);
	LUT3 #(
		.INIT('h08)
	) name2596 (
		decrypt_i_pad,
		\sub1_data_reg_reg[97]/NET0131 ,
		_w995_,
		_w3525_
	);
	LUT4 #(
		.INIT('h5554)
	) name2597 (
		_w2776_,
		_w3523_,
		_w3524_,
		_w3525_,
		_w3526_
	);
	LUT4 #(
		.INIT('h1bbb)
	) name2598 (
		decrypt_i_pad,
		\mix1_ready_o_reg/NET0131 ,
		\sub1_data_reg_reg[97]/NET0131 ,
		\sub1_ready_o_reg/NET0131 ,
		_w3527_
	);
	LUT3 #(
		.INIT('h10)
	) name2599 (
		decrypt_i_pad,
		\mix1_data_o_reg_reg[97]/NET0131 ,
		\mix1_ready_o_reg/NET0131 ,
		_w3528_
	);
	LUT4 #(
		.INIT('haa20)
	) name2600 (
		_w2774_,
		_w3526_,
		_w3527_,
		_w3528_,
		_w3529_
	);
	LUT4 #(
		.INIT('h0545)
	) name2601 (
		\sub1_data_reg_reg[97]/NET0131 ,
		\sub1_ready_o_reg/NET0131 ,
		_w1054_,
		_w2230_,
		_w3530_
	);
	LUT4 #(
		.INIT('h0001)
	) name2602 (
		\state_reg/NET0131 ,
		_w3523_,
		_w3524_,
		_w3525_,
		_w3531_
	);
	LUT4 #(
		.INIT('h0057)
	) name2603 (
		\state_reg/NET0131 ,
		_w3529_,
		_w3530_,
		_w3531_,
		_w3532_
	);
	LUT3 #(
		.INIT('h48)
	) name2604 (
		\key_i[97]_pad ,
		_w931_,
		_w3532_,
		_w3533_
	);
	LUT4 #(
		.INIT('h3222)
	) name2605 (
		\data_o[97]_pad ,
		_w931_,
		_w934_,
		_w2784_,
		_w3534_
	);
	LUT4 #(
		.INIT('h7b00)
	) name2606 (
		\ks1_key_reg_reg[97]/NET0131 ,
		_w2785_,
		_w3532_,
		_w3534_,
		_w3535_
	);
	LUT2 #(
		.INIT('he)
	) name2607 (
		_w3533_,
		_w3535_,
		_w3536_
	);
	LUT4 #(
		.INIT('haab8)
	) name2608 (
		\data_i[98]_pad ,
		decrypt_i_pad,
		\mix1_data_o_reg_reg[98]/NET0131 ,
		_w930_,
		_w3537_
	);
	LUT4 #(
		.INIT('haba8)
	) name2609 (
		\sub1_data_reg_reg[98]/NET0131 ,
		_w996_,
		_w2776_,
		_w3537_,
		_w3538_
	);
	LUT4 #(
		.INIT('h404c)
	) name2610 (
		\mix1_data_o_reg_reg[98]/NET0131 ,
		_w2774_,
		_w2775_,
		_w3538_,
		_w3539_
	);
	LUT4 #(
		.INIT('h0545)
	) name2611 (
		\sub1_data_reg_reg[98]/NET0131 ,
		\sub1_ready_o_reg/NET0131 ,
		_w1054_,
		_w2230_,
		_w3540_
	);
	LUT4 #(
		.INIT('h1015)
	) name2612 (
		\state_reg/NET0131 ,
		\sub1_data_reg_reg[98]/NET0131 ,
		_w996_,
		_w3537_,
		_w3541_
	);
	LUT4 #(
		.INIT('h0057)
	) name2613 (
		\state_reg/NET0131 ,
		_w3539_,
		_w3540_,
		_w3541_,
		_w3542_
	);
	LUT3 #(
		.INIT('h48)
	) name2614 (
		\key_i[98]_pad ,
		_w931_,
		_w3542_,
		_w3543_
	);
	LUT4 #(
		.INIT('h3222)
	) name2615 (
		\data_o[98]_pad ,
		_w931_,
		_w934_,
		_w2784_,
		_w3544_
	);
	LUT4 #(
		.INIT('h7b00)
	) name2616 (
		\ks1_key_reg_reg[98]/NET0131 ,
		_w2785_,
		_w3542_,
		_w3544_,
		_w3545_
	);
	LUT2 #(
		.INIT('he)
	) name2617 (
		_w3543_,
		_w3545_,
		_w3546_
	);
	LUT4 #(
		.INIT('haab8)
	) name2618 (
		\data_i[37]_pad ,
		decrypt_i_pad,
		\mix1_data_o_reg_reg[37]/NET0131 ,
		_w930_,
		_w3547_
	);
	LUT4 #(
		.INIT('haba8)
	) name2619 (
		\sub1_data_reg_reg[37]/NET0131 ,
		_w996_,
		_w2776_,
		_w3547_,
		_w3548_
	);
	LUT4 #(
		.INIT('h404c)
	) name2620 (
		\mix1_data_o_reg_reg[37]/NET0131 ,
		_w2774_,
		_w2775_,
		_w3548_,
		_w3549_
	);
	LUT4 #(
		.INIT('h0545)
	) name2621 (
		\sub1_data_reg_reg[37]/NET0131 ,
		\sub1_ready_o_reg/NET0131 ,
		_w1054_,
		_w2230_,
		_w3550_
	);
	LUT4 #(
		.INIT('h1015)
	) name2622 (
		\state_reg/NET0131 ,
		\sub1_data_reg_reg[37]/NET0131 ,
		_w996_,
		_w3547_,
		_w3551_
	);
	LUT4 #(
		.INIT('h0057)
	) name2623 (
		\state_reg/NET0131 ,
		_w3549_,
		_w3550_,
		_w3551_,
		_w3552_
	);
	LUT3 #(
		.INIT('h48)
	) name2624 (
		\key_i[37]_pad ,
		_w931_,
		_w3552_,
		_w3553_
	);
	LUT4 #(
		.INIT('h3222)
	) name2625 (
		\data_o[37]_pad ,
		_w931_,
		_w934_,
		_w2784_,
		_w3554_
	);
	LUT4 #(
		.INIT('h7b00)
	) name2626 (
		\ks1_key_reg_reg[37]/NET0131 ,
		_w2785_,
		_w3552_,
		_w3554_,
		_w3555_
	);
	LUT2 #(
		.INIT('he)
	) name2627 (
		_w3553_,
		_w3555_,
		_w3556_
	);
	LUT4 #(
		.INIT('haab8)
	) name2628 (
		\data_i[99]_pad ,
		decrypt_i_pad,
		\mix1_data_o_reg_reg[99]/NET0131 ,
		_w930_,
		_w3557_
	);
	LUT4 #(
		.INIT('haba8)
	) name2629 (
		\sub1_data_reg_reg[99]/NET0131 ,
		_w996_,
		_w2776_,
		_w3557_,
		_w3558_
	);
	LUT4 #(
		.INIT('h404c)
	) name2630 (
		\mix1_data_o_reg_reg[99]/NET0131 ,
		_w2774_,
		_w2775_,
		_w3558_,
		_w3559_
	);
	LUT4 #(
		.INIT('h0545)
	) name2631 (
		\sub1_data_reg_reg[99]/NET0131 ,
		\sub1_ready_o_reg/NET0131 ,
		_w1054_,
		_w2230_,
		_w3560_
	);
	LUT4 #(
		.INIT('h1015)
	) name2632 (
		\state_reg/NET0131 ,
		\sub1_data_reg_reg[99]/NET0131 ,
		_w996_,
		_w3557_,
		_w3561_
	);
	LUT4 #(
		.INIT('h0057)
	) name2633 (
		\state_reg/NET0131 ,
		_w3559_,
		_w3560_,
		_w3561_,
		_w3562_
	);
	LUT3 #(
		.INIT('h48)
	) name2634 (
		\key_i[99]_pad ,
		_w931_,
		_w3562_,
		_w3563_
	);
	LUT4 #(
		.INIT('h3222)
	) name2635 (
		\data_o[99]_pad ,
		_w931_,
		_w934_,
		_w2784_,
		_w3564_
	);
	LUT4 #(
		.INIT('h7b00)
	) name2636 (
		\ks1_key_reg_reg[99]/NET0131 ,
		_w2785_,
		_w3562_,
		_w3564_,
		_w3565_
	);
	LUT2 #(
		.INIT('he)
	) name2637 (
		_w3563_,
		_w3565_,
		_w3566_
	);
	LUT4 #(
		.INIT('h5547)
	) name2638 (
		\data_i[121]_pad ,
		decrypt_i_pad,
		\mix1_data_o_reg_reg[121]/NET0131 ,
		_w930_,
		_w3567_
	);
	LUT4 #(
		.INIT('ha8ab)
	) name2639 (
		\sub1_data_reg_reg[121]/NET0131 ,
		_w996_,
		_w2776_,
		_w3567_,
		_w3568_
	);
	LUT4 #(
		.INIT('h404c)
	) name2640 (
		\mix1_data_o_reg_reg[121]/NET0131 ,
		_w2774_,
		_w2775_,
		_w3568_,
		_w3569_
	);
	LUT4 #(
		.INIT('h0545)
	) name2641 (
		\sub1_data_reg_reg[121]/NET0131 ,
		\sub1_ready_o_reg/NET0131 ,
		_w1054_,
		_w2230_,
		_w3570_
	);
	LUT4 #(
		.INIT('h1510)
	) name2642 (
		\state_reg/NET0131 ,
		\sub1_data_reg_reg[121]/NET0131 ,
		_w996_,
		_w3567_,
		_w3571_
	);
	LUT4 #(
		.INIT('h0057)
	) name2643 (
		\state_reg/NET0131 ,
		_w3569_,
		_w3570_,
		_w3571_,
		_w3572_
	);
	LUT3 #(
		.INIT('h48)
	) name2644 (
		\key_i[121]_pad ,
		_w931_,
		_w3572_,
		_w3573_
	);
	LUT4 #(
		.INIT('h3222)
	) name2645 (
		\data_o[121]_pad ,
		_w931_,
		_w934_,
		_w2784_,
		_w3574_
	);
	LUT4 #(
		.INIT('h7b00)
	) name2646 (
		\ks1_key_reg_reg[121]/NET0131 ,
		_w2785_,
		_w3572_,
		_w3574_,
		_w3575_
	);
	LUT2 #(
		.INIT('he)
	) name2647 (
		_w3573_,
		_w3575_,
		_w3576_
	);
	LUT4 #(
		.INIT('h5547)
	) name2648 (
		\data_i[9]_pad ,
		decrypt_i_pad,
		\mix1_data_o_reg_reg[9]/NET0131 ,
		_w930_,
		_w3577_
	);
	LUT4 #(
		.INIT('ha8ab)
	) name2649 (
		\sub1_data_reg_reg[9]/NET0131 ,
		_w996_,
		_w2776_,
		_w3577_,
		_w3578_
	);
	LUT4 #(
		.INIT('h404c)
	) name2650 (
		\mix1_data_o_reg_reg[9]/NET0131 ,
		_w2774_,
		_w2775_,
		_w3578_,
		_w3579_
	);
	LUT4 #(
		.INIT('h0545)
	) name2651 (
		\sub1_data_reg_reg[9]/NET0131 ,
		\sub1_ready_o_reg/NET0131 ,
		_w1054_,
		_w2230_,
		_w3580_
	);
	LUT4 #(
		.INIT('h1510)
	) name2652 (
		\state_reg/NET0131 ,
		\sub1_data_reg_reg[9]/NET0131 ,
		_w996_,
		_w3577_,
		_w3581_
	);
	LUT4 #(
		.INIT('h0057)
	) name2653 (
		\state_reg/NET0131 ,
		_w3579_,
		_w3580_,
		_w3581_,
		_w3582_
	);
	LUT3 #(
		.INIT('h48)
	) name2654 (
		\key_i[9]_pad ,
		_w931_,
		_w3582_,
		_w3583_
	);
	LUT4 #(
		.INIT('h3222)
	) name2655 (
		\data_o[9]_pad ,
		_w931_,
		_w934_,
		_w2784_,
		_w3584_
	);
	LUT4 #(
		.INIT('h7b00)
	) name2656 (
		\ks1_key_reg_reg[9]/NET0131 ,
		_w2785_,
		_w3582_,
		_w3584_,
		_w3585_
	);
	LUT2 #(
		.INIT('he)
	) name2657 (
		_w3583_,
		_w3585_,
		_w3586_
	);
	LUT4 #(
		.INIT('haab8)
	) name2658 (
		\data_i[38]_pad ,
		decrypt_i_pad,
		\mix1_data_o_reg_reg[38]/NET0131 ,
		_w930_,
		_w3587_
	);
	LUT4 #(
		.INIT('haba8)
	) name2659 (
		\sub1_data_reg_reg[38]/NET0131 ,
		_w996_,
		_w2776_,
		_w3587_,
		_w3588_
	);
	LUT4 #(
		.INIT('h404c)
	) name2660 (
		\mix1_data_o_reg_reg[38]/NET0131 ,
		_w2774_,
		_w2775_,
		_w3588_,
		_w3589_
	);
	LUT4 #(
		.INIT('h0545)
	) name2661 (
		\sub1_data_reg_reg[38]/NET0131 ,
		\sub1_ready_o_reg/NET0131 ,
		_w1054_,
		_w2230_,
		_w3590_
	);
	LUT4 #(
		.INIT('h1015)
	) name2662 (
		\state_reg/NET0131 ,
		\sub1_data_reg_reg[38]/NET0131 ,
		_w996_,
		_w3587_,
		_w3591_
	);
	LUT4 #(
		.INIT('h0057)
	) name2663 (
		\state_reg/NET0131 ,
		_w3589_,
		_w3590_,
		_w3591_,
		_w3592_
	);
	LUT3 #(
		.INIT('h48)
	) name2664 (
		\key_i[38]_pad ,
		_w931_,
		_w3592_,
		_w3593_
	);
	LUT4 #(
		.INIT('h3222)
	) name2665 (
		\data_o[38]_pad ,
		_w931_,
		_w934_,
		_w2784_,
		_w3594_
	);
	LUT4 #(
		.INIT('h7b00)
	) name2666 (
		\ks1_key_reg_reg[38]/NET0131 ,
		_w2785_,
		_w3592_,
		_w3594_,
		_w3595_
	);
	LUT2 #(
		.INIT('he)
	) name2667 (
		_w3593_,
		_w3595_,
		_w3596_
	);
	LUT4 #(
		.INIT('h5547)
	) name2668 (
		\data_i[106]_pad ,
		decrypt_i_pad,
		\mix1_data_o_reg_reg[106]/NET0131 ,
		_w930_,
		_w3597_
	);
	LUT4 #(
		.INIT('ha8ab)
	) name2669 (
		\sub1_data_reg_reg[106]/NET0131 ,
		_w996_,
		_w2776_,
		_w3597_,
		_w3598_
	);
	LUT4 #(
		.INIT('h404c)
	) name2670 (
		\mix1_data_o_reg_reg[106]/NET0131 ,
		_w2774_,
		_w2775_,
		_w3598_,
		_w3599_
	);
	LUT4 #(
		.INIT('h0545)
	) name2671 (
		\sub1_data_reg_reg[106]/NET0131 ,
		\sub1_ready_o_reg/NET0131 ,
		_w1054_,
		_w2230_,
		_w3600_
	);
	LUT4 #(
		.INIT('h1510)
	) name2672 (
		\state_reg/NET0131 ,
		\sub1_data_reg_reg[106]/NET0131 ,
		_w996_,
		_w3597_,
		_w3601_
	);
	LUT4 #(
		.INIT('h0057)
	) name2673 (
		\state_reg/NET0131 ,
		_w3599_,
		_w3600_,
		_w3601_,
		_w3602_
	);
	LUT3 #(
		.INIT('h48)
	) name2674 (
		\key_i[106]_pad ,
		_w931_,
		_w3602_,
		_w3603_
	);
	LUT4 #(
		.INIT('h3222)
	) name2675 (
		\data_o[106]_pad ,
		_w931_,
		_w934_,
		_w2784_,
		_w3604_
	);
	LUT4 #(
		.INIT('h7b00)
	) name2676 (
		\ks1_key_reg_reg[106]/NET0131 ,
		_w2785_,
		_w3602_,
		_w3604_,
		_w3605_
	);
	LUT2 #(
		.INIT('he)
	) name2677 (
		_w3603_,
		_w3605_,
		_w3606_
	);
	LUT4 #(
		.INIT('h5547)
	) name2678 (
		\data_i[122]_pad ,
		decrypt_i_pad,
		\mix1_data_o_reg_reg[122]/NET0131 ,
		_w930_,
		_w3607_
	);
	LUT4 #(
		.INIT('ha8ab)
	) name2679 (
		\sub1_data_reg_reg[122]/NET0131 ,
		_w996_,
		_w2776_,
		_w3607_,
		_w3608_
	);
	LUT4 #(
		.INIT('h404c)
	) name2680 (
		\mix1_data_o_reg_reg[122]/NET0131 ,
		_w2774_,
		_w2775_,
		_w3608_,
		_w3609_
	);
	LUT4 #(
		.INIT('h0545)
	) name2681 (
		\sub1_data_reg_reg[122]/NET0131 ,
		\sub1_ready_o_reg/NET0131 ,
		_w1054_,
		_w2230_,
		_w3610_
	);
	LUT4 #(
		.INIT('h1510)
	) name2682 (
		\state_reg/NET0131 ,
		\sub1_data_reg_reg[122]/NET0131 ,
		_w996_,
		_w3607_,
		_w3611_
	);
	LUT4 #(
		.INIT('h0057)
	) name2683 (
		\state_reg/NET0131 ,
		_w3609_,
		_w3610_,
		_w3611_,
		_w3612_
	);
	LUT3 #(
		.INIT('h48)
	) name2684 (
		\key_i[122]_pad ,
		_w931_,
		_w3612_,
		_w3613_
	);
	LUT4 #(
		.INIT('h3222)
	) name2685 (
		\data_o[122]_pad ,
		_w931_,
		_w934_,
		_w2784_,
		_w3614_
	);
	LUT4 #(
		.INIT('h7b00)
	) name2686 (
		\ks1_key_reg_reg[122]/NET0131 ,
		_w2785_,
		_w3612_,
		_w3614_,
		_w3615_
	);
	LUT2 #(
		.INIT('he)
	) name2687 (
		_w3613_,
		_w3615_,
		_w3616_
	);
	LUT4 #(
		.INIT('haab8)
	) name2688 (
		\data_i[39]_pad ,
		decrypt_i_pad,
		\mix1_data_o_reg_reg[39]/NET0131 ,
		_w930_,
		_w3617_
	);
	LUT4 #(
		.INIT('haba8)
	) name2689 (
		\sub1_data_reg_reg[39]/NET0131 ,
		_w996_,
		_w2776_,
		_w3617_,
		_w3618_
	);
	LUT4 #(
		.INIT('h404c)
	) name2690 (
		\mix1_data_o_reg_reg[39]/NET0131 ,
		_w2774_,
		_w2775_,
		_w3618_,
		_w3619_
	);
	LUT4 #(
		.INIT('h0545)
	) name2691 (
		\sub1_data_reg_reg[39]/NET0131 ,
		\sub1_ready_o_reg/NET0131 ,
		_w1054_,
		_w2230_,
		_w3620_
	);
	LUT4 #(
		.INIT('h1015)
	) name2692 (
		\state_reg/NET0131 ,
		\sub1_data_reg_reg[39]/NET0131 ,
		_w996_,
		_w3617_,
		_w3621_
	);
	LUT4 #(
		.INIT('h0057)
	) name2693 (
		\state_reg/NET0131 ,
		_w3619_,
		_w3620_,
		_w3621_,
		_w3622_
	);
	LUT3 #(
		.INIT('h48)
	) name2694 (
		\key_i[39]_pad ,
		_w931_,
		_w3622_,
		_w3623_
	);
	LUT4 #(
		.INIT('h3222)
	) name2695 (
		\data_o[39]_pad ,
		_w931_,
		_w934_,
		_w2784_,
		_w3624_
	);
	LUT4 #(
		.INIT('h7b00)
	) name2696 (
		\ks1_key_reg_reg[39]/NET0131 ,
		_w2785_,
		_w3622_,
		_w3624_,
		_w3625_
	);
	LUT2 #(
		.INIT('he)
	) name2697 (
		_w3623_,
		_w3625_,
		_w3626_
	);
	LUT4 #(
		.INIT('h5547)
	) name2698 (
		\data_i[3]_pad ,
		decrypt_i_pad,
		\mix1_data_o_reg_reg[3]/NET0131 ,
		_w930_,
		_w3627_
	);
	LUT4 #(
		.INIT('ha8ab)
	) name2699 (
		\sub1_data_reg_reg[3]/NET0131 ,
		_w996_,
		_w2776_,
		_w3627_,
		_w3628_
	);
	LUT4 #(
		.INIT('h404c)
	) name2700 (
		\mix1_data_o_reg_reg[3]/NET0131 ,
		_w2774_,
		_w2775_,
		_w3628_,
		_w3629_
	);
	LUT4 #(
		.INIT('h0545)
	) name2701 (
		\sub1_data_reg_reg[3]/NET0131 ,
		\sub1_ready_o_reg/NET0131 ,
		_w1054_,
		_w2230_,
		_w3630_
	);
	LUT4 #(
		.INIT('h1510)
	) name2702 (
		\state_reg/NET0131 ,
		\sub1_data_reg_reg[3]/NET0131 ,
		_w996_,
		_w3627_,
		_w3631_
	);
	LUT4 #(
		.INIT('h0057)
	) name2703 (
		\state_reg/NET0131 ,
		_w3629_,
		_w3630_,
		_w3631_,
		_w3632_
	);
	LUT3 #(
		.INIT('h48)
	) name2704 (
		\key_i[3]_pad ,
		_w931_,
		_w3632_,
		_w3633_
	);
	LUT4 #(
		.INIT('h3222)
	) name2705 (
		\data_o[3]_pad ,
		_w931_,
		_w934_,
		_w2784_,
		_w3634_
	);
	LUT4 #(
		.INIT('h7b00)
	) name2706 (
		\ks1_key_reg_reg[3]/NET0131 ,
		_w2785_,
		_w3632_,
		_w3634_,
		_w3635_
	);
	LUT2 #(
		.INIT('he)
	) name2707 (
		_w3633_,
		_w3635_,
		_w3636_
	);
	LUT4 #(
		.INIT('h5547)
	) name2708 (
		\data_i[0]_pad ,
		decrypt_i_pad,
		\mix1_data_o_reg_reg[0]/NET0131 ,
		_w930_,
		_w3637_
	);
	LUT4 #(
		.INIT('ha8ab)
	) name2709 (
		\sub1_data_reg_reg[0]/NET0131 ,
		_w996_,
		_w2776_,
		_w3637_,
		_w3638_
	);
	LUT4 #(
		.INIT('h404c)
	) name2710 (
		\mix1_data_o_reg_reg[0]/NET0131 ,
		_w2774_,
		_w2775_,
		_w3638_,
		_w3639_
	);
	LUT4 #(
		.INIT('h0545)
	) name2711 (
		\sub1_data_reg_reg[0]/NET0131 ,
		\sub1_ready_o_reg/NET0131 ,
		_w1054_,
		_w2230_,
		_w3640_
	);
	LUT4 #(
		.INIT('h1510)
	) name2712 (
		\state_reg/NET0131 ,
		\sub1_data_reg_reg[0]/NET0131 ,
		_w996_,
		_w3637_,
		_w3641_
	);
	LUT4 #(
		.INIT('h0057)
	) name2713 (
		\state_reg/NET0131 ,
		_w3639_,
		_w3640_,
		_w3641_,
		_w3642_
	);
	LUT3 #(
		.INIT('h48)
	) name2714 (
		\key_i[0]_pad ,
		_w931_,
		_w3642_,
		_w3643_
	);
	LUT4 #(
		.INIT('h3222)
	) name2715 (
		\data_o[0]_pad ,
		_w931_,
		_w934_,
		_w2784_,
		_w3644_
	);
	LUT4 #(
		.INIT('h7b00)
	) name2716 (
		\ks1_key_reg_reg[0]/NET0131 ,
		_w2785_,
		_w3642_,
		_w3644_,
		_w3645_
	);
	LUT2 #(
		.INIT('he)
	) name2717 (
		_w3643_,
		_w3645_,
		_w3646_
	);
	LUT4 #(
		.INIT('h5547)
	) name2718 (
		\data_i[40]_pad ,
		decrypt_i_pad,
		\mix1_data_o_reg_reg[40]/NET0131 ,
		_w930_,
		_w3647_
	);
	LUT4 #(
		.INIT('ha8ab)
	) name2719 (
		\sub1_data_reg_reg[40]/NET0131 ,
		_w996_,
		_w2776_,
		_w3647_,
		_w3648_
	);
	LUT4 #(
		.INIT('h404c)
	) name2720 (
		\mix1_data_o_reg_reg[40]/NET0131 ,
		_w2774_,
		_w2775_,
		_w3648_,
		_w3649_
	);
	LUT4 #(
		.INIT('h0545)
	) name2721 (
		\sub1_data_reg_reg[40]/NET0131 ,
		\sub1_ready_o_reg/NET0131 ,
		_w1054_,
		_w2230_,
		_w3650_
	);
	LUT4 #(
		.INIT('h1510)
	) name2722 (
		\state_reg/NET0131 ,
		\sub1_data_reg_reg[40]/NET0131 ,
		_w996_,
		_w3647_,
		_w3651_
	);
	LUT4 #(
		.INIT('h0057)
	) name2723 (
		\state_reg/NET0131 ,
		_w3649_,
		_w3650_,
		_w3651_,
		_w3652_
	);
	LUT3 #(
		.INIT('h48)
	) name2724 (
		\key_i[40]_pad ,
		_w931_,
		_w3652_,
		_w3653_
	);
	LUT4 #(
		.INIT('h3222)
	) name2725 (
		\data_o[40]_pad ,
		_w931_,
		_w934_,
		_w2784_,
		_w3654_
	);
	LUT4 #(
		.INIT('h7b00)
	) name2726 (
		\ks1_key_reg_reg[40]/P0002 ,
		_w2785_,
		_w3652_,
		_w3654_,
		_w3655_
	);
	LUT2 #(
		.INIT('he)
	) name2727 (
		_w3653_,
		_w3655_,
		_w3656_
	);
	LUT4 #(
		.INIT('h5547)
	) name2728 (
		\data_i[123]_pad ,
		decrypt_i_pad,
		\mix1_data_o_reg_reg[123]/NET0131 ,
		_w930_,
		_w3657_
	);
	LUT4 #(
		.INIT('ha8ab)
	) name2729 (
		\sub1_data_reg_reg[123]/NET0131 ,
		_w996_,
		_w2776_,
		_w3657_,
		_w3658_
	);
	LUT4 #(
		.INIT('h404c)
	) name2730 (
		\mix1_data_o_reg_reg[123]/NET0131 ,
		_w2774_,
		_w2775_,
		_w3658_,
		_w3659_
	);
	LUT4 #(
		.INIT('h0545)
	) name2731 (
		\sub1_data_reg_reg[123]/NET0131 ,
		\sub1_ready_o_reg/NET0131 ,
		_w1054_,
		_w2230_,
		_w3660_
	);
	LUT4 #(
		.INIT('h1510)
	) name2732 (
		\state_reg/NET0131 ,
		\sub1_data_reg_reg[123]/NET0131 ,
		_w996_,
		_w3657_,
		_w3661_
	);
	LUT4 #(
		.INIT('h0057)
	) name2733 (
		\state_reg/NET0131 ,
		_w3659_,
		_w3660_,
		_w3661_,
		_w3662_
	);
	LUT3 #(
		.INIT('h48)
	) name2734 (
		\key_i[123]_pad ,
		_w931_,
		_w3662_,
		_w3663_
	);
	LUT4 #(
		.INIT('h3222)
	) name2735 (
		\data_o[123]_pad ,
		_w931_,
		_w934_,
		_w2784_,
		_w3664_
	);
	LUT4 #(
		.INIT('h7b00)
	) name2736 (
		\ks1_key_reg_reg[123]/NET0131 ,
		_w2785_,
		_w3662_,
		_w3664_,
		_w3665_
	);
	LUT2 #(
		.INIT('he)
	) name2737 (
		_w3663_,
		_w3665_,
		_w3666_
	);
	LUT4 #(
		.INIT('h5547)
	) name2738 (
		\data_i[41]_pad ,
		decrypt_i_pad,
		\mix1_data_o_reg_reg[41]/NET0131 ,
		_w930_,
		_w3667_
	);
	LUT4 #(
		.INIT('ha8ab)
	) name2739 (
		\sub1_data_reg_reg[41]/NET0131 ,
		_w996_,
		_w2776_,
		_w3667_,
		_w3668_
	);
	LUT4 #(
		.INIT('h404c)
	) name2740 (
		\mix1_data_o_reg_reg[41]/NET0131 ,
		_w2774_,
		_w2775_,
		_w3668_,
		_w3669_
	);
	LUT4 #(
		.INIT('h0545)
	) name2741 (
		\sub1_data_reg_reg[41]/NET0131 ,
		\sub1_ready_o_reg/NET0131 ,
		_w1054_,
		_w2230_,
		_w3670_
	);
	LUT4 #(
		.INIT('h1510)
	) name2742 (
		\state_reg/NET0131 ,
		\sub1_data_reg_reg[41]/NET0131 ,
		_w996_,
		_w3667_,
		_w3671_
	);
	LUT4 #(
		.INIT('h0057)
	) name2743 (
		\state_reg/NET0131 ,
		_w3669_,
		_w3670_,
		_w3671_,
		_w3672_
	);
	LUT3 #(
		.INIT('h48)
	) name2744 (
		\key_i[41]_pad ,
		_w931_,
		_w3672_,
		_w3673_
	);
	LUT4 #(
		.INIT('h3222)
	) name2745 (
		\data_o[41]_pad ,
		_w931_,
		_w934_,
		_w2784_,
		_w3674_
	);
	LUT4 #(
		.INIT('h7b00)
	) name2746 (
		\ks1_key_reg_reg[41]/P0002 ,
		_w2785_,
		_w3672_,
		_w3674_,
		_w3675_
	);
	LUT2 #(
		.INIT('he)
	) name2747 (
		_w3673_,
		_w3675_,
		_w3676_
	);
	LUT4 #(
		.INIT('h5547)
	) name2748 (
		\data_i[47]_pad ,
		decrypt_i_pad,
		\mix1_data_o_reg_reg[47]/NET0131 ,
		_w930_,
		_w3677_
	);
	LUT4 #(
		.INIT('ha8ab)
	) name2749 (
		\sub1_data_reg_reg[47]/NET0131 ,
		_w996_,
		_w2776_,
		_w3677_,
		_w3678_
	);
	LUT4 #(
		.INIT('h404c)
	) name2750 (
		\mix1_data_o_reg_reg[47]/NET0131 ,
		_w2774_,
		_w2775_,
		_w3678_,
		_w3679_
	);
	LUT4 #(
		.INIT('h0545)
	) name2751 (
		\sub1_data_reg_reg[47]/NET0131 ,
		\sub1_ready_o_reg/NET0131 ,
		_w1054_,
		_w2230_,
		_w3680_
	);
	LUT4 #(
		.INIT('h1510)
	) name2752 (
		\state_reg/NET0131 ,
		\sub1_data_reg_reg[47]/NET0131 ,
		_w996_,
		_w3677_,
		_w3681_
	);
	LUT4 #(
		.INIT('h0057)
	) name2753 (
		\state_reg/NET0131 ,
		_w3679_,
		_w3680_,
		_w3681_,
		_w3682_
	);
	LUT3 #(
		.INIT('h48)
	) name2754 (
		\key_i[47]_pad ,
		_w931_,
		_w3682_,
		_w3683_
	);
	LUT4 #(
		.INIT('h3222)
	) name2755 (
		\data_o[47]_pad ,
		_w931_,
		_w934_,
		_w2784_,
		_w3684_
	);
	LUT4 #(
		.INIT('h7b00)
	) name2756 (
		\ks1_key_reg_reg[47]/P0002 ,
		_w2785_,
		_w3682_,
		_w3684_,
		_w3685_
	);
	LUT2 #(
		.INIT('he)
	) name2757 (
		_w3683_,
		_w3685_,
		_w3686_
	);
	LUT4 #(
		.INIT('h5547)
	) name2758 (
		\data_i[42]_pad ,
		decrypt_i_pad,
		\mix1_data_o_reg_reg[42]/NET0131 ,
		_w930_,
		_w3687_
	);
	LUT4 #(
		.INIT('ha8ab)
	) name2759 (
		\sub1_data_reg_reg[42]/NET0131 ,
		_w996_,
		_w2776_,
		_w3687_,
		_w3688_
	);
	LUT4 #(
		.INIT('h404c)
	) name2760 (
		\mix1_data_o_reg_reg[42]/NET0131 ,
		_w2774_,
		_w2775_,
		_w3688_,
		_w3689_
	);
	LUT4 #(
		.INIT('h0545)
	) name2761 (
		\sub1_data_reg_reg[42]/NET0131 ,
		\sub1_ready_o_reg/NET0131 ,
		_w1054_,
		_w2230_,
		_w3690_
	);
	LUT4 #(
		.INIT('h1510)
	) name2762 (
		\state_reg/NET0131 ,
		\sub1_data_reg_reg[42]/NET0131 ,
		_w996_,
		_w3687_,
		_w3691_
	);
	LUT4 #(
		.INIT('h0057)
	) name2763 (
		\state_reg/NET0131 ,
		_w3689_,
		_w3690_,
		_w3691_,
		_w3692_
	);
	LUT3 #(
		.INIT('h48)
	) name2764 (
		\key_i[42]_pad ,
		_w931_,
		_w3692_,
		_w3693_
	);
	LUT4 #(
		.INIT('h3222)
	) name2765 (
		\data_o[42]_pad ,
		_w931_,
		_w934_,
		_w2784_,
		_w3694_
	);
	LUT4 #(
		.INIT('h7b00)
	) name2766 (
		\ks1_key_reg_reg[42]/P0002 ,
		_w2785_,
		_w3692_,
		_w3694_,
		_w3695_
	);
	LUT2 #(
		.INIT('he)
	) name2767 (
		_w3693_,
		_w3695_,
		_w3696_
	);
	LUT4 #(
		.INIT('h5547)
	) name2768 (
		\data_i[124]_pad ,
		decrypt_i_pad,
		\mix1_data_o_reg_reg[124]/NET0131 ,
		_w930_,
		_w3697_
	);
	LUT4 #(
		.INIT('ha8ab)
	) name2769 (
		\sub1_data_reg_reg[124]/NET0131 ,
		_w996_,
		_w2776_,
		_w3697_,
		_w3698_
	);
	LUT4 #(
		.INIT('h404c)
	) name2770 (
		\mix1_data_o_reg_reg[124]/NET0131 ,
		_w2774_,
		_w2775_,
		_w3698_,
		_w3699_
	);
	LUT4 #(
		.INIT('h0545)
	) name2771 (
		\sub1_data_reg_reg[124]/NET0131 ,
		\sub1_ready_o_reg/NET0131 ,
		_w1054_,
		_w2230_,
		_w3700_
	);
	LUT4 #(
		.INIT('h1510)
	) name2772 (
		\state_reg/NET0131 ,
		\sub1_data_reg_reg[124]/NET0131 ,
		_w996_,
		_w3697_,
		_w3701_
	);
	LUT4 #(
		.INIT('h0057)
	) name2773 (
		\state_reg/NET0131 ,
		_w3699_,
		_w3700_,
		_w3701_,
		_w3702_
	);
	LUT3 #(
		.INIT('h48)
	) name2774 (
		\key_i[124]_pad ,
		_w931_,
		_w3702_,
		_w3703_
	);
	LUT4 #(
		.INIT('h3222)
	) name2775 (
		\data_o[124]_pad ,
		_w931_,
		_w934_,
		_w2784_,
		_w3704_
	);
	LUT4 #(
		.INIT('h7b00)
	) name2776 (
		\ks1_key_reg_reg[124]/NET0131 ,
		_w2785_,
		_w3702_,
		_w3704_,
		_w3705_
	);
	LUT2 #(
		.INIT('he)
	) name2777 (
		_w3703_,
		_w3705_,
		_w3706_
	);
	LUT4 #(
		.INIT('h5547)
	) name2778 (
		\data_i[43]_pad ,
		decrypt_i_pad,
		\mix1_data_o_reg_reg[43]/NET0131 ,
		_w930_,
		_w3707_
	);
	LUT4 #(
		.INIT('ha8ab)
	) name2779 (
		\sub1_data_reg_reg[43]/NET0131 ,
		_w996_,
		_w2776_,
		_w3707_,
		_w3708_
	);
	LUT4 #(
		.INIT('h404c)
	) name2780 (
		\mix1_data_o_reg_reg[43]/NET0131 ,
		_w2774_,
		_w2775_,
		_w3708_,
		_w3709_
	);
	LUT4 #(
		.INIT('h0545)
	) name2781 (
		\sub1_data_reg_reg[43]/NET0131 ,
		\sub1_ready_o_reg/NET0131 ,
		_w1054_,
		_w2230_,
		_w3710_
	);
	LUT4 #(
		.INIT('h1510)
	) name2782 (
		\state_reg/NET0131 ,
		\sub1_data_reg_reg[43]/NET0131 ,
		_w996_,
		_w3707_,
		_w3711_
	);
	LUT4 #(
		.INIT('h0057)
	) name2783 (
		\state_reg/NET0131 ,
		_w3709_,
		_w3710_,
		_w3711_,
		_w3712_
	);
	LUT3 #(
		.INIT('h48)
	) name2784 (
		\key_i[43]_pad ,
		_w931_,
		_w3712_,
		_w3713_
	);
	LUT4 #(
		.INIT('h3222)
	) name2785 (
		\data_o[43]_pad ,
		_w931_,
		_w934_,
		_w2784_,
		_w3714_
	);
	LUT4 #(
		.INIT('h7b00)
	) name2786 (
		\ks1_key_reg_reg[43]/P0002 ,
		_w2785_,
		_w3712_,
		_w3714_,
		_w3715_
	);
	LUT2 #(
		.INIT('he)
	) name2787 (
		_w3713_,
		_w3715_,
		_w3716_
	);
	LUT4 #(
		.INIT('h5547)
	) name2788 (
		\data_i[107]_pad ,
		decrypt_i_pad,
		\mix1_data_o_reg_reg[107]/NET0131 ,
		_w930_,
		_w3717_
	);
	LUT4 #(
		.INIT('ha8ab)
	) name2789 (
		\sub1_data_reg_reg[107]/NET0131 ,
		_w996_,
		_w2776_,
		_w3717_,
		_w3718_
	);
	LUT4 #(
		.INIT('h404c)
	) name2790 (
		\mix1_data_o_reg_reg[107]/NET0131 ,
		_w2774_,
		_w2775_,
		_w3718_,
		_w3719_
	);
	LUT4 #(
		.INIT('h0545)
	) name2791 (
		\sub1_data_reg_reg[107]/NET0131 ,
		\sub1_ready_o_reg/NET0131 ,
		_w1054_,
		_w2230_,
		_w3720_
	);
	LUT4 #(
		.INIT('h1510)
	) name2792 (
		\state_reg/NET0131 ,
		\sub1_data_reg_reg[107]/NET0131 ,
		_w996_,
		_w3717_,
		_w3721_
	);
	LUT4 #(
		.INIT('h0057)
	) name2793 (
		\state_reg/NET0131 ,
		_w3719_,
		_w3720_,
		_w3721_,
		_w3722_
	);
	LUT3 #(
		.INIT('h48)
	) name2794 (
		\key_i[107]_pad ,
		_w931_,
		_w3722_,
		_w3723_
	);
	LUT4 #(
		.INIT('h3222)
	) name2795 (
		\data_o[107]_pad ,
		_w931_,
		_w934_,
		_w2784_,
		_w3724_
	);
	LUT4 #(
		.INIT('h7b00)
	) name2796 (
		\ks1_key_reg_reg[107]/NET0131 ,
		_w2785_,
		_w3722_,
		_w3724_,
		_w3725_
	);
	LUT2 #(
		.INIT('he)
	) name2797 (
		_w3723_,
		_w3725_,
		_w3726_
	);
	LUT4 #(
		.INIT('h5547)
	) name2798 (
		\data_i[125]_pad ,
		decrypt_i_pad,
		\mix1_data_o_reg_reg[125]/NET0131 ,
		_w930_,
		_w3727_
	);
	LUT4 #(
		.INIT('ha8ab)
	) name2799 (
		\sub1_data_reg_reg[125]/NET0131 ,
		_w996_,
		_w2776_,
		_w3727_,
		_w3728_
	);
	LUT4 #(
		.INIT('h404c)
	) name2800 (
		\mix1_data_o_reg_reg[125]/NET0131 ,
		_w2774_,
		_w2775_,
		_w3728_,
		_w3729_
	);
	LUT4 #(
		.INIT('h0545)
	) name2801 (
		\sub1_data_reg_reg[125]/NET0131 ,
		\sub1_ready_o_reg/NET0131 ,
		_w1054_,
		_w2230_,
		_w3730_
	);
	LUT4 #(
		.INIT('h1510)
	) name2802 (
		\state_reg/NET0131 ,
		\sub1_data_reg_reg[125]/NET0131 ,
		_w996_,
		_w3727_,
		_w3731_
	);
	LUT4 #(
		.INIT('h0057)
	) name2803 (
		\state_reg/NET0131 ,
		_w3729_,
		_w3730_,
		_w3731_,
		_w3732_
	);
	LUT3 #(
		.INIT('h48)
	) name2804 (
		\key_i[125]_pad ,
		_w931_,
		_w3732_,
		_w3733_
	);
	LUT4 #(
		.INIT('h3222)
	) name2805 (
		\data_o[125]_pad ,
		_w931_,
		_w934_,
		_w2784_,
		_w3734_
	);
	LUT4 #(
		.INIT('h7b00)
	) name2806 (
		\ks1_key_reg_reg[125]/NET0131 ,
		_w2785_,
		_w3732_,
		_w3734_,
		_w3735_
	);
	LUT2 #(
		.INIT('he)
	) name2807 (
		_w3733_,
		_w3735_,
		_w3736_
	);
	LUT4 #(
		.INIT('h5547)
	) name2808 (
		\data_i[44]_pad ,
		decrypt_i_pad,
		\mix1_data_o_reg_reg[44]/NET0131 ,
		_w930_,
		_w3737_
	);
	LUT4 #(
		.INIT('ha8ab)
	) name2809 (
		\sub1_data_reg_reg[44]/NET0131 ,
		_w996_,
		_w2776_,
		_w3737_,
		_w3738_
	);
	LUT4 #(
		.INIT('h404c)
	) name2810 (
		\mix1_data_o_reg_reg[44]/NET0131 ,
		_w2774_,
		_w2775_,
		_w3738_,
		_w3739_
	);
	LUT4 #(
		.INIT('h0545)
	) name2811 (
		\sub1_data_reg_reg[44]/NET0131 ,
		\sub1_ready_o_reg/NET0131 ,
		_w1054_,
		_w2230_,
		_w3740_
	);
	LUT4 #(
		.INIT('h1510)
	) name2812 (
		\state_reg/NET0131 ,
		\sub1_data_reg_reg[44]/NET0131 ,
		_w996_,
		_w3737_,
		_w3741_
	);
	LUT4 #(
		.INIT('h0057)
	) name2813 (
		\state_reg/NET0131 ,
		_w3739_,
		_w3740_,
		_w3741_,
		_w3742_
	);
	LUT3 #(
		.INIT('h48)
	) name2814 (
		\key_i[44]_pad ,
		_w931_,
		_w3742_,
		_w3743_
	);
	LUT4 #(
		.INIT('h3222)
	) name2815 (
		\data_o[44]_pad ,
		_w931_,
		_w934_,
		_w2784_,
		_w3744_
	);
	LUT4 #(
		.INIT('h7b00)
	) name2816 (
		\ks1_key_reg_reg[44]/P0002 ,
		_w2785_,
		_w3742_,
		_w3744_,
		_w3745_
	);
	LUT2 #(
		.INIT('he)
	) name2817 (
		_w3743_,
		_w3745_,
		_w3746_
	);
	LUT4 #(
		.INIT('h5547)
	) name2818 (
		\data_i[108]_pad ,
		decrypt_i_pad,
		\mix1_data_o_reg_reg[108]/NET0131 ,
		_w930_,
		_w3747_
	);
	LUT4 #(
		.INIT('ha8ab)
	) name2819 (
		\sub1_data_reg_reg[108]/NET0131 ,
		_w996_,
		_w2776_,
		_w3747_,
		_w3748_
	);
	LUT4 #(
		.INIT('h404c)
	) name2820 (
		\mix1_data_o_reg_reg[108]/NET0131 ,
		_w2774_,
		_w2775_,
		_w3748_,
		_w3749_
	);
	LUT4 #(
		.INIT('h0545)
	) name2821 (
		\sub1_data_reg_reg[108]/NET0131 ,
		\sub1_ready_o_reg/NET0131 ,
		_w1054_,
		_w2230_,
		_w3750_
	);
	LUT4 #(
		.INIT('h1510)
	) name2822 (
		\state_reg/NET0131 ,
		\sub1_data_reg_reg[108]/NET0131 ,
		_w996_,
		_w3747_,
		_w3751_
	);
	LUT4 #(
		.INIT('h0057)
	) name2823 (
		\state_reg/NET0131 ,
		_w3749_,
		_w3750_,
		_w3751_,
		_w3752_
	);
	LUT3 #(
		.INIT('h48)
	) name2824 (
		\key_i[108]_pad ,
		_w931_,
		_w3752_,
		_w3753_
	);
	LUT4 #(
		.INIT('h3222)
	) name2825 (
		\data_o[108]_pad ,
		_w931_,
		_w934_,
		_w2784_,
		_w3754_
	);
	LUT4 #(
		.INIT('h7b00)
	) name2826 (
		\ks1_key_reg_reg[108]/NET0131 ,
		_w2785_,
		_w3752_,
		_w3754_,
		_w3755_
	);
	LUT2 #(
		.INIT('he)
	) name2827 (
		_w3753_,
		_w3755_,
		_w3756_
	);
	LUT4 #(
		.INIT('h5547)
	) name2828 (
		\data_i[45]_pad ,
		decrypt_i_pad,
		\mix1_data_o_reg_reg[45]/NET0131 ,
		_w930_,
		_w3757_
	);
	LUT4 #(
		.INIT('ha8ab)
	) name2829 (
		\sub1_data_reg_reg[45]/NET0131 ,
		_w996_,
		_w2776_,
		_w3757_,
		_w3758_
	);
	LUT4 #(
		.INIT('h404c)
	) name2830 (
		\mix1_data_o_reg_reg[45]/NET0131 ,
		_w2774_,
		_w2775_,
		_w3758_,
		_w3759_
	);
	LUT4 #(
		.INIT('h0545)
	) name2831 (
		\sub1_data_reg_reg[45]/NET0131 ,
		\sub1_ready_o_reg/NET0131 ,
		_w1054_,
		_w2230_,
		_w3760_
	);
	LUT4 #(
		.INIT('h1510)
	) name2832 (
		\state_reg/NET0131 ,
		\sub1_data_reg_reg[45]/NET0131 ,
		_w996_,
		_w3757_,
		_w3761_
	);
	LUT4 #(
		.INIT('h0057)
	) name2833 (
		\state_reg/NET0131 ,
		_w3759_,
		_w3760_,
		_w3761_,
		_w3762_
	);
	LUT3 #(
		.INIT('h48)
	) name2834 (
		\key_i[45]_pad ,
		_w931_,
		_w3762_,
		_w3763_
	);
	LUT4 #(
		.INIT('h3222)
	) name2835 (
		\data_o[45]_pad ,
		_w931_,
		_w934_,
		_w2784_,
		_w3764_
	);
	LUT4 #(
		.INIT('h7b00)
	) name2836 (
		\ks1_key_reg_reg[45]/P0002 ,
		_w2785_,
		_w3762_,
		_w3764_,
		_w3765_
	);
	LUT2 #(
		.INIT('he)
	) name2837 (
		_w3763_,
		_w3765_,
		_w3766_
	);
	LUT4 #(
		.INIT('h5547)
	) name2838 (
		\data_i[46]_pad ,
		decrypt_i_pad,
		\mix1_data_o_reg_reg[46]/NET0131 ,
		_w930_,
		_w3767_
	);
	LUT4 #(
		.INIT('ha8ab)
	) name2839 (
		\sub1_data_reg_reg[46]/NET0131 ,
		_w996_,
		_w2776_,
		_w3767_,
		_w3768_
	);
	LUT4 #(
		.INIT('h404c)
	) name2840 (
		\mix1_data_o_reg_reg[46]/NET0131 ,
		_w2774_,
		_w2775_,
		_w3768_,
		_w3769_
	);
	LUT4 #(
		.INIT('h0545)
	) name2841 (
		\sub1_data_reg_reg[46]/NET0131 ,
		\sub1_ready_o_reg/NET0131 ,
		_w1054_,
		_w2230_,
		_w3770_
	);
	LUT4 #(
		.INIT('h1510)
	) name2842 (
		\state_reg/NET0131 ,
		\sub1_data_reg_reg[46]/NET0131 ,
		_w996_,
		_w3767_,
		_w3771_
	);
	LUT4 #(
		.INIT('h0057)
	) name2843 (
		\state_reg/NET0131 ,
		_w3769_,
		_w3770_,
		_w3771_,
		_w3772_
	);
	LUT3 #(
		.INIT('h48)
	) name2844 (
		\key_i[46]_pad ,
		_w931_,
		_w3772_,
		_w3773_
	);
	LUT4 #(
		.INIT('h3222)
	) name2845 (
		\data_o[46]_pad ,
		_w931_,
		_w934_,
		_w2784_,
		_w3774_
	);
	LUT4 #(
		.INIT('h7b00)
	) name2846 (
		\ks1_key_reg_reg[46]/P0002 ,
		_w2785_,
		_w3772_,
		_w3774_,
		_w3775_
	);
	LUT2 #(
		.INIT('he)
	) name2847 (
		_w3773_,
		_w3775_,
		_w3776_
	);
	LUT4 #(
		.INIT('h5547)
	) name2848 (
		\data_i[126]_pad ,
		decrypt_i_pad,
		\mix1_data_o_reg_reg[126]/NET0131 ,
		_w930_,
		_w3777_
	);
	LUT4 #(
		.INIT('ha8ab)
	) name2849 (
		\sub1_data_reg_reg[126]/NET0131 ,
		_w996_,
		_w2776_,
		_w3777_,
		_w3778_
	);
	LUT4 #(
		.INIT('h404c)
	) name2850 (
		\mix1_data_o_reg_reg[126]/NET0131 ,
		_w2774_,
		_w2775_,
		_w3778_,
		_w3779_
	);
	LUT4 #(
		.INIT('h0545)
	) name2851 (
		\sub1_data_reg_reg[126]/NET0131 ,
		\sub1_ready_o_reg/NET0131 ,
		_w1054_,
		_w2230_,
		_w3780_
	);
	LUT4 #(
		.INIT('h1510)
	) name2852 (
		\state_reg/NET0131 ,
		\sub1_data_reg_reg[126]/NET0131 ,
		_w996_,
		_w3777_,
		_w3781_
	);
	LUT4 #(
		.INIT('h0057)
	) name2853 (
		\state_reg/NET0131 ,
		_w3779_,
		_w3780_,
		_w3781_,
		_w3782_
	);
	LUT3 #(
		.INIT('h48)
	) name2854 (
		\key_i[126]_pad ,
		_w931_,
		_w3782_,
		_w3783_
	);
	LUT4 #(
		.INIT('h3222)
	) name2855 (
		\data_o[126]_pad ,
		_w931_,
		_w934_,
		_w2784_,
		_w3784_
	);
	LUT4 #(
		.INIT('h7b00)
	) name2856 (
		\ks1_key_reg_reg[126]/NET0131 ,
		_w2785_,
		_w3782_,
		_w3784_,
		_w3785_
	);
	LUT2 #(
		.INIT('he)
	) name2857 (
		_w3783_,
		_w3785_,
		_w3786_
	);
	LUT4 #(
		.INIT('haab8)
	) name2858 (
		\data_i[48]_pad ,
		decrypt_i_pad,
		\mix1_data_o_reg_reg[48]/NET0131 ,
		_w930_,
		_w3787_
	);
	LUT4 #(
		.INIT('haba8)
	) name2859 (
		\sub1_data_reg_reg[48]/NET0131 ,
		_w996_,
		_w2776_,
		_w3787_,
		_w3788_
	);
	LUT4 #(
		.INIT('h404c)
	) name2860 (
		\mix1_data_o_reg_reg[48]/NET0131 ,
		_w2774_,
		_w2775_,
		_w3788_,
		_w3789_
	);
	LUT4 #(
		.INIT('h0545)
	) name2861 (
		\sub1_data_reg_reg[48]/NET0131 ,
		\sub1_ready_o_reg/NET0131 ,
		_w1054_,
		_w2230_,
		_w3790_
	);
	LUT4 #(
		.INIT('h1015)
	) name2862 (
		\state_reg/NET0131 ,
		\sub1_data_reg_reg[48]/NET0131 ,
		_w996_,
		_w3787_,
		_w3791_
	);
	LUT4 #(
		.INIT('h0057)
	) name2863 (
		\state_reg/NET0131 ,
		_w3789_,
		_w3790_,
		_w3791_,
		_w3792_
	);
	LUT3 #(
		.INIT('h48)
	) name2864 (
		\key_i[48]_pad ,
		_w931_,
		_w3792_,
		_w3793_
	);
	LUT4 #(
		.INIT('h3222)
	) name2865 (
		\data_o[48]_pad ,
		_w931_,
		_w934_,
		_w2784_,
		_w3794_
	);
	LUT4 #(
		.INIT('h7b00)
	) name2866 (
		\ks1_key_reg_reg[48]/NET0131 ,
		_w2785_,
		_w3792_,
		_w3794_,
		_w3795_
	);
	LUT2 #(
		.INIT('he)
	) name2867 (
		_w3793_,
		_w3795_,
		_w3796_
	);
	LUT4 #(
		.INIT('h5547)
	) name2868 (
		\data_i[127]_pad ,
		decrypt_i_pad,
		\mix1_data_o_reg_reg[127]/NET0131 ,
		_w930_,
		_w3797_
	);
	LUT4 #(
		.INIT('ha8ab)
	) name2869 (
		\sub1_data_reg_reg[127]/NET0131 ,
		_w996_,
		_w2776_,
		_w3797_,
		_w3798_
	);
	LUT4 #(
		.INIT('h404c)
	) name2870 (
		\mix1_data_o_reg_reg[127]/NET0131 ,
		_w2774_,
		_w2775_,
		_w3798_,
		_w3799_
	);
	LUT4 #(
		.INIT('h0545)
	) name2871 (
		\sub1_data_reg_reg[127]/NET0131 ,
		\sub1_ready_o_reg/NET0131 ,
		_w1054_,
		_w2230_,
		_w3800_
	);
	LUT4 #(
		.INIT('h1510)
	) name2872 (
		\state_reg/NET0131 ,
		\sub1_data_reg_reg[127]/NET0131 ,
		_w996_,
		_w3797_,
		_w3801_
	);
	LUT4 #(
		.INIT('h0057)
	) name2873 (
		\state_reg/NET0131 ,
		_w3799_,
		_w3800_,
		_w3801_,
		_w3802_
	);
	LUT3 #(
		.INIT('h48)
	) name2874 (
		\key_i[127]_pad ,
		_w931_,
		_w3802_,
		_w3803_
	);
	LUT4 #(
		.INIT('h3222)
	) name2875 (
		\data_o[127]_pad ,
		_w931_,
		_w934_,
		_w2784_,
		_w3804_
	);
	LUT4 #(
		.INIT('h7b00)
	) name2876 (
		\ks1_key_reg_reg[127]/NET0131 ,
		_w2785_,
		_w3802_,
		_w3804_,
		_w3805_
	);
	LUT2 #(
		.INIT('he)
	) name2877 (
		_w3803_,
		_w3805_,
		_w3806_
	);
	LUT4 #(
		.INIT('haab8)
	) name2878 (
		\data_i[49]_pad ,
		decrypt_i_pad,
		\mix1_data_o_reg_reg[49]/NET0131 ,
		_w930_,
		_w3807_
	);
	LUT4 #(
		.INIT('haba8)
	) name2879 (
		\sub1_data_reg_reg[49]/NET0131 ,
		_w996_,
		_w2776_,
		_w3807_,
		_w3808_
	);
	LUT4 #(
		.INIT('h404c)
	) name2880 (
		\mix1_data_o_reg_reg[49]/NET0131 ,
		_w2774_,
		_w2775_,
		_w3808_,
		_w3809_
	);
	LUT4 #(
		.INIT('h0545)
	) name2881 (
		\sub1_data_reg_reg[49]/NET0131 ,
		\sub1_ready_o_reg/NET0131 ,
		_w1054_,
		_w2230_,
		_w3810_
	);
	LUT4 #(
		.INIT('h1015)
	) name2882 (
		\state_reg/NET0131 ,
		\sub1_data_reg_reg[49]/NET0131 ,
		_w996_,
		_w3807_,
		_w3811_
	);
	LUT4 #(
		.INIT('h0057)
	) name2883 (
		\state_reg/NET0131 ,
		_w3809_,
		_w3810_,
		_w3811_,
		_w3812_
	);
	LUT3 #(
		.INIT('h48)
	) name2884 (
		\key_i[49]_pad ,
		_w931_,
		_w3812_,
		_w3813_
	);
	LUT4 #(
		.INIT('h3222)
	) name2885 (
		\data_o[49]_pad ,
		_w931_,
		_w934_,
		_w2784_,
		_w3814_
	);
	LUT4 #(
		.INIT('h7b00)
	) name2886 (
		\ks1_key_reg_reg[49]/NET0131 ,
		_w2785_,
		_w3812_,
		_w3814_,
		_w3815_
	);
	LUT2 #(
		.INIT('he)
	) name2887 (
		_w3813_,
		_w3815_,
		_w3816_
	);
	LUT4 #(
		.INIT('h5547)
	) name2888 (
		\data_i[109]_pad ,
		decrypt_i_pad,
		\mix1_data_o_reg_reg[109]/NET0131 ,
		_w930_,
		_w3817_
	);
	LUT4 #(
		.INIT('ha8ab)
	) name2889 (
		\sub1_data_reg_reg[109]/NET0131 ,
		_w996_,
		_w2776_,
		_w3817_,
		_w3818_
	);
	LUT4 #(
		.INIT('h404c)
	) name2890 (
		\mix1_data_o_reg_reg[109]/NET0131 ,
		_w2774_,
		_w2775_,
		_w3818_,
		_w3819_
	);
	LUT4 #(
		.INIT('h0545)
	) name2891 (
		\sub1_data_reg_reg[109]/NET0131 ,
		\sub1_ready_o_reg/NET0131 ,
		_w1054_,
		_w2230_,
		_w3820_
	);
	LUT4 #(
		.INIT('h1510)
	) name2892 (
		\state_reg/NET0131 ,
		\sub1_data_reg_reg[109]/NET0131 ,
		_w996_,
		_w3817_,
		_w3821_
	);
	LUT4 #(
		.INIT('h0057)
	) name2893 (
		\state_reg/NET0131 ,
		_w3819_,
		_w3820_,
		_w3821_,
		_w3822_
	);
	LUT3 #(
		.INIT('h48)
	) name2894 (
		\key_i[109]_pad ,
		_w931_,
		_w3822_,
		_w3823_
	);
	LUT4 #(
		.INIT('h3222)
	) name2895 (
		\data_o[109]_pad ,
		_w931_,
		_w934_,
		_w2784_,
		_w3824_
	);
	LUT4 #(
		.INIT('h7b00)
	) name2896 (
		\ks1_key_reg_reg[109]/P0002 ,
		_w2785_,
		_w3822_,
		_w3824_,
		_w3825_
	);
	LUT2 #(
		.INIT('he)
	) name2897 (
		_w3823_,
		_w3825_,
		_w3826_
	);
	LUT4 #(
		.INIT('h5547)
	) name2898 (
		\data_i[4]_pad ,
		decrypt_i_pad,
		\mix1_data_o_reg_reg[4]/NET0131 ,
		_w930_,
		_w3827_
	);
	LUT4 #(
		.INIT('ha8ab)
	) name2899 (
		\sub1_data_reg_reg[4]/NET0131 ,
		_w996_,
		_w2776_,
		_w3827_,
		_w3828_
	);
	LUT4 #(
		.INIT('h404c)
	) name2900 (
		\mix1_data_o_reg_reg[4]/NET0131 ,
		_w2774_,
		_w2775_,
		_w3828_,
		_w3829_
	);
	LUT4 #(
		.INIT('h0545)
	) name2901 (
		\sub1_data_reg_reg[4]/NET0131 ,
		\sub1_ready_o_reg/NET0131 ,
		_w1054_,
		_w2230_,
		_w3830_
	);
	LUT4 #(
		.INIT('h1510)
	) name2902 (
		\state_reg/NET0131 ,
		\sub1_data_reg_reg[4]/NET0131 ,
		_w996_,
		_w3827_,
		_w3831_
	);
	LUT4 #(
		.INIT('h0057)
	) name2903 (
		\state_reg/NET0131 ,
		_w3829_,
		_w3830_,
		_w3831_,
		_w3832_
	);
	LUT3 #(
		.INIT('h48)
	) name2904 (
		\key_i[4]_pad ,
		_w931_,
		_w3832_,
		_w3833_
	);
	LUT4 #(
		.INIT('h3222)
	) name2905 (
		\data_o[4]_pad ,
		_w931_,
		_w934_,
		_w2784_,
		_w3834_
	);
	LUT4 #(
		.INIT('h7b00)
	) name2906 (
		\ks1_key_reg_reg[4]/NET0131 ,
		_w2785_,
		_w3832_,
		_w3834_,
		_w3835_
	);
	LUT2 #(
		.INIT('he)
	) name2907 (
		_w3833_,
		_w3835_,
		_w3836_
	);
	LUT4 #(
		.INIT('h5547)
	) name2908 (
		\data_i[12]_pad ,
		decrypt_i_pad,
		\mix1_data_o_reg_reg[12]/NET0131 ,
		_w930_,
		_w3837_
	);
	LUT4 #(
		.INIT('ha8ab)
	) name2909 (
		\sub1_data_reg_reg[12]/NET0131 ,
		_w996_,
		_w2776_,
		_w3837_,
		_w3838_
	);
	LUT4 #(
		.INIT('h404c)
	) name2910 (
		\mix1_data_o_reg_reg[12]/NET0131 ,
		_w2774_,
		_w2775_,
		_w3838_,
		_w3839_
	);
	LUT4 #(
		.INIT('h0545)
	) name2911 (
		\sub1_data_reg_reg[12]/NET0131 ,
		\sub1_ready_o_reg/NET0131 ,
		_w1054_,
		_w2230_,
		_w3840_
	);
	LUT4 #(
		.INIT('h1510)
	) name2912 (
		\state_reg/NET0131 ,
		\sub1_data_reg_reg[12]/NET0131 ,
		_w996_,
		_w3837_,
		_w3841_
	);
	LUT4 #(
		.INIT('h0057)
	) name2913 (
		\state_reg/NET0131 ,
		_w3839_,
		_w3840_,
		_w3841_,
		_w3842_
	);
	LUT3 #(
		.INIT('h48)
	) name2914 (
		\key_i[12]_pad ,
		_w931_,
		_w3842_,
		_w3843_
	);
	LUT4 #(
		.INIT('h3222)
	) name2915 (
		\data_o[12]_pad ,
		_w931_,
		_w934_,
		_w2784_,
		_w3844_
	);
	LUT4 #(
		.INIT('h7b00)
	) name2916 (
		\ks1_key_reg_reg[12]/NET0131 ,
		_w2785_,
		_w3842_,
		_w3844_,
		_w3845_
	);
	LUT2 #(
		.INIT('he)
	) name2917 (
		_w3843_,
		_w3845_,
		_w3846_
	);
	LUT4 #(
		.INIT('haab8)
	) name2918 (
		\data_i[50]_pad ,
		decrypt_i_pad,
		\mix1_data_o_reg_reg[50]/NET0131 ,
		_w930_,
		_w3847_
	);
	LUT4 #(
		.INIT('haba8)
	) name2919 (
		\sub1_data_reg_reg[50]/NET0131 ,
		_w996_,
		_w2776_,
		_w3847_,
		_w3848_
	);
	LUT4 #(
		.INIT('h404c)
	) name2920 (
		\mix1_data_o_reg_reg[50]/NET0131 ,
		_w2774_,
		_w2775_,
		_w3848_,
		_w3849_
	);
	LUT4 #(
		.INIT('h0545)
	) name2921 (
		\sub1_data_reg_reg[50]/NET0131 ,
		\sub1_ready_o_reg/NET0131 ,
		_w1054_,
		_w2230_,
		_w3850_
	);
	LUT4 #(
		.INIT('h1015)
	) name2922 (
		\state_reg/NET0131 ,
		\sub1_data_reg_reg[50]/NET0131 ,
		_w996_,
		_w3847_,
		_w3851_
	);
	LUT4 #(
		.INIT('h0057)
	) name2923 (
		\state_reg/NET0131 ,
		_w3849_,
		_w3850_,
		_w3851_,
		_w3852_
	);
	LUT3 #(
		.INIT('h48)
	) name2924 (
		\key_i[50]_pad ,
		_w931_,
		_w3852_,
		_w3853_
	);
	LUT4 #(
		.INIT('h3222)
	) name2925 (
		\data_o[50]_pad ,
		_w931_,
		_w934_,
		_w2784_,
		_w3854_
	);
	LUT4 #(
		.INIT('h7b00)
	) name2926 (
		\ks1_key_reg_reg[50]/NET0131 ,
		_w2785_,
		_w3852_,
		_w3854_,
		_w3855_
	);
	LUT2 #(
		.INIT('he)
	) name2927 (
		_w3853_,
		_w3855_,
		_w3856_
	);
	LUT4 #(
		.INIT('h5547)
	) name2928 (
		\data_i[10]_pad ,
		decrypt_i_pad,
		\mix1_data_o_reg_reg[10]/NET0131 ,
		_w930_,
		_w3857_
	);
	LUT4 #(
		.INIT('ha8ab)
	) name2929 (
		\sub1_data_reg_reg[10]/NET0131 ,
		_w996_,
		_w2776_,
		_w3857_,
		_w3858_
	);
	LUT4 #(
		.INIT('h404c)
	) name2930 (
		\mix1_data_o_reg_reg[10]/NET0131 ,
		_w2774_,
		_w2775_,
		_w3858_,
		_w3859_
	);
	LUT4 #(
		.INIT('h0545)
	) name2931 (
		\sub1_data_reg_reg[10]/NET0131 ,
		\sub1_ready_o_reg/NET0131 ,
		_w1054_,
		_w2230_,
		_w3860_
	);
	LUT4 #(
		.INIT('h1510)
	) name2932 (
		\state_reg/NET0131 ,
		\sub1_data_reg_reg[10]/NET0131 ,
		_w996_,
		_w3857_,
		_w3861_
	);
	LUT4 #(
		.INIT('h0057)
	) name2933 (
		\state_reg/NET0131 ,
		_w3859_,
		_w3860_,
		_w3861_,
		_w3862_
	);
	LUT3 #(
		.INIT('h48)
	) name2934 (
		\key_i[10]_pad ,
		_w931_,
		_w3862_,
		_w3863_
	);
	LUT4 #(
		.INIT('h3222)
	) name2935 (
		\data_o[10]_pad ,
		_w931_,
		_w934_,
		_w2784_,
		_w3864_
	);
	LUT4 #(
		.INIT('h7b00)
	) name2936 (
		\ks1_key_reg_reg[10]/NET0131 ,
		_w2785_,
		_w3862_,
		_w3864_,
		_w3865_
	);
	LUT2 #(
		.INIT('he)
	) name2937 (
		_w3863_,
		_w3865_,
		_w3866_
	);
	LUT4 #(
		.INIT('h5547)
	) name2938 (
		\data_i[13]_pad ,
		decrypt_i_pad,
		\mix1_data_o_reg_reg[13]/NET0131 ,
		_w930_,
		_w3867_
	);
	LUT4 #(
		.INIT('ha8ab)
	) name2939 (
		\sub1_data_reg_reg[13]/NET0131 ,
		_w996_,
		_w2776_,
		_w3867_,
		_w3868_
	);
	LUT4 #(
		.INIT('h404c)
	) name2940 (
		\mix1_data_o_reg_reg[13]/NET0131 ,
		_w2774_,
		_w2775_,
		_w3868_,
		_w3869_
	);
	LUT4 #(
		.INIT('h0545)
	) name2941 (
		\sub1_data_reg_reg[13]/NET0131 ,
		\sub1_ready_o_reg/NET0131 ,
		_w1054_,
		_w2230_,
		_w3870_
	);
	LUT4 #(
		.INIT('h1510)
	) name2942 (
		\state_reg/NET0131 ,
		\sub1_data_reg_reg[13]/NET0131 ,
		_w996_,
		_w3867_,
		_w3871_
	);
	LUT4 #(
		.INIT('h0057)
	) name2943 (
		\state_reg/NET0131 ,
		_w3869_,
		_w3870_,
		_w3871_,
		_w3872_
	);
	LUT3 #(
		.INIT('h48)
	) name2944 (
		\key_i[13]_pad ,
		_w931_,
		_w3872_,
		_w3873_
	);
	LUT4 #(
		.INIT('h3222)
	) name2945 (
		\data_o[13]_pad ,
		_w931_,
		_w934_,
		_w2784_,
		_w3874_
	);
	LUT4 #(
		.INIT('h7b00)
	) name2946 (
		\ks1_key_reg_reg[13]/NET0131 ,
		_w2785_,
		_w3872_,
		_w3874_,
		_w3875_
	);
	LUT2 #(
		.INIT('he)
	) name2947 (
		_w3873_,
		_w3875_,
		_w3876_
	);
	LUT4 #(
		.INIT('haab8)
	) name2948 (
		\data_i[51]_pad ,
		decrypt_i_pad,
		\mix1_data_o_reg_reg[51]/NET0131 ,
		_w930_,
		_w3877_
	);
	LUT4 #(
		.INIT('haba8)
	) name2949 (
		\sub1_data_reg_reg[51]/NET0131 ,
		_w996_,
		_w2776_,
		_w3877_,
		_w3878_
	);
	LUT4 #(
		.INIT('h404c)
	) name2950 (
		\mix1_data_o_reg_reg[51]/NET0131 ,
		_w2774_,
		_w2775_,
		_w3878_,
		_w3879_
	);
	LUT4 #(
		.INIT('h0545)
	) name2951 (
		\sub1_data_reg_reg[51]/NET0131 ,
		\sub1_ready_o_reg/NET0131 ,
		_w1054_,
		_w2230_,
		_w3880_
	);
	LUT4 #(
		.INIT('h1015)
	) name2952 (
		\state_reg/NET0131 ,
		\sub1_data_reg_reg[51]/NET0131 ,
		_w996_,
		_w3877_,
		_w3881_
	);
	LUT4 #(
		.INIT('h0057)
	) name2953 (
		\state_reg/NET0131 ,
		_w3879_,
		_w3880_,
		_w3881_,
		_w3882_
	);
	LUT3 #(
		.INIT('h48)
	) name2954 (
		\key_i[51]_pad ,
		_w931_,
		_w3882_,
		_w3883_
	);
	LUT4 #(
		.INIT('h3222)
	) name2955 (
		\data_o[51]_pad ,
		_w931_,
		_w934_,
		_w2784_,
		_w3884_
	);
	LUT4 #(
		.INIT('h7b00)
	) name2956 (
		\ks1_key_reg_reg[51]/NET0131 ,
		_w2785_,
		_w3882_,
		_w3884_,
		_w3885_
	);
	LUT2 #(
		.INIT('he)
	) name2957 (
		_w3883_,
		_w3885_,
		_w3886_
	);
	LUT4 #(
		.INIT('haab8)
	) name2958 (
		\data_i[52]_pad ,
		decrypt_i_pad,
		\mix1_data_o_reg_reg[52]/NET0131 ,
		_w930_,
		_w3887_
	);
	LUT4 #(
		.INIT('haba8)
	) name2959 (
		\sub1_data_reg_reg[52]/NET0131 ,
		_w996_,
		_w2776_,
		_w3887_,
		_w3888_
	);
	LUT4 #(
		.INIT('h404c)
	) name2960 (
		\mix1_data_o_reg_reg[52]/NET0131 ,
		_w2774_,
		_w2775_,
		_w3888_,
		_w3889_
	);
	LUT4 #(
		.INIT('h0545)
	) name2961 (
		\sub1_data_reg_reg[52]/NET0131 ,
		\sub1_ready_o_reg/NET0131 ,
		_w1054_,
		_w2230_,
		_w3890_
	);
	LUT4 #(
		.INIT('h1015)
	) name2962 (
		\state_reg/NET0131 ,
		\sub1_data_reg_reg[52]/NET0131 ,
		_w996_,
		_w3887_,
		_w3891_
	);
	LUT4 #(
		.INIT('h0057)
	) name2963 (
		\state_reg/NET0131 ,
		_w3889_,
		_w3890_,
		_w3891_,
		_w3892_
	);
	LUT3 #(
		.INIT('h48)
	) name2964 (
		\key_i[52]_pad ,
		_w931_,
		_w3892_,
		_w3893_
	);
	LUT4 #(
		.INIT('h3222)
	) name2965 (
		\data_o[52]_pad ,
		_w931_,
		_w934_,
		_w2784_,
		_w3894_
	);
	LUT4 #(
		.INIT('h7b00)
	) name2966 (
		\ks1_key_reg_reg[52]/NET0131 ,
		_w2785_,
		_w3892_,
		_w3894_,
		_w3895_
	);
	LUT2 #(
		.INIT('he)
	) name2967 (
		_w3893_,
		_w3895_,
		_w3896_
	);
	LUT4 #(
		.INIT('haab8)
	) name2968 (
		\data_i[53]_pad ,
		decrypt_i_pad,
		\mix1_data_o_reg_reg[53]/NET0131 ,
		_w930_,
		_w3897_
	);
	LUT4 #(
		.INIT('haba8)
	) name2969 (
		\sub1_data_reg_reg[53]/NET0131 ,
		_w996_,
		_w2776_,
		_w3897_,
		_w3898_
	);
	LUT4 #(
		.INIT('h404c)
	) name2970 (
		\mix1_data_o_reg_reg[53]/NET0131 ,
		_w2774_,
		_w2775_,
		_w3898_,
		_w3899_
	);
	LUT4 #(
		.INIT('h0545)
	) name2971 (
		\sub1_data_reg_reg[53]/NET0131 ,
		\sub1_ready_o_reg/NET0131 ,
		_w1054_,
		_w2230_,
		_w3900_
	);
	LUT4 #(
		.INIT('h1015)
	) name2972 (
		\state_reg/NET0131 ,
		\sub1_data_reg_reg[53]/NET0131 ,
		_w996_,
		_w3897_,
		_w3901_
	);
	LUT4 #(
		.INIT('h0057)
	) name2973 (
		\state_reg/NET0131 ,
		_w3899_,
		_w3900_,
		_w3901_,
		_w3902_
	);
	LUT3 #(
		.INIT('h48)
	) name2974 (
		\key_i[53]_pad ,
		_w931_,
		_w3902_,
		_w3903_
	);
	LUT4 #(
		.INIT('h3222)
	) name2975 (
		\data_o[53]_pad ,
		_w931_,
		_w934_,
		_w2784_,
		_w3904_
	);
	LUT4 #(
		.INIT('h7b00)
	) name2976 (
		\ks1_key_reg_reg[53]/NET0131 ,
		_w2785_,
		_w3902_,
		_w3904_,
		_w3905_
	);
	LUT2 #(
		.INIT('he)
	) name2977 (
		_w3903_,
		_w3905_,
		_w3906_
	);
	LUT4 #(
		.INIT('h5547)
	) name2978 (
		\data_i[14]_pad ,
		decrypt_i_pad,
		\mix1_data_o_reg_reg[14]/NET0131 ,
		_w930_,
		_w3907_
	);
	LUT4 #(
		.INIT('ha8ab)
	) name2979 (
		\sub1_data_reg_reg[14]/NET0131 ,
		_w996_,
		_w2776_,
		_w3907_,
		_w3908_
	);
	LUT4 #(
		.INIT('h404c)
	) name2980 (
		\mix1_data_o_reg_reg[14]/NET0131 ,
		_w2774_,
		_w2775_,
		_w3908_,
		_w3909_
	);
	LUT4 #(
		.INIT('h0545)
	) name2981 (
		\sub1_data_reg_reg[14]/NET0131 ,
		\sub1_ready_o_reg/NET0131 ,
		_w1054_,
		_w2230_,
		_w3910_
	);
	LUT4 #(
		.INIT('h1510)
	) name2982 (
		\state_reg/NET0131 ,
		\sub1_data_reg_reg[14]/NET0131 ,
		_w996_,
		_w3907_,
		_w3911_
	);
	LUT4 #(
		.INIT('h0057)
	) name2983 (
		\state_reg/NET0131 ,
		_w3909_,
		_w3910_,
		_w3911_,
		_w3912_
	);
	LUT3 #(
		.INIT('h48)
	) name2984 (
		\key_i[14]_pad ,
		_w931_,
		_w3912_,
		_w3913_
	);
	LUT4 #(
		.INIT('h3222)
	) name2985 (
		\data_o[14]_pad ,
		_w931_,
		_w934_,
		_w2784_,
		_w3914_
	);
	LUT4 #(
		.INIT('h7b00)
	) name2986 (
		\ks1_key_reg_reg[14]/NET0131 ,
		_w2785_,
		_w3912_,
		_w3914_,
		_w3915_
	);
	LUT2 #(
		.INIT('he)
	) name2987 (
		_w3913_,
		_w3915_,
		_w3916_
	);
	LUT4 #(
		.INIT('haab8)
	) name2988 (
		\data_i[100]_pad ,
		decrypt_i_pad,
		\mix1_data_o_reg_reg[100]/NET0131 ,
		_w930_,
		_w3917_
	);
	LUT4 #(
		.INIT('haba8)
	) name2989 (
		\sub1_data_reg_reg[100]/NET0131 ,
		_w996_,
		_w2776_,
		_w3917_,
		_w3918_
	);
	LUT4 #(
		.INIT('h404c)
	) name2990 (
		\mix1_data_o_reg_reg[100]/NET0131 ,
		_w2774_,
		_w2775_,
		_w3918_,
		_w3919_
	);
	LUT4 #(
		.INIT('h0545)
	) name2991 (
		\sub1_data_reg_reg[100]/NET0131 ,
		\sub1_ready_o_reg/NET0131 ,
		_w1054_,
		_w2230_,
		_w3920_
	);
	LUT4 #(
		.INIT('h1015)
	) name2992 (
		\state_reg/NET0131 ,
		\sub1_data_reg_reg[100]/NET0131 ,
		_w996_,
		_w3917_,
		_w3921_
	);
	LUT4 #(
		.INIT('h0057)
	) name2993 (
		\state_reg/NET0131 ,
		_w3919_,
		_w3920_,
		_w3921_,
		_w3922_
	);
	LUT3 #(
		.INIT('h48)
	) name2994 (
		\key_i[100]_pad ,
		_w931_,
		_w3922_,
		_w3923_
	);
	LUT4 #(
		.INIT('h3222)
	) name2995 (
		\data_o[100]_pad ,
		_w931_,
		_w934_,
		_w2784_,
		_w3924_
	);
	LUT4 #(
		.INIT('h7b00)
	) name2996 (
		\ks1_key_reg_reg[100]/NET0131 ,
		_w2785_,
		_w3922_,
		_w3924_,
		_w3925_
	);
	LUT2 #(
		.INIT('he)
	) name2997 (
		_w3923_,
		_w3925_,
		_w3926_
	);
	LUT4 #(
		.INIT('haab8)
	) name2998 (
		\data_i[54]_pad ,
		decrypt_i_pad,
		\mix1_data_o_reg_reg[54]/NET0131 ,
		_w930_,
		_w3927_
	);
	LUT4 #(
		.INIT('haba8)
	) name2999 (
		\sub1_data_reg_reg[54]/NET0131 ,
		_w996_,
		_w2776_,
		_w3927_,
		_w3928_
	);
	LUT4 #(
		.INIT('h404c)
	) name3000 (
		\mix1_data_o_reg_reg[54]/NET0131 ,
		_w2774_,
		_w2775_,
		_w3928_,
		_w3929_
	);
	LUT4 #(
		.INIT('h0545)
	) name3001 (
		\sub1_data_reg_reg[54]/NET0131 ,
		\sub1_ready_o_reg/NET0131 ,
		_w1054_,
		_w2230_,
		_w3930_
	);
	LUT4 #(
		.INIT('h1015)
	) name3002 (
		\state_reg/NET0131 ,
		\sub1_data_reg_reg[54]/NET0131 ,
		_w996_,
		_w3927_,
		_w3931_
	);
	LUT4 #(
		.INIT('h0057)
	) name3003 (
		\state_reg/NET0131 ,
		_w3929_,
		_w3930_,
		_w3931_,
		_w3932_
	);
	LUT3 #(
		.INIT('h48)
	) name3004 (
		\key_i[54]_pad ,
		_w931_,
		_w3932_,
		_w3933_
	);
	LUT4 #(
		.INIT('h3222)
	) name3005 (
		\data_o[54]_pad ,
		_w931_,
		_w934_,
		_w2784_,
		_w3934_
	);
	LUT4 #(
		.INIT('h7b00)
	) name3006 (
		\ks1_key_reg_reg[54]/NET0131 ,
		_w2785_,
		_w3932_,
		_w3934_,
		_w3935_
	);
	LUT2 #(
		.INIT('he)
	) name3007 (
		_w3933_,
		_w3935_,
		_w3936_
	);
	LUT4 #(
		.INIT('haab8)
	) name3008 (
		\data_i[55]_pad ,
		decrypt_i_pad,
		\mix1_data_o_reg_reg[55]/NET0131 ,
		_w930_,
		_w3937_
	);
	LUT4 #(
		.INIT('haba8)
	) name3009 (
		\sub1_data_reg_reg[55]/NET0131 ,
		_w996_,
		_w2776_,
		_w3937_,
		_w3938_
	);
	LUT4 #(
		.INIT('h404c)
	) name3010 (
		\mix1_data_o_reg_reg[55]/NET0131 ,
		_w2774_,
		_w2775_,
		_w3938_,
		_w3939_
	);
	LUT4 #(
		.INIT('h0545)
	) name3011 (
		\sub1_data_reg_reg[55]/NET0131 ,
		\sub1_ready_o_reg/NET0131 ,
		_w1054_,
		_w2230_,
		_w3940_
	);
	LUT4 #(
		.INIT('h1015)
	) name3012 (
		\state_reg/NET0131 ,
		\sub1_data_reg_reg[55]/NET0131 ,
		_w996_,
		_w3937_,
		_w3941_
	);
	LUT4 #(
		.INIT('h0057)
	) name3013 (
		\state_reg/NET0131 ,
		_w3939_,
		_w3940_,
		_w3941_,
		_w3942_
	);
	LUT3 #(
		.INIT('h48)
	) name3014 (
		\key_i[55]_pad ,
		_w931_,
		_w3942_,
		_w3943_
	);
	LUT4 #(
		.INIT('h3222)
	) name3015 (
		\data_o[55]_pad ,
		_w931_,
		_w934_,
		_w2784_,
		_w3944_
	);
	LUT4 #(
		.INIT('h7b00)
	) name3016 (
		\ks1_key_reg_reg[55]/NET0131 ,
		_w2785_,
		_w3942_,
		_w3944_,
		_w3945_
	);
	LUT2 #(
		.INIT('he)
	) name3017 (
		_w3943_,
		_w3945_,
		_w3946_
	);
	LUT4 #(
		.INIT('h5547)
	) name3018 (
		\data_i[15]_pad ,
		decrypt_i_pad,
		\mix1_data_o_reg_reg[15]/NET0131 ,
		_w930_,
		_w3947_
	);
	LUT4 #(
		.INIT('ha8ab)
	) name3019 (
		\sub1_data_reg_reg[15]/NET0131 ,
		_w996_,
		_w2776_,
		_w3947_,
		_w3948_
	);
	LUT4 #(
		.INIT('h404c)
	) name3020 (
		\mix1_data_o_reg_reg[15]/NET0131 ,
		_w2774_,
		_w2775_,
		_w3948_,
		_w3949_
	);
	LUT4 #(
		.INIT('h0545)
	) name3021 (
		\sub1_data_reg_reg[15]/NET0131 ,
		\sub1_ready_o_reg/NET0131 ,
		_w1054_,
		_w2230_,
		_w3950_
	);
	LUT4 #(
		.INIT('h1510)
	) name3022 (
		\state_reg/NET0131 ,
		\sub1_data_reg_reg[15]/NET0131 ,
		_w996_,
		_w3947_,
		_w3951_
	);
	LUT4 #(
		.INIT('h0057)
	) name3023 (
		\state_reg/NET0131 ,
		_w3949_,
		_w3950_,
		_w3951_,
		_w3952_
	);
	LUT3 #(
		.INIT('h48)
	) name3024 (
		\key_i[15]_pad ,
		_w931_,
		_w3952_,
		_w3953_
	);
	LUT4 #(
		.INIT('h3222)
	) name3025 (
		\data_o[15]_pad ,
		_w931_,
		_w934_,
		_w2784_,
		_w3954_
	);
	LUT4 #(
		.INIT('h7b00)
	) name3026 (
		\ks1_key_reg_reg[15]/NET0131 ,
		_w2785_,
		_w3952_,
		_w3954_,
		_w3955_
	);
	LUT2 #(
		.INIT('he)
	) name3027 (
		_w3953_,
		_w3955_,
		_w3956_
	);
	LUT4 #(
		.INIT('h5547)
	) name3028 (
		\data_i[110]_pad ,
		decrypt_i_pad,
		\mix1_data_o_reg_reg[110]/NET0131 ,
		_w930_,
		_w3957_
	);
	LUT4 #(
		.INIT('ha8ab)
	) name3029 (
		\sub1_data_reg_reg[110]/NET0131 ,
		_w996_,
		_w2776_,
		_w3957_,
		_w3958_
	);
	LUT4 #(
		.INIT('h404c)
	) name3030 (
		\mix1_data_o_reg_reg[110]/NET0131 ,
		_w2774_,
		_w2775_,
		_w3958_,
		_w3959_
	);
	LUT4 #(
		.INIT('h0545)
	) name3031 (
		\sub1_data_reg_reg[110]/NET0131 ,
		\sub1_ready_o_reg/NET0131 ,
		_w1054_,
		_w2230_,
		_w3960_
	);
	LUT4 #(
		.INIT('h1510)
	) name3032 (
		\state_reg/NET0131 ,
		\sub1_data_reg_reg[110]/NET0131 ,
		_w996_,
		_w3957_,
		_w3961_
	);
	LUT4 #(
		.INIT('h0057)
	) name3033 (
		\state_reg/NET0131 ,
		_w3959_,
		_w3960_,
		_w3961_,
		_w3962_
	);
	LUT3 #(
		.INIT('h48)
	) name3034 (
		\key_i[110]_pad ,
		_w931_,
		_w3962_,
		_w3963_
	);
	LUT4 #(
		.INIT('h3222)
	) name3035 (
		\data_o[110]_pad ,
		_w931_,
		_w934_,
		_w2784_,
		_w3964_
	);
	LUT4 #(
		.INIT('h7b00)
	) name3036 (
		\ks1_key_reg_reg[110]/P0002 ,
		_w2785_,
		_w3962_,
		_w3964_,
		_w3965_
	);
	LUT2 #(
		.INIT('he)
	) name3037 (
		_w3963_,
		_w3965_,
		_w3966_
	);
	LUT4 #(
		.INIT('h5547)
	) name3038 (
		\data_i[56]_pad ,
		decrypt_i_pad,
		\mix1_data_o_reg_reg[56]/NET0131 ,
		_w930_,
		_w3967_
	);
	LUT4 #(
		.INIT('ha8ab)
	) name3039 (
		\sub1_data_reg_reg[56]/NET0131 ,
		_w996_,
		_w2776_,
		_w3967_,
		_w3968_
	);
	LUT4 #(
		.INIT('h404c)
	) name3040 (
		\mix1_data_o_reg_reg[56]/NET0131 ,
		_w2774_,
		_w2775_,
		_w3968_,
		_w3969_
	);
	LUT4 #(
		.INIT('h0545)
	) name3041 (
		\sub1_data_reg_reg[56]/NET0131 ,
		\sub1_ready_o_reg/NET0131 ,
		_w1054_,
		_w2230_,
		_w3970_
	);
	LUT4 #(
		.INIT('h1510)
	) name3042 (
		\state_reg/NET0131 ,
		\sub1_data_reg_reg[56]/NET0131 ,
		_w996_,
		_w3967_,
		_w3971_
	);
	LUT4 #(
		.INIT('h0057)
	) name3043 (
		\state_reg/NET0131 ,
		_w3969_,
		_w3970_,
		_w3971_,
		_w3972_
	);
	LUT3 #(
		.INIT('h48)
	) name3044 (
		\key_i[56]_pad ,
		_w931_,
		_w3972_,
		_w3973_
	);
	LUT4 #(
		.INIT('h3222)
	) name3045 (
		\data_o[56]_pad ,
		_w931_,
		_w934_,
		_w2784_,
		_w3974_
	);
	LUT4 #(
		.INIT('h7b00)
	) name3046 (
		\ks1_key_reg_reg[56]/NET0131 ,
		_w2785_,
		_w3972_,
		_w3974_,
		_w3975_
	);
	LUT2 #(
		.INIT('he)
	) name3047 (
		_w3973_,
		_w3975_,
		_w3976_
	);
	LUT4 #(
		.INIT('h5547)
	) name3048 (
		\data_i[57]_pad ,
		decrypt_i_pad,
		\mix1_data_o_reg_reg[57]/NET0131 ,
		_w930_,
		_w3977_
	);
	LUT4 #(
		.INIT('ha8ab)
	) name3049 (
		\sub1_data_reg_reg[57]/NET0131 ,
		_w996_,
		_w2776_,
		_w3977_,
		_w3978_
	);
	LUT4 #(
		.INIT('h404c)
	) name3050 (
		\mix1_data_o_reg_reg[57]/NET0131 ,
		_w2774_,
		_w2775_,
		_w3978_,
		_w3979_
	);
	LUT4 #(
		.INIT('h0545)
	) name3051 (
		\sub1_data_reg_reg[57]/NET0131 ,
		\sub1_ready_o_reg/NET0131 ,
		_w1054_,
		_w2230_,
		_w3980_
	);
	LUT4 #(
		.INIT('h1510)
	) name3052 (
		\state_reg/NET0131 ,
		\sub1_data_reg_reg[57]/NET0131 ,
		_w996_,
		_w3977_,
		_w3981_
	);
	LUT4 #(
		.INIT('h0057)
	) name3053 (
		\state_reg/NET0131 ,
		_w3979_,
		_w3980_,
		_w3981_,
		_w3982_
	);
	LUT3 #(
		.INIT('h48)
	) name3054 (
		\key_i[57]_pad ,
		_w931_,
		_w3982_,
		_w3983_
	);
	LUT4 #(
		.INIT('h3222)
	) name3055 (
		\data_o[57]_pad ,
		_w931_,
		_w934_,
		_w2784_,
		_w3984_
	);
	LUT4 #(
		.INIT('h7b00)
	) name3056 (
		\ks1_key_reg_reg[57]/NET0131 ,
		_w2785_,
		_w3982_,
		_w3984_,
		_w3985_
	);
	LUT2 #(
		.INIT('he)
	) name3057 (
		_w3983_,
		_w3985_,
		_w3986_
	);
	LUT4 #(
		.INIT('haab8)
	) name3058 (
		\data_i[16]_pad ,
		decrypt_i_pad,
		\mix1_data_o_reg_reg[16]/NET0131 ,
		_w930_,
		_w3987_
	);
	LUT4 #(
		.INIT('haba8)
	) name3059 (
		\sub1_data_reg_reg[16]/NET0131 ,
		_w996_,
		_w2776_,
		_w3987_,
		_w3988_
	);
	LUT4 #(
		.INIT('h404c)
	) name3060 (
		\mix1_data_o_reg_reg[16]/NET0131 ,
		_w2774_,
		_w2775_,
		_w3988_,
		_w3989_
	);
	LUT4 #(
		.INIT('h0545)
	) name3061 (
		\sub1_data_reg_reg[16]/NET0131 ,
		\sub1_ready_o_reg/NET0131 ,
		_w1054_,
		_w2230_,
		_w3990_
	);
	LUT4 #(
		.INIT('h1015)
	) name3062 (
		\state_reg/NET0131 ,
		\sub1_data_reg_reg[16]/NET0131 ,
		_w996_,
		_w3987_,
		_w3991_
	);
	LUT4 #(
		.INIT('h0057)
	) name3063 (
		\state_reg/NET0131 ,
		_w3989_,
		_w3990_,
		_w3991_,
		_w3992_
	);
	LUT3 #(
		.INIT('h48)
	) name3064 (
		\key_i[16]_pad ,
		_w931_,
		_w3992_,
		_w3993_
	);
	LUT4 #(
		.INIT('h3222)
	) name3065 (
		\data_o[16]_pad ,
		_w931_,
		_w934_,
		_w2784_,
		_w3994_
	);
	LUT4 #(
		.INIT('h7b00)
	) name3066 (
		\ks1_key_reg_reg[16]/NET0131 ,
		_w2785_,
		_w3992_,
		_w3994_,
		_w3995_
	);
	LUT2 #(
		.INIT('he)
	) name3067 (
		_w3993_,
		_w3995_,
		_w3996_
	);
	LUT4 #(
		.INIT('h5547)
	) name3068 (
		\data_i[58]_pad ,
		decrypt_i_pad,
		\mix1_data_o_reg_reg[58]/NET0131 ,
		_w930_,
		_w3997_
	);
	LUT4 #(
		.INIT('ha8ab)
	) name3069 (
		\sub1_data_reg_reg[58]/NET0131 ,
		_w996_,
		_w2776_,
		_w3997_,
		_w3998_
	);
	LUT4 #(
		.INIT('h404c)
	) name3070 (
		\mix1_data_o_reg_reg[58]/NET0131 ,
		_w2774_,
		_w2775_,
		_w3998_,
		_w3999_
	);
	LUT4 #(
		.INIT('h0545)
	) name3071 (
		\sub1_data_reg_reg[58]/NET0131 ,
		\sub1_ready_o_reg/NET0131 ,
		_w1054_,
		_w2230_,
		_w4000_
	);
	LUT4 #(
		.INIT('h1510)
	) name3072 (
		\state_reg/NET0131 ,
		\sub1_data_reg_reg[58]/NET0131 ,
		_w996_,
		_w3997_,
		_w4001_
	);
	LUT4 #(
		.INIT('h0057)
	) name3073 (
		\state_reg/NET0131 ,
		_w3999_,
		_w4000_,
		_w4001_,
		_w4002_
	);
	LUT3 #(
		.INIT('h48)
	) name3074 (
		\key_i[58]_pad ,
		_w931_,
		_w4002_,
		_w4003_
	);
	LUT4 #(
		.INIT('h3222)
	) name3075 (
		\data_o[58]_pad ,
		_w931_,
		_w934_,
		_w2784_,
		_w4004_
	);
	LUT4 #(
		.INIT('h7b00)
	) name3076 (
		\ks1_key_reg_reg[58]/NET0131 ,
		_w2785_,
		_w4002_,
		_w4004_,
		_w4005_
	);
	LUT2 #(
		.INIT('he)
	) name3077 (
		_w4003_,
		_w4005_,
		_w4006_
	);
	LUT4 #(
		.INIT('h5547)
	) name3078 (
		\data_i[59]_pad ,
		decrypt_i_pad,
		\mix1_data_o_reg_reg[59]/NET0131 ,
		_w930_,
		_w4007_
	);
	LUT4 #(
		.INIT('ha8ab)
	) name3079 (
		\sub1_data_reg_reg[59]/NET0131 ,
		_w996_,
		_w2776_,
		_w4007_,
		_w4008_
	);
	LUT4 #(
		.INIT('h404c)
	) name3080 (
		\mix1_data_o_reg_reg[59]/NET0131 ,
		_w2774_,
		_w2775_,
		_w4008_,
		_w4009_
	);
	LUT4 #(
		.INIT('h0545)
	) name3081 (
		\sub1_data_reg_reg[59]/NET0131 ,
		\sub1_ready_o_reg/NET0131 ,
		_w1054_,
		_w2230_,
		_w4010_
	);
	LUT4 #(
		.INIT('h1510)
	) name3082 (
		\state_reg/NET0131 ,
		\sub1_data_reg_reg[59]/NET0131 ,
		_w996_,
		_w4007_,
		_w4011_
	);
	LUT4 #(
		.INIT('h0057)
	) name3083 (
		\state_reg/NET0131 ,
		_w4009_,
		_w4010_,
		_w4011_,
		_w4012_
	);
	LUT3 #(
		.INIT('h48)
	) name3084 (
		\key_i[59]_pad ,
		_w931_,
		_w4012_,
		_w4013_
	);
	LUT4 #(
		.INIT('h3222)
	) name3085 (
		\data_o[59]_pad ,
		_w931_,
		_w934_,
		_w2784_,
		_w4014_
	);
	LUT4 #(
		.INIT('h7b00)
	) name3086 (
		\ks1_key_reg_reg[59]/NET0131 ,
		_w2785_,
		_w4012_,
		_w4014_,
		_w4015_
	);
	LUT2 #(
		.INIT('he)
	) name3087 (
		_w4013_,
		_w4015_,
		_w4016_
	);
	LUT4 #(
		.INIT('h5547)
	) name3088 (
		\data_i[111]_pad ,
		decrypt_i_pad,
		\mix1_data_o_reg_reg[111]/NET0131 ,
		_w930_,
		_w4017_
	);
	LUT4 #(
		.INIT('ha8ab)
	) name3089 (
		\sub1_data_reg_reg[111]/NET0131 ,
		_w996_,
		_w2776_,
		_w4017_,
		_w4018_
	);
	LUT4 #(
		.INIT('h404c)
	) name3090 (
		\mix1_data_o_reg_reg[111]/NET0131 ,
		_w2774_,
		_w2775_,
		_w4018_,
		_w4019_
	);
	LUT4 #(
		.INIT('h0545)
	) name3091 (
		\sub1_data_reg_reg[111]/NET0131 ,
		\sub1_ready_o_reg/NET0131 ,
		_w1054_,
		_w2230_,
		_w4020_
	);
	LUT4 #(
		.INIT('h1510)
	) name3092 (
		\state_reg/NET0131 ,
		\sub1_data_reg_reg[111]/NET0131 ,
		_w996_,
		_w4017_,
		_w4021_
	);
	LUT4 #(
		.INIT('h0057)
	) name3093 (
		\state_reg/NET0131 ,
		_w4019_,
		_w4020_,
		_w4021_,
		_w4022_
	);
	LUT3 #(
		.INIT('h48)
	) name3094 (
		\key_i[111]_pad ,
		_w931_,
		_w4022_,
		_w4023_
	);
	LUT4 #(
		.INIT('h3222)
	) name3095 (
		\data_o[111]_pad ,
		_w931_,
		_w934_,
		_w2784_,
		_w4024_
	);
	LUT4 #(
		.INIT('h7b00)
	) name3096 (
		\ks1_key_reg_reg[111]/NET0131 ,
		_w2785_,
		_w4022_,
		_w4024_,
		_w4025_
	);
	LUT2 #(
		.INIT('he)
	) name3097 (
		_w4023_,
		_w4025_,
		_w4026_
	);
	LUT4 #(
		.INIT('haab8)
	) name3098 (
		\data_i[17]_pad ,
		decrypt_i_pad,
		\mix1_data_o_reg_reg[17]/NET0131 ,
		_w930_,
		_w4027_
	);
	LUT4 #(
		.INIT('haba8)
	) name3099 (
		\sub1_data_reg_reg[17]/NET0131 ,
		_w996_,
		_w2776_,
		_w4027_,
		_w4028_
	);
	LUT4 #(
		.INIT('h404c)
	) name3100 (
		\mix1_data_o_reg_reg[17]/NET0131 ,
		_w2774_,
		_w2775_,
		_w4028_,
		_w4029_
	);
	LUT4 #(
		.INIT('h0545)
	) name3101 (
		\sub1_data_reg_reg[17]/NET0131 ,
		\sub1_ready_o_reg/NET0131 ,
		_w1054_,
		_w2230_,
		_w4030_
	);
	LUT4 #(
		.INIT('h1015)
	) name3102 (
		\state_reg/NET0131 ,
		\sub1_data_reg_reg[17]/NET0131 ,
		_w996_,
		_w4027_,
		_w4031_
	);
	LUT4 #(
		.INIT('h0057)
	) name3103 (
		\state_reg/NET0131 ,
		_w4029_,
		_w4030_,
		_w4031_,
		_w4032_
	);
	LUT3 #(
		.INIT('h48)
	) name3104 (
		\key_i[17]_pad ,
		_w931_,
		_w4032_,
		_w4033_
	);
	LUT4 #(
		.INIT('h3222)
	) name3105 (
		\data_o[17]_pad ,
		_w931_,
		_w934_,
		_w2784_,
		_w4034_
	);
	LUT4 #(
		.INIT('h7b00)
	) name3106 (
		\ks1_key_reg_reg[17]/NET0131 ,
		_w2785_,
		_w4032_,
		_w4034_,
		_w4035_
	);
	LUT2 #(
		.INIT('he)
	) name3107 (
		_w4033_,
		_w4035_,
		_w4036_
	);
	LUT4 #(
		.INIT('h5547)
	) name3108 (
		\data_i[5]_pad ,
		decrypt_i_pad,
		\mix1_data_o_reg_reg[5]/NET0131 ,
		_w930_,
		_w4037_
	);
	LUT4 #(
		.INIT('ha8ab)
	) name3109 (
		\sub1_data_reg_reg[5]/NET0131 ,
		_w996_,
		_w2776_,
		_w4037_,
		_w4038_
	);
	LUT4 #(
		.INIT('h404c)
	) name3110 (
		\mix1_data_o_reg_reg[5]/NET0131 ,
		_w2774_,
		_w2775_,
		_w4038_,
		_w4039_
	);
	LUT4 #(
		.INIT('h0545)
	) name3111 (
		\sub1_data_reg_reg[5]/NET0131 ,
		\sub1_ready_o_reg/NET0131 ,
		_w1054_,
		_w2230_,
		_w4040_
	);
	LUT4 #(
		.INIT('h1510)
	) name3112 (
		\state_reg/NET0131 ,
		\sub1_data_reg_reg[5]/NET0131 ,
		_w996_,
		_w4037_,
		_w4041_
	);
	LUT4 #(
		.INIT('h0057)
	) name3113 (
		\state_reg/NET0131 ,
		_w4039_,
		_w4040_,
		_w4041_,
		_w4042_
	);
	LUT3 #(
		.INIT('h48)
	) name3114 (
		\key_i[5]_pad ,
		_w931_,
		_w4042_,
		_w4043_
	);
	LUT4 #(
		.INIT('h3222)
	) name3115 (
		\data_o[5]_pad ,
		_w931_,
		_w934_,
		_w2784_,
		_w4044_
	);
	LUT4 #(
		.INIT('h7b00)
	) name3116 (
		\ks1_key_reg_reg[5]/NET0131 ,
		_w2785_,
		_w4042_,
		_w4044_,
		_w4045_
	);
	LUT2 #(
		.INIT('he)
	) name3117 (
		_w4043_,
		_w4045_,
		_w4046_
	);
	LUT4 #(
		.INIT('h5547)
	) name3118 (
		\data_i[60]_pad ,
		decrypt_i_pad,
		\mix1_data_o_reg_reg[60]/NET0131 ,
		_w930_,
		_w4047_
	);
	LUT4 #(
		.INIT('ha8ab)
	) name3119 (
		\sub1_data_reg_reg[60]/NET0131 ,
		_w996_,
		_w2776_,
		_w4047_,
		_w4048_
	);
	LUT4 #(
		.INIT('h404c)
	) name3120 (
		\mix1_data_o_reg_reg[60]/NET0131 ,
		_w2774_,
		_w2775_,
		_w4048_,
		_w4049_
	);
	LUT4 #(
		.INIT('h0545)
	) name3121 (
		\sub1_data_reg_reg[60]/NET0131 ,
		\sub1_ready_o_reg/NET0131 ,
		_w1054_,
		_w2230_,
		_w4050_
	);
	LUT4 #(
		.INIT('h1510)
	) name3122 (
		\state_reg/NET0131 ,
		\sub1_data_reg_reg[60]/NET0131 ,
		_w996_,
		_w4047_,
		_w4051_
	);
	LUT4 #(
		.INIT('h0057)
	) name3123 (
		\state_reg/NET0131 ,
		_w4049_,
		_w4050_,
		_w4051_,
		_w4052_
	);
	LUT3 #(
		.INIT('h48)
	) name3124 (
		\key_i[60]_pad ,
		_w931_,
		_w4052_,
		_w4053_
	);
	LUT4 #(
		.INIT('h3222)
	) name3125 (
		\data_o[60]_pad ,
		_w931_,
		_w934_,
		_w2784_,
		_w4054_
	);
	LUT4 #(
		.INIT('h7b00)
	) name3126 (
		\ks1_key_reg_reg[60]/NET0131 ,
		_w2785_,
		_w4052_,
		_w4054_,
		_w4055_
	);
	LUT2 #(
		.INIT('he)
	) name3127 (
		_w4053_,
		_w4055_,
		_w4056_
	);
	LUT4 #(
		.INIT('haab8)
	) name3128 (
		\data_i[18]_pad ,
		decrypt_i_pad,
		\mix1_data_o_reg_reg[18]/NET0131 ,
		_w930_,
		_w4057_
	);
	LUT4 #(
		.INIT('haba8)
	) name3129 (
		\sub1_data_reg_reg[18]/NET0131 ,
		_w996_,
		_w2776_,
		_w4057_,
		_w4058_
	);
	LUT4 #(
		.INIT('h404c)
	) name3130 (
		\mix1_data_o_reg_reg[18]/NET0131 ,
		_w2774_,
		_w2775_,
		_w4058_,
		_w4059_
	);
	LUT4 #(
		.INIT('h0545)
	) name3131 (
		\sub1_data_reg_reg[18]/NET0131 ,
		\sub1_ready_o_reg/NET0131 ,
		_w1054_,
		_w2230_,
		_w4060_
	);
	LUT4 #(
		.INIT('h1015)
	) name3132 (
		\state_reg/NET0131 ,
		\sub1_data_reg_reg[18]/NET0131 ,
		_w996_,
		_w4057_,
		_w4061_
	);
	LUT4 #(
		.INIT('h0057)
	) name3133 (
		\state_reg/NET0131 ,
		_w4059_,
		_w4060_,
		_w4061_,
		_w4062_
	);
	LUT3 #(
		.INIT('h48)
	) name3134 (
		\key_i[18]_pad ,
		_w931_,
		_w4062_,
		_w4063_
	);
	LUT4 #(
		.INIT('h3222)
	) name3135 (
		\data_o[18]_pad ,
		_w931_,
		_w934_,
		_w2784_,
		_w4064_
	);
	LUT4 #(
		.INIT('h7b00)
	) name3136 (
		\ks1_key_reg_reg[18]/NET0131 ,
		_w2785_,
		_w4062_,
		_w4064_,
		_w4065_
	);
	LUT2 #(
		.INIT('he)
	) name3137 (
		_w4063_,
		_w4065_,
		_w4066_
	);
	LUT3 #(
		.INIT('h2e)
	) name3138 (
		\mix1_data_o_reg_reg[11]/NET0131 ,
		_w2236_,
		_w2585_,
		_w4067_
	);
	LUT3 #(
		.INIT('h2e)
	) name3139 (
		\mix1_data_o_reg_reg[12]/NET0131 ,
		_w2236_,
		_w2604_,
		_w4068_
	);
	LUT4 #(
		.INIT('he22e)
	) name3140 (
		\mix1_data_o_reg_reg[13]/NET0131 ,
		_w2236_,
		_w2612_,
		_w2613_,
		_w4069_
	);
	LUT4 #(
		.INIT('he22e)
	) name3141 (
		\mix1_data_o_reg_reg[19]/NET0131 ,
		_w2236_,
		_w2622_,
		_w2623_,
		_w4070_
	);
	LUT4 #(
		.INIT('h8228)
	) name3142 (
		_w2236_,
		_w2384_,
		_w2625_,
		_w2626_,
		_w4071_
	);
	LUT3 #(
		.INIT('h15)
	) name3143 (
		\mix1_data_o_reg_reg[20]/NET0131 ,
		\mix1_state_reg[0]/NET0131 ,
		\mix1_state_reg[1]/NET0131 ,
		_w4072_
	);
	LUT2 #(
		.INIT('h1)
	) name3144 (
		_w4071_,
		_w4072_,
		_w4073_
	);
	LUT4 #(
		.INIT('h8228)
	) name3145 (
		_w2236_,
		_w2287_,
		_w2308_,
		_w2633_,
		_w4074_
	);
	LUT3 #(
		.INIT('h2a)
	) name3146 (
		\mix1_data_o_reg_reg[21]/NET0131 ,
		\mix1_state_reg[0]/NET0131 ,
		\mix1_state_reg[1]/NET0131 ,
		_w4075_
	);
	LUT2 #(
		.INIT('he)
	) name3147 (
		_w4074_,
		_w4075_,
		_w4076_
	);
	LUT3 #(
		.INIT('h2e)
	) name3148 (
		\mix1_data_o_reg_reg[27]/NET0131 ,
		_w2236_,
		_w2637_,
		_w4077_
	);
	LUT4 #(
		.INIT('h8228)
	) name3149 (
		_w2236_,
		_w2462_,
		_w2591_,
		_w2646_,
		_w4078_
	);
	LUT3 #(
		.INIT('h15)
	) name3150 (
		\mix1_data_o_reg_reg[28]/NET0131 ,
		\mix1_state_reg[0]/NET0131 ,
		\mix1_state_reg[1]/NET0131 ,
		_w4079_
	);
	LUT2 #(
		.INIT('h1)
	) name3151 (
		_w4078_,
		_w4079_,
		_w4080_
	);
	LUT4 #(
		.INIT('he22e)
	) name3152 (
		\mix1_data_o_reg_reg[29]/NET0131 ,
		_w2236_,
		_w2639_,
		_w2642_,
		_w4081_
	);
	LUT4 #(
		.INIT('h2ee2)
	) name3153 (
		\mix1_data_o_reg_reg[3]/NET0131 ,
		_w2236_,
		_w2507_,
		_w2622_,
		_w4082_
	);
	LUT4 #(
		.INIT('he22e)
	) name3154 (
		\mix1_data_o_reg_reg[4]/NET0131 ,
		_w2236_,
		_w2384_,
		_w2450_,
		_w4083_
	);
	LUT4 #(
		.INIT('he22e)
	) name3155 (
		\mix1_data_o_reg_reg[5]/NET0131 ,
		_w2236_,
		_w2452_,
		_w2532_,
		_w4084_
	);
	LUT4 #(
		.INIT('hcbff)
	) name3156 (
		_w2754_,
		_w2759_,
		_w2760_,
		_w2765_,
		_w4085_
	);
	LUT4 #(
		.INIT('haaac)
	) name3157 (
		\key_i[121]_pad ,
		\ks1_key_reg_reg[121]/NET0131 ,
		_w938_,
		_w986_,
		_w4086_
	);
	LUT3 #(
		.INIT('h69)
	) name3158 (
		\ks1_col_reg[25]/NET0131 ,
		_w4085_,
		_w4086_,
		_w4087_
	);
	LUT4 #(
		.INIT('haaac)
	) name3159 (
		\key_i[89]_pad ,
		\ks1_key_reg_reg[89]/NET0131 ,
		_w938_,
		_w986_,
		_w4088_
	);
	LUT4 #(
		.INIT('h9669)
	) name3160 (
		\ks1_col_reg[25]/NET0131 ,
		_w4085_,
		_w4086_,
		_w4088_,
		_w4089_
	);
	LUT4 #(
		.INIT('haaac)
	) name3161 (
		\key_i[57]_pad ,
		\ks1_key_reg_reg[57]/NET0131 ,
		_w938_,
		_w986_,
		_w4090_
	);
	LUT2 #(
		.INIT('h6)
	) name3162 (
		_w4089_,
		_w4090_,
		_w4091_
	);
	LUT3 #(
		.INIT('h69)
	) name3163 (
		_w1287_,
		_w4089_,
		_w4090_,
		_w4092_
	);
	LUT4 #(
		.INIT('hedff)
	) name3164 (
		_w2754_,
		_w2759_,
		_w2760_,
		_w2765_,
		_w4093_
	);
	LUT4 #(
		.INIT('haaac)
	) name3165 (
		\key_i[122]_pad ,
		\ks1_key_reg_reg[122]/NET0131 ,
		_w938_,
		_w986_,
		_w4094_
	);
	LUT3 #(
		.INIT('h69)
	) name3166 (
		\ks1_col_reg[26]/NET0131 ,
		_w4093_,
		_w4094_,
		_w4095_
	);
	LUT4 #(
		.INIT('haaac)
	) name3167 (
		\key_i[90]_pad ,
		\ks1_key_reg_reg[90]/NET0131 ,
		_w938_,
		_w986_,
		_w4096_
	);
	LUT4 #(
		.INIT('h9669)
	) name3168 (
		\ks1_col_reg[26]/NET0131 ,
		_w4093_,
		_w4094_,
		_w4096_,
		_w4097_
	);
	LUT4 #(
		.INIT('haaac)
	) name3169 (
		\key_i[58]_pad ,
		\ks1_key_reg_reg[58]/NET0131 ,
		_w938_,
		_w986_,
		_w4098_
	);
	LUT2 #(
		.INIT('h6)
	) name3170 (
		_w4097_,
		_w4098_,
		_w4099_
	);
	LUT3 #(
		.INIT('h69)
	) name3171 (
		_w1487_,
		_w4097_,
		_w4098_,
		_w4100_
	);
	LUT4 #(
		.INIT('hfb7f)
	) name3172 (
		_w2754_,
		_w2759_,
		_w2760_,
		_w2765_,
		_w4101_
	);
	LUT4 #(
		.INIT('haaac)
	) name3173 (
		\key_i[123]_pad ,
		\ks1_key_reg_reg[123]/NET0131 ,
		_w938_,
		_w986_,
		_w4102_
	);
	LUT3 #(
		.INIT('h69)
	) name3174 (
		\ks1_col_reg[27]/NET0131 ,
		_w4101_,
		_w4102_,
		_w4103_
	);
	LUT4 #(
		.INIT('haaac)
	) name3175 (
		\key_i[91]_pad ,
		\ks1_key_reg_reg[91]/NET0131 ,
		_w938_,
		_w986_,
		_w4104_
	);
	LUT4 #(
		.INIT('h9669)
	) name3176 (
		\ks1_col_reg[27]/NET0131 ,
		_w4101_,
		_w4102_,
		_w4104_,
		_w4105_
	);
	LUT4 #(
		.INIT('haaac)
	) name3177 (
		\key_i[59]_pad ,
		\ks1_key_reg_reg[59]/NET0131 ,
		_w938_,
		_w986_,
		_w4106_
	);
	LUT2 #(
		.INIT('h6)
	) name3178 (
		_w4105_,
		_w4106_,
		_w4107_
	);
	LUT3 #(
		.INIT('h69)
	) name3179 (
		_w1221_,
		_w4105_,
		_w4106_,
		_w4108_
	);
	LUT4 #(
		.INIT('hefdf)
	) name3180 (
		_w2754_,
		_w2759_,
		_w2760_,
		_w2765_,
		_w4109_
	);
	LUT4 #(
		.INIT('haaac)
	) name3181 (
		\key_i[125]_pad ,
		\ks1_key_reg_reg[125]/NET0131 ,
		_w938_,
		_w986_,
		_w4110_
	);
	LUT3 #(
		.INIT('h69)
	) name3182 (
		\ks1_col_reg[29]/NET0131 ,
		_w4109_,
		_w4110_,
		_w4111_
	);
	LUT4 #(
		.INIT('haaac)
	) name3183 (
		\key_i[93]_pad ,
		\ks1_key_reg_reg[93]/NET0131 ,
		_w938_,
		_w986_,
		_w4112_
	);
	LUT4 #(
		.INIT('h9669)
	) name3184 (
		\ks1_col_reg[29]/NET0131 ,
		_w4109_,
		_w4110_,
		_w4112_,
		_w4113_
	);
	LUT4 #(
		.INIT('haaac)
	) name3185 (
		\key_i[61]_pad ,
		\ks1_key_reg_reg[61]/NET0131 ,
		_w938_,
		_w986_,
		_w4114_
	);
	LUT2 #(
		.INIT('h6)
	) name3186 (
		_w4113_,
		_w4114_,
		_w4115_
	);
	LUT3 #(
		.INIT('h69)
	) name3187 (
		_w1425_,
		_w4113_,
		_w4114_,
		_w4116_
	);
	LUT3 #(
		.INIT('hc8)
	) name3188 (
		\addroundkey_start_i_reg/NET0131 ,
		\key_i[94]_pad ,
		_w936_,
		_w4117_
	);
	LUT3 #(
		.INIT('h02)
	) name3189 (
		\ks1_key_reg_reg[94]/NET0131 ,
		_w936_,
		_w938_,
		_w4118_
	);
	LUT4 #(
		.INIT('h0001)
	) name3190 (
		\addroundkey_round_reg[1]/NET0131 ,
		\addroundkey_round_reg[2]/NET0131 ,
		\addroundkey_round_reg[3]/NET0131 ,
		\key_i[94]_pad ,
		_w4119_
	);
	LUT4 #(
		.INIT('h00fe)
	) name3191 (
		\addroundkey_round_reg[1]/NET0131 ,
		\addroundkey_round_reg[2]/NET0131 ,
		\addroundkey_round_reg[3]/NET0131 ,
		\ks1_key_reg_reg[94]/NET0131 ,
		_w4120_
	);
	LUT4 #(
		.INIT('h0008)
	) name3192 (
		\addroundkey_start_i_reg/NET0131 ,
		_w930_,
		_w4120_,
		_w4119_,
		_w4121_
	);
	LUT4 #(
		.INIT('h00ab)
	) name3193 (
		_w931_,
		_w4117_,
		_w4118_,
		_w4121_,
		_w4122_
	);
	LUT4 #(
		.INIT('h0002)
	) name3194 (
		_w2754_,
		_w2759_,
		_w2760_,
		_w2765_,
		_w4123_
	);
	LUT4 #(
		.INIT('haaac)
	) name3195 (
		\key_i[126]_pad ,
		\ks1_key_reg_reg[126]/NET0131 ,
		_w938_,
		_w986_,
		_w4124_
	);
	LUT3 #(
		.INIT('h96)
	) name3196 (
		\ks1_col_reg[30]/NET0131 ,
		_w4123_,
		_w4124_,
		_w4125_
	);
	LUT4 #(
		.INIT('h6996)
	) name3197 (
		\ks1_col_reg[30]/NET0131 ,
		_w4122_,
		_w4123_,
		_w4124_,
		_w4126_
	);
	LUT4 #(
		.INIT('h9669)
	) name3198 (
		\ks1_col_reg[30]/NET0131 ,
		_w4122_,
		_w4123_,
		_w4124_,
		_w4127_
	);
	LUT4 #(
		.INIT('haaac)
	) name3199 (
		\key_i[62]_pad ,
		\ks1_key_reg_reg[62]/NET0131 ,
		_w938_,
		_w986_,
		_w4128_
	);
	LUT2 #(
		.INIT('h9)
	) name3200 (
		_w4126_,
		_w4128_,
		_w4129_
	);
	LUT3 #(
		.INIT('h96)
	) name3201 (
		_w1146_,
		_w4126_,
		_w4128_,
		_w4130_
	);
	LUT3 #(
		.INIT('hc8)
	) name3202 (
		\addroundkey_start_i_reg/NET0131 ,
		\key_i[95]_pad ,
		_w936_,
		_w4131_
	);
	LUT3 #(
		.INIT('h02)
	) name3203 (
		\ks1_key_reg_reg[95]/NET0131 ,
		_w936_,
		_w938_,
		_w4132_
	);
	LUT4 #(
		.INIT('h0001)
	) name3204 (
		\addroundkey_round_reg[1]/NET0131 ,
		\addroundkey_round_reg[2]/NET0131 ,
		\addroundkey_round_reg[3]/NET0131 ,
		\key_i[95]_pad ,
		_w4133_
	);
	LUT4 #(
		.INIT('h00fe)
	) name3205 (
		\addroundkey_round_reg[1]/NET0131 ,
		\addroundkey_round_reg[2]/NET0131 ,
		\addroundkey_round_reg[3]/NET0131 ,
		\ks1_key_reg_reg[95]/NET0131 ,
		_w4134_
	);
	LUT4 #(
		.INIT('h0008)
	) name3206 (
		\addroundkey_start_i_reg/NET0131 ,
		_w930_,
		_w4134_,
		_w4133_,
		_w4135_
	);
	LUT4 #(
		.INIT('h00ab)
	) name3207 (
		_w931_,
		_w4131_,
		_w4132_,
		_w4135_,
		_w4136_
	);
	LUT4 #(
		.INIT('h4000)
	) name3208 (
		_w2754_,
		_w2759_,
		_w2760_,
		_w2765_,
		_w4137_
	);
	LUT4 #(
		.INIT('haaac)
	) name3209 (
		\key_i[127]_pad ,
		\ks1_key_reg_reg[127]/NET0131 ,
		_w938_,
		_w986_,
		_w4138_
	);
	LUT3 #(
		.INIT('h96)
	) name3210 (
		\ks1_col_reg[31]/NET0131 ,
		_w4137_,
		_w4138_,
		_w4139_
	);
	LUT4 #(
		.INIT('h6996)
	) name3211 (
		\ks1_col_reg[31]/NET0131 ,
		_w4136_,
		_w4137_,
		_w4138_,
		_w4140_
	);
	LUT4 #(
		.INIT('h9669)
	) name3212 (
		\ks1_col_reg[31]/NET0131 ,
		_w4136_,
		_w4137_,
		_w4138_,
		_w4141_
	);
	LUT4 #(
		.INIT('haaac)
	) name3213 (
		\key_i[63]_pad ,
		\ks1_key_reg_reg[63]/NET0131 ,
		_w938_,
		_w986_,
		_w4142_
	);
	LUT2 #(
		.INIT('h9)
	) name3214 (
		_w4140_,
		_w4142_,
		_w4143_
	);
	LUT3 #(
		.INIT('h96)
	) name3215 (
		_w1534_,
		_w4140_,
		_w4142_,
		_w4144_
	);
	LUT3 #(
		.INIT('hc8)
	) name3216 (
		\addroundkey_start_i_reg/NET0131 ,
		\key_i[88]_pad ,
		_w936_,
		_w4145_
	);
	LUT3 #(
		.INIT('h02)
	) name3217 (
		\ks1_key_reg_reg[88]/NET0131 ,
		_w936_,
		_w938_,
		_w4146_
	);
	LUT4 #(
		.INIT('h0001)
	) name3218 (
		\addroundkey_round_reg[1]/NET0131 ,
		\addroundkey_round_reg[2]/NET0131 ,
		\addroundkey_round_reg[3]/NET0131 ,
		\key_i[88]_pad ,
		_w4147_
	);
	LUT4 #(
		.INIT('h00fe)
	) name3219 (
		\addroundkey_round_reg[1]/NET0131 ,
		\addroundkey_round_reg[2]/NET0131 ,
		\addroundkey_round_reg[3]/NET0131 ,
		\ks1_key_reg_reg[88]/NET0131 ,
		_w4148_
	);
	LUT4 #(
		.INIT('h0008)
	) name3220 (
		\addroundkey_start_i_reg/NET0131 ,
		_w930_,
		_w4148_,
		_w4147_,
		_w4149_
	);
	LUT4 #(
		.INIT('h00ab)
	) name3221 (
		_w931_,
		_w4145_,
		_w4146_,
		_w4149_,
		_w4150_
	);
	LUT4 #(
		.INIT('h5955)
	) name3222 (
		\ks1_col_reg[24]/NET0131 ,
		_w2759_,
		_w2760_,
		_w2765_,
		_w4151_
	);
	LUT4 #(
		.INIT('haaac)
	) name3223 (
		\key_i[120]_pad ,
		\ks1_key_reg_reg[120]/NET0131 ,
		_w938_,
		_w986_,
		_w4152_
	);
	LUT2 #(
		.INIT('h9)
	) name3224 (
		_w4151_,
		_w4152_,
		_w4153_
	);
	LUT3 #(
		.INIT('h96)
	) name3225 (
		_w4150_,
		_w4151_,
		_w4152_,
		_w4154_
	);
	LUT4 #(
		.INIT('haaac)
	) name3226 (
		\key_i[56]_pad ,
		\ks1_key_reg_reg[56]/NET0131 ,
		_w938_,
		_w986_,
		_w4155_
	);
	LUT4 #(
		.INIT('h6996)
	) name3227 (
		_w4150_,
		_w4151_,
		_w4152_,
		_w4155_,
		_w4156_
	);
	LUT2 #(
		.INIT('h9)
	) name3228 (
		_w1357_,
		_w4156_,
		_w4157_
	);
	LUT4 #(
		.INIT('h827d)
	) name3229 (
		decrypt_i_pad,
		_w2309_,
		_w2330_,
		_w2581_,
		_w4158_
	);
	LUT4 #(
		.INIT('he22e)
	) name3230 (
		\mix1_data_reg_reg[104]/NET0131 ,
		_w2233_,
		_w2557_,
		_w4158_,
		_w4159_
	);
	LUT3 #(
		.INIT('h82)
	) name3231 (
		decrypt_i_pad,
		_w2309_,
		_w2615_,
		_w4160_
	);
	LUT4 #(
		.INIT('h827d)
	) name3232 (
		decrypt_i_pad,
		_w2309_,
		_w2615_,
		_w2663_,
		_w4161_
	);
	LUT4 #(
		.INIT('h2ee2)
	) name3233 (
		\mix1_data_reg_reg[112]/NET0131 ,
		_w2233_,
		_w2619_,
		_w4161_,
		_w4162_
	);
	LUT4 #(
		.INIT('h827d)
	) name3234 (
		decrypt_i_pad,
		_w2309_,
		_w2330_,
		_w2560_,
		_w4163_
	);
	LUT4 #(
		.INIT('h2882)
	) name3235 (
		_w2233_,
		_w2556_,
		_w2618_,
		_w4163_,
		_w4164_
	);
	LUT2 #(
		.INIT('h2)
	) name3236 (
		\mix1_data_reg_reg[120]/NET0131 ,
		_w2233_,
		_w4165_
	);
	LUT2 #(
		.INIT('he)
	) name3237 (
		_w4164_,
		_w4165_,
		_w4166_
	);
	LUT3 #(
		.INIT('h2e)
	) name3238 (
		\mix1_data_reg_reg[33]/NET0131 ,
		_w2243_,
		_w2748_,
		_w4167_
	);
	LUT4 #(
		.INIT('h2882)
	) name3239 (
		_w2243_,
		_w2505_,
		_w2680_,
		_w2743_,
		_w4168_
	);
	LUT3 #(
		.INIT('h8a)
	) name3240 (
		\mix1_data_reg_reg[34]/NET0131 ,
		\mix1_state_reg[0]/NET0131 ,
		\mix1_state_reg[1]/NET0131 ,
		_w4169_
	);
	LUT2 #(
		.INIT('he)
	) name3241 (
		_w4168_,
		_w4169_,
		_w4170_
	);
	LUT4 #(
		.INIT('h8228)
	) name3242 (
		_w2243_,
		_w2330_,
		_w2651_,
		_w2653_,
		_w4171_
	);
	LUT3 #(
		.INIT('h45)
	) name3243 (
		\mix1_data_reg_reg[38]/NET0131 ,
		\mix1_state_reg[0]/NET0131 ,
		\mix1_state_reg[1]/NET0131 ,
		_w4172_
	);
	LUT2 #(
		.INIT('h1)
	) name3244 (
		_w4171_,
		_w4172_,
		_w4173_
	);
	LUT4 #(
		.INIT('h2ee2)
	) name3245 (
		\mix1_data_reg_reg[39]/NET0131 ,
		_w2243_,
		_w2657_,
		_w2658_,
		_w4174_
	);
	LUT4 #(
		.INIT('he22e)
	) name3246 (
		\mix1_data_reg_reg[41]/NET0131 ,
		_w2243_,
		_w2558_,
		_w2660_,
		_w4175_
	);
	LUT4 #(
		.INIT('h2ee2)
	) name3247 (
		\mix1_data_reg_reg[42]/NET0131 ,
		_w2243_,
		_w2662_,
		_w2667_,
		_w4176_
	);
	LUT4 #(
		.INIT('h2882)
	) name3248 (
		_w2243_,
		_w2308_,
		_w2669_,
		_w2672_,
		_w4177_
	);
	LUT3 #(
		.INIT('h8a)
	) name3249 (
		\mix1_data_reg_reg[46]/NET0131 ,
		\mix1_state_reg[0]/NET0131 ,
		\mix1_state_reg[1]/NET0131 ,
		_w4178_
	);
	LUT2 #(
		.INIT('he)
	) name3250 (
		_w4177_,
		_w4178_,
		_w4179_
	);
	LUT4 #(
		.INIT('h2ee2)
	) name3251 (
		\mix1_data_reg_reg[47]/NET0131 ,
		_w2243_,
		_w2448_,
		_w2677_,
		_w4180_
	);
	LUT3 #(
		.INIT('h2e)
	) name3252 (
		\mix1_data_reg_reg[49]/NET0131 ,
		_w2243_,
		_w2682_,
		_w4181_
	);
	LUT4 #(
		.INIT('he22e)
	) name3253 (
		\mix1_data_reg_reg[50]/NET0131 ,
		_w2243_,
		_w2684_,
		_w2688_,
		_w4182_
	);
	LUT4 #(
		.INIT('h8228)
	) name3254 (
		_w2243_,
		_w2473_,
		_w2653_,
		_w2690_,
		_w4183_
	);
	LUT3 #(
		.INIT('h45)
	) name3255 (
		\mix1_data_reg_reg[54]/NET0131 ,
		\mix1_state_reg[0]/NET0131 ,
		\mix1_state_reg[1]/NET0131 ,
		_w4184_
	);
	LUT2 #(
		.INIT('h1)
	) name3256 (
		_w4183_,
		_w4184_,
		_w4185_
	);
	LUT4 #(
		.INIT('he22e)
	) name3257 (
		\mix1_data_reg_reg[55]/NET0131 ,
		_w2243_,
		_w2657_,
		_w2694_,
		_w4186_
	);
	LUT3 #(
		.INIT('he2)
	) name3258 (
		\mix1_data_reg_reg[57]/NET0131 ,
		_w2243_,
		_w2696_,
		_w4187_
	);
	LUT4 #(
		.INIT('h2882)
	) name3259 (
		_w2243_,
		_w2246_,
		_w2698_,
		_w2699_,
		_w4188_
	);
	LUT3 #(
		.INIT('h8a)
	) name3260 (
		\mix1_data_reg_reg[58]/NET0131 ,
		\mix1_state_reg[0]/NET0131 ,
		\mix1_state_reg[1]/NET0131 ,
		_w4189_
	);
	LUT2 #(
		.INIT('he)
	) name3261 (
		_w4188_,
		_w4189_,
		_w4190_
	);
	LUT4 #(
		.INIT('h2ee2)
	) name3262 (
		\mix1_data_reg_reg[62]/NET0131 ,
		_w2243_,
		_w2672_,
		_w2703_,
		_w4191_
	);
	LUT3 #(
		.INIT('he2)
	) name3263 (
		\mix1_data_reg_reg[63]/NET0131 ,
		_w2243_,
		_w2705_,
		_w4192_
	);
	LUT3 #(
		.INIT('h2e)
	) name3264 (
		\mix1_data_reg_reg[65]/NET0131 ,
		_w2240_,
		_w2748_,
		_w4193_
	);
	LUT4 #(
		.INIT('h2882)
	) name3265 (
		_w2240_,
		_w2505_,
		_w2680_,
		_w2743_,
		_w4194_
	);
	LUT3 #(
		.INIT('ha2)
	) name3266 (
		\mix1_data_reg_reg[66]/NET0131 ,
		\mix1_state_reg[0]/NET0131 ,
		\mix1_state_reg[1]/NET0131 ,
		_w4195_
	);
	LUT2 #(
		.INIT('he)
	) name3267 (
		_w4194_,
		_w4195_,
		_w4196_
	);
	LUT4 #(
		.INIT('h8228)
	) name3268 (
		_w2240_,
		_w2330_,
		_w2651_,
		_w2653_,
		_w4197_
	);
	LUT3 #(
		.INIT('h51)
	) name3269 (
		\mix1_data_reg_reg[70]/NET0131 ,
		\mix1_state_reg[0]/NET0131 ,
		\mix1_state_reg[1]/NET0131 ,
		_w4198_
	);
	LUT2 #(
		.INIT('h1)
	) name3270 (
		_w4197_,
		_w4198_,
		_w4199_
	);
	LUT4 #(
		.INIT('h2ee2)
	) name3271 (
		\mix1_data_reg_reg[71]/NET0131 ,
		_w2240_,
		_w2657_,
		_w2658_,
		_w4200_
	);
	LUT4 #(
		.INIT('he22e)
	) name3272 (
		\mix1_data_reg_reg[73]/NET0131 ,
		_w2240_,
		_w2558_,
		_w2660_,
		_w4201_
	);
	LUT4 #(
		.INIT('h2ee2)
	) name3273 (
		\mix1_data_reg_reg[74]/NET0131 ,
		_w2240_,
		_w2662_,
		_w2667_,
		_w4202_
	);
	LUT4 #(
		.INIT('h2882)
	) name3274 (
		_w2240_,
		_w2308_,
		_w2669_,
		_w2672_,
		_w4203_
	);
	LUT3 #(
		.INIT('ha2)
	) name3275 (
		\mix1_data_reg_reg[78]/NET0131 ,
		\mix1_state_reg[0]/NET0131 ,
		\mix1_state_reg[1]/NET0131 ,
		_w4204_
	);
	LUT2 #(
		.INIT('he)
	) name3276 (
		_w4203_,
		_w4204_,
		_w4205_
	);
	LUT4 #(
		.INIT('h2ee2)
	) name3277 (
		\mix1_data_reg_reg[79]/NET0131 ,
		_w2240_,
		_w2448_,
		_w2677_,
		_w4206_
	);
	LUT3 #(
		.INIT('h2e)
	) name3278 (
		\mix1_data_reg_reg[81]/NET0131 ,
		_w2240_,
		_w2682_,
		_w4207_
	);
	LUT4 #(
		.INIT('he22e)
	) name3279 (
		\mix1_data_reg_reg[82]/NET0131 ,
		_w2240_,
		_w2684_,
		_w2688_,
		_w4208_
	);
	LUT4 #(
		.INIT('h8228)
	) name3280 (
		_w2240_,
		_w2473_,
		_w2653_,
		_w2690_,
		_w4209_
	);
	LUT3 #(
		.INIT('h51)
	) name3281 (
		\mix1_data_reg_reg[86]/NET0131 ,
		\mix1_state_reg[0]/NET0131 ,
		\mix1_state_reg[1]/NET0131 ,
		_w4210_
	);
	LUT2 #(
		.INIT('h1)
	) name3282 (
		_w4209_,
		_w4210_,
		_w4211_
	);
	LUT4 #(
		.INIT('he22e)
	) name3283 (
		\mix1_data_reg_reg[87]/NET0131 ,
		_w2240_,
		_w2657_,
		_w2694_,
		_w4212_
	);
	LUT3 #(
		.INIT('he2)
	) name3284 (
		\mix1_data_reg_reg[89]/NET0131 ,
		_w2240_,
		_w2696_,
		_w4213_
	);
	LUT4 #(
		.INIT('h2882)
	) name3285 (
		_w2240_,
		_w2246_,
		_w2698_,
		_w2699_,
		_w4214_
	);
	LUT3 #(
		.INIT('ha2)
	) name3286 (
		\mix1_data_reg_reg[90]/NET0131 ,
		\mix1_state_reg[0]/NET0131 ,
		\mix1_state_reg[1]/NET0131 ,
		_w4215_
	);
	LUT2 #(
		.INIT('he)
	) name3287 (
		_w4214_,
		_w4215_,
		_w4216_
	);
	LUT4 #(
		.INIT('h2ee2)
	) name3288 (
		\mix1_data_reg_reg[94]/NET0131 ,
		_w2240_,
		_w2672_,
		_w2703_,
		_w4217_
	);
	LUT3 #(
		.INIT('he2)
	) name3289 (
		\mix1_data_reg_reg[95]/NET0131 ,
		_w2240_,
		_w2705_,
		_w4218_
	);
	LUT2 #(
		.INIT('h9)
	) name3290 (
		_w2618_,
		_w2664_,
		_w4219_
	);
	LUT4 #(
		.INIT('h2ee2)
	) name3291 (
		\mix1_data_reg_reg[96]/NET0131 ,
		_w2233_,
		_w4160_,
		_w4219_,
		_w4220_
	);
	LUT4 #(
		.INIT('h2ee2)
	) name3292 (
		\mix1_data_o_reg_reg[10]/NET0131 ,
		_w2236_,
		_w2662_,
		_w2667_,
		_w4221_
	);
	LUT4 #(
		.INIT('h2882)
	) name3293 (
		_w2236_,
		_w2308_,
		_w2669_,
		_w2672_,
		_w4222_
	);
	LUT3 #(
		.INIT('h2a)
	) name3294 (
		\mix1_data_o_reg_reg[14]/NET0131 ,
		\mix1_state_reg[0]/NET0131 ,
		\mix1_state_reg[1]/NET0131 ,
		_w4223_
	);
	LUT2 #(
		.INIT('he)
	) name3295 (
		_w4222_,
		_w4223_,
		_w4224_
	);
	LUT4 #(
		.INIT('h2ee2)
	) name3296 (
		\mix1_data_o_reg_reg[15]/NET0131 ,
		_w2236_,
		_w2448_,
		_w2677_,
		_w4225_
	);
	LUT3 #(
		.INIT('h2e)
	) name3297 (
		\mix1_data_o_reg_reg[17]/NET0131 ,
		_w2236_,
		_w2682_,
		_w4226_
	);
	LUT4 #(
		.INIT('he22e)
	) name3298 (
		\mix1_data_o_reg_reg[18]/NET0131 ,
		_w2236_,
		_w2684_,
		_w2688_,
		_w4227_
	);
	LUT3 #(
		.INIT('h2e)
	) name3299 (
		\mix1_data_o_reg_reg[1]/NET0131 ,
		_w2236_,
		_w2748_,
		_w4228_
	);
	LUT4 #(
		.INIT('h8228)
	) name3300 (
		_w2236_,
		_w2473_,
		_w2653_,
		_w2690_,
		_w4229_
	);
	LUT3 #(
		.INIT('h15)
	) name3301 (
		\mix1_data_o_reg_reg[22]/NET0131 ,
		\mix1_state_reg[0]/NET0131 ,
		\mix1_state_reg[1]/NET0131 ,
		_w4230_
	);
	LUT2 #(
		.INIT('h1)
	) name3302 (
		_w4229_,
		_w4230_,
		_w4231_
	);
	LUT4 #(
		.INIT('he22e)
	) name3303 (
		\mix1_data_o_reg_reg[23]/NET0131 ,
		_w2236_,
		_w2657_,
		_w2694_,
		_w4232_
	);
	LUT3 #(
		.INIT('he2)
	) name3304 (
		\mix1_data_o_reg_reg[25]/NET0131 ,
		_w2236_,
		_w2696_,
		_w4233_
	);
	LUT4 #(
		.INIT('h2882)
	) name3305 (
		_w2236_,
		_w2246_,
		_w2698_,
		_w2699_,
		_w4234_
	);
	LUT3 #(
		.INIT('h2a)
	) name3306 (
		\mix1_data_o_reg_reg[26]/NET0131 ,
		\mix1_state_reg[0]/NET0131 ,
		\mix1_state_reg[1]/NET0131 ,
		_w4235_
	);
	LUT2 #(
		.INIT('he)
	) name3307 (
		_w4234_,
		_w4235_,
		_w4236_
	);
	LUT4 #(
		.INIT('h2882)
	) name3308 (
		_w2236_,
		_w2505_,
		_w2680_,
		_w2743_,
		_w4237_
	);
	LUT3 #(
		.INIT('h2a)
	) name3309 (
		\mix1_data_o_reg_reg[2]/NET0131 ,
		\mix1_state_reg[0]/NET0131 ,
		\mix1_state_reg[1]/NET0131 ,
		_w4238_
	);
	LUT2 #(
		.INIT('he)
	) name3310 (
		_w4237_,
		_w4238_,
		_w4239_
	);
	LUT4 #(
		.INIT('h2ee2)
	) name3311 (
		\mix1_data_o_reg_reg[30]/NET0131 ,
		_w2236_,
		_w2672_,
		_w2703_,
		_w4240_
	);
	LUT3 #(
		.INIT('he2)
	) name3312 (
		\mix1_data_o_reg_reg[31]/NET0131 ,
		_w2236_,
		_w2705_,
		_w4241_
	);
	LUT4 #(
		.INIT('h8228)
	) name3313 (
		_w2236_,
		_w2330_,
		_w2651_,
		_w2653_,
		_w4242_
	);
	LUT3 #(
		.INIT('h15)
	) name3314 (
		\mix1_data_o_reg_reg[6]/NET0131 ,
		\mix1_state_reg[0]/NET0131 ,
		\mix1_state_reg[1]/NET0131 ,
		_w4243_
	);
	LUT2 #(
		.INIT('h1)
	) name3315 (
		_w4242_,
		_w4243_,
		_w4244_
	);
	LUT4 #(
		.INIT('h2ee2)
	) name3316 (
		\mix1_data_o_reg_reg[7]/NET0131 ,
		_w2236_,
		_w2657_,
		_w2658_,
		_w4245_
	);
	LUT4 #(
		.INIT('he22e)
	) name3317 (
		\mix1_data_o_reg_reg[9]/NET0131 ,
		_w2236_,
		_w2558_,
		_w2660_,
		_w4246_
	);
	LUT3 #(
		.INIT('he2)
	) name3318 (
		\ks1_key_reg_reg[90]/NET0131 ,
		_w929_,
		_w4097_,
		_w4247_
	);
	LUT3 #(
		.INIT('he2)
	) name3319 (
		\ks1_key_reg_reg[93]/NET0131 ,
		_w929_,
		_w4113_,
		_w4248_
	);
	LUT4 #(
		.INIT('h2ee2)
	) name3320 (
		\mix1_data_reg_reg[32]/NET0131 ,
		_w2243_,
		_w4160_,
		_w4219_,
		_w4249_
	);
	LUT4 #(
		.INIT('he22e)
	) name3321 (
		\mix1_data_reg_reg[40]/NET0131 ,
		_w2243_,
		_w2557_,
		_w4158_,
		_w4250_
	);
	LUT4 #(
		.INIT('h2ee2)
	) name3322 (
		\mix1_data_reg_reg[48]/NET0131 ,
		_w2243_,
		_w2619_,
		_w4161_,
		_w4251_
	);
	LUT4 #(
		.INIT('h2882)
	) name3323 (
		_w2243_,
		_w2556_,
		_w2618_,
		_w4163_,
		_w4252_
	);
	LUT3 #(
		.INIT('h8a)
	) name3324 (
		\mix1_data_reg_reg[56]/NET0131 ,
		\mix1_state_reg[0]/NET0131 ,
		\mix1_state_reg[1]/NET0131 ,
		_w4253_
	);
	LUT2 #(
		.INIT('he)
	) name3325 (
		_w4252_,
		_w4253_,
		_w4254_
	);
	LUT4 #(
		.INIT('h2ee2)
	) name3326 (
		\mix1_data_reg_reg[64]/NET0131 ,
		_w2240_,
		_w4160_,
		_w4219_,
		_w4255_
	);
	LUT4 #(
		.INIT('he22e)
	) name3327 (
		\mix1_data_reg_reg[72]/NET0131 ,
		_w2240_,
		_w2557_,
		_w4158_,
		_w4256_
	);
	LUT4 #(
		.INIT('h2ee2)
	) name3328 (
		\mix1_data_reg_reg[80]/NET0131 ,
		_w2240_,
		_w2619_,
		_w4161_,
		_w4257_
	);
	LUT4 #(
		.INIT('h2882)
	) name3329 (
		_w2240_,
		_w2556_,
		_w2618_,
		_w4163_,
		_w4258_
	);
	LUT3 #(
		.INIT('ha2)
	) name3330 (
		\mix1_data_reg_reg[88]/NET0131 ,
		\mix1_state_reg[0]/NET0131 ,
		\mix1_state_reg[1]/NET0131 ,
		_w4259_
	);
	LUT2 #(
		.INIT('he)
	) name3331 (
		_w4258_,
		_w4259_,
		_w4260_
	);
	LUT3 #(
		.INIT('hc8)
	) name3332 (
		\addroundkey_start_i_reg/NET0131 ,
		\key_i[64]_pad ,
		_w936_,
		_w4261_
	);
	LUT3 #(
		.INIT('h02)
	) name3333 (
		\ks1_key_reg_reg[64]/NET0131 ,
		_w936_,
		_w938_,
		_w4262_
	);
	LUT4 #(
		.INIT('h0001)
	) name3334 (
		\addroundkey_round_reg[1]/NET0131 ,
		\addroundkey_round_reg[2]/NET0131 ,
		\addroundkey_round_reg[3]/NET0131 ,
		\key_i[64]_pad ,
		_w4263_
	);
	LUT4 #(
		.INIT('h00fe)
	) name3335 (
		\addroundkey_round_reg[1]/NET0131 ,
		\addroundkey_round_reg[2]/NET0131 ,
		\addroundkey_round_reg[3]/NET0131 ,
		\ks1_key_reg_reg[64]/NET0131 ,
		_w4264_
	);
	LUT4 #(
		.INIT('h0008)
	) name3336 (
		\addroundkey_start_i_reg/NET0131 ,
		_w930_,
		_w4264_,
		_w4263_,
		_w4265_
	);
	LUT4 #(
		.INIT('h00ab)
	) name3337 (
		_w931_,
		_w4261_,
		_w4262_,
		_w4265_,
		_w4266_
	);
	LUT4 #(
		.INIT('haaac)
	) name3338 (
		\key_i[96]_pad ,
		\ks1_key_reg_reg[96]/NET0131 ,
		_w938_,
		_w986_,
		_w4267_
	);
	LUT2 #(
		.INIT('h9)
	) name3339 (
		\ks1_col_reg[0]/NET0131 ,
		_w4267_,
		_w4268_
	);
	LUT2 #(
		.INIT('h6)
	) name3340 (
		\ks1_col_reg[0]/NET0131 ,
		_w4267_,
		_w4269_
	);
	LUT2 #(
		.INIT('h6)
	) name3341 (
		_w4266_,
		_w4268_,
		_w4270_
	);
	LUT4 #(
		.INIT('haaac)
	) name3342 (
		\key_i[32]_pad ,
		\ks1_key_reg_reg[32]/NET0131 ,
		_w938_,
		_w986_,
		_w4271_
	);
	LUT4 #(
		.INIT('h8228)
	) name3343 (
		_w929_,
		_w4266_,
		_w4268_,
		_w4271_,
		_w4272_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name3344 (
		\ks1_key_reg_reg[32]/NET0131 ,
		\ks1_state_reg[0]/NET0131 ,
		\ks1_state_reg[1]/NET0131 ,
		\ks1_state_reg[2]/NET0131 ,
		_w4273_
	);
	LUT2 #(
		.INIT('he)
	) name3345 (
		_w4272_,
		_w4273_,
		_w4274_
	);
	LUT3 #(
		.INIT('hc8)
	) name3346 (
		\addroundkey_start_i_reg/NET0131 ,
		\key_i[65]_pad ,
		_w936_,
		_w4275_
	);
	LUT3 #(
		.INIT('h02)
	) name3347 (
		\ks1_key_reg_reg[65]/NET0131 ,
		_w936_,
		_w938_,
		_w4276_
	);
	LUT4 #(
		.INIT('h0001)
	) name3348 (
		\addroundkey_round_reg[1]/NET0131 ,
		\addroundkey_round_reg[2]/NET0131 ,
		\addroundkey_round_reg[3]/NET0131 ,
		\key_i[65]_pad ,
		_w4277_
	);
	LUT4 #(
		.INIT('h00fe)
	) name3349 (
		\addroundkey_round_reg[1]/NET0131 ,
		\addroundkey_round_reg[2]/NET0131 ,
		\addroundkey_round_reg[3]/NET0131 ,
		\ks1_key_reg_reg[65]/NET0131 ,
		_w4278_
	);
	LUT4 #(
		.INIT('h0008)
	) name3350 (
		\addroundkey_start_i_reg/NET0131 ,
		_w930_,
		_w4278_,
		_w4277_,
		_w4279_
	);
	LUT4 #(
		.INIT('h00ab)
	) name3351 (
		_w931_,
		_w4275_,
		_w4276_,
		_w4279_,
		_w4280_
	);
	LUT4 #(
		.INIT('haaac)
	) name3352 (
		\key_i[97]_pad ,
		\ks1_key_reg_reg[97]/NET0131 ,
		_w938_,
		_w986_,
		_w4281_
	);
	LUT2 #(
		.INIT('h9)
	) name3353 (
		\ks1_col_reg[1]/NET0131 ,
		_w4281_,
		_w4282_
	);
	LUT2 #(
		.INIT('h6)
	) name3354 (
		\ks1_col_reg[1]/NET0131 ,
		_w4281_,
		_w4283_
	);
	LUT2 #(
		.INIT('h6)
	) name3355 (
		_w4280_,
		_w4282_,
		_w4284_
	);
	LUT4 #(
		.INIT('haaac)
	) name3356 (
		\key_i[33]_pad ,
		\ks1_key_reg_reg[33]/NET0131 ,
		_w938_,
		_w986_,
		_w4285_
	);
	LUT4 #(
		.INIT('h8228)
	) name3357 (
		_w929_,
		_w4280_,
		_w4282_,
		_w4285_,
		_w4286_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name3358 (
		\ks1_key_reg_reg[33]/NET0131 ,
		\ks1_state_reg[0]/NET0131 ,
		\ks1_state_reg[1]/NET0131 ,
		\ks1_state_reg[2]/NET0131 ,
		_w4287_
	);
	LUT2 #(
		.INIT('he)
	) name3359 (
		_w4286_,
		_w4287_,
		_w4288_
	);
	LUT3 #(
		.INIT('hc8)
	) name3360 (
		\addroundkey_start_i_reg/NET0131 ,
		\key_i[66]_pad ,
		_w936_,
		_w4289_
	);
	LUT3 #(
		.INIT('h02)
	) name3361 (
		\ks1_key_reg_reg[66]/NET0131 ,
		_w936_,
		_w938_,
		_w4290_
	);
	LUT4 #(
		.INIT('h0001)
	) name3362 (
		\addroundkey_round_reg[1]/NET0131 ,
		\addroundkey_round_reg[2]/NET0131 ,
		\addroundkey_round_reg[3]/NET0131 ,
		\key_i[66]_pad ,
		_w4291_
	);
	LUT4 #(
		.INIT('h00fe)
	) name3363 (
		\addroundkey_round_reg[1]/NET0131 ,
		\addroundkey_round_reg[2]/NET0131 ,
		\addroundkey_round_reg[3]/NET0131 ,
		\ks1_key_reg_reg[66]/NET0131 ,
		_w4292_
	);
	LUT4 #(
		.INIT('h0008)
	) name3364 (
		\addroundkey_start_i_reg/NET0131 ,
		_w930_,
		_w4292_,
		_w4291_,
		_w4293_
	);
	LUT4 #(
		.INIT('h00ab)
	) name3365 (
		_w931_,
		_w4289_,
		_w4290_,
		_w4293_,
		_w4294_
	);
	LUT4 #(
		.INIT('haaac)
	) name3366 (
		\key_i[98]_pad ,
		\ks1_key_reg_reg[98]/NET0131 ,
		_w938_,
		_w986_,
		_w4295_
	);
	LUT2 #(
		.INIT('h9)
	) name3367 (
		\ks1_col_reg[2]/NET0131 ,
		_w4295_,
		_w4296_
	);
	LUT2 #(
		.INIT('h6)
	) name3368 (
		\ks1_col_reg[2]/NET0131 ,
		_w4295_,
		_w4297_
	);
	LUT2 #(
		.INIT('h6)
	) name3369 (
		_w4294_,
		_w4296_,
		_w4298_
	);
	LUT4 #(
		.INIT('haaac)
	) name3370 (
		\key_i[34]_pad ,
		\ks1_key_reg_reg[34]/NET0131 ,
		_w938_,
		_w986_,
		_w4299_
	);
	LUT4 #(
		.INIT('h8228)
	) name3371 (
		_w929_,
		_w4294_,
		_w4296_,
		_w4299_,
		_w4300_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name3372 (
		\ks1_key_reg_reg[34]/NET0131 ,
		\ks1_state_reg[0]/NET0131 ,
		\ks1_state_reg[1]/NET0131 ,
		\ks1_state_reg[2]/NET0131 ,
		_w4301_
	);
	LUT2 #(
		.INIT('he)
	) name3373 (
		_w4300_,
		_w4301_,
		_w4302_
	);
	LUT4 #(
		.INIT('haaac)
	) name3374 (
		\key_i[99]_pad ,
		\ks1_key_reg_reg[99]/NET0131 ,
		_w938_,
		_w986_,
		_w4303_
	);
	LUT2 #(
		.INIT('h6)
	) name3375 (
		\ks1_col_reg[3]/NET0131 ,
		_w4303_,
		_w4304_
	);
	LUT4 #(
		.INIT('haaac)
	) name3376 (
		\key_i[67]_pad ,
		\ks1_key_reg_reg[67]/NET0131 ,
		_w938_,
		_w986_,
		_w4305_
	);
	LUT3 #(
		.INIT('h96)
	) name3377 (
		\ks1_col_reg[3]/NET0131 ,
		_w4303_,
		_w4305_,
		_w4306_
	);
	LUT4 #(
		.INIT('haaac)
	) name3378 (
		\key_i[35]_pad ,
		\ks1_key_reg_reg[35]/NET0131 ,
		_w938_,
		_w986_,
		_w4307_
	);
	LUT4 #(
		.INIT('h9669)
	) name3379 (
		\ks1_col_reg[3]/NET0131 ,
		_w4303_,
		_w4305_,
		_w4307_,
		_w4308_
	);
	LUT3 #(
		.INIT('h2e)
	) name3380 (
		\ks1_key_reg_reg[35]/NET0131 ,
		_w929_,
		_w4308_,
		_w4309_
	);
	LUT4 #(
		.INIT('haaac)
	) name3381 (
		\key_i[100]_pad ,
		\ks1_key_reg_reg[100]/NET0131 ,
		_w938_,
		_w986_,
		_w4310_
	);
	LUT2 #(
		.INIT('h6)
	) name3382 (
		\ks1_col_reg[4]/NET0131 ,
		_w4310_,
		_w4311_
	);
	LUT4 #(
		.INIT('haaac)
	) name3383 (
		\key_i[68]_pad ,
		\ks1_key_reg_reg[68]/NET0131 ,
		_w938_,
		_w986_,
		_w4312_
	);
	LUT3 #(
		.INIT('h96)
	) name3384 (
		\ks1_col_reg[4]/NET0131 ,
		_w4310_,
		_w4312_,
		_w4313_
	);
	LUT4 #(
		.INIT('haaac)
	) name3385 (
		\key_i[36]_pad ,
		\ks1_key_reg_reg[36]/NET0131 ,
		_w938_,
		_w986_,
		_w4314_
	);
	LUT4 #(
		.INIT('h9669)
	) name3386 (
		\ks1_col_reg[4]/NET0131 ,
		_w4310_,
		_w4312_,
		_w4314_,
		_w4315_
	);
	LUT3 #(
		.INIT('h2e)
	) name3387 (
		\ks1_key_reg_reg[36]/NET0131 ,
		_w929_,
		_w4315_,
		_w4316_
	);
	LUT4 #(
		.INIT('haaac)
	) name3388 (
		\key_i[101]_pad ,
		\ks1_key_reg_reg[101]/NET0131 ,
		_w938_,
		_w986_,
		_w4317_
	);
	LUT2 #(
		.INIT('h6)
	) name3389 (
		\ks1_col_reg[5]/NET0131 ,
		_w4317_,
		_w4318_
	);
	LUT4 #(
		.INIT('haaac)
	) name3390 (
		\key_i[69]_pad ,
		\ks1_key_reg_reg[69]/NET0131 ,
		_w938_,
		_w986_,
		_w4319_
	);
	LUT3 #(
		.INIT('h96)
	) name3391 (
		\ks1_col_reg[5]/NET0131 ,
		_w4317_,
		_w4319_,
		_w4320_
	);
	LUT4 #(
		.INIT('haaac)
	) name3392 (
		\key_i[37]_pad ,
		\ks1_key_reg_reg[37]/NET0131 ,
		_w938_,
		_w986_,
		_w4321_
	);
	LUT4 #(
		.INIT('h9669)
	) name3393 (
		\ks1_col_reg[5]/NET0131 ,
		_w4317_,
		_w4319_,
		_w4321_,
		_w4322_
	);
	LUT3 #(
		.INIT('h2e)
	) name3394 (
		\ks1_key_reg_reg[37]/NET0131 ,
		_w929_,
		_w4322_,
		_w4323_
	);
	LUT4 #(
		.INIT('haaac)
	) name3395 (
		\key_i[102]_pad ,
		\ks1_key_reg_reg[102]/NET0131 ,
		_w938_,
		_w986_,
		_w4324_
	);
	LUT2 #(
		.INIT('h6)
	) name3396 (
		\ks1_col_reg[6]/NET0131 ,
		_w4324_,
		_w4325_
	);
	LUT4 #(
		.INIT('haaac)
	) name3397 (
		\key_i[70]_pad ,
		\ks1_key_reg_reg[70]/NET0131 ,
		_w938_,
		_w986_,
		_w4326_
	);
	LUT3 #(
		.INIT('h96)
	) name3398 (
		\ks1_col_reg[6]/NET0131 ,
		_w4324_,
		_w4326_,
		_w4327_
	);
	LUT4 #(
		.INIT('haaac)
	) name3399 (
		\key_i[38]_pad ,
		\ks1_key_reg_reg[38]/NET0131 ,
		_w938_,
		_w986_,
		_w4328_
	);
	LUT4 #(
		.INIT('h9669)
	) name3400 (
		\ks1_col_reg[6]/NET0131 ,
		_w4324_,
		_w4326_,
		_w4328_,
		_w4329_
	);
	LUT3 #(
		.INIT('h2e)
	) name3401 (
		\ks1_key_reg_reg[38]/NET0131 ,
		_w929_,
		_w4329_,
		_w4330_
	);
	LUT4 #(
		.INIT('haaac)
	) name3402 (
		\key_i[103]_pad ,
		\ks1_key_reg_reg[103]/NET0131 ,
		_w938_,
		_w986_,
		_w4331_
	);
	LUT2 #(
		.INIT('h6)
	) name3403 (
		\ks1_col_reg[7]/NET0131 ,
		_w4331_,
		_w4332_
	);
	LUT4 #(
		.INIT('haaac)
	) name3404 (
		\key_i[71]_pad ,
		\ks1_key_reg_reg[71]/NET0131 ,
		_w938_,
		_w986_,
		_w4333_
	);
	LUT3 #(
		.INIT('h96)
	) name3405 (
		\ks1_col_reg[7]/NET0131 ,
		_w4331_,
		_w4333_,
		_w4334_
	);
	LUT4 #(
		.INIT('haaac)
	) name3406 (
		\key_i[39]_pad ,
		\ks1_key_reg_reg[39]/NET0131 ,
		_w938_,
		_w986_,
		_w4335_
	);
	LUT4 #(
		.INIT('h9669)
	) name3407 (
		\ks1_col_reg[7]/NET0131 ,
		_w4331_,
		_w4333_,
		_w4335_,
		_w4336_
	);
	LUT3 #(
		.INIT('h2e)
	) name3408 (
		\ks1_key_reg_reg[39]/NET0131 ,
		_w929_,
		_w4336_,
		_w4337_
	);
	LUT3 #(
		.INIT('hc8)
	) name3409 (
		\addroundkey_start_i_reg/NET0131 ,
		\key_i[80]_pad ,
		_w936_,
		_w4338_
	);
	LUT3 #(
		.INIT('h02)
	) name3410 (
		\ks1_key_reg_reg[80]/NET0131 ,
		_w936_,
		_w938_,
		_w4339_
	);
	LUT4 #(
		.INIT('h0001)
	) name3411 (
		\addroundkey_round_reg[1]/NET0131 ,
		\addroundkey_round_reg[2]/NET0131 ,
		\addroundkey_round_reg[3]/NET0131 ,
		\key_i[80]_pad ,
		_w4340_
	);
	LUT4 #(
		.INIT('h00fe)
	) name3412 (
		\addroundkey_round_reg[1]/NET0131 ,
		\addroundkey_round_reg[2]/NET0131 ,
		\addroundkey_round_reg[3]/NET0131 ,
		\ks1_key_reg_reg[80]/NET0131 ,
		_w4341_
	);
	LUT4 #(
		.INIT('h0008)
	) name3413 (
		\addroundkey_start_i_reg/NET0131 ,
		_w930_,
		_w4341_,
		_w4340_,
		_w4342_
	);
	LUT4 #(
		.INIT('h00ab)
	) name3414 (
		_w931_,
		_w4338_,
		_w4339_,
		_w4342_,
		_w4343_
	);
	LUT4 #(
		.INIT('haaac)
	) name3415 (
		\key_i[112]_pad ,
		\ks1_key_reg_reg[112]/NET0131 ,
		_w938_,
		_w986_,
		_w4344_
	);
	LUT2 #(
		.INIT('h9)
	) name3416 (
		\ks1_col_reg[16]/NET0131 ,
		_w4344_,
		_w4345_
	);
	LUT2 #(
		.INIT('h6)
	) name3417 (
		\ks1_col_reg[16]/NET0131 ,
		_w4344_,
		_w4346_
	);
	LUT2 #(
		.INIT('h6)
	) name3418 (
		_w4343_,
		_w4345_,
		_w4347_
	);
	LUT4 #(
		.INIT('haaac)
	) name3419 (
		\key_i[48]_pad ,
		\ks1_key_reg_reg[48]/NET0131 ,
		_w938_,
		_w986_,
		_w4348_
	);
	LUT4 #(
		.INIT('h8228)
	) name3420 (
		_w929_,
		_w4343_,
		_w4345_,
		_w4348_,
		_w4349_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name3421 (
		\ks1_key_reg_reg[48]/NET0131 ,
		\ks1_state_reg[0]/NET0131 ,
		\ks1_state_reg[1]/NET0131 ,
		\ks1_state_reg[2]/NET0131 ,
		_w4350_
	);
	LUT2 #(
		.INIT('he)
	) name3422 (
		_w4349_,
		_w4350_,
		_w4351_
	);
	LUT3 #(
		.INIT('hc8)
	) name3423 (
		\addroundkey_start_i_reg/NET0131 ,
		\key_i[81]_pad ,
		_w936_,
		_w4352_
	);
	LUT3 #(
		.INIT('h02)
	) name3424 (
		\ks1_key_reg_reg[81]/NET0131 ,
		_w936_,
		_w938_,
		_w4353_
	);
	LUT4 #(
		.INIT('h0001)
	) name3425 (
		\addroundkey_round_reg[1]/NET0131 ,
		\addroundkey_round_reg[2]/NET0131 ,
		\addroundkey_round_reg[3]/NET0131 ,
		\key_i[81]_pad ,
		_w4354_
	);
	LUT4 #(
		.INIT('h00fe)
	) name3426 (
		\addroundkey_round_reg[1]/NET0131 ,
		\addroundkey_round_reg[2]/NET0131 ,
		\addroundkey_round_reg[3]/NET0131 ,
		\ks1_key_reg_reg[81]/NET0131 ,
		_w4355_
	);
	LUT4 #(
		.INIT('h0008)
	) name3427 (
		\addroundkey_start_i_reg/NET0131 ,
		_w930_,
		_w4355_,
		_w4354_,
		_w4356_
	);
	LUT4 #(
		.INIT('h00ab)
	) name3428 (
		_w931_,
		_w4352_,
		_w4353_,
		_w4356_,
		_w4357_
	);
	LUT4 #(
		.INIT('haaac)
	) name3429 (
		\key_i[113]_pad ,
		\ks1_key_reg_reg[113]/NET0131 ,
		_w938_,
		_w986_,
		_w4358_
	);
	LUT2 #(
		.INIT('h9)
	) name3430 (
		\ks1_col_reg[17]/NET0131 ,
		_w4358_,
		_w4359_
	);
	LUT2 #(
		.INIT('h6)
	) name3431 (
		\ks1_col_reg[17]/NET0131 ,
		_w4358_,
		_w4360_
	);
	LUT2 #(
		.INIT('h6)
	) name3432 (
		_w4357_,
		_w4359_,
		_w4361_
	);
	LUT4 #(
		.INIT('haaac)
	) name3433 (
		\key_i[49]_pad ,
		\ks1_key_reg_reg[49]/NET0131 ,
		_w938_,
		_w986_,
		_w4362_
	);
	LUT4 #(
		.INIT('h8228)
	) name3434 (
		_w929_,
		_w4357_,
		_w4359_,
		_w4362_,
		_w4363_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name3435 (
		\ks1_key_reg_reg[49]/NET0131 ,
		\ks1_state_reg[0]/NET0131 ,
		\ks1_state_reg[1]/NET0131 ,
		\ks1_state_reg[2]/NET0131 ,
		_w4364_
	);
	LUT2 #(
		.INIT('he)
	) name3436 (
		_w4363_,
		_w4364_,
		_w4365_
	);
	LUT3 #(
		.INIT('hc8)
	) name3437 (
		\addroundkey_start_i_reg/NET0131 ,
		\key_i[82]_pad ,
		_w936_,
		_w4366_
	);
	LUT3 #(
		.INIT('h02)
	) name3438 (
		\ks1_key_reg_reg[82]/NET0131 ,
		_w936_,
		_w938_,
		_w4367_
	);
	LUT4 #(
		.INIT('h0001)
	) name3439 (
		\addroundkey_round_reg[1]/NET0131 ,
		\addroundkey_round_reg[2]/NET0131 ,
		\addroundkey_round_reg[3]/NET0131 ,
		\key_i[82]_pad ,
		_w4368_
	);
	LUT4 #(
		.INIT('h00fe)
	) name3440 (
		\addroundkey_round_reg[1]/NET0131 ,
		\addroundkey_round_reg[2]/NET0131 ,
		\addroundkey_round_reg[3]/NET0131 ,
		\ks1_key_reg_reg[82]/NET0131 ,
		_w4369_
	);
	LUT4 #(
		.INIT('h0008)
	) name3441 (
		\addroundkey_start_i_reg/NET0131 ,
		_w930_,
		_w4369_,
		_w4368_,
		_w4370_
	);
	LUT4 #(
		.INIT('h00ab)
	) name3442 (
		_w931_,
		_w4366_,
		_w4367_,
		_w4370_,
		_w4371_
	);
	LUT4 #(
		.INIT('haaac)
	) name3443 (
		\key_i[114]_pad ,
		\ks1_key_reg_reg[114]/NET0131 ,
		_w938_,
		_w986_,
		_w4372_
	);
	LUT2 #(
		.INIT('h9)
	) name3444 (
		\ks1_col_reg[18]/NET0131 ,
		_w4372_,
		_w4373_
	);
	LUT2 #(
		.INIT('h6)
	) name3445 (
		\ks1_col_reg[18]/NET0131 ,
		_w4372_,
		_w4374_
	);
	LUT2 #(
		.INIT('h6)
	) name3446 (
		_w4371_,
		_w4373_,
		_w4375_
	);
	LUT4 #(
		.INIT('haaac)
	) name3447 (
		\key_i[50]_pad ,
		\ks1_key_reg_reg[50]/NET0131 ,
		_w938_,
		_w986_,
		_w4376_
	);
	LUT4 #(
		.INIT('h8228)
	) name3448 (
		_w929_,
		_w4371_,
		_w4373_,
		_w4376_,
		_w4377_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name3449 (
		\ks1_key_reg_reg[50]/NET0131 ,
		\ks1_state_reg[0]/NET0131 ,
		\ks1_state_reg[1]/NET0131 ,
		\ks1_state_reg[2]/NET0131 ,
		_w4378_
	);
	LUT2 #(
		.INIT('he)
	) name3450 (
		_w4377_,
		_w4378_,
		_w4379_
	);
	LUT3 #(
		.INIT('hc8)
	) name3451 (
		\addroundkey_start_i_reg/NET0131 ,
		\key_i[83]_pad ,
		_w936_,
		_w4380_
	);
	LUT3 #(
		.INIT('h02)
	) name3452 (
		\ks1_key_reg_reg[83]/NET0131 ,
		_w936_,
		_w938_,
		_w4381_
	);
	LUT4 #(
		.INIT('h0001)
	) name3453 (
		\addroundkey_round_reg[1]/NET0131 ,
		\addroundkey_round_reg[2]/NET0131 ,
		\addroundkey_round_reg[3]/NET0131 ,
		\key_i[83]_pad ,
		_w4382_
	);
	LUT4 #(
		.INIT('h00fe)
	) name3454 (
		\addroundkey_round_reg[1]/NET0131 ,
		\addroundkey_round_reg[2]/NET0131 ,
		\addroundkey_round_reg[3]/NET0131 ,
		\ks1_key_reg_reg[83]/NET0131 ,
		_w4383_
	);
	LUT4 #(
		.INIT('h0008)
	) name3455 (
		\addroundkey_start_i_reg/NET0131 ,
		_w930_,
		_w4383_,
		_w4382_,
		_w4384_
	);
	LUT4 #(
		.INIT('h00ab)
	) name3456 (
		_w931_,
		_w4380_,
		_w4381_,
		_w4384_,
		_w4385_
	);
	LUT4 #(
		.INIT('haaac)
	) name3457 (
		\key_i[115]_pad ,
		\ks1_key_reg_reg[115]/NET0131 ,
		_w938_,
		_w986_,
		_w4386_
	);
	LUT2 #(
		.INIT('h9)
	) name3458 (
		\ks1_col_reg[19]/NET0131 ,
		_w4386_,
		_w4387_
	);
	LUT2 #(
		.INIT('h6)
	) name3459 (
		\ks1_col_reg[19]/NET0131 ,
		_w4386_,
		_w4388_
	);
	LUT2 #(
		.INIT('h6)
	) name3460 (
		_w4385_,
		_w4387_,
		_w4389_
	);
	LUT4 #(
		.INIT('haaac)
	) name3461 (
		\key_i[51]_pad ,
		\ks1_key_reg_reg[51]/NET0131 ,
		_w938_,
		_w986_,
		_w4390_
	);
	LUT4 #(
		.INIT('h8228)
	) name3462 (
		_w929_,
		_w4385_,
		_w4387_,
		_w4390_,
		_w4391_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name3463 (
		\ks1_key_reg_reg[51]/NET0131 ,
		\ks1_state_reg[0]/NET0131 ,
		\ks1_state_reg[1]/NET0131 ,
		\ks1_state_reg[2]/NET0131 ,
		_w4392_
	);
	LUT2 #(
		.INIT('he)
	) name3464 (
		_w4391_,
		_w4392_,
		_w4393_
	);
	LUT3 #(
		.INIT('hc8)
	) name3465 (
		\addroundkey_start_i_reg/NET0131 ,
		\key_i[84]_pad ,
		_w936_,
		_w4394_
	);
	LUT3 #(
		.INIT('h02)
	) name3466 (
		\ks1_key_reg_reg[84]/NET0131 ,
		_w936_,
		_w938_,
		_w4395_
	);
	LUT4 #(
		.INIT('h0001)
	) name3467 (
		\addroundkey_round_reg[1]/NET0131 ,
		\addroundkey_round_reg[2]/NET0131 ,
		\addroundkey_round_reg[3]/NET0131 ,
		\key_i[84]_pad ,
		_w4396_
	);
	LUT4 #(
		.INIT('h00fe)
	) name3468 (
		\addroundkey_round_reg[1]/NET0131 ,
		\addroundkey_round_reg[2]/NET0131 ,
		\addroundkey_round_reg[3]/NET0131 ,
		\ks1_key_reg_reg[84]/NET0131 ,
		_w4397_
	);
	LUT4 #(
		.INIT('h0008)
	) name3469 (
		\addroundkey_start_i_reg/NET0131 ,
		_w930_,
		_w4397_,
		_w4396_,
		_w4398_
	);
	LUT4 #(
		.INIT('h00ab)
	) name3470 (
		_w931_,
		_w4394_,
		_w4395_,
		_w4398_,
		_w4399_
	);
	LUT4 #(
		.INIT('haaac)
	) name3471 (
		\key_i[116]_pad ,
		\ks1_key_reg_reg[116]/NET0131 ,
		_w938_,
		_w986_,
		_w4400_
	);
	LUT2 #(
		.INIT('h9)
	) name3472 (
		\ks1_col_reg[20]/NET0131 ,
		_w4400_,
		_w4401_
	);
	LUT2 #(
		.INIT('h6)
	) name3473 (
		\ks1_col_reg[20]/NET0131 ,
		_w4400_,
		_w4402_
	);
	LUT2 #(
		.INIT('h6)
	) name3474 (
		_w4399_,
		_w4401_,
		_w4403_
	);
	LUT4 #(
		.INIT('haaac)
	) name3475 (
		\key_i[52]_pad ,
		\ks1_key_reg_reg[52]/NET0131 ,
		_w938_,
		_w986_,
		_w4404_
	);
	LUT4 #(
		.INIT('h8228)
	) name3476 (
		_w929_,
		_w4399_,
		_w4401_,
		_w4404_,
		_w4405_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name3477 (
		\ks1_key_reg_reg[52]/NET0131 ,
		\ks1_state_reg[0]/NET0131 ,
		\ks1_state_reg[1]/NET0131 ,
		\ks1_state_reg[2]/NET0131 ,
		_w4406_
	);
	LUT2 #(
		.INIT('he)
	) name3478 (
		_w4405_,
		_w4406_,
		_w4407_
	);
	LUT3 #(
		.INIT('hc8)
	) name3479 (
		\addroundkey_start_i_reg/NET0131 ,
		\key_i[85]_pad ,
		_w936_,
		_w4408_
	);
	LUT3 #(
		.INIT('h02)
	) name3480 (
		\ks1_key_reg_reg[85]/NET0131 ,
		_w936_,
		_w938_,
		_w4409_
	);
	LUT4 #(
		.INIT('h0001)
	) name3481 (
		\addroundkey_round_reg[1]/NET0131 ,
		\addroundkey_round_reg[2]/NET0131 ,
		\addroundkey_round_reg[3]/NET0131 ,
		\key_i[85]_pad ,
		_w4410_
	);
	LUT4 #(
		.INIT('h00fe)
	) name3482 (
		\addroundkey_round_reg[1]/NET0131 ,
		\addroundkey_round_reg[2]/NET0131 ,
		\addroundkey_round_reg[3]/NET0131 ,
		\ks1_key_reg_reg[85]/NET0131 ,
		_w4411_
	);
	LUT4 #(
		.INIT('h0008)
	) name3483 (
		\addroundkey_start_i_reg/NET0131 ,
		_w930_,
		_w4411_,
		_w4410_,
		_w4412_
	);
	LUT4 #(
		.INIT('h00ab)
	) name3484 (
		_w931_,
		_w4408_,
		_w4409_,
		_w4412_,
		_w4413_
	);
	LUT4 #(
		.INIT('haaac)
	) name3485 (
		\key_i[117]_pad ,
		\ks1_key_reg_reg[117]/NET0131 ,
		_w938_,
		_w986_,
		_w4414_
	);
	LUT2 #(
		.INIT('h9)
	) name3486 (
		\ks1_col_reg[21]/NET0131 ,
		_w4414_,
		_w4415_
	);
	LUT2 #(
		.INIT('h6)
	) name3487 (
		\ks1_col_reg[21]/NET0131 ,
		_w4414_,
		_w4416_
	);
	LUT2 #(
		.INIT('h6)
	) name3488 (
		_w4413_,
		_w4415_,
		_w4417_
	);
	LUT4 #(
		.INIT('haaac)
	) name3489 (
		\key_i[53]_pad ,
		\ks1_key_reg_reg[53]/NET0131 ,
		_w938_,
		_w986_,
		_w4418_
	);
	LUT4 #(
		.INIT('h8228)
	) name3490 (
		_w929_,
		_w4413_,
		_w4415_,
		_w4418_,
		_w4419_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name3491 (
		\ks1_key_reg_reg[53]/NET0131 ,
		\ks1_state_reg[0]/NET0131 ,
		\ks1_state_reg[1]/NET0131 ,
		\ks1_state_reg[2]/NET0131 ,
		_w4420_
	);
	LUT2 #(
		.INIT('he)
	) name3492 (
		_w4419_,
		_w4420_,
		_w4421_
	);
	LUT3 #(
		.INIT('hc8)
	) name3493 (
		\addroundkey_start_i_reg/NET0131 ,
		\key_i[86]_pad ,
		_w936_,
		_w4422_
	);
	LUT3 #(
		.INIT('h02)
	) name3494 (
		\ks1_key_reg_reg[86]/NET0131 ,
		_w936_,
		_w938_,
		_w4423_
	);
	LUT4 #(
		.INIT('h0001)
	) name3495 (
		\addroundkey_round_reg[1]/NET0131 ,
		\addroundkey_round_reg[2]/NET0131 ,
		\addroundkey_round_reg[3]/NET0131 ,
		\key_i[86]_pad ,
		_w4424_
	);
	LUT4 #(
		.INIT('h00fe)
	) name3496 (
		\addroundkey_round_reg[1]/NET0131 ,
		\addroundkey_round_reg[2]/NET0131 ,
		\addroundkey_round_reg[3]/NET0131 ,
		\ks1_key_reg_reg[86]/NET0131 ,
		_w4425_
	);
	LUT4 #(
		.INIT('h0008)
	) name3497 (
		\addroundkey_start_i_reg/NET0131 ,
		_w930_,
		_w4425_,
		_w4424_,
		_w4426_
	);
	LUT4 #(
		.INIT('h00ab)
	) name3498 (
		_w931_,
		_w4422_,
		_w4423_,
		_w4426_,
		_w4427_
	);
	LUT4 #(
		.INIT('haaac)
	) name3499 (
		\key_i[118]_pad ,
		\ks1_key_reg_reg[118]/NET0131 ,
		_w938_,
		_w986_,
		_w4428_
	);
	LUT2 #(
		.INIT('h9)
	) name3500 (
		\ks1_col_reg[22]/NET0131 ,
		_w4428_,
		_w4429_
	);
	LUT2 #(
		.INIT('h6)
	) name3501 (
		\ks1_col_reg[22]/NET0131 ,
		_w4428_,
		_w4430_
	);
	LUT2 #(
		.INIT('h6)
	) name3502 (
		_w4427_,
		_w4429_,
		_w4431_
	);
	LUT4 #(
		.INIT('haaac)
	) name3503 (
		\key_i[54]_pad ,
		\ks1_key_reg_reg[54]/NET0131 ,
		_w938_,
		_w986_,
		_w4432_
	);
	LUT4 #(
		.INIT('h8228)
	) name3504 (
		_w929_,
		_w4427_,
		_w4429_,
		_w4432_,
		_w4433_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name3505 (
		\ks1_key_reg_reg[54]/NET0131 ,
		\ks1_state_reg[0]/NET0131 ,
		\ks1_state_reg[1]/NET0131 ,
		\ks1_state_reg[2]/NET0131 ,
		_w4434_
	);
	LUT2 #(
		.INIT('he)
	) name3506 (
		_w4433_,
		_w4434_,
		_w4435_
	);
	LUT3 #(
		.INIT('hc8)
	) name3507 (
		\addroundkey_start_i_reg/NET0131 ,
		\key_i[87]_pad ,
		_w936_,
		_w4436_
	);
	LUT3 #(
		.INIT('h02)
	) name3508 (
		\ks1_key_reg_reg[87]/NET0131 ,
		_w936_,
		_w938_,
		_w4437_
	);
	LUT4 #(
		.INIT('h0001)
	) name3509 (
		\addroundkey_round_reg[1]/NET0131 ,
		\addroundkey_round_reg[2]/NET0131 ,
		\addroundkey_round_reg[3]/NET0131 ,
		\key_i[87]_pad ,
		_w4438_
	);
	LUT4 #(
		.INIT('h00fe)
	) name3510 (
		\addroundkey_round_reg[1]/NET0131 ,
		\addroundkey_round_reg[2]/NET0131 ,
		\addroundkey_round_reg[3]/NET0131 ,
		\ks1_key_reg_reg[87]/NET0131 ,
		_w4439_
	);
	LUT4 #(
		.INIT('h0008)
	) name3511 (
		\addroundkey_start_i_reg/NET0131 ,
		_w930_,
		_w4439_,
		_w4438_,
		_w4440_
	);
	LUT4 #(
		.INIT('h00ab)
	) name3512 (
		_w931_,
		_w4436_,
		_w4437_,
		_w4440_,
		_w4441_
	);
	LUT4 #(
		.INIT('haaac)
	) name3513 (
		\key_i[119]_pad ,
		\ks1_key_reg_reg[119]/NET0131 ,
		_w938_,
		_w986_,
		_w4442_
	);
	LUT2 #(
		.INIT('h9)
	) name3514 (
		\ks1_col_reg[23]/NET0131 ,
		_w4442_,
		_w4443_
	);
	LUT2 #(
		.INIT('h6)
	) name3515 (
		\ks1_col_reg[23]/NET0131 ,
		_w4442_,
		_w4444_
	);
	LUT2 #(
		.INIT('h6)
	) name3516 (
		_w4441_,
		_w4443_,
		_w4445_
	);
	LUT4 #(
		.INIT('haaac)
	) name3517 (
		\key_i[55]_pad ,
		\ks1_key_reg_reg[55]/NET0131 ,
		_w938_,
		_w986_,
		_w4446_
	);
	LUT4 #(
		.INIT('h8228)
	) name3518 (
		_w929_,
		_w4441_,
		_w4443_,
		_w4446_,
		_w4447_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name3519 (
		\ks1_key_reg_reg[55]/NET0131 ,
		\ks1_state_reg[0]/NET0131 ,
		\ks1_state_reg[1]/NET0131 ,
		\ks1_state_reg[2]/NET0131 ,
		_w4448_
	);
	LUT2 #(
		.INIT('he)
	) name3520 (
		_w4447_,
		_w4448_,
		_w4449_
	);
	LUT2 #(
		.INIT('h6)
	) name3521 (
		_w1202_,
		_w4308_,
		_w4450_
	);
	LUT2 #(
		.INIT('h6)
	) name3522 (
		_w1070_,
		_w4315_,
		_w4451_
	);
	LUT2 #(
		.INIT('h6)
	) name3523 (
		_w1411_,
		_w4322_,
		_w4452_
	);
	LUT2 #(
		.INIT('h6)
	) name3524 (
		_w1147_,
		_w4329_,
		_w4453_
	);
	LUT2 #(
		.INIT('h6)
	) name3525 (
		_w1521_,
		_w4336_,
		_w4454_
	);
	LUT4 #(
		.INIT('h9669)
	) name3526 (
		_w1363_,
		_w4266_,
		_w4268_,
		_w4271_,
		_w4455_
	);
	LUT4 #(
		.INIT('h9669)
	) name3527 (
		_w1343_,
		_w4343_,
		_w4345_,
		_w4348_,
		_w4456_
	);
	LUT4 #(
		.INIT('h9669)
	) name3528 (
		_w1280_,
		_w4357_,
		_w4359_,
		_w4362_,
		_w4457_
	);
	LUT4 #(
		.INIT('h9669)
	) name3529 (
		_w1493_,
		_w4371_,
		_w4373_,
		_w4376_,
		_w4458_
	);
	LUT4 #(
		.INIT('h9669)
	) name3530 (
		_w1208_,
		_w4385_,
		_w4387_,
		_w4390_,
		_w4459_
	);
	LUT4 #(
		.INIT('h9669)
	) name3531 (
		_w1293_,
		_w4280_,
		_w4282_,
		_w4285_,
		_w4460_
	);
	LUT4 #(
		.INIT('h9669)
	) name3532 (
		_w1085_,
		_w4399_,
		_w4401_,
		_w4404_,
		_w4461_
	);
	LUT4 #(
		.INIT('h9669)
	) name3533 (
		_w1418_,
		_w4413_,
		_w4415_,
		_w4418_,
		_w4462_
	);
	LUT4 #(
		.INIT('h9669)
	) name3534 (
		_w1148_,
		_w4427_,
		_w4429_,
		_w4432_,
		_w4463_
	);
	LUT4 #(
		.INIT('h9669)
	) name3535 (
		_w1515_,
		_w4441_,
		_w4443_,
		_w4446_,
		_w4464_
	);
	LUT4 #(
		.INIT('h9669)
	) name3536 (
		_w1506_,
		_w4294_,
		_w4296_,
		_w4299_,
		_w4465_
	);
	LUT4 #(
		.INIT('h2ee2)
	) name3537 (
		\mix1_data_o_reg_reg[0]/NET0131 ,
		_w2236_,
		_w4160_,
		_w4219_,
		_w4466_
	);
	LUT4 #(
		.INIT('h2ee2)
	) name3538 (
		\mix1_data_o_reg_reg[16]/NET0131 ,
		_w2236_,
		_w2619_,
		_w4161_,
		_w4467_
	);
	LUT4 #(
		.INIT('h2882)
	) name3539 (
		_w2236_,
		_w2556_,
		_w2618_,
		_w4163_,
		_w4468_
	);
	LUT3 #(
		.INIT('h2a)
	) name3540 (
		\mix1_data_o_reg_reg[24]/NET0131 ,
		\mix1_state_reg[0]/NET0131 ,
		\mix1_state_reg[1]/NET0131 ,
		_w4469_
	);
	LUT2 #(
		.INIT('he)
	) name3541 (
		_w4468_,
		_w4469_,
		_w4470_
	);
	LUT4 #(
		.INIT('he22e)
	) name3542 (
		\mix1_data_o_reg_reg[8]/NET0131 ,
		_w2236_,
		_w2557_,
		_w4158_,
		_w4471_
	);
	LUT4 #(
		.INIT('hf0e0)
	) name3543 (
		\ks1_state_reg[1]/NET0131 ,
		_w938_,
		_w946_,
		_w945_,
		_w4472_
	);
	LUT4 #(
		.INIT('hf1fa)
	) name3544 (
		\addroundkey_round_reg[0]/NET0131 ,
		_w934_,
		_w938_,
		_w944_,
		_w4473_
	);
	LUT2 #(
		.INIT('h2)
	) name3545 (
		\addroundkey_round_reg[3]/NET0131 ,
		\ks1_ready_o_reg/NET0131 ,
		_w4474_
	);
	LUT4 #(
		.INIT('hf5f4)
	) name3546 (
		\addroundkey_start_i_reg/NET0131 ,
		_w2752_,
		_w2753_,
		_w4474_,
		_w4475_
	);
	LUT2 #(
		.INIT('h2)
	) name3547 (
		\addroundkey_round_reg[1]/NET0131 ,
		\ks1_ready_o_reg/NET0131 ,
		_w4476_
	);
	LUT4 #(
		.INIT('hf5f4)
	) name3548 (
		\addroundkey_start_i_reg/NET0131 ,
		_w2757_,
		_w2758_,
		_w4476_,
		_w4477_
	);
	LUT2 #(
		.INIT('h2)
	) name3549 (
		\addroundkey_round_reg[2]/NET0131 ,
		\ks1_ready_o_reg/NET0131 ,
		_w4478_
	);
	LUT4 #(
		.INIT('hf5f4)
	) name3550 (
		\addroundkey_start_i_reg/NET0131 ,
		_w2763_,
		_w2764_,
		_w4478_,
		_w4479_
	);
	LUT3 #(
		.INIT('hea)
	) name3551 (
		_w931_,
		_w934_,
		_w2784_,
		_w4480_
	);
	LUT3 #(
		.INIT('h0d)
	) name3552 (
		\sub1_ready_o_reg/NET0131 ,
		_w2230_,
		_w2775_,
		_w4481_
	);
	LUT4 #(
		.INIT('h807f)
	) name3553 (
		\round_reg[0]/NET0131 ,
		\round_reg[1]/NET0131 ,
		\round_reg[2]/NET0131 ,
		\round_reg[3]/NET0131 ,
		_w4482_
	);
	LUT4 #(
		.INIT('hf200)
	) name3554 (
		\sub1_ready_o_reg/NET0131 ,
		_w2230_,
		_w2775_,
		_w4482_,
		_w4483_
	);
	LUT4 #(
		.INIT('h0200)
	) name3555 (
		decrypt_i_pad,
		\round_reg[0]/NET0131 ,
		\round_reg[1]/NET0131 ,
		\sub1_ready_o_reg/NET0131 ,
		_w4484_
	);
	LUT3 #(
		.INIT('h8c)
	) name3556 (
		\round_reg[2]/NET0131 ,
		\round_reg[3]/NET0131 ,
		_w4484_,
		_w4485_
	);
	LUT3 #(
		.INIT('h80)
	) name3557 (
		decrypt_i_pad,
		\sub1_ready_o_reg/NET0131 ,
		_w930_,
		_w4486_
	);
	LUT2 #(
		.INIT('h1)
	) name3558 (
		_w4485_,
		_w4486_,
		_w4487_
	);
	LUT4 #(
		.INIT('ha280)
	) name3559 (
		\addroundkey_ready_o_reg/NET0131 ,
		decrypt_i_pad,
		_w930_,
		_w995_,
		_w4488_
	);
	LUT2 #(
		.INIT('h2)
	) name3560 (
		\state_reg/NET0131 ,
		_w4488_,
		_w4489_
	);
	LUT4 #(
		.INIT('h0070)
	) name3561 (
		_w4481_,
		_w4487_,
		_w4489_,
		_w4483_,
		_w4490_
	);
	LUT2 #(
		.INIT('h1)
	) name3562 (
		load_i_pad,
		\state_reg/NET0131 ,
		_w4491_
	);
	LUT2 #(
		.INIT('h2)
	) name3563 (
		load_i_pad,
		\state_reg/NET0131 ,
		_w4492_
	);
	LUT4 #(
		.INIT('hff47)
	) name3564 (
		decrypt_i_pad,
		load_i_pad,
		\round_reg[3]/NET0131 ,
		\state_reg/NET0131 ,
		_w4493_
	);
	LUT2 #(
		.INIT('hb)
	) name3565 (
		_w4490_,
		_w4493_,
		_w4494_
	);
	LUT2 #(
		.INIT('h6)
	) name3566 (
		\round_reg[0]/NET0131 ,
		\round_reg[1]/NET0131 ,
		_w4495_
	);
	LUT3 #(
		.INIT('h13)
	) name3567 (
		decrypt_i_pad,
		\round_reg[0]/NET0131 ,
		\sub1_ready_o_reg/NET0131 ,
		_w4496_
	);
	LUT4 #(
		.INIT('h000d)
	) name3568 (
		\sub1_ready_o_reg/NET0131 ,
		_w2230_,
		_w2775_,
		_w4496_,
		_w4497_
	);
	LUT4 #(
		.INIT('hff47)
	) name3569 (
		decrypt_i_pad,
		load_i_pad,
		\round_reg[1]/NET0131 ,
		\state_reg/NET0131 ,
		_w4498_
	);
	LUT4 #(
		.INIT('h28ff)
	) name3570 (
		_w4489_,
		_w4495_,
		_w4497_,
		_w4498_,
		_w4499_
	);
	LUT2 #(
		.INIT('he)
	) name3571 (
		_w2233_,
		_w2243_,
		_w4500_
	);
	LUT2 #(
		.INIT('h6)
	) name3572 (
		\mix1_state_reg[0]/NET0131 ,
		\mix1_state_reg[1]/NET0131 ,
		_w4501_
	);
	LUT2 #(
		.INIT('h2)
	) name3573 (
		\first_round_reg_reg/NET0131 ,
		\state_reg/NET0131 ,
		_w4502_
	);
	LUT4 #(
		.INIT('h0123)
	) name3574 (
		decrypt_i_pad,
		\first_round_reg_reg/NET0131 ,
		\mix1_ready_o_reg/NET0131 ,
		\sub1_ready_o_reg/NET0131 ,
		_w4503_
	);
	LUT3 #(
		.INIT('hd1)
	) name3575 (
		\sub1_ready_o_reg/NET0131 ,
		_w2230_,
		_w4503_,
		_w4504_
	);
	LUT3 #(
		.INIT('hce)
	) name3576 (
		_w4489_,
		_w4502_,
		_w4504_,
		_w4505_
	);
	LUT4 #(
		.INIT('h5554)
	) name3577 (
		\sub1_state_reg[0]/NET0131 ,
		\sub1_state_reg[1]/NET0131 ,
		\sub1_state_reg[2]/NET0131 ,
		\sub1_state_reg[3]/NET0131 ,
		_w4506_
	);
	LUT4 #(
		.INIT('hab00)
	) name3578 (
		\sub1_state_reg[0]/NET0131 ,
		_w1055_,
		_w1056_,
		_w1060_,
		_w4507_
	);
	LUT2 #(
		.INIT('he)
	) name3579 (
		_w4506_,
		_w4507_,
		_w4508_
	);
	LUT3 #(
		.INIT('h04)
	) name3580 (
		load_i_pad,
		\round_reg[2]/NET0131 ,
		\state_reg/NET0131 ,
		_w4509_
	);
	LUT3 #(
		.INIT('h21)
	) name3581 (
		\round_reg[2]/NET0131 ,
		_w2775_,
		_w4484_,
		_w4510_
	);
	LUT3 #(
		.INIT('h78)
	) name3582 (
		\round_reg[0]/NET0131 ,
		\round_reg[1]/NET0131 ,
		\round_reg[2]/NET0131 ,
		_w4511_
	);
	LUT2 #(
		.INIT('h2)
	) name3583 (
		_w2775_,
		_w4511_,
		_w4512_
	);
	LUT3 #(
		.INIT('h02)
	) name3584 (
		_w2230_,
		_w4510_,
		_w4512_,
		_w4513_
	);
	LUT3 #(
		.INIT('hec)
	) name3585 (
		_w4489_,
		_w4509_,
		_w4513_,
		_w4514_
	);
	LUT3 #(
		.INIT('h46)
	) name3586 (
		\sub1_state_reg[4]/NET0131 ,
		_w1009_,
		_w1053_,
		_w4515_
	);
	LUT3 #(
		.INIT('h78)
	) name3587 (
		\sub1_state_reg[0]/NET0131 ,
		\sub1_state_reg[1]/NET0131 ,
		\sub1_state_reg[2]/NET0131 ,
		_w4516_
	);
	LUT4 #(
		.INIT('h1b0b)
	) name3588 (
		decrypt_i_pad,
		\mix1_ready_o_reg/NET0131 ,
		\sub1_ready_o_reg/NET0131 ,
		_w2230_,
		_w4517_
	);
	LUT4 #(
		.INIT('ha8d8)
	) name3589 (
		\round_reg[0]/NET0131 ,
		_w4491_,
		_w4489_,
		_w4517_,
		_w4518_
	);
	LUT3 #(
		.INIT('h2e)
	) name3590 (
		load_i_pad,
		\state_reg/NET0131 ,
		_w4488_,
		_w4519_
	);
	LUT2 #(
		.INIT('h8)
	) name3591 (
		\addroundkey_ready_o_reg/NET0131 ,
		_w1055_,
		_w4520_
	);
	LUT4 #(
		.INIT('h7f80)
	) name3592 (
		\sub1_state_reg[0]/NET0131 ,
		\sub1_state_reg[1]/NET0131 ,
		\sub1_state_reg[2]/NET0131 ,
		\sub1_state_reg[3]/NET0131 ,
		_w4521_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name3593 (
		\mix1_data_o_reg_reg[89]/NET0131 ,
		\mix1_data_reg_reg[89]/NET0131 ,
		\mix1_state_reg[0]/NET0131 ,
		\mix1_state_reg[1]/NET0131 ,
		_w4522_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name3594 (
		\mix1_data_o_reg_reg[99]/NET0131 ,
		\mix1_data_reg_reg[99]/NET0131 ,
		\mix1_state_reg[0]/NET0131 ,
		\mix1_state_reg[1]/NET0131 ,
		_w4523_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name3595 (
		\mix1_data_o_reg_reg[37]/NET0131 ,
		\mix1_data_reg_reg[37]/NET0131 ,
		\mix1_state_reg[0]/NET0131 ,
		\mix1_state_reg[1]/NET0131 ,
		_w4524_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name3596 (
		\mix1_data_o_reg_reg[110]/NET0131 ,
		\mix1_data_reg_reg[110]/NET0131 ,
		\mix1_state_reg[0]/NET0131 ,
		\mix1_state_reg[1]/NET0131 ,
		_w4525_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name3597 (
		\mix1_data_o_reg_reg[40]/NET0131 ,
		\mix1_data_reg_reg[40]/NET0131 ,
		\mix1_state_reg[0]/NET0131 ,
		\mix1_state_reg[1]/NET0131 ,
		_w4526_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name3598 (
		\mix1_data_o_reg_reg[34]/NET0131 ,
		\mix1_data_reg_reg[34]/NET0131 ,
		\mix1_state_reg[0]/NET0131 ,
		\mix1_state_reg[1]/NET0131 ,
		_w4527_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name3599 (
		\mix1_data_o_reg_reg[48]/NET0131 ,
		\mix1_data_reg_reg[48]/NET0131 ,
		\mix1_state_reg[0]/NET0131 ,
		\mix1_state_reg[1]/NET0131 ,
		_w4528_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name3600 (
		\mix1_data_o_reg_reg[105]/NET0131 ,
		\mix1_data_reg_reg[105]/NET0131 ,
		\mix1_state_reg[0]/NET0131 ,
		\mix1_state_reg[1]/NET0131 ,
		_w4529_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name3601 (
		\mix1_data_o_reg_reg[43]/NET0131 ,
		\mix1_data_reg_reg[43]/NET0131 ,
		\mix1_state_reg[0]/NET0131 ,
		\mix1_state_reg[1]/NET0131 ,
		_w4530_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name3602 (
		\mix1_data_o_reg_reg[95]/NET0131 ,
		\mix1_data_reg_reg[95]/NET0131 ,
		\mix1_state_reg[0]/NET0131 ,
		\mix1_state_reg[1]/NET0131 ,
		_w4531_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name3603 (
		\mix1_data_o_reg_reg[93]/NET0131 ,
		\mix1_data_reg_reg[93]/NET0131 ,
		\mix1_state_reg[0]/NET0131 ,
		\mix1_state_reg[1]/NET0131 ,
		_w4532_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name3604 (
		\mix1_data_o_reg_reg[97]/NET0131 ,
		\mix1_data_reg_reg[97]/NET0131 ,
		\mix1_state_reg[0]/NET0131 ,
		\mix1_state_reg[1]/NET0131 ,
		_w4533_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name3605 (
		\mix1_data_o_reg_reg[35]/NET0131 ,
		\mix1_data_reg_reg[35]/NET0131 ,
		\mix1_state_reg[0]/NET0131 ,
		\mix1_state_reg[1]/NET0131 ,
		_w4534_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name3606 (
		\mix1_data_o_reg_reg[106]/NET0131 ,
		\mix1_data_reg_reg[106]/NET0131 ,
		\mix1_state_reg[0]/NET0131 ,
		\mix1_state_reg[1]/NET0131 ,
		_w4535_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name3607 (
		\mix1_data_o_reg_reg[107]/NET0131 ,
		\mix1_data_reg_reg[107]/NET0131 ,
		\mix1_state_reg[0]/NET0131 ,
		\mix1_state_reg[1]/NET0131 ,
		_w4536_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name3608 (
		\mix1_data_o_reg_reg[108]/NET0131 ,
		\mix1_data_reg_reg[108]/NET0131 ,
		\mix1_state_reg[0]/NET0131 ,
		\mix1_state_reg[1]/NET0131 ,
		_w4537_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name3609 (
		\mix1_data_o_reg_reg[91]/NET0131 ,
		\mix1_data_reg_reg[91]/NET0131 ,
		\mix1_state_reg[0]/NET0131 ,
		\mix1_state_reg[1]/NET0131 ,
		_w4538_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name3610 (
		\mix1_data_o_reg_reg[111]/NET0131 ,
		\mix1_data_reg_reg[111]/NET0131 ,
		\mix1_state_reg[0]/NET0131 ,
		\mix1_state_reg[1]/NET0131 ,
		_w4539_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name3611 (
		\mix1_data_o_reg_reg[33]/NET0131 ,
		\mix1_data_reg_reg[33]/NET0131 ,
		\mix1_state_reg[0]/NET0131 ,
		\mix1_state_reg[1]/NET0131 ,
		_w4540_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name3612 (
		\mix1_data_o_reg_reg[114]/NET0131 ,
		\mix1_data_reg_reg[114]/NET0131 ,
		\mix1_state_reg[0]/NET0131 ,
		\mix1_state_reg[1]/NET0131 ,
		_w4541_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name3613 (
		\mix1_data_o_reg_reg[115]/NET0131 ,
		\mix1_data_reg_reg[115]/NET0131 ,
		\mix1_state_reg[0]/NET0131 ,
		\mix1_state_reg[1]/NET0131 ,
		_w4542_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name3614 (
		\mix1_data_o_reg_reg[116]/NET0131 ,
		\mix1_data_reg_reg[116]/NET0131 ,
		\mix1_state_reg[0]/NET0131 ,
		\mix1_state_reg[1]/NET0131 ,
		_w4543_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name3615 (
		\mix1_data_o_reg_reg[118]/NET0131 ,
		\mix1_data_reg_reg[118]/NET0131 ,
		\mix1_state_reg[0]/NET0131 ,
		\mix1_state_reg[1]/NET0131 ,
		_w4544_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name3616 (
		\mix1_data_o_reg_reg[120]/NET0131 ,
		\mix1_data_reg_reg[120]/NET0131 ,
		\mix1_state_reg[0]/NET0131 ,
		\mix1_state_reg[1]/NET0131 ,
		_w4545_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name3617 (
		\mix1_data_o_reg_reg[112]/NET0131 ,
		\mix1_data_reg_reg[112]/NET0131 ,
		\mix1_state_reg[0]/NET0131 ,
		\mix1_state_reg[1]/NET0131 ,
		_w4546_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name3618 (
		\mix1_data_o_reg_reg[124]/NET0131 ,
		\mix1_data_reg_reg[124]/NET0131 ,
		\mix1_state_reg[0]/NET0131 ,
		\mix1_state_reg[1]/NET0131 ,
		_w4547_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name3619 (
		\mix1_data_o_reg_reg[83]/NET0131 ,
		\mix1_data_reg_reg[83]/NET0131 ,
		\mix1_state_reg[0]/NET0131 ,
		\mix1_state_reg[1]/NET0131 ,
		_w4548_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name3620 (
		\mix1_data_o_reg_reg[81]/NET0131 ,
		\mix1_data_reg_reg[81]/NET0131 ,
		\mix1_state_reg[0]/NET0131 ,
		\mix1_state_reg[1]/NET0131 ,
		_w4549_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name3621 (
		\mix1_data_o_reg_reg[42]/NET0131 ,
		\mix1_data_reg_reg[42]/NET0131 ,
		\mix1_state_reg[0]/NET0131 ,
		\mix1_state_reg[1]/NET0131 ,
		_w4550_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name3622 (
		\mix1_data_o_reg_reg[32]/NET0131 ,
		\mix1_data_reg_reg[32]/NET0131 ,
		\mix1_state_reg[0]/NET0131 ,
		\mix1_state_reg[1]/NET0131 ,
		_w4551_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name3623 (
		\mix1_data_o_reg_reg[113]/NET0131 ,
		\mix1_data_reg_reg[113]/NET0131 ,
		\mix1_state_reg[0]/NET0131 ,
		\mix1_state_reg[1]/NET0131 ,
		_w4552_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name3624 (
		\mix1_data_o_reg_reg[38]/NET0131 ,
		\mix1_data_reg_reg[38]/NET0131 ,
		\mix1_state_reg[0]/NET0131 ,
		\mix1_state_reg[1]/NET0131 ,
		_w4553_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name3625 (
		\mix1_data_o_reg_reg[41]/NET0131 ,
		\mix1_data_reg_reg[41]/NET0131 ,
		\mix1_state_reg[0]/NET0131 ,
		\mix1_state_reg[1]/NET0131 ,
		_w4554_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name3626 (
		\mix1_data_o_reg_reg[45]/NET0131 ,
		\mix1_data_reg_reg[45]/NET0131 ,
		\mix1_state_reg[0]/NET0131 ,
		\mix1_state_reg[1]/NET0131 ,
		_w4555_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name3627 (
		\mix1_data_o_reg_reg[49]/NET0131 ,
		\mix1_data_reg_reg[49]/NET0131 ,
		\mix1_state_reg[0]/NET0131 ,
		\mix1_state_reg[1]/NET0131 ,
		_w4556_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name3628 (
		\mix1_data_o_reg_reg[52]/NET0131 ,
		\mix1_data_reg_reg[52]/NET0131 ,
		\mix1_state_reg[0]/NET0131 ,
		\mix1_state_reg[1]/NET0131 ,
		_w4557_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name3629 (
		\mix1_data_o_reg_reg[56]/NET0131 ,
		\mix1_data_reg_reg[56]/NET0131 ,
		\mix1_state_reg[0]/NET0131 ,
		\mix1_state_reg[1]/NET0131 ,
		_w4558_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name3630 (
		\mix1_data_o_reg_reg[61]/NET0131 ,
		\mix1_data_reg_reg[61]/NET0131 ,
		\mix1_state_reg[0]/NET0131 ,
		\mix1_state_reg[1]/NET0131 ,
		_w4559_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name3631 (
		\mix1_data_o_reg_reg[62]/NET0131 ,
		\mix1_data_reg_reg[62]/NET0131 ,
		\mix1_state_reg[0]/NET0131 ,
		\mix1_state_reg[1]/NET0131 ,
		_w4560_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name3632 (
		\mix1_data_o_reg_reg[64]/NET0131 ,
		\mix1_data_reg_reg[64]/NET0131 ,
		\mix1_state_reg[0]/NET0131 ,
		\mix1_state_reg[1]/NET0131 ,
		_w4561_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name3633 (
		\mix1_data_o_reg_reg[125]/NET0131 ,
		\mix1_data_reg_reg[125]/NET0131 ,
		\mix1_state_reg[0]/NET0131 ,
		\mix1_state_reg[1]/NET0131 ,
		_w4562_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name3634 (
		\mix1_data_o_reg_reg[71]/NET0131 ,
		\mix1_data_reg_reg[71]/NET0131 ,
		\mix1_state_reg[0]/NET0131 ,
		\mix1_state_reg[1]/NET0131 ,
		_w4563_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name3635 (
		\mix1_data_o_reg_reg[75]/NET0131 ,
		\mix1_data_reg_reg[75]/NET0131 ,
		\mix1_state_reg[0]/NET0131 ,
		\mix1_state_reg[1]/NET0131 ,
		_w4564_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name3636 (
		\mix1_data_o_reg_reg[77]/NET0131 ,
		\mix1_data_reg_reg[77]/NET0131 ,
		\mix1_state_reg[0]/NET0131 ,
		\mix1_state_reg[1]/NET0131 ,
		_w4565_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name3637 (
		\mix1_data_o_reg_reg[80]/NET0131 ,
		\mix1_data_reg_reg[80]/NET0131 ,
		\mix1_state_reg[0]/NET0131 ,
		\mix1_state_reg[1]/NET0131 ,
		_w4566_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name3638 (
		\mix1_data_o_reg_reg[98]/NET0131 ,
		\mix1_data_reg_reg[98]/NET0131 ,
		\mix1_state_reg[0]/NET0131 ,
		\mix1_state_reg[1]/NET0131 ,
		_w4567_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name3639 (
		\mix1_data_o_reg_reg[84]/NET0131 ,
		\mix1_data_reg_reg[84]/NET0131 ,
		\mix1_state_reg[0]/NET0131 ,
		\mix1_state_reg[1]/NET0131 ,
		_w4568_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name3640 (
		\mix1_data_o_reg_reg[90]/NET0131 ,
		\mix1_data_reg_reg[90]/NET0131 ,
		\mix1_state_reg[0]/NET0131 ,
		\mix1_state_reg[1]/NET0131 ,
		_w4569_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name3641 (
		\mix1_data_o_reg_reg[92]/NET0131 ,
		\mix1_data_reg_reg[92]/NET0131 ,
		\mix1_state_reg[0]/NET0131 ,
		\mix1_state_reg[1]/NET0131 ,
		_w4570_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name3642 (
		\mix1_data_o_reg_reg[94]/NET0131 ,
		\mix1_data_reg_reg[94]/NET0131 ,
		\mix1_state_reg[0]/NET0131 ,
		\mix1_state_reg[1]/NET0131 ,
		_w4571_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name3643 (
		\mix1_data_o_reg_reg[76]/NET0131 ,
		\mix1_data_reg_reg[76]/NET0131 ,
		\mix1_state_reg[0]/NET0131 ,
		\mix1_state_reg[1]/NET0131 ,
		_w4572_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name3644 (
		\mix1_data_o_reg_reg[127]/NET0131 ,
		\mix1_data_reg_reg[127]/NET0131 ,
		\mix1_state_reg[0]/NET0131 ,
		\mix1_state_reg[1]/NET0131 ,
		_w4573_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name3645 (
		\mix1_data_o_reg_reg[109]/NET0131 ,
		\mix1_data_reg_reg[109]/NET0131 ,
		\mix1_state_reg[0]/NET0131 ,
		\mix1_state_reg[1]/NET0131 ,
		_w4574_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name3646 (
		\mix1_data_o_reg_reg[78]/NET0131 ,
		\mix1_data_reg_reg[78]/NET0131 ,
		\mix1_state_reg[0]/NET0131 ,
		\mix1_state_reg[1]/NET0131 ,
		_w4575_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name3647 (
		\mix1_data_o_reg_reg[72]/NET0131 ,
		\mix1_data_reg_reg[72]/NET0131 ,
		\mix1_state_reg[0]/NET0131 ,
		\mix1_state_reg[1]/NET0131 ,
		_w4576_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name3648 (
		\mix1_data_o_reg_reg[50]/NET0131 ,
		\mix1_data_reg_reg[50]/NET0131 ,
		\mix1_state_reg[0]/NET0131 ,
		\mix1_state_reg[1]/NET0131 ,
		_w4577_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name3649 (
		\mix1_data_o_reg_reg[87]/NET0131 ,
		\mix1_data_reg_reg[87]/NET0131 ,
		\mix1_state_reg[0]/NET0131 ,
		\mix1_state_reg[1]/NET0131 ,
		_w4578_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name3650 (
		\mix1_data_o_reg_reg[123]/NET0131 ,
		\mix1_data_reg_reg[123]/NET0131 ,
		\mix1_state_reg[0]/NET0131 ,
		\mix1_state_reg[1]/NET0131 ,
		_w4579_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name3651 (
		\mix1_data_o_reg_reg[70]/NET0131 ,
		\mix1_data_reg_reg[70]/NET0131 ,
		\mix1_state_reg[0]/NET0131 ,
		\mix1_state_reg[1]/NET0131 ,
		_w4580_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name3652 (
		\mix1_data_o_reg_reg[39]/NET0131 ,
		\mix1_data_reg_reg[39]/NET0131 ,
		\mix1_state_reg[0]/NET0131 ,
		\mix1_state_reg[1]/NET0131 ,
		_w4581_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name3653 (
		\mix1_data_o_reg_reg[122]/NET0131 ,
		\mix1_data_reg_reg[122]/NET0131 ,
		\mix1_state_reg[0]/NET0131 ,
		\mix1_state_reg[1]/NET0131 ,
		_w4582_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name3654 (
		\mix1_data_o_reg_reg[121]/NET0131 ,
		\mix1_data_reg_reg[121]/NET0131 ,
		\mix1_state_reg[0]/NET0131 ,
		\mix1_state_reg[1]/NET0131 ,
		_w4583_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name3655 (
		\mix1_data_o_reg_reg[79]/NET0131 ,
		\mix1_data_reg_reg[79]/NET0131 ,
		\mix1_state_reg[0]/NET0131 ,
		\mix1_state_reg[1]/NET0131 ,
		_w4584_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name3656 (
		\mix1_data_o_reg_reg[88]/NET0131 ,
		\mix1_data_reg_reg[88]/NET0131 ,
		\mix1_state_reg[0]/NET0131 ,
		\mix1_state_reg[1]/NET0131 ,
		_w4585_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name3657 (
		\mix1_data_o_reg_reg[85]/NET0131 ,
		\mix1_data_reg_reg[85]/NET0131 ,
		\mix1_state_reg[0]/NET0131 ,
		\mix1_state_reg[1]/NET0131 ,
		_w4586_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name3658 (
		\mix1_data_o_reg_reg[103]/NET0131 ,
		\mix1_data_reg_reg[103]/NET0131 ,
		\mix1_state_reg[0]/NET0131 ,
		\mix1_state_reg[1]/NET0131 ,
		_w4587_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name3659 (
		\mix1_data_o_reg_reg[69]/NET0131 ,
		\mix1_data_reg_reg[69]/NET0131 ,
		\mix1_state_reg[0]/NET0131 ,
		\mix1_state_reg[1]/NET0131 ,
		_w4588_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name3660 (
		\mix1_data_o_reg_reg[73]/NET0131 ,
		\mix1_data_reg_reg[73]/NET0131 ,
		\mix1_state_reg[0]/NET0131 ,
		\mix1_state_reg[1]/NET0131 ,
		_w4589_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name3661 (
		\mix1_data_o_reg_reg[104]/NET0131 ,
		\mix1_data_reg_reg[104]/NET0131 ,
		\mix1_state_reg[0]/NET0131 ,
		\mix1_state_reg[1]/NET0131 ,
		_w4590_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name3662 (
		\mix1_data_o_reg_reg[68]/NET0131 ,
		\mix1_data_reg_reg[68]/NET0131 ,
		\mix1_state_reg[0]/NET0131 ,
		\mix1_state_reg[1]/NET0131 ,
		_w4591_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name3663 (
		\mix1_data_o_reg_reg[82]/NET0131 ,
		\mix1_data_reg_reg[82]/NET0131 ,
		\mix1_state_reg[0]/NET0131 ,
		\mix1_state_reg[1]/NET0131 ,
		_w4592_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name3664 (
		\mix1_data_o_reg_reg[65]/NET0131 ,
		\mix1_data_reg_reg[65]/NET0131 ,
		\mix1_state_reg[0]/NET0131 ,
		\mix1_state_reg[1]/NET0131 ,
		_w4593_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name3665 (
		\mix1_data_o_reg_reg[66]/NET0131 ,
		\mix1_data_reg_reg[66]/NET0131 ,
		\mix1_state_reg[0]/NET0131 ,
		\mix1_state_reg[1]/NET0131 ,
		_w4594_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name3666 (
		\mix1_data_o_reg_reg[58]/NET0131 ,
		\mix1_data_reg_reg[58]/NET0131 ,
		\mix1_state_reg[0]/NET0131 ,
		\mix1_state_reg[1]/NET0131 ,
		_w4595_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name3667 (
		\mix1_data_o_reg_reg[63]/NET0131 ,
		\mix1_data_reg_reg[63]/NET0131 ,
		\mix1_state_reg[0]/NET0131 ,
		\mix1_state_reg[1]/NET0131 ,
		_w4596_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name3668 (
		\mix1_data_o_reg_reg[36]/NET0131 ,
		\mix1_data_reg_reg[36]/NET0131 ,
		\mix1_state_reg[0]/NET0131 ,
		\mix1_state_reg[1]/NET0131 ,
		_w4597_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name3669 (
		\mix1_data_o_reg_reg[47]/NET0131 ,
		\mix1_data_reg_reg[47]/NET0131 ,
		\mix1_state_reg[0]/NET0131 ,
		\mix1_state_reg[1]/NET0131 ,
		_w4598_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name3670 (
		\mix1_data_o_reg_reg[60]/NET0131 ,
		\mix1_data_reg_reg[60]/NET0131 ,
		\mix1_state_reg[0]/NET0131 ,
		\mix1_state_reg[1]/NET0131 ,
		_w4599_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name3671 (
		\mix1_data_o_reg_reg[86]/NET0131 ,
		\mix1_data_reg_reg[86]/NET0131 ,
		\mix1_state_reg[0]/NET0131 ,
		\mix1_state_reg[1]/NET0131 ,
		_w4600_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name3672 (
		\mix1_data_o_reg_reg[46]/NET0131 ,
		\mix1_data_reg_reg[46]/NET0131 ,
		\mix1_state_reg[0]/NET0131 ,
		\mix1_state_reg[1]/NET0131 ,
		_w4601_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name3673 (
		\mix1_data_o_reg_reg[101]/NET0131 ,
		\mix1_data_reg_reg[101]/NET0131 ,
		\mix1_state_reg[0]/NET0131 ,
		\mix1_state_reg[1]/NET0131 ,
		_w4602_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name3674 (
		\mix1_data_o_reg_reg[44]/NET0131 ,
		\mix1_data_reg_reg[44]/NET0131 ,
		\mix1_state_reg[0]/NET0131 ,
		\mix1_state_reg[1]/NET0131 ,
		_w4603_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name3675 (
		\mix1_data_o_reg_reg[119]/NET0131 ,
		\mix1_data_reg_reg[119]/NET0131 ,
		\mix1_state_reg[0]/NET0131 ,
		\mix1_state_reg[1]/NET0131 ,
		_w4604_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name3676 (
		\mix1_data_o_reg_reg[53]/NET0131 ,
		\mix1_data_reg_reg[53]/NET0131 ,
		\mix1_state_reg[0]/NET0131 ,
		\mix1_state_reg[1]/NET0131 ,
		_w4605_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name3677 (
		\mix1_data_o_reg_reg[100]/NET0131 ,
		\mix1_data_reg_reg[100]/NET0131 ,
		\mix1_state_reg[0]/NET0131 ,
		\mix1_state_reg[1]/NET0131 ,
		_w4606_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name3678 (
		\mix1_data_o_reg_reg[74]/NET0131 ,
		\mix1_data_reg_reg[74]/NET0131 ,
		\mix1_state_reg[0]/NET0131 ,
		\mix1_state_reg[1]/NET0131 ,
		_w4607_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name3679 (
		\mix1_data_o_reg_reg[117]/NET0131 ,
		\mix1_data_reg_reg[117]/NET0131 ,
		\mix1_state_reg[0]/NET0131 ,
		\mix1_state_reg[1]/NET0131 ,
		_w4608_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name3680 (
		\mix1_data_o_reg_reg[67]/NET0131 ,
		\mix1_data_reg_reg[67]/NET0131 ,
		\mix1_state_reg[0]/NET0131 ,
		\mix1_state_reg[1]/NET0131 ,
		_w4609_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name3681 (
		\mix1_data_o_reg_reg[54]/NET0131 ,
		\mix1_data_reg_reg[54]/NET0131 ,
		\mix1_state_reg[0]/NET0131 ,
		\mix1_state_reg[1]/NET0131 ,
		_w4610_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name3682 (
		\mix1_data_o_reg_reg[59]/NET0131 ,
		\mix1_data_reg_reg[59]/NET0131 ,
		\mix1_state_reg[0]/NET0131 ,
		\mix1_state_reg[1]/NET0131 ,
		_w4611_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name3683 (
		\mix1_data_o_reg_reg[51]/NET0131 ,
		\mix1_data_reg_reg[51]/NET0131 ,
		\mix1_state_reg[0]/NET0131 ,
		\mix1_state_reg[1]/NET0131 ,
		_w4612_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name3684 (
		\mix1_data_o_reg_reg[96]/NET0131 ,
		\mix1_data_reg_reg[96]/NET0131 ,
		\mix1_state_reg[0]/NET0131 ,
		\mix1_state_reg[1]/NET0131 ,
		_w4613_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name3685 (
		\mix1_data_o_reg_reg[126]/NET0131 ,
		\mix1_data_reg_reg[126]/NET0131 ,
		\mix1_state_reg[0]/NET0131 ,
		\mix1_state_reg[1]/NET0131 ,
		_w4614_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name3686 (
		\mix1_data_o_reg_reg[57]/NET0131 ,
		\mix1_data_reg_reg[57]/NET0131 ,
		\mix1_state_reg[0]/NET0131 ,
		\mix1_state_reg[1]/NET0131 ,
		_w4615_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name3687 (
		\mix1_data_o_reg_reg[102]/NET0131 ,
		\mix1_data_reg_reg[102]/NET0131 ,
		\mix1_state_reg[0]/NET0131 ,
		\mix1_state_reg[1]/NET0131 ,
		_w4616_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name3688 (
		\mix1_data_o_reg_reg[55]/NET0131 ,
		\mix1_data_reg_reg[55]/NET0131 ,
		\mix1_state_reg[0]/NET0131 ,
		\mix1_state_reg[1]/NET0131 ,
		_w4617_
	);
	LUT3 #(
		.INIT('h06)
	) name3689 (
		\ks1_state_reg[0]/NET0131 ,
		\ks1_state_reg[1]/NET0131 ,
		\ks1_state_reg[2]/NET0131 ,
		_w4618_
	);
	LUT4 #(
		.INIT('h5553)
	) name3690 (
		\key_i[41]_pad ,
		\ks1_key_reg_reg[41]/P0002 ,
		_w938_,
		_w986_,
		_w4619_
	);
	LUT2 #(
		.INIT('h6)
	) name3691 (
		_w2046_,
		_w4619_,
		_w4620_
	);
	LUT4 #(
		.INIT('h2882)
	) name3692 (
		_w929_,
		_w1274_,
		_w2046_,
		_w4619_,
		_w4621_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name3693 (
		\ks1_key_reg_reg[9]/NET0131 ,
		\ks1_state_reg[0]/NET0131 ,
		\ks1_state_reg[1]/NET0131 ,
		\ks1_state_reg[2]/NET0131 ,
		_w4622_
	);
	LUT2 #(
		.INIT('he)
	) name3694 (
		_w4621_,
		_w4622_,
		_w4623_
	);
	LUT4 #(
		.INIT('haaac)
	) name3695 (
		\key_i[108]_pad ,
		\ks1_key_reg_reg[108]/NET0131 ,
		_w938_,
		_w986_,
		_w4624_
	);
	LUT3 #(
		.INIT('h96)
	) name3696 (
		_w1814_,
		_w1816_,
		_w4624_,
		_w4625_
	);
	LUT4 #(
		.INIT('haaac)
	) name3697 (
		\key_i[107]_pad ,
		\ks1_key_reg_reg[107]/NET0131 ,
		_w938_,
		_w986_,
		_w4626_
	);
	LUT2 #(
		.INIT('h6)
	) name3698 (
		_w1809_,
		_w4626_,
		_w4627_
	);
	LUT4 #(
		.INIT('h5553)
	) name3699 (
		\key_i[44]_pad ,
		\ks1_key_reg_reg[44]/P0002 ,
		_w938_,
		_w986_,
		_w4628_
	);
	LUT4 #(
		.INIT('h5553)
	) name3700 (
		\key_i[76]_pad ,
		\ks1_key_reg_reg[76]/P0002 ,
		_w938_,
		_w986_,
		_w4629_
	);
	LUT4 #(
		.INIT('h6996)
	) name3701 (
		_w1814_,
		_w1816_,
		_w4624_,
		_w4629_,
		_w4630_
	);
	LUT4 #(
		.INIT('h9669)
	) name3702 (
		_w1814_,
		_w1816_,
		_w4624_,
		_w4629_,
		_w4631_
	);
	LUT2 #(
		.INIT('h6)
	) name3703 (
		_w4628_,
		_w4630_,
		_w4632_
	);
	LUT4 #(
		.INIT('h2882)
	) name3704 (
		_w929_,
		_w1077_,
		_w4628_,
		_w4630_,
		_w4633_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name3705 (
		\ks1_key_reg_reg[12]/NET0131 ,
		\ks1_state_reg[0]/NET0131 ,
		\ks1_state_reg[1]/NET0131 ,
		\ks1_state_reg[2]/NET0131 ,
		_w4634_
	);
	LUT2 #(
		.INIT('he)
	) name3706 (
		_w4633_,
		_w4634_,
		_w4635_
	);
	LUT4 #(
		.INIT('haaac)
	) name3707 (
		\key_i[75]_pad ,
		\ks1_key_reg_reg[75]/P0002 ,
		_w938_,
		_w986_,
		_w4636_
	);
	LUT3 #(
		.INIT('h96)
	) name3708 (
		_w1809_,
		_w4626_,
		_w4636_,
		_w4637_
	);
	LUT4 #(
		.INIT('haaac)
	) name3709 (
		\key_i[43]_pad ,
		\ks1_key_reg_reg[43]/P0002 ,
		_w938_,
		_w986_,
		_w4638_
	);
	LUT4 #(
		.INIT('h9669)
	) name3710 (
		_w1809_,
		_w4626_,
		_w4636_,
		_w4638_,
		_w4639_
	);
	LUT4 #(
		.INIT('h6996)
	) name3711 (
		_w1809_,
		_w4626_,
		_w4636_,
		_w4638_,
		_w4640_
	);
	LUT4 #(
		.INIT('h2ee2)
	) name3712 (
		\ks1_key_reg_reg[11]/NET0131 ,
		_w929_,
		_w1215_,
		_w4639_,
		_w4641_
	);
	LUT4 #(
		.INIT('haaac)
	) name3713 (
		\key_i[109]_pad ,
		\ks1_key_reg_reg[109]/P0002 ,
		_w938_,
		_w986_,
		_w4642_
	);
	LUT2 #(
		.INIT('h6)
	) name3714 (
		_w1683_,
		_w4642_,
		_w4643_
	);
	LUT4 #(
		.INIT('haaac)
	) name3715 (
		\key_i[77]_pad ,
		\ks1_key_reg_reg[77]/P0002 ,
		_w938_,
		_w986_,
		_w4644_
	);
	LUT3 #(
		.INIT('h96)
	) name3716 (
		_w1683_,
		_w4642_,
		_w4644_,
		_w4645_
	);
	LUT4 #(
		.INIT('haaac)
	) name3717 (
		\key_i[45]_pad ,
		\ks1_key_reg_reg[45]/P0002 ,
		_w938_,
		_w986_,
		_w4646_
	);
	LUT4 #(
		.INIT('h9669)
	) name3718 (
		_w1683_,
		_w4642_,
		_w4644_,
		_w4646_,
		_w4647_
	);
	LUT4 #(
		.INIT('h6996)
	) name3719 (
		_w1683_,
		_w4642_,
		_w4644_,
		_w4646_,
		_w4648_
	);
	LUT4 #(
		.INIT('h2ee2)
	) name3720 (
		\ks1_key_reg_reg[13]/NET0131 ,
		_w929_,
		_w1431_,
		_w4647_,
		_w4649_
	);
	LUT4 #(
		.INIT('haaac)
	) name3721 (
		\key_i[79]_pad ,
		\ks1_key_reg_reg[79]/P0002 ,
		_w938_,
		_w986_,
		_w4650_
	);
	LUT4 #(
		.INIT('h9669)
	) name3722 (
		_w1639_,
		_w1794_,
		_w2196_,
		_w4650_,
		_w4651_
	);
	LUT4 #(
		.INIT('h000e)
	) name3723 (
		_w1585_,
		_w1586_,
		_w1590_,
		_w1591_,
		_w4652_
	);
	LUT3 #(
		.INIT('h0d)
	) name3724 (
		_w1436_,
		_w1592_,
		_w4652_,
		_w4653_
	);
	LUT3 #(
		.INIT('h84)
	) name3725 (
		_w1436_,
		_w1584_,
		_w1600_,
		_w4654_
	);
	LUT4 #(
		.INIT('hf6a3)
	) name3726 (
		_w1600_,
		_w1602_,
		_w1604_,
		_w1608_,
		_w4655_
	);
	LUT3 #(
		.INIT('h69)
	) name3727 (
		_w4653_,
		_w4654_,
		_w4655_,
		_w4656_
	);
	LUT4 #(
		.INIT('haaac)
	) name3728 (
		\key_i[47]_pad ,
		\ks1_key_reg_reg[47]/P0002 ,
		_w938_,
		_w986_,
		_w4657_
	);
	LUT2 #(
		.INIT('h6)
	) name3729 (
		_w4651_,
		_w4657_,
		_w4658_
	);
	LUT4 #(
		.INIT('h2882)
	) name3730 (
		_w929_,
		_w1528_,
		_w4651_,
		_w4657_,
		_w4659_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name3731 (
		\ks1_key_reg_reg[15]/NET0131 ,
		\ks1_state_reg[0]/NET0131 ,
		\ks1_state_reg[1]/NET0131 ,
		\ks1_state_reg[2]/NET0131 ,
		_w4660_
	);
	LUT2 #(
		.INIT('he)
	) name3732 (
		_w4659_,
		_w4660_,
		_w4661_
	);
	assign \_al_n0  = 1'b0;
	assign \_al_n1  = 1'b1;
	assign \g27929/_0_  = _w993_ ;
	assign \g27942/_3_  = _w1613_ ;
	assign \g27943/_3_  = _w1618_ ;
	assign \g27944/_3_  = _w1626_ ;
	assign \g27945/_0_  = _w1649_ ;
	assign \g27995/_0_  = _w1667_ ;
	assign \g27998/_0_  = _w992_ ;
	assign \g28019/_0_  = _w1680_ ;
	assign \g28020/_0_  = _w1691_ ;
	assign \g28021/_0_  = _w1697_ ;
	assign \g28022/_0_  = _w1701_ ;
	assign \g28023/_0_  = _w1708_ ;
	assign \g28024/_0_  = _w1712_ ;
	assign \g28025/_0_  = _w1719_ ;
	assign \g28026/_0_  = _w1726_ ;
	assign \g28027/_0_  = _w1731_ ;
	assign \g28028/_0_  = _w1735_ ;
	assign \g28029/_0_  = _w1739_ ;
	assign \g28030/_0_  = _w1742_ ;
	assign \g28031/_0_  = _w1747_ ;
	assign \g28032/_0_  = _w1751_ ;
	assign \g28033/_0_  = _w1756_ ;
	assign \g28034/_0_  = _w1760_ ;
	assign \g28044/_0_  = _w1765_ ;
	assign \g28045/_0_  = _w1768_ ;
	assign \g28046/_0_  = _w1773_ ;
	assign \g28047/_0_  = _w1776_ ;
	assign \g28048/_0_  = _w1780_ ;
	assign \g28049/_0_  = _w1783_ ;
	assign \g28050/_0_  = _w1787_ ;
	assign \g28051/_0_  = _w1790_ ;
	assign \g28151/_0_  = _w990_ ;
	assign \g28177/_0_  = _w1792_ ;
	assign \g28178/_0_  = _w1802_ ;
	assign \g28179/_0_  = _w1807_ ;
	assign \g28180/_0_  = _w1813_ ;
	assign \g28181/_0_  = _w1821_ ;
	assign \g28182/_0_  = _w1826_ ;
	assign \g28183/_0_  = _w1831_ ;
	assign \g28184/_0_  = _w1835_ ;
	assign \g28185/_0_  = _w1840_ ;
	assign \g28186/_0_  = _w1845_ ;
	assign \g28187/_0_  = _w1853_ ;
	assign \g28188/_0_  = _w1856_ ;
	assign \g28189/_0_  = _w1861_ ;
	assign \g28190/_0_  = _w1864_ ;
	assign \g28191/_0_  = _w1868_ ;
	assign \g28192/_0_  = _w1873_ ;
	assign \g28193/_0_  = _w1878_ ;
	assign \g28194/_0_  = _w1883_ ;
	assign \g28195/_0_  = _w1887_ ;
	assign \g28196/_0_  = _w1892_ ;
	assign \g28197/_0_  = _w1897_ ;
	assign \g28198/_0_  = _w1900_ ;
	assign \g28199/_0_  = _w1905_ ;
	assign \g28200/_0_  = _w1909_ ;
	assign \g28201/_0_  = _w1914_ ;
	assign \g28202/_0_  = _w1919_ ;
	assign \g28203/_0_  = _w1926_ ;
	assign \g28253/_0_  = _w1930_ ;
	assign \g28254/_0_  = _w1933_ ;
	assign \g28255/_0_  = _w1937_ ;
	assign \g28256/_0_  = _w1941_ ;
	assign \g28257/_0_  = _w1944_ ;
	assign \g28258/_0_  = _w1945_ ;
	assign \g28259/_0_  = _w1946_ ;
	assign \g28260/_0_  = _w1950_ ;
	assign \g28261/_0_  = _w1951_ ;
	assign \g28262/_0_  = _w1955_ ;
	assign \g28263/_0_  = _w1956_ ;
	assign \g28264/_0_  = _w1957_ ;
	assign \g28265/_0_  = _w1958_ ;
	assign \g28266/_0_  = _w1962_ ;
	assign \g28267/_0_  = _w1965_ ;
	assign \g28268/_0_  = _w1969_ ;
	assign \g28269/_0_  = _w1973_ ;
	assign \g28270/_0_  = _w1977_ ;
	assign \g28271/_0_  = _w1980_ ;
	assign \g28272/_0_  = _w1984_ ;
	assign \g28273/_0_  = _w1988_ ;
	assign \g28274/_0_  = _w1992_ ;
	assign \g28275/_0_  = _w2000_ ;
	assign \g28276/_0_  = _w2006_ ;
	assign \g28277/_0_  = _w2014_ ;
	assign \g28278/_0_  = _w2022_ ;
	assign \g28279/_0_  = _w2028_ ;
	assign \g28384/_2_  = _w2030_ ;
	assign \g28385/_2_  = _w2031_ ;
	assign \g28388/_2_  = _w2033_ ;
	assign \g28389/_2_  = _w2034_ ;
	assign \g28394/_2_  = _w2036_ ;
	assign \g28395/_2_  = _w2037_ ;
	assign \g28401/_2_  = _w2039_ ;
	assign \g28402/_2_  = _w2040_ ;
	assign \g28403/_0_  = _w2047_ ;
	assign \g28404/_0_  = _w2048_ ;
	assign \g28408/_0_  = _w1666_ ;
	assign \g28410/_0_  = _w1644_ ;
	assign \g28440/_0_  = _w2053_ ;
	assign \g28441/_0_  = _w2058_ ;
	assign \g28442/_0_  = _w2063_ ;
	assign \g28443/_0_  = _w2068_ ;
	assign \g28444/_0_  = _w2070_ ;
	assign \g28445/_0_  = _w2073_ ;
	assign \g28446/_0_  = _w2078_ ;
	assign \g28447/_0_  = _w2083_ ;
	assign \g28448/_0_  = _w2088_ ;
	assign \g28449/_0_  = _w2093_ ;
	assign \g28450/_0_  = _w2098_ ;
	assign \g28451/_0_  = _w2103_ ;
	assign \g28452/_0_  = _w2111_ ;
	assign \g28453/_0_  = _w2119_ ;
	assign \g28538/_0_  = _w2123_ ;
	assign \g28539/_0_  = _w2127_ ;
	assign \g28540/_0_  = _w2128_ ;
	assign \g28541/_0_  = _w2129_ ;
	assign \g28542/_0_  = _w2130_ ;
	assign \g28543/_0_  = _w2131_ ;
	assign \g28544/_0_  = _w2135_ ;
	assign \g28545/_0_  = _w2136_ ;
	assign \g28546/_0_  = _w2137_ ;
	assign \g28547/_0_  = _w2138_ ;
	assign \g28548/_0_  = _w2139_ ;
	assign \g28549/_0_  = _w2140_ ;
	assign \g28550/_0_  = _w2141_ ;
	assign \g28551/_0_  = _w2142_ ;
	assign \g28552/_0_  = _w2143_ ;
	assign \g28557/_0_  = _w2147_ ;
	assign \g28558/_0_  = _w2151_ ;
	assign \g28563/_0_  = _w2155_ ;
	assign \g28564/_0_  = _w2159_ ;
	assign \g28565/_0_  = _w2163_ ;
	assign \g28566/_0_  = _w2171_ ;
	assign \g28567/_0_  = _w2179_ ;
	assign \g28625/_2_  = _w2180_ ;
	assign \g28626/_2_  = _w2181_ ;
	assign \g28633/_2_  = _w2182_ ;
	assign \g28639/_2_  = _w2183_ ;
	assign \g28655/_2_  = _w2184_ ;
	assign \g28656/_2_  = _w2185_ ;
	assign \g28657/_2_  = _w2186_ ;
	assign \g28660/_2_  = _w2187_ ;
	assign \g28661/_2_  = _w2188_ ;
	assign \g28662/_2_  = _w2189_ ;
	assign \g28666/_2_  = _w2190_ ;
	assign \g28667/_2_  = _w2191_ ;
	assign \g28668/_2_  = _w2192_ ;
	assign \g28678/_2_  = _w2193_ ;
	assign \g28679/_2_  = _w2194_ ;
	assign \g28680/_2_  = _w2195_ ;
	assign \g28690/_0_  = _w2197_ ;
	assign \g28710/_0_  = _w1642_ ;
	assign \g28716/_0_  = _w2198_ ;
	assign \g28795/_0_  = _w2201_ ;
	assign \g28796/_0_  = _w2202_ ;
	assign \g28798/_0_  = _w2203_ ;
	assign \g28799/_0_  = _w2204_ ;
	assign \g28800/_0_  = _w2207_ ;
	assign \g28801/_0_  = _w2210_ ;
	assign \g28804/_0_  = _w1592_ ;
	assign \g28825/_2_  = _w2211_ ;
	assign \g28826/_2_  = _w2212_ ;
	assign \g28830/_2_  = _w2213_ ;
	assign \g28834/_2_  = _w2214_ ;
	assign \g28842/_2_  = _w2217_ ;
	assign \g28843/_2_  = _w2220_ ;
	assign \g28845/_2_  = _w2223_ ;
	assign \g28848/_2_  = _w2226_ ;
	assign \g28890/_0_  = _w2045_ ;
	assign \g28936/_0_  = _w2227_ ;
	assign \g28982/_0_  = _w2228_ ;
	assign \g29050/_0_  = _w2451_ ;
	assign \g29051/_0_  = _w2533_ ;
	assign \g29052/_0_  = _w2586_ ;
	assign \g29053/_0_  = _w2605_ ;
	assign \g29054/_0_  = _w2614_ ;
	assign \g29055/_0_  = _w2624_ ;
	assign \g29056/_0_  = _w2629_ ;
	assign \g29057/_0_  = _w2636_ ;
	assign \g29058/_0_  = _w2638_ ;
	assign \g29059/_0_  = _w2643_ ;
	assign \g29060/_0_  = _w2649_ ;
	assign \g29061/_0_  = _w2650_ ;
	assign \g29328/_0_  = _w2656_ ;
	assign \g29329/_0_  = _w2659_ ;
	assign \g29330/_0_  = _w2661_ ;
	assign \g29331/_0_  = _w2668_ ;
	assign \g29332/_0_  = _w2675_ ;
	assign \g29333/_0_  = _w2678_ ;
	assign \g29334/_0_  = _w2683_ ;
	assign \g29335/_0_  = _w2689_ ;
	assign \g29336/_0_  = _w2693_ ;
	assign \g29337/_0_  = _w2695_ ;
	assign \g29338/_0_  = _w2697_ ;
	assign \g29339/_0_  = _w2702_ ;
	assign \g29340/_0_  = _w2704_ ;
	assign \g29341/_0_  = _w2706_ ;
	assign \g29342/_0_  = _w2707_ ;
	assign \g29343/_0_  = _w2708_ ;
	assign \g29344/_0_  = _w2709_ ;
	assign \g29345/_0_  = _w2710_ ;
	assign \g29346/_0_  = _w2711_ ;
	assign \g29347/_0_  = _w2712_ ;
	assign \g29348/_0_  = _w2713_ ;
	assign \g29349/_0_  = _w2716_ ;
	assign \g29350/_0_  = _w2719_ ;
	assign \g29351/_0_  = _w2720_ ;
	assign \g29352/_0_  = _w2723_ ;
	assign \g29353/_0_  = _w2724_ ;
	assign \g29354/_0_  = _w2725_ ;
	assign \g29355/_0_  = _w2726_ ;
	assign \g29356/_0_  = _w2727_ ;
	assign \g29357/_0_  = _w2728_ ;
	assign \g29358/_0_  = _w2729_ ;
	assign \g29359/_0_  = _w2730_ ;
	assign \g29360/_0_  = _w2733_ ;
	assign \g29361/_0_  = _w2736_ ;
	assign \g29362/_0_  = _w2737_ ;
	assign \g29363/_0_  = _w2740_ ;
	assign \g29364/_0_  = _w2741_ ;
	assign \g29365/_0_  = _w2742_ ;
	assign \g29366/_0_  = _w2746_ ;
	assign \g29367/_0_  = _w2749_ ;
	assign \g29395/_0_  = _w2772_ ;
	assign \g29396/_0_  = _w2773_ ;
	assign \g29453/_0_  = _w2788_ ;
	assign \g29454/_0_  = _w2798_ ;
	assign \g29455/_0_  = _w2808_ ;
	assign \g29456/_0_  = _w2818_ ;
	assign \g29457/_0_  = _w2828_ ;
	assign \g29458/_0_  = _w2838_ ;
	assign \g29459/_0_  = _w2848_ ;
	assign \g29460/_0_  = _w2858_ ;
	assign \g29461/_0_  = _w2868_ ;
	assign \g29462/_0_  = _w2878_ ;
	assign \g29463/_0_  = _w2888_ ;
	assign \g29464/_0_  = _w2898_ ;
	assign \g29465/_0_  = _w2908_ ;
	assign \g29466/_0_  = _w2918_ ;
	assign \g29467/_0_  = _w2928_ ;
	assign \g29468/_0_  = _w2938_ ;
	assign \g29469/_0_  = _w2948_ ;
	assign \g29470/_0_  = _w2958_ ;
	assign \g29471/_0_  = _w2968_ ;
	assign \g29472/_0_  = _w2978_ ;
	assign \g29473/_0_  = _w2988_ ;
	assign \g29474/_0_  = _w2998_ ;
	assign \g29475/_0_  = _w3008_ ;
	assign \g29476/_0_  = _w3018_ ;
	assign \g29477/_0_  = _w3028_ ;
	assign \g29478/_0_  = _w3038_ ;
	assign \g29479/_0_  = _w3048_ ;
	assign \g29480/_0_  = _w3058_ ;
	assign \g29481/_0_  = _w3068_ ;
	assign \g29482/_0_  = _w3078_ ;
	assign \g29483/_0_  = _w3088_ ;
	assign \g29484/_0_  = _w3098_ ;
	assign \g29485/_0_  = _w3108_ ;
	assign \g29486/_0_  = _w3118_ ;
	assign \g29487/_0_  = _w3128_ ;
	assign \g29488/_0_  = _w3138_ ;
	assign \g29489/_0_  = _w3148_ ;
	assign \g29490/_0_  = _w3158_ ;
	assign \g29491/_0_  = _w3168_ ;
	assign \g29492/_0_  = _w3178_ ;
	assign \g29493/_0_  = _w3188_ ;
	assign \g29494/_0_  = _w3198_ ;
	assign \g29495/_0_  = _w3208_ ;
	assign \g29496/_0_  = _w3218_ ;
	assign \g29497/_0_  = _w3228_ ;
	assign \g29498/_0_  = _w3238_ ;
	assign \g29499/_0_  = _w3248_ ;
	assign \g29500/_0_  = _w3258_ ;
	assign \g29501/_0_  = _w3268_ ;
	assign \g29502/_0_  = _w3278_ ;
	assign \g29503/_0_  = _w3288_ ;
	assign \g29504/_0_  = _w3298_ ;
	assign \g29505/_0_  = _w3308_ ;
	assign \g29506/_0_  = _w3318_ ;
	assign \g29507/_0_  = _w3328_ ;
	assign \g29508/_0_  = _w3338_ ;
	assign \g29509/_0_  = _w3348_ ;
	assign \g29510/_0_  = _w3358_ ;
	assign \g29511/_0_  = _w3368_ ;
	assign \g29512/_0_  = _w3378_ ;
	assign \g29513/_0_  = _w3388_ ;
	assign \g29514/_0_  = _w3398_ ;
	assign \g29515/_0_  = _w3408_ ;
	assign \g29516/_0_  = _w3418_ ;
	assign \g29517/_0_  = _w3428_ ;
	assign \g29518/_0_  = _w3438_ ;
	assign \g29519/_0_  = _w3448_ ;
	assign \g29520/_0_  = _w3458_ ;
	assign \g29521/_0_  = _w3468_ ;
	assign \g29522/_0_  = _w3478_ ;
	assign \g29523/_0_  = _w3488_ ;
	assign \g29524/_0_  = _w3502_ ;
	assign \g29525/_0_  = _w3512_ ;
	assign \g29526/_0_  = _w3522_ ;
	assign \g29527/_0_  = _w3536_ ;
	assign \g29528/_0_  = _w3546_ ;
	assign \g29529/_0_  = _w3556_ ;
	assign \g29530/_0_  = _w3566_ ;
	assign \g29531/_0_  = _w3576_ ;
	assign \g29532/_0_  = _w3586_ ;
	assign \g29533/_0_  = _w3596_ ;
	assign \g29534/_0_  = _w3606_ ;
	assign \g29535/_0_  = _w3616_ ;
	assign \g29536/_0_  = _w3626_ ;
	assign \g29537/_0_  = _w3636_ ;
	assign \g29538/_0_  = _w3646_ ;
	assign \g29539/_0_  = _w3656_ ;
	assign \g29540/_0_  = _w3666_ ;
	assign \g29541/_0_  = _w3676_ ;
	assign \g29542/_0_  = _w3686_ ;
	assign \g29543/_0_  = _w3696_ ;
	assign \g29544/_0_  = _w3706_ ;
	assign \g29545/_0_  = _w3716_ ;
	assign \g29546/_0_  = _w3726_ ;
	assign \g29547/_0_  = _w3736_ ;
	assign \g29548/_0_  = _w3746_ ;
	assign \g29549/_0_  = _w3756_ ;
	assign \g29550/_0_  = _w3766_ ;
	assign \g29551/_0_  = _w3776_ ;
	assign \g29552/_0_  = _w3786_ ;
	assign \g29553/_0_  = _w3796_ ;
	assign \g29554/_0_  = _w3806_ ;
	assign \g29555/_0_  = _w3816_ ;
	assign \g29556/_0_  = _w3826_ ;
	assign \g29557/_0_  = _w3836_ ;
	assign \g29558/_0_  = _w3846_ ;
	assign \g29559/_0_  = _w3856_ ;
	assign \g29560/_0_  = _w3866_ ;
	assign \g29561/_0_  = _w3876_ ;
	assign \g29562/_0_  = _w3886_ ;
	assign \g29563/_0_  = _w3896_ ;
	assign \g29564/_0_  = _w3906_ ;
	assign \g29565/_0_  = _w3916_ ;
	assign \g29566/_0_  = _w3926_ ;
	assign \g29567/_0_  = _w3936_ ;
	assign \g29568/_0_  = _w3946_ ;
	assign \g29569/_0_  = _w3956_ ;
	assign \g29570/_0_  = _w3966_ ;
	assign \g29571/_0_  = _w3976_ ;
	assign \g29572/_0_  = _w3986_ ;
	assign \g29573/_0_  = _w3996_ ;
	assign \g29574/_0_  = _w4006_ ;
	assign \g29575/_0_  = _w4016_ ;
	assign \g29576/_0_  = _w4026_ ;
	assign \g29577/_0_  = _w4036_ ;
	assign \g29578/_0_  = _w4046_ ;
	assign \g29579/_0_  = _w4056_ ;
	assign \g29580/_0_  = _w4066_ ;
	assign \g29582/_0_  = _w4067_ ;
	assign \g29583/_0_  = _w4068_ ;
	assign \g29584/_0_  = _w4069_ ;
	assign \g29585/_0_  = _w4070_ ;
	assign \g29586/_0_  = _w4073_ ;
	assign \g29587/_0_  = _w4076_ ;
	assign \g29588/_0_  = _w4077_ ;
	assign \g29589/_0_  = _w4080_ ;
	assign \g29590/_0_  = _w4081_ ;
	assign \g29591/_0_  = _w4082_ ;
	assign \g29592/_0_  = _w4083_ ;
	assign \g29593/_0_  = _w4084_ ;
	assign \g29634/_0_  = _w4092_ ;
	assign \g29635/_0_  = _w4100_ ;
	assign \g29636/_0_  = _w4108_ ;
	assign \g29637/_0_  = _w4116_ ;
	assign \g29645/_0_  = _w4130_ ;
	assign \g29646/_0_  = _w4144_ ;
	assign \g29647/_0_  = _w4157_ ;
	assign \g29824/_0_  = _w4159_ ;
	assign \g29828/_0_  = _w4162_ ;
	assign \g29832/_0_  = _w4166_ ;
	assign \g29836/_0_  = _w4167_ ;
	assign \g29837/_0_  = _w4170_ ;
	assign \g29838/_0_  = _w4173_ ;
	assign \g29839/_0_  = _w4174_ ;
	assign \g29840/_0_  = _w4175_ ;
	assign \g29841/_0_  = _w4176_ ;
	assign \g29842/_0_  = _w4179_ ;
	assign \g29843/_0_  = _w4180_ ;
	assign \g29844/_0_  = _w4181_ ;
	assign \g29845/_0_  = _w4182_ ;
	assign \g29846/_0_  = _w4185_ ;
	assign \g29847/_0_  = _w4186_ ;
	assign \g29848/_0_  = _w4187_ ;
	assign \g29849/_0_  = _w4190_ ;
	assign \g29850/_0_  = _w4191_ ;
	assign \g29851/_0_  = _w4192_ ;
	assign \g29852/_0_  = _w4193_ ;
	assign \g29853/_0_  = _w4196_ ;
	assign \g29854/_0_  = _w4199_ ;
	assign \g29855/_0_  = _w4200_ ;
	assign \g29856/_0_  = _w4201_ ;
	assign \g29857/_0_  = _w4202_ ;
	assign \g29858/_0_  = _w4205_ ;
	assign \g29859/_0_  = _w4206_ ;
	assign \g29860/_0_  = _w4207_ ;
	assign \g29861/_0_  = _w4208_ ;
	assign \g29862/_0_  = _w4211_ ;
	assign \g29863/_0_  = _w4212_ ;
	assign \g29864/_0_  = _w4213_ ;
	assign \g29865/_0_  = _w4216_ ;
	assign \g29866/_0_  = _w4217_ ;
	assign \g29867/_0_  = _w4218_ ;
	assign \g29868/_0_  = _w4220_ ;
	assign \g30081/_0_  = _w4221_ ;
	assign \g30082/_0_  = _w4224_ ;
	assign \g30083/_0_  = _w4225_ ;
	assign \g30084/_0_  = _w4226_ ;
	assign \g30085/_0_  = _w4227_ ;
	assign \g30086/_0_  = _w4228_ ;
	assign \g30087/_0_  = _w4231_ ;
	assign \g30088/_0_  = _w4232_ ;
	assign \g30089/_0_  = _w4233_ ;
	assign \g30090/_0_  = _w4236_ ;
	assign \g30091/_0_  = _w4239_ ;
	assign \g30092/_0_  = _w4240_ ;
	assign \g30093/_0_  = _w4241_ ;
	assign \g30094/_0_  = _w4244_ ;
	assign \g30095/_0_  = _w4245_ ;
	assign \g30096/_0_  = _w4246_ ;
	assign \g30135/_0_  = _w4247_ ;
	assign \g30137/_0_  = _w4248_ ;
	assign \g30164/_0_  = _w4129_ ;
	assign \g30165/_0_  = _w4143_ ;
	assign \g30166/_0_  = _w4156_ ;
	assign \g30167/_0_  = _w4091_ ;
	assign \g30168/_0_  = _w4099_ ;
	assign \g30169/_0_  = _w4107_ ;
	assign \g30170/_0_  = _w4115_ ;
	assign \g30231/_0_  = _w4249_ ;
	assign \g30232/_0_  = _w4250_ ;
	assign \g30233/_0_  = _w4251_ ;
	assign \g30234/_0_  = _w4254_ ;
	assign \g30235/_0_  = _w4255_ ;
	assign \g30236/_0_  = _w4256_ ;
	assign \g30237/_0_  = _w4257_ ;
	assign \g30238/_0_  = _w4260_ ;
	assign \g30286/_0_  = _w4274_ ;
	assign \g30287/_0_  = _w4288_ ;
	assign \g30288/_0_  = _w4302_ ;
	assign \g30289/_0_  = _w4309_ ;
	assign \g30290/_0_  = _w4316_ ;
	assign \g30291/_0_  = _w4323_ ;
	assign \g30292/_0_  = _w4330_ ;
	assign \g30293/_0_  = _w4337_ ;
	assign \g30294/_0_  = _w4351_ ;
	assign \g30295/_0_  = _w4365_ ;
	assign \g30296/_0_  = _w4379_ ;
	assign \g30297/_0_  = _w4393_ ;
	assign \g30298/_0_  = _w4407_ ;
	assign \g30299/_0_  = _w4421_ ;
	assign \g30300/_0_  = _w4435_ ;
	assign \g30301/_0_  = _w4449_ ;
	assign \g30303/_0_  = _w4450_ ;
	assign \g30304/_0_  = _w4451_ ;
	assign \g30305/_0_  = _w4452_ ;
	assign \g30306/_0_  = _w4453_ ;
	assign \g30307/_0_  = _w4454_ ;
	assign \g30308/_0_  = _w4455_ ;
	assign \g30309/_0_  = _w4456_ ;
	assign \g30310/_0_  = _w4457_ ;
	assign \g30311/_0_  = _w4458_ ;
	assign \g30312/_0_  = _w4459_ ;
	assign \g30313/_0_  = _w4460_ ;
	assign \g30314/_0_  = _w4461_ ;
	assign \g30315/_0_  = _w4462_ ;
	assign \g30316/_0_  = _w4463_ ;
	assign \g30317/_0_  = _w4464_ ;
	assign \g30318/_0_  = _w2770_ ;
	assign \g30319/_0_  = _w4465_ ;
	assign \g30481/_0_  = _w4466_ ;
	assign \g30482/_0_  = _w4467_ ;
	assign \g30483/_0_  = _w4470_ ;
	assign \g30484/_0_  = _w4471_ ;
	assign \g30493/_0_  = _w4089_ ;
	assign \g30495/_0_  = _w4105_ ;
	assign \g30536/_0_  = _w4127_ ;
	assign \g30537/_0_  = _w4141_ ;
	assign \g30538/_0_  = _w4154_ ;
	assign \g30735/_0_  = _w2768_ ;
	assign \g30927/_0_  = _w4153_ ;
	assign \g30928/_0_  = _w4125_ ;
	assign \g30929/_0_  = _w4139_ ;
	assign \g30971/_0_  = _w4111_ ;
	assign \g30972/_0_  = _w4087_ ;
	assign \g30973/_0_  = _w4095_ ;
	assign \g30974/_0_  = _w4103_ ;
	assign \g31129/_0_  = _w4306_ ;
	assign \g31130/_0_  = _w4313_ ;
	assign \g31131/_0_  = _w4320_ ;
	assign \g31132/_0_  = _w4327_ ;
	assign \g31133/_0_  = _w4334_ ;
	assign \g31134/_0_  = _w4270_ ;
	assign \g31135/_0_  = _w4347_ ;
	assign \g31136/_0_  = _w4361_ ;
	assign \g31137/_0_  = _w4375_ ;
	assign \g31138/_0_  = _w4389_ ;
	assign \g31139/_0_  = _w4284_ ;
	assign \g31140/_0_  = _w4403_ ;
	assign \g31141/_0_  = _w4417_ ;
	assign \g31142/_0_  = _w4431_ ;
	assign \g31143/_0_  = _w4445_ ;
	assign \g31144/_0_  = _w4298_ ;
	assign \g31352/_0_  = _w4304_ ;
	assign \g31353/_0_  = _w4360_ ;
	assign \g31354/_0_  = _w4269_ ;
	assign \g31355/_0_  = _w4416_ ;
	assign \g31356/_0_  = _w4311_ ;
	assign \g31357/_0_  = _w4318_ ;
	assign \g31358/_0_  = _w4325_ ;
	assign \g31359/_0_  = _w4332_ ;
	assign \g31360/_0_  = _w4346_ ;
	assign \g31361/_0_  = _w4374_ ;
	assign \g31362/_0_  = _w4402_ ;
	assign \g31363/_0_  = _w4430_ ;
	assign \g31364/_0_  = _w4444_ ;
	assign \g31365/_0_  = _w4388_ ;
	assign \g31366/_0_  = _w4283_ ;
	assign \g31367/_0_  = _w4297_ ;
	assign \g31706/_0_  = _w4472_ ;
	assign \g32001/_0_  = _w4473_ ;
	assign \g32008/_0_  = _w4475_ ;
	assign \g32009/_0_  = _w4477_ ;
	assign \g32010/_0_  = _w4479_ ;
	assign \g32011/_0_  = _w4480_ ;
	assign \g32118/_0_  = _w4494_ ;
	assign \g33261/_0_  = _w4499_ ;
	assign \g33262/_0_  = _w4500_ ;
	assign \g33263/_0_  = _w4501_ ;
	assign \g33264/_0_  = _w4505_ ;
	assign \g33265/_0_  = _w4508_ ;
	assign \g33266/_0_  = _w4514_ ;
	assign \g33450/_0_  = _w4515_ ;
	assign \g33451/_0_  = _w4516_ ;
	assign \g33453/_0_  = _w4518_ ;
	assign \g33485/_0_  = _w4519_ ;
	assign \g33679/_2_  = _w4520_ ;
	assign \g34838/_2_  = _w4521_ ;
	assign \g34971/_0_  = _w4522_ ;
	assign \g34972/_0_  = _w4523_ ;
	assign \g34973/_0_  = _w4524_ ;
	assign \g34974/_0_  = _w4525_ ;
	assign \g34975/_0_  = _w4526_ ;
	assign \g34976/_0_  = _w4527_ ;
	assign \g34977/_0_  = _w4528_ ;
	assign \g34978/_0_  = _w4529_ ;
	assign \g34979/_0_  = _w4530_ ;
	assign \g34980/_0_  = _w4531_ ;
	assign \g34981/_0_  = _w4532_ ;
	assign \g34982/_0_  = _w4533_ ;
	assign \g34983/_0_  = _w4534_ ;
	assign \g34984/_0_  = _w4535_ ;
	assign \g34985/_0_  = _w4536_ ;
	assign \g34986/_0_  = _w4537_ ;
	assign \g34987/_0_  = _w4538_ ;
	assign \g34988/_0_  = _w4539_ ;
	assign \g34989/_0_  = _w4540_ ;
	assign \g34990/_0_  = _w4541_ ;
	assign \g34991/_0_  = _w4542_ ;
	assign \g34992/_0_  = _w4543_ ;
	assign \g34993/_0_  = _w4544_ ;
	assign \g34994/_0_  = _w4545_ ;
	assign \g34995/_0_  = _w4546_ ;
	assign \g34996/_0_  = _w4547_ ;
	assign \g34997/_0_  = _w4548_ ;
	assign \g34998/_0_  = _w4549_ ;
	assign \g34999/_0_  = _w4550_ ;
	assign \g35000/_0_  = _w4551_ ;
	assign \g35001/_0_  = _w4552_ ;
	assign \g35002/_0_  = _w4553_ ;
	assign \g35003/_0_  = _w4554_ ;
	assign \g35004/_0_  = _w4555_ ;
	assign \g35005/_0_  = _w4556_ ;
	assign \g35006/_0_  = _w4557_ ;
	assign \g35007/_0_  = _w4558_ ;
	assign \g35008/_0_  = _w4559_ ;
	assign \g35009/_0_  = _w4560_ ;
	assign \g35010/_0_  = _w4561_ ;
	assign \g35011/_0_  = _w4562_ ;
	assign \g35012/_0_  = _w4563_ ;
	assign \g35013/_0_  = _w4564_ ;
	assign \g35014/_0_  = _w4565_ ;
	assign \g35015/_0_  = _w4566_ ;
	assign \g35016/_0_  = _w4567_ ;
	assign \g35017/_0_  = _w4568_ ;
	assign \g35018/_0_  = _w4569_ ;
	assign \g35019/_0_  = _w4570_ ;
	assign \g35020/_0_  = _w4571_ ;
	assign \g35021/_0_  = _w4572_ ;
	assign \g35022/_0_  = _w4573_ ;
	assign \g35023/_0_  = _w4574_ ;
	assign \g35024/_0_  = _w4575_ ;
	assign \g35025/_0_  = _w4576_ ;
	assign \g35026/_0_  = _w4577_ ;
	assign \g35027/_0_  = _w4578_ ;
	assign \g35028/_0_  = _w4579_ ;
	assign \g35029/_0_  = _w4580_ ;
	assign \g35030/_0_  = _w4581_ ;
	assign \g35031/_0_  = _w4582_ ;
	assign \g35032/_0_  = _w4583_ ;
	assign \g35033/_0_  = _w4584_ ;
	assign \g35034/_0_  = _w4585_ ;
	assign \g35035/_0_  = _w4586_ ;
	assign \g35036/_0_  = _w4587_ ;
	assign \g35037/_0_  = _w4588_ ;
	assign \g35038/_0_  = _w4589_ ;
	assign \g35039/_0_  = _w4590_ ;
	assign \g35040/_0_  = _w4591_ ;
	assign \g35041/_0_  = _w4592_ ;
	assign \g35042/_0_  = _w4593_ ;
	assign \g35043/_0_  = _w4594_ ;
	assign \g35044/_0_  = _w4595_ ;
	assign \g35045/_0_  = _w4596_ ;
	assign \g35046/_0_  = _w4597_ ;
	assign \g35047/_0_  = _w4598_ ;
	assign \g35048/_0_  = _w4599_ ;
	assign \g35049/_0_  = _w4600_ ;
	assign \g35050/_0_  = _w4601_ ;
	assign \g35051/_0_  = _w4602_ ;
	assign \g35052/_0_  = _w4603_ ;
	assign \g35053/_0_  = _w4604_ ;
	assign \g35054/_0_  = _w4605_ ;
	assign \g35055/_0_  = _w4606_ ;
	assign \g35056/_0_  = _w4607_ ;
	assign \g35057/_0_  = _w4608_ ;
	assign \g35058/_0_  = _w4609_ ;
	assign \g35059/_0_  = _w4610_ ;
	assign \g35060/_0_  = _w4611_ ;
	assign \g35061/_0_  = _w4612_ ;
	assign \g35062/_0_  = _w4613_ ;
	assign \g35063/_0_  = _w4614_ ;
	assign \g35064/_0_  = _w4615_ ;
	assign \g35065/_0_  = _w4616_ ;
	assign \g35066/_0_  = _w4617_ ;
	assign \g35538/_0_  = _w4618_ ;
	assign \g35956/_0_  = _w1677_ ;
	assign \g36298/_1_  = _w4492_ ;
	assign \g36324/_0_  = _w929_ ;
	assign \g36375/_0_  = _w1669_ ;
	assign \g38269/_0_  = _w4623_ ;
	assign \g38473/_0_  = _w4625_ ;
	assign \g38501/_0_  = _w4627_ ;
	assign \g38569/_0_  = _w4635_ ;
	assign \g38629/_0_  = _w4641_ ;
	assign \g38721_dup/_3_  = _w4643_ ;
	assign \g38735/_0_  = _w4649_ ;
	assign \g38753/_0_  = _w1064_ ;
	assign \g38849/_3_  = _w1588_ ;
	assign \g39071/_0_  = _w4648_ ;
	assign \g39073/_0_  = _w4645_ ;
	assign \g39077/_0_  = _w4632_ ;
	assign \g39080/_0_  = _w4631_ ;
	assign \g39135/_0_  = _w4640_ ;
	assign \g39138/_0_  = _w4637_ ;
	assign \g39182/_0_  = _w4651_ ;
	assign \g39197/_3_  = _w4620_ ;
	assign \g39207/_3_  = _w988_ ;
	assign \g39241/_0_  = _w4656_ ;
	assign \g39272/_0_  = _w4661_ ;
	assign \g39307/_0_  = _w1609_ ;
	assign \g39308/_0_  = _w1605_ ;
	assign \g39361/_0_  = _w1624_ ;
	assign \g39494/_0_  = _w2236_ ;
	assign \g39558/_0_  = _w1663_ ;
	assign \g39575/_0_  = _w4658_ ;
	assign \g39583/_0_  = _w1646_ ;
endmodule;