module top( \clgen_cnt_reg[0]/NET0131  , \clgen_cnt_reg[10]/NET0131  , \clgen_cnt_reg[11]/NET0131  , \clgen_cnt_reg[12]/NET0131  , \clgen_cnt_reg[13]/NET0131  , \clgen_cnt_reg[14]/NET0131  , \clgen_cnt_reg[15]/NET0131  , \clgen_cnt_reg[1]/NET0131  , \clgen_cnt_reg[2]/NET0131  , \clgen_cnt_reg[3]/NET0131  , \clgen_cnt_reg[4]/NET0131  , \clgen_cnt_reg[5]/NET0131  , \clgen_cnt_reg[6]/NET0131  , \clgen_cnt_reg[7]/NET0131  , \clgen_cnt_reg[8]/NET0131  , \clgen_cnt_reg[9]/NET0131  , \clgen_neg_edge_reg/NET0131  , \clgen_pos_edge_reg/NET0131  , \ctrl_reg[0]/NET0131  , \ctrl_reg[10]/NET0131  , \ctrl_reg[11]/NET0131  , \ctrl_reg[12]/NET0131  , \ctrl_reg[13]/NET0131  , \ctrl_reg[1]/NET0131  , \ctrl_reg[2]/NET0131  , \ctrl_reg[3]/NET0131  , \ctrl_reg[4]/NET0131  , \ctrl_reg[5]/NET0131  , \ctrl_reg[6]/NET0131  , \ctrl_reg[7]/NET0131  , \ctrl_reg[8]/NET0131  , \ctrl_reg[9]/NET0131  , \divider_reg[0]/NET0131  , \divider_reg[10]/NET0131  , \divider_reg[11]/NET0131  , \divider_reg[12]/NET0131  , \divider_reg[13]/NET0131  , \divider_reg[14]/NET0131  , \divider_reg[15]/NET0131  , \divider_reg[1]/NET0131  , \divider_reg[2]/NET0131  , \divider_reg[3]/NET0131  , \divider_reg[4]/NET0131  , \divider_reg[5]/NET0131  , \divider_reg[6]/NET0131  , \divider_reg[7]/NET0131  , \divider_reg[8]/NET0131  , \divider_reg[9]/NET0131  , miso_pad_i_pad , mosi_pad_o_pad , sclk_pad_o_pad , \shift_cnt_reg[0]/NET0131  , \shift_cnt_reg[1]/NET0131  , \shift_cnt_reg[2]/NET0131  , \shift_cnt_reg[3]/NET0131  , \shift_cnt_reg[4]/NET0131  , \shift_cnt_reg[5]/NET0131  , \shift_cnt_reg[6]/NET0131  , \shift_cnt_reg[7]/NET0131  , \shift_data_reg[0]/NET0131  , \shift_data_reg[100]/NET0131  , \shift_data_reg[101]/NET0131  , \shift_data_reg[102]/NET0131  , \shift_data_reg[103]/NET0131  , \shift_data_reg[104]/NET0131  , \shift_data_reg[105]/NET0131  , \shift_data_reg[106]/NET0131  , \shift_data_reg[107]/NET0131  , \shift_data_reg[108]/NET0131  , \shift_data_reg[109]/NET0131  , \shift_data_reg[10]/NET0131  , \shift_data_reg[110]/NET0131  , \shift_data_reg[111]/NET0131  , \shift_data_reg[112]/NET0131  , \shift_data_reg[113]/NET0131  , \shift_data_reg[114]/NET0131  , \shift_data_reg[115]/NET0131  , \shift_data_reg[116]/NET0131  , \shift_data_reg[117]/NET0131  , \shift_data_reg[118]/NET0131  , \shift_data_reg[119]/NET0131  , \shift_data_reg[11]/NET0131  , \shift_data_reg[120]/NET0131  , \shift_data_reg[121]/NET0131  , \shift_data_reg[122]/NET0131  , \shift_data_reg[123]/NET0131  , \shift_data_reg[124]/NET0131  , \shift_data_reg[125]/NET0131  , \shift_data_reg[126]/NET0131  , \shift_data_reg[127]/NET0131  , \shift_data_reg[12]/NET0131  , \shift_data_reg[13]/NET0131  , \shift_data_reg[14]/NET0131  , \shift_data_reg[15]/NET0131  , \shift_data_reg[16]/NET0131  , \shift_data_reg[17]/NET0131  , \shift_data_reg[18]/NET0131  , \shift_data_reg[19]/NET0131  , \shift_data_reg[1]/NET0131  , \shift_data_reg[20]/NET0131  , \shift_data_reg[21]/NET0131  , \shift_data_reg[22]/NET0131  , \shift_data_reg[23]/NET0131  , \shift_data_reg[24]/NET0131  , \shift_data_reg[25]/NET0131  , \shift_data_reg[26]/NET0131  , \shift_data_reg[27]/NET0131  , \shift_data_reg[28]/NET0131  , \shift_data_reg[29]/NET0131  , \shift_data_reg[2]/NET0131  , \shift_data_reg[30]/NET0131  , \shift_data_reg[31]/NET0131  , \shift_data_reg[32]/NET0131  , \shift_data_reg[33]/NET0131  , \shift_data_reg[34]/NET0131  , \shift_data_reg[35]/NET0131  , \shift_data_reg[36]/NET0131  , \shift_data_reg[37]/NET0131  , \shift_data_reg[38]/NET0131  , \shift_data_reg[39]/NET0131  , \shift_data_reg[3]/NET0131  , \shift_data_reg[40]/NET0131  , \shift_data_reg[41]/NET0131  , \shift_data_reg[42]/NET0131  , \shift_data_reg[43]/NET0131  , \shift_data_reg[44]/NET0131  , \shift_data_reg[45]/NET0131  , \shift_data_reg[46]/NET0131  , \shift_data_reg[47]/NET0131  , \shift_data_reg[48]/NET0131  , \shift_data_reg[49]/NET0131  , \shift_data_reg[4]/NET0131  , \shift_data_reg[50]/NET0131  , \shift_data_reg[51]/NET0131  , \shift_data_reg[52]/NET0131  , \shift_data_reg[53]/NET0131  , \shift_data_reg[54]/NET0131  , \shift_data_reg[55]/NET0131  , \shift_data_reg[56]/NET0131  , \shift_data_reg[57]/NET0131  , \shift_data_reg[58]/NET0131  , \shift_data_reg[59]/NET0131  , \shift_data_reg[5]/NET0131  , \shift_data_reg[60]/NET0131  , \shift_data_reg[61]/NET0131  , \shift_data_reg[62]/NET0131  , \shift_data_reg[63]/NET0131  , \shift_data_reg[64]/NET0131  , \shift_data_reg[65]/NET0131  , \shift_data_reg[66]/NET0131  , \shift_data_reg[67]/NET0131  , \shift_data_reg[68]/NET0131  , \shift_data_reg[69]/NET0131  , \shift_data_reg[6]/NET0131  , \shift_data_reg[70]/NET0131  , \shift_data_reg[71]/NET0131  , \shift_data_reg[72]/NET0131  , \shift_data_reg[73]/NET0131  , \shift_data_reg[74]/NET0131  , \shift_data_reg[75]/NET0131  , \shift_data_reg[76]/NET0131  , \shift_data_reg[77]/NET0131  , \shift_data_reg[78]/NET0131  , \shift_data_reg[79]/NET0131  , \shift_data_reg[7]/NET0131  , \shift_data_reg[80]/NET0131  , \shift_data_reg[81]/NET0131  , \shift_data_reg[82]/NET0131  , \shift_data_reg[83]/NET0131  , \shift_data_reg[84]/NET0131  , \shift_data_reg[85]/NET0131  , \shift_data_reg[86]/NET0131  , \shift_data_reg[87]/NET0131  , \shift_data_reg[88]/NET0131  , \shift_data_reg[89]/NET0131  , \shift_data_reg[8]/NET0131  , \shift_data_reg[90]/NET0131  , \shift_data_reg[91]/NET0131  , \shift_data_reg[92]/NET0131  , \shift_data_reg[93]/NET0131  , \shift_data_reg[94]/NET0131  , \shift_data_reg[95]/NET0131  , \shift_data_reg[96]/NET0131  , \shift_data_reg[97]/NET0131  , \shift_data_reg[98]/NET0131  , \shift_data_reg[99]/NET0131  , \shift_data_reg[9]/NET0131  , \shift_tip_reg/NET0131  , \ss_reg[0]/NET0131  , \ss_reg[1]/NET0131  , \ss_reg[2]/NET0131  , \ss_reg[3]/NET0131  , \ss_reg[4]/NET0131  , \ss_reg[5]/NET0131  , \ss_reg[6]/NET0131  , \ss_reg[7]/NET0131  , wb_ack_o_pad , \wb_adr_i[2]_pad  , \wb_adr_i[3]_pad  , \wb_adr_i[4]_pad  , wb_cyc_i_pad , \wb_dat_i[0]_pad  , \wb_dat_i[10]_pad  , \wb_dat_i[11]_pad  , \wb_dat_i[12]_pad  , \wb_dat_i[13]_pad  , \wb_dat_i[14]_pad  , \wb_dat_i[15]_pad  , \wb_dat_i[16]_pad  , \wb_dat_i[17]_pad  , \wb_dat_i[18]_pad  , \wb_dat_i[19]_pad  , \wb_dat_i[1]_pad  , \wb_dat_i[20]_pad  , \wb_dat_i[21]_pad  , \wb_dat_i[22]_pad  , \wb_dat_i[23]_pad  , \wb_dat_i[24]_pad  , \wb_dat_i[25]_pad  , \wb_dat_i[26]_pad  , \wb_dat_i[27]_pad  , \wb_dat_i[28]_pad  , \wb_dat_i[29]_pad  , \wb_dat_i[2]_pad  , \wb_dat_i[30]_pad  , \wb_dat_i[31]_pad  , \wb_dat_i[3]_pad  , \wb_dat_i[4]_pad  , \wb_dat_i[5]_pad  , \wb_dat_i[6]_pad  , \wb_dat_i[7]_pad  , \wb_dat_i[8]_pad  , \wb_dat_i[9]_pad  , wb_int_o_pad , \wb_sel_i[0]_pad  , \wb_sel_i[1]_pad  , \wb_sel_i[2]_pad  , \wb_sel_i[3]_pad  , wb_stb_i_pad , wb_we_i_pad , \_al_n1  , \g10384/_0_  , \g10421/_0_  , \g10487/_0_  , \g10622/_0_  , \g10625/_0_  , \g10631/_3_  , \g10641/_0_  , \g10677/_3_  , \g10695/_0_  , \g10699/_3_  , \g10796/_0_  , \g10814/_00_  , \g10815/_0_  , \g10819/_0_  , \g10821/_0_  , \g10824/_3_  , \g10858/_0_  , \g11042/_00_  , \g11067/_0_  , \g11071/_00_  , \g11074/_0_  , \g11075/_0_  , \g11076/_0_  , \g11077/_0_  , \g11078/_0_  , \g11079/_0_  , \g11080/_0_  , \g11149/_0_  , \g11151/_0_  , \g11190/_00_  , \g11297/_0_  , \g11298/_0_  , \g11300/_0_  , \g11301/_0_  , \g11303/_0_  , \g11346/_0_  , \g11347/_0_  , \g11348/_0_  , \g11358/_0_  , \g11359/_0_  , \g11360/_0_  , \g11361/_0_  , \g11362/_0_  , \g11363/_0_  , \g11470/_0_  , \g11499/_0_  , \g11501/_0_  , \g11502/_0_  , \g11503/_0_  , \g11504/_0_  , \g11505/_0_  , \g11506/_0_  , \g11507/_0_  , \g11508/_0_  , \g11509/_0_  , \g11510/_0_  , \g11511/_0_  , \g11512/_0_  , \g11513/_0_  , \g11514/_0_  , \g11515/_0_  , \g11516/_0_  , \g11517/_0_  , \g11519/_0_  , \g11520/_0_  , \g11521/_0_  , \g11522/_0_  , \g11523/_0_  , \g11524/_0_  , \g11525/_0_  , \g11526/_0_  , \g11527/_0_  , \g11528/_0_  , \g11529/_0_  , \g11530/_0_  , \g11531/_0_  , \g11532/_0_  , \g11533/_0_  , \g11534/_0_  , \g11535/_0_  , \g11536/_0_  , \g11537/_0_  , \g11538/_0_  , \g11539/_0_  , \g11655/_0_  , \g11658/_0_  , \g11659/_0_  , \g11661/_0_  , \g11662/_0_  , \g11680/_0_  , \g11723/_0_  , \g11726/_0_  , \g11730/_0_  , \g11739/_0_  , \g11750/_0_  , \g11759/_0_  , \g11760/_0_  , \g11761/_0_  , \g11764/_0_  , \g11765/_0_  , \g12212/_0_  , \g13497/_0_  , \g13884/_0_  , \g13982/_0_  , \g13999/_0_  , \g9305/_0_  , \g9306/_0_  , \g9307/_0_  , \g9308/_0_  , \g9309/_0_  , \g9310/_0_  , \g9346/_0_  , \g9347/_0_  , \g9348/_0_  , \g9349/_0_  , \g9350/_0_  , \g9351/_0_  , \g9352/_0_  , \g9353/_0_  , \g9354/_0_  , \g9355/_0_  , \g9356/_0_  , \g9357/_0_  , \g9358/_0_  , \g9359/_0_  , \g9360/_0_  , \g9361/_0_  , \g9362/_0_  , \g9363/_0_  , \g9364/_0_  , \g9365/_0_  , \g9366/_0_  , \g9367/_0_  , \g9368/_0_  , \g9369/_0_  , \g9370/_0_  , \g9371/_0_  , \g9372/_0_  , \g9373/_0_  , \g9374/_0_  , \g9375/_0_  , \g9380/_0_  , \g9381/_0_  , \g9382/_0_  , \g9383/_0_  , \g9384/_0_  , \g9385/_0_  , \g9386/_0_  , \g9387/_0_  , \g9388/_0_  , \g9389/_0_  , \g9390/_0_  , \g9391/_0_  , \g9392/_0_  , \g9393/_0_  , \g9394/_0_  , \g9395/_0_  , \g9396/_0_  , \g9397/_0_  , \g9398/_0_  , \g9399/_0_  , \g9400/_0_  , \g9401/_0_  , \g9402/_0_  , \g9403/_0_  , \g9404/_0_  , \g9405/_0_  , \g9406/_0_  , \g9407/_0_  , \g9408/_0_  , \g9409/_0_  , \g9410/_0_  , \g9411/_0_  , \g9439/_0_  , \g9440/_0_  , \g9441/_0_  , \g9442/_0_  , \g9443/_0_  , \g9444/_0_  , \g9445/_0_  , \g9446/_0_  , \g9447/_0_  , \g9448/_0_  , \g9449/_0_  , \g9450/_0_  , \g9451/_0_  , \g9452/_0_  , \g9453/_0_  , \g9454/_0_  , \g9455/_0_  , \g9456/_0_  , \g9457/_0_  , \g9458/_0_  , \g9459/_0_  , \g9461/_0_  , \g9462/_0_  , \g9463/_0_  , \g9464/_0_  , \g9465/_0_  , \g9466/_0_  , \g9529/_0_  , \g9530/_0_  , \g9531/_0_  , \g9532/_0_  , \g9535/_0_  , \g9542/_0_  , \g9543/_0_  , \g9546/_0_  , \g9547/_0_  , \g9548/_0_  , \g9549/_0_  , \g9550/_0_  , \g9551/_0_  , \g9552/_0_  , \g9553/_0_  , \g9559/_0_  , \g9568/_0_  , \g9571/_0_  , \g9573/_0_  , \g9583/_0_  , \g9589/_0_  , \g9590/_0_  , \g9591/_0_  , \g9592/_0_  , \g9593/_0_  , \g9594/_0_  , \g9595/_0_  , \g9596/_0_  , \g9597/_0_  , \ss_pad_o[0]_pad  , \ss_pad_o[1]_pad  , \ss_pad_o[2]_pad  , \ss_pad_o[3]_pad  , \ss_pad_o[4]_pad  , \ss_pad_o[5]_pad  , \ss_pad_o[6]_pad  , \ss_pad_o[7]_pad  , wb_err_o_pad );
  input \clgen_cnt_reg[0]/NET0131  ;
  input \clgen_cnt_reg[10]/NET0131  ;
  input \clgen_cnt_reg[11]/NET0131  ;
  input \clgen_cnt_reg[12]/NET0131  ;
  input \clgen_cnt_reg[13]/NET0131  ;
  input \clgen_cnt_reg[14]/NET0131  ;
  input \clgen_cnt_reg[15]/NET0131  ;
  input \clgen_cnt_reg[1]/NET0131  ;
  input \clgen_cnt_reg[2]/NET0131  ;
  input \clgen_cnt_reg[3]/NET0131  ;
  input \clgen_cnt_reg[4]/NET0131  ;
  input \clgen_cnt_reg[5]/NET0131  ;
  input \clgen_cnt_reg[6]/NET0131  ;
  input \clgen_cnt_reg[7]/NET0131  ;
  input \clgen_cnt_reg[8]/NET0131  ;
  input \clgen_cnt_reg[9]/NET0131  ;
  input \clgen_neg_edge_reg/NET0131  ;
  input \clgen_pos_edge_reg/NET0131  ;
  input \ctrl_reg[0]/NET0131  ;
  input \ctrl_reg[10]/NET0131  ;
  input \ctrl_reg[11]/NET0131  ;
  input \ctrl_reg[12]/NET0131  ;
  input \ctrl_reg[13]/NET0131  ;
  input \ctrl_reg[1]/NET0131  ;
  input \ctrl_reg[2]/NET0131  ;
  input \ctrl_reg[3]/NET0131  ;
  input \ctrl_reg[4]/NET0131  ;
  input \ctrl_reg[5]/NET0131  ;
  input \ctrl_reg[6]/NET0131  ;
  input \ctrl_reg[7]/NET0131  ;
  input \ctrl_reg[8]/NET0131  ;
  input \ctrl_reg[9]/NET0131  ;
  input \divider_reg[0]/NET0131  ;
  input \divider_reg[10]/NET0131  ;
  input \divider_reg[11]/NET0131  ;
  input \divider_reg[12]/NET0131  ;
  input \divider_reg[13]/NET0131  ;
  input \divider_reg[14]/NET0131  ;
  input \divider_reg[15]/NET0131  ;
  input \divider_reg[1]/NET0131  ;
  input \divider_reg[2]/NET0131  ;
  input \divider_reg[3]/NET0131  ;
  input \divider_reg[4]/NET0131  ;
  input \divider_reg[5]/NET0131  ;
  input \divider_reg[6]/NET0131  ;
  input \divider_reg[7]/NET0131  ;
  input \divider_reg[8]/NET0131  ;
  input \divider_reg[9]/NET0131  ;
  input miso_pad_i_pad ;
  input mosi_pad_o_pad ;
  input sclk_pad_o_pad ;
  input \shift_cnt_reg[0]/NET0131  ;
  input \shift_cnt_reg[1]/NET0131  ;
  input \shift_cnt_reg[2]/NET0131  ;
  input \shift_cnt_reg[3]/NET0131  ;
  input \shift_cnt_reg[4]/NET0131  ;
  input \shift_cnt_reg[5]/NET0131  ;
  input \shift_cnt_reg[6]/NET0131  ;
  input \shift_cnt_reg[7]/NET0131  ;
  input \shift_data_reg[0]/NET0131  ;
  input \shift_data_reg[100]/NET0131  ;
  input \shift_data_reg[101]/NET0131  ;
  input \shift_data_reg[102]/NET0131  ;
  input \shift_data_reg[103]/NET0131  ;
  input \shift_data_reg[104]/NET0131  ;
  input \shift_data_reg[105]/NET0131  ;
  input \shift_data_reg[106]/NET0131  ;
  input \shift_data_reg[107]/NET0131  ;
  input \shift_data_reg[108]/NET0131  ;
  input \shift_data_reg[109]/NET0131  ;
  input \shift_data_reg[10]/NET0131  ;
  input \shift_data_reg[110]/NET0131  ;
  input \shift_data_reg[111]/NET0131  ;
  input \shift_data_reg[112]/NET0131  ;
  input \shift_data_reg[113]/NET0131  ;
  input \shift_data_reg[114]/NET0131  ;
  input \shift_data_reg[115]/NET0131  ;
  input \shift_data_reg[116]/NET0131  ;
  input \shift_data_reg[117]/NET0131  ;
  input \shift_data_reg[118]/NET0131  ;
  input \shift_data_reg[119]/NET0131  ;
  input \shift_data_reg[11]/NET0131  ;
  input \shift_data_reg[120]/NET0131  ;
  input \shift_data_reg[121]/NET0131  ;
  input \shift_data_reg[122]/NET0131  ;
  input \shift_data_reg[123]/NET0131  ;
  input \shift_data_reg[124]/NET0131  ;
  input \shift_data_reg[125]/NET0131  ;
  input \shift_data_reg[126]/NET0131  ;
  input \shift_data_reg[127]/NET0131  ;
  input \shift_data_reg[12]/NET0131  ;
  input \shift_data_reg[13]/NET0131  ;
  input \shift_data_reg[14]/NET0131  ;
  input \shift_data_reg[15]/NET0131  ;
  input \shift_data_reg[16]/NET0131  ;
  input \shift_data_reg[17]/NET0131  ;
  input \shift_data_reg[18]/NET0131  ;
  input \shift_data_reg[19]/NET0131  ;
  input \shift_data_reg[1]/NET0131  ;
  input \shift_data_reg[20]/NET0131  ;
  input \shift_data_reg[21]/NET0131  ;
  input \shift_data_reg[22]/NET0131  ;
  input \shift_data_reg[23]/NET0131  ;
  input \shift_data_reg[24]/NET0131  ;
  input \shift_data_reg[25]/NET0131  ;
  input \shift_data_reg[26]/NET0131  ;
  input \shift_data_reg[27]/NET0131  ;
  input \shift_data_reg[28]/NET0131  ;
  input \shift_data_reg[29]/NET0131  ;
  input \shift_data_reg[2]/NET0131  ;
  input \shift_data_reg[30]/NET0131  ;
  input \shift_data_reg[31]/NET0131  ;
  input \shift_data_reg[32]/NET0131  ;
  input \shift_data_reg[33]/NET0131  ;
  input \shift_data_reg[34]/NET0131  ;
  input \shift_data_reg[35]/NET0131  ;
  input \shift_data_reg[36]/NET0131  ;
  input \shift_data_reg[37]/NET0131  ;
  input \shift_data_reg[38]/NET0131  ;
  input \shift_data_reg[39]/NET0131  ;
  input \shift_data_reg[3]/NET0131  ;
  input \shift_data_reg[40]/NET0131  ;
  input \shift_data_reg[41]/NET0131  ;
  input \shift_data_reg[42]/NET0131  ;
  input \shift_data_reg[43]/NET0131  ;
  input \shift_data_reg[44]/NET0131  ;
  input \shift_data_reg[45]/NET0131  ;
  input \shift_data_reg[46]/NET0131  ;
  input \shift_data_reg[47]/NET0131  ;
  input \shift_data_reg[48]/NET0131  ;
  input \shift_data_reg[49]/NET0131  ;
  input \shift_data_reg[4]/NET0131  ;
  input \shift_data_reg[50]/NET0131  ;
  input \shift_data_reg[51]/NET0131  ;
  input \shift_data_reg[52]/NET0131  ;
  input \shift_data_reg[53]/NET0131  ;
  input \shift_data_reg[54]/NET0131  ;
  input \shift_data_reg[55]/NET0131  ;
  input \shift_data_reg[56]/NET0131  ;
  input \shift_data_reg[57]/NET0131  ;
  input \shift_data_reg[58]/NET0131  ;
  input \shift_data_reg[59]/NET0131  ;
  input \shift_data_reg[5]/NET0131  ;
  input \shift_data_reg[60]/NET0131  ;
  input \shift_data_reg[61]/NET0131  ;
  input \shift_data_reg[62]/NET0131  ;
  input \shift_data_reg[63]/NET0131  ;
  input \shift_data_reg[64]/NET0131  ;
  input \shift_data_reg[65]/NET0131  ;
  input \shift_data_reg[66]/NET0131  ;
  input \shift_data_reg[67]/NET0131  ;
  input \shift_data_reg[68]/NET0131  ;
  input \shift_data_reg[69]/NET0131  ;
  input \shift_data_reg[6]/NET0131  ;
  input \shift_data_reg[70]/NET0131  ;
  input \shift_data_reg[71]/NET0131  ;
  input \shift_data_reg[72]/NET0131  ;
  input \shift_data_reg[73]/NET0131  ;
  input \shift_data_reg[74]/NET0131  ;
  input \shift_data_reg[75]/NET0131  ;
  input \shift_data_reg[76]/NET0131  ;
  input \shift_data_reg[77]/NET0131  ;
  input \shift_data_reg[78]/NET0131  ;
  input \shift_data_reg[79]/NET0131  ;
  input \shift_data_reg[7]/NET0131  ;
  input \shift_data_reg[80]/NET0131  ;
  input \shift_data_reg[81]/NET0131  ;
  input \shift_data_reg[82]/NET0131  ;
  input \shift_data_reg[83]/NET0131  ;
  input \shift_data_reg[84]/NET0131  ;
  input \shift_data_reg[85]/NET0131  ;
  input \shift_data_reg[86]/NET0131  ;
  input \shift_data_reg[87]/NET0131  ;
  input \shift_data_reg[88]/NET0131  ;
  input \shift_data_reg[89]/NET0131  ;
  input \shift_data_reg[8]/NET0131  ;
  input \shift_data_reg[90]/NET0131  ;
  input \shift_data_reg[91]/NET0131  ;
  input \shift_data_reg[92]/NET0131  ;
  input \shift_data_reg[93]/NET0131  ;
  input \shift_data_reg[94]/NET0131  ;
  input \shift_data_reg[95]/NET0131  ;
  input \shift_data_reg[96]/NET0131  ;
  input \shift_data_reg[97]/NET0131  ;
  input \shift_data_reg[98]/NET0131  ;
  input \shift_data_reg[99]/NET0131  ;
  input \shift_data_reg[9]/NET0131  ;
  input \shift_tip_reg/NET0131  ;
  input \ss_reg[0]/NET0131  ;
  input \ss_reg[1]/NET0131  ;
  input \ss_reg[2]/NET0131  ;
  input \ss_reg[3]/NET0131  ;
  input \ss_reg[4]/NET0131  ;
  input \ss_reg[5]/NET0131  ;
  input \ss_reg[6]/NET0131  ;
  input \ss_reg[7]/NET0131  ;
  input wb_ack_o_pad ;
  input \wb_adr_i[2]_pad  ;
  input \wb_adr_i[3]_pad  ;
  input \wb_adr_i[4]_pad  ;
  input wb_cyc_i_pad ;
  input \wb_dat_i[0]_pad  ;
  input \wb_dat_i[10]_pad  ;
  input \wb_dat_i[11]_pad  ;
  input \wb_dat_i[12]_pad  ;
  input \wb_dat_i[13]_pad  ;
  input \wb_dat_i[14]_pad  ;
  input \wb_dat_i[15]_pad  ;
  input \wb_dat_i[16]_pad  ;
  input \wb_dat_i[17]_pad  ;
  input \wb_dat_i[18]_pad  ;
  input \wb_dat_i[19]_pad  ;
  input \wb_dat_i[1]_pad  ;
  input \wb_dat_i[20]_pad  ;
  input \wb_dat_i[21]_pad  ;
  input \wb_dat_i[22]_pad  ;
  input \wb_dat_i[23]_pad  ;
  input \wb_dat_i[24]_pad  ;
  input \wb_dat_i[25]_pad  ;
  input \wb_dat_i[26]_pad  ;
  input \wb_dat_i[27]_pad  ;
  input \wb_dat_i[28]_pad  ;
  input \wb_dat_i[29]_pad  ;
  input \wb_dat_i[2]_pad  ;
  input \wb_dat_i[30]_pad  ;
  input \wb_dat_i[31]_pad  ;
  input \wb_dat_i[3]_pad  ;
  input \wb_dat_i[4]_pad  ;
  input \wb_dat_i[5]_pad  ;
  input \wb_dat_i[6]_pad  ;
  input \wb_dat_i[7]_pad  ;
  input \wb_dat_i[8]_pad  ;
  input \wb_dat_i[9]_pad  ;
  input wb_int_o_pad ;
  input \wb_sel_i[0]_pad  ;
  input \wb_sel_i[1]_pad  ;
  input \wb_sel_i[2]_pad  ;
  input \wb_sel_i[3]_pad  ;
  input wb_stb_i_pad ;
  input wb_we_i_pad ;
  output \_al_n1  ;
  output \g10384/_0_  ;
  output \g10421/_0_  ;
  output \g10487/_0_  ;
  output \g10622/_0_  ;
  output \g10625/_0_  ;
  output \g10631/_3_  ;
  output \g10641/_0_  ;
  output \g10677/_3_  ;
  output \g10695/_0_  ;
  output \g10699/_3_  ;
  output \g10796/_0_  ;
  output \g10814/_00_  ;
  output \g10815/_0_  ;
  output \g10819/_0_  ;
  output \g10821/_0_  ;
  output \g10824/_3_  ;
  output \g10858/_0_  ;
  output \g11042/_00_  ;
  output \g11067/_0_  ;
  output \g11071/_00_  ;
  output \g11074/_0_  ;
  output \g11075/_0_  ;
  output \g11076/_0_  ;
  output \g11077/_0_  ;
  output \g11078/_0_  ;
  output \g11079/_0_  ;
  output \g11080/_0_  ;
  output \g11149/_0_  ;
  output \g11151/_0_  ;
  output \g11190/_00_  ;
  output \g11297/_0_  ;
  output \g11298/_0_  ;
  output \g11300/_0_  ;
  output \g11301/_0_  ;
  output \g11303/_0_  ;
  output \g11346/_0_  ;
  output \g11347/_0_  ;
  output \g11348/_0_  ;
  output \g11358/_0_  ;
  output \g11359/_0_  ;
  output \g11360/_0_  ;
  output \g11361/_0_  ;
  output \g11362/_0_  ;
  output \g11363/_0_  ;
  output \g11470/_0_  ;
  output \g11499/_0_  ;
  output \g11501/_0_  ;
  output \g11502/_0_  ;
  output \g11503/_0_  ;
  output \g11504/_0_  ;
  output \g11505/_0_  ;
  output \g11506/_0_  ;
  output \g11507/_0_  ;
  output \g11508/_0_  ;
  output \g11509/_0_  ;
  output \g11510/_0_  ;
  output \g11511/_0_  ;
  output \g11512/_0_  ;
  output \g11513/_0_  ;
  output \g11514/_0_  ;
  output \g11515/_0_  ;
  output \g11516/_0_  ;
  output \g11517/_0_  ;
  output \g11519/_0_  ;
  output \g11520/_0_  ;
  output \g11521/_0_  ;
  output \g11522/_0_  ;
  output \g11523/_0_  ;
  output \g11524/_0_  ;
  output \g11525/_0_  ;
  output \g11526/_0_  ;
  output \g11527/_0_  ;
  output \g11528/_0_  ;
  output \g11529/_0_  ;
  output \g11530/_0_  ;
  output \g11531/_0_  ;
  output \g11532/_0_  ;
  output \g11533/_0_  ;
  output \g11534/_0_  ;
  output \g11535/_0_  ;
  output \g11536/_0_  ;
  output \g11537/_0_  ;
  output \g11538/_0_  ;
  output \g11539/_0_  ;
  output \g11655/_0_  ;
  output \g11658/_0_  ;
  output \g11659/_0_  ;
  output \g11661/_0_  ;
  output \g11662/_0_  ;
  output \g11680/_0_  ;
  output \g11723/_0_  ;
  output \g11726/_0_  ;
  output \g11730/_0_  ;
  output \g11739/_0_  ;
  output \g11750/_0_  ;
  output \g11759/_0_  ;
  output \g11760/_0_  ;
  output \g11761/_0_  ;
  output \g11764/_0_  ;
  output \g11765/_0_  ;
  output \g12212/_0_  ;
  output \g13497/_0_  ;
  output \g13884/_0_  ;
  output \g13982/_0_  ;
  output \g13999/_0_  ;
  output \g9305/_0_  ;
  output \g9306/_0_  ;
  output \g9307/_0_  ;
  output \g9308/_0_  ;
  output \g9309/_0_  ;
  output \g9310/_0_  ;
  output \g9346/_0_  ;
  output \g9347/_0_  ;
  output \g9348/_0_  ;
  output \g9349/_0_  ;
  output \g9350/_0_  ;
  output \g9351/_0_  ;
  output \g9352/_0_  ;
  output \g9353/_0_  ;
  output \g9354/_0_  ;
  output \g9355/_0_  ;
  output \g9356/_0_  ;
  output \g9357/_0_  ;
  output \g9358/_0_  ;
  output \g9359/_0_  ;
  output \g9360/_0_  ;
  output \g9361/_0_  ;
  output \g9362/_0_  ;
  output \g9363/_0_  ;
  output \g9364/_0_  ;
  output \g9365/_0_  ;
  output \g9366/_0_  ;
  output \g9367/_0_  ;
  output \g9368/_0_  ;
  output \g9369/_0_  ;
  output \g9370/_0_  ;
  output \g9371/_0_  ;
  output \g9372/_0_  ;
  output \g9373/_0_  ;
  output \g9374/_0_  ;
  output \g9375/_0_  ;
  output \g9380/_0_  ;
  output \g9381/_0_  ;
  output \g9382/_0_  ;
  output \g9383/_0_  ;
  output \g9384/_0_  ;
  output \g9385/_0_  ;
  output \g9386/_0_  ;
  output \g9387/_0_  ;
  output \g9388/_0_  ;
  output \g9389/_0_  ;
  output \g9390/_0_  ;
  output \g9391/_0_  ;
  output \g9392/_0_  ;
  output \g9393/_0_  ;
  output \g9394/_0_  ;
  output \g9395/_0_  ;
  output \g9396/_0_  ;
  output \g9397/_0_  ;
  output \g9398/_0_  ;
  output \g9399/_0_  ;
  output \g9400/_0_  ;
  output \g9401/_0_  ;
  output \g9402/_0_  ;
  output \g9403/_0_  ;
  output \g9404/_0_  ;
  output \g9405/_0_  ;
  output \g9406/_0_  ;
  output \g9407/_0_  ;
  output \g9408/_0_  ;
  output \g9409/_0_  ;
  output \g9410/_0_  ;
  output \g9411/_0_  ;
  output \g9439/_0_  ;
  output \g9440/_0_  ;
  output \g9441/_0_  ;
  output \g9442/_0_  ;
  output \g9443/_0_  ;
  output \g9444/_0_  ;
  output \g9445/_0_  ;
  output \g9446/_0_  ;
  output \g9447/_0_  ;
  output \g9448/_0_  ;
  output \g9449/_0_  ;
  output \g9450/_0_  ;
  output \g9451/_0_  ;
  output \g9452/_0_  ;
  output \g9453/_0_  ;
  output \g9454/_0_  ;
  output \g9455/_0_  ;
  output \g9456/_0_  ;
  output \g9457/_0_  ;
  output \g9458/_0_  ;
  output \g9459/_0_  ;
  output \g9461/_0_  ;
  output \g9462/_0_  ;
  output \g9463/_0_  ;
  output \g9464/_0_  ;
  output \g9465/_0_  ;
  output \g9466/_0_  ;
  output \g9529/_0_  ;
  output \g9530/_0_  ;
  output \g9531/_0_  ;
  output \g9532/_0_  ;
  output \g9535/_0_  ;
  output \g9542/_0_  ;
  output \g9543/_0_  ;
  output \g9546/_0_  ;
  output \g9547/_0_  ;
  output \g9548/_0_  ;
  output \g9549/_0_  ;
  output \g9550/_0_  ;
  output \g9551/_0_  ;
  output \g9552/_0_  ;
  output \g9553/_0_  ;
  output \g9559/_0_  ;
  output \g9568/_0_  ;
  output \g9571/_0_  ;
  output \g9573/_0_  ;
  output \g9583/_0_  ;
  output \g9589/_0_  ;
  output \g9590/_0_  ;
  output \g9591/_0_  ;
  output \g9592/_0_  ;
  output \g9593/_0_  ;
  output \g9594/_0_  ;
  output \g9595/_0_  ;
  output \g9596/_0_  ;
  output \g9597/_0_  ;
  output \ss_pad_o[0]_pad  ;
  output \ss_pad_o[1]_pad  ;
  output \ss_pad_o[2]_pad  ;
  output \ss_pad_o[3]_pad  ;
  output \ss_pad_o[4]_pad  ;
  output \ss_pad_o[5]_pad  ;
  output \ss_pad_o[6]_pad  ;
  output \ss_pad_o[7]_pad  ;
  output wb_err_o_pad ;
  wire n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 ;
  assign n330 = ~\ctrl_reg[4]/NET0131  & \shift_cnt_reg[4]/NET0131  ;
  assign n331 = \ctrl_reg[4]/NET0131  & ~\shift_cnt_reg[4]/NET0131  ;
  assign n332 = ~n330 & ~n331 ;
  assign n260 = \ctrl_reg[3]/NET0131  & ~\shift_cnt_reg[3]/NET0131  ;
  assign n259 = ~\ctrl_reg[3]/NET0131  & \shift_cnt_reg[3]/NET0131  ;
  assign n242 = \ctrl_reg[2]/NET0131  & ~\shift_cnt_reg[2]/NET0131  ;
  assign n241 = ~\ctrl_reg[2]/NET0131  & \shift_cnt_reg[2]/NET0131  ;
  assign n244 = \ctrl_reg[1]/NET0131  & ~\shift_cnt_reg[1]/NET0131  ;
  assign n245 = ~\ctrl_reg[1]/NET0131  & \shift_cnt_reg[1]/NET0131  ;
  assign n246 = ~\ctrl_reg[0]/NET0131  & \shift_cnt_reg[0]/NET0131  ;
  assign n247 = ~n245 & ~n246 ;
  assign n248 = ~n244 & ~n247 ;
  assign n262 = ~n241 & ~n248 ;
  assign n263 = ~n242 & ~n262 ;
  assign n333 = ~n259 & ~n263 ;
  assign n334 = ~n260 & ~n333 ;
  assign n335 = ~n332 & ~n334 ;
  assign n336 = n332 & n334 ;
  assign n337 = ~n335 & ~n336 ;
  assign n338 = \ctrl_reg[11]/NET0131  & ~n337 ;
  assign n253 = ~\shift_cnt_reg[0]/NET0131  & ~\shift_cnt_reg[1]/NET0131  ;
  assign n254 = ~\shift_cnt_reg[2]/NET0131  & n253 ;
  assign n268 = ~\shift_cnt_reg[3]/NET0131  & n254 ;
  assign n339 = ~\shift_cnt_reg[4]/NET0131  & n268 ;
  assign n340 = \shift_cnt_reg[4]/NET0131  & ~n268 ;
  assign n341 = ~n339 & ~n340 ;
  assign n342 = ~\ctrl_reg[11]/NET0131  & ~n341 ;
  assign n343 = ~n338 & ~n342 ;
  assign n243 = ~n241 & ~n242 ;
  assign n249 = ~n243 & ~n248 ;
  assign n250 = n243 & n248 ;
  assign n251 = ~n249 & ~n250 ;
  assign n252 = \ctrl_reg[11]/NET0131  & ~n251 ;
  assign n255 = \shift_cnt_reg[2]/NET0131  & ~n253 ;
  assign n256 = ~n254 & ~n255 ;
  assign n257 = ~\ctrl_reg[11]/NET0131  & ~n256 ;
  assign n258 = ~n252 & ~n257 ;
  assign n261 = ~n259 & ~n260 ;
  assign n264 = ~n261 & ~n263 ;
  assign n265 = n261 & n263 ;
  assign n266 = ~n264 & ~n265 ;
  assign n267 = \ctrl_reg[11]/NET0131  & ~n266 ;
  assign n269 = \shift_cnt_reg[3]/NET0131  & ~n254 ;
  assign n270 = ~n268 & ~n269 ;
  assign n271 = ~\ctrl_reg[11]/NET0131  & ~n270 ;
  assign n272 = ~n267 & ~n271 ;
  assign n273 = n258 & n272 ;
  assign n274 = ~n244 & ~n245 ;
  assign n275 = ~n246 & ~n274 ;
  assign n276 = n246 & n274 ;
  assign n277 = ~n275 & ~n276 ;
  assign n278 = \ctrl_reg[11]/NET0131  & ~n277 ;
  assign n279 = \shift_cnt_reg[0]/NET0131  & \shift_cnt_reg[1]/NET0131  ;
  assign n280 = ~n253 & ~n279 ;
  assign n281 = ~\ctrl_reg[11]/NET0131  & ~n280 ;
  assign n282 = ~n278 & ~n281 ;
  assign n283 = \ctrl_reg[11]/NET0131  & n246 ;
  assign n284 = ~\ctrl_reg[0]/NET0131  & \ctrl_reg[11]/NET0131  ;
  assign n285 = ~\shift_cnt_reg[0]/NET0131  & ~n284 ;
  assign n286 = ~n283 & ~n285 ;
  assign n361 = ~\shift_data_reg[51]/NET0131  & ~n286 ;
  assign n362 = ~\shift_data_reg[50]/NET0131  & n286 ;
  assign n363 = ~n361 & ~n362 ;
  assign n364 = ~n282 & n363 ;
  assign n365 = ~\shift_data_reg[49]/NET0131  & ~n286 ;
  assign n366 = ~\shift_data_reg[48]/NET0131  & n286 ;
  assign n367 = ~n365 & ~n366 ;
  assign n368 = n282 & n367 ;
  assign n369 = ~n364 & ~n368 ;
  assign n370 = n273 & ~n369 ;
  assign n403 = ~n343 & ~n370 ;
  assign n385 = ~\shift_data_reg[59]/NET0131  & ~n286 ;
  assign n386 = ~\shift_data_reg[58]/NET0131  & n286 ;
  assign n387 = ~n385 & ~n386 ;
  assign n388 = ~n282 & n387 ;
  assign n381 = ~\shift_data_reg[57]/NET0131  & ~n286 ;
  assign n382 = ~\shift_data_reg[56]/NET0131  & n286 ;
  assign n383 = ~n381 & ~n382 ;
  assign n384 = n282 & n383 ;
  assign n389 = n258 & ~n384 ;
  assign n390 = ~n388 & n389 ;
  assign n375 = ~\shift_data_reg[61]/NET0131  & ~n286 ;
  assign n376 = ~\shift_data_reg[60]/NET0131  & n286 ;
  assign n377 = ~n375 & ~n376 ;
  assign n378 = n282 & n377 ;
  assign n371 = ~\shift_data_reg[63]/NET0131  & ~n286 ;
  assign n372 = ~\shift_data_reg[62]/NET0131  & n286 ;
  assign n373 = ~n371 & ~n372 ;
  assign n374 = ~n282 & n373 ;
  assign n379 = ~n258 & ~n374 ;
  assign n380 = ~n378 & n379 ;
  assign n391 = ~n272 & ~n380 ;
  assign n392 = ~n390 & n391 ;
  assign n297 = ~n258 & n272 ;
  assign n393 = ~\shift_data_reg[55]/NET0131  & ~n286 ;
  assign n394 = ~\shift_data_reg[54]/NET0131  & n286 ;
  assign n395 = ~n393 & ~n394 ;
  assign n396 = ~n282 & n395 ;
  assign n397 = ~\shift_data_reg[53]/NET0131  & ~n286 ;
  assign n398 = ~\shift_data_reg[52]/NET0131  & n286 ;
  assign n399 = ~n397 & ~n398 ;
  assign n400 = n282 & n399 ;
  assign n401 = ~n396 & ~n400 ;
  assign n402 = n297 & ~n401 ;
  assign n404 = ~n392 & ~n402 ;
  assign n405 = n403 & n404 ;
  assign n287 = ~\shift_data_reg[35]/NET0131  & ~n286 ;
  assign n288 = ~\shift_data_reg[34]/NET0131  & n286 ;
  assign n289 = ~n287 & ~n288 ;
  assign n290 = ~n282 & n289 ;
  assign n291 = ~\shift_data_reg[33]/NET0131  & ~n286 ;
  assign n292 = ~\shift_data_reg[32]/NET0131  & n286 ;
  assign n293 = ~n291 & ~n292 ;
  assign n294 = n282 & n293 ;
  assign n295 = ~n290 & ~n294 ;
  assign n296 = n273 & ~n295 ;
  assign n298 = ~\shift_data_reg[39]/NET0131  & ~n286 ;
  assign n299 = ~\shift_data_reg[38]/NET0131  & n286 ;
  assign n300 = ~n298 & ~n299 ;
  assign n301 = ~n282 & n300 ;
  assign n302 = ~\shift_data_reg[37]/NET0131  & ~n286 ;
  assign n303 = ~\shift_data_reg[36]/NET0131  & n286 ;
  assign n304 = ~n302 & ~n303 ;
  assign n305 = n282 & n304 ;
  assign n306 = ~n301 & ~n305 ;
  assign n307 = n297 & ~n306 ;
  assign n344 = ~n296 & ~n307 ;
  assign n322 = ~\shift_data_reg[43]/NET0131  & ~n286 ;
  assign n323 = ~\shift_data_reg[42]/NET0131  & n286 ;
  assign n324 = ~n322 & ~n323 ;
  assign n325 = ~n282 & n324 ;
  assign n318 = ~\shift_data_reg[41]/NET0131  & ~n286 ;
  assign n319 = ~\shift_data_reg[40]/NET0131  & n286 ;
  assign n320 = ~n318 & ~n319 ;
  assign n321 = n282 & n320 ;
  assign n326 = n258 & ~n321 ;
  assign n327 = ~n325 & n326 ;
  assign n312 = ~\shift_data_reg[45]/NET0131  & ~n286 ;
  assign n313 = ~\shift_data_reg[44]/NET0131  & n286 ;
  assign n314 = ~n312 & ~n313 ;
  assign n315 = n282 & n314 ;
  assign n308 = ~\shift_data_reg[47]/NET0131  & ~n286 ;
  assign n309 = ~\shift_data_reg[46]/NET0131  & n286 ;
  assign n310 = ~n308 & ~n309 ;
  assign n311 = ~n282 & n310 ;
  assign n316 = ~n258 & ~n311 ;
  assign n317 = ~n315 & n316 ;
  assign n328 = ~n272 & ~n317 ;
  assign n329 = ~n327 & n328 ;
  assign n345 = ~n329 & n343 ;
  assign n346 = n344 & n345 ;
  assign n347 = ~\ctrl_reg[5]/NET0131  & \shift_cnt_reg[5]/NET0131  ;
  assign n348 = \ctrl_reg[5]/NET0131  & ~\shift_cnt_reg[5]/NET0131  ;
  assign n349 = ~n347 & ~n348 ;
  assign n350 = ~n330 & ~n334 ;
  assign n351 = ~n331 & ~n350 ;
  assign n352 = ~n349 & ~n351 ;
  assign n353 = n349 & n351 ;
  assign n354 = ~n352 & ~n353 ;
  assign n355 = \ctrl_reg[11]/NET0131  & ~n354 ;
  assign n356 = ~\shift_cnt_reg[5]/NET0131  & n339 ;
  assign n357 = \shift_cnt_reg[5]/NET0131  & ~n339 ;
  assign n358 = ~n356 & ~n357 ;
  assign n359 = ~\ctrl_reg[11]/NET0131  & ~n358 ;
  assign n360 = ~n355 & ~n359 ;
  assign n406 = ~n346 & ~n360 ;
  assign n407 = ~n405 & n406 ;
  assign n457 = ~\shift_data_reg[19]/NET0131  & ~n286 ;
  assign n458 = ~\shift_data_reg[18]/NET0131  & n286 ;
  assign n459 = ~n457 & ~n458 ;
  assign n460 = n273 & n459 ;
  assign n453 = ~\shift_data_reg[23]/NET0131  & ~n286 ;
  assign n454 = ~\shift_data_reg[22]/NET0131  & n286 ;
  assign n455 = ~n453 & ~n454 ;
  assign n456 = n297 & n455 ;
  assign n461 = ~n282 & ~n456 ;
  assign n462 = ~n460 & n461 ;
  assign n467 = ~\shift_data_reg[17]/NET0131  & ~n286 ;
  assign n468 = ~\shift_data_reg[16]/NET0131  & n286 ;
  assign n469 = ~n467 & ~n468 ;
  assign n470 = n273 & n469 ;
  assign n463 = ~\shift_data_reg[21]/NET0131  & ~n286 ;
  assign n464 = ~\shift_data_reg[20]/NET0131  & n286 ;
  assign n465 = ~n463 & ~n464 ;
  assign n466 = n297 & n465 ;
  assign n471 = n282 & ~n466 ;
  assign n472 = ~n470 & n471 ;
  assign n473 = ~n462 & ~n472 ;
  assign n488 = ~\shift_data_reg[27]/NET0131  & ~n286 ;
  assign n489 = ~\shift_data_reg[26]/NET0131  & n286 ;
  assign n490 = ~n488 & ~n489 ;
  assign n491 = ~n282 & n490 ;
  assign n484 = ~\shift_data_reg[25]/NET0131  & ~n286 ;
  assign n485 = ~\shift_data_reg[24]/NET0131  & n286 ;
  assign n486 = ~n484 & ~n485 ;
  assign n487 = n282 & n486 ;
  assign n492 = n258 & ~n487 ;
  assign n493 = ~n491 & n492 ;
  assign n478 = ~\shift_data_reg[29]/NET0131  & ~n286 ;
  assign n479 = ~\shift_data_reg[28]/NET0131  & n286 ;
  assign n480 = ~n478 & ~n479 ;
  assign n481 = n282 & n480 ;
  assign n474 = ~\shift_data_reg[31]/NET0131  & ~n286 ;
  assign n475 = ~\shift_data_reg[30]/NET0131  & n286 ;
  assign n476 = ~n474 & ~n475 ;
  assign n477 = ~n282 & n476 ;
  assign n482 = ~n258 & ~n477 ;
  assign n483 = ~n481 & n482 ;
  assign n494 = ~n272 & ~n483 ;
  assign n495 = ~n493 & n494 ;
  assign n496 = ~n343 & ~n495 ;
  assign n497 = ~n473 & n496 ;
  assign n408 = ~\shift_data_reg[3]/NET0131  & ~n286 ;
  assign n409 = ~\shift_data_reg[2]/NET0131  & n286 ;
  assign n410 = ~n408 & ~n409 ;
  assign n411 = ~n282 & n410 ;
  assign n412 = ~\shift_data_reg[1]/NET0131  & ~n286 ;
  assign n413 = ~\shift_data_reg[0]/NET0131  & n286 ;
  assign n414 = ~n412 & ~n413 ;
  assign n415 = n282 & n414 ;
  assign n416 = ~n411 & ~n415 ;
  assign n417 = n273 & ~n416 ;
  assign n450 = n343 & ~n417 ;
  assign n418 = ~\shift_data_reg[7]/NET0131  & ~n286 ;
  assign n419 = ~\shift_data_reg[6]/NET0131  & n286 ;
  assign n420 = ~n418 & ~n419 ;
  assign n421 = ~n282 & n420 ;
  assign n422 = ~\shift_data_reg[5]/NET0131  & ~n286 ;
  assign n423 = ~\shift_data_reg[4]/NET0131  & n286 ;
  assign n424 = ~n422 & ~n423 ;
  assign n425 = n282 & n424 ;
  assign n426 = ~n421 & ~n425 ;
  assign n427 = n297 & ~n426 ;
  assign n442 = ~\shift_data_reg[11]/NET0131  & ~n286 ;
  assign n443 = ~\shift_data_reg[10]/NET0131  & n286 ;
  assign n444 = ~n442 & ~n443 ;
  assign n445 = ~n282 & n444 ;
  assign n438 = ~\shift_data_reg[9]/NET0131  & ~n286 ;
  assign n439 = ~\shift_data_reg[8]/NET0131  & n286 ;
  assign n440 = ~n438 & ~n439 ;
  assign n441 = n282 & n440 ;
  assign n446 = n258 & ~n441 ;
  assign n447 = ~n445 & n446 ;
  assign n432 = ~\shift_data_reg[13]/NET0131  & ~n286 ;
  assign n433 = ~\shift_data_reg[12]/NET0131  & n286 ;
  assign n434 = ~n432 & ~n433 ;
  assign n435 = n282 & n434 ;
  assign n428 = ~\shift_data_reg[15]/NET0131  & ~n286 ;
  assign n429 = ~\shift_data_reg[14]/NET0131  & n286 ;
  assign n430 = ~n428 & ~n429 ;
  assign n431 = ~n282 & n430 ;
  assign n436 = ~n258 & ~n431 ;
  assign n437 = ~n435 & n436 ;
  assign n448 = ~n272 & ~n437 ;
  assign n449 = ~n447 & n448 ;
  assign n451 = ~n427 & ~n449 ;
  assign n452 = n450 & n451 ;
  assign n498 = n360 & ~n452 ;
  assign n499 = ~n497 & n498 ;
  assign n500 = ~n407 & ~n499 ;
  assign n501 = ~\shift_cnt_reg[6]/NET0131  & n356 ;
  assign n502 = \shift_cnt_reg[6]/NET0131  & ~n356 ;
  assign n503 = ~n501 & ~n502 ;
  assign n504 = ~\ctrl_reg[11]/NET0131  & ~n503 ;
  assign n505 = \ctrl_reg[6]/NET0131  & ~\shift_cnt_reg[6]/NET0131  ;
  assign n506 = ~\ctrl_reg[6]/NET0131  & \shift_cnt_reg[6]/NET0131  ;
  assign n507 = ~n505 & ~n506 ;
  assign n508 = ~n347 & ~n351 ;
  assign n509 = ~n348 & ~n508 ;
  assign n510 = n507 & n509 ;
  assign n511 = ~n507 & ~n509 ;
  assign n512 = ~n510 & ~n511 ;
  assign n513 = \ctrl_reg[11]/NET0131  & ~n512 ;
  assign n514 = ~n504 & ~n513 ;
  assign n515 = ~n500 & n514 ;
  assign n608 = ~\shift_data_reg[67]/NET0131  & ~n286 ;
  assign n609 = ~\shift_data_reg[66]/NET0131  & n286 ;
  assign n610 = ~n608 & ~n609 ;
  assign n611 = ~n282 & n610 ;
  assign n612 = ~\shift_data_reg[65]/NET0131  & ~n286 ;
  assign n613 = ~\shift_data_reg[64]/NET0131  & n286 ;
  assign n614 = ~n612 & ~n613 ;
  assign n615 = n282 & n614 ;
  assign n616 = ~n611 & ~n615 ;
  assign n617 = n273 & ~n616 ;
  assign n650 = n343 & ~n617 ;
  assign n618 = ~\shift_data_reg[71]/NET0131  & ~n286 ;
  assign n619 = ~\shift_data_reg[70]/NET0131  & n286 ;
  assign n620 = ~n618 & ~n619 ;
  assign n621 = ~n282 & n620 ;
  assign n622 = ~\shift_data_reg[69]/NET0131  & ~n286 ;
  assign n623 = ~\shift_data_reg[68]/NET0131  & n286 ;
  assign n624 = ~n622 & ~n623 ;
  assign n625 = n282 & n624 ;
  assign n626 = ~n621 & ~n625 ;
  assign n627 = n297 & ~n626 ;
  assign n642 = ~\shift_data_reg[73]/NET0131  & ~n286 ;
  assign n643 = ~\shift_data_reg[72]/NET0131  & n286 ;
  assign n644 = ~n642 & ~n643 ;
  assign n645 = n282 & n644 ;
  assign n638 = ~\shift_data_reg[75]/NET0131  & ~n286 ;
  assign n639 = ~\shift_data_reg[74]/NET0131  & n286 ;
  assign n640 = ~n638 & ~n639 ;
  assign n641 = ~n282 & n640 ;
  assign n646 = n258 & ~n641 ;
  assign n647 = ~n645 & n646 ;
  assign n632 = ~\shift_data_reg[79]/NET0131  & ~n286 ;
  assign n633 = ~\shift_data_reg[78]/NET0131  & n286 ;
  assign n634 = ~n632 & ~n633 ;
  assign n635 = ~n282 & n634 ;
  assign n628 = ~\shift_data_reg[77]/NET0131  & ~n286 ;
  assign n629 = ~\shift_data_reg[76]/NET0131  & n286 ;
  assign n630 = ~n628 & ~n629 ;
  assign n631 = n282 & n630 ;
  assign n636 = ~n258 & ~n631 ;
  assign n637 = ~n635 & n636 ;
  assign n648 = ~n272 & ~n637 ;
  assign n649 = ~n647 & n648 ;
  assign n651 = ~n627 & ~n649 ;
  assign n652 = n650 & n651 ;
  assign n653 = ~\shift_data_reg[83]/NET0131  & ~n286 ;
  assign n654 = ~\shift_data_reg[82]/NET0131  & n286 ;
  assign n655 = ~n653 & ~n654 ;
  assign n656 = ~n282 & n655 ;
  assign n657 = ~\shift_data_reg[81]/NET0131  & ~n286 ;
  assign n658 = ~\shift_data_reg[80]/NET0131  & n286 ;
  assign n659 = ~n657 & ~n658 ;
  assign n660 = n282 & n659 ;
  assign n661 = ~n656 & ~n660 ;
  assign n662 = n273 & ~n661 ;
  assign n695 = ~n343 & ~n662 ;
  assign n663 = ~\shift_data_reg[87]/NET0131  & ~n286 ;
  assign n664 = ~\shift_data_reg[86]/NET0131  & n286 ;
  assign n665 = ~n663 & ~n664 ;
  assign n666 = ~n282 & n665 ;
  assign n667 = ~\shift_data_reg[85]/NET0131  & ~n286 ;
  assign n668 = ~\shift_data_reg[84]/NET0131  & n286 ;
  assign n669 = ~n667 & ~n668 ;
  assign n670 = n282 & n669 ;
  assign n671 = ~n666 & ~n670 ;
  assign n672 = n297 & ~n671 ;
  assign n687 = ~\shift_data_reg[91]/NET0131  & ~n286 ;
  assign n688 = ~\shift_data_reg[90]/NET0131  & n286 ;
  assign n689 = ~n687 & ~n688 ;
  assign n690 = ~n282 & n689 ;
  assign n683 = ~\shift_data_reg[89]/NET0131  & ~n286 ;
  assign n684 = ~\shift_data_reg[88]/NET0131  & n286 ;
  assign n685 = ~n683 & ~n684 ;
  assign n686 = n282 & n685 ;
  assign n691 = n258 & ~n686 ;
  assign n692 = ~n690 & n691 ;
  assign n677 = ~\shift_data_reg[93]/NET0131  & ~n286 ;
  assign n678 = ~\shift_data_reg[92]/NET0131  & n286 ;
  assign n679 = ~n677 & ~n678 ;
  assign n680 = n282 & n679 ;
  assign n673 = ~\shift_data_reg[95]/NET0131  & ~n286 ;
  assign n674 = ~\shift_data_reg[94]/NET0131  & n286 ;
  assign n675 = ~n673 & ~n674 ;
  assign n676 = ~n282 & n675 ;
  assign n681 = ~n258 & ~n676 ;
  assign n682 = ~n680 & n681 ;
  assign n693 = ~n272 & ~n682 ;
  assign n694 = ~n692 & n693 ;
  assign n696 = ~n672 & ~n694 ;
  assign n697 = n695 & n696 ;
  assign n698 = ~n652 & ~n697 ;
  assign n699 = n360 & ~n698 ;
  assign n516 = ~\shift_data_reg[103]/NET0131  & ~n286 ;
  assign n517 = ~\shift_data_reg[102]/NET0131  & n286 ;
  assign n518 = ~n516 & ~n517 ;
  assign n519 = ~n282 & n518 ;
  assign n520 = ~\shift_data_reg[101]/NET0131  & ~n286 ;
  assign n521 = ~\shift_data_reg[100]/NET0131  & n286 ;
  assign n522 = ~n520 & ~n521 ;
  assign n523 = n282 & n522 ;
  assign n524 = ~n519 & ~n523 ;
  assign n525 = n297 & ~n524 ;
  assign n558 = n343 & ~n525 ;
  assign n526 = ~\shift_data_reg[99]/NET0131  & ~n286 ;
  assign n527 = ~\shift_data_reg[98]/NET0131  & n286 ;
  assign n528 = ~n526 & ~n527 ;
  assign n529 = ~n282 & n528 ;
  assign n530 = ~\shift_data_reg[97]/NET0131  & ~n286 ;
  assign n531 = ~\shift_data_reg[96]/NET0131  & n286 ;
  assign n532 = ~n530 & ~n531 ;
  assign n533 = n282 & n532 ;
  assign n534 = ~n529 & ~n533 ;
  assign n535 = n273 & ~n534 ;
  assign n550 = ~\shift_data_reg[107]/NET0131  & ~n286 ;
  assign n551 = ~\shift_data_reg[106]/NET0131  & n286 ;
  assign n552 = ~n550 & ~n551 ;
  assign n553 = ~n282 & n552 ;
  assign n546 = ~\shift_data_reg[105]/NET0131  & ~n286 ;
  assign n547 = ~\shift_data_reg[104]/NET0131  & n286 ;
  assign n548 = ~n546 & ~n547 ;
  assign n549 = n282 & n548 ;
  assign n554 = n258 & ~n549 ;
  assign n555 = ~n553 & n554 ;
  assign n540 = ~\shift_data_reg[109]/NET0131  & ~n286 ;
  assign n541 = ~\shift_data_reg[108]/NET0131  & n286 ;
  assign n542 = ~n540 & ~n541 ;
  assign n543 = n282 & n542 ;
  assign n536 = ~\shift_data_reg[111]/NET0131  & ~n286 ;
  assign n537 = ~\shift_data_reg[110]/NET0131  & n286 ;
  assign n538 = ~n536 & ~n537 ;
  assign n539 = ~n282 & n538 ;
  assign n544 = ~n258 & ~n539 ;
  assign n545 = ~n543 & n544 ;
  assign n556 = ~n272 & ~n545 ;
  assign n557 = ~n555 & n556 ;
  assign n559 = ~n535 & ~n557 ;
  assign n560 = n558 & n559 ;
  assign n561 = ~\shift_data_reg[119]/NET0131  & ~n286 ;
  assign n562 = ~\shift_data_reg[118]/NET0131  & n286 ;
  assign n563 = ~n561 & ~n562 ;
  assign n564 = ~n282 & n563 ;
  assign n565 = ~\shift_data_reg[117]/NET0131  & ~n286 ;
  assign n566 = ~\shift_data_reg[116]/NET0131  & n286 ;
  assign n567 = ~n565 & ~n566 ;
  assign n568 = n282 & n567 ;
  assign n569 = ~n564 & ~n568 ;
  assign n570 = n297 & ~n569 ;
  assign n603 = ~n343 & ~n570 ;
  assign n571 = ~\shift_data_reg[115]/NET0131  & ~n286 ;
  assign n572 = ~\shift_data_reg[114]/NET0131  & n286 ;
  assign n573 = ~n571 & ~n572 ;
  assign n574 = ~n282 & n573 ;
  assign n575 = ~\shift_data_reg[113]/NET0131  & ~n286 ;
  assign n576 = ~\shift_data_reg[112]/NET0131  & n286 ;
  assign n577 = ~n575 & ~n576 ;
  assign n578 = n282 & n577 ;
  assign n579 = ~n574 & ~n578 ;
  assign n580 = n273 & ~n579 ;
  assign n595 = ~\shift_data_reg[123]/NET0131  & ~n286 ;
  assign n596 = ~\shift_data_reg[122]/NET0131  & n286 ;
  assign n597 = ~n595 & ~n596 ;
  assign n598 = ~n282 & n597 ;
  assign n591 = ~\shift_data_reg[121]/NET0131  & ~n286 ;
  assign n592 = ~\shift_data_reg[120]/NET0131  & n286 ;
  assign n593 = ~n591 & ~n592 ;
  assign n594 = n282 & n593 ;
  assign n599 = n258 & ~n594 ;
  assign n600 = ~n598 & n599 ;
  assign n585 = ~\shift_data_reg[125]/NET0131  & ~n286 ;
  assign n586 = ~\shift_data_reg[124]/NET0131  & n286 ;
  assign n587 = ~n585 & ~n586 ;
  assign n588 = n282 & n587 ;
  assign n581 = ~\shift_data_reg[127]/NET0131  & ~n286 ;
  assign n582 = ~\shift_data_reg[126]/NET0131  & n286 ;
  assign n583 = ~n581 & ~n582 ;
  assign n584 = ~n282 & n583 ;
  assign n589 = ~n258 & ~n584 ;
  assign n590 = ~n588 & n589 ;
  assign n601 = ~n272 & ~n590 ;
  assign n602 = ~n600 & n601 ;
  assign n604 = ~n580 & ~n602 ;
  assign n605 = n603 & n604 ;
  assign n606 = ~n560 & ~n605 ;
  assign n607 = ~n360 & ~n606 ;
  assign n700 = ~n514 & ~n607 ;
  assign n701 = ~n699 & n700 ;
  assign n702 = ~n515 & ~n701 ;
  assign n704 = ~\shift_cnt_reg[7]/NET0131  & n501 ;
  assign n703 = ~\clgen_pos_edge_reg/NET0131  & ~\ctrl_reg[10]/NET0131  ;
  assign n705 = ~\clgen_neg_edge_reg/NET0131  & \ctrl_reg[10]/NET0131  ;
  assign n706 = ~n703 & ~n705 ;
  assign n707 = ~n704 & n706 ;
  assign n708 = \shift_tip_reg/NET0131  & ~n707 ;
  assign n709 = ~n702 & ~n708 ;
  assign n710 = mosi_pad_o_pad & n708 ;
  assign n711 = ~n709 & ~n710 ;
  assign n718 = ~\clgen_cnt_reg[7]/NET0131  & ~\clgen_cnt_reg[8]/NET0131  ;
  assign n719 = ~\clgen_cnt_reg[9]/NET0131  & n718 ;
  assign n720 = ~\clgen_cnt_reg[10]/NET0131  & ~\clgen_cnt_reg[11]/NET0131  ;
  assign n721 = ~\clgen_cnt_reg[4]/NET0131  & ~\clgen_cnt_reg[5]/NET0131  ;
  assign n722 = ~\clgen_cnt_reg[6]/NET0131  & n721 ;
  assign n723 = n720 & n722 ;
  assign n724 = n719 & n723 ;
  assign n712 = ~\clgen_cnt_reg[13]/NET0131  & ~\clgen_cnt_reg[14]/NET0131  ;
  assign n713 = ~\clgen_cnt_reg[12]/NET0131  & ~\clgen_cnt_reg[15]/NET0131  ;
  assign n714 = ~\clgen_cnt_reg[2]/NET0131  & ~\clgen_cnt_reg[3]/NET0131  ;
  assign n715 = n713 & n714 ;
  assign n716 = n712 & n715 ;
  assign n717 = ~\clgen_cnt_reg[0]/NET0131  & ~\clgen_cnt_reg[1]/NET0131  ;
  assign n725 = n716 & n717 ;
  assign n726 = n724 & n725 ;
  assign n727 = \shift_tip_reg/NET0131  & ~n726 ;
  assign n728 = ~\clgen_cnt_reg[2]/NET0131  & n717 ;
  assign n729 = ~\clgen_cnt_reg[3]/NET0131  & n728 ;
  assign n730 = ~\clgen_cnt_reg[4]/NET0131  & n729 ;
  assign n731 = ~\clgen_cnt_reg[5]/NET0131  & n730 ;
  assign n732 = ~\clgen_cnt_reg[6]/NET0131  & n731 ;
  assign n733 = n719 & n732 ;
  assign n734 = ~\clgen_cnt_reg[10]/NET0131  & n733 ;
  assign n735 = ~\clgen_cnt_reg[11]/NET0131  & n734 ;
  assign n736 = ~\clgen_cnt_reg[12]/NET0131  & n735 ;
  assign n737 = n712 & n736 ;
  assign n738 = \clgen_cnt_reg[15]/NET0131  & ~n737 ;
  assign n739 = ~\clgen_cnt_reg[15]/NET0131  & n737 ;
  assign n740 = ~n738 & ~n739 ;
  assign n741 = n727 & ~n740 ;
  assign n742 = \divider_reg[15]/NET0131  & ~n727 ;
  assign n743 = ~n741 & ~n742 ;
  assign n744 = \clgen_cnt_reg[11]/NET0131  & ~n734 ;
  assign n745 = ~n735 & ~n744 ;
  assign n746 = n727 & ~n745 ;
  assign n747 = \divider_reg[11]/NET0131  & ~n727 ;
  assign n748 = ~n746 & ~n747 ;
  assign n749 = \clgen_pos_edge_reg/NET0131  & ~n341 ;
  assign n750 = ~\clgen_pos_edge_reg/NET0131  & \shift_cnt_reg[4]/NET0131  ;
  assign n751 = ~n749 & ~n750 ;
  assign n752 = \shift_tip_reg/NET0131  & ~n751 ;
  assign n753 = \ctrl_reg[4]/NET0131  & ~\shift_tip_reg/NET0131  ;
  assign n754 = ~n752 & ~n753 ;
  assign n755 = ~\clgen_cnt_reg[7]/NET0131  & n732 ;
  assign n756 = \clgen_cnt_reg[7]/NET0131  & ~n732 ;
  assign n757 = ~n755 & ~n756 ;
  assign n758 = n727 & ~n757 ;
  assign n759 = \divider_reg[7]/NET0131  & ~n727 ;
  assign n760 = ~n758 & ~n759 ;
  assign n761 = \clgen_cnt_reg[12]/NET0131  & ~n735 ;
  assign n762 = ~n736 & ~n761 ;
  assign n763 = n727 & ~n762 ;
  assign n764 = \divider_reg[12]/NET0131  & ~n727 ;
  assign n765 = ~n763 & ~n764 ;
  assign n766 = \clgen_pos_edge_reg/NET0131  & n704 ;
  assign n767 = \shift_tip_reg/NET0131  & ~n766 ;
  assign n768 = \clgen_pos_edge_reg/NET0131  & n501 ;
  assign n769 = \shift_cnt_reg[7]/NET0131  & ~n768 ;
  assign n770 = n767 & ~n769 ;
  assign n773 = ~\ctrl_reg[4]/NET0131  & ~\ctrl_reg[5]/NET0131  ;
  assign n774 = ~\ctrl_reg[6]/NET0131  & n773 ;
  assign n771 = ~\ctrl_reg[0]/NET0131  & ~\ctrl_reg[1]/NET0131  ;
  assign n772 = ~\ctrl_reg[2]/NET0131  & ~\ctrl_reg[3]/NET0131  ;
  assign n775 = n771 & n772 ;
  assign n776 = n774 & n775 ;
  assign n777 = ~\shift_tip_reg/NET0131  & ~n776 ;
  assign n778 = ~n770 & ~n777 ;
  assign n779 = \clgen_cnt_reg[8]/NET0131  & ~n755 ;
  assign n780 = n718 & n732 ;
  assign n781 = ~n779 & ~n780 ;
  assign n782 = n727 & ~n781 ;
  assign n783 = \divider_reg[8]/NET0131  & ~n727 ;
  assign n784 = ~n782 & ~n783 ;
  assign n785 = \clgen_pos_edge_reg/NET0131  & ~n270 ;
  assign n786 = ~\clgen_pos_edge_reg/NET0131  & \shift_cnt_reg[3]/NET0131  ;
  assign n787 = ~n785 & ~n786 ;
  assign n788 = \shift_tip_reg/NET0131  & ~n787 ;
  assign n789 = \ctrl_reg[3]/NET0131  & ~\shift_tip_reg/NET0131  ;
  assign n790 = ~n788 & ~n789 ;
  assign n791 = \clgen_cnt_reg[4]/NET0131  & ~n729 ;
  assign n792 = ~n730 & ~n791 ;
  assign n793 = n727 & ~n792 ;
  assign n794 = \divider_reg[4]/NET0131  & ~n727 ;
  assign n795 = ~n793 & ~n794 ;
  assign n796 = ~\clgen_cnt_reg[13]/NET0131  & n736 ;
  assign n797 = \clgen_cnt_reg[14]/NET0131  & ~n796 ;
  assign n798 = ~n737 & ~n797 ;
  assign n799 = n727 & ~n798 ;
  assign n800 = \divider_reg[14]/NET0131  & ~n727 ;
  assign n801 = ~n799 & ~n800 ;
  assign n802 = \clgen_pos_edge_reg/NET0131  & ~n503 ;
  assign n803 = ~\clgen_pos_edge_reg/NET0131  & \shift_cnt_reg[6]/NET0131  ;
  assign n804 = ~n802 & ~n803 ;
  assign n805 = \shift_tip_reg/NET0131  & ~n804 ;
  assign n806 = \ctrl_reg[6]/NET0131  & ~\shift_tip_reg/NET0131  ;
  assign n807 = ~n805 & ~n806 ;
  assign n808 = \ctrl_reg[8]/NET0131  & ~\wb_sel_i[1]_pad  ;
  assign n809 = \wb_dat_i[8]_pad  & \wb_sel_i[1]_pad  ;
  assign n810 = ~n808 & ~n809 ;
  assign n811 = ~\wb_adr_i[2]_pad  & wb_stb_i_pad ;
  assign n812 = wb_we_i_pad & n811 ;
  assign n813 = ~\shift_tip_reg/NET0131  & \wb_adr_i[4]_pad  ;
  assign n814 = wb_cyc_i_pad & n813 ;
  assign n815 = ~\wb_adr_i[3]_pad  & n814 ;
  assign n816 = n812 & n815 ;
  assign n817 = ~n810 & n816 ;
  assign n818 = \shift_tip_reg/NET0131  & n766 ;
  assign n819 = \ctrl_reg[8]/NET0131  & ~n816 ;
  assign n820 = ~n818 & n819 ;
  assign n821 = ~n817 & ~n820 ;
  assign n822 = \clgen_cnt_reg[3]/NET0131  & ~n728 ;
  assign n823 = ~n729 & ~n822 ;
  assign n824 = n727 & ~n823 ;
  assign n825 = \divider_reg[3]/NET0131  & ~n727 ;
  assign n826 = ~n824 & ~n825 ;
  assign n827 = \clgen_cnt_reg[13]/NET0131  & ~n736 ;
  assign n828 = ~n796 & ~n827 ;
  assign n829 = n727 & ~n828 ;
  assign n830 = \divider_reg[13]/NET0131  & ~n727 ;
  assign n831 = ~n829 & ~n830 ;
  assign n832 = \clgen_cnt_reg[10]/NET0131  & ~n733 ;
  assign n833 = ~n734 & ~n832 ;
  assign n834 = n727 & ~n833 ;
  assign n835 = \divider_reg[10]/NET0131  & ~n727 ;
  assign n836 = ~n834 & ~n835 ;
  assign n837 = \shift_tip_reg/NET0131  & n726 ;
  assign n838 = sclk_pad_o_pad & ~n837 ;
  assign n839 = ~sclk_pad_o_pad & \shift_tip_reg/NET0131  ;
  assign n840 = n726 & n839 ;
  assign n841 = ~n704 & n840 ;
  assign n842 = ~n838 & ~n841 ;
  assign n843 = ~\clgen_pos_edge_reg/NET0131  & ~\shift_cnt_reg[2]/NET0131  ;
  assign n844 = \clgen_pos_edge_reg/NET0131  & n256 ;
  assign n845 = ~n843 & ~n844 ;
  assign n846 = \shift_tip_reg/NET0131  & ~n845 ;
  assign n847 = ~\ctrl_reg[2]/NET0131  & ~\shift_tip_reg/NET0131  ;
  assign n848 = ~n846 & ~n847 ;
  assign n865 = \clgen_cnt_reg[0]/NET0131  & ~\clgen_cnt_reg[1]/NET0131  ;
  assign n866 = n716 & n865 ;
  assign n867 = n724 & n866 ;
  assign n868 = sclk_pad_o_pad & ~n867 ;
  assign n851 = ~\divider_reg[13]/NET0131  & ~\divider_reg[14]/NET0131  ;
  assign n852 = ~\divider_reg[15]/NET0131  & ~\divider_reg[1]/NET0131  ;
  assign n859 = n851 & n852 ;
  assign n849 = ~\divider_reg[0]/NET0131  & ~\divider_reg[10]/NET0131  ;
  assign n850 = ~\divider_reg[11]/NET0131  & ~\divider_reg[12]/NET0131  ;
  assign n860 = n849 & n850 ;
  assign n861 = n859 & n860 ;
  assign n855 = ~\divider_reg[6]/NET0131  & ~\divider_reg[7]/NET0131  ;
  assign n856 = ~\divider_reg[8]/NET0131  & ~\divider_reg[9]/NET0131  ;
  assign n857 = n855 & n856 ;
  assign n853 = ~\divider_reg[2]/NET0131  & ~\divider_reg[3]/NET0131  ;
  assign n854 = ~\divider_reg[4]/NET0131  & ~\divider_reg[5]/NET0131  ;
  assign n858 = n853 & n854 ;
  assign n862 = n857 & n858 ;
  assign n863 = n861 & n862 ;
  assign n864 = ~sclk_pad_o_pad & ~n863 ;
  assign n869 = \shift_tip_reg/NET0131  & ~n864 ;
  assign n870 = ~n868 & n869 ;
  assign n871 = ~\clgen_pos_edge_reg/NET0131  & ~\shift_cnt_reg[5]/NET0131  ;
  assign n872 = \clgen_pos_edge_reg/NET0131  & n358 ;
  assign n873 = ~n871 & ~n872 ;
  assign n874 = \shift_tip_reg/NET0131  & ~n873 ;
  assign n875 = ~\ctrl_reg[5]/NET0131  & ~\shift_tip_reg/NET0131  ;
  assign n876 = ~n874 & ~n875 ;
  assign n877 = \ctrl_reg[8]/NET0131  & ~\shift_tip_reg/NET0131  ;
  assign n878 = ~n767 & ~n877 ;
  assign n879 = ~sclk_pad_o_pad & ~n877 ;
  assign n880 = n863 & ~n879 ;
  assign n881 = n839 & n867 ;
  assign n882 = ~n880 & ~n881 ;
  assign n883 = ~wb_ack_o_pad & wb_int_o_pad ;
  assign n884 = \ctrl_reg[12]/NET0131  & n818 ;
  assign n885 = ~n883 & ~n884 ;
  assign n886 = \divider_reg[5]/NET0131  & ~n727 ;
  assign n887 = \clgen_cnt_reg[5]/NET0131  & ~n730 ;
  assign n888 = ~n731 & ~n887 ;
  assign n889 = n727 & ~n888 ;
  assign n890 = ~n886 & ~n889 ;
  assign n891 = \divider_reg[6]/NET0131  & ~n727 ;
  assign n892 = \clgen_cnt_reg[6]/NET0131  & ~n731 ;
  assign n893 = ~n732 & ~n892 ;
  assign n894 = n727 & ~n893 ;
  assign n895 = ~n891 & ~n894 ;
  assign n896 = \divider_reg[0]/NET0131  & ~n727 ;
  assign n897 = ~\clgen_cnt_reg[0]/NET0131  & n727 ;
  assign n898 = ~n896 & ~n897 ;
  assign n899 = \clgen_cnt_reg[9]/NET0131  & ~n780 ;
  assign n900 = ~n733 & ~n899 ;
  assign n901 = n727 & ~n900 ;
  assign n902 = \divider_reg[9]/NET0131  & ~n727 ;
  assign n903 = ~n901 & ~n902 ;
  assign n904 = \clgen_cnt_reg[2]/NET0131  & ~n717 ;
  assign n905 = ~n728 & ~n904 ;
  assign n906 = n727 & ~n905 ;
  assign n907 = \divider_reg[2]/NET0131  & ~n727 ;
  assign n908 = ~n906 & ~n907 ;
  assign n909 = \divider_reg[1]/NET0131  & ~n727 ;
  assign n910 = ~\clgen_cnt_reg[0]/NET0131  & \clgen_cnt_reg[1]/NET0131  ;
  assign n911 = ~n865 & ~n910 ;
  assign n912 = n727 & n911 ;
  assign n913 = ~n909 & ~n912 ;
  assign n914 = ~\clgen_pos_edge_reg/NET0131  & ~\shift_cnt_reg[1]/NET0131  ;
  assign n915 = \clgen_pos_edge_reg/NET0131  & n280 ;
  assign n916 = ~n914 & ~n915 ;
  assign n917 = \shift_tip_reg/NET0131  & ~n916 ;
  assign n918 = ~\ctrl_reg[1]/NET0131  & ~\shift_tip_reg/NET0131  ;
  assign n919 = ~n917 & ~n918 ;
  assign n920 = \wb_adr_i[2]_pad  & ~\wb_adr_i[4]_pad  ;
  assign n936 = ~\wb_adr_i[3]_pad  & n920 ;
  assign n937 = \shift_data_reg[35]/NET0131  & n936 ;
  assign n931 = ~\wb_adr_i[2]_pad  & ~\wb_adr_i[4]_pad  ;
  assign n932 = \wb_adr_i[3]_pad  & n931 ;
  assign n933 = \shift_data_reg[67]/NET0131  & n932 ;
  assign n934 = ~\wb_adr_i[3]_pad  & n931 ;
  assign n935 = \shift_data_reg[3]/NET0131  & n934 ;
  assign n940 = ~n933 & ~n935 ;
  assign n941 = ~n937 & n940 ;
  assign n921 = \wb_adr_i[3]_pad  & n920 ;
  assign n922 = \shift_data_reg[99]/NET0131  & n921 ;
  assign n923 = ~\wb_adr_i[2]_pad  & \wb_adr_i[4]_pad  ;
  assign n924 = ~\wb_adr_i[3]_pad  & n923 ;
  assign n925 = \ctrl_reg[3]/NET0131  & n924 ;
  assign n938 = ~n922 & ~n925 ;
  assign n926 = \wb_adr_i[3]_pad  & n923 ;
  assign n927 = \ss_reg[3]/NET0131  & n926 ;
  assign n928 = \wb_adr_i[2]_pad  & ~\wb_adr_i[3]_pad  ;
  assign n929 = \wb_adr_i[4]_pad  & n928 ;
  assign n930 = \divider_reg[3]/NET0131  & n929 ;
  assign n939 = ~n927 & ~n930 ;
  assign n942 = n938 & n939 ;
  assign n943 = n941 & n942 ;
  assign n950 = \shift_data_reg[39]/NET0131  & n936 ;
  assign n948 = \shift_data_reg[71]/NET0131  & n932 ;
  assign n949 = \shift_data_reg[7]/NET0131  & n934 ;
  assign n953 = ~n948 & ~n949 ;
  assign n954 = ~n950 & n953 ;
  assign n944 = \shift_data_reg[103]/NET0131  & n921 ;
  assign n945 = \ctrl_reg[7]/NET0131  & n924 ;
  assign n951 = ~n944 & ~n945 ;
  assign n946 = \ss_reg[7]/NET0131  & n926 ;
  assign n947 = \divider_reg[7]/NET0131  & n929 ;
  assign n952 = ~n946 & ~n947 ;
  assign n955 = n951 & n952 ;
  assign n956 = n954 & n955 ;
  assign n957 = \shift_data_reg[40]/NET0131  & n936 ;
  assign n958 = \shift_data_reg[104]/NET0131  & n921 ;
  assign n963 = ~n957 & ~n958 ;
  assign n959 = \shift_data_reg[8]/NET0131  & n934 ;
  assign n960 = \divider_reg[8]/NET0131  & n929 ;
  assign n964 = ~n959 & ~n960 ;
  assign n961 = \shift_data_reg[72]/NET0131  & n932 ;
  assign n962 = \ctrl_reg[8]/NET0131  & n924 ;
  assign n965 = ~n961 & ~n962 ;
  assign n966 = n964 & n965 ;
  assign n967 = n963 & n966 ;
  assign n968 = \shift_data_reg[41]/NET0131  & n936 ;
  assign n969 = \shift_data_reg[105]/NET0131  & n921 ;
  assign n974 = ~n968 & ~n969 ;
  assign n970 = \shift_data_reg[9]/NET0131  & n934 ;
  assign n971 = \divider_reg[9]/NET0131  & n929 ;
  assign n975 = ~n970 & ~n971 ;
  assign n972 = \shift_data_reg[73]/NET0131  & n932 ;
  assign n973 = \ctrl_reg[9]/NET0131  & n924 ;
  assign n976 = ~n972 & ~n973 ;
  assign n977 = n975 & n976 ;
  assign n978 = n974 & n977 ;
  assign n979 = \shift_data_reg[42]/NET0131  & n936 ;
  assign n980 = \shift_data_reg[106]/NET0131  & n921 ;
  assign n985 = ~n979 & ~n980 ;
  assign n981 = \shift_data_reg[10]/NET0131  & n934 ;
  assign n982 = \divider_reg[10]/NET0131  & n929 ;
  assign n986 = ~n981 & ~n982 ;
  assign n983 = \shift_data_reg[74]/NET0131  & n932 ;
  assign n984 = \ctrl_reg[10]/NET0131  & n924 ;
  assign n987 = ~n983 & ~n984 ;
  assign n988 = n986 & n987 ;
  assign n989 = n985 & n988 ;
  assign n990 = \shift_data_reg[43]/NET0131  & n936 ;
  assign n991 = \shift_data_reg[107]/NET0131  & n921 ;
  assign n996 = ~n990 & ~n991 ;
  assign n992 = \shift_data_reg[11]/NET0131  & n934 ;
  assign n993 = \divider_reg[11]/NET0131  & n929 ;
  assign n997 = ~n992 & ~n993 ;
  assign n994 = \shift_data_reg[75]/NET0131  & n932 ;
  assign n995 = \ctrl_reg[11]/NET0131  & n924 ;
  assign n998 = ~n994 & ~n995 ;
  assign n999 = n997 & n998 ;
  assign n1000 = n996 & n999 ;
  assign n1001 = \shift_data_reg[44]/NET0131  & n936 ;
  assign n1002 = \shift_data_reg[108]/NET0131  & n921 ;
  assign n1007 = ~n1001 & ~n1002 ;
  assign n1003 = \shift_data_reg[12]/NET0131  & n934 ;
  assign n1004 = \divider_reg[12]/NET0131  & n929 ;
  assign n1008 = ~n1003 & ~n1004 ;
  assign n1005 = \shift_data_reg[76]/NET0131  & n932 ;
  assign n1006 = \ctrl_reg[12]/NET0131  & n924 ;
  assign n1009 = ~n1005 & ~n1006 ;
  assign n1010 = n1008 & n1009 ;
  assign n1011 = n1007 & n1010 ;
  assign n1012 = \shift_data_reg[45]/NET0131  & n936 ;
  assign n1013 = \shift_data_reg[109]/NET0131  & n921 ;
  assign n1018 = ~n1012 & ~n1013 ;
  assign n1014 = \shift_data_reg[13]/NET0131  & n934 ;
  assign n1015 = \divider_reg[13]/NET0131  & n929 ;
  assign n1019 = ~n1014 & ~n1015 ;
  assign n1016 = \shift_data_reg[77]/NET0131  & n932 ;
  assign n1017 = \ctrl_reg[13]/NET0131  & n924 ;
  assign n1020 = ~n1016 & ~n1017 ;
  assign n1021 = n1019 & n1020 ;
  assign n1022 = n1018 & n1021 ;
  assign n1029 = \ss_reg[2]/NET0131  & n926 ;
  assign n1027 = \divider_reg[2]/NET0131  & n929 ;
  assign n1028 = \shift_data_reg[98]/NET0131  & n921 ;
  assign n1032 = ~n1027 & ~n1028 ;
  assign n1033 = ~n1029 & n1032 ;
  assign n1023 = \ctrl_reg[2]/NET0131  & n924 ;
  assign n1024 = \shift_data_reg[2]/NET0131  & n934 ;
  assign n1030 = ~n1023 & ~n1024 ;
  assign n1025 = \shift_data_reg[34]/NET0131  & n936 ;
  assign n1026 = \shift_data_reg[66]/NET0131  & n932 ;
  assign n1031 = ~n1025 & ~n1026 ;
  assign n1034 = n1030 & n1031 ;
  assign n1035 = n1033 & n1034 ;
  assign n1042 = \ss_reg[5]/NET0131  & n926 ;
  assign n1040 = \divider_reg[5]/NET0131  & n929 ;
  assign n1041 = \shift_data_reg[101]/NET0131  & n921 ;
  assign n1045 = ~n1040 & ~n1041 ;
  assign n1046 = ~n1042 & n1045 ;
  assign n1036 = \ctrl_reg[5]/NET0131  & n924 ;
  assign n1037 = \shift_data_reg[5]/NET0131  & n934 ;
  assign n1043 = ~n1036 & ~n1037 ;
  assign n1038 = \shift_data_reg[37]/NET0131  & n936 ;
  assign n1039 = \shift_data_reg[69]/NET0131  & n932 ;
  assign n1044 = ~n1038 & ~n1039 ;
  assign n1047 = n1043 & n1044 ;
  assign n1048 = n1046 & n1047 ;
  assign n1055 = \ss_reg[6]/NET0131  & n926 ;
  assign n1053 = \divider_reg[6]/NET0131  & n929 ;
  assign n1054 = \shift_data_reg[102]/NET0131  & n921 ;
  assign n1058 = ~n1053 & ~n1054 ;
  assign n1059 = ~n1055 & n1058 ;
  assign n1049 = \ctrl_reg[6]/NET0131  & n924 ;
  assign n1050 = \shift_data_reg[6]/NET0131  & n934 ;
  assign n1056 = ~n1049 & ~n1050 ;
  assign n1051 = \shift_data_reg[38]/NET0131  & n936 ;
  assign n1052 = \shift_data_reg[70]/NET0131  & n932 ;
  assign n1057 = ~n1051 & ~n1052 ;
  assign n1060 = n1056 & n1057 ;
  assign n1061 = n1059 & n1060 ;
  assign n1068 = \ss_reg[4]/NET0131  & n926 ;
  assign n1066 = \divider_reg[4]/NET0131  & n929 ;
  assign n1067 = \shift_data_reg[100]/NET0131  & n921 ;
  assign n1071 = ~n1066 & ~n1067 ;
  assign n1072 = ~n1068 & n1071 ;
  assign n1062 = \ctrl_reg[4]/NET0131  & n924 ;
  assign n1063 = \shift_data_reg[4]/NET0131  & n934 ;
  assign n1069 = ~n1062 & ~n1063 ;
  assign n1064 = \shift_data_reg[36]/NET0131  & n936 ;
  assign n1065 = \shift_data_reg[68]/NET0131  & n932 ;
  assign n1070 = ~n1064 & ~n1065 ;
  assign n1073 = n1069 & n1070 ;
  assign n1074 = n1072 & n1073 ;
  assign n1081 = \ss_reg[0]/NET0131  & n926 ;
  assign n1079 = \divider_reg[0]/NET0131  & n929 ;
  assign n1080 = \shift_data_reg[96]/NET0131  & n921 ;
  assign n1084 = ~n1079 & ~n1080 ;
  assign n1085 = ~n1081 & n1084 ;
  assign n1075 = \ctrl_reg[0]/NET0131  & n924 ;
  assign n1076 = \shift_data_reg[0]/NET0131  & n934 ;
  assign n1082 = ~n1075 & ~n1076 ;
  assign n1077 = \shift_data_reg[32]/NET0131  & n936 ;
  assign n1078 = \shift_data_reg[64]/NET0131  & n932 ;
  assign n1083 = ~n1077 & ~n1078 ;
  assign n1086 = n1082 & n1083 ;
  assign n1087 = n1085 & n1086 ;
  assign n1094 = \ss_reg[1]/NET0131  & n926 ;
  assign n1092 = \divider_reg[1]/NET0131  & n929 ;
  assign n1093 = \shift_data_reg[97]/NET0131  & n921 ;
  assign n1097 = ~n1092 & ~n1093 ;
  assign n1098 = ~n1094 & n1097 ;
  assign n1088 = \ctrl_reg[1]/NET0131  & n924 ;
  assign n1089 = \shift_data_reg[1]/NET0131  & n934 ;
  assign n1095 = ~n1088 & ~n1089 ;
  assign n1090 = \shift_data_reg[33]/NET0131  & n936 ;
  assign n1091 = \shift_data_reg[65]/NET0131  & n932 ;
  assign n1096 = ~n1090 & ~n1091 ;
  assign n1099 = n1095 & n1096 ;
  assign n1100 = n1098 & n1099 ;
  assign n1101 = \shift_data_reg[78]/NET0131  & n932 ;
  assign n1102 = \shift_data_reg[110]/NET0131  & n921 ;
  assign n1106 = ~n1101 & ~n1102 ;
  assign n1105 = \shift_data_reg[46]/NET0131  & n936 ;
  assign n1103 = \shift_data_reg[14]/NET0131  & n934 ;
  assign n1104 = \divider_reg[14]/NET0131  & n929 ;
  assign n1107 = ~n1103 & ~n1104 ;
  assign n1108 = ~n1105 & n1107 ;
  assign n1109 = n1106 & n1108 ;
  assign n1110 = \shift_data_reg[79]/NET0131  & n932 ;
  assign n1111 = \shift_data_reg[111]/NET0131  & n921 ;
  assign n1115 = ~n1110 & ~n1111 ;
  assign n1114 = \shift_data_reg[47]/NET0131  & n936 ;
  assign n1112 = \shift_data_reg[15]/NET0131  & n934 ;
  assign n1113 = \divider_reg[15]/NET0131  & n929 ;
  assign n1116 = ~n1112 & ~n1113 ;
  assign n1117 = ~n1114 & n1116 ;
  assign n1118 = n1115 & n1117 ;
  assign n1119 = \ctrl_reg[0]/NET0131  & ~\shift_tip_reg/NET0131  ;
  assign n1121 = \clgen_pos_edge_reg/NET0131  & \shift_cnt_reg[0]/NET0131  ;
  assign n1120 = ~\clgen_pos_edge_reg/NET0131  & ~\shift_cnt_reg[0]/NET0131  ;
  assign n1122 = \shift_tip_reg/NET0131  & ~n1120 ;
  assign n1123 = ~n1121 & n1122 ;
  assign n1124 = ~n1119 & ~n1123 ;
  assign n1125 = \wb_sel_i[0]_pad  & n816 ;
  assign n1126 = \wb_dat_i[0]_pad  & n1125 ;
  assign n1127 = ~\ctrl_reg[0]/NET0131  & ~n1126 ;
  assign n1128 = \wb_adr_i[2]_pad  & wb_stb_i_pad ;
  assign n1129 = wb_we_i_pad & n1128 ;
  assign n1130 = n815 & n1129 ;
  assign n1131 = \wb_sel_i[0]_pad  & n1130 ;
  assign n1132 = \divider_reg[4]/NET0131  & ~n1131 ;
  assign n1133 = \wb_dat_i[4]_pad  & \wb_sel_i[0]_pad  ;
  assign n1134 = n1130 & n1133 ;
  assign n1135 = ~n1132 & ~n1134 ;
  assign n1136 = \wb_adr_i[3]_pad  & n812 ;
  assign n1137 = n814 & n1136 ;
  assign n1138 = \wb_sel_i[0]_pad  & n1137 ;
  assign n1139 = \ss_reg[4]/NET0131  & ~n1138 ;
  assign n1140 = n1133 & n1137 ;
  assign n1141 = ~n1139 & ~n1140 ;
  assign n1142 = \wb_sel_i[1]_pad  & n1130 ;
  assign n1143 = \divider_reg[10]/NET0131  & ~n1142 ;
  assign n1144 = \wb_dat_i[10]_pad  & \wb_sel_i[1]_pad  ;
  assign n1145 = n1130 & n1144 ;
  assign n1146 = ~n1143 & ~n1145 ;
  assign n1147 = \ctrl_reg[7]/NET0131  & ~n1125 ;
  assign n1148 = \wb_dat_i[7]_pad  & \wb_sel_i[0]_pad  ;
  assign n1149 = n816 & n1148 ;
  assign n1150 = ~n1147 & ~n1149 ;
  assign n1151 = \divider_reg[13]/NET0131  & ~n1142 ;
  assign n1152 = \wb_dat_i[13]_pad  & \wb_sel_i[1]_pad  ;
  assign n1153 = n1130 & n1152 ;
  assign n1154 = ~n1151 & ~n1153 ;
  assign n1155 = \divider_reg[5]/NET0131  & ~n1131 ;
  assign n1156 = \wb_dat_i[5]_pad  & \wb_sel_i[0]_pad  ;
  assign n1157 = n1130 & n1156 ;
  assign n1158 = ~n1155 & ~n1157 ;
  assign n1159 = \ss_reg[7]/NET0131  & ~n1138 ;
  assign n1160 = n1137 & n1148 ;
  assign n1161 = ~n1159 & ~n1160 ;
  assign n1162 = \divider_reg[2]/NET0131  & ~n1131 ;
  assign n1163 = \wb_dat_i[2]_pad  & \wb_sel_i[0]_pad  ;
  assign n1164 = n1130 & n1163 ;
  assign n1165 = ~n1162 & ~n1164 ;
  assign n1166 = \wb_sel_i[1]_pad  & n816 ;
  assign n1167 = \ctrl_reg[10]/NET0131  & ~n1166 ;
  assign n1168 = n816 & n1144 ;
  assign n1169 = ~n1167 & ~n1168 ;
  assign n1170 = \ctrl_reg[11]/NET0131  & ~n1166 ;
  assign n1171 = \wb_dat_i[11]_pad  & \wb_sel_i[1]_pad  ;
  assign n1172 = n816 & n1171 ;
  assign n1173 = ~n1170 & ~n1172 ;
  assign n1174 = \divider_reg[14]/NET0131  & ~n1142 ;
  assign n1175 = \wb_dat_i[14]_pad  & \wb_sel_i[1]_pad  ;
  assign n1176 = n1130 & n1175 ;
  assign n1177 = ~n1174 & ~n1176 ;
  assign n1178 = \ss_reg[6]/NET0131  & ~n1138 ;
  assign n1179 = \wb_dat_i[6]_pad  & \wb_sel_i[0]_pad  ;
  assign n1180 = n1137 & n1179 ;
  assign n1181 = ~n1178 & ~n1180 ;
  assign n1182 = \ctrl_reg[13]/NET0131  & ~n1166 ;
  assign n1183 = n816 & n1152 ;
  assign n1184 = ~n1182 & ~n1183 ;
  assign n1185 = \ss_reg[5]/NET0131  & ~n1138 ;
  assign n1186 = n1137 & n1156 ;
  assign n1187 = ~n1185 & ~n1186 ;
  assign n1188 = \ctrl_reg[1]/NET0131  & ~n1125 ;
  assign n1189 = \wb_dat_i[1]_pad  & \wb_sel_i[0]_pad  ;
  assign n1190 = n816 & n1189 ;
  assign n1191 = ~n1188 & ~n1190 ;
  assign n1192 = \ctrl_reg[2]/NET0131  & ~n1125 ;
  assign n1193 = n816 & n1163 ;
  assign n1194 = ~n1192 & ~n1193 ;
  assign n1195 = \ss_reg[2]/NET0131  & ~n1138 ;
  assign n1196 = n1137 & n1163 ;
  assign n1197 = ~n1195 & ~n1196 ;
  assign n1198 = \ctrl_reg[3]/NET0131  & ~n1125 ;
  assign n1199 = \wb_dat_i[3]_pad  & \wb_sel_i[0]_pad  ;
  assign n1200 = n816 & n1199 ;
  assign n1201 = ~n1198 & ~n1200 ;
  assign n1202 = \ctrl_reg[4]/NET0131  & ~n1125 ;
  assign n1203 = n816 & n1133 ;
  assign n1204 = ~n1202 & ~n1203 ;
  assign n1205 = \ctrl_reg[5]/NET0131  & ~n1125 ;
  assign n1206 = n816 & n1156 ;
  assign n1207 = ~n1205 & ~n1206 ;
  assign n1208 = \ctrl_reg[12]/NET0131  & ~n1166 ;
  assign n1209 = \wb_dat_i[12]_pad  & \wb_sel_i[1]_pad  ;
  assign n1210 = n816 & n1209 ;
  assign n1211 = ~n1208 & ~n1210 ;
  assign n1212 = \ctrl_reg[6]/NET0131  & ~n1125 ;
  assign n1213 = n816 & n1179 ;
  assign n1214 = ~n1212 & ~n1213 ;
  assign n1215 = \ctrl_reg[9]/NET0131  & ~n1166 ;
  assign n1216 = \wb_dat_i[9]_pad  & \wb_sel_i[1]_pad  ;
  assign n1217 = n816 & n1216 ;
  assign n1218 = ~n1215 & ~n1217 ;
  assign n1219 = \divider_reg[0]/NET0131  & ~n1131 ;
  assign n1220 = \wb_dat_i[0]_pad  & \wb_sel_i[0]_pad  ;
  assign n1221 = n1130 & n1220 ;
  assign n1222 = ~n1219 & ~n1221 ;
  assign n1223 = \divider_reg[11]/NET0131  & ~n1142 ;
  assign n1224 = n1130 & n1171 ;
  assign n1225 = ~n1223 & ~n1224 ;
  assign n1226 = \divider_reg[12]/NET0131  & ~n1142 ;
  assign n1227 = n1130 & n1209 ;
  assign n1228 = ~n1226 & ~n1227 ;
  assign n1229 = \divider_reg[15]/NET0131  & ~n1142 ;
  assign n1230 = \wb_dat_i[15]_pad  & \wb_sel_i[1]_pad  ;
  assign n1231 = n1130 & n1230 ;
  assign n1232 = ~n1229 & ~n1231 ;
  assign n1233 = \divider_reg[8]/NET0131  & ~n1142 ;
  assign n1234 = n809 & n1130 ;
  assign n1235 = ~n1233 & ~n1234 ;
  assign n1236 = \divider_reg[1]/NET0131  & ~n1131 ;
  assign n1237 = n1130 & n1189 ;
  assign n1238 = ~n1236 & ~n1237 ;
  assign n1239 = \divider_reg[6]/NET0131  & ~n1131 ;
  assign n1240 = n1130 & n1179 ;
  assign n1241 = ~n1239 & ~n1240 ;
  assign n1242 = \divider_reg[3]/NET0131  & ~n1131 ;
  assign n1243 = n1130 & n1199 ;
  assign n1244 = ~n1242 & ~n1243 ;
  assign n1245 = \ss_reg[0]/NET0131  & ~n1138 ;
  assign n1246 = n1137 & n1220 ;
  assign n1247 = ~n1245 & ~n1246 ;
  assign n1248 = \ss_reg[1]/NET0131  & ~n1138 ;
  assign n1249 = n1137 & n1189 ;
  assign n1250 = ~n1248 & ~n1249 ;
  assign n1251 = \ss_reg[3]/NET0131  & ~n1138 ;
  assign n1252 = n1137 & n1199 ;
  assign n1253 = ~n1251 & ~n1252 ;
  assign n1254 = \divider_reg[7]/NET0131  & ~n1131 ;
  assign n1255 = n1130 & n1148 ;
  assign n1256 = ~n1254 & ~n1255 ;
  assign n1257 = \divider_reg[9]/NET0131  & ~n1142 ;
  assign n1258 = n1130 & n1216 ;
  assign n1259 = ~n1257 & ~n1258 ;
  assign n1260 = \shift_data_reg[120]/NET0131  & n921 ;
  assign n1261 = \shift_data_reg[56]/NET0131  & n936 ;
  assign n1264 = ~n1260 & ~n1261 ;
  assign n1262 = \shift_data_reg[88]/NET0131  & n932 ;
  assign n1263 = \shift_data_reg[24]/NET0131  & n934 ;
  assign n1265 = ~n1262 & ~n1263 ;
  assign n1266 = n1264 & n1265 ;
  assign n1267 = \shift_data_reg[122]/NET0131  & n921 ;
  assign n1268 = \shift_data_reg[90]/NET0131  & n932 ;
  assign n1271 = ~n1267 & ~n1268 ;
  assign n1269 = \shift_data_reg[26]/NET0131  & n934 ;
  assign n1270 = \shift_data_reg[58]/NET0131  & n936 ;
  assign n1272 = ~n1269 & ~n1270 ;
  assign n1273 = n1271 & n1272 ;
  assign n1274 = \shift_data_reg[125]/NET0131  & n921 ;
  assign n1275 = \shift_data_reg[61]/NET0131  & n936 ;
  assign n1278 = ~n1274 & ~n1275 ;
  assign n1276 = \shift_data_reg[93]/NET0131  & n932 ;
  assign n1277 = \shift_data_reg[29]/NET0131  & n934 ;
  assign n1279 = ~n1276 & ~n1277 ;
  assign n1280 = n1278 & n1279 ;
  assign n1281 = \shift_data_reg[126]/NET0131  & n921 ;
  assign n1282 = \shift_data_reg[62]/NET0131  & n936 ;
  assign n1285 = ~n1281 & ~n1282 ;
  assign n1283 = \shift_data_reg[94]/NET0131  & n932 ;
  assign n1284 = \shift_data_reg[30]/NET0131  & n934 ;
  assign n1286 = ~n1283 & ~n1284 ;
  assign n1287 = n1285 & n1286 ;
  assign n1288 = \shift_data_reg[127]/NET0131  & n921 ;
  assign n1289 = \shift_data_reg[63]/NET0131  & n936 ;
  assign n1292 = ~n1288 & ~n1289 ;
  assign n1290 = \shift_data_reg[95]/NET0131  & n932 ;
  assign n1291 = \shift_data_reg[31]/NET0131  & n934 ;
  assign n1293 = ~n1290 & ~n1291 ;
  assign n1294 = n1292 & n1293 ;
  assign n1295 = \shift_data_reg[121]/NET0131  & n921 ;
  assign n1296 = \shift_data_reg[57]/NET0131  & n936 ;
  assign n1299 = ~n1295 & ~n1296 ;
  assign n1297 = \shift_data_reg[89]/NET0131  & n932 ;
  assign n1298 = \shift_data_reg[25]/NET0131  & n934 ;
  assign n1300 = ~n1297 & ~n1298 ;
  assign n1301 = n1299 & n1300 ;
  assign n1302 = \shift_data_reg[123]/NET0131  & n921 ;
  assign n1303 = \shift_data_reg[59]/NET0131  & n936 ;
  assign n1306 = ~n1302 & ~n1303 ;
  assign n1304 = \shift_data_reg[91]/NET0131  & n932 ;
  assign n1305 = \shift_data_reg[27]/NET0131  & n934 ;
  assign n1307 = ~n1304 & ~n1305 ;
  assign n1308 = n1306 & n1307 ;
  assign n1309 = \shift_data_reg[124]/NET0131  & n921 ;
  assign n1310 = \shift_data_reg[60]/NET0131  & n936 ;
  assign n1313 = ~n1309 & ~n1310 ;
  assign n1311 = \shift_data_reg[92]/NET0131  & n932 ;
  assign n1312 = \shift_data_reg[28]/NET0131  & n934 ;
  assign n1314 = ~n1311 & ~n1312 ;
  assign n1315 = n1313 & n1314 ;
  assign n1316 = \shift_data_reg[114]/NET0131  & n921 ;
  assign n1317 = \shift_data_reg[50]/NET0131  & n936 ;
  assign n1320 = ~n1316 & ~n1317 ;
  assign n1318 = \shift_data_reg[82]/NET0131  & n932 ;
  assign n1319 = \shift_data_reg[18]/NET0131  & n934 ;
  assign n1321 = ~n1318 & ~n1319 ;
  assign n1322 = n1320 & n1321 ;
  assign n1323 = \shift_data_reg[116]/NET0131  & n921 ;
  assign n1324 = \shift_data_reg[52]/NET0131  & n936 ;
  assign n1327 = ~n1323 & ~n1324 ;
  assign n1325 = \shift_data_reg[84]/NET0131  & n932 ;
  assign n1326 = \shift_data_reg[20]/NET0131  & n934 ;
  assign n1328 = ~n1325 & ~n1326 ;
  assign n1329 = n1327 & n1328 ;
  assign n1330 = \shift_data_reg[119]/NET0131  & n921 ;
  assign n1331 = \shift_data_reg[55]/NET0131  & n936 ;
  assign n1334 = ~n1330 & ~n1331 ;
  assign n1332 = \shift_data_reg[87]/NET0131  & n932 ;
  assign n1333 = \shift_data_reg[23]/NET0131  & n934 ;
  assign n1335 = ~n1332 & ~n1333 ;
  assign n1336 = n1334 & n1335 ;
  assign n1337 = \shift_data_reg[16]/NET0131  & n934 ;
  assign n1338 = \shift_data_reg[80]/NET0131  & n932 ;
  assign n1341 = ~n1337 & ~n1338 ;
  assign n1339 = \shift_data_reg[48]/NET0131  & n936 ;
  assign n1340 = \shift_data_reg[112]/NET0131  & n921 ;
  assign n1342 = ~n1339 & ~n1340 ;
  assign n1343 = n1341 & n1342 ;
  assign n1344 = \shift_data_reg[17]/NET0131  & n934 ;
  assign n1345 = \shift_data_reg[81]/NET0131  & n932 ;
  assign n1348 = ~n1344 & ~n1345 ;
  assign n1346 = \shift_data_reg[49]/NET0131  & n936 ;
  assign n1347 = \shift_data_reg[113]/NET0131  & n921 ;
  assign n1349 = ~n1346 & ~n1347 ;
  assign n1350 = n1348 & n1349 ;
  assign n1351 = \shift_data_reg[19]/NET0131  & n934 ;
  assign n1352 = \shift_data_reg[83]/NET0131  & n932 ;
  assign n1355 = ~n1351 & ~n1352 ;
  assign n1353 = \shift_data_reg[51]/NET0131  & n936 ;
  assign n1354 = \shift_data_reg[115]/NET0131  & n921 ;
  assign n1356 = ~n1353 & ~n1354 ;
  assign n1357 = n1355 & n1356 ;
  assign n1358 = \shift_data_reg[117]/NET0131  & n921 ;
  assign n1359 = \shift_data_reg[53]/NET0131  & n936 ;
  assign n1362 = ~n1358 & ~n1359 ;
  assign n1360 = \shift_data_reg[85]/NET0131  & n932 ;
  assign n1361 = \shift_data_reg[21]/NET0131  & n934 ;
  assign n1363 = ~n1360 & ~n1361 ;
  assign n1364 = n1362 & n1363 ;
  assign n1365 = \shift_data_reg[22]/NET0131  & n934 ;
  assign n1366 = \shift_data_reg[86]/NET0131  & n932 ;
  assign n1369 = ~n1365 & ~n1366 ;
  assign n1367 = \shift_data_reg[54]/NET0131  & n936 ;
  assign n1368 = \shift_data_reg[118]/NET0131  & n921 ;
  assign n1370 = ~n1367 & ~n1368 ;
  assign n1371 = n1369 & n1370 ;
  assign n1372 = wb_cyc_i_pad & wb_stb_i_pad ;
  assign n1373 = ~wb_ack_o_pad & n1372 ;
  assign n1385 = ~\ctrl_reg[9]/NET0131  & n280 ;
  assign n1384 = \ctrl_reg[9]/NET0131  & ~\shift_cnt_reg[1]/NET0131  ;
  assign n1386 = ~\ctrl_reg[11]/NET0131  & ~n1384 ;
  assign n1387 = ~n1385 & n1386 ;
  assign n1388 = \ctrl_reg[9]/NET0131  & ~\shift_cnt_reg[0]/NET0131  ;
  assign n1389 = ~\ctrl_reg[9]/NET0131  & \shift_cnt_reg[0]/NET0131  ;
  assign n1390 = ~n1388 & ~n1389 ;
  assign n1391 = ~\ctrl_reg[0]/NET0131  & ~n1390 ;
  assign n1392 = \ctrl_reg[9]/NET0131  & ~n280 ;
  assign n1393 = ~\ctrl_reg[9]/NET0131  & ~\shift_cnt_reg[1]/NET0131  ;
  assign n1394 = ~n1392 & ~n1393 ;
  assign n1395 = \ctrl_reg[1]/NET0131  & ~n1394 ;
  assign n1396 = ~\ctrl_reg[1]/NET0131  & n1394 ;
  assign n1397 = ~n1395 & ~n1396 ;
  assign n1399 = ~n1391 & n1397 ;
  assign n1398 = n1391 & ~n1397 ;
  assign n1400 = \ctrl_reg[11]/NET0131  & ~n1398 ;
  assign n1401 = ~n1399 & n1400 ;
  assign n1402 = ~n1387 & ~n1401 ;
  assign n1403 = ~n284 & n1390 ;
  assign n1404 = n284 & ~n1390 ;
  assign n1405 = ~n1403 & ~n1404 ;
  assign n1406 = ~n1402 & ~n1405 ;
  assign n1407 = ~n1391 & ~n1396 ;
  assign n1408 = ~n1395 & ~n1407 ;
  assign n1409 = \ctrl_reg[9]/NET0131  & n279 ;
  assign n1410 = ~\shift_cnt_reg[2]/NET0131  & ~n1409 ;
  assign n1411 = \shift_cnt_reg[2]/NET0131  & n1409 ;
  assign n1412 = ~n1410 & ~n1411 ;
  assign n1413 = \ctrl_reg[2]/NET0131  & ~n1412 ;
  assign n1414 = ~\ctrl_reg[2]/NET0131  & n1412 ;
  assign n1415 = ~n1413 & ~n1414 ;
  assign n1417 = n1408 & n1415 ;
  assign n1416 = ~n1408 & ~n1415 ;
  assign n1418 = \ctrl_reg[11]/NET0131  & ~n1416 ;
  assign n1419 = ~n1417 & n1418 ;
  assign n1421 = ~\ctrl_reg[9]/NET0131  & ~n256 ;
  assign n1420 = \ctrl_reg[9]/NET0131  & \shift_cnt_reg[2]/NET0131  ;
  assign n1422 = ~\ctrl_reg[11]/NET0131  & ~n1420 ;
  assign n1423 = ~n1421 & n1422 ;
  assign n1424 = ~n1419 & ~n1423 ;
  assign n1425 = n1406 & n1424 ;
  assign n1427 = ~\ctrl_reg[9]/NET0131  & n270 ;
  assign n1426 = \ctrl_reg[9]/NET0131  & ~\shift_cnt_reg[3]/NET0131  ;
  assign n1428 = ~\ctrl_reg[11]/NET0131  & ~n1426 ;
  assign n1429 = ~n1427 & n1428 ;
  assign n1430 = ~n1408 & ~n1414 ;
  assign n1431 = ~n1413 & ~n1430 ;
  assign n1432 = \shift_cnt_reg[3]/NET0131  & n1411 ;
  assign n1433 = ~\shift_cnt_reg[3]/NET0131  & ~n1411 ;
  assign n1434 = ~n1432 & ~n1433 ;
  assign n1435 = ~\ctrl_reg[3]/NET0131  & n1434 ;
  assign n1436 = \ctrl_reg[3]/NET0131  & ~n1434 ;
  assign n1437 = ~n1435 & ~n1436 ;
  assign n1439 = ~n1431 & n1437 ;
  assign n1438 = n1431 & ~n1437 ;
  assign n1440 = \ctrl_reg[11]/NET0131  & ~n1438 ;
  assign n1441 = ~n1439 & n1440 ;
  assign n1442 = ~n1429 & ~n1441 ;
  assign n1443 = n1425 & n1442 ;
  assign n1444 = \shift_cnt_reg[4]/NET0131  & n1432 ;
  assign n1445 = ~\shift_cnt_reg[4]/NET0131  & ~n1432 ;
  assign n1446 = ~n1444 & ~n1445 ;
  assign n1447 = ~\ctrl_reg[4]/NET0131  & n1446 ;
  assign n1450 = ~n1431 & ~n1435 ;
  assign n1448 = \ctrl_reg[4]/NET0131  & ~n1446 ;
  assign n1453 = ~n1436 & ~n1448 ;
  assign n1454 = ~n1450 & n1453 ;
  assign n1455 = ~n1447 & n1454 ;
  assign n1449 = ~n1447 & ~n1448 ;
  assign n1451 = ~n1436 & ~n1450 ;
  assign n1452 = ~n1449 & ~n1451 ;
  assign n1456 = \ctrl_reg[11]/NET0131  & ~n1452 ;
  assign n1457 = ~n1455 & n1456 ;
  assign n1459 = ~\ctrl_reg[9]/NET0131  & ~n341 ;
  assign n1458 = \ctrl_reg[9]/NET0131  & \shift_cnt_reg[4]/NET0131  ;
  assign n1460 = ~\ctrl_reg[11]/NET0131  & ~n1458 ;
  assign n1461 = ~n1459 & n1460 ;
  assign n1462 = ~n1457 & ~n1461 ;
  assign n1464 = ~\shift_cnt_reg[5]/NET0131  & ~n1444 ;
  assign n1465 = \shift_cnt_reg[5]/NET0131  & n1444 ;
  assign n1466 = ~n1464 & ~n1465 ;
  assign n1467 = \ctrl_reg[5]/NET0131  & ~n1466 ;
  assign n1463 = ~n1447 & ~n1454 ;
  assign n1468 = ~\ctrl_reg[5]/NET0131  & n1466 ;
  assign n1471 = n1463 & ~n1468 ;
  assign n1472 = ~n1467 & n1471 ;
  assign n1469 = ~n1467 & ~n1468 ;
  assign n1470 = ~n1463 & ~n1469 ;
  assign n1473 = \ctrl_reg[11]/NET0131  & ~n1470 ;
  assign n1474 = ~n1472 & n1473 ;
  assign n1476 = ~\ctrl_reg[9]/NET0131  & n358 ;
  assign n1475 = \ctrl_reg[9]/NET0131  & ~\shift_cnt_reg[5]/NET0131  ;
  assign n1477 = ~\ctrl_reg[11]/NET0131  & ~n1475 ;
  assign n1478 = ~n1476 & n1477 ;
  assign n1479 = ~n1474 & ~n1478 ;
  assign n1480 = n1462 & ~n1479 ;
  assign n1374 = ~\shift_tip_reg/NET0131  & ~\wb_adr_i[4]_pad  ;
  assign n1481 = \wb_adr_i[3]_pad  & wb_cyc_i_pad ;
  assign n1482 = n1374 & n1481 ;
  assign n1483 = n812 & n1482 ;
  assign n1484 = n1129 & n1482 ;
  assign n1485 = ~n1483 & ~n1484 ;
  assign n1486 = ~n1467 & ~n1471 ;
  assign n1487 = n507 & n1465 ;
  assign n1488 = ~n507 & ~n1465 ;
  assign n1489 = ~n1487 & ~n1488 ;
  assign n1491 = n1486 & ~n1489 ;
  assign n1490 = ~n1486 & n1489 ;
  assign n1492 = \ctrl_reg[11]/NET0131  & ~n1490 ;
  assign n1493 = ~n1491 & n1492 ;
  assign n1495 = ~\ctrl_reg[9]/NET0131  & n503 ;
  assign n1494 = \ctrl_reg[9]/NET0131  & ~\shift_cnt_reg[6]/NET0131  ;
  assign n1496 = ~\ctrl_reg[11]/NET0131  & ~n1494 ;
  assign n1497 = ~n1495 & n1496 ;
  assign n1498 = ~n1493 & ~n1497 ;
  assign n1499 = n1485 & n1498 ;
  assign n1500 = n1480 & n1499 ;
  assign n1501 = n1443 & n1500 ;
  assign n1854 = ~\shift_data_reg[17]/NET0131  & ~n1405 ;
  assign n1855 = ~\shift_data_reg[16]/NET0131  & n1405 ;
  assign n1856 = ~n1854 & ~n1855 ;
  assign n1857 = n1402 & n1856 ;
  assign n1850 = ~\shift_data_reg[19]/NET0131  & ~n1405 ;
  assign n1851 = ~\shift_data_reg[18]/NET0131  & n1405 ;
  assign n1852 = ~n1850 & ~n1851 ;
  assign n1853 = ~n1402 & n1852 ;
  assign n1858 = ~n1424 & ~n1853 ;
  assign n1859 = ~n1857 & n1858 ;
  assign n1844 = ~\shift_data_reg[23]/NET0131  & ~n1405 ;
  assign n1845 = ~\shift_data_reg[22]/NET0131  & n1405 ;
  assign n1846 = ~n1844 & ~n1845 ;
  assign n1847 = ~n1402 & n1846 ;
  assign n1840 = ~\shift_data_reg[21]/NET0131  & ~n1405 ;
  assign n1841 = ~\shift_data_reg[20]/NET0131  & n1405 ;
  assign n1842 = ~n1840 & ~n1841 ;
  assign n1843 = n1402 & n1842 ;
  assign n1848 = n1424 & ~n1843 ;
  assign n1849 = ~n1847 & n1848 ;
  assign n1860 = n1442 & ~n1849 ;
  assign n1861 = ~n1859 & n1860 ;
  assign n1876 = ~\shift_data_reg[25]/NET0131  & ~n1405 ;
  assign n1877 = ~\shift_data_reg[24]/NET0131  & n1405 ;
  assign n1878 = ~n1876 & ~n1877 ;
  assign n1879 = n1402 & n1878 ;
  assign n1872 = ~\shift_data_reg[27]/NET0131  & ~n1405 ;
  assign n1873 = ~\shift_data_reg[26]/NET0131  & n1405 ;
  assign n1874 = ~n1872 & ~n1873 ;
  assign n1875 = ~n1402 & n1874 ;
  assign n1880 = ~n1424 & ~n1875 ;
  assign n1881 = ~n1879 & n1880 ;
  assign n1866 = ~\shift_data_reg[31]/NET0131  & ~n1405 ;
  assign n1867 = ~\shift_data_reg[30]/NET0131  & n1405 ;
  assign n1868 = ~n1866 & ~n1867 ;
  assign n1869 = ~n1402 & n1868 ;
  assign n1862 = ~\shift_data_reg[29]/NET0131  & ~n1405 ;
  assign n1863 = ~\shift_data_reg[28]/NET0131  & n1405 ;
  assign n1864 = ~n1862 & ~n1863 ;
  assign n1865 = n1402 & n1864 ;
  assign n1870 = n1424 & ~n1865 ;
  assign n1871 = ~n1869 & n1870 ;
  assign n1882 = ~n1442 & ~n1871 ;
  assign n1883 = ~n1881 & n1882 ;
  assign n1884 = ~n1861 & ~n1883 ;
  assign n1885 = n1462 & ~n1884 ;
  assign n1808 = ~\shift_data_reg[9]/NET0131  & ~n1405 ;
  assign n1809 = ~\shift_data_reg[8]/NET0131  & n1405 ;
  assign n1810 = ~n1808 & ~n1809 ;
  assign n1811 = n1402 & n1810 ;
  assign n1804 = ~\shift_data_reg[11]/NET0131  & ~n1405 ;
  assign n1805 = ~\shift_data_reg[10]/NET0131  & n1405 ;
  assign n1806 = ~n1804 & ~n1805 ;
  assign n1807 = ~n1402 & n1806 ;
  assign n1812 = ~n1424 & ~n1807 ;
  assign n1813 = ~n1811 & n1812 ;
  assign n1798 = ~\shift_data_reg[15]/NET0131  & ~n1405 ;
  assign n1799 = ~\shift_data_reg[14]/NET0131  & n1405 ;
  assign n1800 = ~n1798 & ~n1799 ;
  assign n1801 = ~n1402 & n1800 ;
  assign n1794 = ~\shift_data_reg[13]/NET0131  & ~n1405 ;
  assign n1795 = ~\shift_data_reg[12]/NET0131  & n1405 ;
  assign n1796 = ~n1794 & ~n1795 ;
  assign n1797 = n1402 & n1796 ;
  assign n1802 = n1424 & ~n1797 ;
  assign n1803 = ~n1801 & n1802 ;
  assign n1814 = ~n1442 & ~n1803 ;
  assign n1815 = ~n1813 & n1814 ;
  assign n1830 = ~\shift_data_reg[1]/NET0131  & ~n1405 ;
  assign n1831 = ~\shift_data_reg[0]/NET0131  & n1405 ;
  assign n1832 = ~n1830 & ~n1831 ;
  assign n1833 = n1402 & n1832 ;
  assign n1826 = ~\shift_data_reg[3]/NET0131  & ~n1405 ;
  assign n1827 = ~\shift_data_reg[2]/NET0131  & n1405 ;
  assign n1828 = ~n1826 & ~n1827 ;
  assign n1829 = ~n1402 & n1828 ;
  assign n1834 = ~n1424 & ~n1829 ;
  assign n1835 = ~n1833 & n1834 ;
  assign n1820 = ~\shift_data_reg[7]/NET0131  & ~n1405 ;
  assign n1821 = ~\shift_data_reg[6]/NET0131  & n1405 ;
  assign n1822 = ~n1820 & ~n1821 ;
  assign n1823 = ~n1402 & n1822 ;
  assign n1816 = ~\shift_data_reg[5]/NET0131  & ~n1405 ;
  assign n1817 = ~\shift_data_reg[4]/NET0131  & n1405 ;
  assign n1818 = ~n1816 & ~n1817 ;
  assign n1819 = n1402 & n1818 ;
  assign n1824 = n1424 & ~n1819 ;
  assign n1825 = ~n1823 & n1824 ;
  assign n1836 = n1442 & ~n1825 ;
  assign n1837 = ~n1835 & n1836 ;
  assign n1838 = ~n1815 & ~n1837 ;
  assign n1839 = ~n1462 & ~n1838 ;
  assign n1886 = n1479 & ~n1839 ;
  assign n1887 = ~n1885 & n1886 ;
  assign n1760 = ~\shift_data_reg[57]/NET0131  & ~n1405 ;
  assign n1761 = ~\shift_data_reg[56]/NET0131  & n1405 ;
  assign n1762 = ~n1760 & ~n1761 ;
  assign n1763 = n1402 & n1762 ;
  assign n1756 = ~\shift_data_reg[59]/NET0131  & ~n1405 ;
  assign n1757 = ~\shift_data_reg[58]/NET0131  & n1405 ;
  assign n1758 = ~n1756 & ~n1757 ;
  assign n1759 = ~n1402 & n1758 ;
  assign n1764 = ~n1424 & ~n1759 ;
  assign n1765 = ~n1763 & n1764 ;
  assign n1750 = ~\shift_data_reg[63]/NET0131  & ~n1405 ;
  assign n1751 = ~\shift_data_reg[62]/NET0131  & n1405 ;
  assign n1752 = ~n1750 & ~n1751 ;
  assign n1753 = ~n1402 & n1752 ;
  assign n1746 = ~\shift_data_reg[61]/NET0131  & ~n1405 ;
  assign n1747 = ~\shift_data_reg[60]/NET0131  & n1405 ;
  assign n1748 = ~n1746 & ~n1747 ;
  assign n1749 = n1402 & n1748 ;
  assign n1754 = n1424 & ~n1749 ;
  assign n1755 = ~n1753 & n1754 ;
  assign n1766 = ~n1442 & ~n1755 ;
  assign n1767 = ~n1765 & n1766 ;
  assign n1782 = ~\shift_data_reg[53]/NET0131  & ~n1405 ;
  assign n1783 = ~\shift_data_reg[52]/NET0131  & n1405 ;
  assign n1784 = ~n1782 & ~n1783 ;
  assign n1785 = n1402 & n1784 ;
  assign n1778 = ~\shift_data_reg[55]/NET0131  & ~n1405 ;
  assign n1779 = ~\shift_data_reg[54]/NET0131  & n1405 ;
  assign n1780 = ~n1778 & ~n1779 ;
  assign n1781 = ~n1402 & n1780 ;
  assign n1786 = n1424 & ~n1781 ;
  assign n1787 = ~n1785 & n1786 ;
  assign n1772 = ~\shift_data_reg[51]/NET0131  & ~n1405 ;
  assign n1773 = ~\shift_data_reg[50]/NET0131  & n1405 ;
  assign n1774 = ~n1772 & ~n1773 ;
  assign n1775 = ~n1402 & n1774 ;
  assign n1768 = ~\shift_data_reg[49]/NET0131  & ~n1405 ;
  assign n1769 = ~\shift_data_reg[48]/NET0131  & n1405 ;
  assign n1770 = ~n1768 & ~n1769 ;
  assign n1771 = n1402 & n1770 ;
  assign n1776 = ~n1424 & ~n1771 ;
  assign n1777 = ~n1775 & n1776 ;
  assign n1788 = n1442 & ~n1777 ;
  assign n1789 = ~n1787 & n1788 ;
  assign n1790 = ~n1767 & ~n1789 ;
  assign n1791 = n1462 & ~n1790 ;
  assign n1714 = ~\shift_data_reg[41]/NET0131  & ~n1405 ;
  assign n1715 = ~\shift_data_reg[40]/NET0131  & n1405 ;
  assign n1716 = ~n1714 & ~n1715 ;
  assign n1717 = n1402 & n1716 ;
  assign n1710 = ~\shift_data_reg[43]/NET0131  & ~n1405 ;
  assign n1711 = ~\shift_data_reg[42]/NET0131  & n1405 ;
  assign n1712 = ~n1710 & ~n1711 ;
  assign n1713 = ~n1402 & n1712 ;
  assign n1718 = ~n1424 & ~n1713 ;
  assign n1719 = ~n1717 & n1718 ;
  assign n1704 = ~\shift_data_reg[47]/NET0131  & ~n1405 ;
  assign n1705 = ~\shift_data_reg[46]/NET0131  & n1405 ;
  assign n1706 = ~n1704 & ~n1705 ;
  assign n1707 = ~n1402 & n1706 ;
  assign n1700 = ~\shift_data_reg[45]/NET0131  & ~n1405 ;
  assign n1701 = ~\shift_data_reg[44]/NET0131  & n1405 ;
  assign n1702 = ~n1700 & ~n1701 ;
  assign n1703 = n1402 & n1702 ;
  assign n1708 = n1424 & ~n1703 ;
  assign n1709 = ~n1707 & n1708 ;
  assign n1720 = ~n1442 & ~n1709 ;
  assign n1721 = ~n1719 & n1720 ;
  assign n1736 = ~\shift_data_reg[39]/NET0131  & ~n1405 ;
  assign n1737 = ~\shift_data_reg[38]/NET0131  & n1405 ;
  assign n1738 = ~n1736 & ~n1737 ;
  assign n1739 = ~n1402 & n1738 ;
  assign n1732 = ~\shift_data_reg[37]/NET0131  & ~n1405 ;
  assign n1733 = ~\shift_data_reg[36]/NET0131  & n1405 ;
  assign n1734 = ~n1732 & ~n1733 ;
  assign n1735 = n1402 & n1734 ;
  assign n1740 = n1424 & ~n1735 ;
  assign n1741 = ~n1739 & n1740 ;
  assign n1726 = ~\shift_data_reg[33]/NET0131  & ~n1405 ;
  assign n1727 = ~\shift_data_reg[32]/NET0131  & n1405 ;
  assign n1728 = ~n1726 & ~n1727 ;
  assign n1729 = n1402 & n1728 ;
  assign n1722 = ~\shift_data_reg[35]/NET0131  & ~n1405 ;
  assign n1723 = ~\shift_data_reg[34]/NET0131  & n1405 ;
  assign n1724 = ~n1722 & ~n1723 ;
  assign n1725 = ~n1402 & n1724 ;
  assign n1730 = ~n1424 & ~n1725 ;
  assign n1731 = ~n1729 & n1730 ;
  assign n1742 = n1442 & ~n1731 ;
  assign n1743 = ~n1741 & n1742 ;
  assign n1744 = ~n1721 & ~n1743 ;
  assign n1745 = ~n1462 & ~n1744 ;
  assign n1792 = ~n1479 & ~n1745 ;
  assign n1793 = ~n1791 & n1792 ;
  assign n1505 = ~sclk_pad_o_pad & n704 ;
  assign n1503 = ~\clgen_pos_edge_reg/NET0131  & ~\ctrl_reg[9]/NET0131  ;
  assign n1504 = ~\clgen_neg_edge_reg/NET0131  & \ctrl_reg[9]/NET0131  ;
  assign n1506 = ~n1503 & ~n1504 ;
  assign n1507 = ~n1505 & n1506 ;
  assign n1888 = n1498 & ~n1507 ;
  assign n1889 = ~n1793 & n1888 ;
  assign n1890 = ~n1887 & n1889 ;
  assign n1508 = miso_pad_i_pad & n1507 ;
  assign n1663 = ~\shift_data_reg[81]/NET0131  & ~n1405 ;
  assign n1664 = ~\shift_data_reg[80]/NET0131  & n1405 ;
  assign n1665 = ~n1663 & ~n1664 ;
  assign n1666 = n1402 & n1665 ;
  assign n1659 = ~\shift_data_reg[83]/NET0131  & ~n1405 ;
  assign n1660 = ~\shift_data_reg[82]/NET0131  & n1405 ;
  assign n1661 = ~n1659 & ~n1660 ;
  assign n1662 = ~n1402 & n1661 ;
  assign n1667 = ~n1424 & ~n1662 ;
  assign n1668 = ~n1666 & n1667 ;
  assign n1653 = ~\shift_data_reg[87]/NET0131  & ~n1405 ;
  assign n1654 = ~\shift_data_reg[86]/NET0131  & n1405 ;
  assign n1655 = ~n1653 & ~n1654 ;
  assign n1656 = ~n1402 & n1655 ;
  assign n1649 = ~\shift_data_reg[85]/NET0131  & ~n1405 ;
  assign n1650 = ~\shift_data_reg[84]/NET0131  & n1405 ;
  assign n1651 = ~n1649 & ~n1650 ;
  assign n1652 = n1402 & n1651 ;
  assign n1657 = n1424 & ~n1652 ;
  assign n1658 = ~n1656 & n1657 ;
  assign n1669 = n1442 & ~n1658 ;
  assign n1670 = ~n1668 & n1669 ;
  assign n1685 = ~\shift_data_reg[89]/NET0131  & ~n1405 ;
  assign n1686 = ~\shift_data_reg[88]/NET0131  & n1405 ;
  assign n1687 = ~n1685 & ~n1686 ;
  assign n1688 = n1402 & n1687 ;
  assign n1681 = ~\shift_data_reg[91]/NET0131  & ~n1405 ;
  assign n1682 = ~\shift_data_reg[90]/NET0131  & n1405 ;
  assign n1683 = ~n1681 & ~n1682 ;
  assign n1684 = ~n1402 & n1683 ;
  assign n1689 = ~n1424 & ~n1684 ;
  assign n1690 = ~n1688 & n1689 ;
  assign n1675 = ~\shift_data_reg[95]/NET0131  & ~n1405 ;
  assign n1676 = ~\shift_data_reg[94]/NET0131  & n1405 ;
  assign n1677 = ~n1675 & ~n1676 ;
  assign n1678 = ~n1402 & n1677 ;
  assign n1671 = ~\shift_data_reg[93]/NET0131  & ~n1405 ;
  assign n1672 = ~\shift_data_reg[92]/NET0131  & n1405 ;
  assign n1673 = ~n1671 & ~n1672 ;
  assign n1674 = n1402 & n1673 ;
  assign n1679 = n1424 & ~n1674 ;
  assign n1680 = ~n1678 & n1679 ;
  assign n1691 = ~n1442 & ~n1680 ;
  assign n1692 = ~n1690 & n1691 ;
  assign n1693 = ~n1670 & ~n1692 ;
  assign n1694 = n1462 & ~n1693 ;
  assign n1617 = ~\shift_data_reg[73]/NET0131  & ~n1405 ;
  assign n1618 = ~\shift_data_reg[72]/NET0131  & n1405 ;
  assign n1619 = ~n1617 & ~n1618 ;
  assign n1620 = n1402 & n1619 ;
  assign n1613 = ~\shift_data_reg[75]/NET0131  & ~n1405 ;
  assign n1614 = ~\shift_data_reg[74]/NET0131  & n1405 ;
  assign n1615 = ~n1613 & ~n1614 ;
  assign n1616 = ~n1402 & n1615 ;
  assign n1621 = ~n1424 & ~n1616 ;
  assign n1622 = ~n1620 & n1621 ;
  assign n1607 = ~\shift_data_reg[79]/NET0131  & ~n1405 ;
  assign n1608 = ~\shift_data_reg[78]/NET0131  & n1405 ;
  assign n1609 = ~n1607 & ~n1608 ;
  assign n1610 = ~n1402 & n1609 ;
  assign n1603 = ~\shift_data_reg[77]/NET0131  & ~n1405 ;
  assign n1604 = ~\shift_data_reg[76]/NET0131  & n1405 ;
  assign n1605 = ~n1603 & ~n1604 ;
  assign n1606 = n1402 & n1605 ;
  assign n1611 = n1424 & ~n1606 ;
  assign n1612 = ~n1610 & n1611 ;
  assign n1623 = ~n1442 & ~n1612 ;
  assign n1624 = ~n1622 & n1623 ;
  assign n1639 = ~\shift_data_reg[65]/NET0131  & ~n1405 ;
  assign n1640 = ~\shift_data_reg[64]/NET0131  & n1405 ;
  assign n1641 = ~n1639 & ~n1640 ;
  assign n1642 = n1402 & n1641 ;
  assign n1635 = ~\shift_data_reg[67]/NET0131  & ~n1405 ;
  assign n1636 = ~\shift_data_reg[66]/NET0131  & n1405 ;
  assign n1637 = ~n1635 & ~n1636 ;
  assign n1638 = ~n1402 & n1637 ;
  assign n1643 = ~n1424 & ~n1638 ;
  assign n1644 = ~n1642 & n1643 ;
  assign n1629 = ~\shift_data_reg[71]/NET0131  & ~n1405 ;
  assign n1630 = ~\shift_data_reg[70]/NET0131  & n1405 ;
  assign n1631 = ~n1629 & ~n1630 ;
  assign n1632 = ~n1402 & n1631 ;
  assign n1625 = ~\shift_data_reg[69]/NET0131  & ~n1405 ;
  assign n1626 = ~\shift_data_reg[68]/NET0131  & n1405 ;
  assign n1627 = ~n1625 & ~n1626 ;
  assign n1628 = n1402 & n1627 ;
  assign n1633 = n1424 & ~n1628 ;
  assign n1634 = ~n1632 & n1633 ;
  assign n1645 = n1442 & ~n1634 ;
  assign n1646 = ~n1644 & n1645 ;
  assign n1647 = ~n1624 & ~n1646 ;
  assign n1648 = ~n1462 & ~n1647 ;
  assign n1695 = n1479 & ~n1648 ;
  assign n1696 = ~n1694 & n1695 ;
  assign n1545 = ~\shift_data_reg[116]/NET0131  & n1405 ;
  assign n1546 = ~\shift_data_reg[117]/NET0131  & ~n1405 ;
  assign n1547 = ~n1545 & ~n1546 ;
  assign n1548 = n1402 & n1547 ;
  assign n1541 = ~\shift_data_reg[118]/NET0131  & n1405 ;
  assign n1542 = ~\shift_data_reg[119]/NET0131  & ~n1405 ;
  assign n1543 = ~n1541 & ~n1542 ;
  assign n1544 = ~n1402 & n1543 ;
  assign n1549 = n1424 & ~n1544 ;
  assign n1550 = ~n1548 & n1549 ;
  assign n1535 = ~\shift_data_reg[114]/NET0131  & n1405 ;
  assign n1536 = ~\shift_data_reg[115]/NET0131  & ~n1405 ;
  assign n1537 = ~n1535 & ~n1536 ;
  assign n1538 = ~n1402 & n1537 ;
  assign n1531 = ~\shift_data_reg[112]/NET0131  & n1405 ;
  assign n1532 = ~\shift_data_reg[113]/NET0131  & ~n1405 ;
  assign n1533 = ~n1531 & ~n1532 ;
  assign n1534 = n1402 & n1533 ;
  assign n1539 = ~n1424 & ~n1534 ;
  assign n1540 = ~n1538 & n1539 ;
  assign n1551 = n1442 & ~n1540 ;
  assign n1552 = ~n1550 & n1551 ;
  assign n1523 = ~\shift_data_reg[124]/NET0131  & n1405 ;
  assign n1524 = ~\shift_data_reg[125]/NET0131  & ~n1405 ;
  assign n1525 = ~n1523 & ~n1524 ;
  assign n1526 = n1402 & n1525 ;
  assign n1519 = ~\shift_data_reg[126]/NET0131  & n1405 ;
  assign n1520 = ~\shift_data_reg[127]/NET0131  & ~n1405 ;
  assign n1521 = ~n1519 & ~n1520 ;
  assign n1522 = ~n1402 & n1521 ;
  assign n1527 = n1424 & ~n1522 ;
  assign n1528 = ~n1526 & n1527 ;
  assign n1513 = ~\shift_data_reg[122]/NET0131  & n1405 ;
  assign n1514 = ~\shift_data_reg[123]/NET0131  & ~n1405 ;
  assign n1515 = ~n1513 & ~n1514 ;
  assign n1516 = ~n1402 & n1515 ;
  assign n1509 = ~\shift_data_reg[120]/NET0131  & n1405 ;
  assign n1510 = ~\shift_data_reg[121]/NET0131  & ~n1405 ;
  assign n1511 = ~n1509 & ~n1510 ;
  assign n1512 = n1402 & n1511 ;
  assign n1517 = ~n1424 & ~n1512 ;
  assign n1518 = ~n1516 & n1517 ;
  assign n1529 = ~n1442 & ~n1518 ;
  assign n1530 = ~n1528 & n1529 ;
  assign n1553 = n1462 & ~n1530 ;
  assign n1554 = ~n1552 & n1553 ;
  assign n1591 = ~\shift_data_reg[108]/NET0131  & n1405 ;
  assign n1592 = ~\shift_data_reg[109]/NET0131  & ~n1405 ;
  assign n1593 = ~n1591 & ~n1592 ;
  assign n1594 = n1402 & n1593 ;
  assign n1587 = ~\shift_data_reg[110]/NET0131  & n1405 ;
  assign n1588 = ~\shift_data_reg[111]/NET0131  & ~n1405 ;
  assign n1589 = ~n1587 & ~n1588 ;
  assign n1590 = ~n1402 & n1589 ;
  assign n1595 = n1424 & ~n1590 ;
  assign n1596 = ~n1594 & n1595 ;
  assign n1581 = ~\shift_data_reg[106]/NET0131  & n1405 ;
  assign n1582 = ~\shift_data_reg[107]/NET0131  & ~n1405 ;
  assign n1583 = ~n1581 & ~n1582 ;
  assign n1584 = ~n1402 & n1583 ;
  assign n1577 = ~\shift_data_reg[104]/NET0131  & n1405 ;
  assign n1578 = ~\shift_data_reg[105]/NET0131  & ~n1405 ;
  assign n1579 = ~n1577 & ~n1578 ;
  assign n1580 = n1402 & n1579 ;
  assign n1585 = ~n1424 & ~n1580 ;
  assign n1586 = ~n1584 & n1585 ;
  assign n1597 = ~n1442 & ~n1586 ;
  assign n1598 = ~n1596 & n1597 ;
  assign n1569 = ~\shift_data_reg[100]/NET0131  & n1405 ;
  assign n1570 = ~\shift_data_reg[101]/NET0131  & ~n1405 ;
  assign n1571 = ~n1569 & ~n1570 ;
  assign n1572 = n1402 & n1571 ;
  assign n1565 = ~\shift_data_reg[102]/NET0131  & n1405 ;
  assign n1566 = ~\shift_data_reg[103]/NET0131  & ~n1405 ;
  assign n1567 = ~n1565 & ~n1566 ;
  assign n1568 = ~n1402 & n1567 ;
  assign n1573 = n1424 & ~n1568 ;
  assign n1574 = ~n1572 & n1573 ;
  assign n1559 = ~\shift_data_reg[98]/NET0131  & n1405 ;
  assign n1560 = ~\shift_data_reg[99]/NET0131  & ~n1405 ;
  assign n1561 = ~n1559 & ~n1560 ;
  assign n1562 = ~n1402 & n1561 ;
  assign n1555 = ~\shift_data_reg[96]/NET0131  & n1405 ;
  assign n1556 = ~\shift_data_reg[97]/NET0131  & ~n1405 ;
  assign n1557 = ~n1555 & ~n1556 ;
  assign n1558 = n1402 & n1557 ;
  assign n1563 = ~n1424 & ~n1558 ;
  assign n1564 = ~n1562 & n1563 ;
  assign n1575 = n1442 & ~n1564 ;
  assign n1576 = ~n1574 & n1575 ;
  assign n1599 = ~n1462 & ~n1576 ;
  assign n1600 = ~n1598 & n1599 ;
  assign n1601 = ~n1554 & ~n1600 ;
  assign n1602 = ~n1479 & ~n1601 ;
  assign n1697 = ~n1498 & ~n1507 ;
  assign n1698 = ~n1602 & n1697 ;
  assign n1699 = ~n1696 & n1698 ;
  assign n1891 = ~n1508 & ~n1699 ;
  assign n1892 = ~n1890 & n1891 ;
  assign n1893 = n1501 & n1892 ;
  assign n1375 = ~\wb_adr_i[3]_pad  & wb_we_i_pad ;
  assign n1376 = n1372 & n1375 ;
  assign n1377 = n1374 & n1376 ;
  assign n1502 = ~\shift_data_reg[55]/NET0131  & ~n1501 ;
  assign n1894 = ~n1377 & ~n1502 ;
  assign n1895 = ~n1893 & n1894 ;
  assign n1378 = \wb_adr_i[2]_pad  & n1377 ;
  assign n1379 = \wb_dat_i[23]_pad  & \wb_sel_i[2]_pad  ;
  assign n1380 = n1378 & n1379 ;
  assign n1381 = \wb_adr_i[2]_pad  & \wb_sel_i[2]_pad  ;
  assign n1382 = n1377 & ~n1381 ;
  assign n1383 = \shift_data_reg[55]/NET0131  & n1382 ;
  assign n1896 = ~n1380 & ~n1383 ;
  assign n1897 = ~n1895 & n1896 ;
  assign n1898 = n1156 & n1484 ;
  assign n1899 = n1485 & ~n1892 ;
  assign n1900 = n1402 & ~n1405 ;
  assign n1901 = n1424 & n1900 ;
  assign n1902 = ~n1462 & ~n1479 ;
  assign n1903 = n1442 & ~n1498 ;
  assign n1904 = n1902 & n1903 ;
  assign n1905 = n1901 & n1904 ;
  assign n1906 = n1899 & n1905 ;
  assign n1907 = ~n1898 & ~n1906 ;
  assign n1908 = ~n1377 & ~n1907 ;
  assign n1909 = ~n1484 & ~n1905 ;
  assign n1910 = ~n1377 & ~n1483 ;
  assign n1911 = ~\wb_sel_i[0]_pad  & n1484 ;
  assign n1912 = n1910 & ~n1911 ;
  assign n1913 = ~n1909 & n1912 ;
  assign n1914 = \shift_data_reg[101]/NET0131  & ~n1913 ;
  assign n1915 = ~n1908 & ~n1914 ;
  assign n1922 = ~n1498 & n1902 ;
  assign n1923 = ~n1442 & n1922 ;
  assign n1924 = n1901 & n1923 ;
  assign n1925 = n1892 & n1924 ;
  assign n1921 = ~n1377 & n1485 ;
  assign n1926 = ~\shift_data_reg[109]/NET0131  & ~n1924 ;
  assign n1927 = n1921 & ~n1926 ;
  assign n1928 = ~n1925 & n1927 ;
  assign n1916 = \shift_data_reg[109]/NET0131  & ~n1910 ;
  assign n1917 = \shift_data_reg[109]/NET0131  & ~\wb_sel_i[1]_pad  ;
  assign n1918 = n1152 & ~n1377 ;
  assign n1919 = ~n1917 & ~n1918 ;
  assign n1920 = n1484 & ~n1919 ;
  assign n1929 = ~n1916 & ~n1920 ;
  assign n1930 = ~n1928 & n1929 ;
  assign n1936 = ~n1402 & n1405 ;
  assign n1937 = n1424 & n1936 ;
  assign n1938 = n1923 & n1937 ;
  assign n1939 = n1892 & n1938 ;
  assign n1940 = ~\shift_data_reg[110]/NET0131  & ~n1938 ;
  assign n1941 = n1921 & ~n1940 ;
  assign n1942 = ~n1939 & n1941 ;
  assign n1931 = \shift_data_reg[110]/NET0131  & ~n1910 ;
  assign n1932 = \shift_data_reg[110]/NET0131  & ~\wb_sel_i[1]_pad  ;
  assign n1933 = n1175 & ~n1377 ;
  assign n1934 = ~n1932 & ~n1933 ;
  assign n1935 = n1484 & ~n1934 ;
  assign n1943 = ~n1931 & ~n1935 ;
  assign n1944 = ~n1942 & n1943 ;
  assign n1949 = n1402 & n1405 ;
  assign n1950 = ~n1424 & n1949 ;
  assign n1951 = n1442 & n1499 ;
  assign n1952 = n1902 & n1951 ;
  assign n1953 = n1950 & n1952 ;
  assign n1955 = n1892 & n1953 ;
  assign n1954 = ~\shift_data_reg[32]/NET0131  & ~n1953 ;
  assign n1956 = ~n1377 & ~n1954 ;
  assign n1957 = ~n1955 & n1956 ;
  assign n1945 = n1220 & n1378 ;
  assign n1946 = \wb_adr_i[2]_pad  & \wb_sel_i[0]_pad  ;
  assign n1947 = n1377 & ~n1946 ;
  assign n1948 = \shift_data_reg[32]/NET0131  & n1947 ;
  assign n1958 = ~n1945 & ~n1948 ;
  assign n1959 = ~n1957 & n1958 ;
  assign n1962 = n1425 & n1952 ;
  assign n1964 = n1892 & n1962 ;
  assign n1963 = ~\shift_data_reg[39]/NET0131  & ~n1962 ;
  assign n1965 = ~n1377 & ~n1963 ;
  assign n1966 = ~n1964 & n1965 ;
  assign n1960 = n1148 & n1378 ;
  assign n1961 = \shift_data_reg[39]/NET0131  & n1947 ;
  assign n1967 = ~n1960 & ~n1961 ;
  assign n1968 = ~n1966 & n1967 ;
  assign n1974 = ~n1442 & n1499 ;
  assign n1975 = n1480 & n1974 ;
  assign n1976 = n1425 & n1975 ;
  assign n1978 = n1892 & n1976 ;
  assign n1977 = ~\shift_data_reg[63]/NET0131  & ~n1976 ;
  assign n1979 = ~n1377 & ~n1977 ;
  assign n1980 = ~n1978 & n1979 ;
  assign n1969 = \wb_dat_i[31]_pad  & \wb_sel_i[3]_pad  ;
  assign n1970 = n1378 & n1969 ;
  assign n1971 = \wb_adr_i[2]_pad  & \wb_sel_i[3]_pad  ;
  assign n1972 = n1377 & ~n1971 ;
  assign n1973 = \shift_data_reg[63]/NET0131  & n1972 ;
  assign n1981 = ~n1970 & ~n1973 ;
  assign n1982 = ~n1980 & n1981 ;
  assign n1986 = n1950 & n1975 ;
  assign n1988 = n1892 & n1986 ;
  assign n1987 = ~\shift_data_reg[56]/NET0131  & ~n1986 ;
  assign n1989 = ~n1377 & ~n1987 ;
  assign n1990 = ~n1988 & n1989 ;
  assign n1983 = \wb_dat_i[24]_pad  & \wb_sel_i[3]_pad  ;
  assign n1984 = n1378 & n1983 ;
  assign n1985 = \shift_data_reg[56]/NET0131  & n1972 ;
  assign n1991 = ~n1984 & ~n1985 ;
  assign n1992 = ~n1990 & n1991 ;
  assign n1993 = \shift_data_reg[89]/NET0131  & n1377 ;
  assign n1994 = ~\wb_adr_i[2]_pad  & n1377 ;
  assign n1995 = \shift_data_reg[89]/NET0131  & ~\wb_sel_i[3]_pad  ;
  assign n1996 = \wb_dat_i[25]_pad  & \wb_sel_i[3]_pad  ;
  assign n1997 = ~n1995 & ~n1996 ;
  assign n1998 = n1483 & ~n1997 ;
  assign n1999 = ~n1484 & ~n1498 ;
  assign n2000 = n1462 & n1479 ;
  assign n2001 = n1999 & n2000 ;
  assign n2002 = ~n1442 & n2001 ;
  assign n2003 = ~n1424 & n1900 ;
  assign n2004 = n2002 & n2003 ;
  assign n2005 = n1892 & n2004 ;
  assign n2006 = ~n1378 & ~n1483 ;
  assign n2007 = ~\shift_data_reg[89]/NET0131  & ~n2004 ;
  assign n2008 = n2006 & ~n2007 ;
  assign n2009 = ~n2005 & n2008 ;
  assign n2010 = ~n1998 & ~n2009 ;
  assign n2011 = ~n1994 & ~n2010 ;
  assign n2012 = ~n1993 & ~n2011 ;
  assign n2013 = \shift_data_reg[92]/NET0131  & ~\wb_sel_i[3]_pad  ;
  assign n2014 = \wb_dat_i[28]_pad  & \wb_sel_i[3]_pad  ;
  assign n2015 = ~n2013 & ~n2014 ;
  assign n2016 = n1483 & ~n2015 ;
  assign n2017 = n1424 & n1949 ;
  assign n2018 = n2002 & n2017 ;
  assign n2019 = n1892 & n2018 ;
  assign n2020 = ~\shift_data_reg[92]/NET0131  & ~n2018 ;
  assign n2021 = n2006 & ~n2020 ;
  assign n2022 = ~n2019 & n2021 ;
  assign n2023 = ~n2016 & ~n2022 ;
  assign n2024 = ~n1994 & ~n2023 ;
  assign n2025 = \shift_data_reg[92]/NET0131  & n1377 ;
  assign n2026 = ~n2024 & ~n2025 ;
  assign n2027 = \shift_data_reg[64]/NET0131  & ~\wb_sel_i[0]_pad  ;
  assign n2028 = ~n1220 & ~n2027 ;
  assign n2029 = n1483 & ~n2028 ;
  assign n2030 = n1442 & n1950 ;
  assign n2031 = ~n1462 & n1479 ;
  assign n2032 = n1999 & n2031 ;
  assign n2033 = n2030 & n2032 ;
  assign n2034 = n1892 & n2033 ;
  assign n2035 = ~\shift_data_reg[64]/NET0131  & ~n2033 ;
  assign n2036 = n2006 & ~n2035 ;
  assign n2037 = ~n2034 & n2036 ;
  assign n2038 = ~n2029 & ~n2037 ;
  assign n2039 = ~n1994 & ~n2038 ;
  assign n2040 = \shift_data_reg[64]/NET0131  & n1377 ;
  assign n2041 = ~n2039 & ~n2040 ;
  assign n2042 = \shift_data_reg[65]/NET0131  & ~\wb_sel_i[0]_pad  ;
  assign n2043 = ~n1189 & ~n2042 ;
  assign n2044 = n1483 & ~n2043 ;
  assign n2045 = n1442 & n2003 ;
  assign n2046 = n2032 & n2045 ;
  assign n2047 = n1892 & n2046 ;
  assign n2048 = ~\shift_data_reg[65]/NET0131  & ~n2046 ;
  assign n2049 = n2006 & ~n2048 ;
  assign n2050 = ~n2047 & n2049 ;
  assign n2051 = ~n2044 & ~n2050 ;
  assign n2052 = ~n1994 & ~n2051 ;
  assign n2053 = \shift_data_reg[65]/NET0131  & n1377 ;
  assign n2054 = ~n2052 & ~n2053 ;
  assign n2055 = \shift_data_reg[66]/NET0131  & ~\wb_sel_i[0]_pad  ;
  assign n2056 = ~n1163 & ~n2055 ;
  assign n2057 = n1483 & ~n2056 ;
  assign n2058 = ~n1424 & n1936 ;
  assign n2059 = n1442 & n2058 ;
  assign n2060 = n2032 & n2059 ;
  assign n2061 = n1892 & n2060 ;
  assign n2062 = ~\shift_data_reg[66]/NET0131  & ~n2060 ;
  assign n2063 = n2006 & ~n2062 ;
  assign n2064 = ~n2061 & n2063 ;
  assign n2065 = ~n2057 & ~n2064 ;
  assign n2066 = ~n1994 & ~n2065 ;
  assign n2067 = \shift_data_reg[66]/NET0131  & n1377 ;
  assign n2068 = ~n2066 & ~n2067 ;
  assign n2069 = \shift_data_reg[67]/NET0131  & ~\wb_sel_i[0]_pad  ;
  assign n2070 = ~n1199 & ~n2069 ;
  assign n2071 = n1483 & ~n2070 ;
  assign n2072 = n1406 & ~n1424 ;
  assign n2073 = n1442 & n2032 ;
  assign n2074 = n2072 & n2073 ;
  assign n2075 = n1892 & n2074 ;
  assign n2076 = ~\shift_data_reg[67]/NET0131  & ~n2074 ;
  assign n2077 = n2006 & ~n2076 ;
  assign n2078 = ~n2075 & n2077 ;
  assign n2079 = ~n2071 & ~n2078 ;
  assign n2080 = ~n1994 & ~n2079 ;
  assign n2081 = \shift_data_reg[67]/NET0131  & n1377 ;
  assign n2082 = ~n2080 & ~n2081 ;
  assign n2083 = \shift_data_reg[68]/NET0131  & ~\wb_sel_i[0]_pad  ;
  assign n2084 = ~n1133 & ~n2083 ;
  assign n2085 = n1483 & ~n2084 ;
  assign n2086 = n1442 & n2017 ;
  assign n2087 = n2032 & n2086 ;
  assign n2088 = n1892 & n2087 ;
  assign n2089 = ~\shift_data_reg[68]/NET0131  & ~n2087 ;
  assign n2090 = n2006 & ~n2089 ;
  assign n2091 = ~n2088 & n2090 ;
  assign n2092 = ~n2085 & ~n2091 ;
  assign n2093 = ~n1994 & ~n2092 ;
  assign n2094 = \shift_data_reg[68]/NET0131  & n1377 ;
  assign n2095 = ~n2093 & ~n2094 ;
  assign n2096 = \shift_data_reg[69]/NET0131  & ~\wb_sel_i[0]_pad  ;
  assign n2097 = ~n1156 & ~n2096 ;
  assign n2098 = n1483 & ~n2097 ;
  assign n2099 = n1901 & n2073 ;
  assign n2100 = n1892 & n2099 ;
  assign n2101 = ~\shift_data_reg[69]/NET0131  & ~n2099 ;
  assign n2102 = n2006 & ~n2101 ;
  assign n2103 = ~n2100 & n2102 ;
  assign n2104 = ~n2098 & ~n2103 ;
  assign n2105 = ~n1994 & ~n2104 ;
  assign n2106 = \shift_data_reg[69]/NET0131  & n1377 ;
  assign n2107 = ~n2105 & ~n2106 ;
  assign n2108 = \shift_data_reg[70]/NET0131  & n1377 ;
  assign n2109 = \shift_data_reg[70]/NET0131  & ~\wb_sel_i[0]_pad  ;
  assign n2110 = ~n1179 & ~n2109 ;
  assign n2111 = n1483 & ~n2110 ;
  assign n2112 = n1937 & n2073 ;
  assign n2113 = n1892 & n2112 ;
  assign n2114 = ~\shift_data_reg[70]/NET0131  & ~n2112 ;
  assign n2115 = n2006 & ~n2114 ;
  assign n2116 = ~n2113 & n2115 ;
  assign n2117 = ~n2111 & ~n2116 ;
  assign n2118 = ~n1994 & ~n2117 ;
  assign n2119 = ~n2108 & ~n2118 ;
  assign n2120 = \shift_data_reg[71]/NET0131  & ~\wb_sel_i[0]_pad  ;
  assign n2121 = ~n1148 & ~n2120 ;
  assign n2122 = n1483 & ~n2121 ;
  assign n2123 = n1442 & n2031 ;
  assign n2124 = n1425 & n2123 ;
  assign n2125 = n1999 & n2124 ;
  assign n2126 = n1892 & n2125 ;
  assign n2127 = ~\shift_data_reg[71]/NET0131  & ~n2125 ;
  assign n2128 = n2006 & ~n2127 ;
  assign n2129 = ~n2126 & n2128 ;
  assign n2130 = ~n2122 & ~n2129 ;
  assign n2131 = ~n1994 & ~n2130 ;
  assign n2132 = \shift_data_reg[71]/NET0131  & n1377 ;
  assign n2133 = ~n2131 & ~n2132 ;
  assign n2134 = \shift_data_reg[72]/NET0131  & ~\wb_sel_i[1]_pad  ;
  assign n2135 = ~n809 & ~n2134 ;
  assign n2136 = n1483 & ~n2135 ;
  assign n2137 = ~n1442 & n2032 ;
  assign n2138 = n1950 & n2137 ;
  assign n2139 = n1892 & n2138 ;
  assign n2140 = ~\shift_data_reg[72]/NET0131  & ~n2138 ;
  assign n2141 = n2006 & ~n2140 ;
  assign n2142 = ~n2139 & n2141 ;
  assign n2143 = ~n2136 & ~n2142 ;
  assign n2144 = ~n1994 & ~n2143 ;
  assign n2145 = \shift_data_reg[72]/NET0131  & n1377 ;
  assign n2146 = ~n2144 & ~n2145 ;
  assign n2147 = \shift_data_reg[74]/NET0131  & ~\wb_sel_i[1]_pad  ;
  assign n2148 = ~n1144 & ~n2147 ;
  assign n2149 = n1483 & ~n2148 ;
  assign n2150 = ~n1442 & n2058 ;
  assign n2151 = n2032 & n2150 ;
  assign n2152 = n1892 & n2151 ;
  assign n2153 = ~\shift_data_reg[74]/NET0131  & ~n2151 ;
  assign n2154 = n2006 & ~n2153 ;
  assign n2155 = ~n2152 & n2154 ;
  assign n2156 = ~n2149 & ~n2155 ;
  assign n2157 = ~n1994 & ~n2156 ;
  assign n2158 = \shift_data_reg[74]/NET0131  & n1377 ;
  assign n2159 = ~n2157 & ~n2158 ;
  assign n2160 = \shift_data_reg[75]/NET0131  & ~\wb_sel_i[1]_pad  ;
  assign n2161 = ~n1171 & ~n2160 ;
  assign n2162 = n1483 & ~n2161 ;
  assign n2163 = n2072 & n2137 ;
  assign n2164 = n1892 & n2163 ;
  assign n2165 = ~\shift_data_reg[75]/NET0131  & ~n2163 ;
  assign n2166 = n2006 & ~n2165 ;
  assign n2167 = ~n2164 & n2166 ;
  assign n2168 = ~n2162 & ~n2167 ;
  assign n2169 = ~n1994 & ~n2168 ;
  assign n2170 = \shift_data_reg[75]/NET0131  & n1377 ;
  assign n2171 = ~n2169 & ~n2170 ;
  assign n2172 = \shift_data_reg[73]/NET0131  & ~\wb_sel_i[1]_pad  ;
  assign n2173 = ~n1216 & ~n2172 ;
  assign n2174 = n1483 & ~n2173 ;
  assign n2175 = ~n1442 & n2031 ;
  assign n2176 = n2003 & n2175 ;
  assign n2177 = n1999 & n2176 ;
  assign n2178 = n1892 & n2177 ;
  assign n2179 = ~\shift_data_reg[73]/NET0131  & ~n2177 ;
  assign n2180 = n2006 & ~n2179 ;
  assign n2181 = ~n2178 & n2180 ;
  assign n2182 = ~n2174 & ~n2181 ;
  assign n2183 = ~n1994 & ~n2182 ;
  assign n2184 = \shift_data_reg[73]/NET0131  & n1377 ;
  assign n2185 = ~n2183 & ~n2184 ;
  assign n2186 = \shift_data_reg[76]/NET0131  & ~\wb_sel_i[1]_pad  ;
  assign n2187 = ~n1209 & ~n2186 ;
  assign n2188 = n1483 & ~n2187 ;
  assign n2189 = n2017 & n2137 ;
  assign n2190 = n1892 & n2189 ;
  assign n2191 = ~\shift_data_reg[76]/NET0131  & ~n2189 ;
  assign n2192 = n2006 & ~n2191 ;
  assign n2193 = ~n2190 & n2192 ;
  assign n2194 = ~n2188 & ~n2193 ;
  assign n2195 = ~n1994 & ~n2194 ;
  assign n2196 = \shift_data_reg[76]/NET0131  & n1377 ;
  assign n2197 = ~n2195 & ~n2196 ;
  assign n2198 = \shift_data_reg[77]/NET0131  & ~\wb_sel_i[1]_pad  ;
  assign n2199 = ~n1152 & ~n2198 ;
  assign n2200 = n1483 & ~n2199 ;
  assign n2201 = n1901 & n2137 ;
  assign n2202 = n1892 & n2201 ;
  assign n2203 = ~\shift_data_reg[77]/NET0131  & ~n2201 ;
  assign n2204 = n2006 & ~n2203 ;
  assign n2205 = ~n2202 & n2204 ;
  assign n2206 = ~n2200 & ~n2205 ;
  assign n2207 = ~n1994 & ~n2206 ;
  assign n2208 = \shift_data_reg[77]/NET0131  & n1377 ;
  assign n2209 = ~n2207 & ~n2208 ;
  assign n2210 = \shift_data_reg[78]/NET0131  & ~\wb_sel_i[1]_pad  ;
  assign n2211 = ~n1175 & ~n2210 ;
  assign n2212 = n1483 & ~n2211 ;
  assign n2213 = n1937 & n2137 ;
  assign n2214 = n1892 & n2213 ;
  assign n2215 = ~\shift_data_reg[78]/NET0131  & ~n2213 ;
  assign n2216 = n2006 & ~n2215 ;
  assign n2217 = ~n2214 & n2216 ;
  assign n2218 = ~n2212 & ~n2217 ;
  assign n2219 = ~n1994 & ~n2218 ;
  assign n2220 = \shift_data_reg[78]/NET0131  & n1377 ;
  assign n2221 = ~n2219 & ~n2220 ;
  assign n2222 = \shift_data_reg[79]/NET0131  & ~\wb_sel_i[1]_pad  ;
  assign n2223 = ~n1230 & ~n2222 ;
  assign n2224 = n1483 & ~n2223 ;
  assign n2225 = n1425 & ~n1442 ;
  assign n2226 = n2032 & n2225 ;
  assign n2227 = n1892 & n2226 ;
  assign n2228 = ~\shift_data_reg[79]/NET0131  & ~n2226 ;
  assign n2229 = n2006 & ~n2228 ;
  assign n2230 = ~n2227 & n2229 ;
  assign n2231 = ~n2224 & ~n2230 ;
  assign n2232 = ~n1994 & ~n2231 ;
  assign n2233 = \shift_data_reg[79]/NET0131  & n1377 ;
  assign n2234 = ~n2232 & ~n2233 ;
  assign n2235 = \shift_data_reg[81]/NET0131  & ~\wb_sel_i[2]_pad  ;
  assign n2236 = \wb_dat_i[17]_pad  & \wb_sel_i[2]_pad  ;
  assign n2237 = ~n2235 & ~n2236 ;
  assign n2238 = n1483 & ~n2237 ;
  assign n2239 = n2001 & n2045 ;
  assign n2240 = n1892 & n2239 ;
  assign n2241 = ~\shift_data_reg[81]/NET0131  & ~n2239 ;
  assign n2242 = n2006 & ~n2241 ;
  assign n2243 = ~n2240 & n2242 ;
  assign n2244 = ~n2238 & ~n2243 ;
  assign n2245 = ~n1994 & ~n2244 ;
  assign n2246 = \shift_data_reg[81]/NET0131  & n1377 ;
  assign n2247 = ~n2245 & ~n2246 ;
  assign n2248 = \shift_data_reg[82]/NET0131  & n1377 ;
  assign n2249 = \shift_data_reg[82]/NET0131  & ~\wb_sel_i[2]_pad  ;
  assign n2250 = \wb_dat_i[18]_pad  & \wb_sel_i[2]_pad  ;
  assign n2251 = ~n2249 & ~n2250 ;
  assign n2252 = n1483 & ~n2251 ;
  assign n2253 = n2001 & n2059 ;
  assign n2254 = n1892 & n2253 ;
  assign n2255 = ~\shift_data_reg[82]/NET0131  & ~n2253 ;
  assign n2256 = n2006 & ~n2255 ;
  assign n2257 = ~n2254 & n2256 ;
  assign n2258 = ~n2252 & ~n2257 ;
  assign n2259 = ~n1994 & ~n2258 ;
  assign n2260 = ~n2248 & ~n2259 ;
  assign n2261 = \shift_data_reg[80]/NET0131  & ~\wb_sel_i[2]_pad  ;
  assign n2262 = \wb_dat_i[16]_pad  & \wb_sel_i[2]_pad  ;
  assign n2263 = ~n2261 & ~n2262 ;
  assign n2264 = n1483 & ~n2263 ;
  assign n2265 = n1442 & n2001 ;
  assign n2266 = n1950 & n2265 ;
  assign n2267 = n1892 & n2266 ;
  assign n2268 = ~\shift_data_reg[80]/NET0131  & ~n2266 ;
  assign n2269 = n2006 & ~n2268 ;
  assign n2270 = ~n2267 & n2269 ;
  assign n2271 = ~n2264 & ~n2270 ;
  assign n2272 = ~n1994 & ~n2271 ;
  assign n2273 = \shift_data_reg[80]/NET0131  & n1377 ;
  assign n2274 = ~n2272 & ~n2273 ;
  assign n2275 = \shift_data_reg[83]/NET0131  & ~\wb_sel_i[2]_pad  ;
  assign n2276 = \wb_dat_i[19]_pad  & \wb_sel_i[2]_pad  ;
  assign n2277 = ~n2275 & ~n2276 ;
  assign n2278 = n1483 & ~n2277 ;
  assign n2279 = n2072 & n2265 ;
  assign n2280 = n1892 & n2279 ;
  assign n2281 = ~\shift_data_reg[83]/NET0131  & ~n2279 ;
  assign n2282 = n2006 & ~n2281 ;
  assign n2283 = ~n2280 & n2282 ;
  assign n2284 = ~n2278 & ~n2283 ;
  assign n2285 = ~n1994 & ~n2284 ;
  assign n2286 = \shift_data_reg[83]/NET0131  & n1377 ;
  assign n2287 = ~n2285 & ~n2286 ;
  assign n2288 = \shift_data_reg[84]/NET0131  & ~\wb_sel_i[2]_pad  ;
  assign n2289 = \wb_dat_i[20]_pad  & \wb_sel_i[2]_pad  ;
  assign n2290 = ~n2288 & ~n2289 ;
  assign n2291 = n1483 & ~n2290 ;
  assign n2292 = n2001 & n2086 ;
  assign n2293 = n1892 & n2292 ;
  assign n2294 = ~\shift_data_reg[84]/NET0131  & ~n2292 ;
  assign n2295 = n2006 & ~n2294 ;
  assign n2296 = ~n2293 & n2295 ;
  assign n2297 = ~n2291 & ~n2296 ;
  assign n2298 = ~n1994 & ~n2297 ;
  assign n2299 = \shift_data_reg[84]/NET0131  & n1377 ;
  assign n2300 = ~n2298 & ~n2299 ;
  assign n2301 = \shift_data_reg[85]/NET0131  & ~\wb_sel_i[2]_pad  ;
  assign n2302 = \wb_dat_i[21]_pad  & \wb_sel_i[2]_pad  ;
  assign n2303 = ~n2301 & ~n2302 ;
  assign n2304 = n1483 & ~n2303 ;
  assign n2305 = n1901 & n2265 ;
  assign n2306 = n1892 & n2305 ;
  assign n2307 = ~\shift_data_reg[85]/NET0131  & ~n2305 ;
  assign n2308 = n2006 & ~n2307 ;
  assign n2309 = ~n2306 & n2308 ;
  assign n2310 = ~n2304 & ~n2309 ;
  assign n2311 = ~n1994 & ~n2310 ;
  assign n2312 = \shift_data_reg[85]/NET0131  & n1377 ;
  assign n2313 = ~n2311 & ~n2312 ;
  assign n2314 = \shift_data_reg[86]/NET0131  & ~\wb_sel_i[2]_pad  ;
  assign n2315 = \wb_dat_i[22]_pad  & \wb_sel_i[2]_pad  ;
  assign n2316 = ~n2314 & ~n2315 ;
  assign n2317 = n1483 & ~n2316 ;
  assign n2318 = n1937 & n2265 ;
  assign n2319 = n1892 & n2318 ;
  assign n2320 = ~\shift_data_reg[86]/NET0131  & ~n2318 ;
  assign n2321 = n2006 & ~n2320 ;
  assign n2322 = ~n2319 & n2321 ;
  assign n2323 = ~n2317 & ~n2322 ;
  assign n2324 = ~n1994 & ~n2323 ;
  assign n2325 = \shift_data_reg[86]/NET0131  & n1377 ;
  assign n2326 = ~n2324 & ~n2325 ;
  assign n2327 = \shift_data_reg[88]/NET0131  & ~\wb_sel_i[3]_pad  ;
  assign n2328 = ~n1983 & ~n2327 ;
  assign n2329 = n1483 & ~n2328 ;
  assign n2330 = n1950 & n2002 ;
  assign n2331 = n1892 & n2330 ;
  assign n2332 = ~\shift_data_reg[88]/NET0131  & ~n2330 ;
  assign n2333 = n2006 & ~n2332 ;
  assign n2334 = ~n2331 & n2333 ;
  assign n2335 = ~n2329 & ~n2334 ;
  assign n2336 = ~n1994 & ~n2335 ;
  assign n2337 = \shift_data_reg[88]/NET0131  & n1377 ;
  assign n2338 = ~n2336 & ~n2337 ;
  assign n2339 = \shift_data_reg[87]/NET0131  & ~\wb_sel_i[2]_pad  ;
  assign n2340 = ~n1379 & ~n2339 ;
  assign n2341 = n1483 & ~n2340 ;
  assign n2342 = n1443 & n2001 ;
  assign n2343 = n1892 & n2342 ;
  assign n2344 = ~\shift_data_reg[87]/NET0131  & ~n2342 ;
  assign n2345 = n2006 & ~n2344 ;
  assign n2346 = ~n2343 & n2345 ;
  assign n2347 = ~n2341 & ~n2346 ;
  assign n2348 = ~n1994 & ~n2347 ;
  assign n2349 = \shift_data_reg[87]/NET0131  & n1377 ;
  assign n2350 = ~n2348 & ~n2349 ;
  assign n2351 = \shift_data_reg[90]/NET0131  & ~\wb_sel_i[3]_pad  ;
  assign n2352 = \wb_dat_i[26]_pad  & \wb_sel_i[3]_pad  ;
  assign n2353 = ~n2351 & ~n2352 ;
  assign n2354 = n1483 & ~n2353 ;
  assign n2355 = n2002 & n2058 ;
  assign n2356 = n1892 & n2355 ;
  assign n2357 = ~\shift_data_reg[90]/NET0131  & ~n2355 ;
  assign n2358 = n2006 & ~n2357 ;
  assign n2359 = ~n2356 & n2358 ;
  assign n2360 = ~n2354 & ~n2359 ;
  assign n2361 = ~n1994 & ~n2360 ;
  assign n2362 = \shift_data_reg[90]/NET0131  & n1377 ;
  assign n2363 = ~n2361 & ~n2362 ;
  assign n2364 = \shift_data_reg[91]/NET0131  & ~\wb_sel_i[3]_pad  ;
  assign n2365 = \wb_dat_i[27]_pad  & \wb_sel_i[3]_pad  ;
  assign n2366 = ~n2364 & ~n2365 ;
  assign n2367 = n1483 & ~n2366 ;
  assign n2368 = n2002 & n2072 ;
  assign n2369 = n1892 & n2368 ;
  assign n2370 = ~\shift_data_reg[91]/NET0131  & ~n2368 ;
  assign n2371 = n2006 & ~n2370 ;
  assign n2372 = ~n2369 & n2371 ;
  assign n2373 = ~n2367 & ~n2372 ;
  assign n2374 = ~n1994 & ~n2373 ;
  assign n2375 = \shift_data_reg[91]/NET0131  & n1377 ;
  assign n2376 = ~n2374 & ~n2375 ;
  assign n2377 = \shift_data_reg[93]/NET0131  & ~\wb_sel_i[3]_pad  ;
  assign n2378 = \wb_dat_i[29]_pad  & \wb_sel_i[3]_pad  ;
  assign n2379 = ~n2377 & ~n2378 ;
  assign n2380 = n1483 & ~n2379 ;
  assign n2381 = n1901 & n2002 ;
  assign n2382 = n1892 & n2381 ;
  assign n2383 = ~\shift_data_reg[93]/NET0131  & ~n2381 ;
  assign n2384 = n2006 & ~n2383 ;
  assign n2385 = ~n2382 & n2384 ;
  assign n2386 = ~n2380 & ~n2385 ;
  assign n2387 = ~n1994 & ~n2386 ;
  assign n2388 = \shift_data_reg[93]/NET0131  & n1377 ;
  assign n2389 = ~n2387 & ~n2388 ;
  assign n2390 = \shift_data_reg[94]/NET0131  & ~\wb_sel_i[3]_pad  ;
  assign n2391 = \wb_dat_i[30]_pad  & \wb_sel_i[3]_pad  ;
  assign n2392 = ~n2390 & ~n2391 ;
  assign n2393 = n1483 & ~n2392 ;
  assign n2394 = n1937 & n2002 ;
  assign n2395 = n1892 & n2394 ;
  assign n2396 = ~\shift_data_reg[94]/NET0131  & ~n2394 ;
  assign n2397 = n2006 & ~n2396 ;
  assign n2398 = ~n2395 & n2397 ;
  assign n2399 = ~n2393 & ~n2398 ;
  assign n2400 = ~n1994 & ~n2399 ;
  assign n2401 = \shift_data_reg[94]/NET0131  & n1377 ;
  assign n2402 = ~n2400 & ~n2401 ;
  assign n2403 = \shift_data_reg[95]/NET0131  & ~\wb_sel_i[3]_pad  ;
  assign n2404 = ~n1969 & ~n2403 ;
  assign n2405 = n1483 & ~n2404 ;
  assign n2406 = n2001 & n2225 ;
  assign n2407 = n1892 & n2406 ;
  assign n2408 = ~\shift_data_reg[95]/NET0131  & ~n2406 ;
  assign n2409 = n2006 & ~n2408 ;
  assign n2410 = ~n2407 & n2409 ;
  assign n2411 = ~n2405 & ~n2410 ;
  assign n2412 = ~n1994 & ~n2411 ;
  assign n2413 = \shift_data_reg[95]/NET0131  & n1377 ;
  assign n2414 = ~n2412 & ~n2413 ;
  assign n2415 = \shift_data_reg[25]/NET0131  & ~\wb_sel_i[3]_pad  ;
  assign n2416 = ~n1996 & ~n2415 ;
  assign n2417 = n1994 & ~n2416 ;
  assign n2418 = n1498 & n2000 ;
  assign n2419 = ~n1378 & n1485 ;
  assign n2420 = n2418 & n2419 ;
  assign n2421 = ~n1442 & n2420 ;
  assign n2422 = n2003 & n2421 ;
  assign n2424 = n1892 & n2422 ;
  assign n2423 = ~\shift_data_reg[25]/NET0131  & ~n2422 ;
  assign n2425 = ~n1994 & ~n2423 ;
  assign n2426 = ~n2424 & n2425 ;
  assign n2427 = ~n2417 & ~n2426 ;
  assign n2428 = \shift_data_reg[27]/NET0131  & ~\wb_sel_i[3]_pad  ;
  assign n2429 = ~n2365 & ~n2428 ;
  assign n2430 = n1994 & ~n2429 ;
  assign n2431 = n2072 & n2421 ;
  assign n2433 = n1892 & n2431 ;
  assign n2432 = ~\shift_data_reg[27]/NET0131  & ~n2431 ;
  assign n2434 = ~n1994 & ~n2432 ;
  assign n2435 = ~n2433 & n2434 ;
  assign n2436 = ~n2430 & ~n2435 ;
  assign n2437 = \shift_data_reg[26]/NET0131  & ~\wb_sel_i[3]_pad  ;
  assign n2438 = ~n2352 & ~n2437 ;
  assign n2439 = n1994 & ~n2438 ;
  assign n2440 = n2150 & n2420 ;
  assign n2442 = n1892 & n2440 ;
  assign n2441 = ~\shift_data_reg[26]/NET0131  & ~n2440 ;
  assign n2443 = ~n1994 & ~n2441 ;
  assign n2444 = ~n2442 & n2443 ;
  assign n2445 = ~n2439 & ~n2444 ;
  assign n2446 = \shift_data_reg[28]/NET0131  & ~\wb_sel_i[3]_pad  ;
  assign n2447 = ~n2014 & ~n2446 ;
  assign n2448 = n1994 & ~n2447 ;
  assign n2449 = n2017 & n2421 ;
  assign n2451 = n1892 & n2449 ;
  assign n2450 = ~\shift_data_reg[28]/NET0131  & ~n2449 ;
  assign n2452 = ~n1994 & ~n2450 ;
  assign n2453 = ~n2451 & n2452 ;
  assign n2454 = ~n2448 & ~n2453 ;
  assign n2455 = \shift_data_reg[29]/NET0131  & ~\wb_sel_i[3]_pad  ;
  assign n2456 = ~n2378 & ~n2455 ;
  assign n2457 = n1994 & ~n2456 ;
  assign n2458 = n1901 & n2421 ;
  assign n2460 = n1892 & n2458 ;
  assign n2459 = ~\shift_data_reg[29]/NET0131  & ~n2458 ;
  assign n2461 = ~n1994 & ~n2459 ;
  assign n2462 = ~n2460 & n2461 ;
  assign n2463 = ~n2457 & ~n2462 ;
  assign n2464 = \shift_data_reg[2]/NET0131  & ~\wb_sel_i[0]_pad  ;
  assign n2465 = ~n1163 & ~n2464 ;
  assign n2466 = n1994 & ~n2465 ;
  assign n2467 = \shift_data_reg[2]/NET0131  & ~n1994 ;
  assign n2468 = ~n1921 & ~n2467 ;
  assign n2469 = n1498 & n2123 ;
  assign n2470 = n2058 & n2469 ;
  assign n2471 = ~n1892 & n2470 ;
  assign n2472 = \shift_data_reg[2]/NET0131  & ~n2470 ;
  assign n2473 = n2419 & ~n2472 ;
  assign n2474 = ~n2471 & n2473 ;
  assign n2475 = ~n2468 & ~n2474 ;
  assign n2476 = ~n2466 & ~n2475 ;
  assign n2477 = \shift_data_reg[30]/NET0131  & ~\wb_sel_i[3]_pad  ;
  assign n2478 = ~n2391 & ~n2477 ;
  assign n2479 = n1994 & ~n2478 ;
  assign n2480 = n1937 & n2421 ;
  assign n2482 = n1892 & n2480 ;
  assign n2481 = ~\shift_data_reg[30]/NET0131  & ~n2480 ;
  assign n2483 = ~n1994 & ~n2481 ;
  assign n2484 = ~n2482 & n2483 ;
  assign n2485 = ~n2479 & ~n2484 ;
  assign n2486 = \shift_data_reg[31]/NET0131  & ~\wb_sel_i[3]_pad  ;
  assign n2487 = ~n1969 & ~n2486 ;
  assign n2488 = n1994 & ~n2487 ;
  assign n2489 = n1425 & n2421 ;
  assign n2491 = n1892 & n2489 ;
  assign n2490 = ~\shift_data_reg[31]/NET0131  & ~n2489 ;
  assign n2492 = ~n1994 & ~n2490 ;
  assign n2493 = ~n2491 & n2492 ;
  assign n2494 = ~n2488 & ~n2493 ;
  assign n2495 = \shift_data_reg[3]/NET0131  & ~\wb_sel_i[0]_pad  ;
  assign n2496 = ~n1199 & ~n2495 ;
  assign n2497 = n1994 & ~n2496 ;
  assign n2498 = n1498 & n2419 ;
  assign n2499 = n2072 & n2498 ;
  assign n2500 = n2123 & n2499 ;
  assign n2502 = n1892 & n2500 ;
  assign n2501 = ~\shift_data_reg[3]/NET0131  & ~n2500 ;
  assign n2503 = ~n1994 & ~n2501 ;
  assign n2504 = ~n2502 & n2503 ;
  assign n2505 = ~n2497 & ~n2504 ;
  assign n2506 = \shift_data_reg[4]/NET0131  & ~\wb_sel_i[0]_pad  ;
  assign n2507 = ~n1133 & ~n2506 ;
  assign n2508 = n1994 & ~n2507 ;
  assign n2509 = \shift_data_reg[4]/NET0131  & ~n1994 ;
  assign n2510 = ~n1921 & ~n2509 ;
  assign n2511 = n2017 & n2469 ;
  assign n2512 = ~n1892 & n2511 ;
  assign n2513 = \shift_data_reg[4]/NET0131  & ~n2511 ;
  assign n2514 = n2419 & ~n2513 ;
  assign n2515 = ~n2512 & n2514 ;
  assign n2516 = ~n2510 & ~n2515 ;
  assign n2517 = ~n2508 & ~n2516 ;
  assign n2518 = \shift_data_reg[5]/NET0131  & ~\wb_sel_i[0]_pad  ;
  assign n2519 = ~n1156 & ~n2518 ;
  assign n2520 = n1994 & ~n2519 ;
  assign n2521 = n1901 & n2419 ;
  assign n2522 = n2469 & n2521 ;
  assign n2524 = n1892 & n2522 ;
  assign n2523 = ~\shift_data_reg[5]/NET0131  & ~n2522 ;
  assign n2525 = ~n1994 & ~n2523 ;
  assign n2526 = ~n2524 & n2525 ;
  assign n2527 = ~n2520 & ~n2526 ;
  assign n2528 = \shift_data_reg[6]/NET0131  & ~\wb_sel_i[0]_pad  ;
  assign n2529 = ~n1179 & ~n2528 ;
  assign n2530 = n1994 & ~n2529 ;
  assign n2531 = n1937 & n2419 ;
  assign n2532 = n2469 & n2531 ;
  assign n2534 = n1892 & n2532 ;
  assign n2533 = ~\shift_data_reg[6]/NET0131  & ~n2532 ;
  assign n2535 = ~n1994 & ~n2533 ;
  assign n2536 = ~n2534 & n2535 ;
  assign n2537 = ~n2530 & ~n2536 ;
  assign n2538 = \shift_data_reg[0]/NET0131  & ~\wb_sel_i[0]_pad  ;
  assign n2539 = ~n1220 & ~n2538 ;
  assign n2540 = n1994 & ~n2539 ;
  assign n2541 = \shift_data_reg[0]/NET0131  & ~n1994 ;
  assign n2542 = ~n1921 & ~n2541 ;
  assign n2543 = n1950 & n2469 ;
  assign n2544 = ~n1892 & n2543 ;
  assign n2545 = \shift_data_reg[0]/NET0131  & ~n2543 ;
  assign n2546 = n2419 & ~n2545 ;
  assign n2547 = ~n2544 & n2546 ;
  assign n2548 = ~n2542 & ~n2547 ;
  assign n2549 = ~n2540 & ~n2548 ;
  assign n2550 = \shift_data_reg[10]/NET0131  & ~\wb_sel_i[1]_pad  ;
  assign n2551 = ~n1144 & ~n2550 ;
  assign n2552 = n1994 & ~n2551 ;
  assign n2553 = \shift_data_reg[10]/NET0131  & \wb_adr_i[2]_pad  ;
  assign n2554 = n1377 & ~n2553 ;
  assign n2555 = n1498 & n2175 ;
  assign n2556 = n2058 & n2555 ;
  assign n2557 = n1899 & n2556 ;
  assign n2558 = n2419 & n2556 ;
  assign n2559 = \shift_data_reg[10]/NET0131  & ~n2558 ;
  assign n2560 = ~n2557 & ~n2559 ;
  assign n2561 = ~n2554 & ~n2560 ;
  assign n2562 = ~n2552 & ~n2561 ;
  assign n2563 = \shift_data_reg[7]/NET0131  & ~\wb_sel_i[0]_pad  ;
  assign n2564 = ~n1148 & ~n2563 ;
  assign n2565 = n1994 & ~n2564 ;
  assign n2566 = n2124 & n2498 ;
  assign n2568 = n1892 & n2566 ;
  assign n2567 = ~\shift_data_reg[7]/NET0131  & ~n2566 ;
  assign n2569 = ~n1994 & ~n2567 ;
  assign n2570 = ~n2568 & n2569 ;
  assign n2571 = ~n2565 & ~n2570 ;
  assign n2572 = \shift_data_reg[11]/NET0131  & ~\wb_sel_i[1]_pad  ;
  assign n2573 = ~n1171 & ~n2572 ;
  assign n2574 = n1994 & ~n2573 ;
  assign n2575 = n2175 & n2499 ;
  assign n2577 = n1892 & n2575 ;
  assign n2576 = ~\shift_data_reg[11]/NET0131  & ~n2575 ;
  assign n2578 = ~n1994 & ~n2576 ;
  assign n2579 = ~n2577 & n2578 ;
  assign n2580 = ~n2574 & ~n2579 ;
  assign n2581 = \shift_data_reg[8]/NET0131  & ~\wb_sel_i[1]_pad  ;
  assign n2582 = ~n809 & ~n2581 ;
  assign n2583 = n1994 & ~n2582 ;
  assign n2584 = \shift_data_reg[8]/NET0131  & ~n1994 ;
  assign n2585 = ~n1921 & ~n2584 ;
  assign n2586 = n1950 & n2555 ;
  assign n2587 = ~n1892 & n2586 ;
  assign n2588 = \shift_data_reg[8]/NET0131  & ~n2586 ;
  assign n2589 = n2419 & ~n2588 ;
  assign n2590 = ~n2587 & n2589 ;
  assign n2591 = ~n2585 & ~n2590 ;
  assign n2592 = ~n2583 & ~n2591 ;
  assign n2593 = \shift_data_reg[9]/NET0131  & ~\wb_sel_i[1]_pad  ;
  assign n2594 = ~n1216 & ~n2593 ;
  assign n2595 = n1994 & ~n2594 ;
  assign n2596 = n2176 & n2498 ;
  assign n2598 = n1892 & n2596 ;
  assign n2597 = ~\shift_data_reg[9]/NET0131  & ~n2596 ;
  assign n2599 = ~n1994 & ~n2597 ;
  assign n2600 = ~n2598 & n2599 ;
  assign n2601 = ~n2595 & ~n2600 ;
  assign n2602 = \shift_data_reg[12]/NET0131  & ~\wb_sel_i[1]_pad  ;
  assign n2603 = ~n1209 & ~n2602 ;
  assign n2604 = n1994 & ~n2603 ;
  assign n2605 = \shift_data_reg[12]/NET0131  & \wb_adr_i[2]_pad  ;
  assign n2606 = n1377 & ~n2605 ;
  assign n2607 = n2017 & n2555 ;
  assign n2608 = n2419 & n2607 ;
  assign n2609 = \shift_data_reg[12]/NET0131  & ~n2608 ;
  assign n2610 = n1899 & n2607 ;
  assign n2611 = ~n2609 & ~n2610 ;
  assign n2612 = ~n2606 & ~n2611 ;
  assign n2613 = ~n2604 & ~n2612 ;
  assign n2614 = \shift_data_reg[14]/NET0131  & ~\wb_sel_i[1]_pad  ;
  assign n2615 = ~n1175 & ~n2614 ;
  assign n2616 = n1994 & ~n2615 ;
  assign n2617 = n2531 & n2555 ;
  assign n2619 = n1892 & n2617 ;
  assign n2618 = ~\shift_data_reg[14]/NET0131  & ~n2617 ;
  assign n2620 = ~n1994 & ~n2618 ;
  assign n2621 = ~n2619 & n2620 ;
  assign n2622 = ~n2616 & ~n2621 ;
  assign n2623 = \shift_data_reg[13]/NET0131  & ~\wb_sel_i[1]_pad  ;
  assign n2624 = ~n1152 & ~n2623 ;
  assign n2625 = n1994 & ~n2624 ;
  assign n2626 = n2521 & n2555 ;
  assign n2628 = n1892 & n2626 ;
  assign n2627 = ~\shift_data_reg[13]/NET0131  & ~n2626 ;
  assign n2629 = ~n1994 & ~n2627 ;
  assign n2630 = ~n2628 & n2629 ;
  assign n2631 = ~n2625 & ~n2630 ;
  assign n2632 = \shift_data_reg[15]/NET0131  & ~\wb_sel_i[1]_pad  ;
  assign n2633 = ~n1230 & ~n2632 ;
  assign n2634 = n1994 & ~n2633 ;
  assign n2635 = \shift_data_reg[15]/NET0131  & ~n1994 ;
  assign n2636 = ~n1921 & ~n2635 ;
  assign n2637 = n1425 & n2555 ;
  assign n2638 = ~n1892 & n2637 ;
  assign n2639 = \shift_data_reg[15]/NET0131  & ~n2637 ;
  assign n2640 = n2419 & ~n2639 ;
  assign n2641 = ~n2638 & n2640 ;
  assign n2642 = ~n2636 & ~n2641 ;
  assign n2643 = ~n2634 & ~n2642 ;
  assign n2644 = \shift_data_reg[16]/NET0131  & ~\wb_sel_i[2]_pad  ;
  assign n2645 = ~n2262 & ~n2644 ;
  assign n2646 = n1994 & ~n2645 ;
  assign n2647 = \shift_data_reg[16]/NET0131  & ~n1994 ;
  assign n2648 = ~n1921 & ~n2647 ;
  assign n2649 = n2030 & n2418 ;
  assign n2650 = ~n1892 & n2649 ;
  assign n2651 = \shift_data_reg[16]/NET0131  & ~n2649 ;
  assign n2652 = n2419 & ~n2651 ;
  assign n2653 = ~n2650 & n2652 ;
  assign n2654 = ~n2648 & ~n2653 ;
  assign n2655 = ~n2646 & ~n2654 ;
  assign n2656 = \shift_data_reg[17]/NET0131  & ~\wb_sel_i[2]_pad  ;
  assign n2657 = ~n2236 & ~n2656 ;
  assign n2658 = n1994 & ~n2657 ;
  assign n2659 = n1442 & n2420 ;
  assign n2660 = n2003 & n2659 ;
  assign n2662 = n1892 & n2660 ;
  assign n2661 = ~\shift_data_reg[17]/NET0131  & ~n2660 ;
  assign n2663 = ~n1994 & ~n2661 ;
  assign n2664 = ~n2662 & n2663 ;
  assign n2665 = ~n2658 & ~n2664 ;
  assign n2666 = \shift_data_reg[18]/NET0131  & ~\wb_sel_i[2]_pad  ;
  assign n2667 = ~n2250 & ~n2666 ;
  assign n2668 = n1994 & ~n2667 ;
  assign n2669 = n2059 & n2420 ;
  assign n2671 = n1892 & n2669 ;
  assign n2670 = ~\shift_data_reg[18]/NET0131  & ~n2669 ;
  assign n2672 = ~n1994 & ~n2670 ;
  assign n2673 = ~n2671 & n2672 ;
  assign n2674 = ~n2668 & ~n2673 ;
  assign n2675 = \shift_data_reg[19]/NET0131  & ~\wb_sel_i[2]_pad  ;
  assign n2676 = ~n2276 & ~n2675 ;
  assign n2677 = n1994 & ~n2676 ;
  assign n2678 = n2072 & n2659 ;
  assign n2680 = n1892 & n2678 ;
  assign n2679 = ~\shift_data_reg[19]/NET0131  & ~n2678 ;
  assign n2681 = ~n1994 & ~n2679 ;
  assign n2682 = ~n2680 & n2681 ;
  assign n2683 = ~n2677 & ~n2682 ;
  assign n2684 = \shift_data_reg[1]/NET0131  & ~\wb_sel_i[0]_pad  ;
  assign n2685 = ~n1189 & ~n2684 ;
  assign n2686 = n1994 & ~n2685 ;
  assign n2687 = \shift_data_reg[1]/NET0131  & ~n1994 ;
  assign n2688 = ~n1921 & ~n2687 ;
  assign n2689 = n2003 & n2469 ;
  assign n2690 = ~n1892 & n2689 ;
  assign n2691 = \shift_data_reg[1]/NET0131  & ~n2689 ;
  assign n2692 = n2419 & ~n2691 ;
  assign n2693 = ~n2690 & n2692 ;
  assign n2694 = ~n2688 & ~n2693 ;
  assign n2695 = ~n2686 & ~n2694 ;
  assign n2696 = \shift_data_reg[20]/NET0131  & ~\wb_sel_i[2]_pad  ;
  assign n2697 = ~n2289 & ~n2696 ;
  assign n2698 = n1994 & ~n2697 ;
  assign n2699 = n2017 & n2659 ;
  assign n2701 = n1892 & n2699 ;
  assign n2700 = ~\shift_data_reg[20]/NET0131  & ~n2699 ;
  assign n2702 = ~n1994 & ~n2700 ;
  assign n2703 = ~n2701 & n2702 ;
  assign n2704 = ~n2698 & ~n2703 ;
  assign n2705 = \shift_data_reg[21]/NET0131  & ~\wb_sel_i[2]_pad  ;
  assign n2706 = ~n2302 & ~n2705 ;
  assign n2707 = n1994 & ~n2706 ;
  assign n2708 = n1901 & n2659 ;
  assign n2710 = n1892 & n2708 ;
  assign n2709 = ~\shift_data_reg[21]/NET0131  & ~n2708 ;
  assign n2711 = ~n1994 & ~n2709 ;
  assign n2712 = ~n2710 & n2711 ;
  assign n2713 = ~n2707 & ~n2712 ;
  assign n2714 = \shift_data_reg[22]/NET0131  & ~\wb_sel_i[2]_pad  ;
  assign n2715 = ~n2315 & ~n2714 ;
  assign n2716 = n1994 & ~n2715 ;
  assign n2717 = n1937 & n2659 ;
  assign n2719 = n1892 & n2717 ;
  assign n2718 = ~\shift_data_reg[22]/NET0131  & ~n2717 ;
  assign n2720 = ~n1994 & ~n2718 ;
  assign n2721 = ~n2719 & n2720 ;
  assign n2722 = ~n2716 & ~n2721 ;
  assign n2723 = \shift_data_reg[23]/NET0131  & ~\wb_sel_i[2]_pad  ;
  assign n2724 = ~n1379 & ~n2723 ;
  assign n2725 = n1994 & ~n2724 ;
  assign n2726 = \shift_data_reg[23]/NET0131  & ~n1994 ;
  assign n2727 = ~n1921 & ~n2726 ;
  assign n2728 = n1443 & n2418 ;
  assign n2729 = ~n1892 & n2728 ;
  assign n2730 = \shift_data_reg[23]/NET0131  & ~n2728 ;
  assign n2731 = n2419 & ~n2730 ;
  assign n2732 = ~n2729 & n2731 ;
  assign n2733 = ~n2727 & ~n2732 ;
  assign n2734 = ~n2725 & ~n2733 ;
  assign n2735 = \shift_data_reg[24]/NET0131  & ~\wb_sel_i[3]_pad  ;
  assign n2736 = ~n1983 & ~n2735 ;
  assign n2737 = n1994 & ~n2736 ;
  assign n2738 = ~n1442 & n1950 ;
  assign n2739 = n2420 & n2738 ;
  assign n2741 = n1892 & n2739 ;
  assign n2740 = ~\shift_data_reg[24]/NET0131  & ~n2739 ;
  assign n2742 = ~n1994 & ~n2740 ;
  assign n2743 = ~n2741 & n2742 ;
  assign n2744 = ~n2737 & ~n2743 ;
  assign n2747 = n1952 & n2003 ;
  assign n2749 = n1892 & n2747 ;
  assign n2748 = ~\shift_data_reg[33]/NET0131  & ~n2747 ;
  assign n2750 = ~n1377 & ~n2748 ;
  assign n2751 = ~n2749 & n2750 ;
  assign n2745 = n1189 & n1378 ;
  assign n2746 = \shift_data_reg[33]/NET0131  & n1947 ;
  assign n2752 = ~n2745 & ~n2746 ;
  assign n2753 = ~n2751 & n2752 ;
  assign n2756 = n1952 & n2058 ;
  assign n2758 = n1892 & n2756 ;
  assign n2757 = ~\shift_data_reg[34]/NET0131  & ~n2756 ;
  assign n2759 = ~n1377 & ~n2757 ;
  assign n2760 = ~n2758 & n2759 ;
  assign n2754 = n1163 & n1378 ;
  assign n2755 = \shift_data_reg[34]/NET0131  & n1947 ;
  assign n2761 = ~n2754 & ~n2755 ;
  assign n2762 = ~n2760 & n2761 ;
  assign n2765 = n1952 & n2072 ;
  assign n2767 = n1892 & n2765 ;
  assign n2766 = ~\shift_data_reg[35]/NET0131  & ~n2765 ;
  assign n2768 = ~n1377 & ~n2766 ;
  assign n2769 = ~n2767 & n2768 ;
  assign n2763 = n1199 & n1378 ;
  assign n2764 = \shift_data_reg[35]/NET0131  & n1947 ;
  assign n2770 = ~n2763 & ~n2764 ;
  assign n2771 = ~n2769 & n2770 ;
  assign n2774 = n1952 & n2017 ;
  assign n2776 = n1892 & n2774 ;
  assign n2775 = ~\shift_data_reg[36]/NET0131  & ~n2774 ;
  assign n2777 = ~n1377 & ~n2775 ;
  assign n2778 = ~n2776 & n2777 ;
  assign n2772 = n1133 & n1378 ;
  assign n2773 = \shift_data_reg[36]/NET0131  & n1947 ;
  assign n2779 = ~n2772 & ~n2773 ;
  assign n2780 = ~n2778 & n2779 ;
  assign n2783 = n1901 & n1952 ;
  assign n2785 = n1892 & n2783 ;
  assign n2784 = ~\shift_data_reg[37]/NET0131  & ~n2783 ;
  assign n2786 = ~n1377 & ~n2784 ;
  assign n2787 = ~n2785 & n2786 ;
  assign n2781 = n1156 & n1378 ;
  assign n2782 = \shift_data_reg[37]/NET0131  & n1947 ;
  assign n2788 = ~n2781 & ~n2782 ;
  assign n2789 = ~n2787 & n2788 ;
  assign n2792 = n1937 & n1952 ;
  assign n2794 = n1892 & n2792 ;
  assign n2793 = ~\shift_data_reg[38]/NET0131  & ~n2792 ;
  assign n2795 = ~n1377 & ~n2793 ;
  assign n2796 = ~n2794 & n2795 ;
  assign n2790 = n1179 & n1378 ;
  assign n2791 = \shift_data_reg[38]/NET0131  & n1947 ;
  assign n2797 = ~n2790 & ~n2791 ;
  assign n2798 = ~n2796 & n2797 ;
  assign n2803 = n1902 & n1974 ;
  assign n2804 = n1950 & n2803 ;
  assign n2806 = n1892 & n2804 ;
  assign n2805 = ~\shift_data_reg[40]/NET0131  & ~n2804 ;
  assign n2807 = ~n1377 & ~n2805 ;
  assign n2808 = ~n2806 & n2807 ;
  assign n2799 = n809 & n1378 ;
  assign n2800 = \wb_adr_i[2]_pad  & \wb_sel_i[1]_pad  ;
  assign n2801 = n1377 & ~n2800 ;
  assign n2802 = \shift_data_reg[40]/NET0131  & n2801 ;
  assign n2809 = ~n2799 & ~n2802 ;
  assign n2810 = ~n2808 & n2809 ;
  assign n2813 = n2003 & n2803 ;
  assign n2815 = n1892 & n2813 ;
  assign n2814 = ~\shift_data_reg[41]/NET0131  & ~n2813 ;
  assign n2816 = ~n1377 & ~n2814 ;
  assign n2817 = ~n2815 & n2816 ;
  assign n2811 = n1216 & n1378 ;
  assign n2812 = \shift_data_reg[41]/NET0131  & n2801 ;
  assign n2818 = ~n2811 & ~n2812 ;
  assign n2819 = ~n2817 & n2818 ;
  assign n2822 = n2058 & n2803 ;
  assign n2824 = n1892 & n2822 ;
  assign n2823 = ~\shift_data_reg[42]/NET0131  & ~n2822 ;
  assign n2825 = ~n1377 & ~n2823 ;
  assign n2826 = ~n2824 & n2825 ;
  assign n2820 = n1144 & n1378 ;
  assign n2821 = \shift_data_reg[42]/NET0131  & n2801 ;
  assign n2827 = ~n2820 & ~n2821 ;
  assign n2828 = ~n2826 & n2827 ;
  assign n2831 = n2072 & n2803 ;
  assign n2833 = n1892 & n2831 ;
  assign n2832 = ~\shift_data_reg[43]/NET0131  & ~n2831 ;
  assign n2834 = ~n1377 & ~n2832 ;
  assign n2835 = ~n2833 & n2834 ;
  assign n2829 = n1171 & n1378 ;
  assign n2830 = \shift_data_reg[43]/NET0131  & n2801 ;
  assign n2836 = ~n2829 & ~n2830 ;
  assign n2837 = ~n2835 & n2836 ;
  assign n2840 = n2017 & n2803 ;
  assign n2842 = n1892 & n2840 ;
  assign n2841 = ~\shift_data_reg[44]/NET0131  & ~n2840 ;
  assign n2843 = ~n1377 & ~n2841 ;
  assign n2844 = ~n2842 & n2843 ;
  assign n2838 = n1209 & n1378 ;
  assign n2839 = \shift_data_reg[44]/NET0131  & n2801 ;
  assign n2845 = ~n2838 & ~n2839 ;
  assign n2846 = ~n2844 & n2845 ;
  assign n2849 = n1901 & n2803 ;
  assign n2851 = n1892 & n2849 ;
  assign n2850 = ~\shift_data_reg[45]/NET0131  & ~n2849 ;
  assign n2852 = ~n1377 & ~n2850 ;
  assign n2853 = ~n2851 & n2852 ;
  assign n2847 = n1152 & n1378 ;
  assign n2848 = \shift_data_reg[45]/NET0131  & n2801 ;
  assign n2854 = ~n2847 & ~n2848 ;
  assign n2855 = ~n2853 & n2854 ;
  assign n2858 = n1937 & n2803 ;
  assign n2860 = n1892 & n2858 ;
  assign n2859 = ~\shift_data_reg[46]/NET0131  & ~n2858 ;
  assign n2861 = ~n1377 & ~n2859 ;
  assign n2862 = ~n2860 & n2861 ;
  assign n2856 = n1175 & n1378 ;
  assign n2857 = \shift_data_reg[46]/NET0131  & n2801 ;
  assign n2863 = ~n2856 & ~n2857 ;
  assign n2864 = ~n2862 & n2863 ;
  assign n2867 = n1425 & n2803 ;
  assign n2869 = n1892 & n2867 ;
  assign n2868 = ~\shift_data_reg[47]/NET0131  & ~n2867 ;
  assign n2870 = ~n1377 & ~n2868 ;
  assign n2871 = ~n2869 & n2870 ;
  assign n2865 = n1230 & n1378 ;
  assign n2866 = \shift_data_reg[47]/NET0131  & n2801 ;
  assign n2872 = ~n2865 & ~n2866 ;
  assign n2873 = ~n2871 & n2872 ;
  assign n2876 = n1500 & n2030 ;
  assign n2878 = n1892 & n2876 ;
  assign n2877 = ~\shift_data_reg[48]/NET0131  & ~n2876 ;
  assign n2879 = ~n1377 & ~n2877 ;
  assign n2880 = ~n2878 & n2879 ;
  assign n2874 = n1378 & n2262 ;
  assign n2875 = \shift_data_reg[48]/NET0131  & n1382 ;
  assign n2881 = ~n2874 & ~n2875 ;
  assign n2882 = ~n2880 & n2881 ;
  assign n2885 = n1500 & n2045 ;
  assign n2887 = n1892 & n2885 ;
  assign n2886 = ~\shift_data_reg[49]/NET0131  & ~n2885 ;
  assign n2888 = ~n1377 & ~n2886 ;
  assign n2889 = ~n2887 & n2888 ;
  assign n2883 = n1378 & n2236 ;
  assign n2884 = \shift_data_reg[49]/NET0131  & n1382 ;
  assign n2890 = ~n2883 & ~n2884 ;
  assign n2891 = ~n2889 & n2890 ;
  assign n2894 = n1500 & n2059 ;
  assign n2896 = n1892 & n2894 ;
  assign n2895 = ~\shift_data_reg[50]/NET0131  & ~n2894 ;
  assign n2897 = ~n1377 & ~n2895 ;
  assign n2898 = ~n2896 & n2897 ;
  assign n2892 = n1378 & n2250 ;
  assign n2893 = \shift_data_reg[50]/NET0131  & n1382 ;
  assign n2899 = ~n2892 & ~n2893 ;
  assign n2900 = ~n2898 & n2899 ;
  assign n2903 = n1480 & n2072 ;
  assign n2904 = n1951 & n2903 ;
  assign n2906 = n1892 & n2904 ;
  assign n2905 = ~\shift_data_reg[51]/NET0131  & ~n2904 ;
  assign n2907 = ~n1377 & ~n2905 ;
  assign n2908 = ~n2906 & n2907 ;
  assign n2901 = n1378 & n2276 ;
  assign n2902 = \shift_data_reg[51]/NET0131  & n1382 ;
  assign n2909 = ~n2901 & ~n2902 ;
  assign n2910 = ~n2908 & n2909 ;
  assign n2913 = n1500 & n2086 ;
  assign n2915 = n1892 & n2913 ;
  assign n2914 = ~\shift_data_reg[52]/NET0131  & ~n2913 ;
  assign n2916 = ~n1377 & ~n2914 ;
  assign n2917 = ~n2915 & n2916 ;
  assign n2911 = n1378 & n2289 ;
  assign n2912 = \shift_data_reg[52]/NET0131  & n1382 ;
  assign n2918 = ~n2911 & ~n2912 ;
  assign n2919 = ~n2917 & n2918 ;
  assign n2922 = n1480 & n1901 ;
  assign n2923 = n1951 & n2922 ;
  assign n2925 = n1892 & n2923 ;
  assign n2924 = ~\shift_data_reg[53]/NET0131  & ~n2923 ;
  assign n2926 = ~n1377 & ~n2924 ;
  assign n2927 = ~n2925 & n2926 ;
  assign n2920 = n1378 & n2302 ;
  assign n2921 = \shift_data_reg[53]/NET0131  & n1382 ;
  assign n2928 = ~n2920 & ~n2921 ;
  assign n2929 = ~n2927 & n2928 ;
  assign n2932 = n1480 & n1937 ;
  assign n2933 = n1951 & n2932 ;
  assign n2935 = n1892 & n2933 ;
  assign n2934 = ~\shift_data_reg[54]/NET0131  & ~n2933 ;
  assign n2936 = ~n1377 & ~n2934 ;
  assign n2937 = ~n2935 & n2936 ;
  assign n2930 = n1378 & n2315 ;
  assign n2931 = \shift_data_reg[54]/NET0131  & n1382 ;
  assign n2938 = ~n2930 & ~n2931 ;
  assign n2939 = ~n2937 & n2938 ;
  assign n2942 = n1975 & n2003 ;
  assign n2944 = n1892 & n2942 ;
  assign n2943 = ~\shift_data_reg[57]/NET0131  & ~n2942 ;
  assign n2945 = ~n1377 & ~n2943 ;
  assign n2946 = ~n2944 & n2945 ;
  assign n2940 = n1378 & n1996 ;
  assign n2941 = \shift_data_reg[57]/NET0131  & n1972 ;
  assign n2947 = ~n2940 & ~n2941 ;
  assign n2948 = ~n2946 & n2947 ;
  assign n2951 = n1975 & n2058 ;
  assign n2953 = n1892 & n2951 ;
  assign n2952 = ~\shift_data_reg[58]/NET0131  & ~n2951 ;
  assign n2954 = ~n1377 & ~n2952 ;
  assign n2955 = ~n2953 & n2954 ;
  assign n2949 = n1378 & n2352 ;
  assign n2950 = \shift_data_reg[58]/NET0131  & n1972 ;
  assign n2956 = ~n2949 & ~n2950 ;
  assign n2957 = ~n2955 & n2956 ;
  assign n2960 = n1974 & n2903 ;
  assign n2962 = n1892 & n2960 ;
  assign n2961 = ~\shift_data_reg[59]/NET0131  & ~n2960 ;
  assign n2963 = ~n1377 & ~n2961 ;
  assign n2964 = ~n2962 & n2963 ;
  assign n2958 = n1378 & n2365 ;
  assign n2959 = \shift_data_reg[59]/NET0131  & n1972 ;
  assign n2965 = ~n2958 & ~n2959 ;
  assign n2966 = ~n2964 & n2965 ;
  assign n2969 = n1975 & n2017 ;
  assign n2971 = n1892 & n2969 ;
  assign n2970 = ~\shift_data_reg[60]/NET0131  & ~n2969 ;
  assign n2972 = ~n1377 & ~n2970 ;
  assign n2973 = ~n2971 & n2972 ;
  assign n2967 = n1378 & n2014 ;
  assign n2968 = \shift_data_reg[60]/NET0131  & n1972 ;
  assign n2974 = ~n2967 & ~n2968 ;
  assign n2975 = ~n2973 & n2974 ;
  assign n2978 = n1974 & n2922 ;
  assign n2980 = n1892 & n2978 ;
  assign n2979 = ~\shift_data_reg[61]/NET0131  & ~n2978 ;
  assign n2981 = ~n1377 & ~n2979 ;
  assign n2982 = ~n2980 & n2981 ;
  assign n2976 = n1378 & n2378 ;
  assign n2977 = \shift_data_reg[61]/NET0131  & n1972 ;
  assign n2983 = ~n2976 & ~n2977 ;
  assign n2984 = ~n2982 & n2983 ;
  assign n2987 = n1974 & n2932 ;
  assign n2989 = n1892 & n2987 ;
  assign n2988 = ~\shift_data_reg[62]/NET0131  & ~n2987 ;
  assign n2990 = ~n1377 & ~n2988 ;
  assign n2991 = ~n2989 & n2990 ;
  assign n2985 = n1378 & n2391 ;
  assign n2986 = \shift_data_reg[62]/NET0131  & n1972 ;
  assign n2992 = ~n2985 & ~n2986 ;
  assign n2993 = ~n2991 & n2992 ;
  assign n2994 = \shift_data_reg[105]/NET0131  & ~\wb_sel_i[1]_pad  ;
  assign n2995 = ~n1216 & ~n2994 ;
  assign n2996 = n1484 & ~n2995 ;
  assign n2997 = n1923 & n2003 ;
  assign n2998 = n1892 & n2997 ;
  assign n2999 = ~\shift_data_reg[105]/NET0131  & ~n2997 ;
  assign n3000 = n1485 & ~n2999 ;
  assign n3001 = ~n2998 & n3000 ;
  assign n3002 = ~n2996 & ~n3001 ;
  assign n3003 = ~n1377 & ~n3002 ;
  assign n3004 = \shift_data_reg[105]/NET0131  & ~n1910 ;
  assign n3005 = ~n3003 & ~n3004 ;
  assign n3006 = \shift_data_reg[113]/NET0131  & ~\wb_sel_i[2]_pad  ;
  assign n3007 = ~n2236 & ~n3006 ;
  assign n3008 = n1484 & ~n3007 ;
  assign n3009 = n1480 & ~n1498 ;
  assign n3010 = n2045 & n3009 ;
  assign n3011 = n1892 & n3010 ;
  assign n3012 = ~\shift_data_reg[113]/NET0131  & ~n3010 ;
  assign n3013 = n1485 & ~n3012 ;
  assign n3014 = ~n3011 & n3013 ;
  assign n3015 = ~n3008 & ~n3014 ;
  assign n3016 = ~n1377 & ~n3015 ;
  assign n3017 = \shift_data_reg[113]/NET0131  & ~n1910 ;
  assign n3018 = ~n3016 & ~n3017 ;
  assign n3019 = \shift_data_reg[108]/NET0131  & ~\wb_sel_i[1]_pad  ;
  assign n3020 = ~n1209 & ~n3019 ;
  assign n3021 = n1484 & ~n3020 ;
  assign n3022 = n1923 & n2017 ;
  assign n3023 = n1892 & n3022 ;
  assign n3024 = ~\shift_data_reg[108]/NET0131  & ~n3022 ;
  assign n3025 = n1485 & ~n3024 ;
  assign n3026 = ~n3023 & n3025 ;
  assign n3027 = ~n3021 & ~n3026 ;
  assign n3028 = ~n1377 & ~n3027 ;
  assign n3029 = \shift_data_reg[108]/NET0131  & ~n1910 ;
  assign n3030 = ~n3028 & ~n3029 ;
  assign n3031 = \shift_data_reg[116]/NET0131  & ~\wb_sel_i[2]_pad  ;
  assign n3032 = ~n2289 & ~n3031 ;
  assign n3033 = n1484 & ~n3032 ;
  assign n3034 = n2086 & n3009 ;
  assign n3035 = n1892 & n3034 ;
  assign n3036 = ~\shift_data_reg[116]/NET0131  & ~n3034 ;
  assign n3037 = n1485 & ~n3036 ;
  assign n3038 = ~n3035 & n3037 ;
  assign n3039 = ~n3033 & ~n3038 ;
  assign n3040 = ~n1377 & ~n3039 ;
  assign n3041 = \shift_data_reg[116]/NET0131  & ~n1910 ;
  assign n3042 = ~n3040 & ~n3041 ;
  assign n3043 = n2738 & n3009 ;
  assign n3044 = n1899 & n3043 ;
  assign n3045 = \shift_data_reg[120]/NET0131  & ~\wb_sel_i[3]_pad  ;
  assign n3046 = ~n1983 & ~n3045 ;
  assign n3047 = n1484 & ~n3046 ;
  assign n3048 = \shift_data_reg[120]/NET0131  & n1485 ;
  assign n3049 = ~n3043 & n3048 ;
  assign n3050 = ~n3047 & ~n3049 ;
  assign n3051 = ~n3044 & n3050 ;
  assign n3052 = ~n1377 & ~n3051 ;
  assign n3053 = \shift_data_reg[120]/NET0131  & ~n1910 ;
  assign n3054 = ~n3052 & ~n3053 ;
  assign n3055 = n1179 & n1484 ;
  assign n3056 = n1904 & n1937 ;
  assign n3057 = n1899 & n3056 ;
  assign n3058 = ~n3055 & ~n3057 ;
  assign n3059 = ~n1377 & ~n3058 ;
  assign n3060 = ~n1484 & ~n3056 ;
  assign n3061 = n1912 & ~n3060 ;
  assign n3062 = \shift_data_reg[102]/NET0131  & ~n3061 ;
  assign n3063 = ~n3059 & ~n3062 ;
  assign n3064 = \shift_data_reg[107]/NET0131  & ~\wb_sel_i[1]_pad  ;
  assign n3065 = ~n1171 & ~n3064 ;
  assign n3066 = n1484 & ~n3065 ;
  assign n3067 = n1923 & n2072 ;
  assign n3068 = n1892 & n3067 ;
  assign n3069 = ~\shift_data_reg[107]/NET0131  & ~n3067 ;
  assign n3070 = n1485 & ~n3069 ;
  assign n3071 = ~n3068 & n3070 ;
  assign n3072 = ~n3066 & ~n3071 ;
  assign n3073 = ~n1377 & ~n3072 ;
  assign n3074 = \shift_data_reg[107]/NET0131  & ~n1910 ;
  assign n3075 = ~n3073 & ~n3074 ;
  assign n3076 = \shift_data_reg[115]/NET0131  & ~n1910 ;
  assign n3077 = n1903 & n2903 ;
  assign n3079 = ~n1892 & n3077 ;
  assign n3078 = \shift_data_reg[115]/NET0131  & ~n3077 ;
  assign n3080 = \shift_data_reg[115]/NET0131  & ~\wb_sel_i[2]_pad  ;
  assign n3081 = ~n2276 & ~n3080 ;
  assign n3082 = n1484 & ~n3081 ;
  assign n3083 = ~n3078 & ~n3082 ;
  assign n3084 = ~n3079 & n3083 ;
  assign n3085 = ~n1485 & ~n3082 ;
  assign n3086 = ~n1377 & ~n3085 ;
  assign n3087 = ~n3084 & n3086 ;
  assign n3088 = ~n3076 & ~n3087 ;
  assign n3089 = \shift_data_reg[118]/NET0131  & ~\wb_sel_i[2]_pad  ;
  assign n3090 = ~n2315 & ~n3089 ;
  assign n3091 = n1484 & ~n3090 ;
  assign n3092 = n1903 & n2932 ;
  assign n3093 = n1892 & n3092 ;
  assign n3094 = ~\shift_data_reg[118]/NET0131  & ~n3092 ;
  assign n3095 = n1485 & ~n3094 ;
  assign n3096 = ~n3093 & n3095 ;
  assign n3097 = ~n3091 & ~n3096 ;
  assign n3098 = ~n1377 & ~n3097 ;
  assign n3099 = \shift_data_reg[118]/NET0131  & ~n1910 ;
  assign n3100 = ~n3098 & ~n3099 ;
  assign n3101 = \shift_data_reg[117]/NET0131  & ~\wb_sel_i[2]_pad  ;
  assign n3102 = ~n2302 & ~n3101 ;
  assign n3103 = n1484 & ~n3102 ;
  assign n3104 = n1903 & n2922 ;
  assign n3105 = n1892 & n3104 ;
  assign n3106 = ~\shift_data_reg[117]/NET0131  & ~n3104 ;
  assign n3107 = n1485 & ~n3106 ;
  assign n3108 = ~n3105 & n3107 ;
  assign n3109 = ~n3103 & ~n3108 ;
  assign n3110 = ~n1377 & ~n3109 ;
  assign n3111 = \shift_data_reg[117]/NET0131  & ~n1910 ;
  assign n3112 = ~n3110 & ~n3111 ;
  assign n3113 = \shift_data_reg[122]/NET0131  & ~\wb_sel_i[3]_pad  ;
  assign n3114 = ~n2352 & ~n3113 ;
  assign n3115 = n1484 & ~n3114 ;
  assign n3116 = n2150 & n3009 ;
  assign n3117 = n1892 & n3116 ;
  assign n3118 = ~\shift_data_reg[122]/NET0131  & ~n3116 ;
  assign n3119 = n1485 & ~n3118 ;
  assign n3120 = ~n3117 & n3119 ;
  assign n3121 = ~n3115 & ~n3120 ;
  assign n3122 = ~n1377 & ~n3121 ;
  assign n3123 = \shift_data_reg[122]/NET0131  & ~n1910 ;
  assign n3124 = ~n3122 & ~n3123 ;
  assign n3125 = \shift_data_reg[127]/NET0131  & ~\wb_sel_i[3]_pad  ;
  assign n3126 = ~n1969 & ~n3125 ;
  assign n3127 = n1484 & ~n3126 ;
  assign n3128 = n2225 & n3009 ;
  assign n3129 = n1892 & n3128 ;
  assign n3130 = ~\shift_data_reg[127]/NET0131  & ~n3128 ;
  assign n3131 = n1485 & ~n3130 ;
  assign n3132 = ~n3129 & n3131 ;
  assign n3133 = ~n3127 & ~n3132 ;
  assign n3134 = ~n1377 & ~n3133 ;
  assign n3135 = \shift_data_reg[127]/NET0131  & ~n1910 ;
  assign n3136 = ~n3134 & ~n3135 ;
  assign n3137 = n1133 & n1484 ;
  assign n3138 = n1904 & n2017 ;
  assign n3139 = n1899 & n3138 ;
  assign n3140 = ~n3137 & ~n3139 ;
  assign n3141 = ~n1377 & ~n3140 ;
  assign n3142 = ~n1484 & ~n3138 ;
  assign n3143 = n1912 & ~n3142 ;
  assign n3144 = \shift_data_reg[100]/NET0131  & ~n3143 ;
  assign n3145 = ~n3141 & ~n3144 ;
  assign n3146 = n1148 & n1484 ;
  assign n3147 = n1443 & n1922 ;
  assign n3148 = n1899 & n3147 ;
  assign n3149 = ~n3146 & ~n3148 ;
  assign n3150 = ~n1377 & ~n3149 ;
  assign n3151 = ~n1484 & ~n3147 ;
  assign n3152 = n1912 & ~n3151 ;
  assign n3153 = \shift_data_reg[103]/NET0131  & ~n3152 ;
  assign n3154 = ~n3150 & ~n3153 ;
  assign n3155 = \shift_data_reg[104]/NET0131  & ~\wb_sel_i[1]_pad  ;
  assign n3156 = ~n809 & ~n3155 ;
  assign n3157 = n1484 & ~n3156 ;
  assign n3158 = n1923 & n1950 ;
  assign n3159 = n1892 & n3158 ;
  assign n3160 = ~\shift_data_reg[104]/NET0131  & ~n3158 ;
  assign n3161 = n1485 & ~n3160 ;
  assign n3162 = ~n3159 & n3161 ;
  assign n3163 = ~n3157 & ~n3162 ;
  assign n3164 = ~n1377 & ~n3163 ;
  assign n3165 = \shift_data_reg[104]/NET0131  & ~n1910 ;
  assign n3166 = ~n3164 & ~n3165 ;
  assign n3167 = \shift_data_reg[106]/NET0131  & ~\wb_sel_i[1]_pad  ;
  assign n3168 = ~n1144 & ~n3167 ;
  assign n3169 = n1484 & ~n3168 ;
  assign n3170 = n1922 & n2150 ;
  assign n3171 = n1892 & n3170 ;
  assign n3172 = ~\shift_data_reg[106]/NET0131  & ~n3170 ;
  assign n3173 = n1485 & ~n3172 ;
  assign n3174 = ~n3171 & n3173 ;
  assign n3175 = ~n3169 & ~n3174 ;
  assign n3176 = ~n1377 & ~n3175 ;
  assign n3177 = \shift_data_reg[106]/NET0131  & ~n1910 ;
  assign n3178 = ~n3176 & ~n3177 ;
  assign n3179 = \shift_data_reg[111]/NET0131  & ~\wb_sel_i[1]_pad  ;
  assign n3180 = ~n1230 & ~n3179 ;
  assign n3181 = n1484 & ~n3180 ;
  assign n3182 = n1425 & n1923 ;
  assign n3183 = n1892 & n3182 ;
  assign n3184 = ~\shift_data_reg[111]/NET0131  & ~n3182 ;
  assign n3185 = n1485 & ~n3184 ;
  assign n3186 = ~n3183 & n3185 ;
  assign n3187 = ~n3181 & ~n3186 ;
  assign n3188 = ~n1377 & ~n3187 ;
  assign n3189 = \shift_data_reg[111]/NET0131  & ~n1910 ;
  assign n3190 = ~n3188 & ~n3189 ;
  assign n3191 = \shift_data_reg[112]/NET0131  & ~\wb_sel_i[2]_pad  ;
  assign n3192 = ~n2262 & ~n3191 ;
  assign n3193 = n1484 & ~n3192 ;
  assign n3194 = n2030 & n3009 ;
  assign n3195 = n1892 & n3194 ;
  assign n3196 = ~\shift_data_reg[112]/NET0131  & ~n3194 ;
  assign n3197 = n1485 & ~n3196 ;
  assign n3198 = ~n3195 & n3197 ;
  assign n3199 = ~n3193 & ~n3198 ;
  assign n3200 = ~n1377 & ~n3199 ;
  assign n3201 = \shift_data_reg[112]/NET0131  & ~n1910 ;
  assign n3202 = ~n3200 & ~n3201 ;
  assign n3203 = \shift_data_reg[114]/NET0131  & ~\wb_sel_i[2]_pad  ;
  assign n3204 = ~n2250 & ~n3203 ;
  assign n3205 = n1484 & ~n3204 ;
  assign n3206 = n2059 & n3009 ;
  assign n3207 = n1892 & n3206 ;
  assign n3208 = ~\shift_data_reg[114]/NET0131  & ~n3206 ;
  assign n3209 = n1485 & ~n3208 ;
  assign n3210 = ~n3207 & n3209 ;
  assign n3211 = ~n3205 & ~n3210 ;
  assign n3212 = ~n1377 & ~n3211 ;
  assign n3213 = \shift_data_reg[114]/NET0131  & ~n1910 ;
  assign n3214 = ~n3212 & ~n3213 ;
  assign n3215 = \shift_data_reg[119]/NET0131  & ~\wb_sel_i[2]_pad  ;
  assign n3216 = ~n1379 & ~n3215 ;
  assign n3217 = n1484 & ~n3216 ;
  assign n3218 = n1443 & n3009 ;
  assign n3219 = n1892 & n3218 ;
  assign n3220 = ~\shift_data_reg[119]/NET0131  & ~n3218 ;
  assign n3221 = n1485 & ~n3220 ;
  assign n3222 = ~n3219 & n3221 ;
  assign n3223 = ~n3217 & ~n3222 ;
  assign n3224 = ~n1377 & ~n3223 ;
  assign n3225 = \shift_data_reg[119]/NET0131  & ~n1910 ;
  assign n3226 = ~n3224 & ~n3225 ;
  assign n3227 = \shift_data_reg[121]/NET0131  & ~\wb_sel_i[3]_pad  ;
  assign n3228 = ~n1996 & ~n3227 ;
  assign n3229 = n1484 & ~n3228 ;
  assign n3230 = ~n1442 & n3009 ;
  assign n3231 = n2003 & n3230 ;
  assign n3232 = n1892 & n3231 ;
  assign n3233 = ~\shift_data_reg[121]/NET0131  & ~n3231 ;
  assign n3234 = n1485 & ~n3233 ;
  assign n3235 = ~n3232 & n3234 ;
  assign n3236 = ~n3229 & ~n3235 ;
  assign n3237 = ~n1377 & ~n3236 ;
  assign n3238 = \shift_data_reg[121]/NET0131  & ~n1910 ;
  assign n3239 = ~n3237 & ~n3238 ;
  assign n3240 = n1220 & n1484 ;
  assign n3241 = n1922 & n2030 ;
  assign n3242 = n1899 & n3241 ;
  assign n3243 = ~n3240 & ~n3242 ;
  assign n3244 = ~n1377 & ~n3243 ;
  assign n3245 = ~n1484 & ~n3241 ;
  assign n3246 = n1912 & ~n3245 ;
  assign n3247 = \shift_data_reg[96]/NET0131  & ~n3246 ;
  assign n3248 = ~n3244 & ~n3247 ;
  assign n3249 = n1189 & n1484 ;
  assign n3250 = n1922 & n2045 ;
  assign n3251 = n1899 & n3250 ;
  assign n3252 = ~n3249 & ~n3251 ;
  assign n3253 = ~n1377 & ~n3252 ;
  assign n3254 = ~n1484 & ~n3250 ;
  assign n3255 = n1912 & ~n3254 ;
  assign n3256 = \shift_data_reg[97]/NET0131  & ~n3255 ;
  assign n3257 = ~n3253 & ~n3256 ;
  assign n3258 = n1163 & n1484 ;
  assign n3259 = n1904 & n2058 ;
  assign n3260 = n1899 & n3259 ;
  assign n3261 = ~n3258 & ~n3260 ;
  assign n3262 = ~n1377 & ~n3261 ;
  assign n3263 = ~n1484 & ~n3259 ;
  assign n3264 = n1912 & ~n3263 ;
  assign n3265 = \shift_data_reg[98]/NET0131  & ~n3264 ;
  assign n3266 = ~n3262 & ~n3265 ;
  assign n3267 = n1199 & n1484 ;
  assign n3268 = n1904 & n2072 ;
  assign n3269 = n1899 & n3268 ;
  assign n3270 = ~n3267 & ~n3269 ;
  assign n3271 = ~n1377 & ~n3270 ;
  assign n3272 = ~n1484 & ~n3268 ;
  assign n3273 = n1912 & ~n3272 ;
  assign n3274 = \shift_data_reg[99]/NET0131  & ~n3273 ;
  assign n3275 = ~n3271 & ~n3274 ;
  assign n3276 = \shift_data_reg[123]/NET0131  & ~\wb_sel_i[3]_pad  ;
  assign n3277 = ~n2365 & ~n3276 ;
  assign n3278 = n1484 & ~n3277 ;
  assign n3279 = ~n1442 & ~n1498 ;
  assign n3280 = n2903 & n3279 ;
  assign n3281 = n1892 & n3280 ;
  assign n3282 = ~\shift_data_reg[123]/NET0131  & ~n3280 ;
  assign n3283 = n1485 & ~n3282 ;
  assign n3284 = ~n3281 & n3283 ;
  assign n3285 = ~n3278 & ~n3284 ;
  assign n3286 = ~n1377 & ~n3285 ;
  assign n3287 = \shift_data_reg[123]/NET0131  & ~n1910 ;
  assign n3288 = ~n3286 & ~n3287 ;
  assign n3289 = \shift_data_reg[124]/NET0131  & ~\wb_sel_i[3]_pad  ;
  assign n3290 = ~n2014 & ~n3289 ;
  assign n3291 = n1484 & ~n3290 ;
  assign n3292 = n2017 & n3230 ;
  assign n3293 = n1892 & n3292 ;
  assign n3294 = ~\shift_data_reg[124]/NET0131  & ~n3292 ;
  assign n3295 = n1485 & ~n3294 ;
  assign n3296 = ~n3293 & n3295 ;
  assign n3297 = ~n3291 & ~n3296 ;
  assign n3298 = ~n1377 & ~n3297 ;
  assign n3299 = \shift_data_reg[124]/NET0131  & ~n1910 ;
  assign n3300 = ~n3298 & ~n3299 ;
  assign n3301 = \shift_data_reg[125]/NET0131  & ~\wb_sel_i[3]_pad  ;
  assign n3302 = ~n2378 & ~n3301 ;
  assign n3303 = n1484 & ~n3302 ;
  assign n3304 = n2922 & n3279 ;
  assign n3305 = n1892 & n3304 ;
  assign n3306 = ~\shift_data_reg[125]/NET0131  & ~n3304 ;
  assign n3307 = n1485 & ~n3306 ;
  assign n3308 = ~n3305 & n3307 ;
  assign n3309 = ~n3303 & ~n3308 ;
  assign n3310 = ~n1377 & ~n3309 ;
  assign n3311 = \shift_data_reg[125]/NET0131  & ~n1910 ;
  assign n3312 = ~n3310 & ~n3311 ;
  assign n3313 = \shift_data_reg[126]/NET0131  & ~\wb_sel_i[3]_pad  ;
  assign n3314 = ~n2391 & ~n3313 ;
  assign n3315 = n1484 & ~n3314 ;
  assign n3316 = n1937 & n3230 ;
  assign n3317 = n1892 & n3316 ;
  assign n3318 = ~\shift_data_reg[126]/NET0131  & ~n3316 ;
  assign n3319 = n1485 & ~n3318 ;
  assign n3320 = ~n3317 & n3319 ;
  assign n3321 = ~n3315 & ~n3320 ;
  assign n3322 = ~n1377 & ~n3321 ;
  assign n3323 = \shift_data_reg[126]/NET0131  & ~n1910 ;
  assign n3324 = ~n3322 & ~n3323 ;
  assign n3325 = \ctrl_reg[13]/NET0131  & ~\shift_tip_reg/NET0131  ;
  assign n3326 = \ss_reg[0]/NET0131  & ~n3325 ;
  assign n3327 = \ss_reg[1]/NET0131  & ~n3325 ;
  assign n3328 = \ss_reg[2]/NET0131  & ~n3325 ;
  assign n3329 = \ss_reg[3]/NET0131  & ~n3325 ;
  assign n3330 = \ss_reg[4]/NET0131  & ~n3325 ;
  assign n3331 = \ss_reg[5]/NET0131  & ~n3325 ;
  assign n3332 = \ss_reg[6]/NET0131  & ~n3325 ;
  assign n3333 = \ss_reg[7]/NET0131  & ~n3325 ;
  assign \_al_n1  = ~1'b0 ;
  assign \g10384/_0_  = ~n711 ;
  assign \g10421/_0_  = ~n743 ;
  assign \g10487/_0_  = ~n748 ;
  assign \g10622/_0_  = ~n754 ;
  assign \g10625/_0_  = ~n760 ;
  assign \g10631/_3_  = ~n765 ;
  assign \g10641/_0_  = n778 ;
  assign \g10677/_3_  = ~n784 ;
  assign \g10695/_0_  = ~n790 ;
  assign \g10699/_3_  = ~n795 ;
  assign \g10796/_0_  = ~n801 ;
  assign \g10814/_00_  = ~n807 ;
  assign \g10815/_0_  = ~n821 ;
  assign \g10819/_0_  = ~n826 ;
  assign \g10821/_0_  = ~n831 ;
  assign \g10824/_3_  = ~n836 ;
  assign \g10858/_0_  = ~n842 ;
  assign \g11042/_00_  = n848 ;
  assign \g11067/_0_  = n870 ;
  assign \g11071/_00_  = n876 ;
  assign \g11074/_0_  = ~n878 ;
  assign \g11075/_0_  = ~n882 ;
  assign \g11076/_0_  = ~n885 ;
  assign \g11077/_0_  = ~n890 ;
  assign \g11078/_0_  = ~n895 ;
  assign \g11079/_0_  = ~n898 ;
  assign \g11080/_0_  = ~n903 ;
  assign \g11149/_0_  = ~n908 ;
  assign \g11151/_0_  = ~n913 ;
  assign \g11190/_00_  = n919 ;
  assign \g11297/_0_  = ~n943 ;
  assign \g11298/_0_  = ~n956 ;
  assign \g11300/_0_  = ~n967 ;
  assign \g11301/_0_  = ~n978 ;
  assign \g11303/_0_  = ~n989 ;
  assign \g11346/_0_  = ~n1000 ;
  assign \g11347/_0_  = ~n1011 ;
  assign \g11348/_0_  = ~n1022 ;
  assign \g11358/_0_  = ~n1035 ;
  assign \g11359/_0_  = ~n1048 ;
  assign \g11360/_0_  = ~n1061 ;
  assign \g11361/_0_  = ~n1074 ;
  assign \g11362/_0_  = ~n1087 ;
  assign \g11363/_0_  = ~n1100 ;
  assign \g11470/_0_  = ~n1109 ;
  assign \g11499/_0_  = ~n1118 ;
  assign \g11501/_0_  = ~n1124 ;
  assign \g11502/_0_  = ~n1127 ;
  assign \g11503/_0_  = ~n1135 ;
  assign \g11504/_0_  = ~n1141 ;
  assign \g11505/_0_  = ~n1146 ;
  assign \g11506/_0_  = ~n1150 ;
  assign \g11507/_0_  = ~n1154 ;
  assign \g11508/_0_  = ~n1158 ;
  assign \g11509/_0_  = ~n1161 ;
  assign \g11510/_0_  = ~n1165 ;
  assign \g11511/_0_  = ~n1169 ;
  assign \g11512/_0_  = ~n1173 ;
  assign \g11513/_0_  = ~n1177 ;
  assign \g11514/_0_  = ~n1181 ;
  assign \g11515/_0_  = ~n1184 ;
  assign \g11516/_0_  = ~n1187 ;
  assign \g11517/_0_  = ~n1191 ;
  assign \g11519/_0_  = ~n1194 ;
  assign \g11520/_0_  = ~n1197 ;
  assign \g11521/_0_  = ~n1201 ;
  assign \g11522/_0_  = ~n1204 ;
  assign \g11523/_0_  = ~n1207 ;
  assign \g11524/_0_  = ~n1211 ;
  assign \g11525/_0_  = ~n1214 ;
  assign \g11526/_0_  = ~n1218 ;
  assign \g11527/_0_  = ~n1222 ;
  assign \g11528/_0_  = ~n1225 ;
  assign \g11529/_0_  = ~n1228 ;
  assign \g11530/_0_  = ~n1232 ;
  assign \g11531/_0_  = ~n1235 ;
  assign \g11532/_0_  = ~n1238 ;
  assign \g11533/_0_  = ~n1241 ;
  assign \g11534/_0_  = ~n1244 ;
  assign \g11535/_0_  = ~n1247 ;
  assign \g11536/_0_  = ~n1250 ;
  assign \g11537/_0_  = ~n1253 ;
  assign \g11538/_0_  = ~n1256 ;
  assign \g11539/_0_  = ~n1259 ;
  assign \g11655/_0_  = ~n1266 ;
  assign \g11658/_0_  = ~n1273 ;
  assign \g11659/_0_  = ~n1280 ;
  assign \g11661/_0_  = ~n1287 ;
  assign \g11662/_0_  = ~n1294 ;
  assign \g11680/_0_  = ~n1301 ;
  assign \g11723/_0_  = ~n1308 ;
  assign \g11726/_0_  = ~n1315 ;
  assign \g11730/_0_  = ~n1322 ;
  assign \g11739/_0_  = ~n1329 ;
  assign \g11750/_0_  = ~n1336 ;
  assign \g11759/_0_  = ~n1343 ;
  assign \g11760/_0_  = ~n1350 ;
  assign \g11761/_0_  = ~n1357 ;
  assign \g11764/_0_  = ~n1364 ;
  assign \g11765/_0_  = ~n1371 ;
  assign \g12212/_0_  = n1373 ;
  assign \g13497/_0_  = ~n1897 ;
  assign \g13884/_0_  = ~n1915 ;
  assign \g13982/_0_  = ~n1930 ;
  assign \g13999/_0_  = ~n1944 ;
  assign \g9305/_0_  = ~n1959 ;
  assign \g9306/_0_  = ~n1968 ;
  assign \g9307/_0_  = ~n1982 ;
  assign \g9308/_0_  = ~n1992 ;
  assign \g9309/_0_  = ~n2012 ;
  assign \g9310/_0_  = ~n2026 ;
  assign \g9346/_0_  = ~n2041 ;
  assign \g9347/_0_  = ~n2054 ;
  assign \g9348/_0_  = ~n2068 ;
  assign \g9349/_0_  = ~n2082 ;
  assign \g9350/_0_  = ~n2095 ;
  assign \g9351/_0_  = ~n2107 ;
  assign \g9352/_0_  = ~n2119 ;
  assign \g9353/_0_  = ~n2133 ;
  assign \g9354/_0_  = ~n2146 ;
  assign \g9355/_0_  = ~n2159 ;
  assign \g9356/_0_  = ~n2171 ;
  assign \g9357/_0_  = ~n2185 ;
  assign \g9358/_0_  = ~n2197 ;
  assign \g9359/_0_  = ~n2209 ;
  assign \g9360/_0_  = ~n2221 ;
  assign \g9361/_0_  = ~n2234 ;
  assign \g9362/_0_  = ~n2247 ;
  assign \g9363/_0_  = ~n2260 ;
  assign \g9364/_0_  = ~n2274 ;
  assign \g9365/_0_  = ~n2287 ;
  assign \g9366/_0_  = ~n2300 ;
  assign \g9367/_0_  = ~n2313 ;
  assign \g9368/_0_  = ~n2326 ;
  assign \g9369/_0_  = ~n2338 ;
  assign \g9370/_0_  = ~n2350 ;
  assign \g9371/_0_  = ~n2363 ;
  assign \g9372/_0_  = ~n2376 ;
  assign \g9373/_0_  = ~n2389 ;
  assign \g9374/_0_  = ~n2402 ;
  assign \g9375/_0_  = ~n2414 ;
  assign \g9380/_0_  = ~n2427 ;
  assign \g9381/_0_  = ~n2436 ;
  assign \g9382/_0_  = ~n2445 ;
  assign \g9383/_0_  = ~n2454 ;
  assign \g9384/_0_  = ~n2463 ;
  assign \g9385/_0_  = ~n2476 ;
  assign \g9386/_0_  = ~n2485 ;
  assign \g9387/_0_  = ~n2494 ;
  assign \g9388/_0_  = ~n2505 ;
  assign \g9389/_0_  = ~n2517 ;
  assign \g9390/_0_  = ~n2527 ;
  assign \g9391/_0_  = ~n2537 ;
  assign \g9392/_0_  = ~n2549 ;
  assign \g9393/_0_  = ~n2562 ;
  assign \g9394/_0_  = ~n2571 ;
  assign \g9395/_0_  = ~n2580 ;
  assign \g9396/_0_  = ~n2592 ;
  assign \g9397/_0_  = ~n2601 ;
  assign \g9398/_0_  = ~n2613 ;
  assign \g9399/_0_  = ~n2622 ;
  assign \g9400/_0_  = ~n2631 ;
  assign \g9401/_0_  = ~n2643 ;
  assign \g9402/_0_  = ~n2655 ;
  assign \g9403/_0_  = ~n2665 ;
  assign \g9404/_0_  = ~n2674 ;
  assign \g9405/_0_  = ~n2683 ;
  assign \g9406/_0_  = ~n2695 ;
  assign \g9407/_0_  = ~n2704 ;
  assign \g9408/_0_  = ~n2713 ;
  assign \g9409/_0_  = ~n2722 ;
  assign \g9410/_0_  = ~n2734 ;
  assign \g9411/_0_  = ~n2744 ;
  assign \g9439/_0_  = ~n2753 ;
  assign \g9440/_0_  = ~n2762 ;
  assign \g9441/_0_  = ~n2771 ;
  assign \g9442/_0_  = ~n2780 ;
  assign \g9443/_0_  = ~n2789 ;
  assign \g9444/_0_  = ~n2798 ;
  assign \g9445/_0_  = ~n2810 ;
  assign \g9446/_0_  = ~n2819 ;
  assign \g9447/_0_  = ~n2828 ;
  assign \g9448/_0_  = ~n2837 ;
  assign \g9449/_0_  = ~n2846 ;
  assign \g9450/_0_  = ~n2855 ;
  assign \g9451/_0_  = ~n2864 ;
  assign \g9452/_0_  = ~n2873 ;
  assign \g9453/_0_  = ~n2882 ;
  assign \g9454/_0_  = ~n2891 ;
  assign \g9455/_0_  = ~n2900 ;
  assign \g9456/_0_  = ~n2910 ;
  assign \g9457/_0_  = ~n2919 ;
  assign \g9458/_0_  = ~n2929 ;
  assign \g9459/_0_  = ~n2939 ;
  assign \g9461/_0_  = ~n2948 ;
  assign \g9462/_0_  = ~n2957 ;
  assign \g9463/_0_  = ~n2966 ;
  assign \g9464/_0_  = ~n2975 ;
  assign \g9465/_0_  = ~n2984 ;
  assign \g9466/_0_  = ~n2993 ;
  assign \g9529/_0_  = ~n3005 ;
  assign \g9530/_0_  = ~n3018 ;
  assign \g9531/_0_  = ~n3030 ;
  assign \g9532/_0_  = ~n3042 ;
  assign \g9535/_0_  = ~n3054 ;
  assign \g9542/_0_  = ~n3063 ;
  assign \g9543/_0_  = ~n3075 ;
  assign \g9546/_0_  = ~n3088 ;
  assign \g9547/_0_  = ~n3100 ;
  assign \g9548/_0_  = ~n3112 ;
  assign \g9549/_0_  = ~n3124 ;
  assign \g9550/_0_  = ~n3136 ;
  assign \g9551/_0_  = ~n3145 ;
  assign \g9552/_0_  = ~n3154 ;
  assign \g9553/_0_  = ~n3166 ;
  assign \g9559/_0_  = ~n3178 ;
  assign \g9568/_0_  = ~n3190 ;
  assign \g9571/_0_  = ~n3202 ;
  assign \g9573/_0_  = ~n3214 ;
  assign \g9583/_0_  = ~n3226 ;
  assign \g9589/_0_  = ~n3239 ;
  assign \g9590/_0_  = ~n3248 ;
  assign \g9591/_0_  = ~n3257 ;
  assign \g9592/_0_  = ~n3266 ;
  assign \g9593/_0_  = ~n3275 ;
  assign \g9594/_0_  = ~n3288 ;
  assign \g9595/_0_  = ~n3300 ;
  assign \g9596/_0_  = ~n3312 ;
  assign \g9597/_0_  = ~n3324 ;
  assign \ss_pad_o[0]_pad  = ~n3326 ;
  assign \ss_pad_o[1]_pad  = ~n3327 ;
  assign \ss_pad_o[2]_pad  = ~n3328 ;
  assign \ss_pad_o[3]_pad  = ~n3329 ;
  assign \ss_pad_o[4]_pad  = ~n3330 ;
  assign \ss_pad_o[5]_pad  = ~n3331 ;
  assign \ss_pad_o[6]_pad  = ~n3332 ;
  assign \ss_pad_o[7]_pad  = ~n3333 ;
  assign wb_err_o_pad = 1'b0 ;
endmodule
