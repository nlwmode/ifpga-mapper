module top( \count[0]  , \count[1]  , \count[2]  , \count[3]  , \count[4]  , \count[5]  , \count[6]  , \count[7]  , \selectp1[0]  , \selectp1[1]  , \selectp1[2]  , \selectp1[3]  , \selectp1[4]  , \selectp1[5]  , \selectp1[6]  , \selectp1[7]  , \selectp1[8]  , \selectp1[9]  , \selectp1[10]  , \selectp1[11]  , \selectp1[12]  , \selectp1[13]  , \selectp1[14]  , \selectp1[15]  , \selectp1[16]  , \selectp1[17]  , \selectp1[18]  , \selectp1[19]  , \selectp1[20]  , \selectp1[21]  , \selectp1[22]  , \selectp1[23]  , \selectp1[24]  , \selectp1[25]  , \selectp1[26]  , \selectp1[27]  , \selectp1[28]  , \selectp1[29]  , \selectp1[30]  , \selectp1[31]  , \selectp1[32]  , \selectp1[33]  , \selectp1[34]  , \selectp1[35]  , \selectp1[36]  , \selectp1[37]  , \selectp1[38]  , \selectp1[39]  , \selectp1[40]  , \selectp1[41]  , \selectp1[42]  , \selectp1[43]  , \selectp1[44]  , \selectp1[45]  , \selectp1[46]  , \selectp1[47]  , \selectp1[48]  , \selectp1[49]  , \selectp1[50]  , \selectp1[51]  , \selectp1[52]  , \selectp1[53]  , \selectp1[54]  , \selectp1[55]  , \selectp1[56]  , \selectp1[57]  , \selectp1[58]  , \selectp1[59]  , \selectp1[60]  , \selectp1[61]  , \selectp1[62]  , \selectp1[63]  , \selectp1[64]  , \selectp1[65]  , \selectp1[66]  , \selectp1[67]  , \selectp1[68]  , \selectp1[69]  , \selectp1[70]  , \selectp1[71]  , \selectp1[72]  , \selectp1[73]  , \selectp1[74]  , \selectp1[75]  , \selectp1[76]  , \selectp1[77]  , \selectp1[78]  , \selectp1[79]  , \selectp1[80]  , \selectp1[81]  , \selectp1[82]  , \selectp1[83]  , \selectp1[84]  , \selectp1[85]  , \selectp1[86]  , \selectp1[87]  , \selectp1[88]  , \selectp1[89]  , \selectp1[90]  , \selectp1[91]  , \selectp1[92]  , \selectp1[93]  , \selectp1[94]  , \selectp1[95]  , \selectp1[96]  , \selectp1[97]  , \selectp1[98]  , \selectp1[99]  , \selectp1[100]  , \selectp1[101]  , \selectp1[102]  , \selectp1[103]  , \selectp1[104]  , \selectp1[105]  , \selectp1[106]  , \selectp1[107]  , \selectp1[108]  , \selectp1[109]  , \selectp1[110]  , \selectp1[111]  , \selectp1[112]  , \selectp1[113]  , \selectp1[114]  , \selectp1[115]  , \selectp1[116]  , \selectp1[117]  , \selectp1[118]  , \selectp1[119]  , \selectp1[120]  , \selectp1[121]  , \selectp1[122]  , \selectp1[123]  , \selectp1[124]  , \selectp1[125]  , \selectp1[126]  , \selectp1[127]  , \selectp2[0]  , \selectp2[1]  , \selectp2[2]  , \selectp2[3]  , \selectp2[4]  , \selectp2[5]  , \selectp2[6]  , \selectp2[7]  , \selectp2[8]  , \selectp2[9]  , \selectp2[10]  , \selectp2[11]  , \selectp2[12]  , \selectp2[13]  , \selectp2[14]  , \selectp2[15]  , \selectp2[16]  , \selectp2[17]  , \selectp2[18]  , \selectp2[19]  , \selectp2[20]  , \selectp2[21]  , \selectp2[22]  , \selectp2[23]  , \selectp2[24]  , \selectp2[25]  , \selectp2[26]  , \selectp2[27]  , \selectp2[28]  , \selectp2[29]  , \selectp2[30]  , \selectp2[31]  , \selectp2[32]  , \selectp2[33]  , \selectp2[34]  , \selectp2[35]  , \selectp2[36]  , \selectp2[37]  , \selectp2[38]  , \selectp2[39]  , \selectp2[40]  , \selectp2[41]  , \selectp2[42]  , \selectp2[43]  , \selectp2[44]  , \selectp2[45]  , \selectp2[46]  , \selectp2[47]  , \selectp2[48]  , \selectp2[49]  , \selectp2[50]  , \selectp2[51]  , \selectp2[52]  , \selectp2[53]  , \selectp2[54]  , \selectp2[55]  , \selectp2[56]  , \selectp2[57]  , \selectp2[58]  , \selectp2[59]  , \selectp2[60]  , \selectp2[61]  , \selectp2[62]  , \selectp2[63]  , \selectp2[64]  , \selectp2[65]  , \selectp2[66]  , \selectp2[67]  , \selectp2[68]  , \selectp2[69]  , \selectp2[70]  , \selectp2[71]  , \selectp2[72]  , \selectp2[73]  , \selectp2[74]  , \selectp2[75]  , \selectp2[76]  , \selectp2[77]  , \selectp2[78]  , \selectp2[79]  , \selectp2[80]  , \selectp2[81]  , \selectp2[82]  , \selectp2[83]  , \selectp2[84]  , \selectp2[85]  , \selectp2[86]  , \selectp2[87]  , \selectp2[88]  , \selectp2[89]  , \selectp2[90]  , \selectp2[91]  , \selectp2[92]  , \selectp2[93]  , \selectp2[94]  , \selectp2[95]  , \selectp2[96]  , \selectp2[97]  , \selectp2[98]  , \selectp2[99]  , \selectp2[100]  , \selectp2[101]  , \selectp2[102]  , \selectp2[103]  , \selectp2[104]  , \selectp2[105]  , \selectp2[106]  , \selectp2[107]  , \selectp2[108]  , \selectp2[109]  , \selectp2[110]  , \selectp2[111]  , \selectp2[112]  , \selectp2[113]  , \selectp2[114]  , \selectp2[115]  , \selectp2[116]  , \selectp2[117]  , \selectp2[118]  , \selectp2[119]  , \selectp2[120]  , \selectp2[121]  , \selectp2[122]  , \selectp2[123]  , \selectp2[124]  , \selectp2[125]  , \selectp2[126]  , \selectp2[127]  );
  input \count[0]  ;
  input \count[1]  ;
  input \count[2]  ;
  input \count[3]  ;
  input \count[4]  ;
  input \count[5]  ;
  input \count[6]  ;
  input \count[7]  ;
  output \selectp1[0]  ;
  output \selectp1[1]  ;
  output \selectp1[2]  ;
  output \selectp1[3]  ;
  output \selectp1[4]  ;
  output \selectp1[5]  ;
  output \selectp1[6]  ;
  output \selectp1[7]  ;
  output \selectp1[8]  ;
  output \selectp1[9]  ;
  output \selectp1[10]  ;
  output \selectp1[11]  ;
  output \selectp1[12]  ;
  output \selectp1[13]  ;
  output \selectp1[14]  ;
  output \selectp1[15]  ;
  output \selectp1[16]  ;
  output \selectp1[17]  ;
  output \selectp1[18]  ;
  output \selectp1[19]  ;
  output \selectp1[20]  ;
  output \selectp1[21]  ;
  output \selectp1[22]  ;
  output \selectp1[23]  ;
  output \selectp1[24]  ;
  output \selectp1[25]  ;
  output \selectp1[26]  ;
  output \selectp1[27]  ;
  output \selectp1[28]  ;
  output \selectp1[29]  ;
  output \selectp1[30]  ;
  output \selectp1[31]  ;
  output \selectp1[32]  ;
  output \selectp1[33]  ;
  output \selectp1[34]  ;
  output \selectp1[35]  ;
  output \selectp1[36]  ;
  output \selectp1[37]  ;
  output \selectp1[38]  ;
  output \selectp1[39]  ;
  output \selectp1[40]  ;
  output \selectp1[41]  ;
  output \selectp1[42]  ;
  output \selectp1[43]  ;
  output \selectp1[44]  ;
  output \selectp1[45]  ;
  output \selectp1[46]  ;
  output \selectp1[47]  ;
  output \selectp1[48]  ;
  output \selectp1[49]  ;
  output \selectp1[50]  ;
  output \selectp1[51]  ;
  output \selectp1[52]  ;
  output \selectp1[53]  ;
  output \selectp1[54]  ;
  output \selectp1[55]  ;
  output \selectp1[56]  ;
  output \selectp1[57]  ;
  output \selectp1[58]  ;
  output \selectp1[59]  ;
  output \selectp1[60]  ;
  output \selectp1[61]  ;
  output \selectp1[62]  ;
  output \selectp1[63]  ;
  output \selectp1[64]  ;
  output \selectp1[65]  ;
  output \selectp1[66]  ;
  output \selectp1[67]  ;
  output \selectp1[68]  ;
  output \selectp1[69]  ;
  output \selectp1[70]  ;
  output \selectp1[71]  ;
  output \selectp1[72]  ;
  output \selectp1[73]  ;
  output \selectp1[74]  ;
  output \selectp1[75]  ;
  output \selectp1[76]  ;
  output \selectp1[77]  ;
  output \selectp1[78]  ;
  output \selectp1[79]  ;
  output \selectp1[80]  ;
  output \selectp1[81]  ;
  output \selectp1[82]  ;
  output \selectp1[83]  ;
  output \selectp1[84]  ;
  output \selectp1[85]  ;
  output \selectp1[86]  ;
  output \selectp1[87]  ;
  output \selectp1[88]  ;
  output \selectp1[89]  ;
  output \selectp1[90]  ;
  output \selectp1[91]  ;
  output \selectp1[92]  ;
  output \selectp1[93]  ;
  output \selectp1[94]  ;
  output \selectp1[95]  ;
  output \selectp1[96]  ;
  output \selectp1[97]  ;
  output \selectp1[98]  ;
  output \selectp1[99]  ;
  output \selectp1[100]  ;
  output \selectp1[101]  ;
  output \selectp1[102]  ;
  output \selectp1[103]  ;
  output \selectp1[104]  ;
  output \selectp1[105]  ;
  output \selectp1[106]  ;
  output \selectp1[107]  ;
  output \selectp1[108]  ;
  output \selectp1[109]  ;
  output \selectp1[110]  ;
  output \selectp1[111]  ;
  output \selectp1[112]  ;
  output \selectp1[113]  ;
  output \selectp1[114]  ;
  output \selectp1[115]  ;
  output \selectp1[116]  ;
  output \selectp1[117]  ;
  output \selectp1[118]  ;
  output \selectp1[119]  ;
  output \selectp1[120]  ;
  output \selectp1[121]  ;
  output \selectp1[122]  ;
  output \selectp1[123]  ;
  output \selectp1[124]  ;
  output \selectp1[125]  ;
  output \selectp1[126]  ;
  output \selectp1[127]  ;
  output \selectp2[0]  ;
  output \selectp2[1]  ;
  output \selectp2[2]  ;
  output \selectp2[3]  ;
  output \selectp2[4]  ;
  output \selectp2[5]  ;
  output \selectp2[6]  ;
  output \selectp2[7]  ;
  output \selectp2[8]  ;
  output \selectp2[9]  ;
  output \selectp2[10]  ;
  output \selectp2[11]  ;
  output \selectp2[12]  ;
  output \selectp2[13]  ;
  output \selectp2[14]  ;
  output \selectp2[15]  ;
  output \selectp2[16]  ;
  output \selectp2[17]  ;
  output \selectp2[18]  ;
  output \selectp2[19]  ;
  output \selectp2[20]  ;
  output \selectp2[21]  ;
  output \selectp2[22]  ;
  output \selectp2[23]  ;
  output \selectp2[24]  ;
  output \selectp2[25]  ;
  output \selectp2[26]  ;
  output \selectp2[27]  ;
  output \selectp2[28]  ;
  output \selectp2[29]  ;
  output \selectp2[30]  ;
  output \selectp2[31]  ;
  output \selectp2[32]  ;
  output \selectp2[33]  ;
  output \selectp2[34]  ;
  output \selectp2[35]  ;
  output \selectp2[36]  ;
  output \selectp2[37]  ;
  output \selectp2[38]  ;
  output \selectp2[39]  ;
  output \selectp2[40]  ;
  output \selectp2[41]  ;
  output \selectp2[42]  ;
  output \selectp2[43]  ;
  output \selectp2[44]  ;
  output \selectp2[45]  ;
  output \selectp2[46]  ;
  output \selectp2[47]  ;
  output \selectp2[48]  ;
  output \selectp2[49]  ;
  output \selectp2[50]  ;
  output \selectp2[51]  ;
  output \selectp2[52]  ;
  output \selectp2[53]  ;
  output \selectp2[54]  ;
  output \selectp2[55]  ;
  output \selectp2[56]  ;
  output \selectp2[57]  ;
  output \selectp2[58]  ;
  output \selectp2[59]  ;
  output \selectp2[60]  ;
  output \selectp2[61]  ;
  output \selectp2[62]  ;
  output \selectp2[63]  ;
  output \selectp2[64]  ;
  output \selectp2[65]  ;
  output \selectp2[66]  ;
  output \selectp2[67]  ;
  output \selectp2[68]  ;
  output \selectp2[69]  ;
  output \selectp2[70]  ;
  output \selectp2[71]  ;
  output \selectp2[72]  ;
  output \selectp2[73]  ;
  output \selectp2[74]  ;
  output \selectp2[75]  ;
  output \selectp2[76]  ;
  output \selectp2[77]  ;
  output \selectp2[78]  ;
  output \selectp2[79]  ;
  output \selectp2[80]  ;
  output \selectp2[81]  ;
  output \selectp2[82]  ;
  output \selectp2[83]  ;
  output \selectp2[84]  ;
  output \selectp2[85]  ;
  output \selectp2[86]  ;
  output \selectp2[87]  ;
  output \selectp2[88]  ;
  output \selectp2[89]  ;
  output \selectp2[90]  ;
  output \selectp2[91]  ;
  output \selectp2[92]  ;
  output \selectp2[93]  ;
  output \selectp2[94]  ;
  output \selectp2[95]  ;
  output \selectp2[96]  ;
  output \selectp2[97]  ;
  output \selectp2[98]  ;
  output \selectp2[99]  ;
  output \selectp2[100]  ;
  output \selectp2[101]  ;
  output \selectp2[102]  ;
  output \selectp2[103]  ;
  output \selectp2[104]  ;
  output \selectp2[105]  ;
  output \selectp2[106]  ;
  output \selectp2[107]  ;
  output \selectp2[108]  ;
  output \selectp2[109]  ;
  output \selectp2[110]  ;
  output \selectp2[111]  ;
  output \selectp2[112]  ;
  output \selectp2[113]  ;
  output \selectp2[114]  ;
  output \selectp2[115]  ;
  output \selectp2[116]  ;
  output \selectp2[117]  ;
  output \selectp2[118]  ;
  output \selectp2[119]  ;
  output \selectp2[120]  ;
  output \selectp2[121]  ;
  output \selectp2[122]  ;
  output \selectp2[123]  ;
  output \selectp2[124]  ;
  output \selectp2[125]  ;
  output \selectp2[126]  ;
  output \selectp2[127]  ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 ;
  assign n9 = ~\count[4]  & ~\count[5]  ;
  assign n10 = ~\count[6]  & \count[7]  ;
  assign n11 = n9 & n10 ;
  assign n12 = ~\count[0]  & ~\count[2]  ;
  assign n13 = ~\count[1]  & ~\count[3]  ;
  assign n14 = n12 & n13 ;
  assign n15 = n11 & n14 ;
  assign n16 = \count[0]  & ~\count[2]  ;
  assign n17 = n13 & n16 ;
  assign n18 = n11 & n17 ;
  assign n19 = \count[1]  & ~\count[3]  ;
  assign n20 = n12 & n19 ;
  assign n21 = n11 & n20 ;
  assign n22 = n16 & n19 ;
  assign n23 = n11 & n22 ;
  assign n24 = ~\count[0]  & \count[2]  ;
  assign n25 = n13 & n24 ;
  assign n26 = n11 & n25 ;
  assign n27 = \count[0]  & \count[2]  ;
  assign n28 = n13 & n27 ;
  assign n29 = n11 & n28 ;
  assign n30 = n19 & n24 ;
  assign n31 = n11 & n30 ;
  assign n32 = n19 & n27 ;
  assign n33 = n11 & n32 ;
  assign n34 = ~\count[1]  & \count[3]  ;
  assign n35 = n12 & n34 ;
  assign n36 = n11 & n35 ;
  assign n37 = n16 & n34 ;
  assign n38 = n11 & n37 ;
  assign n39 = \count[1]  & \count[3]  ;
  assign n40 = n12 & n39 ;
  assign n41 = n11 & n40 ;
  assign n42 = n16 & n39 ;
  assign n43 = n11 & n42 ;
  assign n44 = n24 & n34 ;
  assign n45 = n11 & n44 ;
  assign n46 = n27 & n34 ;
  assign n47 = n11 & n46 ;
  assign n48 = n24 & n39 ;
  assign n49 = n11 & n48 ;
  assign n50 = n27 & n39 ;
  assign n51 = n11 & n50 ;
  assign n52 = \count[4]  & ~\count[5]  ;
  assign n53 = n10 & n52 ;
  assign n54 = n14 & n53 ;
  assign n55 = n17 & n53 ;
  assign n56 = n20 & n53 ;
  assign n57 = n22 & n53 ;
  assign n58 = n25 & n53 ;
  assign n59 = n28 & n53 ;
  assign n60 = n30 & n53 ;
  assign n61 = n32 & n53 ;
  assign n62 = n35 & n53 ;
  assign n63 = n37 & n53 ;
  assign n64 = n40 & n53 ;
  assign n65 = n42 & n53 ;
  assign n66 = n44 & n53 ;
  assign n67 = n46 & n53 ;
  assign n68 = n48 & n53 ;
  assign n69 = n50 & n53 ;
  assign n70 = ~\count[4]  & \count[5]  ;
  assign n71 = n10 & n70 ;
  assign n72 = n14 & n71 ;
  assign n73 = n17 & n71 ;
  assign n74 = n20 & n71 ;
  assign n75 = n22 & n71 ;
  assign n76 = n25 & n71 ;
  assign n77 = n28 & n71 ;
  assign n78 = n30 & n71 ;
  assign n79 = n32 & n71 ;
  assign n80 = n35 & n71 ;
  assign n81 = n37 & n71 ;
  assign n82 = n40 & n71 ;
  assign n83 = n42 & n71 ;
  assign n84 = n44 & n71 ;
  assign n85 = n46 & n71 ;
  assign n86 = n48 & n71 ;
  assign n87 = n50 & n71 ;
  assign n88 = \count[4]  & \count[5]  ;
  assign n89 = n10 & n88 ;
  assign n90 = n14 & n89 ;
  assign n91 = n17 & n89 ;
  assign n92 = n20 & n89 ;
  assign n93 = n22 & n89 ;
  assign n94 = n25 & n89 ;
  assign n95 = n28 & n89 ;
  assign n96 = n30 & n89 ;
  assign n97 = n32 & n89 ;
  assign n98 = n35 & n89 ;
  assign n99 = n37 & n89 ;
  assign n100 = n40 & n89 ;
  assign n101 = n42 & n89 ;
  assign n102 = n44 & n89 ;
  assign n103 = n46 & n89 ;
  assign n104 = n48 & n89 ;
  assign n105 = n50 & n89 ;
  assign n106 = \count[6]  & \count[7]  ;
  assign n107 = n9 & n106 ;
  assign n108 = n14 & n107 ;
  assign n109 = n17 & n107 ;
  assign n110 = n20 & n107 ;
  assign n111 = n22 & n107 ;
  assign n112 = n25 & n107 ;
  assign n113 = n28 & n107 ;
  assign n114 = n30 & n107 ;
  assign n115 = n32 & n107 ;
  assign n116 = n35 & n107 ;
  assign n117 = n37 & n107 ;
  assign n118 = n40 & n107 ;
  assign n119 = n42 & n107 ;
  assign n120 = n44 & n107 ;
  assign n121 = n46 & n107 ;
  assign n122 = n48 & n107 ;
  assign n123 = n50 & n107 ;
  assign n124 = n52 & n106 ;
  assign n125 = n14 & n124 ;
  assign n126 = n17 & n124 ;
  assign n127 = n20 & n124 ;
  assign n128 = n22 & n124 ;
  assign n129 = n25 & n124 ;
  assign n130 = n28 & n124 ;
  assign n131 = n30 & n124 ;
  assign n132 = n32 & n124 ;
  assign n133 = n35 & n124 ;
  assign n134 = n37 & n124 ;
  assign n135 = n40 & n124 ;
  assign n136 = n42 & n124 ;
  assign n137 = n44 & n124 ;
  assign n138 = n46 & n124 ;
  assign n139 = n48 & n124 ;
  assign n140 = n50 & n124 ;
  assign n141 = n70 & n106 ;
  assign n142 = n14 & n141 ;
  assign n143 = n17 & n141 ;
  assign n144 = n20 & n141 ;
  assign n145 = n22 & n141 ;
  assign n146 = n25 & n141 ;
  assign n147 = n28 & n141 ;
  assign n148 = n30 & n141 ;
  assign n149 = n32 & n141 ;
  assign n150 = n35 & n141 ;
  assign n151 = n37 & n141 ;
  assign n152 = n40 & n141 ;
  assign n153 = n42 & n141 ;
  assign n154 = n44 & n141 ;
  assign n155 = n46 & n141 ;
  assign n156 = n48 & n141 ;
  assign n157 = n50 & n141 ;
  assign n158 = n88 & n106 ;
  assign n159 = n14 & n158 ;
  assign n160 = n17 & n158 ;
  assign n161 = n20 & n158 ;
  assign n162 = n22 & n158 ;
  assign n163 = n25 & n158 ;
  assign n164 = n28 & n158 ;
  assign n165 = n30 & n158 ;
  assign n166 = n32 & n158 ;
  assign n167 = n35 & n158 ;
  assign n168 = n37 & n158 ;
  assign n169 = n40 & n158 ;
  assign n170 = n42 & n158 ;
  assign n171 = n44 & n158 ;
  assign n172 = n46 & n158 ;
  assign n173 = n48 & n158 ;
  assign n174 = n50 & n158 ;
  assign n175 = ~\count[6]  & ~\count[7]  ;
  assign n176 = n9 & n175 ;
  assign n177 = n14 & n176 ;
  assign n178 = n17 & n176 ;
  assign n179 = n20 & n176 ;
  assign n180 = n22 & n176 ;
  assign n181 = n25 & n176 ;
  assign n182 = n28 & n176 ;
  assign n183 = n30 & n176 ;
  assign n184 = n32 & n176 ;
  assign n185 = n35 & n176 ;
  assign n186 = n37 & n176 ;
  assign n187 = n40 & n176 ;
  assign n188 = n42 & n176 ;
  assign n189 = n44 & n176 ;
  assign n190 = n46 & n176 ;
  assign n191 = n48 & n176 ;
  assign n192 = n50 & n176 ;
  assign n193 = n52 & n175 ;
  assign n194 = n14 & n193 ;
  assign n195 = n17 & n193 ;
  assign n196 = n20 & n193 ;
  assign n197 = n22 & n193 ;
  assign n198 = n25 & n193 ;
  assign n199 = n28 & n193 ;
  assign n200 = n30 & n193 ;
  assign n201 = n32 & n193 ;
  assign n202 = n35 & n193 ;
  assign n203 = n37 & n193 ;
  assign n204 = n40 & n193 ;
  assign n205 = n42 & n193 ;
  assign n206 = n44 & n193 ;
  assign n207 = n46 & n193 ;
  assign n208 = n48 & n193 ;
  assign n209 = n50 & n193 ;
  assign n210 = n70 & n175 ;
  assign n211 = n14 & n210 ;
  assign n212 = n17 & n210 ;
  assign n213 = n20 & n210 ;
  assign n214 = n22 & n210 ;
  assign n215 = n25 & n210 ;
  assign n216 = n28 & n210 ;
  assign n217 = n30 & n210 ;
  assign n218 = n32 & n210 ;
  assign n219 = n35 & n210 ;
  assign n220 = n37 & n210 ;
  assign n221 = n40 & n210 ;
  assign n222 = n42 & n210 ;
  assign n223 = n44 & n210 ;
  assign n224 = n46 & n210 ;
  assign n225 = n48 & n210 ;
  assign n226 = n50 & n210 ;
  assign n227 = n88 & n175 ;
  assign n228 = n14 & n227 ;
  assign n229 = n17 & n227 ;
  assign n230 = n20 & n227 ;
  assign n231 = n22 & n227 ;
  assign n232 = n25 & n227 ;
  assign n233 = n28 & n227 ;
  assign n234 = n30 & n227 ;
  assign n235 = n32 & n227 ;
  assign n236 = n35 & n227 ;
  assign n237 = n37 & n227 ;
  assign n238 = n40 & n227 ;
  assign n239 = n42 & n227 ;
  assign n240 = n44 & n227 ;
  assign n241 = n46 & n227 ;
  assign n242 = n48 & n227 ;
  assign n243 = n50 & n227 ;
  assign n244 = \count[6]  & ~\count[7]  ;
  assign n245 = n9 & n244 ;
  assign n246 = n14 & n245 ;
  assign n247 = n17 & n245 ;
  assign n248 = n20 & n245 ;
  assign n249 = n22 & n245 ;
  assign n250 = n25 & n245 ;
  assign n251 = n28 & n245 ;
  assign n252 = n30 & n245 ;
  assign n253 = n32 & n245 ;
  assign n254 = n35 & n245 ;
  assign n255 = n37 & n245 ;
  assign n256 = n40 & n245 ;
  assign n257 = n42 & n245 ;
  assign n258 = n44 & n245 ;
  assign n259 = n46 & n245 ;
  assign n260 = n48 & n245 ;
  assign n261 = n50 & n245 ;
  assign n262 = n52 & n244 ;
  assign n263 = n14 & n262 ;
  assign n264 = n17 & n262 ;
  assign n265 = n20 & n262 ;
  assign n266 = n22 & n262 ;
  assign n267 = n25 & n262 ;
  assign n268 = n28 & n262 ;
  assign n269 = n30 & n262 ;
  assign n270 = n32 & n262 ;
  assign n271 = n35 & n262 ;
  assign n272 = n37 & n262 ;
  assign n273 = n40 & n262 ;
  assign n274 = n42 & n262 ;
  assign n275 = n44 & n262 ;
  assign n276 = n46 & n262 ;
  assign n277 = n48 & n262 ;
  assign n278 = n50 & n262 ;
  assign n279 = n70 & n244 ;
  assign n280 = n14 & n279 ;
  assign n281 = n17 & n279 ;
  assign n282 = n20 & n279 ;
  assign n283 = n22 & n279 ;
  assign n284 = n25 & n279 ;
  assign n285 = n28 & n279 ;
  assign n286 = n30 & n279 ;
  assign n287 = n32 & n279 ;
  assign n288 = n35 & n279 ;
  assign n289 = n37 & n279 ;
  assign n290 = n40 & n279 ;
  assign n291 = n42 & n279 ;
  assign n292 = n44 & n279 ;
  assign n293 = n46 & n279 ;
  assign n294 = n48 & n279 ;
  assign n295 = n50 & n279 ;
  assign n296 = n88 & n244 ;
  assign n297 = n14 & n296 ;
  assign n298 = n17 & n296 ;
  assign n299 = n20 & n296 ;
  assign n300 = n22 & n296 ;
  assign n301 = n25 & n296 ;
  assign n302 = n28 & n296 ;
  assign n303 = n30 & n296 ;
  assign n304 = n32 & n296 ;
  assign n305 = n35 & n296 ;
  assign n306 = n37 & n296 ;
  assign n307 = n40 & n296 ;
  assign n308 = n42 & n296 ;
  assign n309 = n44 & n296 ;
  assign n310 = n46 & n296 ;
  assign n311 = n48 & n296 ;
  assign n312 = n50 & n296 ;
  assign \selectp1[0]  = n15 ;
  assign \selectp1[1]  = n18 ;
  assign \selectp1[2]  = n21 ;
  assign \selectp1[3]  = n23 ;
  assign \selectp1[4]  = n26 ;
  assign \selectp1[5]  = n29 ;
  assign \selectp1[6]  = n31 ;
  assign \selectp1[7]  = n33 ;
  assign \selectp1[8]  = n36 ;
  assign \selectp1[9]  = n38 ;
  assign \selectp1[10]  = n41 ;
  assign \selectp1[11]  = n43 ;
  assign \selectp1[12]  = n45 ;
  assign \selectp1[13]  = n47 ;
  assign \selectp1[14]  = n49 ;
  assign \selectp1[15]  = n51 ;
  assign \selectp1[16]  = n54 ;
  assign \selectp1[17]  = n55 ;
  assign \selectp1[18]  = n56 ;
  assign \selectp1[19]  = n57 ;
  assign \selectp1[20]  = n58 ;
  assign \selectp1[21]  = n59 ;
  assign \selectp1[22]  = n60 ;
  assign \selectp1[23]  = n61 ;
  assign \selectp1[24]  = n62 ;
  assign \selectp1[25]  = n63 ;
  assign \selectp1[26]  = n64 ;
  assign \selectp1[27]  = n65 ;
  assign \selectp1[28]  = n66 ;
  assign \selectp1[29]  = n67 ;
  assign \selectp1[30]  = n68 ;
  assign \selectp1[31]  = n69 ;
  assign \selectp1[32]  = n72 ;
  assign \selectp1[33]  = n73 ;
  assign \selectp1[34]  = n74 ;
  assign \selectp1[35]  = n75 ;
  assign \selectp1[36]  = n76 ;
  assign \selectp1[37]  = n77 ;
  assign \selectp1[38]  = n78 ;
  assign \selectp1[39]  = n79 ;
  assign \selectp1[40]  = n80 ;
  assign \selectp1[41]  = n81 ;
  assign \selectp1[42]  = n82 ;
  assign \selectp1[43]  = n83 ;
  assign \selectp1[44]  = n84 ;
  assign \selectp1[45]  = n85 ;
  assign \selectp1[46]  = n86 ;
  assign \selectp1[47]  = n87 ;
  assign \selectp1[48]  = n90 ;
  assign \selectp1[49]  = n91 ;
  assign \selectp1[50]  = n92 ;
  assign \selectp1[51]  = n93 ;
  assign \selectp1[52]  = n94 ;
  assign \selectp1[53]  = n95 ;
  assign \selectp1[54]  = n96 ;
  assign \selectp1[55]  = n97 ;
  assign \selectp1[56]  = n98 ;
  assign \selectp1[57]  = n99 ;
  assign \selectp1[58]  = n100 ;
  assign \selectp1[59]  = n101 ;
  assign \selectp1[60]  = n102 ;
  assign \selectp1[61]  = n103 ;
  assign \selectp1[62]  = n104 ;
  assign \selectp1[63]  = n105 ;
  assign \selectp1[64]  = n108 ;
  assign \selectp1[65]  = n109 ;
  assign \selectp1[66]  = n110 ;
  assign \selectp1[67]  = n111 ;
  assign \selectp1[68]  = n112 ;
  assign \selectp1[69]  = n113 ;
  assign \selectp1[70]  = n114 ;
  assign \selectp1[71]  = n115 ;
  assign \selectp1[72]  = n116 ;
  assign \selectp1[73]  = n117 ;
  assign \selectp1[74]  = n118 ;
  assign \selectp1[75]  = n119 ;
  assign \selectp1[76]  = n120 ;
  assign \selectp1[77]  = n121 ;
  assign \selectp1[78]  = n122 ;
  assign \selectp1[79]  = n123 ;
  assign \selectp1[80]  = n125 ;
  assign \selectp1[81]  = n126 ;
  assign \selectp1[82]  = n127 ;
  assign \selectp1[83]  = n128 ;
  assign \selectp1[84]  = n129 ;
  assign \selectp1[85]  = n130 ;
  assign \selectp1[86]  = n131 ;
  assign \selectp1[87]  = n132 ;
  assign \selectp1[88]  = n133 ;
  assign \selectp1[89]  = n134 ;
  assign \selectp1[90]  = n135 ;
  assign \selectp1[91]  = n136 ;
  assign \selectp1[92]  = n137 ;
  assign \selectp1[93]  = n138 ;
  assign \selectp1[94]  = n139 ;
  assign \selectp1[95]  = n140 ;
  assign \selectp1[96]  = n142 ;
  assign \selectp1[97]  = n143 ;
  assign \selectp1[98]  = n144 ;
  assign \selectp1[99]  = n145 ;
  assign \selectp1[100]  = n146 ;
  assign \selectp1[101]  = n147 ;
  assign \selectp1[102]  = n148 ;
  assign \selectp1[103]  = n149 ;
  assign \selectp1[104]  = n150 ;
  assign \selectp1[105]  = n151 ;
  assign \selectp1[106]  = n152 ;
  assign \selectp1[107]  = n153 ;
  assign \selectp1[108]  = n154 ;
  assign \selectp1[109]  = n155 ;
  assign \selectp1[110]  = n156 ;
  assign \selectp1[111]  = n157 ;
  assign \selectp1[112]  = n159 ;
  assign \selectp1[113]  = n160 ;
  assign \selectp1[114]  = n161 ;
  assign \selectp1[115]  = n162 ;
  assign \selectp1[116]  = n163 ;
  assign \selectp1[117]  = n164 ;
  assign \selectp1[118]  = n165 ;
  assign \selectp1[119]  = n166 ;
  assign \selectp1[120]  = n167 ;
  assign \selectp1[121]  = n168 ;
  assign \selectp1[122]  = n169 ;
  assign \selectp1[123]  = n170 ;
  assign \selectp1[124]  = n171 ;
  assign \selectp1[125]  = n172 ;
  assign \selectp1[126]  = n173 ;
  assign \selectp1[127]  = n174 ;
  assign \selectp2[0]  = n177 ;
  assign \selectp2[1]  = n178 ;
  assign \selectp2[2]  = n179 ;
  assign \selectp2[3]  = n180 ;
  assign \selectp2[4]  = n181 ;
  assign \selectp2[5]  = n182 ;
  assign \selectp2[6]  = n183 ;
  assign \selectp2[7]  = n184 ;
  assign \selectp2[8]  = n185 ;
  assign \selectp2[9]  = n186 ;
  assign \selectp2[10]  = n187 ;
  assign \selectp2[11]  = n188 ;
  assign \selectp2[12]  = n189 ;
  assign \selectp2[13]  = n190 ;
  assign \selectp2[14]  = n191 ;
  assign \selectp2[15]  = n192 ;
  assign \selectp2[16]  = n194 ;
  assign \selectp2[17]  = n195 ;
  assign \selectp2[18]  = n196 ;
  assign \selectp2[19]  = n197 ;
  assign \selectp2[20]  = n198 ;
  assign \selectp2[21]  = n199 ;
  assign \selectp2[22]  = n200 ;
  assign \selectp2[23]  = n201 ;
  assign \selectp2[24]  = n202 ;
  assign \selectp2[25]  = n203 ;
  assign \selectp2[26]  = n204 ;
  assign \selectp2[27]  = n205 ;
  assign \selectp2[28]  = n206 ;
  assign \selectp2[29]  = n207 ;
  assign \selectp2[30]  = n208 ;
  assign \selectp2[31]  = n209 ;
  assign \selectp2[32]  = n211 ;
  assign \selectp2[33]  = n212 ;
  assign \selectp2[34]  = n213 ;
  assign \selectp2[35]  = n214 ;
  assign \selectp2[36]  = n215 ;
  assign \selectp2[37]  = n216 ;
  assign \selectp2[38]  = n217 ;
  assign \selectp2[39]  = n218 ;
  assign \selectp2[40]  = n219 ;
  assign \selectp2[41]  = n220 ;
  assign \selectp2[42]  = n221 ;
  assign \selectp2[43]  = n222 ;
  assign \selectp2[44]  = n223 ;
  assign \selectp2[45]  = n224 ;
  assign \selectp2[46]  = n225 ;
  assign \selectp2[47]  = n226 ;
  assign \selectp2[48]  = n228 ;
  assign \selectp2[49]  = n229 ;
  assign \selectp2[50]  = n230 ;
  assign \selectp2[51]  = n231 ;
  assign \selectp2[52]  = n232 ;
  assign \selectp2[53]  = n233 ;
  assign \selectp2[54]  = n234 ;
  assign \selectp2[55]  = n235 ;
  assign \selectp2[56]  = n236 ;
  assign \selectp2[57]  = n237 ;
  assign \selectp2[58]  = n238 ;
  assign \selectp2[59]  = n239 ;
  assign \selectp2[60]  = n240 ;
  assign \selectp2[61]  = n241 ;
  assign \selectp2[62]  = n242 ;
  assign \selectp2[63]  = n243 ;
  assign \selectp2[64]  = n246 ;
  assign \selectp2[65]  = n247 ;
  assign \selectp2[66]  = n248 ;
  assign \selectp2[67]  = n249 ;
  assign \selectp2[68]  = n250 ;
  assign \selectp2[69]  = n251 ;
  assign \selectp2[70]  = n252 ;
  assign \selectp2[71]  = n253 ;
  assign \selectp2[72]  = n254 ;
  assign \selectp2[73]  = n255 ;
  assign \selectp2[74]  = n256 ;
  assign \selectp2[75]  = n257 ;
  assign \selectp2[76]  = n258 ;
  assign \selectp2[77]  = n259 ;
  assign \selectp2[78]  = n260 ;
  assign \selectp2[79]  = n261 ;
  assign \selectp2[80]  = n263 ;
  assign \selectp2[81]  = n264 ;
  assign \selectp2[82]  = n265 ;
  assign \selectp2[83]  = n266 ;
  assign \selectp2[84]  = n267 ;
  assign \selectp2[85]  = n268 ;
  assign \selectp2[86]  = n269 ;
  assign \selectp2[87]  = n270 ;
  assign \selectp2[88]  = n271 ;
  assign \selectp2[89]  = n272 ;
  assign \selectp2[90]  = n273 ;
  assign \selectp2[91]  = n274 ;
  assign \selectp2[92]  = n275 ;
  assign \selectp2[93]  = n276 ;
  assign \selectp2[94]  = n277 ;
  assign \selectp2[95]  = n278 ;
  assign \selectp2[96]  = n280 ;
  assign \selectp2[97]  = n281 ;
  assign \selectp2[98]  = n282 ;
  assign \selectp2[99]  = n283 ;
  assign \selectp2[100]  = n284 ;
  assign \selectp2[101]  = n285 ;
  assign \selectp2[102]  = n286 ;
  assign \selectp2[103]  = n287 ;
  assign \selectp2[104]  = n288 ;
  assign \selectp2[105]  = n289 ;
  assign \selectp2[106]  = n290 ;
  assign \selectp2[107]  = n291 ;
  assign \selectp2[108]  = n292 ;
  assign \selectp2[109]  = n293 ;
  assign \selectp2[110]  = n294 ;
  assign \selectp2[111]  = n295 ;
  assign \selectp2[112]  = n297 ;
  assign \selectp2[113]  = n298 ;
  assign \selectp2[114]  = n299 ;
  assign \selectp2[115]  = n300 ;
  assign \selectp2[116]  = n301 ;
  assign \selectp2[117]  = n302 ;
  assign \selectp2[118]  = n303 ;
  assign \selectp2[119]  = n304 ;
  assign \selectp2[120]  = n305 ;
  assign \selectp2[121]  = n306 ;
  assign \selectp2[122]  = n307 ;
  assign \selectp2[123]  = n308 ;
  assign \selectp2[124]  = n309 ;
  assign \selectp2[125]  = n310 ;
  assign \selectp2[126]  = n311 ;
  assign \selectp2[127]  = n312 ;
endmodule
