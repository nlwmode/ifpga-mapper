module top (\DataOut_pad_o[0]_pad , \DataOut_pad_o[1]_pad , \DataOut_pad_o[2]_pad , \DataOut_pad_o[3]_pad , \DataOut_pad_o[4]_pad , \DataOut_pad_o[5]_pad , \DataOut_pad_o[6]_pad , \DataOut_pad_o[7]_pad , \LineState_pad_i[0]_pad , \LineState_pad_i[1]_pad , \LineState_r_reg[0]/P0001 , \LineState_r_reg[1]/P0001 , \OpMode_pad_o[1]_pad , RxActive_pad_i_pad, RxError_pad_i_pad, RxValid_pad_i_pad, TermSel_pad_o_pad, TxReady_pad_i_pad, TxValid_pad_o_pad, VControl_Load_pad_o_pad, XcvSelect_pad_o_pad, \dma_ack_i[0]_pad , \dma_ack_i[1]_pad , \dma_ack_i[2]_pad , \dma_ack_i[3]_pad , \dma_req_o[0]_pad , \dma_req_o[1]_pad , \dma_req_o[2]_pad , \dma_req_o[3]_pad , resume_req_i_pad, \resume_req_r_reg/P0001 , rst_i_pad, \sram_data_i[0]_pad , \sram_data_i[10]_pad , \sram_data_i[11]_pad , \sram_data_i[12]_pad , \sram_data_i[13]_pad , \sram_data_i[14]_pad , \sram_data_i[15]_pad , \sram_data_i[16]_pad , \sram_data_i[17]_pad , \sram_data_i[18]_pad , \sram_data_i[19]_pad , \sram_data_i[1]_pad , \sram_data_i[20]_pad , \sram_data_i[21]_pad , \sram_data_i[22]_pad , \sram_data_i[23]_pad , \sram_data_i[24]_pad , \sram_data_i[25]_pad , \sram_data_i[26]_pad , \sram_data_i[27]_pad , \sram_data_i[28]_pad , \sram_data_i[29]_pad , \sram_data_i[2]_pad , \sram_data_i[30]_pad , \sram_data_i[31]_pad , \sram_data_i[3]_pad , \sram_data_i[4]_pad , \sram_data_i[5]_pad , \sram_data_i[6]_pad , \sram_data_i[7]_pad , \sram_data_i[8]_pad , \sram_data_i[9]_pad , susp_o_pad, \suspend_clr_wr_reg/P0001 , \u0_drive_k_r_reg/P0001 , \u0_rx_active_reg/P0001 , \u0_rx_data_reg[0]/P0001 , \u0_rx_data_reg[1]/P0001 , \u0_rx_data_reg[2]/P0001 , \u0_rx_data_reg[3]/P0001 , \u0_rx_data_reg[4]/P0001 , \u0_rx_data_reg[5]/P0001 , \u0_rx_data_reg[6]/P0001 , \u0_rx_data_reg[7]/P0001 , \u0_rx_err_reg/P0001 , \u0_rx_valid_reg/P0001 , \u0_tx_ready_reg/NET0131 , \u0_u0_T1_gt_2_5_uS_reg/P0001 , \u0_u0_T1_gt_3_0_mS_reg/P0001 , \u0_u0_T1_gt_5_0_mS_reg/P0001 , \u0_u0_T1_st_3_0_mS_reg/P0001 , \u0_u0_T2_gt_100_uS_reg/P0001 , \u0_u0_T2_gt_1_0_mS_reg/P0001 , \u0_u0_T2_wakeup_reg/P0001 , \u0_u0_chirp_cnt_is_6_reg/P0001 , \u0_u0_chirp_cnt_reg[0]/P0001 , \u0_u0_chirp_cnt_reg[1]/P0001 , \u0_u0_chirp_cnt_reg[2]/P0001 , \u0_u0_drive_k_reg/P0001 , \u0_u0_idle_cnt1_clr_reg/P0001 , \u0_u0_idle_cnt1_next_reg[0]/P0001 , \u0_u0_idle_cnt1_next_reg[1]/P0001 , \u0_u0_idle_cnt1_next_reg[2]/P0001 , \u0_u0_idle_cnt1_next_reg[3]/P0001 , \u0_u0_idle_cnt1_next_reg[4]/P0001 , \u0_u0_idle_cnt1_next_reg[5]/P0001 , \u0_u0_idle_cnt1_next_reg[6]/P0001 , \u0_u0_idle_cnt1_next_reg[7]/P0001 , \u0_u0_idle_cnt1_reg[0]/P0001 , \u0_u0_idle_cnt1_reg[1]/P0001 , \u0_u0_idle_cnt1_reg[2]/P0001 , \u0_u0_idle_cnt1_reg[3]/P0001 , \u0_u0_idle_cnt1_reg[4]/P0001 , \u0_u0_idle_cnt1_reg[5]/P0001 , \u0_u0_idle_cnt1_reg[6]/P0001 , \u0_u0_idle_cnt1_reg[7]/P0001 , \u0_u0_idle_long_reg/P0001 , \u0_u0_ls_idle_r_reg/P0001 , \u0_u0_ls_j_r_reg/P0001 , \u0_u0_ls_k_r_reg/P0001 , \u0_u0_ls_se0_r_reg/P0001 , \u0_u0_me_cnt_100_ms_reg/P0001 , \u0_u0_me_cnt_reg[0]/P0001 , \u0_u0_me_cnt_reg[1]/P0001 , \u0_u0_me_cnt_reg[2]/P0001 , \u0_u0_me_cnt_reg[3]/P0001 , \u0_u0_me_cnt_reg[4]/P0001 , \u0_u0_me_cnt_reg[5]/P0001 , \u0_u0_me_cnt_reg[6]/P0001 , \u0_u0_me_cnt_reg[7]/P0001 , \u0_u0_me_ps2_0_5_ms_reg/P0001 , \u0_u0_me_ps2_reg[0]/P0001 , \u0_u0_me_ps2_reg[1]/P0001 , \u0_u0_me_ps2_reg[2]/P0001 , \u0_u0_me_ps2_reg[3]/P0001 , \u0_u0_me_ps2_reg[4]/P0001 , \u0_u0_me_ps2_reg[5]/P0001 , \u0_u0_me_ps2_reg[6]/P0001 , \u0_u0_me_ps2_reg[7]/P0001 , \u0_u0_me_ps_2_5_us_reg/P0001 , \u0_u0_me_ps_reg[0]/P0001 , \u0_u0_me_ps_reg[1]/P0001 , \u0_u0_me_ps_reg[2]/P0001 , \u0_u0_me_ps_reg[3]/P0001 , \u0_u0_me_ps_reg[4]/P0001 , \u0_u0_me_ps_reg[5]/P0001 , \u0_u0_me_ps_reg[6]/P0001 , \u0_u0_me_ps_reg[7]/P0001 , \u0_u0_mode_hs_reg/P0001 , \u0_u0_ps_cnt_clr_reg/P0001 , \u0_u0_ps_cnt_reg[0]/P0001 , \u0_u0_ps_cnt_reg[1]/P0001 , \u0_u0_ps_cnt_reg[2]/P0001 , \u0_u0_ps_cnt_reg[3]/P0001 , \u0_u0_resume_req_s_reg/P0001 , \u0_u0_state_reg[0]/NET0131 , \u0_u0_state_reg[10]/P0001 , \u0_u0_state_reg[11]/NET0131 , \u0_u0_state_reg[12]/NET0131 , \u0_u0_state_reg[13]/NET0131 , \u0_u0_state_reg[14]/P0001 , \u0_u0_state_reg[1]/P0001 , \u0_u0_state_reg[2]/NET0131 , \u0_u0_state_reg[3]/P0001 , \u0_u0_state_reg[4]/NET0131 , \u0_u0_state_reg[5]/P0001 , \u0_u0_state_reg[6]/NET0131 , \u0_u0_state_reg[7]/NET0131 , \u0_u0_state_reg[8]/NET0131 , \u0_u0_state_reg[9]/P0001 , \u0_u0_usb_attached_reg/P0001 , \u0_u0_usb_suspend_reg/P0001 , \u1_clr_sof_time_reg/P0001 , \u1_frame_no_r_reg[0]/P0001 , \u1_frame_no_r_reg[10]/P0001 , \u1_frame_no_r_reg[1]/P0001 , \u1_frame_no_r_reg[2]/P0001 , \u1_frame_no_r_reg[3]/P0001 , \u1_frame_no_r_reg[4]/P0001 , \u1_frame_no_r_reg[5]/P0001 , \u1_frame_no_r_reg[6]/P0001 , \u1_frame_no_r_reg[7]/P0001 , \u1_frame_no_r_reg[8]/P0001 , \u1_frame_no_r_reg[9]/P0001 , \u1_frame_no_same_reg/P0001 , \u1_hms_clk_reg/P0001 , \u1_hms_cnt_reg[0]/P0001 , \u1_hms_cnt_reg[1]/P0001 , \u1_hms_cnt_reg[2]/P0001 , \u1_hms_cnt_reg[3]/P0001 , \u1_hms_cnt_reg[4]/P0001 , \u1_mfm_cnt_reg[0]/P0001 , \u1_mfm_cnt_reg[1]/P0001 , \u1_mfm_cnt_reg[2]/P0001 , \u1_mfm_cnt_reg[3]/P0001 , \u1_sof_time_reg[0]/P0001 , \u1_sof_time_reg[10]/P0001 , \u1_sof_time_reg[11]/P0001 , \u1_sof_time_reg[1]/P0001 , \u1_sof_time_reg[2]/P0001 , \u1_sof_time_reg[3]/P0001 , \u1_sof_time_reg[4]/P0001 , \u1_sof_time_reg[5]/P0001 , \u1_sof_time_reg[6]/P0001 , \u1_sof_time_reg[7]/P0001 , \u1_sof_time_reg[8]/P0001 , \u1_sof_time_reg[9]/P0001 , \u1_u0_crc16_sum_reg[0]/P0001 , \u1_u0_crc16_sum_reg[10]/P0001 , \u1_u0_crc16_sum_reg[11]/P0001 , \u1_u0_crc16_sum_reg[12]/P0001 , \u1_u0_crc16_sum_reg[13]/P0001 , \u1_u0_crc16_sum_reg[14]/P0001 , \u1_u0_crc16_sum_reg[15]/P0001 , \u1_u0_crc16_sum_reg[1]/P0001 , \u1_u0_crc16_sum_reg[2]/P0001 , \u1_u0_crc16_sum_reg[3]/P0001 , \u1_u0_crc16_sum_reg[4]/P0001 , \u1_u0_crc16_sum_reg[5]/P0001 , \u1_u0_crc16_sum_reg[6]/P0001 , \u1_u0_crc16_sum_reg[7]/P0001 , \u1_u0_crc16_sum_reg[8]/P0001 , \u1_u0_crc16_sum_reg[9]/P0001 , \u1_u0_data_valid0_reg/P0001 , \u1_u0_pid_reg[0]/NET0131 , \u1_u0_pid_reg[1]/NET0131 , \u1_u0_pid_reg[2]/NET0131 , \u1_u0_pid_reg[3]/NET0131 , \u1_u0_pid_reg[4]/P0001 , \u1_u0_pid_reg[5]/P0001 , \u1_u0_pid_reg[6]/P0001 , \u1_u0_pid_reg[7]/P0001 , \u1_u0_rx_active_r_reg/P0001 , \u1_u0_rxv1_reg/P0001 , \u1_u0_rxv2_reg/P0001 , \u1_u0_state_reg[0]/P0001 , \u1_u0_state_reg[1]/P0001 , \u1_u0_state_reg[2]/P0001 , \u1_u0_state_reg[3]/P0001 , \u1_u0_token0_reg[0]/NET0131 , \u1_u0_token0_reg[1]/P0001 , \u1_u0_token0_reg[2]/NET0131 , \u1_u0_token0_reg[3]/NET0131 , \u1_u0_token0_reg[4]/P0001 , \u1_u0_token0_reg[5]/NET0131 , \u1_u0_token0_reg[6]/P0001 , \u1_u0_token0_reg[7]/P0001 , \u1_u0_token1_reg[0]/P0001 , \u1_u0_token1_reg[1]/P0001 , \u1_u0_token1_reg[2]/P0001 , \u1_u0_token1_reg[3]/P0001 , \u1_u0_token1_reg[4]/P0001 , \u1_u0_token1_reg[5]/P0001 , \u1_u0_token1_reg[6]/P0001 , \u1_u0_token1_reg[7]/P0001 , \u1_u0_token_valid_r1_reg/P0001 , \u1_u0_token_valid_str1_reg/P0001 , \u1_u1_crc16_reg[0]/P0001 , \u1_u1_crc16_reg[10]/P0001 , \u1_u1_crc16_reg[11]/P0001 , \u1_u1_crc16_reg[12]/P0001 , \u1_u1_crc16_reg[13]/P0001 , \u1_u1_crc16_reg[14]/P0001 , \u1_u1_crc16_reg[15]/P0001 , \u1_u1_crc16_reg[1]/P0001 , \u1_u1_crc16_reg[2]/P0001 , \u1_u1_crc16_reg[3]/P0001 , \u1_u1_crc16_reg[4]/P0001 , \u1_u1_crc16_reg[5]/P0001 , \u1_u1_crc16_reg[6]/P0001 , \u1_u1_crc16_reg[7]/P0001 , \u1_u1_crc16_reg[8]/P0001 , \u1_u1_crc16_reg[9]/P0001 , \u1_u1_send_data_r2_reg/P0001 , \u1_u1_send_data_r_reg/P0001 , \u1_u1_send_token_r_reg/P0001 , \u1_u1_send_zero_length_r_reg/P0001 , \u1_u1_state_reg[0]/NET0131 , \u1_u1_state_reg[1]/NET0131 , \u1_u1_state_reg[2]/NET0131 , \u1_u1_state_reg[3]/NET0131 , \u1_u1_state_reg[4]/NET0131 , \u1_u1_tx_first_r_reg/P0001 , \u1_u1_tx_valid_r_reg/NET0131 , \u1_u1_zero_length_r_reg/P0001 , \u1_u2_adr_cb_reg[0]/NET0131 , \u1_u2_adr_cb_reg[1]/NET0131 , \u1_u2_adr_cb_reg[2]/NET0131 , \u1_u2_adr_cw_reg[0]/NET0131 , \u1_u2_adr_cw_reg[10]/P0001 , \u1_u2_adr_cw_reg[11]/P0001 , \u1_u2_adr_cw_reg[12]/P0001 , \u1_u2_adr_cw_reg[13]/P0001 , \u1_u2_adr_cw_reg[14]/P0001 , \u1_u2_adr_cw_reg[1]/P0001 , \u1_u2_adr_cw_reg[2]/P0001 , \u1_u2_adr_cw_reg[3]/NET0131 , \u1_u2_adr_cw_reg[4]/P0001 , \u1_u2_adr_cw_reg[5]/NET0131 , \u1_u2_adr_cw_reg[6]/NET0131 , \u1_u2_adr_cw_reg[7]/NET0131 , \u1_u2_adr_cw_reg[8]/P0001 , \u1_u2_adr_cw_reg[9]/NET0131 , \u1_u2_dout_r_reg[0]/P0001 , \u1_u2_dout_r_reg[10]/P0001 , \u1_u2_dout_r_reg[11]/P0001 , \u1_u2_dout_r_reg[12]/P0001 , \u1_u2_dout_r_reg[13]/P0001 , \u1_u2_dout_r_reg[14]/P0001 , \u1_u2_dout_r_reg[15]/P0001 , \u1_u2_dout_r_reg[16]/P0001 , \u1_u2_dout_r_reg[17]/P0001 , \u1_u2_dout_r_reg[18]/P0001 , \u1_u2_dout_r_reg[19]/P0001 , \u1_u2_dout_r_reg[1]/P0001 , \u1_u2_dout_r_reg[20]/P0001 , \u1_u2_dout_r_reg[21]/P0001 , \u1_u2_dout_r_reg[22]/P0001 , \u1_u2_dout_r_reg[23]/P0001 , \u1_u2_dout_r_reg[24]/P0001 , \u1_u2_dout_r_reg[25]/P0001 , \u1_u2_dout_r_reg[26]/P0001 , \u1_u2_dout_r_reg[27]/P0001 , \u1_u2_dout_r_reg[28]/P0001 , \u1_u2_dout_r_reg[29]/P0001 , \u1_u2_dout_r_reg[2]/P0001 , \u1_u2_dout_r_reg[30]/P0001 , \u1_u2_dout_r_reg[31]/P0001 , \u1_u2_dout_r_reg[3]/P0001 , \u1_u2_dout_r_reg[4]/P0001 , \u1_u2_dout_r_reg[5]/P0001 , \u1_u2_dout_r_reg[6]/P0001 , \u1_u2_dout_r_reg[7]/P0001 , \u1_u2_dout_r_reg[8]/P0001 , \u1_u2_dout_r_reg[9]/P0001 , \u1_u2_dtmp_r_reg[0]/P0001 , \u1_u2_dtmp_r_reg[10]/P0001 , \u1_u2_dtmp_r_reg[11]/P0001 , \u1_u2_dtmp_r_reg[12]/P0001 , \u1_u2_dtmp_r_reg[13]/P0001 , \u1_u2_dtmp_r_reg[14]/P0001 , \u1_u2_dtmp_r_reg[15]/P0001 , \u1_u2_dtmp_r_reg[16]/P0001 , \u1_u2_dtmp_r_reg[17]/P0001 , \u1_u2_dtmp_r_reg[18]/P0001 , \u1_u2_dtmp_r_reg[19]/P0001 , \u1_u2_dtmp_r_reg[1]/P0001 , \u1_u2_dtmp_r_reg[20]/P0001 , \u1_u2_dtmp_r_reg[21]/P0001 , \u1_u2_dtmp_r_reg[22]/P0001 , \u1_u2_dtmp_r_reg[23]/P0001 , \u1_u2_dtmp_r_reg[24]/P0001 , \u1_u2_dtmp_r_reg[25]/P0001 , \u1_u2_dtmp_r_reg[26]/P0001 , \u1_u2_dtmp_r_reg[27]/P0001 , \u1_u2_dtmp_r_reg[28]/P0001 , \u1_u2_dtmp_r_reg[29]/P0001 , \u1_u2_dtmp_r_reg[2]/P0001 , \u1_u2_dtmp_r_reg[30]/P0001 , \u1_u2_dtmp_r_reg[31]/P0001 , \u1_u2_dtmp_r_reg[3]/P0001 , \u1_u2_dtmp_r_reg[4]/P0001 , \u1_u2_dtmp_r_reg[5]/P0001 , \u1_u2_dtmp_r_reg[6]/P0001 , \u1_u2_dtmp_r_reg[7]/P0001 , \u1_u2_dtmp_r_reg[8]/P0001 , \u1_u2_dtmp_r_reg[9]/P0001 , \u1_u2_dtmp_sel_r_reg/P0001 , \u1_u2_idma_done_reg/P0001 , \u1_u2_last_buf_adr_reg[0]/P0001 , \u1_u2_last_buf_adr_reg[10]/P0001 , \u1_u2_last_buf_adr_reg[11]/P0001 , \u1_u2_last_buf_adr_reg[12]/P0001 , \u1_u2_last_buf_adr_reg[13]/P0001 , \u1_u2_last_buf_adr_reg[14]/P0001 , \u1_u2_last_buf_adr_reg[1]/P0001 , \u1_u2_last_buf_adr_reg[2]/P0001 , \u1_u2_last_buf_adr_reg[3]/P0001 , \u1_u2_last_buf_adr_reg[4]/P0001 , \u1_u2_last_buf_adr_reg[5]/P0001 , \u1_u2_last_buf_adr_reg[6]/P0001 , \u1_u2_last_buf_adr_reg[7]/P0001 , \u1_u2_last_buf_adr_reg[8]/P0001 , \u1_u2_last_buf_adr_reg[9]/P0001 , \u1_u2_mack_r_reg/P0001 , \u1_u2_mwe_reg/P0001 , \u1_u2_rd_buf0_reg[0]/NET0131 , \u1_u2_rd_buf0_reg[10]/NET0131 , \u1_u2_rd_buf0_reg[11]/NET0131 , \u1_u2_rd_buf0_reg[12]/P0001 , \u1_u2_rd_buf0_reg[13]/P0001 , \u1_u2_rd_buf0_reg[14]/P0001 , \u1_u2_rd_buf0_reg[15]/P0001 , \u1_u2_rd_buf0_reg[16]/NET0131 , \u1_u2_rd_buf0_reg[17]/NET0131 , \u1_u2_rd_buf0_reg[18]/NET0131 , \u1_u2_rd_buf0_reg[19]/NET0131 , \u1_u2_rd_buf0_reg[1]/NET0131 , \u1_u2_rd_buf0_reg[20]/P0001 , \u1_u2_rd_buf0_reg[21]/P0001 , \u1_u2_rd_buf0_reg[22]/P0001 , \u1_u2_rd_buf0_reg[23]/P0001 , \u1_u2_rd_buf0_reg[24]/NET0131 , \u1_u2_rd_buf0_reg[25]/NET0131 , \u1_u2_rd_buf0_reg[26]/NET0131 , \u1_u2_rd_buf0_reg[27]/NET0131 , \u1_u2_rd_buf0_reg[28]/P0001 , \u1_u2_rd_buf0_reg[29]/P0001 , \u1_u2_rd_buf0_reg[2]/NET0131 , \u1_u2_rd_buf0_reg[30]/P0001 , \u1_u2_rd_buf0_reg[31]/P0001 , \u1_u2_rd_buf0_reg[3]/NET0131 , \u1_u2_rd_buf0_reg[4]/P0001 , \u1_u2_rd_buf0_reg[5]/P0001 , \u1_u2_rd_buf0_reg[6]/P0001 , \u1_u2_rd_buf0_reg[7]/P0001 , \u1_u2_rd_buf0_reg[8]/NET0131 , \u1_u2_rd_buf0_reg[9]/NET0131 , \u1_u2_rd_buf1_reg[0]/NET0131 , \u1_u2_rd_buf1_reg[10]/NET0131 , \u1_u2_rd_buf1_reg[11]/NET0131 , \u1_u2_rd_buf1_reg[12]/P0001 , \u1_u2_rd_buf1_reg[13]/P0001 , \u1_u2_rd_buf1_reg[14]/P0001 , \u1_u2_rd_buf1_reg[15]/P0001 , \u1_u2_rd_buf1_reg[16]/NET0131 , \u1_u2_rd_buf1_reg[17]/NET0131 , \u1_u2_rd_buf1_reg[18]/NET0131 , \u1_u2_rd_buf1_reg[19]/NET0131 , \u1_u2_rd_buf1_reg[1]/NET0131 , \u1_u2_rd_buf1_reg[20]/P0001 , \u1_u2_rd_buf1_reg[21]/P0001 , \u1_u2_rd_buf1_reg[22]/P0001 , \u1_u2_rd_buf1_reg[23]/P0001 , \u1_u2_rd_buf1_reg[24]/NET0131 , \u1_u2_rd_buf1_reg[25]/NET0131 , \u1_u2_rd_buf1_reg[26]/NET0131 , \u1_u2_rd_buf1_reg[27]/NET0131 , \u1_u2_rd_buf1_reg[28]/P0001 , \u1_u2_rd_buf1_reg[29]/P0001 , \u1_u2_rd_buf1_reg[2]/NET0131 , \u1_u2_rd_buf1_reg[30]/P0001 , \u1_u2_rd_buf1_reg[31]/P0001 , \u1_u2_rd_buf1_reg[3]/NET0131 , \u1_u2_rd_buf1_reg[4]/P0001 , \u1_u2_rd_buf1_reg[5]/P0001 , \u1_u2_rd_buf1_reg[6]/P0001 , \u1_u2_rd_buf1_reg[7]/P0001 , \u1_u2_rd_buf1_reg[8]/NET0131 , \u1_u2_rd_buf1_reg[9]/NET0131 , \u1_u2_rx_data_done_r2_reg/P0001 , \u1_u2_rx_data_done_r_reg/P0001 , \u1_u2_rx_data_st_r_reg[0]/P0001 , \u1_u2_rx_data_st_r_reg[1]/P0001 , \u1_u2_rx_data_st_r_reg[2]/P0001 , \u1_u2_rx_data_st_r_reg[3]/P0001 , \u1_u2_rx_data_st_r_reg[4]/P0001 , \u1_u2_rx_data_st_r_reg[5]/P0001 , \u1_u2_rx_data_st_r_reg[6]/P0001 , \u1_u2_rx_data_st_r_reg[7]/P0001 , \u1_u2_rx_data_valid_r_reg/NET0131 , \u1_u2_rx_dma_en_r_reg/P0001 , \u1_u2_send_data_r_reg/NET0131 , \u1_u2_sizd_c_reg[0]/P0001 , \u1_u2_sizd_c_reg[10]/P0001 , \u1_u2_sizd_c_reg[11]/P0001 , \u1_u2_sizd_c_reg[12]/P0001 , \u1_u2_sizd_c_reg[13]/P0001 , \u1_u2_sizd_c_reg[1]/P0001 , \u1_u2_sizd_c_reg[2]/P0001 , \u1_u2_sizd_c_reg[3]/P0001 , \u1_u2_sizd_c_reg[4]/P0001 , \u1_u2_sizd_c_reg[5]/P0001 , \u1_u2_sizd_c_reg[6]/P0001 , \u1_u2_sizd_c_reg[7]/P0001 , \u1_u2_sizd_c_reg[8]/P0001 , \u1_u2_sizd_c_reg[9]/P0001 , \u1_u2_sizd_is_zero_reg/P0001 , \u1_u2_sizu_c_reg[0]/P0001 , \u1_u2_sizu_c_reg[10]/P0001 , \u1_u2_sizu_c_reg[1]/P0001 , \u1_u2_sizu_c_reg[2]/P0001 , \u1_u2_sizu_c_reg[3]/P0001 , \u1_u2_sizu_c_reg[4]/P0001 , \u1_u2_sizu_c_reg[5]/P0001 , \u1_u2_sizu_c_reg[6]/P0001 , \u1_u2_sizu_c_reg[7]/P0001 , \u1_u2_sizu_c_reg[8]/NET0131 , \u1_u2_sizu_c_reg[9]/P0001 , \u1_u2_state_reg[0]/P0001 , \u1_u2_state_reg[1]/NET0131 , \u1_u2_state_reg[2]/NET0131 , \u1_u2_state_reg[3]/NET0131 , \u1_u2_state_reg[4]/NET0131 , \u1_u2_state_reg[5]/NET0131 , \u1_u2_state_reg[6]/NET0131 , \u1_u2_state_reg[7]/NET0131 , \u1_u2_tx_dma_en_r_reg/P0001 , \u1_u2_word_done_r_reg/P0001 , \u1_u2_word_done_reg/NET0131 , \u1_u2_wr_done_reg/P0001 , \u1_u2_wr_last_reg/P0001 , \u1_u3_abort_reg/P0001 , \u1_u3_adr_r_reg[0]/P0001 , \u1_u3_adr_r_reg[10]/P0001 , \u1_u3_adr_r_reg[11]/P0001 , \u1_u3_adr_r_reg[12]/P0001 , \u1_u3_adr_r_reg[13]/P0001 , \u1_u3_adr_r_reg[14]/P0001 , \u1_u3_adr_r_reg[15]/P0001 , \u1_u3_adr_r_reg[16]/P0001 , \u1_u3_adr_r_reg[1]/P0001 , \u1_u3_adr_r_reg[2]/P0001 , \u1_u3_adr_r_reg[3]/P0001 , \u1_u3_adr_r_reg[4]/P0001 , \u1_u3_adr_r_reg[5]/P0001 , \u1_u3_adr_r_reg[6]/P0001 , \u1_u3_adr_r_reg[7]/P0001 , \u1_u3_adr_r_reg[8]/P0001 , \u1_u3_adr_r_reg[9]/P0001 , \u1_u3_adr_reg[0]/P0001 , \u1_u3_adr_reg[10]/P0001 , \u1_u3_adr_reg[11]/P0001 , \u1_u3_adr_reg[12]/P0001 , \u1_u3_adr_reg[13]/P0001 , \u1_u3_adr_reg[14]/P0001 , \u1_u3_adr_reg[15]/P0001 , \u1_u3_adr_reg[16]/P0001 , \u1_u3_adr_reg[1]/P0001 , \u1_u3_adr_reg[2]/P0001 , \u1_u3_adr_reg[3]/P0001 , \u1_u3_adr_reg[4]/P0001 , \u1_u3_adr_reg[5]/P0001 , \u1_u3_adr_reg[6]/P0001 , \u1_u3_adr_reg[7]/P0001 , \u1_u3_adr_reg[8]/P0001 , \u1_u3_adr_reg[9]/P0001 , \u1_u3_buf0_na_reg/NET0131 , \u1_u3_buf0_not_aloc_reg/P0001 , \u1_u3_buf0_rl_reg/P0001 , \u1_u3_buf0_set_reg/P0001 , \u1_u3_buf0_st_max_reg/P0001 , \u1_u3_buf1_na_reg/NET0131 , \u1_u3_buf1_not_aloc_reg/P0001 , \u1_u3_buf1_set_reg/P0001 , \u1_u3_buf1_st_max_reg/P0001 , \u1_u3_buffer_done_reg/P0001 , \u1_u3_buffer_empty_reg/P0001 , \u1_u3_buffer_full_reg/P0001 , \u1_u3_buffer_overflow_reg/P0001 , \u1_u3_idin_reg[0]/P0001 , \u1_u3_idin_reg[10]/P0001 , \u1_u3_idin_reg[11]/P0001 , \u1_u3_idin_reg[12]/P0001 , \u1_u3_idin_reg[13]/P0001 , \u1_u3_idin_reg[14]/P0001 , \u1_u3_idin_reg[15]/P0001 , \u1_u3_idin_reg[16]/P0001 , \u1_u3_idin_reg[17]/P0001 , \u1_u3_idin_reg[18]/P0001 , \u1_u3_idin_reg[19]/P0001 , \u1_u3_idin_reg[1]/P0001 , \u1_u3_idin_reg[20]/P0001 , \u1_u3_idin_reg[21]/P0001 , \u1_u3_idin_reg[22]/P0001 , \u1_u3_idin_reg[23]/P0001 , \u1_u3_idin_reg[24]/P0001 , \u1_u3_idin_reg[25]/P0001 , \u1_u3_idin_reg[26]/P0001 , \u1_u3_idin_reg[27]/P0001 , \u1_u3_idin_reg[28]/P0001 , \u1_u3_idin_reg[29]/P0001 , \u1_u3_idin_reg[2]/P0001 , \u1_u3_idin_reg[30]/P0001 , \u1_u3_idin_reg[31]/P0001 , \u1_u3_idin_reg[3]/P0001 , \u1_u3_idin_reg[4]/P0001 , \u1_u3_idin_reg[5]/P0001 , \u1_u3_idin_reg[6]/P0001 , \u1_u3_idin_reg[7]/P0001 , \u1_u3_idin_reg[8]/P0001 , \u1_u3_idin_reg[9]/P0001 , \u1_u3_in_token_reg/NET0131 , \u1_u3_int_seqerr_set_reg/P0001 , \u1_u3_int_upid_set_reg/P0001 , \u1_u3_match_r_reg/P0001 , \u1_u3_new_size_reg[0]/P0001 , \u1_u3_new_size_reg[10]/P0001 , \u1_u3_new_size_reg[11]/P0001 , \u1_u3_new_size_reg[12]/P0001 , \u1_u3_new_size_reg[13]/P0001 , \u1_u3_new_size_reg[1]/P0001 , \u1_u3_new_size_reg[2]/P0001 , \u1_u3_new_size_reg[3]/P0001 , \u1_u3_new_size_reg[4]/P0001 , \u1_u3_new_size_reg[5]/P0001 , \u1_u3_new_size_reg[6]/P0001 , \u1_u3_new_size_reg[7]/P0001 , \u1_u3_new_size_reg[8]/P0001 , \u1_u3_new_size_reg[9]/P0001 , \u1_u3_new_sizeb_reg[0]/P0001 , \u1_u3_new_sizeb_reg[10]/P0001 , \u1_u3_new_sizeb_reg[1]/P0001 , \u1_u3_new_sizeb_reg[2]/P0001 , \u1_u3_new_sizeb_reg[3]/P0001 , \u1_u3_new_sizeb_reg[4]/P0001 , \u1_u3_new_sizeb_reg[5]/P0001 , \u1_u3_new_sizeb_reg[6]/P0001 , \u1_u3_new_sizeb_reg[7]/P0001 , \u1_u3_new_sizeb_reg[8]/P0001 , \u1_u3_new_sizeb_reg[9]/P0001 , \u1_u3_next_dpid_reg[0]/P0001 , \u1_u3_next_dpid_reg[1]/P0001 , \u1_u3_no_bufs0_reg/P0001 , \u1_u3_no_bufs1_reg/P0001 , \u1_u3_out_to_small_r_reg/P0001 , \u1_u3_out_to_small_reg/P0001 , \u1_u3_out_token_reg/NET0131 , \u1_u3_pid_IN_r_reg/P0001 , \u1_u3_pid_OUT_r_reg/P0001 , \u1_u3_pid_PING_r_reg/P0001 , \u1_u3_pid_SETUP_r_reg/P0001 , \u1_u3_pid_seq_err_reg/P0001 , \u1_u3_rx_ack_to_clr_reg/P0001 , \u1_u3_rx_ack_to_cnt_reg[0]/P0001 , \u1_u3_rx_ack_to_cnt_reg[1]/P0001 , \u1_u3_rx_ack_to_cnt_reg[2]/P0001 , \u1_u3_rx_ack_to_cnt_reg[3]/P0001 , \u1_u3_rx_ack_to_cnt_reg[4]/P0001 , \u1_u3_rx_ack_to_cnt_reg[5]/P0001 , \u1_u3_rx_ack_to_cnt_reg[6]/P0001 , \u1_u3_rx_ack_to_cnt_reg[7]/P0001 , \u1_u3_rx_ack_to_reg/P0001 , \u1_u3_send_token_reg/P0001 , \u1_u3_setup_token_reg/P0001 , \u1_u3_size_next_r_reg[0]/P0001 , \u1_u3_size_next_r_reg[10]/P0001 , \u1_u3_size_next_r_reg[1]/P0001 , \u1_u3_size_next_r_reg[2]/P0001 , \u1_u3_size_next_r_reg[3]/P0001 , \u1_u3_size_next_r_reg[4]/P0001 , \u1_u3_size_next_r_reg[5]/P0001 , \u1_u3_size_next_r_reg[6]/P0001 , \u1_u3_size_next_r_reg[7]/P0001 , \u1_u3_size_next_r_reg[8]/P0001 , \u1_u3_size_next_r_reg[9]/P0001 , \u1_u3_state_reg[0]/P0001 , \u1_u3_state_reg[1]/P0001 , \u1_u3_state_reg[2]/P0001 , \u1_u3_state_reg[3]/P0001 , \u1_u3_state_reg[4]/P0001 , \u1_u3_state_reg[5]/P0001 , \u1_u3_state_reg[6]/P0001 , \u1_u3_state_reg[7]/P0001 , \u1_u3_state_reg[8]/P0001 , \u1_u3_state_reg[9]/P0001 , \u1_u3_this_dpid_reg[0]/P0001 , \u1_u3_this_dpid_reg[1]/P0001 , \u1_u3_to_large_reg/P0001 , \u1_u3_to_small_reg/P0001 , \u1_u3_token_pid_sel_reg[0]/P0001 , \u1_u3_token_pid_sel_reg[1]/P0001 , \u1_u3_tx_data_to_cnt_reg[0]/P0001 , \u1_u3_tx_data_to_cnt_reg[1]/P0001 , \u1_u3_tx_data_to_cnt_reg[2]/P0001 , \u1_u3_tx_data_to_cnt_reg[3]/P0001 , \u1_u3_tx_data_to_cnt_reg[4]/P0001 , \u1_u3_tx_data_to_cnt_reg[5]/P0001 , \u1_u3_tx_data_to_cnt_reg[6]/P0001 , \u1_u3_tx_data_to_cnt_reg[7]/P0001 , \u1_u3_tx_data_to_reg/P0001 , \u1_u3_uc_bsel_set_reg/P0001 , \u2_wack_r_reg/P0001 , \u4_attach_r1_reg/P0001 , \u4_attach_r_reg/P0001 , \u4_buf0_reg[0]/P0001 , \u4_buf0_reg[10]/P0001 , \u4_buf0_reg[11]/P0001 , \u4_buf0_reg[12]/P0001 , \u4_buf0_reg[13]/P0001 , \u4_buf0_reg[14]/P0001 , \u4_buf0_reg[15]/P0001 , \u4_buf0_reg[16]/P0001 , \u4_buf0_reg[17]/NET0131 , \u4_buf0_reg[18]/P0001 , \u4_buf0_reg[19]/NET0131 , \u4_buf0_reg[1]/P0001 , \u4_buf0_reg[20]/NET0131 , \u4_buf0_reg[21]/NET0131 , \u4_buf0_reg[22]/NET0131 , \u4_buf0_reg[23]/NET0131 , \u4_buf0_reg[24]/NET0131 , \u4_buf0_reg[25]/NET0131 , \u4_buf0_reg[26]/NET0131 , \u4_buf0_reg[27]/P0001 , \u4_buf0_reg[28]/P0001 , \u4_buf0_reg[29]/P0001 , \u4_buf0_reg[2]/P0001 , \u4_buf0_reg[30]/P0001 , \u4_buf0_reg[31]/P0001 , \u4_buf0_reg[3]/P0001 , \u4_buf0_reg[4]/P0001 , \u4_buf0_reg[5]/P0001 , \u4_buf0_reg[6]/P0001 , \u4_buf0_reg[7]/P0001 , \u4_buf0_reg[8]/P0001 , \u4_buf0_reg[9]/P0001 , \u4_buf1_reg[0]/P0001 , \u4_buf1_reg[10]/P0001 , \u4_buf1_reg[11]/P0001 , \u4_buf1_reg[12]/P0001 , \u4_buf1_reg[13]/P0001 , \u4_buf1_reg[14]/P0001 , \u4_buf1_reg[15]/P0001 , \u4_buf1_reg[16]/P0001 , \u4_buf1_reg[17]/NET0131 , \u4_buf1_reg[18]/P0001 , \u4_buf1_reg[19]/NET0131 , \u4_buf1_reg[1]/P0001 , \u4_buf1_reg[20]/NET0131 , \u4_buf1_reg[21]/NET0131 , \u4_buf1_reg[22]/NET0131 , \u4_buf1_reg[23]/NET0131 , \u4_buf1_reg[24]/NET0131 , \u4_buf1_reg[25]/NET0131 , \u4_buf1_reg[26]/NET0131 , \u4_buf1_reg[27]/P0001 , \u4_buf1_reg[28]/P0001 , \u4_buf1_reg[29]/P0001 , \u4_buf1_reg[2]/P0001 , \u4_buf1_reg[30]/P0001 , \u4_buf1_reg[31]/P0001 , \u4_buf1_reg[3]/P0001 , \u4_buf1_reg[4]/P0001 , \u4_buf1_reg[5]/P0001 , \u4_buf1_reg[6]/P0001 , \u4_buf1_reg[7]/P0001 , \u4_buf1_reg[8]/P0001 , \u4_buf1_reg[9]/P0001 , \u4_crc5_err_r_reg/P0001 , \u4_csr_reg[0]/P0001 , \u4_csr_reg[10]/P0001 , \u4_csr_reg[11]/P0001 , \u4_csr_reg[12]/P0001 , \u4_csr_reg[15]/NET0131 , \u4_csr_reg[16]/P0001 , \u4_csr_reg[17]/P0001 , \u4_csr_reg[1]/P0001 , \u4_csr_reg[22]/P0001 , \u4_csr_reg[23]/P0001 , \u4_csr_reg[24]/P0001 , \u4_csr_reg[25]/P0001 , \u4_csr_reg[26]/NET0131 , \u4_csr_reg[27]/NET0131 , \u4_csr_reg[28]/P0001 , \u4_csr_reg[29]/P0001 , \u4_csr_reg[2]/NET0131 , \u4_csr_reg[30]/NET0131 , \u4_csr_reg[31]/P0001 , \u4_csr_reg[3]/P0001 , \u4_csr_reg[4]/NET0131 , \u4_csr_reg[5]/NET0131 , \u4_csr_reg[6]/NET0131 , \u4_csr_reg[7]/P0001 , \u4_csr_reg[8]/P0001 , \u4_csr_reg[9]/NET0131 , \u4_dma_in_buf_sz1_reg/P0001 , \u4_dma_out_buf_avail_reg/P0001 , \u4_dout_reg[0]/P0001 , \u4_dout_reg[10]/P0001 , \u4_dout_reg[11]/P0001 , \u4_dout_reg[12]/P0001 , \u4_dout_reg[13]/P0001 , \u4_dout_reg[14]/P0001 , \u4_dout_reg[15]/P0001 , \u4_dout_reg[16]/P0001 , \u4_dout_reg[17]/P0001 , \u4_dout_reg[18]/P0001 , \u4_dout_reg[19]/P0001 , \u4_dout_reg[1]/P0001 , \u4_dout_reg[20]/P0001 , \u4_dout_reg[21]/P0001 , \u4_dout_reg[22]/P0001 , \u4_dout_reg[23]/P0001 , \u4_dout_reg[24]/P0001 , \u4_dout_reg[25]/P0001 , \u4_dout_reg[26]/P0001 , \u4_dout_reg[27]/P0001 , \u4_dout_reg[28]/P0001 , \u4_dout_reg[29]/P0001 , \u4_dout_reg[2]/P0001 , \u4_dout_reg[30]/P0001 , \u4_dout_reg[31]/P0001 , \u4_dout_reg[3]/P0001 , \u4_dout_reg[4]/P0001 , \u4_dout_reg[5]/P0001 , \u4_dout_reg[6]/P0001 , \u4_dout_reg[7]/P0001 , \u4_dout_reg[8]/P0001 , \u4_dout_reg[9]/P0001 , \u4_funct_adr_reg[0]/P0001 , \u4_funct_adr_reg[1]/P0001 , \u4_funct_adr_reg[2]/P0001 , \u4_funct_adr_reg[3]/P0001 , \u4_funct_adr_reg[4]/P0001 , \u4_funct_adr_reg[5]/P0001 , \u4_funct_adr_reg[6]/P0001 , \u4_int_src_re_reg/P0001 , \u4_int_srca_reg[0]/P0001 , \u4_int_srca_reg[1]/P0001 , \u4_int_srca_reg[2]/P0001 , \u4_int_srca_reg[3]/P0001 , \u4_int_srcb_reg[0]/P0001 , \u4_int_srcb_reg[1]/P0001 , \u4_int_srcb_reg[2]/P0001 , \u4_int_srcb_reg[3]/P0001 , \u4_int_srcb_reg[4]/P0001 , \u4_int_srcb_reg[5]/P0001 , \u4_int_srcb_reg[6]/P0001 , \u4_int_srcb_reg[7]/P0001 , \u4_int_srcb_reg[8]/P0001 , \u4_inta_msk_reg[0]/P0001 , \u4_inta_msk_reg[1]/P0001 , \u4_inta_msk_reg[2]/P0001 , \u4_inta_msk_reg[3]/P0001 , \u4_inta_msk_reg[4]/P0001 , \u4_inta_msk_reg[5]/P0001 , \u4_inta_msk_reg[6]/P0001 , \u4_inta_msk_reg[7]/P0001 , \u4_inta_msk_reg[8]/P0001 , \u4_intb_msk_reg[0]/P0001 , \u4_intb_msk_reg[1]/P0001 , \u4_intb_msk_reg[2]/P0001 , \u4_intb_msk_reg[3]/P0001 , \u4_intb_msk_reg[4]/P0001 , \u4_intb_msk_reg[5]/P0001 , \u4_intb_msk_reg[6]/P0001 , \u4_intb_msk_reg[7]/P0001 , \u4_intb_msk_reg[8]/P0001 , \u4_match_r1_reg/P0001 , \u4_nse_err_r_reg/P0001 , \u4_pid_cs_err_r_reg/P0001 , \u4_rx_err_r_reg/P0001 , \u4_suspend_r1_reg/P0001 , \u4_u0_buf0_orig_m3_reg[0]/P0001 , \u4_u0_buf0_orig_m3_reg[10]/P0001 , \u4_u0_buf0_orig_m3_reg[11]/P0001 , \u4_u0_buf0_orig_m3_reg[1]/P0001 , \u4_u0_buf0_orig_m3_reg[2]/P0001 , \u4_u0_buf0_orig_m3_reg[3]/P0001 , \u4_u0_buf0_orig_m3_reg[4]/P0001 , \u4_u0_buf0_orig_m3_reg[5]/P0001 , \u4_u0_buf0_orig_m3_reg[6]/P0001 , \u4_u0_buf0_orig_m3_reg[7]/P0001 , \u4_u0_buf0_orig_m3_reg[8]/P0001 , \u4_u0_buf0_orig_m3_reg[9]/P0001 , \u4_u0_buf0_orig_reg[0]/P0001 , \u4_u0_buf0_orig_reg[10]/P0001 , \u4_u0_buf0_orig_reg[11]/P0001 , \u4_u0_buf0_orig_reg[12]/P0001 , \u4_u0_buf0_orig_reg[13]/P0001 , \u4_u0_buf0_orig_reg[14]/P0001 , \u4_u0_buf0_orig_reg[15]/P0001 , \u4_u0_buf0_orig_reg[16]/P0001 , \u4_u0_buf0_orig_reg[17]/P0001 , \u4_u0_buf0_orig_reg[18]/P0001 , \u4_u0_buf0_orig_reg[19]/P0001 , \u4_u0_buf0_orig_reg[1]/P0001 , \u4_u0_buf0_orig_reg[20]/P0001 , \u4_u0_buf0_orig_reg[21]/P0001 , \u4_u0_buf0_orig_reg[22]/P0001 , \u4_u0_buf0_orig_reg[23]/P0001 , \u4_u0_buf0_orig_reg[24]/P0001 , \u4_u0_buf0_orig_reg[25]/P0001 , \u4_u0_buf0_orig_reg[26]/P0001 , \u4_u0_buf0_orig_reg[27]/P0001 , \u4_u0_buf0_orig_reg[28]/P0001 , \u4_u0_buf0_orig_reg[29]/NET0131 , \u4_u0_buf0_orig_reg[2]/P0001 , \u4_u0_buf0_orig_reg[30]/NET0131 , \u4_u0_buf0_orig_reg[31]/P0001 , \u4_u0_buf0_orig_reg[3]/P0001 , \u4_u0_buf0_orig_reg[4]/P0001 , \u4_u0_buf0_orig_reg[5]/P0001 , \u4_u0_buf0_orig_reg[6]/P0001 , \u4_u0_buf0_orig_reg[7]/P0001 , \u4_u0_buf0_orig_reg[8]/P0001 , \u4_u0_buf0_orig_reg[9]/P0001 , \u4_u0_buf0_reg[0]/P0001 , \u4_u0_buf0_reg[10]/P0001 , \u4_u0_buf0_reg[11]/P0001 , \u4_u0_buf0_reg[12]/P0001 , \u4_u0_buf0_reg[13]/P0001 , \u4_u0_buf0_reg[14]/P0001 , \u4_u0_buf0_reg[15]/P0001 , \u4_u0_buf0_reg[16]/P0001 , \u4_u0_buf0_reg[17]/P0001 , \u4_u0_buf0_reg[18]/P0001 , \u4_u0_buf0_reg[19]/P0001 , \u4_u0_buf0_reg[1]/P0001 , \u4_u0_buf0_reg[20]/P0001 , \u4_u0_buf0_reg[21]/P0001 , \u4_u0_buf0_reg[22]/P0001 , \u4_u0_buf0_reg[23]/P0001 , \u4_u0_buf0_reg[24]/P0001 , \u4_u0_buf0_reg[25]/P0001 , \u4_u0_buf0_reg[26]/P0001 , \u4_u0_buf0_reg[27]/P0001 , \u4_u0_buf0_reg[28]/P0001 , \u4_u0_buf0_reg[29]/P0001 , \u4_u0_buf0_reg[2]/P0001 , \u4_u0_buf0_reg[30]/P0001 , \u4_u0_buf0_reg[31]/P0001 , \u4_u0_buf0_reg[3]/P0001 , \u4_u0_buf0_reg[4]/P0001 , \u4_u0_buf0_reg[5]/P0001 , \u4_u0_buf0_reg[6]/P0001 , \u4_u0_buf0_reg[7]/P0001 , \u4_u0_buf0_reg[8]/P0001 , \u4_u0_buf0_reg[9]/P0001 , \u4_u0_buf1_reg[0]/P0001 , \u4_u0_buf1_reg[10]/P0001 , \u4_u0_buf1_reg[11]/P0001 , \u4_u0_buf1_reg[12]/P0001 , \u4_u0_buf1_reg[13]/P0001 , \u4_u0_buf1_reg[14]/P0001 , \u4_u0_buf1_reg[15]/P0001 , \u4_u0_buf1_reg[16]/P0001 , \u4_u0_buf1_reg[17]/P0001 , \u4_u0_buf1_reg[18]/P0001 , \u4_u0_buf1_reg[19]/P0001 , \u4_u0_buf1_reg[1]/P0001 , \u4_u0_buf1_reg[20]/P0001 , \u4_u0_buf1_reg[21]/P0001 , \u4_u0_buf1_reg[22]/P0001 , \u4_u0_buf1_reg[23]/P0001 , \u4_u0_buf1_reg[24]/P0001 , \u4_u0_buf1_reg[25]/P0001 , \u4_u0_buf1_reg[26]/P0001 , \u4_u0_buf1_reg[27]/P0001 , \u4_u0_buf1_reg[28]/P0001 , \u4_u0_buf1_reg[29]/P0001 , \u4_u0_buf1_reg[2]/P0001 , \u4_u0_buf1_reg[30]/P0001 , \u4_u0_buf1_reg[31]/P0001 , \u4_u0_buf1_reg[3]/P0001 , \u4_u0_buf1_reg[4]/P0001 , \u4_u0_buf1_reg[5]/P0001 , \u4_u0_buf1_reg[6]/P0001 , \u4_u0_buf1_reg[7]/P0001 , \u4_u0_buf1_reg[8]/P0001 , \u4_u0_buf1_reg[9]/P0001 , \u4_u0_csr0_reg[0]/P0001 , \u4_u0_csr0_reg[10]/P0001 , \u4_u0_csr0_reg[11]/P0001 , \u4_u0_csr0_reg[12]/P0001 , \u4_u0_csr0_reg[1]/P0001 , \u4_u0_csr0_reg[2]/P0001 , \u4_u0_csr0_reg[3]/NET0131 , \u4_u0_csr0_reg[4]/P0001 , \u4_u0_csr0_reg[5]/P0001 , \u4_u0_csr0_reg[6]/P0001 , \u4_u0_csr0_reg[7]/P0001 , \u4_u0_csr0_reg[8]/P0001 , \u4_u0_csr0_reg[9]/P0001 , \u4_u0_csr1_reg[0]/P0001 , \u4_u0_csr1_reg[10]/P0001 , \u4_u0_csr1_reg[11]/P0001 , \u4_u0_csr1_reg[12]/P0001 , \u4_u0_csr1_reg[1]/P0001 , \u4_u0_csr1_reg[2]/P0001 , \u4_u0_csr1_reg[3]/P0001 , \u4_u0_csr1_reg[4]/P0001 , \u4_u0_csr1_reg[5]/P0001 , \u4_u0_csr1_reg[6]/P0001 , \u4_u0_csr1_reg[7]/P0001 , \u4_u0_csr1_reg[8]/P0001 , \u4_u0_csr1_reg[9]/P0001 , \u4_u0_dma_ack_clr1_reg/P0001 , \u4_u0_dma_ack_wr1_reg/P0001 , \u4_u0_dma_in_buf_sz1_reg/P0001 , \u4_u0_dma_in_cnt_reg[0]/P0001 , \u4_u0_dma_in_cnt_reg[10]/P0001 , \u4_u0_dma_in_cnt_reg[11]/P0001 , \u4_u0_dma_in_cnt_reg[1]/P0001 , \u4_u0_dma_in_cnt_reg[2]/P0001 , \u4_u0_dma_in_cnt_reg[3]/P0001 , \u4_u0_dma_in_cnt_reg[4]/P0001 , \u4_u0_dma_in_cnt_reg[5]/P0001 , \u4_u0_dma_in_cnt_reg[6]/P0001 , \u4_u0_dma_in_cnt_reg[7]/P0001 , \u4_u0_dma_in_cnt_reg[8]/P0001 , \u4_u0_dma_in_cnt_reg[9]/P0001 , \u4_u0_dma_out_buf_avail_reg/P0001 , \u4_u0_dma_out_cnt_reg[10]/P0001 , \u4_u0_dma_out_cnt_reg[11]/P0001 , \u4_u0_dma_out_cnt_reg[1]/P0001 , \u4_u0_dma_out_cnt_reg[2]/P0001 , \u4_u0_dma_out_cnt_reg[3]/P0001 , \u4_u0_dma_out_cnt_reg[4]/P0001 , \u4_u0_dma_out_cnt_reg[5]/P0001 , \u4_u0_dma_out_cnt_reg[6]/P0001 , \u4_u0_dma_out_cnt_reg[7]/P0001 , \u4_u0_dma_out_cnt_reg[8]/P0001 , \u4_u0_dma_out_cnt_reg[9]/P0001 , \u4_u0_dma_out_left_reg[0]/P0001 , \u4_u0_dma_out_left_reg[10]/P0001 , \u4_u0_dma_out_left_reg[11]/P0001 , \u4_u0_dma_out_left_reg[1]/P0001 , \u4_u0_dma_out_left_reg[2]/P0001 , \u4_u0_dma_out_left_reg[3]/P0001 , \u4_u0_dma_out_left_reg[4]/P0001 , \u4_u0_dma_out_left_reg[5]/P0001 , \u4_u0_dma_out_left_reg[6]/P0001 , \u4_u0_dma_out_left_reg[7]/P0001 , \u4_u0_dma_out_left_reg[8]/P0001 , \u4_u0_dma_out_left_reg[9]/P0001 , \u4_u0_dma_req_in_hold2_reg/P0001 , \u4_u0_dma_req_in_hold_reg/P0001 , \u4_u0_dma_req_out_hold_reg/P0001 , \u4_u0_ep_match_r_reg/P0001 , \u4_u0_iena_reg[0]/P0001 , \u4_u0_iena_reg[1]/P0001 , \u4_u0_iena_reg[2]/P0001 , \u4_u0_iena_reg[3]/P0001 , \u4_u0_iena_reg[4]/P0001 , \u4_u0_iena_reg[5]/P0001 , \u4_u0_ienb_reg[0]/P0001 , \u4_u0_ienb_reg[1]/P0001 , \u4_u0_ienb_reg[2]/P0001 , \u4_u0_ienb_reg[3]/P0001 , \u4_u0_ienb_reg[4]/P0001 , \u4_u0_ienb_reg[5]/P0001 , \u4_u0_int_re_reg/P0001 , \u4_u0_int_stat_reg[0]/P0001 , \u4_u0_int_stat_reg[1]/P0001 , \u4_u0_int_stat_reg[2]/P0001 , \u4_u0_int_stat_reg[3]/P0001 , \u4_u0_int_stat_reg[4]/P0001 , \u4_u0_int_stat_reg[5]/P0001 , \u4_u0_int_stat_reg[6]/P0001 , \u4_u0_inta_reg/P0001 , \u4_u0_intb_reg/P0001 , \u4_u0_ots_stop_reg/P0001 , \u4_u0_r1_reg/P0001 , \u4_u0_r2_reg/P0001 , \u4_u0_r4_reg/P0001 , \u4_u0_r5_reg/NET0131 , \u4_u0_set_r_reg/P0001 , \u4_u0_uc_bsel_reg[0]/P0001 , \u4_u0_uc_bsel_reg[1]/P0001 , \u4_u0_uc_dpd_reg[0]/P0001 , \u4_u0_uc_dpd_reg[1]/P0001 , \u4_u1_buf0_orig_m3_reg[0]/P0001 , \u4_u1_buf0_orig_m3_reg[10]/P0001 , \u4_u1_buf0_orig_m3_reg[11]/P0001 , \u4_u1_buf0_orig_m3_reg[1]/P0001 , \u4_u1_buf0_orig_m3_reg[2]/P0001 , \u4_u1_buf0_orig_m3_reg[3]/P0001 , \u4_u1_buf0_orig_m3_reg[4]/P0001 , \u4_u1_buf0_orig_m3_reg[5]/P0001 , \u4_u1_buf0_orig_m3_reg[6]/P0001 , \u4_u1_buf0_orig_m3_reg[7]/P0001 , \u4_u1_buf0_orig_m3_reg[8]/P0001 , \u4_u1_buf0_orig_m3_reg[9]/P0001 , \u4_u1_buf0_orig_reg[0]/P0001 , \u4_u1_buf0_orig_reg[10]/P0001 , \u4_u1_buf0_orig_reg[11]/P0001 , \u4_u1_buf0_orig_reg[12]/P0001 , \u4_u1_buf0_orig_reg[13]/P0001 , \u4_u1_buf0_orig_reg[14]/P0001 , \u4_u1_buf0_orig_reg[15]/P0001 , \u4_u1_buf0_orig_reg[16]/P0001 , \u4_u1_buf0_orig_reg[17]/P0001 , \u4_u1_buf0_orig_reg[18]/P0001 , \u4_u1_buf0_orig_reg[19]/P0001 , \u4_u1_buf0_orig_reg[1]/P0001 , \u4_u1_buf0_orig_reg[20]/P0001 , \u4_u1_buf0_orig_reg[21]/P0001 , \u4_u1_buf0_orig_reg[22]/P0001 , \u4_u1_buf0_orig_reg[23]/P0001 , \u4_u1_buf0_orig_reg[24]/P0001 , \u4_u1_buf0_orig_reg[25]/P0001 , \u4_u1_buf0_orig_reg[26]/P0001 , \u4_u1_buf0_orig_reg[27]/P0001 , \u4_u1_buf0_orig_reg[28]/P0001 , \u4_u1_buf0_orig_reg[29]/NET0131 , \u4_u1_buf0_orig_reg[2]/P0001 , \u4_u1_buf0_orig_reg[30]/NET0131 , \u4_u1_buf0_orig_reg[31]/P0001 , \u4_u1_buf0_orig_reg[3]/P0001 , \u4_u1_buf0_orig_reg[4]/P0001 , \u4_u1_buf0_orig_reg[5]/P0001 , \u4_u1_buf0_orig_reg[6]/P0001 , \u4_u1_buf0_orig_reg[7]/P0001 , \u4_u1_buf0_orig_reg[8]/P0001 , \u4_u1_buf0_orig_reg[9]/P0001 , \u4_u1_buf0_reg[0]/P0001 , \u4_u1_buf0_reg[10]/P0001 , \u4_u1_buf0_reg[11]/P0001 , \u4_u1_buf0_reg[12]/P0001 , \u4_u1_buf0_reg[13]/P0001 , \u4_u1_buf0_reg[14]/P0001 , \u4_u1_buf0_reg[15]/P0001 , \u4_u1_buf0_reg[16]/P0001 , \u4_u1_buf0_reg[17]/P0001 , \u4_u1_buf0_reg[18]/P0001 , \u4_u1_buf0_reg[19]/P0001 , \u4_u1_buf0_reg[1]/P0001 , \u4_u1_buf0_reg[20]/P0001 , \u4_u1_buf0_reg[21]/P0001 , \u4_u1_buf0_reg[22]/P0001 , \u4_u1_buf0_reg[23]/P0001 , \u4_u1_buf0_reg[24]/P0001 , \u4_u1_buf0_reg[25]/P0001 , \u4_u1_buf0_reg[26]/P0001 , \u4_u1_buf0_reg[27]/P0001 , \u4_u1_buf0_reg[28]/P0001 , \u4_u1_buf0_reg[29]/P0001 , \u4_u1_buf0_reg[2]/P0001 , \u4_u1_buf0_reg[30]/P0001 , \u4_u1_buf0_reg[31]/P0001 , \u4_u1_buf0_reg[3]/P0001 , \u4_u1_buf0_reg[4]/P0001 , \u4_u1_buf0_reg[5]/P0001 , \u4_u1_buf0_reg[6]/P0001 , \u4_u1_buf0_reg[7]/P0001 , \u4_u1_buf0_reg[8]/P0001 , \u4_u1_buf0_reg[9]/P0001 , \u4_u1_buf1_reg[0]/P0001 , \u4_u1_buf1_reg[10]/P0001 , \u4_u1_buf1_reg[11]/P0001 , \u4_u1_buf1_reg[12]/P0001 , \u4_u1_buf1_reg[13]/P0001 , \u4_u1_buf1_reg[14]/P0001 , \u4_u1_buf1_reg[15]/P0001 , \u4_u1_buf1_reg[16]/P0001 , \u4_u1_buf1_reg[17]/P0001 , \u4_u1_buf1_reg[18]/P0001 , \u4_u1_buf1_reg[19]/P0001 , \u4_u1_buf1_reg[1]/P0001 , \u4_u1_buf1_reg[20]/P0001 , \u4_u1_buf1_reg[21]/P0001 , \u4_u1_buf1_reg[22]/P0001 , \u4_u1_buf1_reg[23]/P0001 , \u4_u1_buf1_reg[24]/P0001 , \u4_u1_buf1_reg[25]/P0001 , \u4_u1_buf1_reg[26]/P0001 , \u4_u1_buf1_reg[27]/P0001 , \u4_u1_buf1_reg[28]/P0001 , \u4_u1_buf1_reg[29]/P0001 , \u4_u1_buf1_reg[2]/P0001 , \u4_u1_buf1_reg[30]/P0001 , \u4_u1_buf1_reg[31]/P0001 , \u4_u1_buf1_reg[3]/P0001 , \u4_u1_buf1_reg[4]/P0001 , \u4_u1_buf1_reg[5]/P0001 , \u4_u1_buf1_reg[6]/P0001 , \u4_u1_buf1_reg[7]/P0001 , \u4_u1_buf1_reg[8]/P0001 , \u4_u1_buf1_reg[9]/P0001 , \u4_u1_csr0_reg[0]/P0001 , \u4_u1_csr0_reg[10]/P0001 , \u4_u1_csr0_reg[11]/P0001 , \u4_u1_csr0_reg[12]/P0001 , \u4_u1_csr0_reg[1]/P0001 , \u4_u1_csr0_reg[2]/P0001 , \u4_u1_csr0_reg[3]/NET0131 , \u4_u1_csr0_reg[4]/P0001 , \u4_u1_csr0_reg[5]/P0001 , \u4_u1_csr0_reg[6]/P0001 , \u4_u1_csr0_reg[7]/P0001 , \u4_u1_csr0_reg[8]/P0001 , \u4_u1_csr0_reg[9]/P0001 , \u4_u1_csr1_reg[0]/P0001 , \u4_u1_csr1_reg[10]/P0001 , \u4_u1_csr1_reg[11]/P0001 , \u4_u1_csr1_reg[12]/P0001 , \u4_u1_csr1_reg[1]/P0001 , \u4_u1_csr1_reg[2]/P0001 , \u4_u1_csr1_reg[3]/P0001 , \u4_u1_csr1_reg[4]/P0001 , \u4_u1_csr1_reg[5]/P0001 , \u4_u1_csr1_reg[6]/P0001 , \u4_u1_csr1_reg[7]/P0001 , \u4_u1_csr1_reg[8]/P0001 , \u4_u1_csr1_reg[9]/P0001 , \u4_u1_dma_ack_clr1_reg/P0001 , \u4_u1_dma_ack_wr1_reg/P0001 , \u4_u1_dma_in_buf_sz1_reg/P0001 , \u4_u1_dma_in_cnt_reg[0]/P0001 , \u4_u1_dma_in_cnt_reg[10]/P0001 , \u4_u1_dma_in_cnt_reg[11]/P0001 , \u4_u1_dma_in_cnt_reg[1]/P0001 , \u4_u1_dma_in_cnt_reg[2]/P0001 , \u4_u1_dma_in_cnt_reg[3]/P0001 , \u4_u1_dma_in_cnt_reg[4]/P0001 , \u4_u1_dma_in_cnt_reg[5]/P0001 , \u4_u1_dma_in_cnt_reg[6]/P0001 , \u4_u1_dma_in_cnt_reg[7]/P0001 , \u4_u1_dma_in_cnt_reg[8]/P0001 , \u4_u1_dma_in_cnt_reg[9]/P0001 , \u4_u1_dma_out_buf_avail_reg/P0001 , \u4_u1_dma_out_cnt_reg[10]/P0001 , \u4_u1_dma_out_cnt_reg[11]/P0001 , \u4_u1_dma_out_cnt_reg[1]/P0001 , \u4_u1_dma_out_cnt_reg[2]/P0001 , \u4_u1_dma_out_cnt_reg[3]/P0001 , \u4_u1_dma_out_cnt_reg[4]/P0001 , \u4_u1_dma_out_cnt_reg[5]/P0001 , \u4_u1_dma_out_cnt_reg[6]/P0001 , \u4_u1_dma_out_cnt_reg[7]/P0001 , \u4_u1_dma_out_cnt_reg[8]/P0001 , \u4_u1_dma_out_cnt_reg[9]/P0001 , \u4_u1_dma_out_left_reg[0]/P0001 , \u4_u1_dma_out_left_reg[10]/P0001 , \u4_u1_dma_out_left_reg[11]/P0001 , \u4_u1_dma_out_left_reg[1]/P0001 , \u4_u1_dma_out_left_reg[2]/P0001 , \u4_u1_dma_out_left_reg[3]/P0001 , \u4_u1_dma_out_left_reg[4]/P0001 , \u4_u1_dma_out_left_reg[5]/P0001 , \u4_u1_dma_out_left_reg[6]/P0001 , \u4_u1_dma_out_left_reg[7]/P0001 , \u4_u1_dma_out_left_reg[8]/P0001 , \u4_u1_dma_out_left_reg[9]/P0001 , \u4_u1_dma_req_in_hold2_reg/P0001 , \u4_u1_dma_req_in_hold_reg/P0001 , \u4_u1_dma_req_out_hold_reg/P0001 , \u4_u1_ep_match_r_reg/P0001 , \u4_u1_iena_reg[0]/P0001 , \u4_u1_iena_reg[1]/P0001 , \u4_u1_iena_reg[2]/P0001 , \u4_u1_iena_reg[3]/P0001 , \u4_u1_iena_reg[4]/P0001 , \u4_u1_iena_reg[5]/P0001 , \u4_u1_ienb_reg[0]/P0001 , \u4_u1_ienb_reg[1]/P0001 , \u4_u1_ienb_reg[2]/P0001 , \u4_u1_ienb_reg[3]/P0001 , \u4_u1_ienb_reg[4]/P0001 , \u4_u1_ienb_reg[5]/P0001 , \u4_u1_int_re_reg/P0001 , \u4_u1_int_stat_reg[0]/P0001 , \u4_u1_int_stat_reg[1]/P0001 , \u4_u1_int_stat_reg[2]/P0001 , \u4_u1_int_stat_reg[3]/P0001 , \u4_u1_int_stat_reg[4]/P0001 , \u4_u1_int_stat_reg[5]/P0001 , \u4_u1_int_stat_reg[6]/P0001 , \u4_u1_inta_reg/P0001 , \u4_u1_intb_reg/P0001 , \u4_u1_ots_stop_reg/P0001 , \u4_u1_r1_reg/P0001 , \u4_u1_r2_reg/P0001 , \u4_u1_r4_reg/P0001 , \u4_u1_r5_reg/NET0131 , \u4_u1_set_r_reg/P0001 , \u4_u1_uc_bsel_reg[0]/P0001 , \u4_u1_uc_bsel_reg[1]/P0001 , \u4_u1_uc_dpd_reg[0]/P0001 , \u4_u1_uc_dpd_reg[1]/P0001 , \u4_u2_buf0_orig_m3_reg[0]/P0001 , \u4_u2_buf0_orig_m3_reg[10]/P0001 , \u4_u2_buf0_orig_m3_reg[11]/P0001 , \u4_u2_buf0_orig_m3_reg[1]/P0001 , \u4_u2_buf0_orig_m3_reg[2]/P0001 , \u4_u2_buf0_orig_m3_reg[3]/P0001 , \u4_u2_buf0_orig_m3_reg[4]/P0001 , \u4_u2_buf0_orig_m3_reg[5]/P0001 , \u4_u2_buf0_orig_m3_reg[6]/P0001 , \u4_u2_buf0_orig_m3_reg[7]/P0001 , \u4_u2_buf0_orig_m3_reg[8]/P0001 , \u4_u2_buf0_orig_m3_reg[9]/P0001 , \u4_u2_buf0_orig_reg[0]/P0001 , \u4_u2_buf0_orig_reg[10]/P0001 , \u4_u2_buf0_orig_reg[11]/P0001 , \u4_u2_buf0_orig_reg[12]/P0001 , \u4_u2_buf0_orig_reg[13]/P0001 , \u4_u2_buf0_orig_reg[14]/P0001 , \u4_u2_buf0_orig_reg[15]/P0001 , \u4_u2_buf0_orig_reg[16]/P0001 , \u4_u2_buf0_orig_reg[17]/P0001 , \u4_u2_buf0_orig_reg[18]/P0001 , \u4_u2_buf0_orig_reg[19]/P0001 , \u4_u2_buf0_orig_reg[1]/P0001 , \u4_u2_buf0_orig_reg[20]/P0001 , \u4_u2_buf0_orig_reg[21]/P0001 , \u4_u2_buf0_orig_reg[22]/P0001 , \u4_u2_buf0_orig_reg[23]/P0001 , \u4_u2_buf0_orig_reg[24]/P0001 , \u4_u2_buf0_orig_reg[25]/P0001 , \u4_u2_buf0_orig_reg[26]/P0001 , \u4_u2_buf0_orig_reg[27]/P0001 , \u4_u2_buf0_orig_reg[28]/P0001 , \u4_u2_buf0_orig_reg[29]/NET0131 , \u4_u2_buf0_orig_reg[2]/P0001 , \u4_u2_buf0_orig_reg[30]/NET0131 , \u4_u2_buf0_orig_reg[31]/P0001 , \u4_u2_buf0_orig_reg[3]/P0001 , \u4_u2_buf0_orig_reg[4]/P0001 , \u4_u2_buf0_orig_reg[5]/P0001 , \u4_u2_buf0_orig_reg[6]/P0001 , \u4_u2_buf0_orig_reg[7]/P0001 , \u4_u2_buf0_orig_reg[8]/P0001 , \u4_u2_buf0_orig_reg[9]/P0001 , \u4_u2_buf0_reg[0]/P0001 , \u4_u2_buf0_reg[10]/P0001 , \u4_u2_buf0_reg[11]/P0001 , \u4_u2_buf0_reg[12]/P0001 , \u4_u2_buf0_reg[13]/P0001 , \u4_u2_buf0_reg[14]/P0001 , \u4_u2_buf0_reg[15]/P0001 , \u4_u2_buf0_reg[16]/P0001 , \u4_u2_buf0_reg[17]/P0001 , \u4_u2_buf0_reg[18]/P0001 , \u4_u2_buf0_reg[19]/P0001 , \u4_u2_buf0_reg[1]/P0001 , \u4_u2_buf0_reg[20]/P0001 , \u4_u2_buf0_reg[21]/P0001 , \u4_u2_buf0_reg[22]/P0001 , \u4_u2_buf0_reg[23]/P0001 , \u4_u2_buf0_reg[24]/P0001 , \u4_u2_buf0_reg[25]/P0001 , \u4_u2_buf0_reg[26]/P0001 , \u4_u2_buf0_reg[27]/P0001 , \u4_u2_buf0_reg[28]/P0001 , \u4_u2_buf0_reg[29]/P0001 , \u4_u2_buf0_reg[2]/P0001 , \u4_u2_buf0_reg[30]/P0001 , \u4_u2_buf0_reg[31]/P0001 , \u4_u2_buf0_reg[3]/P0001 , \u4_u2_buf0_reg[4]/P0001 , \u4_u2_buf0_reg[5]/P0001 , \u4_u2_buf0_reg[6]/P0001 , \u4_u2_buf0_reg[7]/P0001 , \u4_u2_buf0_reg[8]/P0001 , \u4_u2_buf0_reg[9]/P0001 , \u4_u2_buf1_reg[0]/P0001 , \u4_u2_buf1_reg[10]/P0001 , \u4_u2_buf1_reg[11]/P0001 , \u4_u2_buf1_reg[12]/P0001 , \u4_u2_buf1_reg[13]/P0001 , \u4_u2_buf1_reg[14]/P0001 , \u4_u2_buf1_reg[15]/P0001 , \u4_u2_buf1_reg[16]/P0001 , \u4_u2_buf1_reg[17]/P0001 , \u4_u2_buf1_reg[18]/P0001 , \u4_u2_buf1_reg[19]/P0001 , \u4_u2_buf1_reg[1]/P0001 , \u4_u2_buf1_reg[20]/P0001 , \u4_u2_buf1_reg[21]/P0001 , \u4_u2_buf1_reg[22]/P0001 , \u4_u2_buf1_reg[23]/P0001 , \u4_u2_buf1_reg[24]/P0001 , \u4_u2_buf1_reg[25]/P0001 , \u4_u2_buf1_reg[26]/P0001 , \u4_u2_buf1_reg[27]/P0001 , \u4_u2_buf1_reg[28]/P0001 , \u4_u2_buf1_reg[29]/P0001 , \u4_u2_buf1_reg[2]/P0001 , \u4_u2_buf1_reg[30]/P0001 , \u4_u2_buf1_reg[31]/P0001 , \u4_u2_buf1_reg[3]/P0001 , \u4_u2_buf1_reg[4]/P0001 , \u4_u2_buf1_reg[5]/P0001 , \u4_u2_buf1_reg[6]/P0001 , \u4_u2_buf1_reg[7]/P0001 , \u4_u2_buf1_reg[8]/P0001 , \u4_u2_buf1_reg[9]/P0001 , \u4_u2_csr0_reg[0]/P0001 , \u4_u2_csr0_reg[10]/P0001 , \u4_u2_csr0_reg[11]/P0001 , \u4_u2_csr0_reg[12]/P0001 , \u4_u2_csr0_reg[1]/P0001 , \u4_u2_csr0_reg[2]/P0001 , \u4_u2_csr0_reg[3]/NET0131 , \u4_u2_csr0_reg[4]/P0001 , \u4_u2_csr0_reg[5]/P0001 , \u4_u2_csr0_reg[6]/P0001 , \u4_u2_csr0_reg[7]/P0001 , \u4_u2_csr0_reg[8]/P0001 , \u4_u2_csr0_reg[9]/P0001 , \u4_u2_csr1_reg[0]/P0001 , \u4_u2_csr1_reg[10]/P0001 , \u4_u2_csr1_reg[11]/P0001 , \u4_u2_csr1_reg[12]/P0001 , \u4_u2_csr1_reg[1]/P0001 , \u4_u2_csr1_reg[2]/P0001 , \u4_u2_csr1_reg[3]/P0001 , \u4_u2_csr1_reg[4]/P0001 , \u4_u2_csr1_reg[5]/P0001 , \u4_u2_csr1_reg[6]/P0001 , \u4_u2_csr1_reg[7]/P0001 , \u4_u2_csr1_reg[8]/P0001 , \u4_u2_csr1_reg[9]/P0001 , \u4_u2_dma_ack_clr1_reg/P0001 , \u4_u2_dma_ack_wr1_reg/P0001 , \u4_u2_dma_in_buf_sz1_reg/P0001 , \u4_u2_dma_in_cnt_reg[0]/P0001 , \u4_u2_dma_in_cnt_reg[10]/P0001 , \u4_u2_dma_in_cnt_reg[11]/P0001 , \u4_u2_dma_in_cnt_reg[1]/P0001 , \u4_u2_dma_in_cnt_reg[2]/P0001 , \u4_u2_dma_in_cnt_reg[3]/P0001 , \u4_u2_dma_in_cnt_reg[4]/P0001 , \u4_u2_dma_in_cnt_reg[5]/P0001 , \u4_u2_dma_in_cnt_reg[6]/P0001 , \u4_u2_dma_in_cnt_reg[7]/P0001 , \u4_u2_dma_in_cnt_reg[8]/P0001 , \u4_u2_dma_in_cnt_reg[9]/P0001 , \u4_u2_dma_out_buf_avail_reg/P0001 , \u4_u2_dma_out_cnt_reg[10]/P0001 , \u4_u2_dma_out_cnt_reg[11]/P0001 , \u4_u2_dma_out_cnt_reg[1]/P0001 , \u4_u2_dma_out_cnt_reg[2]/P0001 , \u4_u2_dma_out_cnt_reg[3]/P0001 , \u4_u2_dma_out_cnt_reg[4]/P0001 , \u4_u2_dma_out_cnt_reg[5]/P0001 , \u4_u2_dma_out_cnt_reg[6]/P0001 , \u4_u2_dma_out_cnt_reg[7]/P0001 , \u4_u2_dma_out_cnt_reg[8]/P0001 , \u4_u2_dma_out_cnt_reg[9]/P0001 , \u4_u2_dma_out_left_reg[0]/P0001 , \u4_u2_dma_out_left_reg[10]/P0001 , \u4_u2_dma_out_left_reg[11]/P0001 , \u4_u2_dma_out_left_reg[1]/P0001 , \u4_u2_dma_out_left_reg[2]/P0001 , \u4_u2_dma_out_left_reg[3]/P0001 , \u4_u2_dma_out_left_reg[4]/P0001 , \u4_u2_dma_out_left_reg[5]/P0001 , \u4_u2_dma_out_left_reg[6]/P0001 , \u4_u2_dma_out_left_reg[7]/P0001 , \u4_u2_dma_out_left_reg[8]/P0001 , \u4_u2_dma_out_left_reg[9]/P0001 , \u4_u2_dma_req_in_hold2_reg/P0001 , \u4_u2_dma_req_in_hold_reg/P0001 , \u4_u2_dma_req_out_hold_reg/P0001 , \u4_u2_ep_match_r_reg/P0001 , \u4_u2_iena_reg[0]/P0001 , \u4_u2_iena_reg[1]/P0001 , \u4_u2_iena_reg[2]/P0001 , \u4_u2_iena_reg[3]/P0001 , \u4_u2_iena_reg[4]/P0001 , \u4_u2_iena_reg[5]/P0001 , \u4_u2_ienb_reg[0]/P0001 , \u4_u2_ienb_reg[1]/P0001 , \u4_u2_ienb_reg[2]/P0001 , \u4_u2_ienb_reg[3]/P0001 , \u4_u2_ienb_reg[4]/P0001 , \u4_u2_ienb_reg[5]/P0001 , \u4_u2_int_re_reg/P0001 , \u4_u2_int_stat_reg[0]/P0001 , \u4_u2_int_stat_reg[1]/P0001 , \u4_u2_int_stat_reg[2]/P0001 , \u4_u2_int_stat_reg[3]/P0001 , \u4_u2_int_stat_reg[4]/P0001 , \u4_u2_int_stat_reg[5]/P0001 , \u4_u2_int_stat_reg[6]/P0001 , \u4_u2_inta_reg/P0001 , \u4_u2_intb_reg/P0001 , \u4_u2_ots_stop_reg/P0001 , \u4_u2_r1_reg/P0001 , \u4_u2_r2_reg/P0001 , \u4_u2_r4_reg/P0001 , \u4_u2_r5_reg/NET0131 , \u4_u2_set_r_reg/P0001 , \u4_u2_uc_bsel_reg[0]/P0001 , \u4_u2_uc_bsel_reg[1]/P0001 , \u4_u2_uc_dpd_reg[0]/P0001 , \u4_u2_uc_dpd_reg[1]/P0001 , \u4_u3_buf0_orig_m3_reg[0]/P0001 , \u4_u3_buf0_orig_m3_reg[10]/P0001 , \u4_u3_buf0_orig_m3_reg[11]/P0001 , \u4_u3_buf0_orig_m3_reg[1]/P0001 , \u4_u3_buf0_orig_m3_reg[2]/P0001 , \u4_u3_buf0_orig_m3_reg[3]/P0001 , \u4_u3_buf0_orig_m3_reg[4]/P0001 , \u4_u3_buf0_orig_m3_reg[5]/P0001 , \u4_u3_buf0_orig_m3_reg[6]/P0001 , \u4_u3_buf0_orig_m3_reg[7]/P0001 , \u4_u3_buf0_orig_m3_reg[8]/P0001 , \u4_u3_buf0_orig_m3_reg[9]/P0001 , \u4_u3_buf0_orig_reg[0]/P0001 , \u4_u3_buf0_orig_reg[10]/P0001 , \u4_u3_buf0_orig_reg[11]/P0001 , \u4_u3_buf0_orig_reg[12]/P0001 , \u4_u3_buf0_orig_reg[13]/P0001 , \u4_u3_buf0_orig_reg[14]/P0001 , \u4_u3_buf0_orig_reg[15]/P0001 , \u4_u3_buf0_orig_reg[16]/P0001 , \u4_u3_buf0_orig_reg[17]/P0001 , \u4_u3_buf0_orig_reg[18]/P0001 , \u4_u3_buf0_orig_reg[19]/P0001 , \u4_u3_buf0_orig_reg[1]/P0001 , \u4_u3_buf0_orig_reg[20]/P0001 , \u4_u3_buf0_orig_reg[21]/P0001 , \u4_u3_buf0_orig_reg[22]/P0001 , \u4_u3_buf0_orig_reg[23]/P0001 , \u4_u3_buf0_orig_reg[24]/P0001 , \u4_u3_buf0_orig_reg[25]/P0001 , \u4_u3_buf0_orig_reg[26]/P0001 , \u4_u3_buf0_orig_reg[27]/P0001 , \u4_u3_buf0_orig_reg[28]/P0001 , \u4_u3_buf0_orig_reg[29]/NET0131 , \u4_u3_buf0_orig_reg[2]/P0001 , \u4_u3_buf0_orig_reg[30]/NET0131 , \u4_u3_buf0_orig_reg[31]/P0001 , \u4_u3_buf0_orig_reg[3]/P0001 , \u4_u3_buf0_orig_reg[4]/P0001 , \u4_u3_buf0_orig_reg[5]/P0001 , \u4_u3_buf0_orig_reg[6]/P0001 , \u4_u3_buf0_orig_reg[7]/P0001 , \u4_u3_buf0_orig_reg[8]/P0001 , \u4_u3_buf0_orig_reg[9]/P0001 , \u4_u3_buf0_reg[0]/P0001 , \u4_u3_buf0_reg[10]/P0001 , \u4_u3_buf0_reg[11]/P0001 , \u4_u3_buf0_reg[12]/P0001 , \u4_u3_buf0_reg[13]/P0001 , \u4_u3_buf0_reg[14]/P0001 , \u4_u3_buf0_reg[15]/P0001 , \u4_u3_buf0_reg[16]/P0001 , \u4_u3_buf0_reg[17]/P0001 , \u4_u3_buf0_reg[18]/P0001 , \u4_u3_buf0_reg[19]/P0001 , \u4_u3_buf0_reg[1]/P0001 , \u4_u3_buf0_reg[20]/P0001 , \u4_u3_buf0_reg[21]/P0001 , \u4_u3_buf0_reg[22]/P0001 , \u4_u3_buf0_reg[23]/P0001 , \u4_u3_buf0_reg[24]/P0001 , \u4_u3_buf0_reg[25]/P0001 , \u4_u3_buf0_reg[26]/P0001 , \u4_u3_buf0_reg[27]/P0001 , \u4_u3_buf0_reg[28]/P0001 , \u4_u3_buf0_reg[29]/P0001 , \u4_u3_buf0_reg[2]/P0001 , \u4_u3_buf0_reg[30]/P0001 , \u4_u3_buf0_reg[31]/P0001 , \u4_u3_buf0_reg[3]/P0001 , \u4_u3_buf0_reg[4]/P0001 , \u4_u3_buf0_reg[5]/P0001 , \u4_u3_buf0_reg[6]/P0001 , \u4_u3_buf0_reg[7]/P0001 , \u4_u3_buf0_reg[8]/P0001 , \u4_u3_buf0_reg[9]/P0001 , \u4_u3_buf1_reg[0]/P0001 , \u4_u3_buf1_reg[10]/P0001 , \u4_u3_buf1_reg[11]/P0001 , \u4_u3_buf1_reg[12]/P0001 , \u4_u3_buf1_reg[13]/P0001 , \u4_u3_buf1_reg[14]/P0001 , \u4_u3_buf1_reg[15]/P0001 , \u4_u3_buf1_reg[16]/P0001 , \u4_u3_buf1_reg[17]/P0001 , \u4_u3_buf1_reg[18]/P0001 , \u4_u3_buf1_reg[19]/P0001 , \u4_u3_buf1_reg[1]/P0001 , \u4_u3_buf1_reg[20]/P0001 , \u4_u3_buf1_reg[21]/P0001 , \u4_u3_buf1_reg[22]/P0001 , \u4_u3_buf1_reg[23]/P0001 , \u4_u3_buf1_reg[24]/P0001 , \u4_u3_buf1_reg[25]/P0001 , \u4_u3_buf1_reg[26]/P0001 , \u4_u3_buf1_reg[27]/P0001 , \u4_u3_buf1_reg[28]/P0001 , \u4_u3_buf1_reg[29]/P0001 , \u4_u3_buf1_reg[2]/P0001 , \u4_u3_buf1_reg[30]/P0001 , \u4_u3_buf1_reg[31]/P0001 , \u4_u3_buf1_reg[3]/P0001 , \u4_u3_buf1_reg[4]/P0001 , \u4_u3_buf1_reg[5]/P0001 , \u4_u3_buf1_reg[6]/P0001 , \u4_u3_buf1_reg[7]/P0001 , \u4_u3_buf1_reg[8]/P0001 , \u4_u3_buf1_reg[9]/P0001 , \u4_u3_csr0_reg[0]/P0001 , \u4_u3_csr0_reg[10]/P0001 , \u4_u3_csr0_reg[11]/P0001 , \u4_u3_csr0_reg[12]/P0001 , \u4_u3_csr0_reg[1]/P0001 , \u4_u3_csr0_reg[2]/P0001 , \u4_u3_csr0_reg[3]/NET0131 , \u4_u3_csr0_reg[4]/P0001 , \u4_u3_csr0_reg[5]/P0001 , \u4_u3_csr0_reg[6]/P0001 , \u4_u3_csr0_reg[7]/P0001 , \u4_u3_csr0_reg[8]/P0001 , \u4_u3_csr0_reg[9]/P0001 , \u4_u3_csr1_reg[0]/P0001 , \u4_u3_csr1_reg[10]/P0001 , \u4_u3_csr1_reg[11]/P0001 , \u4_u3_csr1_reg[12]/P0001 , \u4_u3_csr1_reg[1]/P0001 , \u4_u3_csr1_reg[2]/P0001 , \u4_u3_csr1_reg[3]/P0001 , \u4_u3_csr1_reg[4]/P0001 , \u4_u3_csr1_reg[5]/P0001 , \u4_u3_csr1_reg[6]/P0001 , \u4_u3_csr1_reg[7]/P0001 , \u4_u3_csr1_reg[8]/P0001 , \u4_u3_csr1_reg[9]/P0001 , \u4_u3_dma_ack_clr1_reg/P0001 , \u4_u3_dma_ack_wr1_reg/P0001 , \u4_u3_dma_in_buf_sz1_reg/P0001 , \u4_u3_dma_in_cnt_reg[0]/P0001 , \u4_u3_dma_in_cnt_reg[10]/P0001 , \u4_u3_dma_in_cnt_reg[11]/P0001 , \u4_u3_dma_in_cnt_reg[1]/P0001 , \u4_u3_dma_in_cnt_reg[2]/P0001 , \u4_u3_dma_in_cnt_reg[3]/P0001 , \u4_u3_dma_in_cnt_reg[4]/P0001 , \u4_u3_dma_in_cnt_reg[5]/P0001 , \u4_u3_dma_in_cnt_reg[6]/P0001 , \u4_u3_dma_in_cnt_reg[7]/P0001 , \u4_u3_dma_in_cnt_reg[8]/P0001 , \u4_u3_dma_in_cnt_reg[9]/P0001 , \u4_u3_dma_out_buf_avail_reg/P0001 , \u4_u3_dma_out_cnt_reg[10]/P0001 , \u4_u3_dma_out_cnt_reg[11]/P0001 , \u4_u3_dma_out_cnt_reg[1]/P0001 , \u4_u3_dma_out_cnt_reg[2]/P0001 , \u4_u3_dma_out_cnt_reg[3]/P0001 , \u4_u3_dma_out_cnt_reg[4]/P0001 , \u4_u3_dma_out_cnt_reg[5]/P0001 , \u4_u3_dma_out_cnt_reg[6]/P0001 , \u4_u3_dma_out_cnt_reg[7]/P0001 , \u4_u3_dma_out_cnt_reg[8]/P0001 , \u4_u3_dma_out_cnt_reg[9]/P0001 , \u4_u3_dma_out_left_reg[0]/P0001 , \u4_u3_dma_out_left_reg[10]/P0001 , \u4_u3_dma_out_left_reg[11]/P0001 , \u4_u3_dma_out_left_reg[1]/P0001 , \u4_u3_dma_out_left_reg[2]/P0001 , \u4_u3_dma_out_left_reg[3]/P0001 , \u4_u3_dma_out_left_reg[4]/P0001 , \u4_u3_dma_out_left_reg[5]/P0001 , \u4_u3_dma_out_left_reg[6]/P0001 , \u4_u3_dma_out_left_reg[7]/P0001 , \u4_u3_dma_out_left_reg[8]/P0001 , \u4_u3_dma_out_left_reg[9]/P0001 , \u4_u3_dma_req_in_hold2_reg/P0001 , \u4_u3_dma_req_in_hold_reg/P0001 , \u4_u3_dma_req_out_hold_reg/P0001 , \u4_u3_ep_match_r_reg/P0001 , \u4_u3_iena_reg[0]/P0001 , \u4_u3_iena_reg[1]/P0001 , \u4_u3_iena_reg[2]/P0001 , \u4_u3_iena_reg[3]/P0001 , \u4_u3_iena_reg[4]/P0001 , \u4_u3_iena_reg[5]/P0001 , \u4_u3_ienb_reg[0]/P0001 , \u4_u3_ienb_reg[1]/P0001 , \u4_u3_ienb_reg[2]/P0001 , \u4_u3_ienb_reg[3]/P0001 , \u4_u3_ienb_reg[4]/P0001 , \u4_u3_ienb_reg[5]/P0001 , \u4_u3_int_re_reg/P0001 , \u4_u3_int_stat_reg[0]/P0001 , \u4_u3_int_stat_reg[1]/P0001 , \u4_u3_int_stat_reg[2]/P0001 , \u4_u3_int_stat_reg[3]/P0001 , \u4_u3_int_stat_reg[4]/P0001 , \u4_u3_int_stat_reg[5]/P0001 , \u4_u3_int_stat_reg[6]/P0001 , \u4_u3_inta_reg/P0001 , \u4_u3_intb_reg/P0001 , \u4_u3_ots_stop_reg/P0001 , \u4_u3_r1_reg/P0001 , \u4_u3_r2_reg/P0001 , \u4_u3_r4_reg/P0001 , \u4_u3_r5_reg/NET0131 , \u4_u3_set_r_reg/P0001 , \u4_u3_uc_bsel_reg[0]/P0001 , \u4_u3_uc_bsel_reg[1]/P0001 , \u4_u3_uc_dpd_reg[0]/P0001 , \u4_u3_uc_dpd_reg[1]/P0001 , \u4_usb_reset_r_reg/P0001 , \u4_utmi_vend_ctrl_r_reg[0]/P0001 , \u4_utmi_vend_ctrl_r_reg[1]/P0001 , \u4_utmi_vend_ctrl_r_reg[2]/P0001 , \u4_utmi_vend_ctrl_r_reg[3]/P0001 , \u4_utmi_vend_stat_r_reg[0]/P0001 , \u4_utmi_vend_stat_r_reg[1]/P0001 , \u4_utmi_vend_stat_r_reg[2]/P0001 , \u4_utmi_vend_stat_r_reg[3]/P0001 , \u4_utmi_vend_stat_r_reg[4]/P0001 , \u4_utmi_vend_stat_r_reg[5]/P0001 , \u4_utmi_vend_stat_r_reg[6]/P0001 , \u4_utmi_vend_stat_r_reg[7]/P0001 , \u4_utmi_vend_wr_r_reg/P0001 , \u5_state_reg[0]/P0001 , \u5_state_reg[1]/P0001 , \u5_state_reg[2]/P0001 , \u5_state_reg[3]/P0001 , \u5_state_reg[4]/P0001 , \u5_state_reg[5]/NET0131 , \u5_wb_ack_s1_reg/P0001 , \u5_wb_ack_s2_reg/P0001 , \u5_wb_req_s1_reg/P0001 , usb_vbus_pad_i_pad, wb_ack_o_pad, \wb_addr_i[10]_pad , \wb_addr_i[11]_pad , \wb_addr_i[12]_pad , \wb_addr_i[13]_pad , \wb_addr_i[14]_pad , \wb_addr_i[15]_pad , \wb_addr_i[16]_pad , \wb_addr_i[17]_pad , \wb_addr_i[2]_pad , \wb_addr_i[3]_pad , \wb_addr_i[4]_pad , \wb_addr_i[5]_pad , \wb_addr_i[6]_pad , \wb_addr_i[7]_pad , \wb_addr_i[8]_pad , \wb_addr_i[9]_pad , wb_cyc_i_pad, \wb_data_i[0]_pad , \wb_data_i[10]_pad , \wb_data_i[11]_pad , \wb_data_i[12]_pad , \wb_data_i[13]_pad , \wb_data_i[14]_pad , \wb_data_i[15]_pad , \wb_data_i[16]_pad , \wb_data_i[17]_pad , \wb_data_i[18]_pad , \wb_data_i[19]_pad , \wb_data_i[1]_pad , \wb_data_i[20]_pad , \wb_data_i[21]_pad , \wb_data_i[22]_pad , \wb_data_i[23]_pad , \wb_data_i[24]_pad , \wb_data_i[25]_pad , \wb_data_i[26]_pad , \wb_data_i[27]_pad , \wb_data_i[28]_pad , \wb_data_i[29]_pad , \wb_data_i[2]_pad , \wb_data_i[30]_pad , \wb_data_i[31]_pad , \wb_data_i[3]_pad , \wb_data_i[4]_pad , \wb_data_i[5]_pad , \wb_data_i[6]_pad , \wb_data_i[7]_pad , \wb_data_i[8]_pad , \wb_data_i[9]_pad , wb_stb_i_pad, wb_we_i_pad, \dma_req_o[6]_pad , \g37425/_0_ , \g37426/_0_ , \g37432/_0_ , \g37433/_0_ , \g37439/_0_ , \g37440/_0_ , \g37444/_00_ , \g37448/_0_ , \g37450/_0_ , \g37454/_0_ , \g37473/_0_ , \g37474/_0_ , \g37475/_0_ , \g37476/_0_ , \g37477/_0_ , \g37478/_0_ , \g37479/_0_ , \g37488/_0_ , \g37489/_0_ , \g37490/_0_ , \g37491/_0_ , \g37492/_0_ , \g37517/_0_ , \g37518/_0_ , \g37519/_0_ , \g37520/_0_ , \g37521/_0_ , \g37522/_0_ , \g37540/_0_ , \g37542/_0_ , \g37543/_0_ , \g37545/_0_ , \g37546/_0_ , \g37548/_0_ , \g37549/_0_ , \g37550/_0_ , \g37551/_0_ , \g37556/_0_ , \g37589/_0_ , \g37591/_0_ , \g37592/_0_ , \g37593/_0_ , \g37594/_0_ , \g37596/_0_ , \g37597/_0_ , \g37598/_0_ , \g37599/_0_ , \g37601/_0_ , \g37603/_0_ , \g37604/_0_ , \g37605/_0_ , \g37607/_0_ , \g37608/_0_ , \g37609/_0_ , \g37610/_0_ , \g37645/_0_ , \g37648/_0_ , \g37650/_0_ , \g37653/_0_ , \g37664/_3_ , \g37703/_0_ , \g37704/_0_ , \g37706/_0_ , \g37708/_0_ , \g37709/_0_ , \g37711/_0_ , \g37714/_0_ , \g37715/_0_ , \g37717/_0_ , \g37718/_0_ , \g37719/_0_ , \g37720/_0_ , \g37723/_0_ , \g37724/_0_ , \g37726/_0_ , \g37728/_0_ , \g37729/_0_ , \g37730/_0_ , \g37731/_0_ , \g37732/_0_ , \g37733/_0_ , \g37735/_0_ , \g37736/_0_ , \g37737/_0_ , \g37856/_0_ , \g37857/_0_ , \g37859/_0_ , \g37868/_0_ , \g37869/_0_ , \g37870/_0_ , \g37872/_0_ , \g37886/_0_ , \g37887/_0_ , \g37889/_0_ , \g37897/_0_ , \g37899/_0_ , \g37900/_0_ , \g37907/_0_ , \g37925/_0_ , \g37927/_0_ , \g37928/_0_ , \g37929/_0_ , \g37930/_0_ , \g37932/_0_ , \g37933/_0_ , \g37934/_0_ , \g37935/_0_ , \g37936/_0_ , \g37937/_0_ , \g37938/_0_ , \g37939/_0_ , \g37941/_0_ , \g37942/_0_ , \g37943/_0_ , \g37944/_0_ , \g37945/_0_ , \g38030/_3_ , \g38035/_0_ , \g38036/_0_ , \g38054/_0_ , \g38129/_0_ , \g38130/_0_ , \g38148/_3_ , \g38149/_3_ , \g38150/_3_ , \g38166/_0_ , \g38198/_0_ , \g38201/_0_ , \g38257/_0_ , \g38286/_0_ , \g38294/_3_ , \g38295/_3_ , \g38296/_3_ , \g38297/_3_ , \g38332/_0_ , \g38350/_0_ , \g38365/_3_ , \g38366/_3_ , \g38367/_3_ , \g38389/_0_ , \g38397/_0_ , \g38398/_0_ , \g38399/_0_ , \g38400/_0_ , \g38417/_3_ , \g38418/_3_ , \g38422/_0_ , \g38440/_0_ , \g38443/_0_ , \g38448/_3_ , \g38449/_0_ , \g38450/_0_ , \g38460/_0_ , \g38466/_0_ , \g38467/_0_ , \g38468/_0_ , \g38469/_0_ , \g38470/_0_ , \g38471/_0_ , \g38472/_0_ , \g38473/_0_ , \g38474/_0_ , \g38475/_0_ , \g38476/_0_ , \g38477/_0_ , \g38478/_0_ , \g38479/_0_ , \g38528/_0_ , \g38533/_0_ , \g38534/_0_ , \g38536/_0_ , \g38545/_0_ , \g38551/_0_ , \g38554/_0_ , \g38555/_0_ , \g38556/_0_ , \g38575/_0_ , \g38616/_0_ , \g38653/_0_ , \g38656/_0_ , \g38657/_0_ , \g38658/_0_ , \g38660/_0_ , \g38706/_0_ , \g38716/_0_ , \g38717/_0_ , \g38738/_1_ , \g38763/_0_ , \g38790/_0_ , \g38792/_0_ , \g38801/_0_ , \g38803/_0_ , \g38804/_0_ , \g38805/_0_ , \g38806/_0_ , \g38807/_0_ , \g38808/_0_ , \g38809/_0_ , \g38810/_0_ , \g38814/_0_ , \g38833/_0_ , \g38834/_0_ , \g38839/_0_ , \g38840/_0_ , \g38841/_0_ , \g38842/_0_ , \g38846/_0_ , \g38847/_0_ , \g38848/_0_ , \g38849/_0_ , \g38853/_0_ , \g38857/_0_ , \g38872/_0_ , \g38882/_0_ , \g38884/_0_ , \g38885/_0_ , \g38886/_0_ , \g38887/_0_ , \g38931/_0_ , \g38952/_0_ , \g38960/_0_ , \g38971/_0_ , \g38973/_0_ , \g38974/_0_ , \g38975/_0_ , \g38976/_0_ , \g38978/_0_ , \g38981/_0_ , \g38986/_0_ , \g38987/_0_ , \g39001/_3_ , \g39003/_3_ , \g39009/_3_ , \g39011/_3_ , \g39013/_3_ , \g39015/_2_ , \g39017/_2_ , \g39019/_2_ , \g39021/_2_ , \g39060/_0_ , \g39061/_3_ , \g39062/_0_ , \g39063/_0_ , \g39065/_0_ , \g39066/_0_ , \g39093/_0_ , \g39099/_2_ , \g39118/_0_ , \g39123/_0_ , \g39174/_0_ , \g39175/_0_ , \g39176/_0_ , \g39177/_0_ , \g39178/_0_ , \g39185/_0_ , \g39186/_0_ , \g39187/_0_ , \g39188/_0_ , \g39194/_0_ , \g39195/_0_ , \g39196/_0_ , \g39197/_0_ , \g39198/_0_ , \g39199/_0_ , \g39200/_0_ , \g39201/_0_ , \g39202/_0_ , \g39203/_0_ , \g39204/_0_ , \g39216/_3_ , \g39217/_3_ , \g39218/_0_ , \g39219/_0_ , \g39220/_0_ , \g39221/_0_ , \g39299/_0_ , \g39300/_0_ , \g39301/_0_ , \g39302/_0_ , \g39303/_0_ , \g39304/_0_ , \g39305/_0_ , \g39306/_0_ , \g39307/_0_ , \g39308/_0_ , \g39309/_0_ , \g39310/_0_ , \g39311/_0_ , \g39315/_0_ , \g39318/_0_ , \g39321/_0_ , \g39322/_0_ , \g39323/_0_ , \g39333/_0_ , \g39334/_0_ , \g39336/_0_ , \g39338/_0_ , \g39339/_0_ , \g39340/_0_ , \g39341/_0_ , \g39342/_0_ , \g39343/_0_ , \g39344/_0_ , \g39345/_0_ , \g39346/_0_ , \g39349/_0_ , \g39352/_3_ , \g39354/_3_ , \g39371/_3_ , \g39372/_3_ , \g39373/_3_ , \g39374/_3_ , \g39376/_0_ , \g39377/_0_ , \g39471/_0_ , \g39472/_0_ , \g39473/_0_ , \g39474/_0_ , \g39475/_0_ , \g39476/_0_ , \g39477/_0_ , \g39478/_0_ , \g39479/_0_ , \g39480/_0_ , \g39481/_0_ , \g39482/_0_ , \g39483/_0_ , \g39484/_0_ , \g39485/_0_ , \g39486/_0_ , \g39487/_0_ , \g39488/_0_ , \g39492/_0_ , \g39497/_0_ , \g39501/_0_ , \g39502/_0_ , \g39503/_0_ , \g39504/_0_ , \g39505/_0_ , \g39506/_0_ , \g39539/_0_ , \g39541/_0_ , \g39542/_0_ , \g39543/_0_ , \g39544/_0_ , \g39545/_0_ , \g39546/_0_ , \g39547/_0_ , \g39550/_0_ , \g39551/_0_ , \g39563/_0_ , \g39568/_00_ , \g39617/_0_ , \g39618/_0_ , \g39621/_0_ , \g39622/_0_ , \g39623/_0_ , \g39624/_00_ , \g39685/_0_ , \g39690/_0_ , \g39693/_0_ , \g39695/_0_ , \g39697/_0_ , \g39706/_0_ , \g39749/_0_ , \g39750/_0_ , \g39751/_0_ , \g39752/_0_ , \g39753/_0_ , \g39754/_0_ , \g39755/_0_ , \g39756/_0_ , \g39757/_0_ , \g39758/_0_ , \g39759/_0_ , \g39760/_0_ , \g39761/_0_ , \g39762/_0_ , \g39763/_0_ , \g39764/_0_ , \g39765/_0_ , \g39766/_0_ , \g39767/_0_ , \g39768/_0_ , \g39769/_0_ , \g39770/_0_ , \g39772/_0_ , \g39773/_0_ , \g39775/_3_ , \g39776/_3_ , \g39777/_3_ , \g39778/_3_ , \g39779/_3_ , \g39780/_3_ , \g39781/_3_ , \g39782/_3_ , \g39788/_3_ , \g39799/_0_ , \g39800/_0_ , \g39801/_0_ , \g39802/_0_ , \g39927/_0_ , \g39928/_0_ , \g39929/_0_ , \g39930/_0_ , \g39931/_0_ , \g39932/_0_ , \g39933/_0_ , \g39934/_0_ , \g39935/_0_ , \g39936/_0_ , \g39937/_0_ , \g39938/_0_ , \g39939/_0_ , \g39940/_0_ , \g39942/_0_ , \g39943/_0_ , \g39944/_0_ , \g39945/_0_ , \g39956/_0_ , \g39957/_0_ , \g39958/_0_ , \g39959/_0_ , \g39960/_0_ , \g39961/_0_ , \g39962/_0_ , \g39963/_0_ , \g39964/_0_ , \g39969/_0_ , \g39974/_0_ , \g39975/_0_ , \g39993/_0_ , \g39994/_0_ , \g40003/_0_ , \g40004/_0_ , \g40005/_0_ , \g40006/_0_ , \g40016/_0_ , \g40023/_3_ , \g40033/_0_ , \g40034/_0_ , \g40035/_0_ , \g40036/_0_ , \g40037/_0_ , \g40038/_0_ , \g40199/_0_ , \g40200/_0_ , \g40201/_0_ , \g40202/_0_ , \g40203/_0_ , \g40204/_0_ , \g40205/_0_ , \g40206/_0_ , \g40207/_0_ , \g40208/_0_ , \g40209/_0_ , \g40210/_0_ , \g40224/_0_ , \g40225/_0_ , \g40226/_0_ , \g40227/_0_ , \g40234/_0_ , \g40235/_0_ , \g40236/_0_ , \g40237/_0_ , \g40238/_0_ , \g40239/_0_ , \g40240/_0_ , \g40241/_0_ , \g40242/_0_ , \g40243/_0_ , \g40244/_0_ , \g40246/_0_ , \g40247/_0_ , \g40248/_0_ , \g40249/_0_ , \g40250/_0_ , \g40251/_0_ , \g40252/_0_ , \g40253/_0_ , \g40254/_0_ , \g40255/_0_ , \g40257/_0_ , \g40258/_0_ , \g40262/_0_ , \g40264/_0_ , \g40265/_0_ , \g40266/_0_ , \g40267/_0_ , \g40268/_0_ , \g40269/_0_ , \g40270/_0_ , \g40271/_0_ , \g40272/_0_ , \g40273/_0_ , \g40274/_0_ , \g40275/_0_ , \g40276/_0_ , \g40277/_0_ , \g40278/_0_ , \g40280/_2_ , \g40281/_0_ , \g40282/_0_ , \g40283/_0_ , \g40284/_0_ , \g40285/_0_ , \g40286/_0_ , \g40287/_0_ , \g40288/_0_ , \g40289/_0_ , \g40290/_0_ , \g40291/_0_ , \g40297/_0_ , \g40298/_0_ , \g40299/_0_ , \g40300/_0_ , \g40301/_0_ , \g40302/_0_ , \g40303/_0_ , \g40304/_0_ , \g40306/_0_ , \g40307/_0_ , \g40308/_0_ , \g40309/_0_ , \g40310/_0_ , \g40311/_0_ , \g40312/_0_ , \g40313/_0_ , \g40314/_0_ , \g40315/_0_ , \g40316/_0_ , \g40317/_0_ , \g40318/_0_ , \g40319/_0_ , \g40320/_0_ , \g40324/_0_ , \g40325/_0_ , \g40326/_0_ , \g40327/_0_ , \g40328/_0_ , \g40329/_0_ , \g40330/_0_ , \g40331/_0_ , \g40332/_0_ , \g40333/_0_ , \g40334/_0_ , \g40335/_0_ , \g40336/_0_ , \g40337/_0_ , \g40338/_0_ , \g40339/_0_ , \g40340/_0_ , \g40341/_0_ , \g40342/_0_ , \g40343/_0_ , \g40344/_0_ , \g40345/_0_ , \g40346/_0_ , \g40347/_0_ , \g40350/_0_ , \g40353/_0_ , \g40354/_0_ , \g40355/_0_ , \g40374/_0_ , \g40457/_0_ , \g40458/_0_ , \g40549/_0_ , \g40550/_0_ , \g40551/_0_ , \g40552/_0_ , \g40553/_0_ , \g40554/_0_ , \g40556/_0_ , \g40557/_0_ , \g40558/_0_ , \g40559/_0_ , \g40561/_0_ , \g40562/_0_ , \g40563/_0_ , \g40565/_0_ , \g40566/_0_ , \g40567/_0_ , \g40569/_0_ , \g40570/_0_ , \g40571/_0_ , \g40572/_0_ , \g40573/_0_ , \g40574/_0_ , \g40575/_0_ , \g40576/_0_ , \g40577/_0_ , \g40578/_0_ , \g40579/_0_ , \g40580/_0_ , \g40581/_0_ , \g40582/_0_ , \g40583/_0_ , \g40584/_0_ , \g40586/_0_ , \g40587/_0_ , \g40588/_0_ , \g40589/_0_ , \g40591/_0_ , \g40592/_0_ , \g40593/_0_ , \g40594/_0_ , \g40595/_0_ , \g40596/_0_ , \g40597/_0_ , \g40598/_0_ , \g40599/_0_ , \g40600/_0_ , \g40601/_0_ , \g40602/_0_ , \g40603/_0_ , \g40604/_0_ , \g40605/_0_ , \g40606/_0_ , \g40607/_0_ , \g40608/_0_ , \g40609/_0_ , \g40610/_0_ , \g40611/_0_ , \g40612/_0_ , \g40613/_0_ , \g40614/_0_ , \g40617/_0_ , \g40629/_0_ , \g40632/_0_ , \g40633/_0_ , \g40634/_0_ , \g40635/_0_ , \g40636/_0_ , \g40637/_0_ , \g40638/_0_ , \g40639/_0_ , \g40640/_0_ , \g40641/_0_ , \g40642/_0_ , \g40643/_0_ , \g40644/_0_ , \g40645/_0_ , \g40646/_0_ , \g40647/_0_ , \g40648/_0_ , \g40649/_0_ , \g40650/_0_ , \g40651/_0_ , \g40652/_0_ , \g40653/_0_ , \g40654/_0_ , \g40655/_0_ , \g40661/_0_ , \g40663/_0_ , \g40664/_0_ , \g40665/_0_ , \g40666/_0_ , \g40667/_0_ , \g40668/_0_ , \g40669/_0_ , \g40670/_0_ , \g40671/_0_ , \g40672/_0_ , \g40673/_0_ , \g40674/_0_ , \g40675/_0_ , \g40676/_0_ , \g40677/_0_ , \g40678/_0_ , \g40679/_0_ , \g40680/_0_ , \g40681/_0_ , \g40682/_0_ , \g40683/_0_ , \g40684/_0_ , \g40685/_0_ , \g40689/_0_ , \g40690/_0_ , \g40691/_0_ , \g40692/_0_ , \g40693/_0_ , \g40694/_0_ , \g40695/_0_ , \g40696/_0_ , \g40697/_0_ , \g40698/_0_ , \g40699/_0_ , \g40700/_0_ , \g40701/_0_ , \g40702/_0_ , \g40703/_0_ , \g40704/_0_ , \g40705/_0_ , \g40706/_0_ , \g40707/_0_ , \g40708/_0_ , \g40709/_0_ , \g40710/_0_ , \g40711/_0_ , \g40712/_0_ , \g40758/_00_ , \g40759/_0_ , \g40812/_0_ , \g40816/_0_ , \g40817/_0_ , \g40818/_0_ , \g40819/_0_ , \g40820/_0_ , \g40822/_3_ , \g40823/_3_ , \g40824/_3_ , \g40825/_3_ , \g40849/_3_ , \g40915/_0_ , \g40916/_0_ , \g40917/_0_ , \g40920/_0_ , \g40923/_0_ , \g40926/_0_ , \g40927/_0_ , \g40930/_0_ , \g40931/_0_ , \g41138/_0_ , \g41152/_0_ , \g41180/_0_ , \g41185/_0_ , \g41186/_0_ , \g41187/_0_ , \g41189/_0_ , \g41190/_0_ , \g41191/_0_ , \g41192/_0_ , \g41193/_0_ , \g41195/_0_ , \g41199/_0_ , \g41207/_0_ , \g41221/_0_ , \g41226/_0_ , \g41227/_0_ , \g41230/_0_ , \g41231/_0_ , \g41234/_0_ , \g41238/_0_ , \g41239/_0_ , \g41275/_0_ , \g41277/_0_ , \g41278/_0_ , \g41279/_0_ , \g41280/_0_ , \g41281/_0_ , \g41282/_0_ , \g41283/_0_ , \g41284/_0_ , \g41285/_0_ , \g41286/_0_ , \g41287/_0_ , \g41288/_0_ , \g41289/_0_ , \g41291/_3_ , \g41330/_0_ , \g41332/_0_ , \g41334/_0_ , \g41340/_0_ , \g41343/_0_ , \g41345/_0_ , \g41348/_0_ , \g41349/_0_ , \g41350/_0_ , \g41351/_0_ , \g41356/_0_ , \g41394/_0_ , \g41423/_0_ , \g41426/_3_ , \g41427/_3_ , \g41428/_3_ , \g41429/_3_ , \g41430/_3_ , \g41431/_3_ , \g41432/_3_ , \g41433/_3_ , \g41434/_3_ , \g41435/_3_ , \g41436/_3_ , \g41437/_3_ , \g41438/_3_ , \g41439/_3_ , \g41440/_3_ , \g41441/_3_ , \g41442/_0_ , \g41445/_3_ , \g41446/_0_ , \g41449/_0_ , \g41464/_0_ , \g41466/_0_ , \g41468/_0_ , \g41469/_0_ , \g41471/_0_ , \g41795/_0_ , \g41799/_0_ , \g41800/_0_ , \g41801/_0_ , \g41802/_0_ , \g41803/_0_ , \g41804/_0_ , \g41805/_0_ , \g41806/_0_ , \g41807/_0_ , \g41808/_0_ , \g41809/_0_ , \g41810/_0_ , \g41811/_0_ , \g41812/_0_ , \g41814/_0_ , \g41815/_0_ , \g41816/_0_ , \g41817/_0_ , \g41818/_0_ , \g41819/_0_ , \g41820/_0_ , \g41821/_0_ , \g41822/_0_ , \g41823/_0_ , \g41825/_0_ , \g41826/_0_ , \g41827/_0_ , \g41828/_0_ , \g41829/_0_ , \g41830/_0_ , \g41831/_0_ , \g41832/_0_ , \g41833/_0_ , \g41834/_0_ , \g41835/_0_ , \g41836/_0_ , \g41837/_0_ , \g41838/_0_ , \g41839/_0_ , \g41840/_0_ , \g41841/_0_ , \g41842/_0_ , \g41843/_0_ , \g41844/_0_ , \g41845/_0_ , \g41846/_0_ , \g41847/_0_ , \g41848/_0_ , \g41849/_0_ , \g41850/_0_ , \g41851/_0_ , \g41852/_0_ , \g41853/_0_ , \g41854/_0_ , \g41855/_0_ , \g41856/_0_ , \g41857/_0_ , \g41858/_0_ , \g41859/_0_ , \g41860/_0_ , \g41861/_0_ , \g41862/_0_ , \g41863/_0_ , \g41864/_0_ , \g41865/_0_ , \g41866/_0_ , \g41867/_0_ , \g41868/_0_ , \g41869/_0_ , \g41870/_0_ , \g41871/_0_ , \g41872/_0_ , \g41873/_0_ , \g41874/_0_ , \g41875/_0_ , \g41876/_0_ , \g41877/_0_ , \g41878/_0_ , \g41879/_0_ , \g41880/_0_ , \g41881/_0_ , \g41882/_0_ , \g41883/_0_ , \g41884/_0_ , \g41885/_0_ , \g41886/_0_ , \g41887/_0_ , \g41888/_0_ , \g41889/_0_ , \g41890/_0_ , \g41891/_0_ , \g41902/_0_ , \g41904/_0_ , \g41906/_0_ , \g41907/_0_ , \g41954/_0_ , \g41955/_0_ , \g41956/_0_ , \g41957/_0_ , \g41958/_0_ , \g41959/_0_ , \g41960/_0_ , \g41962/_0_ , \g41963/_0_ , \g41964/_0_ , \g41965/_0_ , \g41966/_0_ , \g41967/_0_ , \g41968/_0_ , \g41969/_0_ , \g41970/_0_ , \g41971/_0_ , \g41972/_0_ , \g41973/_0_ , \g41974/_0_ , \g41975/_0_ , \g41976/_0_ , \g41977/_0_ , \g41978/_0_ , \g41979/_0_ , \g42062/_0_ , \g42079/_0_ , \g42142/_0_ , \g42143/_0_ , \g42144/_0_ , \g42154/_0_ , \g42157/_0_ , \g42160/_0_ , \g42181/_0_ , \g42203/_0_ , \g42204/_3_ , \g42205/_3_ , \g42206/_3_ , \g42208/_0_ , \g42220/_0_ , \g42225/_0_ , \g42251/_0_ , \g42273/_0_ , \g42335/_0_ , \g42357/_0_ , \g42380/_0_ , \g42381/_0_ , \g42383/_0_ , \g42386/_0_ , \g42388/_0_ , \g42475/_0_ , \g42476/_0_ , \g42477/_0_ , \g42478/_0_ , \g42479/_0_ , \g42480/_0_ , \g42481/_0_ , \g42482/_0_ , \g42483/_0_ , \g42484/_0_ , \g42485/_0_ , \g42486/_0_ , \g42487/_0_ , \g42488/_0_ , \g42490/_0_ , \g42491/_0_ , \g42493/_0_ , \g42494/_0_ , \g42495/_0_ , \g42496/_0_ , \g42497/_0_ , \g42498/_0_ , \g42499/_0_ , \g42500/_0_ , \g42501/_0_ , \g42502/_0_ , \g42503/_0_ , \g42504/_0_ , \g42505/_0_ , \g42506/_0_ , \g42507/_0_ , \g42508/_0_ , \g42509/_0_ , \g42510/_0_ , \g42511/_0_ , \g42512/_0_ , \g42513/_0_ , \g42514/_0_ , \g42515/_0_ , \g42516/_0_ , \g42517/_0_ , \g42518/_0_ , \g42519/_0_ , \g42521/_0_ , \g42522/_0_ , \g42523/_0_ , \g42524/_0_ , \g42525/_0_ , \g42526/_0_ , \g42527/_0_ , \g42528/_0_ , \g42529/_0_ , \g42530/_0_ , \g42531/_0_ , \g42532/_0_ , \g42533/_0_ , \g42534/_0_ , \g42535/_0_ , \g42536/_0_ , \g42537/_0_ , \g42538/_0_ , \g42539/_0_ , \g42540/_0_ , \g42541/_0_ , \g42542/_0_ , \g42543/_0_ , \g42544/_0_ , \g42545/_0_ , \g42548/_0_ , \g42557/_0_ , \g42564/_0_ , \g42565/_0_ , \g42566/_0_ , \g42567/_0_ , \g42568/_0_ , \g42569/_0_ , \g42570/_0_ , \g42571/_0_ , \g42572/_0_ , \g42573/_0_ , \g42574/_0_ , \g42575/_0_ , \g42576/_0_ , \g42577/_0_ , \g42578/_0_ , \g42581/_0_ , \g42589/_0_ , \g42590/_0_ , \g42591/_0_ , \g42592/_0_ , \g42593/_0_ , \g42594/_0_ , \g42595/_0_ , \g42596/_0_ , \g42597/_0_ , \g42598/_0_ , \g42599/_0_ , \g42600/_0_ , \g42601/_0_ , \g42602/_0_ , \g42603/_0_ , \g42604/_0_ , \g42605/_0_ , \g42606/_0_ , \g42607/_0_ , \g42608/_0_ , \g42609/_0_ , \g42610/_0_ , \g42611/_0_ , \g42612/_0_ , \g42613/_0_ , \g42614/_0_ , \g42615/_0_ , \g42616/_0_ , \g42617/_0_ , \g42618/_0_ , \g42619/_0_ , \g42620/_0_ , \g42622/_0_ , \g42623/_0_ , \g42627/_0_ , \g42628/_0_ , \g42629/_0_ , \g42630/_0_ , \g42631/_0_ , \g42632/_0_ , \g42633/_0_ , \g42634/_0_ , \g42635/_0_ , \g42636/_0_ , \g42637/_0_ , \g42638/_0_ , \g42639/_0_ , \g42640/_0_ , \g42641/_0_ , \g42642/_0_ , \g42643/_0_ , \g42644/_0_ , \g42645/_0_ , \g42646/_0_ , \g42647/_0_ , \g42648/_0_ , \g42649/_0_ , \g42650/_0_ , \g42666/_0_ , \g42667/_0_ , \g42668/_0_ , \g42669/_0_ , \g42670/_0_ , \g42671/_0_ , \g42672/_0_ , \g42673/_0_ , \g42674/_0_ , \g42675/_0_ , \g42676/_0_ , \g42677/_0_ , \g42678/_0_ , \g42680/_0_ , \g42681/_0_ , \g42685/_0_ , \g42686/_0_ , \g42688/_0_ , \g42689/_0_ , \g42690/_0_ , \g42691/_0_ , \g42692/_0_ , \g42693/_0_ , \g42694/_0_ , \g42695/_0_ , \g42696/_0_ , \g42697/_0_ , \g42698/_0_ , \g42699/_0_ , \g42700/_0_ , \g42701/_0_ , \g42702/_0_ , \g42703/_0_ , \g42704/_0_ , \g42705/_0_ , \g42706/_0_ , \g42707/_0_ , \g42708/_0_ , \g42709/_0_ , \g42710/_0_ , \g42711/_0_ , \g42712/_0_ , \g42713/_0_ , \g42715/_0_ , \g42716/_0_ , \g42717/_0_ , \g42718/_0_ , \g42723/_1_ , \g42727/_0_ , \g42728/_0_ , \g42729/_0_ , \g42730/_0_ , \g42731/_0_ , \g42732/_0_ , \g42733/_0_ , \g42734/_0_ , \g42735/_0_ , \g42736/_0_ , \g42737/_0_ , \g42738/_0_ , \g42739/_0_ , \g42740/_0_ , \g42741/_0_ , \g42742/_0_ , \g42743/_0_ , \g42744/_0_ , \g42745/_0_ , \g42746/_0_ , \g42747/_0_ , \g42748/_0_ , \g42749/_0_ , \g42750/_0_ , \g42751/_0_ , \g42754/_0_ , \g42767/_0_ , \g42768/_0_ , \g42772/_0_ , \g42773/_0_ , \g42774/_0_ , \g42775/_0_ , \g42776/_0_ , \g42777/_0_ , \g42778/_0_ , \g42779/_0_ , \g42780/_0_ , \g42781/_0_ , \g42782/_0_ , \g42783/_0_ , \g42784/_0_ , \g42785/_0_ , \g42790/_0_ , \g42791/_0_ , \g42792/_0_ , \g42793/_0_ , \g42794/_0_ , \g42795/_0_ , \g42796/_0_ , \g42797/_0_ , \g42798/_0_ , \g42799/_0_ , \g42800/_0_ , \g42801/_0_ , \g42802/_0_ , \g42803/_0_ , \g42804/_0_ , \g42805/_0_ , \g42806/_0_ , \g42807/_0_ , \g42808/_0_ , \g42809/_0_ , \g42810/_0_ , \g42811/_0_ , \g42812/_0_ , \g42813/_0_ , \g42814/_0_ , \g42815/_0_ , \g42816/_0_ , \g42817/_0_ , \g42818/_0_ , \g42819/_0_ , \g42820/_0_ , \g42821/_0_ , \g42824/_0_ , \g42825/_0_ , \g42826/_0_ , \g42827/_0_ , \g42828/_0_ , \g42829/_0_ , \g42830/_0_ , \g42831/_0_ , \g42832/_0_ , \g42833/_0_ , \g42834/_0_ , \g42835/_0_ , \g42836/_0_ , \g42837/_0_ , \g42838/_0_ , \g42839/_0_ , \g42840/_0_ , \g42841/_0_ , \g42842/_0_ , \g42843/_0_ , \g42844/_0_ , \g42845/_0_ , \g42846/_0_ , \g42907/_0_ , \g42914/_0_ , \g42924/_0_ , \g42925/_0_ , \g42926/_0_ , \g42927/_0_ , \g42928/_0_ , \g42929/_0_ , \g42930/_0_ , \g42931/_0_ , \g42933/_0_ , \g42941/_0_ , \g42947/_0_ , \g42950/_0_ , \g42955/_0_ , \g42956/_0_ , \g42972/_3_ , \g42973/_3_ , \g42974/_3_ , \g43178/_0_ , \g43179/_0_ , \g43184/_0_ , \g43186/_0_ , \g43187/_0_ , \g43190/_0_ , \g43191/_0_ , \g43192/_0_ , \g43202/_0_ , \g43205/_0_ , \g43206/_0_ , \g43207/_0_ , \g43209/_2_ , \g43228/_0_ , \g43233/_0_ , \g43235/_0_ , \g43236/_0_ , \g43237/_0_ , \g43238/_0_ , \g43280/_0_ , \g43287/_0_ , \g43289/_0_ , \g43290/_0_ , \g43291/_0_ , \g43292/_0_ , \g43303/_0_ , \g43311/_0_ , \g43312/_0_ , \g43363/_0_ , \g43364/_0_ , \g43366/_0_ , \g43367/_0_ , \g43370/_0_ , \g43371/_0_ , \g43374/_0_ , \g43413/_0_ , \g43414/_0_ , \g43415/_0_ , \g43416/_0_ , \g43422/_0_ , \g43427/_0_ , \g43428/_0_ , \g43528/_1__syn_2 , \g43630/_0_ , \g43633/_3_ , \g43647/_0_ , \g43648/_0_ , \g43656/_0_ , \g43657/_0_ , \g43667/_0_ , \g43668/_0_ , \g43675/_0_ , \g43678/_0_ , \g43787/_0_ , \g44055/_0_ , \g44092/_0_ , \g44093/_0_ , \g44176/_0_ , \g44181/_0_ , \g44433/_0_ , \g44510/_0_ , \g44515/_2_ , \g44522/_0_ , \g44529/_2_ , \g44537/_2_ , \g44544/_2_ , \g44594/_0_ , \g44695/_0_ , \g44697/_0_ , \g44699/_0_ , \g44700/_0_ , \g44843/_0_ , \g44844/_0_ , \g44879/_0_ , \g44880/_0_ , \g44881/_0_ , \g44882/_0_ , \g44906/_2_ , \g44910/_0_ , \g44912/_0_ , \g44954/_0_ , \g45000/_0_ , \g45001/_0_ , \g45002/_0_ , \g45003/_0_ , \g45021/_1_ , \g45025/_0_ , \g45051/_0_ , \g45104/_0_ , \g45111/_0_ , \g45112/_0_ , \g45116/_0_ , \g45155/_0_ , \g45238/_0_ , \g45239/_0_ , \g45240/_0_ , \g45241/_0_ , \g45249/_0_ , \g45257/_0_ , \g45332/_0_ , \g45334/_0_ , \g45336/_0_ , \g45337/_0_ , \g45342/_0_ , \g45459/_0_ , \g45460/_0_ , \g45466/_0_ , \g45469/_0_ , \g45470/_0_ , \g45474/_0_ , \g45475/_0_ , \g45477/_0_ , \g45481/_0_ , \g45482/_0_ , \g45487/_0_ , \g45488/_0_ , \g45518/_3_ , \g45519/_3_ , \g45520/_3_ , \g45521/_3_ , \g45522/_3_ , \g45523/_3_ , \g45524/_3_ , \g45525/_3_ , \g45526/_3_ , \g45530/_3_ , \g45531/_3_ , \g45532/_3_ , \g45533/_3_ , \g45534/_3_ , \g45535/_3_ , \g45536/_3_ , \g45559/_3_ , \g45596/_0_ , \g45605/_0_ , \g45622/_0_ , \g45623/_0_ , \g45630/_0_ , \g45747/_0_ , \g45753/_0_ , \g45796/_0_ , \g45837/_0_ , \g45882/_0_ , \g45903/_0_ , \g45912/_0_ , \g45946/_0_ , \g45999/_0_ , \g46000/_0_ , \g46001/_0_ , \g46002/_0_ , \g46012/_0_ , \g46014/_0_ , \g46017/_0_ , \g46018/_0_ , \g46021/_0_ , \g46024/_0_ , \g46026/_0_ , \g46029/_0_ , \g46053/_0_ , \g46083/_0_ , \g46093/_0_ , \g46142/_0_ , \g46154/_1__syn_2 , \g46265/_0_ , \g46266/_0_ , \g46268/_0_ , \g46270/_0_ , \g46273/_0_ , \g46274/_0_ , \g46275/_0_ , \g46276/_0_ , \g46278/_0_ , \g46385/_0_ , \g46411/_0_ , \g46414/_0_ , \g46479/_0_ , \g46520/_0_ , \g46521/_0_ , \g46530/_0_ , \g46531/_0_ , \g46597/_0_ , \g46610/_0_ , \g46617/_0_ , \g46632/_0_ , \g46637/_0_ , \g46722/_0_ , \g46723/_0_ , \g46724/_0_ , \g46725/_0_ , \g46813/_0_ , \g46842/_0_ , \g46888/_0_ , \g46891/_0_ , \g46894/_0_ , \g46905/_0_ , \g46940/_0_ , \g46992/_0_ , \g46995/_0_ , \g47037/_3_ , \g47053/_0_ , \g47140/_0_ , \g47155/_3_ , \g47209/_0_ , \g47211/_0_ , \g47213/_0_ , \g47215/_0_ , \g47337/_0_ , \g47433/_0_ , \g47972/_0_ , \g47976/_0_ , \g48081/_0_ , \g48171/_0_ , \g48227/_0_ , \g48234/_1_ , \g48257/_1_ , \g48266/_0_ , \g48281/_0_ , \g48291/_1_ , \g48322/_0_ , \g48345/_0_ , \g48429/_0_ , \g48495/_1_ , \g48549/_0_ , \g48589/_0_ , \g48642/_0_ , \g48722/_0_ , \g48748/_0_ , \g48749/_0_ , \g48763/_0_ , \g48867/_0_ , \g48876/_0_ , \g48880/_0_ , \g49023/_0_ , \g49205/_0_ , \g49314/_0_ , \g49432/_0__syn_2 , \g49512/_0_ , \g49707/_0_ , \g49737/_0_ , \g49831/_0_ , \g49922/_1_ , \g50132/_0_ , \g51376/_0_ , \g51412/_0_ , \g51822/_0_ , \g52114/_0_ , \g52156/_0_ , \g54427/_0_ , \g54557/_0_ , \g54561/_3_ , \g55079/_0_ , \sram_adr_o[0]_pad , \sram_adr_o[10]_pad , \sram_adr_o[11]_pad , \sram_adr_o[12]_pad , \sram_adr_o[13]_pad , \sram_adr_o[14]_pad , \sram_adr_o[1]_pad , \sram_adr_o[2]_pad , \sram_adr_o[3]_pad , \sram_adr_o[4]_pad , \sram_adr_o[5]_pad , \sram_adr_o[6]_pad , \sram_adr_o[7]_pad , \sram_adr_o[8]_pad , \sram_adr_o[9]_pad , \sram_data_o[0]_pad , \sram_data_o[10]_pad , \sram_data_o[11]_pad , \sram_data_o[12]_pad , \sram_data_o[13]_pad , \sram_data_o[14]_pad , \sram_data_o[15]_pad , \sram_data_o[16]_pad , \sram_data_o[17]_pad , \sram_data_o[18]_pad , \sram_data_o[19]_pad , \sram_data_o[1]_pad , \sram_data_o[20]_pad , \sram_data_o[21]_pad , \sram_data_o[22]_pad , \sram_data_o[23]_pad , \sram_data_o[24]_pad , \sram_data_o[25]_pad , \sram_data_o[26]_pad , \sram_data_o[27]_pad , \sram_data_o[28]_pad , \sram_data_o[29]_pad , \sram_data_o[2]_pad , \sram_data_o[30]_pad , \sram_data_o[31]_pad , \sram_data_o[3]_pad , \sram_data_o[4]_pad , \sram_data_o[5]_pad , \sram_data_o[6]_pad , \sram_data_o[7]_pad , \sram_data_o[8]_pad , \sram_data_o[9]_pad , sram_re_o_pad, sram_we_o_pad, \u4_utmi_vend_ctrl_r_reg[0]/P0001_reg_syn_3 , \u4_utmi_vend_ctrl_r_reg[1]/P0001_reg_syn_3 , \u4_utmi_vend_ctrl_r_reg[2]/P0001_reg_syn_3 , \u4_utmi_vend_ctrl_r_reg[3]/P0001_reg_syn_3 );
	input \DataOut_pad_o[0]_pad  ;
	input \DataOut_pad_o[1]_pad  ;
	input \DataOut_pad_o[2]_pad  ;
	input \DataOut_pad_o[3]_pad  ;
	input \DataOut_pad_o[4]_pad  ;
	input \DataOut_pad_o[5]_pad  ;
	input \DataOut_pad_o[6]_pad  ;
	input \DataOut_pad_o[7]_pad  ;
	input \LineState_pad_i[0]_pad  ;
	input \LineState_pad_i[1]_pad  ;
	input \LineState_r_reg[0]/P0001  ;
	input \LineState_r_reg[1]/P0001  ;
	input \OpMode_pad_o[1]_pad  ;
	input RxActive_pad_i_pad ;
	input RxError_pad_i_pad ;
	input RxValid_pad_i_pad ;
	input TermSel_pad_o_pad ;
	input TxReady_pad_i_pad ;
	input TxValid_pad_o_pad ;
	input VControl_Load_pad_o_pad ;
	input XcvSelect_pad_o_pad ;
	input \dma_ack_i[0]_pad  ;
	input \dma_ack_i[1]_pad  ;
	input \dma_ack_i[2]_pad  ;
	input \dma_ack_i[3]_pad  ;
	input \dma_req_o[0]_pad  ;
	input \dma_req_o[1]_pad  ;
	input \dma_req_o[2]_pad  ;
	input \dma_req_o[3]_pad  ;
	input resume_req_i_pad ;
	input \resume_req_r_reg/P0001  ;
	input rst_i_pad ;
	input \sram_data_i[0]_pad  ;
	input \sram_data_i[10]_pad  ;
	input \sram_data_i[11]_pad  ;
	input \sram_data_i[12]_pad  ;
	input \sram_data_i[13]_pad  ;
	input \sram_data_i[14]_pad  ;
	input \sram_data_i[15]_pad  ;
	input \sram_data_i[16]_pad  ;
	input \sram_data_i[17]_pad  ;
	input \sram_data_i[18]_pad  ;
	input \sram_data_i[19]_pad  ;
	input \sram_data_i[1]_pad  ;
	input \sram_data_i[20]_pad  ;
	input \sram_data_i[21]_pad  ;
	input \sram_data_i[22]_pad  ;
	input \sram_data_i[23]_pad  ;
	input \sram_data_i[24]_pad  ;
	input \sram_data_i[25]_pad  ;
	input \sram_data_i[26]_pad  ;
	input \sram_data_i[27]_pad  ;
	input \sram_data_i[28]_pad  ;
	input \sram_data_i[29]_pad  ;
	input \sram_data_i[2]_pad  ;
	input \sram_data_i[30]_pad  ;
	input \sram_data_i[31]_pad  ;
	input \sram_data_i[3]_pad  ;
	input \sram_data_i[4]_pad  ;
	input \sram_data_i[5]_pad  ;
	input \sram_data_i[6]_pad  ;
	input \sram_data_i[7]_pad  ;
	input \sram_data_i[8]_pad  ;
	input \sram_data_i[9]_pad  ;
	input susp_o_pad ;
	input \suspend_clr_wr_reg/P0001  ;
	input \u0_drive_k_r_reg/P0001  ;
	input \u0_rx_active_reg/P0001  ;
	input \u0_rx_data_reg[0]/P0001  ;
	input \u0_rx_data_reg[1]/P0001  ;
	input \u0_rx_data_reg[2]/P0001  ;
	input \u0_rx_data_reg[3]/P0001  ;
	input \u0_rx_data_reg[4]/P0001  ;
	input \u0_rx_data_reg[5]/P0001  ;
	input \u0_rx_data_reg[6]/P0001  ;
	input \u0_rx_data_reg[7]/P0001  ;
	input \u0_rx_err_reg/P0001  ;
	input \u0_rx_valid_reg/P0001  ;
	input \u0_tx_ready_reg/NET0131  ;
	input \u0_u0_T1_gt_2_5_uS_reg/P0001  ;
	input \u0_u0_T1_gt_3_0_mS_reg/P0001  ;
	input \u0_u0_T1_gt_5_0_mS_reg/P0001  ;
	input \u0_u0_T1_st_3_0_mS_reg/P0001  ;
	input \u0_u0_T2_gt_100_uS_reg/P0001  ;
	input \u0_u0_T2_gt_1_0_mS_reg/P0001  ;
	input \u0_u0_T2_wakeup_reg/P0001  ;
	input \u0_u0_chirp_cnt_is_6_reg/P0001  ;
	input \u0_u0_chirp_cnt_reg[0]/P0001  ;
	input \u0_u0_chirp_cnt_reg[1]/P0001  ;
	input \u0_u0_chirp_cnt_reg[2]/P0001  ;
	input \u0_u0_drive_k_reg/P0001  ;
	input \u0_u0_idle_cnt1_clr_reg/P0001  ;
	input \u0_u0_idle_cnt1_next_reg[0]/P0001  ;
	input \u0_u0_idle_cnt1_next_reg[1]/P0001  ;
	input \u0_u0_idle_cnt1_next_reg[2]/P0001  ;
	input \u0_u0_idle_cnt1_next_reg[3]/P0001  ;
	input \u0_u0_idle_cnt1_next_reg[4]/P0001  ;
	input \u0_u0_idle_cnt1_next_reg[5]/P0001  ;
	input \u0_u0_idle_cnt1_next_reg[6]/P0001  ;
	input \u0_u0_idle_cnt1_next_reg[7]/P0001  ;
	input \u0_u0_idle_cnt1_reg[0]/P0001  ;
	input \u0_u0_idle_cnt1_reg[1]/P0001  ;
	input \u0_u0_idle_cnt1_reg[2]/P0001  ;
	input \u0_u0_idle_cnt1_reg[3]/P0001  ;
	input \u0_u0_idle_cnt1_reg[4]/P0001  ;
	input \u0_u0_idle_cnt1_reg[5]/P0001  ;
	input \u0_u0_idle_cnt1_reg[6]/P0001  ;
	input \u0_u0_idle_cnt1_reg[7]/P0001  ;
	input \u0_u0_idle_long_reg/P0001  ;
	input \u0_u0_ls_idle_r_reg/P0001  ;
	input \u0_u0_ls_j_r_reg/P0001  ;
	input \u0_u0_ls_k_r_reg/P0001  ;
	input \u0_u0_ls_se0_r_reg/P0001  ;
	input \u0_u0_me_cnt_100_ms_reg/P0001  ;
	input \u0_u0_me_cnt_reg[0]/P0001  ;
	input \u0_u0_me_cnt_reg[1]/P0001  ;
	input \u0_u0_me_cnt_reg[2]/P0001  ;
	input \u0_u0_me_cnt_reg[3]/P0001  ;
	input \u0_u0_me_cnt_reg[4]/P0001  ;
	input \u0_u0_me_cnt_reg[5]/P0001  ;
	input \u0_u0_me_cnt_reg[6]/P0001  ;
	input \u0_u0_me_cnt_reg[7]/P0001  ;
	input \u0_u0_me_ps2_0_5_ms_reg/P0001  ;
	input \u0_u0_me_ps2_reg[0]/P0001  ;
	input \u0_u0_me_ps2_reg[1]/P0001  ;
	input \u0_u0_me_ps2_reg[2]/P0001  ;
	input \u0_u0_me_ps2_reg[3]/P0001  ;
	input \u0_u0_me_ps2_reg[4]/P0001  ;
	input \u0_u0_me_ps2_reg[5]/P0001  ;
	input \u0_u0_me_ps2_reg[6]/P0001  ;
	input \u0_u0_me_ps2_reg[7]/P0001  ;
	input \u0_u0_me_ps_2_5_us_reg/P0001  ;
	input \u0_u0_me_ps_reg[0]/P0001  ;
	input \u0_u0_me_ps_reg[1]/P0001  ;
	input \u0_u0_me_ps_reg[2]/P0001  ;
	input \u0_u0_me_ps_reg[3]/P0001  ;
	input \u0_u0_me_ps_reg[4]/P0001  ;
	input \u0_u0_me_ps_reg[5]/P0001  ;
	input \u0_u0_me_ps_reg[6]/P0001  ;
	input \u0_u0_me_ps_reg[7]/P0001  ;
	input \u0_u0_mode_hs_reg/P0001  ;
	input \u0_u0_ps_cnt_clr_reg/P0001  ;
	input \u0_u0_ps_cnt_reg[0]/P0001  ;
	input \u0_u0_ps_cnt_reg[1]/P0001  ;
	input \u0_u0_ps_cnt_reg[2]/P0001  ;
	input \u0_u0_ps_cnt_reg[3]/P0001  ;
	input \u0_u0_resume_req_s_reg/P0001  ;
	input \u0_u0_state_reg[0]/NET0131  ;
	input \u0_u0_state_reg[10]/P0001  ;
	input \u0_u0_state_reg[11]/NET0131  ;
	input \u0_u0_state_reg[12]/NET0131  ;
	input \u0_u0_state_reg[13]/NET0131  ;
	input \u0_u0_state_reg[14]/P0001  ;
	input \u0_u0_state_reg[1]/P0001  ;
	input \u0_u0_state_reg[2]/NET0131  ;
	input \u0_u0_state_reg[3]/P0001  ;
	input \u0_u0_state_reg[4]/NET0131  ;
	input \u0_u0_state_reg[5]/P0001  ;
	input \u0_u0_state_reg[6]/NET0131  ;
	input \u0_u0_state_reg[7]/NET0131  ;
	input \u0_u0_state_reg[8]/NET0131  ;
	input \u0_u0_state_reg[9]/P0001  ;
	input \u0_u0_usb_attached_reg/P0001  ;
	input \u0_u0_usb_suspend_reg/P0001  ;
	input \u1_clr_sof_time_reg/P0001  ;
	input \u1_frame_no_r_reg[0]/P0001  ;
	input \u1_frame_no_r_reg[10]/P0001  ;
	input \u1_frame_no_r_reg[1]/P0001  ;
	input \u1_frame_no_r_reg[2]/P0001  ;
	input \u1_frame_no_r_reg[3]/P0001  ;
	input \u1_frame_no_r_reg[4]/P0001  ;
	input \u1_frame_no_r_reg[5]/P0001  ;
	input \u1_frame_no_r_reg[6]/P0001  ;
	input \u1_frame_no_r_reg[7]/P0001  ;
	input \u1_frame_no_r_reg[8]/P0001  ;
	input \u1_frame_no_r_reg[9]/P0001  ;
	input \u1_frame_no_same_reg/P0001  ;
	input \u1_hms_clk_reg/P0001  ;
	input \u1_hms_cnt_reg[0]/P0001  ;
	input \u1_hms_cnt_reg[1]/P0001  ;
	input \u1_hms_cnt_reg[2]/P0001  ;
	input \u1_hms_cnt_reg[3]/P0001  ;
	input \u1_hms_cnt_reg[4]/P0001  ;
	input \u1_mfm_cnt_reg[0]/P0001  ;
	input \u1_mfm_cnt_reg[1]/P0001  ;
	input \u1_mfm_cnt_reg[2]/P0001  ;
	input \u1_mfm_cnt_reg[3]/P0001  ;
	input \u1_sof_time_reg[0]/P0001  ;
	input \u1_sof_time_reg[10]/P0001  ;
	input \u1_sof_time_reg[11]/P0001  ;
	input \u1_sof_time_reg[1]/P0001  ;
	input \u1_sof_time_reg[2]/P0001  ;
	input \u1_sof_time_reg[3]/P0001  ;
	input \u1_sof_time_reg[4]/P0001  ;
	input \u1_sof_time_reg[5]/P0001  ;
	input \u1_sof_time_reg[6]/P0001  ;
	input \u1_sof_time_reg[7]/P0001  ;
	input \u1_sof_time_reg[8]/P0001  ;
	input \u1_sof_time_reg[9]/P0001  ;
	input \u1_u0_crc16_sum_reg[0]/P0001  ;
	input \u1_u0_crc16_sum_reg[10]/P0001  ;
	input \u1_u0_crc16_sum_reg[11]/P0001  ;
	input \u1_u0_crc16_sum_reg[12]/P0001  ;
	input \u1_u0_crc16_sum_reg[13]/P0001  ;
	input \u1_u0_crc16_sum_reg[14]/P0001  ;
	input \u1_u0_crc16_sum_reg[15]/P0001  ;
	input \u1_u0_crc16_sum_reg[1]/P0001  ;
	input \u1_u0_crc16_sum_reg[2]/P0001  ;
	input \u1_u0_crc16_sum_reg[3]/P0001  ;
	input \u1_u0_crc16_sum_reg[4]/P0001  ;
	input \u1_u0_crc16_sum_reg[5]/P0001  ;
	input \u1_u0_crc16_sum_reg[6]/P0001  ;
	input \u1_u0_crc16_sum_reg[7]/P0001  ;
	input \u1_u0_crc16_sum_reg[8]/P0001  ;
	input \u1_u0_crc16_sum_reg[9]/P0001  ;
	input \u1_u0_data_valid0_reg/P0001  ;
	input \u1_u0_pid_reg[0]/NET0131  ;
	input \u1_u0_pid_reg[1]/NET0131  ;
	input \u1_u0_pid_reg[2]/NET0131  ;
	input \u1_u0_pid_reg[3]/NET0131  ;
	input \u1_u0_pid_reg[4]/P0001  ;
	input \u1_u0_pid_reg[5]/P0001  ;
	input \u1_u0_pid_reg[6]/P0001  ;
	input \u1_u0_pid_reg[7]/P0001  ;
	input \u1_u0_rx_active_r_reg/P0001  ;
	input \u1_u0_rxv1_reg/P0001  ;
	input \u1_u0_rxv2_reg/P0001  ;
	input \u1_u0_state_reg[0]/P0001  ;
	input \u1_u0_state_reg[1]/P0001  ;
	input \u1_u0_state_reg[2]/P0001  ;
	input \u1_u0_state_reg[3]/P0001  ;
	input \u1_u0_token0_reg[0]/NET0131  ;
	input \u1_u0_token0_reg[1]/P0001  ;
	input \u1_u0_token0_reg[2]/NET0131  ;
	input \u1_u0_token0_reg[3]/NET0131  ;
	input \u1_u0_token0_reg[4]/P0001  ;
	input \u1_u0_token0_reg[5]/NET0131  ;
	input \u1_u0_token0_reg[6]/P0001  ;
	input \u1_u0_token0_reg[7]/P0001  ;
	input \u1_u0_token1_reg[0]/P0001  ;
	input \u1_u0_token1_reg[1]/P0001  ;
	input \u1_u0_token1_reg[2]/P0001  ;
	input \u1_u0_token1_reg[3]/P0001  ;
	input \u1_u0_token1_reg[4]/P0001  ;
	input \u1_u0_token1_reg[5]/P0001  ;
	input \u1_u0_token1_reg[6]/P0001  ;
	input \u1_u0_token1_reg[7]/P0001  ;
	input \u1_u0_token_valid_r1_reg/P0001  ;
	input \u1_u0_token_valid_str1_reg/P0001  ;
	input \u1_u1_crc16_reg[0]/P0001  ;
	input \u1_u1_crc16_reg[10]/P0001  ;
	input \u1_u1_crc16_reg[11]/P0001  ;
	input \u1_u1_crc16_reg[12]/P0001  ;
	input \u1_u1_crc16_reg[13]/P0001  ;
	input \u1_u1_crc16_reg[14]/P0001  ;
	input \u1_u1_crc16_reg[15]/P0001  ;
	input \u1_u1_crc16_reg[1]/P0001  ;
	input \u1_u1_crc16_reg[2]/P0001  ;
	input \u1_u1_crc16_reg[3]/P0001  ;
	input \u1_u1_crc16_reg[4]/P0001  ;
	input \u1_u1_crc16_reg[5]/P0001  ;
	input \u1_u1_crc16_reg[6]/P0001  ;
	input \u1_u1_crc16_reg[7]/P0001  ;
	input \u1_u1_crc16_reg[8]/P0001  ;
	input \u1_u1_crc16_reg[9]/P0001  ;
	input \u1_u1_send_data_r2_reg/P0001  ;
	input \u1_u1_send_data_r_reg/P0001  ;
	input \u1_u1_send_token_r_reg/P0001  ;
	input \u1_u1_send_zero_length_r_reg/P0001  ;
	input \u1_u1_state_reg[0]/NET0131  ;
	input \u1_u1_state_reg[1]/NET0131  ;
	input \u1_u1_state_reg[2]/NET0131  ;
	input \u1_u1_state_reg[3]/NET0131  ;
	input \u1_u1_state_reg[4]/NET0131  ;
	input \u1_u1_tx_first_r_reg/P0001  ;
	input \u1_u1_tx_valid_r_reg/NET0131  ;
	input \u1_u1_zero_length_r_reg/P0001  ;
	input \u1_u2_adr_cb_reg[0]/NET0131  ;
	input \u1_u2_adr_cb_reg[1]/NET0131  ;
	input \u1_u2_adr_cb_reg[2]/NET0131  ;
	input \u1_u2_adr_cw_reg[0]/NET0131  ;
	input \u1_u2_adr_cw_reg[10]/P0001  ;
	input \u1_u2_adr_cw_reg[11]/P0001  ;
	input \u1_u2_adr_cw_reg[12]/P0001  ;
	input \u1_u2_adr_cw_reg[13]/P0001  ;
	input \u1_u2_adr_cw_reg[14]/P0001  ;
	input \u1_u2_adr_cw_reg[1]/P0001  ;
	input \u1_u2_adr_cw_reg[2]/P0001  ;
	input \u1_u2_adr_cw_reg[3]/NET0131  ;
	input \u1_u2_adr_cw_reg[4]/P0001  ;
	input \u1_u2_adr_cw_reg[5]/NET0131  ;
	input \u1_u2_adr_cw_reg[6]/NET0131  ;
	input \u1_u2_adr_cw_reg[7]/NET0131  ;
	input \u1_u2_adr_cw_reg[8]/P0001  ;
	input \u1_u2_adr_cw_reg[9]/NET0131  ;
	input \u1_u2_dout_r_reg[0]/P0001  ;
	input \u1_u2_dout_r_reg[10]/P0001  ;
	input \u1_u2_dout_r_reg[11]/P0001  ;
	input \u1_u2_dout_r_reg[12]/P0001  ;
	input \u1_u2_dout_r_reg[13]/P0001  ;
	input \u1_u2_dout_r_reg[14]/P0001  ;
	input \u1_u2_dout_r_reg[15]/P0001  ;
	input \u1_u2_dout_r_reg[16]/P0001  ;
	input \u1_u2_dout_r_reg[17]/P0001  ;
	input \u1_u2_dout_r_reg[18]/P0001  ;
	input \u1_u2_dout_r_reg[19]/P0001  ;
	input \u1_u2_dout_r_reg[1]/P0001  ;
	input \u1_u2_dout_r_reg[20]/P0001  ;
	input \u1_u2_dout_r_reg[21]/P0001  ;
	input \u1_u2_dout_r_reg[22]/P0001  ;
	input \u1_u2_dout_r_reg[23]/P0001  ;
	input \u1_u2_dout_r_reg[24]/P0001  ;
	input \u1_u2_dout_r_reg[25]/P0001  ;
	input \u1_u2_dout_r_reg[26]/P0001  ;
	input \u1_u2_dout_r_reg[27]/P0001  ;
	input \u1_u2_dout_r_reg[28]/P0001  ;
	input \u1_u2_dout_r_reg[29]/P0001  ;
	input \u1_u2_dout_r_reg[2]/P0001  ;
	input \u1_u2_dout_r_reg[30]/P0001  ;
	input \u1_u2_dout_r_reg[31]/P0001  ;
	input \u1_u2_dout_r_reg[3]/P0001  ;
	input \u1_u2_dout_r_reg[4]/P0001  ;
	input \u1_u2_dout_r_reg[5]/P0001  ;
	input \u1_u2_dout_r_reg[6]/P0001  ;
	input \u1_u2_dout_r_reg[7]/P0001  ;
	input \u1_u2_dout_r_reg[8]/P0001  ;
	input \u1_u2_dout_r_reg[9]/P0001  ;
	input \u1_u2_dtmp_r_reg[0]/P0001  ;
	input \u1_u2_dtmp_r_reg[10]/P0001  ;
	input \u1_u2_dtmp_r_reg[11]/P0001  ;
	input \u1_u2_dtmp_r_reg[12]/P0001  ;
	input \u1_u2_dtmp_r_reg[13]/P0001  ;
	input \u1_u2_dtmp_r_reg[14]/P0001  ;
	input \u1_u2_dtmp_r_reg[15]/P0001  ;
	input \u1_u2_dtmp_r_reg[16]/P0001  ;
	input \u1_u2_dtmp_r_reg[17]/P0001  ;
	input \u1_u2_dtmp_r_reg[18]/P0001  ;
	input \u1_u2_dtmp_r_reg[19]/P0001  ;
	input \u1_u2_dtmp_r_reg[1]/P0001  ;
	input \u1_u2_dtmp_r_reg[20]/P0001  ;
	input \u1_u2_dtmp_r_reg[21]/P0001  ;
	input \u1_u2_dtmp_r_reg[22]/P0001  ;
	input \u1_u2_dtmp_r_reg[23]/P0001  ;
	input \u1_u2_dtmp_r_reg[24]/P0001  ;
	input \u1_u2_dtmp_r_reg[25]/P0001  ;
	input \u1_u2_dtmp_r_reg[26]/P0001  ;
	input \u1_u2_dtmp_r_reg[27]/P0001  ;
	input \u1_u2_dtmp_r_reg[28]/P0001  ;
	input \u1_u2_dtmp_r_reg[29]/P0001  ;
	input \u1_u2_dtmp_r_reg[2]/P0001  ;
	input \u1_u2_dtmp_r_reg[30]/P0001  ;
	input \u1_u2_dtmp_r_reg[31]/P0001  ;
	input \u1_u2_dtmp_r_reg[3]/P0001  ;
	input \u1_u2_dtmp_r_reg[4]/P0001  ;
	input \u1_u2_dtmp_r_reg[5]/P0001  ;
	input \u1_u2_dtmp_r_reg[6]/P0001  ;
	input \u1_u2_dtmp_r_reg[7]/P0001  ;
	input \u1_u2_dtmp_r_reg[8]/P0001  ;
	input \u1_u2_dtmp_r_reg[9]/P0001  ;
	input \u1_u2_dtmp_sel_r_reg/P0001  ;
	input \u1_u2_idma_done_reg/P0001  ;
	input \u1_u2_last_buf_adr_reg[0]/P0001  ;
	input \u1_u2_last_buf_adr_reg[10]/P0001  ;
	input \u1_u2_last_buf_adr_reg[11]/P0001  ;
	input \u1_u2_last_buf_adr_reg[12]/P0001  ;
	input \u1_u2_last_buf_adr_reg[13]/P0001  ;
	input \u1_u2_last_buf_adr_reg[14]/P0001  ;
	input \u1_u2_last_buf_adr_reg[1]/P0001  ;
	input \u1_u2_last_buf_adr_reg[2]/P0001  ;
	input \u1_u2_last_buf_adr_reg[3]/P0001  ;
	input \u1_u2_last_buf_adr_reg[4]/P0001  ;
	input \u1_u2_last_buf_adr_reg[5]/P0001  ;
	input \u1_u2_last_buf_adr_reg[6]/P0001  ;
	input \u1_u2_last_buf_adr_reg[7]/P0001  ;
	input \u1_u2_last_buf_adr_reg[8]/P0001  ;
	input \u1_u2_last_buf_adr_reg[9]/P0001  ;
	input \u1_u2_mack_r_reg/P0001  ;
	input \u1_u2_mwe_reg/P0001  ;
	input \u1_u2_rd_buf0_reg[0]/NET0131  ;
	input \u1_u2_rd_buf0_reg[10]/NET0131  ;
	input \u1_u2_rd_buf0_reg[11]/NET0131  ;
	input \u1_u2_rd_buf0_reg[12]/P0001  ;
	input \u1_u2_rd_buf0_reg[13]/P0001  ;
	input \u1_u2_rd_buf0_reg[14]/P0001  ;
	input \u1_u2_rd_buf0_reg[15]/P0001  ;
	input \u1_u2_rd_buf0_reg[16]/NET0131  ;
	input \u1_u2_rd_buf0_reg[17]/NET0131  ;
	input \u1_u2_rd_buf0_reg[18]/NET0131  ;
	input \u1_u2_rd_buf0_reg[19]/NET0131  ;
	input \u1_u2_rd_buf0_reg[1]/NET0131  ;
	input \u1_u2_rd_buf0_reg[20]/P0001  ;
	input \u1_u2_rd_buf0_reg[21]/P0001  ;
	input \u1_u2_rd_buf0_reg[22]/P0001  ;
	input \u1_u2_rd_buf0_reg[23]/P0001  ;
	input \u1_u2_rd_buf0_reg[24]/NET0131  ;
	input \u1_u2_rd_buf0_reg[25]/NET0131  ;
	input \u1_u2_rd_buf0_reg[26]/NET0131  ;
	input \u1_u2_rd_buf0_reg[27]/NET0131  ;
	input \u1_u2_rd_buf0_reg[28]/P0001  ;
	input \u1_u2_rd_buf0_reg[29]/P0001  ;
	input \u1_u2_rd_buf0_reg[2]/NET0131  ;
	input \u1_u2_rd_buf0_reg[30]/P0001  ;
	input \u1_u2_rd_buf0_reg[31]/P0001  ;
	input \u1_u2_rd_buf0_reg[3]/NET0131  ;
	input \u1_u2_rd_buf0_reg[4]/P0001  ;
	input \u1_u2_rd_buf0_reg[5]/P0001  ;
	input \u1_u2_rd_buf0_reg[6]/P0001  ;
	input \u1_u2_rd_buf0_reg[7]/P0001  ;
	input \u1_u2_rd_buf0_reg[8]/NET0131  ;
	input \u1_u2_rd_buf0_reg[9]/NET0131  ;
	input \u1_u2_rd_buf1_reg[0]/NET0131  ;
	input \u1_u2_rd_buf1_reg[10]/NET0131  ;
	input \u1_u2_rd_buf1_reg[11]/NET0131  ;
	input \u1_u2_rd_buf1_reg[12]/P0001  ;
	input \u1_u2_rd_buf1_reg[13]/P0001  ;
	input \u1_u2_rd_buf1_reg[14]/P0001  ;
	input \u1_u2_rd_buf1_reg[15]/P0001  ;
	input \u1_u2_rd_buf1_reg[16]/NET0131  ;
	input \u1_u2_rd_buf1_reg[17]/NET0131  ;
	input \u1_u2_rd_buf1_reg[18]/NET0131  ;
	input \u1_u2_rd_buf1_reg[19]/NET0131  ;
	input \u1_u2_rd_buf1_reg[1]/NET0131  ;
	input \u1_u2_rd_buf1_reg[20]/P0001  ;
	input \u1_u2_rd_buf1_reg[21]/P0001  ;
	input \u1_u2_rd_buf1_reg[22]/P0001  ;
	input \u1_u2_rd_buf1_reg[23]/P0001  ;
	input \u1_u2_rd_buf1_reg[24]/NET0131  ;
	input \u1_u2_rd_buf1_reg[25]/NET0131  ;
	input \u1_u2_rd_buf1_reg[26]/NET0131  ;
	input \u1_u2_rd_buf1_reg[27]/NET0131  ;
	input \u1_u2_rd_buf1_reg[28]/P0001  ;
	input \u1_u2_rd_buf1_reg[29]/P0001  ;
	input \u1_u2_rd_buf1_reg[2]/NET0131  ;
	input \u1_u2_rd_buf1_reg[30]/P0001  ;
	input \u1_u2_rd_buf1_reg[31]/P0001  ;
	input \u1_u2_rd_buf1_reg[3]/NET0131  ;
	input \u1_u2_rd_buf1_reg[4]/P0001  ;
	input \u1_u2_rd_buf1_reg[5]/P0001  ;
	input \u1_u2_rd_buf1_reg[6]/P0001  ;
	input \u1_u2_rd_buf1_reg[7]/P0001  ;
	input \u1_u2_rd_buf1_reg[8]/NET0131  ;
	input \u1_u2_rd_buf1_reg[9]/NET0131  ;
	input \u1_u2_rx_data_done_r2_reg/P0001  ;
	input \u1_u2_rx_data_done_r_reg/P0001  ;
	input \u1_u2_rx_data_st_r_reg[0]/P0001  ;
	input \u1_u2_rx_data_st_r_reg[1]/P0001  ;
	input \u1_u2_rx_data_st_r_reg[2]/P0001  ;
	input \u1_u2_rx_data_st_r_reg[3]/P0001  ;
	input \u1_u2_rx_data_st_r_reg[4]/P0001  ;
	input \u1_u2_rx_data_st_r_reg[5]/P0001  ;
	input \u1_u2_rx_data_st_r_reg[6]/P0001  ;
	input \u1_u2_rx_data_st_r_reg[7]/P0001  ;
	input \u1_u2_rx_data_valid_r_reg/NET0131  ;
	input \u1_u2_rx_dma_en_r_reg/P0001  ;
	input \u1_u2_send_data_r_reg/NET0131  ;
	input \u1_u2_sizd_c_reg[0]/P0001  ;
	input \u1_u2_sizd_c_reg[10]/P0001  ;
	input \u1_u2_sizd_c_reg[11]/P0001  ;
	input \u1_u2_sizd_c_reg[12]/P0001  ;
	input \u1_u2_sizd_c_reg[13]/P0001  ;
	input \u1_u2_sizd_c_reg[1]/P0001  ;
	input \u1_u2_sizd_c_reg[2]/P0001  ;
	input \u1_u2_sizd_c_reg[3]/P0001  ;
	input \u1_u2_sizd_c_reg[4]/P0001  ;
	input \u1_u2_sizd_c_reg[5]/P0001  ;
	input \u1_u2_sizd_c_reg[6]/P0001  ;
	input \u1_u2_sizd_c_reg[7]/P0001  ;
	input \u1_u2_sizd_c_reg[8]/P0001  ;
	input \u1_u2_sizd_c_reg[9]/P0001  ;
	input \u1_u2_sizd_is_zero_reg/P0001  ;
	input \u1_u2_sizu_c_reg[0]/P0001  ;
	input \u1_u2_sizu_c_reg[10]/P0001  ;
	input \u1_u2_sizu_c_reg[1]/P0001  ;
	input \u1_u2_sizu_c_reg[2]/P0001  ;
	input \u1_u2_sizu_c_reg[3]/P0001  ;
	input \u1_u2_sizu_c_reg[4]/P0001  ;
	input \u1_u2_sizu_c_reg[5]/P0001  ;
	input \u1_u2_sizu_c_reg[6]/P0001  ;
	input \u1_u2_sizu_c_reg[7]/P0001  ;
	input \u1_u2_sizu_c_reg[8]/NET0131  ;
	input \u1_u2_sizu_c_reg[9]/P0001  ;
	input \u1_u2_state_reg[0]/P0001  ;
	input \u1_u2_state_reg[1]/NET0131  ;
	input \u1_u2_state_reg[2]/NET0131  ;
	input \u1_u2_state_reg[3]/NET0131  ;
	input \u1_u2_state_reg[4]/NET0131  ;
	input \u1_u2_state_reg[5]/NET0131  ;
	input \u1_u2_state_reg[6]/NET0131  ;
	input \u1_u2_state_reg[7]/NET0131  ;
	input \u1_u2_tx_dma_en_r_reg/P0001  ;
	input \u1_u2_word_done_r_reg/P0001  ;
	input \u1_u2_word_done_reg/NET0131  ;
	input \u1_u2_wr_done_reg/P0001  ;
	input \u1_u2_wr_last_reg/P0001  ;
	input \u1_u3_abort_reg/P0001  ;
	input \u1_u3_adr_r_reg[0]/P0001  ;
	input \u1_u3_adr_r_reg[10]/P0001  ;
	input \u1_u3_adr_r_reg[11]/P0001  ;
	input \u1_u3_adr_r_reg[12]/P0001  ;
	input \u1_u3_adr_r_reg[13]/P0001  ;
	input \u1_u3_adr_r_reg[14]/P0001  ;
	input \u1_u3_adr_r_reg[15]/P0001  ;
	input \u1_u3_adr_r_reg[16]/P0001  ;
	input \u1_u3_adr_r_reg[1]/P0001  ;
	input \u1_u3_adr_r_reg[2]/P0001  ;
	input \u1_u3_adr_r_reg[3]/P0001  ;
	input \u1_u3_adr_r_reg[4]/P0001  ;
	input \u1_u3_adr_r_reg[5]/P0001  ;
	input \u1_u3_adr_r_reg[6]/P0001  ;
	input \u1_u3_adr_r_reg[7]/P0001  ;
	input \u1_u3_adr_r_reg[8]/P0001  ;
	input \u1_u3_adr_r_reg[9]/P0001  ;
	input \u1_u3_adr_reg[0]/P0001  ;
	input \u1_u3_adr_reg[10]/P0001  ;
	input \u1_u3_adr_reg[11]/P0001  ;
	input \u1_u3_adr_reg[12]/P0001  ;
	input \u1_u3_adr_reg[13]/P0001  ;
	input \u1_u3_adr_reg[14]/P0001  ;
	input \u1_u3_adr_reg[15]/P0001  ;
	input \u1_u3_adr_reg[16]/P0001  ;
	input \u1_u3_adr_reg[1]/P0001  ;
	input \u1_u3_adr_reg[2]/P0001  ;
	input \u1_u3_adr_reg[3]/P0001  ;
	input \u1_u3_adr_reg[4]/P0001  ;
	input \u1_u3_adr_reg[5]/P0001  ;
	input \u1_u3_adr_reg[6]/P0001  ;
	input \u1_u3_adr_reg[7]/P0001  ;
	input \u1_u3_adr_reg[8]/P0001  ;
	input \u1_u3_adr_reg[9]/P0001  ;
	input \u1_u3_buf0_na_reg/NET0131  ;
	input \u1_u3_buf0_not_aloc_reg/P0001  ;
	input \u1_u3_buf0_rl_reg/P0001  ;
	input \u1_u3_buf0_set_reg/P0001  ;
	input \u1_u3_buf0_st_max_reg/P0001  ;
	input \u1_u3_buf1_na_reg/NET0131  ;
	input \u1_u3_buf1_not_aloc_reg/P0001  ;
	input \u1_u3_buf1_set_reg/P0001  ;
	input \u1_u3_buf1_st_max_reg/P0001  ;
	input \u1_u3_buffer_done_reg/P0001  ;
	input \u1_u3_buffer_empty_reg/P0001  ;
	input \u1_u3_buffer_full_reg/P0001  ;
	input \u1_u3_buffer_overflow_reg/P0001  ;
	input \u1_u3_idin_reg[0]/P0001  ;
	input \u1_u3_idin_reg[10]/P0001  ;
	input \u1_u3_idin_reg[11]/P0001  ;
	input \u1_u3_idin_reg[12]/P0001  ;
	input \u1_u3_idin_reg[13]/P0001  ;
	input \u1_u3_idin_reg[14]/P0001  ;
	input \u1_u3_idin_reg[15]/P0001  ;
	input \u1_u3_idin_reg[16]/P0001  ;
	input \u1_u3_idin_reg[17]/P0001  ;
	input \u1_u3_idin_reg[18]/P0001  ;
	input \u1_u3_idin_reg[19]/P0001  ;
	input \u1_u3_idin_reg[1]/P0001  ;
	input \u1_u3_idin_reg[20]/P0001  ;
	input \u1_u3_idin_reg[21]/P0001  ;
	input \u1_u3_idin_reg[22]/P0001  ;
	input \u1_u3_idin_reg[23]/P0001  ;
	input \u1_u3_idin_reg[24]/P0001  ;
	input \u1_u3_idin_reg[25]/P0001  ;
	input \u1_u3_idin_reg[26]/P0001  ;
	input \u1_u3_idin_reg[27]/P0001  ;
	input \u1_u3_idin_reg[28]/P0001  ;
	input \u1_u3_idin_reg[29]/P0001  ;
	input \u1_u3_idin_reg[2]/P0001  ;
	input \u1_u3_idin_reg[30]/P0001  ;
	input \u1_u3_idin_reg[31]/P0001  ;
	input \u1_u3_idin_reg[3]/P0001  ;
	input \u1_u3_idin_reg[4]/P0001  ;
	input \u1_u3_idin_reg[5]/P0001  ;
	input \u1_u3_idin_reg[6]/P0001  ;
	input \u1_u3_idin_reg[7]/P0001  ;
	input \u1_u3_idin_reg[8]/P0001  ;
	input \u1_u3_idin_reg[9]/P0001  ;
	input \u1_u3_in_token_reg/NET0131  ;
	input \u1_u3_int_seqerr_set_reg/P0001  ;
	input \u1_u3_int_upid_set_reg/P0001  ;
	input \u1_u3_match_r_reg/P0001  ;
	input \u1_u3_new_size_reg[0]/P0001  ;
	input \u1_u3_new_size_reg[10]/P0001  ;
	input \u1_u3_new_size_reg[11]/P0001  ;
	input \u1_u3_new_size_reg[12]/P0001  ;
	input \u1_u3_new_size_reg[13]/P0001  ;
	input \u1_u3_new_size_reg[1]/P0001  ;
	input \u1_u3_new_size_reg[2]/P0001  ;
	input \u1_u3_new_size_reg[3]/P0001  ;
	input \u1_u3_new_size_reg[4]/P0001  ;
	input \u1_u3_new_size_reg[5]/P0001  ;
	input \u1_u3_new_size_reg[6]/P0001  ;
	input \u1_u3_new_size_reg[7]/P0001  ;
	input \u1_u3_new_size_reg[8]/P0001  ;
	input \u1_u3_new_size_reg[9]/P0001  ;
	input \u1_u3_new_sizeb_reg[0]/P0001  ;
	input \u1_u3_new_sizeb_reg[10]/P0001  ;
	input \u1_u3_new_sizeb_reg[1]/P0001  ;
	input \u1_u3_new_sizeb_reg[2]/P0001  ;
	input \u1_u3_new_sizeb_reg[3]/P0001  ;
	input \u1_u3_new_sizeb_reg[4]/P0001  ;
	input \u1_u3_new_sizeb_reg[5]/P0001  ;
	input \u1_u3_new_sizeb_reg[6]/P0001  ;
	input \u1_u3_new_sizeb_reg[7]/P0001  ;
	input \u1_u3_new_sizeb_reg[8]/P0001  ;
	input \u1_u3_new_sizeb_reg[9]/P0001  ;
	input \u1_u3_next_dpid_reg[0]/P0001  ;
	input \u1_u3_next_dpid_reg[1]/P0001  ;
	input \u1_u3_no_bufs0_reg/P0001  ;
	input \u1_u3_no_bufs1_reg/P0001  ;
	input \u1_u3_out_to_small_r_reg/P0001  ;
	input \u1_u3_out_to_small_reg/P0001  ;
	input \u1_u3_out_token_reg/NET0131  ;
	input \u1_u3_pid_IN_r_reg/P0001  ;
	input \u1_u3_pid_OUT_r_reg/P0001  ;
	input \u1_u3_pid_PING_r_reg/P0001  ;
	input \u1_u3_pid_SETUP_r_reg/P0001  ;
	input \u1_u3_pid_seq_err_reg/P0001  ;
	input \u1_u3_rx_ack_to_clr_reg/P0001  ;
	input \u1_u3_rx_ack_to_cnt_reg[0]/P0001  ;
	input \u1_u3_rx_ack_to_cnt_reg[1]/P0001  ;
	input \u1_u3_rx_ack_to_cnt_reg[2]/P0001  ;
	input \u1_u3_rx_ack_to_cnt_reg[3]/P0001  ;
	input \u1_u3_rx_ack_to_cnt_reg[4]/P0001  ;
	input \u1_u3_rx_ack_to_cnt_reg[5]/P0001  ;
	input \u1_u3_rx_ack_to_cnt_reg[6]/P0001  ;
	input \u1_u3_rx_ack_to_cnt_reg[7]/P0001  ;
	input \u1_u3_rx_ack_to_reg/P0001  ;
	input \u1_u3_send_token_reg/P0001  ;
	input \u1_u3_setup_token_reg/P0001  ;
	input \u1_u3_size_next_r_reg[0]/P0001  ;
	input \u1_u3_size_next_r_reg[10]/P0001  ;
	input \u1_u3_size_next_r_reg[1]/P0001  ;
	input \u1_u3_size_next_r_reg[2]/P0001  ;
	input \u1_u3_size_next_r_reg[3]/P0001  ;
	input \u1_u3_size_next_r_reg[4]/P0001  ;
	input \u1_u3_size_next_r_reg[5]/P0001  ;
	input \u1_u3_size_next_r_reg[6]/P0001  ;
	input \u1_u3_size_next_r_reg[7]/P0001  ;
	input \u1_u3_size_next_r_reg[8]/P0001  ;
	input \u1_u3_size_next_r_reg[9]/P0001  ;
	input \u1_u3_state_reg[0]/P0001  ;
	input \u1_u3_state_reg[1]/P0001  ;
	input \u1_u3_state_reg[2]/P0001  ;
	input \u1_u3_state_reg[3]/P0001  ;
	input \u1_u3_state_reg[4]/P0001  ;
	input \u1_u3_state_reg[5]/P0001  ;
	input \u1_u3_state_reg[6]/P0001  ;
	input \u1_u3_state_reg[7]/P0001  ;
	input \u1_u3_state_reg[8]/P0001  ;
	input \u1_u3_state_reg[9]/P0001  ;
	input \u1_u3_this_dpid_reg[0]/P0001  ;
	input \u1_u3_this_dpid_reg[1]/P0001  ;
	input \u1_u3_to_large_reg/P0001  ;
	input \u1_u3_to_small_reg/P0001  ;
	input \u1_u3_token_pid_sel_reg[0]/P0001  ;
	input \u1_u3_token_pid_sel_reg[1]/P0001  ;
	input \u1_u3_tx_data_to_cnt_reg[0]/P0001  ;
	input \u1_u3_tx_data_to_cnt_reg[1]/P0001  ;
	input \u1_u3_tx_data_to_cnt_reg[2]/P0001  ;
	input \u1_u3_tx_data_to_cnt_reg[3]/P0001  ;
	input \u1_u3_tx_data_to_cnt_reg[4]/P0001  ;
	input \u1_u3_tx_data_to_cnt_reg[5]/P0001  ;
	input \u1_u3_tx_data_to_cnt_reg[6]/P0001  ;
	input \u1_u3_tx_data_to_cnt_reg[7]/P0001  ;
	input \u1_u3_tx_data_to_reg/P0001  ;
	input \u1_u3_uc_bsel_set_reg/P0001  ;
	input \u2_wack_r_reg/P0001  ;
	input \u4_attach_r1_reg/P0001  ;
	input \u4_attach_r_reg/P0001  ;
	input \u4_buf0_reg[0]/P0001  ;
	input \u4_buf0_reg[10]/P0001  ;
	input \u4_buf0_reg[11]/P0001  ;
	input \u4_buf0_reg[12]/P0001  ;
	input \u4_buf0_reg[13]/P0001  ;
	input \u4_buf0_reg[14]/P0001  ;
	input \u4_buf0_reg[15]/P0001  ;
	input \u4_buf0_reg[16]/P0001  ;
	input \u4_buf0_reg[17]/NET0131  ;
	input \u4_buf0_reg[18]/P0001  ;
	input \u4_buf0_reg[19]/NET0131  ;
	input \u4_buf0_reg[1]/P0001  ;
	input \u4_buf0_reg[20]/NET0131  ;
	input \u4_buf0_reg[21]/NET0131  ;
	input \u4_buf0_reg[22]/NET0131  ;
	input \u4_buf0_reg[23]/NET0131  ;
	input \u4_buf0_reg[24]/NET0131  ;
	input \u4_buf0_reg[25]/NET0131  ;
	input \u4_buf0_reg[26]/NET0131  ;
	input \u4_buf0_reg[27]/P0001  ;
	input \u4_buf0_reg[28]/P0001  ;
	input \u4_buf0_reg[29]/P0001  ;
	input \u4_buf0_reg[2]/P0001  ;
	input \u4_buf0_reg[30]/P0001  ;
	input \u4_buf0_reg[31]/P0001  ;
	input \u4_buf0_reg[3]/P0001  ;
	input \u4_buf0_reg[4]/P0001  ;
	input \u4_buf0_reg[5]/P0001  ;
	input \u4_buf0_reg[6]/P0001  ;
	input \u4_buf0_reg[7]/P0001  ;
	input \u4_buf0_reg[8]/P0001  ;
	input \u4_buf0_reg[9]/P0001  ;
	input \u4_buf1_reg[0]/P0001  ;
	input \u4_buf1_reg[10]/P0001  ;
	input \u4_buf1_reg[11]/P0001  ;
	input \u4_buf1_reg[12]/P0001  ;
	input \u4_buf1_reg[13]/P0001  ;
	input \u4_buf1_reg[14]/P0001  ;
	input \u4_buf1_reg[15]/P0001  ;
	input \u4_buf1_reg[16]/P0001  ;
	input \u4_buf1_reg[17]/NET0131  ;
	input \u4_buf1_reg[18]/P0001  ;
	input \u4_buf1_reg[19]/NET0131  ;
	input \u4_buf1_reg[1]/P0001  ;
	input \u4_buf1_reg[20]/NET0131  ;
	input \u4_buf1_reg[21]/NET0131  ;
	input \u4_buf1_reg[22]/NET0131  ;
	input \u4_buf1_reg[23]/NET0131  ;
	input \u4_buf1_reg[24]/NET0131  ;
	input \u4_buf1_reg[25]/NET0131  ;
	input \u4_buf1_reg[26]/NET0131  ;
	input \u4_buf1_reg[27]/P0001  ;
	input \u4_buf1_reg[28]/P0001  ;
	input \u4_buf1_reg[29]/P0001  ;
	input \u4_buf1_reg[2]/P0001  ;
	input \u4_buf1_reg[30]/P0001  ;
	input \u4_buf1_reg[31]/P0001  ;
	input \u4_buf1_reg[3]/P0001  ;
	input \u4_buf1_reg[4]/P0001  ;
	input \u4_buf1_reg[5]/P0001  ;
	input \u4_buf1_reg[6]/P0001  ;
	input \u4_buf1_reg[7]/P0001  ;
	input \u4_buf1_reg[8]/P0001  ;
	input \u4_buf1_reg[9]/P0001  ;
	input \u4_crc5_err_r_reg/P0001  ;
	input \u4_csr_reg[0]/P0001  ;
	input \u4_csr_reg[10]/P0001  ;
	input \u4_csr_reg[11]/P0001  ;
	input \u4_csr_reg[12]/P0001  ;
	input \u4_csr_reg[15]/NET0131  ;
	input \u4_csr_reg[16]/P0001  ;
	input \u4_csr_reg[17]/P0001  ;
	input \u4_csr_reg[1]/P0001  ;
	input \u4_csr_reg[22]/P0001  ;
	input \u4_csr_reg[23]/P0001  ;
	input \u4_csr_reg[24]/P0001  ;
	input \u4_csr_reg[25]/P0001  ;
	input \u4_csr_reg[26]/NET0131  ;
	input \u4_csr_reg[27]/NET0131  ;
	input \u4_csr_reg[28]/P0001  ;
	input \u4_csr_reg[29]/P0001  ;
	input \u4_csr_reg[2]/NET0131  ;
	input \u4_csr_reg[30]/NET0131  ;
	input \u4_csr_reg[31]/P0001  ;
	input \u4_csr_reg[3]/P0001  ;
	input \u4_csr_reg[4]/NET0131  ;
	input \u4_csr_reg[5]/NET0131  ;
	input \u4_csr_reg[6]/NET0131  ;
	input \u4_csr_reg[7]/P0001  ;
	input \u4_csr_reg[8]/P0001  ;
	input \u4_csr_reg[9]/NET0131  ;
	input \u4_dma_in_buf_sz1_reg/P0001  ;
	input \u4_dma_out_buf_avail_reg/P0001  ;
	input \u4_dout_reg[0]/P0001  ;
	input \u4_dout_reg[10]/P0001  ;
	input \u4_dout_reg[11]/P0001  ;
	input \u4_dout_reg[12]/P0001  ;
	input \u4_dout_reg[13]/P0001  ;
	input \u4_dout_reg[14]/P0001  ;
	input \u4_dout_reg[15]/P0001  ;
	input \u4_dout_reg[16]/P0001  ;
	input \u4_dout_reg[17]/P0001  ;
	input \u4_dout_reg[18]/P0001  ;
	input \u4_dout_reg[19]/P0001  ;
	input \u4_dout_reg[1]/P0001  ;
	input \u4_dout_reg[20]/P0001  ;
	input \u4_dout_reg[21]/P0001  ;
	input \u4_dout_reg[22]/P0001  ;
	input \u4_dout_reg[23]/P0001  ;
	input \u4_dout_reg[24]/P0001  ;
	input \u4_dout_reg[25]/P0001  ;
	input \u4_dout_reg[26]/P0001  ;
	input \u4_dout_reg[27]/P0001  ;
	input \u4_dout_reg[28]/P0001  ;
	input \u4_dout_reg[29]/P0001  ;
	input \u4_dout_reg[2]/P0001  ;
	input \u4_dout_reg[30]/P0001  ;
	input \u4_dout_reg[31]/P0001  ;
	input \u4_dout_reg[3]/P0001  ;
	input \u4_dout_reg[4]/P0001  ;
	input \u4_dout_reg[5]/P0001  ;
	input \u4_dout_reg[6]/P0001  ;
	input \u4_dout_reg[7]/P0001  ;
	input \u4_dout_reg[8]/P0001  ;
	input \u4_dout_reg[9]/P0001  ;
	input \u4_funct_adr_reg[0]/P0001  ;
	input \u4_funct_adr_reg[1]/P0001  ;
	input \u4_funct_adr_reg[2]/P0001  ;
	input \u4_funct_adr_reg[3]/P0001  ;
	input \u4_funct_adr_reg[4]/P0001  ;
	input \u4_funct_adr_reg[5]/P0001  ;
	input \u4_funct_adr_reg[6]/P0001  ;
	input \u4_int_src_re_reg/P0001  ;
	input \u4_int_srca_reg[0]/P0001  ;
	input \u4_int_srca_reg[1]/P0001  ;
	input \u4_int_srca_reg[2]/P0001  ;
	input \u4_int_srca_reg[3]/P0001  ;
	input \u4_int_srcb_reg[0]/P0001  ;
	input \u4_int_srcb_reg[1]/P0001  ;
	input \u4_int_srcb_reg[2]/P0001  ;
	input \u4_int_srcb_reg[3]/P0001  ;
	input \u4_int_srcb_reg[4]/P0001  ;
	input \u4_int_srcb_reg[5]/P0001  ;
	input \u4_int_srcb_reg[6]/P0001  ;
	input \u4_int_srcb_reg[7]/P0001  ;
	input \u4_int_srcb_reg[8]/P0001  ;
	input \u4_inta_msk_reg[0]/P0001  ;
	input \u4_inta_msk_reg[1]/P0001  ;
	input \u4_inta_msk_reg[2]/P0001  ;
	input \u4_inta_msk_reg[3]/P0001  ;
	input \u4_inta_msk_reg[4]/P0001  ;
	input \u4_inta_msk_reg[5]/P0001  ;
	input \u4_inta_msk_reg[6]/P0001  ;
	input \u4_inta_msk_reg[7]/P0001  ;
	input \u4_inta_msk_reg[8]/P0001  ;
	input \u4_intb_msk_reg[0]/P0001  ;
	input \u4_intb_msk_reg[1]/P0001  ;
	input \u4_intb_msk_reg[2]/P0001  ;
	input \u4_intb_msk_reg[3]/P0001  ;
	input \u4_intb_msk_reg[4]/P0001  ;
	input \u4_intb_msk_reg[5]/P0001  ;
	input \u4_intb_msk_reg[6]/P0001  ;
	input \u4_intb_msk_reg[7]/P0001  ;
	input \u4_intb_msk_reg[8]/P0001  ;
	input \u4_match_r1_reg/P0001  ;
	input \u4_nse_err_r_reg/P0001  ;
	input \u4_pid_cs_err_r_reg/P0001  ;
	input \u4_rx_err_r_reg/P0001  ;
	input \u4_suspend_r1_reg/P0001  ;
	input \u4_u0_buf0_orig_m3_reg[0]/P0001  ;
	input \u4_u0_buf0_orig_m3_reg[10]/P0001  ;
	input \u4_u0_buf0_orig_m3_reg[11]/P0001  ;
	input \u4_u0_buf0_orig_m3_reg[1]/P0001  ;
	input \u4_u0_buf0_orig_m3_reg[2]/P0001  ;
	input \u4_u0_buf0_orig_m3_reg[3]/P0001  ;
	input \u4_u0_buf0_orig_m3_reg[4]/P0001  ;
	input \u4_u0_buf0_orig_m3_reg[5]/P0001  ;
	input \u4_u0_buf0_orig_m3_reg[6]/P0001  ;
	input \u4_u0_buf0_orig_m3_reg[7]/P0001  ;
	input \u4_u0_buf0_orig_m3_reg[8]/P0001  ;
	input \u4_u0_buf0_orig_m3_reg[9]/P0001  ;
	input \u4_u0_buf0_orig_reg[0]/P0001  ;
	input \u4_u0_buf0_orig_reg[10]/P0001  ;
	input \u4_u0_buf0_orig_reg[11]/P0001  ;
	input \u4_u0_buf0_orig_reg[12]/P0001  ;
	input \u4_u0_buf0_orig_reg[13]/P0001  ;
	input \u4_u0_buf0_orig_reg[14]/P0001  ;
	input \u4_u0_buf0_orig_reg[15]/P0001  ;
	input \u4_u0_buf0_orig_reg[16]/P0001  ;
	input \u4_u0_buf0_orig_reg[17]/P0001  ;
	input \u4_u0_buf0_orig_reg[18]/P0001  ;
	input \u4_u0_buf0_orig_reg[19]/P0001  ;
	input \u4_u0_buf0_orig_reg[1]/P0001  ;
	input \u4_u0_buf0_orig_reg[20]/P0001  ;
	input \u4_u0_buf0_orig_reg[21]/P0001  ;
	input \u4_u0_buf0_orig_reg[22]/P0001  ;
	input \u4_u0_buf0_orig_reg[23]/P0001  ;
	input \u4_u0_buf0_orig_reg[24]/P0001  ;
	input \u4_u0_buf0_orig_reg[25]/P0001  ;
	input \u4_u0_buf0_orig_reg[26]/P0001  ;
	input \u4_u0_buf0_orig_reg[27]/P0001  ;
	input \u4_u0_buf0_orig_reg[28]/P0001  ;
	input \u4_u0_buf0_orig_reg[29]/NET0131  ;
	input \u4_u0_buf0_orig_reg[2]/P0001  ;
	input \u4_u0_buf0_orig_reg[30]/NET0131  ;
	input \u4_u0_buf0_orig_reg[31]/P0001  ;
	input \u4_u0_buf0_orig_reg[3]/P0001  ;
	input \u4_u0_buf0_orig_reg[4]/P0001  ;
	input \u4_u0_buf0_orig_reg[5]/P0001  ;
	input \u4_u0_buf0_orig_reg[6]/P0001  ;
	input \u4_u0_buf0_orig_reg[7]/P0001  ;
	input \u4_u0_buf0_orig_reg[8]/P0001  ;
	input \u4_u0_buf0_orig_reg[9]/P0001  ;
	input \u4_u0_buf0_reg[0]/P0001  ;
	input \u4_u0_buf0_reg[10]/P0001  ;
	input \u4_u0_buf0_reg[11]/P0001  ;
	input \u4_u0_buf0_reg[12]/P0001  ;
	input \u4_u0_buf0_reg[13]/P0001  ;
	input \u4_u0_buf0_reg[14]/P0001  ;
	input \u4_u0_buf0_reg[15]/P0001  ;
	input \u4_u0_buf0_reg[16]/P0001  ;
	input \u4_u0_buf0_reg[17]/P0001  ;
	input \u4_u0_buf0_reg[18]/P0001  ;
	input \u4_u0_buf0_reg[19]/P0001  ;
	input \u4_u0_buf0_reg[1]/P0001  ;
	input \u4_u0_buf0_reg[20]/P0001  ;
	input \u4_u0_buf0_reg[21]/P0001  ;
	input \u4_u0_buf0_reg[22]/P0001  ;
	input \u4_u0_buf0_reg[23]/P0001  ;
	input \u4_u0_buf0_reg[24]/P0001  ;
	input \u4_u0_buf0_reg[25]/P0001  ;
	input \u4_u0_buf0_reg[26]/P0001  ;
	input \u4_u0_buf0_reg[27]/P0001  ;
	input \u4_u0_buf0_reg[28]/P0001  ;
	input \u4_u0_buf0_reg[29]/P0001  ;
	input \u4_u0_buf0_reg[2]/P0001  ;
	input \u4_u0_buf0_reg[30]/P0001  ;
	input \u4_u0_buf0_reg[31]/P0001  ;
	input \u4_u0_buf0_reg[3]/P0001  ;
	input \u4_u0_buf0_reg[4]/P0001  ;
	input \u4_u0_buf0_reg[5]/P0001  ;
	input \u4_u0_buf0_reg[6]/P0001  ;
	input \u4_u0_buf0_reg[7]/P0001  ;
	input \u4_u0_buf0_reg[8]/P0001  ;
	input \u4_u0_buf0_reg[9]/P0001  ;
	input \u4_u0_buf1_reg[0]/P0001  ;
	input \u4_u0_buf1_reg[10]/P0001  ;
	input \u4_u0_buf1_reg[11]/P0001  ;
	input \u4_u0_buf1_reg[12]/P0001  ;
	input \u4_u0_buf1_reg[13]/P0001  ;
	input \u4_u0_buf1_reg[14]/P0001  ;
	input \u4_u0_buf1_reg[15]/P0001  ;
	input \u4_u0_buf1_reg[16]/P0001  ;
	input \u4_u0_buf1_reg[17]/P0001  ;
	input \u4_u0_buf1_reg[18]/P0001  ;
	input \u4_u0_buf1_reg[19]/P0001  ;
	input \u4_u0_buf1_reg[1]/P0001  ;
	input \u4_u0_buf1_reg[20]/P0001  ;
	input \u4_u0_buf1_reg[21]/P0001  ;
	input \u4_u0_buf1_reg[22]/P0001  ;
	input \u4_u0_buf1_reg[23]/P0001  ;
	input \u4_u0_buf1_reg[24]/P0001  ;
	input \u4_u0_buf1_reg[25]/P0001  ;
	input \u4_u0_buf1_reg[26]/P0001  ;
	input \u4_u0_buf1_reg[27]/P0001  ;
	input \u4_u0_buf1_reg[28]/P0001  ;
	input \u4_u0_buf1_reg[29]/P0001  ;
	input \u4_u0_buf1_reg[2]/P0001  ;
	input \u4_u0_buf1_reg[30]/P0001  ;
	input \u4_u0_buf1_reg[31]/P0001  ;
	input \u4_u0_buf1_reg[3]/P0001  ;
	input \u4_u0_buf1_reg[4]/P0001  ;
	input \u4_u0_buf1_reg[5]/P0001  ;
	input \u4_u0_buf1_reg[6]/P0001  ;
	input \u4_u0_buf1_reg[7]/P0001  ;
	input \u4_u0_buf1_reg[8]/P0001  ;
	input \u4_u0_buf1_reg[9]/P0001  ;
	input \u4_u0_csr0_reg[0]/P0001  ;
	input \u4_u0_csr0_reg[10]/P0001  ;
	input \u4_u0_csr0_reg[11]/P0001  ;
	input \u4_u0_csr0_reg[12]/P0001  ;
	input \u4_u0_csr0_reg[1]/P0001  ;
	input \u4_u0_csr0_reg[2]/P0001  ;
	input \u4_u0_csr0_reg[3]/NET0131  ;
	input \u4_u0_csr0_reg[4]/P0001  ;
	input \u4_u0_csr0_reg[5]/P0001  ;
	input \u4_u0_csr0_reg[6]/P0001  ;
	input \u4_u0_csr0_reg[7]/P0001  ;
	input \u4_u0_csr0_reg[8]/P0001  ;
	input \u4_u0_csr0_reg[9]/P0001  ;
	input \u4_u0_csr1_reg[0]/P0001  ;
	input \u4_u0_csr1_reg[10]/P0001  ;
	input \u4_u0_csr1_reg[11]/P0001  ;
	input \u4_u0_csr1_reg[12]/P0001  ;
	input \u4_u0_csr1_reg[1]/P0001  ;
	input \u4_u0_csr1_reg[2]/P0001  ;
	input \u4_u0_csr1_reg[3]/P0001  ;
	input \u4_u0_csr1_reg[4]/P0001  ;
	input \u4_u0_csr1_reg[5]/P0001  ;
	input \u4_u0_csr1_reg[6]/P0001  ;
	input \u4_u0_csr1_reg[7]/P0001  ;
	input \u4_u0_csr1_reg[8]/P0001  ;
	input \u4_u0_csr1_reg[9]/P0001  ;
	input \u4_u0_dma_ack_clr1_reg/P0001  ;
	input \u4_u0_dma_ack_wr1_reg/P0001  ;
	input \u4_u0_dma_in_buf_sz1_reg/P0001  ;
	input \u4_u0_dma_in_cnt_reg[0]/P0001  ;
	input \u4_u0_dma_in_cnt_reg[10]/P0001  ;
	input \u4_u0_dma_in_cnt_reg[11]/P0001  ;
	input \u4_u0_dma_in_cnt_reg[1]/P0001  ;
	input \u4_u0_dma_in_cnt_reg[2]/P0001  ;
	input \u4_u0_dma_in_cnt_reg[3]/P0001  ;
	input \u4_u0_dma_in_cnt_reg[4]/P0001  ;
	input \u4_u0_dma_in_cnt_reg[5]/P0001  ;
	input \u4_u0_dma_in_cnt_reg[6]/P0001  ;
	input \u4_u0_dma_in_cnt_reg[7]/P0001  ;
	input \u4_u0_dma_in_cnt_reg[8]/P0001  ;
	input \u4_u0_dma_in_cnt_reg[9]/P0001  ;
	input \u4_u0_dma_out_buf_avail_reg/P0001  ;
	input \u4_u0_dma_out_cnt_reg[10]/P0001  ;
	input \u4_u0_dma_out_cnt_reg[11]/P0001  ;
	input \u4_u0_dma_out_cnt_reg[1]/P0001  ;
	input \u4_u0_dma_out_cnt_reg[2]/P0001  ;
	input \u4_u0_dma_out_cnt_reg[3]/P0001  ;
	input \u4_u0_dma_out_cnt_reg[4]/P0001  ;
	input \u4_u0_dma_out_cnt_reg[5]/P0001  ;
	input \u4_u0_dma_out_cnt_reg[6]/P0001  ;
	input \u4_u0_dma_out_cnt_reg[7]/P0001  ;
	input \u4_u0_dma_out_cnt_reg[8]/P0001  ;
	input \u4_u0_dma_out_cnt_reg[9]/P0001  ;
	input \u4_u0_dma_out_left_reg[0]/P0001  ;
	input \u4_u0_dma_out_left_reg[10]/P0001  ;
	input \u4_u0_dma_out_left_reg[11]/P0001  ;
	input \u4_u0_dma_out_left_reg[1]/P0001  ;
	input \u4_u0_dma_out_left_reg[2]/P0001  ;
	input \u4_u0_dma_out_left_reg[3]/P0001  ;
	input \u4_u0_dma_out_left_reg[4]/P0001  ;
	input \u4_u0_dma_out_left_reg[5]/P0001  ;
	input \u4_u0_dma_out_left_reg[6]/P0001  ;
	input \u4_u0_dma_out_left_reg[7]/P0001  ;
	input \u4_u0_dma_out_left_reg[8]/P0001  ;
	input \u4_u0_dma_out_left_reg[9]/P0001  ;
	input \u4_u0_dma_req_in_hold2_reg/P0001  ;
	input \u4_u0_dma_req_in_hold_reg/P0001  ;
	input \u4_u0_dma_req_out_hold_reg/P0001  ;
	input \u4_u0_ep_match_r_reg/P0001  ;
	input \u4_u0_iena_reg[0]/P0001  ;
	input \u4_u0_iena_reg[1]/P0001  ;
	input \u4_u0_iena_reg[2]/P0001  ;
	input \u4_u0_iena_reg[3]/P0001  ;
	input \u4_u0_iena_reg[4]/P0001  ;
	input \u4_u0_iena_reg[5]/P0001  ;
	input \u4_u0_ienb_reg[0]/P0001  ;
	input \u4_u0_ienb_reg[1]/P0001  ;
	input \u4_u0_ienb_reg[2]/P0001  ;
	input \u4_u0_ienb_reg[3]/P0001  ;
	input \u4_u0_ienb_reg[4]/P0001  ;
	input \u4_u0_ienb_reg[5]/P0001  ;
	input \u4_u0_int_re_reg/P0001  ;
	input \u4_u0_int_stat_reg[0]/P0001  ;
	input \u4_u0_int_stat_reg[1]/P0001  ;
	input \u4_u0_int_stat_reg[2]/P0001  ;
	input \u4_u0_int_stat_reg[3]/P0001  ;
	input \u4_u0_int_stat_reg[4]/P0001  ;
	input \u4_u0_int_stat_reg[5]/P0001  ;
	input \u4_u0_int_stat_reg[6]/P0001  ;
	input \u4_u0_inta_reg/P0001  ;
	input \u4_u0_intb_reg/P0001  ;
	input \u4_u0_ots_stop_reg/P0001  ;
	input \u4_u0_r1_reg/P0001  ;
	input \u4_u0_r2_reg/P0001  ;
	input \u4_u0_r4_reg/P0001  ;
	input \u4_u0_r5_reg/NET0131  ;
	input \u4_u0_set_r_reg/P0001  ;
	input \u4_u0_uc_bsel_reg[0]/P0001  ;
	input \u4_u0_uc_bsel_reg[1]/P0001  ;
	input \u4_u0_uc_dpd_reg[0]/P0001  ;
	input \u4_u0_uc_dpd_reg[1]/P0001  ;
	input \u4_u1_buf0_orig_m3_reg[0]/P0001  ;
	input \u4_u1_buf0_orig_m3_reg[10]/P0001  ;
	input \u4_u1_buf0_orig_m3_reg[11]/P0001  ;
	input \u4_u1_buf0_orig_m3_reg[1]/P0001  ;
	input \u4_u1_buf0_orig_m3_reg[2]/P0001  ;
	input \u4_u1_buf0_orig_m3_reg[3]/P0001  ;
	input \u4_u1_buf0_orig_m3_reg[4]/P0001  ;
	input \u4_u1_buf0_orig_m3_reg[5]/P0001  ;
	input \u4_u1_buf0_orig_m3_reg[6]/P0001  ;
	input \u4_u1_buf0_orig_m3_reg[7]/P0001  ;
	input \u4_u1_buf0_orig_m3_reg[8]/P0001  ;
	input \u4_u1_buf0_orig_m3_reg[9]/P0001  ;
	input \u4_u1_buf0_orig_reg[0]/P0001  ;
	input \u4_u1_buf0_orig_reg[10]/P0001  ;
	input \u4_u1_buf0_orig_reg[11]/P0001  ;
	input \u4_u1_buf0_orig_reg[12]/P0001  ;
	input \u4_u1_buf0_orig_reg[13]/P0001  ;
	input \u4_u1_buf0_orig_reg[14]/P0001  ;
	input \u4_u1_buf0_orig_reg[15]/P0001  ;
	input \u4_u1_buf0_orig_reg[16]/P0001  ;
	input \u4_u1_buf0_orig_reg[17]/P0001  ;
	input \u4_u1_buf0_orig_reg[18]/P0001  ;
	input \u4_u1_buf0_orig_reg[19]/P0001  ;
	input \u4_u1_buf0_orig_reg[1]/P0001  ;
	input \u4_u1_buf0_orig_reg[20]/P0001  ;
	input \u4_u1_buf0_orig_reg[21]/P0001  ;
	input \u4_u1_buf0_orig_reg[22]/P0001  ;
	input \u4_u1_buf0_orig_reg[23]/P0001  ;
	input \u4_u1_buf0_orig_reg[24]/P0001  ;
	input \u4_u1_buf0_orig_reg[25]/P0001  ;
	input \u4_u1_buf0_orig_reg[26]/P0001  ;
	input \u4_u1_buf0_orig_reg[27]/P0001  ;
	input \u4_u1_buf0_orig_reg[28]/P0001  ;
	input \u4_u1_buf0_orig_reg[29]/NET0131  ;
	input \u4_u1_buf0_orig_reg[2]/P0001  ;
	input \u4_u1_buf0_orig_reg[30]/NET0131  ;
	input \u4_u1_buf0_orig_reg[31]/P0001  ;
	input \u4_u1_buf0_orig_reg[3]/P0001  ;
	input \u4_u1_buf0_orig_reg[4]/P0001  ;
	input \u4_u1_buf0_orig_reg[5]/P0001  ;
	input \u4_u1_buf0_orig_reg[6]/P0001  ;
	input \u4_u1_buf0_orig_reg[7]/P0001  ;
	input \u4_u1_buf0_orig_reg[8]/P0001  ;
	input \u4_u1_buf0_orig_reg[9]/P0001  ;
	input \u4_u1_buf0_reg[0]/P0001  ;
	input \u4_u1_buf0_reg[10]/P0001  ;
	input \u4_u1_buf0_reg[11]/P0001  ;
	input \u4_u1_buf0_reg[12]/P0001  ;
	input \u4_u1_buf0_reg[13]/P0001  ;
	input \u4_u1_buf0_reg[14]/P0001  ;
	input \u4_u1_buf0_reg[15]/P0001  ;
	input \u4_u1_buf0_reg[16]/P0001  ;
	input \u4_u1_buf0_reg[17]/P0001  ;
	input \u4_u1_buf0_reg[18]/P0001  ;
	input \u4_u1_buf0_reg[19]/P0001  ;
	input \u4_u1_buf0_reg[1]/P0001  ;
	input \u4_u1_buf0_reg[20]/P0001  ;
	input \u4_u1_buf0_reg[21]/P0001  ;
	input \u4_u1_buf0_reg[22]/P0001  ;
	input \u4_u1_buf0_reg[23]/P0001  ;
	input \u4_u1_buf0_reg[24]/P0001  ;
	input \u4_u1_buf0_reg[25]/P0001  ;
	input \u4_u1_buf0_reg[26]/P0001  ;
	input \u4_u1_buf0_reg[27]/P0001  ;
	input \u4_u1_buf0_reg[28]/P0001  ;
	input \u4_u1_buf0_reg[29]/P0001  ;
	input \u4_u1_buf0_reg[2]/P0001  ;
	input \u4_u1_buf0_reg[30]/P0001  ;
	input \u4_u1_buf0_reg[31]/P0001  ;
	input \u4_u1_buf0_reg[3]/P0001  ;
	input \u4_u1_buf0_reg[4]/P0001  ;
	input \u4_u1_buf0_reg[5]/P0001  ;
	input \u4_u1_buf0_reg[6]/P0001  ;
	input \u4_u1_buf0_reg[7]/P0001  ;
	input \u4_u1_buf0_reg[8]/P0001  ;
	input \u4_u1_buf0_reg[9]/P0001  ;
	input \u4_u1_buf1_reg[0]/P0001  ;
	input \u4_u1_buf1_reg[10]/P0001  ;
	input \u4_u1_buf1_reg[11]/P0001  ;
	input \u4_u1_buf1_reg[12]/P0001  ;
	input \u4_u1_buf1_reg[13]/P0001  ;
	input \u4_u1_buf1_reg[14]/P0001  ;
	input \u4_u1_buf1_reg[15]/P0001  ;
	input \u4_u1_buf1_reg[16]/P0001  ;
	input \u4_u1_buf1_reg[17]/P0001  ;
	input \u4_u1_buf1_reg[18]/P0001  ;
	input \u4_u1_buf1_reg[19]/P0001  ;
	input \u4_u1_buf1_reg[1]/P0001  ;
	input \u4_u1_buf1_reg[20]/P0001  ;
	input \u4_u1_buf1_reg[21]/P0001  ;
	input \u4_u1_buf1_reg[22]/P0001  ;
	input \u4_u1_buf1_reg[23]/P0001  ;
	input \u4_u1_buf1_reg[24]/P0001  ;
	input \u4_u1_buf1_reg[25]/P0001  ;
	input \u4_u1_buf1_reg[26]/P0001  ;
	input \u4_u1_buf1_reg[27]/P0001  ;
	input \u4_u1_buf1_reg[28]/P0001  ;
	input \u4_u1_buf1_reg[29]/P0001  ;
	input \u4_u1_buf1_reg[2]/P0001  ;
	input \u4_u1_buf1_reg[30]/P0001  ;
	input \u4_u1_buf1_reg[31]/P0001  ;
	input \u4_u1_buf1_reg[3]/P0001  ;
	input \u4_u1_buf1_reg[4]/P0001  ;
	input \u4_u1_buf1_reg[5]/P0001  ;
	input \u4_u1_buf1_reg[6]/P0001  ;
	input \u4_u1_buf1_reg[7]/P0001  ;
	input \u4_u1_buf1_reg[8]/P0001  ;
	input \u4_u1_buf1_reg[9]/P0001  ;
	input \u4_u1_csr0_reg[0]/P0001  ;
	input \u4_u1_csr0_reg[10]/P0001  ;
	input \u4_u1_csr0_reg[11]/P0001  ;
	input \u4_u1_csr0_reg[12]/P0001  ;
	input \u4_u1_csr0_reg[1]/P0001  ;
	input \u4_u1_csr0_reg[2]/P0001  ;
	input \u4_u1_csr0_reg[3]/NET0131  ;
	input \u4_u1_csr0_reg[4]/P0001  ;
	input \u4_u1_csr0_reg[5]/P0001  ;
	input \u4_u1_csr0_reg[6]/P0001  ;
	input \u4_u1_csr0_reg[7]/P0001  ;
	input \u4_u1_csr0_reg[8]/P0001  ;
	input \u4_u1_csr0_reg[9]/P0001  ;
	input \u4_u1_csr1_reg[0]/P0001  ;
	input \u4_u1_csr1_reg[10]/P0001  ;
	input \u4_u1_csr1_reg[11]/P0001  ;
	input \u4_u1_csr1_reg[12]/P0001  ;
	input \u4_u1_csr1_reg[1]/P0001  ;
	input \u4_u1_csr1_reg[2]/P0001  ;
	input \u4_u1_csr1_reg[3]/P0001  ;
	input \u4_u1_csr1_reg[4]/P0001  ;
	input \u4_u1_csr1_reg[5]/P0001  ;
	input \u4_u1_csr1_reg[6]/P0001  ;
	input \u4_u1_csr1_reg[7]/P0001  ;
	input \u4_u1_csr1_reg[8]/P0001  ;
	input \u4_u1_csr1_reg[9]/P0001  ;
	input \u4_u1_dma_ack_clr1_reg/P0001  ;
	input \u4_u1_dma_ack_wr1_reg/P0001  ;
	input \u4_u1_dma_in_buf_sz1_reg/P0001  ;
	input \u4_u1_dma_in_cnt_reg[0]/P0001  ;
	input \u4_u1_dma_in_cnt_reg[10]/P0001  ;
	input \u4_u1_dma_in_cnt_reg[11]/P0001  ;
	input \u4_u1_dma_in_cnt_reg[1]/P0001  ;
	input \u4_u1_dma_in_cnt_reg[2]/P0001  ;
	input \u4_u1_dma_in_cnt_reg[3]/P0001  ;
	input \u4_u1_dma_in_cnt_reg[4]/P0001  ;
	input \u4_u1_dma_in_cnt_reg[5]/P0001  ;
	input \u4_u1_dma_in_cnt_reg[6]/P0001  ;
	input \u4_u1_dma_in_cnt_reg[7]/P0001  ;
	input \u4_u1_dma_in_cnt_reg[8]/P0001  ;
	input \u4_u1_dma_in_cnt_reg[9]/P0001  ;
	input \u4_u1_dma_out_buf_avail_reg/P0001  ;
	input \u4_u1_dma_out_cnt_reg[10]/P0001  ;
	input \u4_u1_dma_out_cnt_reg[11]/P0001  ;
	input \u4_u1_dma_out_cnt_reg[1]/P0001  ;
	input \u4_u1_dma_out_cnt_reg[2]/P0001  ;
	input \u4_u1_dma_out_cnt_reg[3]/P0001  ;
	input \u4_u1_dma_out_cnt_reg[4]/P0001  ;
	input \u4_u1_dma_out_cnt_reg[5]/P0001  ;
	input \u4_u1_dma_out_cnt_reg[6]/P0001  ;
	input \u4_u1_dma_out_cnt_reg[7]/P0001  ;
	input \u4_u1_dma_out_cnt_reg[8]/P0001  ;
	input \u4_u1_dma_out_cnt_reg[9]/P0001  ;
	input \u4_u1_dma_out_left_reg[0]/P0001  ;
	input \u4_u1_dma_out_left_reg[10]/P0001  ;
	input \u4_u1_dma_out_left_reg[11]/P0001  ;
	input \u4_u1_dma_out_left_reg[1]/P0001  ;
	input \u4_u1_dma_out_left_reg[2]/P0001  ;
	input \u4_u1_dma_out_left_reg[3]/P0001  ;
	input \u4_u1_dma_out_left_reg[4]/P0001  ;
	input \u4_u1_dma_out_left_reg[5]/P0001  ;
	input \u4_u1_dma_out_left_reg[6]/P0001  ;
	input \u4_u1_dma_out_left_reg[7]/P0001  ;
	input \u4_u1_dma_out_left_reg[8]/P0001  ;
	input \u4_u1_dma_out_left_reg[9]/P0001  ;
	input \u4_u1_dma_req_in_hold2_reg/P0001  ;
	input \u4_u1_dma_req_in_hold_reg/P0001  ;
	input \u4_u1_dma_req_out_hold_reg/P0001  ;
	input \u4_u1_ep_match_r_reg/P0001  ;
	input \u4_u1_iena_reg[0]/P0001  ;
	input \u4_u1_iena_reg[1]/P0001  ;
	input \u4_u1_iena_reg[2]/P0001  ;
	input \u4_u1_iena_reg[3]/P0001  ;
	input \u4_u1_iena_reg[4]/P0001  ;
	input \u4_u1_iena_reg[5]/P0001  ;
	input \u4_u1_ienb_reg[0]/P0001  ;
	input \u4_u1_ienb_reg[1]/P0001  ;
	input \u4_u1_ienb_reg[2]/P0001  ;
	input \u4_u1_ienb_reg[3]/P0001  ;
	input \u4_u1_ienb_reg[4]/P0001  ;
	input \u4_u1_ienb_reg[5]/P0001  ;
	input \u4_u1_int_re_reg/P0001  ;
	input \u4_u1_int_stat_reg[0]/P0001  ;
	input \u4_u1_int_stat_reg[1]/P0001  ;
	input \u4_u1_int_stat_reg[2]/P0001  ;
	input \u4_u1_int_stat_reg[3]/P0001  ;
	input \u4_u1_int_stat_reg[4]/P0001  ;
	input \u4_u1_int_stat_reg[5]/P0001  ;
	input \u4_u1_int_stat_reg[6]/P0001  ;
	input \u4_u1_inta_reg/P0001  ;
	input \u4_u1_intb_reg/P0001  ;
	input \u4_u1_ots_stop_reg/P0001  ;
	input \u4_u1_r1_reg/P0001  ;
	input \u4_u1_r2_reg/P0001  ;
	input \u4_u1_r4_reg/P0001  ;
	input \u4_u1_r5_reg/NET0131  ;
	input \u4_u1_set_r_reg/P0001  ;
	input \u4_u1_uc_bsel_reg[0]/P0001  ;
	input \u4_u1_uc_bsel_reg[1]/P0001  ;
	input \u4_u1_uc_dpd_reg[0]/P0001  ;
	input \u4_u1_uc_dpd_reg[1]/P0001  ;
	input \u4_u2_buf0_orig_m3_reg[0]/P0001  ;
	input \u4_u2_buf0_orig_m3_reg[10]/P0001  ;
	input \u4_u2_buf0_orig_m3_reg[11]/P0001  ;
	input \u4_u2_buf0_orig_m3_reg[1]/P0001  ;
	input \u4_u2_buf0_orig_m3_reg[2]/P0001  ;
	input \u4_u2_buf0_orig_m3_reg[3]/P0001  ;
	input \u4_u2_buf0_orig_m3_reg[4]/P0001  ;
	input \u4_u2_buf0_orig_m3_reg[5]/P0001  ;
	input \u4_u2_buf0_orig_m3_reg[6]/P0001  ;
	input \u4_u2_buf0_orig_m3_reg[7]/P0001  ;
	input \u4_u2_buf0_orig_m3_reg[8]/P0001  ;
	input \u4_u2_buf0_orig_m3_reg[9]/P0001  ;
	input \u4_u2_buf0_orig_reg[0]/P0001  ;
	input \u4_u2_buf0_orig_reg[10]/P0001  ;
	input \u4_u2_buf0_orig_reg[11]/P0001  ;
	input \u4_u2_buf0_orig_reg[12]/P0001  ;
	input \u4_u2_buf0_orig_reg[13]/P0001  ;
	input \u4_u2_buf0_orig_reg[14]/P0001  ;
	input \u4_u2_buf0_orig_reg[15]/P0001  ;
	input \u4_u2_buf0_orig_reg[16]/P0001  ;
	input \u4_u2_buf0_orig_reg[17]/P0001  ;
	input \u4_u2_buf0_orig_reg[18]/P0001  ;
	input \u4_u2_buf0_orig_reg[19]/P0001  ;
	input \u4_u2_buf0_orig_reg[1]/P0001  ;
	input \u4_u2_buf0_orig_reg[20]/P0001  ;
	input \u4_u2_buf0_orig_reg[21]/P0001  ;
	input \u4_u2_buf0_orig_reg[22]/P0001  ;
	input \u4_u2_buf0_orig_reg[23]/P0001  ;
	input \u4_u2_buf0_orig_reg[24]/P0001  ;
	input \u4_u2_buf0_orig_reg[25]/P0001  ;
	input \u4_u2_buf0_orig_reg[26]/P0001  ;
	input \u4_u2_buf0_orig_reg[27]/P0001  ;
	input \u4_u2_buf0_orig_reg[28]/P0001  ;
	input \u4_u2_buf0_orig_reg[29]/NET0131  ;
	input \u4_u2_buf0_orig_reg[2]/P0001  ;
	input \u4_u2_buf0_orig_reg[30]/NET0131  ;
	input \u4_u2_buf0_orig_reg[31]/P0001  ;
	input \u4_u2_buf0_orig_reg[3]/P0001  ;
	input \u4_u2_buf0_orig_reg[4]/P0001  ;
	input \u4_u2_buf0_orig_reg[5]/P0001  ;
	input \u4_u2_buf0_orig_reg[6]/P0001  ;
	input \u4_u2_buf0_orig_reg[7]/P0001  ;
	input \u4_u2_buf0_orig_reg[8]/P0001  ;
	input \u4_u2_buf0_orig_reg[9]/P0001  ;
	input \u4_u2_buf0_reg[0]/P0001  ;
	input \u4_u2_buf0_reg[10]/P0001  ;
	input \u4_u2_buf0_reg[11]/P0001  ;
	input \u4_u2_buf0_reg[12]/P0001  ;
	input \u4_u2_buf0_reg[13]/P0001  ;
	input \u4_u2_buf0_reg[14]/P0001  ;
	input \u4_u2_buf0_reg[15]/P0001  ;
	input \u4_u2_buf0_reg[16]/P0001  ;
	input \u4_u2_buf0_reg[17]/P0001  ;
	input \u4_u2_buf0_reg[18]/P0001  ;
	input \u4_u2_buf0_reg[19]/P0001  ;
	input \u4_u2_buf0_reg[1]/P0001  ;
	input \u4_u2_buf0_reg[20]/P0001  ;
	input \u4_u2_buf0_reg[21]/P0001  ;
	input \u4_u2_buf0_reg[22]/P0001  ;
	input \u4_u2_buf0_reg[23]/P0001  ;
	input \u4_u2_buf0_reg[24]/P0001  ;
	input \u4_u2_buf0_reg[25]/P0001  ;
	input \u4_u2_buf0_reg[26]/P0001  ;
	input \u4_u2_buf0_reg[27]/P0001  ;
	input \u4_u2_buf0_reg[28]/P0001  ;
	input \u4_u2_buf0_reg[29]/P0001  ;
	input \u4_u2_buf0_reg[2]/P0001  ;
	input \u4_u2_buf0_reg[30]/P0001  ;
	input \u4_u2_buf0_reg[31]/P0001  ;
	input \u4_u2_buf0_reg[3]/P0001  ;
	input \u4_u2_buf0_reg[4]/P0001  ;
	input \u4_u2_buf0_reg[5]/P0001  ;
	input \u4_u2_buf0_reg[6]/P0001  ;
	input \u4_u2_buf0_reg[7]/P0001  ;
	input \u4_u2_buf0_reg[8]/P0001  ;
	input \u4_u2_buf0_reg[9]/P0001  ;
	input \u4_u2_buf1_reg[0]/P0001  ;
	input \u4_u2_buf1_reg[10]/P0001  ;
	input \u4_u2_buf1_reg[11]/P0001  ;
	input \u4_u2_buf1_reg[12]/P0001  ;
	input \u4_u2_buf1_reg[13]/P0001  ;
	input \u4_u2_buf1_reg[14]/P0001  ;
	input \u4_u2_buf1_reg[15]/P0001  ;
	input \u4_u2_buf1_reg[16]/P0001  ;
	input \u4_u2_buf1_reg[17]/P0001  ;
	input \u4_u2_buf1_reg[18]/P0001  ;
	input \u4_u2_buf1_reg[19]/P0001  ;
	input \u4_u2_buf1_reg[1]/P0001  ;
	input \u4_u2_buf1_reg[20]/P0001  ;
	input \u4_u2_buf1_reg[21]/P0001  ;
	input \u4_u2_buf1_reg[22]/P0001  ;
	input \u4_u2_buf1_reg[23]/P0001  ;
	input \u4_u2_buf1_reg[24]/P0001  ;
	input \u4_u2_buf1_reg[25]/P0001  ;
	input \u4_u2_buf1_reg[26]/P0001  ;
	input \u4_u2_buf1_reg[27]/P0001  ;
	input \u4_u2_buf1_reg[28]/P0001  ;
	input \u4_u2_buf1_reg[29]/P0001  ;
	input \u4_u2_buf1_reg[2]/P0001  ;
	input \u4_u2_buf1_reg[30]/P0001  ;
	input \u4_u2_buf1_reg[31]/P0001  ;
	input \u4_u2_buf1_reg[3]/P0001  ;
	input \u4_u2_buf1_reg[4]/P0001  ;
	input \u4_u2_buf1_reg[5]/P0001  ;
	input \u4_u2_buf1_reg[6]/P0001  ;
	input \u4_u2_buf1_reg[7]/P0001  ;
	input \u4_u2_buf1_reg[8]/P0001  ;
	input \u4_u2_buf1_reg[9]/P0001  ;
	input \u4_u2_csr0_reg[0]/P0001  ;
	input \u4_u2_csr0_reg[10]/P0001  ;
	input \u4_u2_csr0_reg[11]/P0001  ;
	input \u4_u2_csr0_reg[12]/P0001  ;
	input \u4_u2_csr0_reg[1]/P0001  ;
	input \u4_u2_csr0_reg[2]/P0001  ;
	input \u4_u2_csr0_reg[3]/NET0131  ;
	input \u4_u2_csr0_reg[4]/P0001  ;
	input \u4_u2_csr0_reg[5]/P0001  ;
	input \u4_u2_csr0_reg[6]/P0001  ;
	input \u4_u2_csr0_reg[7]/P0001  ;
	input \u4_u2_csr0_reg[8]/P0001  ;
	input \u4_u2_csr0_reg[9]/P0001  ;
	input \u4_u2_csr1_reg[0]/P0001  ;
	input \u4_u2_csr1_reg[10]/P0001  ;
	input \u4_u2_csr1_reg[11]/P0001  ;
	input \u4_u2_csr1_reg[12]/P0001  ;
	input \u4_u2_csr1_reg[1]/P0001  ;
	input \u4_u2_csr1_reg[2]/P0001  ;
	input \u4_u2_csr1_reg[3]/P0001  ;
	input \u4_u2_csr1_reg[4]/P0001  ;
	input \u4_u2_csr1_reg[5]/P0001  ;
	input \u4_u2_csr1_reg[6]/P0001  ;
	input \u4_u2_csr1_reg[7]/P0001  ;
	input \u4_u2_csr1_reg[8]/P0001  ;
	input \u4_u2_csr1_reg[9]/P0001  ;
	input \u4_u2_dma_ack_clr1_reg/P0001  ;
	input \u4_u2_dma_ack_wr1_reg/P0001  ;
	input \u4_u2_dma_in_buf_sz1_reg/P0001  ;
	input \u4_u2_dma_in_cnt_reg[0]/P0001  ;
	input \u4_u2_dma_in_cnt_reg[10]/P0001  ;
	input \u4_u2_dma_in_cnt_reg[11]/P0001  ;
	input \u4_u2_dma_in_cnt_reg[1]/P0001  ;
	input \u4_u2_dma_in_cnt_reg[2]/P0001  ;
	input \u4_u2_dma_in_cnt_reg[3]/P0001  ;
	input \u4_u2_dma_in_cnt_reg[4]/P0001  ;
	input \u4_u2_dma_in_cnt_reg[5]/P0001  ;
	input \u4_u2_dma_in_cnt_reg[6]/P0001  ;
	input \u4_u2_dma_in_cnt_reg[7]/P0001  ;
	input \u4_u2_dma_in_cnt_reg[8]/P0001  ;
	input \u4_u2_dma_in_cnt_reg[9]/P0001  ;
	input \u4_u2_dma_out_buf_avail_reg/P0001  ;
	input \u4_u2_dma_out_cnt_reg[10]/P0001  ;
	input \u4_u2_dma_out_cnt_reg[11]/P0001  ;
	input \u4_u2_dma_out_cnt_reg[1]/P0001  ;
	input \u4_u2_dma_out_cnt_reg[2]/P0001  ;
	input \u4_u2_dma_out_cnt_reg[3]/P0001  ;
	input \u4_u2_dma_out_cnt_reg[4]/P0001  ;
	input \u4_u2_dma_out_cnt_reg[5]/P0001  ;
	input \u4_u2_dma_out_cnt_reg[6]/P0001  ;
	input \u4_u2_dma_out_cnt_reg[7]/P0001  ;
	input \u4_u2_dma_out_cnt_reg[8]/P0001  ;
	input \u4_u2_dma_out_cnt_reg[9]/P0001  ;
	input \u4_u2_dma_out_left_reg[0]/P0001  ;
	input \u4_u2_dma_out_left_reg[10]/P0001  ;
	input \u4_u2_dma_out_left_reg[11]/P0001  ;
	input \u4_u2_dma_out_left_reg[1]/P0001  ;
	input \u4_u2_dma_out_left_reg[2]/P0001  ;
	input \u4_u2_dma_out_left_reg[3]/P0001  ;
	input \u4_u2_dma_out_left_reg[4]/P0001  ;
	input \u4_u2_dma_out_left_reg[5]/P0001  ;
	input \u4_u2_dma_out_left_reg[6]/P0001  ;
	input \u4_u2_dma_out_left_reg[7]/P0001  ;
	input \u4_u2_dma_out_left_reg[8]/P0001  ;
	input \u4_u2_dma_out_left_reg[9]/P0001  ;
	input \u4_u2_dma_req_in_hold2_reg/P0001  ;
	input \u4_u2_dma_req_in_hold_reg/P0001  ;
	input \u4_u2_dma_req_out_hold_reg/P0001  ;
	input \u4_u2_ep_match_r_reg/P0001  ;
	input \u4_u2_iena_reg[0]/P0001  ;
	input \u4_u2_iena_reg[1]/P0001  ;
	input \u4_u2_iena_reg[2]/P0001  ;
	input \u4_u2_iena_reg[3]/P0001  ;
	input \u4_u2_iena_reg[4]/P0001  ;
	input \u4_u2_iena_reg[5]/P0001  ;
	input \u4_u2_ienb_reg[0]/P0001  ;
	input \u4_u2_ienb_reg[1]/P0001  ;
	input \u4_u2_ienb_reg[2]/P0001  ;
	input \u4_u2_ienb_reg[3]/P0001  ;
	input \u4_u2_ienb_reg[4]/P0001  ;
	input \u4_u2_ienb_reg[5]/P0001  ;
	input \u4_u2_int_re_reg/P0001  ;
	input \u4_u2_int_stat_reg[0]/P0001  ;
	input \u4_u2_int_stat_reg[1]/P0001  ;
	input \u4_u2_int_stat_reg[2]/P0001  ;
	input \u4_u2_int_stat_reg[3]/P0001  ;
	input \u4_u2_int_stat_reg[4]/P0001  ;
	input \u4_u2_int_stat_reg[5]/P0001  ;
	input \u4_u2_int_stat_reg[6]/P0001  ;
	input \u4_u2_inta_reg/P0001  ;
	input \u4_u2_intb_reg/P0001  ;
	input \u4_u2_ots_stop_reg/P0001  ;
	input \u4_u2_r1_reg/P0001  ;
	input \u4_u2_r2_reg/P0001  ;
	input \u4_u2_r4_reg/P0001  ;
	input \u4_u2_r5_reg/NET0131  ;
	input \u4_u2_set_r_reg/P0001  ;
	input \u4_u2_uc_bsel_reg[0]/P0001  ;
	input \u4_u2_uc_bsel_reg[1]/P0001  ;
	input \u4_u2_uc_dpd_reg[0]/P0001  ;
	input \u4_u2_uc_dpd_reg[1]/P0001  ;
	input \u4_u3_buf0_orig_m3_reg[0]/P0001  ;
	input \u4_u3_buf0_orig_m3_reg[10]/P0001  ;
	input \u4_u3_buf0_orig_m3_reg[11]/P0001  ;
	input \u4_u3_buf0_orig_m3_reg[1]/P0001  ;
	input \u4_u3_buf0_orig_m3_reg[2]/P0001  ;
	input \u4_u3_buf0_orig_m3_reg[3]/P0001  ;
	input \u4_u3_buf0_orig_m3_reg[4]/P0001  ;
	input \u4_u3_buf0_orig_m3_reg[5]/P0001  ;
	input \u4_u3_buf0_orig_m3_reg[6]/P0001  ;
	input \u4_u3_buf0_orig_m3_reg[7]/P0001  ;
	input \u4_u3_buf0_orig_m3_reg[8]/P0001  ;
	input \u4_u3_buf0_orig_m3_reg[9]/P0001  ;
	input \u4_u3_buf0_orig_reg[0]/P0001  ;
	input \u4_u3_buf0_orig_reg[10]/P0001  ;
	input \u4_u3_buf0_orig_reg[11]/P0001  ;
	input \u4_u3_buf0_orig_reg[12]/P0001  ;
	input \u4_u3_buf0_orig_reg[13]/P0001  ;
	input \u4_u3_buf0_orig_reg[14]/P0001  ;
	input \u4_u3_buf0_orig_reg[15]/P0001  ;
	input \u4_u3_buf0_orig_reg[16]/P0001  ;
	input \u4_u3_buf0_orig_reg[17]/P0001  ;
	input \u4_u3_buf0_orig_reg[18]/P0001  ;
	input \u4_u3_buf0_orig_reg[19]/P0001  ;
	input \u4_u3_buf0_orig_reg[1]/P0001  ;
	input \u4_u3_buf0_orig_reg[20]/P0001  ;
	input \u4_u3_buf0_orig_reg[21]/P0001  ;
	input \u4_u3_buf0_orig_reg[22]/P0001  ;
	input \u4_u3_buf0_orig_reg[23]/P0001  ;
	input \u4_u3_buf0_orig_reg[24]/P0001  ;
	input \u4_u3_buf0_orig_reg[25]/P0001  ;
	input \u4_u3_buf0_orig_reg[26]/P0001  ;
	input \u4_u3_buf0_orig_reg[27]/P0001  ;
	input \u4_u3_buf0_orig_reg[28]/P0001  ;
	input \u4_u3_buf0_orig_reg[29]/NET0131  ;
	input \u4_u3_buf0_orig_reg[2]/P0001  ;
	input \u4_u3_buf0_orig_reg[30]/NET0131  ;
	input \u4_u3_buf0_orig_reg[31]/P0001  ;
	input \u4_u3_buf0_orig_reg[3]/P0001  ;
	input \u4_u3_buf0_orig_reg[4]/P0001  ;
	input \u4_u3_buf0_orig_reg[5]/P0001  ;
	input \u4_u3_buf0_orig_reg[6]/P0001  ;
	input \u4_u3_buf0_orig_reg[7]/P0001  ;
	input \u4_u3_buf0_orig_reg[8]/P0001  ;
	input \u4_u3_buf0_orig_reg[9]/P0001  ;
	input \u4_u3_buf0_reg[0]/P0001  ;
	input \u4_u3_buf0_reg[10]/P0001  ;
	input \u4_u3_buf0_reg[11]/P0001  ;
	input \u4_u3_buf0_reg[12]/P0001  ;
	input \u4_u3_buf0_reg[13]/P0001  ;
	input \u4_u3_buf0_reg[14]/P0001  ;
	input \u4_u3_buf0_reg[15]/P0001  ;
	input \u4_u3_buf0_reg[16]/P0001  ;
	input \u4_u3_buf0_reg[17]/P0001  ;
	input \u4_u3_buf0_reg[18]/P0001  ;
	input \u4_u3_buf0_reg[19]/P0001  ;
	input \u4_u3_buf0_reg[1]/P0001  ;
	input \u4_u3_buf0_reg[20]/P0001  ;
	input \u4_u3_buf0_reg[21]/P0001  ;
	input \u4_u3_buf0_reg[22]/P0001  ;
	input \u4_u3_buf0_reg[23]/P0001  ;
	input \u4_u3_buf0_reg[24]/P0001  ;
	input \u4_u3_buf0_reg[25]/P0001  ;
	input \u4_u3_buf0_reg[26]/P0001  ;
	input \u4_u3_buf0_reg[27]/P0001  ;
	input \u4_u3_buf0_reg[28]/P0001  ;
	input \u4_u3_buf0_reg[29]/P0001  ;
	input \u4_u3_buf0_reg[2]/P0001  ;
	input \u4_u3_buf0_reg[30]/P0001  ;
	input \u4_u3_buf0_reg[31]/P0001  ;
	input \u4_u3_buf0_reg[3]/P0001  ;
	input \u4_u3_buf0_reg[4]/P0001  ;
	input \u4_u3_buf0_reg[5]/P0001  ;
	input \u4_u3_buf0_reg[6]/P0001  ;
	input \u4_u3_buf0_reg[7]/P0001  ;
	input \u4_u3_buf0_reg[8]/P0001  ;
	input \u4_u3_buf0_reg[9]/P0001  ;
	input \u4_u3_buf1_reg[0]/P0001  ;
	input \u4_u3_buf1_reg[10]/P0001  ;
	input \u4_u3_buf1_reg[11]/P0001  ;
	input \u4_u3_buf1_reg[12]/P0001  ;
	input \u4_u3_buf1_reg[13]/P0001  ;
	input \u4_u3_buf1_reg[14]/P0001  ;
	input \u4_u3_buf1_reg[15]/P0001  ;
	input \u4_u3_buf1_reg[16]/P0001  ;
	input \u4_u3_buf1_reg[17]/P0001  ;
	input \u4_u3_buf1_reg[18]/P0001  ;
	input \u4_u3_buf1_reg[19]/P0001  ;
	input \u4_u3_buf1_reg[1]/P0001  ;
	input \u4_u3_buf1_reg[20]/P0001  ;
	input \u4_u3_buf1_reg[21]/P0001  ;
	input \u4_u3_buf1_reg[22]/P0001  ;
	input \u4_u3_buf1_reg[23]/P0001  ;
	input \u4_u3_buf1_reg[24]/P0001  ;
	input \u4_u3_buf1_reg[25]/P0001  ;
	input \u4_u3_buf1_reg[26]/P0001  ;
	input \u4_u3_buf1_reg[27]/P0001  ;
	input \u4_u3_buf1_reg[28]/P0001  ;
	input \u4_u3_buf1_reg[29]/P0001  ;
	input \u4_u3_buf1_reg[2]/P0001  ;
	input \u4_u3_buf1_reg[30]/P0001  ;
	input \u4_u3_buf1_reg[31]/P0001  ;
	input \u4_u3_buf1_reg[3]/P0001  ;
	input \u4_u3_buf1_reg[4]/P0001  ;
	input \u4_u3_buf1_reg[5]/P0001  ;
	input \u4_u3_buf1_reg[6]/P0001  ;
	input \u4_u3_buf1_reg[7]/P0001  ;
	input \u4_u3_buf1_reg[8]/P0001  ;
	input \u4_u3_buf1_reg[9]/P0001  ;
	input \u4_u3_csr0_reg[0]/P0001  ;
	input \u4_u3_csr0_reg[10]/P0001  ;
	input \u4_u3_csr0_reg[11]/P0001  ;
	input \u4_u3_csr0_reg[12]/P0001  ;
	input \u4_u3_csr0_reg[1]/P0001  ;
	input \u4_u3_csr0_reg[2]/P0001  ;
	input \u4_u3_csr0_reg[3]/NET0131  ;
	input \u4_u3_csr0_reg[4]/P0001  ;
	input \u4_u3_csr0_reg[5]/P0001  ;
	input \u4_u3_csr0_reg[6]/P0001  ;
	input \u4_u3_csr0_reg[7]/P0001  ;
	input \u4_u3_csr0_reg[8]/P0001  ;
	input \u4_u3_csr0_reg[9]/P0001  ;
	input \u4_u3_csr1_reg[0]/P0001  ;
	input \u4_u3_csr1_reg[10]/P0001  ;
	input \u4_u3_csr1_reg[11]/P0001  ;
	input \u4_u3_csr1_reg[12]/P0001  ;
	input \u4_u3_csr1_reg[1]/P0001  ;
	input \u4_u3_csr1_reg[2]/P0001  ;
	input \u4_u3_csr1_reg[3]/P0001  ;
	input \u4_u3_csr1_reg[4]/P0001  ;
	input \u4_u3_csr1_reg[5]/P0001  ;
	input \u4_u3_csr1_reg[6]/P0001  ;
	input \u4_u3_csr1_reg[7]/P0001  ;
	input \u4_u3_csr1_reg[8]/P0001  ;
	input \u4_u3_csr1_reg[9]/P0001  ;
	input \u4_u3_dma_ack_clr1_reg/P0001  ;
	input \u4_u3_dma_ack_wr1_reg/P0001  ;
	input \u4_u3_dma_in_buf_sz1_reg/P0001  ;
	input \u4_u3_dma_in_cnt_reg[0]/P0001  ;
	input \u4_u3_dma_in_cnt_reg[10]/P0001  ;
	input \u4_u3_dma_in_cnt_reg[11]/P0001  ;
	input \u4_u3_dma_in_cnt_reg[1]/P0001  ;
	input \u4_u3_dma_in_cnt_reg[2]/P0001  ;
	input \u4_u3_dma_in_cnt_reg[3]/P0001  ;
	input \u4_u3_dma_in_cnt_reg[4]/P0001  ;
	input \u4_u3_dma_in_cnt_reg[5]/P0001  ;
	input \u4_u3_dma_in_cnt_reg[6]/P0001  ;
	input \u4_u3_dma_in_cnt_reg[7]/P0001  ;
	input \u4_u3_dma_in_cnt_reg[8]/P0001  ;
	input \u4_u3_dma_in_cnt_reg[9]/P0001  ;
	input \u4_u3_dma_out_buf_avail_reg/P0001  ;
	input \u4_u3_dma_out_cnt_reg[10]/P0001  ;
	input \u4_u3_dma_out_cnt_reg[11]/P0001  ;
	input \u4_u3_dma_out_cnt_reg[1]/P0001  ;
	input \u4_u3_dma_out_cnt_reg[2]/P0001  ;
	input \u4_u3_dma_out_cnt_reg[3]/P0001  ;
	input \u4_u3_dma_out_cnt_reg[4]/P0001  ;
	input \u4_u3_dma_out_cnt_reg[5]/P0001  ;
	input \u4_u3_dma_out_cnt_reg[6]/P0001  ;
	input \u4_u3_dma_out_cnt_reg[7]/P0001  ;
	input \u4_u3_dma_out_cnt_reg[8]/P0001  ;
	input \u4_u3_dma_out_cnt_reg[9]/P0001  ;
	input \u4_u3_dma_out_left_reg[0]/P0001  ;
	input \u4_u3_dma_out_left_reg[10]/P0001  ;
	input \u4_u3_dma_out_left_reg[11]/P0001  ;
	input \u4_u3_dma_out_left_reg[1]/P0001  ;
	input \u4_u3_dma_out_left_reg[2]/P0001  ;
	input \u4_u3_dma_out_left_reg[3]/P0001  ;
	input \u4_u3_dma_out_left_reg[4]/P0001  ;
	input \u4_u3_dma_out_left_reg[5]/P0001  ;
	input \u4_u3_dma_out_left_reg[6]/P0001  ;
	input \u4_u3_dma_out_left_reg[7]/P0001  ;
	input \u4_u3_dma_out_left_reg[8]/P0001  ;
	input \u4_u3_dma_out_left_reg[9]/P0001  ;
	input \u4_u3_dma_req_in_hold2_reg/P0001  ;
	input \u4_u3_dma_req_in_hold_reg/P0001  ;
	input \u4_u3_dma_req_out_hold_reg/P0001  ;
	input \u4_u3_ep_match_r_reg/P0001  ;
	input \u4_u3_iena_reg[0]/P0001  ;
	input \u4_u3_iena_reg[1]/P0001  ;
	input \u4_u3_iena_reg[2]/P0001  ;
	input \u4_u3_iena_reg[3]/P0001  ;
	input \u4_u3_iena_reg[4]/P0001  ;
	input \u4_u3_iena_reg[5]/P0001  ;
	input \u4_u3_ienb_reg[0]/P0001  ;
	input \u4_u3_ienb_reg[1]/P0001  ;
	input \u4_u3_ienb_reg[2]/P0001  ;
	input \u4_u3_ienb_reg[3]/P0001  ;
	input \u4_u3_ienb_reg[4]/P0001  ;
	input \u4_u3_ienb_reg[5]/P0001  ;
	input \u4_u3_int_re_reg/P0001  ;
	input \u4_u3_int_stat_reg[0]/P0001  ;
	input \u4_u3_int_stat_reg[1]/P0001  ;
	input \u4_u3_int_stat_reg[2]/P0001  ;
	input \u4_u3_int_stat_reg[3]/P0001  ;
	input \u4_u3_int_stat_reg[4]/P0001  ;
	input \u4_u3_int_stat_reg[5]/P0001  ;
	input \u4_u3_int_stat_reg[6]/P0001  ;
	input \u4_u3_inta_reg/P0001  ;
	input \u4_u3_intb_reg/P0001  ;
	input \u4_u3_ots_stop_reg/P0001  ;
	input \u4_u3_r1_reg/P0001  ;
	input \u4_u3_r2_reg/P0001  ;
	input \u4_u3_r4_reg/P0001  ;
	input \u4_u3_r5_reg/NET0131  ;
	input \u4_u3_set_r_reg/P0001  ;
	input \u4_u3_uc_bsel_reg[0]/P0001  ;
	input \u4_u3_uc_bsel_reg[1]/P0001  ;
	input \u4_u3_uc_dpd_reg[0]/P0001  ;
	input \u4_u3_uc_dpd_reg[1]/P0001  ;
	input \u4_usb_reset_r_reg/P0001  ;
	input \u4_utmi_vend_ctrl_r_reg[0]/P0001  ;
	input \u4_utmi_vend_ctrl_r_reg[1]/P0001  ;
	input \u4_utmi_vend_ctrl_r_reg[2]/P0001  ;
	input \u4_utmi_vend_ctrl_r_reg[3]/P0001  ;
	input \u4_utmi_vend_stat_r_reg[0]/P0001  ;
	input \u4_utmi_vend_stat_r_reg[1]/P0001  ;
	input \u4_utmi_vend_stat_r_reg[2]/P0001  ;
	input \u4_utmi_vend_stat_r_reg[3]/P0001  ;
	input \u4_utmi_vend_stat_r_reg[4]/P0001  ;
	input \u4_utmi_vend_stat_r_reg[5]/P0001  ;
	input \u4_utmi_vend_stat_r_reg[6]/P0001  ;
	input \u4_utmi_vend_stat_r_reg[7]/P0001  ;
	input \u4_utmi_vend_wr_r_reg/P0001  ;
	input \u5_state_reg[0]/P0001  ;
	input \u5_state_reg[1]/P0001  ;
	input \u5_state_reg[2]/P0001  ;
	input \u5_state_reg[3]/P0001  ;
	input \u5_state_reg[4]/P0001  ;
	input \u5_state_reg[5]/NET0131  ;
	input \u5_wb_ack_s1_reg/P0001  ;
	input \u5_wb_ack_s2_reg/P0001  ;
	input \u5_wb_req_s1_reg/P0001  ;
	input usb_vbus_pad_i_pad ;
	input wb_ack_o_pad ;
	input \wb_addr_i[10]_pad  ;
	input \wb_addr_i[11]_pad  ;
	input \wb_addr_i[12]_pad  ;
	input \wb_addr_i[13]_pad  ;
	input \wb_addr_i[14]_pad  ;
	input \wb_addr_i[15]_pad  ;
	input \wb_addr_i[16]_pad  ;
	input \wb_addr_i[17]_pad  ;
	input \wb_addr_i[2]_pad  ;
	input \wb_addr_i[3]_pad  ;
	input \wb_addr_i[4]_pad  ;
	input \wb_addr_i[5]_pad  ;
	input \wb_addr_i[6]_pad  ;
	input \wb_addr_i[7]_pad  ;
	input \wb_addr_i[8]_pad  ;
	input \wb_addr_i[9]_pad  ;
	input wb_cyc_i_pad ;
	input \wb_data_i[0]_pad  ;
	input \wb_data_i[10]_pad  ;
	input \wb_data_i[11]_pad  ;
	input \wb_data_i[12]_pad  ;
	input \wb_data_i[13]_pad  ;
	input \wb_data_i[14]_pad  ;
	input \wb_data_i[15]_pad  ;
	input \wb_data_i[16]_pad  ;
	input \wb_data_i[17]_pad  ;
	input \wb_data_i[18]_pad  ;
	input \wb_data_i[19]_pad  ;
	input \wb_data_i[1]_pad  ;
	input \wb_data_i[20]_pad  ;
	input \wb_data_i[21]_pad  ;
	input \wb_data_i[22]_pad  ;
	input \wb_data_i[23]_pad  ;
	input \wb_data_i[24]_pad  ;
	input \wb_data_i[25]_pad  ;
	input \wb_data_i[26]_pad  ;
	input \wb_data_i[27]_pad  ;
	input \wb_data_i[28]_pad  ;
	input \wb_data_i[29]_pad  ;
	input \wb_data_i[2]_pad  ;
	input \wb_data_i[30]_pad  ;
	input \wb_data_i[31]_pad  ;
	input \wb_data_i[3]_pad  ;
	input \wb_data_i[4]_pad  ;
	input \wb_data_i[5]_pad  ;
	input \wb_data_i[6]_pad  ;
	input \wb_data_i[7]_pad  ;
	input \wb_data_i[8]_pad  ;
	input \wb_data_i[9]_pad  ;
	input wb_stb_i_pad ;
	input wb_we_i_pad ;
	output \dma_req_o[6]_pad  ;
	output \g37425/_0_  ;
	output \g37426/_0_  ;
	output \g37432/_0_  ;
	output \g37433/_0_  ;
	output \g37439/_0_  ;
	output \g37440/_0_  ;
	output \g37444/_00_  ;
	output \g37448/_0_  ;
	output \g37450/_0_  ;
	output \g37454/_0_  ;
	output \g37473/_0_  ;
	output \g37474/_0_  ;
	output \g37475/_0_  ;
	output \g37476/_0_  ;
	output \g37477/_0_  ;
	output \g37478/_0_  ;
	output \g37479/_0_  ;
	output \g37488/_0_  ;
	output \g37489/_0_  ;
	output \g37490/_0_  ;
	output \g37491/_0_  ;
	output \g37492/_0_  ;
	output \g37517/_0_  ;
	output \g37518/_0_  ;
	output \g37519/_0_  ;
	output \g37520/_0_  ;
	output \g37521/_0_  ;
	output \g37522/_0_  ;
	output \g37540/_0_  ;
	output \g37542/_0_  ;
	output \g37543/_0_  ;
	output \g37545/_0_  ;
	output \g37546/_0_  ;
	output \g37548/_0_  ;
	output \g37549/_0_  ;
	output \g37550/_0_  ;
	output \g37551/_0_  ;
	output \g37556/_0_  ;
	output \g37589/_0_  ;
	output \g37591/_0_  ;
	output \g37592/_0_  ;
	output \g37593/_0_  ;
	output \g37594/_0_  ;
	output \g37596/_0_  ;
	output \g37597/_0_  ;
	output \g37598/_0_  ;
	output \g37599/_0_  ;
	output \g37601/_0_  ;
	output \g37603/_0_  ;
	output \g37604/_0_  ;
	output \g37605/_0_  ;
	output \g37607/_0_  ;
	output \g37608/_0_  ;
	output \g37609/_0_  ;
	output \g37610/_0_  ;
	output \g37645/_0_  ;
	output \g37648/_0_  ;
	output \g37650/_0_  ;
	output \g37653/_0_  ;
	output \g37664/_3_  ;
	output \g37703/_0_  ;
	output \g37704/_0_  ;
	output \g37706/_0_  ;
	output \g37708/_0_  ;
	output \g37709/_0_  ;
	output \g37711/_0_  ;
	output \g37714/_0_  ;
	output \g37715/_0_  ;
	output \g37717/_0_  ;
	output \g37718/_0_  ;
	output \g37719/_0_  ;
	output \g37720/_0_  ;
	output \g37723/_0_  ;
	output \g37724/_0_  ;
	output \g37726/_0_  ;
	output \g37728/_0_  ;
	output \g37729/_0_  ;
	output \g37730/_0_  ;
	output \g37731/_0_  ;
	output \g37732/_0_  ;
	output \g37733/_0_  ;
	output \g37735/_0_  ;
	output \g37736/_0_  ;
	output \g37737/_0_  ;
	output \g37856/_0_  ;
	output \g37857/_0_  ;
	output \g37859/_0_  ;
	output \g37868/_0_  ;
	output \g37869/_0_  ;
	output \g37870/_0_  ;
	output \g37872/_0_  ;
	output \g37886/_0_  ;
	output \g37887/_0_  ;
	output \g37889/_0_  ;
	output \g37897/_0_  ;
	output \g37899/_0_  ;
	output \g37900/_0_  ;
	output \g37907/_0_  ;
	output \g37925/_0_  ;
	output \g37927/_0_  ;
	output \g37928/_0_  ;
	output \g37929/_0_  ;
	output \g37930/_0_  ;
	output \g37932/_0_  ;
	output \g37933/_0_  ;
	output \g37934/_0_  ;
	output \g37935/_0_  ;
	output \g37936/_0_  ;
	output \g37937/_0_  ;
	output \g37938/_0_  ;
	output \g37939/_0_  ;
	output \g37941/_0_  ;
	output \g37942/_0_  ;
	output \g37943/_0_  ;
	output \g37944/_0_  ;
	output \g37945/_0_  ;
	output \g38030/_3_  ;
	output \g38035/_0_  ;
	output \g38036/_0_  ;
	output \g38054/_0_  ;
	output \g38129/_0_  ;
	output \g38130/_0_  ;
	output \g38148/_3_  ;
	output \g38149/_3_  ;
	output \g38150/_3_  ;
	output \g38166/_0_  ;
	output \g38198/_0_  ;
	output \g38201/_0_  ;
	output \g38257/_0_  ;
	output \g38286/_0_  ;
	output \g38294/_3_  ;
	output \g38295/_3_  ;
	output \g38296/_3_  ;
	output \g38297/_3_  ;
	output \g38332/_0_  ;
	output \g38350/_0_  ;
	output \g38365/_3_  ;
	output \g38366/_3_  ;
	output \g38367/_3_  ;
	output \g38389/_0_  ;
	output \g38397/_0_  ;
	output \g38398/_0_  ;
	output \g38399/_0_  ;
	output \g38400/_0_  ;
	output \g38417/_3_  ;
	output \g38418/_3_  ;
	output \g38422/_0_  ;
	output \g38440/_0_  ;
	output \g38443/_0_  ;
	output \g38448/_3_  ;
	output \g38449/_0_  ;
	output \g38450/_0_  ;
	output \g38460/_0_  ;
	output \g38466/_0_  ;
	output \g38467/_0_  ;
	output \g38468/_0_  ;
	output \g38469/_0_  ;
	output \g38470/_0_  ;
	output \g38471/_0_  ;
	output \g38472/_0_  ;
	output \g38473/_0_  ;
	output \g38474/_0_  ;
	output \g38475/_0_  ;
	output \g38476/_0_  ;
	output \g38477/_0_  ;
	output \g38478/_0_  ;
	output \g38479/_0_  ;
	output \g38528/_0_  ;
	output \g38533/_0_  ;
	output \g38534/_0_  ;
	output \g38536/_0_  ;
	output \g38545/_0_  ;
	output \g38551/_0_  ;
	output \g38554/_0_  ;
	output \g38555/_0_  ;
	output \g38556/_0_  ;
	output \g38575/_0_  ;
	output \g38616/_0_  ;
	output \g38653/_0_  ;
	output \g38656/_0_  ;
	output \g38657/_0_  ;
	output \g38658/_0_  ;
	output \g38660/_0_  ;
	output \g38706/_0_  ;
	output \g38716/_0_  ;
	output \g38717/_0_  ;
	output \g38738/_1_  ;
	output \g38763/_0_  ;
	output \g38790/_0_  ;
	output \g38792/_0_  ;
	output \g38801/_0_  ;
	output \g38803/_0_  ;
	output \g38804/_0_  ;
	output \g38805/_0_  ;
	output \g38806/_0_  ;
	output \g38807/_0_  ;
	output \g38808/_0_  ;
	output \g38809/_0_  ;
	output \g38810/_0_  ;
	output \g38814/_0_  ;
	output \g38833/_0_  ;
	output \g38834/_0_  ;
	output \g38839/_0_  ;
	output \g38840/_0_  ;
	output \g38841/_0_  ;
	output \g38842/_0_  ;
	output \g38846/_0_  ;
	output \g38847/_0_  ;
	output \g38848/_0_  ;
	output \g38849/_0_  ;
	output \g38853/_0_  ;
	output \g38857/_0_  ;
	output \g38872/_0_  ;
	output \g38882/_0_  ;
	output \g38884/_0_  ;
	output \g38885/_0_  ;
	output \g38886/_0_  ;
	output \g38887/_0_  ;
	output \g38931/_0_  ;
	output \g38952/_0_  ;
	output \g38960/_0_  ;
	output \g38971/_0_  ;
	output \g38973/_0_  ;
	output \g38974/_0_  ;
	output \g38975/_0_  ;
	output \g38976/_0_  ;
	output \g38978/_0_  ;
	output \g38981/_0_  ;
	output \g38986/_0_  ;
	output \g38987/_0_  ;
	output \g39001/_3_  ;
	output \g39003/_3_  ;
	output \g39009/_3_  ;
	output \g39011/_3_  ;
	output \g39013/_3_  ;
	output \g39015/_2_  ;
	output \g39017/_2_  ;
	output \g39019/_2_  ;
	output \g39021/_2_  ;
	output \g39060/_0_  ;
	output \g39061/_3_  ;
	output \g39062/_0_  ;
	output \g39063/_0_  ;
	output \g39065/_0_  ;
	output \g39066/_0_  ;
	output \g39093/_0_  ;
	output \g39099/_2_  ;
	output \g39118/_0_  ;
	output \g39123/_0_  ;
	output \g39174/_0_  ;
	output \g39175/_0_  ;
	output \g39176/_0_  ;
	output \g39177/_0_  ;
	output \g39178/_0_  ;
	output \g39185/_0_  ;
	output \g39186/_0_  ;
	output \g39187/_0_  ;
	output \g39188/_0_  ;
	output \g39194/_0_  ;
	output \g39195/_0_  ;
	output \g39196/_0_  ;
	output \g39197/_0_  ;
	output \g39198/_0_  ;
	output \g39199/_0_  ;
	output \g39200/_0_  ;
	output \g39201/_0_  ;
	output \g39202/_0_  ;
	output \g39203/_0_  ;
	output \g39204/_0_  ;
	output \g39216/_3_  ;
	output \g39217/_3_  ;
	output \g39218/_0_  ;
	output \g39219/_0_  ;
	output \g39220/_0_  ;
	output \g39221/_0_  ;
	output \g39299/_0_  ;
	output \g39300/_0_  ;
	output \g39301/_0_  ;
	output \g39302/_0_  ;
	output \g39303/_0_  ;
	output \g39304/_0_  ;
	output \g39305/_0_  ;
	output \g39306/_0_  ;
	output \g39307/_0_  ;
	output \g39308/_0_  ;
	output \g39309/_0_  ;
	output \g39310/_0_  ;
	output \g39311/_0_  ;
	output \g39315/_0_  ;
	output \g39318/_0_  ;
	output \g39321/_0_  ;
	output \g39322/_0_  ;
	output \g39323/_0_  ;
	output \g39333/_0_  ;
	output \g39334/_0_  ;
	output \g39336/_0_  ;
	output \g39338/_0_  ;
	output \g39339/_0_  ;
	output \g39340/_0_  ;
	output \g39341/_0_  ;
	output \g39342/_0_  ;
	output \g39343/_0_  ;
	output \g39344/_0_  ;
	output \g39345/_0_  ;
	output \g39346/_0_  ;
	output \g39349/_0_  ;
	output \g39352/_3_  ;
	output \g39354/_3_  ;
	output \g39371/_3_  ;
	output \g39372/_3_  ;
	output \g39373/_3_  ;
	output \g39374/_3_  ;
	output \g39376/_0_  ;
	output \g39377/_0_  ;
	output \g39471/_0_  ;
	output \g39472/_0_  ;
	output \g39473/_0_  ;
	output \g39474/_0_  ;
	output \g39475/_0_  ;
	output \g39476/_0_  ;
	output \g39477/_0_  ;
	output \g39478/_0_  ;
	output \g39479/_0_  ;
	output \g39480/_0_  ;
	output \g39481/_0_  ;
	output \g39482/_0_  ;
	output \g39483/_0_  ;
	output \g39484/_0_  ;
	output \g39485/_0_  ;
	output \g39486/_0_  ;
	output \g39487/_0_  ;
	output \g39488/_0_  ;
	output \g39492/_0_  ;
	output \g39497/_0_  ;
	output \g39501/_0_  ;
	output \g39502/_0_  ;
	output \g39503/_0_  ;
	output \g39504/_0_  ;
	output \g39505/_0_  ;
	output \g39506/_0_  ;
	output \g39539/_0_  ;
	output \g39541/_0_  ;
	output \g39542/_0_  ;
	output \g39543/_0_  ;
	output \g39544/_0_  ;
	output \g39545/_0_  ;
	output \g39546/_0_  ;
	output \g39547/_0_  ;
	output \g39550/_0_  ;
	output \g39551/_0_  ;
	output \g39563/_0_  ;
	output \g39568/_00_  ;
	output \g39617/_0_  ;
	output \g39618/_0_  ;
	output \g39621/_0_  ;
	output \g39622/_0_  ;
	output \g39623/_0_  ;
	output \g39624/_00_  ;
	output \g39685/_0_  ;
	output \g39690/_0_  ;
	output \g39693/_0_  ;
	output \g39695/_0_  ;
	output \g39697/_0_  ;
	output \g39706/_0_  ;
	output \g39749/_0_  ;
	output \g39750/_0_  ;
	output \g39751/_0_  ;
	output \g39752/_0_  ;
	output \g39753/_0_  ;
	output \g39754/_0_  ;
	output \g39755/_0_  ;
	output \g39756/_0_  ;
	output \g39757/_0_  ;
	output \g39758/_0_  ;
	output \g39759/_0_  ;
	output \g39760/_0_  ;
	output \g39761/_0_  ;
	output \g39762/_0_  ;
	output \g39763/_0_  ;
	output \g39764/_0_  ;
	output \g39765/_0_  ;
	output \g39766/_0_  ;
	output \g39767/_0_  ;
	output \g39768/_0_  ;
	output \g39769/_0_  ;
	output \g39770/_0_  ;
	output \g39772/_0_  ;
	output \g39773/_0_  ;
	output \g39775/_3_  ;
	output \g39776/_3_  ;
	output \g39777/_3_  ;
	output \g39778/_3_  ;
	output \g39779/_3_  ;
	output \g39780/_3_  ;
	output \g39781/_3_  ;
	output \g39782/_3_  ;
	output \g39788/_3_  ;
	output \g39799/_0_  ;
	output \g39800/_0_  ;
	output \g39801/_0_  ;
	output \g39802/_0_  ;
	output \g39927/_0_  ;
	output \g39928/_0_  ;
	output \g39929/_0_  ;
	output \g39930/_0_  ;
	output \g39931/_0_  ;
	output \g39932/_0_  ;
	output \g39933/_0_  ;
	output \g39934/_0_  ;
	output \g39935/_0_  ;
	output \g39936/_0_  ;
	output \g39937/_0_  ;
	output \g39938/_0_  ;
	output \g39939/_0_  ;
	output \g39940/_0_  ;
	output \g39942/_0_  ;
	output \g39943/_0_  ;
	output \g39944/_0_  ;
	output \g39945/_0_  ;
	output \g39956/_0_  ;
	output \g39957/_0_  ;
	output \g39958/_0_  ;
	output \g39959/_0_  ;
	output \g39960/_0_  ;
	output \g39961/_0_  ;
	output \g39962/_0_  ;
	output \g39963/_0_  ;
	output \g39964/_0_  ;
	output \g39969/_0_  ;
	output \g39974/_0_  ;
	output \g39975/_0_  ;
	output \g39993/_0_  ;
	output \g39994/_0_  ;
	output \g40003/_0_  ;
	output \g40004/_0_  ;
	output \g40005/_0_  ;
	output \g40006/_0_  ;
	output \g40016/_0_  ;
	output \g40023/_3_  ;
	output \g40033/_0_  ;
	output \g40034/_0_  ;
	output \g40035/_0_  ;
	output \g40036/_0_  ;
	output \g40037/_0_  ;
	output \g40038/_0_  ;
	output \g40199/_0_  ;
	output \g40200/_0_  ;
	output \g40201/_0_  ;
	output \g40202/_0_  ;
	output \g40203/_0_  ;
	output \g40204/_0_  ;
	output \g40205/_0_  ;
	output \g40206/_0_  ;
	output \g40207/_0_  ;
	output \g40208/_0_  ;
	output \g40209/_0_  ;
	output \g40210/_0_  ;
	output \g40224/_0_  ;
	output \g40225/_0_  ;
	output \g40226/_0_  ;
	output \g40227/_0_  ;
	output \g40234/_0_  ;
	output \g40235/_0_  ;
	output \g40236/_0_  ;
	output \g40237/_0_  ;
	output \g40238/_0_  ;
	output \g40239/_0_  ;
	output \g40240/_0_  ;
	output \g40241/_0_  ;
	output \g40242/_0_  ;
	output \g40243/_0_  ;
	output \g40244/_0_  ;
	output \g40246/_0_  ;
	output \g40247/_0_  ;
	output \g40248/_0_  ;
	output \g40249/_0_  ;
	output \g40250/_0_  ;
	output \g40251/_0_  ;
	output \g40252/_0_  ;
	output \g40253/_0_  ;
	output \g40254/_0_  ;
	output \g40255/_0_  ;
	output \g40257/_0_  ;
	output \g40258/_0_  ;
	output \g40262/_0_  ;
	output \g40264/_0_  ;
	output \g40265/_0_  ;
	output \g40266/_0_  ;
	output \g40267/_0_  ;
	output \g40268/_0_  ;
	output \g40269/_0_  ;
	output \g40270/_0_  ;
	output \g40271/_0_  ;
	output \g40272/_0_  ;
	output \g40273/_0_  ;
	output \g40274/_0_  ;
	output \g40275/_0_  ;
	output \g40276/_0_  ;
	output \g40277/_0_  ;
	output \g40278/_0_  ;
	output \g40280/_2_  ;
	output \g40281/_0_  ;
	output \g40282/_0_  ;
	output \g40283/_0_  ;
	output \g40284/_0_  ;
	output \g40285/_0_  ;
	output \g40286/_0_  ;
	output \g40287/_0_  ;
	output \g40288/_0_  ;
	output \g40289/_0_  ;
	output \g40290/_0_  ;
	output \g40291/_0_  ;
	output \g40297/_0_  ;
	output \g40298/_0_  ;
	output \g40299/_0_  ;
	output \g40300/_0_  ;
	output \g40301/_0_  ;
	output \g40302/_0_  ;
	output \g40303/_0_  ;
	output \g40304/_0_  ;
	output \g40306/_0_  ;
	output \g40307/_0_  ;
	output \g40308/_0_  ;
	output \g40309/_0_  ;
	output \g40310/_0_  ;
	output \g40311/_0_  ;
	output \g40312/_0_  ;
	output \g40313/_0_  ;
	output \g40314/_0_  ;
	output \g40315/_0_  ;
	output \g40316/_0_  ;
	output \g40317/_0_  ;
	output \g40318/_0_  ;
	output \g40319/_0_  ;
	output \g40320/_0_  ;
	output \g40324/_0_  ;
	output \g40325/_0_  ;
	output \g40326/_0_  ;
	output \g40327/_0_  ;
	output \g40328/_0_  ;
	output \g40329/_0_  ;
	output \g40330/_0_  ;
	output \g40331/_0_  ;
	output \g40332/_0_  ;
	output \g40333/_0_  ;
	output \g40334/_0_  ;
	output \g40335/_0_  ;
	output \g40336/_0_  ;
	output \g40337/_0_  ;
	output \g40338/_0_  ;
	output \g40339/_0_  ;
	output \g40340/_0_  ;
	output \g40341/_0_  ;
	output \g40342/_0_  ;
	output \g40343/_0_  ;
	output \g40344/_0_  ;
	output \g40345/_0_  ;
	output \g40346/_0_  ;
	output \g40347/_0_  ;
	output \g40350/_0_  ;
	output \g40353/_0_  ;
	output \g40354/_0_  ;
	output \g40355/_0_  ;
	output \g40374/_0_  ;
	output \g40457/_0_  ;
	output \g40458/_0_  ;
	output \g40549/_0_  ;
	output \g40550/_0_  ;
	output \g40551/_0_  ;
	output \g40552/_0_  ;
	output \g40553/_0_  ;
	output \g40554/_0_  ;
	output \g40556/_0_  ;
	output \g40557/_0_  ;
	output \g40558/_0_  ;
	output \g40559/_0_  ;
	output \g40561/_0_  ;
	output \g40562/_0_  ;
	output \g40563/_0_  ;
	output \g40565/_0_  ;
	output \g40566/_0_  ;
	output \g40567/_0_  ;
	output \g40569/_0_  ;
	output \g40570/_0_  ;
	output \g40571/_0_  ;
	output \g40572/_0_  ;
	output \g40573/_0_  ;
	output \g40574/_0_  ;
	output \g40575/_0_  ;
	output \g40576/_0_  ;
	output \g40577/_0_  ;
	output \g40578/_0_  ;
	output \g40579/_0_  ;
	output \g40580/_0_  ;
	output \g40581/_0_  ;
	output \g40582/_0_  ;
	output \g40583/_0_  ;
	output \g40584/_0_  ;
	output \g40586/_0_  ;
	output \g40587/_0_  ;
	output \g40588/_0_  ;
	output \g40589/_0_  ;
	output \g40591/_0_  ;
	output \g40592/_0_  ;
	output \g40593/_0_  ;
	output \g40594/_0_  ;
	output \g40595/_0_  ;
	output \g40596/_0_  ;
	output \g40597/_0_  ;
	output \g40598/_0_  ;
	output \g40599/_0_  ;
	output \g40600/_0_  ;
	output \g40601/_0_  ;
	output \g40602/_0_  ;
	output \g40603/_0_  ;
	output \g40604/_0_  ;
	output \g40605/_0_  ;
	output \g40606/_0_  ;
	output \g40607/_0_  ;
	output \g40608/_0_  ;
	output \g40609/_0_  ;
	output \g40610/_0_  ;
	output \g40611/_0_  ;
	output \g40612/_0_  ;
	output \g40613/_0_  ;
	output \g40614/_0_  ;
	output \g40617/_0_  ;
	output \g40629/_0_  ;
	output \g40632/_0_  ;
	output \g40633/_0_  ;
	output \g40634/_0_  ;
	output \g40635/_0_  ;
	output \g40636/_0_  ;
	output \g40637/_0_  ;
	output \g40638/_0_  ;
	output \g40639/_0_  ;
	output \g40640/_0_  ;
	output \g40641/_0_  ;
	output \g40642/_0_  ;
	output \g40643/_0_  ;
	output \g40644/_0_  ;
	output \g40645/_0_  ;
	output \g40646/_0_  ;
	output \g40647/_0_  ;
	output \g40648/_0_  ;
	output \g40649/_0_  ;
	output \g40650/_0_  ;
	output \g40651/_0_  ;
	output \g40652/_0_  ;
	output \g40653/_0_  ;
	output \g40654/_0_  ;
	output \g40655/_0_  ;
	output \g40661/_0_  ;
	output \g40663/_0_  ;
	output \g40664/_0_  ;
	output \g40665/_0_  ;
	output \g40666/_0_  ;
	output \g40667/_0_  ;
	output \g40668/_0_  ;
	output \g40669/_0_  ;
	output \g40670/_0_  ;
	output \g40671/_0_  ;
	output \g40672/_0_  ;
	output \g40673/_0_  ;
	output \g40674/_0_  ;
	output \g40675/_0_  ;
	output \g40676/_0_  ;
	output \g40677/_0_  ;
	output \g40678/_0_  ;
	output \g40679/_0_  ;
	output \g40680/_0_  ;
	output \g40681/_0_  ;
	output \g40682/_0_  ;
	output \g40683/_0_  ;
	output \g40684/_0_  ;
	output \g40685/_0_  ;
	output \g40689/_0_  ;
	output \g40690/_0_  ;
	output \g40691/_0_  ;
	output \g40692/_0_  ;
	output \g40693/_0_  ;
	output \g40694/_0_  ;
	output \g40695/_0_  ;
	output \g40696/_0_  ;
	output \g40697/_0_  ;
	output \g40698/_0_  ;
	output \g40699/_0_  ;
	output \g40700/_0_  ;
	output \g40701/_0_  ;
	output \g40702/_0_  ;
	output \g40703/_0_  ;
	output \g40704/_0_  ;
	output \g40705/_0_  ;
	output \g40706/_0_  ;
	output \g40707/_0_  ;
	output \g40708/_0_  ;
	output \g40709/_0_  ;
	output \g40710/_0_  ;
	output \g40711/_0_  ;
	output \g40712/_0_  ;
	output \g40758/_00_  ;
	output \g40759/_0_  ;
	output \g40812/_0_  ;
	output \g40816/_0_  ;
	output \g40817/_0_  ;
	output \g40818/_0_  ;
	output \g40819/_0_  ;
	output \g40820/_0_  ;
	output \g40822/_3_  ;
	output \g40823/_3_  ;
	output \g40824/_3_  ;
	output \g40825/_3_  ;
	output \g40849/_3_  ;
	output \g40915/_0_  ;
	output \g40916/_0_  ;
	output \g40917/_0_  ;
	output \g40920/_0_  ;
	output \g40923/_0_  ;
	output \g40926/_0_  ;
	output \g40927/_0_  ;
	output \g40930/_0_  ;
	output \g40931/_0_  ;
	output \g41138/_0_  ;
	output \g41152/_0_  ;
	output \g41180/_0_  ;
	output \g41185/_0_  ;
	output \g41186/_0_  ;
	output \g41187/_0_  ;
	output \g41189/_0_  ;
	output \g41190/_0_  ;
	output \g41191/_0_  ;
	output \g41192/_0_  ;
	output \g41193/_0_  ;
	output \g41195/_0_  ;
	output \g41199/_0_  ;
	output \g41207/_0_  ;
	output \g41221/_0_  ;
	output \g41226/_0_  ;
	output \g41227/_0_  ;
	output \g41230/_0_  ;
	output \g41231/_0_  ;
	output \g41234/_0_  ;
	output \g41238/_0_  ;
	output \g41239/_0_  ;
	output \g41275/_0_  ;
	output \g41277/_0_  ;
	output \g41278/_0_  ;
	output \g41279/_0_  ;
	output \g41280/_0_  ;
	output \g41281/_0_  ;
	output \g41282/_0_  ;
	output \g41283/_0_  ;
	output \g41284/_0_  ;
	output \g41285/_0_  ;
	output \g41286/_0_  ;
	output \g41287/_0_  ;
	output \g41288/_0_  ;
	output \g41289/_0_  ;
	output \g41291/_3_  ;
	output \g41330/_0_  ;
	output \g41332/_0_  ;
	output \g41334/_0_  ;
	output \g41340/_0_  ;
	output \g41343/_0_  ;
	output \g41345/_0_  ;
	output \g41348/_0_  ;
	output \g41349/_0_  ;
	output \g41350/_0_  ;
	output \g41351/_0_  ;
	output \g41356/_0_  ;
	output \g41394/_0_  ;
	output \g41423/_0_  ;
	output \g41426/_3_  ;
	output \g41427/_3_  ;
	output \g41428/_3_  ;
	output \g41429/_3_  ;
	output \g41430/_3_  ;
	output \g41431/_3_  ;
	output \g41432/_3_  ;
	output \g41433/_3_  ;
	output \g41434/_3_  ;
	output \g41435/_3_  ;
	output \g41436/_3_  ;
	output \g41437/_3_  ;
	output \g41438/_3_  ;
	output \g41439/_3_  ;
	output \g41440/_3_  ;
	output \g41441/_3_  ;
	output \g41442/_0_  ;
	output \g41445/_3_  ;
	output \g41446/_0_  ;
	output \g41449/_0_  ;
	output \g41464/_0_  ;
	output \g41466/_0_  ;
	output \g41468/_0_  ;
	output \g41469/_0_  ;
	output \g41471/_0_  ;
	output \g41795/_0_  ;
	output \g41799/_0_  ;
	output \g41800/_0_  ;
	output \g41801/_0_  ;
	output \g41802/_0_  ;
	output \g41803/_0_  ;
	output \g41804/_0_  ;
	output \g41805/_0_  ;
	output \g41806/_0_  ;
	output \g41807/_0_  ;
	output \g41808/_0_  ;
	output \g41809/_0_  ;
	output \g41810/_0_  ;
	output \g41811/_0_  ;
	output \g41812/_0_  ;
	output \g41814/_0_  ;
	output \g41815/_0_  ;
	output \g41816/_0_  ;
	output \g41817/_0_  ;
	output \g41818/_0_  ;
	output \g41819/_0_  ;
	output \g41820/_0_  ;
	output \g41821/_0_  ;
	output \g41822/_0_  ;
	output \g41823/_0_  ;
	output \g41825/_0_  ;
	output \g41826/_0_  ;
	output \g41827/_0_  ;
	output \g41828/_0_  ;
	output \g41829/_0_  ;
	output \g41830/_0_  ;
	output \g41831/_0_  ;
	output \g41832/_0_  ;
	output \g41833/_0_  ;
	output \g41834/_0_  ;
	output \g41835/_0_  ;
	output \g41836/_0_  ;
	output \g41837/_0_  ;
	output \g41838/_0_  ;
	output \g41839/_0_  ;
	output \g41840/_0_  ;
	output \g41841/_0_  ;
	output \g41842/_0_  ;
	output \g41843/_0_  ;
	output \g41844/_0_  ;
	output \g41845/_0_  ;
	output \g41846/_0_  ;
	output \g41847/_0_  ;
	output \g41848/_0_  ;
	output \g41849/_0_  ;
	output \g41850/_0_  ;
	output \g41851/_0_  ;
	output \g41852/_0_  ;
	output \g41853/_0_  ;
	output \g41854/_0_  ;
	output \g41855/_0_  ;
	output \g41856/_0_  ;
	output \g41857/_0_  ;
	output \g41858/_0_  ;
	output \g41859/_0_  ;
	output \g41860/_0_  ;
	output \g41861/_0_  ;
	output \g41862/_0_  ;
	output \g41863/_0_  ;
	output \g41864/_0_  ;
	output \g41865/_0_  ;
	output \g41866/_0_  ;
	output \g41867/_0_  ;
	output \g41868/_0_  ;
	output \g41869/_0_  ;
	output \g41870/_0_  ;
	output \g41871/_0_  ;
	output \g41872/_0_  ;
	output \g41873/_0_  ;
	output \g41874/_0_  ;
	output \g41875/_0_  ;
	output \g41876/_0_  ;
	output \g41877/_0_  ;
	output \g41878/_0_  ;
	output \g41879/_0_  ;
	output \g41880/_0_  ;
	output \g41881/_0_  ;
	output \g41882/_0_  ;
	output \g41883/_0_  ;
	output \g41884/_0_  ;
	output \g41885/_0_  ;
	output \g41886/_0_  ;
	output \g41887/_0_  ;
	output \g41888/_0_  ;
	output \g41889/_0_  ;
	output \g41890/_0_  ;
	output \g41891/_0_  ;
	output \g41902/_0_  ;
	output \g41904/_0_  ;
	output \g41906/_0_  ;
	output \g41907/_0_  ;
	output \g41954/_0_  ;
	output \g41955/_0_  ;
	output \g41956/_0_  ;
	output \g41957/_0_  ;
	output \g41958/_0_  ;
	output \g41959/_0_  ;
	output \g41960/_0_  ;
	output \g41962/_0_  ;
	output \g41963/_0_  ;
	output \g41964/_0_  ;
	output \g41965/_0_  ;
	output \g41966/_0_  ;
	output \g41967/_0_  ;
	output \g41968/_0_  ;
	output \g41969/_0_  ;
	output \g41970/_0_  ;
	output \g41971/_0_  ;
	output \g41972/_0_  ;
	output \g41973/_0_  ;
	output \g41974/_0_  ;
	output \g41975/_0_  ;
	output \g41976/_0_  ;
	output \g41977/_0_  ;
	output \g41978/_0_  ;
	output \g41979/_0_  ;
	output \g42062/_0_  ;
	output \g42079/_0_  ;
	output \g42142/_0_  ;
	output \g42143/_0_  ;
	output \g42144/_0_  ;
	output \g42154/_0_  ;
	output \g42157/_0_  ;
	output \g42160/_0_  ;
	output \g42181/_0_  ;
	output \g42203/_0_  ;
	output \g42204/_3_  ;
	output \g42205/_3_  ;
	output \g42206/_3_  ;
	output \g42208/_0_  ;
	output \g42220/_0_  ;
	output \g42225/_0_  ;
	output \g42251/_0_  ;
	output \g42273/_0_  ;
	output \g42335/_0_  ;
	output \g42357/_0_  ;
	output \g42380/_0_  ;
	output \g42381/_0_  ;
	output \g42383/_0_  ;
	output \g42386/_0_  ;
	output \g42388/_0_  ;
	output \g42475/_0_  ;
	output \g42476/_0_  ;
	output \g42477/_0_  ;
	output \g42478/_0_  ;
	output \g42479/_0_  ;
	output \g42480/_0_  ;
	output \g42481/_0_  ;
	output \g42482/_0_  ;
	output \g42483/_0_  ;
	output \g42484/_0_  ;
	output \g42485/_0_  ;
	output \g42486/_0_  ;
	output \g42487/_0_  ;
	output \g42488/_0_  ;
	output \g42490/_0_  ;
	output \g42491/_0_  ;
	output \g42493/_0_  ;
	output \g42494/_0_  ;
	output \g42495/_0_  ;
	output \g42496/_0_  ;
	output \g42497/_0_  ;
	output \g42498/_0_  ;
	output \g42499/_0_  ;
	output \g42500/_0_  ;
	output \g42501/_0_  ;
	output \g42502/_0_  ;
	output \g42503/_0_  ;
	output \g42504/_0_  ;
	output \g42505/_0_  ;
	output \g42506/_0_  ;
	output \g42507/_0_  ;
	output \g42508/_0_  ;
	output \g42509/_0_  ;
	output \g42510/_0_  ;
	output \g42511/_0_  ;
	output \g42512/_0_  ;
	output \g42513/_0_  ;
	output \g42514/_0_  ;
	output \g42515/_0_  ;
	output \g42516/_0_  ;
	output \g42517/_0_  ;
	output \g42518/_0_  ;
	output \g42519/_0_  ;
	output \g42521/_0_  ;
	output \g42522/_0_  ;
	output \g42523/_0_  ;
	output \g42524/_0_  ;
	output \g42525/_0_  ;
	output \g42526/_0_  ;
	output \g42527/_0_  ;
	output \g42528/_0_  ;
	output \g42529/_0_  ;
	output \g42530/_0_  ;
	output \g42531/_0_  ;
	output \g42532/_0_  ;
	output \g42533/_0_  ;
	output \g42534/_0_  ;
	output \g42535/_0_  ;
	output \g42536/_0_  ;
	output \g42537/_0_  ;
	output \g42538/_0_  ;
	output \g42539/_0_  ;
	output \g42540/_0_  ;
	output \g42541/_0_  ;
	output \g42542/_0_  ;
	output \g42543/_0_  ;
	output \g42544/_0_  ;
	output \g42545/_0_  ;
	output \g42548/_0_  ;
	output \g42557/_0_  ;
	output \g42564/_0_  ;
	output \g42565/_0_  ;
	output \g42566/_0_  ;
	output \g42567/_0_  ;
	output \g42568/_0_  ;
	output \g42569/_0_  ;
	output \g42570/_0_  ;
	output \g42571/_0_  ;
	output \g42572/_0_  ;
	output \g42573/_0_  ;
	output \g42574/_0_  ;
	output \g42575/_0_  ;
	output \g42576/_0_  ;
	output \g42577/_0_  ;
	output \g42578/_0_  ;
	output \g42581/_0_  ;
	output \g42589/_0_  ;
	output \g42590/_0_  ;
	output \g42591/_0_  ;
	output \g42592/_0_  ;
	output \g42593/_0_  ;
	output \g42594/_0_  ;
	output \g42595/_0_  ;
	output \g42596/_0_  ;
	output \g42597/_0_  ;
	output \g42598/_0_  ;
	output \g42599/_0_  ;
	output \g42600/_0_  ;
	output \g42601/_0_  ;
	output \g42602/_0_  ;
	output \g42603/_0_  ;
	output \g42604/_0_  ;
	output \g42605/_0_  ;
	output \g42606/_0_  ;
	output \g42607/_0_  ;
	output \g42608/_0_  ;
	output \g42609/_0_  ;
	output \g42610/_0_  ;
	output \g42611/_0_  ;
	output \g42612/_0_  ;
	output \g42613/_0_  ;
	output \g42614/_0_  ;
	output \g42615/_0_  ;
	output \g42616/_0_  ;
	output \g42617/_0_  ;
	output \g42618/_0_  ;
	output \g42619/_0_  ;
	output \g42620/_0_  ;
	output \g42622/_0_  ;
	output \g42623/_0_  ;
	output \g42627/_0_  ;
	output \g42628/_0_  ;
	output \g42629/_0_  ;
	output \g42630/_0_  ;
	output \g42631/_0_  ;
	output \g42632/_0_  ;
	output \g42633/_0_  ;
	output \g42634/_0_  ;
	output \g42635/_0_  ;
	output \g42636/_0_  ;
	output \g42637/_0_  ;
	output \g42638/_0_  ;
	output \g42639/_0_  ;
	output \g42640/_0_  ;
	output \g42641/_0_  ;
	output \g42642/_0_  ;
	output \g42643/_0_  ;
	output \g42644/_0_  ;
	output \g42645/_0_  ;
	output \g42646/_0_  ;
	output \g42647/_0_  ;
	output \g42648/_0_  ;
	output \g42649/_0_  ;
	output \g42650/_0_  ;
	output \g42666/_0_  ;
	output \g42667/_0_  ;
	output \g42668/_0_  ;
	output \g42669/_0_  ;
	output \g42670/_0_  ;
	output \g42671/_0_  ;
	output \g42672/_0_  ;
	output \g42673/_0_  ;
	output \g42674/_0_  ;
	output \g42675/_0_  ;
	output \g42676/_0_  ;
	output \g42677/_0_  ;
	output \g42678/_0_  ;
	output \g42680/_0_  ;
	output \g42681/_0_  ;
	output \g42685/_0_  ;
	output \g42686/_0_  ;
	output \g42688/_0_  ;
	output \g42689/_0_  ;
	output \g42690/_0_  ;
	output \g42691/_0_  ;
	output \g42692/_0_  ;
	output \g42693/_0_  ;
	output \g42694/_0_  ;
	output \g42695/_0_  ;
	output \g42696/_0_  ;
	output \g42697/_0_  ;
	output \g42698/_0_  ;
	output \g42699/_0_  ;
	output \g42700/_0_  ;
	output \g42701/_0_  ;
	output \g42702/_0_  ;
	output \g42703/_0_  ;
	output \g42704/_0_  ;
	output \g42705/_0_  ;
	output \g42706/_0_  ;
	output \g42707/_0_  ;
	output \g42708/_0_  ;
	output \g42709/_0_  ;
	output \g42710/_0_  ;
	output \g42711/_0_  ;
	output \g42712/_0_  ;
	output \g42713/_0_  ;
	output \g42715/_0_  ;
	output \g42716/_0_  ;
	output \g42717/_0_  ;
	output \g42718/_0_  ;
	output \g42723/_1_  ;
	output \g42727/_0_  ;
	output \g42728/_0_  ;
	output \g42729/_0_  ;
	output \g42730/_0_  ;
	output \g42731/_0_  ;
	output \g42732/_0_  ;
	output \g42733/_0_  ;
	output \g42734/_0_  ;
	output \g42735/_0_  ;
	output \g42736/_0_  ;
	output \g42737/_0_  ;
	output \g42738/_0_  ;
	output \g42739/_0_  ;
	output \g42740/_0_  ;
	output \g42741/_0_  ;
	output \g42742/_0_  ;
	output \g42743/_0_  ;
	output \g42744/_0_  ;
	output \g42745/_0_  ;
	output \g42746/_0_  ;
	output \g42747/_0_  ;
	output \g42748/_0_  ;
	output \g42749/_0_  ;
	output \g42750/_0_  ;
	output \g42751/_0_  ;
	output \g42754/_0_  ;
	output \g42767/_0_  ;
	output \g42768/_0_  ;
	output \g42772/_0_  ;
	output \g42773/_0_  ;
	output \g42774/_0_  ;
	output \g42775/_0_  ;
	output \g42776/_0_  ;
	output \g42777/_0_  ;
	output \g42778/_0_  ;
	output \g42779/_0_  ;
	output \g42780/_0_  ;
	output \g42781/_0_  ;
	output \g42782/_0_  ;
	output \g42783/_0_  ;
	output \g42784/_0_  ;
	output \g42785/_0_  ;
	output \g42790/_0_  ;
	output \g42791/_0_  ;
	output \g42792/_0_  ;
	output \g42793/_0_  ;
	output \g42794/_0_  ;
	output \g42795/_0_  ;
	output \g42796/_0_  ;
	output \g42797/_0_  ;
	output \g42798/_0_  ;
	output \g42799/_0_  ;
	output \g42800/_0_  ;
	output \g42801/_0_  ;
	output \g42802/_0_  ;
	output \g42803/_0_  ;
	output \g42804/_0_  ;
	output \g42805/_0_  ;
	output \g42806/_0_  ;
	output \g42807/_0_  ;
	output \g42808/_0_  ;
	output \g42809/_0_  ;
	output \g42810/_0_  ;
	output \g42811/_0_  ;
	output \g42812/_0_  ;
	output \g42813/_0_  ;
	output \g42814/_0_  ;
	output \g42815/_0_  ;
	output \g42816/_0_  ;
	output \g42817/_0_  ;
	output \g42818/_0_  ;
	output \g42819/_0_  ;
	output \g42820/_0_  ;
	output \g42821/_0_  ;
	output \g42824/_0_  ;
	output \g42825/_0_  ;
	output \g42826/_0_  ;
	output \g42827/_0_  ;
	output \g42828/_0_  ;
	output \g42829/_0_  ;
	output \g42830/_0_  ;
	output \g42831/_0_  ;
	output \g42832/_0_  ;
	output \g42833/_0_  ;
	output \g42834/_0_  ;
	output \g42835/_0_  ;
	output \g42836/_0_  ;
	output \g42837/_0_  ;
	output \g42838/_0_  ;
	output \g42839/_0_  ;
	output \g42840/_0_  ;
	output \g42841/_0_  ;
	output \g42842/_0_  ;
	output \g42843/_0_  ;
	output \g42844/_0_  ;
	output \g42845/_0_  ;
	output \g42846/_0_  ;
	output \g42907/_0_  ;
	output \g42914/_0_  ;
	output \g42924/_0_  ;
	output \g42925/_0_  ;
	output \g42926/_0_  ;
	output \g42927/_0_  ;
	output \g42928/_0_  ;
	output \g42929/_0_  ;
	output \g42930/_0_  ;
	output \g42931/_0_  ;
	output \g42933/_0_  ;
	output \g42941/_0_  ;
	output \g42947/_0_  ;
	output \g42950/_0_  ;
	output \g42955/_0_  ;
	output \g42956/_0_  ;
	output \g42972/_3_  ;
	output \g42973/_3_  ;
	output \g42974/_3_  ;
	output \g43178/_0_  ;
	output \g43179/_0_  ;
	output \g43184/_0_  ;
	output \g43186/_0_  ;
	output \g43187/_0_  ;
	output \g43190/_0_  ;
	output \g43191/_0_  ;
	output \g43192/_0_  ;
	output \g43202/_0_  ;
	output \g43205/_0_  ;
	output \g43206/_0_  ;
	output \g43207/_0_  ;
	output \g43209/_2_  ;
	output \g43228/_0_  ;
	output \g43233/_0_  ;
	output \g43235/_0_  ;
	output \g43236/_0_  ;
	output \g43237/_0_  ;
	output \g43238/_0_  ;
	output \g43280/_0_  ;
	output \g43287/_0_  ;
	output \g43289/_0_  ;
	output \g43290/_0_  ;
	output \g43291/_0_  ;
	output \g43292/_0_  ;
	output \g43303/_0_  ;
	output \g43311/_0_  ;
	output \g43312/_0_  ;
	output \g43363/_0_  ;
	output \g43364/_0_  ;
	output \g43366/_0_  ;
	output \g43367/_0_  ;
	output \g43370/_0_  ;
	output \g43371/_0_  ;
	output \g43374/_0_  ;
	output \g43413/_0_  ;
	output \g43414/_0_  ;
	output \g43415/_0_  ;
	output \g43416/_0_  ;
	output \g43422/_0_  ;
	output \g43427/_0_  ;
	output \g43428/_0_  ;
	output \g43528/_1__syn_2  ;
	output \g43630/_0_  ;
	output \g43633/_3_  ;
	output \g43647/_0_  ;
	output \g43648/_0_  ;
	output \g43656/_0_  ;
	output \g43657/_0_  ;
	output \g43667/_0_  ;
	output \g43668/_0_  ;
	output \g43675/_0_  ;
	output \g43678/_0_  ;
	output \g43787/_0_  ;
	output \g44055/_0_  ;
	output \g44092/_0_  ;
	output \g44093/_0_  ;
	output \g44176/_0_  ;
	output \g44181/_0_  ;
	output \g44433/_0_  ;
	output \g44510/_0_  ;
	output \g44515/_2_  ;
	output \g44522/_0_  ;
	output \g44529/_2_  ;
	output \g44537/_2_  ;
	output \g44544/_2_  ;
	output \g44594/_0_  ;
	output \g44695/_0_  ;
	output \g44697/_0_  ;
	output \g44699/_0_  ;
	output \g44700/_0_  ;
	output \g44843/_0_  ;
	output \g44844/_0_  ;
	output \g44879/_0_  ;
	output \g44880/_0_  ;
	output \g44881/_0_  ;
	output \g44882/_0_  ;
	output \g44906/_2_  ;
	output \g44910/_0_  ;
	output \g44912/_0_  ;
	output \g44954/_0_  ;
	output \g45000/_0_  ;
	output \g45001/_0_  ;
	output \g45002/_0_  ;
	output \g45003/_0_  ;
	output \g45021/_1_  ;
	output \g45025/_0_  ;
	output \g45051/_0_  ;
	output \g45104/_0_  ;
	output \g45111/_0_  ;
	output \g45112/_0_  ;
	output \g45116/_0_  ;
	output \g45155/_0_  ;
	output \g45238/_0_  ;
	output \g45239/_0_  ;
	output \g45240/_0_  ;
	output \g45241/_0_  ;
	output \g45249/_0_  ;
	output \g45257/_0_  ;
	output \g45332/_0_  ;
	output \g45334/_0_  ;
	output \g45336/_0_  ;
	output \g45337/_0_  ;
	output \g45342/_0_  ;
	output \g45459/_0_  ;
	output \g45460/_0_  ;
	output \g45466/_0_  ;
	output \g45469/_0_  ;
	output \g45470/_0_  ;
	output \g45474/_0_  ;
	output \g45475/_0_  ;
	output \g45477/_0_  ;
	output \g45481/_0_  ;
	output \g45482/_0_  ;
	output \g45487/_0_  ;
	output \g45488/_0_  ;
	output \g45518/_3_  ;
	output \g45519/_3_  ;
	output \g45520/_3_  ;
	output \g45521/_3_  ;
	output \g45522/_3_  ;
	output \g45523/_3_  ;
	output \g45524/_3_  ;
	output \g45525/_3_  ;
	output \g45526/_3_  ;
	output \g45530/_3_  ;
	output \g45531/_3_  ;
	output \g45532/_3_  ;
	output \g45533/_3_  ;
	output \g45534/_3_  ;
	output \g45535/_3_  ;
	output \g45536/_3_  ;
	output \g45559/_3_  ;
	output \g45596/_0_  ;
	output \g45605/_0_  ;
	output \g45622/_0_  ;
	output \g45623/_0_  ;
	output \g45630/_0_  ;
	output \g45747/_0_  ;
	output \g45753/_0_  ;
	output \g45796/_0_  ;
	output \g45837/_0_  ;
	output \g45882/_0_  ;
	output \g45903/_0_  ;
	output \g45912/_0_  ;
	output \g45946/_0_  ;
	output \g45999/_0_  ;
	output \g46000/_0_  ;
	output \g46001/_0_  ;
	output \g46002/_0_  ;
	output \g46012/_0_  ;
	output \g46014/_0_  ;
	output \g46017/_0_  ;
	output \g46018/_0_  ;
	output \g46021/_0_  ;
	output \g46024/_0_  ;
	output \g46026/_0_  ;
	output \g46029/_0_  ;
	output \g46053/_0_  ;
	output \g46083/_0_  ;
	output \g46093/_0_  ;
	output \g46142/_0_  ;
	output \g46154/_1__syn_2  ;
	output \g46265/_0_  ;
	output \g46266/_0_  ;
	output \g46268/_0_  ;
	output \g46270/_0_  ;
	output \g46273/_0_  ;
	output \g46274/_0_  ;
	output \g46275/_0_  ;
	output \g46276/_0_  ;
	output \g46278/_0_  ;
	output \g46385/_0_  ;
	output \g46411/_0_  ;
	output \g46414/_0_  ;
	output \g46479/_0_  ;
	output \g46520/_0_  ;
	output \g46521/_0_  ;
	output \g46530/_0_  ;
	output \g46531/_0_  ;
	output \g46597/_0_  ;
	output \g46610/_0_  ;
	output \g46617/_0_  ;
	output \g46632/_0_  ;
	output \g46637/_0_  ;
	output \g46722/_0_  ;
	output \g46723/_0_  ;
	output \g46724/_0_  ;
	output \g46725/_0_  ;
	output \g46813/_0_  ;
	output \g46842/_0_  ;
	output \g46888/_0_  ;
	output \g46891/_0_  ;
	output \g46894/_0_  ;
	output \g46905/_0_  ;
	output \g46940/_0_  ;
	output \g46992/_0_  ;
	output \g46995/_0_  ;
	output \g47037/_3_  ;
	output \g47053/_0_  ;
	output \g47140/_0_  ;
	output \g47155/_3_  ;
	output \g47209/_0_  ;
	output \g47211/_0_  ;
	output \g47213/_0_  ;
	output \g47215/_0_  ;
	output \g47337/_0_  ;
	output \g47433/_0_  ;
	output \g47972/_0_  ;
	output \g47976/_0_  ;
	output \g48081/_0_  ;
	output \g48171/_0_  ;
	output \g48227/_0_  ;
	output \g48234/_1_  ;
	output \g48257/_1_  ;
	output \g48266/_0_  ;
	output \g48281/_0_  ;
	output \g48291/_1_  ;
	output \g48322/_0_  ;
	output \g48345/_0_  ;
	output \g48429/_0_  ;
	output \g48495/_1_  ;
	output \g48549/_0_  ;
	output \g48589/_0_  ;
	output \g48642/_0_  ;
	output \g48722/_0_  ;
	output \g48748/_0_  ;
	output \g48749/_0_  ;
	output \g48763/_0_  ;
	output \g48867/_0_  ;
	output \g48876/_0_  ;
	output \g48880/_0_  ;
	output \g49023/_0_  ;
	output \g49205/_0_  ;
	output \g49314/_0_  ;
	output \g49432/_0__syn_2  ;
	output \g49512/_0_  ;
	output \g49707/_0_  ;
	output \g49737/_0_  ;
	output \g49831/_0_  ;
	output \g49922/_1_  ;
	output \g50132/_0_  ;
	output \g51376/_0_  ;
	output \g51412/_0_  ;
	output \g51822/_0_  ;
	output \g52114/_0_  ;
	output \g52156/_0_  ;
	output \g54427/_0_  ;
	output \g54557/_0_  ;
	output \g54561/_3_  ;
	output \g55079/_0_  ;
	output \sram_adr_o[0]_pad  ;
	output \sram_adr_o[10]_pad  ;
	output \sram_adr_o[11]_pad  ;
	output \sram_adr_o[12]_pad  ;
	output \sram_adr_o[13]_pad  ;
	output \sram_adr_o[14]_pad  ;
	output \sram_adr_o[1]_pad  ;
	output \sram_adr_o[2]_pad  ;
	output \sram_adr_o[3]_pad  ;
	output \sram_adr_o[4]_pad  ;
	output \sram_adr_o[5]_pad  ;
	output \sram_adr_o[6]_pad  ;
	output \sram_adr_o[7]_pad  ;
	output \sram_adr_o[8]_pad  ;
	output \sram_adr_o[9]_pad  ;
	output \sram_data_o[0]_pad  ;
	output \sram_data_o[10]_pad  ;
	output \sram_data_o[11]_pad  ;
	output \sram_data_o[12]_pad  ;
	output \sram_data_o[13]_pad  ;
	output \sram_data_o[14]_pad  ;
	output \sram_data_o[15]_pad  ;
	output \sram_data_o[16]_pad  ;
	output \sram_data_o[17]_pad  ;
	output \sram_data_o[18]_pad  ;
	output \sram_data_o[19]_pad  ;
	output \sram_data_o[1]_pad  ;
	output \sram_data_o[20]_pad  ;
	output \sram_data_o[21]_pad  ;
	output \sram_data_o[22]_pad  ;
	output \sram_data_o[23]_pad  ;
	output \sram_data_o[24]_pad  ;
	output \sram_data_o[25]_pad  ;
	output \sram_data_o[26]_pad  ;
	output \sram_data_o[27]_pad  ;
	output \sram_data_o[28]_pad  ;
	output \sram_data_o[29]_pad  ;
	output \sram_data_o[2]_pad  ;
	output \sram_data_o[30]_pad  ;
	output \sram_data_o[31]_pad  ;
	output \sram_data_o[3]_pad  ;
	output \sram_data_o[4]_pad  ;
	output \sram_data_o[5]_pad  ;
	output \sram_data_o[6]_pad  ;
	output \sram_data_o[7]_pad  ;
	output \sram_data_o[8]_pad  ;
	output \sram_data_o[9]_pad  ;
	output sram_re_o_pad ;
	output sram_we_o_pad ;
	output \u4_utmi_vend_ctrl_r_reg[0]/P0001_reg_syn_3  ;
	output \u4_utmi_vend_ctrl_r_reg[1]/P0001_reg_syn_3  ;
	output \u4_utmi_vend_ctrl_r_reg[2]/P0001_reg_syn_3  ;
	output \u4_utmi_vend_ctrl_r_reg[3]/P0001_reg_syn_3  ;
	wire _w10902_ ;
	wire _w10901_ ;
	wire _w10900_ ;
	wire _w10899_ ;
	wire _w10898_ ;
	wire _w10897_ ;
	wire _w10896_ ;
	wire _w10895_ ;
	wire _w10894_ ;
	wire _w10893_ ;
	wire _w10892_ ;
	wire _w10891_ ;
	wire _w10890_ ;
	wire _w10889_ ;
	wire _w10888_ ;
	wire _w10887_ ;
	wire _w10886_ ;
	wire _w10885_ ;
	wire _w10884_ ;
	wire _w10883_ ;
	wire _w10882_ ;
	wire _w10881_ ;
	wire _w10880_ ;
	wire _w10879_ ;
	wire _w10878_ ;
	wire _w10877_ ;
	wire _w10876_ ;
	wire _w10875_ ;
	wire _w10874_ ;
	wire _w10873_ ;
	wire _w10872_ ;
	wire _w10871_ ;
	wire _w10870_ ;
	wire _w10869_ ;
	wire _w10868_ ;
	wire _w10867_ ;
	wire _w10866_ ;
	wire _w10865_ ;
	wire _w10864_ ;
	wire _w10863_ ;
	wire _w10862_ ;
	wire _w10861_ ;
	wire _w10860_ ;
	wire _w10859_ ;
	wire _w10858_ ;
	wire _w10857_ ;
	wire _w10856_ ;
	wire _w10855_ ;
	wire _w10854_ ;
	wire _w10853_ ;
	wire _w10852_ ;
	wire _w10851_ ;
	wire _w10850_ ;
	wire _w10849_ ;
	wire _w10848_ ;
	wire _w10847_ ;
	wire _w10846_ ;
	wire _w10845_ ;
	wire _w10844_ ;
	wire _w10843_ ;
	wire _w10842_ ;
	wire _w10841_ ;
	wire _w10840_ ;
	wire _w10839_ ;
	wire _w10838_ ;
	wire _w10837_ ;
	wire _w10836_ ;
	wire _w10835_ ;
	wire _w10834_ ;
	wire _w10833_ ;
	wire _w10832_ ;
	wire _w10831_ ;
	wire _w10830_ ;
	wire _w10829_ ;
	wire _w10828_ ;
	wire _w10827_ ;
	wire _w10826_ ;
	wire _w10825_ ;
	wire _w10824_ ;
	wire _w10823_ ;
	wire _w10822_ ;
	wire _w10821_ ;
	wire _w10820_ ;
	wire _w10819_ ;
	wire _w10818_ ;
	wire _w10817_ ;
	wire _w10816_ ;
	wire _w10815_ ;
	wire _w10814_ ;
	wire _w10813_ ;
	wire _w10812_ ;
	wire _w10811_ ;
	wire _w10810_ ;
	wire _w10809_ ;
	wire _w10808_ ;
	wire _w10807_ ;
	wire _w10806_ ;
	wire _w10805_ ;
	wire _w10804_ ;
	wire _w10803_ ;
	wire _w10802_ ;
	wire _w10801_ ;
	wire _w10800_ ;
	wire _w10799_ ;
	wire _w10798_ ;
	wire _w10797_ ;
	wire _w10796_ ;
	wire _w10795_ ;
	wire _w10794_ ;
	wire _w10793_ ;
	wire _w10792_ ;
	wire _w10791_ ;
	wire _w10790_ ;
	wire _w10789_ ;
	wire _w10788_ ;
	wire _w10787_ ;
	wire _w10786_ ;
	wire _w10785_ ;
	wire _w10784_ ;
	wire _w10783_ ;
	wire _w10782_ ;
	wire _w10781_ ;
	wire _w10780_ ;
	wire _w10779_ ;
	wire _w10778_ ;
	wire _w10777_ ;
	wire _w10776_ ;
	wire _w10775_ ;
	wire _w10774_ ;
	wire _w10773_ ;
	wire _w10772_ ;
	wire _w10771_ ;
	wire _w10770_ ;
	wire _w10769_ ;
	wire _w10768_ ;
	wire _w10767_ ;
	wire _w10766_ ;
	wire _w10765_ ;
	wire _w10764_ ;
	wire _w10763_ ;
	wire _w10762_ ;
	wire _w10761_ ;
	wire _w10760_ ;
	wire _w10759_ ;
	wire _w10758_ ;
	wire _w10757_ ;
	wire _w10756_ ;
	wire _w10755_ ;
	wire _w10754_ ;
	wire _w10753_ ;
	wire _w10752_ ;
	wire _w10751_ ;
	wire _w10750_ ;
	wire _w10749_ ;
	wire _w10748_ ;
	wire _w10747_ ;
	wire _w10746_ ;
	wire _w10745_ ;
	wire _w10744_ ;
	wire _w10743_ ;
	wire _w10742_ ;
	wire _w10741_ ;
	wire _w10740_ ;
	wire _w10739_ ;
	wire _w10738_ ;
	wire _w10737_ ;
	wire _w10736_ ;
	wire _w10735_ ;
	wire _w10734_ ;
	wire _w10733_ ;
	wire _w10732_ ;
	wire _w10731_ ;
	wire _w10730_ ;
	wire _w10729_ ;
	wire _w10728_ ;
	wire _w10727_ ;
	wire _w10726_ ;
	wire _w10725_ ;
	wire _w10724_ ;
	wire _w10723_ ;
	wire _w10722_ ;
	wire _w10721_ ;
	wire _w10720_ ;
	wire _w10719_ ;
	wire _w10718_ ;
	wire _w10717_ ;
	wire _w10716_ ;
	wire _w10715_ ;
	wire _w10714_ ;
	wire _w10713_ ;
	wire _w10712_ ;
	wire _w10711_ ;
	wire _w10710_ ;
	wire _w10709_ ;
	wire _w10708_ ;
	wire _w10707_ ;
	wire _w10706_ ;
	wire _w10705_ ;
	wire _w10704_ ;
	wire _w10703_ ;
	wire _w10702_ ;
	wire _w10701_ ;
	wire _w10700_ ;
	wire _w10699_ ;
	wire _w10698_ ;
	wire _w10697_ ;
	wire _w10696_ ;
	wire _w10695_ ;
	wire _w10694_ ;
	wire _w10693_ ;
	wire _w10692_ ;
	wire _w10691_ ;
	wire _w10690_ ;
	wire _w10689_ ;
	wire _w10688_ ;
	wire _w10687_ ;
	wire _w10686_ ;
	wire _w10685_ ;
	wire _w10684_ ;
	wire _w10683_ ;
	wire _w10682_ ;
	wire _w10681_ ;
	wire _w10680_ ;
	wire _w10679_ ;
	wire _w10678_ ;
	wire _w10677_ ;
	wire _w10676_ ;
	wire _w10675_ ;
	wire _w10674_ ;
	wire _w10673_ ;
	wire _w10672_ ;
	wire _w10671_ ;
	wire _w10670_ ;
	wire _w10669_ ;
	wire _w10668_ ;
	wire _w10667_ ;
	wire _w10666_ ;
	wire _w10665_ ;
	wire _w10664_ ;
	wire _w10663_ ;
	wire _w10662_ ;
	wire _w10661_ ;
	wire _w10660_ ;
	wire _w10659_ ;
	wire _w10658_ ;
	wire _w10657_ ;
	wire _w10656_ ;
	wire _w10655_ ;
	wire _w10654_ ;
	wire _w10653_ ;
	wire _w10652_ ;
	wire _w10651_ ;
	wire _w10650_ ;
	wire _w10649_ ;
	wire _w10648_ ;
	wire _w10647_ ;
	wire _w10646_ ;
	wire _w10645_ ;
	wire _w10644_ ;
	wire _w10643_ ;
	wire _w10642_ ;
	wire _w10641_ ;
	wire _w10640_ ;
	wire _w10639_ ;
	wire _w10638_ ;
	wire _w10637_ ;
	wire _w10636_ ;
	wire _w10635_ ;
	wire _w10634_ ;
	wire _w10633_ ;
	wire _w10632_ ;
	wire _w10631_ ;
	wire _w10630_ ;
	wire _w10629_ ;
	wire _w10628_ ;
	wire _w10627_ ;
	wire _w10626_ ;
	wire _w10625_ ;
	wire _w10624_ ;
	wire _w10623_ ;
	wire _w10622_ ;
	wire _w10621_ ;
	wire _w10620_ ;
	wire _w10619_ ;
	wire _w10618_ ;
	wire _w10617_ ;
	wire _w10616_ ;
	wire _w10615_ ;
	wire _w10614_ ;
	wire _w10613_ ;
	wire _w10612_ ;
	wire _w10611_ ;
	wire _w10610_ ;
	wire _w10609_ ;
	wire _w10608_ ;
	wire _w10607_ ;
	wire _w10606_ ;
	wire _w10605_ ;
	wire _w10604_ ;
	wire _w10603_ ;
	wire _w10602_ ;
	wire _w10601_ ;
	wire _w10600_ ;
	wire _w10599_ ;
	wire _w10598_ ;
	wire _w10597_ ;
	wire _w10596_ ;
	wire _w10595_ ;
	wire _w10594_ ;
	wire _w10593_ ;
	wire _w10592_ ;
	wire _w10591_ ;
	wire _w10590_ ;
	wire _w10589_ ;
	wire _w10588_ ;
	wire _w10587_ ;
	wire _w10586_ ;
	wire _w10585_ ;
	wire _w10584_ ;
	wire _w10583_ ;
	wire _w10582_ ;
	wire _w10581_ ;
	wire _w10580_ ;
	wire _w10579_ ;
	wire _w10578_ ;
	wire _w10577_ ;
	wire _w10576_ ;
	wire _w10575_ ;
	wire _w10574_ ;
	wire _w10573_ ;
	wire _w10572_ ;
	wire _w10571_ ;
	wire _w10570_ ;
	wire _w10569_ ;
	wire _w10568_ ;
	wire _w10567_ ;
	wire _w10566_ ;
	wire _w10565_ ;
	wire _w10564_ ;
	wire _w10563_ ;
	wire _w10562_ ;
	wire _w10561_ ;
	wire _w10560_ ;
	wire _w10559_ ;
	wire _w10558_ ;
	wire _w10557_ ;
	wire _w10556_ ;
	wire _w10555_ ;
	wire _w10554_ ;
	wire _w10553_ ;
	wire _w10552_ ;
	wire _w10551_ ;
	wire _w10550_ ;
	wire _w10549_ ;
	wire _w10548_ ;
	wire _w10547_ ;
	wire _w10546_ ;
	wire _w10545_ ;
	wire _w10544_ ;
	wire _w10543_ ;
	wire _w10542_ ;
	wire _w10541_ ;
	wire _w10540_ ;
	wire _w10539_ ;
	wire _w10538_ ;
	wire _w10537_ ;
	wire _w10536_ ;
	wire _w10535_ ;
	wire _w10534_ ;
	wire _w10533_ ;
	wire _w10532_ ;
	wire _w10531_ ;
	wire _w10530_ ;
	wire _w10529_ ;
	wire _w10528_ ;
	wire _w10527_ ;
	wire _w10526_ ;
	wire _w10525_ ;
	wire _w10524_ ;
	wire _w10523_ ;
	wire _w10522_ ;
	wire _w10521_ ;
	wire _w10520_ ;
	wire _w10519_ ;
	wire _w10518_ ;
	wire _w10517_ ;
	wire _w10516_ ;
	wire _w10515_ ;
	wire _w10514_ ;
	wire _w10513_ ;
	wire _w10512_ ;
	wire _w10511_ ;
	wire _w10510_ ;
	wire _w10509_ ;
	wire _w10508_ ;
	wire _w10507_ ;
	wire _w10506_ ;
	wire _w10505_ ;
	wire _w10504_ ;
	wire _w10503_ ;
	wire _w10502_ ;
	wire _w10501_ ;
	wire _w10500_ ;
	wire _w10499_ ;
	wire _w10498_ ;
	wire _w10497_ ;
	wire _w10496_ ;
	wire _w10495_ ;
	wire _w10494_ ;
	wire _w10493_ ;
	wire _w10492_ ;
	wire _w10491_ ;
	wire _w10490_ ;
	wire _w10489_ ;
	wire _w10488_ ;
	wire _w10487_ ;
	wire _w10486_ ;
	wire _w10485_ ;
	wire _w10484_ ;
	wire _w10483_ ;
	wire _w10482_ ;
	wire _w10481_ ;
	wire _w10480_ ;
	wire _w10479_ ;
	wire _w10478_ ;
	wire _w10477_ ;
	wire _w10476_ ;
	wire _w10475_ ;
	wire _w10474_ ;
	wire _w10473_ ;
	wire _w10472_ ;
	wire _w10471_ ;
	wire _w10470_ ;
	wire _w10469_ ;
	wire _w10468_ ;
	wire _w10467_ ;
	wire _w10466_ ;
	wire _w10465_ ;
	wire _w10464_ ;
	wire _w10463_ ;
	wire _w10462_ ;
	wire _w10461_ ;
	wire _w10460_ ;
	wire _w10459_ ;
	wire _w10458_ ;
	wire _w10457_ ;
	wire _w10456_ ;
	wire _w10455_ ;
	wire _w10454_ ;
	wire _w10453_ ;
	wire _w10452_ ;
	wire _w10451_ ;
	wire _w10450_ ;
	wire _w10449_ ;
	wire _w10448_ ;
	wire _w10447_ ;
	wire _w10446_ ;
	wire _w10445_ ;
	wire _w10444_ ;
	wire _w10443_ ;
	wire _w10442_ ;
	wire _w10441_ ;
	wire _w10440_ ;
	wire _w10439_ ;
	wire _w10438_ ;
	wire _w10437_ ;
	wire _w10436_ ;
	wire _w10435_ ;
	wire _w10434_ ;
	wire _w10433_ ;
	wire _w10432_ ;
	wire _w10431_ ;
	wire _w10430_ ;
	wire _w10429_ ;
	wire _w10428_ ;
	wire _w10427_ ;
	wire _w10426_ ;
	wire _w10425_ ;
	wire _w10424_ ;
	wire _w10423_ ;
	wire _w10422_ ;
	wire _w10421_ ;
	wire _w10420_ ;
	wire _w10419_ ;
	wire _w10418_ ;
	wire _w10417_ ;
	wire _w10416_ ;
	wire _w10415_ ;
	wire _w10414_ ;
	wire _w10413_ ;
	wire _w10412_ ;
	wire _w10411_ ;
	wire _w10410_ ;
	wire _w10409_ ;
	wire _w10408_ ;
	wire _w10407_ ;
	wire _w10406_ ;
	wire _w10405_ ;
	wire _w10404_ ;
	wire _w10403_ ;
	wire _w10402_ ;
	wire _w10401_ ;
	wire _w10400_ ;
	wire _w10399_ ;
	wire _w10398_ ;
	wire _w10397_ ;
	wire _w10396_ ;
	wire _w10395_ ;
	wire _w10394_ ;
	wire _w10393_ ;
	wire _w10392_ ;
	wire _w10391_ ;
	wire _w10390_ ;
	wire _w10389_ ;
	wire _w10388_ ;
	wire _w10387_ ;
	wire _w10386_ ;
	wire _w10385_ ;
	wire _w10384_ ;
	wire _w10383_ ;
	wire _w10382_ ;
	wire _w10381_ ;
	wire _w10380_ ;
	wire _w10379_ ;
	wire _w10378_ ;
	wire _w10377_ ;
	wire _w10375_ ;
	wire _w10374_ ;
	wire _w10373_ ;
	wire _w10372_ ;
	wire _w10371_ ;
	wire _w10370_ ;
	wire _w10369_ ;
	wire _w10368_ ;
	wire _w10367_ ;
	wire _w10366_ ;
	wire _w10365_ ;
	wire _w10364_ ;
	wire _w10363_ ;
	wire _w10362_ ;
	wire _w10361_ ;
	wire _w10360_ ;
	wire _w10359_ ;
	wire _w10358_ ;
	wire _w10357_ ;
	wire _w10356_ ;
	wire _w10355_ ;
	wire _w10354_ ;
	wire _w10353_ ;
	wire _w10352_ ;
	wire _w10351_ ;
	wire _w10350_ ;
	wire _w10349_ ;
	wire _w10348_ ;
	wire _w10347_ ;
	wire _w10346_ ;
	wire _w10345_ ;
	wire _w10344_ ;
	wire _w10343_ ;
	wire _w10342_ ;
	wire _w10341_ ;
	wire _w10340_ ;
	wire _w10339_ ;
	wire _w10338_ ;
	wire _w10337_ ;
	wire _w10336_ ;
	wire _w10335_ ;
	wire _w10334_ ;
	wire _w10333_ ;
	wire _w10332_ ;
	wire _w10331_ ;
	wire _w10330_ ;
	wire _w10329_ ;
	wire _w10328_ ;
	wire _w10327_ ;
	wire _w10326_ ;
	wire _w10325_ ;
	wire _w10324_ ;
	wire _w10323_ ;
	wire _w10322_ ;
	wire _w10321_ ;
	wire _w10320_ ;
	wire _w10319_ ;
	wire _w10318_ ;
	wire _w10317_ ;
	wire _w10316_ ;
	wire _w10315_ ;
	wire _w10314_ ;
	wire _w10313_ ;
	wire _w10312_ ;
	wire _w10311_ ;
	wire _w10310_ ;
	wire _w10309_ ;
	wire _w10308_ ;
	wire _w10307_ ;
	wire _w10306_ ;
	wire _w10305_ ;
	wire _w10304_ ;
	wire _w10303_ ;
	wire _w10302_ ;
	wire _w10301_ ;
	wire _w10300_ ;
	wire _w10299_ ;
	wire _w10298_ ;
	wire _w10297_ ;
	wire _w10296_ ;
	wire _w10295_ ;
	wire _w10294_ ;
	wire _w10293_ ;
	wire _w10292_ ;
	wire _w10291_ ;
	wire _w10290_ ;
	wire _w10289_ ;
	wire _w10288_ ;
	wire _w10287_ ;
	wire _w10286_ ;
	wire _w10285_ ;
	wire _w10284_ ;
	wire _w10283_ ;
	wire _w10282_ ;
	wire _w10281_ ;
	wire _w10280_ ;
	wire _w10279_ ;
	wire _w10278_ ;
	wire _w10277_ ;
	wire _w10276_ ;
	wire _w10275_ ;
	wire _w10274_ ;
	wire _w10273_ ;
	wire _w10272_ ;
	wire _w10271_ ;
	wire _w10270_ ;
	wire _w10269_ ;
	wire _w10268_ ;
	wire _w10267_ ;
	wire _w10266_ ;
	wire _w10265_ ;
	wire _w10264_ ;
	wire _w10263_ ;
	wire _w10262_ ;
	wire _w10261_ ;
	wire _w10260_ ;
	wire _w10259_ ;
	wire _w10258_ ;
	wire _w10257_ ;
	wire _w10256_ ;
	wire _w10255_ ;
	wire _w10254_ ;
	wire _w10253_ ;
	wire _w10252_ ;
	wire _w10251_ ;
	wire _w10250_ ;
	wire _w10249_ ;
	wire _w10248_ ;
	wire _w10247_ ;
	wire _w10246_ ;
	wire _w10245_ ;
	wire _w10244_ ;
	wire _w10243_ ;
	wire _w10242_ ;
	wire _w10241_ ;
	wire _w10240_ ;
	wire _w10239_ ;
	wire _w10238_ ;
	wire _w10237_ ;
	wire _w10236_ ;
	wire _w10235_ ;
	wire _w10234_ ;
	wire _w10233_ ;
	wire _w10232_ ;
	wire _w10231_ ;
	wire _w10230_ ;
	wire _w10229_ ;
	wire _w10228_ ;
	wire _w10227_ ;
	wire _w10226_ ;
	wire _w10225_ ;
	wire _w10224_ ;
	wire _w10223_ ;
	wire _w10222_ ;
	wire _w10221_ ;
	wire _w10220_ ;
	wire _w10219_ ;
	wire _w10218_ ;
	wire _w10217_ ;
	wire _w10216_ ;
	wire _w10215_ ;
	wire _w10214_ ;
	wire _w10213_ ;
	wire _w10212_ ;
	wire _w10211_ ;
	wire _w10210_ ;
	wire _w10209_ ;
	wire _w10208_ ;
	wire _w10207_ ;
	wire _w10206_ ;
	wire _w10205_ ;
	wire _w10204_ ;
	wire _w10203_ ;
	wire _w10202_ ;
	wire _w10201_ ;
	wire _w10200_ ;
	wire _w10199_ ;
	wire _w10198_ ;
	wire _w10197_ ;
	wire _w10196_ ;
	wire _w10195_ ;
	wire _w10194_ ;
	wire _w10193_ ;
	wire _w10192_ ;
	wire _w10191_ ;
	wire _w10190_ ;
	wire _w10189_ ;
	wire _w10188_ ;
	wire _w10187_ ;
	wire _w10186_ ;
	wire _w10185_ ;
	wire _w10184_ ;
	wire _w10183_ ;
	wire _w10182_ ;
	wire _w10181_ ;
	wire _w10180_ ;
	wire _w10179_ ;
	wire _w10178_ ;
	wire _w10177_ ;
	wire _w10176_ ;
	wire _w10175_ ;
	wire _w10174_ ;
	wire _w10173_ ;
	wire _w10172_ ;
	wire _w10171_ ;
	wire _w10170_ ;
	wire _w10169_ ;
	wire _w10168_ ;
	wire _w10167_ ;
	wire _w10166_ ;
	wire _w10165_ ;
	wire _w10164_ ;
	wire _w10163_ ;
	wire _w10162_ ;
	wire _w10161_ ;
	wire _w10160_ ;
	wire _w10159_ ;
	wire _w10158_ ;
	wire _w10157_ ;
	wire _w10156_ ;
	wire _w10155_ ;
	wire _w10154_ ;
	wire _w10153_ ;
	wire _w10152_ ;
	wire _w10151_ ;
	wire _w10150_ ;
	wire _w10149_ ;
	wire _w10148_ ;
	wire _w10147_ ;
	wire _w10146_ ;
	wire _w10145_ ;
	wire _w10144_ ;
	wire _w10143_ ;
	wire _w10142_ ;
	wire _w10141_ ;
	wire _w10140_ ;
	wire _w10139_ ;
	wire _w10138_ ;
	wire _w10137_ ;
	wire _w10136_ ;
	wire _w10135_ ;
	wire _w10134_ ;
	wire _w10133_ ;
	wire _w10132_ ;
	wire _w10131_ ;
	wire _w10130_ ;
	wire _w10129_ ;
	wire _w10128_ ;
	wire _w10127_ ;
	wire _w10126_ ;
	wire _w10125_ ;
	wire _w10124_ ;
	wire _w10123_ ;
	wire _w10122_ ;
	wire _w10121_ ;
	wire _w10120_ ;
	wire _w10119_ ;
	wire _w10118_ ;
	wire _w10117_ ;
	wire _w10116_ ;
	wire _w10115_ ;
	wire _w10114_ ;
	wire _w10113_ ;
	wire _w10112_ ;
	wire _w10111_ ;
	wire _w10110_ ;
	wire _w10109_ ;
	wire _w10108_ ;
	wire _w10107_ ;
	wire _w10106_ ;
	wire _w10105_ ;
	wire _w10104_ ;
	wire _w10103_ ;
	wire _w10102_ ;
	wire _w10101_ ;
	wire _w10100_ ;
	wire _w10099_ ;
	wire _w10098_ ;
	wire _w10097_ ;
	wire _w10096_ ;
	wire _w10095_ ;
	wire _w10094_ ;
	wire _w10093_ ;
	wire _w10092_ ;
	wire _w10091_ ;
	wire _w10090_ ;
	wire _w10089_ ;
	wire _w10088_ ;
	wire _w10087_ ;
	wire _w10086_ ;
	wire _w10085_ ;
	wire _w10084_ ;
	wire _w10083_ ;
	wire _w10082_ ;
	wire _w10081_ ;
	wire _w10080_ ;
	wire _w10079_ ;
	wire _w10078_ ;
	wire _w10077_ ;
	wire _w10076_ ;
	wire _w10075_ ;
	wire _w10074_ ;
	wire _w10073_ ;
	wire _w10072_ ;
	wire _w10071_ ;
	wire _w10070_ ;
	wire _w10069_ ;
	wire _w10068_ ;
	wire _w10067_ ;
	wire _w10066_ ;
	wire _w10065_ ;
	wire _w10064_ ;
	wire _w10063_ ;
	wire _w10062_ ;
	wire _w10061_ ;
	wire _w10060_ ;
	wire _w10059_ ;
	wire _w10058_ ;
	wire _w10057_ ;
	wire _w10056_ ;
	wire _w10055_ ;
	wire _w10054_ ;
	wire _w10053_ ;
	wire _w10052_ ;
	wire _w10051_ ;
	wire _w10050_ ;
	wire _w10049_ ;
	wire _w10048_ ;
	wire _w10047_ ;
	wire _w10046_ ;
	wire _w10045_ ;
	wire _w10044_ ;
	wire _w10043_ ;
	wire _w10042_ ;
	wire _w10041_ ;
	wire _w10040_ ;
	wire _w10039_ ;
	wire _w10038_ ;
	wire _w10037_ ;
	wire _w10036_ ;
	wire _w10035_ ;
	wire _w10034_ ;
	wire _w10033_ ;
	wire _w10032_ ;
	wire _w10031_ ;
	wire _w10030_ ;
	wire _w10029_ ;
	wire _w10028_ ;
	wire _w10027_ ;
	wire _w10026_ ;
	wire _w10025_ ;
	wire _w10024_ ;
	wire _w10023_ ;
	wire _w10022_ ;
	wire _w10021_ ;
	wire _w10020_ ;
	wire _w10019_ ;
	wire _w10018_ ;
	wire _w10017_ ;
	wire _w10016_ ;
	wire _w10015_ ;
	wire _w10014_ ;
	wire _w10013_ ;
	wire _w10012_ ;
	wire _w10011_ ;
	wire _w10010_ ;
	wire _w10009_ ;
	wire _w10008_ ;
	wire _w10007_ ;
	wire _w10006_ ;
	wire _w10005_ ;
	wire _w10004_ ;
	wire _w10003_ ;
	wire _w10002_ ;
	wire _w10001_ ;
	wire _w10000_ ;
	wire _w9999_ ;
	wire _w9998_ ;
	wire _w9997_ ;
	wire _w9996_ ;
	wire _w9995_ ;
	wire _w9994_ ;
	wire _w9993_ ;
	wire _w9992_ ;
	wire _w9991_ ;
	wire _w9990_ ;
	wire _w9989_ ;
	wire _w9988_ ;
	wire _w9987_ ;
	wire _w9986_ ;
	wire _w9985_ ;
	wire _w9984_ ;
	wire _w9983_ ;
	wire _w9982_ ;
	wire _w9981_ ;
	wire _w9980_ ;
	wire _w9979_ ;
	wire _w9978_ ;
	wire _w9977_ ;
	wire _w9976_ ;
	wire _w9975_ ;
	wire _w9974_ ;
	wire _w9973_ ;
	wire _w9972_ ;
	wire _w9971_ ;
	wire _w9970_ ;
	wire _w9969_ ;
	wire _w9968_ ;
	wire _w9967_ ;
	wire _w9966_ ;
	wire _w9965_ ;
	wire _w9964_ ;
	wire _w9963_ ;
	wire _w9962_ ;
	wire _w9961_ ;
	wire _w9960_ ;
	wire _w9959_ ;
	wire _w9958_ ;
	wire _w9957_ ;
	wire _w9956_ ;
	wire _w9955_ ;
	wire _w9954_ ;
	wire _w9953_ ;
	wire _w9952_ ;
	wire _w9951_ ;
	wire _w9950_ ;
	wire _w9949_ ;
	wire _w9948_ ;
	wire _w9947_ ;
	wire _w9946_ ;
	wire _w9945_ ;
	wire _w9944_ ;
	wire _w9943_ ;
	wire _w9942_ ;
	wire _w9941_ ;
	wire _w9940_ ;
	wire _w9939_ ;
	wire _w9938_ ;
	wire _w9937_ ;
	wire _w9936_ ;
	wire _w9935_ ;
	wire _w9934_ ;
	wire _w9933_ ;
	wire _w9932_ ;
	wire _w9931_ ;
	wire _w9930_ ;
	wire _w9929_ ;
	wire _w9928_ ;
	wire _w9927_ ;
	wire _w9926_ ;
	wire _w9925_ ;
	wire _w9924_ ;
	wire _w9923_ ;
	wire _w9922_ ;
	wire _w9921_ ;
	wire _w9920_ ;
	wire _w9919_ ;
	wire _w9918_ ;
	wire _w9917_ ;
	wire _w9916_ ;
	wire _w9915_ ;
	wire _w9914_ ;
	wire _w9913_ ;
	wire _w9912_ ;
	wire _w9911_ ;
	wire _w9910_ ;
	wire _w9909_ ;
	wire _w9908_ ;
	wire _w9907_ ;
	wire _w9906_ ;
	wire _w9905_ ;
	wire _w9904_ ;
	wire _w9903_ ;
	wire _w9902_ ;
	wire _w9901_ ;
	wire _w9900_ ;
	wire _w9899_ ;
	wire _w9898_ ;
	wire _w9897_ ;
	wire _w9896_ ;
	wire _w9895_ ;
	wire _w9894_ ;
	wire _w9893_ ;
	wire _w9892_ ;
	wire _w9891_ ;
	wire _w9890_ ;
	wire _w9889_ ;
	wire _w9888_ ;
	wire _w9887_ ;
	wire _w9886_ ;
	wire _w9885_ ;
	wire _w9884_ ;
	wire _w9883_ ;
	wire _w9882_ ;
	wire _w9881_ ;
	wire _w9880_ ;
	wire _w9879_ ;
	wire _w9878_ ;
	wire _w9877_ ;
	wire _w9876_ ;
	wire _w9875_ ;
	wire _w9874_ ;
	wire _w9873_ ;
	wire _w9872_ ;
	wire _w9871_ ;
	wire _w9870_ ;
	wire _w9869_ ;
	wire _w9868_ ;
	wire _w9867_ ;
	wire _w9866_ ;
	wire _w9865_ ;
	wire _w9864_ ;
	wire _w9863_ ;
	wire _w9862_ ;
	wire _w9861_ ;
	wire _w9860_ ;
	wire _w9859_ ;
	wire _w9858_ ;
	wire _w9857_ ;
	wire _w9856_ ;
	wire _w9855_ ;
	wire _w9854_ ;
	wire _w9853_ ;
	wire _w9852_ ;
	wire _w9851_ ;
	wire _w9850_ ;
	wire _w9849_ ;
	wire _w9848_ ;
	wire _w9847_ ;
	wire _w9846_ ;
	wire _w9845_ ;
	wire _w9844_ ;
	wire _w9843_ ;
	wire _w9842_ ;
	wire _w9841_ ;
	wire _w9840_ ;
	wire _w9839_ ;
	wire _w9838_ ;
	wire _w9837_ ;
	wire _w9836_ ;
	wire _w9835_ ;
	wire _w9834_ ;
	wire _w9833_ ;
	wire _w9832_ ;
	wire _w9831_ ;
	wire _w9830_ ;
	wire _w9829_ ;
	wire _w9828_ ;
	wire _w9827_ ;
	wire _w9826_ ;
	wire _w9825_ ;
	wire _w9824_ ;
	wire _w9823_ ;
	wire _w9822_ ;
	wire _w9821_ ;
	wire _w9820_ ;
	wire _w9819_ ;
	wire _w9818_ ;
	wire _w9817_ ;
	wire _w9816_ ;
	wire _w9815_ ;
	wire _w9814_ ;
	wire _w9813_ ;
	wire _w9812_ ;
	wire _w9811_ ;
	wire _w9810_ ;
	wire _w9809_ ;
	wire _w9808_ ;
	wire _w9807_ ;
	wire _w9806_ ;
	wire _w9805_ ;
	wire _w9804_ ;
	wire _w9803_ ;
	wire _w9802_ ;
	wire _w9801_ ;
	wire _w9800_ ;
	wire _w9799_ ;
	wire _w9798_ ;
	wire _w9797_ ;
	wire _w9796_ ;
	wire _w9795_ ;
	wire _w9794_ ;
	wire _w9793_ ;
	wire _w9792_ ;
	wire _w9791_ ;
	wire _w9790_ ;
	wire _w9789_ ;
	wire _w9788_ ;
	wire _w9787_ ;
	wire _w9786_ ;
	wire _w9785_ ;
	wire _w9784_ ;
	wire _w9783_ ;
	wire _w9782_ ;
	wire _w9781_ ;
	wire _w9780_ ;
	wire _w9779_ ;
	wire _w9778_ ;
	wire _w9777_ ;
	wire _w9776_ ;
	wire _w9775_ ;
	wire _w9774_ ;
	wire _w9773_ ;
	wire _w9772_ ;
	wire _w9771_ ;
	wire _w9770_ ;
	wire _w9769_ ;
	wire _w9768_ ;
	wire _w9767_ ;
	wire _w9766_ ;
	wire _w9765_ ;
	wire _w9764_ ;
	wire _w9763_ ;
	wire _w9762_ ;
	wire _w9761_ ;
	wire _w9760_ ;
	wire _w9759_ ;
	wire _w9758_ ;
	wire _w9757_ ;
	wire _w9756_ ;
	wire _w9755_ ;
	wire _w9754_ ;
	wire _w9753_ ;
	wire _w9752_ ;
	wire _w9751_ ;
	wire _w9750_ ;
	wire _w9749_ ;
	wire _w9748_ ;
	wire _w9747_ ;
	wire _w9746_ ;
	wire _w9745_ ;
	wire _w9744_ ;
	wire _w9743_ ;
	wire _w9742_ ;
	wire _w9741_ ;
	wire _w9740_ ;
	wire _w9739_ ;
	wire _w9738_ ;
	wire _w9737_ ;
	wire _w9736_ ;
	wire _w9735_ ;
	wire _w9734_ ;
	wire _w9733_ ;
	wire _w9732_ ;
	wire _w9731_ ;
	wire _w9730_ ;
	wire _w9729_ ;
	wire _w9728_ ;
	wire _w9727_ ;
	wire _w9726_ ;
	wire _w9725_ ;
	wire _w9724_ ;
	wire _w9723_ ;
	wire _w9722_ ;
	wire _w9721_ ;
	wire _w9720_ ;
	wire _w9719_ ;
	wire _w9718_ ;
	wire _w9717_ ;
	wire _w9716_ ;
	wire _w9715_ ;
	wire _w9714_ ;
	wire _w9713_ ;
	wire _w9712_ ;
	wire _w9711_ ;
	wire _w9710_ ;
	wire _w9709_ ;
	wire _w9708_ ;
	wire _w9707_ ;
	wire _w9706_ ;
	wire _w9705_ ;
	wire _w9704_ ;
	wire _w9703_ ;
	wire _w9702_ ;
	wire _w9701_ ;
	wire _w9700_ ;
	wire _w9699_ ;
	wire _w9698_ ;
	wire _w9697_ ;
	wire _w9696_ ;
	wire _w9695_ ;
	wire _w9694_ ;
	wire _w9693_ ;
	wire _w9692_ ;
	wire _w9691_ ;
	wire _w9690_ ;
	wire _w9689_ ;
	wire _w9688_ ;
	wire _w9687_ ;
	wire _w9686_ ;
	wire _w9685_ ;
	wire _w9684_ ;
	wire _w9683_ ;
	wire _w9682_ ;
	wire _w9681_ ;
	wire _w9680_ ;
	wire _w9679_ ;
	wire _w9678_ ;
	wire _w9677_ ;
	wire _w9676_ ;
	wire _w9675_ ;
	wire _w9674_ ;
	wire _w9673_ ;
	wire _w9672_ ;
	wire _w9671_ ;
	wire _w9670_ ;
	wire _w9669_ ;
	wire _w9668_ ;
	wire _w9667_ ;
	wire _w9666_ ;
	wire _w9665_ ;
	wire _w9664_ ;
	wire _w9663_ ;
	wire _w9662_ ;
	wire _w9661_ ;
	wire _w9660_ ;
	wire _w9659_ ;
	wire _w9658_ ;
	wire _w9657_ ;
	wire _w9656_ ;
	wire _w9655_ ;
	wire _w9654_ ;
	wire _w9653_ ;
	wire _w9652_ ;
	wire _w9651_ ;
	wire _w9650_ ;
	wire _w9649_ ;
	wire _w9648_ ;
	wire _w9647_ ;
	wire _w9646_ ;
	wire _w9645_ ;
	wire _w9644_ ;
	wire _w9643_ ;
	wire _w9642_ ;
	wire _w9641_ ;
	wire _w9640_ ;
	wire _w9639_ ;
	wire _w9638_ ;
	wire _w9637_ ;
	wire _w9636_ ;
	wire _w9635_ ;
	wire _w9634_ ;
	wire _w9633_ ;
	wire _w9632_ ;
	wire _w9631_ ;
	wire _w9630_ ;
	wire _w9629_ ;
	wire _w9628_ ;
	wire _w9627_ ;
	wire _w9626_ ;
	wire _w9625_ ;
	wire _w9624_ ;
	wire _w9623_ ;
	wire _w9622_ ;
	wire _w9621_ ;
	wire _w9620_ ;
	wire _w9619_ ;
	wire _w9618_ ;
	wire _w9617_ ;
	wire _w9616_ ;
	wire _w9615_ ;
	wire _w9614_ ;
	wire _w9613_ ;
	wire _w9612_ ;
	wire _w9611_ ;
	wire _w9610_ ;
	wire _w9609_ ;
	wire _w9608_ ;
	wire _w9607_ ;
	wire _w9606_ ;
	wire _w9605_ ;
	wire _w9604_ ;
	wire _w9603_ ;
	wire _w9602_ ;
	wire _w9601_ ;
	wire _w9600_ ;
	wire _w9599_ ;
	wire _w9598_ ;
	wire _w9597_ ;
	wire _w9596_ ;
	wire _w9595_ ;
	wire _w9594_ ;
	wire _w9593_ ;
	wire _w9592_ ;
	wire _w9591_ ;
	wire _w9590_ ;
	wire _w9589_ ;
	wire _w9588_ ;
	wire _w9587_ ;
	wire _w9586_ ;
	wire _w9585_ ;
	wire _w9584_ ;
	wire _w9583_ ;
	wire _w9582_ ;
	wire _w9581_ ;
	wire _w9580_ ;
	wire _w9579_ ;
	wire _w9578_ ;
	wire _w9577_ ;
	wire _w9576_ ;
	wire _w9575_ ;
	wire _w9574_ ;
	wire _w9573_ ;
	wire _w9572_ ;
	wire _w9571_ ;
	wire _w9570_ ;
	wire _w9569_ ;
	wire _w9568_ ;
	wire _w9567_ ;
	wire _w9566_ ;
	wire _w9565_ ;
	wire _w9564_ ;
	wire _w9563_ ;
	wire _w9562_ ;
	wire _w9561_ ;
	wire _w9560_ ;
	wire _w9559_ ;
	wire _w9558_ ;
	wire _w9557_ ;
	wire _w9556_ ;
	wire _w9555_ ;
	wire _w9554_ ;
	wire _w9553_ ;
	wire _w9552_ ;
	wire _w9551_ ;
	wire _w9550_ ;
	wire _w9549_ ;
	wire _w9548_ ;
	wire _w9547_ ;
	wire _w9546_ ;
	wire _w9545_ ;
	wire _w9544_ ;
	wire _w9543_ ;
	wire _w9542_ ;
	wire _w9541_ ;
	wire _w9540_ ;
	wire _w9539_ ;
	wire _w9538_ ;
	wire _w9537_ ;
	wire _w9536_ ;
	wire _w9535_ ;
	wire _w9534_ ;
	wire _w9533_ ;
	wire _w9532_ ;
	wire _w9531_ ;
	wire _w9530_ ;
	wire _w9529_ ;
	wire _w9528_ ;
	wire _w9527_ ;
	wire _w9526_ ;
	wire _w9525_ ;
	wire _w9524_ ;
	wire _w9523_ ;
	wire _w9522_ ;
	wire _w9521_ ;
	wire _w9520_ ;
	wire _w9519_ ;
	wire _w9518_ ;
	wire _w9517_ ;
	wire _w9516_ ;
	wire _w9515_ ;
	wire _w9514_ ;
	wire _w9513_ ;
	wire _w9512_ ;
	wire _w9511_ ;
	wire _w9510_ ;
	wire _w9509_ ;
	wire _w9508_ ;
	wire _w9507_ ;
	wire _w9506_ ;
	wire _w9505_ ;
	wire _w9504_ ;
	wire _w9503_ ;
	wire _w9502_ ;
	wire _w9501_ ;
	wire _w9500_ ;
	wire _w9499_ ;
	wire _w9498_ ;
	wire _w9497_ ;
	wire _w9496_ ;
	wire _w9495_ ;
	wire _w9494_ ;
	wire _w9493_ ;
	wire _w9492_ ;
	wire _w9491_ ;
	wire _w9490_ ;
	wire _w9489_ ;
	wire _w9488_ ;
	wire _w9487_ ;
	wire _w9486_ ;
	wire _w9485_ ;
	wire _w9484_ ;
	wire _w9483_ ;
	wire _w9482_ ;
	wire _w9481_ ;
	wire _w9480_ ;
	wire _w9479_ ;
	wire _w9478_ ;
	wire _w9477_ ;
	wire _w9476_ ;
	wire _w9475_ ;
	wire _w9474_ ;
	wire _w9473_ ;
	wire _w9472_ ;
	wire _w9471_ ;
	wire _w9470_ ;
	wire _w9469_ ;
	wire _w9468_ ;
	wire _w9467_ ;
	wire _w9466_ ;
	wire _w9465_ ;
	wire _w9464_ ;
	wire _w9463_ ;
	wire _w9462_ ;
	wire _w9461_ ;
	wire _w9460_ ;
	wire _w9459_ ;
	wire _w9458_ ;
	wire _w9457_ ;
	wire _w9456_ ;
	wire _w9455_ ;
	wire _w9454_ ;
	wire _w9453_ ;
	wire _w9452_ ;
	wire _w9451_ ;
	wire _w9450_ ;
	wire _w9449_ ;
	wire _w9448_ ;
	wire _w9447_ ;
	wire _w9446_ ;
	wire _w9445_ ;
	wire _w9444_ ;
	wire _w9443_ ;
	wire _w9442_ ;
	wire _w9441_ ;
	wire _w9440_ ;
	wire _w9439_ ;
	wire _w9438_ ;
	wire _w9437_ ;
	wire _w9436_ ;
	wire _w9435_ ;
	wire _w9434_ ;
	wire _w9433_ ;
	wire _w9432_ ;
	wire _w9431_ ;
	wire _w9430_ ;
	wire _w9429_ ;
	wire _w9428_ ;
	wire _w9427_ ;
	wire _w9426_ ;
	wire _w9425_ ;
	wire _w9424_ ;
	wire _w9423_ ;
	wire _w9422_ ;
	wire _w9421_ ;
	wire _w9420_ ;
	wire _w9419_ ;
	wire _w9418_ ;
	wire _w9417_ ;
	wire _w9416_ ;
	wire _w9415_ ;
	wire _w9414_ ;
	wire _w9413_ ;
	wire _w9412_ ;
	wire _w9411_ ;
	wire _w9410_ ;
	wire _w9409_ ;
	wire _w9408_ ;
	wire _w9407_ ;
	wire _w9406_ ;
	wire _w9405_ ;
	wire _w9404_ ;
	wire _w9403_ ;
	wire _w9402_ ;
	wire _w9401_ ;
	wire _w9400_ ;
	wire _w9399_ ;
	wire _w9398_ ;
	wire _w9397_ ;
	wire _w9396_ ;
	wire _w9395_ ;
	wire _w9394_ ;
	wire _w9393_ ;
	wire _w9392_ ;
	wire _w9391_ ;
	wire _w9390_ ;
	wire _w9389_ ;
	wire _w9388_ ;
	wire _w9387_ ;
	wire _w9386_ ;
	wire _w9385_ ;
	wire _w9384_ ;
	wire _w9383_ ;
	wire _w9382_ ;
	wire _w9381_ ;
	wire _w9380_ ;
	wire _w9379_ ;
	wire _w9378_ ;
	wire _w9377_ ;
	wire _w9376_ ;
	wire _w9375_ ;
	wire _w9374_ ;
	wire _w9373_ ;
	wire _w9372_ ;
	wire _w9371_ ;
	wire _w9370_ ;
	wire _w9369_ ;
	wire _w9368_ ;
	wire _w9367_ ;
	wire _w9366_ ;
	wire _w9365_ ;
	wire _w9364_ ;
	wire _w9363_ ;
	wire _w9362_ ;
	wire _w9361_ ;
	wire _w9360_ ;
	wire _w9359_ ;
	wire _w9358_ ;
	wire _w9357_ ;
	wire _w9356_ ;
	wire _w9355_ ;
	wire _w9354_ ;
	wire _w9353_ ;
	wire _w9352_ ;
	wire _w9351_ ;
	wire _w9350_ ;
	wire _w9349_ ;
	wire _w9348_ ;
	wire _w9347_ ;
	wire _w9346_ ;
	wire _w9345_ ;
	wire _w9344_ ;
	wire _w9343_ ;
	wire _w9342_ ;
	wire _w9341_ ;
	wire _w9340_ ;
	wire _w9339_ ;
	wire _w9338_ ;
	wire _w9337_ ;
	wire _w9336_ ;
	wire _w9335_ ;
	wire _w9334_ ;
	wire _w9333_ ;
	wire _w9332_ ;
	wire _w9331_ ;
	wire _w9330_ ;
	wire _w9329_ ;
	wire _w9328_ ;
	wire _w9327_ ;
	wire _w9326_ ;
	wire _w9325_ ;
	wire _w9324_ ;
	wire _w9323_ ;
	wire _w9322_ ;
	wire _w9321_ ;
	wire _w9320_ ;
	wire _w9319_ ;
	wire _w9318_ ;
	wire _w9317_ ;
	wire _w9316_ ;
	wire _w9315_ ;
	wire _w9314_ ;
	wire _w9313_ ;
	wire _w9312_ ;
	wire _w9311_ ;
	wire _w9310_ ;
	wire _w9309_ ;
	wire _w9308_ ;
	wire _w9307_ ;
	wire _w9306_ ;
	wire _w9305_ ;
	wire _w9304_ ;
	wire _w9303_ ;
	wire _w9302_ ;
	wire _w9301_ ;
	wire _w9300_ ;
	wire _w9299_ ;
	wire _w9298_ ;
	wire _w9297_ ;
	wire _w9296_ ;
	wire _w9295_ ;
	wire _w9294_ ;
	wire _w9293_ ;
	wire _w9292_ ;
	wire _w9291_ ;
	wire _w9290_ ;
	wire _w9289_ ;
	wire _w9288_ ;
	wire _w9287_ ;
	wire _w9286_ ;
	wire _w9285_ ;
	wire _w9284_ ;
	wire _w9283_ ;
	wire _w9282_ ;
	wire _w9281_ ;
	wire _w9280_ ;
	wire _w9279_ ;
	wire _w9278_ ;
	wire _w9277_ ;
	wire _w9276_ ;
	wire _w9275_ ;
	wire _w9274_ ;
	wire _w9273_ ;
	wire _w9272_ ;
	wire _w9271_ ;
	wire _w9270_ ;
	wire _w9269_ ;
	wire _w9268_ ;
	wire _w9267_ ;
	wire _w9266_ ;
	wire _w9265_ ;
	wire _w9264_ ;
	wire _w9263_ ;
	wire _w9262_ ;
	wire _w9261_ ;
	wire _w9260_ ;
	wire _w9259_ ;
	wire _w9258_ ;
	wire _w9257_ ;
	wire _w9256_ ;
	wire _w9255_ ;
	wire _w9254_ ;
	wire _w9253_ ;
	wire _w9252_ ;
	wire _w9251_ ;
	wire _w9250_ ;
	wire _w9249_ ;
	wire _w9248_ ;
	wire _w9247_ ;
	wire _w9246_ ;
	wire _w9245_ ;
	wire _w9244_ ;
	wire _w9243_ ;
	wire _w9242_ ;
	wire _w9241_ ;
	wire _w9240_ ;
	wire _w9239_ ;
	wire _w9238_ ;
	wire _w9237_ ;
	wire _w9236_ ;
	wire _w9235_ ;
	wire _w9234_ ;
	wire _w9233_ ;
	wire _w9232_ ;
	wire _w9231_ ;
	wire _w9230_ ;
	wire _w9229_ ;
	wire _w9228_ ;
	wire _w9227_ ;
	wire _w9226_ ;
	wire _w9225_ ;
	wire _w9224_ ;
	wire _w9223_ ;
	wire _w9222_ ;
	wire _w9221_ ;
	wire _w9220_ ;
	wire _w9219_ ;
	wire _w9218_ ;
	wire _w9217_ ;
	wire _w9216_ ;
	wire _w9215_ ;
	wire _w9214_ ;
	wire _w9213_ ;
	wire _w9212_ ;
	wire _w9211_ ;
	wire _w9210_ ;
	wire _w9209_ ;
	wire _w9208_ ;
	wire _w9207_ ;
	wire _w9206_ ;
	wire _w9205_ ;
	wire _w9204_ ;
	wire _w9203_ ;
	wire _w9202_ ;
	wire _w9201_ ;
	wire _w9200_ ;
	wire _w9199_ ;
	wire _w9198_ ;
	wire _w9197_ ;
	wire _w9196_ ;
	wire _w9195_ ;
	wire _w9194_ ;
	wire _w9193_ ;
	wire _w9192_ ;
	wire _w9191_ ;
	wire _w9190_ ;
	wire _w9189_ ;
	wire _w9188_ ;
	wire _w9187_ ;
	wire _w9186_ ;
	wire _w9185_ ;
	wire _w9184_ ;
	wire _w9183_ ;
	wire _w9182_ ;
	wire _w9181_ ;
	wire _w9180_ ;
	wire _w9179_ ;
	wire _w9178_ ;
	wire _w9177_ ;
	wire _w9176_ ;
	wire _w9175_ ;
	wire _w9174_ ;
	wire _w9173_ ;
	wire _w9172_ ;
	wire _w9171_ ;
	wire _w9170_ ;
	wire _w9169_ ;
	wire _w9168_ ;
	wire _w9167_ ;
	wire _w9166_ ;
	wire _w9165_ ;
	wire _w9164_ ;
	wire _w9163_ ;
	wire _w9162_ ;
	wire _w9161_ ;
	wire _w9160_ ;
	wire _w9159_ ;
	wire _w9158_ ;
	wire _w9157_ ;
	wire _w9156_ ;
	wire _w9155_ ;
	wire _w9154_ ;
	wire _w9153_ ;
	wire _w9152_ ;
	wire _w9151_ ;
	wire _w9150_ ;
	wire _w9149_ ;
	wire _w9148_ ;
	wire _w9147_ ;
	wire _w9146_ ;
	wire _w9145_ ;
	wire _w9144_ ;
	wire _w9143_ ;
	wire _w9142_ ;
	wire _w9141_ ;
	wire _w9140_ ;
	wire _w9139_ ;
	wire _w9138_ ;
	wire _w9137_ ;
	wire _w9136_ ;
	wire _w9135_ ;
	wire _w9134_ ;
	wire _w9133_ ;
	wire _w9132_ ;
	wire _w9131_ ;
	wire _w9130_ ;
	wire _w9129_ ;
	wire _w9128_ ;
	wire _w9127_ ;
	wire _w9126_ ;
	wire _w9125_ ;
	wire _w9124_ ;
	wire _w9123_ ;
	wire _w9122_ ;
	wire _w9121_ ;
	wire _w9120_ ;
	wire _w9119_ ;
	wire _w9118_ ;
	wire _w9117_ ;
	wire _w9116_ ;
	wire _w9115_ ;
	wire _w9114_ ;
	wire _w9113_ ;
	wire _w9112_ ;
	wire _w9111_ ;
	wire _w9110_ ;
	wire _w9109_ ;
	wire _w9108_ ;
	wire _w9107_ ;
	wire _w9106_ ;
	wire _w9105_ ;
	wire _w9104_ ;
	wire _w9103_ ;
	wire _w9102_ ;
	wire _w9101_ ;
	wire _w9100_ ;
	wire _w9099_ ;
	wire _w9098_ ;
	wire _w9097_ ;
	wire _w9096_ ;
	wire _w9095_ ;
	wire _w9094_ ;
	wire _w9093_ ;
	wire _w9092_ ;
	wire _w9091_ ;
	wire _w9090_ ;
	wire _w9089_ ;
	wire _w9088_ ;
	wire _w9087_ ;
	wire _w9086_ ;
	wire _w9085_ ;
	wire _w9084_ ;
	wire _w9083_ ;
	wire _w9082_ ;
	wire _w9081_ ;
	wire _w9080_ ;
	wire _w9079_ ;
	wire _w9078_ ;
	wire _w9077_ ;
	wire _w9076_ ;
	wire _w9075_ ;
	wire _w9074_ ;
	wire _w9073_ ;
	wire _w9072_ ;
	wire _w9071_ ;
	wire _w9070_ ;
	wire _w9069_ ;
	wire _w9068_ ;
	wire _w9067_ ;
	wire _w9066_ ;
	wire _w9065_ ;
	wire _w9064_ ;
	wire _w9063_ ;
	wire _w9062_ ;
	wire _w9061_ ;
	wire _w9060_ ;
	wire _w9059_ ;
	wire _w9058_ ;
	wire _w9057_ ;
	wire _w9056_ ;
	wire _w9055_ ;
	wire _w9054_ ;
	wire _w9053_ ;
	wire _w9052_ ;
	wire _w9051_ ;
	wire _w9050_ ;
	wire _w9049_ ;
	wire _w9048_ ;
	wire _w9047_ ;
	wire _w9046_ ;
	wire _w9045_ ;
	wire _w9044_ ;
	wire _w9043_ ;
	wire _w9042_ ;
	wire _w9041_ ;
	wire _w9040_ ;
	wire _w9039_ ;
	wire _w9038_ ;
	wire _w9037_ ;
	wire _w9036_ ;
	wire _w9035_ ;
	wire _w9034_ ;
	wire _w9033_ ;
	wire _w9032_ ;
	wire _w9031_ ;
	wire _w9030_ ;
	wire _w9029_ ;
	wire _w9028_ ;
	wire _w9027_ ;
	wire _w9026_ ;
	wire _w9025_ ;
	wire _w9024_ ;
	wire _w9023_ ;
	wire _w9022_ ;
	wire _w9021_ ;
	wire _w9020_ ;
	wire _w9019_ ;
	wire _w9018_ ;
	wire _w9017_ ;
	wire _w9016_ ;
	wire _w9015_ ;
	wire _w9014_ ;
	wire _w9013_ ;
	wire _w9012_ ;
	wire _w9011_ ;
	wire _w9010_ ;
	wire _w9009_ ;
	wire _w9008_ ;
	wire _w9007_ ;
	wire _w9006_ ;
	wire _w9005_ ;
	wire _w9004_ ;
	wire _w9003_ ;
	wire _w9002_ ;
	wire _w9001_ ;
	wire _w9000_ ;
	wire _w8999_ ;
	wire _w8998_ ;
	wire _w8997_ ;
	wire _w8996_ ;
	wire _w8995_ ;
	wire _w8994_ ;
	wire _w8993_ ;
	wire _w8992_ ;
	wire _w8991_ ;
	wire _w8990_ ;
	wire _w8989_ ;
	wire _w8988_ ;
	wire _w8987_ ;
	wire _w8986_ ;
	wire _w8985_ ;
	wire _w8984_ ;
	wire _w8983_ ;
	wire _w8982_ ;
	wire _w8981_ ;
	wire _w8980_ ;
	wire _w8979_ ;
	wire _w8978_ ;
	wire _w8977_ ;
	wire _w8976_ ;
	wire _w8975_ ;
	wire _w8974_ ;
	wire _w8973_ ;
	wire _w8972_ ;
	wire _w8971_ ;
	wire _w8970_ ;
	wire _w8969_ ;
	wire _w8968_ ;
	wire _w8967_ ;
	wire _w8966_ ;
	wire _w8965_ ;
	wire _w8964_ ;
	wire _w8963_ ;
	wire _w8962_ ;
	wire _w8961_ ;
	wire _w8960_ ;
	wire _w8959_ ;
	wire _w8958_ ;
	wire _w8957_ ;
	wire _w8956_ ;
	wire _w8955_ ;
	wire _w8954_ ;
	wire _w8953_ ;
	wire _w8952_ ;
	wire _w8951_ ;
	wire _w8950_ ;
	wire _w8949_ ;
	wire _w8948_ ;
	wire _w8947_ ;
	wire _w8946_ ;
	wire _w8945_ ;
	wire _w8944_ ;
	wire _w8943_ ;
	wire _w8942_ ;
	wire _w8941_ ;
	wire _w8940_ ;
	wire _w8939_ ;
	wire _w8938_ ;
	wire _w8937_ ;
	wire _w8936_ ;
	wire _w8935_ ;
	wire _w8934_ ;
	wire _w8933_ ;
	wire _w8932_ ;
	wire _w8931_ ;
	wire _w8930_ ;
	wire _w8929_ ;
	wire _w8928_ ;
	wire _w8927_ ;
	wire _w8926_ ;
	wire _w8925_ ;
	wire _w8924_ ;
	wire _w8923_ ;
	wire _w8922_ ;
	wire _w8921_ ;
	wire _w8920_ ;
	wire _w8919_ ;
	wire _w8918_ ;
	wire _w8917_ ;
	wire _w8916_ ;
	wire _w8915_ ;
	wire _w8914_ ;
	wire _w8913_ ;
	wire _w8912_ ;
	wire _w8911_ ;
	wire _w8910_ ;
	wire _w8909_ ;
	wire _w8908_ ;
	wire _w8907_ ;
	wire _w8906_ ;
	wire _w8905_ ;
	wire _w8904_ ;
	wire _w8903_ ;
	wire _w8902_ ;
	wire _w8901_ ;
	wire _w8900_ ;
	wire _w8899_ ;
	wire _w8898_ ;
	wire _w8897_ ;
	wire _w8896_ ;
	wire _w8895_ ;
	wire _w8894_ ;
	wire _w8893_ ;
	wire _w8892_ ;
	wire _w8891_ ;
	wire _w8890_ ;
	wire _w8889_ ;
	wire _w8888_ ;
	wire _w8887_ ;
	wire _w8886_ ;
	wire _w8885_ ;
	wire _w8884_ ;
	wire _w8883_ ;
	wire _w8882_ ;
	wire _w8881_ ;
	wire _w8880_ ;
	wire _w8879_ ;
	wire _w8878_ ;
	wire _w8877_ ;
	wire _w8876_ ;
	wire _w8875_ ;
	wire _w8874_ ;
	wire _w8873_ ;
	wire _w8872_ ;
	wire _w8871_ ;
	wire _w8870_ ;
	wire _w8869_ ;
	wire _w8868_ ;
	wire _w8867_ ;
	wire _w8866_ ;
	wire _w8865_ ;
	wire _w8864_ ;
	wire _w8863_ ;
	wire _w8862_ ;
	wire _w8861_ ;
	wire _w8860_ ;
	wire _w8859_ ;
	wire _w8858_ ;
	wire _w8857_ ;
	wire _w8856_ ;
	wire _w8855_ ;
	wire _w8854_ ;
	wire _w8853_ ;
	wire _w8852_ ;
	wire _w8851_ ;
	wire _w8850_ ;
	wire _w8849_ ;
	wire _w8848_ ;
	wire _w8847_ ;
	wire _w8846_ ;
	wire _w8845_ ;
	wire _w8844_ ;
	wire _w8843_ ;
	wire _w8842_ ;
	wire _w8841_ ;
	wire _w8840_ ;
	wire _w8839_ ;
	wire _w8838_ ;
	wire _w8837_ ;
	wire _w8836_ ;
	wire _w8835_ ;
	wire _w8834_ ;
	wire _w8833_ ;
	wire _w8832_ ;
	wire _w8831_ ;
	wire _w8830_ ;
	wire _w8829_ ;
	wire _w8828_ ;
	wire _w8827_ ;
	wire _w8826_ ;
	wire _w8825_ ;
	wire _w8824_ ;
	wire _w8823_ ;
	wire _w8822_ ;
	wire _w8821_ ;
	wire _w8820_ ;
	wire _w8819_ ;
	wire _w8818_ ;
	wire _w8817_ ;
	wire _w8816_ ;
	wire _w8815_ ;
	wire _w8814_ ;
	wire _w8813_ ;
	wire _w8812_ ;
	wire _w8811_ ;
	wire _w8810_ ;
	wire _w8809_ ;
	wire _w8808_ ;
	wire _w8807_ ;
	wire _w8806_ ;
	wire _w8805_ ;
	wire _w8804_ ;
	wire _w8803_ ;
	wire _w8802_ ;
	wire _w8801_ ;
	wire _w8800_ ;
	wire _w8799_ ;
	wire _w8798_ ;
	wire _w8797_ ;
	wire _w8796_ ;
	wire _w8795_ ;
	wire _w8794_ ;
	wire _w8793_ ;
	wire _w8792_ ;
	wire _w8791_ ;
	wire _w8790_ ;
	wire _w8789_ ;
	wire _w8788_ ;
	wire _w8787_ ;
	wire _w8786_ ;
	wire _w8785_ ;
	wire _w8784_ ;
	wire _w8783_ ;
	wire _w8782_ ;
	wire _w8781_ ;
	wire _w8780_ ;
	wire _w8779_ ;
	wire _w8778_ ;
	wire _w8777_ ;
	wire _w8776_ ;
	wire _w8775_ ;
	wire _w8774_ ;
	wire _w8773_ ;
	wire _w8772_ ;
	wire _w8771_ ;
	wire _w8770_ ;
	wire _w8769_ ;
	wire _w8768_ ;
	wire _w8767_ ;
	wire _w8766_ ;
	wire _w8765_ ;
	wire _w8764_ ;
	wire _w8763_ ;
	wire _w8762_ ;
	wire _w8761_ ;
	wire _w8760_ ;
	wire _w8759_ ;
	wire _w8758_ ;
	wire _w8757_ ;
	wire _w8756_ ;
	wire _w8755_ ;
	wire _w8754_ ;
	wire _w8753_ ;
	wire _w8752_ ;
	wire _w8751_ ;
	wire _w8750_ ;
	wire _w8749_ ;
	wire _w8748_ ;
	wire _w8747_ ;
	wire _w8746_ ;
	wire _w8745_ ;
	wire _w8744_ ;
	wire _w8743_ ;
	wire _w8742_ ;
	wire _w8741_ ;
	wire _w8740_ ;
	wire _w8739_ ;
	wire _w8738_ ;
	wire _w8737_ ;
	wire _w8736_ ;
	wire _w8735_ ;
	wire _w8734_ ;
	wire _w8733_ ;
	wire _w8732_ ;
	wire _w8731_ ;
	wire _w8730_ ;
	wire _w8729_ ;
	wire _w8728_ ;
	wire _w8727_ ;
	wire _w8726_ ;
	wire _w8725_ ;
	wire _w8724_ ;
	wire _w8723_ ;
	wire _w8722_ ;
	wire _w8721_ ;
	wire _w8720_ ;
	wire _w8719_ ;
	wire _w8718_ ;
	wire _w8717_ ;
	wire _w8716_ ;
	wire _w8715_ ;
	wire _w8714_ ;
	wire _w8713_ ;
	wire _w8712_ ;
	wire _w8711_ ;
	wire _w8710_ ;
	wire _w8709_ ;
	wire _w8708_ ;
	wire _w8707_ ;
	wire _w8706_ ;
	wire _w8705_ ;
	wire _w8704_ ;
	wire _w8703_ ;
	wire _w8702_ ;
	wire _w8701_ ;
	wire _w8700_ ;
	wire _w8699_ ;
	wire _w8698_ ;
	wire _w8697_ ;
	wire _w8696_ ;
	wire _w8695_ ;
	wire _w8694_ ;
	wire _w8693_ ;
	wire _w8692_ ;
	wire _w8691_ ;
	wire _w8690_ ;
	wire _w8689_ ;
	wire _w8688_ ;
	wire _w8687_ ;
	wire _w8686_ ;
	wire _w8685_ ;
	wire _w8684_ ;
	wire _w8683_ ;
	wire _w8682_ ;
	wire _w8681_ ;
	wire _w8680_ ;
	wire _w8679_ ;
	wire _w8678_ ;
	wire _w8677_ ;
	wire _w8676_ ;
	wire _w8675_ ;
	wire _w8674_ ;
	wire _w8673_ ;
	wire _w8672_ ;
	wire _w8671_ ;
	wire _w8670_ ;
	wire _w8669_ ;
	wire _w8668_ ;
	wire _w8667_ ;
	wire _w8666_ ;
	wire _w8665_ ;
	wire _w8664_ ;
	wire _w8663_ ;
	wire _w8662_ ;
	wire _w8661_ ;
	wire _w8660_ ;
	wire _w8659_ ;
	wire _w8658_ ;
	wire _w8657_ ;
	wire _w8656_ ;
	wire _w8655_ ;
	wire _w8654_ ;
	wire _w8653_ ;
	wire _w8652_ ;
	wire _w8651_ ;
	wire _w8650_ ;
	wire _w8649_ ;
	wire _w8648_ ;
	wire _w8647_ ;
	wire _w8646_ ;
	wire _w8645_ ;
	wire _w8644_ ;
	wire _w8643_ ;
	wire _w8642_ ;
	wire _w8641_ ;
	wire _w8640_ ;
	wire _w8639_ ;
	wire _w8638_ ;
	wire _w8637_ ;
	wire _w8636_ ;
	wire _w8635_ ;
	wire _w8634_ ;
	wire _w8633_ ;
	wire _w8632_ ;
	wire _w8631_ ;
	wire _w8630_ ;
	wire _w8629_ ;
	wire _w8628_ ;
	wire _w8627_ ;
	wire _w8626_ ;
	wire _w8625_ ;
	wire _w8624_ ;
	wire _w8623_ ;
	wire _w8622_ ;
	wire _w8621_ ;
	wire _w8620_ ;
	wire _w8619_ ;
	wire _w8618_ ;
	wire _w8617_ ;
	wire _w8616_ ;
	wire _w8615_ ;
	wire _w8614_ ;
	wire _w8613_ ;
	wire _w8612_ ;
	wire _w8611_ ;
	wire _w8610_ ;
	wire _w8609_ ;
	wire _w8608_ ;
	wire _w8607_ ;
	wire _w8606_ ;
	wire _w8605_ ;
	wire _w8604_ ;
	wire _w8603_ ;
	wire _w8602_ ;
	wire _w8601_ ;
	wire _w8600_ ;
	wire _w8599_ ;
	wire _w8598_ ;
	wire _w8597_ ;
	wire _w8596_ ;
	wire _w8595_ ;
	wire _w8594_ ;
	wire _w8593_ ;
	wire _w8592_ ;
	wire _w8591_ ;
	wire _w8590_ ;
	wire _w8589_ ;
	wire _w8588_ ;
	wire _w8587_ ;
	wire _w8586_ ;
	wire _w8585_ ;
	wire _w8584_ ;
	wire _w8583_ ;
	wire _w8582_ ;
	wire _w8581_ ;
	wire _w8580_ ;
	wire _w8579_ ;
	wire _w8578_ ;
	wire _w8577_ ;
	wire _w8576_ ;
	wire _w8575_ ;
	wire _w8574_ ;
	wire _w8573_ ;
	wire _w8572_ ;
	wire _w8571_ ;
	wire _w8570_ ;
	wire _w8569_ ;
	wire _w8568_ ;
	wire _w8567_ ;
	wire _w8566_ ;
	wire _w8565_ ;
	wire _w8564_ ;
	wire _w8563_ ;
	wire _w8562_ ;
	wire _w8561_ ;
	wire _w8560_ ;
	wire _w8559_ ;
	wire _w8558_ ;
	wire _w8557_ ;
	wire _w8556_ ;
	wire _w8555_ ;
	wire _w8554_ ;
	wire _w8553_ ;
	wire _w8552_ ;
	wire _w8551_ ;
	wire _w8550_ ;
	wire _w8549_ ;
	wire _w8548_ ;
	wire _w8547_ ;
	wire _w8546_ ;
	wire _w8545_ ;
	wire _w8544_ ;
	wire _w8543_ ;
	wire _w8542_ ;
	wire _w8541_ ;
	wire _w8540_ ;
	wire _w8539_ ;
	wire _w8538_ ;
	wire _w8537_ ;
	wire _w8536_ ;
	wire _w8535_ ;
	wire _w8534_ ;
	wire _w8533_ ;
	wire _w8532_ ;
	wire _w8531_ ;
	wire _w8530_ ;
	wire _w8529_ ;
	wire _w8528_ ;
	wire _w8527_ ;
	wire _w8526_ ;
	wire _w8525_ ;
	wire _w8524_ ;
	wire _w8523_ ;
	wire _w8522_ ;
	wire _w8521_ ;
	wire _w8520_ ;
	wire _w8519_ ;
	wire _w8518_ ;
	wire _w8517_ ;
	wire _w8516_ ;
	wire _w8515_ ;
	wire _w8514_ ;
	wire _w8513_ ;
	wire _w8512_ ;
	wire _w8511_ ;
	wire _w8510_ ;
	wire _w8509_ ;
	wire _w8508_ ;
	wire _w8507_ ;
	wire _w8506_ ;
	wire _w8505_ ;
	wire _w8504_ ;
	wire _w8503_ ;
	wire _w8502_ ;
	wire _w8501_ ;
	wire _w8500_ ;
	wire _w8499_ ;
	wire _w8498_ ;
	wire _w8497_ ;
	wire _w8496_ ;
	wire _w8495_ ;
	wire _w8494_ ;
	wire _w8493_ ;
	wire _w8492_ ;
	wire _w8491_ ;
	wire _w8490_ ;
	wire _w8489_ ;
	wire _w8488_ ;
	wire _w8487_ ;
	wire _w8486_ ;
	wire _w8485_ ;
	wire _w8484_ ;
	wire _w8483_ ;
	wire _w8482_ ;
	wire _w8481_ ;
	wire _w8480_ ;
	wire _w8479_ ;
	wire _w8478_ ;
	wire _w8477_ ;
	wire _w8476_ ;
	wire _w8475_ ;
	wire _w8474_ ;
	wire _w8473_ ;
	wire _w8472_ ;
	wire _w8471_ ;
	wire _w8470_ ;
	wire _w8469_ ;
	wire _w8468_ ;
	wire _w8467_ ;
	wire _w8466_ ;
	wire _w8465_ ;
	wire _w8464_ ;
	wire _w8463_ ;
	wire _w8462_ ;
	wire _w8461_ ;
	wire _w8460_ ;
	wire _w8459_ ;
	wire _w8458_ ;
	wire _w8457_ ;
	wire _w8456_ ;
	wire _w8455_ ;
	wire _w8454_ ;
	wire _w8453_ ;
	wire _w8452_ ;
	wire _w8451_ ;
	wire _w8450_ ;
	wire _w8449_ ;
	wire _w8448_ ;
	wire _w8447_ ;
	wire _w8446_ ;
	wire _w8445_ ;
	wire _w8444_ ;
	wire _w8443_ ;
	wire _w8442_ ;
	wire _w8441_ ;
	wire _w8440_ ;
	wire _w8439_ ;
	wire _w8438_ ;
	wire _w8437_ ;
	wire _w8436_ ;
	wire _w8435_ ;
	wire _w8434_ ;
	wire _w8433_ ;
	wire _w8432_ ;
	wire _w8431_ ;
	wire _w8430_ ;
	wire _w8429_ ;
	wire _w8428_ ;
	wire _w8427_ ;
	wire _w8426_ ;
	wire _w8425_ ;
	wire _w8424_ ;
	wire _w8423_ ;
	wire _w8422_ ;
	wire _w8421_ ;
	wire _w8420_ ;
	wire _w8419_ ;
	wire _w8418_ ;
	wire _w8417_ ;
	wire _w8416_ ;
	wire _w8415_ ;
	wire _w8414_ ;
	wire _w8413_ ;
	wire _w8412_ ;
	wire _w8411_ ;
	wire _w8410_ ;
	wire _w8409_ ;
	wire _w8408_ ;
	wire _w8407_ ;
	wire _w8406_ ;
	wire _w8405_ ;
	wire _w8404_ ;
	wire _w8403_ ;
	wire _w8402_ ;
	wire _w8401_ ;
	wire _w8400_ ;
	wire _w8399_ ;
	wire _w8398_ ;
	wire _w8397_ ;
	wire _w8396_ ;
	wire _w8395_ ;
	wire _w8394_ ;
	wire _w8393_ ;
	wire _w8392_ ;
	wire _w8391_ ;
	wire _w8390_ ;
	wire _w8389_ ;
	wire _w8388_ ;
	wire _w8387_ ;
	wire _w8386_ ;
	wire _w8385_ ;
	wire _w8384_ ;
	wire _w8383_ ;
	wire _w8382_ ;
	wire _w8381_ ;
	wire _w8380_ ;
	wire _w8379_ ;
	wire _w8378_ ;
	wire _w8377_ ;
	wire _w8376_ ;
	wire _w8375_ ;
	wire _w8374_ ;
	wire _w8373_ ;
	wire _w8372_ ;
	wire _w8371_ ;
	wire _w8370_ ;
	wire _w8369_ ;
	wire _w8368_ ;
	wire _w8367_ ;
	wire _w8366_ ;
	wire _w8365_ ;
	wire _w8364_ ;
	wire _w8363_ ;
	wire _w8362_ ;
	wire _w8361_ ;
	wire _w8360_ ;
	wire _w8359_ ;
	wire _w8358_ ;
	wire _w8357_ ;
	wire _w8356_ ;
	wire _w8355_ ;
	wire _w8354_ ;
	wire _w8353_ ;
	wire _w8352_ ;
	wire _w8351_ ;
	wire _w8350_ ;
	wire _w8349_ ;
	wire _w8348_ ;
	wire _w8347_ ;
	wire _w8346_ ;
	wire _w8345_ ;
	wire _w8344_ ;
	wire _w8343_ ;
	wire _w8342_ ;
	wire _w8341_ ;
	wire _w8340_ ;
	wire _w8339_ ;
	wire _w8338_ ;
	wire _w8337_ ;
	wire _w8336_ ;
	wire _w8335_ ;
	wire _w8334_ ;
	wire _w8333_ ;
	wire _w8332_ ;
	wire _w8331_ ;
	wire _w8330_ ;
	wire _w8329_ ;
	wire _w8328_ ;
	wire _w8327_ ;
	wire _w8326_ ;
	wire _w8325_ ;
	wire _w8324_ ;
	wire _w8323_ ;
	wire _w8322_ ;
	wire _w8321_ ;
	wire _w8320_ ;
	wire _w8319_ ;
	wire _w8318_ ;
	wire _w8317_ ;
	wire _w8316_ ;
	wire _w8315_ ;
	wire _w8314_ ;
	wire _w8313_ ;
	wire _w8312_ ;
	wire _w8311_ ;
	wire _w8310_ ;
	wire _w8309_ ;
	wire _w8308_ ;
	wire _w8307_ ;
	wire _w8306_ ;
	wire _w8305_ ;
	wire _w8304_ ;
	wire _w8303_ ;
	wire _w8302_ ;
	wire _w8301_ ;
	wire _w8300_ ;
	wire _w8299_ ;
	wire _w8298_ ;
	wire _w8297_ ;
	wire _w8296_ ;
	wire _w8295_ ;
	wire _w8294_ ;
	wire _w8293_ ;
	wire _w8292_ ;
	wire _w8291_ ;
	wire _w8290_ ;
	wire _w8289_ ;
	wire _w8288_ ;
	wire _w8287_ ;
	wire _w8286_ ;
	wire _w8285_ ;
	wire _w8284_ ;
	wire _w8283_ ;
	wire _w8282_ ;
	wire _w8281_ ;
	wire _w8280_ ;
	wire _w8279_ ;
	wire _w8278_ ;
	wire _w8277_ ;
	wire _w8276_ ;
	wire _w8275_ ;
	wire _w8274_ ;
	wire _w8273_ ;
	wire _w8272_ ;
	wire _w8271_ ;
	wire _w8270_ ;
	wire _w8269_ ;
	wire _w8268_ ;
	wire _w8267_ ;
	wire _w8266_ ;
	wire _w8265_ ;
	wire _w8264_ ;
	wire _w8263_ ;
	wire _w8262_ ;
	wire _w8261_ ;
	wire _w8260_ ;
	wire _w8259_ ;
	wire _w8258_ ;
	wire _w8257_ ;
	wire _w8256_ ;
	wire _w8255_ ;
	wire _w8254_ ;
	wire _w8253_ ;
	wire _w8252_ ;
	wire _w8251_ ;
	wire _w8250_ ;
	wire _w8249_ ;
	wire _w8248_ ;
	wire _w8247_ ;
	wire _w8246_ ;
	wire _w8245_ ;
	wire _w8244_ ;
	wire _w8243_ ;
	wire _w8242_ ;
	wire _w8241_ ;
	wire _w8240_ ;
	wire _w8239_ ;
	wire _w8238_ ;
	wire _w8237_ ;
	wire _w8236_ ;
	wire _w8235_ ;
	wire _w8234_ ;
	wire _w8233_ ;
	wire _w8232_ ;
	wire _w8231_ ;
	wire _w8230_ ;
	wire _w8229_ ;
	wire _w8228_ ;
	wire _w8227_ ;
	wire _w8226_ ;
	wire _w8225_ ;
	wire _w8224_ ;
	wire _w8223_ ;
	wire _w8222_ ;
	wire _w8221_ ;
	wire _w8220_ ;
	wire _w8219_ ;
	wire _w8218_ ;
	wire _w8217_ ;
	wire _w8216_ ;
	wire _w8215_ ;
	wire _w8214_ ;
	wire _w8213_ ;
	wire _w8212_ ;
	wire _w8211_ ;
	wire _w8210_ ;
	wire _w8209_ ;
	wire _w8208_ ;
	wire _w8207_ ;
	wire _w8206_ ;
	wire _w8205_ ;
	wire _w8204_ ;
	wire _w8203_ ;
	wire _w8202_ ;
	wire _w8201_ ;
	wire _w8200_ ;
	wire _w8199_ ;
	wire _w8198_ ;
	wire _w8197_ ;
	wire _w8196_ ;
	wire _w8195_ ;
	wire _w8194_ ;
	wire _w8193_ ;
	wire _w8192_ ;
	wire _w8191_ ;
	wire _w8190_ ;
	wire _w8189_ ;
	wire _w8188_ ;
	wire _w8187_ ;
	wire _w8186_ ;
	wire _w8185_ ;
	wire _w8184_ ;
	wire _w8183_ ;
	wire _w8182_ ;
	wire _w8181_ ;
	wire _w8180_ ;
	wire _w8179_ ;
	wire _w8178_ ;
	wire _w8177_ ;
	wire _w8176_ ;
	wire _w8175_ ;
	wire _w8174_ ;
	wire _w8173_ ;
	wire _w8172_ ;
	wire _w8171_ ;
	wire _w8170_ ;
	wire _w8169_ ;
	wire _w8168_ ;
	wire _w8167_ ;
	wire _w8166_ ;
	wire _w8165_ ;
	wire _w8164_ ;
	wire _w8163_ ;
	wire _w8162_ ;
	wire _w8161_ ;
	wire _w8160_ ;
	wire _w8159_ ;
	wire _w8158_ ;
	wire _w8157_ ;
	wire _w8156_ ;
	wire _w8155_ ;
	wire _w8154_ ;
	wire _w8153_ ;
	wire _w8152_ ;
	wire _w8151_ ;
	wire _w8150_ ;
	wire _w8149_ ;
	wire _w8148_ ;
	wire _w8147_ ;
	wire _w8146_ ;
	wire _w8145_ ;
	wire _w8144_ ;
	wire _w8143_ ;
	wire _w8142_ ;
	wire _w8141_ ;
	wire _w8140_ ;
	wire _w8139_ ;
	wire _w8138_ ;
	wire _w8137_ ;
	wire _w8136_ ;
	wire _w8135_ ;
	wire _w8134_ ;
	wire _w8133_ ;
	wire _w8132_ ;
	wire _w8131_ ;
	wire _w8130_ ;
	wire _w8129_ ;
	wire _w8128_ ;
	wire _w8127_ ;
	wire _w8126_ ;
	wire _w8125_ ;
	wire _w8124_ ;
	wire _w8123_ ;
	wire _w8122_ ;
	wire _w8121_ ;
	wire _w8120_ ;
	wire _w8119_ ;
	wire _w8118_ ;
	wire _w8117_ ;
	wire _w8116_ ;
	wire _w8115_ ;
	wire _w8114_ ;
	wire _w8113_ ;
	wire _w8112_ ;
	wire _w8111_ ;
	wire _w8110_ ;
	wire _w8109_ ;
	wire _w8108_ ;
	wire _w8107_ ;
	wire _w8106_ ;
	wire _w8105_ ;
	wire _w8104_ ;
	wire _w8103_ ;
	wire _w8102_ ;
	wire _w8101_ ;
	wire _w8100_ ;
	wire _w8099_ ;
	wire _w8098_ ;
	wire _w8097_ ;
	wire _w8096_ ;
	wire _w8095_ ;
	wire _w8094_ ;
	wire _w8093_ ;
	wire _w8092_ ;
	wire _w8091_ ;
	wire _w8090_ ;
	wire _w8089_ ;
	wire _w8088_ ;
	wire _w8087_ ;
	wire _w8086_ ;
	wire _w8085_ ;
	wire _w8084_ ;
	wire _w8083_ ;
	wire _w8082_ ;
	wire _w8081_ ;
	wire _w8080_ ;
	wire _w8079_ ;
	wire _w8078_ ;
	wire _w8077_ ;
	wire _w8076_ ;
	wire _w8075_ ;
	wire _w8074_ ;
	wire _w8073_ ;
	wire _w8072_ ;
	wire _w8071_ ;
	wire _w8070_ ;
	wire _w8069_ ;
	wire _w8068_ ;
	wire _w8067_ ;
	wire _w8066_ ;
	wire _w8065_ ;
	wire _w8064_ ;
	wire _w8063_ ;
	wire _w8062_ ;
	wire _w8061_ ;
	wire _w8060_ ;
	wire _w8059_ ;
	wire _w8058_ ;
	wire _w8057_ ;
	wire _w8056_ ;
	wire _w8055_ ;
	wire _w8054_ ;
	wire _w8053_ ;
	wire _w8052_ ;
	wire _w8051_ ;
	wire _w8050_ ;
	wire _w8049_ ;
	wire _w8048_ ;
	wire _w8047_ ;
	wire _w8046_ ;
	wire _w8045_ ;
	wire _w8044_ ;
	wire _w8043_ ;
	wire _w8042_ ;
	wire _w8041_ ;
	wire _w8040_ ;
	wire _w8039_ ;
	wire _w8038_ ;
	wire _w8037_ ;
	wire _w8036_ ;
	wire _w8035_ ;
	wire _w8034_ ;
	wire _w8033_ ;
	wire _w8032_ ;
	wire _w8031_ ;
	wire _w8030_ ;
	wire _w8029_ ;
	wire _w8028_ ;
	wire _w8027_ ;
	wire _w8026_ ;
	wire _w8025_ ;
	wire _w8024_ ;
	wire _w8023_ ;
	wire _w8022_ ;
	wire _w8021_ ;
	wire _w8020_ ;
	wire _w8019_ ;
	wire _w8018_ ;
	wire _w8017_ ;
	wire _w8016_ ;
	wire _w8015_ ;
	wire _w8014_ ;
	wire _w8013_ ;
	wire _w8012_ ;
	wire _w8011_ ;
	wire _w8010_ ;
	wire _w8009_ ;
	wire _w8008_ ;
	wire _w8007_ ;
	wire _w8006_ ;
	wire _w8005_ ;
	wire _w8004_ ;
	wire _w8003_ ;
	wire _w8002_ ;
	wire _w8001_ ;
	wire _w8000_ ;
	wire _w7999_ ;
	wire _w7998_ ;
	wire _w7997_ ;
	wire _w7996_ ;
	wire _w7995_ ;
	wire _w7994_ ;
	wire _w7993_ ;
	wire _w7992_ ;
	wire _w7991_ ;
	wire _w7990_ ;
	wire _w7989_ ;
	wire _w7988_ ;
	wire _w7987_ ;
	wire _w7986_ ;
	wire _w7985_ ;
	wire _w7984_ ;
	wire _w7983_ ;
	wire _w7982_ ;
	wire _w7981_ ;
	wire _w7980_ ;
	wire _w7979_ ;
	wire _w7978_ ;
	wire _w7977_ ;
	wire _w7976_ ;
	wire _w7975_ ;
	wire _w7974_ ;
	wire _w7973_ ;
	wire _w7972_ ;
	wire _w7971_ ;
	wire _w7970_ ;
	wire _w7969_ ;
	wire _w7968_ ;
	wire _w7967_ ;
	wire _w7966_ ;
	wire _w7965_ ;
	wire _w7964_ ;
	wire _w7963_ ;
	wire _w7962_ ;
	wire _w7961_ ;
	wire _w7960_ ;
	wire _w7959_ ;
	wire _w7958_ ;
	wire _w7957_ ;
	wire _w7956_ ;
	wire _w7955_ ;
	wire _w7954_ ;
	wire _w7953_ ;
	wire _w7952_ ;
	wire _w7951_ ;
	wire _w7950_ ;
	wire _w7949_ ;
	wire _w7948_ ;
	wire _w7947_ ;
	wire _w7946_ ;
	wire _w7945_ ;
	wire _w7944_ ;
	wire _w7943_ ;
	wire _w7942_ ;
	wire _w7941_ ;
	wire _w7940_ ;
	wire _w7939_ ;
	wire _w7938_ ;
	wire _w7937_ ;
	wire _w7936_ ;
	wire _w7935_ ;
	wire _w7934_ ;
	wire _w7933_ ;
	wire _w7932_ ;
	wire _w7931_ ;
	wire _w7930_ ;
	wire _w7929_ ;
	wire _w7928_ ;
	wire _w7927_ ;
	wire _w7926_ ;
	wire _w7925_ ;
	wire _w7924_ ;
	wire _w7923_ ;
	wire _w7922_ ;
	wire _w7921_ ;
	wire _w7920_ ;
	wire _w7919_ ;
	wire _w7918_ ;
	wire _w7917_ ;
	wire _w7916_ ;
	wire _w7915_ ;
	wire _w7914_ ;
	wire _w7913_ ;
	wire _w7912_ ;
	wire _w7911_ ;
	wire _w7910_ ;
	wire _w7909_ ;
	wire _w7908_ ;
	wire _w7907_ ;
	wire _w7906_ ;
	wire _w7905_ ;
	wire _w7904_ ;
	wire _w7903_ ;
	wire _w7902_ ;
	wire _w7901_ ;
	wire _w7900_ ;
	wire _w7899_ ;
	wire _w7898_ ;
	wire _w7897_ ;
	wire _w7896_ ;
	wire _w7895_ ;
	wire _w7894_ ;
	wire _w7893_ ;
	wire _w7892_ ;
	wire _w7891_ ;
	wire _w7890_ ;
	wire _w7889_ ;
	wire _w7888_ ;
	wire _w7887_ ;
	wire _w7886_ ;
	wire _w7885_ ;
	wire _w7884_ ;
	wire _w7883_ ;
	wire _w7882_ ;
	wire _w7881_ ;
	wire _w7880_ ;
	wire _w7879_ ;
	wire _w7878_ ;
	wire _w7877_ ;
	wire _w7876_ ;
	wire _w7875_ ;
	wire _w7874_ ;
	wire _w7873_ ;
	wire _w7872_ ;
	wire _w7871_ ;
	wire _w7870_ ;
	wire _w7869_ ;
	wire _w7868_ ;
	wire _w7867_ ;
	wire _w7866_ ;
	wire _w7865_ ;
	wire _w7864_ ;
	wire _w7863_ ;
	wire _w7862_ ;
	wire _w7861_ ;
	wire _w7860_ ;
	wire _w7859_ ;
	wire _w7858_ ;
	wire _w7857_ ;
	wire _w7856_ ;
	wire _w7855_ ;
	wire _w7854_ ;
	wire _w7853_ ;
	wire _w7852_ ;
	wire _w7851_ ;
	wire _w7850_ ;
	wire _w7849_ ;
	wire _w7848_ ;
	wire _w7847_ ;
	wire _w7846_ ;
	wire _w7845_ ;
	wire _w7844_ ;
	wire _w7843_ ;
	wire _w7842_ ;
	wire _w7841_ ;
	wire _w7840_ ;
	wire _w7839_ ;
	wire _w7838_ ;
	wire _w7837_ ;
	wire _w7836_ ;
	wire _w7835_ ;
	wire _w7834_ ;
	wire _w7833_ ;
	wire _w7832_ ;
	wire _w7831_ ;
	wire _w7830_ ;
	wire _w7829_ ;
	wire _w7828_ ;
	wire _w7827_ ;
	wire _w7826_ ;
	wire _w7825_ ;
	wire _w7824_ ;
	wire _w7823_ ;
	wire _w7822_ ;
	wire _w7821_ ;
	wire _w7820_ ;
	wire _w7819_ ;
	wire _w7818_ ;
	wire _w7817_ ;
	wire _w7816_ ;
	wire _w7815_ ;
	wire _w7814_ ;
	wire _w7813_ ;
	wire _w7812_ ;
	wire _w7811_ ;
	wire _w7810_ ;
	wire _w7809_ ;
	wire _w7808_ ;
	wire _w7807_ ;
	wire _w7806_ ;
	wire _w7805_ ;
	wire _w7804_ ;
	wire _w7803_ ;
	wire _w7802_ ;
	wire _w7801_ ;
	wire _w7800_ ;
	wire _w7799_ ;
	wire _w7798_ ;
	wire _w7797_ ;
	wire _w7796_ ;
	wire _w7795_ ;
	wire _w7794_ ;
	wire _w7793_ ;
	wire _w7792_ ;
	wire _w7791_ ;
	wire _w7790_ ;
	wire _w7789_ ;
	wire _w7788_ ;
	wire _w7787_ ;
	wire _w7786_ ;
	wire _w7785_ ;
	wire _w7784_ ;
	wire _w7783_ ;
	wire _w7782_ ;
	wire _w7781_ ;
	wire _w7780_ ;
	wire _w7779_ ;
	wire _w7778_ ;
	wire _w7777_ ;
	wire _w7776_ ;
	wire _w7775_ ;
	wire _w7774_ ;
	wire _w7773_ ;
	wire _w7772_ ;
	wire _w7771_ ;
	wire _w7770_ ;
	wire _w7769_ ;
	wire _w7768_ ;
	wire _w7767_ ;
	wire _w7766_ ;
	wire _w7765_ ;
	wire _w7764_ ;
	wire _w7763_ ;
	wire _w7762_ ;
	wire _w7761_ ;
	wire _w7760_ ;
	wire _w7759_ ;
	wire _w7758_ ;
	wire _w7757_ ;
	wire _w7756_ ;
	wire _w7755_ ;
	wire _w7754_ ;
	wire _w7753_ ;
	wire _w7752_ ;
	wire _w7751_ ;
	wire _w7750_ ;
	wire _w7749_ ;
	wire _w7748_ ;
	wire _w7747_ ;
	wire _w7746_ ;
	wire _w7745_ ;
	wire _w7744_ ;
	wire _w7743_ ;
	wire _w7742_ ;
	wire _w7741_ ;
	wire _w7740_ ;
	wire _w7739_ ;
	wire _w7738_ ;
	wire _w7737_ ;
	wire _w7736_ ;
	wire _w7735_ ;
	wire _w7734_ ;
	wire _w7733_ ;
	wire _w7732_ ;
	wire _w7731_ ;
	wire _w7730_ ;
	wire _w7729_ ;
	wire _w7728_ ;
	wire _w7727_ ;
	wire _w7726_ ;
	wire _w7725_ ;
	wire _w7724_ ;
	wire _w7723_ ;
	wire _w7722_ ;
	wire _w7721_ ;
	wire _w7720_ ;
	wire _w7719_ ;
	wire _w7718_ ;
	wire _w7717_ ;
	wire _w7716_ ;
	wire _w7715_ ;
	wire _w7714_ ;
	wire _w7713_ ;
	wire _w7712_ ;
	wire _w7711_ ;
	wire _w7710_ ;
	wire _w7709_ ;
	wire _w7708_ ;
	wire _w7707_ ;
	wire _w7706_ ;
	wire _w7705_ ;
	wire _w7704_ ;
	wire _w7703_ ;
	wire _w7702_ ;
	wire _w7701_ ;
	wire _w7700_ ;
	wire _w7699_ ;
	wire _w7698_ ;
	wire _w7697_ ;
	wire _w7696_ ;
	wire _w7695_ ;
	wire _w7694_ ;
	wire _w7693_ ;
	wire _w7692_ ;
	wire _w7691_ ;
	wire _w7690_ ;
	wire _w7689_ ;
	wire _w7688_ ;
	wire _w7687_ ;
	wire _w7686_ ;
	wire _w7685_ ;
	wire _w7684_ ;
	wire _w7683_ ;
	wire _w7682_ ;
	wire _w7681_ ;
	wire _w7680_ ;
	wire _w7679_ ;
	wire _w7678_ ;
	wire _w7677_ ;
	wire _w7676_ ;
	wire _w7675_ ;
	wire _w7674_ ;
	wire _w7673_ ;
	wire _w7672_ ;
	wire _w7671_ ;
	wire _w7670_ ;
	wire _w7669_ ;
	wire _w7668_ ;
	wire _w7667_ ;
	wire _w7666_ ;
	wire _w7665_ ;
	wire _w7664_ ;
	wire _w7663_ ;
	wire _w7662_ ;
	wire _w7661_ ;
	wire _w7660_ ;
	wire _w7659_ ;
	wire _w7658_ ;
	wire _w7657_ ;
	wire _w7656_ ;
	wire _w7655_ ;
	wire _w7654_ ;
	wire _w7653_ ;
	wire _w7652_ ;
	wire _w7651_ ;
	wire _w7650_ ;
	wire _w7649_ ;
	wire _w7648_ ;
	wire _w7647_ ;
	wire _w7646_ ;
	wire _w7645_ ;
	wire _w7644_ ;
	wire _w7643_ ;
	wire _w7642_ ;
	wire _w7641_ ;
	wire _w7640_ ;
	wire _w7639_ ;
	wire _w7638_ ;
	wire _w7637_ ;
	wire _w7636_ ;
	wire _w7635_ ;
	wire _w7634_ ;
	wire _w7633_ ;
	wire _w7632_ ;
	wire _w7631_ ;
	wire _w7630_ ;
	wire _w7629_ ;
	wire _w7628_ ;
	wire _w7627_ ;
	wire _w7626_ ;
	wire _w7625_ ;
	wire _w7624_ ;
	wire _w7623_ ;
	wire _w7622_ ;
	wire _w7621_ ;
	wire _w7620_ ;
	wire _w7619_ ;
	wire _w7618_ ;
	wire _w7617_ ;
	wire _w7616_ ;
	wire _w7615_ ;
	wire _w7614_ ;
	wire _w7613_ ;
	wire _w7612_ ;
	wire _w7611_ ;
	wire _w7610_ ;
	wire _w7609_ ;
	wire _w7608_ ;
	wire _w7607_ ;
	wire _w7606_ ;
	wire _w7605_ ;
	wire _w7604_ ;
	wire _w7603_ ;
	wire _w7602_ ;
	wire _w7601_ ;
	wire _w7600_ ;
	wire _w7599_ ;
	wire _w7598_ ;
	wire _w7597_ ;
	wire _w7596_ ;
	wire _w7595_ ;
	wire _w7594_ ;
	wire _w7593_ ;
	wire _w7592_ ;
	wire _w7591_ ;
	wire _w7590_ ;
	wire _w7589_ ;
	wire _w7588_ ;
	wire _w7587_ ;
	wire _w7586_ ;
	wire _w7585_ ;
	wire _w7584_ ;
	wire _w7583_ ;
	wire _w7582_ ;
	wire _w7581_ ;
	wire _w7580_ ;
	wire _w7579_ ;
	wire _w7578_ ;
	wire _w7577_ ;
	wire _w7576_ ;
	wire _w7575_ ;
	wire _w7574_ ;
	wire _w7573_ ;
	wire _w7572_ ;
	wire _w7571_ ;
	wire _w7570_ ;
	wire _w7569_ ;
	wire _w7568_ ;
	wire _w7567_ ;
	wire _w7566_ ;
	wire _w7565_ ;
	wire _w7564_ ;
	wire _w7563_ ;
	wire _w7562_ ;
	wire _w7561_ ;
	wire _w7560_ ;
	wire _w7559_ ;
	wire _w7558_ ;
	wire _w7557_ ;
	wire _w7556_ ;
	wire _w7555_ ;
	wire _w7554_ ;
	wire _w7553_ ;
	wire _w7552_ ;
	wire _w7551_ ;
	wire _w7550_ ;
	wire _w7549_ ;
	wire _w7548_ ;
	wire _w7547_ ;
	wire _w7546_ ;
	wire _w7545_ ;
	wire _w7544_ ;
	wire _w7543_ ;
	wire _w7542_ ;
	wire _w7541_ ;
	wire _w7540_ ;
	wire _w7539_ ;
	wire _w7538_ ;
	wire _w7537_ ;
	wire _w7536_ ;
	wire _w7535_ ;
	wire _w7534_ ;
	wire _w7533_ ;
	wire _w7532_ ;
	wire _w7531_ ;
	wire _w7530_ ;
	wire _w7529_ ;
	wire _w7528_ ;
	wire _w7527_ ;
	wire _w7526_ ;
	wire _w7525_ ;
	wire _w7524_ ;
	wire _w7523_ ;
	wire _w7522_ ;
	wire _w7521_ ;
	wire _w7520_ ;
	wire _w7519_ ;
	wire _w7518_ ;
	wire _w7517_ ;
	wire _w7516_ ;
	wire _w7515_ ;
	wire _w7514_ ;
	wire _w7513_ ;
	wire _w7512_ ;
	wire _w7511_ ;
	wire _w7510_ ;
	wire _w7509_ ;
	wire _w7508_ ;
	wire _w7507_ ;
	wire _w7506_ ;
	wire _w7505_ ;
	wire _w7504_ ;
	wire _w7503_ ;
	wire _w7502_ ;
	wire _w7501_ ;
	wire _w7500_ ;
	wire _w7499_ ;
	wire _w7498_ ;
	wire _w7497_ ;
	wire _w7496_ ;
	wire _w7495_ ;
	wire _w7494_ ;
	wire _w7493_ ;
	wire _w7492_ ;
	wire _w7491_ ;
	wire _w7490_ ;
	wire _w7489_ ;
	wire _w7488_ ;
	wire _w7487_ ;
	wire _w7486_ ;
	wire _w7485_ ;
	wire _w7484_ ;
	wire _w7483_ ;
	wire _w7482_ ;
	wire _w7481_ ;
	wire _w7480_ ;
	wire _w7479_ ;
	wire _w7478_ ;
	wire _w7477_ ;
	wire _w7476_ ;
	wire _w7475_ ;
	wire _w7474_ ;
	wire _w7473_ ;
	wire _w7472_ ;
	wire _w7471_ ;
	wire _w7470_ ;
	wire _w7469_ ;
	wire _w7468_ ;
	wire _w7467_ ;
	wire _w7466_ ;
	wire _w7465_ ;
	wire _w7464_ ;
	wire _w7463_ ;
	wire _w7462_ ;
	wire _w7461_ ;
	wire _w7460_ ;
	wire _w7459_ ;
	wire _w7458_ ;
	wire _w7457_ ;
	wire _w7456_ ;
	wire _w7455_ ;
	wire _w7454_ ;
	wire _w7453_ ;
	wire _w7452_ ;
	wire _w7451_ ;
	wire _w7450_ ;
	wire _w7449_ ;
	wire _w7448_ ;
	wire _w7447_ ;
	wire _w7446_ ;
	wire _w7445_ ;
	wire _w7444_ ;
	wire _w7443_ ;
	wire _w7442_ ;
	wire _w7441_ ;
	wire _w7440_ ;
	wire _w7439_ ;
	wire _w7438_ ;
	wire _w7437_ ;
	wire _w7436_ ;
	wire _w7435_ ;
	wire _w7434_ ;
	wire _w7433_ ;
	wire _w7432_ ;
	wire _w7431_ ;
	wire _w7430_ ;
	wire _w7429_ ;
	wire _w7428_ ;
	wire _w7427_ ;
	wire _w7426_ ;
	wire _w7425_ ;
	wire _w7424_ ;
	wire _w7423_ ;
	wire _w7422_ ;
	wire _w7421_ ;
	wire _w7420_ ;
	wire _w7419_ ;
	wire _w7418_ ;
	wire _w7417_ ;
	wire _w7416_ ;
	wire _w7415_ ;
	wire _w7414_ ;
	wire _w7413_ ;
	wire _w7412_ ;
	wire _w7411_ ;
	wire _w7410_ ;
	wire _w7409_ ;
	wire _w7408_ ;
	wire _w7407_ ;
	wire _w7406_ ;
	wire _w7405_ ;
	wire _w7404_ ;
	wire _w7403_ ;
	wire _w7402_ ;
	wire _w7401_ ;
	wire _w7400_ ;
	wire _w7399_ ;
	wire _w7398_ ;
	wire _w7397_ ;
	wire _w7396_ ;
	wire _w7395_ ;
	wire _w7394_ ;
	wire _w7393_ ;
	wire _w7392_ ;
	wire _w7391_ ;
	wire _w7390_ ;
	wire _w7389_ ;
	wire _w7388_ ;
	wire _w7387_ ;
	wire _w7386_ ;
	wire _w7385_ ;
	wire _w7384_ ;
	wire _w7383_ ;
	wire _w7382_ ;
	wire _w7381_ ;
	wire _w7380_ ;
	wire _w7379_ ;
	wire _w7378_ ;
	wire _w7377_ ;
	wire _w7376_ ;
	wire _w7375_ ;
	wire _w7374_ ;
	wire _w7373_ ;
	wire _w7372_ ;
	wire _w7371_ ;
	wire _w7370_ ;
	wire _w7369_ ;
	wire _w7368_ ;
	wire _w7367_ ;
	wire _w7366_ ;
	wire _w7365_ ;
	wire _w7364_ ;
	wire _w7363_ ;
	wire _w7362_ ;
	wire _w7361_ ;
	wire _w7360_ ;
	wire _w7359_ ;
	wire _w7358_ ;
	wire _w7357_ ;
	wire _w7356_ ;
	wire _w7355_ ;
	wire _w7354_ ;
	wire _w7353_ ;
	wire _w7352_ ;
	wire _w7351_ ;
	wire _w7350_ ;
	wire _w7349_ ;
	wire _w7348_ ;
	wire _w7347_ ;
	wire _w7346_ ;
	wire _w7345_ ;
	wire _w7344_ ;
	wire _w7343_ ;
	wire _w7342_ ;
	wire _w7341_ ;
	wire _w7340_ ;
	wire _w7339_ ;
	wire _w7338_ ;
	wire _w7337_ ;
	wire _w7336_ ;
	wire _w7335_ ;
	wire _w7334_ ;
	wire _w7333_ ;
	wire _w7332_ ;
	wire _w7331_ ;
	wire _w7330_ ;
	wire _w7329_ ;
	wire _w7328_ ;
	wire _w7327_ ;
	wire _w7326_ ;
	wire _w7325_ ;
	wire _w7324_ ;
	wire _w7323_ ;
	wire _w7322_ ;
	wire _w7321_ ;
	wire _w7320_ ;
	wire _w7319_ ;
	wire _w7318_ ;
	wire _w7317_ ;
	wire _w7316_ ;
	wire _w7315_ ;
	wire _w7314_ ;
	wire _w7313_ ;
	wire _w7312_ ;
	wire _w7311_ ;
	wire _w7310_ ;
	wire _w7309_ ;
	wire _w7308_ ;
	wire _w7307_ ;
	wire _w7306_ ;
	wire _w7305_ ;
	wire _w7304_ ;
	wire _w7303_ ;
	wire _w7302_ ;
	wire _w7301_ ;
	wire _w7300_ ;
	wire _w7299_ ;
	wire _w7298_ ;
	wire _w7297_ ;
	wire _w7296_ ;
	wire _w7295_ ;
	wire _w7294_ ;
	wire _w7293_ ;
	wire _w7292_ ;
	wire _w7291_ ;
	wire _w7290_ ;
	wire _w7289_ ;
	wire _w7288_ ;
	wire _w7287_ ;
	wire _w7286_ ;
	wire _w7285_ ;
	wire _w7284_ ;
	wire _w7283_ ;
	wire _w7282_ ;
	wire _w7281_ ;
	wire _w7280_ ;
	wire _w7279_ ;
	wire _w7278_ ;
	wire _w7277_ ;
	wire _w7276_ ;
	wire _w7275_ ;
	wire _w7274_ ;
	wire _w7273_ ;
	wire _w7272_ ;
	wire _w7271_ ;
	wire _w7270_ ;
	wire _w7269_ ;
	wire _w7268_ ;
	wire _w7267_ ;
	wire _w7266_ ;
	wire _w7265_ ;
	wire _w7264_ ;
	wire _w7263_ ;
	wire _w7262_ ;
	wire _w7261_ ;
	wire _w7260_ ;
	wire _w7259_ ;
	wire _w7258_ ;
	wire _w7257_ ;
	wire _w7256_ ;
	wire _w7255_ ;
	wire _w7254_ ;
	wire _w7253_ ;
	wire _w7252_ ;
	wire _w7251_ ;
	wire _w7250_ ;
	wire _w7249_ ;
	wire _w7248_ ;
	wire _w7247_ ;
	wire _w7246_ ;
	wire _w7245_ ;
	wire _w7244_ ;
	wire _w7243_ ;
	wire _w7242_ ;
	wire _w7241_ ;
	wire _w7240_ ;
	wire _w7239_ ;
	wire _w7238_ ;
	wire _w7237_ ;
	wire _w7236_ ;
	wire _w7235_ ;
	wire _w7234_ ;
	wire _w7233_ ;
	wire _w7232_ ;
	wire _w7231_ ;
	wire _w7230_ ;
	wire _w7229_ ;
	wire _w7228_ ;
	wire _w7227_ ;
	wire _w7226_ ;
	wire _w7225_ ;
	wire _w7224_ ;
	wire _w7223_ ;
	wire _w7222_ ;
	wire _w7221_ ;
	wire _w7220_ ;
	wire _w7219_ ;
	wire _w7218_ ;
	wire _w7217_ ;
	wire _w7216_ ;
	wire _w7215_ ;
	wire _w7214_ ;
	wire _w7213_ ;
	wire _w7212_ ;
	wire _w7211_ ;
	wire _w7210_ ;
	wire _w7209_ ;
	wire _w7208_ ;
	wire _w7207_ ;
	wire _w7206_ ;
	wire _w7205_ ;
	wire _w7204_ ;
	wire _w7203_ ;
	wire _w7202_ ;
	wire _w7201_ ;
	wire _w7200_ ;
	wire _w7199_ ;
	wire _w7198_ ;
	wire _w7197_ ;
	wire _w7196_ ;
	wire _w7195_ ;
	wire _w7194_ ;
	wire _w7193_ ;
	wire _w7192_ ;
	wire _w7191_ ;
	wire _w7190_ ;
	wire _w7189_ ;
	wire _w7188_ ;
	wire _w7187_ ;
	wire _w7186_ ;
	wire _w7185_ ;
	wire _w7184_ ;
	wire _w7183_ ;
	wire _w7182_ ;
	wire _w7181_ ;
	wire _w7180_ ;
	wire _w7179_ ;
	wire _w7178_ ;
	wire _w7177_ ;
	wire _w7176_ ;
	wire _w7175_ ;
	wire _w7174_ ;
	wire _w7173_ ;
	wire _w7172_ ;
	wire _w7171_ ;
	wire _w7170_ ;
	wire _w7169_ ;
	wire _w7168_ ;
	wire _w7167_ ;
	wire _w7166_ ;
	wire _w7165_ ;
	wire _w7164_ ;
	wire _w7163_ ;
	wire _w7162_ ;
	wire _w7161_ ;
	wire _w7160_ ;
	wire _w7159_ ;
	wire _w7158_ ;
	wire _w7157_ ;
	wire _w7156_ ;
	wire _w7155_ ;
	wire _w7154_ ;
	wire _w7153_ ;
	wire _w7152_ ;
	wire _w7151_ ;
	wire _w7150_ ;
	wire _w7149_ ;
	wire _w7148_ ;
	wire _w7147_ ;
	wire _w7146_ ;
	wire _w7145_ ;
	wire _w7144_ ;
	wire _w7143_ ;
	wire _w7142_ ;
	wire _w7141_ ;
	wire _w7140_ ;
	wire _w7139_ ;
	wire _w7138_ ;
	wire _w7137_ ;
	wire _w7136_ ;
	wire _w7135_ ;
	wire _w7134_ ;
	wire _w7133_ ;
	wire _w7132_ ;
	wire _w7131_ ;
	wire _w7130_ ;
	wire _w7129_ ;
	wire _w7128_ ;
	wire _w7127_ ;
	wire _w7126_ ;
	wire _w7125_ ;
	wire _w7124_ ;
	wire _w7123_ ;
	wire _w7122_ ;
	wire _w7121_ ;
	wire _w7120_ ;
	wire _w7119_ ;
	wire _w7118_ ;
	wire _w7117_ ;
	wire _w7116_ ;
	wire _w7115_ ;
	wire _w7114_ ;
	wire _w7113_ ;
	wire _w7112_ ;
	wire _w7111_ ;
	wire _w7110_ ;
	wire _w7109_ ;
	wire _w7108_ ;
	wire _w7107_ ;
	wire _w7106_ ;
	wire _w7105_ ;
	wire _w7104_ ;
	wire _w7103_ ;
	wire _w7102_ ;
	wire _w7101_ ;
	wire _w7100_ ;
	wire _w7099_ ;
	wire _w7098_ ;
	wire _w7097_ ;
	wire _w7096_ ;
	wire _w7095_ ;
	wire _w7094_ ;
	wire _w7093_ ;
	wire _w7092_ ;
	wire _w7091_ ;
	wire _w7090_ ;
	wire _w7089_ ;
	wire _w7088_ ;
	wire _w7087_ ;
	wire _w7086_ ;
	wire _w7085_ ;
	wire _w7084_ ;
	wire _w7083_ ;
	wire _w7082_ ;
	wire _w7081_ ;
	wire _w7080_ ;
	wire _w7079_ ;
	wire _w7078_ ;
	wire _w7077_ ;
	wire _w7076_ ;
	wire _w7075_ ;
	wire _w7074_ ;
	wire _w7073_ ;
	wire _w7072_ ;
	wire _w7071_ ;
	wire _w7070_ ;
	wire _w7069_ ;
	wire _w7068_ ;
	wire _w7067_ ;
	wire _w7066_ ;
	wire _w7065_ ;
	wire _w7064_ ;
	wire _w7063_ ;
	wire _w7062_ ;
	wire _w7061_ ;
	wire _w7060_ ;
	wire _w7059_ ;
	wire _w7058_ ;
	wire _w7057_ ;
	wire _w7056_ ;
	wire _w7055_ ;
	wire _w7054_ ;
	wire _w7053_ ;
	wire _w7052_ ;
	wire _w7051_ ;
	wire _w7050_ ;
	wire _w7049_ ;
	wire _w7048_ ;
	wire _w7047_ ;
	wire _w7046_ ;
	wire _w7045_ ;
	wire _w7044_ ;
	wire _w7043_ ;
	wire _w7042_ ;
	wire _w7041_ ;
	wire _w7040_ ;
	wire _w7039_ ;
	wire _w7038_ ;
	wire _w7037_ ;
	wire _w7036_ ;
	wire _w7035_ ;
	wire _w7034_ ;
	wire _w7033_ ;
	wire _w7032_ ;
	wire _w7031_ ;
	wire _w7030_ ;
	wire _w7029_ ;
	wire _w7028_ ;
	wire _w7027_ ;
	wire _w7026_ ;
	wire _w7025_ ;
	wire _w7024_ ;
	wire _w7023_ ;
	wire _w7022_ ;
	wire _w7021_ ;
	wire _w7020_ ;
	wire _w7019_ ;
	wire _w7018_ ;
	wire _w7017_ ;
	wire _w7016_ ;
	wire _w7015_ ;
	wire _w7014_ ;
	wire _w7013_ ;
	wire _w7012_ ;
	wire _w7011_ ;
	wire _w7010_ ;
	wire _w7009_ ;
	wire _w7008_ ;
	wire _w7007_ ;
	wire _w7006_ ;
	wire _w7005_ ;
	wire _w7004_ ;
	wire _w7003_ ;
	wire _w7002_ ;
	wire _w7001_ ;
	wire _w7000_ ;
	wire _w6999_ ;
	wire _w6998_ ;
	wire _w6997_ ;
	wire _w6996_ ;
	wire _w6995_ ;
	wire _w6994_ ;
	wire _w6993_ ;
	wire _w6992_ ;
	wire _w6991_ ;
	wire _w6990_ ;
	wire _w6989_ ;
	wire _w6988_ ;
	wire _w6987_ ;
	wire _w6986_ ;
	wire _w6985_ ;
	wire _w6984_ ;
	wire _w6983_ ;
	wire _w6982_ ;
	wire _w6981_ ;
	wire _w6980_ ;
	wire _w6979_ ;
	wire _w6978_ ;
	wire _w6977_ ;
	wire _w6976_ ;
	wire _w6975_ ;
	wire _w6974_ ;
	wire _w6973_ ;
	wire _w6972_ ;
	wire _w6971_ ;
	wire _w6970_ ;
	wire _w6969_ ;
	wire _w6968_ ;
	wire _w6967_ ;
	wire _w6966_ ;
	wire _w6965_ ;
	wire _w6964_ ;
	wire _w6963_ ;
	wire _w6962_ ;
	wire _w6961_ ;
	wire _w6960_ ;
	wire _w6959_ ;
	wire _w6958_ ;
	wire _w6957_ ;
	wire _w6956_ ;
	wire _w6955_ ;
	wire _w6954_ ;
	wire _w6953_ ;
	wire _w6952_ ;
	wire _w6951_ ;
	wire _w6950_ ;
	wire _w6949_ ;
	wire _w6948_ ;
	wire _w6947_ ;
	wire _w6946_ ;
	wire _w6945_ ;
	wire _w6944_ ;
	wire _w6943_ ;
	wire _w6942_ ;
	wire _w6941_ ;
	wire _w6940_ ;
	wire _w6939_ ;
	wire _w6938_ ;
	wire _w6937_ ;
	wire _w6936_ ;
	wire _w6935_ ;
	wire _w6934_ ;
	wire _w6933_ ;
	wire _w6932_ ;
	wire _w6931_ ;
	wire _w6930_ ;
	wire _w6929_ ;
	wire _w6928_ ;
	wire _w6927_ ;
	wire _w6926_ ;
	wire _w6925_ ;
	wire _w6924_ ;
	wire _w6923_ ;
	wire _w6922_ ;
	wire _w6921_ ;
	wire _w6920_ ;
	wire _w6919_ ;
	wire _w6918_ ;
	wire _w6917_ ;
	wire _w6916_ ;
	wire _w6915_ ;
	wire _w6914_ ;
	wire _w6913_ ;
	wire _w6912_ ;
	wire _w6911_ ;
	wire _w6910_ ;
	wire _w6909_ ;
	wire _w6908_ ;
	wire _w6907_ ;
	wire _w6906_ ;
	wire _w6905_ ;
	wire _w6904_ ;
	wire _w6903_ ;
	wire _w6902_ ;
	wire _w6901_ ;
	wire _w6900_ ;
	wire _w6899_ ;
	wire _w6898_ ;
	wire _w6897_ ;
	wire _w6896_ ;
	wire _w6895_ ;
	wire _w6894_ ;
	wire _w6893_ ;
	wire _w6892_ ;
	wire _w6891_ ;
	wire _w6890_ ;
	wire _w6889_ ;
	wire _w6888_ ;
	wire _w6887_ ;
	wire _w6886_ ;
	wire _w6885_ ;
	wire _w6884_ ;
	wire _w6883_ ;
	wire _w6882_ ;
	wire _w6881_ ;
	wire _w6880_ ;
	wire _w6879_ ;
	wire _w6878_ ;
	wire _w6877_ ;
	wire _w6876_ ;
	wire _w6875_ ;
	wire _w6874_ ;
	wire _w6873_ ;
	wire _w6872_ ;
	wire _w6871_ ;
	wire _w6870_ ;
	wire _w6869_ ;
	wire _w6868_ ;
	wire _w6867_ ;
	wire _w6866_ ;
	wire _w6865_ ;
	wire _w6864_ ;
	wire _w6863_ ;
	wire _w6862_ ;
	wire _w6861_ ;
	wire _w6860_ ;
	wire _w6859_ ;
	wire _w6858_ ;
	wire _w6857_ ;
	wire _w6856_ ;
	wire _w6855_ ;
	wire _w6854_ ;
	wire _w6853_ ;
	wire _w6852_ ;
	wire _w6851_ ;
	wire _w6850_ ;
	wire _w6849_ ;
	wire _w6848_ ;
	wire _w6847_ ;
	wire _w6846_ ;
	wire _w6845_ ;
	wire _w6844_ ;
	wire _w6843_ ;
	wire _w6842_ ;
	wire _w6841_ ;
	wire _w6840_ ;
	wire _w6839_ ;
	wire _w6838_ ;
	wire _w6837_ ;
	wire _w4106_ ;
	wire _w4105_ ;
	wire _w4104_ ;
	wire _w4103_ ;
	wire _w4102_ ;
	wire _w4101_ ;
	wire _w4100_ ;
	wire _w4099_ ;
	wire _w4098_ ;
	wire _w4097_ ;
	wire _w4096_ ;
	wire _w4095_ ;
	wire _w4094_ ;
	wire _w4093_ ;
	wire _w4092_ ;
	wire _w4091_ ;
	wire _w4090_ ;
	wire _w4089_ ;
	wire _w4088_ ;
	wire _w4087_ ;
	wire _w4086_ ;
	wire _w4085_ ;
	wire _w4084_ ;
	wire _w4083_ ;
	wire _w4082_ ;
	wire _w4081_ ;
	wire _w4080_ ;
	wire _w4079_ ;
	wire _w4078_ ;
	wire _w4077_ ;
	wire _w4076_ ;
	wire _w4075_ ;
	wire _w4074_ ;
	wire _w4073_ ;
	wire _w4072_ ;
	wire _w4071_ ;
	wire _w4070_ ;
	wire _w4069_ ;
	wire _w4068_ ;
	wire _w4067_ ;
	wire _w4066_ ;
	wire _w4065_ ;
	wire _w4064_ ;
	wire _w4063_ ;
	wire _w4062_ ;
	wire _w4061_ ;
	wire _w4060_ ;
	wire _w4059_ ;
	wire _w4058_ ;
	wire _w4057_ ;
	wire _w4056_ ;
	wire _w4055_ ;
	wire _w4054_ ;
	wire _w4053_ ;
	wire _w4052_ ;
	wire _w4051_ ;
	wire _w4050_ ;
	wire _w4049_ ;
	wire _w4048_ ;
	wire _w4047_ ;
	wire _w4046_ ;
	wire _w4045_ ;
	wire _w4044_ ;
	wire _w4043_ ;
	wire _w4042_ ;
	wire _w4041_ ;
	wire _w4040_ ;
	wire _w4039_ ;
	wire _w4038_ ;
	wire _w4037_ ;
	wire _w4036_ ;
	wire _w4035_ ;
	wire _w4034_ ;
	wire _w4033_ ;
	wire _w4032_ ;
	wire _w4031_ ;
	wire _w4030_ ;
	wire _w4029_ ;
	wire _w4028_ ;
	wire _w4027_ ;
	wire _w4026_ ;
	wire _w4025_ ;
	wire _w4024_ ;
	wire _w4023_ ;
	wire _w4022_ ;
	wire _w4021_ ;
	wire _w4020_ ;
	wire _w4019_ ;
	wire _w4018_ ;
	wire _w4017_ ;
	wire _w4016_ ;
	wire _w4015_ ;
	wire _w4014_ ;
	wire _w4013_ ;
	wire _w4012_ ;
	wire _w4011_ ;
	wire _w4010_ ;
	wire _w4009_ ;
	wire _w4008_ ;
	wire _w4007_ ;
	wire _w4006_ ;
	wire _w4005_ ;
	wire _w4004_ ;
	wire _w4003_ ;
	wire _w4002_ ;
	wire _w4001_ ;
	wire _w4000_ ;
	wire _w3999_ ;
	wire _w3998_ ;
	wire _w3997_ ;
	wire _w3996_ ;
	wire _w3995_ ;
	wire _w3994_ ;
	wire _w3993_ ;
	wire _w3992_ ;
	wire _w3991_ ;
	wire _w3990_ ;
	wire _w3989_ ;
	wire _w3988_ ;
	wire _w3987_ ;
	wire _w3986_ ;
	wire _w3985_ ;
	wire _w3984_ ;
	wire _w3983_ ;
	wire _w3982_ ;
	wire _w3981_ ;
	wire _w3980_ ;
	wire _w3979_ ;
	wire _w3978_ ;
	wire _w3977_ ;
	wire _w3976_ ;
	wire _w3975_ ;
	wire _w3974_ ;
	wire _w3973_ ;
	wire _w3972_ ;
	wire _w3971_ ;
	wire _w3970_ ;
	wire _w3969_ ;
	wire _w3968_ ;
	wire _w3967_ ;
	wire _w3966_ ;
	wire _w3965_ ;
	wire _w3964_ ;
	wire _w3963_ ;
	wire _w3962_ ;
	wire _w3961_ ;
	wire _w3960_ ;
	wire _w3959_ ;
	wire _w3958_ ;
	wire _w3957_ ;
	wire _w3956_ ;
	wire _w3955_ ;
	wire _w3954_ ;
	wire _w3953_ ;
	wire _w3952_ ;
	wire _w3951_ ;
	wire _w3950_ ;
	wire _w3949_ ;
	wire _w3948_ ;
	wire _w3947_ ;
	wire _w3946_ ;
	wire _w3945_ ;
	wire _w3944_ ;
	wire _w3943_ ;
	wire _w3942_ ;
	wire _w3941_ ;
	wire _w3940_ ;
	wire _w3939_ ;
	wire _w3938_ ;
	wire _w3937_ ;
	wire _w3936_ ;
	wire _w3935_ ;
	wire _w3934_ ;
	wire _w3933_ ;
	wire _w3932_ ;
	wire _w3931_ ;
	wire _w3930_ ;
	wire _w3929_ ;
	wire _w3928_ ;
	wire _w3927_ ;
	wire _w3926_ ;
	wire _w3925_ ;
	wire _w3924_ ;
	wire _w3923_ ;
	wire _w3922_ ;
	wire _w3921_ ;
	wire _w3920_ ;
	wire _w3919_ ;
	wire _w3918_ ;
	wire _w3917_ ;
	wire _w3916_ ;
	wire _w3915_ ;
	wire _w3914_ ;
	wire _w3913_ ;
	wire _w3912_ ;
	wire _w3911_ ;
	wire _w3910_ ;
	wire _w3909_ ;
	wire _w3908_ ;
	wire _w3907_ ;
	wire _w3906_ ;
	wire _w3905_ ;
	wire _w3904_ ;
	wire _w3903_ ;
	wire _w3902_ ;
	wire _w3901_ ;
	wire _w3900_ ;
	wire _w3899_ ;
	wire _w3898_ ;
	wire _w3897_ ;
	wire _w3896_ ;
	wire _w3895_ ;
	wire _w3894_ ;
	wire _w3893_ ;
	wire _w3892_ ;
	wire _w3891_ ;
	wire _w3890_ ;
	wire _w3889_ ;
	wire _w3888_ ;
	wire _w3887_ ;
	wire _w3886_ ;
	wire _w3885_ ;
	wire _w3884_ ;
	wire _w3883_ ;
	wire _w3882_ ;
	wire _w3881_ ;
	wire _w3880_ ;
	wire _w3879_ ;
	wire _w3878_ ;
	wire _w3877_ ;
	wire _w3876_ ;
	wire _w3875_ ;
	wire _w3874_ ;
	wire _w3873_ ;
	wire _w3872_ ;
	wire _w3871_ ;
	wire _w3870_ ;
	wire _w3869_ ;
	wire _w3868_ ;
	wire _w3867_ ;
	wire _w3866_ ;
	wire _w3865_ ;
	wire _w3864_ ;
	wire _w3863_ ;
	wire _w3862_ ;
	wire _w3861_ ;
	wire _w3860_ ;
	wire _w3859_ ;
	wire _w3858_ ;
	wire _w3857_ ;
	wire _w3856_ ;
	wire _w3855_ ;
	wire _w3854_ ;
	wire _w3853_ ;
	wire _w3852_ ;
	wire _w3851_ ;
	wire _w3850_ ;
	wire _w3848_ ;
	wire _w3847_ ;
	wire _w3846_ ;
	wire _w3845_ ;
	wire _w3844_ ;
	wire _w3843_ ;
	wire _w3842_ ;
	wire _w3841_ ;
	wire _w3840_ ;
	wire _w3839_ ;
	wire _w3838_ ;
	wire _w3837_ ;
	wire _w3836_ ;
	wire _w3835_ ;
	wire _w3834_ ;
	wire _w3833_ ;
	wire _w3832_ ;
	wire _w3831_ ;
	wire _w3830_ ;
	wire _w3829_ ;
	wire _w3828_ ;
	wire _w3827_ ;
	wire _w3826_ ;
	wire _w3825_ ;
	wire _w3824_ ;
	wire _w3823_ ;
	wire _w3822_ ;
	wire _w3821_ ;
	wire _w3820_ ;
	wire _w3819_ ;
	wire _w3818_ ;
	wire _w3817_ ;
	wire _w3816_ ;
	wire _w3815_ ;
	wire _w3814_ ;
	wire _w3813_ ;
	wire _w3812_ ;
	wire _w3811_ ;
	wire _w3810_ ;
	wire _w3809_ ;
	wire _w3808_ ;
	wire _w3807_ ;
	wire _w3806_ ;
	wire _w3805_ ;
	wire _w3804_ ;
	wire _w3803_ ;
	wire _w3802_ ;
	wire _w3801_ ;
	wire _w3800_ ;
	wire _w3799_ ;
	wire _w3798_ ;
	wire _w3797_ ;
	wire _w3796_ ;
	wire _w3795_ ;
	wire _w3794_ ;
	wire _w3793_ ;
	wire _w3792_ ;
	wire _w3791_ ;
	wire _w3790_ ;
	wire _w3789_ ;
	wire _w3788_ ;
	wire _w3787_ ;
	wire _w3786_ ;
	wire _w3785_ ;
	wire _w3784_ ;
	wire _w3783_ ;
	wire _w3782_ ;
	wire _w3781_ ;
	wire _w3780_ ;
	wire _w3779_ ;
	wire _w3778_ ;
	wire _w3777_ ;
	wire _w3776_ ;
	wire _w3775_ ;
	wire _w3774_ ;
	wire _w3773_ ;
	wire _w3772_ ;
	wire _w3771_ ;
	wire _w3770_ ;
	wire _w3769_ ;
	wire _w3768_ ;
	wire _w3767_ ;
	wire _w3766_ ;
	wire _w3765_ ;
	wire _w3764_ ;
	wire _w3763_ ;
	wire _w3762_ ;
	wire _w3761_ ;
	wire _w3760_ ;
	wire _w3759_ ;
	wire _w3758_ ;
	wire _w3757_ ;
	wire _w3756_ ;
	wire _w3755_ ;
	wire _w3754_ ;
	wire _w3753_ ;
	wire _w3752_ ;
	wire _w3751_ ;
	wire _w3750_ ;
	wire _w3749_ ;
	wire _w3748_ ;
	wire _w3747_ ;
	wire _w3746_ ;
	wire _w3745_ ;
	wire _w3744_ ;
	wire _w3743_ ;
	wire _w3742_ ;
	wire _w3741_ ;
	wire _w3740_ ;
	wire _w3739_ ;
	wire _w3738_ ;
	wire _w3737_ ;
	wire _w3736_ ;
	wire _w3735_ ;
	wire _w3734_ ;
	wire _w3733_ ;
	wire _w3732_ ;
	wire _w3731_ ;
	wire _w3730_ ;
	wire _w3729_ ;
	wire _w3728_ ;
	wire _w3727_ ;
	wire _w3726_ ;
	wire _w3725_ ;
	wire _w3724_ ;
	wire _w3723_ ;
	wire _w3722_ ;
	wire _w3721_ ;
	wire _w3720_ ;
	wire _w3719_ ;
	wire _w3718_ ;
	wire _w3717_ ;
	wire _w3716_ ;
	wire _w3715_ ;
	wire _w3714_ ;
	wire _w3713_ ;
	wire _w3712_ ;
	wire _w3711_ ;
	wire _w3710_ ;
	wire _w3709_ ;
	wire _w3708_ ;
	wire _w3707_ ;
	wire _w3706_ ;
	wire _w3705_ ;
	wire _w3704_ ;
	wire _w3703_ ;
	wire _w3702_ ;
	wire _w3701_ ;
	wire _w3700_ ;
	wire _w3699_ ;
	wire _w3698_ ;
	wire _w3697_ ;
	wire _w3696_ ;
	wire _w3695_ ;
	wire _w3694_ ;
	wire _w3693_ ;
	wire _w3692_ ;
	wire _w3691_ ;
	wire _w3690_ ;
	wire _w3689_ ;
	wire _w3688_ ;
	wire _w3687_ ;
	wire _w3686_ ;
	wire _w3685_ ;
	wire _w3684_ ;
	wire _w3683_ ;
	wire _w3682_ ;
	wire _w3681_ ;
	wire _w3680_ ;
	wire _w3679_ ;
	wire _w3678_ ;
	wire _w3677_ ;
	wire _w3676_ ;
	wire _w3675_ ;
	wire _w3674_ ;
	wire _w3673_ ;
	wire _w3672_ ;
	wire _w3671_ ;
	wire _w3670_ ;
	wire _w3669_ ;
	wire _w3668_ ;
	wire _w3667_ ;
	wire _w3666_ ;
	wire _w3665_ ;
	wire _w3664_ ;
	wire _w3663_ ;
	wire _w3662_ ;
	wire _w3661_ ;
	wire _w3660_ ;
	wire _w3659_ ;
	wire _w3658_ ;
	wire _w3657_ ;
	wire _w3656_ ;
	wire _w3655_ ;
	wire _w3654_ ;
	wire _w3653_ ;
	wire _w3652_ ;
	wire _w3651_ ;
	wire _w3650_ ;
	wire _w3649_ ;
	wire _w3648_ ;
	wire _w3647_ ;
	wire _w3646_ ;
	wire _w3645_ ;
	wire _w3644_ ;
	wire _w3643_ ;
	wire _w3642_ ;
	wire _w3641_ ;
	wire _w3640_ ;
	wire _w3638_ ;
	wire _w3637_ ;
	wire _w3636_ ;
	wire _w3635_ ;
	wire _w3634_ ;
	wire _w3633_ ;
	wire _w3632_ ;
	wire _w3631_ ;
	wire _w3630_ ;
	wire _w3629_ ;
	wire _w3628_ ;
	wire _w3627_ ;
	wire _w3626_ ;
	wire _w3625_ ;
	wire _w3624_ ;
	wire _w3623_ ;
	wire _w3622_ ;
	wire _w3621_ ;
	wire _w3620_ ;
	wire _w3619_ ;
	wire _w3618_ ;
	wire _w3617_ ;
	wire _w3616_ ;
	wire _w3615_ ;
	wire _w3614_ ;
	wire _w3613_ ;
	wire _w3612_ ;
	wire _w3611_ ;
	wire _w3610_ ;
	wire _w3609_ ;
	wire _w3608_ ;
	wire _w3607_ ;
	wire _w3606_ ;
	wire _w3605_ ;
	wire _w3604_ ;
	wire _w3603_ ;
	wire _w3602_ ;
	wire _w3601_ ;
	wire _w3600_ ;
	wire _w3599_ ;
	wire _w3598_ ;
	wire _w3597_ ;
	wire _w3596_ ;
	wire _w3595_ ;
	wire _w3594_ ;
	wire _w3593_ ;
	wire _w3592_ ;
	wire _w3591_ ;
	wire _w3590_ ;
	wire _w3589_ ;
	wire _w3588_ ;
	wire _w3587_ ;
	wire _w3586_ ;
	wire _w3585_ ;
	wire _w3584_ ;
	wire _w3583_ ;
	wire _w3582_ ;
	wire _w3581_ ;
	wire _w3580_ ;
	wire _w3579_ ;
	wire _w3578_ ;
	wire _w3577_ ;
	wire _w3576_ ;
	wire _w3575_ ;
	wire _w3574_ ;
	wire _w3573_ ;
	wire _w3572_ ;
	wire _w3571_ ;
	wire _w3570_ ;
	wire _w3569_ ;
	wire _w3568_ ;
	wire _w3567_ ;
	wire _w3566_ ;
	wire _w3565_ ;
	wire _w3564_ ;
	wire _w3563_ ;
	wire _w3562_ ;
	wire _w3561_ ;
	wire _w3560_ ;
	wire _w3559_ ;
	wire _w3558_ ;
	wire _w3557_ ;
	wire _w3556_ ;
	wire _w3555_ ;
	wire _w3554_ ;
	wire _w3553_ ;
	wire _w3552_ ;
	wire _w3551_ ;
	wire _w3550_ ;
	wire _w3549_ ;
	wire _w3548_ ;
	wire _w3547_ ;
	wire _w3546_ ;
	wire _w3545_ ;
	wire _w3544_ ;
	wire _w3543_ ;
	wire _w3542_ ;
	wire _w3541_ ;
	wire _w3540_ ;
	wire _w3539_ ;
	wire _w3538_ ;
	wire _w3537_ ;
	wire _w3536_ ;
	wire _w3535_ ;
	wire _w3534_ ;
	wire _w3533_ ;
	wire _w3532_ ;
	wire _w3531_ ;
	wire _w3530_ ;
	wire _w3529_ ;
	wire _w3528_ ;
	wire _w3527_ ;
	wire _w3526_ ;
	wire _w3525_ ;
	wire _w3524_ ;
	wire _w3523_ ;
	wire _w3522_ ;
	wire _w3521_ ;
	wire _w3520_ ;
	wire _w3519_ ;
	wire _w3518_ ;
	wire _w3517_ ;
	wire _w3516_ ;
	wire _w3515_ ;
	wire _w3514_ ;
	wire _w3513_ ;
	wire _w3512_ ;
	wire _w3511_ ;
	wire _w3510_ ;
	wire _w3509_ ;
	wire _w3508_ ;
	wire _w3507_ ;
	wire _w3506_ ;
	wire _w3505_ ;
	wire _w3504_ ;
	wire _w3503_ ;
	wire _w3502_ ;
	wire _w3501_ ;
	wire _w3500_ ;
	wire _w3499_ ;
	wire _w3498_ ;
	wire _w3497_ ;
	wire _w3496_ ;
	wire _w3495_ ;
	wire _w3494_ ;
	wire _w3493_ ;
	wire _w3492_ ;
	wire _w3491_ ;
	wire _w3490_ ;
	wire _w3489_ ;
	wire _w3488_ ;
	wire _w3487_ ;
	wire _w3486_ ;
	wire _w3485_ ;
	wire _w3484_ ;
	wire _w3483_ ;
	wire _w3482_ ;
	wire _w3481_ ;
	wire _w3480_ ;
	wire _w3479_ ;
	wire _w3478_ ;
	wire _w3477_ ;
	wire _w3476_ ;
	wire _w3475_ ;
	wire _w3474_ ;
	wire _w3473_ ;
	wire _w3472_ ;
	wire _w3471_ ;
	wire _w3470_ ;
	wire _w3469_ ;
	wire _w3468_ ;
	wire _w3467_ ;
	wire _w3466_ ;
	wire _w3465_ ;
	wire _w3464_ ;
	wire _w3463_ ;
	wire _w3462_ ;
	wire _w3461_ ;
	wire _w3460_ ;
	wire _w3459_ ;
	wire _w3458_ ;
	wire _w3457_ ;
	wire _w3456_ ;
	wire _w3455_ ;
	wire _w3454_ ;
	wire _w3453_ ;
	wire _w3452_ ;
	wire _w3451_ ;
	wire _w3450_ ;
	wire _w3449_ ;
	wire _w3448_ ;
	wire _w3447_ ;
	wire _w3446_ ;
	wire _w3445_ ;
	wire _w3444_ ;
	wire _w3443_ ;
	wire _w3442_ ;
	wire _w3441_ ;
	wire _w3440_ ;
	wire _w3439_ ;
	wire _w3438_ ;
	wire _w3437_ ;
	wire _w3436_ ;
	wire _w3435_ ;
	wire _w3434_ ;
	wire _w3433_ ;
	wire _w3432_ ;
	wire _w3431_ ;
	wire _w3430_ ;
	wire _w3428_ ;
	wire _w3427_ ;
	wire _w3426_ ;
	wire _w3425_ ;
	wire _w3424_ ;
	wire _w3423_ ;
	wire _w3422_ ;
	wire _w3421_ ;
	wire _w3420_ ;
	wire _w3419_ ;
	wire _w3418_ ;
	wire _w3417_ ;
	wire _w3416_ ;
	wire _w3415_ ;
	wire _w3414_ ;
	wire _w3413_ ;
	wire _w3412_ ;
	wire _w3411_ ;
	wire _w3410_ ;
	wire _w3409_ ;
	wire _w3408_ ;
	wire _w3407_ ;
	wire _w3406_ ;
	wire _w3405_ ;
	wire _w3404_ ;
	wire _w3403_ ;
	wire _w3402_ ;
	wire _w3401_ ;
	wire _w3400_ ;
	wire _w3399_ ;
	wire _w3398_ ;
	wire _w3397_ ;
	wire _w3396_ ;
	wire _w3395_ ;
	wire _w3394_ ;
	wire _w3393_ ;
	wire _w3392_ ;
	wire _w3391_ ;
	wire _w3390_ ;
	wire _w3389_ ;
	wire _w3388_ ;
	wire _w3387_ ;
	wire _w3386_ ;
	wire _w3385_ ;
	wire _w3384_ ;
	wire _w3383_ ;
	wire _w3382_ ;
	wire _w3381_ ;
	wire _w3380_ ;
	wire _w3379_ ;
	wire _w3378_ ;
	wire _w3377_ ;
	wire _w3376_ ;
	wire _w3375_ ;
	wire _w3374_ ;
	wire _w3373_ ;
	wire _w3372_ ;
	wire _w3371_ ;
	wire _w3370_ ;
	wire _w3369_ ;
	wire _w3368_ ;
	wire _w3367_ ;
	wire _w3366_ ;
	wire _w3365_ ;
	wire _w3364_ ;
	wire _w3363_ ;
	wire _w3362_ ;
	wire _w3361_ ;
	wire _w3360_ ;
	wire _w3359_ ;
	wire _w3358_ ;
	wire _w3357_ ;
	wire _w3356_ ;
	wire _w3355_ ;
	wire _w3354_ ;
	wire _w3353_ ;
	wire _w3352_ ;
	wire _w3351_ ;
	wire _w3350_ ;
	wire _w3349_ ;
	wire _w3348_ ;
	wire _w3347_ ;
	wire _w3346_ ;
	wire _w3345_ ;
	wire _w3344_ ;
	wire _w3343_ ;
	wire _w3342_ ;
	wire _w3341_ ;
	wire _w3340_ ;
	wire _w3339_ ;
	wire _w3338_ ;
	wire _w3337_ ;
	wire _w3336_ ;
	wire _w3335_ ;
	wire _w3334_ ;
	wire _w3333_ ;
	wire _w3332_ ;
	wire _w3331_ ;
	wire _w3330_ ;
	wire _w3329_ ;
	wire _w3328_ ;
	wire _w3327_ ;
	wire _w3326_ ;
	wire _w3325_ ;
	wire _w3324_ ;
	wire _w3323_ ;
	wire _w3322_ ;
	wire _w3321_ ;
	wire _w3320_ ;
	wire _w3319_ ;
	wire _w3318_ ;
	wire _w3317_ ;
	wire _w3316_ ;
	wire _w3315_ ;
	wire _w3314_ ;
	wire _w3313_ ;
	wire _w3312_ ;
	wire _w3311_ ;
	wire _w3310_ ;
	wire _w3309_ ;
	wire _w3308_ ;
	wire _w3307_ ;
	wire _w3306_ ;
	wire _w3305_ ;
	wire _w3304_ ;
	wire _w3303_ ;
	wire _w3302_ ;
	wire _w3301_ ;
	wire _w3300_ ;
	wire _w3299_ ;
	wire _w3298_ ;
	wire _w3297_ ;
	wire _w3296_ ;
	wire _w3295_ ;
	wire _w3294_ ;
	wire _w3293_ ;
	wire _w3292_ ;
	wire _w3291_ ;
	wire _w3290_ ;
	wire _w3289_ ;
	wire _w3288_ ;
	wire _w3287_ ;
	wire _w3286_ ;
	wire _w3285_ ;
	wire _w3284_ ;
	wire _w3283_ ;
	wire _w3282_ ;
	wire _w3281_ ;
	wire _w3280_ ;
	wire _w3279_ ;
	wire _w3278_ ;
	wire _w3277_ ;
	wire _w3276_ ;
	wire _w3275_ ;
	wire _w3274_ ;
	wire _w3273_ ;
	wire _w3272_ ;
	wire _w3271_ ;
	wire _w3270_ ;
	wire _w3269_ ;
	wire _w3268_ ;
	wire _w3267_ ;
	wire _w3266_ ;
	wire _w3265_ ;
	wire _w3264_ ;
	wire _w3263_ ;
	wire _w3262_ ;
	wire _w3261_ ;
	wire _w3260_ ;
	wire _w3259_ ;
	wire _w3258_ ;
	wire _w3257_ ;
	wire _w3256_ ;
	wire _w3255_ ;
	wire _w3254_ ;
	wire _w3253_ ;
	wire _w3252_ ;
	wire _w3251_ ;
	wire _w3250_ ;
	wire _w3249_ ;
	wire _w3248_ ;
	wire _w3247_ ;
	wire _w3246_ ;
	wire _w3245_ ;
	wire _w3244_ ;
	wire _w3243_ ;
	wire _w3242_ ;
	wire _w3241_ ;
	wire _w3240_ ;
	wire _w3239_ ;
	wire _w3238_ ;
	wire _w3237_ ;
	wire _w3236_ ;
	wire _w3235_ ;
	wire _w3234_ ;
	wire _w3233_ ;
	wire _w3232_ ;
	wire _w3231_ ;
	wire _w3230_ ;
	wire _w3229_ ;
	wire _w3228_ ;
	wire _w3227_ ;
	wire _w3226_ ;
	wire _w3225_ ;
	wire _w3224_ ;
	wire _w3223_ ;
	wire _w3222_ ;
	wire _w3221_ ;
	wire _w3220_ ;
	wire _w3218_ ;
	wire _w3217_ ;
	wire _w3216_ ;
	wire _w3215_ ;
	wire _w3214_ ;
	wire _w3213_ ;
	wire _w3212_ ;
	wire _w3211_ ;
	wire _w3210_ ;
	wire _w3209_ ;
	wire _w3208_ ;
	wire _w3207_ ;
	wire _w3206_ ;
	wire _w3205_ ;
	wire _w3204_ ;
	wire _w3203_ ;
	wire _w3202_ ;
	wire _w3201_ ;
	wire _w3200_ ;
	wire _w3199_ ;
	wire _w3198_ ;
	wire _w3197_ ;
	wire _w3196_ ;
	wire _w3195_ ;
	wire _w3194_ ;
	wire _w3193_ ;
	wire _w3192_ ;
	wire _w3191_ ;
	wire _w3190_ ;
	wire _w3189_ ;
	wire _w3188_ ;
	wire _w3187_ ;
	wire _w3186_ ;
	wire _w3185_ ;
	wire _w3184_ ;
	wire _w3183_ ;
	wire _w3182_ ;
	wire _w3181_ ;
	wire _w3180_ ;
	wire _w3179_ ;
	wire _w3178_ ;
	wire _w3177_ ;
	wire _w3176_ ;
	wire _w3175_ ;
	wire _w3174_ ;
	wire _w3173_ ;
	wire _w3172_ ;
	wire _w3171_ ;
	wire _w3170_ ;
	wire _w3169_ ;
	wire _w3168_ ;
	wire _w3167_ ;
	wire _w3166_ ;
	wire _w3165_ ;
	wire _w3164_ ;
	wire _w3163_ ;
	wire _w3162_ ;
	wire _w3161_ ;
	wire _w3160_ ;
	wire _w3159_ ;
	wire _w3158_ ;
	wire _w3157_ ;
	wire _w3156_ ;
	wire _w3155_ ;
	wire _w3154_ ;
	wire _w3153_ ;
	wire _w3152_ ;
	wire _w3151_ ;
	wire _w3150_ ;
	wire _w3149_ ;
	wire _w3148_ ;
	wire _w3147_ ;
	wire _w3146_ ;
	wire _w3145_ ;
	wire _w3144_ ;
	wire _w3143_ ;
	wire _w3142_ ;
	wire _w3141_ ;
	wire _w3140_ ;
	wire _w3139_ ;
	wire _w3138_ ;
	wire _w3137_ ;
	wire _w3136_ ;
	wire _w3135_ ;
	wire _w3134_ ;
	wire _w3133_ ;
	wire _w3132_ ;
	wire _w3131_ ;
	wire _w3130_ ;
	wire _w3129_ ;
	wire _w3128_ ;
	wire _w3127_ ;
	wire _w3126_ ;
	wire _w3125_ ;
	wire _w3124_ ;
	wire _w3123_ ;
	wire _w3122_ ;
	wire _w3121_ ;
	wire _w3120_ ;
	wire _w3119_ ;
	wire _w3118_ ;
	wire _w3117_ ;
	wire _w3116_ ;
	wire _w3115_ ;
	wire _w3114_ ;
	wire _w3113_ ;
	wire _w3112_ ;
	wire _w3111_ ;
	wire _w3110_ ;
	wire _w3109_ ;
	wire _w3108_ ;
	wire _w3107_ ;
	wire _w3106_ ;
	wire _w3105_ ;
	wire _w3104_ ;
	wire _w3103_ ;
	wire _w3102_ ;
	wire _w3101_ ;
	wire _w3100_ ;
	wire _w3099_ ;
	wire _w3098_ ;
	wire _w3097_ ;
	wire _w3096_ ;
	wire _w3095_ ;
	wire _w3094_ ;
	wire _w3093_ ;
	wire _w3092_ ;
	wire _w3091_ ;
	wire _w3090_ ;
	wire _w3089_ ;
	wire _w3088_ ;
	wire _w3087_ ;
	wire _w3086_ ;
	wire _w3085_ ;
	wire _w3084_ ;
	wire _w3083_ ;
	wire _w3082_ ;
	wire _w3081_ ;
	wire _w3080_ ;
	wire _w3079_ ;
	wire _w3078_ ;
	wire _w3077_ ;
	wire _w3076_ ;
	wire _w3075_ ;
	wire _w3074_ ;
	wire _w3073_ ;
	wire _w3072_ ;
	wire _w3071_ ;
	wire _w3070_ ;
	wire _w3069_ ;
	wire _w3068_ ;
	wire _w3067_ ;
	wire _w3066_ ;
	wire _w3065_ ;
	wire _w3064_ ;
	wire _w3063_ ;
	wire _w3062_ ;
	wire _w3061_ ;
	wire _w3060_ ;
	wire _w3059_ ;
	wire _w3058_ ;
	wire _w3057_ ;
	wire _w3056_ ;
	wire _w3055_ ;
	wire _w3054_ ;
	wire _w3053_ ;
	wire _w3052_ ;
	wire _w3051_ ;
	wire _w3050_ ;
	wire _w3049_ ;
	wire _w3048_ ;
	wire _w3047_ ;
	wire _w3046_ ;
	wire _w3045_ ;
	wire _w3044_ ;
	wire _w3043_ ;
	wire _w3042_ ;
	wire _w3041_ ;
	wire _w3040_ ;
	wire _w3039_ ;
	wire _w3038_ ;
	wire _w3037_ ;
	wire _w3036_ ;
	wire _w3035_ ;
	wire _w3034_ ;
	wire _w3033_ ;
	wire _w3032_ ;
	wire _w3031_ ;
	wire _w3030_ ;
	wire _w3029_ ;
	wire _w3028_ ;
	wire _w3027_ ;
	wire _w3026_ ;
	wire _w3025_ ;
	wire _w3024_ ;
	wire _w3023_ ;
	wire _w3022_ ;
	wire _w3021_ ;
	wire _w3020_ ;
	wire _w3019_ ;
	wire _w3018_ ;
	wire _w3017_ ;
	wire _w3016_ ;
	wire _w3015_ ;
	wire _w3014_ ;
	wire _w3013_ ;
	wire _w3012_ ;
	wire _w3011_ ;
	wire _w3010_ ;
	wire _w3009_ ;
	wire _w3008_ ;
	wire _w3007_ ;
	wire _w3006_ ;
	wire _w3005_ ;
	wire _w3004_ ;
	wire _w3003_ ;
	wire _w3002_ ;
	wire _w3001_ ;
	wire _w3000_ ;
	wire _w2999_ ;
	wire _w2998_ ;
	wire _w2997_ ;
	wire _w2996_ ;
	wire _w2995_ ;
	wire _w2994_ ;
	wire _w2993_ ;
	wire _w2992_ ;
	wire _w2991_ ;
	wire _w2990_ ;
	wire _w2989_ ;
	wire _w2988_ ;
	wire _w2987_ ;
	wire _w2986_ ;
	wire _w2985_ ;
	wire _w2984_ ;
	wire _w2983_ ;
	wire _w2982_ ;
	wire _w2981_ ;
	wire _w2980_ ;
	wire _w2979_ ;
	wire _w2978_ ;
	wire _w2977_ ;
	wire _w2976_ ;
	wire _w2975_ ;
	wire _w2974_ ;
	wire _w2973_ ;
	wire _w2972_ ;
	wire _w2971_ ;
	wire _w2970_ ;
	wire _w2969_ ;
	wire _w2968_ ;
	wire _w2967_ ;
	wire _w2966_ ;
	wire _w2965_ ;
	wire _w2964_ ;
	wire _w2963_ ;
	wire _w2962_ ;
	wire _w2961_ ;
	wire _w2960_ ;
	wire _w2959_ ;
	wire _w2958_ ;
	wire _w2957_ ;
	wire _w2956_ ;
	wire _w2955_ ;
	wire _w2954_ ;
	wire _w2953_ ;
	wire _w2952_ ;
	wire _w2951_ ;
	wire _w2950_ ;
	wire _w2949_ ;
	wire _w2948_ ;
	wire _w2947_ ;
	wire _w2946_ ;
	wire _w2945_ ;
	wire _w2944_ ;
	wire _w2943_ ;
	wire _w2942_ ;
	wire _w2941_ ;
	wire _w2940_ ;
	wire _w2939_ ;
	wire _w2938_ ;
	wire _w2937_ ;
	wire _w2936_ ;
	wire _w2935_ ;
	wire _w2934_ ;
	wire _w2933_ ;
	wire _w2932_ ;
	wire _w2931_ ;
	wire _w2930_ ;
	wire _w2929_ ;
	wire _w2928_ ;
	wire _w2927_ ;
	wire _w2926_ ;
	wire _w2925_ ;
	wire _w2924_ ;
	wire _w2923_ ;
	wire _w2922_ ;
	wire _w2921_ ;
	wire _w2920_ ;
	wire _w2919_ ;
	wire _w2918_ ;
	wire _w2917_ ;
	wire _w2916_ ;
	wire _w2915_ ;
	wire _w2914_ ;
	wire _w2913_ ;
	wire _w2912_ ;
	wire _w2911_ ;
	wire _w2910_ ;
	wire _w2909_ ;
	wire _w2908_ ;
	wire _w2907_ ;
	wire _w2906_ ;
	wire _w2905_ ;
	wire _w2904_ ;
	wire _w2903_ ;
	wire _w2902_ ;
	wire _w2901_ ;
	wire _w2900_ ;
	wire _w2899_ ;
	wire _w2898_ ;
	wire _w2897_ ;
	wire _w2896_ ;
	wire _w2895_ ;
	wire _w2894_ ;
	wire _w2893_ ;
	wire _w2892_ ;
	wire _w2891_ ;
	wire _w2890_ ;
	wire _w2889_ ;
	wire _w2888_ ;
	wire _w2887_ ;
	wire _w2886_ ;
	wire _w2885_ ;
	wire _w2884_ ;
	wire _w2883_ ;
	wire _w2882_ ;
	wire _w2881_ ;
	wire _w2880_ ;
	wire _w2879_ ;
	wire _w2878_ ;
	wire _w2877_ ;
	wire _w2876_ ;
	wire _w2875_ ;
	wire _w2874_ ;
	wire _w2873_ ;
	wire _w2872_ ;
	wire _w2871_ ;
	wire _w2870_ ;
	wire _w2869_ ;
	wire _w2868_ ;
	wire _w2867_ ;
	wire _w2866_ ;
	wire _w2865_ ;
	wire _w2864_ ;
	wire _w2863_ ;
	wire _w2862_ ;
	wire _w2861_ ;
	wire _w2860_ ;
	wire _w2859_ ;
	wire _w2290_ ;
	wire _w2289_ ;
	wire _w2288_ ;
	wire _w2287_ ;
	wire _w2286_ ;
	wire _w2285_ ;
	wire _w2284_ ;
	wire _w2283_ ;
	wire _w2282_ ;
	wire _w2281_ ;
	wire _w2280_ ;
	wire _w2279_ ;
	wire _w2278_ ;
	wire _w2277_ ;
	wire _w2276_ ;
	wire _w2275_ ;
	wire _w2274_ ;
	wire _w2273_ ;
	wire _w2272_ ;
	wire _w2271_ ;
	wire _w2270_ ;
	wire _w2269_ ;
	wire _w2268_ ;
	wire _w2266_ ;
	wire _w2265_ ;
	wire _w2264_ ;
	wire _w2263_ ;
	wire _w2262_ ;
	wire _w2261_ ;
	wire _w2260_ ;
	wire _w2259_ ;
	wire _w2258_ ;
	wire _w2257_ ;
	wire _w2256_ ;
	wire _w2255_ ;
	wire _w2254_ ;
	wire _w2253_ ;
	wire _w2252_ ;
	wire _w2251_ ;
	wire _w2250_ ;
	wire _w2249_ ;
	wire _w2248_ ;
	wire _w2247_ ;
	wire _w2246_ ;
	wire _w2245_ ;
	wire _w2244_ ;
	wire _w2243_ ;
	wire _w2242_ ;
	wire _w2241_ ;
	wire _w2240_ ;
	wire _w2239_ ;
	wire _w2238_ ;
	wire _w2237_ ;
	wire _w2236_ ;
	wire _w2235_ ;
	wire _w2234_ ;
	wire _w2233_ ;
	wire _w2232_ ;
	wire _w2231_ ;
	wire _w2230_ ;
	wire _w2229_ ;
	wire _w2228_ ;
	wire _w2227_ ;
	wire _w2226_ ;
	wire _w2225_ ;
	wire _w2224_ ;
	wire _w2223_ ;
	wire _w2222_ ;
	wire _w2221_ ;
	wire _w2220_ ;
	wire _w2219_ ;
	wire _w2218_ ;
	wire _w2217_ ;
	wire _w2216_ ;
	wire _w2215_ ;
	wire _w2214_ ;
	wire _w2213_ ;
	wire _w2212_ ;
	wire _w2211_ ;
	wire _w2210_ ;
	wire _w2209_ ;
	wire _w2208_ ;
	wire _w2207_ ;
	wire _w2206_ ;
	wire _w2205_ ;
	wire _w2204_ ;
	wire _w2203_ ;
	wire _w2202_ ;
	wire _w2201_ ;
	wire _w2200_ ;
	wire _w2199_ ;
	wire _w2198_ ;
	wire _w2197_ ;
	wire _w2196_ ;
	wire _w2195_ ;
	wire _w2194_ ;
	wire _w2193_ ;
	wire _w2192_ ;
	wire _w2191_ ;
	wire _w2190_ ;
	wire _w2189_ ;
	wire _w2188_ ;
	wire _w2187_ ;
	wire _w2186_ ;
	wire _w2185_ ;
	wire _w2184_ ;
	wire _w2183_ ;
	wire _w2182_ ;
	wire _w2181_ ;
	wire _w3429_ ;
	wire _w1072_ ;
	wire _w6159_ ;
	wire _w2180_ ;
	wire _w2179_ ;
	wire _w2178_ ;
	wire _w2177_ ;
	wire _w2176_ ;
	wire _w2175_ ;
	wire _w2174_ ;
	wire _w2173_ ;
	wire _w2172_ ;
	wire _w2171_ ;
	wire _w2170_ ;
	wire _w2169_ ;
	wire _w2168_ ;
	wire _w2167_ ;
	wire _w2166_ ;
	wire _w2165_ ;
	wire _w2164_ ;
	wire _w2163_ ;
	wire _w2162_ ;
	wire _w2161_ ;
	wire _w2160_ ;
	wire _w2159_ ;
	wire _w2158_ ;
	wire _w2157_ ;
	wire _w2156_ ;
	wire _w2155_ ;
	wire _w2153_ ;
	wire _w2152_ ;
	wire _w2151_ ;
	wire _w2150_ ;
	wire _w2149_ ;
	wire _w2148_ ;
	wire _w2147_ ;
	wire _w2146_ ;
	wire _w2145_ ;
	wire _w2144_ ;
	wire _w2143_ ;
	wire _w2142_ ;
	wire _w2141_ ;
	wire _w2140_ ;
	wire _w2139_ ;
	wire _w2138_ ;
	wire _w2137_ ;
	wire _w2136_ ;
	wire _w2135_ ;
	wire _w2134_ ;
	wire _w2133_ ;
	wire _w2132_ ;
	wire _w2131_ ;
	wire _w2130_ ;
	wire _w2129_ ;
	wire _w2128_ ;
	wire _w2127_ ;
	wire _w2126_ ;
	wire _w2125_ ;
	wire _w2124_ ;
	wire _w2123_ ;
	wire _w2122_ ;
	wire _w2121_ ;
	wire _w2120_ ;
	wire _w2119_ ;
	wire _w2118_ ;
	wire _w2117_ ;
	wire _w2116_ ;
	wire _w2115_ ;
	wire _w2114_ ;
	wire _w2113_ ;
	wire _w2112_ ;
	wire _w2111_ ;
	wire _w2110_ ;
	wire _w2109_ ;
	wire _w2108_ ;
	wire _w2107_ ;
	wire _w2106_ ;
	wire _w2105_ ;
	wire _w2104_ ;
	wire _w2103_ ;
	wire _w2102_ ;
	wire _w2101_ ;
	wire _w2100_ ;
	wire _w2099_ ;
	wire _w2098_ ;
	wire _w2097_ ;
	wire _w2096_ ;
	wire _w2095_ ;
	wire _w2094_ ;
	wire _w2093_ ;
	wire _w2092_ ;
	wire _w2091_ ;
	wire _w2090_ ;
	wire _w2089_ ;
	wire _w2088_ ;
	wire _w2087_ ;
	wire _w2086_ ;
	wire _w2085_ ;
	wire _w2084_ ;
	wire _w2083_ ;
	wire _w2082_ ;
	wire _w2081_ ;
	wire _w2080_ ;
	wire _w2079_ ;
	wire _w2078_ ;
	wire _w2077_ ;
	wire _w2076_ ;
	wire _w2075_ ;
	wire _w2074_ ;
	wire _w2073_ ;
	wire _w2072_ ;
	wire _w2071_ ;
	wire _w2070_ ;
	wire _w2069_ ;
	wire _w2068_ ;
	wire _w2067_ ;
	wire _w2066_ ;
	wire _w2065_ ;
	wire _w2064_ ;
	wire _w2063_ ;
	wire _w2062_ ;
	wire _w2061_ ;
	wire _w2060_ ;
	wire _w2059_ ;
	wire _w2058_ ;
	wire _w2057_ ;
	wire _w2056_ ;
	wire _w2055_ ;
	wire _w2054_ ;
	wire _w2053_ ;
	wire _w2052_ ;
	wire _w2051_ ;
	wire _w2050_ ;
	wire _w2049_ ;
	wire _w2048_ ;
	wire _w2047_ ;
	wire _w2046_ ;
	wire _w2045_ ;
	wire _w2044_ ;
	wire _w2043_ ;
	wire _w2042_ ;
	wire _w2041_ ;
	wire _w2040_ ;
	wire _w2039_ ;
	wire _w2038_ ;
	wire _w2037_ ;
	wire _w2036_ ;
	wire _w2035_ ;
	wire _w2034_ ;
	wire _w2032_ ;
	wire _w2031_ ;
	wire _w2030_ ;
	wire _w2029_ ;
	wire _w2028_ ;
	wire _w2027_ ;
	wire _w2026_ ;
	wire _w2025_ ;
	wire _w2024_ ;
	wire _w2023_ ;
	wire _w2022_ ;
	wire _w2021_ ;
	wire _w2020_ ;
	wire _w2019_ ;
	wire _w2018_ ;
	wire _w2017_ ;
	wire _w2016_ ;
	wire _w2015_ ;
	wire _w2014_ ;
	wire _w2013_ ;
	wire _w2012_ ;
	wire _w2011_ ;
	wire _w2010_ ;
	wire _w2009_ ;
	wire _w2008_ ;
	wire _w2007_ ;
	wire _w1876_ ;
	wire _w1875_ ;
	wire _w1874_ ;
	wire _w1872_ ;
	wire _w1871_ ;
	wire _w1870_ ;
	wire _w1869_ ;
	wire _w1868_ ;
	wire _w1867_ ;
	wire _w1866_ ;
	wire _w1865_ ;
	wire _w1864_ ;
	wire _w1863_ ;
	wire _w1862_ ;
	wire _w1861_ ;
	wire _w1860_ ;
	wire _w1859_ ;
	wire _w1858_ ;
	wire _w1857_ ;
	wire _w1856_ ;
	wire _w1855_ ;
	wire _w1854_ ;
	wire _w1853_ ;
	wire _w1852_ ;
	wire _w1851_ ;
	wire _w1850_ ;
	wire _w1849_ ;
	wire _w1848_ ;
	wire _w1847_ ;
	wire _w1846_ ;
	wire _w1845_ ;
	wire _w1844_ ;
	wire _w1843_ ;
	wire _w2154_ ;
	wire _w1842_ ;
	wire _w1841_ ;
	wire _w1840_ ;
	wire _w1839_ ;
	wire _w1838_ ;
	wire _w1837_ ;
	wire _w1836_ ;
	wire _w1835_ ;
	wire _w1833_ ;
	wire _w1832_ ;
	wire _w1831_ ;
	wire _w1830_ ;
	wire _w1829_ ;
	wire _w1828_ ;
	wire _w1827_ ;
	wire _w1826_ ;
	wire _w1825_ ;
	wire _w1824_ ;
	wire _w1822_ ;
	wire _w1821_ ;
	wire _w1820_ ;
	wire _w1819_ ;
	wire _w1818_ ;
	wire _w1817_ ;
	wire _w1816_ ;
	wire _w1815_ ;
	wire _w1814_ ;
	wire _w1813_ ;
	wire _w1812_ ;
	wire _w1811_ ;
	wire _w1810_ ;
	wire _w1809_ ;
	wire _w1778_ ;
	wire _w1777_ ;
	wire _w1776_ ;
	wire _w1774_ ;
	wire _w1773_ ;
	wire _w1772_ ;
	wire _w1771_ ;
	wire _w1770_ ;
	wire _w1769_ ;
	wire _w1767_ ;
	wire _w1766_ ;
	wire _w1765_ ;
	wire _w1764_ ;
	wire _w1763_ ;
	wire _w1759_ ;
	wire _w1768_ ;
	wire _w1834_ ;
	wire _w1780_ ;
	wire _w1890_ ;
	wire _w1806_ ;
	wire _w1761_ ;
	wire _w1775_ ;
	wire _w1873_ ;
	wire _w2033_ ;
	wire _w3849_ ;
	wire _w1492_ ;
	wire _w6579_ ;
	wire _w2601_ ;
	wire _w2006_ ;
	wire _w1787_ ;
	wire _w1755_ ;
	wire _w2267_ ;
	wire _w2321_ ;
	wire _w1902_ ;
	wire _w1756_ ;
	wire _w1757_ ;
	wire _w1758_ ;
	wire _w1760_ ;
	wire _w1762_ ;
	wire _w1779_ ;
	wire _w1781_ ;
	wire _w1782_ ;
	wire _w1783_ ;
	wire _w1784_ ;
	wire _w1785_ ;
	wire _w1786_ ;
	wire _w1788_ ;
	wire _w1789_ ;
	wire _w1823_ ;
	wire _w3639_ ;
	wire _w1282_ ;
	wire _w6369_ ;
	wire _w2391_ ;
	wire _w1796_ ;
	wire _w1790_ ;
	wire _w1791_ ;
	wire _w1792_ ;
	wire _w1793_ ;
	wire _w1794_ ;
	wire _w1795_ ;
	wire _w1797_ ;
	wire _w1798_ ;
	wire _w1799_ ;
	wire _w1800_ ;
	wire _w1801_ ;
	wire _w1802_ ;
	wire _w1803_ ;
	wire _w1804_ ;
	wire _w1805_ ;
	wire _w1807_ ;
	wire _w1808_ ;
	wire _w1877_ ;
	wire _w1878_ ;
	wire _w1879_ ;
	wire _w1880_ ;
	wire _w1881_ ;
	wire _w1882_ ;
	wire _w1883_ ;
	wire _w1884_ ;
	wire _w1885_ ;
	wire _w1886_ ;
	wire _w1887_ ;
	wire _w1888_ ;
	wire _w1889_ ;
	wire _w1891_ ;
	wire _w1892_ ;
	wire _w1893_ ;
	wire _w1894_ ;
	wire _w1895_ ;
	wire _w1896_ ;
	wire _w1897_ ;
	wire _w1898_ ;
	wire _w1899_ ;
	wire _w1900_ ;
	wire _w1901_ ;
	wire _w1903_ ;
	wire _w1904_ ;
	wire _w1905_ ;
	wire _w1906_ ;
	wire _w1907_ ;
	wire _w1908_ ;
	wire _w1909_ ;
	wire _w1910_ ;
	wire _w1911_ ;
	wire _w1912_ ;
	wire _w1913_ ;
	wire _w1914_ ;
	wire _w1915_ ;
	wire _w1916_ ;
	wire _w1917_ ;
	wire _w1918_ ;
	wire _w1919_ ;
	wire _w1920_ ;
	wire _w1921_ ;
	wire _w1922_ ;
	wire _w1923_ ;
	wire _w1924_ ;
	wire _w1925_ ;
	wire _w1926_ ;
	wire _w1927_ ;
	wire _w1928_ ;
	wire _w1929_ ;
	wire _w1930_ ;
	wire _w1931_ ;
	wire _w1932_ ;
	wire _w1933_ ;
	wire _w1934_ ;
	wire _w1935_ ;
	wire _w1936_ ;
	wire _w1937_ ;
	wire _w1938_ ;
	wire _w1939_ ;
	wire _w1940_ ;
	wire _w1941_ ;
	wire _w1942_ ;
	wire _w1943_ ;
	wire _w3219_ ;
	wire _w862_ ;
	wire _w5949_ ;
	wire _w1971_ ;
	wire _w1944_ ;
	wire _w1945_ ;
	wire _w1946_ ;
	wire _w1947_ ;
	wire _w1948_ ;
	wire _w1949_ ;
	wire _w1950_ ;
	wire _w1951_ ;
	wire _w1952_ ;
	wire _w1953_ ;
	wire _w1954_ ;
	wire _w1955_ ;
	wire _w1956_ ;
	wire _w1957_ ;
	wire _w1958_ ;
	wire _w1959_ ;
	wire _w1960_ ;
	wire _w1961_ ;
	wire _w1962_ ;
	wire _w1963_ ;
	wire _w1964_ ;
	wire _w1965_ ;
	wire _w1966_ ;
	wire _w1967_ ;
	wire _w1968_ ;
	wire _w1969_ ;
	wire _w1970_ ;
	wire _w1972_ ;
	wire _w1973_ ;
	wire _w1974_ ;
	wire _w1975_ ;
	wire _w1976_ ;
	wire _w1977_ ;
	wire _w1978_ ;
	wire _w1979_ ;
	wire _w1980_ ;
	wire _w1981_ ;
	wire _w1982_ ;
	wire _w1983_ ;
	wire _w1984_ ;
	wire _w1985_ ;
	wire _w1986_ ;
	wire _w1987_ ;
	wire _w1988_ ;
	wire _w1989_ ;
	wire _w1990_ ;
	wire _w1991_ ;
	wire _w1992_ ;
	wire _w1993_ ;
	wire _w1994_ ;
	wire _w1995_ ;
	wire _w1996_ ;
	wire _w1997_ ;
	wire _w1998_ ;
	wire _w1999_ ;
	wire _w2000_ ;
	wire _w2001_ ;
	wire _w2002_ ;
	wire _w2003_ ;
	wire _w2004_ ;
	wire _w2005_ ;
	wire _w2291_ ;
	wire _w2292_ ;
	wire _w2293_ ;
	wire _w2294_ ;
	wire _w2295_ ;
	wire _w2296_ ;
	wire _w2297_ ;
	wire _w2298_ ;
	wire _w2299_ ;
	wire _w2300_ ;
	wire _w2301_ ;
	wire _w2302_ ;
	wire _w2303_ ;
	wire _w2304_ ;
	wire _w2305_ ;
	wire _w2306_ ;
	wire _w2307_ ;
	wire _w2308_ ;
	wire _w2309_ ;
	wire _w2310_ ;
	wire _w2311_ ;
	wire _w2312_ ;
	wire _w2313_ ;
	wire _w2314_ ;
	wire _w2315_ ;
	wire _w2316_ ;
	wire _w2317_ ;
	wire _w2318_ ;
	wire _w2319_ ;
	wire _w2320_ ;
	wire _w2322_ ;
	wire _w2323_ ;
	wire _w2324_ ;
	wire _w2325_ ;
	wire _w2326_ ;
	wire _w2327_ ;
	wire _w2328_ ;
	wire _w2329_ ;
	wire _w2330_ ;
	wire _w2331_ ;
	wire _w2332_ ;
	wire _w2333_ ;
	wire _w2334_ ;
	wire _w2335_ ;
	wire _w2336_ ;
	wire _w2337_ ;
	wire _w2338_ ;
	wire _w2339_ ;
	wire _w2340_ ;
	wire _w2341_ ;
	wire _w2342_ ;
	wire _w2343_ ;
	wire _w2344_ ;
	wire _w2345_ ;
	wire _w2346_ ;
	wire _w2347_ ;
	wire _w2348_ ;
	wire _w2349_ ;
	wire _w2350_ ;
	wire _w2351_ ;
	wire _w2352_ ;
	wire _w2353_ ;
	wire _w2354_ ;
	wire _w2355_ ;
	wire _w2356_ ;
	wire _w2357_ ;
	wire _w2358_ ;
	wire _w2359_ ;
	wire _w2360_ ;
	wire _w2361_ ;
	wire _w2362_ ;
	wire _w2363_ ;
	wire _w2364_ ;
	wire _w2365_ ;
	wire _w2366_ ;
	wire _w2367_ ;
	wire _w2368_ ;
	wire _w2369_ ;
	wire _w2370_ ;
	wire _w2371_ ;
	wire _w2372_ ;
	wire _w2373_ ;
	wire _w2374_ ;
	wire _w2375_ ;
	wire _w2376_ ;
	wire _w2377_ ;
	wire _w2378_ ;
	wire _w2379_ ;
	wire _w2380_ ;
	wire _w2381_ ;
	wire _w2382_ ;
	wire _w2383_ ;
	wire _w2384_ ;
	wire _w2385_ ;
	wire _w2386_ ;
	wire _w2387_ ;
	wire _w2388_ ;
	wire _w2389_ ;
	wire _w2390_ ;
	wire _w2392_ ;
	wire _w2393_ ;
	wire _w2394_ ;
	wire _w2395_ ;
	wire _w2396_ ;
	wire _w2397_ ;
	wire _w2398_ ;
	wire _w2399_ ;
	wire _w2400_ ;
	wire _w2401_ ;
	wire _w2402_ ;
	wire _w2403_ ;
	wire _w2404_ ;
	wire _w2405_ ;
	wire _w2406_ ;
	wire _w2407_ ;
	wire _w2408_ ;
	wire _w2409_ ;
	wire _w2410_ ;
	wire _w2411_ ;
	wire _w2412_ ;
	wire _w2413_ ;
	wire _w2414_ ;
	wire _w2415_ ;
	wire _w2416_ ;
	wire _w2417_ ;
	wire _w2418_ ;
	wire _w2419_ ;
	wire _w2420_ ;
	wire _w2421_ ;
	wire _w2422_ ;
	wire _w2423_ ;
	wire _w2424_ ;
	wire _w2425_ ;
	wire _w2426_ ;
	wire _w2427_ ;
	wire _w2428_ ;
	wire _w2429_ ;
	wire _w2430_ ;
	wire _w2431_ ;
	wire _w2432_ ;
	wire _w2433_ ;
	wire _w2434_ ;
	wire _w2435_ ;
	wire _w2436_ ;
	wire _w2437_ ;
	wire _w2438_ ;
	wire _w2439_ ;
	wire _w2440_ ;
	wire _w2441_ ;
	wire _w2442_ ;
	wire _w2443_ ;
	wire _w2444_ ;
	wire _w2445_ ;
	wire _w2446_ ;
	wire _w2447_ ;
	wire _w2448_ ;
	wire _w2449_ ;
	wire _w2450_ ;
	wire _w2451_ ;
	wire _w2452_ ;
	wire _w2453_ ;
	wire _w2454_ ;
	wire _w2455_ ;
	wire _w2456_ ;
	wire _w2457_ ;
	wire _w2458_ ;
	wire _w2459_ ;
	wire _w10376_ ;
	wire _w103_ ;
	wire _w5190_ ;
	wire _w2460_ ;
	wire _w2461_ ;
	wire _w2462_ ;
	wire _w2463_ ;
	wire _w2464_ ;
	wire _w2465_ ;
	wire _w2466_ ;
	wire _w2467_ ;
	wire _w2468_ ;
	wire _w2469_ ;
	wire _w2470_ ;
	wire _w2471_ ;
	wire _w2472_ ;
	wire _w2473_ ;
	wire _w2474_ ;
	wire _w2475_ ;
	wire _w2476_ ;
	wire _w2477_ ;
	wire _w2478_ ;
	wire _w2479_ ;
	wire _w2480_ ;
	wire _w2481_ ;
	wire _w2482_ ;
	wire _w2483_ ;
	wire _w2484_ ;
	wire _w2485_ ;
	wire _w2486_ ;
	wire _w2487_ ;
	wire _w2488_ ;
	wire _w2489_ ;
	wire _w2490_ ;
	wire _w2491_ ;
	wire _w2492_ ;
	wire _w2493_ ;
	wire _w2494_ ;
	wire _w2495_ ;
	wire _w2496_ ;
	wire _w2497_ ;
	wire _w2498_ ;
	wire _w2499_ ;
	wire _w2500_ ;
	wire _w2501_ ;
	wire _w2502_ ;
	wire _w2503_ ;
	wire _w2504_ ;
	wire _w2505_ ;
	wire _w2506_ ;
	wire _w2507_ ;
	wire _w2508_ ;
	wire _w2509_ ;
	wire _w2510_ ;
	wire _w2511_ ;
	wire _w2512_ ;
	wire _w2513_ ;
	wire _w2514_ ;
	wire _w2515_ ;
	wire _w2516_ ;
	wire _w2517_ ;
	wire _w2518_ ;
	wire _w2519_ ;
	wire _w2520_ ;
	wire _w2521_ ;
	wire _w2522_ ;
	wire _w2523_ ;
	wire _w2524_ ;
	wire _w2525_ ;
	wire _w2526_ ;
	wire _w2527_ ;
	wire _w2528_ ;
	wire _w2529_ ;
	wire _w2530_ ;
	wire _w2531_ ;
	wire _w2532_ ;
	wire _w2533_ ;
	wire _w2534_ ;
	wire _w2535_ ;
	wire _w2536_ ;
	wire _w2537_ ;
	wire _w2538_ ;
	wire _w2539_ ;
	wire _w2540_ ;
	wire _w2541_ ;
	wire _w2542_ ;
	wire _w2543_ ;
	wire _w2544_ ;
	wire _w2545_ ;
	wire _w2546_ ;
	wire _w2547_ ;
	wire _w2548_ ;
	wire _w2549_ ;
	wire _w2550_ ;
	wire _w2551_ ;
	wire _w2552_ ;
	wire _w2553_ ;
	wire _w2554_ ;
	wire _w2555_ ;
	wire _w2556_ ;
	wire _w2557_ ;
	wire _w2558_ ;
	wire _w2559_ ;
	wire _w2560_ ;
	wire _w2561_ ;
	wire _w2562_ ;
	wire _w2563_ ;
	wire _w2564_ ;
	wire _w2565_ ;
	wire _w2566_ ;
	wire _w2567_ ;
	wire _w2568_ ;
	wire _w2569_ ;
	wire _w2570_ ;
	wire _w2571_ ;
	wire _w2572_ ;
	wire _w2573_ ;
	wire _w2574_ ;
	wire _w2575_ ;
	wire _w2576_ ;
	wire _w2577_ ;
	wire _w2578_ ;
	wire _w2579_ ;
	wire _w2580_ ;
	wire _w2581_ ;
	wire _w2582_ ;
	wire _w2583_ ;
	wire _w2584_ ;
	wire _w2585_ ;
	wire _w2586_ ;
	wire _w2587_ ;
	wire _w2588_ ;
	wire _w2589_ ;
	wire _w2590_ ;
	wire _w2591_ ;
	wire _w2592_ ;
	wire _w2593_ ;
	wire _w2594_ ;
	wire _w2595_ ;
	wire _w2596_ ;
	wire _w2597_ ;
	wire _w2598_ ;
	wire _w2599_ ;
	wire _w2600_ ;
	wire _w2602_ ;
	wire _w2603_ ;
	wire _w2604_ ;
	wire _w2605_ ;
	wire _w2606_ ;
	wire _w2607_ ;
	wire _w2608_ ;
	wire _w2609_ ;
	wire _w2610_ ;
	wire _w2611_ ;
	wire _w2612_ ;
	wire _w2613_ ;
	wire _w2614_ ;
	wire _w2615_ ;
	wire _w2616_ ;
	wire _w2617_ ;
	wire _w2618_ ;
	wire _w2619_ ;
	wire _w2620_ ;
	wire _w2621_ ;
	wire _w2622_ ;
	wire _w2623_ ;
	wire _w2624_ ;
	wire _w2625_ ;
	wire _w2626_ ;
	wire _w2627_ ;
	wire _w2628_ ;
	wire _w2629_ ;
	wire _w2630_ ;
	wire _w2631_ ;
	wire _w2632_ ;
	wire _w2633_ ;
	wire _w2634_ ;
	wire _w2635_ ;
	wire _w2636_ ;
	wire _w2637_ ;
	wire _w2638_ ;
	wire _w2639_ ;
	wire _w2640_ ;
	wire _w2641_ ;
	wire _w2642_ ;
	wire _w2643_ ;
	wire _w2644_ ;
	wire _w2645_ ;
	wire _w2646_ ;
	wire _w2647_ ;
	wire _w2648_ ;
	wire _w2649_ ;
	wire _w2650_ ;
	wire _w2651_ ;
	wire _w2652_ ;
	wire _w2653_ ;
	wire _w2654_ ;
	wire _w2655_ ;
	wire _w2656_ ;
	wire _w2657_ ;
	wire _w2658_ ;
	wire _w2659_ ;
	wire _w2660_ ;
	wire _w2661_ ;
	wire _w2662_ ;
	wire _w2663_ ;
	wire _w2664_ ;
	wire _w2665_ ;
	wire _w2666_ ;
	wire _w2667_ ;
	wire _w2668_ ;
	wire _w2669_ ;
	wire _w2670_ ;
	wire _w2671_ ;
	wire _w2672_ ;
	wire _w2673_ ;
	wire _w2674_ ;
	wire _w2675_ ;
	wire _w2676_ ;
	wire _w2677_ ;
	wire _w2678_ ;
	wire _w2679_ ;
	wire _w2680_ ;
	wire _w2681_ ;
	wire _w2682_ ;
	wire _w2683_ ;
	wire _w2684_ ;
	wire _w2685_ ;
	wire _w2686_ ;
	wire _w2687_ ;
	wire _w2688_ ;
	wire _w2689_ ;
	wire _w2690_ ;
	wire _w2691_ ;
	wire _w2692_ ;
	wire _w2693_ ;
	wire _w2694_ ;
	wire _w2695_ ;
	wire _w2696_ ;
	wire _w2697_ ;
	wire _w2698_ ;
	wire _w2699_ ;
	wire _w2700_ ;
	wire _w2701_ ;
	wire _w2702_ ;
	wire _w2703_ ;
	wire _w2704_ ;
	wire _w2705_ ;
	wire _w2706_ ;
	wire _w2707_ ;
	wire _w2708_ ;
	wire _w2709_ ;
	wire _w2710_ ;
	wire _w2711_ ;
	wire _w2712_ ;
	wire _w2713_ ;
	wire _w2714_ ;
	wire _w2715_ ;
	wire _w2716_ ;
	wire _w2717_ ;
	wire _w2718_ ;
	wire _w2719_ ;
	wire _w2720_ ;
	wire _w2721_ ;
	wire _w2722_ ;
	wire _w2723_ ;
	wire _w2724_ ;
	wire _w2725_ ;
	wire _w2726_ ;
	wire _w2727_ ;
	wire _w2728_ ;
	wire _w2729_ ;
	wire _w2730_ ;
	wire _w2731_ ;
	wire _w2732_ ;
	wire _w2733_ ;
	wire _w2734_ ;
	wire _w2735_ ;
	wire _w2736_ ;
	wire _w2737_ ;
	wire _w2738_ ;
	wire _w2739_ ;
	wire _w2740_ ;
	wire _w2741_ ;
	wire _w2742_ ;
	wire _w2743_ ;
	wire _w2744_ ;
	wire _w2745_ ;
	wire _w2746_ ;
	wire _w2747_ ;
	wire _w2748_ ;
	wire _w2749_ ;
	wire _w2750_ ;
	wire _w2751_ ;
	wire _w2752_ ;
	wire _w2753_ ;
	wire _w2754_ ;
	wire _w2755_ ;
	wire _w2756_ ;
	wire _w2757_ ;
	wire _w2758_ ;
	wire _w2759_ ;
	wire _w2760_ ;
	wire _w2761_ ;
	wire _w2762_ ;
	wire _w2763_ ;
	wire _w2764_ ;
	wire _w2765_ ;
	wire _w2766_ ;
	wire _w2767_ ;
	wire _w2768_ ;
	wire _w2769_ ;
	wire _w2770_ ;
	wire _w2771_ ;
	wire _w2772_ ;
	wire _w2773_ ;
	wire _w2774_ ;
	wire _w2775_ ;
	wire _w2776_ ;
	wire _w2777_ ;
	wire _w2778_ ;
	wire _w2779_ ;
	wire _w2780_ ;
	wire _w2781_ ;
	wire _w2782_ ;
	wire _w2783_ ;
	wire _w2784_ ;
	wire _w2785_ ;
	wire _w2786_ ;
	wire _w2787_ ;
	wire _w2788_ ;
	wire _w2789_ ;
	wire _w2790_ ;
	wire _w2791_ ;
	wire _w2792_ ;
	wire _w2793_ ;
	wire _w2794_ ;
	wire _w2795_ ;
	wire _w2796_ ;
	wire _w2797_ ;
	wire _w2798_ ;
	wire _w2799_ ;
	wire _w2800_ ;
	wire _w2801_ ;
	wire _w2802_ ;
	wire _w2803_ ;
	wire _w2804_ ;
	wire _w2805_ ;
	wire _w2806_ ;
	wire _w2807_ ;
	wire _w2808_ ;
	wire _w2809_ ;
	wire _w2810_ ;
	wire _w2811_ ;
	wire _w2812_ ;
	wire _w2813_ ;
	wire _w2814_ ;
	wire _w2815_ ;
	wire _w2816_ ;
	wire _w2817_ ;
	wire _w2818_ ;
	wire _w2819_ ;
	wire _w2820_ ;
	wire _w2821_ ;
	wire _w2822_ ;
	wire _w2823_ ;
	wire _w2824_ ;
	wire _w2825_ ;
	wire _w2826_ ;
	wire _w2827_ ;
	wire _w2828_ ;
	wire _w2829_ ;
	wire _w2830_ ;
	wire _w2831_ ;
	wire _w2832_ ;
	wire _w2833_ ;
	wire _w2834_ ;
	wire _w2835_ ;
	wire _w2836_ ;
	wire _w2837_ ;
	wire _w2838_ ;
	wire _w2839_ ;
	wire _w2840_ ;
	wire _w2841_ ;
	wire _w2842_ ;
	wire _w2843_ ;
	wire _w2844_ ;
	wire _w2845_ ;
	wire _w2846_ ;
	wire _w2847_ ;
	wire _w2848_ ;
	wire _w2849_ ;
	wire _w2850_ ;
	wire _w2851_ ;
	wire _w2852_ ;
	wire _w2853_ ;
	wire _w2854_ ;
	wire _w2855_ ;
	wire _w2856_ ;
	wire _w2857_ ;
	wire _w2858_ ;
	wire _w4107_ ;
	wire _w4108_ ;
	wire _w4109_ ;
	wire _w4110_ ;
	wire _w4111_ ;
	wire _w4112_ ;
	wire _w4113_ ;
	wire _w4114_ ;
	wire _w4115_ ;
	wire _w4116_ ;
	wire _w4117_ ;
	wire _w4118_ ;
	wire _w4119_ ;
	wire _w4120_ ;
	wire _w4121_ ;
	wire _w4122_ ;
	wire _w4123_ ;
	wire _w4124_ ;
	wire _w4125_ ;
	wire _w4126_ ;
	wire _w4127_ ;
	wire _w4128_ ;
	wire _w4129_ ;
	wire _w4130_ ;
	wire _w4131_ ;
	wire _w4132_ ;
	wire _w4133_ ;
	wire _w4134_ ;
	wire _w4135_ ;
	wire _w4136_ ;
	wire _w4137_ ;
	wire _w4138_ ;
	wire _w4139_ ;
	wire _w4140_ ;
	wire _w4141_ ;
	wire _w4142_ ;
	wire _w4143_ ;
	wire _w4144_ ;
	wire _w4145_ ;
	wire _w4146_ ;
	wire _w4147_ ;
	wire _w4148_ ;
	wire _w4149_ ;
	wire _w4150_ ;
	wire _w4151_ ;
	wire _w4152_ ;
	wire _w4153_ ;
	wire _w4154_ ;
	wire _w4155_ ;
	wire _w4156_ ;
	wire _w4157_ ;
	wire _w4158_ ;
	wire _w4159_ ;
	wire _w4160_ ;
	wire _w4161_ ;
	wire _w4162_ ;
	wire _w4163_ ;
	wire _w4164_ ;
	wire _w4165_ ;
	wire _w4166_ ;
	wire _w4167_ ;
	wire _w4168_ ;
	wire _w4169_ ;
	wire _w4170_ ;
	wire _w4171_ ;
	wire _w4172_ ;
	wire _w4173_ ;
	wire _w4174_ ;
	wire _w4175_ ;
	wire _w4176_ ;
	wire _w4177_ ;
	wire _w4178_ ;
	wire _w4179_ ;
	wire _w4180_ ;
	wire _w4181_ ;
	wire _w4182_ ;
	wire _w4183_ ;
	wire _w4184_ ;
	wire _w4185_ ;
	wire _w4186_ ;
	wire _w4187_ ;
	wire _w4188_ ;
	wire _w4189_ ;
	wire _w4190_ ;
	wire _w4191_ ;
	wire _w4192_ ;
	wire _w4193_ ;
	wire _w4194_ ;
	wire _w4195_ ;
	wire _w4196_ ;
	wire _w4197_ ;
	wire _w4198_ ;
	wire _w4199_ ;
	wire _w4200_ ;
	wire _w4201_ ;
	wire _w4202_ ;
	wire _w4203_ ;
	wire _w4204_ ;
	wire _w4205_ ;
	wire _w4206_ ;
	wire _w4207_ ;
	wire _w4208_ ;
	wire _w4209_ ;
	wire _w4210_ ;
	wire _w4211_ ;
	wire _w4212_ ;
	wire _w4213_ ;
	wire _w4214_ ;
	wire _w4215_ ;
	wire _w4216_ ;
	wire _w4217_ ;
	wire _w4218_ ;
	wire _w4219_ ;
	wire _w4220_ ;
	wire _w4221_ ;
	wire _w4222_ ;
	wire _w4223_ ;
	wire _w4224_ ;
	wire _w4225_ ;
	wire _w4226_ ;
	wire _w4227_ ;
	wire _w4228_ ;
	wire _w4229_ ;
	wire _w4230_ ;
	wire _w4231_ ;
	wire _w4232_ ;
	wire _w4233_ ;
	wire _w4234_ ;
	wire _w4235_ ;
	wire _w4236_ ;
	wire _w4237_ ;
	wire _w4238_ ;
	wire _w4239_ ;
	wire _w4240_ ;
	wire _w4241_ ;
	wire _w4242_ ;
	wire _w4243_ ;
	wire _w4244_ ;
	wire _w4245_ ;
	wire _w4246_ ;
	wire _w4247_ ;
	wire _w4248_ ;
	wire _w4249_ ;
	wire _w4250_ ;
	wire _w4251_ ;
	wire _w4252_ ;
	wire _w4253_ ;
	wire _w4254_ ;
	wire _w4255_ ;
	wire _w4256_ ;
	wire _w4257_ ;
	wire _w4258_ ;
	wire _w4259_ ;
	wire _w4260_ ;
	wire _w4261_ ;
	wire _w4262_ ;
	wire _w4263_ ;
	wire _w4264_ ;
	wire _w4265_ ;
	wire _w4266_ ;
	wire _w4267_ ;
	wire _w4268_ ;
	wire _w4269_ ;
	wire _w4270_ ;
	wire _w4271_ ;
	wire _w4272_ ;
	wire _w4273_ ;
	wire _w4274_ ;
	wire _w4275_ ;
	wire _w4276_ ;
	wire _w4277_ ;
	wire _w4278_ ;
	wire _w4279_ ;
	wire _w4280_ ;
	wire _w4281_ ;
	wire _w4282_ ;
	wire _w4283_ ;
	wire _w4284_ ;
	wire _w4285_ ;
	wire _w4286_ ;
	wire _w4287_ ;
	wire _w4288_ ;
	wire _w4289_ ;
	wire _w4290_ ;
	wire _w4291_ ;
	wire _w4292_ ;
	wire _w4293_ ;
	wire _w4294_ ;
	wire _w4295_ ;
	wire _w4296_ ;
	wire _w4297_ ;
	wire _w4298_ ;
	wire _w4299_ ;
	wire _w4300_ ;
	wire _w4301_ ;
	wire _w4302_ ;
	wire _w4303_ ;
	wire _w4304_ ;
	wire _w4305_ ;
	wire _w4306_ ;
	wire _w4307_ ;
	wire _w4308_ ;
	wire _w4309_ ;
	wire _w4310_ ;
	wire _w4311_ ;
	wire _w4312_ ;
	wire _w4313_ ;
	wire _w4314_ ;
	wire _w4315_ ;
	wire _w4316_ ;
	wire _w4317_ ;
	wire _w4318_ ;
	wire _w4319_ ;
	wire _w4320_ ;
	wire _w4321_ ;
	wire _w4322_ ;
	wire _w4323_ ;
	wire _w4324_ ;
	wire _w4325_ ;
	wire _w4326_ ;
	wire _w4327_ ;
	wire _w4328_ ;
	wire _w4329_ ;
	wire _w4330_ ;
	wire _w4331_ ;
	wire _w4332_ ;
	wire _w4333_ ;
	wire _w4334_ ;
	wire _w4335_ ;
	wire _w4336_ ;
	wire _w4337_ ;
	wire _w4338_ ;
	wire _w4339_ ;
	wire _w4340_ ;
	wire _w4341_ ;
	wire _w4342_ ;
	wire _w4343_ ;
	wire _w4344_ ;
	wire _w4345_ ;
	wire _w4346_ ;
	wire _w4347_ ;
	wire _w4348_ ;
	wire _w4349_ ;
	wire _w4350_ ;
	wire _w4351_ ;
	wire _w4352_ ;
	wire _w4353_ ;
	wire _w4354_ ;
	wire _w4355_ ;
	wire _w4356_ ;
	wire _w4357_ ;
	wire _w4358_ ;
	wire _w4359_ ;
	wire _w4360_ ;
	wire _w4361_ ;
	wire _w4362_ ;
	wire _w4363_ ;
	wire _w4364_ ;
	wire _w4365_ ;
	wire _w4366_ ;
	wire _w4367_ ;
	wire _w4368_ ;
	wire _w4369_ ;
	wire _w4370_ ;
	wire _w4371_ ;
	wire _w4372_ ;
	wire _w4373_ ;
	wire _w4374_ ;
	wire _w4375_ ;
	wire _w4376_ ;
	wire _w4377_ ;
	wire _w4378_ ;
	wire _w4379_ ;
	wire _w4380_ ;
	wire _w4381_ ;
	wire _w4382_ ;
	wire _w4383_ ;
	wire _w4384_ ;
	wire _w4385_ ;
	wire _w4386_ ;
	wire _w4387_ ;
	wire _w4388_ ;
	wire _w4389_ ;
	wire _w4390_ ;
	wire _w4391_ ;
	wire _w4392_ ;
	wire _w4393_ ;
	wire _w4394_ ;
	wire _w4395_ ;
	wire _w4396_ ;
	wire _w4397_ ;
	wire _w4398_ ;
	wire _w4399_ ;
	wire _w4400_ ;
	wire _w4401_ ;
	wire _w4402_ ;
	wire _w4403_ ;
	wire _w4404_ ;
	wire _w4405_ ;
	wire _w4406_ ;
	wire _w4407_ ;
	wire _w4408_ ;
	wire _w4409_ ;
	wire _w4410_ ;
	wire _w4411_ ;
	wire _w4412_ ;
	wire _w4413_ ;
	wire _w4414_ ;
	wire _w4415_ ;
	wire _w4416_ ;
	wire _w4417_ ;
	wire _w4418_ ;
	wire _w4419_ ;
	wire _w4420_ ;
	wire _w4421_ ;
	wire _w4422_ ;
	wire _w4423_ ;
	wire _w4424_ ;
	wire _w4425_ ;
	wire _w4426_ ;
	wire _w4427_ ;
	wire _w4428_ ;
	wire _w4429_ ;
	wire _w4430_ ;
	wire _w4431_ ;
	wire _w4432_ ;
	wire _w4433_ ;
	wire _w4434_ ;
	wire _w4435_ ;
	wire _w4436_ ;
	wire _w4437_ ;
	wire _w4438_ ;
	wire _w4439_ ;
	wire _w4440_ ;
	wire _w4441_ ;
	wire _w4442_ ;
	wire _w4443_ ;
	wire _w4444_ ;
	wire _w4445_ ;
	wire _w4446_ ;
	wire _w4447_ ;
	wire _w4448_ ;
	wire _w4449_ ;
	wire _w4450_ ;
	wire _w4451_ ;
	wire _w4452_ ;
	wire _w4453_ ;
	wire _w4454_ ;
	wire _w4455_ ;
	wire _w4456_ ;
	wire _w4457_ ;
	wire _w4458_ ;
	wire _w4459_ ;
	wire _w4460_ ;
	wire _w4461_ ;
	wire _w4462_ ;
	wire _w4463_ ;
	wire _w4464_ ;
	wire _w4465_ ;
	wire _w4466_ ;
	wire _w4467_ ;
	wire _w4468_ ;
	wire _w4469_ ;
	wire _w4470_ ;
	wire _w4471_ ;
	wire _w4472_ ;
	wire _w4473_ ;
	wire _w4474_ ;
	wire _w4475_ ;
	wire _w4476_ ;
	wire _w4477_ ;
	wire _w4478_ ;
	wire _w4479_ ;
	wire _w4480_ ;
	wire _w4481_ ;
	wire _w4482_ ;
	wire _w4483_ ;
	wire _w4484_ ;
	wire _w4485_ ;
	wire _w4486_ ;
	wire _w4487_ ;
	wire _w4488_ ;
	wire _w4489_ ;
	wire _w4490_ ;
	wire _w4491_ ;
	wire _w4492_ ;
	wire _w4493_ ;
	wire _w4494_ ;
	wire _w4495_ ;
	wire _w4496_ ;
	wire _w4497_ ;
	wire _w4498_ ;
	wire _w4499_ ;
	wire _w4500_ ;
	wire _w4501_ ;
	wire _w4502_ ;
	wire _w4503_ ;
	wire _w4504_ ;
	wire _w4505_ ;
	wire _w4506_ ;
	wire _w4507_ ;
	wire _w4508_ ;
	wire _w4509_ ;
	wire _w4510_ ;
	wire _w4511_ ;
	wire _w4512_ ;
	wire _w4513_ ;
	wire _w4514_ ;
	wire _w4515_ ;
	wire _w4516_ ;
	wire _w4517_ ;
	wire _w4518_ ;
	wire _w4519_ ;
	wire _w4520_ ;
	wire _w4521_ ;
	wire _w4522_ ;
	wire _w4523_ ;
	wire _w4524_ ;
	wire _w4525_ ;
	wire _w4526_ ;
	wire _w4527_ ;
	wire _w4528_ ;
	wire _w4529_ ;
	wire _w4530_ ;
	wire _w4531_ ;
	wire _w4532_ ;
	wire _w4533_ ;
	wire _w4534_ ;
	wire _w4535_ ;
	wire _w4536_ ;
	wire _w4537_ ;
	wire _w4538_ ;
	wire _w4539_ ;
	wire _w4540_ ;
	wire _w4541_ ;
	wire _w4542_ ;
	wire _w4543_ ;
	wire _w4544_ ;
	wire _w4545_ ;
	wire _w4546_ ;
	wire _w4547_ ;
	wire _w4548_ ;
	wire _w4549_ ;
	wire _w4550_ ;
	wire _w4551_ ;
	wire _w4552_ ;
	wire _w4553_ ;
	wire _w4554_ ;
	wire _w4555_ ;
	wire _w4556_ ;
	wire _w4557_ ;
	wire _w4558_ ;
	wire _w4559_ ;
	wire _w4560_ ;
	wire _w4561_ ;
	wire _w4562_ ;
	wire _w4563_ ;
	wire _w4564_ ;
	wire _w4565_ ;
	wire _w4566_ ;
	wire _w4567_ ;
	wire _w4568_ ;
	wire _w4569_ ;
	wire _w4570_ ;
	wire _w4571_ ;
	wire _w4572_ ;
	wire _w4573_ ;
	wire _w4574_ ;
	wire _w4575_ ;
	wire _w4576_ ;
	wire _w4577_ ;
	wire _w4578_ ;
	wire _w4579_ ;
	wire _w4580_ ;
	wire _w4581_ ;
	wire _w4582_ ;
	wire _w4583_ ;
	wire _w4584_ ;
	wire _w4585_ ;
	wire _w4586_ ;
	wire _w4587_ ;
	wire _w4588_ ;
	wire _w4589_ ;
	wire _w4590_ ;
	wire _w4591_ ;
	wire _w4592_ ;
	wire _w4593_ ;
	wire _w4594_ ;
	wire _w4595_ ;
	wire _w4596_ ;
	wire _w4597_ ;
	wire _w4598_ ;
	wire _w4599_ ;
	wire _w4600_ ;
	wire _w4601_ ;
	wire _w4602_ ;
	wire _w4603_ ;
	wire _w4604_ ;
	wire _w4605_ ;
	wire _w4606_ ;
	wire _w4607_ ;
	wire _w4608_ ;
	wire _w4609_ ;
	wire _w4610_ ;
	wire _w4611_ ;
	wire _w4612_ ;
	wire _w4613_ ;
	wire _w4614_ ;
	wire _w4615_ ;
	wire _w4616_ ;
	wire _w4617_ ;
	wire _w4618_ ;
	wire _w4619_ ;
	wire _w4620_ ;
	wire _w4621_ ;
	wire _w4622_ ;
	wire _w4623_ ;
	wire _w4624_ ;
	wire _w4625_ ;
	wire _w4626_ ;
	wire _w4627_ ;
	wire _w4628_ ;
	wire _w4629_ ;
	wire _w4630_ ;
	wire _w4631_ ;
	wire _w4632_ ;
	wire _w4633_ ;
	wire _w4634_ ;
	wire _w4635_ ;
	wire _w4636_ ;
	wire _w4637_ ;
	wire _w4638_ ;
	wire _w4639_ ;
	wire _w4640_ ;
	wire _w4641_ ;
	wire _w4642_ ;
	wire _w4643_ ;
	wire _w4644_ ;
	wire _w4645_ ;
	wire _w4646_ ;
	wire _w4647_ ;
	wire _w4648_ ;
	wire _w4649_ ;
	wire _w4650_ ;
	wire _w4651_ ;
	wire _w4652_ ;
	wire _w4653_ ;
	wire _w4654_ ;
	wire _w4655_ ;
	wire _w4656_ ;
	wire _w4657_ ;
	wire _w4658_ ;
	wire _w4659_ ;
	wire _w4660_ ;
	wire _w4661_ ;
	wire _w4662_ ;
	wire _w4663_ ;
	wire _w4664_ ;
	wire _w4665_ ;
	wire _w4666_ ;
	wire _w4667_ ;
	wire _w4668_ ;
	wire _w4669_ ;
	wire _w4670_ ;
	wire _w4671_ ;
	wire _w4672_ ;
	wire _w4673_ ;
	wire _w4674_ ;
	wire _w4675_ ;
	wire _w4676_ ;
	wire _w4677_ ;
	wire _w4678_ ;
	wire _w4679_ ;
	wire _w4680_ ;
	wire _w4681_ ;
	wire _w4682_ ;
	wire _w4683_ ;
	wire _w4684_ ;
	wire _w4685_ ;
	wire _w4686_ ;
	wire _w4687_ ;
	wire _w4688_ ;
	wire _w4689_ ;
	wire _w4690_ ;
	wire _w4691_ ;
	wire _w4692_ ;
	wire _w4693_ ;
	wire _w4694_ ;
	wire _w4695_ ;
	wire _w4696_ ;
	wire _w4697_ ;
	wire _w4698_ ;
	wire _w4699_ ;
	wire _w4700_ ;
	wire _w4701_ ;
	wire _w4702_ ;
	wire _w4703_ ;
	wire _w4704_ ;
	wire _w4705_ ;
	wire _w4706_ ;
	wire _w4707_ ;
	wire _w4708_ ;
	wire _w4709_ ;
	wire _w4710_ ;
	wire _w4711_ ;
	wire _w4712_ ;
	wire _w4713_ ;
	wire _w4714_ ;
	wire _w4715_ ;
	wire _w4716_ ;
	wire _w4717_ ;
	wire _w4718_ ;
	wire _w4719_ ;
	wire _w4720_ ;
	wire _w4721_ ;
	wire _w4722_ ;
	wire _w4723_ ;
	wire _w4724_ ;
	wire _w4725_ ;
	wire _w4726_ ;
	wire _w4727_ ;
	wire _w4728_ ;
	wire _w4729_ ;
	wire _w4730_ ;
	wire _w4731_ ;
	wire _w4732_ ;
	wire _w4733_ ;
	wire _w4734_ ;
	wire _w4735_ ;
	wire _w4736_ ;
	wire _w4737_ ;
	wire _w4738_ ;
	wire _w4739_ ;
	wire _w4740_ ;
	wire _w4741_ ;
	wire _w4742_ ;
	wire _w4743_ ;
	wire _w4744_ ;
	wire _w4745_ ;
	wire _w4746_ ;
	wire _w4747_ ;
	wire _w4748_ ;
	wire _w4749_ ;
	wire _w4750_ ;
	wire _w4751_ ;
	wire _w4752_ ;
	wire _w4753_ ;
	wire _w4754_ ;
	wire _w4755_ ;
	wire _w4756_ ;
	wire _w4757_ ;
	wire _w4758_ ;
	wire _w4759_ ;
	wire _w4760_ ;
	wire _w4761_ ;
	wire _w4762_ ;
	wire _w4763_ ;
	wire _w4764_ ;
	wire _w4765_ ;
	wire _w4766_ ;
	wire _w4767_ ;
	wire _w4768_ ;
	wire _w4769_ ;
	wire _w4770_ ;
	wire _w4771_ ;
	wire _w4772_ ;
	wire _w4773_ ;
	wire _w4774_ ;
	wire _w4775_ ;
	wire _w4776_ ;
	wire _w4777_ ;
	wire _w4778_ ;
	wire _w4779_ ;
	wire _w4780_ ;
	wire _w4781_ ;
	wire _w4782_ ;
	wire _w4783_ ;
	wire _w4784_ ;
	wire _w4785_ ;
	wire _w4786_ ;
	wire _w4787_ ;
	wire _w4788_ ;
	wire _w4789_ ;
	wire _w4790_ ;
	wire _w4791_ ;
	wire _w4792_ ;
	wire _w4793_ ;
	wire _w4794_ ;
	wire _w4795_ ;
	wire _w4796_ ;
	wire _w4797_ ;
	wire _w4798_ ;
	wire _w4799_ ;
	wire _w4800_ ;
	wire _w4801_ ;
	wire _w4802_ ;
	wire _w4803_ ;
	wire _w4804_ ;
	wire _w4805_ ;
	wire _w4806_ ;
	wire _w4807_ ;
	wire _w4808_ ;
	wire _w4809_ ;
	wire _w4810_ ;
	wire _w4811_ ;
	wire _w4812_ ;
	wire _w4813_ ;
	wire _w4814_ ;
	wire _w4815_ ;
	wire _w4816_ ;
	wire _w4817_ ;
	wire _w4818_ ;
	wire _w4819_ ;
	wire _w4820_ ;
	wire _w4821_ ;
	wire _w4822_ ;
	wire _w4823_ ;
	wire _w4824_ ;
	wire _w4825_ ;
	wire _w4826_ ;
	wire _w4827_ ;
	wire _w4828_ ;
	wire _w4829_ ;
	wire _w4830_ ;
	wire _w4831_ ;
	wire _w4832_ ;
	wire _w4833_ ;
	wire _w4834_ ;
	wire _w4835_ ;
	wire _w4836_ ;
	wire _w4837_ ;
	wire _w4838_ ;
	wire _w4839_ ;
	wire _w4840_ ;
	wire _w4841_ ;
	wire _w4842_ ;
	wire _w4843_ ;
	wire _w4844_ ;
	wire _w4845_ ;
	wire _w4846_ ;
	wire _w4847_ ;
	wire _w4848_ ;
	wire _w4849_ ;
	wire _w4850_ ;
	wire _w4851_ ;
	wire _w4852_ ;
	wire _w4853_ ;
	wire _w4854_ ;
	wire _w4855_ ;
	wire _w4856_ ;
	wire _w4857_ ;
	wire _w4858_ ;
	wire _w4859_ ;
	wire _w4860_ ;
	wire _w4861_ ;
	wire _w4862_ ;
	wire _w4863_ ;
	wire _w4864_ ;
	wire _w4865_ ;
	wire _w4866_ ;
	wire _w4867_ ;
	wire _w4868_ ;
	wire _w4869_ ;
	wire _w4870_ ;
	wire _w4871_ ;
	wire _w4872_ ;
	wire _w4873_ ;
	wire _w4874_ ;
	wire _w4875_ ;
	wire _w4876_ ;
	wire _w4877_ ;
	wire _w4878_ ;
	wire _w4879_ ;
	wire _w4880_ ;
	wire _w4881_ ;
	wire _w4882_ ;
	wire _w4883_ ;
	wire _w4884_ ;
	wire _w4885_ ;
	wire _w4886_ ;
	wire _w4887_ ;
	wire _w4888_ ;
	wire _w4889_ ;
	wire _w4890_ ;
	wire _w4891_ ;
	wire _w4892_ ;
	wire _w4893_ ;
	wire _w4894_ ;
	wire _w4895_ ;
	wire _w4896_ ;
	wire _w4897_ ;
	wire _w4898_ ;
	wire _w4899_ ;
	wire _w4900_ ;
	wire _w4901_ ;
	wire _w4902_ ;
	wire _w4903_ ;
	wire _w4904_ ;
	wire _w4905_ ;
	wire _w4906_ ;
	wire _w4907_ ;
	wire _w4908_ ;
	wire _w4909_ ;
	wire _w4910_ ;
	wire _w4911_ ;
	wire _w4912_ ;
	wire _w4913_ ;
	wire _w4914_ ;
	wire _w4915_ ;
	wire _w4916_ ;
	wire _w4917_ ;
	wire _w4918_ ;
	wire _w4919_ ;
	wire _w4920_ ;
	wire _w4921_ ;
	wire _w4922_ ;
	wire _w4923_ ;
	wire _w4924_ ;
	wire _w4925_ ;
	wire _w4926_ ;
	wire _w4927_ ;
	wire _w4928_ ;
	wire _w4929_ ;
	wire _w4930_ ;
	wire _w4931_ ;
	wire _w4932_ ;
	wire _w4933_ ;
	wire _w4934_ ;
	wire _w4935_ ;
	wire _w4936_ ;
	wire _w4937_ ;
	wire _w4938_ ;
	wire _w4939_ ;
	wire _w4940_ ;
	wire _w4941_ ;
	wire _w4942_ ;
	wire _w4943_ ;
	wire _w4944_ ;
	wire _w4945_ ;
	wire _w4946_ ;
	wire _w4947_ ;
	wire _w4948_ ;
	wire _w4949_ ;
	wire _w4950_ ;
	wire _w4951_ ;
	wire _w4952_ ;
	wire _w4953_ ;
	wire _w4954_ ;
	wire _w4955_ ;
	wire _w4956_ ;
	wire _w4957_ ;
	wire _w4958_ ;
	wire _w4959_ ;
	wire _w4960_ ;
	wire _w4961_ ;
	wire _w4962_ ;
	wire _w4963_ ;
	wire _w4964_ ;
	wire _w4965_ ;
	wire _w4966_ ;
	wire _w4967_ ;
	wire _w4968_ ;
	wire _w4969_ ;
	wire _w4970_ ;
	wire _w4971_ ;
	wire _w4972_ ;
	wire _w4973_ ;
	wire _w4974_ ;
	wire _w4975_ ;
	wire _w4976_ ;
	wire _w4977_ ;
	wire _w4978_ ;
	wire _w4979_ ;
	wire _w4980_ ;
	wire _w4981_ ;
	wire _w4982_ ;
	wire _w4983_ ;
	wire _w4984_ ;
	wire _w4985_ ;
	wire _w4986_ ;
	wire _w4987_ ;
	wire _w4988_ ;
	wire _w4989_ ;
	wire _w4990_ ;
	wire _w4991_ ;
	wire _w4992_ ;
	wire _w4993_ ;
	wire _w4994_ ;
	wire _w4995_ ;
	wire _w4996_ ;
	wire _w4997_ ;
	wire _w4998_ ;
	wire _w4999_ ;
	wire _w5000_ ;
	wire _w5001_ ;
	wire _w5002_ ;
	wire _w5003_ ;
	wire _w5004_ ;
	wire _w5005_ ;
	wire _w5006_ ;
	wire _w5007_ ;
	wire _w5008_ ;
	wire _w5009_ ;
	wire _w5010_ ;
	wire _w5011_ ;
	wire _w5012_ ;
	wire _w5013_ ;
	wire _w5014_ ;
	wire _w5015_ ;
	wire _w5016_ ;
	wire _w5017_ ;
	wire _w5018_ ;
	wire _w5019_ ;
	wire _w5020_ ;
	wire _w5021_ ;
	wire _w5022_ ;
	wire _w5023_ ;
	wire _w5024_ ;
	wire _w5025_ ;
	wire _w5026_ ;
	wire _w5027_ ;
	wire _w5028_ ;
	wire _w5029_ ;
	wire _w5030_ ;
	wire _w5031_ ;
	wire _w5032_ ;
	wire _w5033_ ;
	wire _w5034_ ;
	wire _w5035_ ;
	wire _w5036_ ;
	wire _w5037_ ;
	wire _w5038_ ;
	wire _w5039_ ;
	wire _w5040_ ;
	wire _w5041_ ;
	wire _w5042_ ;
	wire _w5043_ ;
	wire _w5044_ ;
	wire _w5045_ ;
	wire _w5046_ ;
	wire _w5047_ ;
	wire _w5048_ ;
	wire _w5049_ ;
	wire _w5050_ ;
	wire _w5051_ ;
	wire _w5052_ ;
	wire _w5053_ ;
	wire _w5054_ ;
	wire _w5055_ ;
	wire _w5056_ ;
	wire _w5057_ ;
	wire _w5058_ ;
	wire _w5059_ ;
	wire _w5060_ ;
	wire _w5061_ ;
	wire _w5062_ ;
	wire _w5063_ ;
	wire _w5064_ ;
	wire _w5065_ ;
	wire _w5066_ ;
	wire _w5067_ ;
	wire _w5068_ ;
	wire _w5069_ ;
	wire _w5070_ ;
	wire _w5071_ ;
	wire _w5072_ ;
	wire _w5073_ ;
	wire _w5074_ ;
	wire _w5075_ ;
	wire _w5076_ ;
	wire _w5077_ ;
	wire _w5078_ ;
	wire _w5079_ ;
	wire _w5080_ ;
	wire _w5081_ ;
	wire _w5082_ ;
	wire _w5083_ ;
	wire _w5084_ ;
	wire _w5085_ ;
	wire _w5086_ ;
	wire _w5087_ ;
	wire _w5088_ ;
	wire _w5089_ ;
	wire _w5090_ ;
	wire _w5091_ ;
	wire _w5092_ ;
	wire _w5093_ ;
	wire _w5094_ ;
	wire _w5095_ ;
	wire _w5096_ ;
	wire _w5097_ ;
	wire _w5098_ ;
	wire _w5099_ ;
	wire _w5100_ ;
	wire _w5101_ ;
	wire _w5102_ ;
	wire _w5103_ ;
	wire _w5104_ ;
	wire _w5105_ ;
	wire _w5106_ ;
	wire _w5107_ ;
	wire _w5108_ ;
	wire _w5109_ ;
	wire _w5110_ ;
	wire _w5111_ ;
	wire _w5112_ ;
	wire _w5113_ ;
	wire _w5114_ ;
	wire _w5115_ ;
	wire _w5116_ ;
	wire _w5117_ ;
	wire _w5118_ ;
	wire _w5119_ ;
	wire _w5120_ ;
	wire _w5121_ ;
	wire _w5122_ ;
	wire _w5123_ ;
	wire _w5124_ ;
	wire _w5125_ ;
	wire _w5126_ ;
	wire _w5127_ ;
	wire _w5128_ ;
	wire _w5129_ ;
	wire _w5130_ ;
	wire _w5131_ ;
	wire _w5132_ ;
	wire _w5133_ ;
	wire _w5134_ ;
	wire _w5135_ ;
	wire _w5136_ ;
	wire _w5137_ ;
	wire _w5138_ ;
	wire _w5139_ ;
	wire _w5140_ ;
	wire _w5141_ ;
	wire _w5142_ ;
	wire _w5143_ ;
	wire _w5144_ ;
	wire _w5145_ ;
	wire _w5146_ ;
	wire _w5147_ ;
	wire _w5148_ ;
	wire _w5149_ ;
	wire _w5150_ ;
	wire _w5151_ ;
	wire _w5152_ ;
	wire _w5153_ ;
	wire _w5154_ ;
	wire _w5155_ ;
	wire _w5156_ ;
	wire _w5157_ ;
	wire _w5158_ ;
	wire _w5159_ ;
	wire _w5160_ ;
	wire _w5161_ ;
	wire _w5162_ ;
	wire _w5163_ ;
	wire _w5164_ ;
	wire _w5165_ ;
	wire _w5166_ ;
	wire _w5167_ ;
	wire _w5168_ ;
	wire _w5169_ ;
	wire _w5170_ ;
	wire _w5171_ ;
	wire _w5172_ ;
	wire _w5173_ ;
	wire _w5174_ ;
	wire _w5175_ ;
	wire _w5176_ ;
	wire _w5177_ ;
	wire _w5178_ ;
	wire _w5179_ ;
	wire _w5180_ ;
	wire _w5181_ ;
	wire _w5182_ ;
	wire _w5183_ ;
	wire _w5184_ ;
	wire _w5185_ ;
	wire _w5186_ ;
	wire _w5187_ ;
	wire _w5188_ ;
	wire _w5189_ ;
	wire _w5191_ ;
	wire _w5192_ ;
	wire _w5193_ ;
	wire _w5194_ ;
	wire _w5195_ ;
	wire _w5196_ ;
	wire _w5197_ ;
	wire _w5198_ ;
	wire _w5199_ ;
	wire _w5200_ ;
	wire _w5201_ ;
	wire _w5202_ ;
	wire _w5203_ ;
	wire _w5204_ ;
	wire _w5205_ ;
	wire _w5206_ ;
	wire _w5207_ ;
	wire _w5208_ ;
	wire _w5209_ ;
	wire _w5210_ ;
	wire _w5211_ ;
	wire _w5212_ ;
	wire _w5213_ ;
	wire _w5214_ ;
	wire _w5215_ ;
	wire _w5216_ ;
	wire _w5217_ ;
	wire _w5218_ ;
	wire _w5219_ ;
	wire _w5220_ ;
	wire _w5221_ ;
	wire _w5222_ ;
	wire _w5223_ ;
	wire _w5224_ ;
	wire _w5225_ ;
	wire _w5226_ ;
	wire _w5227_ ;
	wire _w5228_ ;
	wire _w5229_ ;
	wire _w5230_ ;
	wire _w5231_ ;
	wire _w5232_ ;
	wire _w5233_ ;
	wire _w5234_ ;
	wire _w5235_ ;
	wire _w5236_ ;
	wire _w5237_ ;
	wire _w5238_ ;
	wire _w5239_ ;
	wire _w5240_ ;
	wire _w5241_ ;
	wire _w5242_ ;
	wire _w5243_ ;
	wire _w5244_ ;
	wire _w5245_ ;
	wire _w5246_ ;
	wire _w5247_ ;
	wire _w5248_ ;
	wire _w5249_ ;
	wire _w5250_ ;
	wire _w5251_ ;
	wire _w5252_ ;
	wire _w5253_ ;
	wire _w5254_ ;
	wire _w5255_ ;
	wire _w5256_ ;
	wire _w5257_ ;
	wire _w5258_ ;
	wire _w5259_ ;
	wire _w5260_ ;
	wire _w5261_ ;
	wire _w5262_ ;
	wire _w5263_ ;
	wire _w5264_ ;
	wire _w5265_ ;
	wire _w5266_ ;
	wire _w5267_ ;
	wire _w5268_ ;
	wire _w5269_ ;
	wire _w5270_ ;
	wire _w5271_ ;
	wire _w5272_ ;
	wire _w5273_ ;
	wire _w5274_ ;
	wire _w5275_ ;
	wire _w5276_ ;
	wire _w5277_ ;
	wire _w5278_ ;
	wire _w5279_ ;
	wire _w5280_ ;
	wire _w5281_ ;
	wire _w5282_ ;
	wire _w5283_ ;
	wire _w5284_ ;
	wire _w5285_ ;
	wire _w5286_ ;
	wire _w5287_ ;
	wire _w5288_ ;
	wire _w5289_ ;
	wire _w5290_ ;
	wire _w5291_ ;
	wire _w5292_ ;
	wire _w5293_ ;
	wire _w5294_ ;
	wire _w5295_ ;
	wire _w5296_ ;
	wire _w5297_ ;
	wire _w5298_ ;
	wire _w5299_ ;
	wire _w5300_ ;
	wire _w5301_ ;
	wire _w5302_ ;
	wire _w5303_ ;
	wire _w5304_ ;
	wire _w5305_ ;
	wire _w5306_ ;
	wire _w5307_ ;
	wire _w5308_ ;
	wire _w5309_ ;
	wire _w5310_ ;
	wire _w5311_ ;
	wire _w5312_ ;
	wire _w5313_ ;
	wire _w5314_ ;
	wire _w5315_ ;
	wire _w5316_ ;
	wire _w5317_ ;
	wire _w5318_ ;
	wire _w5319_ ;
	wire _w5320_ ;
	wire _w5321_ ;
	wire _w5322_ ;
	wire _w5323_ ;
	wire _w5324_ ;
	wire _w5325_ ;
	wire _w5326_ ;
	wire _w5327_ ;
	wire _w5328_ ;
	wire _w5329_ ;
	wire _w5330_ ;
	wire _w5331_ ;
	wire _w5332_ ;
	wire _w5333_ ;
	wire _w5334_ ;
	wire _w5335_ ;
	wire _w5336_ ;
	wire _w5337_ ;
	wire _w5338_ ;
	wire _w5339_ ;
	wire _w5340_ ;
	wire _w5341_ ;
	wire _w5342_ ;
	wire _w5343_ ;
	wire _w5344_ ;
	wire _w5345_ ;
	wire _w5346_ ;
	wire _w5347_ ;
	wire _w5348_ ;
	wire _w5349_ ;
	wire _w5350_ ;
	wire _w5351_ ;
	wire _w5352_ ;
	wire _w5353_ ;
	wire _w5354_ ;
	wire _w5355_ ;
	wire _w5356_ ;
	wire _w5357_ ;
	wire _w5358_ ;
	wire _w5359_ ;
	wire _w5360_ ;
	wire _w5361_ ;
	wire _w5362_ ;
	wire _w5363_ ;
	wire _w5364_ ;
	wire _w5365_ ;
	wire _w5366_ ;
	wire _w5367_ ;
	wire _w5368_ ;
	wire _w5369_ ;
	wire _w5370_ ;
	wire _w5371_ ;
	wire _w5372_ ;
	wire _w5373_ ;
	wire _w5374_ ;
	wire _w5375_ ;
	wire _w5376_ ;
	wire _w5377_ ;
	wire _w5378_ ;
	wire _w5379_ ;
	wire _w5380_ ;
	wire _w5381_ ;
	wire _w5382_ ;
	wire _w5383_ ;
	wire _w5384_ ;
	wire _w5385_ ;
	wire _w5386_ ;
	wire _w5387_ ;
	wire _w5388_ ;
	wire _w5389_ ;
	wire _w5390_ ;
	wire _w5391_ ;
	wire _w5392_ ;
	wire _w5393_ ;
	wire _w5394_ ;
	wire _w5395_ ;
	wire _w5396_ ;
	wire _w5397_ ;
	wire _w5398_ ;
	wire _w5399_ ;
	wire _w5400_ ;
	wire _w5401_ ;
	wire _w5402_ ;
	wire _w5403_ ;
	wire _w5404_ ;
	wire _w5405_ ;
	wire _w5406_ ;
	wire _w5407_ ;
	wire _w5408_ ;
	wire _w5409_ ;
	wire _w5410_ ;
	wire _w5411_ ;
	wire _w5412_ ;
	wire _w5413_ ;
	wire _w5414_ ;
	wire _w5415_ ;
	wire _w5416_ ;
	wire _w5417_ ;
	wire _w5418_ ;
	wire _w5419_ ;
	wire _w5420_ ;
	wire _w5421_ ;
	wire _w5422_ ;
	wire _w5423_ ;
	wire _w5424_ ;
	wire _w5425_ ;
	wire _w5426_ ;
	wire _w5427_ ;
	wire _w5428_ ;
	wire _w5429_ ;
	wire _w5430_ ;
	wire _w5431_ ;
	wire _w5432_ ;
	wire _w5433_ ;
	wire _w5434_ ;
	wire _w5435_ ;
	wire _w5436_ ;
	wire _w5437_ ;
	wire _w5438_ ;
	wire _w5439_ ;
	wire _w5440_ ;
	wire _w5441_ ;
	wire _w5442_ ;
	wire _w5443_ ;
	wire _w5444_ ;
	wire _w5445_ ;
	wire _w5446_ ;
	wire _w5447_ ;
	wire _w5448_ ;
	wire _w5449_ ;
	wire _w5450_ ;
	wire _w5451_ ;
	wire _w5452_ ;
	wire _w5453_ ;
	wire _w5454_ ;
	wire _w5455_ ;
	wire _w5456_ ;
	wire _w5457_ ;
	wire _w5458_ ;
	wire _w5459_ ;
	wire _w5460_ ;
	wire _w5461_ ;
	wire _w5462_ ;
	wire _w5463_ ;
	wire _w5464_ ;
	wire _w5465_ ;
	wire _w5466_ ;
	wire _w5467_ ;
	wire _w5468_ ;
	wire _w5469_ ;
	wire _w5470_ ;
	wire _w5471_ ;
	wire _w5472_ ;
	wire _w5473_ ;
	wire _w5474_ ;
	wire _w5475_ ;
	wire _w5476_ ;
	wire _w5477_ ;
	wire _w5478_ ;
	wire _w5479_ ;
	wire _w5480_ ;
	wire _w5481_ ;
	wire _w5482_ ;
	wire _w5483_ ;
	wire _w5484_ ;
	wire _w5485_ ;
	wire _w5486_ ;
	wire _w5487_ ;
	wire _w5488_ ;
	wire _w5489_ ;
	wire _w5490_ ;
	wire _w5491_ ;
	wire _w5492_ ;
	wire _w5493_ ;
	wire _w5494_ ;
	wire _w5495_ ;
	wire _w5496_ ;
	wire _w5497_ ;
	wire _w5498_ ;
	wire _w5499_ ;
	wire _w5500_ ;
	wire _w5501_ ;
	wire _w5502_ ;
	wire _w5503_ ;
	wire _w5504_ ;
	wire _w5505_ ;
	wire _w5506_ ;
	wire _w5507_ ;
	wire _w5508_ ;
	wire _w5509_ ;
	wire _w5510_ ;
	wire _w5511_ ;
	wire _w5512_ ;
	wire _w5513_ ;
	wire _w5514_ ;
	wire _w5515_ ;
	wire _w5516_ ;
	wire _w5517_ ;
	wire _w5518_ ;
	wire _w5519_ ;
	wire _w5520_ ;
	wire _w5521_ ;
	wire _w5522_ ;
	wire _w5523_ ;
	wire _w5524_ ;
	wire _w5525_ ;
	wire _w5526_ ;
	wire _w5527_ ;
	wire _w5528_ ;
	wire _w5529_ ;
	wire _w5530_ ;
	wire _w5531_ ;
	wire _w5532_ ;
	wire _w5533_ ;
	wire _w5534_ ;
	wire _w5535_ ;
	wire _w5536_ ;
	wire _w5537_ ;
	wire _w5538_ ;
	wire _w5539_ ;
	wire _w5540_ ;
	wire _w5541_ ;
	wire _w5542_ ;
	wire _w5543_ ;
	wire _w5544_ ;
	wire _w5545_ ;
	wire _w5546_ ;
	wire _w5547_ ;
	wire _w5548_ ;
	wire _w5549_ ;
	wire _w5550_ ;
	wire _w5551_ ;
	wire _w5552_ ;
	wire _w5553_ ;
	wire _w5554_ ;
	wire _w5555_ ;
	wire _w5556_ ;
	wire _w5557_ ;
	wire _w5558_ ;
	wire _w5559_ ;
	wire _w5560_ ;
	wire _w5561_ ;
	wire _w5562_ ;
	wire _w5563_ ;
	wire _w5564_ ;
	wire _w5565_ ;
	wire _w5566_ ;
	wire _w5567_ ;
	wire _w5568_ ;
	wire _w5569_ ;
	wire _w5570_ ;
	wire _w5571_ ;
	wire _w5572_ ;
	wire _w5573_ ;
	wire _w5574_ ;
	wire _w5575_ ;
	wire _w5576_ ;
	wire _w5577_ ;
	wire _w5578_ ;
	wire _w5579_ ;
	wire _w5580_ ;
	wire _w5581_ ;
	wire _w5582_ ;
	wire _w5583_ ;
	wire _w5584_ ;
	wire _w5585_ ;
	wire _w5586_ ;
	wire _w5587_ ;
	wire _w5588_ ;
	wire _w5589_ ;
	wire _w5590_ ;
	wire _w5591_ ;
	wire _w5592_ ;
	wire _w5593_ ;
	wire _w5594_ ;
	wire _w5595_ ;
	wire _w5596_ ;
	wire _w5597_ ;
	wire _w5598_ ;
	wire _w5599_ ;
	wire _w5600_ ;
	wire _w5601_ ;
	wire _w5602_ ;
	wire _w5603_ ;
	wire _w5604_ ;
	wire _w5605_ ;
	wire _w5606_ ;
	wire _w5607_ ;
	wire _w5608_ ;
	wire _w5609_ ;
	wire _w5610_ ;
	wire _w5611_ ;
	wire _w5612_ ;
	wire _w5613_ ;
	wire _w5614_ ;
	wire _w5615_ ;
	wire _w5616_ ;
	wire _w5617_ ;
	wire _w5618_ ;
	wire _w5619_ ;
	wire _w5620_ ;
	wire _w5621_ ;
	wire _w5622_ ;
	wire _w5623_ ;
	wire _w5624_ ;
	wire _w5625_ ;
	wire _w5626_ ;
	wire _w5627_ ;
	wire _w5628_ ;
	wire _w5629_ ;
	wire _w5630_ ;
	wire _w5631_ ;
	wire _w5632_ ;
	wire _w5633_ ;
	wire _w5634_ ;
	wire _w5635_ ;
	wire _w5636_ ;
	wire _w5637_ ;
	wire _w5638_ ;
	wire _w5639_ ;
	wire _w5640_ ;
	wire _w5641_ ;
	wire _w5642_ ;
	wire _w5643_ ;
	wire _w5644_ ;
	wire _w5645_ ;
	wire _w5646_ ;
	wire _w5647_ ;
	wire _w5648_ ;
	wire _w5649_ ;
	wire _w5650_ ;
	wire _w5651_ ;
	wire _w5652_ ;
	wire _w5653_ ;
	wire _w5654_ ;
	wire _w5655_ ;
	wire _w5656_ ;
	wire _w5657_ ;
	wire _w5658_ ;
	wire _w5659_ ;
	wire _w5660_ ;
	wire _w5661_ ;
	wire _w5662_ ;
	wire _w5663_ ;
	wire _w5664_ ;
	wire _w5665_ ;
	wire _w5666_ ;
	wire _w5667_ ;
	wire _w5668_ ;
	wire _w5669_ ;
	wire _w5670_ ;
	wire _w5671_ ;
	wire _w5672_ ;
	wire _w5673_ ;
	wire _w5674_ ;
	wire _w5675_ ;
	wire _w5676_ ;
	wire _w5677_ ;
	wire _w5678_ ;
	wire _w5679_ ;
	wire _w5680_ ;
	wire _w5681_ ;
	wire _w5682_ ;
	wire _w5683_ ;
	wire _w5684_ ;
	wire _w5685_ ;
	wire _w5686_ ;
	wire _w5687_ ;
	wire _w5688_ ;
	wire _w5689_ ;
	wire _w5690_ ;
	wire _w5691_ ;
	wire _w5692_ ;
	wire _w5693_ ;
	wire _w5694_ ;
	wire _w5695_ ;
	wire _w5696_ ;
	wire _w5697_ ;
	wire _w5698_ ;
	wire _w5699_ ;
	wire _w5700_ ;
	wire _w5701_ ;
	wire _w5702_ ;
	wire _w5703_ ;
	wire _w5704_ ;
	wire _w5705_ ;
	wire _w5706_ ;
	wire _w5707_ ;
	wire _w5708_ ;
	wire _w5709_ ;
	wire _w5710_ ;
	wire _w5711_ ;
	wire _w5712_ ;
	wire _w5713_ ;
	wire _w5714_ ;
	wire _w5715_ ;
	wire _w5716_ ;
	wire _w5717_ ;
	wire _w5718_ ;
	wire _w5719_ ;
	wire _w5720_ ;
	wire _w5721_ ;
	wire _w5722_ ;
	wire _w5723_ ;
	wire _w5724_ ;
	wire _w5725_ ;
	wire _w5726_ ;
	wire _w5727_ ;
	wire _w5728_ ;
	wire _w5729_ ;
	wire _w5730_ ;
	wire _w5731_ ;
	wire _w5732_ ;
	wire _w5733_ ;
	wire _w5734_ ;
	wire _w5735_ ;
	wire _w5736_ ;
	wire _w5737_ ;
	wire _w5738_ ;
	wire _w5739_ ;
	wire _w5740_ ;
	wire _w5741_ ;
	wire _w5742_ ;
	wire _w5743_ ;
	wire _w5744_ ;
	wire _w5745_ ;
	wire _w5746_ ;
	wire _w5747_ ;
	wire _w5748_ ;
	wire _w5749_ ;
	wire _w5750_ ;
	wire _w5751_ ;
	wire _w5752_ ;
	wire _w5753_ ;
	wire _w5754_ ;
	wire _w5755_ ;
	wire _w5756_ ;
	wire _w5757_ ;
	wire _w5758_ ;
	wire _w5759_ ;
	wire _w5760_ ;
	wire _w5761_ ;
	wire _w5762_ ;
	wire _w5763_ ;
	wire _w5764_ ;
	wire _w5765_ ;
	wire _w5766_ ;
	wire _w5767_ ;
	wire _w5768_ ;
	wire _w5769_ ;
	wire _w5770_ ;
	wire _w5771_ ;
	wire _w5772_ ;
	wire _w5773_ ;
	wire _w5774_ ;
	wire _w5775_ ;
	wire _w5776_ ;
	wire _w5777_ ;
	wire _w5778_ ;
	wire _w5779_ ;
	wire _w5780_ ;
	wire _w5781_ ;
	wire _w5782_ ;
	wire _w5783_ ;
	wire _w5784_ ;
	wire _w5785_ ;
	wire _w5786_ ;
	wire _w5787_ ;
	wire _w5788_ ;
	wire _w5789_ ;
	wire _w5790_ ;
	wire _w5791_ ;
	wire _w5792_ ;
	wire _w5793_ ;
	wire _w5794_ ;
	wire _w5795_ ;
	wire _w5796_ ;
	wire _w5797_ ;
	wire _w5798_ ;
	wire _w5799_ ;
	wire _w5800_ ;
	wire _w5801_ ;
	wire _w5802_ ;
	wire _w5803_ ;
	wire _w5804_ ;
	wire _w5805_ ;
	wire _w5806_ ;
	wire _w5807_ ;
	wire _w5808_ ;
	wire _w5809_ ;
	wire _w5810_ ;
	wire _w5811_ ;
	wire _w5812_ ;
	wire _w5813_ ;
	wire _w5814_ ;
	wire _w5815_ ;
	wire _w5816_ ;
	wire _w5817_ ;
	wire _w5818_ ;
	wire _w5819_ ;
	wire _w5820_ ;
	wire _w5821_ ;
	wire _w5822_ ;
	wire _w5823_ ;
	wire _w5824_ ;
	wire _w5825_ ;
	wire _w5826_ ;
	wire _w5827_ ;
	wire _w5828_ ;
	wire _w5829_ ;
	wire _w5830_ ;
	wire _w5831_ ;
	wire _w5832_ ;
	wire _w5833_ ;
	wire _w5834_ ;
	wire _w5835_ ;
	wire _w5836_ ;
	wire _w5837_ ;
	wire _w5838_ ;
	wire _w5839_ ;
	wire _w5840_ ;
	wire _w5841_ ;
	wire _w5842_ ;
	wire _w5843_ ;
	wire _w5844_ ;
	wire _w5845_ ;
	wire _w5846_ ;
	wire _w5847_ ;
	wire _w5848_ ;
	wire _w5849_ ;
	wire _w5850_ ;
	wire _w5851_ ;
	wire _w5852_ ;
	wire _w5853_ ;
	wire _w5854_ ;
	wire _w5855_ ;
	wire _w5856_ ;
	wire _w5857_ ;
	wire _w5858_ ;
	wire _w5859_ ;
	wire _w5860_ ;
	wire _w5861_ ;
	wire _w5862_ ;
	wire _w5863_ ;
	wire _w5864_ ;
	wire _w5865_ ;
	wire _w5866_ ;
	wire _w5867_ ;
	wire _w5868_ ;
	wire _w5869_ ;
	wire _w5870_ ;
	wire _w5871_ ;
	wire _w5872_ ;
	wire _w5873_ ;
	wire _w5874_ ;
	wire _w5875_ ;
	wire _w5876_ ;
	wire _w5877_ ;
	wire _w5878_ ;
	wire _w5879_ ;
	wire _w5880_ ;
	wire _w5881_ ;
	wire _w5882_ ;
	wire _w5883_ ;
	wire _w5884_ ;
	wire _w5885_ ;
	wire _w5886_ ;
	wire _w5887_ ;
	wire _w5888_ ;
	wire _w5889_ ;
	wire _w5890_ ;
	wire _w5891_ ;
	wire _w5892_ ;
	wire _w5893_ ;
	wire _w5894_ ;
	wire _w5895_ ;
	wire _w5896_ ;
	wire _w5897_ ;
	wire _w5898_ ;
	wire _w5899_ ;
	wire _w5900_ ;
	wire _w5901_ ;
	wire _w5902_ ;
	wire _w5903_ ;
	wire _w5904_ ;
	wire _w5905_ ;
	wire _w5906_ ;
	wire _w5907_ ;
	wire _w5908_ ;
	wire _w5909_ ;
	wire _w5910_ ;
	wire _w5911_ ;
	wire _w5912_ ;
	wire _w5913_ ;
	wire _w5914_ ;
	wire _w5915_ ;
	wire _w5916_ ;
	wire _w5917_ ;
	wire _w5918_ ;
	wire _w5919_ ;
	wire _w5920_ ;
	wire _w5921_ ;
	wire _w5922_ ;
	wire _w5923_ ;
	wire _w5924_ ;
	wire _w5925_ ;
	wire _w5926_ ;
	wire _w5927_ ;
	wire _w5928_ ;
	wire _w5929_ ;
	wire _w5930_ ;
	wire _w5931_ ;
	wire _w5932_ ;
	wire _w5933_ ;
	wire _w5934_ ;
	wire _w5935_ ;
	wire _w5936_ ;
	wire _w5937_ ;
	wire _w5938_ ;
	wire _w5939_ ;
	wire _w5940_ ;
	wire _w5941_ ;
	wire _w5942_ ;
	wire _w5943_ ;
	wire _w5944_ ;
	wire _w5945_ ;
	wire _w5946_ ;
	wire _w5947_ ;
	wire _w5948_ ;
	wire _w5950_ ;
	wire _w5951_ ;
	wire _w5952_ ;
	wire _w5953_ ;
	wire _w5954_ ;
	wire _w5955_ ;
	wire _w5956_ ;
	wire _w5957_ ;
	wire _w5958_ ;
	wire _w5959_ ;
	wire _w5960_ ;
	wire _w5961_ ;
	wire _w5962_ ;
	wire _w5963_ ;
	wire _w5964_ ;
	wire _w5965_ ;
	wire _w5966_ ;
	wire _w5967_ ;
	wire _w5968_ ;
	wire _w5969_ ;
	wire _w5970_ ;
	wire _w5971_ ;
	wire _w5972_ ;
	wire _w5973_ ;
	wire _w5974_ ;
	wire _w5975_ ;
	wire _w5976_ ;
	wire _w5977_ ;
	wire _w5978_ ;
	wire _w5979_ ;
	wire _w5980_ ;
	wire _w5981_ ;
	wire _w5982_ ;
	wire _w5983_ ;
	wire _w5984_ ;
	wire _w5985_ ;
	wire _w5986_ ;
	wire _w5987_ ;
	wire _w5988_ ;
	wire _w5989_ ;
	wire _w5990_ ;
	wire _w5991_ ;
	wire _w5992_ ;
	wire _w5993_ ;
	wire _w5994_ ;
	wire _w5995_ ;
	wire _w5996_ ;
	wire _w5997_ ;
	wire _w5998_ ;
	wire _w5999_ ;
	wire _w6000_ ;
	wire _w6001_ ;
	wire _w6002_ ;
	wire _w6003_ ;
	wire _w6004_ ;
	wire _w6005_ ;
	wire _w6006_ ;
	wire _w6007_ ;
	wire _w6008_ ;
	wire _w6009_ ;
	wire _w6010_ ;
	wire _w6011_ ;
	wire _w6012_ ;
	wire _w6013_ ;
	wire _w6014_ ;
	wire _w6015_ ;
	wire _w6016_ ;
	wire _w6017_ ;
	wire _w6018_ ;
	wire _w6019_ ;
	wire _w6020_ ;
	wire _w6021_ ;
	wire _w6022_ ;
	wire _w6023_ ;
	wire _w6024_ ;
	wire _w6025_ ;
	wire _w6026_ ;
	wire _w6027_ ;
	wire _w6028_ ;
	wire _w6029_ ;
	wire _w6030_ ;
	wire _w6031_ ;
	wire _w6032_ ;
	wire _w6033_ ;
	wire _w6034_ ;
	wire _w6035_ ;
	wire _w6036_ ;
	wire _w6037_ ;
	wire _w6038_ ;
	wire _w6039_ ;
	wire _w6040_ ;
	wire _w6041_ ;
	wire _w6042_ ;
	wire _w6043_ ;
	wire _w6044_ ;
	wire _w6045_ ;
	wire _w6046_ ;
	wire _w6047_ ;
	wire _w6048_ ;
	wire _w6049_ ;
	wire _w6050_ ;
	wire _w6051_ ;
	wire _w6052_ ;
	wire _w6053_ ;
	wire _w6054_ ;
	wire _w6055_ ;
	wire _w6056_ ;
	wire _w6057_ ;
	wire _w6058_ ;
	wire _w6059_ ;
	wire _w6060_ ;
	wire _w6061_ ;
	wire _w6062_ ;
	wire _w6063_ ;
	wire _w6064_ ;
	wire _w6065_ ;
	wire _w6066_ ;
	wire _w6067_ ;
	wire _w6068_ ;
	wire _w6069_ ;
	wire _w6070_ ;
	wire _w6071_ ;
	wire _w6072_ ;
	wire _w6073_ ;
	wire _w6074_ ;
	wire _w6075_ ;
	wire _w6076_ ;
	wire _w6077_ ;
	wire _w6078_ ;
	wire _w6079_ ;
	wire _w6080_ ;
	wire _w6081_ ;
	wire _w6082_ ;
	wire _w6083_ ;
	wire _w6084_ ;
	wire _w6085_ ;
	wire _w6086_ ;
	wire _w6087_ ;
	wire _w6088_ ;
	wire _w6089_ ;
	wire _w6090_ ;
	wire _w6091_ ;
	wire _w6092_ ;
	wire _w6093_ ;
	wire _w6094_ ;
	wire _w6095_ ;
	wire _w6096_ ;
	wire _w6097_ ;
	wire _w6098_ ;
	wire _w6099_ ;
	wire _w6100_ ;
	wire _w6101_ ;
	wire _w6102_ ;
	wire _w6103_ ;
	wire _w6104_ ;
	wire _w6105_ ;
	wire _w6106_ ;
	wire _w6107_ ;
	wire _w6108_ ;
	wire _w6109_ ;
	wire _w6110_ ;
	wire _w6111_ ;
	wire _w6112_ ;
	wire _w6113_ ;
	wire _w6114_ ;
	wire _w6115_ ;
	wire _w6116_ ;
	wire _w6117_ ;
	wire _w6118_ ;
	wire _w6119_ ;
	wire _w6120_ ;
	wire _w6121_ ;
	wire _w6122_ ;
	wire _w6123_ ;
	wire _w6124_ ;
	wire _w6125_ ;
	wire _w6126_ ;
	wire _w6127_ ;
	wire _w6128_ ;
	wire _w6129_ ;
	wire _w6130_ ;
	wire _w6131_ ;
	wire _w6132_ ;
	wire _w6133_ ;
	wire _w6134_ ;
	wire _w6135_ ;
	wire _w6136_ ;
	wire _w6137_ ;
	wire _w6138_ ;
	wire _w6139_ ;
	wire _w6140_ ;
	wire _w6141_ ;
	wire _w6142_ ;
	wire _w6143_ ;
	wire _w6144_ ;
	wire _w6145_ ;
	wire _w6146_ ;
	wire _w6147_ ;
	wire _w6148_ ;
	wire _w6149_ ;
	wire _w6150_ ;
	wire _w6151_ ;
	wire _w6152_ ;
	wire _w6153_ ;
	wire _w6154_ ;
	wire _w6155_ ;
	wire _w6156_ ;
	wire _w6157_ ;
	wire _w6158_ ;
	wire _w6160_ ;
	wire _w6161_ ;
	wire _w6162_ ;
	wire _w6163_ ;
	wire _w6164_ ;
	wire _w6165_ ;
	wire _w6166_ ;
	wire _w6167_ ;
	wire _w6168_ ;
	wire _w6169_ ;
	wire _w6170_ ;
	wire _w6171_ ;
	wire _w6172_ ;
	wire _w6173_ ;
	wire _w6174_ ;
	wire _w6175_ ;
	wire _w6176_ ;
	wire _w6177_ ;
	wire _w6178_ ;
	wire _w6179_ ;
	wire _w6180_ ;
	wire _w6181_ ;
	wire _w6182_ ;
	wire _w6183_ ;
	wire _w6184_ ;
	wire _w6185_ ;
	wire _w6186_ ;
	wire _w6187_ ;
	wire _w6188_ ;
	wire _w6189_ ;
	wire _w6190_ ;
	wire _w6191_ ;
	wire _w6192_ ;
	wire _w6193_ ;
	wire _w6194_ ;
	wire _w6195_ ;
	wire _w6196_ ;
	wire _w6197_ ;
	wire _w6198_ ;
	wire _w6199_ ;
	wire _w6200_ ;
	wire _w6201_ ;
	wire _w6202_ ;
	wire _w6203_ ;
	wire _w6204_ ;
	wire _w6205_ ;
	wire _w6206_ ;
	wire _w6207_ ;
	wire _w6208_ ;
	wire _w6209_ ;
	wire _w6210_ ;
	wire _w6211_ ;
	wire _w6212_ ;
	wire _w6213_ ;
	wire _w6214_ ;
	wire _w6215_ ;
	wire _w6216_ ;
	wire _w6217_ ;
	wire _w6218_ ;
	wire _w6219_ ;
	wire _w6220_ ;
	wire _w6221_ ;
	wire _w6222_ ;
	wire _w6223_ ;
	wire _w6224_ ;
	wire _w6225_ ;
	wire _w6226_ ;
	wire _w6227_ ;
	wire _w6228_ ;
	wire _w6229_ ;
	wire _w6230_ ;
	wire _w6231_ ;
	wire _w6232_ ;
	wire _w6233_ ;
	wire _w6234_ ;
	wire _w6235_ ;
	wire _w6236_ ;
	wire _w6237_ ;
	wire _w6238_ ;
	wire _w6239_ ;
	wire _w6240_ ;
	wire _w6241_ ;
	wire _w6242_ ;
	wire _w6243_ ;
	wire _w6244_ ;
	wire _w6245_ ;
	wire _w6246_ ;
	wire _w6247_ ;
	wire _w6248_ ;
	wire _w6249_ ;
	wire _w6250_ ;
	wire _w6251_ ;
	wire _w6252_ ;
	wire _w6253_ ;
	wire _w6254_ ;
	wire _w6255_ ;
	wire _w6256_ ;
	wire _w6257_ ;
	wire _w6258_ ;
	wire _w6259_ ;
	wire _w6260_ ;
	wire _w6261_ ;
	wire _w6262_ ;
	wire _w6263_ ;
	wire _w6264_ ;
	wire _w6265_ ;
	wire _w6266_ ;
	wire _w6267_ ;
	wire _w6268_ ;
	wire _w6269_ ;
	wire _w6270_ ;
	wire _w6271_ ;
	wire _w6272_ ;
	wire _w6273_ ;
	wire _w6274_ ;
	wire _w6275_ ;
	wire _w6276_ ;
	wire _w6277_ ;
	wire _w6278_ ;
	wire _w6279_ ;
	wire _w6280_ ;
	wire _w6281_ ;
	wire _w6282_ ;
	wire _w6283_ ;
	wire _w6284_ ;
	wire _w6285_ ;
	wire _w6286_ ;
	wire _w6287_ ;
	wire _w6288_ ;
	wire _w6289_ ;
	wire _w6290_ ;
	wire _w6291_ ;
	wire _w6292_ ;
	wire _w6293_ ;
	wire _w6294_ ;
	wire _w6295_ ;
	wire _w6296_ ;
	wire _w6297_ ;
	wire _w6298_ ;
	wire _w6299_ ;
	wire _w6300_ ;
	wire _w6301_ ;
	wire _w6302_ ;
	wire _w6303_ ;
	wire _w6304_ ;
	wire _w6305_ ;
	wire _w6306_ ;
	wire _w6307_ ;
	wire _w6308_ ;
	wire _w6309_ ;
	wire _w6310_ ;
	wire _w6311_ ;
	wire _w6312_ ;
	wire _w6313_ ;
	wire _w6314_ ;
	wire _w6315_ ;
	wire _w6316_ ;
	wire _w6317_ ;
	wire _w6318_ ;
	wire _w6319_ ;
	wire _w6320_ ;
	wire _w6321_ ;
	wire _w6322_ ;
	wire _w6323_ ;
	wire _w6324_ ;
	wire _w6325_ ;
	wire _w6326_ ;
	wire _w6327_ ;
	wire _w6328_ ;
	wire _w6329_ ;
	wire _w6330_ ;
	wire _w6331_ ;
	wire _w6332_ ;
	wire _w6333_ ;
	wire _w6334_ ;
	wire _w6335_ ;
	wire _w6336_ ;
	wire _w6337_ ;
	wire _w6338_ ;
	wire _w6339_ ;
	wire _w6340_ ;
	wire _w6341_ ;
	wire _w6342_ ;
	wire _w6343_ ;
	wire _w6344_ ;
	wire _w6345_ ;
	wire _w6346_ ;
	wire _w6347_ ;
	wire _w6348_ ;
	wire _w6349_ ;
	wire _w6350_ ;
	wire _w6351_ ;
	wire _w6352_ ;
	wire _w6353_ ;
	wire _w6354_ ;
	wire _w6355_ ;
	wire _w6356_ ;
	wire _w6357_ ;
	wire _w6358_ ;
	wire _w6359_ ;
	wire _w6360_ ;
	wire _w6361_ ;
	wire _w6362_ ;
	wire _w6363_ ;
	wire _w6364_ ;
	wire _w6365_ ;
	wire _w6366_ ;
	wire _w6367_ ;
	wire _w6368_ ;
	wire _w6370_ ;
	wire _w6371_ ;
	wire _w6372_ ;
	wire _w6373_ ;
	wire _w6374_ ;
	wire _w6375_ ;
	wire _w6376_ ;
	wire _w6377_ ;
	wire _w6378_ ;
	wire _w6379_ ;
	wire _w6380_ ;
	wire _w6381_ ;
	wire _w6382_ ;
	wire _w6383_ ;
	wire _w6384_ ;
	wire _w6385_ ;
	wire _w6386_ ;
	wire _w6387_ ;
	wire _w6388_ ;
	wire _w6389_ ;
	wire _w6390_ ;
	wire _w6391_ ;
	wire _w6392_ ;
	wire _w6393_ ;
	wire _w6394_ ;
	wire _w6395_ ;
	wire _w6396_ ;
	wire _w6397_ ;
	wire _w6398_ ;
	wire _w6399_ ;
	wire _w6400_ ;
	wire _w6401_ ;
	wire _w6402_ ;
	wire _w6403_ ;
	wire _w6404_ ;
	wire _w6405_ ;
	wire _w6406_ ;
	wire _w6407_ ;
	wire _w6408_ ;
	wire _w6409_ ;
	wire _w6410_ ;
	wire _w6411_ ;
	wire _w6412_ ;
	wire _w6413_ ;
	wire _w6414_ ;
	wire _w6415_ ;
	wire _w6416_ ;
	wire _w6417_ ;
	wire _w6418_ ;
	wire _w6419_ ;
	wire _w6420_ ;
	wire _w6421_ ;
	wire _w6422_ ;
	wire _w6423_ ;
	wire _w6424_ ;
	wire _w6425_ ;
	wire _w6426_ ;
	wire _w6427_ ;
	wire _w6428_ ;
	wire _w6429_ ;
	wire _w6430_ ;
	wire _w6431_ ;
	wire _w6432_ ;
	wire _w6433_ ;
	wire _w6434_ ;
	wire _w6435_ ;
	wire _w6436_ ;
	wire _w6437_ ;
	wire _w6438_ ;
	wire _w6439_ ;
	wire _w6440_ ;
	wire _w6441_ ;
	wire _w6442_ ;
	wire _w6443_ ;
	wire _w6444_ ;
	wire _w6445_ ;
	wire _w6446_ ;
	wire _w6447_ ;
	wire _w6448_ ;
	wire _w6449_ ;
	wire _w6450_ ;
	wire _w6451_ ;
	wire _w6452_ ;
	wire _w6453_ ;
	wire _w6454_ ;
	wire _w6455_ ;
	wire _w6456_ ;
	wire _w6457_ ;
	wire _w6458_ ;
	wire _w6459_ ;
	wire _w6460_ ;
	wire _w6461_ ;
	wire _w6462_ ;
	wire _w6463_ ;
	wire _w6464_ ;
	wire _w6465_ ;
	wire _w6466_ ;
	wire _w6467_ ;
	wire _w6468_ ;
	wire _w6469_ ;
	wire _w6470_ ;
	wire _w6471_ ;
	wire _w6472_ ;
	wire _w6473_ ;
	wire _w6474_ ;
	wire _w6475_ ;
	wire _w6476_ ;
	wire _w6477_ ;
	wire _w6478_ ;
	wire _w6479_ ;
	wire _w6480_ ;
	wire _w6481_ ;
	wire _w6482_ ;
	wire _w6483_ ;
	wire _w6484_ ;
	wire _w6485_ ;
	wire _w6486_ ;
	wire _w6487_ ;
	wire _w6488_ ;
	wire _w6489_ ;
	wire _w6490_ ;
	wire _w6491_ ;
	wire _w6492_ ;
	wire _w6493_ ;
	wire _w6494_ ;
	wire _w6495_ ;
	wire _w6496_ ;
	wire _w6497_ ;
	wire _w6498_ ;
	wire _w6499_ ;
	wire _w6500_ ;
	wire _w6501_ ;
	wire _w6502_ ;
	wire _w6503_ ;
	wire _w6504_ ;
	wire _w6505_ ;
	wire _w6506_ ;
	wire _w6507_ ;
	wire _w6508_ ;
	wire _w6509_ ;
	wire _w6510_ ;
	wire _w6511_ ;
	wire _w6512_ ;
	wire _w6513_ ;
	wire _w6514_ ;
	wire _w6515_ ;
	wire _w6516_ ;
	wire _w6517_ ;
	wire _w6518_ ;
	wire _w6519_ ;
	wire _w6520_ ;
	wire _w6521_ ;
	wire _w6522_ ;
	wire _w6523_ ;
	wire _w6524_ ;
	wire _w6525_ ;
	wire _w6526_ ;
	wire _w6527_ ;
	wire _w6528_ ;
	wire _w6529_ ;
	wire _w6530_ ;
	wire _w6531_ ;
	wire _w6532_ ;
	wire _w6533_ ;
	wire _w6534_ ;
	wire _w6535_ ;
	wire _w6536_ ;
	wire _w6537_ ;
	wire _w6538_ ;
	wire _w6539_ ;
	wire _w6540_ ;
	wire _w6541_ ;
	wire _w6542_ ;
	wire _w6543_ ;
	wire _w6544_ ;
	wire _w6545_ ;
	wire _w6546_ ;
	wire _w6547_ ;
	wire _w6548_ ;
	wire _w6549_ ;
	wire _w6550_ ;
	wire _w6551_ ;
	wire _w6552_ ;
	wire _w6553_ ;
	wire _w6554_ ;
	wire _w6555_ ;
	wire _w6556_ ;
	wire _w6557_ ;
	wire _w6558_ ;
	wire _w6559_ ;
	wire _w6560_ ;
	wire _w6561_ ;
	wire _w6562_ ;
	wire _w6563_ ;
	wire _w6564_ ;
	wire _w6565_ ;
	wire _w6566_ ;
	wire _w6567_ ;
	wire _w6568_ ;
	wire _w6569_ ;
	wire _w6570_ ;
	wire _w6571_ ;
	wire _w6572_ ;
	wire _w6573_ ;
	wire _w6574_ ;
	wire _w6575_ ;
	wire _w6576_ ;
	wire _w6577_ ;
	wire _w6578_ ;
	wire _w6580_ ;
	wire _w6581_ ;
	wire _w6582_ ;
	wire _w6583_ ;
	wire _w6584_ ;
	wire _w6585_ ;
	wire _w6586_ ;
	wire _w6587_ ;
	wire _w6588_ ;
	wire _w6589_ ;
	wire _w6590_ ;
	wire _w6591_ ;
	wire _w6592_ ;
	wire _w6593_ ;
	wire _w6594_ ;
	wire _w6595_ ;
	wire _w6596_ ;
	wire _w6597_ ;
	wire _w6598_ ;
	wire _w6599_ ;
	wire _w6600_ ;
	wire _w6601_ ;
	wire _w6602_ ;
	wire _w6603_ ;
	wire _w6604_ ;
	wire _w6605_ ;
	wire _w6606_ ;
	wire _w6607_ ;
	wire _w6608_ ;
	wire _w6609_ ;
	wire _w6610_ ;
	wire _w6611_ ;
	wire _w6612_ ;
	wire _w6613_ ;
	wire _w6614_ ;
	wire _w6615_ ;
	wire _w6616_ ;
	wire _w6617_ ;
	wire _w6618_ ;
	wire _w6619_ ;
	wire _w6620_ ;
	wire _w6621_ ;
	wire _w6622_ ;
	wire _w6623_ ;
	wire _w6624_ ;
	wire _w6625_ ;
	wire _w6626_ ;
	wire _w6627_ ;
	wire _w6628_ ;
	wire _w6629_ ;
	wire _w6630_ ;
	wire _w6631_ ;
	wire _w6632_ ;
	wire _w6633_ ;
	wire _w6634_ ;
	wire _w6635_ ;
	wire _w6636_ ;
	wire _w6637_ ;
	wire _w6638_ ;
	wire _w6639_ ;
	wire _w6640_ ;
	wire _w6641_ ;
	wire _w6642_ ;
	wire _w6643_ ;
	wire _w6644_ ;
	wire _w6645_ ;
	wire _w6646_ ;
	wire _w6647_ ;
	wire _w6648_ ;
	wire _w6649_ ;
	wire _w6650_ ;
	wire _w6651_ ;
	wire _w6652_ ;
	wire _w6653_ ;
	wire _w6654_ ;
	wire _w6655_ ;
	wire _w6656_ ;
	wire _w6657_ ;
	wire _w6658_ ;
	wire _w6659_ ;
	wire _w6660_ ;
	wire _w6661_ ;
	wire _w6662_ ;
	wire _w6663_ ;
	wire _w6664_ ;
	wire _w6665_ ;
	wire _w6666_ ;
	wire _w6667_ ;
	wire _w6668_ ;
	wire _w6669_ ;
	wire _w6670_ ;
	wire _w6671_ ;
	wire _w6672_ ;
	wire _w6673_ ;
	wire _w6674_ ;
	wire _w6675_ ;
	wire _w6676_ ;
	wire _w6677_ ;
	wire _w6678_ ;
	wire _w6679_ ;
	wire _w6680_ ;
	wire _w6681_ ;
	wire _w6682_ ;
	wire _w6683_ ;
	wire _w6684_ ;
	wire _w6685_ ;
	wire _w6686_ ;
	wire _w6687_ ;
	wire _w6688_ ;
	wire _w6689_ ;
	wire _w6690_ ;
	wire _w6691_ ;
	wire _w6692_ ;
	wire _w6693_ ;
	wire _w6694_ ;
	wire _w6695_ ;
	wire _w6696_ ;
	wire _w6697_ ;
	wire _w6698_ ;
	wire _w6699_ ;
	wire _w6700_ ;
	wire _w6701_ ;
	wire _w6702_ ;
	wire _w6703_ ;
	wire _w6704_ ;
	wire _w6705_ ;
	wire _w6706_ ;
	wire _w6707_ ;
	wire _w6708_ ;
	wire _w6709_ ;
	wire _w6710_ ;
	wire _w6711_ ;
	wire _w6712_ ;
	wire _w6713_ ;
	wire _w6714_ ;
	wire _w6715_ ;
	wire _w6716_ ;
	wire _w6717_ ;
	wire _w6718_ ;
	wire _w6719_ ;
	wire _w6720_ ;
	wire _w6721_ ;
	wire _w6722_ ;
	wire _w6723_ ;
	wire _w6724_ ;
	wire _w6725_ ;
	wire _w6726_ ;
	wire _w6727_ ;
	wire _w6728_ ;
	wire _w6729_ ;
	wire _w6730_ ;
	wire _w6731_ ;
	wire _w6732_ ;
	wire _w6733_ ;
	wire _w6734_ ;
	wire _w6735_ ;
	wire _w6736_ ;
	wire _w6737_ ;
	wire _w6738_ ;
	wire _w6739_ ;
	wire _w6740_ ;
	wire _w6741_ ;
	wire _w6742_ ;
	wire _w6743_ ;
	wire _w6744_ ;
	wire _w6745_ ;
	wire _w6746_ ;
	wire _w6747_ ;
	wire _w6748_ ;
	wire _w6749_ ;
	wire _w6750_ ;
	wire _w6751_ ;
	wire _w6752_ ;
	wire _w6753_ ;
	wire _w6754_ ;
	wire _w6755_ ;
	wire _w6756_ ;
	wire _w6757_ ;
	wire _w6758_ ;
	wire _w6759_ ;
	wire _w6760_ ;
	wire _w6761_ ;
	wire _w6762_ ;
	wire _w6763_ ;
	wire _w6764_ ;
	wire _w6765_ ;
	wire _w6766_ ;
	wire _w6767_ ;
	wire _w6768_ ;
	wire _w6769_ ;
	wire _w6770_ ;
	wire _w6771_ ;
	wire _w6772_ ;
	wire _w6773_ ;
	wire _w6774_ ;
	wire _w6775_ ;
	wire _w6776_ ;
	wire _w6777_ ;
	wire _w6778_ ;
	wire _w6779_ ;
	wire _w6780_ ;
	wire _w6781_ ;
	wire _w6782_ ;
	wire _w6783_ ;
	wire _w6784_ ;
	wire _w6785_ ;
	wire _w6786_ ;
	wire _w6787_ ;
	wire _w6788_ ;
	wire _w6789_ ;
	wire _w6790_ ;
	wire _w6791_ ;
	wire _w6792_ ;
	wire _w6793_ ;
	wire _w6794_ ;
	wire _w6795_ ;
	wire _w6796_ ;
	wire _w6797_ ;
	wire _w6798_ ;
	wire _w6799_ ;
	wire _w6800_ ;
	wire _w6801_ ;
	wire _w6802_ ;
	wire _w6803_ ;
	wire _w6804_ ;
	wire _w6805_ ;
	wire _w6806_ ;
	wire _w6807_ ;
	wire _w6808_ ;
	wire _w6809_ ;
	wire _w6810_ ;
	wire _w6811_ ;
	wire _w6812_ ;
	wire _w6813_ ;
	wire _w6814_ ;
	wire _w6815_ ;
	wire _w6816_ ;
	wire _w6817_ ;
	wire _w6818_ ;
	wire _w6819_ ;
	wire _w6820_ ;
	wire _w6821_ ;
	wire _w6822_ ;
	wire _w6823_ ;
	wire _w6824_ ;
	wire _w6825_ ;
	wire _w6826_ ;
	wire _w6827_ ;
	wire _w6828_ ;
	wire _w6829_ ;
	wire _w6830_ ;
	wire _w6831_ ;
	wire _w6832_ ;
	wire _w6833_ ;
	wire _w6834_ ;
	wire _w6835_ ;
	wire _w6836_ ;
	LUT1 #(
		.INIT('h1)
	) name0 (
		\u0_u0_idle_cnt1_reg[0]/P0001 ,
		_w103_
	);
	LUT1 #(
		.INIT('h1)
	) name1 (
		\u4_u0_buf0_orig_reg[19]/P0001 ,
		_w862_
	);
	LUT1 #(
		.INIT('h1)
	) name2 (
		\u4_u1_buf0_orig_reg[19]/P0001 ,
		_w1072_
	);
	LUT1 #(
		.INIT('h1)
	) name3 (
		\u4_u2_buf0_orig_reg[19]/P0001 ,
		_w1282_
	);
	LUT1 #(
		.INIT('h1)
	) name4 (
		\u4_u3_buf0_orig_reg[19]/P0001 ,
		_w1492_
	);
	LUT2 #(
		.INIT('h4)
	) name5 (
		TxReady_pad_i_pad,
		\u1_u1_tx_first_r_reg/P0001 ,
		_w1755_
	);
	LUT2 #(
		.INIT('he)
	) name6 (
		\u1_u1_send_zero_length_r_reg/P0001 ,
		\u1_u2_send_data_r_reg/NET0131 ,
		_w1756_
	);
	LUT4 #(
		.INIT('h0001)
	) name7 (
		TxReady_pad_i_pad,
		\u1_u1_send_zero_length_r_reg/P0001 ,
		\u1_u2_send_data_r_reg/NET0131 ,
		\u1_u3_send_token_reg/P0001 ,
		_w1757_
	);
	LUT2 #(
		.INIT('h1)
	) name8 (
		_w1755_,
		_w1757_,
		_w1758_
	);
	LUT2 #(
		.INIT('h2)
	) name9 (
		\DataOut_pad_o[3]_pad ,
		\u0_u0_drive_k_reg/P0001 ,
		_w1759_
	);
	LUT3 #(
		.INIT('he0)
	) name10 (
		_w1755_,
		_w1757_,
		_w1759_,
		_w1760_
	);
	LUT2 #(
		.INIT('h8)
	) name11 (
		\u0_tx_ready_reg/NET0131 ,
		\u1_u1_tx_valid_r_reg/NET0131 ,
		_w1761_
	);
	LUT3 #(
		.INIT('h80)
	) name12 (
		\u0_tx_ready_reg/NET0131 ,
		\u1_u1_state_reg[1]/NET0131 ,
		\u1_u1_tx_valid_r_reg/NET0131 ,
		_w1762_
	);
	LUT4 #(
		.INIT('h0080)
	) name13 (
		\u1_u2_adr_cb_reg[0]/NET0131 ,
		\u1_u2_adr_cb_reg[1]/NET0131 ,
		\u1_u2_adr_cb_reg[2]/NET0131 ,
		\u1_u2_rx_data_valid_r_reg/NET0131 ,
		_w1763_
	);
	LUT3 #(
		.INIT('h20)
	) name14 (
		\u1_u2_rd_buf1_reg[27]/NET0131 ,
		_w1762_,
		_w1763_,
		_w1764_
	);
	LUT4 #(
		.INIT('h007f)
	) name15 (
		\u0_tx_ready_reg/NET0131 ,
		\u1_u1_state_reg[1]/NET0131 ,
		\u1_u1_tx_valid_r_reg/NET0131 ,
		\u1_u2_rx_data_valid_r_reg/NET0131 ,
		_w1765_
	);
	LUT4 #(
		.INIT('h4000)
	) name16 (
		\u1_u2_adr_cb_reg[0]/NET0131 ,
		\u1_u2_adr_cb_reg[1]/NET0131 ,
		\u1_u2_adr_cb_reg[2]/NET0131 ,
		\u1_u2_rd_buf1_reg[27]/NET0131 ,
		_w1766_
	);
	LUT2 #(
		.INIT('h4)
	) name17 (
		_w1765_,
		_w1766_,
		_w1767_
	);
	LUT2 #(
		.INIT('h1)
	) name18 (
		\u1_u2_adr_cb_reg[1]/NET0131 ,
		\u1_u2_rx_data_valid_r_reg/NET0131 ,
		_w1768_
	);
	LUT4 #(
		.INIT('h0020)
	) name19 (
		\u1_u2_adr_cb_reg[0]/NET0131 ,
		\u1_u2_adr_cb_reg[1]/NET0131 ,
		\u1_u2_adr_cb_reg[2]/NET0131 ,
		\u1_u2_rx_data_valid_r_reg/NET0131 ,
		_w1769_
	);
	LUT3 #(
		.INIT('h20)
	) name20 (
		\u1_u2_rd_buf1_reg[11]/NET0131 ,
		_w1762_,
		_w1769_,
		_w1770_
	);
	LUT4 #(
		.INIT('h1000)
	) name21 (
		\u1_u2_adr_cb_reg[0]/NET0131 ,
		\u1_u2_adr_cb_reg[1]/NET0131 ,
		\u1_u2_adr_cb_reg[2]/NET0131 ,
		\u1_u2_rd_buf1_reg[11]/NET0131 ,
		_w1771_
	);
	LUT2 #(
		.INIT('h4)
	) name22 (
		_w1765_,
		_w1771_,
		_w1772_
	);
	LUT4 #(
		.INIT('h0001)
	) name23 (
		_w1764_,
		_w1767_,
		_w1770_,
		_w1772_,
		_w1773_
	);
	LUT4 #(
		.INIT('h0010)
	) name24 (
		\u1_u2_adr_cb_reg[0]/NET0131 ,
		\u1_u2_adr_cb_reg[1]/NET0131 ,
		\u1_u2_adr_cb_reg[2]/NET0131 ,
		\u1_u2_rx_data_valid_r_reg/NET0131 ,
		_w1774_
	);
	LUT3 #(
		.INIT('h20)
	) name25 (
		\u1_u2_rd_buf1_reg[3]/NET0131 ,
		_w1762_,
		_w1774_,
		_w1775_
	);
	LUT4 #(
		.INIT('h0800)
	) name26 (
		\u1_u2_adr_cb_reg[0]/NET0131 ,
		\u1_u2_adr_cb_reg[1]/NET0131 ,
		\u1_u2_adr_cb_reg[2]/NET0131 ,
		\u1_u2_rd_buf1_reg[3]/NET0131 ,
		_w1776_
	);
	LUT2 #(
		.INIT('h4)
	) name27 (
		_w1765_,
		_w1776_,
		_w1777_
	);
	LUT4 #(
		.INIT('h0040)
	) name28 (
		\u1_u2_adr_cb_reg[0]/NET0131 ,
		\u1_u2_adr_cb_reg[1]/NET0131 ,
		\u1_u2_adr_cb_reg[2]/NET0131 ,
		\u1_u2_rx_data_valid_r_reg/NET0131 ,
		_w1778_
	);
	LUT3 #(
		.INIT('h20)
	) name29 (
		\u1_u2_rd_buf1_reg[19]/NET0131 ,
		_w1762_,
		_w1778_,
		_w1779_
	);
	LUT4 #(
		.INIT('h2000)
	) name30 (
		\u1_u2_adr_cb_reg[0]/NET0131 ,
		\u1_u2_adr_cb_reg[1]/NET0131 ,
		\u1_u2_adr_cb_reg[2]/NET0131 ,
		\u1_u2_rd_buf1_reg[19]/NET0131 ,
		_w1780_
	);
	LUT2 #(
		.INIT('h4)
	) name31 (
		_w1765_,
		_w1780_,
		_w1781_
	);
	LUT4 #(
		.INIT('h0001)
	) name32 (
		_w1775_,
		_w1777_,
		_w1779_,
		_w1781_,
		_w1782_
	);
	LUT4 #(
		.INIT('h0008)
	) name33 (
		\u1_u2_adr_cb_reg[0]/NET0131 ,
		\u1_u2_adr_cb_reg[1]/NET0131 ,
		\u1_u2_adr_cb_reg[2]/NET0131 ,
		\u1_u2_rx_data_valid_r_reg/NET0131 ,
		_w1783_
	);
	LUT3 #(
		.INIT('h20)
	) name34 (
		\u1_u2_rd_buf0_reg[27]/NET0131 ,
		_w1762_,
		_w1783_,
		_w1784_
	);
	LUT4 #(
		.INIT('h0400)
	) name35 (
		\u1_u2_adr_cb_reg[0]/NET0131 ,
		\u1_u2_adr_cb_reg[1]/NET0131 ,
		\u1_u2_adr_cb_reg[2]/NET0131 ,
		\u1_u2_rd_buf0_reg[27]/NET0131 ,
		_w1785_
	);
	LUT2 #(
		.INIT('h4)
	) name36 (
		_w1765_,
		_w1785_,
		_w1786_
	);
	LUT4 #(
		.INIT('h0002)
	) name37 (
		\u1_u2_adr_cb_reg[0]/NET0131 ,
		\u1_u2_adr_cb_reg[1]/NET0131 ,
		\u1_u2_adr_cb_reg[2]/NET0131 ,
		\u1_u2_rx_data_valid_r_reg/NET0131 ,
		_w1787_
	);
	LUT3 #(
		.INIT('h20)
	) name38 (
		\u1_u2_rd_buf0_reg[11]/NET0131 ,
		_w1762_,
		_w1787_,
		_w1788_
	);
	LUT4 #(
		.INIT('h0100)
	) name39 (
		\u1_u2_adr_cb_reg[0]/NET0131 ,
		\u1_u2_adr_cb_reg[1]/NET0131 ,
		\u1_u2_adr_cb_reg[2]/NET0131 ,
		\u1_u2_rd_buf0_reg[11]/NET0131 ,
		_w1789_
	);
	LUT2 #(
		.INIT('h4)
	) name40 (
		_w1765_,
		_w1789_,
		_w1790_
	);
	LUT4 #(
		.INIT('h0001)
	) name41 (
		_w1784_,
		_w1786_,
		_w1788_,
		_w1790_,
		_w1791_
	);
	LUT4 #(
		.INIT('h0004)
	) name42 (
		\u1_u2_adr_cb_reg[0]/NET0131 ,
		\u1_u2_adr_cb_reg[1]/NET0131 ,
		\u1_u2_adr_cb_reg[2]/NET0131 ,
		\u1_u2_rx_data_valid_r_reg/NET0131 ,
		_w1792_
	);
	LUT3 #(
		.INIT('h20)
	) name43 (
		\u1_u2_rd_buf0_reg[19]/NET0131 ,
		_w1762_,
		_w1792_,
		_w1793_
	);
	LUT4 #(
		.INIT('h0200)
	) name44 (
		\u1_u2_adr_cb_reg[0]/NET0131 ,
		\u1_u2_adr_cb_reg[1]/NET0131 ,
		\u1_u2_adr_cb_reg[2]/NET0131 ,
		\u1_u2_rd_buf0_reg[19]/NET0131 ,
		_w1794_
	);
	LUT2 #(
		.INIT('h4)
	) name45 (
		_w1765_,
		_w1794_,
		_w1795_
	);
	LUT4 #(
		.INIT('h0001)
	) name46 (
		\u1_u2_adr_cb_reg[0]/NET0131 ,
		\u1_u2_adr_cb_reg[1]/NET0131 ,
		\u1_u2_adr_cb_reg[2]/NET0131 ,
		\u1_u2_rx_data_valid_r_reg/NET0131 ,
		_w1796_
	);
	LUT3 #(
		.INIT('h20)
	) name47 (
		\u1_u2_rd_buf0_reg[3]/NET0131 ,
		_w1762_,
		_w1796_,
		_w1797_
	);
	LUT4 #(
		.INIT('h8000)
	) name48 (
		\u1_u2_adr_cb_reg[0]/NET0131 ,
		\u1_u2_adr_cb_reg[1]/NET0131 ,
		\u1_u2_adr_cb_reg[2]/NET0131 ,
		\u1_u2_rd_buf0_reg[3]/NET0131 ,
		_w1798_
	);
	LUT2 #(
		.INIT('h4)
	) name49 (
		_w1765_,
		_w1798_,
		_w1799_
	);
	LUT4 #(
		.INIT('h0001)
	) name50 (
		_w1793_,
		_w1795_,
		_w1797_,
		_w1799_,
		_w1800_
	);
	LUT4 #(
		.INIT('h8000)
	) name51 (
		_w1773_,
		_w1782_,
		_w1791_,
		_w1800_,
		_w1801_
	);
	LUT4 #(
		.INIT('h0020)
	) name52 (
		\u0_tx_ready_reg/NET0131 ,
		\u1_u1_send_zero_length_r_reg/P0001 ,
		\u1_u1_tx_valid_r_reg/NET0131 ,
		\u1_u2_send_data_r_reg/NET0131 ,
		_w1802_
	);
	LUT3 #(
		.INIT('h01)
	) name53 (
		\u1_u1_state_reg[2]/NET0131 ,
		\u1_u1_state_reg[3]/NET0131 ,
		\u1_u1_state_reg[4]/NET0131 ,
		_w1803_
	);
	LUT2 #(
		.INIT('h4)
	) name54 (
		\u1_u1_state_reg[0]/NET0131 ,
		\u1_u1_state_reg[1]/NET0131 ,
		_w1804_
	);
	LUT3 #(
		.INIT('h80)
	) name55 (
		_w1802_,
		_w1803_,
		_w1804_,
		_w1805_
	);
	LUT2 #(
		.INIT('h1)
	) name56 (
		\u1_u1_state_reg[0]/NET0131 ,
		\u1_u1_state_reg[1]/NET0131 ,
		_w1806_
	);
	LUT3 #(
		.INIT('h01)
	) name57 (
		\u1_u1_state_reg[0]/NET0131 ,
		\u1_u1_state_reg[1]/NET0131 ,
		\u1_u1_state_reg[3]/NET0131 ,
		_w1807_
	);
	LUT2 #(
		.INIT('h4)
	) name58 (
		\u1_u1_state_reg[2]/NET0131 ,
		\u1_u1_state_reg[4]/NET0131 ,
		_w1808_
	);
	LUT3 #(
		.INIT('h04)
	) name59 (
		\u1_u1_state_reg[2]/NET0131 ,
		\u1_u1_state_reg[3]/NET0131 ,
		\u1_u1_state_reg[4]/NET0131 ,
		_w1809_
	);
	LUT4 #(
		.INIT('hebff)
	) name60 (
		\u1_u1_state_reg[2]/NET0131 ,
		\u1_u1_state_reg[3]/NET0131 ,
		\u1_u1_state_reg[4]/NET0131 ,
		_w1806_,
		_w1810_
	);
	LUT2 #(
		.INIT('h1)
	) name61 (
		\u1_u1_send_token_r_reg/P0001 ,
		\u1_u3_send_token_reg/P0001 ,
		_w1811_
	);
	LUT4 #(
		.INIT('h0ee0)
	) name62 (
		\u1_u1_send_token_r_reg/P0001 ,
		\u1_u3_send_token_reg/P0001 ,
		\u1_u3_token_pid_sel_reg[0]/P0001 ,
		\u1_u3_token_pid_sel_reg[1]/P0001 ,
		_w1812_
	);
	LUT4 #(
		.INIT('h0c08)
	) name63 (
		\u1_u1_send_zero_length_r_reg/P0001 ,
		\u1_u1_state_reg[0]/NET0131 ,
		\u1_u1_state_reg[1]/NET0131 ,
		\u1_u2_send_data_r_reg/NET0131 ,
		_w1813_
	);
	LUT2 #(
		.INIT('h8)
	) name64 (
		_w1803_,
		_w1813_,
		_w1814_
	);
	LUT2 #(
		.INIT('h2)
	) name65 (
		\u1_u1_state_reg[2]/NET0131 ,
		\u1_u1_state_reg[4]/NET0131 ,
		_w1815_
	);
	LUT4 #(
		.INIT('h135f)
	) name66 (
		_w1803_,
		_w1807_,
		_w1813_,
		_w1815_,
		_w1816_
	);
	LUT4 #(
		.INIT('h0400)
	) name67 (
		_w1805_,
		_w1810_,
		_w1812_,
		_w1816_,
		_w1817_
	);
	LUT4 #(
		.INIT('he00e)
	) name68 (
		\u1_u1_send_token_r_reg/P0001 ,
		\u1_u3_send_token_reg/P0001 ,
		\u1_u3_token_pid_sel_reg[0]/P0001 ,
		\u1_u3_token_pid_sel_reg[1]/P0001 ,
		_w1818_
	);
	LUT3 #(
		.INIT('h04)
	) name69 (
		\u0_tx_ready_reg/NET0131 ,
		\u1_u1_state_reg[2]/NET0131 ,
		\u1_u1_state_reg[4]/NET0131 ,
		_w1819_
	);
	LUT3 #(
		.INIT('h57)
	) name70 (
		_w1807_,
		_w1808_,
		_w1819_,
		_w1820_
	);
	LUT3 #(
		.INIT('h45)
	) name71 (
		\u1_u1_crc16_reg[12]/P0001 ,
		_w1805_,
		_w1820_,
		_w1821_
	);
	LUT3 #(
		.INIT('h07)
	) name72 (
		\u0_tx_ready_reg/NET0131 ,
		\u1_u1_state_reg[2]/NET0131 ,
		\u1_u3_this_dpid_reg[0]/P0001 ,
		_w1822_
	);
	LUT3 #(
		.INIT('h70)
	) name73 (
		_w1806_,
		_w1809_,
		_w1822_,
		_w1823_
	);
	LUT3 #(
		.INIT('h80)
	) name74 (
		\u0_tx_ready_reg/NET0131 ,
		\u1_u1_crc16_reg[4]/P0001 ,
		\u1_u1_state_reg[2]/NET0131 ,
		_w1824_
	);
	LUT3 #(
		.INIT('h02)
	) name75 (
		\u1_u1_crc16_reg[4]/P0001 ,
		\u1_u1_state_reg[0]/NET0131 ,
		\u1_u1_state_reg[1]/NET0131 ,
		_w1825_
	);
	LUT3 #(
		.INIT('h13)
	) name76 (
		_w1809_,
		_w1824_,
		_w1825_,
		_w1826_
	);
	LUT4 #(
		.INIT('h0400)
	) name77 (
		_w1805_,
		_w1820_,
		_w1823_,
		_w1826_,
		_w1827_
	);
	LUT3 #(
		.INIT('h40)
	) name78 (
		_w1805_,
		_w1810_,
		_w1816_,
		_w1828_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name79 (
		_w1805_,
		_w1810_,
		_w1812_,
		_w1816_,
		_w1829_
	);
	LUT4 #(
		.INIT('h5455)
	) name80 (
		_w1818_,
		_w1821_,
		_w1827_,
		_w1829_,
		_w1830_
	);
	LUT4 #(
		.INIT('h2a00)
	) name81 (
		_w1758_,
		_w1801_,
		_w1817_,
		_w1830_,
		_w1831_
	);
	LUT2 #(
		.INIT('he)
	) name82 (
		_w1760_,
		_w1831_,
		_w1832_
	);
	LUT3 #(
		.INIT('h8a)
	) name83 (
		\u1_u1_crc16_reg[8]/P0001 ,
		_w1805_,
		_w1820_,
		_w1833_
	);
	LUT3 #(
		.INIT('h20)
	) name84 (
		\u0_tx_ready_reg/NET0131 ,
		\u1_u1_crc16_reg[0]/P0001 ,
		\u1_u1_state_reg[2]/NET0131 ,
		_w1834_
	);
	LUT3 #(
		.INIT('h01)
	) name85 (
		\u1_u1_crc16_reg[0]/P0001 ,
		\u1_u1_state_reg[0]/NET0131 ,
		\u1_u1_state_reg[1]/NET0131 ,
		_w1835_
	);
	LUT3 #(
		.INIT('h13)
	) name86 (
		_w1809_,
		_w1834_,
		_w1835_,
		_w1836_
	);
	LUT4 #(
		.INIT('h0400)
	) name87 (
		_w1805_,
		_w1820_,
		_w1823_,
		_w1836_,
		_w1837_
	);
	LUT4 #(
		.INIT('h5551)
	) name88 (
		_w1818_,
		_w1829_,
		_w1833_,
		_w1837_,
		_w1838_
	);
	LUT2 #(
		.INIT('h2)
	) name89 (
		_w1758_,
		_w1838_,
		_w1839_
	);
	LUT2 #(
		.INIT('h2)
	) name90 (
		\DataOut_pad_o[7]_pad ,
		\u0_u0_drive_k_reg/P0001 ,
		_w1840_
	);
	LUT3 #(
		.INIT('he0)
	) name91 (
		_w1755_,
		_w1757_,
		_w1840_,
		_w1841_
	);
	LUT3 #(
		.INIT('h20)
	) name92 (
		\u1_u2_rd_buf0_reg[15]/P0001 ,
		_w1762_,
		_w1787_,
		_w1842_
	);
	LUT4 #(
		.INIT('h0100)
	) name93 (
		\u1_u2_adr_cb_reg[0]/NET0131 ,
		\u1_u2_adr_cb_reg[1]/NET0131 ,
		\u1_u2_adr_cb_reg[2]/NET0131 ,
		\u1_u2_rd_buf0_reg[15]/P0001 ,
		_w1843_
	);
	LUT2 #(
		.INIT('h4)
	) name94 (
		_w1765_,
		_w1843_,
		_w1844_
	);
	LUT3 #(
		.INIT('h20)
	) name95 (
		\u1_u2_rd_buf0_reg[23]/P0001 ,
		_w1762_,
		_w1792_,
		_w1845_
	);
	LUT4 #(
		.INIT('h0200)
	) name96 (
		\u1_u2_adr_cb_reg[0]/NET0131 ,
		\u1_u2_adr_cb_reg[1]/NET0131 ,
		\u1_u2_adr_cb_reg[2]/NET0131 ,
		\u1_u2_rd_buf0_reg[23]/P0001 ,
		_w1846_
	);
	LUT2 #(
		.INIT('h4)
	) name97 (
		_w1765_,
		_w1846_,
		_w1847_
	);
	LUT4 #(
		.INIT('h0001)
	) name98 (
		_w1842_,
		_w1844_,
		_w1845_,
		_w1847_,
		_w1848_
	);
	LUT3 #(
		.INIT('h20)
	) name99 (
		\u1_u2_rd_buf1_reg[7]/P0001 ,
		_w1762_,
		_w1774_,
		_w1849_
	);
	LUT4 #(
		.INIT('h0800)
	) name100 (
		\u1_u2_adr_cb_reg[0]/NET0131 ,
		\u1_u2_adr_cb_reg[1]/NET0131 ,
		\u1_u2_adr_cb_reg[2]/NET0131 ,
		\u1_u2_rd_buf1_reg[7]/P0001 ,
		_w1850_
	);
	LUT2 #(
		.INIT('h4)
	) name101 (
		_w1765_,
		_w1850_,
		_w1851_
	);
	LUT3 #(
		.INIT('h20)
	) name102 (
		\u1_u2_rd_buf1_reg[15]/P0001 ,
		_w1762_,
		_w1769_,
		_w1852_
	);
	LUT4 #(
		.INIT('h1000)
	) name103 (
		\u1_u2_adr_cb_reg[0]/NET0131 ,
		\u1_u2_adr_cb_reg[1]/NET0131 ,
		\u1_u2_adr_cb_reg[2]/NET0131 ,
		\u1_u2_rd_buf1_reg[15]/P0001 ,
		_w1853_
	);
	LUT2 #(
		.INIT('h4)
	) name104 (
		_w1765_,
		_w1853_,
		_w1854_
	);
	LUT4 #(
		.INIT('h0001)
	) name105 (
		_w1849_,
		_w1851_,
		_w1852_,
		_w1854_,
		_w1855_
	);
	LUT3 #(
		.INIT('h20)
	) name106 (
		\u1_u2_rd_buf1_reg[23]/P0001 ,
		_w1762_,
		_w1778_,
		_w1856_
	);
	LUT4 #(
		.INIT('h2000)
	) name107 (
		\u1_u2_adr_cb_reg[0]/NET0131 ,
		\u1_u2_adr_cb_reg[1]/NET0131 ,
		\u1_u2_adr_cb_reg[2]/NET0131 ,
		\u1_u2_rd_buf1_reg[23]/P0001 ,
		_w1857_
	);
	LUT2 #(
		.INIT('h4)
	) name108 (
		_w1765_,
		_w1857_,
		_w1858_
	);
	LUT3 #(
		.INIT('h20)
	) name109 (
		\u1_u2_rd_buf1_reg[31]/P0001 ,
		_w1762_,
		_w1763_,
		_w1859_
	);
	LUT4 #(
		.INIT('h4000)
	) name110 (
		\u1_u2_adr_cb_reg[0]/NET0131 ,
		\u1_u2_adr_cb_reg[1]/NET0131 ,
		\u1_u2_adr_cb_reg[2]/NET0131 ,
		\u1_u2_rd_buf1_reg[31]/P0001 ,
		_w1860_
	);
	LUT2 #(
		.INIT('h4)
	) name111 (
		_w1765_,
		_w1860_,
		_w1861_
	);
	LUT4 #(
		.INIT('h0001)
	) name112 (
		_w1856_,
		_w1858_,
		_w1859_,
		_w1861_,
		_w1862_
	);
	LUT3 #(
		.INIT('h20)
	) name113 (
		\u1_u2_rd_buf0_reg[7]/P0001 ,
		_w1762_,
		_w1796_,
		_w1863_
	);
	LUT4 #(
		.INIT('h8000)
	) name114 (
		\u1_u2_adr_cb_reg[0]/NET0131 ,
		\u1_u2_adr_cb_reg[1]/NET0131 ,
		\u1_u2_adr_cb_reg[2]/NET0131 ,
		\u1_u2_rd_buf0_reg[7]/P0001 ,
		_w1864_
	);
	LUT2 #(
		.INIT('h4)
	) name115 (
		_w1765_,
		_w1864_,
		_w1865_
	);
	LUT3 #(
		.INIT('h20)
	) name116 (
		\u1_u2_rd_buf0_reg[31]/P0001 ,
		_w1762_,
		_w1783_,
		_w1866_
	);
	LUT4 #(
		.INIT('h0400)
	) name117 (
		\u1_u2_adr_cb_reg[0]/NET0131 ,
		\u1_u2_adr_cb_reg[1]/NET0131 ,
		\u1_u2_adr_cb_reg[2]/NET0131 ,
		\u1_u2_rd_buf0_reg[31]/P0001 ,
		_w1867_
	);
	LUT2 #(
		.INIT('h4)
	) name118 (
		_w1765_,
		_w1867_,
		_w1868_
	);
	LUT4 #(
		.INIT('h0001)
	) name119 (
		_w1863_,
		_w1865_,
		_w1866_,
		_w1868_,
		_w1869_
	);
	LUT4 #(
		.INIT('h8000)
	) name120 (
		_w1848_,
		_w1855_,
		_w1862_,
		_w1869_,
		_w1870_
	);
	LUT3 #(
		.INIT('h01)
	) name121 (
		_w1755_,
		_w1757_,
		_w1812_,
		_w1871_
	);
	LUT4 #(
		.INIT('h4000)
	) name122 (
		_w1805_,
		_w1810_,
		_w1816_,
		_w1871_,
		_w1872_
	);
	LUT3 #(
		.INIT('h45)
	) name123 (
		_w1841_,
		_w1870_,
		_w1872_,
		_w1873_
	);
	LUT2 #(
		.INIT('hb)
	) name124 (
		_w1839_,
		_w1873_,
		_w1874_
	);
	LUT2 #(
		.INIT('h2)
	) name125 (
		\DataOut_pad_o[2]_pad ,
		\u0_u0_drive_k_reg/P0001 ,
		_w1875_
	);
	LUT3 #(
		.INIT('he0)
	) name126 (
		_w1755_,
		_w1757_,
		_w1875_,
		_w1876_
	);
	LUT3 #(
		.INIT('h20)
	) name127 (
		\u1_u2_rd_buf0_reg[2]/NET0131 ,
		_w1762_,
		_w1796_,
		_w1877_
	);
	LUT4 #(
		.INIT('h8000)
	) name128 (
		\u1_u2_adr_cb_reg[0]/NET0131 ,
		\u1_u2_adr_cb_reg[1]/NET0131 ,
		\u1_u2_adr_cb_reg[2]/NET0131 ,
		\u1_u2_rd_buf0_reg[2]/NET0131 ,
		_w1878_
	);
	LUT2 #(
		.INIT('h4)
	) name129 (
		_w1765_,
		_w1878_,
		_w1879_
	);
	LUT3 #(
		.INIT('h20)
	) name130 (
		\u1_u2_rd_buf1_reg[18]/NET0131 ,
		_w1762_,
		_w1778_,
		_w1880_
	);
	LUT4 #(
		.INIT('h2000)
	) name131 (
		\u1_u2_adr_cb_reg[0]/NET0131 ,
		\u1_u2_adr_cb_reg[1]/NET0131 ,
		\u1_u2_adr_cb_reg[2]/NET0131 ,
		\u1_u2_rd_buf1_reg[18]/NET0131 ,
		_w1881_
	);
	LUT2 #(
		.INIT('h4)
	) name132 (
		_w1765_,
		_w1881_,
		_w1882_
	);
	LUT4 #(
		.INIT('h0001)
	) name133 (
		_w1877_,
		_w1879_,
		_w1880_,
		_w1882_,
		_w1883_
	);
	LUT3 #(
		.INIT('h20)
	) name134 (
		\u1_u2_rd_buf0_reg[18]/NET0131 ,
		_w1762_,
		_w1792_,
		_w1884_
	);
	LUT4 #(
		.INIT('h0200)
	) name135 (
		\u1_u2_adr_cb_reg[0]/NET0131 ,
		\u1_u2_adr_cb_reg[1]/NET0131 ,
		\u1_u2_adr_cb_reg[2]/NET0131 ,
		\u1_u2_rd_buf0_reg[18]/NET0131 ,
		_w1885_
	);
	LUT2 #(
		.INIT('h4)
	) name136 (
		_w1765_,
		_w1885_,
		_w1886_
	);
	LUT3 #(
		.INIT('h20)
	) name137 (
		\u1_u2_rd_buf1_reg[2]/NET0131 ,
		_w1762_,
		_w1774_,
		_w1887_
	);
	LUT4 #(
		.INIT('h0800)
	) name138 (
		\u1_u2_adr_cb_reg[0]/NET0131 ,
		\u1_u2_adr_cb_reg[1]/NET0131 ,
		\u1_u2_adr_cb_reg[2]/NET0131 ,
		\u1_u2_rd_buf1_reg[2]/NET0131 ,
		_w1888_
	);
	LUT2 #(
		.INIT('h4)
	) name139 (
		_w1765_,
		_w1888_,
		_w1889_
	);
	LUT4 #(
		.INIT('h0001)
	) name140 (
		_w1884_,
		_w1886_,
		_w1887_,
		_w1889_,
		_w1890_
	);
	LUT3 #(
		.INIT('h20)
	) name141 (
		\u1_u2_rd_buf0_reg[10]/NET0131 ,
		_w1762_,
		_w1787_,
		_w1891_
	);
	LUT4 #(
		.INIT('h0100)
	) name142 (
		\u1_u2_adr_cb_reg[0]/NET0131 ,
		\u1_u2_adr_cb_reg[1]/NET0131 ,
		\u1_u2_adr_cb_reg[2]/NET0131 ,
		\u1_u2_rd_buf0_reg[10]/NET0131 ,
		_w1892_
	);
	LUT2 #(
		.INIT('h4)
	) name143 (
		_w1765_,
		_w1892_,
		_w1893_
	);
	LUT3 #(
		.INIT('h20)
	) name144 (
		\u1_u2_rd_buf0_reg[26]/NET0131 ,
		_w1762_,
		_w1783_,
		_w1894_
	);
	LUT4 #(
		.INIT('h0400)
	) name145 (
		\u1_u2_adr_cb_reg[0]/NET0131 ,
		\u1_u2_adr_cb_reg[1]/NET0131 ,
		\u1_u2_adr_cb_reg[2]/NET0131 ,
		\u1_u2_rd_buf0_reg[26]/NET0131 ,
		_w1895_
	);
	LUT2 #(
		.INIT('h4)
	) name146 (
		_w1765_,
		_w1895_,
		_w1896_
	);
	LUT4 #(
		.INIT('h0001)
	) name147 (
		_w1891_,
		_w1893_,
		_w1894_,
		_w1896_,
		_w1897_
	);
	LUT3 #(
		.INIT('h20)
	) name148 (
		\u1_u2_rd_buf1_reg[26]/NET0131 ,
		_w1762_,
		_w1763_,
		_w1898_
	);
	LUT4 #(
		.INIT('h4000)
	) name149 (
		\u1_u2_adr_cb_reg[0]/NET0131 ,
		\u1_u2_adr_cb_reg[1]/NET0131 ,
		\u1_u2_adr_cb_reg[2]/NET0131 ,
		\u1_u2_rd_buf1_reg[26]/NET0131 ,
		_w1899_
	);
	LUT2 #(
		.INIT('h4)
	) name150 (
		_w1765_,
		_w1899_,
		_w1900_
	);
	LUT3 #(
		.INIT('h20)
	) name151 (
		\u1_u2_rd_buf1_reg[10]/NET0131 ,
		_w1762_,
		_w1769_,
		_w1901_
	);
	LUT4 #(
		.INIT('h1000)
	) name152 (
		\u1_u2_adr_cb_reg[0]/NET0131 ,
		\u1_u2_adr_cb_reg[1]/NET0131 ,
		\u1_u2_adr_cb_reg[2]/NET0131 ,
		\u1_u2_rd_buf1_reg[10]/NET0131 ,
		_w1902_
	);
	LUT2 #(
		.INIT('h4)
	) name153 (
		_w1765_,
		_w1902_,
		_w1903_
	);
	LUT4 #(
		.INIT('h0001)
	) name154 (
		_w1898_,
		_w1900_,
		_w1901_,
		_w1903_,
		_w1904_
	);
	LUT4 #(
		.INIT('h8000)
	) name155 (
		_w1883_,
		_w1890_,
		_w1897_,
		_w1904_,
		_w1905_
	);
	LUT3 #(
		.INIT('he0)
	) name156 (
		\u1_u1_send_token_r_reg/P0001 ,
		\u1_u3_send_token_reg/P0001 ,
		\u1_u3_token_pid_sel_reg[1]/P0001 ,
		_w1906_
	);
	LUT4 #(
		.INIT('h0040)
	) name157 (
		_w1805_,
		_w1810_,
		_w1816_,
		_w1906_,
		_w1907_
	);
	LUT3 #(
		.INIT('h0e)
	) name158 (
		\u1_u1_send_token_r_reg/P0001 ,
		\u1_u3_send_token_reg/P0001 ,
		\u1_u3_token_pid_sel_reg[1]/P0001 ,
		_w1908_
	);
	LUT3 #(
		.INIT('h45)
	) name159 (
		\u1_u1_crc16_reg[13]/P0001 ,
		_w1805_,
		_w1820_,
		_w1909_
	);
	LUT3 #(
		.INIT('h80)
	) name160 (
		\u0_tx_ready_reg/NET0131 ,
		\u1_u1_crc16_reg[5]/P0001 ,
		\u1_u1_state_reg[2]/NET0131 ,
		_w1910_
	);
	LUT3 #(
		.INIT('h02)
	) name161 (
		\u1_u1_crc16_reg[5]/P0001 ,
		\u1_u1_state_reg[0]/NET0131 ,
		\u1_u1_state_reg[1]/NET0131 ,
		_w1911_
	);
	LUT3 #(
		.INIT('h13)
	) name162 (
		_w1809_,
		_w1910_,
		_w1911_,
		_w1912_
	);
	LUT3 #(
		.INIT('h07)
	) name163 (
		\u0_tx_ready_reg/NET0131 ,
		\u1_u1_state_reg[2]/NET0131 ,
		\u1_u3_this_dpid_reg[1]/P0001 ,
		_w1913_
	);
	LUT3 #(
		.INIT('h70)
	) name164 (
		_w1806_,
		_w1809_,
		_w1913_,
		_w1914_
	);
	LUT4 #(
		.INIT('h0040)
	) name165 (
		_w1805_,
		_w1820_,
		_w1912_,
		_w1914_,
		_w1915_
	);
	LUT4 #(
		.INIT('h00bf)
	) name166 (
		_w1805_,
		_w1810_,
		_w1816_,
		_w1906_,
		_w1916_
	);
	LUT4 #(
		.INIT('h5455)
	) name167 (
		_w1908_,
		_w1909_,
		_w1915_,
		_w1916_,
		_w1917_
	);
	LUT4 #(
		.INIT('h2a00)
	) name168 (
		_w1758_,
		_w1905_,
		_w1907_,
		_w1917_,
		_w1918_
	);
	LUT2 #(
		.INIT('he)
	) name169 (
		_w1876_,
		_w1918_,
		_w1919_
	);
	LUT3 #(
		.INIT('h8a)
	) name170 (
		\u1_u1_crc16_reg[9]/P0001 ,
		_w1805_,
		_w1820_,
		_w1920_
	);
	LUT3 #(
		.INIT('h20)
	) name171 (
		\u0_tx_ready_reg/NET0131 ,
		\u1_u1_crc16_reg[1]/P0001 ,
		\u1_u1_state_reg[2]/NET0131 ,
		_w1921_
	);
	LUT3 #(
		.INIT('h01)
	) name172 (
		\u1_u1_crc16_reg[1]/P0001 ,
		\u1_u1_state_reg[0]/NET0131 ,
		\u1_u1_state_reg[1]/NET0131 ,
		_w1922_
	);
	LUT3 #(
		.INIT('h13)
	) name173 (
		_w1809_,
		_w1921_,
		_w1922_,
		_w1923_
	);
	LUT4 #(
		.INIT('h0400)
	) name174 (
		_w1805_,
		_w1820_,
		_w1914_,
		_w1923_,
		_w1924_
	);
	LUT4 #(
		.INIT('h5551)
	) name175 (
		_w1908_,
		_w1916_,
		_w1920_,
		_w1924_,
		_w1925_
	);
	LUT2 #(
		.INIT('h2)
	) name176 (
		_w1758_,
		_w1925_,
		_w1926_
	);
	LUT2 #(
		.INIT('h2)
	) name177 (
		\DataOut_pad_o[6]_pad ,
		\u0_u0_drive_k_reg/P0001 ,
		_w1927_
	);
	LUT3 #(
		.INIT('he0)
	) name178 (
		_w1755_,
		_w1757_,
		_w1927_,
		_w1928_
	);
	LUT3 #(
		.INIT('h20)
	) name179 (
		\u1_u2_rd_buf1_reg[6]/P0001 ,
		_w1762_,
		_w1774_,
		_w1929_
	);
	LUT4 #(
		.INIT('h0800)
	) name180 (
		\u1_u2_adr_cb_reg[0]/NET0131 ,
		\u1_u2_adr_cb_reg[1]/NET0131 ,
		\u1_u2_adr_cb_reg[2]/NET0131 ,
		\u1_u2_rd_buf1_reg[6]/P0001 ,
		_w1930_
	);
	LUT2 #(
		.INIT('h4)
	) name181 (
		_w1765_,
		_w1930_,
		_w1931_
	);
	LUT3 #(
		.INIT('h20)
	) name182 (
		\u1_u2_rd_buf1_reg[14]/P0001 ,
		_w1762_,
		_w1769_,
		_w1932_
	);
	LUT4 #(
		.INIT('h1000)
	) name183 (
		\u1_u2_adr_cb_reg[0]/NET0131 ,
		\u1_u2_adr_cb_reg[1]/NET0131 ,
		\u1_u2_adr_cb_reg[2]/NET0131 ,
		\u1_u2_rd_buf1_reg[14]/P0001 ,
		_w1933_
	);
	LUT2 #(
		.INIT('h4)
	) name184 (
		_w1765_,
		_w1933_,
		_w1934_
	);
	LUT4 #(
		.INIT('h0001)
	) name185 (
		_w1929_,
		_w1931_,
		_w1932_,
		_w1934_,
		_w1935_
	);
	LUT3 #(
		.INIT('h20)
	) name186 (
		\u1_u2_rd_buf0_reg[14]/P0001 ,
		_w1762_,
		_w1787_,
		_w1936_
	);
	LUT4 #(
		.INIT('h0100)
	) name187 (
		\u1_u2_adr_cb_reg[0]/NET0131 ,
		\u1_u2_adr_cb_reg[1]/NET0131 ,
		\u1_u2_adr_cb_reg[2]/NET0131 ,
		\u1_u2_rd_buf0_reg[14]/P0001 ,
		_w1937_
	);
	LUT2 #(
		.INIT('h4)
	) name188 (
		_w1765_,
		_w1937_,
		_w1938_
	);
	LUT3 #(
		.INIT('h20)
	) name189 (
		\u1_u2_rd_buf1_reg[22]/P0001 ,
		_w1762_,
		_w1778_,
		_w1939_
	);
	LUT4 #(
		.INIT('h2000)
	) name190 (
		\u1_u2_adr_cb_reg[0]/NET0131 ,
		\u1_u2_adr_cb_reg[1]/NET0131 ,
		\u1_u2_adr_cb_reg[2]/NET0131 ,
		\u1_u2_rd_buf1_reg[22]/P0001 ,
		_w1940_
	);
	LUT2 #(
		.INIT('h4)
	) name191 (
		_w1765_,
		_w1940_,
		_w1941_
	);
	LUT4 #(
		.INIT('h0001)
	) name192 (
		_w1936_,
		_w1938_,
		_w1939_,
		_w1941_,
		_w1942_
	);
	LUT3 #(
		.INIT('h20)
	) name193 (
		\u1_u2_rd_buf1_reg[30]/P0001 ,
		_w1762_,
		_w1763_,
		_w1943_
	);
	LUT4 #(
		.INIT('h4000)
	) name194 (
		\u1_u2_adr_cb_reg[0]/NET0131 ,
		\u1_u2_adr_cb_reg[1]/NET0131 ,
		\u1_u2_adr_cb_reg[2]/NET0131 ,
		\u1_u2_rd_buf1_reg[30]/P0001 ,
		_w1944_
	);
	LUT2 #(
		.INIT('h4)
	) name195 (
		_w1765_,
		_w1944_,
		_w1945_
	);
	LUT3 #(
		.INIT('h20)
	) name196 (
		\u1_u2_rd_buf0_reg[30]/P0001 ,
		_w1762_,
		_w1783_,
		_w1946_
	);
	LUT4 #(
		.INIT('h0400)
	) name197 (
		\u1_u2_adr_cb_reg[0]/NET0131 ,
		\u1_u2_adr_cb_reg[1]/NET0131 ,
		\u1_u2_adr_cb_reg[2]/NET0131 ,
		\u1_u2_rd_buf0_reg[30]/P0001 ,
		_w1947_
	);
	LUT2 #(
		.INIT('h4)
	) name198 (
		_w1765_,
		_w1947_,
		_w1948_
	);
	LUT4 #(
		.INIT('h0001)
	) name199 (
		_w1943_,
		_w1945_,
		_w1946_,
		_w1948_,
		_w1949_
	);
	LUT3 #(
		.INIT('h20)
	) name200 (
		\u1_u2_rd_buf0_reg[6]/P0001 ,
		_w1762_,
		_w1796_,
		_w1950_
	);
	LUT4 #(
		.INIT('h8000)
	) name201 (
		\u1_u2_adr_cb_reg[0]/NET0131 ,
		\u1_u2_adr_cb_reg[1]/NET0131 ,
		\u1_u2_adr_cb_reg[2]/NET0131 ,
		\u1_u2_rd_buf0_reg[6]/P0001 ,
		_w1951_
	);
	LUT2 #(
		.INIT('h4)
	) name202 (
		_w1765_,
		_w1951_,
		_w1952_
	);
	LUT3 #(
		.INIT('h20)
	) name203 (
		\u1_u2_rd_buf0_reg[22]/P0001 ,
		_w1762_,
		_w1792_,
		_w1953_
	);
	LUT4 #(
		.INIT('h0200)
	) name204 (
		\u1_u2_adr_cb_reg[0]/NET0131 ,
		\u1_u2_adr_cb_reg[1]/NET0131 ,
		\u1_u2_adr_cb_reg[2]/NET0131 ,
		\u1_u2_rd_buf0_reg[22]/P0001 ,
		_w1954_
	);
	LUT2 #(
		.INIT('h4)
	) name205 (
		_w1765_,
		_w1954_,
		_w1955_
	);
	LUT4 #(
		.INIT('h0001)
	) name206 (
		_w1950_,
		_w1952_,
		_w1953_,
		_w1955_,
		_w1956_
	);
	LUT4 #(
		.INIT('h8000)
	) name207 (
		_w1935_,
		_w1942_,
		_w1949_,
		_w1956_,
		_w1957_
	);
	LUT3 #(
		.INIT('h01)
	) name208 (
		_w1755_,
		_w1757_,
		_w1906_,
		_w1958_
	);
	LUT4 #(
		.INIT('h4000)
	) name209 (
		_w1805_,
		_w1810_,
		_w1816_,
		_w1958_,
		_w1959_
	);
	LUT3 #(
		.INIT('h45)
	) name210 (
		_w1928_,
		_w1957_,
		_w1959_,
		_w1960_
	);
	LUT2 #(
		.INIT('hb)
	) name211 (
		_w1926_,
		_w1960_,
		_w1961_
	);
	LUT3 #(
		.INIT('h20)
	) name212 (
		\u1_u2_rd_buf0_reg[4]/P0001 ,
		_w1762_,
		_w1796_,
		_w1962_
	);
	LUT4 #(
		.INIT('h8000)
	) name213 (
		\u1_u2_adr_cb_reg[0]/NET0131 ,
		\u1_u2_adr_cb_reg[1]/NET0131 ,
		\u1_u2_adr_cb_reg[2]/NET0131 ,
		\u1_u2_rd_buf0_reg[4]/P0001 ,
		_w1963_
	);
	LUT2 #(
		.INIT('h4)
	) name214 (
		_w1765_,
		_w1963_,
		_w1964_
	);
	LUT3 #(
		.INIT('h20)
	) name215 (
		\u1_u2_rd_buf0_reg[12]/P0001 ,
		_w1762_,
		_w1787_,
		_w1965_
	);
	LUT4 #(
		.INIT('h0100)
	) name216 (
		\u1_u2_adr_cb_reg[0]/NET0131 ,
		\u1_u2_adr_cb_reg[1]/NET0131 ,
		\u1_u2_adr_cb_reg[2]/NET0131 ,
		\u1_u2_rd_buf0_reg[12]/P0001 ,
		_w1966_
	);
	LUT2 #(
		.INIT('h4)
	) name217 (
		_w1765_,
		_w1966_,
		_w1967_
	);
	LUT4 #(
		.INIT('h0001)
	) name218 (
		_w1962_,
		_w1964_,
		_w1965_,
		_w1967_,
		_w1968_
	);
	LUT3 #(
		.INIT('h20)
	) name219 (
		\u1_u2_rd_buf1_reg[20]/P0001 ,
		_w1762_,
		_w1778_,
		_w1969_
	);
	LUT4 #(
		.INIT('h2000)
	) name220 (
		\u1_u2_adr_cb_reg[0]/NET0131 ,
		\u1_u2_adr_cb_reg[1]/NET0131 ,
		\u1_u2_adr_cb_reg[2]/NET0131 ,
		\u1_u2_rd_buf1_reg[20]/P0001 ,
		_w1970_
	);
	LUT2 #(
		.INIT('h4)
	) name221 (
		_w1765_,
		_w1970_,
		_w1971_
	);
	LUT3 #(
		.INIT('h20)
	) name222 (
		\u1_u2_rd_buf1_reg[28]/P0001 ,
		_w1762_,
		_w1763_,
		_w1972_
	);
	LUT4 #(
		.INIT('h4000)
	) name223 (
		\u1_u2_adr_cb_reg[0]/NET0131 ,
		\u1_u2_adr_cb_reg[1]/NET0131 ,
		\u1_u2_adr_cb_reg[2]/NET0131 ,
		\u1_u2_rd_buf1_reg[28]/P0001 ,
		_w1973_
	);
	LUT2 #(
		.INIT('h4)
	) name224 (
		_w1765_,
		_w1973_,
		_w1974_
	);
	LUT4 #(
		.INIT('h0001)
	) name225 (
		_w1969_,
		_w1971_,
		_w1972_,
		_w1974_,
		_w1975_
	);
	LUT3 #(
		.INIT('h20)
	) name226 (
		\u1_u2_rd_buf0_reg[20]/P0001 ,
		_w1762_,
		_w1792_,
		_w1976_
	);
	LUT4 #(
		.INIT('h0200)
	) name227 (
		\u1_u2_adr_cb_reg[0]/NET0131 ,
		\u1_u2_adr_cb_reg[1]/NET0131 ,
		\u1_u2_adr_cb_reg[2]/NET0131 ,
		\u1_u2_rd_buf0_reg[20]/P0001 ,
		_w1977_
	);
	LUT2 #(
		.INIT('h4)
	) name228 (
		_w1765_,
		_w1977_,
		_w1978_
	);
	LUT3 #(
		.INIT('h20)
	) name229 (
		\u1_u2_rd_buf0_reg[28]/P0001 ,
		_w1762_,
		_w1783_,
		_w1979_
	);
	LUT4 #(
		.INIT('h0400)
	) name230 (
		\u1_u2_adr_cb_reg[0]/NET0131 ,
		\u1_u2_adr_cb_reg[1]/NET0131 ,
		\u1_u2_adr_cb_reg[2]/NET0131 ,
		\u1_u2_rd_buf0_reg[28]/P0001 ,
		_w1980_
	);
	LUT2 #(
		.INIT('h4)
	) name231 (
		_w1765_,
		_w1980_,
		_w1981_
	);
	LUT4 #(
		.INIT('h0001)
	) name232 (
		_w1976_,
		_w1978_,
		_w1979_,
		_w1981_,
		_w1982_
	);
	LUT3 #(
		.INIT('h20)
	) name233 (
		\u1_u2_rd_buf1_reg[4]/P0001 ,
		_w1762_,
		_w1774_,
		_w1983_
	);
	LUT4 #(
		.INIT('h0800)
	) name234 (
		\u1_u2_adr_cb_reg[0]/NET0131 ,
		\u1_u2_adr_cb_reg[1]/NET0131 ,
		\u1_u2_adr_cb_reg[2]/NET0131 ,
		\u1_u2_rd_buf1_reg[4]/P0001 ,
		_w1984_
	);
	LUT2 #(
		.INIT('h4)
	) name235 (
		_w1765_,
		_w1984_,
		_w1985_
	);
	LUT3 #(
		.INIT('h20)
	) name236 (
		\u1_u2_rd_buf1_reg[12]/P0001 ,
		_w1762_,
		_w1769_,
		_w1986_
	);
	LUT4 #(
		.INIT('h1000)
	) name237 (
		\u1_u2_adr_cb_reg[0]/NET0131 ,
		\u1_u2_adr_cb_reg[1]/NET0131 ,
		\u1_u2_adr_cb_reg[2]/NET0131 ,
		\u1_u2_rd_buf1_reg[12]/P0001 ,
		_w1987_
	);
	LUT2 #(
		.INIT('h4)
	) name238 (
		_w1765_,
		_w1987_,
		_w1988_
	);
	LUT4 #(
		.INIT('h0001)
	) name239 (
		_w1983_,
		_w1985_,
		_w1986_,
		_w1988_,
		_w1989_
	);
	LUT4 #(
		.INIT('h8000)
	) name240 (
		_w1968_,
		_w1975_,
		_w1982_,
		_w1989_,
		_w1990_
	);
	LUT3 #(
		.INIT('h20)
	) name241 (
		\u1_u2_rd_buf1_reg[5]/P0001 ,
		_w1762_,
		_w1774_,
		_w1991_
	);
	LUT4 #(
		.INIT('h0800)
	) name242 (
		\u1_u2_adr_cb_reg[0]/NET0131 ,
		\u1_u2_adr_cb_reg[1]/NET0131 ,
		\u1_u2_adr_cb_reg[2]/NET0131 ,
		\u1_u2_rd_buf1_reg[5]/P0001 ,
		_w1992_
	);
	LUT2 #(
		.INIT('h4)
	) name243 (
		_w1765_,
		_w1992_,
		_w1993_
	);
	LUT3 #(
		.INIT('h20)
	) name244 (
		\u1_u2_rd_buf1_reg[13]/P0001 ,
		_w1762_,
		_w1769_,
		_w1994_
	);
	LUT4 #(
		.INIT('h1000)
	) name245 (
		\u1_u2_adr_cb_reg[0]/NET0131 ,
		\u1_u2_adr_cb_reg[1]/NET0131 ,
		\u1_u2_adr_cb_reg[2]/NET0131 ,
		\u1_u2_rd_buf1_reg[13]/P0001 ,
		_w1995_
	);
	LUT2 #(
		.INIT('h4)
	) name246 (
		_w1765_,
		_w1995_,
		_w1996_
	);
	LUT4 #(
		.INIT('h0001)
	) name247 (
		_w1991_,
		_w1993_,
		_w1994_,
		_w1996_,
		_w1997_
	);
	LUT3 #(
		.INIT('h20)
	) name248 (
		\u1_u2_rd_buf1_reg[21]/P0001 ,
		_w1762_,
		_w1778_,
		_w1998_
	);
	LUT4 #(
		.INIT('h2000)
	) name249 (
		\u1_u2_adr_cb_reg[0]/NET0131 ,
		\u1_u2_adr_cb_reg[1]/NET0131 ,
		\u1_u2_adr_cb_reg[2]/NET0131 ,
		\u1_u2_rd_buf1_reg[21]/P0001 ,
		_w1999_
	);
	LUT2 #(
		.INIT('h4)
	) name250 (
		_w1765_,
		_w1999_,
		_w2000_
	);
	LUT3 #(
		.INIT('h20)
	) name251 (
		\u1_u2_rd_buf1_reg[29]/P0001 ,
		_w1762_,
		_w1763_,
		_w2001_
	);
	LUT4 #(
		.INIT('h4000)
	) name252 (
		\u1_u2_adr_cb_reg[0]/NET0131 ,
		\u1_u2_adr_cb_reg[1]/NET0131 ,
		\u1_u2_adr_cb_reg[2]/NET0131 ,
		\u1_u2_rd_buf1_reg[29]/P0001 ,
		_w2002_
	);
	LUT2 #(
		.INIT('h4)
	) name253 (
		_w1765_,
		_w2002_,
		_w2003_
	);
	LUT4 #(
		.INIT('h0001)
	) name254 (
		_w1998_,
		_w2000_,
		_w2001_,
		_w2003_,
		_w2004_
	);
	LUT3 #(
		.INIT('h20)
	) name255 (
		\u1_u2_rd_buf0_reg[29]/P0001 ,
		_w1762_,
		_w1783_,
		_w2005_
	);
	LUT4 #(
		.INIT('h0400)
	) name256 (
		\u1_u2_adr_cb_reg[0]/NET0131 ,
		\u1_u2_adr_cb_reg[1]/NET0131 ,
		\u1_u2_adr_cb_reg[2]/NET0131 ,
		\u1_u2_rd_buf0_reg[29]/P0001 ,
		_w2006_
	);
	LUT2 #(
		.INIT('h4)
	) name257 (
		_w1765_,
		_w2006_,
		_w2007_
	);
	LUT3 #(
		.INIT('h20)
	) name258 (
		\u1_u2_rd_buf0_reg[21]/P0001 ,
		_w1762_,
		_w1792_,
		_w2008_
	);
	LUT4 #(
		.INIT('h0200)
	) name259 (
		\u1_u2_adr_cb_reg[0]/NET0131 ,
		\u1_u2_adr_cb_reg[1]/NET0131 ,
		\u1_u2_adr_cb_reg[2]/NET0131 ,
		\u1_u2_rd_buf0_reg[21]/P0001 ,
		_w2009_
	);
	LUT2 #(
		.INIT('h4)
	) name260 (
		_w1765_,
		_w2009_,
		_w2010_
	);
	LUT4 #(
		.INIT('h0001)
	) name261 (
		_w2005_,
		_w2007_,
		_w2008_,
		_w2010_,
		_w2011_
	);
	LUT3 #(
		.INIT('h20)
	) name262 (
		\u1_u2_rd_buf0_reg[13]/P0001 ,
		_w1762_,
		_w1787_,
		_w2012_
	);
	LUT4 #(
		.INIT('h0100)
	) name263 (
		\u1_u2_adr_cb_reg[0]/NET0131 ,
		\u1_u2_adr_cb_reg[1]/NET0131 ,
		\u1_u2_adr_cb_reg[2]/NET0131 ,
		\u1_u2_rd_buf0_reg[13]/P0001 ,
		_w2013_
	);
	LUT2 #(
		.INIT('h4)
	) name264 (
		_w1765_,
		_w2013_,
		_w2014_
	);
	LUT3 #(
		.INIT('h20)
	) name265 (
		\u1_u2_rd_buf0_reg[5]/P0001 ,
		_w1762_,
		_w1796_,
		_w2015_
	);
	LUT4 #(
		.INIT('h8000)
	) name266 (
		\u1_u2_adr_cb_reg[0]/NET0131 ,
		\u1_u2_adr_cb_reg[1]/NET0131 ,
		\u1_u2_adr_cb_reg[2]/NET0131 ,
		\u1_u2_rd_buf0_reg[5]/P0001 ,
		_w2016_
	);
	LUT2 #(
		.INIT('h4)
	) name267 (
		_w1765_,
		_w2016_,
		_w2017_
	);
	LUT4 #(
		.INIT('h0001)
	) name268 (
		_w2012_,
		_w2014_,
		_w2015_,
		_w2017_,
		_w2018_
	);
	LUT4 #(
		.INIT('h8000)
	) name269 (
		_w1997_,
		_w2004_,
		_w2011_,
		_w2018_,
		_w2019_
	);
	LUT4 #(
		.INIT('h6996)
	) name270 (
		_w1870_,
		_w1957_,
		_w1990_,
		_w2019_,
		_w2020_
	);
	LUT2 #(
		.INIT('h9)
	) name271 (
		\u1_u1_crc16_reg[7]/P0001 ,
		\u1_u1_crc16_reg[8]/P0001 ,
		_w2021_
	);
	LUT2 #(
		.INIT('h9)
	) name272 (
		_w1801_,
		_w1905_,
		_w2022_
	);
	LUT3 #(
		.INIT('h69)
	) name273 (
		_w2020_,
		_w2021_,
		_w2022_,
		_w2023_
	);
	LUT2 #(
		.INIT('h6)
	) name274 (
		\u1_u1_crc16_reg[13]/P0001 ,
		\u1_u1_crc16_reg[14]/P0001 ,
		_w2024_
	);
	LUT3 #(
		.INIT('h20)
	) name275 (
		\u1_u2_rd_buf0_reg[16]/NET0131 ,
		_w1762_,
		_w1792_,
		_w2025_
	);
	LUT4 #(
		.INIT('h0200)
	) name276 (
		\u1_u2_adr_cb_reg[0]/NET0131 ,
		\u1_u2_adr_cb_reg[1]/NET0131 ,
		\u1_u2_adr_cb_reg[2]/NET0131 ,
		\u1_u2_rd_buf0_reg[16]/NET0131 ,
		_w2026_
	);
	LUT2 #(
		.INIT('h4)
	) name277 (
		_w1765_,
		_w2026_,
		_w2027_
	);
	LUT3 #(
		.INIT('h20)
	) name278 (
		\u1_u2_rd_buf1_reg[8]/NET0131 ,
		_w1762_,
		_w1769_,
		_w2028_
	);
	LUT4 #(
		.INIT('h1000)
	) name279 (
		\u1_u2_adr_cb_reg[0]/NET0131 ,
		\u1_u2_adr_cb_reg[1]/NET0131 ,
		\u1_u2_adr_cb_reg[2]/NET0131 ,
		\u1_u2_rd_buf1_reg[8]/NET0131 ,
		_w2029_
	);
	LUT2 #(
		.INIT('h4)
	) name280 (
		_w1765_,
		_w2029_,
		_w2030_
	);
	LUT4 #(
		.INIT('h0001)
	) name281 (
		_w2025_,
		_w2027_,
		_w2028_,
		_w2030_,
		_w2031_
	);
	LUT3 #(
		.INIT('h20)
	) name282 (
		\u1_u2_rd_buf1_reg[0]/NET0131 ,
		_w1762_,
		_w1774_,
		_w2032_
	);
	LUT4 #(
		.INIT('h0800)
	) name283 (
		\u1_u2_adr_cb_reg[0]/NET0131 ,
		\u1_u2_adr_cb_reg[1]/NET0131 ,
		\u1_u2_adr_cb_reg[2]/NET0131 ,
		\u1_u2_rd_buf1_reg[0]/NET0131 ,
		_w2033_
	);
	LUT2 #(
		.INIT('h4)
	) name284 (
		_w1765_,
		_w2033_,
		_w2034_
	);
	LUT3 #(
		.INIT('h20)
	) name285 (
		\u1_u2_rd_buf0_reg[24]/NET0131 ,
		_w1762_,
		_w1783_,
		_w2035_
	);
	LUT4 #(
		.INIT('h0400)
	) name286 (
		\u1_u2_adr_cb_reg[0]/NET0131 ,
		\u1_u2_adr_cb_reg[1]/NET0131 ,
		\u1_u2_adr_cb_reg[2]/NET0131 ,
		\u1_u2_rd_buf0_reg[24]/NET0131 ,
		_w2036_
	);
	LUT2 #(
		.INIT('h4)
	) name287 (
		_w1765_,
		_w2036_,
		_w2037_
	);
	LUT4 #(
		.INIT('h0001)
	) name288 (
		_w2032_,
		_w2034_,
		_w2035_,
		_w2037_,
		_w2038_
	);
	LUT3 #(
		.INIT('h20)
	) name289 (
		\u1_u2_rd_buf0_reg[8]/NET0131 ,
		_w1762_,
		_w1787_,
		_w2039_
	);
	LUT4 #(
		.INIT('h0100)
	) name290 (
		\u1_u2_adr_cb_reg[0]/NET0131 ,
		\u1_u2_adr_cb_reg[1]/NET0131 ,
		\u1_u2_adr_cb_reg[2]/NET0131 ,
		\u1_u2_rd_buf0_reg[8]/NET0131 ,
		_w2040_
	);
	LUT2 #(
		.INIT('h4)
	) name291 (
		_w1765_,
		_w2040_,
		_w2041_
	);
	LUT3 #(
		.INIT('h20)
	) name292 (
		\u1_u2_rd_buf1_reg[24]/NET0131 ,
		_w1762_,
		_w1763_,
		_w2042_
	);
	LUT4 #(
		.INIT('h4000)
	) name293 (
		\u1_u2_adr_cb_reg[0]/NET0131 ,
		\u1_u2_adr_cb_reg[1]/NET0131 ,
		\u1_u2_adr_cb_reg[2]/NET0131 ,
		\u1_u2_rd_buf1_reg[24]/NET0131 ,
		_w2043_
	);
	LUT2 #(
		.INIT('h4)
	) name294 (
		_w1765_,
		_w2043_,
		_w2044_
	);
	LUT4 #(
		.INIT('h0001)
	) name295 (
		_w2039_,
		_w2041_,
		_w2042_,
		_w2044_,
		_w2045_
	);
	LUT3 #(
		.INIT('h20)
	) name296 (
		\u1_u2_rd_buf0_reg[0]/NET0131 ,
		_w1762_,
		_w1796_,
		_w2046_
	);
	LUT4 #(
		.INIT('h8000)
	) name297 (
		\u1_u2_adr_cb_reg[0]/NET0131 ,
		\u1_u2_adr_cb_reg[1]/NET0131 ,
		\u1_u2_adr_cb_reg[2]/NET0131 ,
		\u1_u2_rd_buf0_reg[0]/NET0131 ,
		_w2047_
	);
	LUT2 #(
		.INIT('h4)
	) name298 (
		_w1765_,
		_w2047_,
		_w2048_
	);
	LUT3 #(
		.INIT('h20)
	) name299 (
		\u1_u2_rd_buf1_reg[16]/NET0131 ,
		_w1762_,
		_w1778_,
		_w2049_
	);
	LUT4 #(
		.INIT('h2000)
	) name300 (
		\u1_u2_adr_cb_reg[0]/NET0131 ,
		\u1_u2_adr_cb_reg[1]/NET0131 ,
		\u1_u2_adr_cb_reg[2]/NET0131 ,
		\u1_u2_rd_buf1_reg[16]/NET0131 ,
		_w2050_
	);
	LUT2 #(
		.INIT('h4)
	) name301 (
		_w1765_,
		_w2050_,
		_w2051_
	);
	LUT4 #(
		.INIT('h0001)
	) name302 (
		_w2046_,
		_w2048_,
		_w2049_,
		_w2051_,
		_w2052_
	);
	LUT4 #(
		.INIT('h8000)
	) name303 (
		_w2031_,
		_w2038_,
		_w2045_,
		_w2052_,
		_w2053_
	);
	LUT2 #(
		.INIT('h9)
	) name304 (
		\u1_u1_crc16_reg[15]/P0001 ,
		_w2053_,
		_w2054_
	);
	LUT4 #(
		.INIT('h4000)
	) name305 (
		\u1_u2_adr_cb_reg[0]/NET0131 ,
		\u1_u2_adr_cb_reg[1]/NET0131 ,
		\u1_u2_adr_cb_reg[2]/NET0131 ,
		\u1_u2_rd_buf1_reg[25]/NET0131 ,
		_w2055_
	);
	LUT2 #(
		.INIT('h4)
	) name306 (
		_w1765_,
		_w2055_,
		_w2056_
	);
	LUT3 #(
		.INIT('h20)
	) name307 (
		\u1_u2_rd_buf1_reg[25]/NET0131 ,
		_w1762_,
		_w1763_,
		_w2057_
	);
	LUT3 #(
		.INIT('h20)
	) name308 (
		\u1_u2_rd_buf1_reg[9]/NET0131 ,
		_w1762_,
		_w1769_,
		_w2058_
	);
	LUT4 #(
		.INIT('h1000)
	) name309 (
		\u1_u2_adr_cb_reg[0]/NET0131 ,
		\u1_u2_adr_cb_reg[1]/NET0131 ,
		\u1_u2_adr_cb_reg[2]/NET0131 ,
		\u1_u2_rd_buf1_reg[9]/NET0131 ,
		_w2059_
	);
	LUT2 #(
		.INIT('h4)
	) name310 (
		_w1765_,
		_w2059_,
		_w2060_
	);
	LUT4 #(
		.INIT('h0001)
	) name311 (
		_w2056_,
		_w2057_,
		_w2058_,
		_w2060_,
		_w2061_
	);
	LUT3 #(
		.INIT('h20)
	) name312 (
		\u1_u2_rd_buf1_reg[17]/NET0131 ,
		_w1762_,
		_w1778_,
		_w2062_
	);
	LUT4 #(
		.INIT('h2000)
	) name313 (
		\u1_u2_adr_cb_reg[0]/NET0131 ,
		\u1_u2_adr_cb_reg[1]/NET0131 ,
		\u1_u2_adr_cb_reg[2]/NET0131 ,
		\u1_u2_rd_buf1_reg[17]/NET0131 ,
		_w2063_
	);
	LUT2 #(
		.INIT('h4)
	) name314 (
		_w1765_,
		_w2063_,
		_w2064_
	);
	LUT3 #(
		.INIT('h20)
	) name315 (
		\u1_u2_rd_buf1_reg[1]/NET0131 ,
		_w1762_,
		_w1774_,
		_w2065_
	);
	LUT4 #(
		.INIT('h0800)
	) name316 (
		\u1_u2_adr_cb_reg[0]/NET0131 ,
		\u1_u2_adr_cb_reg[1]/NET0131 ,
		\u1_u2_adr_cb_reg[2]/NET0131 ,
		\u1_u2_rd_buf1_reg[1]/NET0131 ,
		_w2066_
	);
	LUT2 #(
		.INIT('h4)
	) name317 (
		_w1765_,
		_w2066_,
		_w2067_
	);
	LUT4 #(
		.INIT('h0001)
	) name318 (
		_w2062_,
		_w2064_,
		_w2065_,
		_w2067_,
		_w2068_
	);
	LUT3 #(
		.INIT('h20)
	) name319 (
		\u1_u2_rd_buf0_reg[9]/NET0131 ,
		_w1762_,
		_w1787_,
		_w2069_
	);
	LUT4 #(
		.INIT('h0100)
	) name320 (
		\u1_u2_adr_cb_reg[0]/NET0131 ,
		\u1_u2_adr_cb_reg[1]/NET0131 ,
		\u1_u2_adr_cb_reg[2]/NET0131 ,
		\u1_u2_rd_buf0_reg[9]/NET0131 ,
		_w2070_
	);
	LUT2 #(
		.INIT('h4)
	) name321 (
		_w1765_,
		_w2070_,
		_w2071_
	);
	LUT3 #(
		.INIT('h20)
	) name322 (
		\u1_u2_rd_buf0_reg[25]/NET0131 ,
		_w1762_,
		_w1783_,
		_w2072_
	);
	LUT4 #(
		.INIT('h0400)
	) name323 (
		\u1_u2_adr_cb_reg[0]/NET0131 ,
		\u1_u2_adr_cb_reg[1]/NET0131 ,
		\u1_u2_adr_cb_reg[2]/NET0131 ,
		\u1_u2_rd_buf0_reg[25]/NET0131 ,
		_w2073_
	);
	LUT2 #(
		.INIT('h4)
	) name324 (
		_w1765_,
		_w2073_,
		_w2074_
	);
	LUT4 #(
		.INIT('h0001)
	) name325 (
		_w2069_,
		_w2071_,
		_w2072_,
		_w2074_,
		_w2075_
	);
	LUT3 #(
		.INIT('h20)
	) name326 (
		\u1_u2_rd_buf0_reg[17]/NET0131 ,
		_w1762_,
		_w1792_,
		_w2076_
	);
	LUT4 #(
		.INIT('h0200)
	) name327 (
		\u1_u2_adr_cb_reg[0]/NET0131 ,
		\u1_u2_adr_cb_reg[1]/NET0131 ,
		\u1_u2_adr_cb_reg[2]/NET0131 ,
		\u1_u2_rd_buf0_reg[17]/NET0131 ,
		_w2077_
	);
	LUT2 #(
		.INIT('h4)
	) name328 (
		_w1765_,
		_w2077_,
		_w2078_
	);
	LUT3 #(
		.INIT('h20)
	) name329 (
		\u1_u2_rd_buf0_reg[1]/NET0131 ,
		_w1762_,
		_w1796_,
		_w2079_
	);
	LUT4 #(
		.INIT('h8000)
	) name330 (
		\u1_u2_adr_cb_reg[0]/NET0131 ,
		\u1_u2_adr_cb_reg[1]/NET0131 ,
		\u1_u2_adr_cb_reg[2]/NET0131 ,
		\u1_u2_rd_buf0_reg[1]/NET0131 ,
		_w2080_
	);
	LUT2 #(
		.INIT('h4)
	) name331 (
		_w1765_,
		_w2080_,
		_w2081_
	);
	LUT4 #(
		.INIT('h0001)
	) name332 (
		_w2076_,
		_w2078_,
		_w2079_,
		_w2081_,
		_w2082_
	);
	LUT4 #(
		.INIT('h8000)
	) name333 (
		_w2061_,
		_w2068_,
		_w2075_,
		_w2082_,
		_w2083_
	);
	LUT2 #(
		.INIT('h9)
	) name334 (
		\u1_u1_crc16_reg[10]/P0001 ,
		\u1_u1_crc16_reg[9]/P0001 ,
		_w2084_
	);
	LUT2 #(
		.INIT('h9)
	) name335 (
		\u1_u1_crc16_reg[11]/P0001 ,
		\u1_u1_crc16_reg[12]/P0001 ,
		_w2085_
	);
	LUT4 #(
		.INIT('h4182)
	) name336 (
		\u1_u1_crc16_reg[10]/P0001 ,
		\u1_u1_crc16_reg[11]/P0001 ,
		\u1_u1_crc16_reg[12]/P0001 ,
		\u1_u1_crc16_reg[9]/P0001 ,
		_w2086_
	);
	LUT4 #(
		.INIT('h69ff)
	) name337 (
		\u1_u1_crc16_reg[15]/P0001 ,
		_w2053_,
		_w2083_,
		_w2086_,
		_w2087_
	);
	LUT4 #(
		.INIT('h8241)
	) name338 (
		\u1_u1_crc16_reg[10]/P0001 ,
		\u1_u1_crc16_reg[11]/P0001 ,
		\u1_u1_crc16_reg[12]/P0001 ,
		\u1_u1_crc16_reg[9]/P0001 ,
		_w2088_
	);
	LUT4 #(
		.INIT('h96ff)
	) name339 (
		\u1_u1_crc16_reg[15]/P0001 ,
		_w2053_,
		_w2083_,
		_w2088_,
		_w2089_
	);
	LUT4 #(
		.INIT('h1428)
	) name340 (
		\u1_u1_crc16_reg[10]/P0001 ,
		\u1_u1_crc16_reg[11]/P0001 ,
		\u1_u1_crc16_reg[12]/P0001 ,
		\u1_u1_crc16_reg[9]/P0001 ,
		_w2090_
	);
	LUT4 #(
		.INIT('h96ff)
	) name341 (
		\u1_u1_crc16_reg[15]/P0001 ,
		_w2053_,
		_w2083_,
		_w2090_,
		_w2091_
	);
	LUT4 #(
		.INIT('h2814)
	) name342 (
		\u1_u1_crc16_reg[10]/P0001 ,
		\u1_u1_crc16_reg[11]/P0001 ,
		\u1_u1_crc16_reg[12]/P0001 ,
		\u1_u1_crc16_reg[9]/P0001 ,
		_w2092_
	);
	LUT4 #(
		.INIT('h69ff)
	) name343 (
		\u1_u1_crc16_reg[15]/P0001 ,
		_w2053_,
		_w2083_,
		_w2092_,
		_w2093_
	);
	LUT4 #(
		.INIT('h8000)
	) name344 (
		_w2087_,
		_w2089_,
		_w2091_,
		_w2093_,
		_w2094_
	);
	LUT3 #(
		.INIT('h04)
	) name345 (
		\u1_u1_send_data_r2_reg/P0001 ,
		\u1_u1_send_data_r_reg/P0001 ,
		\u1_u1_zero_length_r_reg/P0001 ,
		_w2095_
	);
	LUT4 #(
		.INIT('h00df)
	) name346 (
		_w1762_,
		_w1805_,
		_w1820_,
		_w2095_,
		_w2096_
	);
	LUT4 #(
		.INIT('h0069)
	) name347 (
		_w2023_,
		_w2024_,
		_w2094_,
		_w2096_,
		_w2097_
	);
	LUT3 #(
		.INIT('h54)
	) name348 (
		\u1_u1_send_data_r_reg/P0001 ,
		\u1_u1_send_zero_length_r_reg/P0001 ,
		\u1_u2_send_data_r_reg/NET0131 ,
		_w2098_
	);
	LUT4 #(
		.INIT('haa8a)
	) name349 (
		\u1_u1_crc16_reg[15]/P0001 ,
		\u1_u1_send_data_r2_reg/P0001 ,
		\u1_u1_send_data_r_reg/P0001 ,
		\u1_u1_zero_length_r_reg/P0001 ,
		_w2099_
	);
	LUT4 #(
		.INIT('hdf00)
	) name350 (
		_w1762_,
		_w1805_,
		_w1820_,
		_w2099_,
		_w2100_
	);
	LUT2 #(
		.INIT('h1)
	) name351 (
		_w2098_,
		_w2100_,
		_w2101_
	);
	LUT2 #(
		.INIT('hb)
	) name352 (
		_w2097_,
		_w2101_,
		_w2102_
	);
	LUT4 #(
		.INIT('h6996)
	) name353 (
		_w1801_,
		_w1905_,
		_w2053_,
		_w2083_,
		_w2103_
	);
	LUT2 #(
		.INIT('h9)
	) name354 (
		\u1_u1_crc16_reg[10]/P0001 ,
		\u1_u1_crc16_reg[11]/P0001 ,
		_w2104_
	);
	LUT3 #(
		.INIT('h96)
	) name355 (
		\u1_u1_crc16_reg[10]/P0001 ,
		\u1_u1_crc16_reg[11]/P0001 ,
		\u1_u1_crc16_reg[9]/P0001 ,
		_w2105_
	);
	LUT2 #(
		.INIT('h6)
	) name356 (
		_w1990_,
		_w2105_,
		_w2106_
	);
	LUT2 #(
		.INIT('h9)
	) name357 (
		\u1_u1_crc16_reg[12]/P0001 ,
		\u1_u1_crc16_reg[13]/P0001 ,
		_w2107_
	);
	LUT4 #(
		.INIT('h6996)
	) name358 (
		\u1_u1_crc16_reg[12]/P0001 ,
		\u1_u1_crc16_reg[13]/P0001 ,
		\u1_u1_crc16_reg[14]/P0001 ,
		\u1_u1_crc16_reg[15]/P0001 ,
		_w2108_
	);
	LUT3 #(
		.INIT('h96)
	) name359 (
		_w1957_,
		_w2019_,
		_w2108_,
		_w2109_
	);
	LUT4 #(
		.INIT('h1441)
	) name360 (
		_w2096_,
		_w2103_,
		_w2106_,
		_w2109_,
		_w2110_
	);
	LUT4 #(
		.INIT('haa8a)
	) name361 (
		\u1_u1_crc16_reg[1]/P0001 ,
		\u1_u1_send_data_r2_reg/P0001 ,
		\u1_u1_send_data_r_reg/P0001 ,
		\u1_u1_zero_length_r_reg/P0001 ,
		_w2111_
	);
	LUT4 #(
		.INIT('hdf00)
	) name362 (
		_w1762_,
		_w1805_,
		_w1820_,
		_w2111_,
		_w2112_
	);
	LUT2 #(
		.INIT('h1)
	) name363 (
		_w2098_,
		_w2112_,
		_w2113_
	);
	LUT2 #(
		.INIT('hb)
	) name364 (
		_w2110_,
		_w2113_,
		_w2114_
	);
	LUT4 #(
		.INIT('h0200)
	) name365 (
		\u1_u0_pid_reg[0]/NET0131 ,
		\u1_u0_pid_reg[1]/NET0131 ,
		\u1_u0_pid_reg[2]/NET0131 ,
		\u1_u0_pid_reg[3]/NET0131 ,
		_w2115_
	);
	LUT4 #(
		.INIT('h0002)
	) name366 (
		\u1_u0_pid_reg[0]/NET0131 ,
		\u1_u0_pid_reg[1]/NET0131 ,
		\u1_u0_pid_reg[2]/NET0131 ,
		\u1_u0_pid_reg[3]/NET0131 ,
		_w2116_
	);
	LUT4 #(
		.INIT('h153f)
	) name367 (
		\u1_u3_buf0_na_reg/NET0131 ,
		\u1_u3_buf1_na_reg/NET0131 ,
		_w2115_,
		_w2116_,
		_w2117_
	);
	LUT2 #(
		.INIT('h1)
	) name368 (
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		_w2118_
	);
	LUT2 #(
		.INIT('h8)
	) name369 (
		\u1_u3_buf0_na_reg/NET0131 ,
		\u1_u3_buf1_na_reg/NET0131 ,
		_w2119_
	);
	LUT2 #(
		.INIT('h4)
	) name370 (
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		_w2120_
	);
	LUT4 #(
		.INIT('hfdb9)
	) name371 (
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		\u4_dma_in_buf_sz1_reg/P0001 ,
		\u4_dma_out_buf_avail_reg/P0001 ,
		_w2121_
	);
	LUT3 #(
		.INIT('ha8)
	) name372 (
		\u4_csr_reg[15]/NET0131 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		_w2122_
	);
	LUT2 #(
		.INIT('h4)
	) name373 (
		_w2121_,
		_w2122_,
		_w2123_
	);
	LUT3 #(
		.INIT('h45)
	) name374 (
		_w2119_,
		_w2121_,
		_w2122_,
		_w2124_
	);
	LUT3 #(
		.INIT('hb0)
	) name375 (
		_w2117_,
		_w2118_,
		_w2124_,
		_w2125_
	);
	LUT2 #(
		.INIT('h1)
	) name376 (
		\u1_u3_state_reg[7]/P0001 ,
		\u1_u3_state_reg[9]/P0001 ,
		_w2126_
	);
	LUT4 #(
		.INIT('h0001)
	) name377 (
		\u1_u3_state_reg[6]/P0001 ,
		\u1_u3_state_reg[7]/P0001 ,
		\u1_u3_state_reg[8]/P0001 ,
		\u1_u3_state_reg[9]/P0001 ,
		_w2127_
	);
	LUT4 #(
		.INIT('h0001)
	) name378 (
		\u1_u3_state_reg[2]/P0001 ,
		\u1_u3_state_reg[3]/P0001 ,
		\u1_u3_state_reg[4]/P0001 ,
		\u1_u3_state_reg[5]/P0001 ,
		_w2128_
	);
	LUT2 #(
		.INIT('h8)
	) name379 (
		_w2127_,
		_w2128_,
		_w2129_
	);
	LUT2 #(
		.INIT('h2)
	) name380 (
		\u1_u3_match_r_reg/P0001 ,
		\u1_u3_state_reg[1]/P0001 ,
		_w2130_
	);
	LUT4 #(
		.INIT('h0020)
	) name381 (
		\u1_u0_pid_reg[0]/NET0131 ,
		\u1_u0_pid_reg[1]/NET0131 ,
		\u1_u0_pid_reg[2]/NET0131 ,
		\u1_u0_pid_reg[3]/NET0131 ,
		_w2131_
	);
	LUT4 #(
		.INIT('h0080)
	) name382 (
		_w2127_,
		_w2128_,
		_w2130_,
		_w2131_,
		_w2132_
	);
	LUT2 #(
		.INIT('h4)
	) name383 (
		\u4_csr_reg[22]/P0001 ,
		\u4_csr_reg[23]/P0001 ,
		_w2133_
	);
	LUT3 #(
		.INIT('h51)
	) name384 (
		\u1_u3_state_reg[6]/P0001 ,
		\u4_csr_reg[22]/P0001 ,
		\u4_csr_reg[23]/P0001 ,
		_w2134_
	);
	LUT3 #(
		.INIT('h41)
	) name385 (
		\u1_u3_state_reg[6]/P0001 ,
		\u4_csr_reg[22]/P0001 ,
		\u4_csr_reg[23]/P0001 ,
		_w2135_
	);
	LUT2 #(
		.INIT('h8)
	) name386 (
		_w2132_,
		_w2135_,
		_w2136_
	);
	LUT2 #(
		.INIT('h1)
	) name387 (
		\u1_u3_to_large_reg/P0001 ,
		\u1_u3_to_small_reg/P0001 ,
		_w2137_
	);
	LUT4 #(
		.INIT('h0080)
	) name388 (
		\u0_u0_mode_hs_reg/P0001 ,
		\u1_u3_no_bufs0_reg/P0001 ,
		\u1_u3_no_bufs1_reg/P0001 ,
		\u1_u3_pid_seq_err_reg/P0001 ,
		_w2138_
	);
	LUT2 #(
		.INIT('h4)
	) name389 (
		\u1_u3_abort_reg/P0001 ,
		\u1_u3_state_reg[6]/P0001 ,
		_w2139_
	);
	LUT3 #(
		.INIT('hd0)
	) name390 (
		_w2137_,
		_w2138_,
		_w2139_,
		_w2140_
	);
	LUT3 #(
		.INIT('hf4)
	) name391 (
		_w2125_,
		_w2136_,
		_w2140_,
		_w2141_
	);
	LUT4 #(
		.INIT('h6996)
	) name392 (
		\u1_u1_crc16_reg[10]/P0001 ,
		\u1_u1_crc16_reg[11]/P0001 ,
		\u1_u1_crc16_reg[8]/P0001 ,
		\u1_u1_crc16_reg[9]/P0001 ,
		_w2142_
	);
	LUT4 #(
		.INIT('h9009)
	) name393 (
		_w2020_,
		_w2103_,
		_w2108_,
		_w2142_,
		_w2143_
	);
	LUT2 #(
		.INIT('h9)
	) name394 (
		_w2108_,
		_w2142_,
		_w2144_
	);
	LUT4 #(
		.INIT('h3321)
	) name395 (
		_w2020_,
		_w2096_,
		_w2103_,
		_w2144_,
		_w2145_
	);
	LUT4 #(
		.INIT('haa8a)
	) name396 (
		\u1_u1_crc16_reg[0]/P0001 ,
		\u1_u1_send_data_r2_reg/P0001 ,
		\u1_u1_send_data_r_reg/P0001 ,
		\u1_u1_zero_length_r_reg/P0001 ,
		_w2146_
	);
	LUT4 #(
		.INIT('hdf00)
	) name397 (
		_w1762_,
		_w1805_,
		_w1820_,
		_w2146_,
		_w2147_
	);
	LUT2 #(
		.INIT('h1)
	) name398 (
		_w2098_,
		_w2147_,
		_w2148_
	);
	LUT3 #(
		.INIT('h4f)
	) name399 (
		_w2143_,
		_w2145_,
		_w2148_,
		_w2149_
	);
	LUT4 #(
		.INIT('h0200)
	) name400 (
		\u1_u3_match_r_reg/P0001 ,
		\u1_u3_state_reg[1]/P0001 ,
		\u4_csr_reg[22]/P0001 ,
		\u4_csr_reg[23]/P0001 ,
		_w2150_
	);
	LUT4 #(
		.INIT('h0800)
	) name401 (
		_w2127_,
		_w2128_,
		_w2131_,
		_w2150_,
		_w2151_
	);
	LUT4 #(
		.INIT('h0004)
	) name402 (
		\u1_u3_abort_reg/P0001 ,
		\u1_u3_state_reg[6]/P0001 ,
		\u1_u3_to_large_reg/P0001 ,
		\u1_u3_to_small_reg/P0001 ,
		_w2152_
	);
	LUT2 #(
		.INIT('h8)
	) name403 (
		_w2138_,
		_w2152_,
		_w2153_
	);
	LUT2 #(
		.INIT('he)
	) name404 (
		_w2151_,
		_w2153_,
		_w2154_
	);
	LUT4 #(
		.INIT('hdeed)
	) name405 (
		\u1_u1_crc16_reg[0]/P0001 ,
		\u1_u1_crc16_reg[14]/P0001 ,
		_w2054_,
		_w2083_,
		_w2155_
	);
	LUT4 #(
		.INIT('hb77b)
	) name406 (
		\u1_u1_crc16_reg[0]/P0001 ,
		\u1_u1_crc16_reg[14]/P0001 ,
		_w2054_,
		_w2083_,
		_w2156_
	);
	LUT4 #(
		.INIT('haa8a)
	) name407 (
		\u1_u1_crc16_reg[8]/P0001 ,
		\u1_u1_send_data_r2_reg/P0001 ,
		\u1_u1_send_data_r_reg/P0001 ,
		\u1_u1_zero_length_r_reg/P0001 ,
		_w2157_
	);
	LUT4 #(
		.INIT('hdf00)
	) name408 (
		_w1762_,
		_w1805_,
		_w1820_,
		_w2157_,
		_w2158_
	);
	LUT2 #(
		.INIT('h1)
	) name409 (
		_w2098_,
		_w2158_,
		_w2159_
	);
	LUT4 #(
		.INIT('h40ff)
	) name410 (
		_w2096_,
		_w2155_,
		_w2156_,
		_w2159_,
		_w2160_
	);
	LUT2 #(
		.INIT('h8)
	) name411 (
		\u1_u1_crc16_reg[8]/P0001 ,
		\u1_u1_crc16_reg[9]/P0001 ,
		_w2161_
	);
	LUT3 #(
		.INIT('h90)
	) name412 (
		_w1870_,
		_w1957_,
		_w2161_,
		_w2162_
	);
	LUT2 #(
		.INIT('h1)
	) name413 (
		\u1_u1_crc16_reg[8]/P0001 ,
		\u1_u1_crc16_reg[9]/P0001 ,
		_w2163_
	);
	LUT4 #(
		.INIT('h060f)
	) name414 (
		_w1870_,
		_w1957_,
		_w2096_,
		_w2163_,
		_w2164_
	);
	LUT4 #(
		.INIT('hf99f)
	) name415 (
		\u1_u1_crc16_reg[8]/P0001 ,
		\u1_u1_crc16_reg[9]/P0001 ,
		_w1870_,
		_w1957_,
		_w2165_
	);
	LUT4 #(
		.INIT('haa8a)
	) name416 (
		\u1_u1_crc16_reg[2]/P0001 ,
		\u1_u1_send_data_r2_reg/P0001 ,
		\u1_u1_send_data_r_reg/P0001 ,
		\u1_u1_zero_length_r_reg/P0001 ,
		_w2166_
	);
	LUT4 #(
		.INIT('hdf00)
	) name417 (
		_w1762_,
		_w1805_,
		_w1820_,
		_w2166_,
		_w2167_
	);
	LUT2 #(
		.INIT('h1)
	) name418 (
		_w2098_,
		_w2167_,
		_w2168_
	);
	LUT4 #(
		.INIT('h40ff)
	) name419 (
		_w2162_,
		_w2164_,
		_w2165_,
		_w2168_,
		_w2169_
	);
	LUT2 #(
		.INIT('h8)
	) name420 (
		_w2084_,
		_w2095_,
		_w2170_
	);
	LUT2 #(
		.INIT('h8)
	) name421 (
		_w1762_,
		_w2084_,
		_w2171_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name422 (
		_w1805_,
		_w1820_,
		_w2170_,
		_w2171_,
		_w2172_
	);
	LUT3 #(
		.INIT('h06)
	) name423 (
		_w1957_,
		_w2019_,
		_w2172_,
		_w2173_
	);
	LUT2 #(
		.INIT('h4)
	) name424 (
		_w2084_,
		_w2095_,
		_w2174_
	);
	LUT2 #(
		.INIT('h2)
	) name425 (
		_w1762_,
		_w2084_,
		_w2175_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name426 (
		_w1805_,
		_w1820_,
		_w2174_,
		_w2175_,
		_w2176_
	);
	LUT4 #(
		.INIT('haa8a)
	) name427 (
		\u1_u1_crc16_reg[3]/P0001 ,
		\u1_u1_send_data_r2_reg/P0001 ,
		\u1_u1_send_data_r_reg/P0001 ,
		\u1_u1_zero_length_r_reg/P0001 ,
		_w2177_
	);
	LUT4 #(
		.INIT('hdf00)
	) name428 (
		_w1762_,
		_w1805_,
		_w1820_,
		_w2177_,
		_w2178_
	);
	LUT2 #(
		.INIT('h1)
	) name429 (
		_w2098_,
		_w2178_,
		_w2179_
	);
	LUT4 #(
		.INIT('hf600)
	) name430 (
		_w1957_,
		_w2019_,
		_w2176_,
		_w2179_,
		_w2180_
	);
	LUT2 #(
		.INIT('hb)
	) name431 (
		_w2173_,
		_w2180_,
		_w2181_
	);
	LUT2 #(
		.INIT('h1)
	) name432 (
		_w2096_,
		_w2104_,
		_w2182_
	);
	LUT2 #(
		.INIT('h8)
	) name433 (
		_w2095_,
		_w2104_,
		_w2183_
	);
	LUT2 #(
		.INIT('h8)
	) name434 (
		_w1762_,
		_w2104_,
		_w2184_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name435 (
		_w1805_,
		_w1820_,
		_w2183_,
		_w2184_,
		_w2185_
	);
	LUT4 #(
		.INIT('h6f09)
	) name436 (
		_w1990_,
		_w2019_,
		_w2182_,
		_w2185_,
		_w2186_
	);
	LUT4 #(
		.INIT('haa8a)
	) name437 (
		\u1_u1_crc16_reg[4]/P0001 ,
		\u1_u1_send_data_r2_reg/P0001 ,
		\u1_u1_send_data_r_reg/P0001 ,
		\u1_u1_zero_length_r_reg/P0001 ,
		_w2187_
	);
	LUT4 #(
		.INIT('hdf00)
	) name438 (
		_w1762_,
		_w1805_,
		_w1820_,
		_w2187_,
		_w2188_
	);
	LUT2 #(
		.INIT('h1)
	) name439 (
		_w2098_,
		_w2188_,
		_w2189_
	);
	LUT2 #(
		.INIT('h7)
	) name440 (
		_w2186_,
		_w2189_,
		_w2190_
	);
	LUT2 #(
		.INIT('h8)
	) name441 (
		_w2085_,
		_w2095_,
		_w2191_
	);
	LUT2 #(
		.INIT('h8)
	) name442 (
		_w1762_,
		_w2085_,
		_w2192_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name443 (
		_w1805_,
		_w1820_,
		_w2191_,
		_w2192_,
		_w2193_
	);
	LUT3 #(
		.INIT('h06)
	) name444 (
		_w1801_,
		_w1990_,
		_w2193_,
		_w2194_
	);
	LUT2 #(
		.INIT('h4)
	) name445 (
		_w2085_,
		_w2095_,
		_w2195_
	);
	LUT2 #(
		.INIT('h2)
	) name446 (
		_w1762_,
		_w2085_,
		_w2196_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name447 (
		_w1805_,
		_w1820_,
		_w2195_,
		_w2196_,
		_w2197_
	);
	LUT4 #(
		.INIT('haa8a)
	) name448 (
		\u1_u1_crc16_reg[5]/P0001 ,
		\u1_u1_send_data_r2_reg/P0001 ,
		\u1_u1_send_data_r_reg/P0001 ,
		\u1_u1_zero_length_r_reg/P0001 ,
		_w2198_
	);
	LUT4 #(
		.INIT('hdf00)
	) name449 (
		_w1762_,
		_w1805_,
		_w1820_,
		_w2198_,
		_w2199_
	);
	LUT2 #(
		.INIT('h1)
	) name450 (
		_w2098_,
		_w2199_,
		_w2200_
	);
	LUT4 #(
		.INIT('hf600)
	) name451 (
		_w1801_,
		_w1990_,
		_w2197_,
		_w2200_,
		_w2201_
	);
	LUT2 #(
		.INIT('hb)
	) name452 (
		_w2194_,
		_w2201_,
		_w2202_
	);
	LUT2 #(
		.INIT('h1)
	) name453 (
		_w2096_,
		_w2107_,
		_w2203_
	);
	LUT2 #(
		.INIT('h8)
	) name454 (
		_w2095_,
		_w2107_,
		_w2204_
	);
	LUT2 #(
		.INIT('h8)
	) name455 (
		_w1762_,
		_w2107_,
		_w2205_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name456 (
		_w1805_,
		_w1820_,
		_w2204_,
		_w2205_,
		_w2206_
	);
	LUT4 #(
		.INIT('h6f09)
	) name457 (
		_w1801_,
		_w1905_,
		_w2203_,
		_w2206_,
		_w2207_
	);
	LUT4 #(
		.INIT('haa8a)
	) name458 (
		\u1_u1_crc16_reg[6]/P0001 ,
		\u1_u1_send_data_r2_reg/P0001 ,
		\u1_u1_send_data_r_reg/P0001 ,
		\u1_u1_zero_length_r_reg/P0001 ,
		_w2208_
	);
	LUT4 #(
		.INIT('hdf00)
	) name459 (
		_w1762_,
		_w1805_,
		_w1820_,
		_w2208_,
		_w2209_
	);
	LUT2 #(
		.INIT('h1)
	) name460 (
		_w2098_,
		_w2209_,
		_w2210_
	);
	LUT2 #(
		.INIT('h7)
	) name461 (
		_w2207_,
		_w2210_,
		_w2211_
	);
	LUT4 #(
		.INIT('h0096)
	) name462 (
		_w1905_,
		_w2024_,
		_w2083_,
		_w2096_,
		_w2212_
	);
	LUT4 #(
		.INIT('haa8a)
	) name463 (
		\u1_u1_crc16_reg[7]/P0001 ,
		\u1_u1_send_data_r2_reg/P0001 ,
		\u1_u1_send_data_r_reg/P0001 ,
		\u1_u1_zero_length_r_reg/P0001 ,
		_w2213_
	);
	LUT4 #(
		.INIT('hdf00)
	) name464 (
		_w1762_,
		_w1805_,
		_w1820_,
		_w2213_,
		_w2214_
	);
	LUT2 #(
		.INIT('h1)
	) name465 (
		_w2098_,
		_w2214_,
		_w2215_
	);
	LUT2 #(
		.INIT('hb)
	) name466 (
		_w2212_,
		_w2215_,
		_w2216_
	);
	LUT2 #(
		.INIT('h6)
	) name467 (
		\u1_u1_crc16_reg[15]/P0001 ,
		\u1_u1_crc16_reg[1]/P0001 ,
		_w2217_
	);
	LUT2 #(
		.INIT('h1)
	) name468 (
		_w2096_,
		_w2217_,
		_w2218_
	);
	LUT2 #(
		.INIT('h4)
	) name469 (
		_w2096_,
		_w2217_,
		_w2219_
	);
	LUT4 #(
		.INIT('haa8a)
	) name470 (
		\u1_u1_crc16_reg[9]/P0001 ,
		\u1_u1_send_data_r2_reg/P0001 ,
		\u1_u1_send_data_r_reg/P0001 ,
		\u1_u1_zero_length_r_reg/P0001 ,
		_w2220_
	);
	LUT4 #(
		.INIT('hdf00)
	) name471 (
		_w1762_,
		_w1805_,
		_w1820_,
		_w2220_,
		_w2221_
	);
	LUT2 #(
		.INIT('h1)
	) name472 (
		_w2098_,
		_w2221_,
		_w2222_
	);
	LUT4 #(
		.INIT('he4ff)
	) name473 (
		_w2053_,
		_w2218_,
		_w2219_,
		_w2222_,
		_w2223_
	);
	LUT3 #(
		.INIT('h01)
	) name474 (
		\u5_state_reg[3]/P0001 ,
		\u5_state_reg[4]/P0001 ,
		\u5_state_reg[5]/NET0131 ,
		_w2224_
	);
	LUT2 #(
		.INIT('h1)
	) name475 (
		\u5_state_reg[1]/P0001 ,
		\u5_state_reg[2]/P0001 ,
		_w2225_
	);
	LUT3 #(
		.INIT('h01)
	) name476 (
		\u5_state_reg[1]/P0001 ,
		\u5_state_reg[2]/P0001 ,
		\wb_addr_i[17]_pad ,
		_w2226_
	);
	LUT3 #(
		.INIT('h02)
	) name477 (
		\wb_addr_i[4]_pad ,
		\wb_addr_i[7]_pad ,
		\wb_addr_i[8]_pad ,
		_w2227_
	);
	LUT2 #(
		.INIT('h8)
	) name478 (
		\wb_addr_i[5]_pad ,
		\wb_addr_i[6]_pad ,
		_w2228_
	);
	LUT2 #(
		.INIT('h8)
	) name479 (
		\u5_wb_req_s1_reg/P0001 ,
		wb_we_i_pad,
		_w2229_
	);
	LUT4 #(
		.INIT('h8000)
	) name480 (
		\u5_wb_req_s1_reg/P0001 ,
		\wb_addr_i[5]_pad ,
		\wb_addr_i[6]_pad ,
		wb_we_i_pad,
		_w2230_
	);
	LUT4 #(
		.INIT('h8000)
	) name481 (
		_w2224_,
		_w2226_,
		_w2227_,
		_w2230_,
		_w2231_
	);
	LUT2 #(
		.INIT('h4)
	) name482 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w2232_
	);
	LUT3 #(
		.INIT('h40)
	) name483 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_data_i[14]_pad ,
		_w2233_
	);
	LUT3 #(
		.INIT('h2a)
	) name484 (
		rst_i_pad,
		_w2231_,
		_w2233_,
		_w2234_
	);
	LUT2 #(
		.INIT('h8)
	) name485 (
		\u1_u3_buf0_rl_reg/P0001 ,
		\u4_u3_ep_match_r_reg/P0001 ,
		_w2235_
	);
	LUT4 #(
		.INIT('hd8f0)
	) name486 (
		\u1_u3_buf0_set_reg/P0001 ,
		\u1_u3_idin_reg[14]/P0001 ,
		\u4_u3_buf0_reg[14]/P0001 ,
		\u4_u3_ep_match_r_reg/P0001 ,
		_w2236_
	);
	LUT3 #(
		.INIT('hb8)
	) name487 (
		\u4_u3_buf0_orig_reg[14]/P0001 ,
		_w2235_,
		_w2236_,
		_w2237_
	);
	LUT3 #(
		.INIT('h70)
	) name488 (
		_w2231_,
		_w2232_,
		_w2237_,
		_w2238_
	);
	LUT2 #(
		.INIT('hd)
	) name489 (
		_w2234_,
		_w2238_,
		_w2239_
	);
	LUT3 #(
		.INIT('h01)
	) name490 (
		\wb_addr_i[4]_pad ,
		\wb_addr_i[7]_pad ,
		\wb_addr_i[8]_pad ,
		_w2240_
	);
	LUT2 #(
		.INIT('h4)
	) name491 (
		\wb_addr_i[5]_pad ,
		\wb_addr_i[6]_pad ,
		_w2241_
	);
	LUT4 #(
		.INIT('h2000)
	) name492 (
		\u5_wb_req_s1_reg/P0001 ,
		\wb_addr_i[5]_pad ,
		\wb_addr_i[6]_pad ,
		wb_we_i_pad,
		_w2242_
	);
	LUT4 #(
		.INIT('h8000)
	) name493 (
		_w2224_,
		_w2226_,
		_w2240_,
		_w2242_,
		_w2243_
	);
	LUT3 #(
		.INIT('h2a)
	) name494 (
		rst_i_pad,
		_w2233_,
		_w2243_,
		_w2244_
	);
	LUT2 #(
		.INIT('h8)
	) name495 (
		\u1_u3_buf0_rl_reg/P0001 ,
		\u4_u0_ep_match_r_reg/P0001 ,
		_w2245_
	);
	LUT4 #(
		.INIT('hd8f0)
	) name496 (
		\u1_u3_buf0_set_reg/P0001 ,
		\u1_u3_idin_reg[14]/P0001 ,
		\u4_u0_buf0_reg[14]/P0001 ,
		\u4_u0_ep_match_r_reg/P0001 ,
		_w2246_
	);
	LUT3 #(
		.INIT('h20)
	) name497 (
		\u1_u3_buf0_rl_reg/P0001 ,
		\u4_u0_buf0_orig_reg[14]/P0001 ,
		\u4_u0_ep_match_r_reg/P0001 ,
		_w2247_
	);
	LUT3 #(
		.INIT('h0e)
	) name498 (
		_w2245_,
		_w2246_,
		_w2247_,
		_w2248_
	);
	LUT3 #(
		.INIT('h70)
	) name499 (
		_w2232_,
		_w2243_,
		_w2248_,
		_w2249_
	);
	LUT2 #(
		.INIT('hd)
	) name500 (
		_w2244_,
		_w2249_,
		_w2250_
	);
	LUT4 #(
		.INIT('h1000)
	) name501 (
		_w1755_,
		_w1757_,
		_w1803_,
		_w1813_,
		_w2251_
	);
	LUT4 #(
		.INIT('hacaa)
	) name502 (
		\u1_u1_crc16_reg[14]/P0001 ,
		\u1_u1_crc16_reg[6]/P0001 ,
		_w1805_,
		_w1820_,
		_w2252_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name503 (
		_w1758_,
		_w1805_,
		_w1810_,
		_w1816_,
		_w2253_
	);
	LUT3 #(
		.INIT('h45)
	) name504 (
		_w2251_,
		_w2252_,
		_w2253_,
		_w2254_
	);
	LUT4 #(
		.INIT('h2000)
	) name505 (
		_w1758_,
		_w1805_,
		_w1810_,
		_w1816_,
		_w2255_
	);
	LUT4 #(
		.INIT('haf8c)
	) name506 (
		TxReady_pad_i_pad,
		\u1_u1_send_token_r_reg/P0001 ,
		\u1_u1_tx_first_r_reg/P0001 ,
		\u1_u3_send_token_reg/P0001 ,
		_w2256_
	);
	LUT2 #(
		.INIT('h2)
	) name507 (
		\DataOut_pad_o[1]_pad ,
		\u0_u0_drive_k_reg/P0001 ,
		_w2257_
	);
	LUT4 #(
		.INIT('h10fe)
	) name508 (
		_w1755_,
		_w1757_,
		_w1811_,
		_w2257_,
		_w2258_
	);
	LUT4 #(
		.INIT('h73ff)
	) name509 (
		_w2083_,
		_w2254_,
		_w2255_,
		_w2258_,
		_w2259_
	);
	LUT4 #(
		.INIT('h8000)
	) name510 (
		_w2224_,
		_w2226_,
		_w2227_,
		_w2242_,
		_w2260_
	);
	LUT3 #(
		.INIT('h2a)
	) name511 (
		rst_i_pad,
		_w2233_,
		_w2260_,
		_w2261_
	);
	LUT2 #(
		.INIT('h8)
	) name512 (
		\u1_u3_buf0_rl_reg/P0001 ,
		\u4_u1_ep_match_r_reg/P0001 ,
		_w2262_
	);
	LUT4 #(
		.INIT('hd8f0)
	) name513 (
		\u1_u3_buf0_set_reg/P0001 ,
		\u1_u3_idin_reg[14]/P0001 ,
		\u4_u1_buf0_reg[14]/P0001 ,
		\u4_u1_ep_match_r_reg/P0001 ,
		_w2263_
	);
	LUT3 #(
		.INIT('hb8)
	) name514 (
		\u4_u1_buf0_orig_reg[14]/P0001 ,
		_w2262_,
		_w2263_,
		_w2264_
	);
	LUT3 #(
		.INIT('h70)
	) name515 (
		_w2232_,
		_w2260_,
		_w2264_,
		_w2265_
	);
	LUT2 #(
		.INIT('hd)
	) name516 (
		_w2261_,
		_w2265_,
		_w2266_
	);
	LUT4 #(
		.INIT('h8000)
	) name517 (
		_w2224_,
		_w2226_,
		_w2230_,
		_w2240_,
		_w2267_
	);
	LUT3 #(
		.INIT('h2a)
	) name518 (
		rst_i_pad,
		_w2233_,
		_w2267_,
		_w2268_
	);
	LUT2 #(
		.INIT('h8)
	) name519 (
		\u1_u3_buf0_rl_reg/P0001 ,
		\u4_u2_ep_match_r_reg/P0001 ,
		_w2269_
	);
	LUT4 #(
		.INIT('hd8f0)
	) name520 (
		\u1_u3_buf0_set_reg/P0001 ,
		\u1_u3_idin_reg[14]/P0001 ,
		\u4_u2_buf0_reg[14]/P0001 ,
		\u4_u2_ep_match_r_reg/P0001 ,
		_w2270_
	);
	LUT3 #(
		.INIT('hb8)
	) name521 (
		\u4_u2_buf0_orig_reg[14]/P0001 ,
		_w2269_,
		_w2270_,
		_w2271_
	);
	LUT3 #(
		.INIT('h70)
	) name522 (
		_w2232_,
		_w2267_,
		_w2271_,
		_w2272_
	);
	LUT2 #(
		.INIT('hd)
	) name523 (
		_w2268_,
		_w2272_,
		_w2273_
	);
	LUT3 #(
		.INIT('h40)
	) name524 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_data_i[10]_pad ,
		_w2274_
	);
	LUT3 #(
		.INIT('h2a)
	) name525 (
		rst_i_pad,
		_w2231_,
		_w2274_,
		_w2275_
	);
	LUT4 #(
		.INIT('hd8f0)
	) name526 (
		\u1_u3_buf0_set_reg/P0001 ,
		\u1_u3_idin_reg[10]/P0001 ,
		\u4_u3_buf0_reg[10]/P0001 ,
		\u4_u3_ep_match_r_reg/P0001 ,
		_w2276_
	);
	LUT3 #(
		.INIT('hb8)
	) name527 (
		\u4_u3_buf0_orig_reg[10]/P0001 ,
		_w2235_,
		_w2276_,
		_w2277_
	);
	LUT3 #(
		.INIT('h70)
	) name528 (
		_w2231_,
		_w2232_,
		_w2277_,
		_w2278_
	);
	LUT2 #(
		.INIT('hd)
	) name529 (
		_w2275_,
		_w2278_,
		_w2279_
	);
	LUT3 #(
		.INIT('h2a)
	) name530 (
		rst_i_pad,
		_w2243_,
		_w2274_,
		_w2280_
	);
	LUT4 #(
		.INIT('hd8f0)
	) name531 (
		\u1_u3_buf0_set_reg/P0001 ,
		\u1_u3_idin_reg[10]/P0001 ,
		\u4_u0_buf0_reg[10]/P0001 ,
		\u4_u0_ep_match_r_reg/P0001 ,
		_w2281_
	);
	LUT3 #(
		.INIT('hb8)
	) name532 (
		\u4_u0_buf0_orig_reg[10]/P0001 ,
		_w2245_,
		_w2281_,
		_w2282_
	);
	LUT3 #(
		.INIT('h70)
	) name533 (
		_w2232_,
		_w2243_,
		_w2282_,
		_w2283_
	);
	LUT2 #(
		.INIT('hd)
	) name534 (
		_w2280_,
		_w2283_,
		_w2284_
	);
	LUT3 #(
		.INIT('h2a)
	) name535 (
		rst_i_pad,
		_w2260_,
		_w2274_,
		_w2285_
	);
	LUT4 #(
		.INIT('hd8f0)
	) name536 (
		\u1_u3_buf0_set_reg/P0001 ,
		\u1_u3_idin_reg[10]/P0001 ,
		\u4_u1_buf0_reg[10]/P0001 ,
		\u4_u1_ep_match_r_reg/P0001 ,
		_w2286_
	);
	LUT3 #(
		.INIT('hb8)
	) name537 (
		\u4_u1_buf0_orig_reg[10]/P0001 ,
		_w2262_,
		_w2286_,
		_w2287_
	);
	LUT3 #(
		.INIT('h70)
	) name538 (
		_w2232_,
		_w2260_,
		_w2287_,
		_w2288_
	);
	LUT2 #(
		.INIT('hd)
	) name539 (
		_w2285_,
		_w2288_,
		_w2289_
	);
	LUT3 #(
		.INIT('h2a)
	) name540 (
		rst_i_pad,
		_w2267_,
		_w2274_,
		_w2290_
	);
	LUT4 #(
		.INIT('hd8f0)
	) name541 (
		\u1_u3_buf0_set_reg/P0001 ,
		\u1_u3_idin_reg[10]/P0001 ,
		\u4_u2_buf0_reg[10]/P0001 ,
		\u4_u2_ep_match_r_reg/P0001 ,
		_w2291_
	);
	LUT3 #(
		.INIT('hb8)
	) name542 (
		\u4_u2_buf0_orig_reg[10]/P0001 ,
		_w2269_,
		_w2291_,
		_w2292_
	);
	LUT3 #(
		.INIT('h70)
	) name543 (
		_w2232_,
		_w2267_,
		_w2292_,
		_w2293_
	);
	LUT2 #(
		.INIT('hd)
	) name544 (
		_w2290_,
		_w2293_,
		_w2294_
	);
	LUT2 #(
		.INIT('h2)
	) name545 (
		\DataOut_pad_o[0]_pad ,
		\u0_u0_drive_k_reg/P0001 ,
		_w2295_
	);
	LUT3 #(
		.INIT('he0)
	) name546 (
		_w1755_,
		_w1757_,
		_w2295_,
		_w2296_
	);
	LUT4 #(
		.INIT('h0023)
	) name547 (
		TxReady_pad_i_pad,
		\u1_u1_send_token_r_reg/P0001 ,
		\u1_u1_tx_first_r_reg/P0001 ,
		\u1_u3_send_token_reg/P0001 ,
		_w2297_
	);
	LUT2 #(
		.INIT('h4)
	) name548 (
		_w1757_,
		_w2297_,
		_w2298_
	);
	LUT4 #(
		.INIT('hacaa)
	) name549 (
		\u1_u1_crc16_reg[15]/P0001 ,
		\u1_u1_crc16_reg[7]/P0001 ,
		_w1805_,
		_w1820_,
		_w2299_
	);
	LUT3 #(
		.INIT('h54)
	) name550 (
		_w1814_,
		_w1828_,
		_w2299_,
		_w2300_
	);
	LUT4 #(
		.INIT('h20f0)
	) name551 (
		_w1828_,
		_w2053_,
		_w2298_,
		_w2300_,
		_w2301_
	);
	LUT2 #(
		.INIT('he)
	) name552 (
		_w2296_,
		_w2301_,
		_w2302_
	);
	LUT2 #(
		.INIT('h2)
	) name553 (
		\DataOut_pad_o[4]_pad ,
		\u0_u0_drive_k_reg/P0001 ,
		_w2303_
	);
	LUT4 #(
		.INIT('h10fe)
	) name554 (
		_w1755_,
		_w1757_,
		_w1811_,
		_w2303_,
		_w2304_
	);
	LUT4 #(
		.INIT('h4000)
	) name555 (
		_w1805_,
		_w1810_,
		_w1816_,
		_w2304_,
		_w2305_
	);
	LUT4 #(
		.INIT('h00ce)
	) name556 (
		_w1755_,
		_w1757_,
		_w2256_,
		_w2303_,
		_w2306_
	);
	LUT3 #(
		.INIT('h45)
	) name557 (
		\u1_u1_crc16_reg[11]/P0001 ,
		_w1805_,
		_w1820_,
		_w2307_
	);
	LUT3 #(
		.INIT('h20)
	) name558 (
		\u0_tx_ready_reg/NET0131 ,
		\u1_u1_crc16_reg[3]/P0001 ,
		\u1_u1_state_reg[2]/NET0131 ,
		_w2308_
	);
	LUT3 #(
		.INIT('h01)
	) name559 (
		\u1_u1_crc16_reg[3]/P0001 ,
		\u1_u1_state_reg[0]/NET0131 ,
		\u1_u1_state_reg[1]/NET0131 ,
		_w2309_
	);
	LUT3 #(
		.INIT('h13)
	) name560 (
		_w1809_,
		_w2308_,
		_w2309_,
		_w2310_
	);
	LUT4 #(
		.INIT('hf0b0)
	) name561 (
		_w1805_,
		_w1820_,
		_w2304_,
		_w2310_,
		_w2311_
	);
	LUT4 #(
		.INIT('h3233)
	) name562 (
		_w1828_,
		_w2306_,
		_w2307_,
		_w2311_,
		_w2312_
	);
	LUT3 #(
		.INIT('h70)
	) name563 (
		_w1990_,
		_w2305_,
		_w2312_,
		_w2313_
	);
	LUT3 #(
		.INIT('h40)
	) name564 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_data_i[13]_pad ,
		_w2314_
	);
	LUT3 #(
		.INIT('h2a)
	) name565 (
		rst_i_pad,
		_w2231_,
		_w2314_,
		_w2315_
	);
	LUT4 #(
		.INIT('hd8f0)
	) name566 (
		\u1_u3_buf0_set_reg/P0001 ,
		\u1_u3_idin_reg[13]/P0001 ,
		\u4_u3_buf0_reg[13]/P0001 ,
		\u4_u3_ep_match_r_reg/P0001 ,
		_w2316_
	);
	LUT3 #(
		.INIT('hb8)
	) name567 (
		\u4_u3_buf0_orig_reg[13]/P0001 ,
		_w2235_,
		_w2316_,
		_w2317_
	);
	LUT3 #(
		.INIT('h70)
	) name568 (
		_w2231_,
		_w2232_,
		_w2317_,
		_w2318_
	);
	LUT2 #(
		.INIT('hd)
	) name569 (
		_w2315_,
		_w2318_,
		_w2319_
	);
	LUT2 #(
		.INIT('h8)
	) name570 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w2320_
	);
	LUT4 #(
		.INIT('h10f0)
	) name571 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u3_buf1_reg[14]/P0001 ,
		\u4_u3_ep_match_r_reg/P0001 ,
		_w2321_
	);
	LUT4 #(
		.INIT('hc800)
	) name572 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_idin_reg[14]/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u3_ep_match_r_reg/P0001 ,
		_w2322_
	);
	LUT2 #(
		.INIT('h1)
	) name573 (
		_w2321_,
		_w2322_,
		_w2323_
	);
	LUT3 #(
		.INIT('h07)
	) name574 (
		_w2231_,
		_w2320_,
		_w2323_,
		_w2324_
	);
	LUT3 #(
		.INIT('h80)
	) name575 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_data_i[14]_pad ,
		_w2325_
	);
	LUT3 #(
		.INIT('h2a)
	) name576 (
		rst_i_pad,
		_w2231_,
		_w2325_,
		_w2326_
	);
	LUT2 #(
		.INIT('hb)
	) name577 (
		_w2324_,
		_w2326_,
		_w2327_
	);
	LUT3 #(
		.INIT('h2a)
	) name578 (
		rst_i_pad,
		_w2243_,
		_w2314_,
		_w2328_
	);
	LUT4 #(
		.INIT('hd8f0)
	) name579 (
		\u1_u3_buf0_set_reg/P0001 ,
		\u1_u3_idin_reg[13]/P0001 ,
		\u4_u0_buf0_reg[13]/P0001 ,
		\u4_u0_ep_match_r_reg/P0001 ,
		_w2329_
	);
	LUT3 #(
		.INIT('hb8)
	) name580 (
		\u4_u0_buf0_orig_reg[13]/P0001 ,
		_w2245_,
		_w2329_,
		_w2330_
	);
	LUT3 #(
		.INIT('h70)
	) name581 (
		_w2232_,
		_w2243_,
		_w2330_,
		_w2331_
	);
	LUT2 #(
		.INIT('hd)
	) name582 (
		_w2328_,
		_w2331_,
		_w2332_
	);
	LUT4 #(
		.INIT('h10f0)
	) name583 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u0_buf1_reg[14]/P0001 ,
		\u4_u0_ep_match_r_reg/P0001 ,
		_w2333_
	);
	LUT4 #(
		.INIT('hc800)
	) name584 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_idin_reg[14]/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u0_ep_match_r_reg/P0001 ,
		_w2334_
	);
	LUT2 #(
		.INIT('h1)
	) name585 (
		_w2333_,
		_w2334_,
		_w2335_
	);
	LUT3 #(
		.INIT('h07)
	) name586 (
		_w2243_,
		_w2320_,
		_w2335_,
		_w2336_
	);
	LUT3 #(
		.INIT('h2a)
	) name587 (
		rst_i_pad,
		_w2243_,
		_w2325_,
		_w2337_
	);
	LUT2 #(
		.INIT('hb)
	) name588 (
		_w2336_,
		_w2337_,
		_w2338_
	);
	LUT3 #(
		.INIT('h2a)
	) name589 (
		rst_i_pad,
		_w2260_,
		_w2314_,
		_w2339_
	);
	LUT4 #(
		.INIT('hd8f0)
	) name590 (
		\u1_u3_buf0_set_reg/P0001 ,
		\u1_u3_idin_reg[13]/P0001 ,
		\u4_u1_buf0_reg[13]/P0001 ,
		\u4_u1_ep_match_r_reg/P0001 ,
		_w2340_
	);
	LUT3 #(
		.INIT('hb8)
	) name591 (
		\u4_u1_buf0_orig_reg[13]/P0001 ,
		_w2262_,
		_w2340_,
		_w2341_
	);
	LUT3 #(
		.INIT('h70)
	) name592 (
		_w2232_,
		_w2260_,
		_w2341_,
		_w2342_
	);
	LUT2 #(
		.INIT('hd)
	) name593 (
		_w2339_,
		_w2342_,
		_w2343_
	);
	LUT4 #(
		.INIT('h10f0)
	) name594 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u1_buf1_reg[14]/P0001 ,
		\u4_u1_ep_match_r_reg/P0001 ,
		_w2344_
	);
	LUT4 #(
		.INIT('hc800)
	) name595 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_idin_reg[14]/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u1_ep_match_r_reg/P0001 ,
		_w2345_
	);
	LUT2 #(
		.INIT('h1)
	) name596 (
		_w2344_,
		_w2345_,
		_w2346_
	);
	LUT3 #(
		.INIT('h07)
	) name597 (
		_w2260_,
		_w2320_,
		_w2346_,
		_w2347_
	);
	LUT3 #(
		.INIT('h2a)
	) name598 (
		rst_i_pad,
		_w2260_,
		_w2325_,
		_w2348_
	);
	LUT2 #(
		.INIT('hb)
	) name599 (
		_w2347_,
		_w2348_,
		_w2349_
	);
	LUT3 #(
		.INIT('h45)
	) name600 (
		\u1_u3_buf0_na_reg/NET0131 ,
		_w2121_,
		_w2122_,
		_w2350_
	);
	LUT4 #(
		.INIT('h0008)
	) name601 (
		\u1_u3_buf0_st_max_reg/P0001 ,
		\u1_u3_in_token_reg/NET0131 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		_w2351_
	);
	LUT4 #(
		.INIT('h1110)
	) name602 (
		\u1_u3_buf1_na_reg/NET0131 ,
		\u4_csr_reg[15]/NET0131 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		_w2352_
	);
	LUT2 #(
		.INIT('h1)
	) name603 (
		\u1_u3_buf0_na_reg/NET0131 ,
		\u4_csr_reg[30]/NET0131 ,
		_w2353_
	);
	LUT3 #(
		.INIT('hc8)
	) name604 (
		\u1_u3_buf0_na_reg/NET0131 ,
		\u1_u3_buf0_st_max_reg/P0001 ,
		\u4_csr_reg[30]/NET0131 ,
		_w2354_
	);
	LUT3 #(
		.INIT('h15)
	) name605 (
		_w2351_,
		_w2352_,
		_w2354_,
		_w2355_
	);
	LUT3 #(
		.INIT('h02)
	) name606 (
		\u1_u3_in_token_reg/NET0131 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		_w2356_
	);
	LUT3 #(
		.INIT('h0d)
	) name607 (
		_w2352_,
		_w2353_,
		_w2356_,
		_w2357_
	);
	LUT4 #(
		.INIT('h222a)
	) name608 (
		\u1_u3_buffer_full_reg/P0001 ,
		\u4_csr_reg[15]/NET0131 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		_w2358_
	);
	LUT4 #(
		.INIT('h0d00)
	) name609 (
		_w2352_,
		_w2353_,
		_w2356_,
		_w2358_,
		_w2359_
	);
	LUT3 #(
		.INIT('hf7)
	) name610 (
		_w2350_,
		_w2355_,
		_w2359_,
		_w2360_
	);
	LUT3 #(
		.INIT('h2a)
	) name611 (
		rst_i_pad,
		_w2267_,
		_w2314_,
		_w2361_
	);
	LUT4 #(
		.INIT('hd8f0)
	) name612 (
		\u1_u3_buf0_set_reg/P0001 ,
		\u1_u3_idin_reg[13]/P0001 ,
		\u4_u2_buf0_reg[13]/P0001 ,
		\u4_u2_ep_match_r_reg/P0001 ,
		_w2362_
	);
	LUT3 #(
		.INIT('hb8)
	) name613 (
		\u4_u2_buf0_orig_reg[13]/P0001 ,
		_w2269_,
		_w2362_,
		_w2363_
	);
	LUT3 #(
		.INIT('h70)
	) name614 (
		_w2232_,
		_w2267_,
		_w2363_,
		_w2364_
	);
	LUT2 #(
		.INIT('hd)
	) name615 (
		_w2361_,
		_w2364_,
		_w2365_
	);
	LUT4 #(
		.INIT('h10f0)
	) name616 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u2_buf1_reg[14]/P0001 ,
		\u4_u2_ep_match_r_reg/P0001 ,
		_w2366_
	);
	LUT4 #(
		.INIT('hc800)
	) name617 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_idin_reg[14]/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u2_ep_match_r_reg/P0001 ,
		_w2367_
	);
	LUT2 #(
		.INIT('h1)
	) name618 (
		_w2366_,
		_w2367_,
		_w2368_
	);
	LUT3 #(
		.INIT('h07)
	) name619 (
		_w2267_,
		_w2320_,
		_w2368_,
		_w2369_
	);
	LUT3 #(
		.INIT('h2a)
	) name620 (
		rst_i_pad,
		_w2267_,
		_w2325_,
		_w2370_
	);
	LUT2 #(
		.INIT('hb)
	) name621 (
		_w2369_,
		_w2370_,
		_w2371_
	);
	LUT2 #(
		.INIT('h2)
	) name622 (
		\DataOut_pad_o[5]_pad ,
		\u0_u0_drive_k_reg/P0001 ,
		_w2372_
	);
	LUT3 #(
		.INIT('he0)
	) name623 (
		_w1755_,
		_w1757_,
		_w2372_,
		_w2373_
	);
	LUT4 #(
		.INIT('h01ef)
	) name624 (
		_w1755_,
		_w1757_,
		_w1811_,
		_w2372_,
		_w2374_
	);
	LUT3 #(
		.INIT('h45)
	) name625 (
		\u1_u1_crc16_reg[10]/P0001 ,
		_w1805_,
		_w1820_,
		_w2375_
	);
	LUT3 #(
		.INIT('h20)
	) name626 (
		\u0_tx_ready_reg/NET0131 ,
		\u1_u1_crc16_reg[2]/P0001 ,
		\u1_u1_state_reg[2]/NET0131 ,
		_w2376_
	);
	LUT3 #(
		.INIT('h01)
	) name627 (
		\u1_u1_crc16_reg[2]/P0001 ,
		\u1_u1_state_reg[0]/NET0131 ,
		\u1_u1_state_reg[1]/NET0131 ,
		_w2377_
	);
	LUT3 #(
		.INIT('h13)
	) name628 (
		_w1809_,
		_w2376_,
		_w2377_,
		_w2378_
	);
	LUT4 #(
		.INIT('h0f0b)
	) name629 (
		_w1805_,
		_w1820_,
		_w2373_,
		_w2378_,
		_w2379_
	);
	LUT4 #(
		.INIT('h3233)
	) name630 (
		_w1828_,
		_w2374_,
		_w2375_,
		_w2379_,
		_w2380_
	);
	LUT4 #(
		.INIT('h0040)
	) name631 (
		_w1805_,
		_w1810_,
		_w1816_,
		_w2373_,
		_w2381_
	);
	LUT3 #(
		.INIT('h4c)
	) name632 (
		_w2019_,
		_w2380_,
		_w2381_,
		_w2382_
	);
	LUT4 #(
		.INIT('h0008)
	) name633 (
		\u1_u3_buffer_full_reg/P0001 ,
		\u1_u3_in_token_reg/NET0131 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		_w2383_
	);
	LUT3 #(
		.INIT('hc8)
	) name634 (
		\u1_u3_buf0_na_reg/NET0131 ,
		\u1_u3_buffer_full_reg/P0001 ,
		\u4_csr_reg[30]/NET0131 ,
		_w2384_
	);
	LUT3 #(
		.INIT('h13)
	) name635 (
		_w2352_,
		_w2383_,
		_w2384_,
		_w2385_
	);
	LUT4 #(
		.INIT('haaa2)
	) name636 (
		\u1_u3_buf1_st_max_reg/P0001 ,
		\u1_u3_in_token_reg/NET0131 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		_w2386_
	);
	LUT4 #(
		.INIT('h0455)
	) name637 (
		\u1_u3_buf1_na_reg/NET0131 ,
		_w2352_,
		_w2353_,
		_w2386_,
		_w2387_
	);
	LUT2 #(
		.INIT('h7)
	) name638 (
		_w2385_,
		_w2387_,
		_w2388_
	);
	LUT3 #(
		.INIT('h40)
	) name639 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_data_i[11]_pad ,
		_w2389_
	);
	LUT3 #(
		.INIT('h2a)
	) name640 (
		rst_i_pad,
		_w2231_,
		_w2389_,
		_w2390_
	);
	LUT4 #(
		.INIT('hd8f0)
	) name641 (
		\u1_u3_buf0_set_reg/P0001 ,
		\u1_u3_idin_reg[11]/P0001 ,
		\u4_u3_buf0_reg[11]/P0001 ,
		\u4_u3_ep_match_r_reg/P0001 ,
		_w2391_
	);
	LUT3 #(
		.INIT('hb8)
	) name642 (
		\u4_u3_buf0_orig_reg[11]/P0001 ,
		_w2235_,
		_w2391_,
		_w2392_
	);
	LUT3 #(
		.INIT('h70)
	) name643 (
		_w2231_,
		_w2232_,
		_w2392_,
		_w2393_
	);
	LUT2 #(
		.INIT('hd)
	) name644 (
		_w2390_,
		_w2393_,
		_w2394_
	);
	LUT3 #(
		.INIT('h40)
	) name645 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_data_i[15]_pad ,
		_w2395_
	);
	LUT3 #(
		.INIT('h2a)
	) name646 (
		rst_i_pad,
		_w2231_,
		_w2395_,
		_w2396_
	);
	LUT4 #(
		.INIT('hd8f0)
	) name647 (
		\u1_u3_buf0_set_reg/P0001 ,
		\u1_u3_idin_reg[15]/P0001 ,
		\u4_u3_buf0_reg[15]/P0001 ,
		\u4_u3_ep_match_r_reg/P0001 ,
		_w2397_
	);
	LUT3 #(
		.INIT('hb8)
	) name648 (
		\u4_u3_buf0_orig_reg[15]/P0001 ,
		_w2235_,
		_w2397_,
		_w2398_
	);
	LUT3 #(
		.INIT('h70)
	) name649 (
		_w2231_,
		_w2232_,
		_w2398_,
		_w2399_
	);
	LUT2 #(
		.INIT('hd)
	) name650 (
		_w2396_,
		_w2399_,
		_w2400_
	);
	LUT4 #(
		.INIT('h10f0)
	) name651 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u3_buf1_reg[10]/P0001 ,
		\u4_u3_ep_match_r_reg/P0001 ,
		_w2401_
	);
	LUT4 #(
		.INIT('hc800)
	) name652 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_idin_reg[10]/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u3_ep_match_r_reg/P0001 ,
		_w2402_
	);
	LUT2 #(
		.INIT('h1)
	) name653 (
		_w2401_,
		_w2402_,
		_w2403_
	);
	LUT3 #(
		.INIT('h07)
	) name654 (
		_w2231_,
		_w2320_,
		_w2403_,
		_w2404_
	);
	LUT3 #(
		.INIT('h80)
	) name655 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_data_i[10]_pad ,
		_w2405_
	);
	LUT3 #(
		.INIT('h2a)
	) name656 (
		rst_i_pad,
		_w2231_,
		_w2405_,
		_w2406_
	);
	LUT2 #(
		.INIT('hb)
	) name657 (
		_w2404_,
		_w2406_,
		_w2407_
	);
	LUT3 #(
		.INIT('h40)
	) name658 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_data_i[6]_pad ,
		_w2408_
	);
	LUT3 #(
		.INIT('h2a)
	) name659 (
		rst_i_pad,
		_w2231_,
		_w2408_,
		_w2409_
	);
	LUT4 #(
		.INIT('hd8f0)
	) name660 (
		\u1_u3_buf0_set_reg/P0001 ,
		\u1_u3_idin_reg[6]/P0001 ,
		\u4_u3_buf0_reg[6]/P0001 ,
		\u4_u3_ep_match_r_reg/P0001 ,
		_w2410_
	);
	LUT3 #(
		.INIT('hb8)
	) name661 (
		\u4_u3_buf0_orig_reg[6]/P0001 ,
		_w2235_,
		_w2410_,
		_w2411_
	);
	LUT3 #(
		.INIT('h70)
	) name662 (
		_w2231_,
		_w2232_,
		_w2411_,
		_w2412_
	);
	LUT2 #(
		.INIT('hd)
	) name663 (
		_w2409_,
		_w2412_,
		_w2413_
	);
	LUT3 #(
		.INIT('h2a)
	) name664 (
		rst_i_pad,
		_w2243_,
		_w2389_,
		_w2414_
	);
	LUT4 #(
		.INIT('hd8f0)
	) name665 (
		\u1_u3_buf0_set_reg/P0001 ,
		\u1_u3_idin_reg[11]/P0001 ,
		\u4_u0_buf0_reg[11]/P0001 ,
		\u4_u0_ep_match_r_reg/P0001 ,
		_w2415_
	);
	LUT3 #(
		.INIT('hb8)
	) name666 (
		\u4_u0_buf0_orig_reg[11]/P0001 ,
		_w2245_,
		_w2415_,
		_w2416_
	);
	LUT3 #(
		.INIT('h70)
	) name667 (
		_w2232_,
		_w2243_,
		_w2416_,
		_w2417_
	);
	LUT2 #(
		.INIT('hd)
	) name668 (
		_w2414_,
		_w2417_,
		_w2418_
	);
	LUT3 #(
		.INIT('h2a)
	) name669 (
		rst_i_pad,
		_w2243_,
		_w2395_,
		_w2419_
	);
	LUT4 #(
		.INIT('hd8f0)
	) name670 (
		\u1_u3_buf0_set_reg/P0001 ,
		\u1_u3_idin_reg[15]/P0001 ,
		\u4_u0_buf0_reg[15]/P0001 ,
		\u4_u0_ep_match_r_reg/P0001 ,
		_w2420_
	);
	LUT3 #(
		.INIT('hb8)
	) name671 (
		\u4_u0_buf0_orig_reg[15]/P0001 ,
		_w2245_,
		_w2420_,
		_w2421_
	);
	LUT3 #(
		.INIT('h70)
	) name672 (
		_w2232_,
		_w2243_,
		_w2421_,
		_w2422_
	);
	LUT2 #(
		.INIT('hd)
	) name673 (
		_w2419_,
		_w2422_,
		_w2423_
	);
	LUT3 #(
		.INIT('h2a)
	) name674 (
		rst_i_pad,
		_w2243_,
		_w2408_,
		_w2424_
	);
	LUT4 #(
		.INIT('hd8f0)
	) name675 (
		\u1_u3_buf0_set_reg/P0001 ,
		\u1_u3_idin_reg[6]/P0001 ,
		\u4_u0_buf0_reg[6]/P0001 ,
		\u4_u0_ep_match_r_reg/P0001 ,
		_w2425_
	);
	LUT3 #(
		.INIT('hb8)
	) name676 (
		\u4_u0_buf0_orig_reg[6]/P0001 ,
		_w2245_,
		_w2425_,
		_w2426_
	);
	LUT3 #(
		.INIT('h70)
	) name677 (
		_w2232_,
		_w2243_,
		_w2426_,
		_w2427_
	);
	LUT2 #(
		.INIT('hd)
	) name678 (
		_w2424_,
		_w2427_,
		_w2428_
	);
	LUT4 #(
		.INIT('h10f0)
	) name679 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u0_buf1_reg[10]/P0001 ,
		\u4_u0_ep_match_r_reg/P0001 ,
		_w2429_
	);
	LUT4 #(
		.INIT('hc800)
	) name680 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_idin_reg[10]/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u0_ep_match_r_reg/P0001 ,
		_w2430_
	);
	LUT2 #(
		.INIT('h1)
	) name681 (
		_w2429_,
		_w2430_,
		_w2431_
	);
	LUT3 #(
		.INIT('h07)
	) name682 (
		_w2243_,
		_w2320_,
		_w2431_,
		_w2432_
	);
	LUT3 #(
		.INIT('h2a)
	) name683 (
		rst_i_pad,
		_w2243_,
		_w2405_,
		_w2433_
	);
	LUT2 #(
		.INIT('hb)
	) name684 (
		_w2432_,
		_w2433_,
		_w2434_
	);
	LUT3 #(
		.INIT('h2a)
	) name685 (
		rst_i_pad,
		_w2260_,
		_w2389_,
		_w2435_
	);
	LUT4 #(
		.INIT('hd8f0)
	) name686 (
		\u1_u3_buf0_set_reg/P0001 ,
		\u1_u3_idin_reg[11]/P0001 ,
		\u4_u1_buf0_reg[11]/P0001 ,
		\u4_u1_ep_match_r_reg/P0001 ,
		_w2436_
	);
	LUT3 #(
		.INIT('hb8)
	) name687 (
		\u4_u1_buf0_orig_reg[11]/P0001 ,
		_w2262_,
		_w2436_,
		_w2437_
	);
	LUT3 #(
		.INIT('h70)
	) name688 (
		_w2232_,
		_w2260_,
		_w2437_,
		_w2438_
	);
	LUT2 #(
		.INIT('hd)
	) name689 (
		_w2435_,
		_w2438_,
		_w2439_
	);
	LUT3 #(
		.INIT('h2a)
	) name690 (
		rst_i_pad,
		_w2260_,
		_w2395_,
		_w2440_
	);
	LUT4 #(
		.INIT('hd8f0)
	) name691 (
		\u1_u3_buf0_set_reg/P0001 ,
		\u1_u3_idin_reg[15]/P0001 ,
		\u4_u1_buf0_reg[15]/P0001 ,
		\u4_u1_ep_match_r_reg/P0001 ,
		_w2441_
	);
	LUT3 #(
		.INIT('hb8)
	) name692 (
		\u4_u1_buf0_orig_reg[15]/P0001 ,
		_w2262_,
		_w2441_,
		_w2442_
	);
	LUT3 #(
		.INIT('h70)
	) name693 (
		_w2232_,
		_w2260_,
		_w2442_,
		_w2443_
	);
	LUT2 #(
		.INIT('hd)
	) name694 (
		_w2440_,
		_w2443_,
		_w2444_
	);
	LUT4 #(
		.INIT('h10f0)
	) name695 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u1_buf1_reg[10]/P0001 ,
		\u4_u1_ep_match_r_reg/P0001 ,
		_w2445_
	);
	LUT4 #(
		.INIT('hc800)
	) name696 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_idin_reg[10]/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u1_ep_match_r_reg/P0001 ,
		_w2446_
	);
	LUT2 #(
		.INIT('h1)
	) name697 (
		_w2445_,
		_w2446_,
		_w2447_
	);
	LUT3 #(
		.INIT('h07)
	) name698 (
		_w2260_,
		_w2320_,
		_w2447_,
		_w2448_
	);
	LUT3 #(
		.INIT('h2a)
	) name699 (
		rst_i_pad,
		_w2260_,
		_w2405_,
		_w2449_
	);
	LUT2 #(
		.INIT('hb)
	) name700 (
		_w2448_,
		_w2449_,
		_w2450_
	);
	LUT3 #(
		.INIT('h2a)
	) name701 (
		rst_i_pad,
		_w2260_,
		_w2408_,
		_w2451_
	);
	LUT4 #(
		.INIT('hd8f0)
	) name702 (
		\u1_u3_buf0_set_reg/P0001 ,
		\u1_u3_idin_reg[6]/P0001 ,
		\u4_u1_buf0_reg[6]/P0001 ,
		\u4_u1_ep_match_r_reg/P0001 ,
		_w2452_
	);
	LUT3 #(
		.INIT('hb8)
	) name703 (
		\u4_u1_buf0_orig_reg[6]/P0001 ,
		_w2262_,
		_w2452_,
		_w2453_
	);
	LUT3 #(
		.INIT('h70)
	) name704 (
		_w2232_,
		_w2260_,
		_w2453_,
		_w2454_
	);
	LUT2 #(
		.INIT('hd)
	) name705 (
		_w2451_,
		_w2454_,
		_w2455_
	);
	LUT3 #(
		.INIT('h2a)
	) name706 (
		rst_i_pad,
		_w2267_,
		_w2389_,
		_w2456_
	);
	LUT4 #(
		.INIT('hd8f0)
	) name707 (
		\u1_u3_buf0_set_reg/P0001 ,
		\u1_u3_idin_reg[11]/P0001 ,
		\u4_u2_buf0_reg[11]/P0001 ,
		\u4_u2_ep_match_r_reg/P0001 ,
		_w2457_
	);
	LUT3 #(
		.INIT('hb8)
	) name708 (
		\u4_u2_buf0_orig_reg[11]/P0001 ,
		_w2269_,
		_w2457_,
		_w2458_
	);
	LUT3 #(
		.INIT('h70)
	) name709 (
		_w2232_,
		_w2267_,
		_w2458_,
		_w2459_
	);
	LUT2 #(
		.INIT('hd)
	) name710 (
		_w2456_,
		_w2459_,
		_w2460_
	);
	LUT3 #(
		.INIT('h2a)
	) name711 (
		rst_i_pad,
		_w2267_,
		_w2395_,
		_w2461_
	);
	LUT4 #(
		.INIT('hd8f0)
	) name712 (
		\u1_u3_buf0_set_reg/P0001 ,
		\u1_u3_idin_reg[15]/P0001 ,
		\u4_u2_buf0_reg[15]/P0001 ,
		\u4_u2_ep_match_r_reg/P0001 ,
		_w2462_
	);
	LUT3 #(
		.INIT('hb8)
	) name713 (
		\u4_u2_buf0_orig_reg[15]/P0001 ,
		_w2269_,
		_w2462_,
		_w2463_
	);
	LUT3 #(
		.INIT('h70)
	) name714 (
		_w2232_,
		_w2267_,
		_w2463_,
		_w2464_
	);
	LUT2 #(
		.INIT('hd)
	) name715 (
		_w2461_,
		_w2464_,
		_w2465_
	);
	LUT4 #(
		.INIT('h10f0)
	) name716 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u2_buf1_reg[10]/P0001 ,
		\u4_u2_ep_match_r_reg/P0001 ,
		_w2466_
	);
	LUT4 #(
		.INIT('hc800)
	) name717 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_idin_reg[10]/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u2_ep_match_r_reg/P0001 ,
		_w2467_
	);
	LUT2 #(
		.INIT('h1)
	) name718 (
		_w2466_,
		_w2467_,
		_w2468_
	);
	LUT3 #(
		.INIT('h07)
	) name719 (
		_w2267_,
		_w2320_,
		_w2468_,
		_w2469_
	);
	LUT3 #(
		.INIT('h2a)
	) name720 (
		rst_i_pad,
		_w2267_,
		_w2405_,
		_w2470_
	);
	LUT2 #(
		.INIT('hb)
	) name721 (
		_w2469_,
		_w2470_,
		_w2471_
	);
	LUT3 #(
		.INIT('h2a)
	) name722 (
		rst_i_pad,
		_w2267_,
		_w2408_,
		_w2472_
	);
	LUT4 #(
		.INIT('hd8f0)
	) name723 (
		\u1_u3_buf0_set_reg/P0001 ,
		\u1_u3_idin_reg[6]/P0001 ,
		\u4_u2_buf0_reg[6]/P0001 ,
		\u4_u2_ep_match_r_reg/P0001 ,
		_w2473_
	);
	LUT3 #(
		.INIT('hb8)
	) name724 (
		\u4_u2_buf0_orig_reg[6]/P0001 ,
		_w2269_,
		_w2473_,
		_w2474_
	);
	LUT3 #(
		.INIT('h70)
	) name725 (
		_w2232_,
		_w2267_,
		_w2474_,
		_w2475_
	);
	LUT2 #(
		.INIT('hd)
	) name726 (
		_w2472_,
		_w2475_,
		_w2476_
	);
	LUT4 #(
		.INIT('h10f0)
	) name727 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u3_buf1_reg[13]/P0001 ,
		\u4_u3_ep_match_r_reg/P0001 ,
		_w2477_
	);
	LUT4 #(
		.INIT('hc800)
	) name728 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_idin_reg[13]/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u3_ep_match_r_reg/P0001 ,
		_w2478_
	);
	LUT2 #(
		.INIT('h1)
	) name729 (
		_w2477_,
		_w2478_,
		_w2479_
	);
	LUT3 #(
		.INIT('h07)
	) name730 (
		_w2231_,
		_w2320_,
		_w2479_,
		_w2480_
	);
	LUT3 #(
		.INIT('h80)
	) name731 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_data_i[13]_pad ,
		_w2481_
	);
	LUT3 #(
		.INIT('h2a)
	) name732 (
		rst_i_pad,
		_w2231_,
		_w2481_,
		_w2482_
	);
	LUT2 #(
		.INIT('hb)
	) name733 (
		_w2480_,
		_w2482_,
		_w2483_
	);
	LUT4 #(
		.INIT('h10f0)
	) name734 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u0_buf1_reg[13]/P0001 ,
		\u4_u0_ep_match_r_reg/P0001 ,
		_w2484_
	);
	LUT4 #(
		.INIT('hc800)
	) name735 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_idin_reg[13]/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u0_ep_match_r_reg/P0001 ,
		_w2485_
	);
	LUT2 #(
		.INIT('h1)
	) name736 (
		_w2484_,
		_w2485_,
		_w2486_
	);
	LUT3 #(
		.INIT('h07)
	) name737 (
		_w2243_,
		_w2320_,
		_w2486_,
		_w2487_
	);
	LUT3 #(
		.INIT('h2a)
	) name738 (
		rst_i_pad,
		_w2243_,
		_w2481_,
		_w2488_
	);
	LUT2 #(
		.INIT('hb)
	) name739 (
		_w2487_,
		_w2488_,
		_w2489_
	);
	LUT4 #(
		.INIT('h10f0)
	) name740 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u1_buf1_reg[13]/P0001 ,
		\u4_u1_ep_match_r_reg/P0001 ,
		_w2490_
	);
	LUT4 #(
		.INIT('hc800)
	) name741 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_idin_reg[13]/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u1_ep_match_r_reg/P0001 ,
		_w2491_
	);
	LUT2 #(
		.INIT('h1)
	) name742 (
		_w2490_,
		_w2491_,
		_w2492_
	);
	LUT3 #(
		.INIT('h07)
	) name743 (
		_w2260_,
		_w2320_,
		_w2492_,
		_w2493_
	);
	LUT3 #(
		.INIT('h2a)
	) name744 (
		rst_i_pad,
		_w2260_,
		_w2481_,
		_w2494_
	);
	LUT2 #(
		.INIT('hb)
	) name745 (
		_w2493_,
		_w2494_,
		_w2495_
	);
	LUT4 #(
		.INIT('h10f0)
	) name746 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u2_buf1_reg[13]/P0001 ,
		\u4_u2_ep_match_r_reg/P0001 ,
		_w2496_
	);
	LUT4 #(
		.INIT('hc800)
	) name747 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_idin_reg[13]/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u2_ep_match_r_reg/P0001 ,
		_w2497_
	);
	LUT2 #(
		.INIT('h1)
	) name748 (
		_w2496_,
		_w2497_,
		_w2498_
	);
	LUT3 #(
		.INIT('h07)
	) name749 (
		_w2267_,
		_w2320_,
		_w2498_,
		_w2499_
	);
	LUT3 #(
		.INIT('h2a)
	) name750 (
		rst_i_pad,
		_w2267_,
		_w2481_,
		_w2500_
	);
	LUT2 #(
		.INIT('hb)
	) name751 (
		_w2499_,
		_w2500_,
		_w2501_
	);
	LUT4 #(
		.INIT('h00a8)
	) name752 (
		\u1_u3_buffer_empty_reg/P0001 ,
		\u1_u3_in_token_reg/NET0131 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		_w2502_
	);
	LUT3 #(
		.INIT('h0e)
	) name753 (
		\u1_u3_in_token_reg/NET0131 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		_w2503_
	);
	LUT4 #(
		.INIT('haa02)
	) name754 (
		\u1_u3_buffer_full_reg/P0001 ,
		\u1_u3_in_token_reg/NET0131 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		_w2504_
	);
	LUT2 #(
		.INIT('he)
	) name755 (
		_w2502_,
		_w2504_,
		_w2505_
	);
	LUT3 #(
		.INIT('h40)
	) name756 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_data_i[4]_pad ,
		_w2506_
	);
	LUT3 #(
		.INIT('h2a)
	) name757 (
		rst_i_pad,
		_w2231_,
		_w2506_,
		_w2507_
	);
	LUT4 #(
		.INIT('hd8f0)
	) name758 (
		\u1_u3_buf0_set_reg/P0001 ,
		\u1_u3_idin_reg[4]/P0001 ,
		\u4_u3_buf0_reg[4]/P0001 ,
		\u4_u3_ep_match_r_reg/P0001 ,
		_w2508_
	);
	LUT3 #(
		.INIT('hb8)
	) name759 (
		\u4_u3_buf0_orig_reg[4]/P0001 ,
		_w2235_,
		_w2508_,
		_w2509_
	);
	LUT3 #(
		.INIT('h70)
	) name760 (
		_w2231_,
		_w2232_,
		_w2509_,
		_w2510_
	);
	LUT2 #(
		.INIT('hd)
	) name761 (
		_w2507_,
		_w2510_,
		_w2511_
	);
	LUT3 #(
		.INIT('h40)
	) name762 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_data_i[5]_pad ,
		_w2512_
	);
	LUT3 #(
		.INIT('h2a)
	) name763 (
		rst_i_pad,
		_w2231_,
		_w2512_,
		_w2513_
	);
	LUT4 #(
		.INIT('hd8f0)
	) name764 (
		\u1_u3_buf0_set_reg/P0001 ,
		\u1_u3_idin_reg[5]/P0001 ,
		\u4_u3_buf0_reg[5]/P0001 ,
		\u4_u3_ep_match_r_reg/P0001 ,
		_w2514_
	);
	LUT3 #(
		.INIT('hb8)
	) name765 (
		\u4_u3_buf0_orig_reg[5]/P0001 ,
		_w2235_,
		_w2514_,
		_w2515_
	);
	LUT3 #(
		.INIT('h70)
	) name766 (
		_w2231_,
		_w2232_,
		_w2515_,
		_w2516_
	);
	LUT2 #(
		.INIT('hd)
	) name767 (
		_w2513_,
		_w2516_,
		_w2517_
	);
	LUT3 #(
		.INIT('h40)
	) name768 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_data_i[7]_pad ,
		_w2518_
	);
	LUT3 #(
		.INIT('h2a)
	) name769 (
		rst_i_pad,
		_w2231_,
		_w2518_,
		_w2519_
	);
	LUT4 #(
		.INIT('hd8f0)
	) name770 (
		\u1_u3_buf0_set_reg/P0001 ,
		\u1_u3_idin_reg[7]/P0001 ,
		\u4_u3_buf0_reg[7]/P0001 ,
		\u4_u3_ep_match_r_reg/P0001 ,
		_w2520_
	);
	LUT3 #(
		.INIT('hb8)
	) name771 (
		\u4_u3_buf0_orig_reg[7]/P0001 ,
		_w2235_,
		_w2520_,
		_w2521_
	);
	LUT3 #(
		.INIT('h70)
	) name772 (
		_w2231_,
		_w2232_,
		_w2521_,
		_w2522_
	);
	LUT2 #(
		.INIT('hd)
	) name773 (
		_w2519_,
		_w2522_,
		_w2523_
	);
	LUT4 #(
		.INIT('h10f0)
	) name774 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u3_buf1_reg[11]/P0001 ,
		\u4_u3_ep_match_r_reg/P0001 ,
		_w2524_
	);
	LUT4 #(
		.INIT('hc800)
	) name775 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_idin_reg[11]/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u3_ep_match_r_reg/P0001 ,
		_w2525_
	);
	LUT2 #(
		.INIT('h1)
	) name776 (
		_w2524_,
		_w2525_,
		_w2526_
	);
	LUT3 #(
		.INIT('h07)
	) name777 (
		_w2231_,
		_w2320_,
		_w2526_,
		_w2527_
	);
	LUT3 #(
		.INIT('h80)
	) name778 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_data_i[11]_pad ,
		_w2528_
	);
	LUT3 #(
		.INIT('h2a)
	) name779 (
		rst_i_pad,
		_w2231_,
		_w2528_,
		_w2529_
	);
	LUT2 #(
		.INIT('hb)
	) name780 (
		_w2527_,
		_w2529_,
		_w2530_
	);
	LUT4 #(
		.INIT('h10f0)
	) name781 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u3_buf1_reg[15]/P0001 ,
		\u4_u3_ep_match_r_reg/P0001 ,
		_w2531_
	);
	LUT4 #(
		.INIT('hc800)
	) name782 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_idin_reg[15]/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u3_ep_match_r_reg/P0001 ,
		_w2532_
	);
	LUT2 #(
		.INIT('h1)
	) name783 (
		_w2531_,
		_w2532_,
		_w2533_
	);
	LUT3 #(
		.INIT('h07)
	) name784 (
		_w2231_,
		_w2320_,
		_w2533_,
		_w2534_
	);
	LUT3 #(
		.INIT('h80)
	) name785 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_data_i[15]_pad ,
		_w2535_
	);
	LUT3 #(
		.INIT('h2a)
	) name786 (
		rst_i_pad,
		_w2231_,
		_w2535_,
		_w2536_
	);
	LUT2 #(
		.INIT('hb)
	) name787 (
		_w2534_,
		_w2536_,
		_w2537_
	);
	LUT4 #(
		.INIT('h10f0)
	) name788 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u3_buf1_reg[6]/P0001 ,
		\u4_u3_ep_match_r_reg/P0001 ,
		_w2538_
	);
	LUT4 #(
		.INIT('hc800)
	) name789 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_idin_reg[6]/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u3_ep_match_r_reg/P0001 ,
		_w2539_
	);
	LUT2 #(
		.INIT('h1)
	) name790 (
		_w2538_,
		_w2539_,
		_w2540_
	);
	LUT3 #(
		.INIT('h07)
	) name791 (
		_w2231_,
		_w2320_,
		_w2540_,
		_w2541_
	);
	LUT3 #(
		.INIT('h80)
	) name792 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_data_i[6]_pad ,
		_w2542_
	);
	LUT3 #(
		.INIT('h2a)
	) name793 (
		rst_i_pad,
		_w2231_,
		_w2542_,
		_w2543_
	);
	LUT2 #(
		.INIT('hb)
	) name794 (
		_w2541_,
		_w2543_,
		_w2544_
	);
	LUT3 #(
		.INIT('h2a)
	) name795 (
		rst_i_pad,
		_w2243_,
		_w2506_,
		_w2545_
	);
	LUT4 #(
		.INIT('hd8f0)
	) name796 (
		\u1_u3_buf0_set_reg/P0001 ,
		\u1_u3_idin_reg[4]/P0001 ,
		\u4_u0_buf0_reg[4]/P0001 ,
		\u4_u0_ep_match_r_reg/P0001 ,
		_w2546_
	);
	LUT3 #(
		.INIT('hb8)
	) name797 (
		\u4_u0_buf0_orig_reg[4]/P0001 ,
		_w2245_,
		_w2546_,
		_w2547_
	);
	LUT3 #(
		.INIT('h70)
	) name798 (
		_w2232_,
		_w2243_,
		_w2547_,
		_w2548_
	);
	LUT2 #(
		.INIT('hd)
	) name799 (
		_w2545_,
		_w2548_,
		_w2549_
	);
	LUT3 #(
		.INIT('h2a)
	) name800 (
		rst_i_pad,
		_w2243_,
		_w2512_,
		_w2550_
	);
	LUT4 #(
		.INIT('hd8f0)
	) name801 (
		\u1_u3_buf0_set_reg/P0001 ,
		\u1_u3_idin_reg[5]/P0001 ,
		\u4_u0_buf0_reg[5]/P0001 ,
		\u4_u0_ep_match_r_reg/P0001 ,
		_w2551_
	);
	LUT3 #(
		.INIT('hb8)
	) name802 (
		\u4_u0_buf0_orig_reg[5]/P0001 ,
		_w2245_,
		_w2551_,
		_w2552_
	);
	LUT3 #(
		.INIT('h70)
	) name803 (
		_w2232_,
		_w2243_,
		_w2552_,
		_w2553_
	);
	LUT2 #(
		.INIT('hd)
	) name804 (
		_w2550_,
		_w2553_,
		_w2554_
	);
	LUT3 #(
		.INIT('h2a)
	) name805 (
		rst_i_pad,
		_w2243_,
		_w2518_,
		_w2555_
	);
	LUT4 #(
		.INIT('hd8f0)
	) name806 (
		\u1_u3_buf0_set_reg/P0001 ,
		\u1_u3_idin_reg[7]/P0001 ,
		\u4_u0_buf0_reg[7]/P0001 ,
		\u4_u0_ep_match_r_reg/P0001 ,
		_w2556_
	);
	LUT3 #(
		.INIT('hb8)
	) name807 (
		\u4_u0_buf0_orig_reg[7]/P0001 ,
		_w2245_,
		_w2556_,
		_w2557_
	);
	LUT3 #(
		.INIT('h70)
	) name808 (
		_w2232_,
		_w2243_,
		_w2557_,
		_w2558_
	);
	LUT2 #(
		.INIT('hd)
	) name809 (
		_w2555_,
		_w2558_,
		_w2559_
	);
	LUT4 #(
		.INIT('h10f0)
	) name810 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u0_buf1_reg[11]/P0001 ,
		\u4_u0_ep_match_r_reg/P0001 ,
		_w2560_
	);
	LUT4 #(
		.INIT('hc800)
	) name811 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_idin_reg[11]/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u0_ep_match_r_reg/P0001 ,
		_w2561_
	);
	LUT2 #(
		.INIT('h1)
	) name812 (
		_w2560_,
		_w2561_,
		_w2562_
	);
	LUT3 #(
		.INIT('h07)
	) name813 (
		_w2243_,
		_w2320_,
		_w2562_,
		_w2563_
	);
	LUT3 #(
		.INIT('h2a)
	) name814 (
		rst_i_pad,
		_w2243_,
		_w2528_,
		_w2564_
	);
	LUT2 #(
		.INIT('hb)
	) name815 (
		_w2563_,
		_w2564_,
		_w2565_
	);
	LUT4 #(
		.INIT('h10f0)
	) name816 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u0_buf1_reg[15]/P0001 ,
		\u4_u0_ep_match_r_reg/P0001 ,
		_w2566_
	);
	LUT4 #(
		.INIT('hc800)
	) name817 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_idin_reg[15]/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u0_ep_match_r_reg/P0001 ,
		_w2567_
	);
	LUT2 #(
		.INIT('h1)
	) name818 (
		_w2566_,
		_w2567_,
		_w2568_
	);
	LUT3 #(
		.INIT('h07)
	) name819 (
		_w2243_,
		_w2320_,
		_w2568_,
		_w2569_
	);
	LUT3 #(
		.INIT('h2a)
	) name820 (
		rst_i_pad,
		_w2243_,
		_w2535_,
		_w2570_
	);
	LUT2 #(
		.INIT('hb)
	) name821 (
		_w2569_,
		_w2570_,
		_w2571_
	);
	LUT4 #(
		.INIT('h10f0)
	) name822 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u0_buf1_reg[6]/P0001 ,
		\u4_u0_ep_match_r_reg/P0001 ,
		_w2572_
	);
	LUT4 #(
		.INIT('hc800)
	) name823 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_idin_reg[6]/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u0_ep_match_r_reg/P0001 ,
		_w2573_
	);
	LUT2 #(
		.INIT('h1)
	) name824 (
		_w2572_,
		_w2573_,
		_w2574_
	);
	LUT3 #(
		.INIT('h07)
	) name825 (
		_w2243_,
		_w2320_,
		_w2574_,
		_w2575_
	);
	LUT3 #(
		.INIT('h2a)
	) name826 (
		rst_i_pad,
		_w2243_,
		_w2542_,
		_w2576_
	);
	LUT2 #(
		.INIT('hb)
	) name827 (
		_w2575_,
		_w2576_,
		_w2577_
	);
	LUT3 #(
		.INIT('h2a)
	) name828 (
		rst_i_pad,
		_w2260_,
		_w2506_,
		_w2578_
	);
	LUT4 #(
		.INIT('hd8f0)
	) name829 (
		\u1_u3_buf0_set_reg/P0001 ,
		\u1_u3_idin_reg[4]/P0001 ,
		\u4_u1_buf0_reg[4]/P0001 ,
		\u4_u1_ep_match_r_reg/P0001 ,
		_w2579_
	);
	LUT3 #(
		.INIT('hb8)
	) name830 (
		\u4_u1_buf0_orig_reg[4]/P0001 ,
		_w2262_,
		_w2579_,
		_w2580_
	);
	LUT3 #(
		.INIT('h70)
	) name831 (
		_w2232_,
		_w2260_,
		_w2580_,
		_w2581_
	);
	LUT2 #(
		.INIT('hd)
	) name832 (
		_w2578_,
		_w2581_,
		_w2582_
	);
	LUT3 #(
		.INIT('h2a)
	) name833 (
		rst_i_pad,
		_w2260_,
		_w2512_,
		_w2583_
	);
	LUT4 #(
		.INIT('hd8f0)
	) name834 (
		\u1_u3_buf0_set_reg/P0001 ,
		\u1_u3_idin_reg[5]/P0001 ,
		\u4_u1_buf0_reg[5]/P0001 ,
		\u4_u1_ep_match_r_reg/P0001 ,
		_w2584_
	);
	LUT3 #(
		.INIT('hb8)
	) name835 (
		\u4_u1_buf0_orig_reg[5]/P0001 ,
		_w2262_,
		_w2584_,
		_w2585_
	);
	LUT3 #(
		.INIT('h70)
	) name836 (
		_w2232_,
		_w2260_,
		_w2585_,
		_w2586_
	);
	LUT2 #(
		.INIT('hd)
	) name837 (
		_w2583_,
		_w2586_,
		_w2587_
	);
	LUT3 #(
		.INIT('h2a)
	) name838 (
		rst_i_pad,
		_w2260_,
		_w2518_,
		_w2588_
	);
	LUT4 #(
		.INIT('hd8f0)
	) name839 (
		\u1_u3_buf0_set_reg/P0001 ,
		\u1_u3_idin_reg[7]/P0001 ,
		\u4_u1_buf0_reg[7]/P0001 ,
		\u4_u1_ep_match_r_reg/P0001 ,
		_w2589_
	);
	LUT3 #(
		.INIT('hb8)
	) name840 (
		\u4_u1_buf0_orig_reg[7]/P0001 ,
		_w2262_,
		_w2589_,
		_w2590_
	);
	LUT3 #(
		.INIT('h70)
	) name841 (
		_w2232_,
		_w2260_,
		_w2590_,
		_w2591_
	);
	LUT2 #(
		.INIT('hd)
	) name842 (
		_w2588_,
		_w2591_,
		_w2592_
	);
	LUT4 #(
		.INIT('h10f0)
	) name843 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u1_buf1_reg[11]/P0001 ,
		\u4_u1_ep_match_r_reg/P0001 ,
		_w2593_
	);
	LUT4 #(
		.INIT('hc800)
	) name844 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_idin_reg[11]/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u1_ep_match_r_reg/P0001 ,
		_w2594_
	);
	LUT2 #(
		.INIT('h1)
	) name845 (
		_w2593_,
		_w2594_,
		_w2595_
	);
	LUT3 #(
		.INIT('h07)
	) name846 (
		_w2260_,
		_w2320_,
		_w2595_,
		_w2596_
	);
	LUT3 #(
		.INIT('h2a)
	) name847 (
		rst_i_pad,
		_w2260_,
		_w2528_,
		_w2597_
	);
	LUT2 #(
		.INIT('hb)
	) name848 (
		_w2596_,
		_w2597_,
		_w2598_
	);
	LUT4 #(
		.INIT('h10f0)
	) name849 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u1_buf1_reg[15]/P0001 ,
		\u4_u1_ep_match_r_reg/P0001 ,
		_w2599_
	);
	LUT4 #(
		.INIT('hc800)
	) name850 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_idin_reg[15]/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u1_ep_match_r_reg/P0001 ,
		_w2600_
	);
	LUT2 #(
		.INIT('h1)
	) name851 (
		_w2599_,
		_w2600_,
		_w2601_
	);
	LUT3 #(
		.INIT('h07)
	) name852 (
		_w2260_,
		_w2320_,
		_w2601_,
		_w2602_
	);
	LUT3 #(
		.INIT('h2a)
	) name853 (
		rst_i_pad,
		_w2260_,
		_w2535_,
		_w2603_
	);
	LUT2 #(
		.INIT('hb)
	) name854 (
		_w2602_,
		_w2603_,
		_w2604_
	);
	LUT4 #(
		.INIT('h10f0)
	) name855 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u1_buf1_reg[6]/P0001 ,
		\u4_u1_ep_match_r_reg/P0001 ,
		_w2605_
	);
	LUT4 #(
		.INIT('hc800)
	) name856 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_idin_reg[6]/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u1_ep_match_r_reg/P0001 ,
		_w2606_
	);
	LUT2 #(
		.INIT('h1)
	) name857 (
		_w2605_,
		_w2606_,
		_w2607_
	);
	LUT3 #(
		.INIT('h07)
	) name858 (
		_w2260_,
		_w2320_,
		_w2607_,
		_w2608_
	);
	LUT3 #(
		.INIT('h2a)
	) name859 (
		rst_i_pad,
		_w2260_,
		_w2542_,
		_w2609_
	);
	LUT2 #(
		.INIT('hb)
	) name860 (
		_w2608_,
		_w2609_,
		_w2610_
	);
	LUT3 #(
		.INIT('h2a)
	) name861 (
		rst_i_pad,
		_w2267_,
		_w2506_,
		_w2611_
	);
	LUT4 #(
		.INIT('hd8f0)
	) name862 (
		\u1_u3_buf0_set_reg/P0001 ,
		\u1_u3_idin_reg[4]/P0001 ,
		\u4_u2_buf0_reg[4]/P0001 ,
		\u4_u2_ep_match_r_reg/P0001 ,
		_w2612_
	);
	LUT3 #(
		.INIT('hb8)
	) name863 (
		\u4_u2_buf0_orig_reg[4]/P0001 ,
		_w2269_,
		_w2612_,
		_w2613_
	);
	LUT3 #(
		.INIT('h70)
	) name864 (
		_w2232_,
		_w2267_,
		_w2613_,
		_w2614_
	);
	LUT2 #(
		.INIT('hd)
	) name865 (
		_w2611_,
		_w2614_,
		_w2615_
	);
	LUT3 #(
		.INIT('h2a)
	) name866 (
		rst_i_pad,
		_w2267_,
		_w2512_,
		_w2616_
	);
	LUT4 #(
		.INIT('hd8f0)
	) name867 (
		\u1_u3_buf0_set_reg/P0001 ,
		\u1_u3_idin_reg[5]/P0001 ,
		\u4_u2_buf0_reg[5]/P0001 ,
		\u4_u2_ep_match_r_reg/P0001 ,
		_w2617_
	);
	LUT3 #(
		.INIT('hb8)
	) name868 (
		\u4_u2_buf0_orig_reg[5]/P0001 ,
		_w2269_,
		_w2617_,
		_w2618_
	);
	LUT3 #(
		.INIT('h70)
	) name869 (
		_w2232_,
		_w2267_,
		_w2618_,
		_w2619_
	);
	LUT2 #(
		.INIT('hd)
	) name870 (
		_w2616_,
		_w2619_,
		_w2620_
	);
	LUT3 #(
		.INIT('h2a)
	) name871 (
		rst_i_pad,
		_w2267_,
		_w2518_,
		_w2621_
	);
	LUT4 #(
		.INIT('hd8f0)
	) name872 (
		\u1_u3_buf0_set_reg/P0001 ,
		\u1_u3_idin_reg[7]/P0001 ,
		\u4_u2_buf0_reg[7]/P0001 ,
		\u4_u2_ep_match_r_reg/P0001 ,
		_w2622_
	);
	LUT3 #(
		.INIT('hb8)
	) name873 (
		\u4_u2_buf0_orig_reg[7]/P0001 ,
		_w2269_,
		_w2622_,
		_w2623_
	);
	LUT3 #(
		.INIT('h70)
	) name874 (
		_w2232_,
		_w2267_,
		_w2623_,
		_w2624_
	);
	LUT2 #(
		.INIT('hd)
	) name875 (
		_w2621_,
		_w2624_,
		_w2625_
	);
	LUT4 #(
		.INIT('h10f0)
	) name876 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u2_buf1_reg[11]/P0001 ,
		\u4_u2_ep_match_r_reg/P0001 ,
		_w2626_
	);
	LUT4 #(
		.INIT('hc800)
	) name877 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_idin_reg[11]/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u2_ep_match_r_reg/P0001 ,
		_w2627_
	);
	LUT2 #(
		.INIT('h1)
	) name878 (
		_w2626_,
		_w2627_,
		_w2628_
	);
	LUT3 #(
		.INIT('h07)
	) name879 (
		_w2267_,
		_w2320_,
		_w2628_,
		_w2629_
	);
	LUT3 #(
		.INIT('h2a)
	) name880 (
		rst_i_pad,
		_w2267_,
		_w2528_,
		_w2630_
	);
	LUT2 #(
		.INIT('hb)
	) name881 (
		_w2629_,
		_w2630_,
		_w2631_
	);
	LUT4 #(
		.INIT('h10f0)
	) name882 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u2_buf1_reg[15]/P0001 ,
		\u4_u2_ep_match_r_reg/P0001 ,
		_w2632_
	);
	LUT4 #(
		.INIT('hc800)
	) name883 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_idin_reg[15]/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u2_ep_match_r_reg/P0001 ,
		_w2633_
	);
	LUT2 #(
		.INIT('h1)
	) name884 (
		_w2632_,
		_w2633_,
		_w2634_
	);
	LUT3 #(
		.INIT('h07)
	) name885 (
		_w2267_,
		_w2320_,
		_w2634_,
		_w2635_
	);
	LUT3 #(
		.INIT('h2a)
	) name886 (
		rst_i_pad,
		_w2267_,
		_w2535_,
		_w2636_
	);
	LUT2 #(
		.INIT('hb)
	) name887 (
		_w2635_,
		_w2636_,
		_w2637_
	);
	LUT4 #(
		.INIT('h10f0)
	) name888 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u2_buf1_reg[6]/P0001 ,
		\u4_u2_ep_match_r_reg/P0001 ,
		_w2638_
	);
	LUT4 #(
		.INIT('hc800)
	) name889 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_idin_reg[6]/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u2_ep_match_r_reg/P0001 ,
		_w2639_
	);
	LUT2 #(
		.INIT('h1)
	) name890 (
		_w2638_,
		_w2639_,
		_w2640_
	);
	LUT3 #(
		.INIT('h07)
	) name891 (
		_w2267_,
		_w2320_,
		_w2640_,
		_w2641_
	);
	LUT3 #(
		.INIT('h2a)
	) name892 (
		rst_i_pad,
		_w2267_,
		_w2542_,
		_w2642_
	);
	LUT2 #(
		.INIT('hb)
	) name893 (
		_w2641_,
		_w2642_,
		_w2643_
	);
	LUT4 #(
		.INIT('h10f0)
	) name894 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u3_buf1_reg[4]/P0001 ,
		\u4_u3_ep_match_r_reg/P0001 ,
		_w2644_
	);
	LUT4 #(
		.INIT('hc800)
	) name895 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_idin_reg[4]/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u3_ep_match_r_reg/P0001 ,
		_w2645_
	);
	LUT2 #(
		.INIT('h1)
	) name896 (
		_w2644_,
		_w2645_,
		_w2646_
	);
	LUT3 #(
		.INIT('h07)
	) name897 (
		_w2231_,
		_w2320_,
		_w2646_,
		_w2647_
	);
	LUT3 #(
		.INIT('h80)
	) name898 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_data_i[4]_pad ,
		_w2648_
	);
	LUT3 #(
		.INIT('h2a)
	) name899 (
		rst_i_pad,
		_w2231_,
		_w2648_,
		_w2649_
	);
	LUT2 #(
		.INIT('hb)
	) name900 (
		_w2647_,
		_w2649_,
		_w2650_
	);
	LUT4 #(
		.INIT('h10f0)
	) name901 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u3_buf1_reg[5]/P0001 ,
		\u4_u3_ep_match_r_reg/P0001 ,
		_w2651_
	);
	LUT4 #(
		.INIT('hc800)
	) name902 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_idin_reg[5]/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u3_ep_match_r_reg/P0001 ,
		_w2652_
	);
	LUT2 #(
		.INIT('h1)
	) name903 (
		_w2651_,
		_w2652_,
		_w2653_
	);
	LUT3 #(
		.INIT('h07)
	) name904 (
		_w2231_,
		_w2320_,
		_w2653_,
		_w2654_
	);
	LUT3 #(
		.INIT('h80)
	) name905 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_data_i[5]_pad ,
		_w2655_
	);
	LUT3 #(
		.INIT('h2a)
	) name906 (
		rst_i_pad,
		_w2231_,
		_w2655_,
		_w2656_
	);
	LUT2 #(
		.INIT('hb)
	) name907 (
		_w2654_,
		_w2656_,
		_w2657_
	);
	LUT4 #(
		.INIT('h10f0)
	) name908 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u3_buf1_reg[7]/P0001 ,
		\u4_u3_ep_match_r_reg/P0001 ,
		_w2658_
	);
	LUT4 #(
		.INIT('hc800)
	) name909 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_idin_reg[7]/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u3_ep_match_r_reg/P0001 ,
		_w2659_
	);
	LUT2 #(
		.INIT('h1)
	) name910 (
		_w2658_,
		_w2659_,
		_w2660_
	);
	LUT3 #(
		.INIT('h07)
	) name911 (
		_w2231_,
		_w2320_,
		_w2660_,
		_w2661_
	);
	LUT3 #(
		.INIT('h80)
	) name912 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_data_i[7]_pad ,
		_w2662_
	);
	LUT3 #(
		.INIT('h2a)
	) name913 (
		rst_i_pad,
		_w2231_,
		_w2662_,
		_w2663_
	);
	LUT2 #(
		.INIT('hb)
	) name914 (
		_w2661_,
		_w2663_,
		_w2664_
	);
	LUT4 #(
		.INIT('h10f0)
	) name915 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u0_buf1_reg[4]/P0001 ,
		\u4_u0_ep_match_r_reg/P0001 ,
		_w2665_
	);
	LUT4 #(
		.INIT('hc800)
	) name916 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_idin_reg[4]/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u0_ep_match_r_reg/P0001 ,
		_w2666_
	);
	LUT2 #(
		.INIT('h1)
	) name917 (
		_w2665_,
		_w2666_,
		_w2667_
	);
	LUT3 #(
		.INIT('h07)
	) name918 (
		_w2243_,
		_w2320_,
		_w2667_,
		_w2668_
	);
	LUT3 #(
		.INIT('h2a)
	) name919 (
		rst_i_pad,
		_w2243_,
		_w2648_,
		_w2669_
	);
	LUT2 #(
		.INIT('hb)
	) name920 (
		_w2668_,
		_w2669_,
		_w2670_
	);
	LUT4 #(
		.INIT('h10f0)
	) name921 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u0_buf1_reg[5]/P0001 ,
		\u4_u0_ep_match_r_reg/P0001 ,
		_w2671_
	);
	LUT4 #(
		.INIT('hc800)
	) name922 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_idin_reg[5]/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u0_ep_match_r_reg/P0001 ,
		_w2672_
	);
	LUT2 #(
		.INIT('h1)
	) name923 (
		_w2671_,
		_w2672_,
		_w2673_
	);
	LUT3 #(
		.INIT('h07)
	) name924 (
		_w2243_,
		_w2320_,
		_w2673_,
		_w2674_
	);
	LUT3 #(
		.INIT('h2a)
	) name925 (
		rst_i_pad,
		_w2243_,
		_w2655_,
		_w2675_
	);
	LUT2 #(
		.INIT('hb)
	) name926 (
		_w2674_,
		_w2675_,
		_w2676_
	);
	LUT4 #(
		.INIT('h10f0)
	) name927 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u0_buf1_reg[7]/P0001 ,
		\u4_u0_ep_match_r_reg/P0001 ,
		_w2677_
	);
	LUT4 #(
		.INIT('hc800)
	) name928 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_idin_reg[7]/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u0_ep_match_r_reg/P0001 ,
		_w2678_
	);
	LUT2 #(
		.INIT('h1)
	) name929 (
		_w2677_,
		_w2678_,
		_w2679_
	);
	LUT3 #(
		.INIT('h07)
	) name930 (
		_w2243_,
		_w2320_,
		_w2679_,
		_w2680_
	);
	LUT3 #(
		.INIT('h2a)
	) name931 (
		rst_i_pad,
		_w2243_,
		_w2662_,
		_w2681_
	);
	LUT2 #(
		.INIT('hb)
	) name932 (
		_w2680_,
		_w2681_,
		_w2682_
	);
	LUT4 #(
		.INIT('hf531)
	) name933 (
		\u1_u3_new_size_reg[4]/P0001 ,
		\u1_u3_new_size_reg[5]/P0001 ,
		\u4_csr_reg[4]/NET0131 ,
		\u4_csr_reg[5]/NET0131 ,
		_w2683_
	);
	LUT4 #(
		.INIT('h8caf)
	) name934 (
		\u1_u3_new_size_reg[3]/P0001 ,
		\u1_u3_new_size_reg[4]/P0001 ,
		\u4_csr_reg[3]/P0001 ,
		\u4_csr_reg[4]/NET0131 ,
		_w2684_
	);
	LUT2 #(
		.INIT('h2)
	) name935 (
		_w2683_,
		_w2684_,
		_w2685_
	);
	LUT4 #(
		.INIT('h5010)
	) name936 (
		\u1_u3_new_size_reg[0]/P0001 ,
		\u1_u3_new_size_reg[1]/P0001 ,
		\u4_csr_reg[0]/P0001 ,
		\u4_csr_reg[1]/P0001 ,
		_w2686_
	);
	LUT4 #(
		.INIT('h8caf)
	) name937 (
		\u1_u3_new_size_reg[1]/P0001 ,
		\u1_u3_new_size_reg[2]/P0001 ,
		\u4_csr_reg[1]/P0001 ,
		\u4_csr_reg[2]/NET0131 ,
		_w2687_
	);
	LUT4 #(
		.INIT('hf531)
	) name938 (
		\u1_u3_new_size_reg[2]/P0001 ,
		\u1_u3_new_size_reg[3]/P0001 ,
		\u4_csr_reg[2]/NET0131 ,
		\u4_csr_reg[3]/P0001 ,
		_w2688_
	);
	LUT4 #(
		.INIT('h8a00)
	) name939 (
		_w2683_,
		_w2686_,
		_w2687_,
		_w2688_,
		_w2689_
	);
	LUT4 #(
		.INIT('h8caf)
	) name940 (
		\u1_u3_new_size_reg[8]/P0001 ,
		\u1_u3_new_size_reg[9]/P0001 ,
		\u4_csr_reg[8]/P0001 ,
		\u4_csr_reg[9]/NET0131 ,
		_w2690_
	);
	LUT2 #(
		.INIT('h4)
	) name941 (
		\u1_u3_new_size_reg[10]/P0001 ,
		\u4_csr_reg[10]/P0001 ,
		_w2691_
	);
	LUT4 #(
		.INIT('h8caf)
	) name942 (
		\u1_u3_new_size_reg[10]/P0001 ,
		\u1_u3_new_size_reg[7]/P0001 ,
		\u4_csr_reg[10]/P0001 ,
		\u4_csr_reg[7]/P0001 ,
		_w2692_
	);
	LUT4 #(
		.INIT('h8caf)
	) name943 (
		\u1_u3_new_size_reg[5]/P0001 ,
		\u1_u3_new_size_reg[6]/P0001 ,
		\u4_csr_reg[5]/NET0131 ,
		\u4_csr_reg[6]/NET0131 ,
		_w2693_
	);
	LUT3 #(
		.INIT('h80)
	) name944 (
		_w2690_,
		_w2692_,
		_w2693_,
		_w2694_
	);
	LUT3 #(
		.INIT('h10)
	) name945 (
		_w2685_,
		_w2689_,
		_w2694_,
		_w2695_
	);
	LUT4 #(
		.INIT('h008c)
	) name946 (
		\u1_u3_new_size_reg[10]/P0001 ,
		\u1_u3_new_size_reg[9]/P0001 ,
		\u4_csr_reg[10]/P0001 ,
		\u4_csr_reg[9]/NET0131 ,
		_w2696_
	);
	LUT4 #(
		.INIT('h080a)
	) name947 (
		\u1_u3_new_size_reg[6]/P0001 ,
		\u1_u3_new_size_reg[7]/P0001 ,
		\u4_csr_reg[6]/NET0131 ,
		\u4_csr_reg[7]/P0001 ,
		_w2697_
	);
	LUT4 #(
		.INIT('hf531)
	) name948 (
		\u1_u3_new_size_reg[7]/P0001 ,
		\u1_u3_new_size_reg[8]/P0001 ,
		\u4_csr_reg[7]/P0001 ,
		\u4_csr_reg[8]/P0001 ,
		_w2698_
	);
	LUT4 #(
		.INIT('h2022)
	) name949 (
		_w2690_,
		_w2691_,
		_w2697_,
		_w2698_,
		_w2699_
	);
	LUT2 #(
		.INIT('h2)
	) name950 (
		\u1_u3_new_size_reg[10]/P0001 ,
		\u4_csr_reg[10]/P0001 ,
		_w2700_
	);
	LUT3 #(
		.INIT('h01)
	) name951 (
		\u1_u3_new_size_reg[11]/P0001 ,
		\u1_u3_new_size_reg[12]/P0001 ,
		\u1_u3_new_size_reg[13]/P0001 ,
		_w2701_
	);
	LUT2 #(
		.INIT('h4)
	) name952 (
		_w2700_,
		_w2701_,
		_w2702_
	);
	LUT3 #(
		.INIT('h10)
	) name953 (
		_w2696_,
		_w2699_,
		_w2702_,
		_w2703_
	);
	LUT2 #(
		.INIT('h4)
	) name954 (
		_w2695_,
		_w2703_,
		_w2704_
	);
	LUT4 #(
		.INIT('h10f0)
	) name955 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u1_buf1_reg[4]/P0001 ,
		\u4_u1_ep_match_r_reg/P0001 ,
		_w2705_
	);
	LUT4 #(
		.INIT('hc800)
	) name956 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_idin_reg[4]/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u1_ep_match_r_reg/P0001 ,
		_w2706_
	);
	LUT2 #(
		.INIT('h1)
	) name957 (
		_w2705_,
		_w2706_,
		_w2707_
	);
	LUT3 #(
		.INIT('h07)
	) name958 (
		_w2260_,
		_w2320_,
		_w2707_,
		_w2708_
	);
	LUT3 #(
		.INIT('h2a)
	) name959 (
		rst_i_pad,
		_w2260_,
		_w2648_,
		_w2709_
	);
	LUT2 #(
		.INIT('hb)
	) name960 (
		_w2708_,
		_w2709_,
		_w2710_
	);
	LUT4 #(
		.INIT('h10f0)
	) name961 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u1_buf1_reg[5]/P0001 ,
		\u4_u1_ep_match_r_reg/P0001 ,
		_w2711_
	);
	LUT4 #(
		.INIT('hc800)
	) name962 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_idin_reg[5]/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u1_ep_match_r_reg/P0001 ,
		_w2712_
	);
	LUT2 #(
		.INIT('h1)
	) name963 (
		_w2711_,
		_w2712_,
		_w2713_
	);
	LUT3 #(
		.INIT('h07)
	) name964 (
		_w2260_,
		_w2320_,
		_w2713_,
		_w2714_
	);
	LUT3 #(
		.INIT('h2a)
	) name965 (
		rst_i_pad,
		_w2260_,
		_w2655_,
		_w2715_
	);
	LUT2 #(
		.INIT('hb)
	) name966 (
		_w2714_,
		_w2715_,
		_w2716_
	);
	LUT4 #(
		.INIT('h10f0)
	) name967 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u1_buf1_reg[7]/P0001 ,
		\u4_u1_ep_match_r_reg/P0001 ,
		_w2717_
	);
	LUT4 #(
		.INIT('hc800)
	) name968 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_idin_reg[7]/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u1_ep_match_r_reg/P0001 ,
		_w2718_
	);
	LUT2 #(
		.INIT('h1)
	) name969 (
		_w2717_,
		_w2718_,
		_w2719_
	);
	LUT3 #(
		.INIT('h07)
	) name970 (
		_w2260_,
		_w2320_,
		_w2719_,
		_w2720_
	);
	LUT3 #(
		.INIT('h2a)
	) name971 (
		rst_i_pad,
		_w2260_,
		_w2662_,
		_w2721_
	);
	LUT2 #(
		.INIT('hb)
	) name972 (
		_w2720_,
		_w2721_,
		_w2722_
	);
	LUT4 #(
		.INIT('h10f0)
	) name973 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u2_buf1_reg[5]/P0001 ,
		\u4_u2_ep_match_r_reg/P0001 ,
		_w2723_
	);
	LUT4 #(
		.INIT('hc800)
	) name974 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_idin_reg[5]/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u2_ep_match_r_reg/P0001 ,
		_w2724_
	);
	LUT2 #(
		.INIT('h1)
	) name975 (
		_w2723_,
		_w2724_,
		_w2725_
	);
	LUT3 #(
		.INIT('h07)
	) name976 (
		_w2267_,
		_w2320_,
		_w2725_,
		_w2726_
	);
	LUT3 #(
		.INIT('h2a)
	) name977 (
		rst_i_pad,
		_w2267_,
		_w2655_,
		_w2727_
	);
	LUT2 #(
		.INIT('hb)
	) name978 (
		_w2726_,
		_w2727_,
		_w2728_
	);
	LUT4 #(
		.INIT('h10f0)
	) name979 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u2_buf1_reg[7]/P0001 ,
		\u4_u2_ep_match_r_reg/P0001 ,
		_w2729_
	);
	LUT4 #(
		.INIT('hc800)
	) name980 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_idin_reg[7]/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u2_ep_match_r_reg/P0001 ,
		_w2730_
	);
	LUT2 #(
		.INIT('h1)
	) name981 (
		_w2729_,
		_w2730_,
		_w2731_
	);
	LUT3 #(
		.INIT('h07)
	) name982 (
		_w2267_,
		_w2320_,
		_w2731_,
		_w2732_
	);
	LUT3 #(
		.INIT('h2a)
	) name983 (
		rst_i_pad,
		_w2267_,
		_w2662_,
		_w2733_
	);
	LUT2 #(
		.INIT('hb)
	) name984 (
		_w2732_,
		_w2733_,
		_w2734_
	);
	LUT4 #(
		.INIT('h10f0)
	) name985 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u2_buf1_reg[4]/P0001 ,
		\u4_u2_ep_match_r_reg/P0001 ,
		_w2735_
	);
	LUT4 #(
		.INIT('hc800)
	) name986 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_idin_reg[4]/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u2_ep_match_r_reg/P0001 ,
		_w2736_
	);
	LUT2 #(
		.INIT('h1)
	) name987 (
		_w2735_,
		_w2736_,
		_w2737_
	);
	LUT3 #(
		.INIT('h07)
	) name988 (
		_w2267_,
		_w2320_,
		_w2737_,
		_w2738_
	);
	LUT3 #(
		.INIT('h2a)
	) name989 (
		rst_i_pad,
		_w2267_,
		_w2648_,
		_w2739_
	);
	LUT2 #(
		.INIT('hb)
	) name990 (
		_w2738_,
		_w2739_,
		_w2740_
	);
	LUT4 #(
		.INIT('h0001)
	) name991 (
		\u1_u3_new_size_reg[3]/P0001 ,
		\u1_u3_new_size_reg[4]/P0001 ,
		\u1_u3_new_size_reg[5]/P0001 ,
		\u1_u3_new_size_reg[6]/P0001 ,
		_w2741_
	);
	LUT4 #(
		.INIT('h0001)
	) name992 (
		\u1_u3_new_size_reg[0]/P0001 ,
		\u1_u3_new_size_reg[10]/P0001 ,
		\u1_u3_new_size_reg[1]/P0001 ,
		\u1_u3_new_size_reg[2]/P0001 ,
		_w2742_
	);
	LUT4 #(
		.INIT('h0001)
	) name993 (
		\u1_u3_new_size_reg[11]/P0001 ,
		\u1_u3_new_size_reg[12]/P0001 ,
		\u1_u3_new_size_reg[13]/P0001 ,
		\u1_u3_new_size_reg[9]/P0001 ,
		_w2743_
	);
	LUT2 #(
		.INIT('h1)
	) name994 (
		\u1_u3_new_size_reg[7]/P0001 ,
		\u1_u3_new_size_reg[8]/P0001 ,
		_w2744_
	);
	LUT4 #(
		.INIT('h8000)
	) name995 (
		_w2741_,
		_w2742_,
		_w2743_,
		_w2744_,
		_w2745_
	);
	LUT2 #(
		.INIT('h1)
	) name996 (
		\u1_u2_sizd_c_reg[12]/P0001 ,
		\u1_u2_tx_dma_en_r_reg/P0001 ,
		_w2746_
	);
	LUT2 #(
		.INIT('h8)
	) name997 (
		\u1_u2_mack_r_reg/P0001 ,
		\u1_u2_state_reg[5]/NET0131 ,
		_w2747_
	);
	LUT3 #(
		.INIT('h20)
	) name998 (
		\u1_u2_mack_r_reg/P0001 ,
		\u1_u2_sizd_c_reg[0]/P0001 ,
		\u1_u2_state_reg[5]/NET0131 ,
		_w2748_
	);
	LUT2 #(
		.INIT('h1)
	) name999 (
		\u1_u2_sizd_c_reg[1]/P0001 ,
		\u1_u2_sizd_c_reg[2]/P0001 ,
		_w2749_
	);
	LUT4 #(
		.INIT('h0001)
	) name1000 (
		\u1_u2_sizd_c_reg[1]/P0001 ,
		\u1_u2_sizd_c_reg[2]/P0001 ,
		\u1_u2_sizd_c_reg[3]/P0001 ,
		\u1_u2_sizd_c_reg[4]/P0001 ,
		_w2750_
	);
	LUT2 #(
		.INIT('h1)
	) name1001 (
		\u1_u2_sizd_c_reg[5]/P0001 ,
		\u1_u2_sizd_c_reg[6]/P0001 ,
		_w2751_
	);
	LUT3 #(
		.INIT('h80)
	) name1002 (
		_w2748_,
		_w2750_,
		_w2751_,
		_w2752_
	);
	LUT4 #(
		.INIT('h0001)
	) name1003 (
		\u1_u2_sizd_c_reg[5]/P0001 ,
		\u1_u2_sizd_c_reg[6]/P0001 ,
		\u1_u2_sizd_c_reg[7]/P0001 ,
		\u1_u2_sizd_c_reg[8]/P0001 ,
		_w2753_
	);
	LUT2 #(
		.INIT('h8)
	) name1004 (
		_w2750_,
		_w2753_,
		_w2754_
	);
	LUT2 #(
		.INIT('h1)
	) name1005 (
		\u1_u2_sizd_c_reg[10]/P0001 ,
		\u1_u2_sizd_c_reg[11]/P0001 ,
		_w2755_
	);
	LUT3 #(
		.INIT('h01)
	) name1006 (
		\u1_u2_sizd_c_reg[12]/P0001 ,
		\u1_u2_sizd_c_reg[13]/P0001 ,
		\u1_u2_sizd_c_reg[9]/P0001 ,
		_w2756_
	);
	LUT4 #(
		.INIT('h8000)
	) name1007 (
		_w2750_,
		_w2753_,
		_w2755_,
		_w2756_,
		_w2757_
	);
	LUT4 #(
		.INIT('h0080)
	) name1008 (
		\u0_tx_ready_reg/NET0131 ,
		\u1_u1_state_reg[1]/NET0131 ,
		\u1_u1_tx_valid_r_reg/NET0131 ,
		\u1_u2_sizd_c_reg[0]/P0001 ,
		_w2758_
	);
	LUT3 #(
		.INIT('h80)
	) name1009 (
		_w2750_,
		_w2751_,
		_w2758_,
		_w2759_
	);
	LUT3 #(
		.INIT('h45)
	) name1010 (
		_w2752_,
		_w2757_,
		_w2759_,
		_w2760_
	);
	LUT3 #(
		.INIT('h01)
	) name1011 (
		\u1_u2_sizd_c_reg[7]/P0001 ,
		\u1_u2_sizd_c_reg[8]/P0001 ,
		\u1_u2_sizd_c_reg[9]/P0001 ,
		_w2761_
	);
	LUT2 #(
		.INIT('h8)
	) name1012 (
		_w2755_,
		_w2761_,
		_w2762_
	);
	LUT4 #(
		.INIT('hba00)
	) name1013 (
		_w2752_,
		_w2757_,
		_w2759_,
		_w2762_,
		_w2763_
	);
	LUT4 #(
		.INIT('h0010)
	) name1014 (
		\u1_u0_pid_reg[0]/NET0131 ,
		\u1_u0_pid_reg[1]/NET0131 ,
		\u1_u0_pid_reg[2]/NET0131 ,
		\u1_u0_pid_reg[3]/NET0131 ,
		_w2764_
	);
	LUT3 #(
		.INIT('h13)
	) name1015 (
		\u0_u0_mode_hs_reg/P0001 ,
		_w2119_,
		_w2764_,
		_w2765_
	);
	LUT4 #(
		.INIT('h0b00)
	) name1016 (
		_w2117_,
		_w2118_,
		_w2123_,
		_w2765_,
		_w2766_
	);
	LUT3 #(
		.INIT('h40)
	) name1017 (
		\u1_u3_state_reg[1]/P0001 ,
		_w2127_,
		_w2128_,
		_w2767_
	);
	LUT3 #(
		.INIT('ha2)
	) name1018 (
		\u1_u3_match_r_reg/P0001 ,
		\u4_csr_reg[22]/P0001 ,
		\u4_csr_reg[23]/P0001 ,
		_w2768_
	);
	LUT2 #(
		.INIT('h4)
	) name1019 (
		_w2131_,
		_w2768_,
		_w2769_
	);
	LUT3 #(
		.INIT('h10)
	) name1020 (
		_w2131_,
		_w2133_,
		_w2768_,
		_w2770_
	);
	LUT3 #(
		.INIT('h32)
	) name1021 (
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		_w2115_,
		_w2771_
	);
	LUT2 #(
		.INIT('h8)
	) name1022 (
		_w2770_,
		_w2771_,
		_w2772_
	);
	LUT3 #(
		.INIT('h80)
	) name1023 (
		_w2767_,
		_w2770_,
		_w2771_,
		_w2773_
	);
	LUT2 #(
		.INIT('h8)
	) name1024 (
		_w2766_,
		_w2773_,
		_w2774_
	);
	LUT4 #(
		.INIT('h0888)
	) name1025 (
		_w2746_,
		_w2763_,
		_w2766_,
		_w2773_,
		_w2775_
	);
	LUT2 #(
		.INIT('h2)
	) name1026 (
		\u1_u2_sizd_c_reg[12]/P0001 ,
		\u1_u2_tx_dma_en_r_reg/P0001 ,
		_w2776_
	);
	LUT4 #(
		.INIT('h1500)
	) name1027 (
		_w2763_,
		_w2766_,
		_w2773_,
		_w2776_,
		_w2777_
	);
	LUT3 #(
		.INIT('hfd)
	) name1028 (
		rst_i_pad,
		_w2775_,
		_w2777_,
		_w2778_
	);
	LUT3 #(
		.INIT('h15)
	) name1029 (
		\u1_u2_tx_dma_en_r_reg/P0001 ,
		_w2766_,
		_w2773_,
		_w2779_
	);
	LUT4 #(
		.INIT('h0008)
	) name1030 (
		\u1_u3_in_token_reg/NET0131 ,
		\u4_buf1_reg[18]/P0001 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		_w2780_
	);
	LUT3 #(
		.INIT('hc8)
	) name1031 (
		\u1_u3_buf0_na_reg/NET0131 ,
		\u4_buf1_reg[18]/P0001 ,
		\u4_csr_reg[30]/NET0131 ,
		_w2781_
	);
	LUT3 #(
		.INIT('h13)
	) name1032 (
		_w2352_,
		_w2780_,
		_w2781_,
		_w2782_
	);
	LUT4 #(
		.INIT('hccc4)
	) name1033 (
		\u1_u3_in_token_reg/NET0131 ,
		\u4_buf0_reg[18]/P0001 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		_w2783_
	);
	LUT3 #(
		.INIT('hd0)
	) name1034 (
		_w2352_,
		_w2353_,
		_w2783_,
		_w2784_
	);
	LUT2 #(
		.INIT('h2)
	) name1035 (
		_w2782_,
		_w2784_,
		_w2785_
	);
	LUT4 #(
		.INIT('h0008)
	) name1036 (
		\u1_u3_in_token_reg/NET0131 ,
		\u4_buf1_reg[17]/NET0131 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		_w2786_
	);
	LUT3 #(
		.INIT('hc8)
	) name1037 (
		\u1_u3_buf0_na_reg/NET0131 ,
		\u4_buf1_reg[17]/NET0131 ,
		\u4_csr_reg[30]/NET0131 ,
		_w2787_
	);
	LUT3 #(
		.INIT('h13)
	) name1038 (
		_w2352_,
		_w2786_,
		_w2787_,
		_w2788_
	);
	LUT4 #(
		.INIT('hccc4)
	) name1039 (
		\u1_u3_in_token_reg/NET0131 ,
		\u4_buf0_reg[17]/NET0131 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		_w2789_
	);
	LUT3 #(
		.INIT('hd0)
	) name1040 (
		_w2352_,
		_w2353_,
		_w2789_,
		_w2790_
	);
	LUT2 #(
		.INIT('h2)
	) name1041 (
		_w2788_,
		_w2790_,
		_w2791_
	);
	LUT3 #(
		.INIT('h08)
	) name1042 (
		\u4_csr_reg[0]/P0001 ,
		_w2788_,
		_w2790_,
		_w2792_
	);
	LUT4 #(
		.INIT('h0008)
	) name1043 (
		\u1_u3_in_token_reg/NET0131 ,
		\u4_buf1_reg[19]/NET0131 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		_w2793_
	);
	LUT3 #(
		.INIT('hc8)
	) name1044 (
		\u1_u3_buf0_na_reg/NET0131 ,
		\u4_buf1_reg[19]/NET0131 ,
		\u4_csr_reg[30]/NET0131 ,
		_w2794_
	);
	LUT3 #(
		.INIT('h13)
	) name1045 (
		_w2352_,
		_w2793_,
		_w2794_,
		_w2795_
	);
	LUT4 #(
		.INIT('hccc4)
	) name1046 (
		\u1_u3_in_token_reg/NET0131 ,
		\u4_buf0_reg[19]/NET0131 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		_w2796_
	);
	LUT3 #(
		.INIT('hd0)
	) name1047 (
		_w2352_,
		_w2353_,
		_w2796_,
		_w2797_
	);
	LUT2 #(
		.INIT('h2)
	) name1048 (
		_w2795_,
		_w2797_,
		_w2798_
	);
	LUT3 #(
		.INIT('h51)
	) name1049 (
		\u4_csr_reg[2]/NET0131 ,
		_w2795_,
		_w2797_,
		_w2799_
	);
	LUT4 #(
		.INIT('h00e8)
	) name1050 (
		\u4_csr_reg[1]/P0001 ,
		_w2785_,
		_w2792_,
		_w2799_,
		_w2800_
	);
	LUT4 #(
		.INIT('h0008)
	) name1051 (
		\u1_u3_in_token_reg/NET0131 ,
		\u4_buf1_reg[21]/NET0131 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		_w2801_
	);
	LUT3 #(
		.INIT('hc8)
	) name1052 (
		\u1_u3_buf0_na_reg/NET0131 ,
		\u4_buf1_reg[21]/NET0131 ,
		\u4_csr_reg[30]/NET0131 ,
		_w2802_
	);
	LUT3 #(
		.INIT('h13)
	) name1053 (
		_w2352_,
		_w2801_,
		_w2802_,
		_w2803_
	);
	LUT4 #(
		.INIT('hccc4)
	) name1054 (
		\u1_u3_in_token_reg/NET0131 ,
		\u4_buf0_reg[21]/NET0131 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		_w2804_
	);
	LUT3 #(
		.INIT('hd0)
	) name1055 (
		_w2352_,
		_w2353_,
		_w2804_,
		_w2805_
	);
	LUT2 #(
		.INIT('h2)
	) name1056 (
		_w2803_,
		_w2805_,
		_w2806_
	);
	LUT3 #(
		.INIT('h08)
	) name1057 (
		\u4_csr_reg[4]/NET0131 ,
		_w2803_,
		_w2805_,
		_w2807_
	);
	LUT4 #(
		.INIT('h0008)
	) name1058 (
		\u1_u3_in_token_reg/NET0131 ,
		\u4_buf1_reg[20]/NET0131 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		_w2808_
	);
	LUT3 #(
		.INIT('hc8)
	) name1059 (
		\u1_u3_buf0_na_reg/NET0131 ,
		\u4_buf1_reg[20]/NET0131 ,
		\u4_csr_reg[30]/NET0131 ,
		_w2809_
	);
	LUT3 #(
		.INIT('h13)
	) name1060 (
		_w2352_,
		_w2808_,
		_w2809_,
		_w2810_
	);
	LUT4 #(
		.INIT('hccc4)
	) name1061 (
		\u1_u3_in_token_reg/NET0131 ,
		\u4_buf0_reg[20]/NET0131 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		_w2811_
	);
	LUT3 #(
		.INIT('hd0)
	) name1062 (
		_w2352_,
		_w2353_,
		_w2811_,
		_w2812_
	);
	LUT2 #(
		.INIT('h2)
	) name1063 (
		_w2810_,
		_w2812_,
		_w2813_
	);
	LUT3 #(
		.INIT('h08)
	) name1064 (
		\u4_csr_reg[3]/P0001 ,
		_w2810_,
		_w2812_,
		_w2814_
	);
	LUT3 #(
		.INIT('h08)
	) name1065 (
		\u4_csr_reg[2]/NET0131 ,
		_w2795_,
		_w2797_,
		_w2815_
	);
	LUT3 #(
		.INIT('h01)
	) name1066 (
		_w2807_,
		_w2814_,
		_w2815_,
		_w2816_
	);
	LUT3 #(
		.INIT('h51)
	) name1067 (
		\u4_csr_reg[3]/P0001 ,
		_w2810_,
		_w2812_,
		_w2817_
	);
	LUT4 #(
		.INIT('h0008)
	) name1068 (
		\u1_u3_in_token_reg/NET0131 ,
		\u4_buf1_reg[22]/NET0131 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		_w2818_
	);
	LUT3 #(
		.INIT('hc8)
	) name1069 (
		\u1_u3_buf0_na_reg/NET0131 ,
		\u4_buf1_reg[22]/NET0131 ,
		\u4_csr_reg[30]/NET0131 ,
		_w2819_
	);
	LUT3 #(
		.INIT('h13)
	) name1070 (
		_w2352_,
		_w2818_,
		_w2819_,
		_w2820_
	);
	LUT4 #(
		.INIT('hccc4)
	) name1071 (
		\u1_u3_in_token_reg/NET0131 ,
		\u4_buf0_reg[22]/NET0131 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		_w2821_
	);
	LUT3 #(
		.INIT('hd0)
	) name1072 (
		_w2352_,
		_w2353_,
		_w2821_,
		_w2822_
	);
	LUT2 #(
		.INIT('h2)
	) name1073 (
		_w2820_,
		_w2822_,
		_w2823_
	);
	LUT3 #(
		.INIT('h51)
	) name1074 (
		\u4_csr_reg[5]/NET0131 ,
		_w2820_,
		_w2822_,
		_w2824_
	);
	LUT4 #(
		.INIT('h008e)
	) name1075 (
		\u4_csr_reg[4]/NET0131 ,
		_w2806_,
		_w2817_,
		_w2824_,
		_w2825_
	);
	LUT3 #(
		.INIT('hb0)
	) name1076 (
		_w2800_,
		_w2816_,
		_w2825_,
		_w2826_
	);
	LUT3 #(
		.INIT('h08)
	) name1077 (
		\u4_csr_reg[5]/NET0131 ,
		_w2820_,
		_w2822_,
		_w2827_
	);
	LUT4 #(
		.INIT('h0008)
	) name1078 (
		\u1_u3_in_token_reg/NET0131 ,
		\u4_buf1_reg[24]/NET0131 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		_w2828_
	);
	LUT3 #(
		.INIT('hc8)
	) name1079 (
		\u1_u3_buf0_na_reg/NET0131 ,
		\u4_buf1_reg[24]/NET0131 ,
		\u4_csr_reg[30]/NET0131 ,
		_w2829_
	);
	LUT3 #(
		.INIT('h13)
	) name1080 (
		_w2352_,
		_w2828_,
		_w2829_,
		_w2830_
	);
	LUT4 #(
		.INIT('hccc4)
	) name1081 (
		\u1_u3_in_token_reg/NET0131 ,
		\u4_buf0_reg[24]/NET0131 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		_w2831_
	);
	LUT3 #(
		.INIT('hd0)
	) name1082 (
		_w2352_,
		_w2353_,
		_w2831_,
		_w2832_
	);
	LUT2 #(
		.INIT('h2)
	) name1083 (
		_w2830_,
		_w2832_,
		_w2833_
	);
	LUT3 #(
		.INIT('h08)
	) name1084 (
		\u4_csr_reg[7]/P0001 ,
		_w2830_,
		_w2832_,
		_w2834_
	);
	LUT4 #(
		.INIT('h0008)
	) name1085 (
		\u1_u3_in_token_reg/NET0131 ,
		\u4_buf1_reg[25]/NET0131 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		_w2835_
	);
	LUT3 #(
		.INIT('hc8)
	) name1086 (
		\u1_u3_buf0_na_reg/NET0131 ,
		\u4_buf1_reg[25]/NET0131 ,
		\u4_csr_reg[30]/NET0131 ,
		_w2836_
	);
	LUT3 #(
		.INIT('h13)
	) name1087 (
		_w2352_,
		_w2835_,
		_w2836_,
		_w2837_
	);
	LUT4 #(
		.INIT('hccc4)
	) name1088 (
		\u1_u3_in_token_reg/NET0131 ,
		\u4_buf0_reg[25]/NET0131 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		_w2838_
	);
	LUT3 #(
		.INIT('hd0)
	) name1089 (
		_w2352_,
		_w2353_,
		_w2838_,
		_w2839_
	);
	LUT2 #(
		.INIT('h2)
	) name1090 (
		_w2837_,
		_w2839_,
		_w2840_
	);
	LUT3 #(
		.INIT('h08)
	) name1091 (
		\u4_csr_reg[8]/P0001 ,
		_w2837_,
		_w2839_,
		_w2841_
	);
	LUT2 #(
		.INIT('h1)
	) name1092 (
		_w2834_,
		_w2841_,
		_w2842_
	);
	LUT4 #(
		.INIT('h0008)
	) name1093 (
		\u1_u3_in_token_reg/NET0131 ,
		\u4_buf1_reg[27]/P0001 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		_w2843_
	);
	LUT3 #(
		.INIT('hc8)
	) name1094 (
		\u1_u3_buf0_na_reg/NET0131 ,
		\u4_buf1_reg[27]/P0001 ,
		\u4_csr_reg[30]/NET0131 ,
		_w2844_
	);
	LUT3 #(
		.INIT('h13)
	) name1095 (
		_w2352_,
		_w2843_,
		_w2844_,
		_w2845_
	);
	LUT4 #(
		.INIT('hccc4)
	) name1096 (
		\u1_u3_in_token_reg/NET0131 ,
		\u4_buf0_reg[27]/P0001 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		_w2846_
	);
	LUT3 #(
		.INIT('hd0)
	) name1097 (
		_w2352_,
		_w2353_,
		_w2846_,
		_w2847_
	);
	LUT2 #(
		.INIT('h2)
	) name1098 (
		_w2845_,
		_w2847_,
		_w2848_
	);
	LUT3 #(
		.INIT('h08)
	) name1099 (
		\u4_csr_reg[10]/P0001 ,
		_w2845_,
		_w2847_,
		_w2849_
	);
	LUT4 #(
		.INIT('h0008)
	) name1100 (
		\u1_u3_in_token_reg/NET0131 ,
		\u4_buf1_reg[26]/NET0131 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		_w2850_
	);
	LUT3 #(
		.INIT('hc8)
	) name1101 (
		\u1_u3_buf0_na_reg/NET0131 ,
		\u4_buf1_reg[26]/NET0131 ,
		\u4_csr_reg[30]/NET0131 ,
		_w2851_
	);
	LUT3 #(
		.INIT('h13)
	) name1102 (
		_w2352_,
		_w2850_,
		_w2851_,
		_w2852_
	);
	LUT4 #(
		.INIT('hccc4)
	) name1103 (
		\u1_u3_in_token_reg/NET0131 ,
		\u4_buf0_reg[26]/NET0131 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		_w2853_
	);
	LUT3 #(
		.INIT('hd0)
	) name1104 (
		_w2352_,
		_w2353_,
		_w2853_,
		_w2854_
	);
	LUT2 #(
		.INIT('h2)
	) name1105 (
		_w2852_,
		_w2854_,
		_w2855_
	);
	LUT3 #(
		.INIT('h08)
	) name1106 (
		\u4_csr_reg[9]/NET0131 ,
		_w2852_,
		_w2854_,
		_w2856_
	);
	LUT2 #(
		.INIT('h1)
	) name1107 (
		_w2849_,
		_w2856_,
		_w2857_
	);
	LUT4 #(
		.INIT('h0008)
	) name1108 (
		\u1_u3_in_token_reg/NET0131 ,
		\u4_buf1_reg[23]/NET0131 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		_w2858_
	);
	LUT3 #(
		.INIT('hc8)
	) name1109 (
		\u1_u3_buf0_na_reg/NET0131 ,
		\u4_buf1_reg[23]/NET0131 ,
		\u4_csr_reg[30]/NET0131 ,
		_w2859_
	);
	LUT3 #(
		.INIT('h13)
	) name1110 (
		_w2352_,
		_w2858_,
		_w2859_,
		_w2860_
	);
	LUT4 #(
		.INIT('hccc4)
	) name1111 (
		\u1_u3_in_token_reg/NET0131 ,
		\u4_buf0_reg[23]/NET0131 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		_w2861_
	);
	LUT3 #(
		.INIT('hd0)
	) name1112 (
		_w2352_,
		_w2353_,
		_w2861_,
		_w2862_
	);
	LUT2 #(
		.INIT('h2)
	) name1113 (
		_w2860_,
		_w2862_,
		_w2863_
	);
	LUT3 #(
		.INIT('h08)
	) name1114 (
		\u4_csr_reg[6]/NET0131 ,
		_w2860_,
		_w2862_,
		_w2864_
	);
	LUT3 #(
		.INIT('h01)
	) name1115 (
		_w2849_,
		_w2856_,
		_w2864_,
		_w2865_
	);
	LUT3 #(
		.INIT('h40)
	) name1116 (
		_w2827_,
		_w2842_,
		_w2865_,
		_w2866_
	);
	LUT3 #(
		.INIT('h51)
	) name1117 (
		\u4_csr_reg[6]/NET0131 ,
		_w2860_,
		_w2862_,
		_w2867_
	);
	LUT4 #(
		.INIT('h0701)
	) name1118 (
		\u4_csr_reg[7]/P0001 ,
		_w2833_,
		_w2841_,
		_w2867_,
		_w2868_
	);
	LUT3 #(
		.INIT('h51)
	) name1119 (
		\u4_csr_reg[9]/NET0131 ,
		_w2852_,
		_w2854_,
		_w2869_
	);
	LUT3 #(
		.INIT('h51)
	) name1120 (
		\u4_csr_reg[8]/P0001 ,
		_w2837_,
		_w2839_,
		_w2870_
	);
	LUT2 #(
		.INIT('h1)
	) name1121 (
		_w2869_,
		_w2870_,
		_w2871_
	);
	LUT3 #(
		.INIT('h51)
	) name1122 (
		\u4_csr_reg[10]/P0001 ,
		_w2845_,
		_w2847_,
		_w2872_
	);
	LUT4 #(
		.INIT('h0008)
	) name1123 (
		\u1_u3_in_token_reg/NET0131 ,
		\u4_buf1_reg[29]/P0001 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		_w2873_
	);
	LUT3 #(
		.INIT('hc8)
	) name1124 (
		\u1_u3_buf0_na_reg/NET0131 ,
		\u4_buf1_reg[29]/P0001 ,
		\u4_csr_reg[30]/NET0131 ,
		_w2874_
	);
	LUT3 #(
		.INIT('h13)
	) name1125 (
		_w2352_,
		_w2873_,
		_w2874_,
		_w2875_
	);
	LUT4 #(
		.INIT('hccc4)
	) name1126 (
		\u1_u3_in_token_reg/NET0131 ,
		\u4_buf0_reg[29]/P0001 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		_w2876_
	);
	LUT3 #(
		.INIT('hd0)
	) name1127 (
		_w2352_,
		_w2353_,
		_w2876_,
		_w2877_
	);
	LUT2 #(
		.INIT('h2)
	) name1128 (
		_w2875_,
		_w2877_,
		_w2878_
	);
	LUT4 #(
		.INIT('h0008)
	) name1129 (
		\u1_u3_in_token_reg/NET0131 ,
		\u4_buf1_reg[28]/P0001 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		_w2879_
	);
	LUT3 #(
		.INIT('hc8)
	) name1130 (
		\u1_u3_buf0_na_reg/NET0131 ,
		\u4_buf1_reg[28]/P0001 ,
		\u4_csr_reg[30]/NET0131 ,
		_w2880_
	);
	LUT3 #(
		.INIT('h13)
	) name1131 (
		_w2352_,
		_w2879_,
		_w2880_,
		_w2881_
	);
	LUT4 #(
		.INIT('hccc4)
	) name1132 (
		\u1_u3_in_token_reg/NET0131 ,
		\u4_buf0_reg[28]/P0001 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		_w2882_
	);
	LUT3 #(
		.INIT('hd0)
	) name1133 (
		_w2352_,
		_w2353_,
		_w2882_,
		_w2883_
	);
	LUT2 #(
		.INIT('h2)
	) name1134 (
		_w2881_,
		_w2883_,
		_w2884_
	);
	LUT4 #(
		.INIT('h0020)
	) name1135 (
		_w2875_,
		_w2877_,
		_w2881_,
		_w2883_,
		_w2885_
	);
	LUT4 #(
		.INIT('h0008)
	) name1136 (
		\u1_u3_in_token_reg/NET0131 ,
		\u4_buf1_reg[30]/P0001 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		_w2886_
	);
	LUT3 #(
		.INIT('hc8)
	) name1137 (
		\u1_u3_buf0_na_reg/NET0131 ,
		\u4_buf1_reg[30]/P0001 ,
		\u4_csr_reg[30]/NET0131 ,
		_w2887_
	);
	LUT3 #(
		.INIT('h13)
	) name1138 (
		_w2352_,
		_w2886_,
		_w2887_,
		_w2888_
	);
	LUT4 #(
		.INIT('hccc4)
	) name1139 (
		\u1_u3_in_token_reg/NET0131 ,
		\u4_buf0_reg[30]/P0001 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		_w2889_
	);
	LUT3 #(
		.INIT('hd0)
	) name1140 (
		_w2352_,
		_w2353_,
		_w2889_,
		_w2890_
	);
	LUT2 #(
		.INIT('h2)
	) name1141 (
		_w2888_,
		_w2890_,
		_w2891_
	);
	LUT2 #(
		.INIT('h8)
	) name1142 (
		_w2885_,
		_w2891_,
		_w2892_
	);
	LUT3 #(
		.INIT('h40)
	) name1143 (
		_w2872_,
		_w2885_,
		_w2891_,
		_w2893_
	);
	LUT4 #(
		.INIT('h1000)
	) name1144 (
		_w2791_,
		_w2872_,
		_w2885_,
		_w2891_,
		_w2894_
	);
	LUT4 #(
		.INIT('h7500)
	) name1145 (
		_w2857_,
		_w2868_,
		_w2871_,
		_w2894_,
		_w2895_
	);
	LUT3 #(
		.INIT('hb0)
	) name1146 (
		_w2826_,
		_w2866_,
		_w2895_,
		_w2896_
	);
	LUT4 #(
		.INIT('h4500)
	) name1147 (
		_w2779_,
		_w2826_,
		_w2866_,
		_w2895_,
		_w2897_
	);
	LUT4 #(
		.INIT('h7500)
	) name1148 (
		_w2857_,
		_w2868_,
		_w2871_,
		_w2893_,
		_w2898_
	);
	LUT4 #(
		.INIT('hc888)
	) name1149 (
		\u1_u2_tx_dma_en_r_reg/P0001 ,
		\u4_csr_reg[0]/P0001 ,
		_w2766_,
		_w2773_,
		_w2899_
	);
	LUT4 #(
		.INIT('h4f00)
	) name1150 (
		_w2826_,
		_w2866_,
		_w2898_,
		_w2899_,
		_w2900_
	);
	LUT3 #(
		.INIT('h13)
	) name1151 (
		\u1_u2_mack_r_reg/P0001 ,
		\u1_u2_sizd_c_reg[0]/P0001 ,
		\u1_u2_state_reg[5]/NET0131 ,
		_w2901_
	);
	LUT4 #(
		.INIT('h8000)
	) name1152 (
		\u0_tx_ready_reg/NET0131 ,
		\u1_u1_state_reg[1]/NET0131 ,
		\u1_u1_tx_valid_r_reg/NET0131 ,
		\u1_u2_sizd_c_reg[0]/P0001 ,
		_w2902_
	);
	LUT4 #(
		.INIT('h005e)
	) name1153 (
		\u1_u2_sizd_c_reg[0]/P0001 ,
		_w1762_,
		_w2747_,
		_w2902_,
		_w2903_
	);
	LUT4 #(
		.INIT('h1500)
	) name1154 (
		\u1_u2_tx_dma_en_r_reg/P0001 ,
		_w2757_,
		_w2901_,
		_w2903_,
		_w2904_
	);
	LUT4 #(
		.INIT('h80aa)
	) name1155 (
		rst_i_pad,
		_w2766_,
		_w2773_,
		_w2904_,
		_w2905_
	);
	LUT3 #(
		.INIT('hef)
	) name1156 (
		_w2897_,
		_w2900_,
		_w2905_,
		_w2906_
	);
	LUT4 #(
		.INIT('h0020)
	) name1157 (
		_w2845_,
		_w2847_,
		_w2888_,
		_w2890_,
		_w2907_
	);
	LUT2 #(
		.INIT('h8)
	) name1158 (
		_w2885_,
		_w2907_,
		_w2908_
	);
	LUT4 #(
		.INIT('hc888)
	) name1159 (
		\u1_u2_tx_dma_en_r_reg/P0001 ,
		\u4_csr_reg[10]/P0001 ,
		_w2766_,
		_w2773_,
		_w2909_
	);
	LUT4 #(
		.INIT('h4f00)
	) name1160 (
		_w2826_,
		_w2866_,
		_w2908_,
		_w2909_,
		_w2910_
	);
	LUT4 #(
		.INIT('ha888)
	) name1161 (
		rst_i_pad,
		\u1_u2_tx_dma_en_r_reg/P0001 ,
		_w2766_,
		_w2773_,
		_w2911_
	);
	LUT2 #(
		.INIT('h8)
	) name1162 (
		rst_i_pad,
		\u1_u2_sizd_c_reg[10]/P0001 ,
		_w2912_
	);
	LUT2 #(
		.INIT('h8)
	) name1163 (
		_w2761_,
		_w2912_,
		_w2913_
	);
	LUT4 #(
		.INIT('hba00)
	) name1164 (
		_w2752_,
		_w2757_,
		_w2759_,
		_w2913_,
		_w2914_
	);
	LUT4 #(
		.INIT('hba00)
	) name1165 (
		_w2752_,
		_w2757_,
		_w2759_,
		_w2761_,
		_w2915_
	);
	LUT2 #(
		.INIT('h2)
	) name1166 (
		rst_i_pad,
		\u1_u2_sizd_c_reg[10]/P0001 ,
		_w2916_
	);
	LUT3 #(
		.INIT('h45)
	) name1167 (
		_w2914_,
		_w2915_,
		_w2916_,
		_w2917_
	);
	LUT2 #(
		.INIT('h4)
	) name1168 (
		_w2911_,
		_w2917_,
		_w2918_
	);
	LUT2 #(
		.INIT('he)
	) name1169 (
		_w2910_,
		_w2918_,
		_w2919_
	);
	LUT4 #(
		.INIT('h0001)
	) name1170 (
		\u1_u2_sizd_c_reg[10]/P0001 ,
		\u1_u2_sizd_c_reg[7]/P0001 ,
		\u1_u2_sizd_c_reg[8]/P0001 ,
		\u1_u2_sizd_c_reg[9]/P0001 ,
		_w2920_
	);
	LUT4 #(
		.INIT('hba00)
	) name1171 (
		_w2752_,
		_w2757_,
		_w2759_,
		_w2920_,
		_w2921_
	);
	LUT3 #(
		.INIT('h7d)
	) name1172 (
		rst_i_pad,
		\u1_u2_sizd_c_reg[11]/P0001 ,
		_w2921_,
		_w2922_
	);
	LUT2 #(
		.INIT('h4)
	) name1173 (
		_w2911_,
		_w2922_,
		_w2923_
	);
	LUT3 #(
		.INIT('h01)
	) name1174 (
		\u1_u2_sizd_c_reg[11]/P0001 ,
		\u1_u2_sizd_c_reg[12]/P0001 ,
		\u1_u2_sizd_c_reg[13]/P0001 ,
		_w2924_
	);
	LUT2 #(
		.INIT('h8)
	) name1175 (
		_w2921_,
		_w2924_,
		_w2925_
	);
	LUT2 #(
		.INIT('h8)
	) name1176 (
		_w2779_,
		_w2925_,
		_w2926_
	);
	LUT2 #(
		.INIT('h1)
	) name1177 (
		\u1_u2_sizd_c_reg[11]/P0001 ,
		\u1_u2_sizd_c_reg[12]/P0001 ,
		_w2927_
	);
	LUT2 #(
		.INIT('h8)
	) name1178 (
		_w2921_,
		_w2927_,
		_w2928_
	);
	LUT2 #(
		.INIT('h2)
	) name1179 (
		\u1_u2_sizd_c_reg[13]/P0001 ,
		\u1_u2_tx_dma_en_r_reg/P0001 ,
		_w2929_
	);
	LUT3 #(
		.INIT('h70)
	) name1180 (
		_w2766_,
		_w2773_,
		_w2929_,
		_w2930_
	);
	LUT3 #(
		.INIT('h8a)
	) name1181 (
		rst_i_pad,
		_w2928_,
		_w2930_,
		_w2931_
	);
	LUT2 #(
		.INIT('hb)
	) name1182 (
		_w2926_,
		_w2931_,
		_w2932_
	);
	LUT4 #(
		.INIT('h1000)
	) name1183 (
		_w2798_,
		_w2872_,
		_w2885_,
		_w2891_,
		_w2933_
	);
	LUT4 #(
		.INIT('h7500)
	) name1184 (
		_w2857_,
		_w2868_,
		_w2871_,
		_w2933_,
		_w2934_
	);
	LUT3 #(
		.INIT('hb0)
	) name1185 (
		_w2826_,
		_w2866_,
		_w2934_,
		_w2935_
	);
	LUT4 #(
		.INIT('h4500)
	) name1186 (
		_w2779_,
		_w2826_,
		_w2866_,
		_w2934_,
		_w2936_
	);
	LUT4 #(
		.INIT('hc888)
	) name1187 (
		\u1_u2_tx_dma_en_r_reg/P0001 ,
		\u4_csr_reg[2]/NET0131 ,
		_w2766_,
		_w2773_,
		_w2937_
	);
	LUT4 #(
		.INIT('h4f00)
	) name1188 (
		_w2826_,
		_w2866_,
		_w2898_,
		_w2937_,
		_w2938_
	);
	LUT4 #(
		.INIT('h0200)
	) name1189 (
		\u1_u2_mack_r_reg/P0001 ,
		\u1_u2_sizd_c_reg[0]/P0001 ,
		\u1_u2_sizd_c_reg[1]/P0001 ,
		\u1_u2_state_reg[5]/NET0131 ,
		_w2939_
	);
	LUT2 #(
		.INIT('h4)
	) name1190 (
		\u1_u2_sizd_c_reg[1]/P0001 ,
		_w2758_,
		_w2940_
	);
	LUT4 #(
		.INIT('h080a)
	) name1191 (
		\u1_u2_sizd_c_reg[2]/P0001 ,
		_w2757_,
		_w2939_,
		_w2940_,
		_w2941_
	);
	LUT2 #(
		.INIT('h8)
	) name1192 (
		_w2748_,
		_w2749_,
		_w2942_
	);
	LUT2 #(
		.INIT('h8)
	) name1193 (
		_w2749_,
		_w2758_,
		_w2943_
	);
	LUT3 #(
		.INIT('h23)
	) name1194 (
		_w2757_,
		_w2942_,
		_w2943_,
		_w2944_
	);
	LUT2 #(
		.INIT('h4)
	) name1195 (
		_w2941_,
		_w2944_,
		_w2945_
	);
	LUT3 #(
		.INIT('ha2)
	) name1196 (
		rst_i_pad,
		_w2779_,
		_w2945_,
		_w2946_
	);
	LUT3 #(
		.INIT('hef)
	) name1197 (
		_w2936_,
		_w2938_,
		_w2946_,
		_w2947_
	);
	LUT4 #(
		.INIT('h1000)
	) name1198 (
		_w2813_,
		_w2872_,
		_w2885_,
		_w2891_,
		_w2948_
	);
	LUT4 #(
		.INIT('h7500)
	) name1199 (
		_w2857_,
		_w2868_,
		_w2871_,
		_w2948_,
		_w2949_
	);
	LUT3 #(
		.INIT('hb0)
	) name1200 (
		_w2826_,
		_w2866_,
		_w2949_,
		_w2950_
	);
	LUT4 #(
		.INIT('h4500)
	) name1201 (
		_w2779_,
		_w2826_,
		_w2866_,
		_w2949_,
		_w2951_
	);
	LUT4 #(
		.INIT('hc888)
	) name1202 (
		\u1_u2_tx_dma_en_r_reg/P0001 ,
		\u4_csr_reg[3]/P0001 ,
		_w2766_,
		_w2773_,
		_w2952_
	);
	LUT4 #(
		.INIT('h4f00)
	) name1203 (
		_w2826_,
		_w2866_,
		_w2898_,
		_w2952_,
		_w2953_
	);
	LUT4 #(
		.INIT('h5150)
	) name1204 (
		\u1_u2_sizd_c_reg[3]/P0001 ,
		_w2757_,
		_w2942_,
		_w2943_,
		_w2954_
	);
	LUT4 #(
		.INIT('ha6a5)
	) name1205 (
		\u1_u2_sizd_c_reg[3]/P0001 ,
		_w2757_,
		_w2942_,
		_w2943_,
		_w2955_
	);
	LUT4 #(
		.INIT('h0015)
	) name1206 (
		\u1_u2_tx_dma_en_r_reg/P0001 ,
		_w2766_,
		_w2773_,
		_w2955_,
		_w2956_
	);
	LUT2 #(
		.INIT('h2)
	) name1207 (
		rst_i_pad,
		_w2956_,
		_w2957_
	);
	LUT3 #(
		.INIT('hef)
	) name1208 (
		_w2951_,
		_w2953_,
		_w2957_,
		_w2958_
	);
	LUT4 #(
		.INIT('h1000)
	) name1209 (
		_w2806_,
		_w2872_,
		_w2885_,
		_w2891_,
		_w2959_
	);
	LUT4 #(
		.INIT('h7500)
	) name1210 (
		_w2857_,
		_w2868_,
		_w2871_,
		_w2959_,
		_w2960_
	);
	LUT3 #(
		.INIT('hb0)
	) name1211 (
		_w2826_,
		_w2866_,
		_w2960_,
		_w2961_
	);
	LUT4 #(
		.INIT('h4500)
	) name1212 (
		_w2779_,
		_w2826_,
		_w2866_,
		_w2960_,
		_w2962_
	);
	LUT4 #(
		.INIT('hc888)
	) name1213 (
		\u1_u2_tx_dma_en_r_reg/P0001 ,
		\u4_csr_reg[4]/NET0131 ,
		_w2766_,
		_w2773_,
		_w2963_
	);
	LUT4 #(
		.INIT('h4f00)
	) name1214 (
		_w2826_,
		_w2866_,
		_w2898_,
		_w2963_,
		_w2964_
	);
	LUT2 #(
		.INIT('h8)
	) name1215 (
		_w2748_,
		_w2750_,
		_w2965_
	);
	LUT2 #(
		.INIT('h8)
	) name1216 (
		_w2750_,
		_w2758_,
		_w2966_
	);
	LUT4 #(
		.INIT('h080a)
	) name1217 (
		rst_i_pad,
		_w2757_,
		_w2965_,
		_w2966_,
		_w2967_
	);
	LUT3 #(
		.INIT('hd0)
	) name1218 (
		\u1_u2_sizd_c_reg[4]/P0001 ,
		_w2954_,
		_w2967_,
		_w2968_
	);
	LUT2 #(
		.INIT('h1)
	) name1219 (
		_w2911_,
		_w2968_,
		_w2969_
	);
	LUT3 #(
		.INIT('hfe)
	) name1220 (
		_w2962_,
		_w2964_,
		_w2969_,
		_w2970_
	);
	LUT4 #(
		.INIT('h1000)
	) name1221 (
		_w2823_,
		_w2872_,
		_w2885_,
		_w2891_,
		_w2971_
	);
	LUT4 #(
		.INIT('h7500)
	) name1222 (
		_w2857_,
		_w2868_,
		_w2871_,
		_w2971_,
		_w2972_
	);
	LUT3 #(
		.INIT('hb0)
	) name1223 (
		_w2826_,
		_w2866_,
		_w2972_,
		_w2973_
	);
	LUT4 #(
		.INIT('h4500)
	) name1224 (
		_w2779_,
		_w2826_,
		_w2866_,
		_w2972_,
		_w2974_
	);
	LUT4 #(
		.INIT('hc888)
	) name1225 (
		\u1_u2_tx_dma_en_r_reg/P0001 ,
		\u4_csr_reg[5]/NET0131 ,
		_w2766_,
		_w2773_,
		_w2975_
	);
	LUT4 #(
		.INIT('h4f00)
	) name1226 (
		_w2826_,
		_w2866_,
		_w2898_,
		_w2975_,
		_w2976_
	);
	LUT4 #(
		.INIT('h5150)
	) name1227 (
		\u1_u2_sizd_c_reg[5]/P0001 ,
		_w2757_,
		_w2965_,
		_w2966_,
		_w2977_
	);
	LUT4 #(
		.INIT('ha6a5)
	) name1228 (
		\u1_u2_sizd_c_reg[5]/P0001 ,
		_w2757_,
		_w2965_,
		_w2966_,
		_w2978_
	);
	LUT4 #(
		.INIT('h0015)
	) name1229 (
		\u1_u2_tx_dma_en_r_reg/P0001 ,
		_w2766_,
		_w2773_,
		_w2978_,
		_w2979_
	);
	LUT2 #(
		.INIT('h2)
	) name1230 (
		rst_i_pad,
		_w2979_,
		_w2980_
	);
	LUT3 #(
		.INIT('hef)
	) name1231 (
		_w2974_,
		_w2976_,
		_w2980_,
		_w2981_
	);
	LUT4 #(
		.INIT('h1000)
	) name1232 (
		_w2863_,
		_w2872_,
		_w2885_,
		_w2891_,
		_w2982_
	);
	LUT4 #(
		.INIT('h7500)
	) name1233 (
		_w2857_,
		_w2868_,
		_w2871_,
		_w2982_,
		_w2983_
	);
	LUT3 #(
		.INIT('hb0)
	) name1234 (
		_w2826_,
		_w2866_,
		_w2983_,
		_w2984_
	);
	LUT4 #(
		.INIT('h4500)
	) name1235 (
		_w2779_,
		_w2826_,
		_w2866_,
		_w2983_,
		_w2985_
	);
	LUT4 #(
		.INIT('hc888)
	) name1236 (
		\u1_u2_tx_dma_en_r_reg/P0001 ,
		\u4_csr_reg[6]/NET0131 ,
		_w2766_,
		_w2773_,
		_w2986_
	);
	LUT4 #(
		.INIT('h4f00)
	) name1237 (
		_w2826_,
		_w2866_,
		_w2898_,
		_w2986_,
		_w2987_
	);
	LUT4 #(
		.INIT('h2022)
	) name1238 (
		rst_i_pad,
		_w2752_,
		_w2757_,
		_w2759_,
		_w2988_
	);
	LUT3 #(
		.INIT('hd0)
	) name1239 (
		\u1_u2_sizd_c_reg[6]/P0001 ,
		_w2977_,
		_w2988_,
		_w2989_
	);
	LUT2 #(
		.INIT('h1)
	) name1240 (
		_w2911_,
		_w2989_,
		_w2990_
	);
	LUT3 #(
		.INIT('hfe)
	) name1241 (
		_w2985_,
		_w2987_,
		_w2990_,
		_w2991_
	);
	LUT4 #(
		.INIT('h1000)
	) name1242 (
		_w2833_,
		_w2872_,
		_w2885_,
		_w2891_,
		_w2992_
	);
	LUT4 #(
		.INIT('h7500)
	) name1243 (
		_w2857_,
		_w2868_,
		_w2871_,
		_w2992_,
		_w2993_
	);
	LUT3 #(
		.INIT('hb0)
	) name1244 (
		_w2826_,
		_w2866_,
		_w2993_,
		_w2994_
	);
	LUT4 #(
		.INIT('h4500)
	) name1245 (
		_w2779_,
		_w2826_,
		_w2866_,
		_w2993_,
		_w2995_
	);
	LUT4 #(
		.INIT('hc888)
	) name1246 (
		\u1_u2_tx_dma_en_r_reg/P0001 ,
		\u4_csr_reg[7]/P0001 ,
		_w2766_,
		_w2773_,
		_w2996_
	);
	LUT4 #(
		.INIT('h4f00)
	) name1247 (
		_w2826_,
		_w2866_,
		_w2898_,
		_w2996_,
		_w2997_
	);
	LUT4 #(
		.INIT('h9a99)
	) name1248 (
		\u1_u2_sizd_c_reg[7]/P0001 ,
		_w2752_,
		_w2757_,
		_w2759_,
		_w2998_
	);
	LUT4 #(
		.INIT('h0015)
	) name1249 (
		\u1_u2_tx_dma_en_r_reg/P0001 ,
		_w2766_,
		_w2773_,
		_w2998_,
		_w2999_
	);
	LUT2 #(
		.INIT('h2)
	) name1250 (
		rst_i_pad,
		_w2999_,
		_w3000_
	);
	LUT3 #(
		.INIT('hef)
	) name1251 (
		_w2995_,
		_w2997_,
		_w3000_,
		_w3001_
	);
	LUT4 #(
		.INIT('h1000)
	) name1252 (
		_w2840_,
		_w2872_,
		_w2885_,
		_w2891_,
		_w3002_
	);
	LUT4 #(
		.INIT('h7500)
	) name1253 (
		_w2857_,
		_w2868_,
		_w2871_,
		_w3002_,
		_w3003_
	);
	LUT3 #(
		.INIT('hb0)
	) name1254 (
		_w2826_,
		_w2866_,
		_w3003_,
		_w3004_
	);
	LUT4 #(
		.INIT('h4500)
	) name1255 (
		_w2779_,
		_w2826_,
		_w2866_,
		_w3003_,
		_w3005_
	);
	LUT4 #(
		.INIT('hc888)
	) name1256 (
		\u1_u2_tx_dma_en_r_reg/P0001 ,
		\u4_csr_reg[8]/P0001 ,
		_w2766_,
		_w2773_,
		_w3006_
	);
	LUT4 #(
		.INIT('h4f00)
	) name1257 (
		_w2826_,
		_w2866_,
		_w2898_,
		_w3006_,
		_w3007_
	);
	LUT4 #(
		.INIT('h0a28)
	) name1258 (
		rst_i_pad,
		\u1_u2_sizd_c_reg[7]/P0001 ,
		\u1_u2_sizd_c_reg[8]/P0001 ,
		_w2760_,
		_w3008_
	);
	LUT2 #(
		.INIT('h1)
	) name1259 (
		_w2911_,
		_w3008_,
		_w3009_
	);
	LUT3 #(
		.INIT('hfe)
	) name1260 (
		_w3005_,
		_w3007_,
		_w3009_,
		_w3010_
	);
	LUT4 #(
		.INIT('h1000)
	) name1261 (
		_w2855_,
		_w2872_,
		_w2885_,
		_w2891_,
		_w3011_
	);
	LUT4 #(
		.INIT('h7500)
	) name1262 (
		_w2857_,
		_w2868_,
		_w2871_,
		_w3011_,
		_w3012_
	);
	LUT3 #(
		.INIT('hb0)
	) name1263 (
		_w2826_,
		_w2866_,
		_w3012_,
		_w3013_
	);
	LUT4 #(
		.INIT('h4500)
	) name1264 (
		_w2779_,
		_w2826_,
		_w2866_,
		_w3012_,
		_w3014_
	);
	LUT4 #(
		.INIT('hc888)
	) name1265 (
		\u1_u2_tx_dma_en_r_reg/P0001 ,
		\u4_csr_reg[9]/NET0131 ,
		_w2766_,
		_w2773_,
		_w3015_
	);
	LUT4 #(
		.INIT('h4f00)
	) name1266 (
		_w2826_,
		_w2866_,
		_w2898_,
		_w3015_,
		_w3016_
	);
	LUT3 #(
		.INIT('h80)
	) name1267 (
		_w2748_,
		_w2750_,
		_w2753_,
		_w3017_
	);
	LUT3 #(
		.INIT('h70)
	) name1268 (
		_w2755_,
		_w2756_,
		_w2758_,
		_w3018_
	);
	LUT4 #(
		.INIT('ha9a5)
	) name1269 (
		\u1_u2_sizd_c_reg[9]/P0001 ,
		_w2754_,
		_w3017_,
		_w3018_,
		_w3019_
	);
	LUT4 #(
		.INIT('h0015)
	) name1270 (
		\u1_u2_tx_dma_en_r_reg/P0001 ,
		_w2766_,
		_w2773_,
		_w3019_,
		_w3020_
	);
	LUT2 #(
		.INIT('h2)
	) name1271 (
		rst_i_pad,
		_w3020_,
		_w3021_
	);
	LUT3 #(
		.INIT('hef)
	) name1272 (
		_w3014_,
		_w3016_,
		_w3021_,
		_w3022_
	);
	LUT4 #(
		.INIT('h0020)
	) name1273 (
		\u1_u1_crc16_reg[2]/P0001 ,
		\u1_u1_send_data_r2_reg/P0001 ,
		\u1_u1_send_data_r_reg/P0001 ,
		\u1_u1_zero_length_r_reg/P0001 ,
		_w3023_
	);
	LUT4 #(
		.INIT('h8000)
	) name1274 (
		\u0_tx_ready_reg/NET0131 ,
		\u1_u1_crc16_reg[2]/P0001 ,
		\u1_u1_state_reg[1]/NET0131 ,
		\u1_u1_tx_valid_r_reg/NET0131 ,
		_w3024_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name1275 (
		_w1805_,
		_w1820_,
		_w3023_,
		_w3024_,
		_w3025_
	);
	LUT4 #(
		.INIT('haa8a)
	) name1276 (
		\u1_u1_crc16_reg[10]/P0001 ,
		\u1_u1_send_data_r2_reg/P0001 ,
		\u1_u1_send_data_r_reg/P0001 ,
		\u1_u1_zero_length_r_reg/P0001 ,
		_w3026_
	);
	LUT2 #(
		.INIT('h1)
	) name1277 (
		_w2098_,
		_w3026_,
		_w3027_
	);
	LUT2 #(
		.INIT('h2)
	) name1278 (
		_w1762_,
		_w2098_,
		_w3028_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name1279 (
		_w1805_,
		_w1820_,
		_w3027_,
		_w3028_,
		_w3029_
	);
	LUT2 #(
		.INIT('hd)
	) name1280 (
		_w3025_,
		_w3029_,
		_w3030_
	);
	LUT4 #(
		.INIT('h0020)
	) name1281 (
		\u1_u1_crc16_reg[3]/P0001 ,
		\u1_u1_send_data_r2_reg/P0001 ,
		\u1_u1_send_data_r_reg/P0001 ,
		\u1_u1_zero_length_r_reg/P0001 ,
		_w3031_
	);
	LUT4 #(
		.INIT('h8000)
	) name1282 (
		\u0_tx_ready_reg/NET0131 ,
		\u1_u1_crc16_reg[3]/P0001 ,
		\u1_u1_state_reg[1]/NET0131 ,
		\u1_u1_tx_valid_r_reg/NET0131 ,
		_w3032_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name1283 (
		_w1805_,
		_w1820_,
		_w3031_,
		_w3032_,
		_w3033_
	);
	LUT4 #(
		.INIT('haa8a)
	) name1284 (
		\u1_u1_crc16_reg[11]/P0001 ,
		\u1_u1_send_data_r2_reg/P0001 ,
		\u1_u1_send_data_r_reg/P0001 ,
		\u1_u1_zero_length_r_reg/P0001 ,
		_w3034_
	);
	LUT4 #(
		.INIT('hdf00)
	) name1285 (
		_w1762_,
		_w1805_,
		_w1820_,
		_w3034_,
		_w3035_
	);
	LUT3 #(
		.INIT('hfb)
	) name1286 (
		_w2098_,
		_w3033_,
		_w3035_,
		_w3036_
	);
	LUT4 #(
		.INIT('h0020)
	) name1287 (
		\u1_u1_crc16_reg[4]/P0001 ,
		\u1_u1_send_data_r2_reg/P0001 ,
		\u1_u1_send_data_r_reg/P0001 ,
		\u1_u1_zero_length_r_reg/P0001 ,
		_w3037_
	);
	LUT4 #(
		.INIT('h8000)
	) name1288 (
		\u0_tx_ready_reg/NET0131 ,
		\u1_u1_crc16_reg[4]/P0001 ,
		\u1_u1_state_reg[1]/NET0131 ,
		\u1_u1_tx_valid_r_reg/NET0131 ,
		_w3038_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name1289 (
		_w1805_,
		_w1820_,
		_w3037_,
		_w3038_,
		_w3039_
	);
	LUT4 #(
		.INIT('haa8a)
	) name1290 (
		\u1_u1_crc16_reg[12]/P0001 ,
		\u1_u1_send_data_r2_reg/P0001 ,
		\u1_u1_send_data_r_reg/P0001 ,
		\u1_u1_zero_length_r_reg/P0001 ,
		_w3040_
	);
	LUT4 #(
		.INIT('hdf00)
	) name1291 (
		_w1762_,
		_w1805_,
		_w1820_,
		_w3040_,
		_w3041_
	);
	LUT3 #(
		.INIT('hfb)
	) name1292 (
		_w2098_,
		_w3039_,
		_w3041_,
		_w3042_
	);
	LUT4 #(
		.INIT('h0020)
	) name1293 (
		\u1_u1_crc16_reg[5]/P0001 ,
		\u1_u1_send_data_r2_reg/P0001 ,
		\u1_u1_send_data_r_reg/P0001 ,
		\u1_u1_zero_length_r_reg/P0001 ,
		_w3043_
	);
	LUT4 #(
		.INIT('h8000)
	) name1294 (
		\u0_tx_ready_reg/NET0131 ,
		\u1_u1_crc16_reg[5]/P0001 ,
		\u1_u1_state_reg[1]/NET0131 ,
		\u1_u1_tx_valid_r_reg/NET0131 ,
		_w3044_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name1295 (
		_w1805_,
		_w1820_,
		_w3043_,
		_w3044_,
		_w3045_
	);
	LUT4 #(
		.INIT('haa8a)
	) name1296 (
		\u1_u1_crc16_reg[13]/P0001 ,
		\u1_u1_send_data_r2_reg/P0001 ,
		\u1_u1_send_data_r_reg/P0001 ,
		\u1_u1_zero_length_r_reg/P0001 ,
		_w3046_
	);
	LUT4 #(
		.INIT('hdf00)
	) name1297 (
		_w1762_,
		_w1805_,
		_w1820_,
		_w3046_,
		_w3047_
	);
	LUT3 #(
		.INIT('hfb)
	) name1298 (
		_w2098_,
		_w3045_,
		_w3047_,
		_w3048_
	);
	LUT4 #(
		.INIT('h0020)
	) name1299 (
		\u1_u1_crc16_reg[6]/P0001 ,
		\u1_u1_send_data_r2_reg/P0001 ,
		\u1_u1_send_data_r_reg/P0001 ,
		\u1_u1_zero_length_r_reg/P0001 ,
		_w3049_
	);
	LUT4 #(
		.INIT('h8000)
	) name1300 (
		\u0_tx_ready_reg/NET0131 ,
		\u1_u1_crc16_reg[6]/P0001 ,
		\u1_u1_state_reg[1]/NET0131 ,
		\u1_u1_tx_valid_r_reg/NET0131 ,
		_w3050_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name1301 (
		_w1805_,
		_w1820_,
		_w3049_,
		_w3050_,
		_w3051_
	);
	LUT4 #(
		.INIT('haa8a)
	) name1302 (
		\u1_u1_crc16_reg[14]/P0001 ,
		\u1_u1_send_data_r2_reg/P0001 ,
		\u1_u1_send_data_r_reg/P0001 ,
		\u1_u1_zero_length_r_reg/P0001 ,
		_w3052_
	);
	LUT4 #(
		.INIT('hdf00)
	) name1303 (
		_w1762_,
		_w1805_,
		_w1820_,
		_w3052_,
		_w3053_
	);
	LUT3 #(
		.INIT('hfb)
	) name1304 (
		_w2098_,
		_w3051_,
		_w3053_,
		_w3054_
	);
	LUT4 #(
		.INIT('h2000)
	) name1305 (
		\u4_csr_reg[15]/NET0131 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		\u4_csr_reg[8]/P0001 ,
		_w3055_
	);
	LUT2 #(
		.INIT('h1)
	) name1306 (
		\u1_u3_adr_r_reg[8]/P0001 ,
		_w3055_,
		_w3056_
	);
	LUT4 #(
		.INIT('ha200)
	) name1307 (
		\u1_u2_sizu_c_reg[8]/NET0131 ,
		\u4_csr_reg[15]/NET0131 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		_w3057_
	);
	LUT4 #(
		.INIT('h0002)
	) name1308 (
		\u1_u2_sizu_c_reg[8]/NET0131 ,
		\u1_u3_in_token_reg/NET0131 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		_w3058_
	);
	LUT3 #(
		.INIT('hf1)
	) name1309 (
		\u1_u3_in_token_reg/NET0131 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		_w3059_
	);
	LUT4 #(
		.INIT('h00c8)
	) name1310 (
		\u1_u3_in_token_reg/NET0131 ,
		\u1_u3_size_next_r_reg[8]/P0001 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		_w3060_
	);
	LUT3 #(
		.INIT('h01)
	) name1311 (
		_w3057_,
		_w3058_,
		_w3060_,
		_w3061_
	);
	LUT4 #(
		.INIT('ha200)
	) name1312 (
		\u1_u2_sizu_c_reg[9]/P0001 ,
		\u4_csr_reg[15]/NET0131 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		_w3062_
	);
	LUT4 #(
		.INIT('h0002)
	) name1313 (
		\u1_u2_sizu_c_reg[9]/P0001 ,
		\u1_u3_in_token_reg/NET0131 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		_w3063_
	);
	LUT2 #(
		.INIT('h1)
	) name1314 (
		_w3062_,
		_w3063_,
		_w3064_
	);
	LUT4 #(
		.INIT('h00c8)
	) name1315 (
		\u1_u3_in_token_reg/NET0131 ,
		\u1_u3_size_next_r_reg[9]/P0001 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		_w3065_
	);
	LUT4 #(
		.INIT('h2000)
	) name1316 (
		\u4_csr_reg[15]/NET0131 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		\u4_csr_reg[9]/NET0131 ,
		_w3066_
	);
	LUT3 #(
		.INIT('h01)
	) name1317 (
		\u1_u3_adr_r_reg[9]/P0001 ,
		_w3065_,
		_w3066_,
		_w3067_
	);
	LUT4 #(
		.INIT('h0777)
	) name1318 (
		_w3056_,
		_w3061_,
		_w3064_,
		_w3067_,
		_w3068_
	);
	LUT4 #(
		.INIT('ha200)
	) name1319 (
		\u1_u2_sizu_c_reg[7]/P0001 ,
		\u4_csr_reg[15]/NET0131 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		_w3069_
	);
	LUT4 #(
		.INIT('h0002)
	) name1320 (
		\u1_u2_sizu_c_reg[7]/P0001 ,
		\u1_u3_in_token_reg/NET0131 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		_w3070_
	);
	LUT2 #(
		.INIT('h1)
	) name1321 (
		_w3069_,
		_w3070_,
		_w3071_
	);
	LUT4 #(
		.INIT('h00c8)
	) name1322 (
		\u1_u3_in_token_reg/NET0131 ,
		\u1_u3_size_next_r_reg[7]/P0001 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		_w3072_
	);
	LUT4 #(
		.INIT('h2000)
	) name1323 (
		\u4_csr_reg[15]/NET0131 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		\u4_csr_reg[7]/P0001 ,
		_w3073_
	);
	LUT3 #(
		.INIT('h01)
	) name1324 (
		\u1_u3_adr_r_reg[7]/P0001 ,
		_w3072_,
		_w3073_,
		_w3074_
	);
	LUT4 #(
		.INIT('ha200)
	) name1325 (
		\u1_u2_sizu_c_reg[6]/P0001 ,
		\u4_csr_reg[15]/NET0131 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		_w3075_
	);
	LUT4 #(
		.INIT('h0002)
	) name1326 (
		\u1_u2_sizu_c_reg[6]/P0001 ,
		\u1_u3_in_token_reg/NET0131 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		_w3076_
	);
	LUT2 #(
		.INIT('h1)
	) name1327 (
		_w3075_,
		_w3076_,
		_w3077_
	);
	LUT4 #(
		.INIT('h00c8)
	) name1328 (
		\u1_u3_in_token_reg/NET0131 ,
		\u1_u3_size_next_r_reg[6]/P0001 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		_w3078_
	);
	LUT4 #(
		.INIT('h2000)
	) name1329 (
		\u4_csr_reg[15]/NET0131 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		\u4_csr_reg[6]/NET0131 ,
		_w3079_
	);
	LUT4 #(
		.INIT('h0001)
	) name1330 (
		_w3075_,
		_w3076_,
		_w3078_,
		_w3079_,
		_w3080_
	);
	LUT2 #(
		.INIT('h2)
	) name1331 (
		\u1_u3_adr_r_reg[6]/P0001 ,
		_w3080_,
		_w3081_
	);
	LUT4 #(
		.INIT('h002a)
	) name1332 (
		\u1_u3_adr_r_reg[6]/P0001 ,
		_w3071_,
		_w3074_,
		_w3080_,
		_w3082_
	);
	LUT4 #(
		.INIT('h0001)
	) name1333 (
		_w3055_,
		_w3057_,
		_w3058_,
		_w3060_,
		_w3083_
	);
	LUT2 #(
		.INIT('h2)
	) name1334 (
		\u1_u3_adr_r_reg[8]/P0001 ,
		_w3083_,
		_w3084_
	);
	LUT4 #(
		.INIT('h0001)
	) name1335 (
		_w3069_,
		_w3070_,
		_w3072_,
		_w3073_,
		_w3085_
	);
	LUT2 #(
		.INIT('h2)
	) name1336 (
		\u1_u3_adr_r_reg[7]/P0001 ,
		_w3085_,
		_w3086_
	);
	LUT4 #(
		.INIT('hf351)
	) name1337 (
		\u1_u3_adr_r_reg[7]/P0001 ,
		\u1_u3_adr_r_reg[8]/P0001 ,
		_w3083_,
		_w3085_,
		_w3087_
	);
	LUT4 #(
		.INIT('h0800)
	) name1338 (
		\u4_csr_reg[10]/P0001 ,
		\u4_csr_reg[15]/NET0131 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		_w3088_
	);
	LUT2 #(
		.INIT('h8)
	) name1339 (
		\u1_u3_adr_r_reg[10]/P0001 ,
		_w3088_,
		_w3089_
	);
	LUT4 #(
		.INIT('h00c8)
	) name1340 (
		\u1_u3_in_token_reg/NET0131 ,
		\u1_u3_size_next_r_reg[10]/P0001 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		_w3090_
	);
	LUT4 #(
		.INIT('haa02)
	) name1341 (
		\u1_u2_sizu_c_reg[10]/P0001 ,
		\u1_u3_in_token_reg/NET0131 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		_w3091_
	);
	LUT2 #(
		.INIT('h1)
	) name1342 (
		_w3090_,
		_w3091_,
		_w3092_
	);
	LUT3 #(
		.INIT('h20)
	) name1343 (
		\u4_csr_reg[15]/NET0131 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		_w3093_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name1344 (
		\u1_u3_adr_r_reg[10]/P0001 ,
		\u4_csr_reg[15]/NET0131 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		_w3094_
	);
	LUT3 #(
		.INIT('he0)
	) name1345 (
		_w3090_,
		_w3091_,
		_w3094_,
		_w3095_
	);
	LUT2 #(
		.INIT('h1)
	) name1346 (
		_w3089_,
		_w3095_,
		_w3096_
	);
	LUT4 #(
		.INIT('h0001)
	) name1347 (
		_w3062_,
		_w3063_,
		_w3065_,
		_w3066_,
		_w3097_
	);
	LUT2 #(
		.INIT('h2)
	) name1348 (
		\u1_u3_adr_r_reg[9]/P0001 ,
		_w3097_,
		_w3098_
	);
	LUT4 #(
		.INIT('h0301)
	) name1349 (
		\u1_u3_adr_r_reg[9]/P0001 ,
		_w3089_,
		_w3095_,
		_w3097_,
		_w3099_
	);
	LUT4 #(
		.INIT('h7500)
	) name1350 (
		_w3068_,
		_w3082_,
		_w3087_,
		_w3099_,
		_w3100_
	);
	LUT3 #(
		.INIT('h0e)
	) name1351 (
		_w3090_,
		_w3091_,
		_w3093_,
		_w3101_
	);
	LUT2 #(
		.INIT('h1)
	) name1352 (
		\u1_u3_adr_r_reg[10]/P0001 ,
		_w3088_,
		_w3102_
	);
	LUT2 #(
		.INIT('h4)
	) name1353 (
		_w3101_,
		_w3102_,
		_w3103_
	);
	LUT2 #(
		.INIT('h1)
	) name1354 (
		_w3100_,
		_w3103_,
		_w3104_
	);
	LUT4 #(
		.INIT('h00c8)
	) name1355 (
		\u1_u3_in_token_reg/NET0131 ,
		\u1_u3_size_next_r_reg[5]/P0001 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		_w3105_
	);
	LUT4 #(
		.INIT('haa02)
	) name1356 (
		\u1_u2_sizu_c_reg[5]/P0001 ,
		\u1_u3_in_token_reg/NET0131 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		_w3106_
	);
	LUT3 #(
		.INIT('h54)
	) name1357 (
		_w3093_,
		_w3105_,
		_w3106_,
		_w3107_
	);
	LUT4 #(
		.INIT('h2000)
	) name1358 (
		\u4_csr_reg[15]/NET0131 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		\u4_csr_reg[5]/NET0131 ,
		_w3108_
	);
	LUT2 #(
		.INIT('h1)
	) name1359 (
		\u1_u3_adr_r_reg[5]/P0001 ,
		_w3108_,
		_w3109_
	);
	LUT4 #(
		.INIT('haa02)
	) name1360 (
		\u1_u2_sizu_c_reg[4]/P0001 ,
		\u1_u3_in_token_reg/NET0131 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		_w3110_
	);
	LUT4 #(
		.INIT('h00c8)
	) name1361 (
		\u1_u3_in_token_reg/NET0131 ,
		\u1_u3_size_next_r_reg[4]/P0001 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		_w3111_
	);
	LUT3 #(
		.INIT('h54)
	) name1362 (
		_w3093_,
		_w3110_,
		_w3111_,
		_w3112_
	);
	LUT4 #(
		.INIT('h2000)
	) name1363 (
		\u4_csr_reg[15]/NET0131 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		\u4_csr_reg[4]/NET0131 ,
		_w3113_
	);
	LUT2 #(
		.INIT('h1)
	) name1364 (
		\u1_u3_adr_r_reg[4]/P0001 ,
		_w3113_,
		_w3114_
	);
	LUT2 #(
		.INIT('h4)
	) name1365 (
		_w3112_,
		_w3114_,
		_w3115_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name1366 (
		_w3107_,
		_w3109_,
		_w3112_,
		_w3114_,
		_w3116_
	);
	LUT4 #(
		.INIT('h2000)
	) name1367 (
		\u4_csr_reg[15]/NET0131 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		\u4_csr_reg[3]/P0001 ,
		_w3117_
	);
	LUT2 #(
		.INIT('h8)
	) name1368 (
		\u1_u3_adr_r_reg[3]/P0001 ,
		_w3117_,
		_w3118_
	);
	LUT4 #(
		.INIT('h00c8)
	) name1369 (
		\u1_u3_in_token_reg/NET0131 ,
		\u1_u3_size_next_r_reg[3]/P0001 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		_w3119_
	);
	LUT4 #(
		.INIT('haa02)
	) name1370 (
		\u1_u2_sizu_c_reg[3]/P0001 ,
		\u1_u3_in_token_reg/NET0131 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		_w3120_
	);
	LUT2 #(
		.INIT('h1)
	) name1371 (
		_w3119_,
		_w3120_,
		_w3121_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name1372 (
		\u1_u3_adr_r_reg[3]/P0001 ,
		\u4_csr_reg[15]/NET0131 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		_w3122_
	);
	LUT3 #(
		.INIT('he0)
	) name1373 (
		_w3119_,
		_w3120_,
		_w3122_,
		_w3123_
	);
	LUT2 #(
		.INIT('h1)
	) name1374 (
		_w3118_,
		_w3123_,
		_w3124_
	);
	LUT3 #(
		.INIT('h54)
	) name1375 (
		_w3093_,
		_w3119_,
		_w3120_,
		_w3125_
	);
	LUT2 #(
		.INIT('h1)
	) name1376 (
		\u1_u3_adr_r_reg[3]/P0001 ,
		_w3117_,
		_w3126_
	);
	LUT4 #(
		.INIT('h2000)
	) name1377 (
		\u4_csr_reg[15]/NET0131 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		\u4_csr_reg[2]/NET0131 ,
		_w3127_
	);
	LUT2 #(
		.INIT('h8)
	) name1378 (
		\u1_u3_adr_r_reg[2]/P0001 ,
		_w3127_,
		_w3128_
	);
	LUT4 #(
		.INIT('h00c8)
	) name1379 (
		\u1_u3_in_token_reg/NET0131 ,
		\u1_u3_size_next_r_reg[2]/P0001 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		_w3129_
	);
	LUT4 #(
		.INIT('haa02)
	) name1380 (
		\u1_u2_sizu_c_reg[2]/P0001 ,
		\u1_u3_in_token_reg/NET0131 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		_w3130_
	);
	LUT2 #(
		.INIT('h1)
	) name1381 (
		_w3129_,
		_w3130_,
		_w3131_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name1382 (
		\u1_u3_adr_r_reg[2]/P0001 ,
		\u4_csr_reg[15]/NET0131 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		_w3132_
	);
	LUT3 #(
		.INIT('he0)
	) name1383 (
		_w3129_,
		_w3130_,
		_w3132_,
		_w3133_
	);
	LUT4 #(
		.INIT('hbbb0)
	) name1384 (
		_w3125_,
		_w3126_,
		_w3128_,
		_w3133_,
		_w3134_
	);
	LUT2 #(
		.INIT('h2)
	) name1385 (
		_w3124_,
		_w3134_,
		_w3135_
	);
	LUT3 #(
		.INIT('ha2)
	) name1386 (
		_w3116_,
		_w3124_,
		_w3134_,
		_w3136_
	);
	LUT4 #(
		.INIT('h0800)
	) name1387 (
		\u4_csr_reg[15]/NET0131 ,
		\u4_csr_reg[1]/P0001 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		_w3137_
	);
	LUT2 #(
		.INIT('h8)
	) name1388 (
		\u1_u3_adr_r_reg[1]/P0001 ,
		_w3137_,
		_w3138_
	);
	LUT4 #(
		.INIT('h00c8)
	) name1389 (
		\u1_u3_in_token_reg/NET0131 ,
		\u1_u3_size_next_r_reg[1]/P0001 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		_w3139_
	);
	LUT4 #(
		.INIT('haa02)
	) name1390 (
		\u1_u2_sizu_c_reg[1]/P0001 ,
		\u1_u3_in_token_reg/NET0131 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		_w3140_
	);
	LUT2 #(
		.INIT('h1)
	) name1391 (
		_w3139_,
		_w3140_,
		_w3141_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name1392 (
		\u1_u3_adr_r_reg[1]/P0001 ,
		\u4_csr_reg[15]/NET0131 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		_w3142_
	);
	LUT3 #(
		.INIT('he0)
	) name1393 (
		_w3139_,
		_w3140_,
		_w3142_,
		_w3143_
	);
	LUT2 #(
		.INIT('h1)
	) name1394 (
		_w3138_,
		_w3143_,
		_w3144_
	);
	LUT3 #(
		.INIT('h54)
	) name1395 (
		_w3093_,
		_w3139_,
		_w3140_,
		_w3145_
	);
	LUT2 #(
		.INIT('h1)
	) name1396 (
		\u1_u3_adr_r_reg[1]/P0001 ,
		_w3137_,
		_w3146_
	);
	LUT4 #(
		.INIT('h0800)
	) name1397 (
		\u4_csr_reg[0]/P0001 ,
		\u4_csr_reg[15]/NET0131 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		_w3147_
	);
	LUT2 #(
		.INIT('h8)
	) name1398 (
		\u1_u3_adr_r_reg[0]/P0001 ,
		_w3147_,
		_w3148_
	);
	LUT4 #(
		.INIT('h00c8)
	) name1399 (
		\u1_u3_in_token_reg/NET0131 ,
		\u1_u3_size_next_r_reg[0]/P0001 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		_w3149_
	);
	LUT4 #(
		.INIT('haa02)
	) name1400 (
		\u1_u2_sizu_c_reg[0]/P0001 ,
		\u1_u3_in_token_reg/NET0131 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		_w3150_
	);
	LUT2 #(
		.INIT('h1)
	) name1401 (
		_w3149_,
		_w3150_,
		_w3151_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name1402 (
		\u1_u3_adr_r_reg[0]/P0001 ,
		\u4_csr_reg[15]/NET0131 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		_w3152_
	);
	LUT3 #(
		.INIT('he0)
	) name1403 (
		_w3149_,
		_w3150_,
		_w3152_,
		_w3153_
	);
	LUT4 #(
		.INIT('hbbb0)
	) name1404 (
		_w3145_,
		_w3146_,
		_w3148_,
		_w3153_,
		_w3154_
	);
	LUT3 #(
		.INIT('h54)
	) name1405 (
		_w3093_,
		_w3129_,
		_w3130_,
		_w3155_
	);
	LUT2 #(
		.INIT('h1)
	) name1406 (
		\u1_u3_adr_r_reg[2]/P0001 ,
		_w3127_,
		_w3156_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name1407 (
		_w3125_,
		_w3126_,
		_w3155_,
		_w3156_,
		_w3157_
	);
	LUT4 #(
		.INIT('ha200)
	) name1408 (
		_w3116_,
		_w3144_,
		_w3154_,
		_w3157_,
		_w3158_
	);
	LUT4 #(
		.INIT('h0020)
	) name1409 (
		\u4_csr_reg[15]/NET0131 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		\u4_csr_reg[5]/NET0131 ,
		_w3159_
	);
	LUT4 #(
		.INIT('h00fe)
	) name1410 (
		_w3105_,
		_w3106_,
		_w3108_,
		_w3159_,
		_w3160_
	);
	LUT2 #(
		.INIT('h8)
	) name1411 (
		\u1_u3_adr_r_reg[5]/P0001 ,
		_w3160_,
		_w3161_
	);
	LUT4 #(
		.INIT('h0020)
	) name1412 (
		\u4_csr_reg[15]/NET0131 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		\u4_csr_reg[4]/NET0131 ,
		_w3162_
	);
	LUT4 #(
		.INIT('h00fe)
	) name1413 (
		_w3110_,
		_w3111_,
		_w3113_,
		_w3162_,
		_w3163_
	);
	LUT4 #(
		.INIT('h8a00)
	) name1414 (
		\u1_u3_adr_r_reg[4]/P0001 ,
		_w3107_,
		_w3109_,
		_w3163_,
		_w3164_
	);
	LUT2 #(
		.INIT('h1)
	) name1415 (
		_w3161_,
		_w3164_,
		_w3165_
	);
	LUT3 #(
		.INIT('h01)
	) name1416 (
		\u1_u3_adr_r_reg[6]/P0001 ,
		_w3078_,
		_w3079_,
		_w3166_
	);
	LUT2 #(
		.INIT('h8)
	) name1417 (
		_w3077_,
		_w3166_,
		_w3167_
	);
	LUT4 #(
		.INIT('h0777)
	) name1418 (
		_w3071_,
		_w3074_,
		_w3077_,
		_w3166_,
		_w3168_
	);
	LUT2 #(
		.INIT('h8)
	) name1419 (
		_w3068_,
		_w3168_,
		_w3169_
	);
	LUT3 #(
		.INIT('h20)
	) name1420 (
		_w3068_,
		_w3103_,
		_w3168_,
		_w3170_
	);
	LUT4 #(
		.INIT('hef00)
	) name1421 (
		_w3136_,
		_w3158_,
		_w3165_,
		_w3170_,
		_w3171_
	);
	LUT2 #(
		.INIT('h8)
	) name1422 (
		\u1_u3_adr_r_reg[11]/P0001 ,
		\u1_u3_adr_r_reg[12]/P0001 ,
		_w3172_
	);
	LUT3 #(
		.INIT('h80)
	) name1423 (
		\u1_u3_adr_r_reg[11]/P0001 ,
		\u1_u3_adr_r_reg[12]/P0001 ,
		\u1_u3_adr_r_reg[13]/P0001 ,
		_w3173_
	);
	LUT2 #(
		.INIT('h1)
	) name1424 (
		\u1_u3_adr_r_reg[14]/P0001 ,
		\u1_u3_out_to_small_r_reg/P0001 ,
		_w3174_
	);
	LUT2 #(
		.INIT('h8)
	) name1425 (
		_w3173_,
		_w3174_,
		_w3175_
	);
	LUT3 #(
		.INIT('he0)
	) name1426 (
		_w3104_,
		_w3171_,
		_w3175_,
		_w3176_
	);
	LUT2 #(
		.INIT('h8)
	) name1427 (
		\u1_u3_out_to_small_r_reg/P0001 ,
		\u4_buf0_reg[14]/P0001 ,
		_w3177_
	);
	LUT3 #(
		.INIT('h1d)
	) name1428 (
		\u1_u3_adr_r_reg[14]/P0001 ,
		\u1_u3_out_to_small_r_reg/P0001 ,
		\u4_buf0_reg[14]/P0001 ,
		_w3178_
	);
	LUT2 #(
		.INIT('h2)
	) name1429 (
		_w3173_,
		_w3177_,
		_w3179_
	);
	LUT4 #(
		.INIT('h010f)
	) name1430 (
		_w3104_,
		_w3171_,
		_w3178_,
		_w3179_,
		_w3180_
	);
	LUT2 #(
		.INIT('he)
	) name1431 (
		_w3176_,
		_w3180_,
		_w3181_
	);
	LUT2 #(
		.INIT('h8)
	) name1432 (
		\u1_u2_adr_cb_reg[0]/NET0131 ,
		\u1_u2_adr_cb_reg[1]/NET0131 ,
		_w3182_
	);
	LUT3 #(
		.INIT('h78)
	) name1433 (
		\u1_u2_adr_cb_reg[0]/NET0131 ,
		\u1_u2_adr_cb_reg[1]/NET0131 ,
		\u1_u2_adr_cb_reg[2]/NET0131 ,
		_w3183_
	);
	LUT2 #(
		.INIT('h1)
	) name1434 (
		_w1765_,
		_w3183_,
		_w3184_
	);
	LUT2 #(
		.INIT('h1)
	) name1435 (
		\u1_u2_rx_dma_en_r_reg/P0001 ,
		\u1_u2_tx_dma_en_r_reg/P0001 ,
		_w3185_
	);
	LUT2 #(
		.INIT('h1)
	) name1436 (
		\u1_u2_adr_cb_reg[2]/NET0131 ,
		\u1_u2_rx_data_valid_r_reg/NET0131 ,
		_w3186_
	);
	LUT3 #(
		.INIT('h8c)
	) name1437 (
		_w1762_,
		_w3185_,
		_w3186_,
		_w3187_
	);
	LUT3 #(
		.INIT('he0)
	) name1438 (
		\u1_u2_rx_dma_en_r_reg/P0001 ,
		\u1_u2_tx_dma_en_r_reg/P0001 ,
		\u1_u3_adr_reg[2]/P0001 ,
		_w3188_
	);
	LUT4 #(
		.INIT('haa20)
	) name1439 (
		rst_i_pad,
		_w3184_,
		_w3187_,
		_w3188_,
		_w3189_
	);
	LUT3 #(
		.INIT('h40)
	) name1440 (
		_w1762_,
		_w1768_,
		_w3185_,
		_w3190_
	);
	LUT2 #(
		.INIT('h4)
	) name1441 (
		\u1_u2_adr_cb_reg[0]/NET0131 ,
		\u1_u2_adr_cb_reg[1]/NET0131 ,
		_w3191_
	);
	LUT4 #(
		.INIT('h0009)
	) name1442 (
		\u1_u2_adr_cb_reg[0]/NET0131 ,
		\u1_u2_adr_cb_reg[1]/NET0131 ,
		\u1_u2_rx_dma_en_r_reg/P0001 ,
		\u1_u2_tx_dma_en_r_reg/P0001 ,
		_w3192_
	);
	LUT2 #(
		.INIT('h4)
	) name1443 (
		_w1765_,
		_w3192_,
		_w3193_
	);
	LUT4 #(
		.INIT('haa02)
	) name1444 (
		rst_i_pad,
		\u1_u2_rx_dma_en_r_reg/P0001 ,
		\u1_u2_tx_dma_en_r_reg/P0001 ,
		\u1_u3_adr_reg[1]/P0001 ,
		_w3194_
	);
	LUT3 #(
		.INIT('h10)
	) name1445 (
		_w3190_,
		_w3193_,
		_w3194_,
		_w3195_
	);
	LUT4 #(
		.INIT('h363c)
	) name1446 (
		\u1_u1_state_reg[1]/NET0131 ,
		\u1_u2_adr_cb_reg[0]/NET0131 ,
		\u1_u2_rx_data_valid_r_reg/NET0131 ,
		_w1761_,
		_w3196_
	);
	LUT4 #(
		.INIT('haa02)
	) name1447 (
		rst_i_pad,
		\u1_u2_rx_dma_en_r_reg/P0001 ,
		\u1_u2_tx_dma_en_r_reg/P0001 ,
		\u1_u3_adr_reg[0]/P0001 ,
		_w3197_
	);
	LUT3 #(
		.INIT('hd0)
	) name1448 (
		_w3185_,
		_w3196_,
		_w3197_,
		_w3198_
	);
	LUT4 #(
		.INIT('h7f00)
	) name1449 (
		\u0_tx_ready_reg/NET0131 ,
		\u1_u1_state_reg[1]/NET0131 ,
		\u1_u1_tx_valid_r_reg/NET0131 ,
		\u1_u2_sizd_c_reg[0]/P0001 ,
		_w3199_
	);
	LUT2 #(
		.INIT('h1)
	) name1450 (
		_w2747_,
		_w3199_,
		_w3200_
	);
	LUT4 #(
		.INIT('ha8a0)
	) name1451 (
		rst_i_pad,
		\u1_u2_mack_r_reg/P0001 ,
		\u1_u2_send_data_r_reg/NET0131 ,
		\u1_u2_state_reg[5]/NET0131 ,
		_w3201_
	);
	LUT3 #(
		.INIT('h70)
	) name1452 (
		_w2757_,
		_w3200_,
		_w3201_,
		_w3202_
	);
	LUT2 #(
		.INIT('h1)
	) name1453 (
		\u1_u2_mack_r_reg/P0001 ,
		\u1_u2_state_reg[0]/P0001 ,
		_w3203_
	);
	LUT2 #(
		.INIT('h1)
	) name1454 (
		\u1_u2_state_reg[0]/P0001 ,
		\u1_u2_state_reg[1]/NET0131 ,
		_w3204_
	);
	LUT4 #(
		.INIT('h0001)
	) name1455 (
		\u1_u2_state_reg[0]/P0001 ,
		\u1_u2_state_reg[1]/NET0131 ,
		\u1_u2_state_reg[2]/NET0131 ,
		\u1_u2_state_reg[3]/NET0131 ,
		_w3205_
	);
	LUT4 #(
		.INIT('h0002)
	) name1456 (
		\u1_u2_state_reg[4]/NET0131 ,
		\u1_u2_state_reg[5]/NET0131 ,
		\u1_u2_state_reg[6]/NET0131 ,
		\u1_u2_state_reg[7]/NET0131 ,
		_w3206_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name1457 (
		rst_i_pad,
		_w3203_,
		_w3205_,
		_w3206_,
		_w3207_
	);
	LUT2 #(
		.INIT('h1)
	) name1458 (
		\u1_u2_state_reg[4]/NET0131 ,
		\u1_u2_state_reg[6]/NET0131 ,
		_w3208_
	);
	LUT4 #(
		.INIT('h0001)
	) name1459 (
		\u1_u2_state_reg[4]/NET0131 ,
		\u1_u2_state_reg[5]/NET0131 ,
		\u1_u2_state_reg[6]/NET0131 ,
		\u1_u2_state_reg[7]/NET0131 ,
		_w3209_
	);
	LUT3 #(
		.INIT('h0b)
	) name1460 (
		\u1_u2_rx_data_done_r2_reg/P0001 ,
		\u1_u2_state_reg[0]/P0001 ,
		\u1_u3_abort_reg/P0001 ,
		_w3210_
	);
	LUT2 #(
		.INIT('h2)
	) name1461 (
		\u1_u2_state_reg[2]/NET0131 ,
		\u1_u2_state_reg[3]/NET0131 ,
		_w3211_
	);
	LUT4 #(
		.INIT('h0800)
	) name1462 (
		_w3204_,
		_w3209_,
		_w3210_,
		_w3211_,
		_w3212_
	);
	LUT4 #(
		.INIT('h00f1)
	) name1463 (
		\u1_u2_state_reg[0]/P0001 ,
		\u1_u2_wr_done_reg/P0001 ,
		\u1_u2_wr_last_reg/P0001 ,
		\u1_u3_abort_reg/P0001 ,
		_w3213_
	);
	LUT4 #(
		.INIT('h0100)
	) name1464 (
		\u1_u2_state_reg[0]/P0001 ,
		\u1_u2_state_reg[1]/NET0131 ,
		\u1_u2_state_reg[2]/NET0131 ,
		\u1_u2_state_reg[3]/NET0131 ,
		_w3214_
	);
	LUT3 #(
		.INIT('h20)
	) name1465 (
		_w3209_,
		_w3213_,
		_w3214_,
		_w3215_
	);
	LUT4 #(
		.INIT('h0002)
	) name1466 (
		\u1_u2_state_reg[0]/P0001 ,
		\u1_u2_state_reg[1]/NET0131 ,
		\u1_u2_state_reg[2]/NET0131 ,
		\u1_u2_state_reg[3]/NET0131 ,
		_w3216_
	);
	LUT3 #(
		.INIT('h04)
	) name1467 (
		\u1_u1_send_zero_length_r_reg/P0001 ,
		\u1_u2_tx_dma_en_r_reg/P0001 ,
		\u1_u3_abort_reg/P0001 ,
		_w3217_
	);
	LUT4 #(
		.INIT('hff23)
	) name1468 (
		\u1_u1_send_zero_length_r_reg/P0001 ,
		\u1_u2_rx_dma_en_r_reg/P0001 ,
		\u1_u2_tx_dma_en_r_reg/P0001 ,
		\u1_u3_abort_reg/P0001 ,
		_w3218_
	);
	LUT3 #(
		.INIT('h80)
	) name1469 (
		_w3209_,
		_w3216_,
		_w3218_,
		_w3219_
	);
	LUT4 #(
		.INIT('h0002)
	) name1470 (
		_w3207_,
		_w3212_,
		_w3215_,
		_w3219_,
		_w3220_
	);
	LUT3 #(
		.INIT('h0b)
	) name1471 (
		\u1_u2_mack_r_reg/P0001 ,
		\u1_u2_state_reg[0]/P0001 ,
		\u1_u3_abort_reg/P0001 ,
		_w3221_
	);
	LUT4 #(
		.INIT('h0004)
	) name1472 (
		\u1_u2_state_reg[4]/NET0131 ,
		\u1_u2_state_reg[5]/NET0131 ,
		\u1_u2_state_reg[6]/NET0131 ,
		\u1_u2_state_reg[7]/NET0131 ,
		_w3222_
	);
	LUT4 #(
		.INIT('h0010)
	) name1473 (
		\u1_u2_state_reg[4]/NET0131 ,
		\u1_u2_state_reg[5]/NET0131 ,
		\u1_u2_state_reg[6]/NET0131 ,
		\u1_u2_state_reg[7]/NET0131 ,
		_w3223_
	);
	LUT3 #(
		.INIT('h57)
	) name1474 (
		_w3205_,
		_w3222_,
		_w3223_,
		_w3224_
	);
	LUT4 #(
		.INIT('h0004)
	) name1475 (
		\u1_u2_state_reg[0]/P0001 ,
		\u1_u2_state_reg[1]/NET0131 ,
		\u1_u2_state_reg[2]/NET0131 ,
		\u1_u2_state_reg[3]/NET0131 ,
		_w3225_
	);
	LUT2 #(
		.INIT('h8)
	) name1476 (
		_w3209_,
		_w3225_,
		_w3226_
	);
	LUT3 #(
		.INIT('h51)
	) name1477 (
		_w3221_,
		_w3224_,
		_w3226_,
		_w3227_
	);
	LUT2 #(
		.INIT('h1)
	) name1478 (
		\u1_u2_sizd_is_zero_reg/P0001 ,
		\u1_u3_abort_reg/P0001 ,
		_w3228_
	);
	LUT3 #(
		.INIT('h01)
	) name1479 (
		\u1_u2_sizd_is_zero_reg/P0001 ,
		\u1_u2_state_reg[0]/P0001 ,
		\u1_u3_abort_reg/P0001 ,
		_w3229_
	);
	LUT4 #(
		.INIT('h0008)
	) name1480 (
		\u1_u2_adr_cb_reg[0]/NET0131 ,
		\u1_u2_adr_cb_reg[1]/NET0131 ,
		\u1_u2_sizd_is_zero_reg/P0001 ,
		\u1_u3_abort_reg/P0001 ,
		_w3230_
	);
	LUT3 #(
		.INIT('h13)
	) name1481 (
		_w1762_,
		_w3229_,
		_w3230_,
		_w3231_
	);
	LUT2 #(
		.INIT('h4)
	) name1482 (
		\u1_u2_state_reg[5]/NET0131 ,
		\u1_u2_state_reg[7]/NET0131 ,
		_w3232_
	);
	LUT3 #(
		.INIT('h80)
	) name1483 (
		_w3205_,
		_w3208_,
		_w3232_,
		_w3233_
	);
	LUT2 #(
		.INIT('h8)
	) name1484 (
		_w3231_,
		_w3233_,
		_w3234_
	);
	LUT3 #(
		.INIT('hfd)
	) name1485 (
		_w3220_,
		_w3227_,
		_w3234_,
		_w3235_
	);
	LUT4 #(
		.INIT('hef00)
	) name1486 (
		_w3136_,
		_w3158_,
		_w3165_,
		_w3169_,
		_w3236_
	);
	LUT4 #(
		.INIT('h0075)
	) name1487 (
		_w3068_,
		_w3082_,
		_w3087_,
		_w3098_,
		_w3237_
	);
	LUT3 #(
		.INIT('h13)
	) name1488 (
		\u1_u3_adr_r_reg[10]/P0001 ,
		\u1_u3_out_to_small_r_reg/P0001 ,
		_w3088_,
		_w3238_
	);
	LUT4 #(
		.INIT('h4500)
	) name1489 (
		_w3095_,
		_w3101_,
		_w3102_,
		_w3238_,
		_w3239_
	);
	LUT2 #(
		.INIT('h8)
	) name1490 (
		_w3237_,
		_w3239_,
		_w3240_
	);
	LUT2 #(
		.INIT('h4)
	) name1491 (
		_w3236_,
		_w3240_,
		_w3241_
	);
	LUT4 #(
		.INIT('h6665)
	) name1492 (
		\u1_u3_adr_r_reg[10]/P0001 ,
		_w3088_,
		_w3092_,
		_w3093_,
		_w3242_
	);
	LUT2 #(
		.INIT('h1)
	) name1493 (
		\u1_u3_out_to_small_r_reg/P0001 ,
		_w3242_,
		_w3243_
	);
	LUT2 #(
		.INIT('h4)
	) name1494 (
		_w3237_,
		_w3243_,
		_w3244_
	);
	LUT4 #(
		.INIT('h0040)
	) name1495 (
		\u1_u3_out_to_small_r_reg/P0001 ,
		_w3068_,
		_w3168_,
		_w3242_,
		_w3245_
	);
	LUT4 #(
		.INIT('hef00)
	) name1496 (
		_w3136_,
		_w3158_,
		_w3165_,
		_w3245_,
		_w3246_
	);
	LUT2 #(
		.INIT('h8)
	) name1497 (
		\u1_u3_out_to_small_r_reg/P0001 ,
		\u4_buf0_reg[10]/P0001 ,
		_w3247_
	);
	LUT3 #(
		.INIT('h01)
	) name1498 (
		_w3244_,
		_w3246_,
		_w3247_,
		_w3248_
	);
	LUT2 #(
		.INIT('hb)
	) name1499 (
		_w3241_,
		_w3248_,
		_w3249_
	);
	LUT4 #(
		.INIT('hf531)
	) name1500 (
		\u1_u3_adr_r_reg[8]/P0001 ,
		\u1_u3_adr_r_reg[9]/P0001 ,
		_w3083_,
		_w3097_,
		_w3250_
	);
	LUT4 #(
		.INIT('h7077)
	) name1501 (
		_w3064_,
		_w3067_,
		_w3101_,
		_w3102_,
		_w3251_
	);
	LUT2 #(
		.INIT('h2)
	) name1502 (
		\u1_u3_adr_r_reg[11]/P0001 ,
		\u1_u3_adr_r_reg[12]/P0001 ,
		_w3252_
	);
	LUT4 #(
		.INIT('h7500)
	) name1503 (
		_w3096_,
		_w3250_,
		_w3251_,
		_w3252_,
		_w3253_
	);
	LUT4 #(
		.INIT('h0001)
	) name1504 (
		_w3082_,
		_w3086_,
		_w3161_,
		_w3164_,
		_w3254_
	);
	LUT3 #(
		.INIT('h10)
	) name1505 (
		_w3136_,
		_w3158_,
		_w3254_,
		_w3255_
	);
	LUT3 #(
		.INIT('h01)
	) name1506 (
		_w3082_,
		_w3086_,
		_w3168_,
		_w3256_
	);
	LUT3 #(
		.INIT('h20)
	) name1507 (
		_w3068_,
		_w3103_,
		_w3252_,
		_w3257_
	);
	LUT2 #(
		.INIT('h4)
	) name1508 (
		_w3256_,
		_w3257_,
		_w3258_
	);
	LUT3 #(
		.INIT('h45)
	) name1509 (
		_w3253_,
		_w3255_,
		_w3258_,
		_w3259_
	);
	LUT3 #(
		.INIT('h08)
	) name1510 (
		\u1_u3_adr_r_reg[11]/P0001 ,
		_w3068_,
		_w3103_,
		_w3260_
	);
	LUT2 #(
		.INIT('h4)
	) name1511 (
		_w3256_,
		_w3260_,
		_w3261_
	);
	LUT2 #(
		.INIT('h4)
	) name1512 (
		\u1_u3_adr_r_reg[11]/P0001 ,
		\u1_u3_adr_r_reg[12]/P0001 ,
		_w3262_
	);
	LUT3 #(
		.INIT('h02)
	) name1513 (
		\u1_u3_adr_r_reg[12]/P0001 ,
		_w3089_,
		_w3095_,
		_w3263_
	);
	LUT4 #(
		.INIT('h040f)
	) name1514 (
		_w3250_,
		_w3251_,
		_w3262_,
		_w3263_,
		_w3264_
	);
	LUT3 #(
		.INIT('h0b)
	) name1515 (
		_w3255_,
		_w3261_,
		_w3264_,
		_w3265_
	);
	LUT4 #(
		.INIT('hdd8d)
	) name1516 (
		\u1_u3_out_to_small_r_reg/P0001 ,
		\u4_buf0_reg[12]/P0001 ,
		_w3259_,
		_w3265_,
		_w3266_
	);
	LUT4 #(
		.INIT('h8000)
	) name1517 (
		\u1_u3_adr_r_reg[12]/P0001 ,
		\u1_u3_adr_r_reg[13]/P0001 ,
		\u1_u3_adr_r_reg[14]/P0001 ,
		\u1_u3_adr_r_reg[15]/P0001 ,
		_w3267_
	);
	LUT2 #(
		.INIT('h2)
	) name1518 (
		\u1_u3_adr_r_reg[16]/P0001 ,
		\u1_u3_out_to_small_r_reg/P0001 ,
		_w3268_
	);
	LUT2 #(
		.INIT('h4)
	) name1519 (
		_w3267_,
		_w3268_,
		_w3269_
	);
	LUT4 #(
		.INIT('h2a22)
	) name1520 (
		\u1_u3_adr_r_reg[11]/P0001 ,
		_w3096_,
		_w3250_,
		_w3251_,
		_w3270_
	);
	LUT2 #(
		.INIT('h2)
	) name1521 (
		_w3268_,
		_w3270_,
		_w3271_
	);
	LUT4 #(
		.INIT('h040f)
	) name1522 (
		_w3255_,
		_w3261_,
		_w3269_,
		_w3271_,
		_w3272_
	);
	LUT2 #(
		.INIT('h1)
	) name1523 (
		\u1_u3_adr_r_reg[16]/P0001 ,
		\u1_u3_out_to_small_r_reg/P0001 ,
		_w3273_
	);
	LUT2 #(
		.INIT('h8)
	) name1524 (
		_w3267_,
		_w3273_,
		_w3274_
	);
	LUT4 #(
		.INIT('hf400)
	) name1525 (
		_w3255_,
		_w3261_,
		_w3270_,
		_w3274_,
		_w3275_
	);
	LUT2 #(
		.INIT('h8)
	) name1526 (
		\u1_u3_out_to_small_r_reg/P0001 ,
		\u4_buf0_reg[16]/P0001 ,
		_w3276_
	);
	LUT3 #(
		.INIT('hfd)
	) name1527 (
		_w3272_,
		_w3275_,
		_w3276_,
		_w3277_
	);
	LUT3 #(
		.INIT('h15)
	) name1528 (
		\u1_u2_state_reg[6]/NET0131 ,
		_w1762_,
		_w3182_,
		_w3278_
	);
	LUT4 #(
		.INIT('h0100)
	) name1529 (
		\u1_u2_state_reg[4]/NET0131 ,
		\u1_u2_state_reg[5]/NET0131 ,
		\u1_u2_state_reg[6]/NET0131 ,
		\u1_u2_state_reg[7]/NET0131 ,
		_w3279_
	);
	LUT3 #(
		.INIT('h80)
	) name1530 (
		_w3205_,
		_w3228_,
		_w3279_,
		_w3280_
	);
	LUT3 #(
		.INIT('h0e)
	) name1531 (
		\u1_u2_mack_r_reg/P0001 ,
		\u1_u2_state_reg[6]/NET0131 ,
		\u1_u3_abort_reg/P0001 ,
		_w3281_
	);
	LUT3 #(
		.INIT('h80)
	) name1532 (
		_w3205_,
		_w3222_,
		_w3281_,
		_w3282_
	);
	LUT2 #(
		.INIT('h1)
	) name1533 (
		\u1_u2_mack_r_reg/P0001 ,
		\u1_u3_abort_reg/P0001 ,
		_w3283_
	);
	LUT3 #(
		.INIT('h80)
	) name1534 (
		_w3205_,
		_w3223_,
		_w3283_,
		_w3284_
	);
	LUT4 #(
		.INIT('h000b)
	) name1535 (
		_w3278_,
		_w3280_,
		_w3282_,
		_w3284_,
		_w3285_
	);
	LUT2 #(
		.INIT('h2)
	) name1536 (
		rst_i_pad,
		_w3285_,
		_w3286_
	);
	LUT4 #(
		.INIT('h00a8)
	) name1537 (
		rst_i_pad,
		\u1_u2_mack_r_reg/P0001 ,
		\u1_u2_state_reg[7]/NET0131 ,
		\u1_u3_abort_reg/P0001 ,
		_w3287_
	);
	LUT3 #(
		.INIT('h80)
	) name1538 (
		_w3205_,
		_w3223_,
		_w3287_,
		_w3288_
	);
	LUT3 #(
		.INIT('h2a)
	) name1539 (
		rst_i_pad,
		_w1762_,
		_w3182_,
		_w3289_
	);
	LUT3 #(
		.INIT('hec)
	) name1540 (
		_w3280_,
		_w3288_,
		_w3289_,
		_w3290_
	);
	LUT4 #(
		.INIT('h0001)
	) name1541 (
		_w3128_,
		_w3133_,
		_w3138_,
		_w3143_,
		_w3291_
	);
	LUT3 #(
		.INIT('h8c)
	) name1542 (
		_w3154_,
		_w3157_,
		_w3291_,
		_w3292_
	);
	LUT4 #(
		.INIT('h0103)
	) name1543 (
		\u1_u3_adr_r_reg[4]/P0001 ,
		_w3118_,
		_w3123_,
		_w3163_,
		_w3293_
	);
	LUT4 #(
		.INIT('h7300)
	) name1544 (
		_w3154_,
		_w3157_,
		_w3291_,
		_w3293_,
		_w3294_
	);
	LUT4 #(
		.INIT('h0777)
	) name1545 (
		_w3056_,
		_w3061_,
		_w3071_,
		_w3074_,
		_w3295_
	);
	LUT3 #(
		.INIT('h20)
	) name1546 (
		_w3116_,
		_w3167_,
		_w3295_,
		_w3296_
	);
	LUT2 #(
		.INIT('h4)
	) name1547 (
		_w3294_,
		_w3296_,
		_w3297_
	);
	LUT4 #(
		.INIT('h20a0)
	) name1548 (
		\u1_u3_adr_r_reg[5]/P0001 ,
		_w3077_,
		_w3160_,
		_w3166_,
		_w3298_
	);
	LUT3 #(
		.INIT('hc8)
	) name1549 (
		_w3081_,
		_w3295_,
		_w3298_,
		_w3299_
	);
	LUT4 #(
		.INIT('h2022)
	) name1550 (
		\u1_u3_adr_r_reg[9]/P0001 ,
		_w3097_,
		_w3101_,
		_w3102_,
		_w3300_
	);
	LUT2 #(
		.INIT('h2)
	) name1551 (
		_w3096_,
		_w3300_,
		_w3301_
	);
	LUT4 #(
		.INIT('h002a)
	) name1552 (
		\u1_u3_adr_r_reg[7]/P0001 ,
		_w3056_,
		_w3061_,
		_w3085_,
		_w3302_
	);
	LUT2 #(
		.INIT('h1)
	) name1553 (
		_w3084_,
		_w3302_,
		_w3303_
	);
	LUT4 #(
		.INIT('h0004)
	) name1554 (
		_w3084_,
		_w3096_,
		_w3300_,
		_w3302_,
		_w3304_
	);
	LUT4 #(
		.INIT('h0b00)
	) name1555 (
		_w3294_,
		_w3296_,
		_w3299_,
		_w3304_,
		_w3305_
	);
	LUT4 #(
		.INIT('h0004)
	) name1556 (
		\u1_u3_adr_r_reg[9]/P0001 ,
		_w3064_,
		_w3065_,
		_w3066_,
		_w3306_
	);
	LUT4 #(
		.INIT('h5070)
	) name1557 (
		_w3096_,
		_w3103_,
		_w3172_,
		_w3306_,
		_w3307_
	);
	LUT2 #(
		.INIT('h1)
	) name1558 (
		\u1_u3_adr_r_reg[13]/P0001 ,
		\u1_u3_out_to_small_r_reg/P0001 ,
		_w3308_
	);
	LUT2 #(
		.INIT('h8)
	) name1559 (
		_w3307_,
		_w3308_,
		_w3309_
	);
	LUT2 #(
		.INIT('h4)
	) name1560 (
		_w3305_,
		_w3309_,
		_w3310_
	);
	LUT2 #(
		.INIT('h2)
	) name1561 (
		\u1_u3_adr_r_reg[13]/P0001 ,
		\u1_u3_out_to_small_r_reg/P0001 ,
		_w3311_
	);
	LUT2 #(
		.INIT('h4)
	) name1562 (
		_w3307_,
		_w3311_,
		_w3312_
	);
	LUT3 #(
		.INIT('h40)
	) name1563 (
		_w3299_,
		_w3304_,
		_w3311_,
		_w3313_
	);
	LUT2 #(
		.INIT('h8)
	) name1564 (
		\u1_u3_out_to_small_r_reg/P0001 ,
		\u4_buf0_reg[13]/P0001 ,
		_w3314_
	);
	LUT4 #(
		.INIT('h0023)
	) name1565 (
		_w3297_,
		_w3312_,
		_w3313_,
		_w3314_,
		_w3315_
	);
	LUT2 #(
		.INIT('hb)
	) name1566 (
		_w3310_,
		_w3315_,
		_w3316_
	);
	LUT4 #(
		.INIT('h0400)
	) name1567 (
		\u1_u1_send_zero_length_r_reg/P0001 ,
		\u1_u1_state_reg[0]/NET0131 ,
		\u1_u1_state_reg[1]/NET0131 ,
		\u1_u2_send_data_r_reg/NET0131 ,
		_w3317_
	);
	LUT4 #(
		.INIT('h0002)
	) name1568 (
		rst_i_pad,
		\u1_u1_state_reg[2]/NET0131 ,
		\u1_u1_state_reg[3]/NET0131 ,
		\u1_u1_state_reg[4]/NET0131 ,
		_w3318_
	);
	LUT2 #(
		.INIT('h8)
	) name1569 (
		_w3317_,
		_w3318_,
		_w3319_
	);
	LUT4 #(
		.INIT('h2000)
	) name1570 (
		rst_i_pad,
		_w1802_,
		_w1803_,
		_w1804_,
		_w3320_
	);
	LUT2 #(
		.INIT('he)
	) name1571 (
		_w3319_,
		_w3320_,
		_w3321_
	);
	LUT4 #(
		.INIT('h5501)
	) name1572 (
		_w3081_,
		_w3116_,
		_w3161_,
		_w3167_,
		_w3322_
	);
	LUT3 #(
		.INIT('h04)
	) name1573 (
		_w3081_,
		_w3293_,
		_w3298_,
		_w3323_
	);
	LUT4 #(
		.INIT('h8000)
	) name1574 (
		\u1_u3_adr_r_reg[11]/P0001 ,
		\u1_u3_adr_r_reg[12]/P0001 ,
		\u1_u3_adr_r_reg[13]/P0001 ,
		\u1_u3_adr_r_reg[14]/P0001 ,
		_w3324_
	);
	LUT3 #(
		.INIT('h80)
	) name1575 (
		_w3251_,
		_w3295_,
		_w3324_,
		_w3325_
	);
	LUT4 #(
		.INIT('h2300)
	) name1576 (
		_w3292_,
		_w3322_,
		_w3323_,
		_w3325_,
		_w3326_
	);
	LUT3 #(
		.INIT('hd0)
	) name1577 (
		_w3096_,
		_w3300_,
		_w3324_,
		_w3327_
	);
	LUT4 #(
		.INIT('hc800)
	) name1578 (
		_w3084_,
		_w3251_,
		_w3302_,
		_w3324_,
		_w3328_
	);
	LUT2 #(
		.INIT('h2)
	) name1579 (
		\u1_u3_adr_r_reg[15]/P0001 ,
		\u1_u3_out_to_small_r_reg/P0001 ,
		_w3329_
	);
	LUT3 #(
		.INIT('h10)
	) name1580 (
		_w3327_,
		_w3328_,
		_w3329_,
		_w3330_
	);
	LUT2 #(
		.INIT('h4)
	) name1581 (
		_w3326_,
		_w3330_,
		_w3331_
	);
	LUT2 #(
		.INIT('h1)
	) name1582 (
		\u1_u3_adr_r_reg[15]/P0001 ,
		\u1_u3_out_to_small_r_reg/P0001 ,
		_w3332_
	);
	LUT3 #(
		.INIT('he0)
	) name1583 (
		_w3327_,
		_w3328_,
		_w3332_,
		_w3333_
	);
	LUT4 #(
		.INIT('h8000)
	) name1584 (
		_w3251_,
		_w3295_,
		_w3324_,
		_w3332_,
		_w3334_
	);
	LUT4 #(
		.INIT('h2300)
	) name1585 (
		_w3292_,
		_w3322_,
		_w3323_,
		_w3334_,
		_w3335_
	);
	LUT2 #(
		.INIT('h8)
	) name1586 (
		\u1_u3_out_to_small_r_reg/P0001 ,
		\u4_buf0_reg[15]/P0001 ,
		_w3336_
	);
	LUT3 #(
		.INIT('h01)
	) name1587 (
		_w3333_,
		_w3335_,
		_w3336_,
		_w3337_
	);
	LUT2 #(
		.INIT('hb)
	) name1588 (
		_w3331_,
		_w3337_,
		_w3338_
	);
	LUT3 #(
		.INIT('h51)
	) name1589 (
		\u1_u3_adr_r_reg[11]/P0001 ,
		_w3096_,
		_w3300_,
		_w3339_
	);
	LUT4 #(
		.INIT('h5040)
	) name1590 (
		\u1_u3_adr_r_reg[11]/P0001 ,
		_w3084_,
		_w3251_,
		_w3302_,
		_w3340_
	);
	LUT2 #(
		.INIT('h1)
	) name1591 (
		_w3339_,
		_w3340_,
		_w3341_
	);
	LUT2 #(
		.INIT('h8)
	) name1592 (
		_w3251_,
		_w3295_,
		_w3342_
	);
	LUT3 #(
		.INIT('h40)
	) name1593 (
		\u1_u3_adr_r_reg[11]/P0001 ,
		_w3251_,
		_w3295_,
		_w3343_
	);
	LUT4 #(
		.INIT('h2300)
	) name1594 (
		_w3292_,
		_w3322_,
		_w3323_,
		_w3343_,
		_w3344_
	);
	LUT4 #(
		.INIT('h2300)
	) name1595 (
		_w3292_,
		_w3322_,
		_w3323_,
		_w3342_,
		_w3345_
	);
	LUT3 #(
		.INIT('hc8)
	) name1596 (
		_w3084_,
		_w3251_,
		_w3302_,
		_w3346_
	);
	LUT3 #(
		.INIT('h08)
	) name1597 (
		\u1_u3_adr_r_reg[11]/P0001 ,
		_w3301_,
		_w3346_,
		_w3347_
	);
	LUT4 #(
		.INIT('h2022)
	) name1598 (
		_w3341_,
		_w3344_,
		_w3345_,
		_w3347_,
		_w3348_
	);
	LUT3 #(
		.INIT('h8d)
	) name1599 (
		\u1_u3_out_to_small_r_reg/P0001 ,
		\u4_buf0_reg[11]/P0001 ,
		_w3348_,
		_w3349_
	);
	LUT4 #(
		.INIT('h5559)
	) name1600 (
		\u1_u3_adr_r_reg[6]/P0001 ,
		_w3077_,
		_w3078_,
		_w3079_,
		_w3350_
	);
	LUT2 #(
		.INIT('h1)
	) name1601 (
		\u1_u3_out_to_small_r_reg/P0001 ,
		_w3350_,
		_w3351_
	);
	LUT4 #(
		.INIT('hef00)
	) name1602 (
		_w3136_,
		_w3158_,
		_w3165_,
		_w3351_,
		_w3352_
	);
	LUT3 #(
		.INIT('h15)
	) name1603 (
		\u1_u3_out_to_small_r_reg/P0001 ,
		_w3077_,
		_w3166_,
		_w3353_
	);
	LUT4 #(
		.INIT('h0100)
	) name1604 (
		_w3081_,
		_w3161_,
		_w3164_,
		_w3353_,
		_w3354_
	);
	LUT2 #(
		.INIT('h8)
	) name1605 (
		\u1_u3_out_to_small_r_reg/P0001 ,
		\u4_buf0_reg[6]/P0001 ,
		_w3355_
	);
	LUT4 #(
		.INIT('h00ef)
	) name1606 (
		_w3136_,
		_w3158_,
		_w3354_,
		_w3355_,
		_w3356_
	);
	LUT2 #(
		.INIT('hb)
	) name1607 (
		_w3352_,
		_w3356_,
		_w3357_
	);
	LUT4 #(
		.INIT('hdedd)
	) name1608 (
		\u1_u3_adr_r_reg[8]/P0001 ,
		\u1_u3_out_to_small_r_reg/P0001 ,
		_w3055_,
		_w3061_,
		_w3358_
	);
	LUT4 #(
		.INIT('h00fe)
	) name1609 (
		_w3082_,
		_w3086_,
		_w3168_,
		_w3358_,
		_w3359_
	);
	LUT4 #(
		.INIT('hef00)
	) name1610 (
		_w3136_,
		_w3158_,
		_w3254_,
		_w3359_,
		_w3360_
	);
	LUT4 #(
		.INIT('h1211)
	) name1611 (
		\u1_u3_adr_r_reg[8]/P0001 ,
		\u1_u3_out_to_small_r_reg/P0001 ,
		_w3055_,
		_w3061_,
		_w3361_
	);
	LUT2 #(
		.INIT('h8)
	) name1612 (
		\u1_u3_out_to_small_r_reg/P0001 ,
		\u4_buf0_reg[8]/P0001 ,
		_w3362_
	);
	LUT2 #(
		.INIT('h1)
	) name1613 (
		_w3361_,
		_w3362_,
		_w3363_
	);
	LUT4 #(
		.INIT('h00fe)
	) name1614 (
		_w3082_,
		_w3086_,
		_w3168_,
		_w3362_,
		_w3364_
	);
	LUT4 #(
		.INIT('hef00)
	) name1615 (
		_w3136_,
		_w3158_,
		_w3254_,
		_w3364_,
		_w3365_
	);
	LUT3 #(
		.INIT('hab)
	) name1616 (
		_w3360_,
		_w3363_,
		_w3365_,
		_w3366_
	);
	LUT4 #(
		.INIT('h5559)
	) name1617 (
		\u1_u3_adr_r_reg[9]/P0001 ,
		_w3064_,
		_w3065_,
		_w3066_,
		_w3367_
	);
	LUT2 #(
		.INIT('h4)
	) name1618 (
		\u1_u3_out_to_small_r_reg/P0001 ,
		_w3367_,
		_w3368_
	);
	LUT3 #(
		.INIT('h40)
	) name1619 (
		_w3299_,
		_w3303_,
		_w3368_,
		_w3369_
	);
	LUT2 #(
		.INIT('h8)
	) name1620 (
		\u1_u3_out_to_small_r_reg/P0001 ,
		\u4_buf0_reg[9]/P0001 ,
		_w3370_
	);
	LUT3 #(
		.INIT('h72)
	) name1621 (
		\u1_u3_out_to_small_r_reg/P0001 ,
		\u4_buf0_reg[9]/P0001 ,
		_w3367_,
		_w3371_
	);
	LUT3 #(
		.INIT('h04)
	) name1622 (
		_w3299_,
		_w3303_,
		_w3370_,
		_w3372_
	);
	LUT4 #(
		.INIT('h4e4f)
	) name1623 (
		_w3297_,
		_w3369_,
		_w3371_,
		_w3372_,
		_w3373_
	);
	LUT3 #(
		.INIT('h8a)
	) name1624 (
		rst_i_pad,
		_w1805_,
		_w1820_,
		_w3374_
	);
	LUT2 #(
		.INIT('h2)
	) name1625 (
		\u1_u3_new_size_reg[12]/P0001 ,
		\u1_u3_out_to_small_r_reg/P0001 ,
		_w3375_
	);
	LUT3 #(
		.INIT('hd0)
	) name1626 (
		_w3144_,
		_w3154_,
		_w3157_,
		_w3376_
	);
	LUT4 #(
		.INIT('h54fe)
	) name1627 (
		\u1_u3_adr_r_reg[4]/P0001 ,
		_w3112_,
		_w3113_,
		_w3163_,
		_w3377_
	);
	LUT4 #(
		.INIT('h00d0)
	) name1628 (
		_w3144_,
		_w3154_,
		_w3157_,
		_w3377_,
		_w3378_
	);
	LUT4 #(
		.INIT('h00da)
	) name1629 (
		_w3135_,
		_w3376_,
		_w3377_,
		_w3378_,
		_w3379_
	);
	LUT3 #(
		.INIT('h8d)
	) name1630 (
		\u1_u3_out_to_small_r_reg/P0001 ,
		\u4_buf0_reg[4]/P0001 ,
		_w3379_,
		_w3380_
	);
	LUT2 #(
		.INIT('h1)
	) name1631 (
		_w3115_,
		_w3293_,
		_w3381_
	);
	LUT4 #(
		.INIT('h4050)
	) name1632 (
		_w3115_,
		_w3154_,
		_w3157_,
		_w3291_,
		_w3382_
	);
	LUT4 #(
		.INIT('h54fe)
	) name1633 (
		\u1_u3_adr_r_reg[5]/P0001 ,
		_w3107_,
		_w3108_,
		_w3160_,
		_w3383_
	);
	LUT4 #(
		.INIT('hfeab)
	) name1634 (
		\u1_u3_out_to_small_r_reg/P0001 ,
		_w3381_,
		_w3382_,
		_w3383_,
		_w3384_
	);
	LUT2 #(
		.INIT('h8)
	) name1635 (
		\u1_u3_out_to_small_r_reg/P0001 ,
		\u4_buf0_reg[5]/P0001 ,
		_w3385_
	);
	LUT2 #(
		.INIT('hd)
	) name1636 (
		_w3384_,
		_w3385_,
		_w3386_
	);
	LUT4 #(
		.INIT('h5559)
	) name1637 (
		\u1_u3_adr_r_reg[7]/P0001 ,
		_w3071_,
		_w3072_,
		_w3073_,
		_w3387_
	);
	LUT2 #(
		.INIT('h1)
	) name1638 (
		\u1_u3_out_to_small_r_reg/P0001 ,
		_w3387_,
		_w3388_
	);
	LUT4 #(
		.INIT('h2300)
	) name1639 (
		_w3292_,
		_w3322_,
		_w3323_,
		_w3388_,
		_w3389_
	);
	LUT2 #(
		.INIT('h4)
	) name1640 (
		\u1_u3_out_to_small_r_reg/P0001 ,
		_w3387_,
		_w3390_
	);
	LUT4 #(
		.INIT('hdc00)
	) name1641 (
		_w3292_,
		_w3322_,
		_w3323_,
		_w3390_,
		_w3391_
	);
	LUT2 #(
		.INIT('h8)
	) name1642 (
		\u1_u3_out_to_small_r_reg/P0001 ,
		\u4_buf0_reg[7]/P0001 ,
		_w3392_
	);
	LUT3 #(
		.INIT('hfe)
	) name1643 (
		_w3389_,
		_w3391_,
		_w3392_,
		_w3393_
	);
	LUT2 #(
		.INIT('h2)
	) name1644 (
		\u1_u3_new_size_reg[13]/P0001 ,
		\u1_u3_out_to_small_r_reg/P0001 ,
		_w3394_
	);
	LUT2 #(
		.INIT('h4)
	) name1645 (
		\u4_u2_csr1_reg[11]/P0001 ,
		\u4_u2_csr1_reg[12]/P0001 ,
		_w3395_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name1646 (
		\dma_ack_i[2]_pad ,
		\u4_u2_csr1_reg[11]/P0001 ,
		\u4_u2_csr1_reg[12]/P0001 ,
		\u4_u2_dma_req_out_hold_reg/P0001 ,
		_w3396_
	);
	LUT2 #(
		.INIT('h2)
	) name1647 (
		\u4_u2_r1_reg/P0001 ,
		\u4_u2_r2_reg/P0001 ,
		_w3397_
	);
	LUT4 #(
		.INIT('hb000)
	) name1648 (
		\u4_u2_csr1_reg[11]/P0001 ,
		\u4_u2_csr1_reg[12]/P0001 ,
		\u4_u2_dma_req_in_hold2_reg/P0001 ,
		\u4_u2_dma_req_in_hold_reg/P0001 ,
		_w3398_
	);
	LUT4 #(
		.INIT('h88c8)
	) name1649 (
		\dma_req_o[2]_pad ,
		rst_i_pad,
		\u4_u2_r1_reg/P0001 ,
		\u4_u2_r2_reg/P0001 ,
		_w3399_
	);
	LUT4 #(
		.INIT('hfd00)
	) name1650 (
		_w3396_,
		_w3397_,
		_w3398_,
		_w3399_,
		_w3400_
	);
	LUT2 #(
		.INIT('h4)
	) name1651 (
		\u4_u3_csr1_reg[11]/P0001 ,
		\u4_u3_csr1_reg[12]/P0001 ,
		_w3401_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name1652 (
		\dma_ack_i[3]_pad ,
		\u4_u3_csr1_reg[11]/P0001 ,
		\u4_u3_csr1_reg[12]/P0001 ,
		\u4_u3_dma_req_out_hold_reg/P0001 ,
		_w3402_
	);
	LUT2 #(
		.INIT('h2)
	) name1653 (
		\u4_u3_r1_reg/P0001 ,
		\u4_u3_r2_reg/P0001 ,
		_w3403_
	);
	LUT4 #(
		.INIT('hb000)
	) name1654 (
		\u4_u3_csr1_reg[11]/P0001 ,
		\u4_u3_csr1_reg[12]/P0001 ,
		\u4_u3_dma_req_in_hold2_reg/P0001 ,
		\u4_u3_dma_req_in_hold_reg/P0001 ,
		_w3404_
	);
	LUT4 #(
		.INIT('h88c8)
	) name1655 (
		\dma_req_o[3]_pad ,
		rst_i_pad,
		\u4_u3_r1_reg/P0001 ,
		\u4_u3_r2_reg/P0001 ,
		_w3405_
	);
	LUT4 #(
		.INIT('hfd00)
	) name1656 (
		_w3402_,
		_w3403_,
		_w3404_,
		_w3405_,
		_w3406_
	);
	LUT2 #(
		.INIT('h4)
	) name1657 (
		\u4_u0_csr1_reg[11]/P0001 ,
		\u4_u0_csr1_reg[12]/P0001 ,
		_w3407_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name1658 (
		\dma_ack_i[0]_pad ,
		\u4_u0_csr1_reg[11]/P0001 ,
		\u4_u0_csr1_reg[12]/P0001 ,
		\u4_u0_dma_req_out_hold_reg/P0001 ,
		_w3408_
	);
	LUT2 #(
		.INIT('h2)
	) name1659 (
		\u4_u0_r1_reg/P0001 ,
		\u4_u0_r2_reg/P0001 ,
		_w3409_
	);
	LUT4 #(
		.INIT('hb000)
	) name1660 (
		\u4_u0_csr1_reg[11]/P0001 ,
		\u4_u0_csr1_reg[12]/P0001 ,
		\u4_u0_dma_req_in_hold2_reg/P0001 ,
		\u4_u0_dma_req_in_hold_reg/P0001 ,
		_w3410_
	);
	LUT4 #(
		.INIT('h88c8)
	) name1661 (
		\dma_req_o[0]_pad ,
		rst_i_pad,
		\u4_u0_r1_reg/P0001 ,
		\u4_u0_r2_reg/P0001 ,
		_w3411_
	);
	LUT4 #(
		.INIT('hfd00)
	) name1662 (
		_w3408_,
		_w3409_,
		_w3410_,
		_w3411_,
		_w3412_
	);
	LUT2 #(
		.INIT('h4)
	) name1663 (
		\u4_u1_csr1_reg[11]/P0001 ,
		\u4_u1_csr1_reg[12]/P0001 ,
		_w3413_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name1664 (
		\dma_ack_i[1]_pad ,
		\u4_u1_csr1_reg[11]/P0001 ,
		\u4_u1_csr1_reg[12]/P0001 ,
		\u4_u1_dma_req_out_hold_reg/P0001 ,
		_w3414_
	);
	LUT2 #(
		.INIT('h2)
	) name1665 (
		\u4_u1_r1_reg/P0001 ,
		\u4_u1_r2_reg/P0001 ,
		_w3415_
	);
	LUT4 #(
		.INIT('hb000)
	) name1666 (
		\u4_u1_csr1_reg[11]/P0001 ,
		\u4_u1_csr1_reg[12]/P0001 ,
		\u4_u1_dma_req_in_hold2_reg/P0001 ,
		\u4_u1_dma_req_in_hold_reg/P0001 ,
		_w3416_
	);
	LUT4 #(
		.INIT('h88c8)
	) name1667 (
		\dma_req_o[1]_pad ,
		rst_i_pad,
		\u4_u1_r1_reg/P0001 ,
		\u4_u1_r2_reg/P0001 ,
		_w3417_
	);
	LUT4 #(
		.INIT('hfd00)
	) name1668 (
		_w3414_,
		_w3415_,
		_w3416_,
		_w3417_,
		_w3418_
	);
	LUT4 #(
		.INIT('h8880)
	) name1669 (
		\u1_u3_buffer_done_reg/P0001 ,
		\u4_csr_reg[15]/NET0131 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		_w3419_
	);
	LUT2 #(
		.INIT('h2)
	) name1670 (
		\u1_u3_state_reg[8]/P0001 ,
		_w3419_,
		_w3420_
	);
	LUT3 #(
		.INIT('he2)
	) name1671 (
		\u1_u3_next_dpid_reg[0]/P0001 ,
		\u1_u3_out_to_small_r_reg/P0001 ,
		\u4_buf0_reg[2]/P0001 ,
		_w3421_
	);
	LUT3 #(
		.INIT('hd0)
	) name1672 (
		\u1_u3_state_reg[8]/P0001 ,
		_w3419_,
		_w3421_,
		_w3422_
	);
	LUT4 #(
		.INIT('h5a59)
	) name1673 (
		\u1_u3_adr_r_reg[2]/P0001 ,
		_w3093_,
		_w3127_,
		_w3131_,
		_w3423_
	);
	LUT4 #(
		.INIT('h20d0)
	) name1674 (
		_w3144_,
		_w3154_,
		_w3420_,
		_w3423_,
		_w3424_
	);
	LUT2 #(
		.INIT('he)
	) name1675 (
		_w3422_,
		_w3424_,
		_w3425_
	);
	LUT3 #(
		.INIT('he2)
	) name1676 (
		\u1_u3_next_dpid_reg[1]/P0001 ,
		\u1_u3_out_to_small_r_reg/P0001 ,
		\u4_buf0_reg[3]/P0001 ,
		_w3426_
	);
	LUT3 #(
		.INIT('hd0)
	) name1677 (
		\u1_u3_state_reg[8]/P0001 ,
		_w3419_,
		_w3426_,
		_w3427_
	);
	LUT4 #(
		.INIT('h80a0)
	) name1678 (
		_w3124_,
		_w3154_,
		_w3157_,
		_w3291_,
		_w3428_
	);
	LUT4 #(
		.INIT('h00c8)
	) name1679 (
		\u1_u3_adr_r_reg[2]/P0001 ,
		\u1_u3_state_reg[8]/P0001 ,
		_w3127_,
		_w3419_,
		_w3429_
	);
	LUT3 #(
		.INIT('h02)
	) name1680 (
		\u1_u3_state_reg[8]/P0001 ,
		_w3093_,
		_w3419_,
		_w3430_
	);
	LUT3 #(
		.INIT('h23)
	) name1681 (
		_w3131_,
		_w3429_,
		_w3430_,
		_w3431_
	);
	LUT3 #(
		.INIT('h0b)
	) name1682 (
		_w3154_,
		_w3291_,
		_w3431_,
		_w3432_
	);
	LUT4 #(
		.INIT('h00c8)
	) name1683 (
		\u1_u3_adr_r_reg[3]/P0001 ,
		\u1_u3_state_reg[8]/P0001 ,
		_w3117_,
		_w3419_,
		_w3433_
	);
	LUT3 #(
		.INIT('h0b)
	) name1684 (
		_w3121_,
		_w3430_,
		_w3433_,
		_w3434_
	);
	LUT2 #(
		.INIT('h2)
	) name1685 (
		_w3124_,
		_w3434_,
		_w3435_
	);
	LUT4 #(
		.INIT('hbbba)
	) name1686 (
		_w3427_,
		_w3428_,
		_w3432_,
		_w3435_,
		_w3436_
	);
	LUT3 #(
		.INIT('h08)
	) name1687 (
		\u1_u3_new_sizeb_reg[3]/P0001 ,
		_w2810_,
		_w2812_,
		_w3437_
	);
	LUT3 #(
		.INIT('h51)
	) name1688 (
		\u1_u3_new_sizeb_reg[2]/P0001 ,
		_w2795_,
		_w2797_,
		_w3438_
	);
	LUT3 #(
		.INIT('h71)
	) name1689 (
		\u1_u3_new_sizeb_reg[3]/P0001 ,
		_w2813_,
		_w3438_,
		_w3439_
	);
	LUT3 #(
		.INIT('h08)
	) name1690 (
		\u1_u3_new_sizeb_reg[0]/P0001 ,
		_w2788_,
		_w2790_,
		_w3440_
	);
	LUT3 #(
		.INIT('he8)
	) name1691 (
		\u1_u3_new_sizeb_reg[1]/P0001 ,
		_w2785_,
		_w3440_,
		_w3441_
	);
	LUT3 #(
		.INIT('h08)
	) name1692 (
		\u1_u3_new_sizeb_reg[2]/P0001 ,
		_w2795_,
		_w2797_,
		_w3442_
	);
	LUT2 #(
		.INIT('h1)
	) name1693 (
		_w3437_,
		_w3442_,
		_w3443_
	);
	LUT3 #(
		.INIT('h08)
	) name1694 (
		\u1_u3_new_sizeb_reg[7]/P0001 ,
		_w2830_,
		_w2832_,
		_w3444_
	);
	LUT3 #(
		.INIT('h08)
	) name1695 (
		\u1_u3_new_sizeb_reg[6]/P0001 ,
		_w2860_,
		_w2862_,
		_w3445_
	);
	LUT2 #(
		.INIT('h1)
	) name1696 (
		_w3444_,
		_w3445_,
		_w3446_
	);
	LUT3 #(
		.INIT('h08)
	) name1697 (
		\u1_u3_new_sizeb_reg[5]/P0001 ,
		_w2820_,
		_w2822_,
		_w3447_
	);
	LUT3 #(
		.INIT('h08)
	) name1698 (
		\u1_u3_new_sizeb_reg[4]/P0001 ,
		_w2803_,
		_w2805_,
		_w3448_
	);
	LUT2 #(
		.INIT('h1)
	) name1699 (
		_w3447_,
		_w3448_,
		_w3449_
	);
	LUT4 #(
		.INIT('h0001)
	) name1700 (
		_w3444_,
		_w3445_,
		_w3447_,
		_w3448_,
		_w3450_
	);
	LUT4 #(
		.INIT('hba00)
	) name1701 (
		_w3439_,
		_w3441_,
		_w3443_,
		_w3450_,
		_w3451_
	);
	LUT3 #(
		.INIT('h51)
	) name1702 (
		\u1_u3_new_sizeb_reg[5]/P0001 ,
		_w2820_,
		_w2822_,
		_w3452_
	);
	LUT3 #(
		.INIT('h51)
	) name1703 (
		\u1_u3_new_sizeb_reg[4]/P0001 ,
		_w2803_,
		_w2805_,
		_w3453_
	);
	LUT3 #(
		.INIT('h8e)
	) name1704 (
		\u1_u3_new_sizeb_reg[5]/P0001 ,
		_w2823_,
		_w3453_,
		_w3454_
	);
	LUT2 #(
		.INIT('h2)
	) name1705 (
		_w3446_,
		_w3454_,
		_w3455_
	);
	LUT3 #(
		.INIT('h51)
	) name1706 (
		\u1_u3_new_sizeb_reg[9]/P0001 ,
		_w2852_,
		_w2854_,
		_w3456_
	);
	LUT3 #(
		.INIT('h08)
	) name1707 (
		\u1_u3_new_sizeb_reg[9]/P0001 ,
		_w2852_,
		_w2854_,
		_w3457_
	);
	LUT3 #(
		.INIT('h51)
	) name1708 (
		\u1_u3_new_sizeb_reg[8]/P0001 ,
		_w2837_,
		_w2839_,
		_w3458_
	);
	LUT3 #(
		.INIT('h8e)
	) name1709 (
		\u1_u3_new_sizeb_reg[9]/P0001 ,
		_w2855_,
		_w3458_,
		_w3459_
	);
	LUT3 #(
		.INIT('h51)
	) name1710 (
		\u1_u3_new_sizeb_reg[7]/P0001 ,
		_w2830_,
		_w2832_,
		_w3460_
	);
	LUT3 #(
		.INIT('h51)
	) name1711 (
		\u1_u3_new_sizeb_reg[6]/P0001 ,
		_w2860_,
		_w2862_,
		_w3461_
	);
	LUT3 #(
		.INIT('h8e)
	) name1712 (
		\u1_u3_new_sizeb_reg[7]/P0001 ,
		_w2833_,
		_w3461_,
		_w3462_
	);
	LUT4 #(
		.INIT('hd000)
	) name1713 (
		_w3446_,
		_w3454_,
		_w3459_,
		_w3462_,
		_w3463_
	);
	LUT3 #(
		.INIT('h08)
	) name1714 (
		\u1_u3_new_sizeb_reg[10]/P0001 ,
		_w2845_,
		_w2847_,
		_w3464_
	);
	LUT3 #(
		.INIT('h08)
	) name1715 (
		\u1_u3_new_sizeb_reg[8]/P0001 ,
		_w2837_,
		_w2839_,
		_w3465_
	);
	LUT4 #(
		.INIT('h137f)
	) name1716 (
		\u1_u3_new_sizeb_reg[8]/P0001 ,
		\u1_u3_new_sizeb_reg[9]/P0001 ,
		_w2840_,
		_w2855_,
		_w3466_
	);
	LUT2 #(
		.INIT('h4)
	) name1717 (
		_w3464_,
		_w3466_,
		_w3467_
	);
	LUT3 #(
		.INIT('h51)
	) name1718 (
		\u1_u3_new_sizeb_reg[10]/P0001 ,
		_w2845_,
		_w2847_,
		_w3468_
	);
	LUT2 #(
		.INIT('h2)
	) name1719 (
		_w2884_,
		_w3468_,
		_w3469_
	);
	LUT4 #(
		.INIT('h4f00)
	) name1720 (
		_w3451_,
		_w3463_,
		_w3467_,
		_w3469_,
		_w3470_
	);
	LUT2 #(
		.INIT('h2)
	) name1721 (
		_w2885_,
		_w3468_,
		_w3471_
	);
	LUT4 #(
		.INIT('h4f00)
	) name1722 (
		_w3451_,
		_w3463_,
		_w3467_,
		_w3471_,
		_w3472_
	);
	LUT3 #(
		.INIT('hf1)
	) name1723 (
		_w2878_,
		_w3470_,
		_w3472_,
		_w3473_
	);
	LUT4 #(
		.INIT('h0777)
	) name1724 (
		_w1803_,
		_w1804_,
		_w1807_,
		_w1808_,
		_w3474_
	);
	LUT2 #(
		.INIT('h8)
	) name1725 (
		_w1816_,
		_w3474_,
		_w3475_
	);
	LUT2 #(
		.INIT('h7)
	) name1726 (
		_w1816_,
		_w3474_,
		_w3476_
	);
	LUT2 #(
		.INIT('h1)
	) name1727 (
		\u0_u0_drive_k_reg/P0001 ,
		\u1_u3_send_token_reg/P0001 ,
		_w3477_
	);
	LUT4 #(
		.INIT('h00fb)
	) name1728 (
		TxReady_pad_i_pad,
		TxValid_pad_o_pad,
		\u0_drive_k_r_reg/P0001 ,
		\u0_tx_ready_reg/NET0131 ,
		_w3478_
	);
	LUT3 #(
		.INIT('h70)
	) name1729 (
		_w1806_,
		_w1809_,
		_w3478_,
		_w3479_
	);
	LUT4 #(
		.INIT('hfb00)
	) name1730 (
		TxReady_pad_i_pad,
		TxValid_pad_o_pad,
		\u0_drive_k_r_reg/P0001 ,
		\u0_tx_ready_reg/NET0131 ,
		_w3480_
	);
	LUT3 #(
		.INIT('h70)
	) name1731 (
		_w1807_,
		_w1815_,
		_w3480_,
		_w3481_
	);
	LUT3 #(
		.INIT('ha8)
	) name1732 (
		_w3477_,
		_w3479_,
		_w3481_,
		_w3482_
	);
	LUT3 #(
		.INIT('h2a)
	) name1733 (
		rst_i_pad,
		_w3475_,
		_w3482_,
		_w3483_
	);
	LUT4 #(
		.INIT('h5a59)
	) name1734 (
		\u1_u3_adr_r_reg[1]/P0001 ,
		_w3093_,
		_w3137_,
		_w3141_,
		_w3484_
	);
	LUT4 #(
		.INIT('h004c)
	) name1735 (
		\u1_u3_adr_r_reg[0]/P0001 ,
		\u1_u3_state_reg[8]/P0001 ,
		_w3147_,
		_w3419_,
		_w3485_
	);
	LUT2 #(
		.INIT('h4)
	) name1736 (
		_w3153_,
		_w3485_,
		_w3486_
	);
	LUT2 #(
		.INIT('h8)
	) name1737 (
		\u1_u3_out_to_small_r_reg/P0001 ,
		\u4_buf0_reg[1]/P0001 ,
		_w3487_
	);
	LUT4 #(
		.INIT('h1115)
	) name1738 (
		\u1_u3_out_to_small_r_reg/P0001 ,
		\u4_csr_reg[15]/NET0131 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		_w3488_
	);
	LUT3 #(
		.INIT('h78)
	) name1739 (
		\u1_u3_buffer_done_reg/P0001 ,
		\u4_csr_reg[30]/NET0131 ,
		\u4_csr_reg[31]/P0001 ,
		_w3489_
	);
	LUT3 #(
		.INIT('h15)
	) name1740 (
		_w3487_,
		_w3488_,
		_w3489_,
		_w3490_
	);
	LUT2 #(
		.INIT('h1)
	) name1741 (
		_w3420_,
		_w3490_,
		_w3491_
	);
	LUT4 #(
		.INIT('h0080)
	) name1742 (
		\u1_u3_adr_r_reg[0]/P0001 ,
		\u1_u3_state_reg[8]/P0001 ,
		_w3147_,
		_w3419_,
		_w3492_
	);
	LUT3 #(
		.INIT('h08)
	) name1743 (
		\u1_u3_state_reg[8]/P0001 ,
		_w3152_,
		_w3419_,
		_w3493_
	);
	LUT3 #(
		.INIT('h23)
	) name1744 (
		_w3151_,
		_w3492_,
		_w3493_,
		_w3494_
	);
	LUT4 #(
		.INIT('hf8fd)
	) name1745 (
		_w3484_,
		_w3486_,
		_w3491_,
		_w3494_,
		_w3495_
	);
	LUT3 #(
		.INIT('hac)
	) name1746 (
		\u1_u2_sizu_c_reg[10]/P0001 ,
		\u1_u3_new_size_reg[10]/P0001 ,
		\u1_u3_out_to_small_r_reg/P0001 ,
		_w3496_
	);
	LUT2 #(
		.INIT('h4)
	) name1747 (
		_w2884_,
		_w3468_,
		_w3497_
	);
	LUT2 #(
		.INIT('h1)
	) name1748 (
		_w2884_,
		_w3464_,
		_w3498_
	);
	LUT2 #(
		.INIT('h8)
	) name1749 (
		_w3466_,
		_w3498_,
		_w3499_
	);
	LUT4 #(
		.INIT('h040f)
	) name1750 (
		_w3451_,
		_w3463_,
		_w3497_,
		_w3499_,
		_w3500_
	);
	LUT2 #(
		.INIT('hb)
	) name1751 (
		_w3470_,
		_w3500_,
		_w3501_
	);
	LUT4 #(
		.INIT('he080)
	) name1752 (
		\u1_u3_new_sizeb_reg[10]/P0001 ,
		_w2848_,
		_w2885_,
		_w3457_,
		_w3502_
	);
	LUT3 #(
		.INIT('h01)
	) name1753 (
		_w3444_,
		_w3445_,
		_w3465_,
		_w3503_
	);
	LUT4 #(
		.INIT('h0001)
	) name1754 (
		\u1_u3_new_sizeb_reg[6]/P0001 ,
		_w2863_,
		_w3444_,
		_w3465_,
		_w3504_
	);
	LUT2 #(
		.INIT('h1)
	) name1755 (
		_w3452_,
		_w3453_,
		_w3505_
	);
	LUT4 #(
		.INIT('h4500)
	) name1756 (
		_w3439_,
		_w3441_,
		_w3443_,
		_w3505_,
		_w3506_
	);
	LUT3 #(
		.INIT('he8)
	) name1757 (
		\u1_u3_new_sizeb_reg[5]/P0001 ,
		_w2823_,
		_w3448_,
		_w3507_
	);
	LUT2 #(
		.INIT('h2)
	) name1758 (
		_w3503_,
		_w3507_,
		_w3508_
	);
	LUT3 #(
		.INIT('h45)
	) name1759 (
		_w3504_,
		_w3506_,
		_w3508_,
		_w3509_
	);
	LUT4 #(
		.INIT('h80e0)
	) name1760 (
		\u1_u3_new_sizeb_reg[10]/P0001 ,
		_w2848_,
		_w2885_,
		_w3456_,
		_w3510_
	);
	LUT3 #(
		.INIT('h8e)
	) name1761 (
		\u1_u3_new_sizeb_reg[8]/P0001 ,
		_w2840_,
		_w3460_,
		_w3511_
	);
	LUT2 #(
		.INIT('h8)
	) name1762 (
		_w3510_,
		_w3511_,
		_w3512_
	);
	LUT3 #(
		.INIT('h40)
	) name1763 (
		_w2891_,
		_w3510_,
		_w3511_,
		_w3513_
	);
	LUT4 #(
		.INIT('h4500)
	) name1764 (
		_w3504_,
		_w3506_,
		_w3508_,
		_w3513_,
		_w3514_
	);
	LUT4 #(
		.INIT('h4500)
	) name1765 (
		_w3504_,
		_w3506_,
		_w3508_,
		_w3512_,
		_w3515_
	);
	LUT4 #(
		.INIT('h0b09)
	) name1766 (
		_w2891_,
		_w3502_,
		_w3514_,
		_w3515_,
		_w3516_
	);
	LUT2 #(
		.INIT('h4)
	) name1767 (
		\u1_u2_dtmp_sel_r_reg/P0001 ,
		\u1_u2_mack_r_reg/P0001 ,
		_w3517_
	);
	LUT4 #(
		.INIT('h0800)
	) name1768 (
		\u1_u2_adr_cw_reg[0]/NET0131 ,
		\u1_u2_adr_cw_reg[1]/P0001 ,
		\u1_u2_dtmp_sel_r_reg/P0001 ,
		\u1_u2_mack_r_reg/P0001 ,
		_w3518_
	);
	LUT2 #(
		.INIT('h8)
	) name1769 (
		\u1_u2_adr_cw_reg[2]/P0001 ,
		\u1_u2_adr_cw_reg[3]/NET0131 ,
		_w3519_
	);
	LUT4 #(
		.INIT('hdeee)
	) name1770 (
		\u1_u2_adr_cw_reg[4]/P0001 ,
		\u1_u2_last_buf_adr_reg[4]/P0001 ,
		_w3518_,
		_w3519_,
		_w3520_
	);
	LUT3 #(
		.INIT('h15)
	) name1771 (
		\u1_u2_adr_cw_reg[4]/P0001 ,
		_w3518_,
		_w3519_,
		_w3521_
	);
	LUT3 #(
		.INIT('h80)
	) name1772 (
		\u1_u2_adr_cw_reg[2]/P0001 ,
		\u1_u2_adr_cw_reg[3]/NET0131 ,
		\u1_u2_adr_cw_reg[4]/P0001 ,
		_w3522_
	);
	LUT2 #(
		.INIT('h8)
	) name1773 (
		_w3518_,
		_w3522_,
		_w3523_
	);
	LUT3 #(
		.INIT('h2a)
	) name1774 (
		\u1_u2_last_buf_adr_reg[4]/P0001 ,
		_w3518_,
		_w3522_,
		_w3524_
	);
	LUT4 #(
		.INIT('h060c)
	) name1775 (
		\u1_u2_adr_cw_reg[2]/P0001 ,
		\u1_u2_adr_cw_reg[3]/NET0131 ,
		\u1_u2_last_buf_adr_reg[3]/P0001 ,
		_w3518_,
		_w3525_
	);
	LUT4 #(
		.INIT('h0075)
	) name1776 (
		_w3520_,
		_w3521_,
		_w3524_,
		_w3525_,
		_w3526_
	);
	LUT4 #(
		.INIT('h963c)
	) name1777 (
		\u1_u2_adr_cw_reg[0]/NET0131 ,
		\u1_u2_adr_cw_reg[1]/P0001 ,
		\u1_u2_last_buf_adr_reg[1]/P0001 ,
		_w3517_,
		_w3527_
	);
	LUT4 #(
		.INIT('h695a)
	) name1778 (
		\u1_u2_adr_cw_reg[0]/NET0131 ,
		\u1_u2_dtmp_sel_r_reg/P0001 ,
		\u1_u2_last_buf_adr_reg[0]/P0001 ,
		\u1_u2_mack_r_reg/P0001 ,
		_w3528_
	);
	LUT2 #(
		.INIT('h2)
	) name1779 (
		_w2122_,
		_w3528_,
		_w3529_
	);
	LUT4 #(
		.INIT('h6fcf)
	) name1780 (
		\u1_u2_adr_cw_reg[2]/P0001 ,
		\u1_u2_adr_cw_reg[3]/NET0131 ,
		\u1_u2_last_buf_adr_reg[3]/P0001 ,
		_w3518_,
		_w3530_
	);
	LUT3 #(
		.INIT('h96)
	) name1781 (
		\u1_u2_adr_cw_reg[2]/P0001 ,
		\u1_u2_last_buf_adr_reg[2]/P0001 ,
		_w3518_,
		_w3531_
	);
	LUT4 #(
		.INIT('h0040)
	) name1782 (
		_w3527_,
		_w3529_,
		_w3530_,
		_w3531_,
		_w3532_
	);
	LUT4 #(
		.INIT('h7bbb)
	) name1783 (
		\u1_u2_adr_cw_reg[5]/NET0131 ,
		\u1_u2_last_buf_adr_reg[5]/P0001 ,
		_w3518_,
		_w3522_,
		_w3533_
	);
	LUT4 #(
		.INIT('h0080)
	) name1784 (
		\u1_u2_adr_cw_reg[2]/P0001 ,
		\u1_u2_adr_cw_reg[3]/NET0131 ,
		\u1_u2_adr_cw_reg[4]/P0001 ,
		\u1_u2_adr_cw_reg[5]/NET0131 ,
		_w3534_
	);
	LUT3 #(
		.INIT('h40)
	) name1785 (
		\u1_u2_last_buf_adr_reg[5]/P0001 ,
		_w3518_,
		_w3534_,
		_w3535_
	);
	LUT2 #(
		.INIT('h2)
	) name1786 (
		\u1_u2_adr_cw_reg[5]/NET0131 ,
		\u1_u2_last_buf_adr_reg[5]/P0001 ,
		_w3536_
	);
	LUT3 #(
		.INIT('h70)
	) name1787 (
		_w3518_,
		_w3522_,
		_w3536_,
		_w3537_
	);
	LUT3 #(
		.INIT('h02)
	) name1788 (
		_w3533_,
		_w3535_,
		_w3537_,
		_w3538_
	);
	LUT2 #(
		.INIT('h8)
	) name1789 (
		\u1_u2_adr_cw_reg[5]/NET0131 ,
		\u1_u2_adr_cw_reg[6]/NET0131 ,
		_w3539_
	);
	LUT4 #(
		.INIT('h1555)
	) name1790 (
		\u1_u2_adr_cw_reg[7]/NET0131 ,
		_w3518_,
		_w3522_,
		_w3539_,
		_w3540_
	);
	LUT3 #(
		.INIT('h80)
	) name1791 (
		\u1_u2_adr_cw_reg[5]/NET0131 ,
		\u1_u2_adr_cw_reg[6]/NET0131 ,
		\u1_u2_adr_cw_reg[7]/NET0131 ,
		_w3541_
	);
	LUT4 #(
		.INIT('h1555)
	) name1792 (
		\u1_u2_last_buf_adr_reg[7]/P0001 ,
		_w3518_,
		_w3522_,
		_w3541_,
		_w3542_
	);
	LUT2 #(
		.INIT('h4)
	) name1793 (
		_w3540_,
		_w3542_,
		_w3543_
	);
	LUT4 #(
		.INIT('h0080)
	) name1794 (
		_w3526_,
		_w3532_,
		_w3538_,
		_w3543_,
		_w3544_
	);
	LUT2 #(
		.INIT('h4)
	) name1795 (
		\u1_u2_adr_cw_reg[7]/NET0131 ,
		\u1_u2_last_buf_adr_reg[7]/P0001 ,
		_w3545_
	);
	LUT4 #(
		.INIT('h7f00)
	) name1796 (
		_w3518_,
		_w3522_,
		_w3539_,
		_w3545_,
		_w3546_
	);
	LUT4 #(
		.INIT('h8000)
	) name1797 (
		\u1_u2_adr_cw_reg[5]/NET0131 ,
		\u1_u2_adr_cw_reg[6]/NET0131 ,
		\u1_u2_adr_cw_reg[7]/NET0131 ,
		\u1_u2_last_buf_adr_reg[7]/P0001 ,
		_w3547_
	);
	LUT3 #(
		.INIT('h80)
	) name1798 (
		_w3518_,
		_w3522_,
		_w3547_,
		_w3548_
	);
	LUT2 #(
		.INIT('h1)
	) name1799 (
		_w3546_,
		_w3548_,
		_w3549_
	);
	LUT4 #(
		.INIT('h963c)
	) name1800 (
		\u1_u2_adr_cw_reg[5]/NET0131 ,
		\u1_u2_adr_cw_reg[6]/NET0131 ,
		\u1_u2_last_buf_adr_reg[6]/P0001 ,
		_w3523_,
		_w3550_
	);
	LUT2 #(
		.INIT('h1)
	) name1801 (
		\u1_u2_adr_cw_reg[8]/P0001 ,
		\u1_u2_last_buf_adr_reg[8]/P0001 ,
		_w3551_
	);
	LUT4 #(
		.INIT('h7f00)
	) name1802 (
		_w3518_,
		_w3522_,
		_w3541_,
		_w3551_,
		_w3552_
	);
	LUT2 #(
		.INIT('h2)
	) name1803 (
		\u1_u2_adr_cw_reg[8]/P0001 ,
		\u1_u2_last_buf_adr_reg[8]/P0001 ,
		_w3553_
	);
	LUT4 #(
		.INIT('h8000)
	) name1804 (
		_w3518_,
		_w3522_,
		_w3541_,
		_w3553_,
		_w3554_
	);
	LUT2 #(
		.INIT('h8)
	) name1805 (
		\u1_u2_adr_cw_reg[8]/P0001 ,
		\u1_u2_last_buf_adr_reg[8]/P0001 ,
		_w3555_
	);
	LUT4 #(
		.INIT('h7f00)
	) name1806 (
		_w3518_,
		_w3522_,
		_w3541_,
		_w3555_,
		_w3556_
	);
	LUT2 #(
		.INIT('h4)
	) name1807 (
		\u1_u2_adr_cw_reg[8]/P0001 ,
		\u1_u2_last_buf_adr_reg[8]/P0001 ,
		_w3557_
	);
	LUT4 #(
		.INIT('h8000)
	) name1808 (
		_w3518_,
		_w3522_,
		_w3541_,
		_w3557_,
		_w3558_
	);
	LUT4 #(
		.INIT('h0001)
	) name1809 (
		_w3552_,
		_w3554_,
		_w3556_,
		_w3558_,
		_w3559_
	);
	LUT4 #(
		.INIT('h8000)
	) name1810 (
		\u1_u2_adr_cw_reg[5]/NET0131 ,
		\u1_u2_adr_cw_reg[6]/NET0131 ,
		\u1_u2_adr_cw_reg[7]/NET0131 ,
		\u1_u2_adr_cw_reg[8]/P0001 ,
		_w3560_
	);
	LUT3 #(
		.INIT('h80)
	) name1811 (
		_w3518_,
		_w3522_,
		_w3560_,
		_w3561_
	);
	LUT4 #(
		.INIT('h1555)
	) name1812 (
		\u1_u2_adr_cw_reg[9]/NET0131 ,
		_w3518_,
		_w3522_,
		_w3560_,
		_w3562_
	);
	LUT2 #(
		.INIT('h8)
	) name1813 (
		\u1_u2_adr_cw_reg[8]/P0001 ,
		\u1_u2_adr_cw_reg[9]/NET0131 ,
		_w3563_
	);
	LUT4 #(
		.INIT('h8000)
	) name1814 (
		_w3518_,
		_w3522_,
		_w3541_,
		_w3563_,
		_w3564_
	);
	LUT4 #(
		.INIT('h7b49)
	) name1815 (
		\u1_u2_adr_cw_reg[9]/NET0131 ,
		\u1_u2_last_buf_adr_reg[9]/P0001 ,
		_w3561_,
		_w3564_,
		_w3565_
	);
	LUT4 #(
		.INIT('h0200)
	) name1816 (
		_w3549_,
		_w3550_,
		_w3559_,
		_w3565_,
		_w3566_
	);
	LUT3 #(
		.INIT('h80)
	) name1817 (
		\u1_u2_adr_cw_reg[10]/P0001 ,
		\u1_u2_adr_cw_reg[8]/P0001 ,
		\u1_u2_adr_cw_reg[9]/NET0131 ,
		_w3567_
	);
	LUT4 #(
		.INIT('h8000)
	) name1818 (
		_w3518_,
		_w3522_,
		_w3541_,
		_w3567_,
		_w3568_
	);
	LUT2 #(
		.INIT('h8)
	) name1819 (
		\u1_u2_adr_cw_reg[11]/P0001 ,
		\u1_u2_adr_cw_reg[12]/P0001 ,
		_w3569_
	);
	LUT4 #(
		.INIT('h963c)
	) name1820 (
		\u1_u2_adr_cw_reg[11]/P0001 ,
		\u1_u2_adr_cw_reg[12]/P0001 ,
		\u1_u2_last_buf_adr_reg[12]/P0001 ,
		_w3568_,
		_w3570_
	);
	LUT4 #(
		.INIT('hecfd)
	) name1821 (
		\u1_u2_adr_cw_reg[11]/P0001 ,
		\u1_u2_last_buf_adr_reg[11]/P0001 ,
		_w3568_,
		_w3568_,
		_w3571_
	);
	LUT4 #(
		.INIT('hdcfe)
	) name1822 (
		\u1_u2_adr_cw_reg[10]/P0001 ,
		\u1_u2_last_buf_adr_reg[10]/P0001 ,
		_w3564_,
		_w3564_,
		_w3572_
	);
	LUT4 #(
		.INIT('h00c8)
	) name1823 (
		\u1_u2_adr_cw_reg[10]/P0001 ,
		\u1_u2_last_buf_adr_reg[10]/P0001 ,
		_w3564_,
		_w3568_,
		_w3573_
	);
	LUT4 #(
		.INIT('h73fb)
	) name1824 (
		\u1_u2_adr_cw_reg[11]/P0001 ,
		\u1_u2_last_buf_adr_reg[11]/P0001 ,
		_w3568_,
		_w3568_,
		_w3574_
	);
	LUT4 #(
		.INIT('ha200)
	) name1825 (
		_w3571_,
		_w3572_,
		_w3573_,
		_w3574_,
		_w3575_
	);
	LUT4 #(
		.INIT('h0800)
	) name1826 (
		_w3544_,
		_w3566_,
		_w3570_,
		_w3575_,
		_w3576_
	);
	LUT4 #(
		.INIT('h7bbb)
	) name1827 (
		\u1_u2_adr_cw_reg[13]/P0001 ,
		\u1_u2_last_buf_adr_reg[13]/P0001 ,
		_w3568_,
		_w3569_,
		_w3577_
	);
	LUT3 #(
		.INIT('h15)
	) name1828 (
		\u1_u2_adr_cw_reg[13]/P0001 ,
		_w3568_,
		_w3569_,
		_w3578_
	);
	LUT3 #(
		.INIT('h80)
	) name1829 (
		\u1_u2_adr_cw_reg[11]/P0001 ,
		\u1_u2_adr_cw_reg[12]/P0001 ,
		\u1_u2_adr_cw_reg[13]/P0001 ,
		_w3579_
	);
	LUT3 #(
		.INIT('h15)
	) name1830 (
		\u1_u2_last_buf_adr_reg[13]/P0001 ,
		_w3568_,
		_w3579_,
		_w3580_
	);
	LUT4 #(
		.INIT('h6999)
	) name1831 (
		\u1_u2_adr_cw_reg[14]/P0001 ,
		\u1_u2_last_buf_adr_reg[14]/P0001 ,
		_w3568_,
		_w3579_,
		_w3581_
	);
	LUT4 #(
		.INIT('h8a00)
	) name1832 (
		_w3577_,
		_w3578_,
		_w3580_,
		_w3581_,
		_w3582_
	);
	LUT3 #(
		.INIT('h9a)
	) name1833 (
		\u1_u2_adr_cw_reg[0]/NET0131 ,
		\u1_u2_dtmp_sel_r_reg/P0001 ,
		\u1_u2_mack_r_reg/P0001 ,
		_w3583_
	);
	LUT2 #(
		.INIT('h8)
	) name1834 (
		_w3185_,
		_w3583_,
		_w3584_
	);
	LUT4 #(
		.INIT('hbfaa)
	) name1835 (
		_w3188_,
		_w3576_,
		_w3582_,
		_w3584_,
		_w3585_
	);
	LUT3 #(
		.INIT('he0)
	) name1836 (
		\u1_u2_rx_dma_en_r_reg/P0001 ,
		\u1_u2_tx_dma_en_r_reg/P0001 ,
		\u1_u3_adr_reg[12]/P0001 ,
		_w3586_
	);
	LUT4 #(
		.INIT('h00c8)
	) name1837 (
		\u1_u2_adr_cw_reg[10]/P0001 ,
		_w3185_,
		_w3564_,
		_w3568_,
		_w3587_
	);
	LUT4 #(
		.INIT('hf7f0)
	) name1838 (
		_w3576_,
		_w3582_,
		_w3586_,
		_w3587_,
		_w3588_
	);
	LUT3 #(
		.INIT('he0)
	) name1839 (
		\u1_u2_rx_dma_en_r_reg/P0001 ,
		\u1_u2_tx_dma_en_r_reg/P0001 ,
		\u1_u3_adr_reg[13]/P0001 ,
		_w3589_
	);
	LUT3 #(
		.INIT('h48)
	) name1840 (
		\u1_u2_adr_cw_reg[11]/P0001 ,
		_w3185_,
		_w3568_,
		_w3590_
	);
	LUT4 #(
		.INIT('hf7f0)
	) name1841 (
		_w3576_,
		_w3582_,
		_w3589_,
		_w3590_,
		_w3591_
	);
	LUT3 #(
		.INIT('he0)
	) name1842 (
		\u1_u2_rx_dma_en_r_reg/P0001 ,
		\u1_u2_tx_dma_en_r_reg/P0001 ,
		\u1_u3_adr_reg[14]/P0001 ,
		_w3592_
	);
	LUT4 #(
		.INIT('h60c0)
	) name1843 (
		\u1_u2_adr_cw_reg[11]/P0001 ,
		\u1_u2_adr_cw_reg[12]/P0001 ,
		_w3185_,
		_w3568_,
		_w3593_
	);
	LUT4 #(
		.INIT('hf7f0)
	) name1844 (
		_w3576_,
		_w3582_,
		_w3592_,
		_w3593_,
		_w3594_
	);
	LUT3 #(
		.INIT('he0)
	) name1845 (
		\u1_u2_rx_dma_en_r_reg/P0001 ,
		\u1_u2_tx_dma_en_r_reg/P0001 ,
		\u1_u3_adr_reg[15]/P0001 ,
		_w3595_
	);
	LUT4 #(
		.INIT('h78f0)
	) name1846 (
		\u1_u2_adr_cw_reg[11]/P0001 ,
		\u1_u2_adr_cw_reg[12]/P0001 ,
		\u1_u2_adr_cw_reg[13]/P0001 ,
		_w3568_,
		_w3596_
	);
	LUT2 #(
		.INIT('h8)
	) name1847 (
		_w3185_,
		_w3596_,
		_w3597_
	);
	LUT4 #(
		.INIT('hf7f0)
	) name1848 (
		_w3576_,
		_w3582_,
		_w3595_,
		_w3597_,
		_w3598_
	);
	LUT3 #(
		.INIT('he0)
	) name1849 (
		\u1_u2_rx_dma_en_r_reg/P0001 ,
		\u1_u2_tx_dma_en_r_reg/P0001 ,
		\u1_u3_adr_reg[16]/P0001 ,
		_w3599_
	);
	LUT4 #(
		.INIT('h4888)
	) name1850 (
		\u1_u2_adr_cw_reg[14]/P0001 ,
		_w3185_,
		_w3568_,
		_w3579_,
		_w3600_
	);
	LUT4 #(
		.INIT('hf7f0)
	) name1851 (
		_w3576_,
		_w3582_,
		_w3599_,
		_w3600_,
		_w3601_
	);
	LUT3 #(
		.INIT('he0)
	) name1852 (
		\u1_u2_rx_dma_en_r_reg/P0001 ,
		\u1_u2_tx_dma_en_r_reg/P0001 ,
		\u1_u3_adr_reg[3]/P0001 ,
		_w3602_
	);
	LUT4 #(
		.INIT('hc6cc)
	) name1853 (
		\u1_u2_adr_cw_reg[0]/NET0131 ,
		\u1_u2_adr_cw_reg[1]/P0001 ,
		\u1_u2_dtmp_sel_r_reg/P0001 ,
		\u1_u2_mack_r_reg/P0001 ,
		_w3603_
	);
	LUT2 #(
		.INIT('h8)
	) name1854 (
		_w3185_,
		_w3603_,
		_w3604_
	);
	LUT4 #(
		.INIT('hf7f0)
	) name1855 (
		_w3576_,
		_w3582_,
		_w3602_,
		_w3604_,
		_w3605_
	);
	LUT3 #(
		.INIT('he0)
	) name1856 (
		\u1_u2_rx_dma_en_r_reg/P0001 ,
		\u1_u2_tx_dma_en_r_reg/P0001 ,
		\u1_u3_adr_reg[4]/P0001 ,
		_w3606_
	);
	LUT3 #(
		.INIT('h48)
	) name1857 (
		\u1_u2_adr_cw_reg[2]/P0001 ,
		_w3185_,
		_w3518_,
		_w3607_
	);
	LUT4 #(
		.INIT('hf7f0)
	) name1858 (
		_w3576_,
		_w3582_,
		_w3606_,
		_w3607_,
		_w3608_
	);
	LUT3 #(
		.INIT('he0)
	) name1859 (
		\u1_u2_rx_dma_en_r_reg/P0001 ,
		\u1_u2_tx_dma_en_r_reg/P0001 ,
		\u1_u3_adr_reg[5]/P0001 ,
		_w3609_
	);
	LUT4 #(
		.INIT('h60c0)
	) name1860 (
		\u1_u2_adr_cw_reg[2]/P0001 ,
		\u1_u2_adr_cw_reg[3]/NET0131 ,
		_w3185_,
		_w3518_,
		_w3610_
	);
	LUT4 #(
		.INIT('hf7f0)
	) name1861 (
		_w3576_,
		_w3582_,
		_w3609_,
		_w3610_,
		_w3611_
	);
	LUT3 #(
		.INIT('he0)
	) name1862 (
		\u1_u2_rx_dma_en_r_reg/P0001 ,
		\u1_u2_tx_dma_en_r_reg/P0001 ,
		\u1_u3_adr_reg[6]/P0001 ,
		_w3612_
	);
	LUT4 #(
		.INIT('h78f0)
	) name1863 (
		\u1_u2_adr_cw_reg[2]/P0001 ,
		\u1_u2_adr_cw_reg[3]/NET0131 ,
		\u1_u2_adr_cw_reg[4]/P0001 ,
		_w3518_,
		_w3613_
	);
	LUT2 #(
		.INIT('h8)
	) name1864 (
		_w3185_,
		_w3613_,
		_w3614_
	);
	LUT4 #(
		.INIT('hf7f0)
	) name1865 (
		_w3576_,
		_w3582_,
		_w3612_,
		_w3614_,
		_w3615_
	);
	LUT3 #(
		.INIT('he0)
	) name1866 (
		\u1_u2_rx_dma_en_r_reg/P0001 ,
		\u1_u2_tx_dma_en_r_reg/P0001 ,
		\u1_u3_adr_reg[7]/P0001 ,
		_w3616_
	);
	LUT4 #(
		.INIT('h4888)
	) name1867 (
		\u1_u2_adr_cw_reg[5]/NET0131 ,
		_w3185_,
		_w3518_,
		_w3522_,
		_w3617_
	);
	LUT4 #(
		.INIT('hf7f0)
	) name1868 (
		_w3576_,
		_w3582_,
		_w3616_,
		_w3617_,
		_w3618_
	);
	LUT3 #(
		.INIT('he0)
	) name1869 (
		\u1_u2_rx_dma_en_r_reg/P0001 ,
		\u1_u2_tx_dma_en_r_reg/P0001 ,
		\u1_u3_adr_reg[8]/P0001 ,
		_w3619_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name1870 (
		\u1_u2_adr_cw_reg[5]/NET0131 ,
		\u1_u2_adr_cw_reg[6]/NET0131 ,
		_w3518_,
		_w3522_,
		_w3620_
	);
	LUT2 #(
		.INIT('h8)
	) name1871 (
		_w3185_,
		_w3620_,
		_w3621_
	);
	LUT4 #(
		.INIT('hf7f0)
	) name1872 (
		_w3576_,
		_w3582_,
		_w3619_,
		_w3621_,
		_w3622_
	);
	LUT3 #(
		.INIT('he0)
	) name1873 (
		\u1_u2_rx_dma_en_r_reg/P0001 ,
		\u1_u2_tx_dma_en_r_reg/P0001 ,
		\u1_u3_adr_reg[9]/P0001 ,
		_w3623_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name1874 (
		\u1_u2_adr_cw_reg[7]/NET0131 ,
		_w3518_,
		_w3522_,
		_w3539_,
		_w3624_
	);
	LUT2 #(
		.INIT('h8)
	) name1875 (
		_w3185_,
		_w3624_,
		_w3625_
	);
	LUT4 #(
		.INIT('hf7f0)
	) name1876 (
		_w3576_,
		_w3582_,
		_w3623_,
		_w3625_,
		_w3626_
	);
	LUT3 #(
		.INIT('he0)
	) name1877 (
		\u1_u2_rx_dma_en_r_reg/P0001 ,
		\u1_u2_tx_dma_en_r_reg/P0001 ,
		\u1_u3_adr_reg[10]/P0001 ,
		_w3627_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name1878 (
		\u1_u2_adr_cw_reg[8]/P0001 ,
		_w3518_,
		_w3522_,
		_w3541_,
		_w3628_
	);
	LUT4 #(
		.INIT('h0080)
	) name1879 (
		\u1_u2_adr_cw_reg[5]/NET0131 ,
		\u1_u2_adr_cw_reg[6]/NET0131 ,
		\u1_u2_adr_cw_reg[7]/NET0131 ,
		\u1_u2_adr_cw_reg[8]/P0001 ,
		_w3629_
	);
	LUT3 #(
		.INIT('h80)
	) name1880 (
		_w3518_,
		_w3522_,
		_w3629_,
		_w3630_
	);
	LUT3 #(
		.INIT('ha8)
	) name1881 (
		_w3185_,
		_w3628_,
		_w3630_,
		_w3631_
	);
	LUT4 #(
		.INIT('hf7f0)
	) name1882 (
		_w3576_,
		_w3582_,
		_w3627_,
		_w3631_,
		_w3632_
	);
	LUT3 #(
		.INIT('he0)
	) name1883 (
		\u1_u2_rx_dma_en_r_reg/P0001 ,
		\u1_u2_tx_dma_en_r_reg/P0001 ,
		\u1_u3_adr_reg[11]/P0001 ,
		_w3633_
	);
	LUT3 #(
		.INIT('h02)
	) name1884 (
		_w3185_,
		_w3562_,
		_w3564_,
		_w3634_
	);
	LUT4 #(
		.INIT('hf7f0)
	) name1885 (
		_w3576_,
		_w3582_,
		_w3633_,
		_w3634_,
		_w3635_
	);
	LUT3 #(
		.INIT('ha6)
	) name1886 (
		\u1_u3_new_sizeb_reg[10]/P0001 ,
		_w2845_,
		_w2847_,
		_w3636_
	);
	LUT4 #(
		.INIT('h4fb0)
	) name1887 (
		_w3451_,
		_w3463_,
		_w3466_,
		_w3636_,
		_w3637_
	);
	LUT3 #(
		.INIT('h02)
	) name1888 (
		\u0_tx_ready_reg/NET0131 ,
		\u1_u1_state_reg[0]/NET0131 ,
		\u1_u1_state_reg[1]/NET0131 ,
		_w3638_
	);
	LUT3 #(
		.INIT('h2a)
	) name1889 (
		rst_i_pad,
		_w1809_,
		_w3638_,
		_w3639_
	);
	LUT4 #(
		.INIT('h0001)
	) name1890 (
		\u1_u1_send_zero_length_r_reg/P0001 ,
		\u1_u1_state_reg[2]/NET0131 ,
		\u1_u1_state_reg[3]/NET0131 ,
		\u1_u1_state_reg[4]/NET0131 ,
		_w3640_
	);
	LUT4 #(
		.INIT('h0004)
	) name1891 (
		\u1_u1_send_zero_length_r_reg/P0001 ,
		\u1_u1_state_reg[0]/NET0131 ,
		\u1_u1_state_reg[1]/NET0131 ,
		\u1_u2_send_data_r_reg/NET0131 ,
		_w3641_
	);
	LUT2 #(
		.INIT('h8)
	) name1892 (
		_w3640_,
		_w3641_,
		_w3642_
	);
	LUT2 #(
		.INIT('hd)
	) name1893 (
		_w3639_,
		_w3642_,
		_w3643_
	);
	LUT3 #(
		.INIT('h80)
	) name1894 (
		\u1_u1_send_zero_length_r_reg/P0001 ,
		_w1813_,
		_w3318_,
		_w3644_
	);
	LUT3 #(
		.INIT('h15)
	) name1895 (
		\u0_tx_ready_reg/NET0131 ,
		_w1806_,
		_w1809_,
		_w3645_
	);
	LUT3 #(
		.INIT('h2a)
	) name1896 (
		\u0_tx_ready_reg/NET0131 ,
		_w1807_,
		_w1815_,
		_w3646_
	);
	LUT3 #(
		.INIT('hf4)
	) name1897 (
		\u1_u1_send_data_r_reg/P0001 ,
		\u1_u1_send_zero_length_r_reg/P0001 ,
		\u1_u1_zero_length_r_reg/P0001 ,
		_w3647_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name1898 (
		rst_i_pad,
		\u1_u1_send_data_r_reg/P0001 ,
		\u1_u1_send_zero_length_r_reg/P0001 ,
		\u1_u2_send_data_r_reg/NET0131 ,
		_w3648_
	);
	LUT2 #(
		.INIT('h8)
	) name1899 (
		_w3647_,
		_w3648_,
		_w3649_
	);
	LUT3 #(
		.INIT('he0)
	) name1900 (
		_w3645_,
		_w3646_,
		_w3649_,
		_w3650_
	);
	LUT2 #(
		.INIT('h8)
	) name1901 (
		\u1_u3_out_to_small_r_reg/P0001 ,
		\u4_buf0_reg[0]/P0001 ,
		_w3651_
	);
	LUT2 #(
		.INIT('h6)
	) name1902 (
		\u1_u3_buffer_done_reg/P0001 ,
		\u4_csr_reg[30]/NET0131 ,
		_w3652_
	);
	LUT3 #(
		.INIT('h13)
	) name1903 (
		_w3488_,
		_w3651_,
		_w3652_,
		_w3653_
	);
	LUT2 #(
		.INIT('h1)
	) name1904 (
		_w3420_,
		_w3653_,
		_w3654_
	);
	LUT3 #(
		.INIT('h54)
	) name1905 (
		_w3093_,
		_w3149_,
		_w3150_,
		_w3655_
	);
	LUT2 #(
		.INIT('h1)
	) name1906 (
		\u1_u3_adr_r_reg[0]/P0001 ,
		_w3147_,
		_w3656_
	);
	LUT4 #(
		.INIT('h4044)
	) name1907 (
		_w3153_,
		_w3485_,
		_w3655_,
		_w3656_,
		_w3657_
	);
	LUT2 #(
		.INIT('he)
	) name1908 (
		_w3654_,
		_w3657_,
		_w3658_
	);
	LUT3 #(
		.INIT('h08)
	) name1909 (
		rst_i_pad,
		\u1_u2_rx_dma_en_r_reg/P0001 ,
		\u1_u3_abort_reg/P0001 ,
		_w3659_
	);
	LUT4 #(
		.INIT('h0800)
	) name1910 (
		_w3209_,
		_w3216_,
		_w3217_,
		_w3659_,
		_w3660_
	);
	LUT4 #(
		.INIT('h0020)
	) name1911 (
		rst_i_pad,
		\u1_u2_mack_r_reg/P0001 ,
		\u1_u2_state_reg[1]/NET0131 ,
		\u1_u3_abort_reg/P0001 ,
		_w3661_
	);
	LUT4 #(
		.INIT('hfdf0)
	) name1912 (
		_w3224_,
		_w3226_,
		_w3660_,
		_w3661_,
		_w3662_
	);
	LUT3 #(
		.INIT('hc4)
	) name1913 (
		\u1_u2_rx_dma_en_r_reg/P0001 ,
		\u1_u2_state_reg[5]/NET0131 ,
		\u1_u3_abort_reg/P0001 ,
		_w3663_
	);
	LUT4 #(
		.INIT('h8880)
	) name1914 (
		_w3209_,
		_w3216_,
		_w3217_,
		_w3663_,
		_w3664_
	);
	LUT4 #(
		.INIT('h0020)
	) name1915 (
		rst_i_pad,
		\u1_u2_mack_r_reg/P0001 ,
		\u1_u2_state_reg[5]/NET0131 ,
		\u1_u3_abort_reg/P0001 ,
		_w3665_
	);
	LUT4 #(
		.INIT('ha800)
	) name1916 (
		_w3205_,
		_w3222_,
		_w3223_,
		_w3665_,
		_w3666_
	);
	LUT3 #(
		.INIT('hf8)
	) name1917 (
		rst_i_pad,
		_w3664_,
		_w3666_,
		_w3667_
	);
	LUT2 #(
		.INIT('h4)
	) name1918 (
		\u1_u3_state_reg[2]/P0001 ,
		_w2127_,
		_w3668_
	);
	LUT2 #(
		.INIT('h1)
	) name1919 (
		\u1_u3_abort_reg/P0001 ,
		\u1_u3_tx_data_to_reg/P0001 ,
		_w3669_
	);
	LUT3 #(
		.INIT('h01)
	) name1920 (
		\u1_u3_abort_reg/P0001 ,
		\u1_u3_state_reg[0]/P0001 ,
		\u1_u3_tx_data_to_reg/P0001 ,
		_w3670_
	);
	LUT4 #(
		.INIT('h0100)
	) name1921 (
		\u1_u0_state_reg[0]/P0001 ,
		\u1_u0_state_reg[1]/P0001 ,
		\u1_u0_state_reg[2]/P0001 ,
		\u1_u0_state_reg[3]/P0001 ,
		_w3671_
	);
	LUT2 #(
		.INIT('h2)
	) name1922 (
		\u0_rx_active_reg/P0001 ,
		\u0_rx_err_reg/P0001 ,
		_w3672_
	);
	LUT4 #(
		.INIT('h000d)
	) name1923 (
		\u0_rx_active_reg/P0001 ,
		\u0_rx_err_reg/P0001 ,
		\u1_u3_abort_reg/P0001 ,
		\u1_u3_tx_data_to_reg/P0001 ,
		_w3673_
	);
	LUT3 #(
		.INIT('h15)
	) name1924 (
		_w3670_,
		_w3671_,
		_w3673_,
		_w3674_
	);
	LUT2 #(
		.INIT('h1)
	) name1925 (
		\u1_u3_state_reg[0]/P0001 ,
		\u1_u3_state_reg[1]/P0001 ,
		_w3675_
	);
	LUT4 #(
		.INIT('h0001)
	) name1926 (
		\u1_u3_state_reg[0]/P0001 ,
		\u1_u3_state_reg[1]/P0001 ,
		\u1_u3_state_reg[3]/P0001 ,
		\u1_u3_state_reg[5]/P0001 ,
		_w3676_
	);
	LUT2 #(
		.INIT('h8)
	) name1927 (
		\u1_u3_state_reg[4]/P0001 ,
		_w3676_,
		_w3677_
	);
	LUT4 #(
		.INIT('h0020)
	) name1928 (
		\u1_u0_crc16_sum_reg[0]/P0001 ,
		\u1_u0_crc16_sum_reg[14]/P0001 ,
		\u1_u0_crc16_sum_reg[15]/P0001 ,
		\u1_u0_crc16_sum_reg[1]/P0001 ,
		_w3678_
	);
	LUT4 #(
		.INIT('h0001)
	) name1929 (
		\u1_u0_crc16_sum_reg[10]/P0001 ,
		\u1_u0_crc16_sum_reg[11]/P0001 ,
		\u1_u0_crc16_sum_reg[12]/P0001 ,
		\u1_u0_crc16_sum_reg[13]/P0001 ,
		_w3679_
	);
	LUT4 #(
		.INIT('h0001)
	) name1930 (
		\u1_u0_crc16_sum_reg[6]/P0001 ,
		\u1_u0_crc16_sum_reg[7]/P0001 ,
		\u1_u0_crc16_sum_reg[8]/P0001 ,
		\u1_u0_crc16_sum_reg[9]/P0001 ,
		_w3680_
	);
	LUT4 #(
		.INIT('h0008)
	) name1931 (
		\u1_u0_crc16_sum_reg[2]/P0001 ,
		\u1_u0_crc16_sum_reg[3]/P0001 ,
		\u1_u0_crc16_sum_reg[4]/P0001 ,
		\u1_u0_crc16_sum_reg[5]/P0001 ,
		_w3681_
	);
	LUT4 #(
		.INIT('h8000)
	) name1932 (
		_w3678_,
		_w3679_,
		_w3680_,
		_w3681_,
		_w3682_
	);
	LUT2 #(
		.INIT('h2)
	) name1933 (
		_w3671_,
		_w3672_,
		_w3683_
	);
	LUT4 #(
		.INIT('h7377)
	) name1934 (
		_w3674_,
		_w3677_,
		_w3682_,
		_w3683_,
		_w3684_
	);
	LUT2 #(
		.INIT('h4)
	) name1935 (
		\u1_u3_state_reg[0]/P0001 ,
		\u1_u3_state_reg[1]/P0001 ,
		_w3685_
	);
	LUT3 #(
		.INIT('h80)
	) name1936 (
		_w2127_,
		_w2128_,
		_w3685_,
		_w3686_
	);
	LUT4 #(
		.INIT('h0001)
	) name1937 (
		\u1_u3_state_reg[0]/P0001 ,
		\u1_u3_state_reg[1]/P0001 ,
		\u1_u3_state_reg[6]/P0001 ,
		\u1_u3_state_reg[8]/P0001 ,
		_w3687_
	);
	LUT2 #(
		.INIT('h4)
	) name1938 (
		\u1_u3_state_reg[7]/P0001 ,
		\u1_u3_state_reg[9]/P0001 ,
		_w3688_
	);
	LUT3 #(
		.INIT('h80)
	) name1939 (
		_w2128_,
		_w3687_,
		_w3688_,
		_w3689_
	);
	LUT4 #(
		.INIT('h0001)
	) name1940 (
		\u1_u3_abort_reg/P0001 ,
		\u1_u3_pid_seq_err_reg/P0001 ,
		\u1_u3_to_large_reg/P0001 ,
		\u1_u3_to_small_reg/P0001 ,
		_w3690_
	);
	LUT4 #(
		.INIT('h0010)
	) name1941 (
		\u1_u3_state_reg[0]/P0001 ,
		\u1_u3_state_reg[1]/P0001 ,
		\u1_u3_state_reg[6]/P0001 ,
		\u1_u3_state_reg[8]/P0001 ,
		_w3691_
	);
	LUT4 #(
		.INIT('h0800)
	) name1942 (
		_w2126_,
		_w2128_,
		_w3690_,
		_w3691_,
		_w3692_
	);
	LUT3 #(
		.INIT('h01)
	) name1943 (
		_w3686_,
		_w3689_,
		_w3692_,
		_w3693_
	);
	LUT2 #(
		.INIT('h1)
	) name1944 (
		\u1_u3_rx_ack_to_reg/P0001 ,
		\u1_u3_state_reg[0]/P0001 ,
		_w3694_
	);
	LUT4 #(
		.INIT('h0004)
	) name1945 (
		\u1_u0_pid_reg[0]/NET0131 ,
		\u1_u0_pid_reg[1]/NET0131 ,
		\u1_u0_pid_reg[2]/NET0131 ,
		\u1_u0_pid_reg[3]/NET0131 ,
		_w3695_
	);
	LUT2 #(
		.INIT('h2)
	) name1946 (
		\u1_u0_token_valid_str1_reg/P0001 ,
		\u1_u3_rx_ack_to_reg/P0001 ,
		_w3696_
	);
	LUT3 #(
		.INIT('h15)
	) name1947 (
		_w3694_,
		_w3695_,
		_w3696_,
		_w3697_
	);
	LUT2 #(
		.INIT('h2)
	) name1948 (
		\u1_u3_state_reg[3]/P0001 ,
		\u1_u3_state_reg[5]/P0001 ,
		_w3698_
	);
	LUT4 #(
		.INIT('h0001)
	) name1949 (
		\u1_u3_state_reg[0]/P0001 ,
		\u1_u3_state_reg[1]/P0001 ,
		\u1_u3_state_reg[2]/P0001 ,
		\u1_u3_state_reg[4]/P0001 ,
		_w3699_
	);
	LUT3 #(
		.INIT('h80)
	) name1950 (
		_w2127_,
		_w3698_,
		_w3699_,
		_w3700_
	);
	LUT3 #(
		.INIT('h20)
	) name1951 (
		\u1_u3_abort_reg/P0001 ,
		\u1_u3_state_reg[3]/P0001 ,
		\u1_u3_state_reg[5]/P0001 ,
		_w3701_
	);
	LUT3 #(
		.INIT('h80)
	) name1952 (
		_w2127_,
		_w3699_,
		_w3701_,
		_w3702_
	);
	LUT3 #(
		.INIT('h07)
	) name1953 (
		_w3697_,
		_w3700_,
		_w3702_,
		_w3703_
	);
	LUT4 #(
		.INIT('hd000)
	) name1954 (
		_w3668_,
		_w3684_,
		_w3693_,
		_w3703_,
		_w3704_
	);
	LUT2 #(
		.INIT('h6)
	) name1955 (
		\u1_u0_token0_reg[2]/NET0131 ,
		\u4_funct_adr_reg[2]/P0001 ,
		_w3705_
	);
	LUT4 #(
		.INIT('hc400)
	) name1956 (
		\u1_u0_token0_reg[3]/NET0131 ,
		\u1_u0_token_valid_str1_reg/P0001 ,
		\u4_funct_adr_reg[3]/P0001 ,
		\u4_match_r1_reg/P0001 ,
		_w3706_
	);
	LUT4 #(
		.INIT('hfefb)
	) name1957 (
		\u1_u0_pid_reg[0]/NET0131 ,
		\u1_u0_pid_reg[1]/NET0131 ,
		\u1_u0_pid_reg[2]/NET0131 ,
		\u1_u0_pid_reg[3]/NET0131 ,
		_w3707_
	);
	LUT3 #(
		.INIT('h40)
	) name1958 (
		_w3705_,
		_w3706_,
		_w3707_,
		_w3708_
	);
	LUT2 #(
		.INIT('h9)
	) name1959 (
		\u1_u0_token0_reg[5]/NET0131 ,
		\u4_funct_adr_reg[5]/P0001 ,
		_w3709_
	);
	LUT4 #(
		.INIT('haf23)
	) name1960 (
		\u1_u0_token0_reg[0]/NET0131 ,
		\u1_u0_token0_reg[4]/P0001 ,
		\u4_funct_adr_reg[0]/P0001 ,
		\u4_funct_adr_reg[4]/P0001 ,
		_w3710_
	);
	LUT4 #(
		.INIT('h8421)
	) name1961 (
		\u1_u0_token0_reg[1]/P0001 ,
		\u1_u0_token0_reg[6]/P0001 ,
		\u4_funct_adr_reg[1]/P0001 ,
		\u4_funct_adr_reg[6]/P0001 ,
		_w3711_
	);
	LUT3 #(
		.INIT('h80)
	) name1962 (
		_w3709_,
		_w3710_,
		_w3711_,
		_w3712_
	);
	LUT2 #(
		.INIT('h2)
	) name1963 (
		\u1_u0_token0_reg[0]/NET0131 ,
		\u4_funct_adr_reg[0]/P0001 ,
		_w3713_
	);
	LUT4 #(
		.INIT('h8caf)
	) name1964 (
		\u1_u0_token0_reg[3]/NET0131 ,
		\u1_u0_token0_reg[4]/P0001 ,
		\u4_funct_adr_reg[3]/P0001 ,
		\u4_funct_adr_reg[4]/P0001 ,
		_w3714_
	);
	LUT4 #(
		.INIT('h0b00)
	) name1965 (
		\u0_u0_mode_hs_reg/P0001 ,
		_w2764_,
		_w3713_,
		_w3714_,
		_w3715_
	);
	LUT4 #(
		.INIT('h5440)
	) name1966 (
		\u1_u0_pid_reg[0]/NET0131 ,
		\u1_u0_pid_reg[1]/NET0131 ,
		\u1_u0_pid_reg[2]/NET0131 ,
		\u1_u0_pid_reg[3]/NET0131 ,
		_w3716_
	);
	LUT4 #(
		.INIT('h0080)
	) name1967 (
		_w3708_,
		_w3712_,
		_w3715_,
		_w3716_,
		_w3717_
	);
	LUT2 #(
		.INIT('h2)
	) name1968 (
		rst_i_pad,
		_w3717_,
		_w3718_
	);
	LUT2 #(
		.INIT('h2)
	) name1969 (
		\u1_u3_state_reg[0]/P0001 ,
		\u1_u3_state_reg[1]/P0001 ,
		_w3719_
	);
	LUT3 #(
		.INIT('h80)
	) name1970 (
		_w2127_,
		_w2128_,
		_w3719_,
		_w3720_
	);
	LUT4 #(
		.INIT('h2000)
	) name1971 (
		\u1_u0_pid_reg[0]/NET0131 ,
		\u1_u0_pid_reg[1]/NET0131 ,
		\u1_u0_pid_reg[2]/NET0131 ,
		\u1_u0_pid_reg[3]/NET0131 ,
		_w3721_
	);
	LUT4 #(
		.INIT('hdffd)
	) name1972 (
		\u1_u0_pid_reg[0]/NET0131 ,
		\u1_u0_pid_reg[1]/NET0131 ,
		\u1_u0_pid_reg[2]/NET0131 ,
		\u1_u0_pid_reg[3]/NET0131 ,
		_w3722_
	);
	LUT4 #(
		.INIT('h7677)
	) name1973 (
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		_w2115_,
		_w3722_,
		_w3723_
	);
	LUT2 #(
		.INIT('h1)
	) name1974 (
		_w2133_,
		_w3723_,
		_w3724_
	);
	LUT4 #(
		.INIT('hb030)
	) name1975 (
		_w2766_,
		_w2769_,
		_w3720_,
		_w3724_,
		_w3725_
	);
	LUT2 #(
		.INIT('h9)
	) name1976 (
		\u1_u0_token0_reg[7]/P0001 ,
		\u1_u0_token1_reg[2]/P0001 ,
		_w3726_
	);
	LUT3 #(
		.INIT('h96)
	) name1977 (
		\u1_u0_token0_reg[4]/P0001 ,
		\u1_u0_token1_reg[0]/P0001 ,
		\u1_u0_token1_reg[5]/P0001 ,
		_w3727_
	);
	LUT2 #(
		.INIT('h9)
	) name1978 (
		\u1_u0_token0_reg[0]/NET0131 ,
		\u1_u0_token0_reg[1]/P0001 ,
		_w3728_
	);
	LUT4 #(
		.INIT('h6996)
	) name1979 (
		\u1_u0_token0_reg[0]/NET0131 ,
		\u1_u0_token0_reg[1]/P0001 ,
		\u1_u0_token0_reg[2]/NET0131 ,
		\u1_u0_token0_reg[3]/NET0131 ,
		_w3729_
	);
	LUT3 #(
		.INIT('h09)
	) name1980 (
		_w3726_,
		_w3727_,
		_w3729_,
		_w3730_
	);
	LUT3 #(
		.INIT('h96)
	) name1981 (
		\u1_u0_token0_reg[0]/NET0131 ,
		\u1_u0_token0_reg[1]/P0001 ,
		\u1_u0_token0_reg[2]/NET0131 ,
		_w3731_
	);
	LUT2 #(
		.INIT('h6)
	) name1982 (
		\u1_u0_token0_reg[6]/P0001 ,
		\u1_u0_token1_reg[0]/P0001 ,
		_w3732_
	);
	LUT2 #(
		.INIT('h9)
	) name1983 (
		\u1_u0_token0_reg[5]/NET0131 ,
		\u1_u0_token1_reg[3]/P0001 ,
		_w3733_
	);
	LUT3 #(
		.INIT('hb7)
	) name1984 (
		_w3731_,
		_w3732_,
		_w3733_,
		_w3734_
	);
	LUT2 #(
		.INIT('h4)
	) name1985 (
		_w3730_,
		_w3734_,
		_w3735_
	);
	LUT4 #(
		.INIT('h9669)
	) name1986 (
		\u1_u0_token0_reg[6]/P0001 ,
		\u1_u0_token0_reg[7]/P0001 ,
		\u1_u0_token1_reg[1]/P0001 ,
		\u1_u0_token1_reg[4]/P0001 ,
		_w3736_
	);
	LUT2 #(
		.INIT('h2)
	) name1987 (
		_w3729_,
		_w3736_,
		_w3737_
	);
	LUT3 #(
		.INIT('hde)
	) name1988 (
		_w3731_,
		_w3732_,
		_w3733_,
		_w3738_
	);
	LUT2 #(
		.INIT('h4)
	) name1989 (
		_w3737_,
		_w3738_,
		_w3739_
	);
	LUT4 #(
		.INIT('h0400)
	) name1990 (
		_w3730_,
		_w3734_,
		_w3737_,
		_w3738_,
		_w3740_
	);
	LUT3 #(
		.INIT('h69)
	) name1991 (
		\u1_u0_token0_reg[4]/P0001 ,
		\u1_u0_token0_reg[7]/P0001 ,
		\u1_u0_token1_reg[2]/P0001 ,
		_w3741_
	);
	LUT2 #(
		.INIT('h9)
	) name1992 (
		\u1_u0_token0_reg[5]/NET0131 ,
		\u1_u0_token1_reg[7]/P0001 ,
		_w3742_
	);
	LUT3 #(
		.INIT('h69)
	) name1993 (
		_w3728_,
		_w3741_,
		_w3742_,
		_w3743_
	);
	LUT2 #(
		.INIT('h9)
	) name1994 (
		\u1_u0_token1_reg[1]/P0001 ,
		\u1_u0_token1_reg[6]/P0001 ,
		_w3744_
	);
	LUT4 #(
		.INIT('h9669)
	) name1995 (
		\u1_u0_token0_reg[0]/NET0131 ,
		\u1_u0_token0_reg[3]/NET0131 ,
		\u1_u0_token0_reg[4]/P0001 ,
		\u1_u0_token0_reg[6]/P0001 ,
		_w3745_
	);
	LUT2 #(
		.INIT('h6)
	) name1996 (
		_w3744_,
		_w3745_,
		_w3746_
	);
	LUT3 #(
		.INIT('h60)
	) name1997 (
		_w3726_,
		_w3727_,
		_w3736_,
		_w3747_
	);
	LUT3 #(
		.INIT('h01)
	) name1998 (
		_w3743_,
		_w3746_,
		_w3747_,
		_w3748_
	);
	LUT2 #(
		.INIT('h8)
	) name1999 (
		_w3740_,
		_w3748_,
		_w3749_
	);
	LUT2 #(
		.INIT('h8)
	) name2000 (
		rst_i_pad,
		\u1_u0_token_valid_str1_reg/P0001 ,
		_w3750_
	);
	LUT4 #(
		.INIT('hdcdd)
	) name2001 (
		_w3718_,
		_w3725_,
		_w3749_,
		_w3750_,
		_w3751_
	);
	LUT2 #(
		.INIT('hd)
	) name2002 (
		_w3704_,
		_w3751_,
		_w3752_
	);
	LUT4 #(
		.INIT('haa20)
	) name2003 (
		rst_i_pad,
		\u0_tx_ready_reg/NET0131 ,
		\u1_u1_send_token_r_reg/P0001 ,
		\u1_u3_send_token_reg/P0001 ,
		_w3753_
	);
	LUT3 #(
		.INIT('hfe)
	) name2004 (
		\u1_u1_send_zero_length_r_reg/P0001 ,
		\u1_u2_send_data_r_reg/NET0131 ,
		\u1_u3_send_token_reg/P0001 ,
		_w3754_
	);
	LUT4 #(
		.INIT('h8421)
	) name2005 (
		\u1_u0_token0_reg[7]/P0001 ,
		\u1_u0_token1_reg[1]/P0001 ,
		\u4_u0_csr1_reg[3]/P0001 ,
		\u4_u0_csr1_reg[5]/P0001 ,
		_w3755_
	);
	LUT4 #(
		.INIT('h8421)
	) name2006 (
		\u1_u0_token1_reg[0]/P0001 ,
		\u1_u0_token1_reg[2]/P0001 ,
		\u4_u0_csr1_reg[4]/P0001 ,
		\u4_u0_csr1_reg[6]/P0001 ,
		_w3756_
	);
	LUT2 #(
		.INIT('h8)
	) name2007 (
		_w3755_,
		_w3756_,
		_w3757_
	);
	LUT4 #(
		.INIT('h8421)
	) name2008 (
		\u1_u0_token0_reg[7]/P0001 ,
		\u1_u0_token1_reg[2]/P0001 ,
		\u4_u1_csr1_reg[3]/P0001 ,
		\u4_u1_csr1_reg[6]/P0001 ,
		_w3758_
	);
	LUT4 #(
		.INIT('h8421)
	) name2009 (
		\u1_u0_token1_reg[0]/P0001 ,
		\u1_u0_token1_reg[1]/P0001 ,
		\u4_u1_csr1_reg[4]/P0001 ,
		\u4_u1_csr1_reg[5]/P0001 ,
		_w3759_
	);
	LUT2 #(
		.INIT('h8)
	) name2010 (
		_w3758_,
		_w3759_,
		_w3760_
	);
	LUT4 #(
		.INIT('h0777)
	) name2011 (
		_w3755_,
		_w3756_,
		_w3758_,
		_w3759_,
		_w3761_
	);
	LUT4 #(
		.INIT('h8421)
	) name2012 (
		\u1_u0_token0_reg[7]/P0001 ,
		\u1_u0_token1_reg[2]/P0001 ,
		\u4_u2_csr1_reg[3]/P0001 ,
		\u4_u2_csr1_reg[6]/P0001 ,
		_w3762_
	);
	LUT4 #(
		.INIT('h8421)
	) name2013 (
		\u1_u0_token1_reg[0]/P0001 ,
		\u1_u0_token1_reg[1]/P0001 ,
		\u4_u2_csr1_reg[4]/P0001 ,
		\u4_u2_csr1_reg[5]/P0001 ,
		_w3763_
	);
	LUT2 #(
		.INIT('h8)
	) name2014 (
		_w3762_,
		_w3763_,
		_w3764_
	);
	LUT3 #(
		.INIT('h80)
	) name2015 (
		\u4_u2_dma_out_buf_avail_reg/P0001 ,
		_w3762_,
		_w3763_,
		_w3765_
	);
	LUT2 #(
		.INIT('h8)
	) name2016 (
		_w3761_,
		_w3765_,
		_w3766_
	);
	LUT3 #(
		.INIT('h80)
	) name2017 (
		\u4_u0_dma_out_buf_avail_reg/P0001 ,
		_w3755_,
		_w3756_,
		_w3767_
	);
	LUT4 #(
		.INIT('h7000)
	) name2018 (
		_w3755_,
		_w3756_,
		_w3758_,
		_w3759_,
		_w3768_
	);
	LUT3 #(
		.INIT('h13)
	) name2019 (
		\u4_u1_dma_out_buf_avail_reg/P0001 ,
		_w3767_,
		_w3768_,
		_w3769_
	);
	LUT4 #(
		.INIT('h8421)
	) name2020 (
		\u1_u0_token0_reg[7]/P0001 ,
		\u1_u0_token1_reg[2]/P0001 ,
		\u4_u3_csr1_reg[3]/P0001 ,
		\u4_u3_csr1_reg[6]/P0001 ,
		_w3770_
	);
	LUT4 #(
		.INIT('h8421)
	) name2021 (
		\u1_u0_token1_reg[0]/P0001 ,
		\u1_u0_token1_reg[1]/P0001 ,
		\u4_u3_csr1_reg[4]/P0001 ,
		\u4_u3_csr1_reg[5]/P0001 ,
		_w3771_
	);
	LUT2 #(
		.INIT('h8)
	) name2022 (
		_w3770_,
		_w3771_,
		_w3772_
	);
	LUT4 #(
		.INIT('h7000)
	) name2023 (
		_w3762_,
		_w3763_,
		_w3770_,
		_w3771_,
		_w3773_
	);
	LUT3 #(
		.INIT('h80)
	) name2024 (
		\u4_u3_dma_out_buf_avail_reg/P0001 ,
		_w3761_,
		_w3773_,
		_w3774_
	);
	LUT4 #(
		.INIT('h0777)
	) name2025 (
		_w3762_,
		_w3763_,
		_w3770_,
		_w3771_,
		_w3775_
	);
	LUT2 #(
		.INIT('h7)
	) name2026 (
		_w3761_,
		_w3775_,
		_w3776_
	);
	LUT3 #(
		.INIT('h80)
	) name2027 (
		\u4_dma_out_buf_avail_reg/P0001 ,
		_w3761_,
		_w3775_,
		_w3777_
	);
	LUT4 #(
		.INIT('hfffb)
	) name2028 (
		_w3766_,
		_w3769_,
		_w3774_,
		_w3777_,
		_w3778_
	);
	LUT2 #(
		.INIT('h2)
	) name2029 (
		\u4_u2_buf0_orig_m3_reg[11]/P0001 ,
		\u4_u2_dma_in_cnt_reg[11]/P0001 ,
		_w3779_
	);
	LUT4 #(
		.INIT('h8cef)
	) name2030 (
		\u4_u2_buf0_orig_m3_reg[10]/P0001 ,
		\u4_u2_buf0_orig_m3_reg[11]/P0001 ,
		\u4_u2_dma_in_cnt_reg[10]/P0001 ,
		\u4_u2_dma_in_cnt_reg[11]/P0001 ,
		_w3780_
	);
	LUT4 #(
		.INIT('hf531)
	) name2031 (
		\u4_u2_buf0_orig_m3_reg[10]/P0001 ,
		\u4_u2_buf0_orig_m3_reg[9]/P0001 ,
		\u4_u2_dma_in_cnt_reg[10]/P0001 ,
		\u4_u2_dma_in_cnt_reg[9]/P0001 ,
		_w3781_
	);
	LUT3 #(
		.INIT('h8c)
	) name2032 (
		_w3779_,
		_w3780_,
		_w3781_,
		_w3782_
	);
	LUT4 #(
		.INIT('hf531)
	) name2033 (
		\u4_u2_buf0_orig_m3_reg[7]/P0001 ,
		\u4_u2_buf0_orig_m3_reg[8]/P0001 ,
		\u4_u2_dma_in_cnt_reg[7]/P0001 ,
		\u4_u2_dma_in_cnt_reg[8]/P0001 ,
		_w3783_
	);
	LUT4 #(
		.INIT('h8caf)
	) name2034 (
		\u4_u2_buf0_orig_m3_reg[6]/P0001 ,
		\u4_u2_buf0_orig_m3_reg[7]/P0001 ,
		\u4_u2_dma_in_cnt_reg[6]/P0001 ,
		\u4_u2_dma_in_cnt_reg[7]/P0001 ,
		_w3784_
	);
	LUT2 #(
		.INIT('h2)
	) name2035 (
		_w3783_,
		_w3784_,
		_w3785_
	);
	LUT4 #(
		.INIT('h8caf)
	) name2036 (
		\u4_u2_buf0_orig_m3_reg[4]/P0001 ,
		\u4_u2_buf0_orig_m3_reg[5]/P0001 ,
		\u4_u2_dma_in_cnt_reg[4]/P0001 ,
		\u4_u2_dma_in_cnt_reg[5]/P0001 ,
		_w3786_
	);
	LUT4 #(
		.INIT('hf531)
	) name2037 (
		\u4_u2_buf0_orig_m3_reg[3]/P0001 ,
		\u4_u2_buf0_orig_m3_reg[4]/P0001 ,
		\u4_u2_dma_in_cnt_reg[3]/P0001 ,
		\u4_u2_dma_in_cnt_reg[4]/P0001 ,
		_w3787_
	);
	LUT2 #(
		.INIT('h2)
	) name2038 (
		_w3786_,
		_w3787_,
		_w3788_
	);
	LUT4 #(
		.INIT('h080a)
	) name2039 (
		\u4_u2_buf0_orig_m3_reg[0]/P0001 ,
		\u4_u2_buf0_orig_m3_reg[1]/P0001 ,
		\u4_u2_dma_in_cnt_reg[0]/P0001 ,
		\u4_u2_dma_in_cnt_reg[1]/P0001 ,
		_w3789_
	);
	LUT4 #(
		.INIT('hf531)
	) name2040 (
		\u4_u2_buf0_orig_m3_reg[1]/P0001 ,
		\u4_u2_buf0_orig_m3_reg[2]/P0001 ,
		\u4_u2_dma_in_cnt_reg[1]/P0001 ,
		\u4_u2_dma_in_cnt_reg[2]/P0001 ,
		_w3790_
	);
	LUT4 #(
		.INIT('h8caf)
	) name2041 (
		\u4_u2_buf0_orig_m3_reg[2]/P0001 ,
		\u4_u2_buf0_orig_m3_reg[3]/P0001 ,
		\u4_u2_dma_in_cnt_reg[2]/P0001 ,
		\u4_u2_dma_in_cnt_reg[3]/P0001 ,
		_w3791_
	);
	LUT4 #(
		.INIT('h8a00)
	) name2042 (
		_w3786_,
		_w3789_,
		_w3790_,
		_w3791_,
		_w3792_
	);
	LUT4 #(
		.INIT('hf531)
	) name2043 (
		\u4_u2_buf0_orig_m3_reg[5]/P0001 ,
		\u4_u2_buf0_orig_m3_reg[6]/P0001 ,
		\u4_u2_dma_in_cnt_reg[5]/P0001 ,
		\u4_u2_dma_in_cnt_reg[6]/P0001 ,
		_w3793_
	);
	LUT2 #(
		.INIT('h8)
	) name2044 (
		_w3783_,
		_w3793_,
		_w3794_
	);
	LUT4 #(
		.INIT('h5455)
	) name2045 (
		_w3785_,
		_w3788_,
		_w3792_,
		_w3794_,
		_w3795_
	);
	LUT4 #(
		.INIT('h8caf)
	) name2046 (
		\u4_u2_buf0_orig_m3_reg[8]/P0001 ,
		\u4_u2_buf0_orig_m3_reg[9]/P0001 ,
		\u4_u2_dma_in_cnt_reg[8]/P0001 ,
		\u4_u2_dma_in_cnt_reg[9]/P0001 ,
		_w3796_
	);
	LUT2 #(
		.INIT('h8)
	) name2047 (
		_w3780_,
		_w3796_,
		_w3797_
	);
	LUT3 #(
		.INIT('hea)
	) name2048 (
		_w3782_,
		_w3795_,
		_w3797_,
		_w3798_
	);
	LUT2 #(
		.INIT('h2)
	) name2049 (
		\u4_u3_buf0_orig_m3_reg[11]/P0001 ,
		\u4_u3_dma_in_cnt_reg[11]/P0001 ,
		_w3799_
	);
	LUT4 #(
		.INIT('h8cef)
	) name2050 (
		\u4_u3_buf0_orig_m3_reg[10]/P0001 ,
		\u4_u3_buf0_orig_m3_reg[11]/P0001 ,
		\u4_u3_dma_in_cnt_reg[10]/P0001 ,
		\u4_u3_dma_in_cnt_reg[11]/P0001 ,
		_w3800_
	);
	LUT4 #(
		.INIT('hf531)
	) name2051 (
		\u4_u3_buf0_orig_m3_reg[10]/P0001 ,
		\u4_u3_buf0_orig_m3_reg[9]/P0001 ,
		\u4_u3_dma_in_cnt_reg[10]/P0001 ,
		\u4_u3_dma_in_cnt_reg[9]/P0001 ,
		_w3801_
	);
	LUT3 #(
		.INIT('h8c)
	) name2052 (
		_w3799_,
		_w3800_,
		_w3801_,
		_w3802_
	);
	LUT4 #(
		.INIT('hf531)
	) name2053 (
		\u4_u3_buf0_orig_m3_reg[7]/P0001 ,
		\u4_u3_buf0_orig_m3_reg[8]/P0001 ,
		\u4_u3_dma_in_cnt_reg[7]/P0001 ,
		\u4_u3_dma_in_cnt_reg[8]/P0001 ,
		_w3803_
	);
	LUT4 #(
		.INIT('h8caf)
	) name2054 (
		\u4_u3_buf0_orig_m3_reg[6]/P0001 ,
		\u4_u3_buf0_orig_m3_reg[7]/P0001 ,
		\u4_u3_dma_in_cnt_reg[6]/P0001 ,
		\u4_u3_dma_in_cnt_reg[7]/P0001 ,
		_w3804_
	);
	LUT2 #(
		.INIT('h2)
	) name2055 (
		_w3803_,
		_w3804_,
		_w3805_
	);
	LUT4 #(
		.INIT('h8caf)
	) name2056 (
		\u4_u3_buf0_orig_m3_reg[4]/P0001 ,
		\u4_u3_buf0_orig_m3_reg[5]/P0001 ,
		\u4_u3_dma_in_cnt_reg[4]/P0001 ,
		\u4_u3_dma_in_cnt_reg[5]/P0001 ,
		_w3806_
	);
	LUT4 #(
		.INIT('hf531)
	) name2057 (
		\u4_u3_buf0_orig_m3_reg[3]/P0001 ,
		\u4_u3_buf0_orig_m3_reg[4]/P0001 ,
		\u4_u3_dma_in_cnt_reg[3]/P0001 ,
		\u4_u3_dma_in_cnt_reg[4]/P0001 ,
		_w3807_
	);
	LUT2 #(
		.INIT('h2)
	) name2058 (
		_w3806_,
		_w3807_,
		_w3808_
	);
	LUT4 #(
		.INIT('h080a)
	) name2059 (
		\u4_u3_buf0_orig_m3_reg[0]/P0001 ,
		\u4_u3_buf0_orig_m3_reg[1]/P0001 ,
		\u4_u3_dma_in_cnt_reg[0]/P0001 ,
		\u4_u3_dma_in_cnt_reg[1]/P0001 ,
		_w3809_
	);
	LUT4 #(
		.INIT('hf531)
	) name2060 (
		\u4_u3_buf0_orig_m3_reg[1]/P0001 ,
		\u4_u3_buf0_orig_m3_reg[2]/P0001 ,
		\u4_u3_dma_in_cnt_reg[1]/P0001 ,
		\u4_u3_dma_in_cnt_reg[2]/P0001 ,
		_w3810_
	);
	LUT4 #(
		.INIT('h8caf)
	) name2061 (
		\u4_u3_buf0_orig_m3_reg[2]/P0001 ,
		\u4_u3_buf0_orig_m3_reg[3]/P0001 ,
		\u4_u3_dma_in_cnt_reg[2]/P0001 ,
		\u4_u3_dma_in_cnt_reg[3]/P0001 ,
		_w3811_
	);
	LUT4 #(
		.INIT('h8a00)
	) name2062 (
		_w3806_,
		_w3809_,
		_w3810_,
		_w3811_,
		_w3812_
	);
	LUT4 #(
		.INIT('hf531)
	) name2063 (
		\u4_u3_buf0_orig_m3_reg[5]/P0001 ,
		\u4_u3_buf0_orig_m3_reg[6]/P0001 ,
		\u4_u3_dma_in_cnt_reg[5]/P0001 ,
		\u4_u3_dma_in_cnt_reg[6]/P0001 ,
		_w3813_
	);
	LUT2 #(
		.INIT('h8)
	) name2064 (
		_w3803_,
		_w3813_,
		_w3814_
	);
	LUT4 #(
		.INIT('h5455)
	) name2065 (
		_w3805_,
		_w3808_,
		_w3812_,
		_w3814_,
		_w3815_
	);
	LUT4 #(
		.INIT('h8caf)
	) name2066 (
		\u4_u3_buf0_orig_m3_reg[8]/P0001 ,
		\u4_u3_buf0_orig_m3_reg[9]/P0001 ,
		\u4_u3_dma_in_cnt_reg[8]/P0001 ,
		\u4_u3_dma_in_cnt_reg[9]/P0001 ,
		_w3816_
	);
	LUT2 #(
		.INIT('h8)
	) name2067 (
		_w3800_,
		_w3816_,
		_w3817_
	);
	LUT3 #(
		.INIT('hea)
	) name2068 (
		_w3802_,
		_w3815_,
		_w3817_,
		_w3818_
	);
	LUT2 #(
		.INIT('h2)
	) name2069 (
		\u4_u0_buf0_orig_m3_reg[11]/P0001 ,
		\u4_u0_dma_in_cnt_reg[11]/P0001 ,
		_w3819_
	);
	LUT4 #(
		.INIT('h8cef)
	) name2070 (
		\u4_u0_buf0_orig_m3_reg[10]/P0001 ,
		\u4_u0_buf0_orig_m3_reg[11]/P0001 ,
		\u4_u0_dma_in_cnt_reg[10]/P0001 ,
		\u4_u0_dma_in_cnt_reg[11]/P0001 ,
		_w3820_
	);
	LUT4 #(
		.INIT('hf531)
	) name2071 (
		\u4_u0_buf0_orig_m3_reg[10]/P0001 ,
		\u4_u0_buf0_orig_m3_reg[9]/P0001 ,
		\u4_u0_dma_in_cnt_reg[10]/P0001 ,
		\u4_u0_dma_in_cnt_reg[9]/P0001 ,
		_w3821_
	);
	LUT3 #(
		.INIT('h8c)
	) name2072 (
		_w3819_,
		_w3820_,
		_w3821_,
		_w3822_
	);
	LUT4 #(
		.INIT('hf531)
	) name2073 (
		\u4_u0_buf0_orig_m3_reg[7]/P0001 ,
		\u4_u0_buf0_orig_m3_reg[8]/P0001 ,
		\u4_u0_dma_in_cnt_reg[7]/P0001 ,
		\u4_u0_dma_in_cnt_reg[8]/P0001 ,
		_w3823_
	);
	LUT4 #(
		.INIT('h8caf)
	) name2074 (
		\u4_u0_buf0_orig_m3_reg[6]/P0001 ,
		\u4_u0_buf0_orig_m3_reg[7]/P0001 ,
		\u4_u0_dma_in_cnt_reg[6]/P0001 ,
		\u4_u0_dma_in_cnt_reg[7]/P0001 ,
		_w3824_
	);
	LUT2 #(
		.INIT('h2)
	) name2075 (
		_w3823_,
		_w3824_,
		_w3825_
	);
	LUT4 #(
		.INIT('h8caf)
	) name2076 (
		\u4_u0_buf0_orig_m3_reg[4]/P0001 ,
		\u4_u0_buf0_orig_m3_reg[5]/P0001 ,
		\u4_u0_dma_in_cnt_reg[4]/P0001 ,
		\u4_u0_dma_in_cnt_reg[5]/P0001 ,
		_w3826_
	);
	LUT4 #(
		.INIT('hf531)
	) name2077 (
		\u4_u0_buf0_orig_m3_reg[3]/P0001 ,
		\u4_u0_buf0_orig_m3_reg[4]/P0001 ,
		\u4_u0_dma_in_cnt_reg[3]/P0001 ,
		\u4_u0_dma_in_cnt_reg[4]/P0001 ,
		_w3827_
	);
	LUT2 #(
		.INIT('h2)
	) name2078 (
		_w3826_,
		_w3827_,
		_w3828_
	);
	LUT4 #(
		.INIT('h080a)
	) name2079 (
		\u4_u0_buf0_orig_m3_reg[0]/P0001 ,
		\u4_u0_buf0_orig_m3_reg[1]/P0001 ,
		\u4_u0_dma_in_cnt_reg[0]/P0001 ,
		\u4_u0_dma_in_cnt_reg[1]/P0001 ,
		_w3829_
	);
	LUT4 #(
		.INIT('hf531)
	) name2080 (
		\u4_u0_buf0_orig_m3_reg[1]/P0001 ,
		\u4_u0_buf0_orig_m3_reg[2]/P0001 ,
		\u4_u0_dma_in_cnt_reg[1]/P0001 ,
		\u4_u0_dma_in_cnt_reg[2]/P0001 ,
		_w3830_
	);
	LUT4 #(
		.INIT('h8caf)
	) name2081 (
		\u4_u0_buf0_orig_m3_reg[2]/P0001 ,
		\u4_u0_buf0_orig_m3_reg[3]/P0001 ,
		\u4_u0_dma_in_cnt_reg[2]/P0001 ,
		\u4_u0_dma_in_cnt_reg[3]/P0001 ,
		_w3831_
	);
	LUT4 #(
		.INIT('h8a00)
	) name2082 (
		_w3826_,
		_w3829_,
		_w3830_,
		_w3831_,
		_w3832_
	);
	LUT4 #(
		.INIT('hf531)
	) name2083 (
		\u4_u0_buf0_orig_m3_reg[5]/P0001 ,
		\u4_u0_buf0_orig_m3_reg[6]/P0001 ,
		\u4_u0_dma_in_cnt_reg[5]/P0001 ,
		\u4_u0_dma_in_cnt_reg[6]/P0001 ,
		_w3833_
	);
	LUT2 #(
		.INIT('h8)
	) name2084 (
		_w3823_,
		_w3833_,
		_w3834_
	);
	LUT4 #(
		.INIT('h5455)
	) name2085 (
		_w3825_,
		_w3828_,
		_w3832_,
		_w3834_,
		_w3835_
	);
	LUT4 #(
		.INIT('h8caf)
	) name2086 (
		\u4_u0_buf0_orig_m3_reg[8]/P0001 ,
		\u4_u0_buf0_orig_m3_reg[9]/P0001 ,
		\u4_u0_dma_in_cnt_reg[8]/P0001 ,
		\u4_u0_dma_in_cnt_reg[9]/P0001 ,
		_w3836_
	);
	LUT2 #(
		.INIT('h8)
	) name2087 (
		_w3820_,
		_w3836_,
		_w3837_
	);
	LUT3 #(
		.INIT('hea)
	) name2088 (
		_w3822_,
		_w3835_,
		_w3837_,
		_w3838_
	);
	LUT2 #(
		.INIT('h2)
	) name2089 (
		\u4_u1_buf0_orig_m3_reg[11]/P0001 ,
		\u4_u1_dma_in_cnt_reg[11]/P0001 ,
		_w3839_
	);
	LUT4 #(
		.INIT('h8cef)
	) name2090 (
		\u4_u1_buf0_orig_m3_reg[10]/P0001 ,
		\u4_u1_buf0_orig_m3_reg[11]/P0001 ,
		\u4_u1_dma_in_cnt_reg[10]/P0001 ,
		\u4_u1_dma_in_cnt_reg[11]/P0001 ,
		_w3840_
	);
	LUT4 #(
		.INIT('hf531)
	) name2091 (
		\u4_u1_buf0_orig_m3_reg[10]/P0001 ,
		\u4_u1_buf0_orig_m3_reg[9]/P0001 ,
		\u4_u1_dma_in_cnt_reg[10]/P0001 ,
		\u4_u1_dma_in_cnt_reg[9]/P0001 ,
		_w3841_
	);
	LUT3 #(
		.INIT('h8c)
	) name2092 (
		_w3839_,
		_w3840_,
		_w3841_,
		_w3842_
	);
	LUT4 #(
		.INIT('hf531)
	) name2093 (
		\u4_u1_buf0_orig_m3_reg[7]/P0001 ,
		\u4_u1_buf0_orig_m3_reg[8]/P0001 ,
		\u4_u1_dma_in_cnt_reg[7]/P0001 ,
		\u4_u1_dma_in_cnt_reg[8]/P0001 ,
		_w3843_
	);
	LUT4 #(
		.INIT('h8caf)
	) name2094 (
		\u4_u1_buf0_orig_m3_reg[6]/P0001 ,
		\u4_u1_buf0_orig_m3_reg[7]/P0001 ,
		\u4_u1_dma_in_cnt_reg[6]/P0001 ,
		\u4_u1_dma_in_cnt_reg[7]/P0001 ,
		_w3844_
	);
	LUT2 #(
		.INIT('h2)
	) name2095 (
		_w3843_,
		_w3844_,
		_w3845_
	);
	LUT4 #(
		.INIT('h8caf)
	) name2096 (
		\u4_u1_buf0_orig_m3_reg[4]/P0001 ,
		\u4_u1_buf0_orig_m3_reg[5]/P0001 ,
		\u4_u1_dma_in_cnt_reg[4]/P0001 ,
		\u4_u1_dma_in_cnt_reg[5]/P0001 ,
		_w3846_
	);
	LUT4 #(
		.INIT('hf531)
	) name2097 (
		\u4_u1_buf0_orig_m3_reg[3]/P0001 ,
		\u4_u1_buf0_orig_m3_reg[4]/P0001 ,
		\u4_u1_dma_in_cnt_reg[3]/P0001 ,
		\u4_u1_dma_in_cnt_reg[4]/P0001 ,
		_w3847_
	);
	LUT2 #(
		.INIT('h2)
	) name2098 (
		_w3846_,
		_w3847_,
		_w3848_
	);
	LUT4 #(
		.INIT('h080a)
	) name2099 (
		\u4_u1_buf0_orig_m3_reg[0]/P0001 ,
		\u4_u1_buf0_orig_m3_reg[1]/P0001 ,
		\u4_u1_dma_in_cnt_reg[0]/P0001 ,
		\u4_u1_dma_in_cnt_reg[1]/P0001 ,
		_w3849_
	);
	LUT4 #(
		.INIT('hf531)
	) name2100 (
		\u4_u1_buf0_orig_m3_reg[1]/P0001 ,
		\u4_u1_buf0_orig_m3_reg[2]/P0001 ,
		\u4_u1_dma_in_cnt_reg[1]/P0001 ,
		\u4_u1_dma_in_cnt_reg[2]/P0001 ,
		_w3850_
	);
	LUT4 #(
		.INIT('h8caf)
	) name2101 (
		\u4_u1_buf0_orig_m3_reg[2]/P0001 ,
		\u4_u1_buf0_orig_m3_reg[3]/P0001 ,
		\u4_u1_dma_in_cnt_reg[2]/P0001 ,
		\u4_u1_dma_in_cnt_reg[3]/P0001 ,
		_w3851_
	);
	LUT4 #(
		.INIT('h8a00)
	) name2102 (
		_w3846_,
		_w3849_,
		_w3850_,
		_w3851_,
		_w3852_
	);
	LUT4 #(
		.INIT('hf531)
	) name2103 (
		\u4_u1_buf0_orig_m3_reg[5]/P0001 ,
		\u4_u1_buf0_orig_m3_reg[6]/P0001 ,
		\u4_u1_dma_in_cnt_reg[5]/P0001 ,
		\u4_u1_dma_in_cnt_reg[6]/P0001 ,
		_w3853_
	);
	LUT2 #(
		.INIT('h8)
	) name2104 (
		_w3843_,
		_w3853_,
		_w3854_
	);
	LUT4 #(
		.INIT('h5455)
	) name2105 (
		_w3845_,
		_w3848_,
		_w3852_,
		_w3854_,
		_w3855_
	);
	LUT4 #(
		.INIT('h8caf)
	) name2106 (
		\u4_u1_buf0_orig_m3_reg[8]/P0001 ,
		\u4_u1_buf0_orig_m3_reg[9]/P0001 ,
		\u4_u1_dma_in_cnt_reg[8]/P0001 ,
		\u4_u1_dma_in_cnt_reg[9]/P0001 ,
		_w3856_
	);
	LUT2 #(
		.INIT('h8)
	) name2107 (
		_w3840_,
		_w3856_,
		_w3857_
	);
	LUT3 #(
		.INIT('hea)
	) name2108 (
		_w3842_,
		_w3855_,
		_w3857_,
		_w3858_
	);
	LUT3 #(
		.INIT('h70)
	) name2109 (
		_w3740_,
		_w3748_,
		_w3750_,
		_w3859_
	);
	LUT2 #(
		.INIT('h1)
	) name2110 (
		_w3718_,
		_w3859_,
		_w3860_
	);
	LUT2 #(
		.INIT('h2)
	) name2111 (
		\u1_u3_state_reg[2]/P0001 ,
		\u1_u3_state_reg[4]/P0001 ,
		_w3861_
	);
	LUT4 #(
		.INIT('h4000)
	) name2112 (
		\u1_u2_idma_done_reg/P0001 ,
		_w2127_,
		_w3676_,
		_w3861_,
		_w3862_
	);
	LUT3 #(
		.INIT('h80)
	) name2113 (
		_w2766_,
		_w2772_,
		_w3720_,
		_w3863_
	);
	LUT2 #(
		.INIT('h4)
	) name2114 (
		\u4_csr_reg[27]/NET0131 ,
		_w3722_,
		_w3864_
	);
	LUT4 #(
		.INIT('h0b0a)
	) name2115 (
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		_w2133_,
		_w3722_,
		_w3865_
	);
	LUT4 #(
		.INIT('h8000)
	) name2116 (
		\u1_u3_state_reg[2]/P0001 ,
		_w2127_,
		_w2128_,
		_w3719_,
		_w3866_
	);
	LUT4 #(
		.INIT('hb300)
	) name2117 (
		_w2766_,
		_w2769_,
		_w3865_,
		_w3866_,
		_w3867_
	);
	LUT3 #(
		.INIT('h01)
	) name2118 (
		_w3862_,
		_w3863_,
		_w3867_,
		_w3868_
	);
	LUT2 #(
		.INIT('h1)
	) name2119 (
		_w3860_,
		_w3868_,
		_w3869_
	);
	LUT4 #(
		.INIT('h00cd)
	) name2120 (
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		_w2115_,
		_w2133_,
		_w3870_
	);
	LUT4 #(
		.INIT('h00a2)
	) name2121 (
		\u1_u3_match_r_reg/P0001 ,
		\u4_csr_reg[22]/P0001 ,
		\u4_csr_reg[23]/P0001 ,
		\u4_csr_reg[26]/NET0131 ,
		_w3871_
	);
	LUT3 #(
		.INIT('h45)
	) name2122 (
		\u1_u3_state_reg[4]/P0001 ,
		_w2131_,
		_w3871_,
		_w3872_
	);
	LUT2 #(
		.INIT('h1)
	) name2123 (
		\u1_u3_state_reg[4]/P0001 ,
		\u4_csr_reg[27]/NET0131 ,
		_w3873_
	);
	LUT2 #(
		.INIT('h8)
	) name2124 (
		_w3722_,
		_w3873_,
		_w3874_
	);
	LUT3 #(
		.INIT('h02)
	) name2125 (
		_w3720_,
		_w3872_,
		_w3874_,
		_w3875_
	);
	LUT4 #(
		.INIT('hb300)
	) name2126 (
		_w2766_,
		_w2769_,
		_w3870_,
		_w3875_,
		_w3876_
	);
	LUT4 #(
		.INIT('h4000)
	) name2127 (
		\u1_u3_state_reg[2]/P0001 ,
		\u1_u3_state_reg[4]/P0001 ,
		_w2127_,
		_w3676_,
		_w3877_
	);
	LUT4 #(
		.INIT('h8a00)
	) name2128 (
		_w3669_,
		_w3682_,
		_w3683_,
		_w3877_,
		_w3878_
	);
	LUT3 #(
		.INIT('ha2)
	) name2129 (
		\u1_u3_state_reg[4]/P0001 ,
		_w3671_,
		_w3672_,
		_w3879_
	);
	LUT2 #(
		.INIT('h8)
	) name2130 (
		_w3878_,
		_w3879_,
		_w3880_
	);
	LUT4 #(
		.INIT('heee0)
	) name2131 (
		_w3718_,
		_w3859_,
		_w3876_,
		_w3880_,
		_w3881_
	);
	LUT2 #(
		.INIT('h2)
	) name2132 (
		\u1_u3_state_reg[1]/P0001 ,
		_w3723_,
		_w3882_
	);
	LUT2 #(
		.INIT('h8)
	) name2133 (
		_w2769_,
		_w3720_,
		_w3883_
	);
	LUT4 #(
		.INIT('hfb00)
	) name2134 (
		_w2133_,
		_w2766_,
		_w3882_,
		_w3883_,
		_w3884_
	);
	LUT4 #(
		.INIT('hba00)
	) name2135 (
		_w3718_,
		_w3749_,
		_w3750_,
		_w3884_,
		_w3885_
	);
	LUT2 #(
		.INIT('h1)
	) name2136 (
		_w2151_,
		_w2152_,
		_w3886_
	);
	LUT2 #(
		.INIT('h8)
	) name2137 (
		_w2132_,
		_w2134_,
		_w3887_
	);
	LUT3 #(
		.INIT('h73)
	) name2138 (
		_w2766_,
		_w3886_,
		_w3887_,
		_w3888_
	);
	LUT3 #(
		.INIT('h07)
	) name2139 (
		\u1_u3_int_upid_set_reg/P0001 ,
		\u4_u2_ep_match_r_reg/P0001 ,
		\u4_u2_int_stat_reg[2]/P0001 ,
		_w3889_
	);
	LUT2 #(
		.INIT('h2)
	) name2140 (
		rst_i_pad,
		\u4_u2_int_re_reg/P0001 ,
		_w3890_
	);
	LUT2 #(
		.INIT('h4)
	) name2141 (
		_w3889_,
		_w3890_,
		_w3891_
	);
	LUT3 #(
		.INIT('h07)
	) name2142 (
		\u1_u3_int_upid_set_reg/P0001 ,
		\u4_u3_ep_match_r_reg/P0001 ,
		\u4_u3_int_stat_reg[2]/P0001 ,
		_w3892_
	);
	LUT2 #(
		.INIT('h2)
	) name2143 (
		rst_i_pad,
		\u4_u3_int_re_reg/P0001 ,
		_w3893_
	);
	LUT2 #(
		.INIT('h4)
	) name2144 (
		_w3892_,
		_w3893_,
		_w3894_
	);
	LUT3 #(
		.INIT('h07)
	) name2145 (
		\u1_u3_int_upid_set_reg/P0001 ,
		\u4_u0_ep_match_r_reg/P0001 ,
		\u4_u0_int_stat_reg[2]/P0001 ,
		_w3895_
	);
	LUT2 #(
		.INIT('h2)
	) name2146 (
		rst_i_pad,
		\u4_u0_int_re_reg/P0001 ,
		_w3896_
	);
	LUT2 #(
		.INIT('h4)
	) name2147 (
		_w3895_,
		_w3896_,
		_w3897_
	);
	LUT3 #(
		.INIT('h07)
	) name2148 (
		\u1_u3_int_upid_set_reg/P0001 ,
		\u4_u1_ep_match_r_reg/P0001 ,
		\u4_u1_int_stat_reg[2]/P0001 ,
		_w3898_
	);
	LUT2 #(
		.INIT('h2)
	) name2149 (
		rst_i_pad,
		\u4_u1_int_re_reg/P0001 ,
		_w3899_
	);
	LUT2 #(
		.INIT('h4)
	) name2150 (
		_w3898_,
		_w3899_,
		_w3900_
	);
	LUT4 #(
		.INIT('h8a00)
	) name2151 (
		_w2503_,
		_w2826_,
		_w2866_,
		_w2895_,
		_w3901_
	);
	LUT4 #(
		.INIT('h00c8)
	) name2152 (
		\u1_u3_in_token_reg/NET0131 ,
		\u4_csr_reg[0]/P0001 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		_w3902_
	);
	LUT4 #(
		.INIT('h4f00)
	) name2153 (
		_w2826_,
		_w2866_,
		_w2898_,
		_w3902_,
		_w3903_
	);
	LUT4 #(
		.INIT('ha200)
	) name2154 (
		\u1_u2_sizu_c_reg[0]/P0001 ,
		\u4_csr_reg[15]/NET0131 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		_w3904_
	);
	LUT4 #(
		.INIT('h0002)
	) name2155 (
		\u1_u2_sizu_c_reg[0]/P0001 ,
		\u1_u3_in_token_reg/NET0131 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		_w3905_
	);
	LUT3 #(
		.INIT('h01)
	) name2156 (
		_w3147_,
		_w3904_,
		_w3905_,
		_w3906_
	);
	LUT3 #(
		.INIT('hef)
	) name2157 (
		_w3901_,
		_w3903_,
		_w3906_,
		_w3907_
	);
	LUT4 #(
		.INIT('h00c8)
	) name2158 (
		\u1_u3_in_token_reg/NET0131 ,
		\u4_csr_reg[10]/P0001 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		_w3908_
	);
	LUT4 #(
		.INIT('h4f00)
	) name2159 (
		_w2826_,
		_w2866_,
		_w2908_,
		_w3908_,
		_w3909_
	);
	LUT4 #(
		.INIT('ha200)
	) name2160 (
		\u1_u2_sizu_c_reg[10]/P0001 ,
		\u4_csr_reg[15]/NET0131 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		_w3910_
	);
	LUT4 #(
		.INIT('h0002)
	) name2161 (
		\u1_u2_sizu_c_reg[10]/P0001 ,
		\u1_u3_in_token_reg/NET0131 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		_w3911_
	);
	LUT3 #(
		.INIT('h01)
	) name2162 (
		_w3088_,
		_w3910_,
		_w3911_,
		_w3912_
	);
	LUT2 #(
		.INIT('hb)
	) name2163 (
		_w3909_,
		_w3912_,
		_w3913_
	);
	LUT4 #(
		.INIT('h1000)
	) name2164 (
		_w2785_,
		_w2872_,
		_w2885_,
		_w2891_,
		_w3914_
	);
	LUT4 #(
		.INIT('h7500)
	) name2165 (
		_w2857_,
		_w2868_,
		_w2871_,
		_w3914_,
		_w3915_
	);
	LUT3 #(
		.INIT('hb0)
	) name2166 (
		_w2826_,
		_w2866_,
		_w3915_,
		_w3916_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name2167 (
		\u4_csr_reg[1]/P0001 ,
		_w2872_,
		_w2885_,
		_w2891_,
		_w3917_
	);
	LUT3 #(
		.INIT('h02)
	) name2168 (
		\u4_csr_reg[1]/P0001 ,
		_w2849_,
		_w2856_,
		_w3918_
	);
	LUT4 #(
		.INIT('h040f)
	) name2169 (
		_w2868_,
		_w2871_,
		_w3917_,
		_w3918_,
		_w3919_
	);
	LUT3 #(
		.INIT('h02)
	) name2170 (
		\u4_csr_reg[1]/P0001 ,
		_w2834_,
		_w2841_,
		_w3920_
	);
	LUT3 #(
		.INIT('h40)
	) name2171 (
		_w2827_,
		_w2865_,
		_w3920_,
		_w3921_
	);
	LUT3 #(
		.INIT('h8c)
	) name2172 (
		_w2826_,
		_w3919_,
		_w3921_,
		_w3922_
	);
	LUT2 #(
		.INIT('hb)
	) name2173 (
		_w3916_,
		_w3922_,
		_w3923_
	);
	LUT4 #(
		.INIT('ha200)
	) name2174 (
		\u1_u2_sizu_c_reg[1]/P0001 ,
		\u4_csr_reg[15]/NET0131 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		_w3924_
	);
	LUT4 #(
		.INIT('h0002)
	) name2175 (
		\u1_u2_sizu_c_reg[1]/P0001 ,
		\u1_u3_in_token_reg/NET0131 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		_w3925_
	);
	LUT3 #(
		.INIT('h01)
	) name2176 (
		_w3137_,
		_w3924_,
		_w3925_,
		_w3926_
	);
	LUT4 #(
		.INIT('h8aff)
	) name2177 (
		_w2503_,
		_w3916_,
		_w3922_,
		_w3926_,
		_w3927_
	);
	LUT4 #(
		.INIT('h0e00)
	) name2178 (
		\u1_u3_in_token_reg/NET0131 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		\u4_csr_reg[2]/NET0131 ,
		_w3928_
	);
	LUT4 #(
		.INIT('h4f00)
	) name2179 (
		_w2826_,
		_w2866_,
		_w2898_,
		_w3928_,
		_w3929_
	);
	LUT3 #(
		.INIT('ha2)
	) name2180 (
		_w2503_,
		_w2795_,
		_w2797_,
		_w3930_
	);
	LUT4 #(
		.INIT('hb000)
	) name2181 (
		_w2826_,
		_w2866_,
		_w2898_,
		_w3930_,
		_w3931_
	);
	LUT4 #(
		.INIT('ha200)
	) name2182 (
		\u1_u2_sizu_c_reg[2]/P0001 ,
		\u4_csr_reg[15]/NET0131 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		_w3932_
	);
	LUT4 #(
		.INIT('h0002)
	) name2183 (
		\u1_u2_sizu_c_reg[2]/P0001 ,
		\u1_u3_in_token_reg/NET0131 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		_w3933_
	);
	LUT3 #(
		.INIT('h01)
	) name2184 (
		_w3127_,
		_w3932_,
		_w3933_,
		_w3934_
	);
	LUT3 #(
		.INIT('hef)
	) name2185 (
		_w3929_,
		_w3931_,
		_w3934_,
		_w3935_
	);
	LUT4 #(
		.INIT('h0e00)
	) name2186 (
		\u1_u3_in_token_reg/NET0131 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		\u4_csr_reg[3]/P0001 ,
		_w3936_
	);
	LUT4 #(
		.INIT('h4f00)
	) name2187 (
		_w2826_,
		_w2866_,
		_w2898_,
		_w3936_,
		_w3937_
	);
	LUT3 #(
		.INIT('ha2)
	) name2188 (
		_w2503_,
		_w2810_,
		_w2812_,
		_w3938_
	);
	LUT4 #(
		.INIT('hb000)
	) name2189 (
		_w2826_,
		_w2866_,
		_w2898_,
		_w3938_,
		_w3939_
	);
	LUT4 #(
		.INIT('ha200)
	) name2190 (
		\u1_u2_sizu_c_reg[3]/P0001 ,
		\u4_csr_reg[15]/NET0131 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		_w3940_
	);
	LUT4 #(
		.INIT('h0002)
	) name2191 (
		\u1_u2_sizu_c_reg[3]/P0001 ,
		\u1_u3_in_token_reg/NET0131 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		_w3941_
	);
	LUT3 #(
		.INIT('h01)
	) name2192 (
		_w3117_,
		_w3940_,
		_w3941_,
		_w3942_
	);
	LUT3 #(
		.INIT('hef)
	) name2193 (
		_w3937_,
		_w3939_,
		_w3942_,
		_w3943_
	);
	LUT4 #(
		.INIT('h0e00)
	) name2194 (
		\u1_u3_in_token_reg/NET0131 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		\u4_csr_reg[4]/NET0131 ,
		_w3944_
	);
	LUT4 #(
		.INIT('h4f00)
	) name2195 (
		_w2826_,
		_w2866_,
		_w2898_,
		_w3944_,
		_w3945_
	);
	LUT3 #(
		.INIT('ha2)
	) name2196 (
		_w2503_,
		_w2803_,
		_w2805_,
		_w3946_
	);
	LUT4 #(
		.INIT('hb000)
	) name2197 (
		_w2826_,
		_w2866_,
		_w2898_,
		_w3946_,
		_w3947_
	);
	LUT4 #(
		.INIT('ha200)
	) name2198 (
		\u1_u2_sizu_c_reg[4]/P0001 ,
		\u4_csr_reg[15]/NET0131 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		_w3948_
	);
	LUT4 #(
		.INIT('h0002)
	) name2199 (
		\u1_u2_sizu_c_reg[4]/P0001 ,
		\u1_u3_in_token_reg/NET0131 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		_w3949_
	);
	LUT3 #(
		.INIT('h01)
	) name2200 (
		_w3113_,
		_w3948_,
		_w3949_,
		_w3950_
	);
	LUT3 #(
		.INIT('hef)
	) name2201 (
		_w3945_,
		_w3947_,
		_w3950_,
		_w3951_
	);
	LUT4 #(
		.INIT('h0e00)
	) name2202 (
		\u1_u3_in_token_reg/NET0131 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		\u4_csr_reg[5]/NET0131 ,
		_w3952_
	);
	LUT4 #(
		.INIT('h4f00)
	) name2203 (
		_w2826_,
		_w2866_,
		_w2898_,
		_w3952_,
		_w3953_
	);
	LUT3 #(
		.INIT('ha2)
	) name2204 (
		_w2503_,
		_w2820_,
		_w2822_,
		_w3954_
	);
	LUT4 #(
		.INIT('hb000)
	) name2205 (
		_w2826_,
		_w2866_,
		_w2898_,
		_w3954_,
		_w3955_
	);
	LUT4 #(
		.INIT('ha200)
	) name2206 (
		\u1_u2_sizu_c_reg[5]/P0001 ,
		\u4_csr_reg[15]/NET0131 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		_w3956_
	);
	LUT4 #(
		.INIT('h0002)
	) name2207 (
		\u1_u2_sizu_c_reg[5]/P0001 ,
		\u1_u3_in_token_reg/NET0131 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		_w3957_
	);
	LUT3 #(
		.INIT('h01)
	) name2208 (
		_w3108_,
		_w3956_,
		_w3957_,
		_w3958_
	);
	LUT3 #(
		.INIT('hef)
	) name2209 (
		_w3953_,
		_w3955_,
		_w3958_,
		_w3959_
	);
	LUT2 #(
		.INIT('h1)
	) name2210 (
		\u1_u2_idma_done_reg/P0001 ,
		\u1_u3_state_reg[8]/P0001 ,
		_w3960_
	);
	LUT2 #(
		.INIT('h2)
	) name2211 (
		\u4_csr_reg[24]/P0001 ,
		\u4_csr_reg[25]/P0001 ,
		_w3961_
	);
	LUT3 #(
		.INIT('ha2)
	) name2212 (
		\u1_u2_idma_done_reg/P0001 ,
		\u4_csr_reg[24]/P0001 ,
		\u4_csr_reg[25]/P0001 ,
		_w3962_
	);
	LUT4 #(
		.INIT('h0080)
	) name2213 (
		_w2127_,
		_w3676_,
		_w3861_,
		_w3962_,
		_w3963_
	);
	LUT4 #(
		.INIT('h8000)
	) name2214 (
		_w2126_,
		_w2128_,
		_w3690_,
		_w3691_,
		_w3964_
	);
	LUT3 #(
		.INIT('h0b)
	) name2215 (
		_w3960_,
		_w3963_,
		_w3964_,
		_w3965_
	);
	LUT3 #(
		.INIT('h13)
	) name2216 (
		\u1_u0_token_valid_str1_reg/P0001 ,
		\u1_u3_state_reg[8]/P0001 ,
		_w3695_,
		_w3966_
	);
	LUT3 #(
		.INIT('h04)
	) name2217 (
		\u1_u3_rx_ack_to_reg/P0001 ,
		\u1_u3_state_reg[3]/P0001 ,
		\u1_u3_state_reg[5]/P0001 ,
		_w3967_
	);
	LUT3 #(
		.INIT('h80)
	) name2218 (
		_w2127_,
		_w3699_,
		_w3967_,
		_w3968_
	);
	LUT2 #(
		.INIT('h2)
	) name2219 (
		\u1_u3_state_reg[7]/P0001 ,
		\u1_u3_state_reg[9]/P0001 ,
		_w3969_
	);
	LUT3 #(
		.INIT('h80)
	) name2220 (
		_w2128_,
		_w3687_,
		_w3969_,
		_w3970_
	);
	LUT3 #(
		.INIT('h0b)
	) name2221 (
		_w3966_,
		_w3968_,
		_w3970_,
		_w3971_
	);
	LUT4 #(
		.INIT('h0222)
	) name2222 (
		rst_i_pad,
		_w3717_,
		_w3965_,
		_w3971_,
		_w3972_
	);
	LUT3 #(
		.INIT('h2a)
	) name2223 (
		_w3750_,
		_w3965_,
		_w3971_,
		_w3973_
	);
	LUT3 #(
		.INIT('hdc)
	) name2224 (
		_w3749_,
		_w3972_,
		_w3973_,
		_w3974_
	);
	LUT4 #(
		.INIT('h0001)
	) name2225 (
		\u4_csr_reg[3]/P0001 ,
		\u4_csr_reg[4]/NET0131 ,
		\u4_csr_reg[5]/NET0131 ,
		\u4_csr_reg[6]/NET0131 ,
		_w3975_
	);
	LUT4 #(
		.INIT('h0001)
	) name2226 (
		\u4_csr_reg[0]/P0001 ,
		\u4_csr_reg[10]/P0001 ,
		\u4_csr_reg[1]/P0001 ,
		\u4_csr_reg[2]/NET0131 ,
		_w3976_
	);
	LUT3 #(
		.INIT('h01)
	) name2227 (
		\u4_csr_reg[7]/P0001 ,
		\u4_csr_reg[8]/P0001 ,
		\u4_csr_reg[9]/NET0131 ,
		_w3977_
	);
	LUT4 #(
		.INIT('h4000)
	) name2228 (
		\u1_u3_state_reg[1]/P0001 ,
		_w3975_,
		_w3976_,
		_w3977_,
		_w3978_
	);
	LUT3 #(
		.INIT('h80)
	) name2229 (
		_w2770_,
		_w2771_,
		_w3978_,
		_w3979_
	);
	LUT3 #(
		.INIT('h80)
	) name2230 (
		_w2129_,
		_w2766_,
		_w3979_,
		_w3980_
	);
	LUT2 #(
		.INIT('h1)
	) name2231 (
		\u1_u3_state_reg[1]/P0001 ,
		\u4_csr_reg[26]/NET0131 ,
		_w3981_
	);
	LUT3 #(
		.INIT('h80)
	) name2232 (
		_w2127_,
		_w2128_,
		_w3981_,
		_w3982_
	);
	LUT3 #(
		.INIT('h20)
	) name2233 (
		_w2770_,
		_w3864_,
		_w3982_,
		_w3983_
	);
	LUT2 #(
		.INIT('h8)
	) name2234 (
		_w2766_,
		_w3983_,
		_w3984_
	);
	LUT4 #(
		.INIT('h0e00)
	) name2235 (
		\u1_u3_in_token_reg/NET0131 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		\u4_csr_reg[6]/NET0131 ,
		_w3985_
	);
	LUT4 #(
		.INIT('h4f00)
	) name2236 (
		_w2826_,
		_w2866_,
		_w2898_,
		_w3985_,
		_w3986_
	);
	LUT3 #(
		.INIT('h0d)
	) name2237 (
		_w2860_,
		_w2862_,
		_w3059_,
		_w3987_
	);
	LUT4 #(
		.INIT('hb000)
	) name2238 (
		_w2826_,
		_w2866_,
		_w2898_,
		_w3987_,
		_w3988_
	);
	LUT3 #(
		.INIT('h01)
	) name2239 (
		_w3075_,
		_w3076_,
		_w3079_,
		_w3989_
	);
	LUT3 #(
		.INIT('hef)
	) name2240 (
		_w3986_,
		_w3988_,
		_w3989_,
		_w3990_
	);
	LUT3 #(
		.INIT('h01)
	) name2241 (
		_w3069_,
		_w3070_,
		_w3073_,
		_w3991_
	);
	LUT4 #(
		.INIT('h0e00)
	) name2242 (
		\u1_u3_in_token_reg/NET0131 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		\u4_csr_reg[7]/P0001 ,
		_w3992_
	);
	LUT4 #(
		.INIT('h4f00)
	) name2243 (
		_w2826_,
		_w2866_,
		_w2898_,
		_w3992_,
		_w3993_
	);
	LUT3 #(
		.INIT('h0d)
	) name2244 (
		_w2830_,
		_w2832_,
		_w3059_,
		_w3994_
	);
	LUT4 #(
		.INIT('hb000)
	) name2245 (
		_w2826_,
		_w2866_,
		_w2898_,
		_w3994_,
		_w3995_
	);
	LUT3 #(
		.INIT('hfd)
	) name2246 (
		_w3991_,
		_w3993_,
		_w3995_,
		_w3996_
	);
	LUT3 #(
		.INIT('h01)
	) name2247 (
		_w3055_,
		_w3057_,
		_w3058_,
		_w3997_
	);
	LUT4 #(
		.INIT('h0e00)
	) name2248 (
		\u1_u3_in_token_reg/NET0131 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		\u4_csr_reg[8]/P0001 ,
		_w3998_
	);
	LUT4 #(
		.INIT('h4f00)
	) name2249 (
		_w2826_,
		_w2866_,
		_w2898_,
		_w3998_,
		_w3999_
	);
	LUT3 #(
		.INIT('h0d)
	) name2250 (
		_w2837_,
		_w2839_,
		_w3059_,
		_w4000_
	);
	LUT4 #(
		.INIT('hb000)
	) name2251 (
		_w2826_,
		_w2866_,
		_w2898_,
		_w4000_,
		_w4001_
	);
	LUT3 #(
		.INIT('hfd)
	) name2252 (
		_w3997_,
		_w3999_,
		_w4001_,
		_w4002_
	);
	LUT4 #(
		.INIT('h0e00)
	) name2253 (
		\u1_u3_in_token_reg/NET0131 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		\u4_csr_reg[9]/NET0131 ,
		_w4003_
	);
	LUT4 #(
		.INIT('h4f00)
	) name2254 (
		_w2826_,
		_w2866_,
		_w2898_,
		_w4003_,
		_w4004_
	);
	LUT3 #(
		.INIT('h0d)
	) name2255 (
		_w2852_,
		_w2854_,
		_w3059_,
		_w4005_
	);
	LUT4 #(
		.INIT('hb000)
	) name2256 (
		_w2826_,
		_w2866_,
		_w2898_,
		_w4005_,
		_w4006_
	);
	LUT3 #(
		.INIT('h01)
	) name2257 (
		_w3062_,
		_w3063_,
		_w3066_,
		_w4007_
	);
	LUT3 #(
		.INIT('hef)
	) name2258 (
		_w4004_,
		_w4006_,
		_w4007_,
		_w4008_
	);
	LUT4 #(
		.INIT('hdd0d)
	) name2259 (
		\u0_rx_active_reg/P0001 ,
		\u0_rx_err_reg/P0001 ,
		\u4_csr_reg[24]/P0001 ,
		\u4_csr_reg[25]/P0001 ,
		_w4009_
	);
	LUT4 #(
		.INIT('h5d51)
	) name2260 (
		\u1_u3_state_reg[5]/P0001 ,
		_w3671_,
		_w3672_,
		_w3961_,
		_w4010_
	);
	LUT4 #(
		.INIT('h0020)
	) name2261 (
		rst_i_pad,
		_w3717_,
		_w3878_,
		_w4010_,
		_w4011_
	);
	LUT3 #(
		.INIT('h08)
	) name2262 (
		_w3750_,
		_w3878_,
		_w4010_,
		_w4012_
	);
	LUT3 #(
		.INIT('hdc)
	) name2263 (
		_w3749_,
		_w4011_,
		_w4012_,
		_w4013_
	);
	LUT3 #(
		.INIT('h10)
	) name2264 (
		\u1_u3_abort_reg/P0001 ,
		\u1_u3_state_reg[3]/P0001 ,
		\u1_u3_state_reg[5]/P0001 ,
		_w4014_
	);
	LUT3 #(
		.INIT('h80)
	) name2265 (
		_w2127_,
		_w3699_,
		_w4014_,
		_w4015_
	);
	LUT3 #(
		.INIT('h20)
	) name2266 (
		rst_i_pad,
		_w3717_,
		_w4015_,
		_w4016_
	);
	LUT4 #(
		.INIT('h8000)
	) name2267 (
		_w2127_,
		_w3699_,
		_w3750_,
		_w4014_,
		_w4017_
	);
	LUT3 #(
		.INIT('h70)
	) name2268 (
		_w3740_,
		_w3748_,
		_w4017_,
		_w4018_
	);
	LUT2 #(
		.INIT('he)
	) name2269 (
		_w4016_,
		_w4018_,
		_w4019_
	);
	LUT3 #(
		.INIT('h2a)
	) name2270 (
		_w3669_,
		_w3671_,
		_w4009_,
		_w4020_
	);
	LUT4 #(
		.INIT('hb000)
	) name2271 (
		_w3682_,
		_w3683_,
		_w3877_,
		_w4020_,
		_w4021_
	);
	LUT3 #(
		.INIT('h51)
	) name2272 (
		\u1_u3_state_reg[7]/P0001 ,
		_w3671_,
		_w3672_,
		_w4022_
	);
	LUT3 #(
		.INIT('h02)
	) name2273 (
		rst_i_pad,
		_w3717_,
		_w4022_,
		_w4023_
	);
	LUT4 #(
		.INIT('hae00)
	) name2274 (
		\u1_u3_state_reg[7]/P0001 ,
		_w3671_,
		_w3672_,
		_w3750_,
		_w4024_
	);
	LUT3 #(
		.INIT('h70)
	) name2275 (
		_w3740_,
		_w3748_,
		_w4024_,
		_w4025_
	);
	LUT3 #(
		.INIT('ha8)
	) name2276 (
		_w4021_,
		_w4023_,
		_w4025_,
		_w4026_
	);
	LUT4 #(
		.INIT('h0010)
	) name2277 (
		\u1_u3_state_reg[6]/P0001 ,
		\u1_u3_state_reg[7]/P0001 ,
		\u1_u3_state_reg[8]/P0001 ,
		\u1_u3_state_reg[9]/P0001 ,
		_w4027_
	);
	LUT2 #(
		.INIT('h8)
	) name2278 (
		_w2128_,
		_w4027_,
		_w4028_
	);
	LUT3 #(
		.INIT('h20)
	) name2279 (
		rst_i_pad,
		_w3717_,
		_w4028_,
		_w4029_
	);
	LUT3 #(
		.INIT('h80)
	) name2280 (
		_w2128_,
		_w3750_,
		_w4027_,
		_w4030_
	);
	LUT3 #(
		.INIT('h70)
	) name2281 (
		_w3740_,
		_w3748_,
		_w4030_,
		_w4031_
	);
	LUT3 #(
		.INIT('ha8)
	) name2282 (
		_w3675_,
		_w4029_,
		_w4031_,
		_w4032_
	);
	LUT4 #(
		.INIT('h11b1)
	) name2283 (
		\u1_u2_idma_done_reg/P0001 ,
		\u1_u3_state_reg[3]/P0001 ,
		\u4_csr_reg[24]/P0001 ,
		\u4_csr_reg[25]/P0001 ,
		_w4033_
	);
	LUT4 #(
		.INIT('h0080)
	) name2284 (
		_w2127_,
		_w3676_,
		_w3861_,
		_w4033_,
		_w4034_
	);
	LUT3 #(
		.INIT('h4c)
	) name2285 (
		\u1_u0_token_valid_str1_reg/P0001 ,
		\u1_u3_state_reg[3]/P0001 ,
		_w3695_,
		_w4035_
	);
	LUT3 #(
		.INIT('h13)
	) name2286 (
		_w3968_,
		_w4034_,
		_w4035_,
		_w4036_
	);
	LUT3 #(
		.INIT('h02)
	) name2287 (
		rst_i_pad,
		_w3717_,
		_w4036_,
		_w4037_
	);
	LUT4 #(
		.INIT('ha8a0)
	) name2288 (
		_w3750_,
		_w3968_,
		_w4034_,
		_w4035_,
		_w4038_
	);
	LUT3 #(
		.INIT('h70)
	) name2289 (
		_w3740_,
		_w3748_,
		_w4038_,
		_w4039_
	);
	LUT2 #(
		.INIT('he)
	) name2290 (
		_w4037_,
		_w4039_,
		_w4040_
	);
	LUT2 #(
		.INIT('h2)
	) name2291 (
		rst_i_pad,
		\u4_int_src_re_reg/P0001 ,
		_w4041_
	);
	LUT4 #(
		.INIT('h2220)
	) name2292 (
		rst_i_pad,
		\u4_int_src_re_reg/P0001 ,
		\u4_int_srcb_reg[2]/P0001 ,
		\u4_nse_err_r_reg/P0001 ,
		_w4042_
	);
	LUT3 #(
		.INIT('h04)
	) name2293 (
		\u1_u3_adr_reg[8]/P0001 ,
		_w2837_,
		_w2839_,
		_w4043_
	);
	LUT3 #(
		.INIT('h04)
	) name2294 (
		\u1_u3_adr_reg[11]/P0001 ,
		_w2881_,
		_w2883_,
		_w4044_
	);
	LUT3 #(
		.INIT('h04)
	) name2295 (
		\u1_u3_adr_reg[12]/P0001 ,
		_w2875_,
		_w2877_,
		_w4045_
	);
	LUT2 #(
		.INIT('h1)
	) name2296 (
		_w4044_,
		_w4045_,
		_w4046_
	);
	LUT3 #(
		.INIT('h04)
	) name2297 (
		\u1_u3_adr_reg[10]/P0001 ,
		_w2845_,
		_w2847_,
		_w4047_
	);
	LUT3 #(
		.INIT('h04)
	) name2298 (
		\u1_u3_adr_reg[9]/P0001 ,
		_w2852_,
		_w2854_,
		_w4048_
	);
	LUT4 #(
		.INIT('h0001)
	) name2299 (
		_w4044_,
		_w4045_,
		_w4047_,
		_w4048_,
		_w4049_
	);
	LUT2 #(
		.INIT('h4)
	) name2300 (
		_w4043_,
		_w4049_,
		_w4050_
	);
	LUT3 #(
		.INIT('ha2)
	) name2301 (
		\u1_u3_adr_reg[9]/P0001 ,
		_w2852_,
		_w2854_,
		_w4051_
	);
	LUT3 #(
		.INIT('ha2)
	) name2302 (
		\u1_u3_adr_reg[11]/P0001 ,
		_w2881_,
		_w2883_,
		_w4052_
	);
	LUT3 #(
		.INIT('ha2)
	) name2303 (
		\u1_u3_adr_reg[10]/P0001 ,
		_w2845_,
		_w2847_,
		_w4053_
	);
	LUT4 #(
		.INIT('h004d)
	) name2304 (
		\u1_u3_adr_reg[10]/P0001 ,
		_w2848_,
		_w4051_,
		_w4052_,
		_w4054_
	);
	LUT3 #(
		.INIT('ha2)
	) name2305 (
		\u1_u3_adr_reg[13]/P0001 ,
		_w2888_,
		_w2890_,
		_w4055_
	);
	LUT3 #(
		.INIT('h04)
	) name2306 (
		\u1_u3_adr_reg[13]/P0001 ,
		_w2888_,
		_w2890_,
		_w4056_
	);
	LUT3 #(
		.INIT('h59)
	) name2307 (
		\u1_u3_adr_reg[13]/P0001 ,
		_w2888_,
		_w2890_,
		_w4057_
	);
	LUT3 #(
		.INIT('ha2)
	) name2308 (
		\u1_u3_adr_reg[12]/P0001 ,
		_w2875_,
		_w2877_,
		_w4058_
	);
	LUT2 #(
		.INIT('h2)
	) name2309 (
		_w4057_,
		_w4058_,
		_w4059_
	);
	LUT3 #(
		.INIT('hd0)
	) name2310 (
		_w4046_,
		_w4054_,
		_w4059_,
		_w4060_
	);
	LUT2 #(
		.INIT('h4)
	) name2311 (
		_w4050_,
		_w4060_,
		_w4061_
	);
	LUT3 #(
		.INIT('h04)
	) name2312 (
		\u1_u3_adr_reg[6]/P0001 ,
		_w2860_,
		_w2862_,
		_w4062_
	);
	LUT3 #(
		.INIT('h04)
	) name2313 (
		\u1_u3_adr_reg[7]/P0001 ,
		_w2830_,
		_w2832_,
		_w4063_
	);
	LUT3 #(
		.INIT('ha2)
	) name2314 (
		\u1_u3_adr_reg[6]/P0001 ,
		_w2860_,
		_w2862_,
		_w4064_
	);
	LUT3 #(
		.INIT('ha2)
	) name2315 (
		\u1_u3_adr_reg[5]/P0001 ,
		_w2820_,
		_w2822_,
		_w4065_
	);
	LUT4 #(
		.INIT('h0b02)
	) name2316 (
		\u1_u3_adr_reg[6]/P0001 ,
		_w2863_,
		_w4063_,
		_w4065_,
		_w4066_
	);
	LUT3 #(
		.INIT('h04)
	) name2317 (
		\u1_u3_adr_reg[5]/P0001 ,
		_w2820_,
		_w2822_,
		_w4067_
	);
	LUT3 #(
		.INIT('h04)
	) name2318 (
		\u1_u3_adr_reg[4]/P0001 ,
		_w2803_,
		_w2805_,
		_w4068_
	);
	LUT4 #(
		.INIT('h0001)
	) name2319 (
		_w4062_,
		_w4063_,
		_w4067_,
		_w4068_,
		_w4069_
	);
	LUT2 #(
		.INIT('h1)
	) name2320 (
		_w4066_,
		_w4069_,
		_w4070_
	);
	LUT3 #(
		.INIT('ha2)
	) name2321 (
		\u1_u3_adr_reg[0]/P0001 ,
		_w2788_,
		_w2790_,
		_w4071_
	);
	LUT3 #(
		.INIT('ha2)
	) name2322 (
		\u1_u3_adr_reg[2]/P0001 ,
		_w2795_,
		_w2797_,
		_w4072_
	);
	LUT4 #(
		.INIT('h004d)
	) name2323 (
		\u1_u3_adr_reg[1]/P0001 ,
		_w2785_,
		_w4071_,
		_w4072_,
		_w4073_
	);
	LUT3 #(
		.INIT('h04)
	) name2324 (
		\u1_u3_adr_reg[3]/P0001 ,
		_w2810_,
		_w2812_,
		_w4074_
	);
	LUT3 #(
		.INIT('h04)
	) name2325 (
		\u1_u3_adr_reg[2]/P0001 ,
		_w2795_,
		_w2797_,
		_w4075_
	);
	LUT2 #(
		.INIT('h1)
	) name2326 (
		_w4074_,
		_w4075_,
		_w4076_
	);
	LUT3 #(
		.INIT('ha2)
	) name2327 (
		\u1_u3_adr_reg[4]/P0001 ,
		_w2803_,
		_w2805_,
		_w4077_
	);
	LUT3 #(
		.INIT('ha2)
	) name2328 (
		\u1_u3_adr_reg[3]/P0001 ,
		_w2810_,
		_w2812_,
		_w4078_
	);
	LUT2 #(
		.INIT('h1)
	) name2329 (
		_w4077_,
		_w4078_,
		_w4079_
	);
	LUT4 #(
		.INIT('h4500)
	) name2330 (
		_w4066_,
		_w4073_,
		_w4076_,
		_w4079_,
		_w4080_
	);
	LUT3 #(
		.INIT('ha2)
	) name2331 (
		\u1_u3_adr_reg[8]/P0001 ,
		_w2837_,
		_w2839_,
		_w4081_
	);
	LUT3 #(
		.INIT('ha2)
	) name2332 (
		\u1_u3_adr_reg[7]/P0001 ,
		_w2830_,
		_w2832_,
		_w4082_
	);
	LUT2 #(
		.INIT('h1)
	) name2333 (
		_w4081_,
		_w4082_,
		_w4083_
	);
	LUT4 #(
		.INIT('hd000)
	) name2334 (
		_w4046_,
		_w4054_,
		_w4059_,
		_w4083_,
		_w4084_
	);
	LUT3 #(
		.INIT('he0)
	) name2335 (
		_w4070_,
		_w4080_,
		_w4084_,
		_w4085_
	);
	LUT2 #(
		.INIT('h1)
	) name2336 (
		_w4061_,
		_w4085_,
		_w4086_
	);
	LUT3 #(
		.INIT('h0d)
	) name2337 (
		_w4046_,
		_w4054_,
		_w4058_,
		_w4087_
	);
	LUT2 #(
		.INIT('h4)
	) name2338 (
		_w4050_,
		_w4087_,
		_w4088_
	);
	LUT4 #(
		.INIT('h0d00)
	) name2339 (
		_w4046_,
		_w4054_,
		_w4058_,
		_w4083_,
		_w4089_
	);
	LUT3 #(
		.INIT('he0)
	) name2340 (
		_w4070_,
		_w4080_,
		_w4089_,
		_w4090_
	);
	LUT3 #(
		.INIT('h01)
	) name2341 (
		_w4057_,
		_w4088_,
		_w4090_,
		_w4091_
	);
	LUT2 #(
		.INIT('hd)
	) name2342 (
		_w4086_,
		_w4091_,
		_w4092_
	);
	LUT2 #(
		.INIT('h1)
	) name2343 (
		\u0_u0_state_reg[13]/NET0131 ,
		\u0_u0_state_reg[14]/P0001 ,
		_w4093_
	);
	LUT3 #(
		.INIT('h01)
	) name2344 (
		\u0_u0_state_reg[0]/NET0131 ,
		\u0_u0_state_reg[13]/NET0131 ,
		\u0_u0_state_reg[14]/P0001 ,
		_w4094_
	);
	LUT4 #(
		.INIT('h0002)
	) name2345 (
		\u0_u0_state_reg[10]/P0001 ,
		\u0_u0_state_reg[7]/NET0131 ,
		\u0_u0_state_reg[8]/NET0131 ,
		\u0_u0_state_reg[9]/P0001 ,
		_w4095_
	);
	LUT2 #(
		.INIT('h1)
	) name2346 (
		\u0_u0_state_reg[4]/NET0131 ,
		\u0_u0_state_reg[5]/P0001 ,
		_w4096_
	);
	LUT2 #(
		.INIT('h1)
	) name2347 (
		\u0_u0_state_reg[3]/P0001 ,
		\u0_u0_state_reg[6]/NET0131 ,
		_w4097_
	);
	LUT4 #(
		.INIT('h0001)
	) name2348 (
		\u0_u0_state_reg[3]/P0001 ,
		\u0_u0_state_reg[4]/NET0131 ,
		\u0_u0_state_reg[5]/P0001 ,
		\u0_u0_state_reg[6]/NET0131 ,
		_w4098_
	);
	LUT2 #(
		.INIT('h1)
	) name2349 (
		\u0_u0_state_reg[1]/P0001 ,
		\u0_u0_state_reg[2]/NET0131 ,
		_w4099_
	);
	LUT2 #(
		.INIT('h1)
	) name2350 (
		\u0_u0_state_reg[11]/NET0131 ,
		\u0_u0_state_reg[12]/NET0131 ,
		_w4100_
	);
	LUT4 #(
		.INIT('h0001)
	) name2351 (
		\u0_u0_state_reg[11]/NET0131 ,
		\u0_u0_state_reg[12]/NET0131 ,
		\u0_u0_state_reg[1]/P0001 ,
		\u0_u0_state_reg[2]/NET0131 ,
		_w4101_
	);
	LUT4 #(
		.INIT('h8000)
	) name2352 (
		_w4094_,
		_w4095_,
		_w4098_,
		_w4101_,
		_w4102_
	);
	LUT2 #(
		.INIT('h2)
	) name2353 (
		rst_i_pad,
		usb_vbus_pad_i_pad,
		_w4103_
	);
	LUT2 #(
		.INIT('hd)
	) name2354 (
		rst_i_pad,
		usb_vbus_pad_i_pad,
		_w4104_
	);
	LUT4 #(
		.INIT('h00a8)
	) name2355 (
		rst_i_pad,
		\u0_u0_T2_gt_1_0_mS_reg/P0001 ,
		\u0_u0_state_reg[11]/NET0131 ,
		usb_vbus_pad_i_pad,
		_w4105_
	);
	LUT2 #(
		.INIT('h8)
	) name2356 (
		_w4102_,
		_w4105_,
		_w4106_
	);
	LUT2 #(
		.INIT('he)
	) name2357 (
		\u0_u0_state_reg[10]/P0001 ,
		\u0_u0_state_reg[7]/NET0131 ,
		_w4107_
	);
	LUT3 #(
		.INIT('h01)
	) name2358 (
		\u0_u0_state_reg[10]/P0001 ,
		\u0_u0_state_reg[7]/NET0131 ,
		\u0_u0_state_reg[8]/NET0131 ,
		_w4108_
	);
	LUT4 #(
		.INIT('h0001)
	) name2359 (
		\u0_u0_state_reg[0]/NET0131 ,
		\u0_u0_state_reg[13]/NET0131 ,
		\u0_u0_state_reg[14]/P0001 ,
		\u0_u0_state_reg[9]/P0001 ,
		_w4109_
	);
	LUT4 #(
		.INIT('h8000)
	) name2360 (
		_w4098_,
		_w4099_,
		_w4108_,
		_w4109_,
		_w4110_
	);
	LUT2 #(
		.INIT('h2)
	) name2361 (
		\LineState_r_reg[0]/P0001 ,
		\LineState_r_reg[1]/P0001 ,
		_w4111_
	);
	LUT3 #(
		.INIT('h20)
	) name2362 (
		\LineState_r_reg[0]/P0001 ,
		\LineState_r_reg[1]/P0001 ,
		\u0_u0_ls_j_r_reg/P0001 ,
		_w4112_
	);
	LUT2 #(
		.INIT('h4)
	) name2363 (
		\u0_u0_state_reg[11]/NET0131 ,
		\u0_u0_state_reg[12]/NET0131 ,
		_w4113_
	);
	LUT2 #(
		.INIT('h8)
	) name2364 (
		_w4112_,
		_w4113_,
		_w4114_
	);
	LUT2 #(
		.INIT('h2)
	) name2365 (
		\u0_u0_state_reg[11]/NET0131 ,
		\u0_u0_state_reg[12]/NET0131 ,
		_w4115_
	);
	LUT2 #(
		.INIT('h1)
	) name2366 (
		\LineState_r_reg[0]/P0001 ,
		\LineState_r_reg[1]/P0001 ,
		_w4116_
	);
	LUT3 #(
		.INIT('h10)
	) name2367 (
		\LineState_r_reg[0]/P0001 ,
		\LineState_r_reg[1]/P0001 ,
		\u0_u0_ls_se0_r_reg/P0001 ,
		_w4117_
	);
	LUT2 #(
		.INIT('h4)
	) name2368 (
		\LineState_r_reg[0]/P0001 ,
		\LineState_r_reg[1]/P0001 ,
		_w4118_
	);
	LUT3 #(
		.INIT('h40)
	) name2369 (
		\LineState_r_reg[0]/P0001 ,
		\LineState_r_reg[1]/P0001 ,
		\u0_u0_ls_k_r_reg/P0001 ,
		_w4119_
	);
	LUT4 #(
		.INIT('haebf)
	) name2370 (
		\LineState_r_reg[0]/P0001 ,
		\LineState_r_reg[1]/P0001 ,
		\u0_u0_ls_k_r_reg/P0001 ,
		\u0_u0_ls_se0_r_reg/P0001 ,
		_w4120_
	);
	LUT2 #(
		.INIT('h8)
	) name2371 (
		_w4115_,
		_w4120_,
		_w4121_
	);
	LUT3 #(
		.INIT('h02)
	) name2372 (
		rst_i_pad,
		\u0_u0_chirp_cnt_is_6_reg/P0001 ,
		usb_vbus_pad_i_pad,
		_w4122_
	);
	LUT4 #(
		.INIT('ha800)
	) name2373 (
		_w4110_,
		_w4114_,
		_w4121_,
		_w4122_,
		_w4123_
	);
	LUT2 #(
		.INIT('he)
	) name2374 (
		_w4106_,
		_w4123_,
		_w4124_
	);
	LUT4 #(
		.INIT('hf351)
	) name2375 (
		\u4_u3_csr0_reg[10]/P0001 ,
		\u4_u3_csr0_reg[9]/P0001 ,
		\u4_u3_dma_out_left_reg[7]/P0001 ,
		\u4_u3_dma_out_left_reg[8]/P0001 ,
		_w4125_
	);
	LUT4 #(
		.INIT('h8caf)
	) name2376 (
		\u4_u3_csr0_reg[8]/P0001 ,
		\u4_u3_csr0_reg[9]/P0001 ,
		\u4_u3_dma_out_left_reg[6]/P0001 ,
		\u4_u3_dma_out_left_reg[7]/P0001 ,
		_w4126_
	);
	LUT2 #(
		.INIT('h2)
	) name2377 (
		_w4125_,
		_w4126_,
		_w4127_
	);
	LUT4 #(
		.INIT('h8caf)
	) name2378 (
		\u4_u3_csr0_reg[6]/P0001 ,
		\u4_u3_csr0_reg[7]/P0001 ,
		\u4_u3_dma_out_left_reg[4]/P0001 ,
		\u4_u3_dma_out_left_reg[5]/P0001 ,
		_w4128_
	);
	LUT4 #(
		.INIT('hf531)
	) name2379 (
		\u4_u3_csr0_reg[5]/P0001 ,
		\u4_u3_csr0_reg[6]/P0001 ,
		\u4_u3_dma_out_left_reg[3]/P0001 ,
		\u4_u3_dma_out_left_reg[4]/P0001 ,
		_w4129_
	);
	LUT2 #(
		.INIT('h2)
	) name2380 (
		_w4128_,
		_w4129_,
		_w4130_
	);
	LUT4 #(
		.INIT('h080a)
	) name2381 (
		\u4_u3_csr0_reg[2]/P0001 ,
		\u4_u3_csr0_reg[3]/NET0131 ,
		\u4_u3_dma_out_left_reg[0]/P0001 ,
		\u4_u3_dma_out_left_reg[1]/P0001 ,
		_w4131_
	);
	LUT4 #(
		.INIT('hf531)
	) name2382 (
		\u4_u3_csr0_reg[3]/NET0131 ,
		\u4_u3_csr0_reg[4]/P0001 ,
		\u4_u3_dma_out_left_reg[1]/P0001 ,
		\u4_u3_dma_out_left_reg[2]/P0001 ,
		_w4132_
	);
	LUT4 #(
		.INIT('h8caf)
	) name2383 (
		\u4_u3_csr0_reg[4]/P0001 ,
		\u4_u3_csr0_reg[5]/P0001 ,
		\u4_u3_dma_out_left_reg[2]/P0001 ,
		\u4_u3_dma_out_left_reg[3]/P0001 ,
		_w4133_
	);
	LUT4 #(
		.INIT('h8a00)
	) name2384 (
		_w4128_,
		_w4131_,
		_w4132_,
		_w4133_,
		_w4134_
	);
	LUT4 #(
		.INIT('hf531)
	) name2385 (
		\u4_u3_csr0_reg[7]/P0001 ,
		\u4_u3_csr0_reg[8]/P0001 ,
		\u4_u3_dma_out_left_reg[5]/P0001 ,
		\u4_u3_dma_out_left_reg[6]/P0001 ,
		_w4135_
	);
	LUT2 #(
		.INIT('h8)
	) name2386 (
		_w4125_,
		_w4135_,
		_w4136_
	);
	LUT4 #(
		.INIT('h5455)
	) name2387 (
		_w4127_,
		_w4130_,
		_w4134_,
		_w4136_,
		_w4137_
	);
	LUT2 #(
		.INIT('h4)
	) name2388 (
		\u4_u3_csr0_reg[10]/P0001 ,
		\u4_u3_dma_out_left_reg[8]/P0001 ,
		_w4138_
	);
	LUT3 #(
		.INIT('h01)
	) name2389 (
		\u4_u3_dma_out_left_reg[10]/P0001 ,
		\u4_u3_dma_out_left_reg[11]/P0001 ,
		\u4_u3_dma_out_left_reg[9]/P0001 ,
		_w4139_
	);
	LUT2 #(
		.INIT('h4)
	) name2390 (
		_w4138_,
		_w4139_,
		_w4140_
	);
	LUT2 #(
		.INIT('h7)
	) name2391 (
		_w4137_,
		_w4140_,
		_w4141_
	);
	LUT4 #(
		.INIT('hf351)
	) name2392 (
		\u4_u0_csr0_reg[10]/P0001 ,
		\u4_u0_csr0_reg[9]/P0001 ,
		\u4_u0_dma_out_left_reg[7]/P0001 ,
		\u4_u0_dma_out_left_reg[8]/P0001 ,
		_w4142_
	);
	LUT4 #(
		.INIT('h8caf)
	) name2393 (
		\u4_u0_csr0_reg[8]/P0001 ,
		\u4_u0_csr0_reg[9]/P0001 ,
		\u4_u0_dma_out_left_reg[6]/P0001 ,
		\u4_u0_dma_out_left_reg[7]/P0001 ,
		_w4143_
	);
	LUT2 #(
		.INIT('h2)
	) name2394 (
		_w4142_,
		_w4143_,
		_w4144_
	);
	LUT4 #(
		.INIT('h8caf)
	) name2395 (
		\u4_u0_csr0_reg[6]/P0001 ,
		\u4_u0_csr0_reg[7]/P0001 ,
		\u4_u0_dma_out_left_reg[4]/P0001 ,
		\u4_u0_dma_out_left_reg[5]/P0001 ,
		_w4145_
	);
	LUT4 #(
		.INIT('hf531)
	) name2396 (
		\u4_u0_csr0_reg[5]/P0001 ,
		\u4_u0_csr0_reg[6]/P0001 ,
		\u4_u0_dma_out_left_reg[3]/P0001 ,
		\u4_u0_dma_out_left_reg[4]/P0001 ,
		_w4146_
	);
	LUT2 #(
		.INIT('h2)
	) name2397 (
		_w4145_,
		_w4146_,
		_w4147_
	);
	LUT4 #(
		.INIT('h080a)
	) name2398 (
		\u4_u0_csr0_reg[2]/P0001 ,
		\u4_u0_csr0_reg[3]/NET0131 ,
		\u4_u0_dma_out_left_reg[0]/P0001 ,
		\u4_u0_dma_out_left_reg[1]/P0001 ,
		_w4148_
	);
	LUT4 #(
		.INIT('hf531)
	) name2399 (
		\u4_u0_csr0_reg[3]/NET0131 ,
		\u4_u0_csr0_reg[4]/P0001 ,
		\u4_u0_dma_out_left_reg[1]/P0001 ,
		\u4_u0_dma_out_left_reg[2]/P0001 ,
		_w4149_
	);
	LUT4 #(
		.INIT('h8caf)
	) name2400 (
		\u4_u0_csr0_reg[4]/P0001 ,
		\u4_u0_csr0_reg[5]/P0001 ,
		\u4_u0_dma_out_left_reg[2]/P0001 ,
		\u4_u0_dma_out_left_reg[3]/P0001 ,
		_w4150_
	);
	LUT4 #(
		.INIT('h8a00)
	) name2401 (
		_w4145_,
		_w4148_,
		_w4149_,
		_w4150_,
		_w4151_
	);
	LUT4 #(
		.INIT('hf531)
	) name2402 (
		\u4_u0_csr0_reg[7]/P0001 ,
		\u4_u0_csr0_reg[8]/P0001 ,
		\u4_u0_dma_out_left_reg[5]/P0001 ,
		\u4_u0_dma_out_left_reg[6]/P0001 ,
		_w4152_
	);
	LUT2 #(
		.INIT('h8)
	) name2403 (
		_w4142_,
		_w4152_,
		_w4153_
	);
	LUT4 #(
		.INIT('h5455)
	) name2404 (
		_w4144_,
		_w4147_,
		_w4151_,
		_w4153_,
		_w4154_
	);
	LUT2 #(
		.INIT('h4)
	) name2405 (
		\u4_u0_csr0_reg[10]/P0001 ,
		\u4_u0_dma_out_left_reg[8]/P0001 ,
		_w4155_
	);
	LUT3 #(
		.INIT('h01)
	) name2406 (
		\u4_u0_dma_out_left_reg[10]/P0001 ,
		\u4_u0_dma_out_left_reg[11]/P0001 ,
		\u4_u0_dma_out_left_reg[9]/P0001 ,
		_w4156_
	);
	LUT2 #(
		.INIT('h4)
	) name2407 (
		_w4155_,
		_w4156_,
		_w4157_
	);
	LUT2 #(
		.INIT('h7)
	) name2408 (
		_w4154_,
		_w4157_,
		_w4158_
	);
	LUT4 #(
		.INIT('hf351)
	) name2409 (
		\u4_u1_csr0_reg[10]/P0001 ,
		\u4_u1_csr0_reg[9]/P0001 ,
		\u4_u1_dma_out_left_reg[7]/P0001 ,
		\u4_u1_dma_out_left_reg[8]/P0001 ,
		_w4159_
	);
	LUT4 #(
		.INIT('h8caf)
	) name2410 (
		\u4_u1_csr0_reg[8]/P0001 ,
		\u4_u1_csr0_reg[9]/P0001 ,
		\u4_u1_dma_out_left_reg[6]/P0001 ,
		\u4_u1_dma_out_left_reg[7]/P0001 ,
		_w4160_
	);
	LUT2 #(
		.INIT('h2)
	) name2411 (
		_w4159_,
		_w4160_,
		_w4161_
	);
	LUT4 #(
		.INIT('h8caf)
	) name2412 (
		\u4_u1_csr0_reg[6]/P0001 ,
		\u4_u1_csr0_reg[7]/P0001 ,
		\u4_u1_dma_out_left_reg[4]/P0001 ,
		\u4_u1_dma_out_left_reg[5]/P0001 ,
		_w4162_
	);
	LUT4 #(
		.INIT('hf531)
	) name2413 (
		\u4_u1_csr0_reg[5]/P0001 ,
		\u4_u1_csr0_reg[6]/P0001 ,
		\u4_u1_dma_out_left_reg[3]/P0001 ,
		\u4_u1_dma_out_left_reg[4]/P0001 ,
		_w4163_
	);
	LUT2 #(
		.INIT('h2)
	) name2414 (
		_w4162_,
		_w4163_,
		_w4164_
	);
	LUT4 #(
		.INIT('h080a)
	) name2415 (
		\u4_u1_csr0_reg[2]/P0001 ,
		\u4_u1_csr0_reg[3]/NET0131 ,
		\u4_u1_dma_out_left_reg[0]/P0001 ,
		\u4_u1_dma_out_left_reg[1]/P0001 ,
		_w4165_
	);
	LUT4 #(
		.INIT('hf531)
	) name2416 (
		\u4_u1_csr0_reg[3]/NET0131 ,
		\u4_u1_csr0_reg[4]/P0001 ,
		\u4_u1_dma_out_left_reg[1]/P0001 ,
		\u4_u1_dma_out_left_reg[2]/P0001 ,
		_w4166_
	);
	LUT4 #(
		.INIT('h8caf)
	) name2417 (
		\u4_u1_csr0_reg[4]/P0001 ,
		\u4_u1_csr0_reg[5]/P0001 ,
		\u4_u1_dma_out_left_reg[2]/P0001 ,
		\u4_u1_dma_out_left_reg[3]/P0001 ,
		_w4167_
	);
	LUT4 #(
		.INIT('h8a00)
	) name2418 (
		_w4162_,
		_w4165_,
		_w4166_,
		_w4167_,
		_w4168_
	);
	LUT4 #(
		.INIT('hf531)
	) name2419 (
		\u4_u1_csr0_reg[7]/P0001 ,
		\u4_u1_csr0_reg[8]/P0001 ,
		\u4_u1_dma_out_left_reg[5]/P0001 ,
		\u4_u1_dma_out_left_reg[6]/P0001 ,
		_w4169_
	);
	LUT2 #(
		.INIT('h8)
	) name2420 (
		_w4159_,
		_w4169_,
		_w4170_
	);
	LUT4 #(
		.INIT('h5455)
	) name2421 (
		_w4161_,
		_w4164_,
		_w4168_,
		_w4170_,
		_w4171_
	);
	LUT2 #(
		.INIT('h4)
	) name2422 (
		\u4_u1_csr0_reg[10]/P0001 ,
		\u4_u1_dma_out_left_reg[8]/P0001 ,
		_w4172_
	);
	LUT3 #(
		.INIT('h01)
	) name2423 (
		\u4_u1_dma_out_left_reg[10]/P0001 ,
		\u4_u1_dma_out_left_reg[11]/P0001 ,
		\u4_u1_dma_out_left_reg[9]/P0001 ,
		_w4173_
	);
	LUT2 #(
		.INIT('h4)
	) name2424 (
		_w4172_,
		_w4173_,
		_w4174_
	);
	LUT2 #(
		.INIT('h7)
	) name2425 (
		_w4171_,
		_w4174_,
		_w4175_
	);
	LUT4 #(
		.INIT('hf351)
	) name2426 (
		\u4_u2_csr0_reg[10]/P0001 ,
		\u4_u2_csr0_reg[9]/P0001 ,
		\u4_u2_dma_out_left_reg[7]/P0001 ,
		\u4_u2_dma_out_left_reg[8]/P0001 ,
		_w4176_
	);
	LUT4 #(
		.INIT('h8caf)
	) name2427 (
		\u4_u2_csr0_reg[8]/P0001 ,
		\u4_u2_csr0_reg[9]/P0001 ,
		\u4_u2_dma_out_left_reg[6]/P0001 ,
		\u4_u2_dma_out_left_reg[7]/P0001 ,
		_w4177_
	);
	LUT2 #(
		.INIT('h2)
	) name2428 (
		_w4176_,
		_w4177_,
		_w4178_
	);
	LUT4 #(
		.INIT('h8caf)
	) name2429 (
		\u4_u2_csr0_reg[6]/P0001 ,
		\u4_u2_csr0_reg[7]/P0001 ,
		\u4_u2_dma_out_left_reg[4]/P0001 ,
		\u4_u2_dma_out_left_reg[5]/P0001 ,
		_w4179_
	);
	LUT4 #(
		.INIT('hf531)
	) name2430 (
		\u4_u2_csr0_reg[5]/P0001 ,
		\u4_u2_csr0_reg[6]/P0001 ,
		\u4_u2_dma_out_left_reg[3]/P0001 ,
		\u4_u2_dma_out_left_reg[4]/P0001 ,
		_w4180_
	);
	LUT2 #(
		.INIT('h2)
	) name2431 (
		_w4179_,
		_w4180_,
		_w4181_
	);
	LUT4 #(
		.INIT('h080a)
	) name2432 (
		\u4_u2_csr0_reg[2]/P0001 ,
		\u4_u2_csr0_reg[3]/NET0131 ,
		\u4_u2_dma_out_left_reg[0]/P0001 ,
		\u4_u2_dma_out_left_reg[1]/P0001 ,
		_w4182_
	);
	LUT4 #(
		.INIT('hf531)
	) name2433 (
		\u4_u2_csr0_reg[3]/NET0131 ,
		\u4_u2_csr0_reg[4]/P0001 ,
		\u4_u2_dma_out_left_reg[1]/P0001 ,
		\u4_u2_dma_out_left_reg[2]/P0001 ,
		_w4183_
	);
	LUT4 #(
		.INIT('h8caf)
	) name2434 (
		\u4_u2_csr0_reg[4]/P0001 ,
		\u4_u2_csr0_reg[5]/P0001 ,
		\u4_u2_dma_out_left_reg[2]/P0001 ,
		\u4_u2_dma_out_left_reg[3]/P0001 ,
		_w4184_
	);
	LUT4 #(
		.INIT('h8a00)
	) name2435 (
		_w4179_,
		_w4182_,
		_w4183_,
		_w4184_,
		_w4185_
	);
	LUT4 #(
		.INIT('hf531)
	) name2436 (
		\u4_u2_csr0_reg[7]/P0001 ,
		\u4_u2_csr0_reg[8]/P0001 ,
		\u4_u2_dma_out_left_reg[5]/P0001 ,
		\u4_u2_dma_out_left_reg[6]/P0001 ,
		_w4186_
	);
	LUT2 #(
		.INIT('h8)
	) name2437 (
		_w4176_,
		_w4186_,
		_w4187_
	);
	LUT4 #(
		.INIT('h5455)
	) name2438 (
		_w4178_,
		_w4181_,
		_w4185_,
		_w4187_,
		_w4188_
	);
	LUT2 #(
		.INIT('h4)
	) name2439 (
		\u4_u2_csr0_reg[10]/P0001 ,
		\u4_u2_dma_out_left_reg[8]/P0001 ,
		_w4189_
	);
	LUT3 #(
		.INIT('h01)
	) name2440 (
		\u4_u2_dma_out_left_reg[10]/P0001 ,
		\u4_u2_dma_out_left_reg[11]/P0001 ,
		\u4_u2_dma_out_left_reg[9]/P0001 ,
		_w4190_
	);
	LUT2 #(
		.INIT('h4)
	) name2441 (
		_w4189_,
		_w4190_,
		_w4191_
	);
	LUT2 #(
		.INIT('h7)
	) name2442 (
		_w4188_,
		_w4191_,
		_w4192_
	);
	LUT3 #(
		.INIT('h15)
	) name2443 (
		\u1_u3_buffer_overflow_reg/P0001 ,
		\u1_u3_match_r_reg/P0001 ,
		\u1_u3_to_large_reg/P0001 ,
		_w4193_
	);
	LUT3 #(
		.INIT('hd0)
	) name2444 (
		_w3717_,
		_w3720_,
		_w4193_,
		_w4194_
	);
	LUT4 #(
		.INIT('h0222)
	) name2445 (
		\u1_u0_token_valid_str1_reg/P0001 ,
		\u1_u3_buffer_overflow_reg/P0001 ,
		\u1_u3_match_r_reg/P0001 ,
		\u1_u3_to_large_reg/P0001 ,
		_w4195_
	);
	LUT3 #(
		.INIT('h70)
	) name2446 (
		_w3740_,
		_w3748_,
		_w4195_,
		_w4196_
	);
	LUT2 #(
		.INIT('h1)
	) name2447 (
		_w4194_,
		_w4196_,
		_w4197_
	);
	LUT4 #(
		.INIT('h0100)
	) name2448 (
		\u0_u0_state_reg[10]/P0001 ,
		\u0_u0_state_reg[7]/NET0131 ,
		\u0_u0_state_reg[8]/NET0131 ,
		\u0_u0_state_reg[9]/P0001 ,
		_w4198_
	);
	LUT4 #(
		.INIT('h8000)
	) name2449 (
		_w4094_,
		_w4098_,
		_w4101_,
		_w4198_,
		_w4199_
	);
	LUT4 #(
		.INIT('h01af)
	) name2450 (
		\u0_u0_T2_gt_1_0_mS_reg/P0001 ,
		\u0_u0_state_reg[10]/P0001 ,
		_w4102_,
		_w4199_,
		_w4200_
	);
	LUT2 #(
		.INIT('h2)
	) name2451 (
		_w4103_,
		_w4200_,
		_w4201_
	);
	LUT4 #(
		.INIT('h8ecf)
	) name2452 (
		\u1_u3_adr_reg[6]/P0001 ,
		\u1_u3_adr_reg[7]/P0001 ,
		_w2833_,
		_w2863_,
		_w4202_
	);
	LUT3 #(
		.INIT('h4d)
	) name2453 (
		\u1_u3_adr_reg[7]/P0001 ,
		_w2833_,
		_w4064_,
		_w4203_
	);
	LUT3 #(
		.INIT('h4d)
	) name2454 (
		\u1_u3_adr_reg[5]/P0001 ,
		_w2823_,
		_w4077_,
		_w4204_
	);
	LUT3 #(
		.INIT('h2a)
	) name2455 (
		_w4202_,
		_w4203_,
		_w4204_,
		_w4205_
	);
	LUT3 #(
		.INIT('h0e)
	) name2456 (
		_w4073_,
		_w4075_,
		_w4078_,
		_w4206_
	);
	LUT3 #(
		.INIT('h01)
	) name2457 (
		_w4067_,
		_w4068_,
		_w4074_,
		_w4207_
	);
	LUT2 #(
		.INIT('h8)
	) name2458 (
		_w4202_,
		_w4207_,
		_w4208_
	);
	LUT4 #(
		.INIT('h0001)
	) name2459 (
		_w4044_,
		_w4045_,
		_w4047_,
		_w4056_,
		_w4209_
	);
	LUT2 #(
		.INIT('h1)
	) name2460 (
		_w4043_,
		_w4048_,
		_w4210_
	);
	LUT2 #(
		.INIT('h8)
	) name2461 (
		_w4209_,
		_w4210_,
		_w4211_
	);
	LUT4 #(
		.INIT('hba00)
	) name2462 (
		_w4205_,
		_w4206_,
		_w4208_,
		_w4211_,
		_w4212_
	);
	LUT4 #(
		.INIT('h0b02)
	) name2463 (
		\u1_u3_adr_reg[11]/P0001 ,
		_w2884_,
		_w4045_,
		_w4053_,
		_w4213_
	);
	LUT2 #(
		.INIT('h1)
	) name2464 (
		_w4055_,
		_w4058_,
		_w4214_
	);
	LUT3 #(
		.INIT('h45)
	) name2465 (
		_w4056_,
		_w4213_,
		_w4214_,
		_w4215_
	);
	LUT3 #(
		.INIT('h4d)
	) name2466 (
		\u1_u3_adr_reg[9]/P0001 ,
		_w2855_,
		_w4081_,
		_w4216_
	);
	LUT2 #(
		.INIT('h2)
	) name2467 (
		_w4209_,
		_w4216_,
		_w4217_
	);
	LUT4 #(
		.INIT('h5556)
	) name2468 (
		\u1_u3_adr_reg[14]/P0001 ,
		_w4212_,
		_w4215_,
		_w4217_,
		_w4218_
	);
	LUT2 #(
		.INIT('h8)
	) name2469 (
		\u1_frame_no_same_reg/P0001 ,
		\u1_mfm_cnt_reg[0]/P0001 ,
		_w4219_
	);
	LUT3 #(
		.INIT('ha2)
	) name2470 (
		rst_i_pad,
		\u1_clr_sof_time_reg/P0001 ,
		\u1_frame_no_same_reg/P0001 ,
		_w4220_
	);
	LUT3 #(
		.INIT('h60)
	) name2471 (
		\u1_mfm_cnt_reg[1]/P0001 ,
		_w4219_,
		_w4220_,
		_w4221_
	);
	LUT3 #(
		.INIT('h07)
	) name2472 (
		\u1_u3_int_seqerr_set_reg/P0001 ,
		\u4_u2_ep_match_r_reg/P0001 ,
		\u4_u2_int_stat_reg[5]/P0001 ,
		_w4222_
	);
	LUT2 #(
		.INIT('h2)
	) name2473 (
		_w3890_,
		_w4222_,
		_w4223_
	);
	LUT4 #(
		.INIT('h02a0)
	) name2474 (
		rst_i_pad,
		\u1_clr_sof_time_reg/P0001 ,
		\u1_frame_no_same_reg/P0001 ,
		\u1_mfm_cnt_reg[0]/P0001 ,
		_w4224_
	);
	LUT4 #(
		.INIT('h007f)
	) name2475 (
		\u1_frame_no_same_reg/P0001 ,
		\u1_mfm_cnt_reg[0]/P0001 ,
		\u1_mfm_cnt_reg[1]/P0001 ,
		\u1_mfm_cnt_reg[2]/P0001 ,
		_w4225_
	);
	LUT4 #(
		.INIT('h8000)
	) name2476 (
		\u1_frame_no_same_reg/P0001 ,
		\u1_mfm_cnt_reg[0]/P0001 ,
		\u1_mfm_cnt_reg[1]/P0001 ,
		\u1_mfm_cnt_reg[2]/P0001 ,
		_w4226_
	);
	LUT3 #(
		.INIT('h02)
	) name2477 (
		_w4220_,
		_w4225_,
		_w4226_,
		_w4227_
	);
	LUT4 #(
		.INIT('ha200)
	) name2478 (
		rst_i_pad,
		\u1_clr_sof_time_reg/P0001 ,
		\u1_frame_no_same_reg/P0001 ,
		\u1_mfm_cnt_reg[3]/P0001 ,
		_w4228_
	);
	LUT4 #(
		.INIT('h00a2)
	) name2479 (
		rst_i_pad,
		\u1_clr_sof_time_reg/P0001 ,
		\u1_frame_no_same_reg/P0001 ,
		\u1_mfm_cnt_reg[3]/P0001 ,
		_w4229_
	);
	LUT3 #(
		.INIT('he4)
	) name2480 (
		_w4226_,
		_w4228_,
		_w4229_,
		_w4230_
	);
	LUT3 #(
		.INIT('h07)
	) name2481 (
		\u1_u3_int_seqerr_set_reg/P0001 ,
		\u4_u3_ep_match_r_reg/P0001 ,
		\u4_u3_int_stat_reg[5]/P0001 ,
		_w4231_
	);
	LUT2 #(
		.INIT('h2)
	) name2482 (
		_w3893_,
		_w4231_,
		_w4232_
	);
	LUT3 #(
		.INIT('h07)
	) name2483 (
		\u1_u3_int_seqerr_set_reg/P0001 ,
		\u4_u0_ep_match_r_reg/P0001 ,
		\u4_u0_int_stat_reg[5]/P0001 ,
		_w4233_
	);
	LUT2 #(
		.INIT('h2)
	) name2484 (
		_w3896_,
		_w4233_,
		_w4234_
	);
	LUT3 #(
		.INIT('h07)
	) name2485 (
		\u1_u3_int_seqerr_set_reg/P0001 ,
		\u4_u1_ep_match_r_reg/P0001 ,
		\u4_u1_int_stat_reg[5]/P0001 ,
		_w4235_
	);
	LUT2 #(
		.INIT('h2)
	) name2486 (
		_w3899_,
		_w4235_,
		_w4236_
	);
	LUT2 #(
		.INIT('h2)
	) name2487 (
		\u1_u3_match_r_reg/P0001 ,
		_w2131_,
		_w4237_
	);
	LUT3 #(
		.INIT('h04)
	) name2488 (
		\u1_u3_pid_IN_r_reg/P0001 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		_w4238_
	);
	LUT3 #(
		.INIT('h0e)
	) name2489 (
		\u1_u3_pid_IN_r_reg/P0001 ,
		\u1_u3_pid_SETUP_r_reg/P0001 ,
		\u4_csr_reg[27]/NET0131 ,
		_w4239_
	);
	LUT3 #(
		.INIT('h01)
	) name2490 (
		\u1_u3_pid_OUT_r_reg/P0001 ,
		\u1_u3_pid_PING_r_reg/P0001 ,
		\u4_csr_reg[26]/NET0131 ,
		_w4240_
	);
	LUT3 #(
		.INIT('h45)
	) name2491 (
		_w4238_,
		_w4239_,
		_w4240_,
		_w4241_
	);
	LUT2 #(
		.INIT('h2)
	) name2492 (
		_w4237_,
		_w4241_,
		_w4242_
	);
	LUT4 #(
		.INIT('h20aa)
	) name2493 (
		\u4_csr_reg[0]/P0001 ,
		_w2826_,
		_w2866_,
		_w2898_,
		_w4243_
	);
	LUT2 #(
		.INIT('he)
	) name2494 (
		_w2896_,
		_w4243_,
		_w4244_
	);
	LUT4 #(
		.INIT('h20aa)
	) name2495 (
		\u4_csr_reg[10]/P0001 ,
		_w2826_,
		_w2866_,
		_w2908_,
		_w4245_
	);
	LUT4 #(
		.INIT('h20aa)
	) name2496 (
		\u4_csr_reg[3]/P0001 ,
		_w2826_,
		_w2866_,
		_w2898_,
		_w4246_
	);
	LUT2 #(
		.INIT('he)
	) name2497 (
		_w2950_,
		_w4246_,
		_w4247_
	);
	LUT4 #(
		.INIT('h20aa)
	) name2498 (
		\u4_csr_reg[4]/NET0131 ,
		_w2826_,
		_w2866_,
		_w2898_,
		_w4248_
	);
	LUT2 #(
		.INIT('he)
	) name2499 (
		_w2961_,
		_w4248_,
		_w4249_
	);
	LUT4 #(
		.INIT('h20aa)
	) name2500 (
		\u4_csr_reg[5]/NET0131 ,
		_w2826_,
		_w2866_,
		_w2898_,
		_w4250_
	);
	LUT2 #(
		.INIT('he)
	) name2501 (
		_w2973_,
		_w4250_,
		_w4251_
	);
	LUT4 #(
		.INIT('h20aa)
	) name2502 (
		\u4_csr_reg[6]/NET0131 ,
		_w2826_,
		_w2866_,
		_w2898_,
		_w4252_
	);
	LUT2 #(
		.INIT('he)
	) name2503 (
		_w2984_,
		_w4252_,
		_w4253_
	);
	LUT4 #(
		.INIT('h20aa)
	) name2504 (
		\u4_csr_reg[7]/P0001 ,
		_w2826_,
		_w2866_,
		_w2898_,
		_w4254_
	);
	LUT2 #(
		.INIT('he)
	) name2505 (
		_w2994_,
		_w4254_,
		_w4255_
	);
	LUT4 #(
		.INIT('h20aa)
	) name2506 (
		\u4_csr_reg[8]/P0001 ,
		_w2826_,
		_w2866_,
		_w2898_,
		_w4256_
	);
	LUT2 #(
		.INIT('he)
	) name2507 (
		_w3004_,
		_w4256_,
		_w4257_
	);
	LUT4 #(
		.INIT('h20aa)
	) name2508 (
		\u4_csr_reg[9]/NET0131 ,
		_w2826_,
		_w2866_,
		_w2898_,
		_w4258_
	);
	LUT2 #(
		.INIT('he)
	) name2509 (
		_w3013_,
		_w4258_,
		_w4259_
	);
	LUT4 #(
		.INIT('h2202)
	) name2510 (
		\u1_u0_pid_reg[0]/NET0131 ,
		\u1_u0_pid_reg[1]/NET0131 ,
		\u1_u0_pid_reg[2]/NET0131 ,
		\u1_u0_pid_reg[3]/NET0131 ,
		_w4260_
	);
	LUT2 #(
		.INIT('h8)
	) name2511 (
		\u1_u0_token_valid_str1_reg/P0001 ,
		_w4260_,
		_w4261_
	);
	LUT2 #(
		.INIT('h4)
	) name2512 (
		_w3717_,
		_w4261_,
		_w4262_
	);
	LUT3 #(
		.INIT('h70)
	) name2513 (
		_w3740_,
		_w3748_,
		_w4261_,
		_w4263_
	);
	LUT2 #(
		.INIT('he)
	) name2514 (
		_w4262_,
		_w4263_,
		_w4264_
	);
	LUT3 #(
		.INIT('hac)
	) name2515 (
		\u1_u2_sizu_c_reg[8]/NET0131 ,
		\u1_u3_new_size_reg[8]/P0001 ,
		\u1_u3_out_to_small_r_reg/P0001 ,
		_w4265_
	);
	LUT3 #(
		.INIT('hac)
	) name2516 (
		\u1_u2_sizu_c_reg[9]/P0001 ,
		\u1_u3_new_size_reg[9]/P0001 ,
		\u1_u3_out_to_small_r_reg/P0001 ,
		_w4266_
	);
	LUT4 #(
		.INIT('hba00)
	) name2517 (
		_w4205_,
		_w4206_,
		_w4208_,
		_w4210_,
		_w4267_
	);
	LUT3 #(
		.INIT('h59)
	) name2518 (
		\u1_u3_adr_reg[10]/P0001 ,
		_w2845_,
		_w2847_,
		_w4268_
	);
	LUT3 #(
		.INIT('h01)
	) name2519 (
		_w4043_,
		_w4048_,
		_w4268_,
		_w4269_
	);
	LUT4 #(
		.INIT('hba00)
	) name2520 (
		_w4205_,
		_w4206_,
		_w4208_,
		_w4269_,
		_w4270_
	);
	LUT4 #(
		.INIT('hff25)
	) name2521 (
		_w4216_,
		_w4267_,
		_w4268_,
		_w4270_,
		_w4271_
	);
	LUT3 #(
		.INIT('h59)
	) name2522 (
		\u1_u3_adr_reg[12]/P0001 ,
		_w2875_,
		_w2877_,
		_w4272_
	);
	LUT3 #(
		.INIT('hb2)
	) name2523 (
		\u1_u3_adr_reg[11]/P0001 ,
		_w2884_,
		_w4053_,
		_w4273_
	);
	LUT2 #(
		.INIT('h1)
	) name2524 (
		_w4044_,
		_w4047_,
		_w4274_
	);
	LUT2 #(
		.INIT('h4)
	) name2525 (
		_w4216_,
		_w4274_,
		_w4275_
	);
	LUT4 #(
		.INIT('h0001)
	) name2526 (
		_w4043_,
		_w4044_,
		_w4047_,
		_w4048_,
		_w4276_
	);
	LUT4 #(
		.INIT('hba00)
	) name2527 (
		_w4205_,
		_w4206_,
		_w4208_,
		_w4276_,
		_w4277_
	);
	LUT4 #(
		.INIT('h5556)
	) name2528 (
		_w4272_,
		_w4273_,
		_w4275_,
		_w4277_,
		_w4278_
	);
	LUT3 #(
		.INIT('h59)
	) name2529 (
		\u1_u3_adr_reg[9]/P0001 ,
		_w2852_,
		_w2854_,
		_w4279_
	);
	LUT2 #(
		.INIT('h1)
	) name2530 (
		_w4043_,
		_w4279_,
		_w4280_
	);
	LUT4 #(
		.INIT('h1f00)
	) name2531 (
		_w4070_,
		_w4080_,
		_w4083_,
		_w4280_,
		_w4281_
	);
	LUT2 #(
		.INIT('h8)
	) name2532 (
		_w4043_,
		_w4279_,
		_w4282_
	);
	LUT3 #(
		.INIT('h10)
	) name2533 (
		_w4081_,
		_w4082_,
		_w4279_,
		_w4283_
	);
	LUT4 #(
		.INIT('h010f)
	) name2534 (
		_w4070_,
		_w4080_,
		_w4282_,
		_w4283_,
		_w4284_
	);
	LUT2 #(
		.INIT('hb)
	) name2535 (
		_w4281_,
		_w4284_,
		_w4285_
	);
	LUT3 #(
		.INIT('h08)
	) name2536 (
		\u1_u2_sizu_c_reg[10]/P0001 ,
		_w2845_,
		_w2847_,
		_w4286_
	);
	LUT3 #(
		.INIT('h51)
	) name2537 (
		\u1_u2_sizu_c_reg[9]/P0001 ,
		_w2852_,
		_w2854_,
		_w4287_
	);
	LUT3 #(
		.INIT('h08)
	) name2538 (
		\u1_u2_sizu_c_reg[8]/NET0131 ,
		_w2837_,
		_w2839_,
		_w4288_
	);
	LUT4 #(
		.INIT('h0107)
	) name2539 (
		\u1_u2_sizu_c_reg[9]/P0001 ,
		_w2855_,
		_w4286_,
		_w4288_,
		_w4289_
	);
	LUT4 #(
		.INIT('h88a8)
	) name2540 (
		\u1_u0_data_valid0_reg/P0001 ,
		\u1_u2_sizu_c_reg[10]/P0001 ,
		_w2845_,
		_w2847_,
		_w4290_
	);
	LUT2 #(
		.INIT('h4)
	) name2541 (
		_w4289_,
		_w4290_,
		_w4291_
	);
	LUT3 #(
		.INIT('h08)
	) name2542 (
		\u1_u2_sizu_c_reg[7]/P0001 ,
		_w2830_,
		_w2832_,
		_w4292_
	);
	LUT3 #(
		.INIT('h08)
	) name2543 (
		\u1_u2_sizu_c_reg[6]/P0001 ,
		_w2860_,
		_w2862_,
		_w4293_
	);
	LUT3 #(
		.INIT('h51)
	) name2544 (
		\u1_u2_sizu_c_reg[5]/P0001 ,
		_w2820_,
		_w2822_,
		_w4294_
	);
	LUT4 #(
		.INIT('h0701)
	) name2545 (
		\u1_u2_sizu_c_reg[6]/P0001 ,
		_w2863_,
		_w4292_,
		_w4294_,
		_w4295_
	);
	LUT3 #(
		.INIT('h51)
	) name2546 (
		\u1_u2_sizu_c_reg[3]/P0001 ,
		_w2810_,
		_w2812_,
		_w4296_
	);
	LUT3 #(
		.INIT('h51)
	) name2547 (
		\u1_u2_sizu_c_reg[4]/P0001 ,
		_w2803_,
		_w2805_,
		_w4297_
	);
	LUT3 #(
		.INIT('h08)
	) name2548 (
		\u1_u2_sizu_c_reg[2]/P0001 ,
		_w2795_,
		_w2797_,
		_w4298_
	);
	LUT4 #(
		.INIT('h0e08)
	) name2549 (
		\u1_u2_sizu_c_reg[3]/P0001 ,
		_w2813_,
		_w4297_,
		_w4298_,
		_w4299_
	);
	LUT4 #(
		.INIT('h3313)
	) name2550 (
		\u1_u2_sizu_c_reg[0]/P0001 ,
		\u1_u2_sizu_c_reg[1]/P0001 ,
		_w2788_,
		_w2790_,
		_w4300_
	);
	LUT3 #(
		.INIT('h51)
	) name2551 (
		\u1_u2_sizu_c_reg[2]/P0001 ,
		_w2795_,
		_w2797_,
		_w4301_
	);
	LUT2 #(
		.INIT('h1)
	) name2552 (
		_w4300_,
		_w4301_,
		_w4302_
	);
	LUT2 #(
		.INIT('h8)
	) name2553 (
		\u1_u2_sizu_c_reg[0]/P0001 ,
		\u1_u2_sizu_c_reg[1]/P0001 ,
		_w4303_
	);
	LUT3 #(
		.INIT('h20)
	) name2554 (
		_w2788_,
		_w2790_,
		_w4303_,
		_w4304_
	);
	LUT4 #(
		.INIT('h0302)
	) name2555 (
		_w2785_,
		_w4296_,
		_w4297_,
		_w4304_,
		_w4305_
	);
	LUT3 #(
		.INIT('h08)
	) name2556 (
		\u1_u2_sizu_c_reg[5]/P0001 ,
		_w2820_,
		_w2822_,
		_w4306_
	);
	LUT3 #(
		.INIT('h08)
	) name2557 (
		\u1_u2_sizu_c_reg[4]/P0001 ,
		_w2803_,
		_w2805_,
		_w4307_
	);
	LUT4 #(
		.INIT('h0001)
	) name2558 (
		_w4292_,
		_w4293_,
		_w4306_,
		_w4307_,
		_w4308_
	);
	LUT4 #(
		.INIT('h1500)
	) name2559 (
		_w4299_,
		_w4302_,
		_w4305_,
		_w4308_,
		_w4309_
	);
	LUT3 #(
		.INIT('h51)
	) name2560 (
		\u1_u2_sizu_c_reg[8]/NET0131 ,
		_w2837_,
		_w2839_,
		_w4310_
	);
	LUT3 #(
		.INIT('h51)
	) name2561 (
		\u1_u2_sizu_c_reg[7]/P0001 ,
		_w2830_,
		_w2832_,
		_w4311_
	);
	LUT4 #(
		.INIT('h0004)
	) name2562 (
		_w4287_,
		_w4290_,
		_w4310_,
		_w4311_,
		_w4312_
	);
	LUT4 #(
		.INIT('h5455)
	) name2563 (
		_w4291_,
		_w4295_,
		_w4309_,
		_w4312_,
		_w4313_
	);
	LUT2 #(
		.INIT('h2)
	) name2564 (
		_w2892_,
		_w4313_,
		_w4314_
	);
	LUT2 #(
		.INIT('h8)
	) name2565 (
		\u0_u0_T1_gt_3_0_mS_reg/P0001 ,
		\u0_u0_mode_hs_reg/P0001 ,
		_w4315_
	);
	LUT4 #(
		.INIT('h0008)
	) name2566 (
		\u0_u0_T1_gt_2_5_uS_reg/P0001 ,
		\u0_u0_T1_st_3_0_mS_reg/P0001 ,
		\u0_u0_idle_long_reg/P0001 ,
		\u0_u0_mode_hs_reg/P0001 ,
		_w4316_
	);
	LUT2 #(
		.INIT('h1)
	) name2567 (
		_w4315_,
		_w4316_,
		_w4317_
	);
	LUT4 #(
		.INIT('h0001)
	) name2568 (
		\u0_u0_state_reg[11]/NET0131 ,
		\u0_u0_state_reg[12]/NET0131 ,
		\u0_u0_state_reg[3]/P0001 ,
		\u0_u0_state_reg[6]/NET0131 ,
		_w4318_
	);
	LUT4 #(
		.INIT('h8000)
	) name2569 (
		_w4099_,
		_w4108_,
		_w4109_,
		_w4318_,
		_w4319_
	);
	LUT2 #(
		.INIT('h4)
	) name2570 (
		\u0_u0_state_reg[4]/NET0131 ,
		\u0_u0_state_reg[5]/P0001 ,
		_w4320_
	);
	LUT2 #(
		.INIT('h2)
	) name2571 (
		\u0_u0_state_reg[4]/NET0131 ,
		\u0_u0_state_reg[5]/P0001 ,
		_w4321_
	);
	LUT2 #(
		.INIT('h9)
	) name2572 (
		\u0_u0_state_reg[4]/NET0131 ,
		\u0_u0_state_reg[5]/P0001 ,
		_w4322_
	);
	LUT4 #(
		.INIT('h0001)
	) name2573 (
		\u0_u0_state_reg[11]/NET0131 ,
		\u0_u0_state_reg[12]/NET0131 ,
		\u0_u0_state_reg[4]/NET0131 ,
		\u0_u0_state_reg[5]/P0001 ,
		_w4323_
	);
	LUT2 #(
		.INIT('h2)
	) name2574 (
		\u0_u0_state_reg[1]/P0001 ,
		\u0_u0_state_reg[2]/NET0131 ,
		_w4324_
	);
	LUT4 #(
		.INIT('h0002)
	) name2575 (
		\u0_u0_state_reg[1]/P0001 ,
		\u0_u0_state_reg[2]/NET0131 ,
		\u0_u0_state_reg[3]/P0001 ,
		\u0_u0_state_reg[6]/NET0131 ,
		_w4325_
	);
	LUT4 #(
		.INIT('h8000)
	) name2576 (
		_w4108_,
		_w4109_,
		_w4323_,
		_w4325_,
		_w4326_
	);
	LUT4 #(
		.INIT('h0100)
	) name2577 (
		\u0_u0_state_reg[1]/P0001 ,
		\u0_u0_state_reg[2]/NET0131 ,
		\u0_u0_state_reg[4]/NET0131 ,
		\u0_u0_state_reg[5]/P0001 ,
		_w4327_
	);
	LUT4 #(
		.INIT('h8000)
	) name2578 (
		_w4108_,
		_w4109_,
		_w4318_,
		_w4327_,
		_w4328_
	);
	LUT4 #(
		.INIT('hddd0)
	) name2579 (
		_w4319_,
		_w4322_,
		_w4326_,
		_w4328_,
		_w4329_
	);
	LUT2 #(
		.INIT('h4)
	) name2580 (
		_w4317_,
		_w4329_,
		_w4330_
	);
	LUT4 #(
		.INIT('h0001)
	) name2581 (
		\u0_u0_state_reg[10]/P0001 ,
		\u0_u0_state_reg[7]/NET0131 ,
		\u0_u0_state_reg[8]/NET0131 ,
		\u0_u0_state_reg[9]/P0001 ,
		_w4331_
	);
	LUT3 #(
		.INIT('h02)
	) name2582 (
		\u0_u0_state_reg[0]/NET0131 ,
		\u0_u0_state_reg[13]/NET0131 ,
		\u0_u0_state_reg[14]/P0001 ,
		_w4332_
	);
	LUT4 #(
		.INIT('h8000)
	) name2583 (
		_w4098_,
		_w4101_,
		_w4331_,
		_w4332_,
		_w4333_
	);
	LUT4 #(
		.INIT('h000d)
	) name2584 (
		_w4319_,
		_w4322_,
		_w4326_,
		_w4328_,
		_w4334_
	);
	LUT4 #(
		.INIT('h0010)
	) name2585 (
		\LineState_r_reg[0]/P0001 ,
		\LineState_r_reg[1]/P0001 ,
		\u0_u0_state_reg[4]/NET0131 ,
		\u0_u0_state_reg[5]/P0001 ,
		_w4335_
	);
	LUT3 #(
		.INIT('h20)
	) name2586 (
		_w4319_,
		_w4326_,
		_w4335_,
		_w4336_
	);
	LUT4 #(
		.INIT('h0302)
	) name2587 (
		\u0_u0_T2_wakeup_reg/P0001 ,
		\u0_u0_state_reg[1]/P0001 ,
		\u0_u0_state_reg[2]/NET0131 ,
		\u0_u0_state_reg[7]/NET0131 ,
		_w4337_
	);
	LUT4 #(
		.INIT('h8000)
	) name2588 (
		_w4108_,
		_w4109_,
		_w4318_,
		_w4337_,
		_w4338_
	);
	LUT2 #(
		.INIT('h8)
	) name2589 (
		_w4320_,
		_w4338_,
		_w4339_
	);
	LUT4 #(
		.INIT('h0007)
	) name2590 (
		_w4333_,
		_w4334_,
		_w4336_,
		_w4339_,
		_w4340_
	);
	LUT2 #(
		.INIT('h2)
	) name2591 (
		\u0_u0_state_reg[3]/P0001 ,
		\u0_u0_state_reg[6]/NET0131 ,
		_w4341_
	);
	LUT4 #(
		.INIT('h0010)
	) name2592 (
		\u0_u0_state_reg[1]/P0001 ,
		\u0_u0_state_reg[2]/NET0131 ,
		\u0_u0_state_reg[3]/P0001 ,
		\u0_u0_state_reg[6]/NET0131 ,
		_w4342_
	);
	LUT4 #(
		.INIT('h8000)
	) name2593 (
		_w4108_,
		_w4109_,
		_w4323_,
		_w4342_,
		_w4343_
	);
	LUT4 #(
		.INIT('hdf00)
	) name2594 (
		_w4319_,
		_w4326_,
		_w4335_,
		_w4343_,
		_w4344_
	);
	LUT2 #(
		.INIT('h4)
	) name2595 (
		\u0_u0_state_reg[1]/P0001 ,
		\u0_u0_state_reg[2]/NET0131 ,
		_w4345_
	);
	LUT4 #(
		.INIT('h0004)
	) name2596 (
		\u0_u0_state_reg[1]/P0001 ,
		\u0_u0_state_reg[2]/NET0131 ,
		\u0_u0_state_reg[3]/P0001 ,
		\u0_u0_state_reg[6]/NET0131 ,
		_w4346_
	);
	LUT4 #(
		.INIT('h8000)
	) name2597 (
		_w4108_,
		_w4109_,
		_w4323_,
		_w4346_,
		_w4347_
	);
	LUT2 #(
		.INIT('h1)
	) name2598 (
		_w4199_,
		_w4347_,
		_w4348_
	);
	LUT2 #(
		.INIT('h4)
	) name2599 (
		_w4344_,
		_w4348_,
		_w4349_
	);
	LUT3 #(
		.INIT('hb0)
	) name2600 (
		_w4330_,
		_w4340_,
		_w4349_,
		_w4350_
	);
	LUT4 #(
		.INIT('h2220)
	) name2601 (
		_w4319_,
		_w4322_,
		_w4343_,
		_w4347_,
		_w4351_
	);
	LUT4 #(
		.INIT('h00fd)
	) name2602 (
		\u0_u0_T2_gt_1_0_mS_reg/P0001 ,
		_w4326_,
		_w4328_,
		_w4343_,
		_w4352_
	);
	LUT3 #(
		.INIT('h0e)
	) name2603 (
		_w4199_,
		_w4351_,
		_w4352_,
		_w4353_
	);
	LUT4 #(
		.INIT('h1000)
	) name2604 (
		\LineState_r_reg[0]/P0001 ,
		\LineState_r_reg[1]/P0001 ,
		\u0_u0_T1_gt_2_5_uS_reg/P0001 ,
		\u0_u0_ls_se0_r_reg/P0001 ,
		_w4354_
	);
	LUT4 #(
		.INIT('h2000)
	) name2605 (
		\LineState_r_reg[0]/P0001 ,
		\LineState_r_reg[1]/P0001 ,
		\u0_u0_T2_gt_100_uS_reg/P0001 ,
		\u0_u0_ls_j_r_reg/P0001 ,
		_w4355_
	);
	LUT4 #(
		.INIT('h1000)
	) name2606 (
		\LineState_r_reg[0]/P0001 ,
		\LineState_r_reg[1]/P0001 ,
		\u0_u0_T2_gt_100_uS_reg/P0001 ,
		\u0_u0_ls_se0_r_reg/P0001 ,
		_w4356_
	);
	LUT3 #(
		.INIT('h0d)
	) name2607 (
		\u0_u0_state_reg[9]/P0001 ,
		_w4355_,
		_w4356_,
		_w4357_
	);
	LUT4 #(
		.INIT('h5f13)
	) name2608 (
		_w4343_,
		_w4347_,
		_w4354_,
		_w4357_,
		_w4358_
	);
	LUT4 #(
		.INIT('h4000)
	) name2609 (
		\u0_u0_me_cnt_reg[2]/P0001 ,
		\u0_u0_me_cnt_reg[3]/P0001 ,
		\u0_u0_me_cnt_reg[6]/P0001 ,
		\u0_u0_me_cnt_reg[7]/P0001 ,
		_w4359_
	);
	LUT4 #(
		.INIT('h0001)
	) name2610 (
		\u0_u0_me_cnt_reg[0]/P0001 ,
		\u0_u0_me_cnt_reg[1]/P0001 ,
		\u0_u0_me_cnt_reg[4]/P0001 ,
		\u0_u0_me_cnt_reg[5]/P0001 ,
		_w4360_
	);
	LUT2 #(
		.INIT('h8)
	) name2611 (
		_w4359_,
		_w4360_,
		_w4361_
	);
	LUT2 #(
		.INIT('h8)
	) name2612 (
		_w4358_,
		_w4361_,
		_w4362_
	);
	LUT2 #(
		.INIT('h4)
	) name2613 (
		_w4353_,
		_w4362_,
		_w4363_
	);
	LUT2 #(
		.INIT('h4)
	) name2614 (
		_w4350_,
		_w4363_,
		_w4364_
	);
	LUT2 #(
		.INIT('h8)
	) name2615 (
		\u1_hms_clk_reg/P0001 ,
		\u1_sof_time_reg[0]/P0001 ,
		_w4365_
	);
	LUT3 #(
		.INIT('h80)
	) name2616 (
		\u1_sof_time_reg[6]/P0001 ,
		\u1_sof_time_reg[7]/P0001 ,
		\u1_sof_time_reg[8]/P0001 ,
		_w4366_
	);
	LUT3 #(
		.INIT('h80)
	) name2617 (
		\u1_sof_time_reg[3]/P0001 ,
		\u1_sof_time_reg[4]/P0001 ,
		\u1_sof_time_reg[5]/P0001 ,
		_w4367_
	);
	LUT2 #(
		.INIT('h8)
	) name2618 (
		\u1_sof_time_reg[1]/P0001 ,
		\u1_sof_time_reg[2]/P0001 ,
		_w4368_
	);
	LUT4 #(
		.INIT('h8000)
	) name2619 (
		\u1_sof_time_reg[10]/P0001 ,
		\u1_sof_time_reg[1]/P0001 ,
		\u1_sof_time_reg[2]/P0001 ,
		\u1_sof_time_reg[9]/P0001 ,
		_w4369_
	);
	LUT4 #(
		.INIT('h8000)
	) name2620 (
		_w4365_,
		_w4366_,
		_w4367_,
		_w4369_,
		_w4370_
	);
	LUT3 #(
		.INIT('h14)
	) name2621 (
		\u1_clr_sof_time_reg/P0001 ,
		\u1_sof_time_reg[11]/P0001 ,
		_w4370_,
		_w4371_
	);
	LUT3 #(
		.INIT('h01)
	) name2622 (
		_w4043_,
		_w4047_,
		_w4048_,
		_w4372_
	);
	LUT3 #(
		.INIT('h4d)
	) name2623 (
		\u1_u3_adr_reg[10]/P0001 ,
		_w2848_,
		_w4051_,
		_w4373_
	);
	LUT3 #(
		.INIT('h59)
	) name2624 (
		\u1_u3_adr_reg[11]/P0001 ,
		_w2881_,
		_w2883_,
		_w4374_
	);
	LUT4 #(
		.INIT('h4d00)
	) name2625 (
		\u1_u3_adr_reg[10]/P0001 ,
		_w2848_,
		_w4051_,
		_w4374_,
		_w4375_
	);
	LUT2 #(
		.INIT('h4)
	) name2626 (
		_w4372_,
		_w4375_,
		_w4376_
	);
	LUT2 #(
		.INIT('h8)
	) name2627 (
		_w4083_,
		_w4375_,
		_w4377_
	);
	LUT4 #(
		.INIT('h010f)
	) name2628 (
		_w4070_,
		_w4080_,
		_w4376_,
		_w4377_,
		_w4378_
	);
	LUT2 #(
		.INIT('h4)
	) name2629 (
		_w4372_,
		_w4373_,
		_w4379_
	);
	LUT2 #(
		.INIT('h8)
	) name2630 (
		_w4083_,
		_w4373_,
		_w4380_
	);
	LUT4 #(
		.INIT('h010f)
	) name2631 (
		_w4070_,
		_w4080_,
		_w4379_,
		_w4380_,
		_w4381_
	);
	LUT3 #(
		.INIT('h73)
	) name2632 (
		_w4374_,
		_w4378_,
		_w4381_,
		_w4382_
	);
	LUT2 #(
		.INIT('h2)
	) name2633 (
		\u4_u3_csr0_reg[2]/P0001 ,
		\u4_u3_dma_in_cnt_reg[0]/P0001 ,
		_w4383_
	);
	LUT4 #(
		.INIT('hf531)
	) name2634 (
		\u4_u3_csr0_reg[2]/P0001 ,
		\u4_u3_csr0_reg[3]/NET0131 ,
		\u4_u3_dma_in_cnt_reg[0]/P0001 ,
		\u4_u3_dma_in_cnt_reg[1]/P0001 ,
		_w4384_
	);
	LUT4 #(
		.INIT('h8caf)
	) name2635 (
		\u4_u3_csr0_reg[3]/NET0131 ,
		\u4_u3_csr0_reg[4]/P0001 ,
		\u4_u3_dma_in_cnt_reg[1]/P0001 ,
		\u4_u3_dma_in_cnt_reg[2]/P0001 ,
		_w4385_
	);
	LUT2 #(
		.INIT('h2)
	) name2636 (
		\u4_u3_csr0_reg[6]/P0001 ,
		\u4_u3_dma_in_cnt_reg[4]/P0001 ,
		_w4386_
	);
	LUT4 #(
		.INIT('hf531)
	) name2637 (
		\u4_u3_csr0_reg[6]/P0001 ,
		\u4_u3_csr0_reg[7]/P0001 ,
		\u4_u3_dma_in_cnt_reg[4]/P0001 ,
		\u4_u3_dma_in_cnt_reg[5]/P0001 ,
		_w4387_
	);
	LUT2 #(
		.INIT('h2)
	) name2638 (
		\u4_u3_csr0_reg[4]/P0001 ,
		\u4_u3_dma_in_cnt_reg[2]/P0001 ,
		_w4388_
	);
	LUT4 #(
		.INIT('hf531)
	) name2639 (
		\u4_u3_csr0_reg[4]/P0001 ,
		\u4_u3_csr0_reg[5]/P0001 ,
		\u4_u3_dma_in_cnt_reg[2]/P0001 ,
		\u4_u3_dma_in_cnt_reg[3]/P0001 ,
		_w4389_
	);
	LUT4 #(
		.INIT('hb000)
	) name2640 (
		_w4384_,
		_w4385_,
		_w4387_,
		_w4389_,
		_w4390_
	);
	LUT4 #(
		.INIT('h8caf)
	) name2641 (
		\u4_u3_csr0_reg[5]/P0001 ,
		\u4_u3_csr0_reg[6]/P0001 ,
		\u4_u3_dma_in_cnt_reg[3]/P0001 ,
		\u4_u3_dma_in_cnt_reg[4]/P0001 ,
		_w4391_
	);
	LUT4 #(
		.INIT('h8caf)
	) name2642 (
		\u4_u3_csr0_reg[7]/P0001 ,
		\u4_u3_csr0_reg[8]/P0001 ,
		\u4_u3_dma_in_cnt_reg[5]/P0001 ,
		\u4_u3_dma_in_cnt_reg[6]/P0001 ,
		_w4392_
	);
	LUT3 #(
		.INIT('hd0)
	) name2643 (
		_w4387_,
		_w4391_,
		_w4392_,
		_w4393_
	);
	LUT4 #(
		.INIT('hf351)
	) name2644 (
		\u4_u3_csr0_reg[10]/P0001 ,
		\u4_u3_csr0_reg[9]/P0001 ,
		\u4_u3_dma_in_cnt_reg[7]/P0001 ,
		\u4_u3_dma_in_cnt_reg[8]/P0001 ,
		_w4394_
	);
	LUT2 #(
		.INIT('h2)
	) name2645 (
		\u4_u3_csr0_reg[8]/P0001 ,
		\u4_u3_dma_in_cnt_reg[6]/P0001 ,
		_w4395_
	);
	LUT2 #(
		.INIT('h2)
	) name2646 (
		_w4394_,
		_w4395_,
		_w4396_
	);
	LUT3 #(
		.INIT('hb0)
	) name2647 (
		_w4390_,
		_w4393_,
		_w4396_,
		_w4397_
	);
	LUT3 #(
		.INIT('h80)
	) name2648 (
		\u4_u3_dma_in_cnt_reg[4]/P0001 ,
		\u4_u3_dma_in_cnt_reg[5]/P0001 ,
		\u4_u3_dma_in_cnt_reg[6]/P0001 ,
		_w4398_
	);
	LUT4 #(
		.INIT('h8000)
	) name2649 (
		\u4_u3_dma_in_cnt_reg[0]/P0001 ,
		\u4_u3_dma_in_cnt_reg[1]/P0001 ,
		\u4_u3_dma_in_cnt_reg[2]/P0001 ,
		\u4_u3_dma_in_cnt_reg[3]/P0001 ,
		_w4399_
	);
	LUT2 #(
		.INIT('h8)
	) name2650 (
		\u4_u3_dma_in_cnt_reg[7]/P0001 ,
		\u4_u3_dma_in_cnt_reg[8]/P0001 ,
		_w4400_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name2651 (
		\u4_u3_r5_reg/NET0131 ,
		_w4398_,
		_w4399_,
		_w4400_,
		_w4401_
	);
	LUT3 #(
		.INIT('h01)
	) name2652 (
		\u1_u3_buf0_rl_reg/P0001 ,
		\u1_u3_buf0_set_reg/P0001 ,
		\u4_u3_set_r_reg/P0001 ,
		_w4402_
	);
	LUT3 #(
		.INIT('hb0)
	) name2653 (
		\u4_u3_csr0_reg[10]/P0001 ,
		\u4_u3_dma_in_cnt_reg[8]/P0001 ,
		\u4_u3_ep_match_r_reg/P0001 ,
		_w4403_
	);
	LUT4 #(
		.INIT('h3010)
	) name2654 (
		\u4_u3_csr0_reg[10]/P0001 ,
		\u4_u3_csr0_reg[9]/P0001 ,
		\u4_u3_dma_in_cnt_reg[7]/P0001 ,
		\u4_u3_dma_in_cnt_reg[8]/P0001 ,
		_w4404_
	);
	LUT3 #(
		.INIT('h04)
	) name2655 (
		_w4402_,
		_w4403_,
		_w4404_,
		_w4405_
	);
	LUT2 #(
		.INIT('h4)
	) name2656 (
		_w4401_,
		_w4405_,
		_w4406_
	);
	LUT3 #(
		.INIT('h80)
	) name2657 (
		\u4_u3_dma_in_cnt_reg[7]/P0001 ,
		\u4_u3_dma_in_cnt_reg[8]/P0001 ,
		\u4_u3_r5_reg/NET0131 ,
		_w4407_
	);
	LUT3 #(
		.INIT('h80)
	) name2658 (
		_w4398_,
		_w4399_,
		_w4407_,
		_w4408_
	);
	LUT2 #(
		.INIT('h8)
	) name2659 (
		\u4_u3_csr1_reg[0]/P0001 ,
		\u4_u3_dma_in_cnt_reg[9]/P0001 ,
		_w4409_
	);
	LUT4 #(
		.INIT('h7f00)
	) name2660 (
		_w4398_,
		_w4399_,
		_w4407_,
		_w4409_,
		_w4410_
	);
	LUT3 #(
		.INIT('hb0)
	) name2661 (
		_w4397_,
		_w4406_,
		_w4410_,
		_w4411_
	);
	LUT2 #(
		.INIT('h2)
	) name2662 (
		\u4_u3_csr1_reg[0]/P0001 ,
		\u4_u3_dma_in_cnt_reg[9]/P0001 ,
		_w4412_
	);
	LUT4 #(
		.INIT('hf400)
	) name2663 (
		_w4397_,
		_w4406_,
		_w4408_,
		_w4412_,
		_w4413_
	);
	LUT2 #(
		.INIT('he)
	) name2664 (
		_w4411_,
		_w4413_,
		_w4414_
	);
	LUT2 #(
		.INIT('h2)
	) name2665 (
		\u4_u0_csr0_reg[2]/P0001 ,
		\u4_u0_dma_in_cnt_reg[0]/P0001 ,
		_w4415_
	);
	LUT4 #(
		.INIT('hf531)
	) name2666 (
		\u4_u0_csr0_reg[2]/P0001 ,
		\u4_u0_csr0_reg[3]/NET0131 ,
		\u4_u0_dma_in_cnt_reg[0]/P0001 ,
		\u4_u0_dma_in_cnt_reg[1]/P0001 ,
		_w4416_
	);
	LUT4 #(
		.INIT('h8caf)
	) name2667 (
		\u4_u0_csr0_reg[3]/NET0131 ,
		\u4_u0_csr0_reg[4]/P0001 ,
		\u4_u0_dma_in_cnt_reg[1]/P0001 ,
		\u4_u0_dma_in_cnt_reg[2]/P0001 ,
		_w4417_
	);
	LUT2 #(
		.INIT('h2)
	) name2668 (
		\u4_u0_csr0_reg[6]/P0001 ,
		\u4_u0_dma_in_cnt_reg[4]/P0001 ,
		_w4418_
	);
	LUT4 #(
		.INIT('hf531)
	) name2669 (
		\u4_u0_csr0_reg[6]/P0001 ,
		\u4_u0_csr0_reg[7]/P0001 ,
		\u4_u0_dma_in_cnt_reg[4]/P0001 ,
		\u4_u0_dma_in_cnt_reg[5]/P0001 ,
		_w4419_
	);
	LUT2 #(
		.INIT('h2)
	) name2670 (
		\u4_u0_csr0_reg[4]/P0001 ,
		\u4_u0_dma_in_cnt_reg[2]/P0001 ,
		_w4420_
	);
	LUT4 #(
		.INIT('hf531)
	) name2671 (
		\u4_u0_csr0_reg[4]/P0001 ,
		\u4_u0_csr0_reg[5]/P0001 ,
		\u4_u0_dma_in_cnt_reg[2]/P0001 ,
		\u4_u0_dma_in_cnt_reg[3]/P0001 ,
		_w4421_
	);
	LUT4 #(
		.INIT('hb000)
	) name2672 (
		_w4416_,
		_w4417_,
		_w4419_,
		_w4421_,
		_w4422_
	);
	LUT4 #(
		.INIT('h8caf)
	) name2673 (
		\u4_u0_csr0_reg[5]/P0001 ,
		\u4_u0_csr0_reg[6]/P0001 ,
		\u4_u0_dma_in_cnt_reg[3]/P0001 ,
		\u4_u0_dma_in_cnt_reg[4]/P0001 ,
		_w4423_
	);
	LUT4 #(
		.INIT('h8caf)
	) name2674 (
		\u4_u0_csr0_reg[7]/P0001 ,
		\u4_u0_csr0_reg[8]/P0001 ,
		\u4_u0_dma_in_cnt_reg[5]/P0001 ,
		\u4_u0_dma_in_cnt_reg[6]/P0001 ,
		_w4424_
	);
	LUT3 #(
		.INIT('hd0)
	) name2675 (
		_w4419_,
		_w4423_,
		_w4424_,
		_w4425_
	);
	LUT4 #(
		.INIT('hf351)
	) name2676 (
		\u4_u0_csr0_reg[10]/P0001 ,
		\u4_u0_csr0_reg[9]/P0001 ,
		\u4_u0_dma_in_cnt_reg[7]/P0001 ,
		\u4_u0_dma_in_cnt_reg[8]/P0001 ,
		_w4426_
	);
	LUT2 #(
		.INIT('h2)
	) name2677 (
		\u4_u0_csr0_reg[8]/P0001 ,
		\u4_u0_dma_in_cnt_reg[6]/P0001 ,
		_w4427_
	);
	LUT2 #(
		.INIT('h2)
	) name2678 (
		_w4426_,
		_w4427_,
		_w4428_
	);
	LUT3 #(
		.INIT('hb0)
	) name2679 (
		_w4422_,
		_w4425_,
		_w4428_,
		_w4429_
	);
	LUT3 #(
		.INIT('h80)
	) name2680 (
		\u4_u0_dma_in_cnt_reg[4]/P0001 ,
		\u4_u0_dma_in_cnt_reg[5]/P0001 ,
		\u4_u0_dma_in_cnt_reg[6]/P0001 ,
		_w4430_
	);
	LUT4 #(
		.INIT('h8000)
	) name2681 (
		\u4_u0_dma_in_cnt_reg[0]/P0001 ,
		\u4_u0_dma_in_cnt_reg[1]/P0001 ,
		\u4_u0_dma_in_cnt_reg[2]/P0001 ,
		\u4_u0_dma_in_cnt_reg[3]/P0001 ,
		_w4431_
	);
	LUT2 #(
		.INIT('h8)
	) name2682 (
		\u4_u0_dma_in_cnt_reg[7]/P0001 ,
		\u4_u0_dma_in_cnt_reg[8]/P0001 ,
		_w4432_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name2683 (
		\u4_u0_r5_reg/NET0131 ,
		_w4430_,
		_w4431_,
		_w4432_,
		_w4433_
	);
	LUT3 #(
		.INIT('h01)
	) name2684 (
		\u1_u3_buf0_rl_reg/P0001 ,
		\u1_u3_buf0_set_reg/P0001 ,
		\u4_u0_set_r_reg/P0001 ,
		_w4434_
	);
	LUT3 #(
		.INIT('hb0)
	) name2685 (
		\u4_u0_csr0_reg[10]/P0001 ,
		\u4_u0_dma_in_cnt_reg[8]/P0001 ,
		\u4_u0_ep_match_r_reg/P0001 ,
		_w4435_
	);
	LUT4 #(
		.INIT('h3010)
	) name2686 (
		\u4_u0_csr0_reg[10]/P0001 ,
		\u4_u0_csr0_reg[9]/P0001 ,
		\u4_u0_dma_in_cnt_reg[7]/P0001 ,
		\u4_u0_dma_in_cnt_reg[8]/P0001 ,
		_w4436_
	);
	LUT3 #(
		.INIT('h04)
	) name2687 (
		_w4434_,
		_w4435_,
		_w4436_,
		_w4437_
	);
	LUT2 #(
		.INIT('h4)
	) name2688 (
		_w4433_,
		_w4437_,
		_w4438_
	);
	LUT3 #(
		.INIT('h80)
	) name2689 (
		\u4_u0_dma_in_cnt_reg[7]/P0001 ,
		\u4_u0_dma_in_cnt_reg[8]/P0001 ,
		\u4_u0_r5_reg/NET0131 ,
		_w4439_
	);
	LUT3 #(
		.INIT('h80)
	) name2690 (
		_w4430_,
		_w4431_,
		_w4439_,
		_w4440_
	);
	LUT2 #(
		.INIT('h8)
	) name2691 (
		\u4_u0_csr1_reg[0]/P0001 ,
		\u4_u0_dma_in_cnt_reg[9]/P0001 ,
		_w4441_
	);
	LUT4 #(
		.INIT('h7f00)
	) name2692 (
		_w4430_,
		_w4431_,
		_w4439_,
		_w4441_,
		_w4442_
	);
	LUT3 #(
		.INIT('hb0)
	) name2693 (
		_w4429_,
		_w4438_,
		_w4442_,
		_w4443_
	);
	LUT2 #(
		.INIT('h2)
	) name2694 (
		\u4_u0_csr1_reg[0]/P0001 ,
		\u4_u0_dma_in_cnt_reg[9]/P0001 ,
		_w4444_
	);
	LUT4 #(
		.INIT('hf400)
	) name2695 (
		_w4429_,
		_w4438_,
		_w4440_,
		_w4444_,
		_w4445_
	);
	LUT2 #(
		.INIT('he)
	) name2696 (
		_w4443_,
		_w4445_,
		_w4446_
	);
	LUT3 #(
		.INIT('h80)
	) name2697 (
		\u4_u1_dma_in_cnt_reg[4]/P0001 ,
		\u4_u1_dma_in_cnt_reg[5]/P0001 ,
		\u4_u1_dma_in_cnt_reg[6]/P0001 ,
		_w4447_
	);
	LUT4 #(
		.INIT('h8000)
	) name2698 (
		\u4_u1_dma_in_cnt_reg[0]/P0001 ,
		\u4_u1_dma_in_cnt_reg[1]/P0001 ,
		\u4_u1_dma_in_cnt_reg[2]/P0001 ,
		\u4_u1_dma_in_cnt_reg[3]/P0001 ,
		_w4448_
	);
	LUT2 #(
		.INIT('h8)
	) name2699 (
		\u4_u1_dma_in_cnt_reg[7]/P0001 ,
		\u4_u1_dma_in_cnt_reg[8]/P0001 ,
		_w4449_
	);
	LUT3 #(
		.INIT('h80)
	) name2700 (
		\u4_u1_dma_in_cnt_reg[7]/P0001 ,
		\u4_u1_dma_in_cnt_reg[8]/P0001 ,
		\u4_u1_r5_reg/NET0131 ,
		_w4450_
	);
	LUT3 #(
		.INIT('h80)
	) name2701 (
		_w4447_,
		_w4448_,
		_w4450_,
		_w4451_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name2702 (
		\u4_u1_r5_reg/NET0131 ,
		_w4447_,
		_w4448_,
		_w4449_,
		_w4452_
	);
	LUT3 #(
		.INIT('h01)
	) name2703 (
		\u1_u3_buf0_rl_reg/P0001 ,
		\u1_u3_buf0_set_reg/P0001 ,
		\u4_u1_set_r_reg/P0001 ,
		_w4453_
	);
	LUT4 #(
		.INIT('hf0e0)
	) name2704 (
		\u1_u3_buf0_rl_reg/P0001 ,
		\u1_u3_buf0_set_reg/P0001 ,
		\u4_u1_ep_match_r_reg/P0001 ,
		\u4_u1_set_r_reg/P0001 ,
		_w4454_
	);
	LUT4 #(
		.INIT('h3010)
	) name2705 (
		\u4_u1_csr0_reg[10]/P0001 ,
		\u4_u1_csr0_reg[9]/P0001 ,
		\u4_u1_dma_in_cnt_reg[7]/P0001 ,
		\u4_u1_dma_in_cnt_reg[8]/P0001 ,
		_w4455_
	);
	LUT4 #(
		.INIT('h8aef)
	) name2706 (
		\u4_u1_csr0_reg[10]/P0001 ,
		\u4_u1_csr0_reg[9]/P0001 ,
		\u4_u1_dma_in_cnt_reg[7]/P0001 ,
		\u4_u1_dma_in_cnt_reg[8]/P0001 ,
		_w4456_
	);
	LUT2 #(
		.INIT('h8)
	) name2707 (
		_w4454_,
		_w4456_,
		_w4457_
	);
	LUT3 #(
		.INIT('h45)
	) name2708 (
		_w4451_,
		_w4452_,
		_w4457_,
		_w4458_
	);
	LUT2 #(
		.INIT('h4)
	) name2709 (
		\u4_u1_csr0_reg[8]/P0001 ,
		\u4_u1_dma_in_cnt_reg[6]/P0001 ,
		_w4459_
	);
	LUT2 #(
		.INIT('h2)
	) name2710 (
		\u4_u1_csr0_reg[7]/P0001 ,
		\u4_u1_dma_in_cnt_reg[5]/P0001 ,
		_w4460_
	);
	LUT4 #(
		.INIT('h080a)
	) name2711 (
		\u4_u1_csr0_reg[7]/P0001 ,
		\u4_u1_csr0_reg[8]/P0001 ,
		\u4_u1_dma_in_cnt_reg[5]/P0001 ,
		\u4_u1_dma_in_cnt_reg[6]/P0001 ,
		_w4461_
	);
	LUT4 #(
		.INIT('hf531)
	) name2712 (
		\u4_u1_csr0_reg[5]/P0001 ,
		\u4_u1_csr0_reg[6]/P0001 ,
		\u4_u1_dma_in_cnt_reg[3]/P0001 ,
		\u4_u1_dma_in_cnt_reg[4]/P0001 ,
		_w4462_
	);
	LUT4 #(
		.INIT('h5010)
	) name2713 (
		\u4_u1_csr0_reg[5]/P0001 ,
		\u4_u1_csr0_reg[6]/P0001 ,
		\u4_u1_dma_in_cnt_reg[3]/P0001 ,
		\u4_u1_dma_in_cnt_reg[4]/P0001 ,
		_w4463_
	);
	LUT2 #(
		.INIT('h2)
	) name2714 (
		\u4_u1_csr0_reg[2]/P0001 ,
		\u4_u1_dma_in_cnt_reg[0]/P0001 ,
		_w4464_
	);
	LUT4 #(
		.INIT('hf531)
	) name2715 (
		\u4_u1_csr0_reg[2]/P0001 ,
		\u4_u1_csr0_reg[3]/NET0131 ,
		\u4_u1_dma_in_cnt_reg[0]/P0001 ,
		\u4_u1_dma_in_cnt_reg[1]/P0001 ,
		_w4465_
	);
	LUT4 #(
		.INIT('h8caf)
	) name2716 (
		\u4_u1_csr0_reg[3]/NET0131 ,
		\u4_u1_csr0_reg[4]/P0001 ,
		\u4_u1_dma_in_cnt_reg[1]/P0001 ,
		\u4_u1_dma_in_cnt_reg[2]/P0001 ,
		_w4466_
	);
	LUT2 #(
		.INIT('h2)
	) name2717 (
		\u4_u1_csr0_reg[4]/P0001 ,
		\u4_u1_dma_in_cnt_reg[2]/P0001 ,
		_w4467_
	);
	LUT4 #(
		.INIT('h008a)
	) name2718 (
		_w4462_,
		_w4465_,
		_w4466_,
		_w4467_,
		_w4468_
	);
	LUT4 #(
		.INIT('h8caf)
	) name2719 (
		\u4_u1_csr0_reg[6]/P0001 ,
		\u4_u1_csr0_reg[7]/P0001 ,
		\u4_u1_dma_in_cnt_reg[4]/P0001 ,
		\u4_u1_dma_in_cnt_reg[5]/P0001 ,
		_w4469_
	);
	LUT2 #(
		.INIT('h4)
	) name2720 (
		_w4459_,
		_w4469_,
		_w4470_
	);
	LUT4 #(
		.INIT('h5455)
	) name2721 (
		_w4461_,
		_w4463_,
		_w4468_,
		_w4470_,
		_w4471_
	);
	LUT2 #(
		.INIT('h2)
	) name2722 (
		\u4_u1_csr0_reg[9]/P0001 ,
		\u4_u1_dma_in_cnt_reg[7]/P0001 ,
		_w4472_
	);
	LUT4 #(
		.INIT('hf351)
	) name2723 (
		\u4_u1_csr0_reg[10]/P0001 ,
		\u4_u1_csr0_reg[9]/P0001 ,
		\u4_u1_dma_in_cnt_reg[7]/P0001 ,
		\u4_u1_dma_in_cnt_reg[8]/P0001 ,
		_w4473_
	);
	LUT2 #(
		.INIT('h2)
	) name2724 (
		\u4_u1_csr0_reg[8]/P0001 ,
		\u4_u1_dma_in_cnt_reg[6]/P0001 ,
		_w4474_
	);
	LUT2 #(
		.INIT('h2)
	) name2725 (
		_w4473_,
		_w4474_,
		_w4475_
	);
	LUT2 #(
		.INIT('h4)
	) name2726 (
		_w4451_,
		_w4475_,
		_w4476_
	);
	LUT2 #(
		.INIT('h8)
	) name2727 (
		\u4_u1_csr1_reg[0]/P0001 ,
		\u4_u1_dma_in_cnt_reg[9]/P0001 ,
		_w4477_
	);
	LUT4 #(
		.INIT('hea00)
	) name2728 (
		_w4458_,
		_w4471_,
		_w4476_,
		_w4477_,
		_w4478_
	);
	LUT2 #(
		.INIT('h2)
	) name2729 (
		\u4_u1_csr1_reg[0]/P0001 ,
		\u4_u1_dma_in_cnt_reg[9]/P0001 ,
		_w4479_
	);
	LUT4 #(
		.INIT('h1500)
	) name2730 (
		_w4458_,
		_w4471_,
		_w4476_,
		_w4479_,
		_w4480_
	);
	LUT2 #(
		.INIT('he)
	) name2731 (
		_w4478_,
		_w4480_,
		_w4481_
	);
	LUT3 #(
		.INIT('h01)
	) name2732 (
		\u1_u3_buf0_rl_reg/P0001 ,
		\u1_u3_buf0_set_reg/P0001 ,
		\u4_u2_set_r_reg/P0001 ,
		_w4482_
	);
	LUT3 #(
		.INIT('h20)
	) name2733 (
		\u4_u2_csr0_reg[10]/P0001 ,
		\u4_u2_dma_in_cnt_reg[8]/P0001 ,
		\u4_u2_ep_match_r_reg/P0001 ,
		_w4483_
	);
	LUT3 #(
		.INIT('hb0)
	) name2734 (
		\u4_u2_csr0_reg[10]/P0001 ,
		\u4_u2_dma_in_cnt_reg[8]/P0001 ,
		\u4_u2_ep_match_r_reg/P0001 ,
		_w4484_
	);
	LUT2 #(
		.INIT('h4)
	) name2735 (
		\u4_u2_csr0_reg[9]/P0001 ,
		\u4_u2_dma_in_cnt_reg[7]/P0001 ,
		_w4485_
	);
	LUT4 #(
		.INIT('hbbab)
	) name2736 (
		_w4482_,
		_w4483_,
		_w4484_,
		_w4485_,
		_w4486_
	);
	LUT2 #(
		.INIT('h4)
	) name2737 (
		\u4_u2_csr0_reg[8]/P0001 ,
		\u4_u2_dma_in_cnt_reg[6]/P0001 ,
		_w4487_
	);
	LUT2 #(
		.INIT('h2)
	) name2738 (
		\u4_u2_csr0_reg[7]/P0001 ,
		\u4_u2_dma_in_cnt_reg[5]/P0001 ,
		_w4488_
	);
	LUT4 #(
		.INIT('h080a)
	) name2739 (
		\u4_u2_csr0_reg[7]/P0001 ,
		\u4_u2_csr0_reg[8]/P0001 ,
		\u4_u2_dma_in_cnt_reg[5]/P0001 ,
		\u4_u2_dma_in_cnt_reg[6]/P0001 ,
		_w4489_
	);
	LUT4 #(
		.INIT('hf531)
	) name2740 (
		\u4_u2_csr0_reg[5]/P0001 ,
		\u4_u2_csr0_reg[6]/P0001 ,
		\u4_u2_dma_in_cnt_reg[3]/P0001 ,
		\u4_u2_dma_in_cnt_reg[4]/P0001 ,
		_w4490_
	);
	LUT4 #(
		.INIT('h5010)
	) name2741 (
		\u4_u2_csr0_reg[5]/P0001 ,
		\u4_u2_csr0_reg[6]/P0001 ,
		\u4_u2_dma_in_cnt_reg[3]/P0001 ,
		\u4_u2_dma_in_cnt_reg[4]/P0001 ,
		_w4491_
	);
	LUT2 #(
		.INIT('h2)
	) name2742 (
		\u4_u2_csr0_reg[2]/P0001 ,
		\u4_u2_dma_in_cnt_reg[0]/P0001 ,
		_w4492_
	);
	LUT4 #(
		.INIT('hf531)
	) name2743 (
		\u4_u2_csr0_reg[2]/P0001 ,
		\u4_u2_csr0_reg[3]/NET0131 ,
		\u4_u2_dma_in_cnt_reg[0]/P0001 ,
		\u4_u2_dma_in_cnt_reg[1]/P0001 ,
		_w4493_
	);
	LUT4 #(
		.INIT('h8caf)
	) name2744 (
		\u4_u2_csr0_reg[3]/NET0131 ,
		\u4_u2_csr0_reg[4]/P0001 ,
		\u4_u2_dma_in_cnt_reg[1]/P0001 ,
		\u4_u2_dma_in_cnt_reg[2]/P0001 ,
		_w4494_
	);
	LUT2 #(
		.INIT('h2)
	) name2745 (
		\u4_u2_csr0_reg[4]/P0001 ,
		\u4_u2_dma_in_cnt_reg[2]/P0001 ,
		_w4495_
	);
	LUT4 #(
		.INIT('h008a)
	) name2746 (
		_w4490_,
		_w4493_,
		_w4494_,
		_w4495_,
		_w4496_
	);
	LUT4 #(
		.INIT('h8caf)
	) name2747 (
		\u4_u2_csr0_reg[6]/P0001 ,
		\u4_u2_csr0_reg[7]/P0001 ,
		\u4_u2_dma_in_cnt_reg[4]/P0001 ,
		\u4_u2_dma_in_cnt_reg[5]/P0001 ,
		_w4497_
	);
	LUT2 #(
		.INIT('h4)
	) name2748 (
		_w4487_,
		_w4497_,
		_w4498_
	);
	LUT4 #(
		.INIT('h5455)
	) name2749 (
		_w4489_,
		_w4491_,
		_w4496_,
		_w4498_,
		_w4499_
	);
	LUT4 #(
		.INIT('hf531)
	) name2750 (
		\u4_u2_csr0_reg[8]/P0001 ,
		\u4_u2_csr0_reg[9]/P0001 ,
		\u4_u2_dma_in_cnt_reg[6]/P0001 ,
		\u4_u2_dma_in_cnt_reg[7]/P0001 ,
		_w4500_
	);
	LUT3 #(
		.INIT('hb0)
	) name2751 (
		_w4482_,
		_w4483_,
		_w4500_,
		_w4501_
	);
	LUT4 #(
		.INIT('h5444)
	) name2752 (
		\u4_u2_r5_reg/NET0131 ,
		_w4486_,
		_w4499_,
		_w4501_,
		_w4502_
	);
	LUT2 #(
		.INIT('h2)
	) name2753 (
		\u4_u2_dma_in_cnt_reg[9]/P0001 ,
		\u4_u2_r5_reg/NET0131 ,
		_w4503_
	);
	LUT3 #(
		.INIT('h80)
	) name2754 (
		\u4_u2_dma_in_cnt_reg[4]/P0001 ,
		\u4_u2_dma_in_cnt_reg[5]/P0001 ,
		\u4_u2_dma_in_cnt_reg[6]/P0001 ,
		_w4504_
	);
	LUT4 #(
		.INIT('h8000)
	) name2755 (
		\u4_u2_dma_in_cnt_reg[0]/P0001 ,
		\u4_u2_dma_in_cnt_reg[1]/P0001 ,
		\u4_u2_dma_in_cnt_reg[2]/P0001 ,
		\u4_u2_dma_in_cnt_reg[3]/P0001 ,
		_w4505_
	);
	LUT2 #(
		.INIT('h8)
	) name2756 (
		\u4_u2_dma_in_cnt_reg[7]/P0001 ,
		\u4_u2_dma_in_cnt_reg[8]/P0001 ,
		_w4506_
	);
	LUT3 #(
		.INIT('h80)
	) name2757 (
		\u4_u2_dma_in_cnt_reg[7]/P0001 ,
		\u4_u2_dma_in_cnt_reg[8]/P0001 ,
		\u4_u2_dma_in_cnt_reg[9]/P0001 ,
		_w4507_
	);
	LUT4 #(
		.INIT('h1555)
	) name2758 (
		_w4503_,
		_w4504_,
		_w4505_,
		_w4507_,
		_w4508_
	);
	LUT2 #(
		.INIT('h1)
	) name2759 (
		\u4_u2_dma_in_cnt_reg[9]/P0001 ,
		\u4_u2_r5_reg/NET0131 ,
		_w4509_
	);
	LUT4 #(
		.INIT('hea00)
	) name2760 (
		_w4486_,
		_w4499_,
		_w4501_,
		_w4509_,
		_w4510_
	);
	LUT2 #(
		.INIT('h4)
	) name2761 (
		\u4_u2_dma_in_cnt_reg[9]/P0001 ,
		\u4_u2_r5_reg/NET0131 ,
		_w4511_
	);
	LUT4 #(
		.INIT('h7f00)
	) name2762 (
		_w4504_,
		_w4505_,
		_w4506_,
		_w4511_,
		_w4512_
	);
	LUT2 #(
		.INIT('h2)
	) name2763 (
		\u4_u2_csr1_reg[0]/P0001 ,
		_w4512_,
		_w4513_
	);
	LUT4 #(
		.INIT('h0e00)
	) name2764 (
		_w4502_,
		_w4508_,
		_w4510_,
		_w4513_,
		_w4514_
	);
	LUT3 #(
		.INIT('h02)
	) name2765 (
		rst_i_pad,
		\u1_clr_sof_time_reg/P0001 ,
		\u1_hms_clk_reg/P0001 ,
		_w4515_
	);
	LUT2 #(
		.INIT('h1)
	) name2766 (
		\u1_hms_cnt_reg[0]/P0001 ,
		\u1_hms_cnt_reg[1]/P0001 ,
		_w4516_
	);
	LUT2 #(
		.INIT('h6)
	) name2767 (
		\u1_hms_cnt_reg[0]/P0001 ,
		\u1_hms_cnt_reg[1]/P0001 ,
		_w4517_
	);
	LUT2 #(
		.INIT('h8)
	) name2768 (
		_w4515_,
		_w4517_,
		_w4518_
	);
	LUT3 #(
		.INIT('h78)
	) name2769 (
		\u1_hms_cnt_reg[0]/P0001 ,
		\u1_hms_cnt_reg[1]/P0001 ,
		\u1_hms_cnt_reg[2]/P0001 ,
		_w4519_
	);
	LUT2 #(
		.INIT('h8)
	) name2770 (
		_w4515_,
		_w4519_,
		_w4520_
	);
	LUT4 #(
		.INIT('h007f)
	) name2771 (
		\u1_hms_cnt_reg[0]/P0001 ,
		\u1_hms_cnt_reg[1]/P0001 ,
		\u1_hms_cnt_reg[2]/P0001 ,
		\u1_hms_cnt_reg[3]/P0001 ,
		_w4521_
	);
	LUT4 #(
		.INIT('h8000)
	) name2772 (
		\u1_hms_cnt_reg[0]/P0001 ,
		\u1_hms_cnt_reg[1]/P0001 ,
		\u1_hms_cnt_reg[2]/P0001 ,
		\u1_hms_cnt_reg[3]/P0001 ,
		_w4522_
	);
	LUT3 #(
		.INIT('h02)
	) name2773 (
		_w4515_,
		_w4521_,
		_w4522_,
		_w4523_
	);
	LUT4 #(
		.INIT('h0200)
	) name2774 (
		rst_i_pad,
		\u1_clr_sof_time_reg/P0001 ,
		\u1_hms_clk_reg/P0001 ,
		\u1_hms_cnt_reg[4]/P0001 ,
		_w4524_
	);
	LUT4 #(
		.INIT('h0002)
	) name2775 (
		rst_i_pad,
		\u1_clr_sof_time_reg/P0001 ,
		\u1_hms_clk_reg/P0001 ,
		\u1_hms_cnt_reg[4]/P0001 ,
		_w4525_
	);
	LUT3 #(
		.INIT('he4)
	) name2776 (
		_w4522_,
		_w4524_,
		_w4525_,
		_w4526_
	);
	LUT3 #(
		.INIT('h2a)
	) name2777 (
		\u1_u0_token_valid_str1_reg/P0001 ,
		_w3740_,
		_w3748_,
		_w4527_
	);
	LUT4 #(
		.INIT('hc444)
	) name2778 (
		\u1_u0_token_valid_str1_reg/P0001 ,
		_w3717_,
		_w3740_,
		_w3748_,
		_w4528_
	);
	LUT4 #(
		.INIT('ha820)
	) name2779 (
		rst_i_pad,
		\u1_clr_sof_time_reg/P0001 ,
		\u1_frame_no_r_reg[0]/P0001 ,
		\u1_u0_token0_reg[0]/NET0131 ,
		_w4529_
	);
	LUT4 #(
		.INIT('ha820)
	) name2780 (
		rst_i_pad,
		\u1_clr_sof_time_reg/P0001 ,
		\u1_frame_no_r_reg[10]/P0001 ,
		\u1_u0_token1_reg[2]/P0001 ,
		_w4530_
	);
	LUT4 #(
		.INIT('ha820)
	) name2781 (
		rst_i_pad,
		\u1_clr_sof_time_reg/P0001 ,
		\u1_frame_no_r_reg[1]/P0001 ,
		\u1_u0_token0_reg[1]/P0001 ,
		_w4531_
	);
	LUT4 #(
		.INIT('ha820)
	) name2782 (
		rst_i_pad,
		\u1_clr_sof_time_reg/P0001 ,
		\u1_frame_no_r_reg[3]/P0001 ,
		\u1_u0_token0_reg[3]/NET0131 ,
		_w4532_
	);
	LUT4 #(
		.INIT('ha820)
	) name2783 (
		rst_i_pad,
		\u1_clr_sof_time_reg/P0001 ,
		\u1_frame_no_r_reg[2]/P0001 ,
		\u1_u0_token0_reg[2]/NET0131 ,
		_w4533_
	);
	LUT4 #(
		.INIT('ha820)
	) name2784 (
		rst_i_pad,
		\u1_clr_sof_time_reg/P0001 ,
		\u1_frame_no_r_reg[4]/P0001 ,
		\u1_u0_token0_reg[4]/P0001 ,
		_w4534_
	);
	LUT4 #(
		.INIT('ha820)
	) name2785 (
		rst_i_pad,
		\u1_clr_sof_time_reg/P0001 ,
		\u1_frame_no_r_reg[5]/P0001 ,
		\u1_u0_token0_reg[5]/NET0131 ,
		_w4535_
	);
	LUT4 #(
		.INIT('ha820)
	) name2786 (
		rst_i_pad,
		\u1_clr_sof_time_reg/P0001 ,
		\u1_frame_no_r_reg[6]/P0001 ,
		\u1_u0_token0_reg[6]/P0001 ,
		_w4536_
	);
	LUT4 #(
		.INIT('ha820)
	) name2787 (
		rst_i_pad,
		\u1_clr_sof_time_reg/P0001 ,
		\u1_frame_no_r_reg[7]/P0001 ,
		\u1_u0_token0_reg[7]/P0001 ,
		_w4537_
	);
	LUT4 #(
		.INIT('ha820)
	) name2788 (
		rst_i_pad,
		\u1_clr_sof_time_reg/P0001 ,
		\u1_frame_no_r_reg[8]/P0001 ,
		\u1_u0_token1_reg[0]/P0001 ,
		_w4538_
	);
	LUT4 #(
		.INIT('ha820)
	) name2789 (
		rst_i_pad,
		\u1_clr_sof_time_reg/P0001 ,
		\u1_frame_no_r_reg[9]/P0001 ,
		\u1_u0_token1_reg[1]/P0001 ,
		_w4539_
	);
	LUT3 #(
		.INIT('hac)
	) name2790 (
		\u1_u2_sizu_c_reg[4]/P0001 ,
		\u1_u3_new_size_reg[4]/P0001 ,
		\u1_u3_out_to_small_r_reg/P0001 ,
		_w4540_
	);
	LUT3 #(
		.INIT('hac)
	) name2791 (
		\u1_u2_sizu_c_reg[5]/P0001 ,
		\u1_u3_new_size_reg[5]/P0001 ,
		\u1_u3_out_to_small_r_reg/P0001 ,
		_w4541_
	);
	LUT3 #(
		.INIT('hac)
	) name2792 (
		\u1_u2_sizu_c_reg[6]/P0001 ,
		\u1_u3_new_size_reg[6]/P0001 ,
		\u1_u3_out_to_small_r_reg/P0001 ,
		_w4542_
	);
	LUT3 #(
		.INIT('hac)
	) name2793 (
		\u1_u2_sizu_c_reg[7]/P0001 ,
		\u1_u3_new_size_reg[7]/P0001 ,
		\u1_u3_out_to_small_r_reg/P0001 ,
		_w4543_
	);
	LUT3 #(
		.INIT('h59)
	) name2794 (
		\u1_u3_adr_reg[6]/P0001 ,
		_w2860_,
		_w2862_,
		_w4544_
	);
	LUT2 #(
		.INIT('h2)
	) name2795 (
		_w4204_,
		_w4207_,
		_w4545_
	);
	LUT4 #(
		.INIT('h004d)
	) name2796 (
		\u1_u3_adr_reg[5]/P0001 ,
		_w2823_,
		_w4077_,
		_w4078_,
		_w4546_
	);
	LUT3 #(
		.INIT('he0)
	) name2797 (
		_w4073_,
		_w4075_,
		_w4546_,
		_w4547_
	);
	LUT3 #(
		.INIT('ha9)
	) name2798 (
		_w4544_,
		_w4545_,
		_w4547_,
		_w4548_
	);
	LUT3 #(
		.INIT('h59)
	) name2799 (
		\u1_u3_adr_reg[8]/P0001 ,
		_w2837_,
		_w2839_,
		_w4549_
	);
	LUT4 #(
		.INIT('h45ba)
	) name2800 (
		_w4205_,
		_w4206_,
		_w4208_,
		_w4549_,
		_w4550_
	);
	LUT2 #(
		.INIT('h8)
	) name2801 (
		\u4_u3_csr1_reg[0]/P0001 ,
		\u4_u3_dma_in_cnt_reg[8]/P0001 ,
		_w4551_
	);
	LUT2 #(
		.INIT('h8)
	) name2802 (
		\u4_u3_csr1_reg[0]/P0001 ,
		\u4_u3_dma_in_cnt_reg[7]/P0001 ,
		_w4552_
	);
	LUT4 #(
		.INIT('h070f)
	) name2803 (
		_w4398_,
		_w4399_,
		_w4551_,
		_w4552_,
		_w4553_
	);
	LUT2 #(
		.INIT('h2)
	) name2804 (
		_w4401_,
		_w4553_,
		_w4554_
	);
	LUT4 #(
		.INIT('h0001)
	) name2805 (
		\u1_u3_buf0_rl_reg/P0001 ,
		\u1_u3_buf0_set_reg/P0001 ,
		\u4_u3_dma_in_cnt_reg[8]/P0001 ,
		\u4_u3_set_r_reg/P0001 ,
		_w4555_
	);
	LUT4 #(
		.INIT('h00a8)
	) name2806 (
		\u4_u3_csr1_reg[0]/P0001 ,
		\u4_u3_dma_in_cnt_reg[8]/P0001 ,
		\u4_u3_ep_match_r_reg/P0001 ,
		\u4_u3_r5_reg/NET0131 ,
		_w4556_
	);
	LUT2 #(
		.INIT('h4)
	) name2807 (
		_w4555_,
		_w4556_,
		_w4557_
	);
	LUT2 #(
		.INIT('h9)
	) name2808 (
		\u4_u3_csr0_reg[10]/P0001 ,
		\u4_u3_dma_in_cnt_reg[8]/P0001 ,
		_w4558_
	);
	LUT4 #(
		.INIT('h7310)
	) name2809 (
		\u4_u3_csr0_reg[4]/P0001 ,
		\u4_u3_csr0_reg[5]/P0001 ,
		\u4_u3_dma_in_cnt_reg[2]/P0001 ,
		\u4_u3_dma_in_cnt_reg[3]/P0001 ,
		_w4559_
	);
	LUT4 #(
		.INIT('h08ce)
	) name2810 (
		\u4_u3_csr0_reg[2]/P0001 ,
		\u4_u3_csr0_reg[3]/NET0131 ,
		\u4_u3_dma_in_cnt_reg[0]/P0001 ,
		\u4_u3_dma_in_cnt_reg[1]/P0001 ,
		_w4560_
	);
	LUT4 #(
		.INIT('h5f57)
	) name2811 (
		_w4387_,
		_w4389_,
		_w4559_,
		_w4560_,
		_w4561_
	);
	LUT4 #(
		.INIT('h8caf)
	) name2812 (
		\u4_u3_csr0_reg[8]/P0001 ,
		\u4_u3_csr0_reg[9]/P0001 ,
		\u4_u3_dma_in_cnt_reg[6]/P0001 ,
		\u4_u3_dma_in_cnt_reg[7]/P0001 ,
		_w4562_
	);
	LUT4 #(
		.INIT('h8caf)
	) name2813 (
		\u4_u3_csr0_reg[6]/P0001 ,
		\u4_u3_csr0_reg[7]/P0001 ,
		\u4_u3_dma_in_cnt_reg[4]/P0001 ,
		\u4_u3_dma_in_cnt_reg[5]/P0001 ,
		_w4563_
	);
	LUT4 #(
		.INIT('h7310)
	) name2814 (
		\u4_u3_csr0_reg[6]/P0001 ,
		\u4_u3_csr0_reg[7]/P0001 ,
		\u4_u3_dma_in_cnt_reg[4]/P0001 ,
		\u4_u3_dma_in_cnt_reg[5]/P0001 ,
		_w4564_
	);
	LUT2 #(
		.INIT('h2)
	) name2815 (
		_w4562_,
		_w4564_,
		_w4565_
	);
	LUT4 #(
		.INIT('h080a)
	) name2816 (
		\u4_u3_csr0_reg[8]/P0001 ,
		\u4_u3_csr0_reg[9]/P0001 ,
		\u4_u3_dma_in_cnt_reg[6]/P0001 ,
		\u4_u3_dma_in_cnt_reg[7]/P0001 ,
		_w4566_
	);
	LUT4 #(
		.INIT('hf731)
	) name2817 (
		\u4_u3_csr0_reg[8]/P0001 ,
		\u4_u3_csr0_reg[9]/P0001 ,
		\u4_u3_dma_in_cnt_reg[6]/P0001 ,
		\u4_u3_dma_in_cnt_reg[7]/P0001 ,
		_w4567_
	);
	LUT4 #(
		.INIT('h80aa)
	) name2818 (
		_w4558_,
		_w4561_,
		_w4565_,
		_w4567_,
		_w4568_
	);
	LUT4 #(
		.INIT('hf0e0)
	) name2819 (
		\u1_u3_buf0_rl_reg/P0001 ,
		\u1_u3_buf0_set_reg/P0001 ,
		\u4_u3_ep_match_r_reg/P0001 ,
		\u4_u3_set_r_reg/P0001 ,
		_w4569_
	);
	LUT2 #(
		.INIT('h4)
	) name2820 (
		_w4558_,
		_w4567_,
		_w4570_
	);
	LUT4 #(
		.INIT('h80f0)
	) name2821 (
		_w4561_,
		_w4565_,
		_w4569_,
		_w4570_,
		_w4571_
	);
	LUT4 #(
		.INIT('heaee)
	) name2822 (
		_w4554_,
		_w4557_,
		_w4568_,
		_w4571_,
		_w4572_
	);
	LUT2 #(
		.INIT('h8)
	) name2823 (
		\u4_u0_csr1_reg[0]/P0001 ,
		\u4_u0_dma_in_cnt_reg[8]/P0001 ,
		_w4573_
	);
	LUT2 #(
		.INIT('h8)
	) name2824 (
		\u4_u0_csr1_reg[0]/P0001 ,
		\u4_u0_dma_in_cnt_reg[7]/P0001 ,
		_w4574_
	);
	LUT4 #(
		.INIT('h070f)
	) name2825 (
		_w4430_,
		_w4431_,
		_w4573_,
		_w4574_,
		_w4575_
	);
	LUT2 #(
		.INIT('h2)
	) name2826 (
		_w4433_,
		_w4575_,
		_w4576_
	);
	LUT4 #(
		.INIT('h0001)
	) name2827 (
		\u1_u3_buf0_rl_reg/P0001 ,
		\u1_u3_buf0_set_reg/P0001 ,
		\u4_u0_dma_in_cnt_reg[8]/P0001 ,
		\u4_u0_set_r_reg/P0001 ,
		_w4577_
	);
	LUT2 #(
		.INIT('h2)
	) name2828 (
		\u4_u0_csr1_reg[0]/P0001 ,
		\u4_u0_r5_reg/NET0131 ,
		_w4578_
	);
	LUT4 #(
		.INIT('h00a8)
	) name2829 (
		\u4_u0_csr1_reg[0]/P0001 ,
		\u4_u0_dma_in_cnt_reg[8]/P0001 ,
		\u4_u0_ep_match_r_reg/P0001 ,
		\u4_u0_r5_reg/NET0131 ,
		_w4579_
	);
	LUT2 #(
		.INIT('h4)
	) name2830 (
		_w4577_,
		_w4579_,
		_w4580_
	);
	LUT2 #(
		.INIT('h9)
	) name2831 (
		\u4_u0_csr0_reg[10]/P0001 ,
		\u4_u0_dma_in_cnt_reg[8]/P0001 ,
		_w4581_
	);
	LUT4 #(
		.INIT('h7310)
	) name2832 (
		\u4_u0_csr0_reg[4]/P0001 ,
		\u4_u0_csr0_reg[5]/P0001 ,
		\u4_u0_dma_in_cnt_reg[2]/P0001 ,
		\u4_u0_dma_in_cnt_reg[3]/P0001 ,
		_w4582_
	);
	LUT4 #(
		.INIT('h08ce)
	) name2833 (
		\u4_u0_csr0_reg[2]/P0001 ,
		\u4_u0_csr0_reg[3]/NET0131 ,
		\u4_u0_dma_in_cnt_reg[0]/P0001 ,
		\u4_u0_dma_in_cnt_reg[1]/P0001 ,
		_w4583_
	);
	LUT4 #(
		.INIT('h5f57)
	) name2834 (
		_w4419_,
		_w4421_,
		_w4582_,
		_w4583_,
		_w4584_
	);
	LUT4 #(
		.INIT('h8caf)
	) name2835 (
		\u4_u0_csr0_reg[8]/P0001 ,
		\u4_u0_csr0_reg[9]/P0001 ,
		\u4_u0_dma_in_cnt_reg[6]/P0001 ,
		\u4_u0_dma_in_cnt_reg[7]/P0001 ,
		_w4585_
	);
	LUT4 #(
		.INIT('h8caf)
	) name2836 (
		\u4_u0_csr0_reg[6]/P0001 ,
		\u4_u0_csr0_reg[7]/P0001 ,
		\u4_u0_dma_in_cnt_reg[4]/P0001 ,
		\u4_u0_dma_in_cnt_reg[5]/P0001 ,
		_w4586_
	);
	LUT4 #(
		.INIT('h7310)
	) name2837 (
		\u4_u0_csr0_reg[6]/P0001 ,
		\u4_u0_csr0_reg[7]/P0001 ,
		\u4_u0_dma_in_cnt_reg[4]/P0001 ,
		\u4_u0_dma_in_cnt_reg[5]/P0001 ,
		_w4587_
	);
	LUT2 #(
		.INIT('h2)
	) name2838 (
		_w4585_,
		_w4587_,
		_w4588_
	);
	LUT4 #(
		.INIT('h080a)
	) name2839 (
		\u4_u0_csr0_reg[8]/P0001 ,
		\u4_u0_csr0_reg[9]/P0001 ,
		\u4_u0_dma_in_cnt_reg[6]/P0001 ,
		\u4_u0_dma_in_cnt_reg[7]/P0001 ,
		_w4589_
	);
	LUT4 #(
		.INIT('hf731)
	) name2840 (
		\u4_u0_csr0_reg[8]/P0001 ,
		\u4_u0_csr0_reg[9]/P0001 ,
		\u4_u0_dma_in_cnt_reg[6]/P0001 ,
		\u4_u0_dma_in_cnt_reg[7]/P0001 ,
		_w4590_
	);
	LUT4 #(
		.INIT('h80aa)
	) name2841 (
		_w4581_,
		_w4584_,
		_w4588_,
		_w4590_,
		_w4591_
	);
	LUT4 #(
		.INIT('hf0e0)
	) name2842 (
		\u1_u3_buf0_rl_reg/P0001 ,
		\u1_u3_buf0_set_reg/P0001 ,
		\u4_u0_ep_match_r_reg/P0001 ,
		\u4_u0_set_r_reg/P0001 ,
		_w4592_
	);
	LUT2 #(
		.INIT('h4)
	) name2843 (
		_w4581_,
		_w4590_,
		_w4593_
	);
	LUT4 #(
		.INIT('h80f0)
	) name2844 (
		_w4584_,
		_w4588_,
		_w4592_,
		_w4593_,
		_w4594_
	);
	LUT4 #(
		.INIT('heaee)
	) name2845 (
		_w4576_,
		_w4580_,
		_w4591_,
		_w4594_,
		_w4595_
	);
	LUT4 #(
		.INIT('h0001)
	) name2846 (
		\u1_u3_buf0_rl_reg/P0001 ,
		\u1_u3_buf0_set_reg/P0001 ,
		\u4_u1_dma_in_cnt_reg[8]/P0001 ,
		\u4_u1_set_r_reg/P0001 ,
		_w4596_
	);
	LUT4 #(
		.INIT('h00a8)
	) name2847 (
		\u4_u1_csr1_reg[0]/P0001 ,
		\u4_u1_dma_in_cnt_reg[8]/P0001 ,
		\u4_u1_ep_match_r_reg/P0001 ,
		\u4_u1_r5_reg/NET0131 ,
		_w4597_
	);
	LUT2 #(
		.INIT('h4)
	) name2848 (
		_w4596_,
		_w4597_,
		_w4598_
	);
	LUT4 #(
		.INIT('h1333)
	) name2849 (
		\u4_u1_dma_in_cnt_reg[7]/P0001 ,
		\u4_u1_dma_in_cnt_reg[8]/P0001 ,
		_w4447_,
		_w4448_,
		_w4599_
	);
	LUT2 #(
		.INIT('h8)
	) name2850 (
		\u4_u1_csr1_reg[0]/P0001 ,
		\u4_u1_r5_reg/NET0131 ,
		_w4600_
	);
	LUT4 #(
		.INIT('h7f00)
	) name2851 (
		_w4447_,
		_w4448_,
		_w4449_,
		_w4600_,
		_w4601_
	);
	LUT3 #(
		.INIT('h45)
	) name2852 (
		_w4598_,
		_w4599_,
		_w4601_,
		_w4602_
	);
	LUT2 #(
		.INIT('h9)
	) name2853 (
		\u4_u1_csr0_reg[10]/P0001 ,
		\u4_u1_dma_in_cnt_reg[8]/P0001 ,
		_w4603_
	);
	LUT4 #(
		.INIT('hf531)
	) name2854 (
		\u4_u1_csr0_reg[7]/P0001 ,
		\u4_u1_csr0_reg[8]/P0001 ,
		\u4_u1_dma_in_cnt_reg[5]/P0001 ,
		\u4_u1_dma_in_cnt_reg[6]/P0001 ,
		_w4604_
	);
	LUT4 #(
		.INIT('hef00)
	) name2855 (
		_w4463_,
		_w4468_,
		_w4469_,
		_w4604_,
		_w4605_
	);
	LUT4 #(
		.INIT('h8caf)
	) name2856 (
		\u4_u1_csr0_reg[8]/P0001 ,
		\u4_u1_csr0_reg[9]/P0001 ,
		\u4_u1_dma_in_cnt_reg[6]/P0001 ,
		\u4_u1_dma_in_cnt_reg[7]/P0001 ,
		_w4606_
	);
	LUT4 #(
		.INIT('h6366)
	) name2857 (
		_w4472_,
		_w4603_,
		_w4605_,
		_w4606_,
		_w4607_
	);
	LUT3 #(
		.INIT('h8a)
	) name2858 (
		_w4454_,
		_w4599_,
		_w4601_,
		_w4608_
	);
	LUT3 #(
		.INIT('h15)
	) name2859 (
		_w4602_,
		_w4607_,
		_w4608_,
		_w4609_
	);
	LUT4 #(
		.INIT('hf0e0)
	) name2860 (
		\u1_u3_buf0_rl_reg/P0001 ,
		\u1_u3_buf0_set_reg/P0001 ,
		\u4_u2_ep_match_r_reg/P0001 ,
		\u4_u2_set_r_reg/P0001 ,
		_w4610_
	);
	LUT2 #(
		.INIT('h9)
	) name2861 (
		\u4_u2_csr0_reg[10]/P0001 ,
		\u4_u2_dma_in_cnt_reg[8]/P0001 ,
		_w4611_
	);
	LUT4 #(
		.INIT('hddfd)
	) name2862 (
		\u4_u2_ep_match_r_reg/P0001 ,
		_w4482_,
		_w4485_,
		_w4611_,
		_w4612_
	);
	LUT3 #(
		.INIT('h2a)
	) name2863 (
		_w4500_,
		_w4610_,
		_w4611_,
		_w4613_
	);
	LUT3 #(
		.INIT('h13)
	) name2864 (
		_w4499_,
		_w4612_,
		_w4613_,
		_w4614_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name2865 (
		\u4_u2_r5_reg/NET0131 ,
		_w4504_,
		_w4505_,
		_w4506_,
		_w4615_
	);
	LUT4 #(
		.INIT('h1333)
	) name2866 (
		\u4_u2_dma_in_cnt_reg[7]/P0001 ,
		\u4_u2_dma_in_cnt_reg[8]/P0001 ,
		_w4504_,
		_w4505_,
		_w4616_
	);
	LUT4 #(
		.INIT('h8a45)
	) name2867 (
		\u4_u2_csr0_reg[10]/P0001 ,
		\u4_u2_csr0_reg[9]/P0001 ,
		\u4_u2_dma_in_cnt_reg[7]/P0001 ,
		\u4_u2_dma_in_cnt_reg[8]/P0001 ,
		_w4617_
	);
	LUT3 #(
		.INIT('h0d)
	) name2868 (
		_w4615_,
		_w4616_,
		_w4617_,
		_w4618_
	);
	LUT3 #(
		.INIT('ha2)
	) name2869 (
		_w4500_,
		_w4615_,
		_w4616_,
		_w4619_
	);
	LUT3 #(
		.INIT('h13)
	) name2870 (
		_w4499_,
		_w4618_,
		_w4619_,
		_w4620_
	);
	LUT4 #(
		.INIT('h0001)
	) name2871 (
		\u1_u3_buf0_rl_reg/P0001 ,
		\u1_u3_buf0_set_reg/P0001 ,
		\u4_u2_dma_in_cnt_reg[8]/P0001 ,
		\u4_u2_set_r_reg/P0001 ,
		_w4621_
	);
	LUT3 #(
		.INIT('h0e)
	) name2872 (
		\u4_u2_dma_in_cnt_reg[8]/P0001 ,
		\u4_u2_ep_match_r_reg/P0001 ,
		\u4_u2_r5_reg/NET0131 ,
		_w4622_
	);
	LUT2 #(
		.INIT('h4)
	) name2873 (
		_w4621_,
		_w4622_,
		_w4623_
	);
	LUT4 #(
		.INIT('haa08)
	) name2874 (
		\u4_u2_csr1_reg[0]/P0001 ,
		_w4615_,
		_w4616_,
		_w4623_,
		_w4624_
	);
	LUT3 #(
		.INIT('hd0)
	) name2875 (
		_w4614_,
		_w4620_,
		_w4624_,
		_w4625_
	);
	LUT4 #(
		.INIT('hf100)
	) name2876 (
		_w4199_,
		_w4351_,
		_w4352_,
		_w4358_,
		_w4626_
	);
	LUT4 #(
		.INIT('h0001)
	) name2877 (
		\u0_u0_me_ps2_reg[0]/P0001 ,
		\u0_u0_me_ps2_reg[1]/P0001 ,
		\u0_u0_me_ps2_reg[2]/P0001 ,
		\u0_u0_me_ps2_reg[4]/P0001 ,
		_w4627_
	);
	LUT3 #(
		.INIT('he0)
	) name2878 (
		\u0_u0_me_ps2_reg[3]/P0001 ,
		\u0_u0_me_ps2_reg[4]/P0001 ,
		\u0_u0_me_ps2_reg[5]/P0001 ,
		_w4628_
	);
	LUT2 #(
		.INIT('h1)
	) name2879 (
		\u0_u0_me_ps2_reg[6]/P0001 ,
		\u0_u0_me_ps2_reg[7]/P0001 ,
		_w4629_
	);
	LUT3 #(
		.INIT('hb0)
	) name2880 (
		_w4627_,
		_w4628_,
		_w4629_,
		_w4630_
	);
	LUT2 #(
		.INIT('h2)
	) name2881 (
		_w4626_,
		_w4630_,
		_w4631_
	);
	LUT2 #(
		.INIT('h4)
	) name2882 (
		_w4350_,
		_w4631_,
		_w4632_
	);
	LUT2 #(
		.INIT('h1)
	) name2883 (
		\u0_u0_me_ps_2_5_us_reg/P0001 ,
		\u0_u0_me_ps_reg[0]/P0001 ,
		_w4633_
	);
	LUT2 #(
		.INIT('h8)
	) name2884 (
		_w4626_,
		_w4633_,
		_w4634_
	);
	LUT2 #(
		.INIT('h4)
	) name2885 (
		_w4350_,
		_w4634_,
		_w4635_
	);
	LUT4 #(
		.INIT('h8000)
	) name2886 (
		\u0_u0_me_ps_reg[0]/P0001 ,
		\u0_u0_me_ps_reg[1]/P0001 ,
		\u0_u0_me_ps_reg[2]/P0001 ,
		\u0_u0_me_ps_reg[3]/P0001 ,
		_w4636_
	);
	LUT2 #(
		.INIT('h8)
	) name2887 (
		\u0_u0_me_ps_reg[4]/P0001 ,
		\u0_u0_me_ps_reg[5]/P0001 ,
		_w4637_
	);
	LUT4 #(
		.INIT('h1450)
	) name2888 (
		\u0_u0_me_ps_2_5_us_reg/P0001 ,
		\u0_u0_me_ps_reg[4]/P0001 ,
		\u0_u0_me_ps_reg[5]/P0001 ,
		_w4636_,
		_w4638_
	);
	LUT2 #(
		.INIT('h8)
	) name2889 (
		_w4626_,
		_w4638_,
		_w4639_
	);
	LUT2 #(
		.INIT('h4)
	) name2890 (
		_w4350_,
		_w4639_,
		_w4640_
	);
	LUT3 #(
		.INIT('h15)
	) name2891 (
		\u0_u0_me_ps_reg[6]/P0001 ,
		_w4636_,
		_w4637_,
		_w4641_
	);
	LUT3 #(
		.INIT('h80)
	) name2892 (
		\u0_u0_me_ps_reg[4]/P0001 ,
		\u0_u0_me_ps_reg[5]/P0001 ,
		\u0_u0_me_ps_reg[6]/P0001 ,
		_w4642_
	);
	LUT3 #(
		.INIT('h15)
	) name2893 (
		\u0_u0_me_ps_2_5_us_reg/P0001 ,
		_w4636_,
		_w4642_,
		_w4643_
	);
	LUT2 #(
		.INIT('h4)
	) name2894 (
		_w4641_,
		_w4643_,
		_w4644_
	);
	LUT2 #(
		.INIT('h8)
	) name2895 (
		_w4626_,
		_w4644_,
		_w4645_
	);
	LUT2 #(
		.INIT('h4)
	) name2896 (
		_w4350_,
		_w4645_,
		_w4646_
	);
	LUT4 #(
		.INIT('hebbb)
	) name2897 (
		\u0_u0_me_ps_2_5_us_reg/P0001 ,
		\u0_u0_me_ps_reg[7]/P0001 ,
		_w4636_,
		_w4642_,
		_w4647_
	);
	LUT2 #(
		.INIT('h2)
	) name2898 (
		_w4626_,
		_w4647_,
		_w4648_
	);
	LUT2 #(
		.INIT('h4)
	) name2899 (
		_w4350_,
		_w4648_,
		_w4649_
	);
	LUT3 #(
		.INIT('h01)
	) name2900 (
		\u4_u3_dma_out_cnt_reg[4]/P0001 ,
		\u4_u3_dma_out_cnt_reg[5]/P0001 ,
		\u4_u3_dma_out_cnt_reg[6]/P0001 ,
		_w4650_
	);
	LUT2 #(
		.INIT('h1)
	) name2901 (
		\u4_u3_dma_in_cnt_reg[0]/P0001 ,
		\u4_u3_dma_out_cnt_reg[1]/P0001 ,
		_w4651_
	);
	LUT4 #(
		.INIT('h0001)
	) name2902 (
		\u4_u3_dma_in_cnt_reg[0]/P0001 ,
		\u4_u3_dma_out_cnt_reg[1]/P0001 ,
		\u4_u3_dma_out_cnt_reg[2]/P0001 ,
		\u4_u3_dma_out_cnt_reg[3]/P0001 ,
		_w4652_
	);
	LUT3 #(
		.INIT('h10)
	) name2903 (
		\u4_u3_dma_out_cnt_reg[7]/P0001 ,
		\u4_u3_dma_out_cnt_reg[8]/P0001 ,
		\u4_u3_r5_reg/NET0131 ,
		_w4653_
	);
	LUT4 #(
		.INIT('h8000)
	) name2904 (
		\u4_u3_csr1_reg[0]/P0001 ,
		_w4650_,
		_w4652_,
		_w4653_,
		_w4654_
	);
	LUT3 #(
		.INIT('h80)
	) name2905 (
		\u4_u3_csr1_reg[0]/P0001 ,
		\u4_u3_dma_out_cnt_reg[8]/P0001 ,
		\u4_u3_r5_reg/NET0131 ,
		_w4655_
	);
	LUT4 #(
		.INIT('hbf00)
	) name2906 (
		\u4_u3_dma_out_cnt_reg[7]/P0001 ,
		_w4650_,
		_w4652_,
		_w4655_,
		_w4656_
	);
	LUT4 #(
		.INIT('h0001)
	) name2907 (
		\u1_u3_buf0_rl_reg/P0001 ,
		\u1_u3_buf0_set_reg/P0001 ,
		\u4_u3_dma_out_cnt_reg[8]/P0001 ,
		\u4_u3_set_r_reg/P0001 ,
		_w4657_
	);
	LUT4 #(
		.INIT('h00a8)
	) name2908 (
		\u4_u3_csr1_reg[0]/P0001 ,
		\u4_u3_dma_out_cnt_reg[8]/P0001 ,
		\u4_u3_ep_match_r_reg/P0001 ,
		\u4_u3_r5_reg/NET0131 ,
		_w4658_
	);
	LUT2 #(
		.INIT('h4)
	) name2909 (
		_w4657_,
		_w4658_,
		_w4659_
	);
	LUT3 #(
		.INIT('h01)
	) name2910 (
		_w4654_,
		_w4656_,
		_w4659_,
		_w4660_
	);
	LUT2 #(
		.INIT('h8)
	) name2911 (
		\u4_u3_csr0_reg[10]/P0001 ,
		\u4_u3_dma_out_cnt_reg[8]/P0001 ,
		_w4661_
	);
	LUT2 #(
		.INIT('h6)
	) name2912 (
		\u4_u3_csr0_reg[10]/P0001 ,
		\u4_u3_dma_out_cnt_reg[8]/P0001 ,
		_w4662_
	);
	LUT2 #(
		.INIT('h1)
	) name2913 (
		\u4_u3_csr0_reg[9]/P0001 ,
		\u4_u3_dma_out_cnt_reg[7]/P0001 ,
		_w4663_
	);
	LUT2 #(
		.INIT('h1)
	) name2914 (
		\u4_u3_csr0_reg[8]/P0001 ,
		\u4_u3_dma_out_cnt_reg[6]/P0001 ,
		_w4664_
	);
	LUT4 #(
		.INIT('ha080)
	) name2915 (
		\u4_u3_csr0_reg[7]/P0001 ,
		\u4_u3_csr0_reg[8]/P0001 ,
		\u4_u3_dma_out_cnt_reg[5]/P0001 ,
		\u4_u3_dma_out_cnt_reg[6]/P0001 ,
		_w4665_
	);
	LUT4 #(
		.INIT('h135f)
	) name2916 (
		\u4_u3_csr0_reg[5]/P0001 ,
		\u4_u3_csr0_reg[6]/P0001 ,
		\u4_u3_dma_out_cnt_reg[3]/P0001 ,
		\u4_u3_dma_out_cnt_reg[4]/P0001 ,
		_w4666_
	);
	LUT4 #(
		.INIT('h0105)
	) name2917 (
		\u4_u3_csr0_reg[5]/P0001 ,
		\u4_u3_csr0_reg[6]/P0001 ,
		\u4_u3_dma_out_cnt_reg[3]/P0001 ,
		\u4_u3_dma_out_cnt_reg[4]/P0001 ,
		_w4667_
	);
	LUT2 #(
		.INIT('h8)
	) name2918 (
		\u4_u3_csr0_reg[2]/P0001 ,
		\u4_u3_dma_in_cnt_reg[0]/P0001 ,
		_w4668_
	);
	LUT4 #(
		.INIT('h135f)
	) name2919 (
		\u4_u3_csr0_reg[2]/P0001 ,
		\u4_u3_csr0_reg[3]/NET0131 ,
		\u4_u3_dma_in_cnt_reg[0]/P0001 ,
		\u4_u3_dma_out_cnt_reg[1]/P0001 ,
		_w4669_
	);
	LUT4 #(
		.INIT('hfac8)
	) name2920 (
		\u4_u3_csr0_reg[3]/NET0131 ,
		\u4_u3_csr0_reg[4]/P0001 ,
		\u4_u3_dma_out_cnt_reg[1]/P0001 ,
		\u4_u3_dma_out_cnt_reg[2]/P0001 ,
		_w4670_
	);
	LUT2 #(
		.INIT('h8)
	) name2921 (
		\u4_u3_csr0_reg[4]/P0001 ,
		\u4_u3_dma_out_cnt_reg[2]/P0001 ,
		_w4671_
	);
	LUT4 #(
		.INIT('h008a)
	) name2922 (
		_w4666_,
		_w4669_,
		_w4670_,
		_w4671_,
		_w4672_
	);
	LUT2 #(
		.INIT('h1)
	) name2923 (
		\u4_u3_csr0_reg[6]/P0001 ,
		\u4_u3_dma_out_cnt_reg[4]/P0001 ,
		_w4673_
	);
	LUT4 #(
		.INIT('hfac8)
	) name2924 (
		\u4_u3_csr0_reg[6]/P0001 ,
		\u4_u3_csr0_reg[7]/P0001 ,
		\u4_u3_dma_out_cnt_reg[4]/P0001 ,
		\u4_u3_dma_out_cnt_reg[5]/P0001 ,
		_w4674_
	);
	LUT2 #(
		.INIT('h4)
	) name2925 (
		_w4664_,
		_w4674_,
		_w4675_
	);
	LUT4 #(
		.INIT('h5455)
	) name2926 (
		_w4665_,
		_w4667_,
		_w4672_,
		_w4675_,
		_w4676_
	);
	LUT4 #(
		.INIT('h135f)
	) name2927 (
		\u4_u3_csr0_reg[8]/P0001 ,
		\u4_u3_csr0_reg[9]/P0001 ,
		\u4_u3_dma_out_cnt_reg[6]/P0001 ,
		\u4_u3_dma_out_cnt_reg[7]/P0001 ,
		_w4677_
	);
	LUT4 #(
		.INIT('h5666)
	) name2928 (
		_w4662_,
		_w4663_,
		_w4676_,
		_w4677_,
		_w4678_
	);
	LUT3 #(
		.INIT('h02)
	) name2929 (
		_w4569_,
		_w4654_,
		_w4656_,
		_w4679_
	);
	LUT3 #(
		.INIT('h15)
	) name2930 (
		_w4660_,
		_w4678_,
		_w4679_,
		_w4680_
	);
	LUT3 #(
		.INIT('h01)
	) name2931 (
		\u4_u0_dma_out_cnt_reg[4]/P0001 ,
		\u4_u0_dma_out_cnt_reg[5]/P0001 ,
		\u4_u0_dma_out_cnt_reg[6]/P0001 ,
		_w4681_
	);
	LUT2 #(
		.INIT('h1)
	) name2932 (
		\u4_u0_dma_in_cnt_reg[0]/P0001 ,
		\u4_u0_dma_out_cnt_reg[1]/P0001 ,
		_w4682_
	);
	LUT4 #(
		.INIT('h0001)
	) name2933 (
		\u4_u0_dma_in_cnt_reg[0]/P0001 ,
		\u4_u0_dma_out_cnt_reg[1]/P0001 ,
		\u4_u0_dma_out_cnt_reg[2]/P0001 ,
		\u4_u0_dma_out_cnt_reg[3]/P0001 ,
		_w4683_
	);
	LUT3 #(
		.INIT('h10)
	) name2934 (
		\u4_u0_dma_out_cnt_reg[7]/P0001 ,
		\u4_u0_dma_out_cnt_reg[8]/P0001 ,
		\u4_u0_r5_reg/NET0131 ,
		_w4684_
	);
	LUT4 #(
		.INIT('h8000)
	) name2935 (
		\u4_u0_csr1_reg[0]/P0001 ,
		_w4681_,
		_w4683_,
		_w4684_,
		_w4685_
	);
	LUT3 #(
		.INIT('h80)
	) name2936 (
		\u4_u0_csr1_reg[0]/P0001 ,
		\u4_u0_dma_out_cnt_reg[8]/P0001 ,
		\u4_u0_r5_reg/NET0131 ,
		_w4686_
	);
	LUT4 #(
		.INIT('hbf00)
	) name2937 (
		\u4_u0_dma_out_cnt_reg[7]/P0001 ,
		_w4681_,
		_w4683_,
		_w4686_,
		_w4687_
	);
	LUT4 #(
		.INIT('h0001)
	) name2938 (
		\u1_u3_buf0_rl_reg/P0001 ,
		\u1_u3_buf0_set_reg/P0001 ,
		\u4_u0_dma_out_cnt_reg[8]/P0001 ,
		\u4_u0_set_r_reg/P0001 ,
		_w4688_
	);
	LUT4 #(
		.INIT('h00a8)
	) name2939 (
		\u4_u0_csr1_reg[0]/P0001 ,
		\u4_u0_dma_out_cnt_reg[8]/P0001 ,
		\u4_u0_ep_match_r_reg/P0001 ,
		\u4_u0_r5_reg/NET0131 ,
		_w4689_
	);
	LUT2 #(
		.INIT('h4)
	) name2940 (
		_w4688_,
		_w4689_,
		_w4690_
	);
	LUT3 #(
		.INIT('h01)
	) name2941 (
		_w4685_,
		_w4687_,
		_w4690_,
		_w4691_
	);
	LUT2 #(
		.INIT('h6)
	) name2942 (
		\u4_u0_csr0_reg[10]/P0001 ,
		\u4_u0_dma_out_cnt_reg[8]/P0001 ,
		_w4692_
	);
	LUT2 #(
		.INIT('h1)
	) name2943 (
		\u4_u0_csr0_reg[9]/P0001 ,
		\u4_u0_dma_out_cnt_reg[7]/P0001 ,
		_w4693_
	);
	LUT2 #(
		.INIT('h1)
	) name2944 (
		\u4_u0_csr0_reg[8]/P0001 ,
		\u4_u0_dma_out_cnt_reg[6]/P0001 ,
		_w4694_
	);
	LUT4 #(
		.INIT('ha080)
	) name2945 (
		\u4_u0_csr0_reg[7]/P0001 ,
		\u4_u0_csr0_reg[8]/P0001 ,
		\u4_u0_dma_out_cnt_reg[5]/P0001 ,
		\u4_u0_dma_out_cnt_reg[6]/P0001 ,
		_w4695_
	);
	LUT4 #(
		.INIT('h135f)
	) name2946 (
		\u4_u0_csr0_reg[5]/P0001 ,
		\u4_u0_csr0_reg[6]/P0001 ,
		\u4_u0_dma_out_cnt_reg[3]/P0001 ,
		\u4_u0_dma_out_cnt_reg[4]/P0001 ,
		_w4696_
	);
	LUT4 #(
		.INIT('h0105)
	) name2947 (
		\u4_u0_csr0_reg[5]/P0001 ,
		\u4_u0_csr0_reg[6]/P0001 ,
		\u4_u0_dma_out_cnt_reg[3]/P0001 ,
		\u4_u0_dma_out_cnt_reg[4]/P0001 ,
		_w4697_
	);
	LUT2 #(
		.INIT('h8)
	) name2948 (
		\u4_u0_csr0_reg[2]/P0001 ,
		\u4_u0_dma_in_cnt_reg[0]/P0001 ,
		_w4698_
	);
	LUT4 #(
		.INIT('h135f)
	) name2949 (
		\u4_u0_csr0_reg[2]/P0001 ,
		\u4_u0_csr0_reg[3]/NET0131 ,
		\u4_u0_dma_in_cnt_reg[0]/P0001 ,
		\u4_u0_dma_out_cnt_reg[1]/P0001 ,
		_w4699_
	);
	LUT4 #(
		.INIT('hfac8)
	) name2950 (
		\u4_u0_csr0_reg[3]/NET0131 ,
		\u4_u0_csr0_reg[4]/P0001 ,
		\u4_u0_dma_out_cnt_reg[1]/P0001 ,
		\u4_u0_dma_out_cnt_reg[2]/P0001 ,
		_w4700_
	);
	LUT2 #(
		.INIT('h8)
	) name2951 (
		\u4_u0_csr0_reg[4]/P0001 ,
		\u4_u0_dma_out_cnt_reg[2]/P0001 ,
		_w4701_
	);
	LUT4 #(
		.INIT('h008a)
	) name2952 (
		_w4696_,
		_w4699_,
		_w4700_,
		_w4701_,
		_w4702_
	);
	LUT2 #(
		.INIT('h1)
	) name2953 (
		\u4_u0_csr0_reg[6]/P0001 ,
		\u4_u0_dma_out_cnt_reg[4]/P0001 ,
		_w4703_
	);
	LUT4 #(
		.INIT('hfac8)
	) name2954 (
		\u4_u0_csr0_reg[6]/P0001 ,
		\u4_u0_csr0_reg[7]/P0001 ,
		\u4_u0_dma_out_cnt_reg[4]/P0001 ,
		\u4_u0_dma_out_cnt_reg[5]/P0001 ,
		_w4704_
	);
	LUT2 #(
		.INIT('h4)
	) name2955 (
		_w4694_,
		_w4704_,
		_w4705_
	);
	LUT4 #(
		.INIT('h5455)
	) name2956 (
		_w4695_,
		_w4697_,
		_w4702_,
		_w4705_,
		_w4706_
	);
	LUT4 #(
		.INIT('h135f)
	) name2957 (
		\u4_u0_csr0_reg[8]/P0001 ,
		\u4_u0_csr0_reg[9]/P0001 ,
		\u4_u0_dma_out_cnt_reg[6]/P0001 ,
		\u4_u0_dma_out_cnt_reg[7]/P0001 ,
		_w4707_
	);
	LUT4 #(
		.INIT('h5666)
	) name2958 (
		_w4692_,
		_w4693_,
		_w4706_,
		_w4707_,
		_w4708_
	);
	LUT3 #(
		.INIT('h02)
	) name2959 (
		_w4592_,
		_w4685_,
		_w4687_,
		_w4709_
	);
	LUT3 #(
		.INIT('h15)
	) name2960 (
		_w4691_,
		_w4708_,
		_w4709_,
		_w4710_
	);
	LUT3 #(
		.INIT('h01)
	) name2961 (
		\u4_u1_dma_out_cnt_reg[4]/P0001 ,
		\u4_u1_dma_out_cnt_reg[5]/P0001 ,
		\u4_u1_dma_out_cnt_reg[6]/P0001 ,
		_w4711_
	);
	LUT2 #(
		.INIT('h1)
	) name2962 (
		\u4_u1_dma_in_cnt_reg[0]/P0001 ,
		\u4_u1_dma_out_cnt_reg[1]/P0001 ,
		_w4712_
	);
	LUT4 #(
		.INIT('h0001)
	) name2963 (
		\u4_u1_dma_in_cnt_reg[0]/P0001 ,
		\u4_u1_dma_out_cnt_reg[1]/P0001 ,
		\u4_u1_dma_out_cnt_reg[2]/P0001 ,
		\u4_u1_dma_out_cnt_reg[3]/P0001 ,
		_w4713_
	);
	LUT3 #(
		.INIT('h10)
	) name2964 (
		\u4_u1_dma_out_cnt_reg[7]/P0001 ,
		\u4_u1_dma_out_cnt_reg[8]/P0001 ,
		\u4_u1_r5_reg/NET0131 ,
		_w4714_
	);
	LUT4 #(
		.INIT('h8000)
	) name2965 (
		\u4_u1_csr1_reg[0]/P0001 ,
		_w4711_,
		_w4713_,
		_w4714_,
		_w4715_
	);
	LUT3 #(
		.INIT('h80)
	) name2966 (
		\u4_u1_csr1_reg[0]/P0001 ,
		\u4_u1_dma_out_cnt_reg[8]/P0001 ,
		\u4_u1_r5_reg/NET0131 ,
		_w4716_
	);
	LUT4 #(
		.INIT('hbf00)
	) name2967 (
		\u4_u1_dma_out_cnt_reg[7]/P0001 ,
		_w4711_,
		_w4713_,
		_w4716_,
		_w4717_
	);
	LUT4 #(
		.INIT('h0001)
	) name2968 (
		\u1_u3_buf0_rl_reg/P0001 ,
		\u1_u3_buf0_set_reg/P0001 ,
		\u4_u1_dma_out_cnt_reg[8]/P0001 ,
		\u4_u1_set_r_reg/P0001 ,
		_w4718_
	);
	LUT4 #(
		.INIT('h00a8)
	) name2969 (
		\u4_u1_csr1_reg[0]/P0001 ,
		\u4_u1_dma_out_cnt_reg[8]/P0001 ,
		\u4_u1_ep_match_r_reg/P0001 ,
		\u4_u1_r5_reg/NET0131 ,
		_w4719_
	);
	LUT2 #(
		.INIT('h4)
	) name2970 (
		_w4718_,
		_w4719_,
		_w4720_
	);
	LUT3 #(
		.INIT('h01)
	) name2971 (
		_w4715_,
		_w4717_,
		_w4720_,
		_w4721_
	);
	LUT2 #(
		.INIT('h8)
	) name2972 (
		\u4_u1_csr0_reg[10]/P0001 ,
		\u4_u1_dma_out_cnt_reg[8]/P0001 ,
		_w4722_
	);
	LUT2 #(
		.INIT('h6)
	) name2973 (
		\u4_u1_csr0_reg[10]/P0001 ,
		\u4_u1_dma_out_cnt_reg[8]/P0001 ,
		_w4723_
	);
	LUT2 #(
		.INIT('h1)
	) name2974 (
		\u4_u1_csr0_reg[9]/P0001 ,
		\u4_u1_dma_out_cnt_reg[7]/P0001 ,
		_w4724_
	);
	LUT2 #(
		.INIT('h1)
	) name2975 (
		\u4_u1_csr0_reg[8]/P0001 ,
		\u4_u1_dma_out_cnt_reg[6]/P0001 ,
		_w4725_
	);
	LUT4 #(
		.INIT('ha080)
	) name2976 (
		\u4_u1_csr0_reg[7]/P0001 ,
		\u4_u1_csr0_reg[8]/P0001 ,
		\u4_u1_dma_out_cnt_reg[5]/P0001 ,
		\u4_u1_dma_out_cnt_reg[6]/P0001 ,
		_w4726_
	);
	LUT4 #(
		.INIT('h135f)
	) name2977 (
		\u4_u1_csr0_reg[5]/P0001 ,
		\u4_u1_csr0_reg[6]/P0001 ,
		\u4_u1_dma_out_cnt_reg[3]/P0001 ,
		\u4_u1_dma_out_cnt_reg[4]/P0001 ,
		_w4727_
	);
	LUT4 #(
		.INIT('h0105)
	) name2978 (
		\u4_u1_csr0_reg[5]/P0001 ,
		\u4_u1_csr0_reg[6]/P0001 ,
		\u4_u1_dma_out_cnt_reg[3]/P0001 ,
		\u4_u1_dma_out_cnt_reg[4]/P0001 ,
		_w4728_
	);
	LUT2 #(
		.INIT('h8)
	) name2979 (
		\u4_u1_csr0_reg[2]/P0001 ,
		\u4_u1_dma_in_cnt_reg[0]/P0001 ,
		_w4729_
	);
	LUT4 #(
		.INIT('h135f)
	) name2980 (
		\u4_u1_csr0_reg[2]/P0001 ,
		\u4_u1_csr0_reg[3]/NET0131 ,
		\u4_u1_dma_in_cnt_reg[0]/P0001 ,
		\u4_u1_dma_out_cnt_reg[1]/P0001 ,
		_w4730_
	);
	LUT4 #(
		.INIT('hfac8)
	) name2981 (
		\u4_u1_csr0_reg[3]/NET0131 ,
		\u4_u1_csr0_reg[4]/P0001 ,
		\u4_u1_dma_out_cnt_reg[1]/P0001 ,
		\u4_u1_dma_out_cnt_reg[2]/P0001 ,
		_w4731_
	);
	LUT2 #(
		.INIT('h8)
	) name2982 (
		\u4_u1_csr0_reg[4]/P0001 ,
		\u4_u1_dma_out_cnt_reg[2]/P0001 ,
		_w4732_
	);
	LUT4 #(
		.INIT('h008a)
	) name2983 (
		_w4727_,
		_w4730_,
		_w4731_,
		_w4732_,
		_w4733_
	);
	LUT2 #(
		.INIT('h1)
	) name2984 (
		\u4_u1_csr0_reg[6]/P0001 ,
		\u4_u1_dma_out_cnt_reg[4]/P0001 ,
		_w4734_
	);
	LUT4 #(
		.INIT('hfac8)
	) name2985 (
		\u4_u1_csr0_reg[6]/P0001 ,
		\u4_u1_csr0_reg[7]/P0001 ,
		\u4_u1_dma_out_cnt_reg[4]/P0001 ,
		\u4_u1_dma_out_cnt_reg[5]/P0001 ,
		_w4735_
	);
	LUT2 #(
		.INIT('h4)
	) name2986 (
		_w4725_,
		_w4735_,
		_w4736_
	);
	LUT4 #(
		.INIT('h5455)
	) name2987 (
		_w4726_,
		_w4728_,
		_w4733_,
		_w4736_,
		_w4737_
	);
	LUT4 #(
		.INIT('h135f)
	) name2988 (
		\u4_u1_csr0_reg[8]/P0001 ,
		\u4_u1_csr0_reg[9]/P0001 ,
		\u4_u1_dma_out_cnt_reg[6]/P0001 ,
		\u4_u1_dma_out_cnt_reg[7]/P0001 ,
		_w4738_
	);
	LUT4 #(
		.INIT('h5666)
	) name2989 (
		_w4723_,
		_w4724_,
		_w4737_,
		_w4738_,
		_w4739_
	);
	LUT3 #(
		.INIT('h02)
	) name2990 (
		_w4454_,
		_w4715_,
		_w4717_,
		_w4740_
	);
	LUT3 #(
		.INIT('h15)
	) name2991 (
		_w4721_,
		_w4739_,
		_w4740_,
		_w4741_
	);
	LUT3 #(
		.INIT('h01)
	) name2992 (
		\u4_u2_dma_out_cnt_reg[4]/P0001 ,
		\u4_u2_dma_out_cnt_reg[5]/P0001 ,
		\u4_u2_dma_out_cnt_reg[6]/P0001 ,
		_w4742_
	);
	LUT2 #(
		.INIT('h1)
	) name2993 (
		\u4_u2_dma_in_cnt_reg[0]/P0001 ,
		\u4_u2_dma_out_cnt_reg[1]/P0001 ,
		_w4743_
	);
	LUT4 #(
		.INIT('h0001)
	) name2994 (
		\u4_u2_dma_in_cnt_reg[0]/P0001 ,
		\u4_u2_dma_out_cnt_reg[1]/P0001 ,
		\u4_u2_dma_out_cnt_reg[2]/P0001 ,
		\u4_u2_dma_out_cnt_reg[3]/P0001 ,
		_w4744_
	);
	LUT3 #(
		.INIT('h10)
	) name2995 (
		\u4_u2_dma_out_cnt_reg[7]/P0001 ,
		\u4_u2_dma_out_cnt_reg[8]/P0001 ,
		\u4_u2_r5_reg/NET0131 ,
		_w4745_
	);
	LUT4 #(
		.INIT('h8000)
	) name2996 (
		\u4_u2_csr1_reg[0]/P0001 ,
		_w4742_,
		_w4744_,
		_w4745_,
		_w4746_
	);
	LUT3 #(
		.INIT('h80)
	) name2997 (
		\u4_u2_csr1_reg[0]/P0001 ,
		\u4_u2_dma_out_cnt_reg[8]/P0001 ,
		\u4_u2_r5_reg/NET0131 ,
		_w4747_
	);
	LUT4 #(
		.INIT('hbf00)
	) name2998 (
		\u4_u2_dma_out_cnt_reg[7]/P0001 ,
		_w4742_,
		_w4744_,
		_w4747_,
		_w4748_
	);
	LUT4 #(
		.INIT('h0001)
	) name2999 (
		\u1_u3_buf0_rl_reg/P0001 ,
		\u1_u3_buf0_set_reg/P0001 ,
		\u4_u2_dma_out_cnt_reg[8]/P0001 ,
		\u4_u2_set_r_reg/P0001 ,
		_w4749_
	);
	LUT4 #(
		.INIT('h00a8)
	) name3000 (
		\u4_u2_csr1_reg[0]/P0001 ,
		\u4_u2_dma_out_cnt_reg[8]/P0001 ,
		\u4_u2_ep_match_r_reg/P0001 ,
		\u4_u2_r5_reg/NET0131 ,
		_w4750_
	);
	LUT2 #(
		.INIT('h4)
	) name3001 (
		_w4749_,
		_w4750_,
		_w4751_
	);
	LUT3 #(
		.INIT('h01)
	) name3002 (
		_w4746_,
		_w4748_,
		_w4751_,
		_w4752_
	);
	LUT2 #(
		.INIT('h6)
	) name3003 (
		\u4_u2_csr0_reg[10]/P0001 ,
		\u4_u2_dma_out_cnt_reg[8]/P0001 ,
		_w4753_
	);
	LUT2 #(
		.INIT('h1)
	) name3004 (
		\u4_u2_csr0_reg[9]/P0001 ,
		\u4_u2_dma_out_cnt_reg[7]/P0001 ,
		_w4754_
	);
	LUT2 #(
		.INIT('h1)
	) name3005 (
		\u4_u2_csr0_reg[8]/P0001 ,
		\u4_u2_dma_out_cnt_reg[6]/P0001 ,
		_w4755_
	);
	LUT4 #(
		.INIT('ha080)
	) name3006 (
		\u4_u2_csr0_reg[7]/P0001 ,
		\u4_u2_csr0_reg[8]/P0001 ,
		\u4_u2_dma_out_cnt_reg[5]/P0001 ,
		\u4_u2_dma_out_cnt_reg[6]/P0001 ,
		_w4756_
	);
	LUT4 #(
		.INIT('h135f)
	) name3007 (
		\u4_u2_csr0_reg[5]/P0001 ,
		\u4_u2_csr0_reg[6]/P0001 ,
		\u4_u2_dma_out_cnt_reg[3]/P0001 ,
		\u4_u2_dma_out_cnt_reg[4]/P0001 ,
		_w4757_
	);
	LUT4 #(
		.INIT('h0105)
	) name3008 (
		\u4_u2_csr0_reg[5]/P0001 ,
		\u4_u2_csr0_reg[6]/P0001 ,
		\u4_u2_dma_out_cnt_reg[3]/P0001 ,
		\u4_u2_dma_out_cnt_reg[4]/P0001 ,
		_w4758_
	);
	LUT2 #(
		.INIT('h8)
	) name3009 (
		\u4_u2_csr0_reg[2]/P0001 ,
		\u4_u2_dma_in_cnt_reg[0]/P0001 ,
		_w4759_
	);
	LUT4 #(
		.INIT('h135f)
	) name3010 (
		\u4_u2_csr0_reg[2]/P0001 ,
		\u4_u2_csr0_reg[3]/NET0131 ,
		\u4_u2_dma_in_cnt_reg[0]/P0001 ,
		\u4_u2_dma_out_cnt_reg[1]/P0001 ,
		_w4760_
	);
	LUT4 #(
		.INIT('hfac8)
	) name3011 (
		\u4_u2_csr0_reg[3]/NET0131 ,
		\u4_u2_csr0_reg[4]/P0001 ,
		\u4_u2_dma_out_cnt_reg[1]/P0001 ,
		\u4_u2_dma_out_cnt_reg[2]/P0001 ,
		_w4761_
	);
	LUT2 #(
		.INIT('h8)
	) name3012 (
		\u4_u2_csr0_reg[4]/P0001 ,
		\u4_u2_dma_out_cnt_reg[2]/P0001 ,
		_w4762_
	);
	LUT4 #(
		.INIT('h008a)
	) name3013 (
		_w4757_,
		_w4760_,
		_w4761_,
		_w4762_,
		_w4763_
	);
	LUT2 #(
		.INIT('h1)
	) name3014 (
		\u4_u2_csr0_reg[6]/P0001 ,
		\u4_u2_dma_out_cnt_reg[4]/P0001 ,
		_w4764_
	);
	LUT4 #(
		.INIT('hfac8)
	) name3015 (
		\u4_u2_csr0_reg[6]/P0001 ,
		\u4_u2_csr0_reg[7]/P0001 ,
		\u4_u2_dma_out_cnt_reg[4]/P0001 ,
		\u4_u2_dma_out_cnt_reg[5]/P0001 ,
		_w4765_
	);
	LUT2 #(
		.INIT('h4)
	) name3016 (
		_w4755_,
		_w4765_,
		_w4766_
	);
	LUT4 #(
		.INIT('h5455)
	) name3017 (
		_w4756_,
		_w4758_,
		_w4763_,
		_w4766_,
		_w4767_
	);
	LUT4 #(
		.INIT('h135f)
	) name3018 (
		\u4_u2_csr0_reg[8]/P0001 ,
		\u4_u2_csr0_reg[9]/P0001 ,
		\u4_u2_dma_out_cnt_reg[6]/P0001 ,
		\u4_u2_dma_out_cnt_reg[7]/P0001 ,
		_w4768_
	);
	LUT4 #(
		.INIT('h5666)
	) name3019 (
		_w4753_,
		_w4754_,
		_w4767_,
		_w4768_,
		_w4769_
	);
	LUT3 #(
		.INIT('h02)
	) name3020 (
		_w4610_,
		_w4746_,
		_w4748_,
		_w4770_
	);
	LUT3 #(
		.INIT('h15)
	) name3021 (
		_w4752_,
		_w4769_,
		_w4770_,
		_w4771_
	);
	LUT4 #(
		.INIT('h0002)
	) name3022 (
		rst_i_pad,
		\u1_clr_sof_time_reg/P0001 ,
		\u1_hms_clk_reg/P0001 ,
		\u1_hms_cnt_reg[0]/P0001 ,
		_w4772_
	);
	LUT4 #(
		.INIT('h0001)
	) name3023 (
		\u0_u0_me_cnt_reg[4]/P0001 ,
		\u0_u0_me_cnt_reg[5]/P0001 ,
		\u0_u0_me_cnt_reg[6]/P0001 ,
		\u0_u0_me_cnt_reg[7]/P0001 ,
		_w4773_
	);
	LUT4 #(
		.INIT('h0007)
	) name3024 (
		\u0_u0_me_cnt_reg[0]/P0001 ,
		\u0_u0_me_cnt_reg[1]/P0001 ,
		\u0_u0_me_cnt_reg[2]/P0001 ,
		\u0_u0_me_cnt_reg[3]/P0001 ,
		_w4774_
	);
	LUT2 #(
		.INIT('h8)
	) name3025 (
		_w4773_,
		_w4774_,
		_w4775_
	);
	LUT2 #(
		.INIT('h2)
	) name3026 (
		_w4626_,
		_w4775_,
		_w4776_
	);
	LUT2 #(
		.INIT('h4)
	) name3027 (
		_w4350_,
		_w4776_,
		_w4777_
	);
	LUT4 #(
		.INIT('hf800)
	) name3028 (
		\u0_u0_me_cnt_reg[0]/P0001 ,
		\u0_u0_me_cnt_reg[1]/P0001 ,
		\u0_u0_me_cnt_reg[2]/P0001 ,
		\u0_u0_me_cnt_reg[3]/P0001 ,
		_w4778_
	);
	LUT2 #(
		.INIT('h2)
	) name3029 (
		_w4773_,
		_w4778_,
		_w4779_
	);
	LUT2 #(
		.INIT('h2)
	) name3030 (
		_w4626_,
		_w4779_,
		_w4780_
	);
	LUT2 #(
		.INIT('h4)
	) name3031 (
		_w4350_,
		_w4780_,
		_w4781_
	);
	LUT3 #(
		.INIT('h02)
	) name3032 (
		\u5_wb_ack_s1_reg/P0001 ,
		\u5_wb_ack_s2_reg/P0001 ,
		wb_ack_o_pad,
		_w4782_
	);
	LUT4 #(
		.INIT('h8000)
	) name3033 (
		\u1_u2_rx_data_valid_r_reg/NET0131 ,
		\u1_u2_sizu_c_reg[0]/P0001 ,
		\u1_u2_sizu_c_reg[1]/P0001 ,
		\u1_u2_sizu_c_reg[2]/P0001 ,
		_w4783_
	);
	LUT3 #(
		.INIT('h80)
	) name3034 (
		\u1_u2_sizu_c_reg[3]/P0001 ,
		\u1_u2_sizu_c_reg[4]/P0001 ,
		\u1_u2_sizu_c_reg[5]/P0001 ,
		_w4784_
	);
	LUT2 #(
		.INIT('h8)
	) name3035 (
		\u1_u2_sizu_c_reg[6]/P0001 ,
		\u1_u2_sizu_c_reg[7]/P0001 ,
		_w4785_
	);
	LUT4 #(
		.INIT('h1555)
	) name3036 (
		\u1_u2_sizu_c_reg[8]/NET0131 ,
		_w4783_,
		_w4784_,
		_w4785_,
		_w4786_
	);
	LUT2 #(
		.INIT('h2)
	) name3037 (
		rst_i_pad,
		\u1_u2_rx_dma_en_r_reg/P0001 ,
		_w4787_
	);
	LUT4 #(
		.INIT('h8000)
	) name3038 (
		\u1_u2_sizu_c_reg[3]/P0001 ,
		\u1_u2_sizu_c_reg[4]/P0001 ,
		\u1_u2_sizu_c_reg[5]/P0001 ,
		\u1_u2_sizu_c_reg[8]/NET0131 ,
		_w4788_
	);
	LUT4 #(
		.INIT('h70f0)
	) name3039 (
		_w4783_,
		_w4785_,
		_w4787_,
		_w4788_,
		_w4789_
	);
	LUT2 #(
		.INIT('h4)
	) name3040 (
		_w4786_,
		_w4789_,
		_w4790_
	);
	LUT3 #(
		.INIT('h14)
	) name3041 (
		\u0_u0_me_ps2_0_5_ms_reg/P0001 ,
		\u0_u0_me_ps2_reg[0]/P0001 ,
		\u0_u0_me_ps_2_5_us_reg/P0001 ,
		_w4791_
	);
	LUT2 #(
		.INIT('h8)
	) name3042 (
		_w4626_,
		_w4791_,
		_w4792_
	);
	LUT2 #(
		.INIT('h4)
	) name3043 (
		_w4350_,
		_w4792_,
		_w4793_
	);
	LUT4 #(
		.INIT('hebaf)
	) name3044 (
		\u0_u0_me_ps2_0_5_ms_reg/P0001 ,
		\u0_u0_me_ps2_reg[0]/P0001 ,
		\u0_u0_me_ps2_reg[1]/P0001 ,
		\u0_u0_me_ps_2_5_us_reg/P0001 ,
		_w4794_
	);
	LUT2 #(
		.INIT('h2)
	) name3045 (
		_w4626_,
		_w4794_,
		_w4795_
	);
	LUT2 #(
		.INIT('h4)
	) name3046 (
		_w4350_,
		_w4795_,
		_w4796_
	);
	LUT4 #(
		.INIT('h8000)
	) name3047 (
		\u0_u0_me_ps2_reg[0]/P0001 ,
		\u0_u0_me_ps2_reg[1]/P0001 ,
		\u0_u0_me_ps2_reg[2]/P0001 ,
		\u0_u0_me_ps_2_5_us_reg/P0001 ,
		_w4797_
	);
	LUT2 #(
		.INIT('h4)
	) name3048 (
		\u0_u0_me_ps2_0_5_ms_reg/P0001 ,
		\u0_u0_me_ps2_reg[2]/P0001 ,
		_w4798_
	);
	LUT4 #(
		.INIT('h4000)
	) name3049 (
		\u0_u0_me_ps2_0_5_ms_reg/P0001 ,
		\u0_u0_me_ps2_reg[0]/P0001 ,
		\u0_u0_me_ps2_reg[1]/P0001 ,
		\u0_u0_me_ps_2_5_us_reg/P0001 ,
		_w4799_
	);
	LUT3 #(
		.INIT('h54)
	) name3050 (
		_w4797_,
		_w4798_,
		_w4799_,
		_w4800_
	);
	LUT2 #(
		.INIT('h8)
	) name3051 (
		_w4626_,
		_w4800_,
		_w4801_
	);
	LUT2 #(
		.INIT('h4)
	) name3052 (
		_w4350_,
		_w4801_,
		_w4802_
	);
	LUT3 #(
		.INIT('heb)
	) name3053 (
		\u0_u0_me_ps2_0_5_ms_reg/P0001 ,
		\u0_u0_me_ps2_reg[3]/P0001 ,
		_w4797_,
		_w4803_
	);
	LUT2 #(
		.INIT('h2)
	) name3054 (
		_w4626_,
		_w4803_,
		_w4804_
	);
	LUT2 #(
		.INIT('h4)
	) name3055 (
		_w4350_,
		_w4804_,
		_w4805_
	);
	LUT2 #(
		.INIT('h8)
	) name3056 (
		\u0_u0_me_ps2_reg[3]/P0001 ,
		\u0_u0_me_ps2_reg[4]/P0001 ,
		_w4806_
	);
	LUT4 #(
		.INIT('h1450)
	) name3057 (
		\u0_u0_me_ps2_0_5_ms_reg/P0001 ,
		\u0_u0_me_ps2_reg[3]/P0001 ,
		\u0_u0_me_ps2_reg[4]/P0001 ,
		_w4797_,
		_w4807_
	);
	LUT2 #(
		.INIT('h8)
	) name3058 (
		_w4626_,
		_w4807_,
		_w4808_
	);
	LUT2 #(
		.INIT('h4)
	) name3059 (
		_w4350_,
		_w4808_,
		_w4809_
	);
	LUT3 #(
		.INIT('h15)
	) name3060 (
		\u0_u0_me_ps2_reg[5]/P0001 ,
		_w4797_,
		_w4806_,
		_w4810_
	);
	LUT3 #(
		.INIT('h80)
	) name3061 (
		\u0_u0_me_ps2_reg[3]/P0001 ,
		\u0_u0_me_ps2_reg[4]/P0001 ,
		\u0_u0_me_ps2_reg[5]/P0001 ,
		_w4811_
	);
	LUT3 #(
		.INIT('h15)
	) name3062 (
		\u0_u0_me_ps2_0_5_ms_reg/P0001 ,
		_w4797_,
		_w4811_,
		_w4812_
	);
	LUT2 #(
		.INIT('h4)
	) name3063 (
		_w4810_,
		_w4812_,
		_w4813_
	);
	LUT2 #(
		.INIT('h8)
	) name3064 (
		_w4358_,
		_w4813_,
		_w4814_
	);
	LUT2 #(
		.INIT('h4)
	) name3065 (
		_w4353_,
		_w4814_,
		_w4815_
	);
	LUT2 #(
		.INIT('h4)
	) name3066 (
		_w4350_,
		_w4815_,
		_w4816_
	);
	LUT4 #(
		.INIT('hebbb)
	) name3067 (
		\u0_u0_me_ps2_0_5_ms_reg/P0001 ,
		\u0_u0_me_ps2_reg[6]/P0001 ,
		_w4797_,
		_w4811_,
		_w4817_
	);
	LUT2 #(
		.INIT('h2)
	) name3068 (
		_w4358_,
		_w4817_,
		_w4818_
	);
	LUT2 #(
		.INIT('h4)
	) name3069 (
		_w4353_,
		_w4818_,
		_w4819_
	);
	LUT2 #(
		.INIT('h4)
	) name3070 (
		_w4350_,
		_w4819_,
		_w4820_
	);
	LUT4 #(
		.INIT('h1333)
	) name3071 (
		\u0_u0_me_ps2_reg[6]/P0001 ,
		\u0_u0_me_ps2_reg[7]/P0001 ,
		_w4797_,
		_w4811_,
		_w4821_
	);
	LUT2 #(
		.INIT('h8)
	) name3072 (
		\u0_u0_me_ps2_reg[6]/P0001 ,
		\u0_u0_me_ps2_reg[7]/P0001 ,
		_w4822_
	);
	LUT4 #(
		.INIT('h1555)
	) name3073 (
		\u0_u0_me_ps2_0_5_ms_reg/P0001 ,
		_w4797_,
		_w4811_,
		_w4822_,
		_w4823_
	);
	LUT2 #(
		.INIT('h4)
	) name3074 (
		_w4821_,
		_w4823_,
		_w4824_
	);
	LUT2 #(
		.INIT('h8)
	) name3075 (
		_w4358_,
		_w4824_,
		_w4825_
	);
	LUT2 #(
		.INIT('h4)
	) name3076 (
		_w4353_,
		_w4825_,
		_w4826_
	);
	LUT2 #(
		.INIT('h4)
	) name3077 (
		_w4350_,
		_w4826_,
		_w4827_
	);
	LUT3 #(
		.INIT('h14)
	) name3078 (
		\u0_u0_me_ps_2_5_us_reg/P0001 ,
		\u0_u0_me_ps_reg[0]/P0001 ,
		\u0_u0_me_ps_reg[1]/P0001 ,
		_w4828_
	);
	LUT2 #(
		.INIT('h8)
	) name3079 (
		_w4358_,
		_w4828_,
		_w4829_
	);
	LUT2 #(
		.INIT('h4)
	) name3080 (
		_w4353_,
		_w4829_,
		_w4830_
	);
	LUT2 #(
		.INIT('h4)
	) name3081 (
		_w4350_,
		_w4830_,
		_w4831_
	);
	LUT4 #(
		.INIT('heabf)
	) name3082 (
		\u0_u0_me_ps_2_5_us_reg/P0001 ,
		\u0_u0_me_ps_reg[0]/P0001 ,
		\u0_u0_me_ps_reg[1]/P0001 ,
		\u0_u0_me_ps_reg[2]/P0001 ,
		_w4832_
	);
	LUT2 #(
		.INIT('h2)
	) name3083 (
		_w4358_,
		_w4832_,
		_w4833_
	);
	LUT2 #(
		.INIT('h4)
	) name3084 (
		_w4353_,
		_w4833_,
		_w4834_
	);
	LUT2 #(
		.INIT('h4)
	) name3085 (
		_w4350_,
		_w4834_,
		_w4835_
	);
	LUT4 #(
		.INIT('h007f)
	) name3086 (
		\u0_u0_me_ps_reg[0]/P0001 ,
		\u0_u0_me_ps_reg[1]/P0001 ,
		\u0_u0_me_ps_reg[2]/P0001 ,
		\u0_u0_me_ps_reg[3]/P0001 ,
		_w4836_
	);
	LUT3 #(
		.INIT('h01)
	) name3087 (
		\u0_u0_me_ps_2_5_us_reg/P0001 ,
		_w4636_,
		_w4836_,
		_w4837_
	);
	LUT2 #(
		.INIT('h8)
	) name3088 (
		_w4358_,
		_w4837_,
		_w4838_
	);
	LUT2 #(
		.INIT('h4)
	) name3089 (
		_w4353_,
		_w4838_,
		_w4839_
	);
	LUT2 #(
		.INIT('h4)
	) name3090 (
		_w4350_,
		_w4839_,
		_w4840_
	);
	LUT3 #(
		.INIT('heb)
	) name3091 (
		\u0_u0_me_ps_2_5_us_reg/P0001 ,
		\u0_u0_me_ps_reg[4]/P0001 ,
		_w4636_,
		_w4841_
	);
	LUT2 #(
		.INIT('h2)
	) name3092 (
		_w4358_,
		_w4841_,
		_w4842_
	);
	LUT2 #(
		.INIT('h4)
	) name3093 (
		_w4353_,
		_w4842_,
		_w4843_
	);
	LUT2 #(
		.INIT('h4)
	) name3094 (
		_w4350_,
		_w4843_,
		_w4844_
	);
	LUT4 #(
		.INIT('h8000)
	) name3095 (
		\u1_hms_clk_reg/P0001 ,
		\u1_sof_time_reg[0]/P0001 ,
		\u1_sof_time_reg[1]/P0001 ,
		\u1_sof_time_reg[2]/P0001 ,
		_w4845_
	);
	LUT4 #(
		.INIT('h1333)
	) name3096 (
		\u1_sof_time_reg[6]/P0001 ,
		\u1_sof_time_reg[7]/P0001 ,
		_w4367_,
		_w4845_,
		_w4846_
	);
	LUT2 #(
		.INIT('h8)
	) name3097 (
		\u1_sof_time_reg[6]/P0001 ,
		\u1_sof_time_reg[7]/P0001 ,
		_w4847_
	);
	LUT4 #(
		.INIT('h1555)
	) name3098 (
		\u1_clr_sof_time_reg/P0001 ,
		_w4367_,
		_w4845_,
		_w4847_,
		_w4848_
	);
	LUT2 #(
		.INIT('h4)
	) name3099 (
		_w4846_,
		_w4848_,
		_w4849_
	);
	LUT2 #(
		.INIT('h8)
	) name3100 (
		\u1_u3_pid_seq_err_reg/P0001 ,
		\u1_u3_state_reg[4]/P0001 ,
		_w4850_
	);
	LUT4 #(
		.INIT('h0010)
	) name3101 (
		\u1_u3_abort_reg/P0001 ,
		\u1_u3_tx_data_to_reg/P0001 ,
		\u4_csr_reg[24]/P0001 ,
		\u4_csr_reg[25]/P0001 ,
		_w4851_
	);
	LUT4 #(
		.INIT('h2000)
	) name3102 (
		_w3671_,
		_w3672_,
		_w4850_,
		_w4851_,
		_w4852_
	);
	LUT2 #(
		.INIT('h8)
	) name3103 (
		_w3682_,
		_w4852_,
		_w4853_
	);
	LUT2 #(
		.INIT('h6)
	) name3104 (
		\u1_frame_no_r_reg[8]/P0001 ,
		\u1_u0_token1_reg[0]/P0001 ,
		_w4854_
	);
	LUT2 #(
		.INIT('h8)
	) name3105 (
		\u1_u0_token_valid_str1_reg/P0001 ,
		_w2131_,
		_w4855_
	);
	LUT4 #(
		.INIT('h0100)
	) name3106 (
		_w3743_,
		_w3746_,
		_w3747_,
		_w4855_,
		_w4856_
	);
	LUT2 #(
		.INIT('h6)
	) name3107 (
		\u1_frame_no_r_reg[7]/P0001 ,
		\u1_u0_token0_reg[7]/P0001 ,
		_w4857_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name3108 (
		\u1_frame_no_r_reg[4]/P0001 ,
		\u1_frame_no_r_reg[9]/P0001 ,
		\u1_u0_token0_reg[4]/P0001 ,
		\u1_u0_token1_reg[1]/P0001 ,
		_w4858_
	);
	LUT2 #(
		.INIT('h4)
	) name3109 (
		_w4857_,
		_w4858_,
		_w4859_
	);
	LUT4 #(
		.INIT('hcf45)
	) name3110 (
		\u1_frame_no_r_reg[10]/P0001 ,
		\u1_frame_no_r_reg[6]/P0001 ,
		\u1_u0_token0_reg[6]/P0001 ,
		\u1_u0_token1_reg[2]/P0001 ,
		_w4860_
	);
	LUT4 #(
		.INIT('h8acf)
	) name3111 (
		\u1_frame_no_r_reg[10]/P0001 ,
		\u1_frame_no_r_reg[1]/P0001 ,
		\u1_u0_token0_reg[1]/P0001 ,
		\u1_u0_token1_reg[2]/P0001 ,
		_w4861_
	);
	LUT4 #(
		.INIT('hf531)
	) name3112 (
		\u1_frame_no_r_reg[1]/P0001 ,
		\u1_frame_no_r_reg[2]/P0001 ,
		\u1_u0_token0_reg[1]/P0001 ,
		\u1_u0_token0_reg[2]/NET0131 ,
		_w4862_
	);
	LUT4 #(
		.INIT('h8caf)
	) name3113 (
		\u1_frame_no_r_reg[2]/P0001 ,
		\u1_frame_no_r_reg[5]/P0001 ,
		\u1_u0_token0_reg[2]/NET0131 ,
		\u1_u0_token0_reg[5]/NET0131 ,
		_w4863_
	);
	LUT4 #(
		.INIT('h8000)
	) name3114 (
		_w4860_,
		_w4861_,
		_w4862_,
		_w4863_,
		_w4864_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name3115 (
		\u1_frame_no_r_reg[0]/P0001 ,
		\u1_frame_no_r_reg[3]/P0001 ,
		\u1_u0_token0_reg[0]/NET0131 ,
		\u1_u0_token0_reg[3]/NET0131 ,
		_w4865_
	);
	LUT4 #(
		.INIT('haf23)
	) name3116 (
		\u1_frame_no_r_reg[0]/P0001 ,
		\u1_frame_no_r_reg[9]/P0001 ,
		\u1_u0_token0_reg[0]/NET0131 ,
		\u1_u0_token1_reg[1]/P0001 ,
		_w4866_
	);
	LUT4 #(
		.INIT('hf531)
	) name3117 (
		\u1_frame_no_r_reg[5]/P0001 ,
		\u1_frame_no_r_reg[6]/P0001 ,
		\u1_u0_token0_reg[5]/NET0131 ,
		\u1_u0_token0_reg[6]/P0001 ,
		_w4867_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name3118 (
		\u1_frame_no_r_reg[3]/P0001 ,
		\u1_frame_no_r_reg[4]/P0001 ,
		\u1_u0_token0_reg[3]/NET0131 ,
		\u1_u0_token0_reg[4]/P0001 ,
		_w4868_
	);
	LUT4 #(
		.INIT('h8000)
	) name3119 (
		_w4865_,
		_w4866_,
		_w4867_,
		_w4868_,
		_w4869_
	);
	LUT3 #(
		.INIT('h80)
	) name3120 (
		_w4859_,
		_w4864_,
		_w4869_,
		_w4870_
	);
	LUT4 #(
		.INIT('h8000)
	) name3121 (
		_w3735_,
		_w3739_,
		_w4856_,
		_w4870_,
		_w4871_
	);
	LUT2 #(
		.INIT('h4)
	) name3122 (
		_w4854_,
		_w4871_,
		_w4872_
	);
	LUT3 #(
		.INIT('hac)
	) name3123 (
		\sram_data_i[0]_pad ,
		\u4_dout_reg[0]/P0001 ,
		\wb_addr_i[17]_pad ,
		_w4873_
	);
	LUT3 #(
		.INIT('hac)
	) name3124 (
		\sram_data_i[1]_pad ,
		\u4_dout_reg[1]/P0001 ,
		\wb_addr_i[17]_pad ,
		_w4874_
	);
	LUT3 #(
		.INIT('hac)
	) name3125 (
		\sram_data_i[2]_pad ,
		\u4_dout_reg[2]/P0001 ,
		\wb_addr_i[17]_pad ,
		_w4875_
	);
	LUT3 #(
		.INIT('hac)
	) name3126 (
		\sram_data_i[3]_pad ,
		\u4_dout_reg[3]/P0001 ,
		\wb_addr_i[17]_pad ,
		_w4876_
	);
	LUT3 #(
		.INIT('ha6)
	) name3127 (
		\u1_u3_new_sizeb_reg[8]/P0001 ,
		_w2837_,
		_w2839_,
		_w4877_
	);
	LUT4 #(
		.INIT('h10ef)
	) name3128 (
		_w3451_,
		_w3455_,
		_w3462_,
		_w4877_,
		_w4878_
	);
	LUT3 #(
		.INIT('ha6)
	) name3129 (
		\u1_u3_new_sizeb_reg[9]/P0001 ,
		_w2852_,
		_w2854_,
		_w4879_
	);
	LUT3 #(
		.INIT('h87)
	) name3130 (
		_w3509_,
		_w3511_,
		_w4879_,
		_w4880_
	);
	LUT4 #(
		.INIT('h0004)
	) name3131 (
		\u1_u0_state_reg[0]/P0001 ,
		\u1_u0_state_reg[1]/P0001 ,
		\u1_u0_state_reg[2]/P0001 ,
		\u1_u0_state_reg[3]/P0001 ,
		_w4881_
	);
	LUT3 #(
		.INIT('hb0)
	) name3132 (
		\u0_rx_err_reg/P0001 ,
		_w3695_,
		_w4881_,
		_w4882_
	);
	LUT2 #(
		.INIT('h8)
	) name3133 (
		\u0_rx_active_reg/P0001 ,
		\u0_rx_valid_reg/P0001 ,
		_w4883_
	);
	LUT3 #(
		.INIT('h20)
	) name3134 (
		\u0_rx_active_reg/P0001 ,
		\u0_rx_err_reg/P0001 ,
		\u0_rx_valid_reg/P0001 ,
		_w4884_
	);
	LUT4 #(
		.INIT('hddcd)
	) name3135 (
		\u1_u0_pid_reg[0]/NET0131 ,
		\u1_u0_pid_reg[1]/NET0131 ,
		\u1_u0_pid_reg[2]/NET0131 ,
		\u1_u0_pid_reg[3]/NET0131 ,
		_w4885_
	);
	LUT2 #(
		.INIT('h2)
	) name3136 (
		_w4884_,
		_w4885_,
		_w4886_
	);
	LUT2 #(
		.INIT('h8)
	) name3137 (
		_w4882_,
		_w4886_,
		_w4887_
	);
	LUT4 #(
		.INIT('h0010)
	) name3138 (
		\u1_u0_state_reg[0]/P0001 ,
		\u1_u0_state_reg[1]/P0001 ,
		\u1_u0_state_reg[2]/P0001 ,
		\u1_u0_state_reg[3]/P0001 ,
		_w4888_
	);
	LUT2 #(
		.INIT('h8)
	) name3139 (
		\u0_rx_active_reg/P0001 ,
		\u1_u0_state_reg[2]/P0001 ,
		_w4889_
	);
	LUT4 #(
		.INIT('hba00)
	) name3140 (
		_w3671_,
		_w4884_,
		_w4888_,
		_w4889_,
		_w4890_
	);
	LUT4 #(
		.INIT('haa80)
	) name3141 (
		rst_i_pad,
		_w4882_,
		_w4886_,
		_w4890_,
		_w4891_
	);
	LUT4 #(
		.INIT('h0010)
	) name3142 (
		\u4_u3_r5_reg/NET0131 ,
		_w4402_,
		_w4403_,
		_w4404_,
		_w4892_
	);
	LUT2 #(
		.INIT('h1)
	) name3143 (
		\u4_u3_dma_in_cnt_reg[10]/P0001 ,
		_w4892_,
		_w4893_
	);
	LUT3 #(
		.INIT('h04)
	) name3144 (
		\u4_u3_dma_in_cnt_reg[10]/P0001 ,
		_w4394_,
		_w4395_,
		_w4894_
	);
	LUT3 #(
		.INIT('hb0)
	) name3145 (
		_w4390_,
		_w4393_,
		_w4894_,
		_w4895_
	);
	LUT2 #(
		.INIT('h1)
	) name3146 (
		\u4_u3_dma_in_cnt_reg[10]/P0001 ,
		\u4_u3_dma_in_cnt_reg[9]/P0001 ,
		_w4896_
	);
	LUT3 #(
		.INIT('h0e)
	) name3147 (
		\u4_u3_dma_in_cnt_reg[10]/P0001 ,
		\u4_u3_dma_in_cnt_reg[9]/P0001 ,
		\u4_u3_r5_reg/NET0131 ,
		_w4897_
	);
	LUT3 #(
		.INIT('h01)
	) name3148 (
		\u4_u3_dma_in_cnt_reg[10]/P0001 ,
		\u4_u3_dma_in_cnt_reg[9]/P0001 ,
		\u4_u3_r5_reg/NET0131 ,
		_w4898_
	);
	LUT3 #(
		.INIT('h80)
	) name3149 (
		\u4_u3_dma_in_cnt_reg[7]/P0001 ,
		\u4_u3_dma_in_cnt_reg[8]/P0001 ,
		\u4_u3_dma_in_cnt_reg[9]/P0001 ,
		_w4899_
	);
	LUT4 #(
		.INIT('h0800)
	) name3150 (
		_w4398_,
		_w4399_,
		_w4897_,
		_w4899_,
		_w4900_
	);
	LUT3 #(
		.INIT('ha8)
	) name3151 (
		\u4_u3_dma_in_cnt_reg[11]/P0001 ,
		_w4898_,
		_w4900_,
		_w4901_
	);
	LUT3 #(
		.INIT('h10)
	) name3152 (
		_w4893_,
		_w4895_,
		_w4901_,
		_w4902_
	);
	LUT4 #(
		.INIT('haaa8)
	) name3153 (
		\u4_u3_csr1_reg[0]/P0001 ,
		\u4_u3_dma_in_cnt_reg[11]/P0001 ,
		_w4898_,
		_w4900_,
		_w4903_
	);
	LUT4 #(
		.INIT('hab00)
	) name3154 (
		\u4_u3_dma_in_cnt_reg[11]/P0001 ,
		_w4893_,
		_w4895_,
		_w4903_,
		_w4904_
	);
	LUT2 #(
		.INIT('h4)
	) name3155 (
		_w4902_,
		_w4904_,
		_w4905_
	);
	LUT4 #(
		.INIT('h0010)
	) name3156 (
		\u4_u0_r5_reg/NET0131 ,
		_w4434_,
		_w4435_,
		_w4436_,
		_w4906_
	);
	LUT2 #(
		.INIT('h1)
	) name3157 (
		\u4_u0_dma_in_cnt_reg[10]/P0001 ,
		_w4906_,
		_w4907_
	);
	LUT3 #(
		.INIT('h04)
	) name3158 (
		\u4_u0_dma_in_cnt_reg[10]/P0001 ,
		_w4426_,
		_w4427_,
		_w4908_
	);
	LUT3 #(
		.INIT('hb0)
	) name3159 (
		_w4422_,
		_w4425_,
		_w4908_,
		_w4909_
	);
	LUT2 #(
		.INIT('h1)
	) name3160 (
		\u4_u0_dma_in_cnt_reg[10]/P0001 ,
		\u4_u0_dma_in_cnt_reg[9]/P0001 ,
		_w4910_
	);
	LUT3 #(
		.INIT('h0e)
	) name3161 (
		\u4_u0_dma_in_cnt_reg[10]/P0001 ,
		\u4_u0_dma_in_cnt_reg[9]/P0001 ,
		\u4_u0_r5_reg/NET0131 ,
		_w4911_
	);
	LUT3 #(
		.INIT('h01)
	) name3162 (
		\u4_u0_dma_in_cnt_reg[10]/P0001 ,
		\u4_u0_dma_in_cnt_reg[9]/P0001 ,
		\u4_u0_r5_reg/NET0131 ,
		_w4912_
	);
	LUT3 #(
		.INIT('h80)
	) name3163 (
		\u4_u0_dma_in_cnt_reg[7]/P0001 ,
		\u4_u0_dma_in_cnt_reg[8]/P0001 ,
		\u4_u0_dma_in_cnt_reg[9]/P0001 ,
		_w4913_
	);
	LUT4 #(
		.INIT('h0800)
	) name3164 (
		_w4430_,
		_w4431_,
		_w4911_,
		_w4913_,
		_w4914_
	);
	LUT3 #(
		.INIT('ha8)
	) name3165 (
		\u4_u0_dma_in_cnt_reg[11]/P0001 ,
		_w4912_,
		_w4914_,
		_w4915_
	);
	LUT3 #(
		.INIT('h10)
	) name3166 (
		_w4907_,
		_w4909_,
		_w4915_,
		_w4916_
	);
	LUT4 #(
		.INIT('haaa8)
	) name3167 (
		\u4_u0_csr1_reg[0]/P0001 ,
		\u4_u0_dma_in_cnt_reg[11]/P0001 ,
		_w4912_,
		_w4914_,
		_w4917_
	);
	LUT4 #(
		.INIT('hab00)
	) name3168 (
		\u4_u0_dma_in_cnt_reg[11]/P0001 ,
		_w4907_,
		_w4909_,
		_w4917_,
		_w4918_
	);
	LUT2 #(
		.INIT('h4)
	) name3169 (
		_w4916_,
		_w4918_,
		_w4919_
	);
	LUT3 #(
		.INIT('h0b)
	) name3170 (
		\u4_u1_csr0_reg[10]/P0001 ,
		\u4_u1_dma_in_cnt_reg[8]/P0001 ,
		\u4_u1_r5_reg/NET0131 ,
		_w4920_
	);
	LUT4 #(
		.INIT('h5155)
	) name3171 (
		\u4_u1_dma_in_cnt_reg[10]/P0001 ,
		_w4454_,
		_w4455_,
		_w4920_,
		_w4921_
	);
	LUT3 #(
		.INIT('h04)
	) name3172 (
		\u4_u1_dma_in_cnt_reg[10]/P0001 ,
		_w4473_,
		_w4474_,
		_w4922_
	);
	LUT3 #(
		.INIT('h0e)
	) name3173 (
		\u4_u1_dma_in_cnt_reg[10]/P0001 ,
		\u4_u1_dma_in_cnt_reg[9]/P0001 ,
		\u4_u1_r5_reg/NET0131 ,
		_w4923_
	);
	LUT3 #(
		.INIT('h01)
	) name3174 (
		\u4_u1_dma_in_cnt_reg[10]/P0001 ,
		\u4_u1_dma_in_cnt_reg[9]/P0001 ,
		\u4_u1_r5_reg/NET0131 ,
		_w4924_
	);
	LUT3 #(
		.INIT('h80)
	) name3175 (
		\u4_u1_dma_in_cnt_reg[7]/P0001 ,
		\u4_u1_dma_in_cnt_reg[8]/P0001 ,
		\u4_u1_dma_in_cnt_reg[9]/P0001 ,
		_w4925_
	);
	LUT4 #(
		.INIT('h0800)
	) name3176 (
		_w4447_,
		_w4448_,
		_w4923_,
		_w4925_,
		_w4926_
	);
	LUT3 #(
		.INIT('ha8)
	) name3177 (
		\u4_u1_dma_in_cnt_reg[11]/P0001 ,
		_w4924_,
		_w4926_,
		_w4927_
	);
	LUT4 #(
		.INIT('h1300)
	) name3178 (
		_w4471_,
		_w4921_,
		_w4922_,
		_w4927_,
		_w4928_
	);
	LUT2 #(
		.INIT('h1)
	) name3179 (
		\u4_u1_dma_in_cnt_reg[10]/P0001 ,
		\u4_u1_dma_in_cnt_reg[11]/P0001 ,
		_w4929_
	);
	LUT4 #(
		.INIT('hdf00)
	) name3180 (
		_w4454_,
		_w4455_,
		_w4920_,
		_w4929_,
		_w4930_
	);
	LUT3 #(
		.INIT('h20)
	) name3181 (
		_w4473_,
		_w4474_,
		_w4929_,
		_w4931_
	);
	LUT4 #(
		.INIT('haaa8)
	) name3182 (
		\u4_u1_csr1_reg[0]/P0001 ,
		\u4_u1_dma_in_cnt_reg[11]/P0001 ,
		_w4924_,
		_w4926_,
		_w4932_
	);
	LUT4 #(
		.INIT('h1300)
	) name3183 (
		_w4471_,
		_w4930_,
		_w4931_,
		_w4932_,
		_w4933_
	);
	LUT2 #(
		.INIT('h4)
	) name3184 (
		_w4928_,
		_w4933_,
		_w4934_
	);
	LUT3 #(
		.INIT('h0e)
	) name3185 (
		\u4_u2_dma_in_cnt_reg[10]/P0001 ,
		\u4_u2_dma_in_cnt_reg[9]/P0001 ,
		\u4_u2_r5_reg/NET0131 ,
		_w4935_
	);
	LUT4 #(
		.INIT('h0800)
	) name3186 (
		_w4504_,
		_w4505_,
		_w4935_,
		_w4507_,
		_w4936_
	);
	LUT3 #(
		.INIT('h51)
	) name3187 (
		\u4_u2_r5_reg/NET0131 ,
		_w4935_,
		_w4936_,
		_w4937_
	);
	LUT4 #(
		.INIT('h1500)
	) name3188 (
		_w4486_,
		_w4499_,
		_w4501_,
		_w4937_,
		_w4938_
	);
	LUT2 #(
		.INIT('h8)
	) name3189 (
		\u4_u2_dma_in_cnt_reg[10]/P0001 ,
		\u4_u2_r5_reg/NET0131 ,
		_w4939_
	);
	LUT4 #(
		.INIT('h8000)
	) name3190 (
		_w4504_,
		_w4505_,
		_w4507_,
		_w4939_,
		_w4940_
	);
	LUT2 #(
		.INIT('h8)
	) name3191 (
		\u4_u2_csr1_reg[0]/P0001 ,
		\u4_u2_dma_in_cnt_reg[11]/P0001 ,
		_w4941_
	);
	LUT2 #(
		.INIT('h4)
	) name3192 (
		_w4940_,
		_w4941_,
		_w4942_
	);
	LUT2 #(
		.INIT('h4)
	) name3193 (
		_w4938_,
		_w4942_,
		_w4943_
	);
	LUT2 #(
		.INIT('h2)
	) name3194 (
		\u4_u2_csr1_reg[0]/P0001 ,
		\u4_u2_dma_in_cnt_reg[11]/P0001 ,
		_w4944_
	);
	LUT3 #(
		.INIT('h01)
	) name3195 (
		\u4_u2_dma_in_cnt_reg[10]/P0001 ,
		\u4_u2_dma_in_cnt_reg[9]/P0001 ,
		\u4_u2_r5_reg/NET0131 ,
		_w4945_
	);
	LUT4 #(
		.INIT('h1500)
	) name3196 (
		_w4486_,
		_w4499_,
		_w4501_,
		_w4945_,
		_w4946_
	);
	LUT3 #(
		.INIT('hc8)
	) name3197 (
		_w4940_,
		_w4944_,
		_w4946_,
		_w4947_
	);
	LUT2 #(
		.INIT('he)
	) name3198 (
		_w4943_,
		_w4947_,
		_w4948_
	);
	LUT3 #(
		.INIT('he0)
	) name3199 (
		\u4_u3_csr0_reg[10]/P0001 ,
		\u4_u3_dma_out_cnt_reg[8]/P0001 ,
		\u4_u3_dma_out_cnt_reg[9]/P0001 ,
		_w4949_
	);
	LUT3 #(
		.INIT('h80)
	) name3200 (
		\u4_u3_csr0_reg[10]/P0001 ,
		\u4_u3_dma_out_cnt_reg[8]/P0001 ,
		\u4_u3_dma_out_cnt_reg[9]/P0001 ,
		_w4950_
	);
	LUT3 #(
		.INIT('h0b)
	) name3201 (
		_w4663_,
		_w4949_,
		_w4950_,
		_w4951_
	);
	LUT2 #(
		.INIT('h2)
	) name3202 (
		_w4677_,
		_w4950_,
		_w4952_
	);
	LUT2 #(
		.INIT('h1)
	) name3203 (
		\u4_u3_dma_out_cnt_reg[4]/P0001 ,
		\u4_u3_dma_out_cnt_reg[5]/P0001 ,
		_w4953_
	);
	LUT4 #(
		.INIT('h0001)
	) name3204 (
		\u4_u3_dma_out_cnt_reg[6]/P0001 ,
		\u4_u3_dma_out_cnt_reg[7]/P0001 ,
		\u4_u3_dma_out_cnt_reg[8]/P0001 ,
		\u4_u3_dma_out_cnt_reg[9]/P0001 ,
		_w4954_
	);
	LUT4 #(
		.INIT('h4000)
	) name3205 (
		\u4_u3_dma_out_cnt_reg[10]/P0001 ,
		_w4652_,
		_w4953_,
		_w4954_,
		_w4955_
	);
	LUT2 #(
		.INIT('h8)
	) name3206 (
		\u4_u3_dma_out_cnt_reg[10]/P0001 ,
		\u4_u3_ep_match_r_reg/P0001 ,
		_w4956_
	);
	LUT2 #(
		.INIT('h4)
	) name3207 (
		_w4402_,
		_w4956_,
		_w4957_
	);
	LUT3 #(
		.INIT('hd0)
	) name3208 (
		\u4_u3_r5_reg/NET0131 ,
		_w4955_,
		_w4957_,
		_w4958_
	);
	LUT4 #(
		.INIT('h1300)
	) name3209 (
		_w4676_,
		_w4951_,
		_w4952_,
		_w4958_,
		_w4959_
	);
	LUT2 #(
		.INIT('h4)
	) name3210 (
		\u4_u3_dma_out_cnt_reg[10]/P0001 ,
		\u4_u3_r5_reg/NET0131 ,
		_w4960_
	);
	LUT4 #(
		.INIT('h8000)
	) name3211 (
		_w4652_,
		_w4953_,
		_w4954_,
		_w4960_,
		_w4961_
	);
	LUT2 #(
		.INIT('h8)
	) name3212 (
		\u4_u3_csr1_reg[0]/P0001 ,
		\u4_u3_dma_out_cnt_reg[11]/P0001 ,
		_w4962_
	);
	LUT2 #(
		.INIT('h4)
	) name3213 (
		_w4961_,
		_w4962_,
		_w4963_
	);
	LUT2 #(
		.INIT('h2)
	) name3214 (
		\u4_u3_csr1_reg[0]/P0001 ,
		\u4_u3_dma_out_cnt_reg[11]/P0001 ,
		_w4964_
	);
	LUT2 #(
		.INIT('h8)
	) name3215 (
		_w4961_,
		_w4964_,
		_w4965_
	);
	LUT4 #(
		.INIT('hd000)
	) name3216 (
		\u4_u3_r5_reg/NET0131 ,
		_w4955_,
		_w4957_,
		_w4964_,
		_w4966_
	);
	LUT4 #(
		.INIT('h1300)
	) name3217 (
		_w4676_,
		_w4951_,
		_w4952_,
		_w4966_,
		_w4967_
	);
	LUT4 #(
		.INIT('hfff4)
	) name3218 (
		_w4959_,
		_w4963_,
		_w4965_,
		_w4967_,
		_w4968_
	);
	LUT4 #(
		.INIT('h0157)
	) name3219 (
		\u4_u3_csr0_reg[10]/P0001 ,
		\u4_u3_csr0_reg[9]/P0001 ,
		\u4_u3_dma_out_cnt_reg[7]/P0001 ,
		\u4_u3_dma_out_cnt_reg[8]/P0001 ,
		_w4969_
	);
	LUT2 #(
		.INIT('h4)
	) name3220 (
		_w4661_,
		_w4677_,
		_w4970_
	);
	LUT4 #(
		.INIT('h5450)
	) name3221 (
		\u4_u3_r5_reg/NET0131 ,
		_w4676_,
		_w4969_,
		_w4970_,
		_w4971_
	);
	LUT2 #(
		.INIT('h4)
	) name3222 (
		\u4_u3_r5_reg/NET0131 ,
		_w4569_,
		_w4972_
	);
	LUT3 #(
		.INIT('h80)
	) name3223 (
		_w4650_,
		_w4652_,
		_w4653_,
		_w4973_
	);
	LUT3 #(
		.INIT('ha8)
	) name3224 (
		\u4_u3_dma_out_cnt_reg[9]/P0001 ,
		_w4972_,
		_w4973_,
		_w4974_
	);
	LUT2 #(
		.INIT('h1)
	) name3225 (
		\u4_u3_dma_out_cnt_reg[9]/P0001 ,
		\u4_u3_r5_reg/NET0131 ,
		_w4975_
	);
	LUT4 #(
		.INIT('hec00)
	) name3226 (
		_w4676_,
		_w4969_,
		_w4970_,
		_w4975_,
		_w4976_
	);
	LUT4 #(
		.INIT('haaa8)
	) name3227 (
		\u4_u3_csr1_reg[0]/P0001 ,
		\u4_u3_dma_out_cnt_reg[9]/P0001 ,
		_w4972_,
		_w4973_,
		_w4977_
	);
	LUT4 #(
		.INIT('h0b00)
	) name3228 (
		_w4971_,
		_w4974_,
		_w4976_,
		_w4977_,
		_w4978_
	);
	LUT3 #(
		.INIT('he0)
	) name3229 (
		\u4_u0_csr0_reg[10]/P0001 ,
		\u4_u0_dma_out_cnt_reg[8]/P0001 ,
		\u4_u0_dma_out_cnt_reg[9]/P0001 ,
		_w4979_
	);
	LUT3 #(
		.INIT('h80)
	) name3230 (
		\u4_u0_csr0_reg[10]/P0001 ,
		\u4_u0_dma_out_cnt_reg[8]/P0001 ,
		\u4_u0_dma_out_cnt_reg[9]/P0001 ,
		_w4980_
	);
	LUT3 #(
		.INIT('h0b)
	) name3231 (
		_w4693_,
		_w4979_,
		_w4980_,
		_w4981_
	);
	LUT2 #(
		.INIT('h2)
	) name3232 (
		_w4707_,
		_w4980_,
		_w4982_
	);
	LUT2 #(
		.INIT('h1)
	) name3233 (
		\u4_u0_dma_out_cnt_reg[4]/P0001 ,
		\u4_u0_dma_out_cnt_reg[5]/P0001 ,
		_w4983_
	);
	LUT4 #(
		.INIT('h0001)
	) name3234 (
		\u4_u0_dma_out_cnt_reg[6]/P0001 ,
		\u4_u0_dma_out_cnt_reg[7]/P0001 ,
		\u4_u0_dma_out_cnt_reg[8]/P0001 ,
		\u4_u0_dma_out_cnt_reg[9]/P0001 ,
		_w4984_
	);
	LUT4 #(
		.INIT('h4000)
	) name3235 (
		\u4_u0_dma_out_cnt_reg[10]/P0001 ,
		_w4683_,
		_w4983_,
		_w4984_,
		_w4985_
	);
	LUT2 #(
		.INIT('h8)
	) name3236 (
		\u4_u0_dma_out_cnt_reg[10]/P0001 ,
		\u4_u0_ep_match_r_reg/P0001 ,
		_w4986_
	);
	LUT4 #(
		.INIT('h3100)
	) name3237 (
		\u4_u0_r5_reg/NET0131 ,
		_w4434_,
		_w4985_,
		_w4986_,
		_w4987_
	);
	LUT4 #(
		.INIT('h1300)
	) name3238 (
		_w4706_,
		_w4981_,
		_w4982_,
		_w4987_,
		_w4988_
	);
	LUT3 #(
		.INIT('h10)
	) name3239 (
		\u4_u0_dma_out_cnt_reg[4]/P0001 ,
		\u4_u0_dma_out_cnt_reg[5]/P0001 ,
		\u4_u0_r5_reg/NET0131 ,
		_w4989_
	);
	LUT4 #(
		.INIT('h4000)
	) name3240 (
		\u4_u0_dma_out_cnt_reg[10]/P0001 ,
		_w4683_,
		_w4984_,
		_w4989_,
		_w4990_
	);
	LUT2 #(
		.INIT('h8)
	) name3241 (
		\u4_u0_csr1_reg[0]/P0001 ,
		\u4_u0_dma_out_cnt_reg[11]/P0001 ,
		_w4991_
	);
	LUT2 #(
		.INIT('h4)
	) name3242 (
		_w4990_,
		_w4991_,
		_w4992_
	);
	LUT2 #(
		.INIT('h2)
	) name3243 (
		\u4_u0_csr1_reg[0]/P0001 ,
		\u4_u0_dma_out_cnt_reg[11]/P0001 ,
		_w4993_
	);
	LUT2 #(
		.INIT('h4)
	) name3244 (
		\u4_u0_dma_out_cnt_reg[10]/P0001 ,
		\u4_u0_r5_reg/NET0131 ,
		_w4994_
	);
	LUT4 #(
		.INIT('h8000)
	) name3245 (
		_w4683_,
		_w4983_,
		_w4984_,
		_w4994_,
		_w4995_
	);
	LUT4 #(
		.INIT('hf4e4)
	) name3246 (
		_w4988_,
		_w4992_,
		_w4993_,
		_w4995_,
		_w4996_
	);
	LUT4 #(
		.INIT('hfca8)
	) name3247 (
		\u4_u0_csr0_reg[10]/P0001 ,
		\u4_u0_csr0_reg[9]/P0001 ,
		\u4_u0_dma_out_cnt_reg[7]/P0001 ,
		\u4_u0_dma_out_cnt_reg[8]/P0001 ,
		_w4997_
	);
	LUT3 #(
		.INIT('h07)
	) name3248 (
		\u4_u0_csr0_reg[10]/P0001 ,
		\u4_u0_dma_out_cnt_reg[8]/P0001 ,
		\u4_u0_r5_reg/NET0131 ,
		_w4998_
	);
	LUT4 #(
		.INIT('h8f00)
	) name3249 (
		_w4706_,
		_w4707_,
		_w4997_,
		_w4998_,
		_w4999_
	);
	LUT2 #(
		.INIT('h1)
	) name3250 (
		\u4_u0_dma_out_cnt_reg[7]/P0001 ,
		\u4_u0_dma_out_cnt_reg[8]/P0001 ,
		_w5000_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name3251 (
		\u4_u0_r5_reg/NET0131 ,
		_w4681_,
		_w4683_,
		_w5000_,
		_w5001_
	);
	LUT2 #(
		.INIT('h1)
	) name3252 (
		\u4_u0_ep_match_r_reg/P0001 ,
		\u4_u0_r5_reg/NET0131 ,
		_w5002_
	);
	LUT4 #(
		.INIT('h0001)
	) name3253 (
		\u1_u3_buf0_rl_reg/P0001 ,
		\u1_u3_buf0_set_reg/P0001 ,
		\u4_u0_r5_reg/NET0131 ,
		\u4_u0_set_r_reg/P0001 ,
		_w5003_
	);
	LUT3 #(
		.INIT('h02)
	) name3254 (
		\u4_u0_dma_out_cnt_reg[9]/P0001 ,
		_w5002_,
		_w5003_,
		_w5004_
	);
	LUT2 #(
		.INIT('h4)
	) name3255 (
		_w5001_,
		_w5004_,
		_w5005_
	);
	LUT4 #(
		.INIT('h0007)
	) name3256 (
		\u4_u0_csr0_reg[10]/P0001 ,
		\u4_u0_dma_out_cnt_reg[8]/P0001 ,
		\u4_u0_dma_out_cnt_reg[9]/P0001 ,
		\u4_u0_r5_reg/NET0131 ,
		_w5006_
	);
	LUT4 #(
		.INIT('h8f00)
	) name3257 (
		_w4706_,
		_w4707_,
		_w4997_,
		_w5006_,
		_w5007_
	);
	LUT3 #(
		.INIT('h54)
	) name3258 (
		\u4_u0_dma_out_cnt_reg[9]/P0001 ,
		_w5002_,
		_w5003_,
		_w5008_
	);
	LUT2 #(
		.INIT('h4)
	) name3259 (
		\u4_u0_dma_out_cnt_reg[9]/P0001 ,
		\u4_u0_r5_reg/NET0131 ,
		_w5009_
	);
	LUT4 #(
		.INIT('h7f00)
	) name3260 (
		_w4681_,
		_w4683_,
		_w5000_,
		_w5009_,
		_w5010_
	);
	LUT3 #(
		.INIT('h02)
	) name3261 (
		\u4_u0_csr1_reg[0]/P0001 ,
		_w5008_,
		_w5010_,
		_w5011_
	);
	LUT4 #(
		.INIT('h0b00)
	) name3262 (
		_w4999_,
		_w5005_,
		_w5007_,
		_w5011_,
		_w5012_
	);
	LUT3 #(
		.INIT('he0)
	) name3263 (
		\u4_u1_csr0_reg[10]/P0001 ,
		\u4_u1_dma_out_cnt_reg[8]/P0001 ,
		\u4_u1_dma_out_cnt_reg[9]/P0001 ,
		_w5013_
	);
	LUT3 #(
		.INIT('h80)
	) name3264 (
		\u4_u1_csr0_reg[10]/P0001 ,
		\u4_u1_dma_out_cnt_reg[8]/P0001 ,
		\u4_u1_dma_out_cnt_reg[9]/P0001 ,
		_w5014_
	);
	LUT3 #(
		.INIT('h0b)
	) name3265 (
		_w4724_,
		_w5013_,
		_w5014_,
		_w5015_
	);
	LUT2 #(
		.INIT('h2)
	) name3266 (
		_w4738_,
		_w5014_,
		_w5016_
	);
	LUT2 #(
		.INIT('h1)
	) name3267 (
		\u4_u1_dma_out_cnt_reg[4]/P0001 ,
		\u4_u1_dma_out_cnt_reg[5]/P0001 ,
		_w5017_
	);
	LUT4 #(
		.INIT('h0001)
	) name3268 (
		\u4_u1_dma_out_cnt_reg[6]/P0001 ,
		\u4_u1_dma_out_cnt_reg[7]/P0001 ,
		\u4_u1_dma_out_cnt_reg[8]/P0001 ,
		\u4_u1_dma_out_cnt_reg[9]/P0001 ,
		_w5018_
	);
	LUT4 #(
		.INIT('h4000)
	) name3269 (
		\u4_u1_dma_out_cnt_reg[10]/P0001 ,
		_w4713_,
		_w5017_,
		_w5018_,
		_w5019_
	);
	LUT2 #(
		.INIT('h8)
	) name3270 (
		\u4_u1_dma_out_cnt_reg[10]/P0001 ,
		\u4_u1_ep_match_r_reg/P0001 ,
		_w5020_
	);
	LUT4 #(
		.INIT('h3100)
	) name3271 (
		\u4_u1_r5_reg/NET0131 ,
		_w4453_,
		_w5019_,
		_w5020_,
		_w5021_
	);
	LUT4 #(
		.INIT('h1300)
	) name3272 (
		_w4737_,
		_w5015_,
		_w5016_,
		_w5021_,
		_w5022_
	);
	LUT3 #(
		.INIT('h10)
	) name3273 (
		\u4_u1_dma_out_cnt_reg[4]/P0001 ,
		\u4_u1_dma_out_cnt_reg[5]/P0001 ,
		\u4_u1_r5_reg/NET0131 ,
		_w5023_
	);
	LUT4 #(
		.INIT('h4000)
	) name3274 (
		\u4_u1_dma_out_cnt_reg[10]/P0001 ,
		_w4713_,
		_w5018_,
		_w5023_,
		_w5024_
	);
	LUT2 #(
		.INIT('h8)
	) name3275 (
		\u4_u1_csr1_reg[0]/P0001 ,
		\u4_u1_dma_out_cnt_reg[11]/P0001 ,
		_w5025_
	);
	LUT2 #(
		.INIT('h4)
	) name3276 (
		_w5024_,
		_w5025_,
		_w5026_
	);
	LUT2 #(
		.INIT('h2)
	) name3277 (
		\u4_u1_csr1_reg[0]/P0001 ,
		\u4_u1_dma_out_cnt_reg[11]/P0001 ,
		_w5027_
	);
	LUT2 #(
		.INIT('h4)
	) name3278 (
		\u4_u1_dma_out_cnt_reg[10]/P0001 ,
		\u4_u1_r5_reg/NET0131 ,
		_w5028_
	);
	LUT4 #(
		.INIT('h8000)
	) name3279 (
		_w4713_,
		_w5017_,
		_w5018_,
		_w5028_,
		_w5029_
	);
	LUT4 #(
		.INIT('hf4e4)
	) name3280 (
		_w5022_,
		_w5026_,
		_w5027_,
		_w5029_,
		_w5030_
	);
	LUT4 #(
		.INIT('h0157)
	) name3281 (
		\u4_u1_csr0_reg[10]/P0001 ,
		\u4_u1_csr0_reg[9]/P0001 ,
		\u4_u1_dma_out_cnt_reg[7]/P0001 ,
		\u4_u1_dma_out_cnt_reg[8]/P0001 ,
		_w5031_
	);
	LUT2 #(
		.INIT('h4)
	) name3282 (
		_w4722_,
		_w4738_,
		_w5032_
	);
	LUT4 #(
		.INIT('h5450)
	) name3283 (
		\u4_u1_r5_reg/NET0131 ,
		_w4737_,
		_w5031_,
		_w5032_,
		_w5033_
	);
	LUT2 #(
		.INIT('h1)
	) name3284 (
		\u4_u1_dma_out_cnt_reg[7]/P0001 ,
		\u4_u1_dma_out_cnt_reg[8]/P0001 ,
		_w5034_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name3285 (
		\u4_u1_r5_reg/NET0131 ,
		_w4711_,
		_w4713_,
		_w5034_,
		_w5035_
	);
	LUT2 #(
		.INIT('h1)
	) name3286 (
		\u4_u1_ep_match_r_reg/P0001 ,
		\u4_u1_r5_reg/NET0131 ,
		_w5036_
	);
	LUT4 #(
		.INIT('h0001)
	) name3287 (
		\u1_u3_buf0_rl_reg/P0001 ,
		\u1_u3_buf0_set_reg/P0001 ,
		\u4_u1_r5_reg/NET0131 ,
		\u4_u1_set_r_reg/P0001 ,
		_w5037_
	);
	LUT3 #(
		.INIT('h02)
	) name3288 (
		\u4_u1_dma_out_cnt_reg[9]/P0001 ,
		_w5036_,
		_w5037_,
		_w5038_
	);
	LUT2 #(
		.INIT('h4)
	) name3289 (
		_w5035_,
		_w5038_,
		_w5039_
	);
	LUT2 #(
		.INIT('h1)
	) name3290 (
		\u4_u1_dma_out_cnt_reg[9]/P0001 ,
		\u4_u1_r5_reg/NET0131 ,
		_w5040_
	);
	LUT4 #(
		.INIT('hec00)
	) name3291 (
		_w4737_,
		_w5031_,
		_w5032_,
		_w5040_,
		_w5041_
	);
	LUT3 #(
		.INIT('h54)
	) name3292 (
		\u4_u1_dma_out_cnt_reg[9]/P0001 ,
		_w5036_,
		_w5037_,
		_w5042_
	);
	LUT2 #(
		.INIT('h4)
	) name3293 (
		\u4_u1_dma_out_cnt_reg[9]/P0001 ,
		\u4_u1_r5_reg/NET0131 ,
		_w5043_
	);
	LUT4 #(
		.INIT('h7f00)
	) name3294 (
		_w4711_,
		_w4713_,
		_w5034_,
		_w5043_,
		_w5044_
	);
	LUT3 #(
		.INIT('h02)
	) name3295 (
		\u4_u1_csr1_reg[0]/P0001 ,
		_w5042_,
		_w5044_,
		_w5045_
	);
	LUT4 #(
		.INIT('h0b00)
	) name3296 (
		_w5033_,
		_w5039_,
		_w5041_,
		_w5045_,
		_w5046_
	);
	LUT2 #(
		.INIT('h1)
	) name3297 (
		\u4_u2_dma_out_cnt_reg[4]/P0001 ,
		\u4_u2_dma_out_cnt_reg[5]/P0001 ,
		_w5047_
	);
	LUT4 #(
		.INIT('h0001)
	) name3298 (
		\u4_u2_dma_out_cnt_reg[6]/P0001 ,
		\u4_u2_dma_out_cnt_reg[7]/P0001 ,
		\u4_u2_dma_out_cnt_reg[8]/P0001 ,
		\u4_u2_dma_out_cnt_reg[9]/P0001 ,
		_w5048_
	);
	LUT2 #(
		.INIT('h4)
	) name3299 (
		\u4_u2_dma_out_cnt_reg[10]/P0001 ,
		\u4_u2_r5_reg/NET0131 ,
		_w5049_
	);
	LUT4 #(
		.INIT('h8000)
	) name3300 (
		_w4744_,
		_w5047_,
		_w5048_,
		_w5049_,
		_w5050_
	);
	LUT4 #(
		.INIT('h4000)
	) name3301 (
		\u4_u2_dma_out_cnt_reg[10]/P0001 ,
		_w4744_,
		_w5047_,
		_w5048_,
		_w5051_
	);
	LUT2 #(
		.INIT('h8)
	) name3302 (
		\u4_u2_dma_out_cnt_reg[10]/P0001 ,
		\u4_u2_ep_match_r_reg/P0001 ,
		_w5052_
	);
	LUT2 #(
		.INIT('h4)
	) name3303 (
		_w4482_,
		_w5052_,
		_w5053_
	);
	LUT4 #(
		.INIT('h0233)
	) name3304 (
		\u4_u2_r5_reg/NET0131 ,
		_w5050_,
		_w5051_,
		_w5053_,
		_w5054_
	);
	LUT3 #(
		.INIT('he0)
	) name3305 (
		\u4_u2_csr0_reg[10]/P0001 ,
		\u4_u2_dma_out_cnt_reg[8]/P0001 ,
		\u4_u2_dma_out_cnt_reg[9]/P0001 ,
		_w5055_
	);
	LUT2 #(
		.INIT('h4)
	) name3306 (
		_w4754_,
		_w5055_,
		_w5056_
	);
	LUT3 #(
		.INIT('h80)
	) name3307 (
		\u4_u2_csr0_reg[10]/P0001 ,
		\u4_u2_dma_out_cnt_reg[8]/P0001 ,
		\u4_u2_dma_out_cnt_reg[9]/P0001 ,
		_w5057_
	);
	LUT2 #(
		.INIT('h1)
	) name3308 (
		_w5050_,
		_w5057_,
		_w5058_
	);
	LUT4 #(
		.INIT('h8f00)
	) name3309 (
		_w4767_,
		_w4768_,
		_w5056_,
		_w5058_,
		_w5059_
	);
	LUT4 #(
		.INIT('h8882)
	) name3310 (
		\u4_u2_csr1_reg[0]/P0001 ,
		\u4_u2_dma_out_cnt_reg[11]/P0001 ,
		_w5054_,
		_w5059_,
		_w5060_
	);
	LUT4 #(
		.INIT('hfca8)
	) name3311 (
		\u4_u2_csr0_reg[10]/P0001 ,
		\u4_u2_csr0_reg[9]/P0001 ,
		\u4_u2_dma_out_cnt_reg[7]/P0001 ,
		\u4_u2_dma_out_cnt_reg[8]/P0001 ,
		_w5061_
	);
	LUT3 #(
		.INIT('h07)
	) name3312 (
		\u4_u2_csr0_reg[10]/P0001 ,
		\u4_u2_dma_out_cnt_reg[8]/P0001 ,
		\u4_u2_r5_reg/NET0131 ,
		_w5062_
	);
	LUT4 #(
		.INIT('h8f00)
	) name3313 (
		_w4767_,
		_w4768_,
		_w5061_,
		_w5062_,
		_w5063_
	);
	LUT2 #(
		.INIT('h4)
	) name3314 (
		\u4_u2_r5_reg/NET0131 ,
		_w4610_,
		_w5064_
	);
	LUT3 #(
		.INIT('h80)
	) name3315 (
		_w4742_,
		_w4744_,
		_w4745_,
		_w5065_
	);
	LUT3 #(
		.INIT('ha8)
	) name3316 (
		\u4_u2_dma_out_cnt_reg[9]/P0001 ,
		_w5064_,
		_w5065_,
		_w5066_
	);
	LUT4 #(
		.INIT('h0007)
	) name3317 (
		\u4_u2_csr0_reg[10]/P0001 ,
		\u4_u2_dma_out_cnt_reg[8]/P0001 ,
		\u4_u2_dma_out_cnt_reg[9]/P0001 ,
		\u4_u2_r5_reg/NET0131 ,
		_w5067_
	);
	LUT4 #(
		.INIT('h8f00)
	) name3318 (
		_w4767_,
		_w4768_,
		_w5061_,
		_w5067_,
		_w5068_
	);
	LUT4 #(
		.INIT('haaa8)
	) name3319 (
		\u4_u2_csr1_reg[0]/P0001 ,
		\u4_u2_dma_out_cnt_reg[9]/P0001 ,
		_w5064_,
		_w5065_,
		_w5069_
	);
	LUT4 #(
		.INIT('h0b00)
	) name3320 (
		_w5063_,
		_w5066_,
		_w5068_,
		_w5069_,
		_w5070_
	);
	LUT2 #(
		.INIT('h2)
	) name3321 (
		_w4389_,
		_w4560_,
		_w5071_
	);
	LUT3 #(
		.INIT('h08)
	) name3322 (
		_w4387_,
		_w4394_,
		_w4395_,
		_w5072_
	);
	LUT4 #(
		.INIT('h0b00)
	) name3323 (
		\u4_u3_csr0_reg[10]/P0001 ,
		\u4_u3_dma_in_cnt_reg[8]/P0001 ,
		\u4_u3_dma_in_cnt_reg[9]/P0001 ,
		\u4_u3_ep_match_r_reg/P0001 ,
		_w5073_
	);
	LUT2 #(
		.INIT('h4)
	) name3324 (
		_w4402_,
		_w5073_,
		_w5074_
	);
	LUT4 #(
		.INIT('h4055)
	) name3325 (
		\u4_u3_r5_reg/NET0131 ,
		_w5071_,
		_w5072_,
		_w5074_,
		_w5075_
	);
	LUT3 #(
		.INIT('h20)
	) name3326 (
		_w4387_,
		_w4395_,
		_w4559_,
		_w5076_
	);
	LUT4 #(
		.INIT('hf531)
	) name3327 (
		\u4_u3_csr0_reg[7]/P0001 ,
		\u4_u3_csr0_reg[8]/P0001 ,
		\u4_u3_dma_in_cnt_reg[5]/P0001 ,
		\u4_u3_dma_in_cnt_reg[6]/P0001 ,
		_w5077_
	);
	LUT3 #(
		.INIT('h8a)
	) name3328 (
		_w4562_,
		_w4563_,
		_w5077_,
		_w5078_
	);
	LUT2 #(
		.INIT('h4)
	) name3329 (
		\u4_u3_r5_reg/NET0131 ,
		_w4394_,
		_w5079_
	);
	LUT2 #(
		.INIT('h2)
	) name3330 (
		\u4_u3_dma_in_cnt_reg[10]/P0001 ,
		\u4_u3_r5_reg/NET0131 ,
		_w5080_
	);
	LUT4 #(
		.INIT('h8000)
	) name3331 (
		\u4_u3_dma_in_cnt_reg[10]/P0001 ,
		\u4_u3_dma_in_cnt_reg[7]/P0001 ,
		\u4_u3_dma_in_cnt_reg[8]/P0001 ,
		\u4_u3_dma_in_cnt_reg[9]/P0001 ,
		_w5081_
	);
	LUT4 #(
		.INIT('h070f)
	) name3332 (
		_w4398_,
		_w4399_,
		_w5080_,
		_w5081_,
		_w5082_
	);
	LUT4 #(
		.INIT('h004f)
	) name3333 (
		_w5076_,
		_w5078_,
		_w5079_,
		_w5082_,
		_w5083_
	);
	LUT2 #(
		.INIT('h8)
	) name3334 (
		\u4_u3_csr1_reg[0]/P0001 ,
		\u4_u3_dma_in_cnt_reg[10]/P0001 ,
		_w5084_
	);
	LUT2 #(
		.INIT('h2)
	) name3335 (
		\u4_u3_csr1_reg[0]/P0001 ,
		\u4_u3_r5_reg/NET0131 ,
		_w5085_
	);
	LUT4 #(
		.INIT('h8000)
	) name3336 (
		\u4_u3_csr1_reg[0]/P0001 ,
		\u4_u3_dma_in_cnt_reg[7]/P0001 ,
		\u4_u3_dma_in_cnt_reg[8]/P0001 ,
		\u4_u3_dma_in_cnt_reg[9]/P0001 ,
		_w5086_
	);
	LUT4 #(
		.INIT('h070f)
	) name3337 (
		_w4398_,
		_w4399_,
		_w5085_,
		_w5086_,
		_w5087_
	);
	LUT4 #(
		.INIT('h004f)
	) name3338 (
		_w5076_,
		_w5078_,
		_w5079_,
		_w5087_,
		_w5088_
	);
	LUT4 #(
		.INIT('hb1b0)
	) name3339 (
		_w5075_,
		_w5083_,
		_w5084_,
		_w5088_,
		_w5089_
	);
	LUT2 #(
		.INIT('h2)
	) name3340 (
		_w4421_,
		_w4583_,
		_w5090_
	);
	LUT3 #(
		.INIT('h08)
	) name3341 (
		_w4419_,
		_w4426_,
		_w4427_,
		_w5091_
	);
	LUT4 #(
		.INIT('h0b00)
	) name3342 (
		\u4_u0_csr0_reg[10]/P0001 ,
		\u4_u0_dma_in_cnt_reg[8]/P0001 ,
		\u4_u0_dma_in_cnt_reg[9]/P0001 ,
		\u4_u0_ep_match_r_reg/P0001 ,
		_w5092_
	);
	LUT2 #(
		.INIT('h4)
	) name3343 (
		_w4434_,
		_w5092_,
		_w5093_
	);
	LUT4 #(
		.INIT('h4055)
	) name3344 (
		\u4_u0_r5_reg/NET0131 ,
		_w5090_,
		_w5091_,
		_w5093_,
		_w5094_
	);
	LUT3 #(
		.INIT('h20)
	) name3345 (
		_w4419_,
		_w4427_,
		_w4582_,
		_w5095_
	);
	LUT4 #(
		.INIT('hf531)
	) name3346 (
		\u4_u0_csr0_reg[7]/P0001 ,
		\u4_u0_csr0_reg[8]/P0001 ,
		\u4_u0_dma_in_cnt_reg[5]/P0001 ,
		\u4_u0_dma_in_cnt_reg[6]/P0001 ,
		_w5096_
	);
	LUT3 #(
		.INIT('h8a)
	) name3347 (
		_w4585_,
		_w4586_,
		_w5096_,
		_w5097_
	);
	LUT2 #(
		.INIT('h4)
	) name3348 (
		\u4_u0_r5_reg/NET0131 ,
		_w4426_,
		_w5098_
	);
	LUT2 #(
		.INIT('h2)
	) name3349 (
		\u4_u0_dma_in_cnt_reg[10]/P0001 ,
		\u4_u0_r5_reg/NET0131 ,
		_w5099_
	);
	LUT4 #(
		.INIT('h8000)
	) name3350 (
		\u4_u0_dma_in_cnt_reg[10]/P0001 ,
		\u4_u0_dma_in_cnt_reg[7]/P0001 ,
		\u4_u0_dma_in_cnt_reg[8]/P0001 ,
		\u4_u0_dma_in_cnt_reg[9]/P0001 ,
		_w5100_
	);
	LUT4 #(
		.INIT('h070f)
	) name3351 (
		_w4430_,
		_w4431_,
		_w5099_,
		_w5100_,
		_w5101_
	);
	LUT4 #(
		.INIT('h004f)
	) name3352 (
		_w5095_,
		_w5097_,
		_w5098_,
		_w5101_,
		_w5102_
	);
	LUT2 #(
		.INIT('h8)
	) name3353 (
		\u4_u0_csr1_reg[0]/P0001 ,
		\u4_u0_dma_in_cnt_reg[10]/P0001 ,
		_w5103_
	);
	LUT4 #(
		.INIT('h8000)
	) name3354 (
		\u4_u0_csr1_reg[0]/P0001 ,
		\u4_u0_dma_in_cnt_reg[7]/P0001 ,
		\u4_u0_dma_in_cnt_reg[8]/P0001 ,
		\u4_u0_dma_in_cnt_reg[9]/P0001 ,
		_w5104_
	);
	LUT4 #(
		.INIT('h070f)
	) name3355 (
		_w4430_,
		_w4431_,
		_w4578_,
		_w5104_,
		_w5105_
	);
	LUT4 #(
		.INIT('h004f)
	) name3356 (
		_w5095_,
		_w5097_,
		_w5098_,
		_w5105_,
		_w5106_
	);
	LUT4 #(
		.INIT('hb1b0)
	) name3357 (
		_w5094_,
		_w5102_,
		_w5103_,
		_w5106_,
		_w5107_
	);
	LUT3 #(
		.INIT('h80)
	) name3358 (
		_w4447_,
		_w4448_,
		_w4925_,
		_w5108_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name3359 (
		\u4_u1_r5_reg/NET0131 ,
		_w4447_,
		_w4448_,
		_w4925_,
		_w5109_
	);
	LUT3 #(
		.INIT('h0b)
	) name3360 (
		\u4_u1_csr0_reg[10]/P0001 ,
		\u4_u1_dma_in_cnt_reg[8]/P0001 ,
		\u4_u1_dma_in_cnt_reg[9]/P0001 ,
		_w5110_
	);
	LUT3 #(
		.INIT('h10)
	) name3361 (
		_w5036_,
		_w5037_,
		_w5110_,
		_w5111_
	);
	LUT3 #(
		.INIT('h10)
	) name3362 (
		_w4473_,
		_w5109_,
		_w5111_,
		_w5112_
	);
	LUT3 #(
		.INIT('h20)
	) name3363 (
		_w4606_,
		_w5109_,
		_w5111_,
		_w5113_
	);
	LUT3 #(
		.INIT('h0c)
	) name3364 (
		\u4_u1_ep_match_r_reg/P0001 ,
		\u4_u1_r5_reg/NET0131 ,
		_w5037_,
		_w5114_
	);
	LUT2 #(
		.INIT('h8)
	) name3365 (
		_w5108_,
		_w5114_,
		_w5115_
	);
	LUT2 #(
		.INIT('h8)
	) name3366 (
		\u4_u1_csr1_reg[0]/P0001 ,
		\u4_u1_dma_in_cnt_reg[10]/P0001 ,
		_w5116_
	);
	LUT3 #(
		.INIT('h70)
	) name3367 (
		_w5108_,
		_w5114_,
		_w5116_,
		_w5117_
	);
	LUT4 #(
		.INIT('h2300)
	) name3368 (
		_w4605_,
		_w5112_,
		_w5113_,
		_w5117_,
		_w5118_
	);
	LUT4 #(
		.INIT('h0023)
	) name3369 (
		_w4605_,
		_w5112_,
		_w5113_,
		_w5115_,
		_w5119_
	);
	LUT2 #(
		.INIT('h2)
	) name3370 (
		\u4_u1_csr1_reg[0]/P0001 ,
		\u4_u1_dma_in_cnt_reg[10]/P0001 ,
		_w5120_
	);
	LUT3 #(
		.INIT('hba)
	) name3371 (
		_w5118_,
		_w5119_,
		_w5120_,
		_w5121_
	);
	LUT4 #(
		.INIT('h8000)
	) name3372 (
		\u4_u2_dma_in_cnt_reg[7]/P0001 ,
		\u4_u2_dma_in_cnt_reg[8]/P0001 ,
		\u4_u2_dma_in_cnt_reg[9]/P0001 ,
		\u4_u2_r5_reg/NET0131 ,
		_w5122_
	);
	LUT4 #(
		.INIT('h070f)
	) name3373 (
		_w4504_,
		_w4505_,
		_w4509_,
		_w5122_,
		_w5123_
	);
	LUT2 #(
		.INIT('h2)
	) name3374 (
		\u4_u2_dma_in_cnt_reg[10]/P0001 ,
		_w5123_,
		_w5124_
	);
	LUT2 #(
		.INIT('h1)
	) name3375 (
		\u4_u2_dma_in_cnt_reg[10]/P0001 ,
		\u4_u2_r5_reg/NET0131 ,
		_w5125_
	);
	LUT4 #(
		.INIT('hea00)
	) name3376 (
		_w4486_,
		_w4499_,
		_w4501_,
		_w5125_,
		_w5126_
	);
	LUT3 #(
		.INIT('h8a)
	) name3377 (
		\u4_u2_csr1_reg[0]/P0001 ,
		\u4_u2_dma_in_cnt_reg[10]/P0001 ,
		_w5123_,
		_w5127_
	);
	LUT4 #(
		.INIT('h0b00)
	) name3378 (
		_w4502_,
		_w5124_,
		_w5126_,
		_w5127_,
		_w5128_
	);
	LUT4 #(
		.INIT('h4000)
	) name3379 (
		\u0_u0_me_cnt_100_ms_reg/P0001 ,
		\u0_u0_me_cnt_reg[0]/P0001 ,
		\u0_u0_me_cnt_reg[1]/P0001 ,
		\u0_u0_me_ps2_0_5_ms_reg/P0001 ,
		_w5129_
	);
	LUT4 #(
		.INIT('hb4f0)
	) name3380 (
		\u0_u0_me_cnt_100_ms_reg/P0001 ,
		\u0_u0_me_cnt_reg[0]/P0001 ,
		\u0_u0_me_cnt_reg[1]/P0001 ,
		\u0_u0_me_ps2_0_5_ms_reg/P0001 ,
		_w5130_
	);
	LUT2 #(
		.INIT('h8)
	) name3381 (
		_w4358_,
		_w5130_,
		_w5131_
	);
	LUT2 #(
		.INIT('h4)
	) name3382 (
		_w4353_,
		_w5131_,
		_w5132_
	);
	LUT2 #(
		.INIT('h4)
	) name3383 (
		_w4350_,
		_w5132_,
		_w5133_
	);
	LUT3 #(
		.INIT('h14)
	) name3384 (
		\u1_clr_sof_time_reg/P0001 ,
		\u1_hms_clk_reg/P0001 ,
		\u1_sof_time_reg[0]/P0001 ,
		_w5134_
	);
	LUT3 #(
		.INIT('h9c)
	) name3385 (
		\u0_u0_me_cnt_100_ms_reg/P0001 ,
		\u0_u0_me_cnt_reg[0]/P0001 ,
		\u0_u0_me_ps2_0_5_ms_reg/P0001 ,
		_w5135_
	);
	LUT2 #(
		.INIT('h8)
	) name3386 (
		_w4626_,
		_w5135_,
		_w5136_
	);
	LUT2 #(
		.INIT('h4)
	) name3387 (
		_w4350_,
		_w5136_,
		_w5137_
	);
	LUT2 #(
		.INIT('h6)
	) name3388 (
		\u0_u0_me_cnt_reg[2]/P0001 ,
		_w5129_,
		_w5138_
	);
	LUT2 #(
		.INIT('h8)
	) name3389 (
		_w4626_,
		_w5138_,
		_w5139_
	);
	LUT2 #(
		.INIT('h4)
	) name3390 (
		_w4350_,
		_w5139_,
		_w5140_
	);
	LUT3 #(
		.INIT('h6c)
	) name3391 (
		\u0_u0_me_cnt_reg[2]/P0001 ,
		\u0_u0_me_cnt_reg[3]/P0001 ,
		_w5129_,
		_w5141_
	);
	LUT2 #(
		.INIT('h8)
	) name3392 (
		_w4626_,
		_w5141_,
		_w5142_
	);
	LUT2 #(
		.INIT('h4)
	) name3393 (
		_w4350_,
		_w5142_,
		_w5143_
	);
	LUT3 #(
		.INIT('h80)
	) name3394 (
		\u0_u0_me_cnt_reg[2]/P0001 ,
		\u0_u0_me_cnt_reg[3]/P0001 ,
		\u0_u0_me_cnt_reg[4]/P0001 ,
		_w5144_
	);
	LUT4 #(
		.INIT('h78f0)
	) name3395 (
		\u0_u0_me_cnt_reg[2]/P0001 ,
		\u0_u0_me_cnt_reg[3]/P0001 ,
		\u0_u0_me_cnt_reg[4]/P0001 ,
		_w5129_,
		_w5145_
	);
	LUT2 #(
		.INIT('h8)
	) name3396 (
		_w4358_,
		_w5145_,
		_w5146_
	);
	LUT2 #(
		.INIT('h4)
	) name3397 (
		_w4353_,
		_w5146_,
		_w5147_
	);
	LUT2 #(
		.INIT('h4)
	) name3398 (
		_w4350_,
		_w5147_,
		_w5148_
	);
	LUT3 #(
		.INIT('h6a)
	) name3399 (
		\u0_u0_me_cnt_reg[5]/P0001 ,
		_w5129_,
		_w5144_,
		_w5149_
	);
	LUT2 #(
		.INIT('h8)
	) name3400 (
		_w4626_,
		_w5149_,
		_w5150_
	);
	LUT2 #(
		.INIT('h4)
	) name3401 (
		_w4350_,
		_w5150_,
		_w5151_
	);
	LUT2 #(
		.INIT('h8)
	) name3402 (
		\u0_u0_me_cnt_reg[5]/P0001 ,
		\u0_u0_me_cnt_reg[6]/P0001 ,
		_w5152_
	);
	LUT3 #(
		.INIT('h80)
	) name3403 (
		_w5129_,
		_w5144_,
		_w5152_,
		_w5153_
	);
	LUT2 #(
		.INIT('h2)
	) name3404 (
		_w4358_,
		_w5153_,
		_w5154_
	);
	LUT4 #(
		.INIT('h1333)
	) name3405 (
		\u0_u0_me_cnt_reg[5]/P0001 ,
		\u0_u0_me_cnt_reg[6]/P0001 ,
		_w5129_,
		_w5144_,
		_w5155_
	);
	LUT3 #(
		.INIT('h04)
	) name3406 (
		_w4353_,
		_w5154_,
		_w5155_,
		_w5156_
	);
	LUT2 #(
		.INIT('h4)
	) name3407 (
		_w4350_,
		_w5156_,
		_w5157_
	);
	LUT4 #(
		.INIT('h9555)
	) name3408 (
		\u0_u0_me_cnt_reg[7]/P0001 ,
		_w5129_,
		_w5144_,
		_w5152_,
		_w5158_
	);
	LUT2 #(
		.INIT('h2)
	) name3409 (
		_w4358_,
		_w5158_,
		_w5159_
	);
	LUT2 #(
		.INIT('h4)
	) name3410 (
		_w4353_,
		_w5159_,
		_w5160_
	);
	LUT2 #(
		.INIT('h4)
	) name3411 (
		_w4350_,
		_w5160_,
		_w5161_
	);
	LUT3 #(
		.INIT('h80)
	) name3412 (
		\u4_u2_dma_in_buf_sz1_reg/P0001 ,
		_w3762_,
		_w3763_,
		_w5162_
	);
	LUT2 #(
		.INIT('h8)
	) name3413 (
		_w3761_,
		_w5162_,
		_w5163_
	);
	LUT3 #(
		.INIT('h80)
	) name3414 (
		\u4_u0_dma_in_buf_sz1_reg/P0001 ,
		_w3755_,
		_w3756_,
		_w5164_
	);
	LUT3 #(
		.INIT('h07)
	) name3415 (
		\u4_u1_dma_in_buf_sz1_reg/P0001 ,
		_w3768_,
		_w5164_,
		_w5165_
	);
	LUT3 #(
		.INIT('h80)
	) name3416 (
		\u4_dma_in_buf_sz1_reg/P0001 ,
		_w3761_,
		_w3775_,
		_w5166_
	);
	LUT3 #(
		.INIT('h80)
	) name3417 (
		\u4_u3_dma_in_buf_sz1_reg/P0001 ,
		_w3761_,
		_w3773_,
		_w5167_
	);
	LUT4 #(
		.INIT('hfffb)
	) name3418 (
		_w5163_,
		_w5165_,
		_w5166_,
		_w5167_,
		_w5168_
	);
	LUT3 #(
		.INIT('h80)
	) name3419 (
		\u1_sof_time_reg[1]/P0001 ,
		\u1_sof_time_reg[2]/P0001 ,
		\u1_sof_time_reg[9]/P0001 ,
		_w5169_
	);
	LUT4 #(
		.INIT('h8000)
	) name3420 (
		_w4365_,
		_w4366_,
		_w4367_,
		_w5169_,
		_w5170_
	);
	LUT4 #(
		.INIT('h0504)
	) name3421 (
		\u1_clr_sof_time_reg/P0001 ,
		\u1_sof_time_reg[10]/P0001 ,
		_w4370_,
		_w5170_,
		_w5171_
	);
	LUT4 #(
		.INIT('h1540)
	) name3422 (
		\u1_clr_sof_time_reg/P0001 ,
		\u1_hms_clk_reg/P0001 ,
		\u1_sof_time_reg[0]/P0001 ,
		\u1_sof_time_reg[1]/P0001 ,
		_w5172_
	);
	LUT4 #(
		.INIT('h007f)
	) name3423 (
		\u1_hms_clk_reg/P0001 ,
		\u1_sof_time_reg[0]/P0001 ,
		\u1_sof_time_reg[1]/P0001 ,
		\u1_sof_time_reg[2]/P0001 ,
		_w5173_
	);
	LUT3 #(
		.INIT('h01)
	) name3424 (
		\u1_clr_sof_time_reg/P0001 ,
		_w4845_,
		_w5173_,
		_w5174_
	);
	LUT3 #(
		.INIT('h14)
	) name3425 (
		\u1_clr_sof_time_reg/P0001 ,
		\u1_sof_time_reg[3]/P0001 ,
		_w4845_,
		_w5175_
	);
	LUT2 #(
		.INIT('h8)
	) name3426 (
		\u1_sof_time_reg[3]/P0001 ,
		\u1_sof_time_reg[4]/P0001 ,
		_w5176_
	);
	LUT4 #(
		.INIT('h1450)
	) name3427 (
		\u1_clr_sof_time_reg/P0001 ,
		\u1_sof_time_reg[3]/P0001 ,
		\u1_sof_time_reg[4]/P0001 ,
		_w4845_,
		_w5177_
	);
	LUT3 #(
		.INIT('h15)
	) name3428 (
		\u1_sof_time_reg[5]/P0001 ,
		_w4845_,
		_w5176_,
		_w5178_
	);
	LUT3 #(
		.INIT('h15)
	) name3429 (
		\u1_clr_sof_time_reg/P0001 ,
		_w4367_,
		_w4845_,
		_w5179_
	);
	LUT2 #(
		.INIT('h4)
	) name3430 (
		_w5178_,
		_w5179_,
		_w5180_
	);
	LUT4 #(
		.INIT('h1444)
	) name3431 (
		\u1_clr_sof_time_reg/P0001 ,
		\u1_sof_time_reg[6]/P0001 ,
		_w4367_,
		_w4845_,
		_w5181_
	);
	LUT4 #(
		.INIT('h1555)
	) name3432 (
		\u1_sof_time_reg[8]/P0001 ,
		_w4367_,
		_w4845_,
		_w4847_,
		_w5182_
	);
	LUT4 #(
		.INIT('h8000)
	) name3433 (
		_w4365_,
		_w4366_,
		_w4367_,
		_w4368_,
		_w5183_
	);
	LUT3 #(
		.INIT('h01)
	) name3434 (
		\u1_clr_sof_time_reg/P0001 ,
		_w5182_,
		_w5183_,
		_w5184_
	);
	LUT2 #(
		.INIT('h4)
	) name3435 (
		\u1_clr_sof_time_reg/P0001 ,
		\u1_sof_time_reg[9]/P0001 ,
		_w5185_
	);
	LUT2 #(
		.INIT('h1)
	) name3436 (
		\u1_clr_sof_time_reg/P0001 ,
		\u1_sof_time_reg[9]/P0001 ,
		_w5186_
	);
	LUT4 #(
		.INIT('h8000)
	) name3437 (
		_w4366_,
		_w4367_,
		_w4845_,
		_w5186_,
		_w5187_
	);
	LUT3 #(
		.INIT('hf4)
	) name3438 (
		_w5183_,
		_w5185_,
		_w5187_,
		_w5188_
	);
	LUT4 #(
		.INIT('h0a08)
	) name3439 (
		rst_i_pad,
		\u4_crc5_err_r_reg/P0001 ,
		\u4_int_src_re_reg/P0001 ,
		\u4_int_srcb_reg[0]/P0001 ,
		_w5189_
	);
	LUT2 #(
		.INIT('h4)
	) name3440 (
		\u1_u2_sizu_c_reg[10]/P0001 ,
		\u4_csr_reg[10]/P0001 ,
		_w5190_
	);
	LUT4 #(
		.INIT('hf531)
	) name3441 (
		\u1_u2_sizu_c_reg[10]/P0001 ,
		\u1_u2_sizu_c_reg[9]/P0001 ,
		\u4_csr_reg[10]/P0001 ,
		\u4_csr_reg[9]/NET0131 ,
		_w5191_
	);
	LUT2 #(
		.INIT('h2)
	) name3442 (
		\u1_u2_sizu_c_reg[8]/NET0131 ,
		\u4_csr_reg[8]/P0001 ,
		_w5192_
	);
	LUT2 #(
		.INIT('h2)
	) name3443 (
		\u1_u2_sizu_c_reg[7]/P0001 ,
		\u4_csr_reg[7]/P0001 ,
		_w5193_
	);
	LUT4 #(
		.INIT('hf531)
	) name3444 (
		\u1_u2_sizu_c_reg[7]/P0001 ,
		\u1_u2_sizu_c_reg[8]/NET0131 ,
		\u4_csr_reg[7]/P0001 ,
		\u4_csr_reg[8]/P0001 ,
		_w5194_
	);
	LUT4 #(
		.INIT('h8caf)
	) name3445 (
		\u1_u2_sizu_c_reg[8]/NET0131 ,
		\u1_u2_sizu_c_reg[9]/P0001 ,
		\u4_csr_reg[8]/P0001 ,
		\u4_csr_reg[9]/NET0131 ,
		_w5195_
	);
	LUT4 #(
		.INIT('h1511)
	) name3446 (
		_w5190_,
		_w5191_,
		_w5194_,
		_w5195_,
		_w5196_
	);
	LUT4 #(
		.INIT('h8caf)
	) name3447 (
		\u1_u2_sizu_c_reg[3]/P0001 ,
		\u1_u2_sizu_c_reg[4]/P0001 ,
		\u4_csr_reg[3]/P0001 ,
		\u4_csr_reg[4]/NET0131 ,
		_w5197_
	);
	LUT4 #(
		.INIT('hf531)
	) name3448 (
		\u1_u2_sizu_c_reg[5]/P0001 ,
		\u1_u2_sizu_c_reg[6]/P0001 ,
		\u4_csr_reg[5]/NET0131 ,
		\u4_csr_reg[6]/NET0131 ,
		_w5198_
	);
	LUT2 #(
		.INIT('h2)
	) name3449 (
		\u1_u2_sizu_c_reg[4]/P0001 ,
		\u4_csr_reg[4]/NET0131 ,
		_w5199_
	);
	LUT3 #(
		.INIT('h04)
	) name3450 (
		_w5197_,
		_w5198_,
		_w5199_,
		_w5200_
	);
	LUT4 #(
		.INIT('h8caf)
	) name3451 (
		\u1_u2_sizu_c_reg[7]/P0001 ,
		\u1_u2_sizu_c_reg[8]/NET0131 ,
		\u4_csr_reg[7]/P0001 ,
		\u4_csr_reg[8]/P0001 ,
		_w5201_
	);
	LUT3 #(
		.INIT('h02)
	) name3452 (
		_w5191_,
		_w5192_,
		_w5201_,
		_w5202_
	);
	LUT4 #(
		.INIT('h8caf)
	) name3453 (
		\u1_u2_sizu_c_reg[10]/P0001 ,
		\u1_u2_sizu_c_reg[9]/P0001 ,
		\u4_csr_reg[10]/P0001 ,
		\u4_csr_reg[9]/NET0131 ,
		_w5203_
	);
	LUT4 #(
		.INIT('h7150)
	) name3454 (
		\u1_u2_sizu_c_reg[10]/P0001 ,
		\u1_u2_sizu_c_reg[9]/P0001 ,
		\u4_csr_reg[10]/P0001 ,
		\u4_csr_reg[9]/NET0131 ,
		_w5204_
	);
	LUT2 #(
		.INIT('h4)
	) name3455 (
		\u1_u2_sizu_c_reg[6]/P0001 ,
		\u4_csr_reg[6]/NET0131 ,
		_w5205_
	);
	LUT4 #(
		.INIT('h8caf)
	) name3456 (
		\u1_u2_sizu_c_reg[5]/P0001 ,
		\u1_u2_sizu_c_reg[6]/P0001 ,
		\u4_csr_reg[5]/NET0131 ,
		\u4_csr_reg[6]/NET0131 ,
		_w5206_
	);
	LUT4 #(
		.INIT('h7310)
	) name3457 (
		\u1_u2_sizu_c_reg[5]/P0001 ,
		\u1_u2_sizu_c_reg[6]/P0001 ,
		\u4_csr_reg[5]/NET0131 ,
		\u4_csr_reg[6]/NET0131 ,
		_w5207_
	);
	LUT2 #(
		.INIT('h1)
	) name3458 (
		_w5204_,
		_w5207_,
		_w5208_
	);
	LUT4 #(
		.INIT('h5455)
	) name3459 (
		_w5196_,
		_w5200_,
		_w5202_,
		_w5208_,
		_w5209_
	);
	LUT4 #(
		.INIT('h00fd)
	) name3460 (
		_w5191_,
		_w5192_,
		_w5201_,
		_w5204_,
		_w5210_
	);
	LUT4 #(
		.INIT('hf531)
	) name3461 (
		\u1_u2_sizu_c_reg[3]/P0001 ,
		\u1_u2_sizu_c_reg[4]/P0001 ,
		\u4_csr_reg[3]/P0001 ,
		\u4_csr_reg[4]/NET0131 ,
		_w5211_
	);
	LUT4 #(
		.INIT('h8caf)
	) name3462 (
		\u1_u2_sizu_c_reg[4]/P0001 ,
		\u1_u2_sizu_c_reg[5]/P0001 ,
		\u4_csr_reg[4]/NET0131 ,
		\u4_csr_reg[5]/NET0131 ,
		_w5212_
	);
	LUT4 #(
		.INIT('h1311)
	) name3463 (
		_w5198_,
		_w5205_,
		_w5211_,
		_w5212_,
		_w5213_
	);
	LUT2 #(
		.INIT('h4)
	) name3464 (
		\u1_u2_sizu_c_reg[2]/P0001 ,
		\u4_csr_reg[2]/NET0131 ,
		_w5214_
	);
	LUT4 #(
		.INIT('h8caf)
	) name3465 (
		\u1_u2_sizu_c_reg[0]/P0001 ,
		\u1_u2_sizu_c_reg[1]/P0001 ,
		\u4_csr_reg[0]/P0001 ,
		\u4_csr_reg[1]/P0001 ,
		_w5215_
	);
	LUT4 #(
		.INIT('hf531)
	) name3466 (
		\u1_u2_sizu_c_reg[1]/P0001 ,
		\u1_u2_sizu_c_reg[2]/P0001 ,
		\u4_csr_reg[1]/P0001 ,
		\u4_csr_reg[2]/NET0131 ,
		_w5216_
	);
	LUT4 #(
		.INIT('h4544)
	) name3467 (
		\u4_csr_reg[16]/P0001 ,
		_w5214_,
		_w5215_,
		_w5216_,
		_w5217_
	);
	LUT4 #(
		.INIT('h3700)
	) name3468 (
		_w5196_,
		_w5210_,
		_w5213_,
		_w5217_,
		_w5218_
	);
	LUT3 #(
		.INIT('hf4)
	) name3469 (
		\u4_csr_reg[16]/P0001 ,
		_w5209_,
		_w5218_,
		_w5219_
	);
	LUT3 #(
		.INIT('hac)
	) name3470 (
		\u1_u2_sizu_c_reg[2]/P0001 ,
		\u1_u3_new_size_reg[2]/P0001 ,
		\u1_u3_out_to_small_r_reg/P0001 ,
		_w5220_
	);
	LUT3 #(
		.INIT('hac)
	) name3471 (
		\u1_u2_sizu_c_reg[3]/P0001 ,
		\u1_u3_new_size_reg[3]/P0001 ,
		\u1_u3_out_to_small_r_reg/P0001 ,
		_w5221_
	);
	LUT3 #(
		.INIT('h59)
	) name3472 (
		\u1_u3_adr_reg[4]/P0001 ,
		_w2803_,
		_w2805_,
		_w5222_
	);
	LUT4 #(
		.INIT('h0bf4)
	) name3473 (
		_w4073_,
		_w4076_,
		_w4078_,
		_w5222_,
		_w5223_
	);
	LUT3 #(
		.INIT('h59)
	) name3474 (
		\u1_u3_adr_reg[5]/P0001 ,
		_w2820_,
		_w2822_,
		_w5224_
	);
	LUT2 #(
		.INIT('h1)
	) name3475 (
		_w4068_,
		_w5224_,
		_w5225_
	);
	LUT4 #(
		.INIT('h4f00)
	) name3476 (
		_w4073_,
		_w4076_,
		_w4079_,
		_w5225_,
		_w5226_
	);
	LUT2 #(
		.INIT('h8)
	) name3477 (
		_w4068_,
		_w5224_,
		_w5227_
	);
	LUT3 #(
		.INIT('h10)
	) name3478 (
		_w4077_,
		_w4078_,
		_w5224_,
		_w5228_
	);
	LUT4 #(
		.INIT('h040f)
	) name3479 (
		_w4073_,
		_w4076_,
		_w5227_,
		_w5228_,
		_w5229_
	);
	LUT2 #(
		.INIT('hb)
	) name3480 (
		_w5226_,
		_w5229_,
		_w5230_
	);
	LUT3 #(
		.INIT('h59)
	) name3481 (
		\u1_u3_adr_reg[7]/P0001 ,
		_w2830_,
		_w2832_,
		_w5231_
	);
	LUT3 #(
		.INIT('hb2)
	) name3482 (
		\u1_u3_adr_reg[6]/P0001 ,
		_w2863_,
		_w4065_,
		_w5232_
	);
	LUT3 #(
		.INIT('h01)
	) name3483 (
		_w4062_,
		_w4067_,
		_w4068_,
		_w5233_
	);
	LUT2 #(
		.INIT('h1)
	) name3484 (
		_w5232_,
		_w5233_,
		_w5234_
	);
	LUT4 #(
		.INIT('h00b0)
	) name3485 (
		_w4073_,
		_w4076_,
		_w4079_,
		_w5232_,
		_w5235_
	);
	LUT3 #(
		.INIT('ha9)
	) name3486 (
		_w5231_,
		_w5234_,
		_w5235_,
		_w5236_
	);
	LUT4 #(
		.INIT('h0200)
	) name3487 (
		_w5191_,
		_w5192_,
		_w5193_,
		_w5198_,
		_w5237_
	);
	LUT2 #(
		.INIT('h2)
	) name3488 (
		\u1_u2_sizu_c_reg[0]/P0001 ,
		\u4_csr_reg[0]/P0001 ,
		_w5238_
	);
	LUT2 #(
		.INIT('h2)
	) name3489 (
		_w5216_,
		_w5238_,
		_w5239_
	);
	LUT4 #(
		.INIT('h5010)
	) name3490 (
		\u1_u2_sizu_c_reg[1]/P0001 ,
		\u1_u2_sizu_c_reg[2]/P0001 ,
		\u4_csr_reg[1]/P0001 ,
		\u4_csr_reg[2]/NET0131 ,
		_w5240_
	);
	LUT3 #(
		.INIT('h23)
	) name3491 (
		\u1_u2_sizu_c_reg[2]/P0001 ,
		\u4_csr_reg[17]/P0001 ,
		\u4_csr_reg[2]/NET0131 ,
		_w5241_
	);
	LUT4 #(
		.INIT('h0d00)
	) name3492 (
		_w5216_,
		_w5238_,
		_w5240_,
		_w5241_,
		_w5242_
	);
	LUT4 #(
		.INIT('h00ea)
	) name3493 (
		\u4_csr_reg[17]/P0001 ,
		_w5211_,
		_w5237_,
		_w5242_,
		_w5243_
	);
	LUT2 #(
		.INIT('h1)
	) name3494 (
		_w5209_,
		_w5243_,
		_w5244_
	);
	LUT2 #(
		.INIT('h8)
	) name3495 (
		\u1_u0_pid_reg[0]/NET0131 ,
		\u1_u0_pid_reg[1]/NET0131 ,
		_w5245_
	);
	LUT4 #(
		.INIT('h8000)
	) name3496 (
		rst_i_pad,
		_w4881_,
		_w4884_,
		_w5245_,
		_w5246_
	);
	LUT3 #(
		.INIT('h80)
	) name3497 (
		rst_i_pad,
		\u0_rx_active_reg/P0001 ,
		\u1_u0_state_reg[3]/P0001 ,
		_w5247_
	);
	LUT4 #(
		.INIT('hba00)
	) name3498 (
		_w3671_,
		_w4884_,
		_w4888_,
		_w5247_,
		_w5248_
	);
	LUT2 #(
		.INIT('he)
	) name3499 (
		_w5246_,
		_w5248_,
		_w5249_
	);
	LUT4 #(
		.INIT('hf531)
	) name3500 (
		\u4_u2_buf0_orig_reg[26]/P0001 ,
		\u4_u2_buf0_orig_reg[27]/P0001 ,
		\u4_u2_dma_in_cnt_reg[7]/P0001 ,
		\u4_u2_dma_in_cnt_reg[8]/P0001 ,
		_w5250_
	);
	LUT4 #(
		.INIT('h8caf)
	) name3501 (
		\u4_u2_buf0_orig_reg[25]/P0001 ,
		\u4_u2_buf0_orig_reg[26]/P0001 ,
		\u4_u2_dma_in_cnt_reg[6]/P0001 ,
		\u4_u2_dma_in_cnt_reg[7]/P0001 ,
		_w5251_
	);
	LUT2 #(
		.INIT('h2)
	) name3502 (
		_w5250_,
		_w5251_,
		_w5252_
	);
	LUT4 #(
		.INIT('h8caf)
	) name3503 (
		\u4_u2_buf0_orig_reg[23]/P0001 ,
		\u4_u2_buf0_orig_reg[24]/P0001 ,
		\u4_u2_dma_in_cnt_reg[4]/P0001 ,
		\u4_u2_dma_in_cnt_reg[5]/P0001 ,
		_w5253_
	);
	LUT4 #(
		.INIT('hf531)
	) name3504 (
		\u4_u2_buf0_orig_reg[22]/P0001 ,
		\u4_u2_buf0_orig_reg[23]/P0001 ,
		\u4_u2_dma_in_cnt_reg[3]/P0001 ,
		\u4_u2_dma_in_cnt_reg[4]/P0001 ,
		_w5254_
	);
	LUT2 #(
		.INIT('h2)
	) name3505 (
		_w5253_,
		_w5254_,
		_w5255_
	);
	LUT4 #(
		.INIT('h080a)
	) name3506 (
		\u4_u2_buf0_orig_reg[19]/P0001 ,
		\u4_u2_buf0_orig_reg[20]/P0001 ,
		\u4_u2_dma_in_cnt_reg[0]/P0001 ,
		\u4_u2_dma_in_cnt_reg[1]/P0001 ,
		_w5256_
	);
	LUT4 #(
		.INIT('hf531)
	) name3507 (
		\u4_u2_buf0_orig_reg[20]/P0001 ,
		\u4_u2_buf0_orig_reg[21]/P0001 ,
		\u4_u2_dma_in_cnt_reg[1]/P0001 ,
		\u4_u2_dma_in_cnt_reg[2]/P0001 ,
		_w5257_
	);
	LUT4 #(
		.INIT('h8caf)
	) name3508 (
		\u4_u2_buf0_orig_reg[21]/P0001 ,
		\u4_u2_buf0_orig_reg[22]/P0001 ,
		\u4_u2_dma_in_cnt_reg[2]/P0001 ,
		\u4_u2_dma_in_cnt_reg[3]/P0001 ,
		_w5258_
	);
	LUT4 #(
		.INIT('h8a00)
	) name3509 (
		_w5253_,
		_w5256_,
		_w5257_,
		_w5258_,
		_w5259_
	);
	LUT4 #(
		.INIT('hf531)
	) name3510 (
		\u4_u2_buf0_orig_reg[24]/P0001 ,
		\u4_u2_buf0_orig_reg[25]/P0001 ,
		\u4_u2_dma_in_cnt_reg[5]/P0001 ,
		\u4_u2_dma_in_cnt_reg[6]/P0001 ,
		_w5260_
	);
	LUT2 #(
		.INIT('h8)
	) name3511 (
		_w5250_,
		_w5260_,
		_w5261_
	);
	LUT4 #(
		.INIT('h5455)
	) name3512 (
		_w5252_,
		_w5255_,
		_w5259_,
		_w5261_,
		_w5262_
	);
	LUT2 #(
		.INIT('h4)
	) name3513 (
		\u4_u2_buf0_orig_reg[30]/NET0131 ,
		\u4_u2_dma_in_cnt_reg[11]/P0001 ,
		_w5263_
	);
	LUT2 #(
		.INIT('h2)
	) name3514 (
		\u4_u2_csr1_reg[11]/P0001 ,
		\u4_u2_csr1_reg[12]/P0001 ,
		_w5264_
	);
	LUT3 #(
		.INIT('h08)
	) name3515 (
		\u4_u2_csr1_reg[0]/P0001 ,
		\u4_u2_csr1_reg[11]/P0001 ,
		\u4_u2_csr1_reg[12]/P0001 ,
		_w5265_
	);
	LUT4 #(
		.INIT('h5010)
	) name3516 (
		\u4_u2_buf0_orig_reg[29]/NET0131 ,
		\u4_u2_buf0_orig_reg[30]/NET0131 ,
		\u4_u2_dma_in_cnt_reg[10]/P0001 ,
		\u4_u2_dma_in_cnt_reg[11]/P0001 ,
		_w5266_
	);
	LUT4 #(
		.INIT('h8caf)
	) name3517 (
		\u4_u2_buf0_orig_reg[27]/P0001 ,
		\u4_u2_buf0_orig_reg[28]/P0001 ,
		\u4_u2_dma_in_cnt_reg[8]/P0001 ,
		\u4_u2_dma_in_cnt_reg[9]/P0001 ,
		_w5267_
	);
	LUT4 #(
		.INIT('h0400)
	) name3518 (
		_w5263_,
		_w5265_,
		_w5266_,
		_w5267_,
		_w5268_
	);
	LUT2 #(
		.INIT('h2)
	) name3519 (
		\u4_u2_buf0_orig_reg[28]/P0001 ,
		\u4_u2_dma_in_cnt_reg[9]/P0001 ,
		_w5269_
	);
	LUT4 #(
		.INIT('hf531)
	) name3520 (
		\u4_u2_buf0_orig_reg[29]/NET0131 ,
		\u4_u2_buf0_orig_reg[30]/NET0131 ,
		\u4_u2_dma_in_cnt_reg[10]/P0001 ,
		\u4_u2_dma_in_cnt_reg[11]/P0001 ,
		_w5270_
	);
	LUT4 #(
		.INIT('h4044)
	) name3521 (
		_w5263_,
		_w5265_,
		_w5269_,
		_w5270_,
		_w5271_
	);
	LUT3 #(
		.INIT('h01)
	) name3522 (
		\u4_u2_dma_out_cnt_reg[10]/P0001 ,
		\u4_u2_dma_out_cnt_reg[4]/P0001 ,
		\u4_u2_dma_out_cnt_reg[5]/P0001 ,
		_w5272_
	);
	LUT3 #(
		.INIT('h01)
	) name3523 (
		\u4_u2_dma_out_cnt_reg[11]/P0001 ,
		\u4_u2_dma_out_cnt_reg[2]/P0001 ,
		\u4_u2_dma_out_cnt_reg[3]/P0001 ,
		_w5273_
	);
	LUT4 #(
		.INIT('h8000)
	) name3524 (
		_w4743_,
		_w5048_,
		_w5272_,
		_w5273_,
		_w5274_
	);
	LUT3 #(
		.INIT('h20)
	) name3525 (
		\u4_u2_csr1_reg[0]/P0001 ,
		\u4_u2_csr1_reg[11]/P0001 ,
		\u4_u2_csr1_reg[12]/P0001 ,
		_w5275_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name3526 (
		_w5266_,
		_w5271_,
		_w5274_,
		_w5275_,
		_w5276_
	);
	LUT3 #(
		.INIT('h01)
	) name3527 (
		\u4_u2_r2_reg/P0001 ,
		\u4_u2_r4_reg/P0001 ,
		\u4_u2_r5_reg/NET0131 ,
		_w5277_
	);
	LUT4 #(
		.INIT('h8f00)
	) name3528 (
		_w5262_,
		_w5268_,
		_w5276_,
		_w5277_,
		_w5278_
	);
	LUT2 #(
		.INIT('h2)
	) name3529 (
		\u4_u3_buf0_orig_reg[26]/P0001 ,
		\u4_u3_dma_in_cnt_reg[7]/P0001 ,
		_w5279_
	);
	LUT4 #(
		.INIT('hf531)
	) name3530 (
		\u4_u3_buf0_orig_reg[27]/P0001 ,
		\u4_u3_buf0_orig_reg[28]/P0001 ,
		\u4_u3_dma_in_cnt_reg[8]/P0001 ,
		\u4_u3_dma_in_cnt_reg[9]/P0001 ,
		_w5280_
	);
	LUT4 #(
		.INIT('h8caf)
	) name3531 (
		\u4_u3_buf0_orig_reg[25]/P0001 ,
		\u4_u3_buf0_orig_reg[26]/P0001 ,
		\u4_u3_dma_in_cnt_reg[6]/P0001 ,
		\u4_u3_dma_in_cnt_reg[7]/P0001 ,
		_w5281_
	);
	LUT3 #(
		.INIT('h04)
	) name3532 (
		_w5279_,
		_w5280_,
		_w5281_,
		_w5282_
	);
	LUT4 #(
		.INIT('h8caf)
	) name3533 (
		\u4_u3_buf0_orig_reg[23]/P0001 ,
		\u4_u3_buf0_orig_reg[24]/P0001 ,
		\u4_u3_dma_in_cnt_reg[4]/P0001 ,
		\u4_u3_dma_in_cnt_reg[5]/P0001 ,
		_w5283_
	);
	LUT4 #(
		.INIT('hf531)
	) name3534 (
		\u4_u3_buf0_orig_reg[22]/P0001 ,
		\u4_u3_buf0_orig_reg[23]/P0001 ,
		\u4_u3_dma_in_cnt_reg[3]/P0001 ,
		\u4_u3_dma_in_cnt_reg[4]/P0001 ,
		_w5284_
	);
	LUT2 #(
		.INIT('h2)
	) name3535 (
		_w5283_,
		_w5284_,
		_w5285_
	);
	LUT4 #(
		.INIT('h08cc)
	) name3536 (
		\u4_u3_buf0_orig_reg[19]/P0001 ,
		\u4_u3_buf0_orig_reg[20]/P0001 ,
		\u4_u3_dma_in_cnt_reg[0]/P0001 ,
		\u4_u3_dma_in_cnt_reg[1]/P0001 ,
		_w5286_
	);
	LUT2 #(
		.INIT('h2)
	) name3537 (
		\u4_u3_buf0_orig_reg[21]/P0001 ,
		\u4_u3_dma_in_cnt_reg[2]/P0001 ,
		_w5287_
	);
	LUT3 #(
		.INIT('h02)
	) name3538 (
		\u4_u3_buf0_orig_reg[19]/P0001 ,
		\u4_u3_dma_in_cnt_reg[0]/P0001 ,
		\u4_u3_dma_in_cnt_reg[1]/P0001 ,
		_w5288_
	);
	LUT3 #(
		.INIT('h01)
	) name3539 (
		_w5286_,
		_w5287_,
		_w5288_,
		_w5289_
	);
	LUT4 #(
		.INIT('h8caf)
	) name3540 (
		\u4_u3_buf0_orig_reg[21]/P0001 ,
		\u4_u3_buf0_orig_reg[22]/P0001 ,
		\u4_u3_dma_in_cnt_reg[2]/P0001 ,
		\u4_u3_dma_in_cnt_reg[3]/P0001 ,
		_w5290_
	);
	LUT2 #(
		.INIT('h8)
	) name3541 (
		_w5283_,
		_w5290_,
		_w5291_
	);
	LUT4 #(
		.INIT('hf531)
	) name3542 (
		\u4_u3_buf0_orig_reg[24]/P0001 ,
		\u4_u3_buf0_orig_reg[25]/P0001 ,
		\u4_u3_dma_in_cnt_reg[5]/P0001 ,
		\u4_u3_dma_in_cnt_reg[6]/P0001 ,
		_w5292_
	);
	LUT3 #(
		.INIT('h40)
	) name3543 (
		_w5279_,
		_w5280_,
		_w5292_,
		_w5293_
	);
	LUT4 #(
		.INIT('h4500)
	) name3544 (
		_w5285_,
		_w5289_,
		_w5291_,
		_w5293_,
		_w5294_
	);
	LUT4 #(
		.INIT('h5010)
	) name3545 (
		\u4_u3_buf0_orig_reg[29]/NET0131 ,
		\u4_u3_buf0_orig_reg[30]/NET0131 ,
		\u4_u3_dma_in_cnt_reg[10]/P0001 ,
		\u4_u3_dma_in_cnt_reg[11]/P0001 ,
		_w5295_
	);
	LUT2 #(
		.INIT('h4)
	) name3546 (
		\u4_u3_buf0_orig_reg[30]/NET0131 ,
		\u4_u3_dma_in_cnt_reg[11]/P0001 ,
		_w5296_
	);
	LUT2 #(
		.INIT('h2)
	) name3547 (
		\u4_u3_csr1_reg[11]/P0001 ,
		\u4_u3_csr1_reg[12]/P0001 ,
		_w5297_
	);
	LUT3 #(
		.INIT('h08)
	) name3548 (
		\u4_u3_csr1_reg[0]/P0001 ,
		\u4_u3_csr1_reg[11]/P0001 ,
		\u4_u3_csr1_reg[12]/P0001 ,
		_w5298_
	);
	LUT4 #(
		.INIT('h8cef)
	) name3549 (
		\u4_u3_buf0_orig_reg[27]/P0001 ,
		\u4_u3_buf0_orig_reg[28]/P0001 ,
		\u4_u3_dma_in_cnt_reg[8]/P0001 ,
		\u4_u3_dma_in_cnt_reg[9]/P0001 ,
		_w5299_
	);
	LUT4 #(
		.INIT('h1000)
	) name3550 (
		_w5295_,
		_w5296_,
		_w5298_,
		_w5299_,
		_w5300_
	);
	LUT4 #(
		.INIT('h0ace)
	) name3551 (
		\u4_u3_buf0_orig_reg[29]/NET0131 ,
		\u4_u3_buf0_orig_reg[30]/NET0131 ,
		\u4_u3_dma_in_cnt_reg[10]/P0001 ,
		\u4_u3_dma_in_cnt_reg[11]/P0001 ,
		_w5301_
	);
	LUT3 #(
		.INIT('h40)
	) name3552 (
		_w5296_,
		_w5298_,
		_w5301_,
		_w5302_
	);
	LUT3 #(
		.INIT('h01)
	) name3553 (
		\u4_u3_dma_out_cnt_reg[10]/P0001 ,
		\u4_u3_dma_out_cnt_reg[4]/P0001 ,
		\u4_u3_dma_out_cnt_reg[5]/P0001 ,
		_w5303_
	);
	LUT3 #(
		.INIT('h01)
	) name3554 (
		\u4_u3_dma_out_cnt_reg[11]/P0001 ,
		\u4_u3_dma_out_cnt_reg[2]/P0001 ,
		\u4_u3_dma_out_cnt_reg[3]/P0001 ,
		_w5304_
	);
	LUT4 #(
		.INIT('h8000)
	) name3555 (
		_w4651_,
		_w4954_,
		_w5303_,
		_w5304_,
		_w5305_
	);
	LUT3 #(
		.INIT('h20)
	) name3556 (
		\u4_u3_csr1_reg[0]/P0001 ,
		\u4_u3_csr1_reg[11]/P0001 ,
		\u4_u3_csr1_reg[12]/P0001 ,
		_w5306_
	);
	LUT3 #(
		.INIT('h45)
	) name3557 (
		_w5302_,
		_w5305_,
		_w5306_,
		_w5307_
	);
	LUT4 #(
		.INIT('hef00)
	) name3558 (
		_w5282_,
		_w5294_,
		_w5300_,
		_w5307_,
		_w5308_
	);
	LUT3 #(
		.INIT('h01)
	) name3559 (
		\u4_u3_r2_reg/P0001 ,
		\u4_u3_r4_reg/P0001 ,
		\u4_u3_r5_reg/NET0131 ,
		_w5309_
	);
	LUT2 #(
		.INIT('h4)
	) name3560 (
		_w5308_,
		_w5309_,
		_w5310_
	);
	LUT4 #(
		.INIT('h8000)
	) name3561 (
		\u1_u2_sizu_c_reg[10]/P0001 ,
		\u1_u2_sizu_c_reg[6]/P0001 ,
		\u1_u2_sizu_c_reg[7]/P0001 ,
		\u1_u2_sizu_c_reg[9]/P0001 ,
		_w5311_
	);
	LUT3 #(
		.INIT('h80)
	) name3562 (
		_w4783_,
		_w4788_,
		_w5311_,
		_w5312_
	);
	LUT3 #(
		.INIT('h20)
	) name3563 (
		rst_i_pad,
		\u1_u2_rx_dma_en_r_reg/P0001 ,
		\u1_u2_sizu_c_reg[10]/P0001 ,
		_w5313_
	);
	LUT3 #(
		.INIT('h20)
	) name3564 (
		rst_i_pad,
		\u1_u2_rx_dma_en_r_reg/P0001 ,
		\u1_u2_sizu_c_reg[9]/P0001 ,
		_w5314_
	);
	LUT4 #(
		.INIT('h8000)
	) name3565 (
		_w4783_,
		_w4785_,
		_w4788_,
		_w5314_,
		_w5315_
	);
	LUT3 #(
		.INIT('h54)
	) name3566 (
		_w5312_,
		_w5313_,
		_w5315_,
		_w5316_
	);
	LUT2 #(
		.INIT('h4)
	) name3567 (
		\u1_u2_word_done_r_reg/P0001 ,
		\u1_u2_word_done_reg/NET0131 ,
		_w5317_
	);
	LUT4 #(
		.INIT('h0002)
	) name3568 (
		\u5_state_reg[0]/P0001 ,
		\u5_state_reg[1]/P0001 ,
		\u5_state_reg[2]/P0001 ,
		\u5_wb_req_s1_reg/P0001 ,
		_w5318_
	);
	LUT2 #(
		.INIT('h8)
	) name3569 (
		_w2224_,
		_w5318_,
		_w5319_
	);
	LUT2 #(
		.INIT('h1)
	) name3570 (
		\u5_state_reg[3]/P0001 ,
		\u5_state_reg[4]/P0001 ,
		_w5320_
	);
	LUT4 #(
		.INIT('h0100)
	) name3571 (
		\u5_state_reg[0]/P0001 ,
		\u5_state_reg[1]/P0001 ,
		\u5_state_reg[2]/P0001 ,
		\u5_state_reg[5]/NET0131 ,
		_w5321_
	);
	LUT3 #(
		.INIT('h2a)
	) name3572 (
		rst_i_pad,
		_w5320_,
		_w5321_,
		_w5322_
	);
	LUT2 #(
		.INIT('hb)
	) name3573 (
		_w5319_,
		_w5322_,
		_w5323_
	);
	LUT2 #(
		.INIT('h8)
	) name3574 (
		\u1_u2_rx_data_st_r_reg[2]/P0001 ,
		\u1_u2_rx_data_valid_r_reg/NET0131 ,
		_w5324_
	);
	LUT3 #(
		.INIT('h02)
	) name3575 (
		\u1_u2_adr_cb_reg[0]/NET0131 ,
		\u1_u2_adr_cb_reg[1]/NET0131 ,
		\u1_u2_dtmp_sel_r_reg/P0001 ,
		_w5325_
	);
	LUT3 #(
		.INIT('h20)
	) name3576 (
		\u1_u2_adr_cb_reg[0]/NET0131 ,
		\u1_u2_adr_cb_reg[1]/NET0131 ,
		\u1_u2_rx_data_valid_r_reg/NET0131 ,
		_w5326_
	);
	LUT2 #(
		.INIT('h2)
	) name3577 (
		\u1_u2_dtmp_r_reg[10]/P0001 ,
		\u1_u2_dtmp_sel_r_reg/P0001 ,
		_w5327_
	);
	LUT4 #(
		.INIT('h7077)
	) name3578 (
		_w5324_,
		_w5325_,
		_w5326_,
		_w5327_,
		_w5328_
	);
	LUT2 #(
		.INIT('h8)
	) name3579 (
		\sram_data_i[10]_pad ,
		\u1_u2_dtmp_sel_r_reg/P0001 ,
		_w5329_
	);
	LUT2 #(
		.INIT('hd)
	) name3580 (
		_w5328_,
		_w5329_,
		_w5330_
	);
	LUT2 #(
		.INIT('h8)
	) name3581 (
		\u1_u2_rx_data_st_r_reg[3]/P0001 ,
		\u1_u2_rx_data_valid_r_reg/NET0131 ,
		_w5331_
	);
	LUT2 #(
		.INIT('h8)
	) name3582 (
		_w5325_,
		_w5331_,
		_w5332_
	);
	LUT2 #(
		.INIT('h2)
	) name3583 (
		\u1_u2_dtmp_r_reg[11]/P0001 ,
		\u1_u2_dtmp_sel_r_reg/P0001 ,
		_w5333_
	);
	LUT2 #(
		.INIT('h8)
	) name3584 (
		\sram_data_i[11]_pad ,
		\u1_u2_dtmp_sel_r_reg/P0001 ,
		_w5334_
	);
	LUT3 #(
		.INIT('h0b)
	) name3585 (
		_w5326_,
		_w5333_,
		_w5334_,
		_w5335_
	);
	LUT2 #(
		.INIT('hb)
	) name3586 (
		_w5332_,
		_w5335_,
		_w5336_
	);
	LUT2 #(
		.INIT('h8)
	) name3587 (
		\u1_u2_rx_data_st_r_reg[4]/P0001 ,
		\u1_u2_rx_data_valid_r_reg/NET0131 ,
		_w5337_
	);
	LUT2 #(
		.INIT('h8)
	) name3588 (
		_w5325_,
		_w5337_,
		_w5338_
	);
	LUT2 #(
		.INIT('h2)
	) name3589 (
		\u1_u2_dtmp_r_reg[12]/P0001 ,
		\u1_u2_dtmp_sel_r_reg/P0001 ,
		_w5339_
	);
	LUT2 #(
		.INIT('h8)
	) name3590 (
		\sram_data_i[12]_pad ,
		\u1_u2_dtmp_sel_r_reg/P0001 ,
		_w5340_
	);
	LUT3 #(
		.INIT('h0b)
	) name3591 (
		_w5326_,
		_w5339_,
		_w5340_,
		_w5341_
	);
	LUT2 #(
		.INIT('hb)
	) name3592 (
		_w5338_,
		_w5341_,
		_w5342_
	);
	LUT2 #(
		.INIT('h8)
	) name3593 (
		\u1_u2_rx_data_st_r_reg[5]/P0001 ,
		\u1_u2_rx_data_valid_r_reg/NET0131 ,
		_w5343_
	);
	LUT2 #(
		.INIT('h8)
	) name3594 (
		_w5325_,
		_w5343_,
		_w5344_
	);
	LUT2 #(
		.INIT('h2)
	) name3595 (
		\u1_u2_dtmp_r_reg[13]/P0001 ,
		\u1_u2_dtmp_sel_r_reg/P0001 ,
		_w5345_
	);
	LUT2 #(
		.INIT('h8)
	) name3596 (
		\sram_data_i[13]_pad ,
		\u1_u2_dtmp_sel_r_reg/P0001 ,
		_w5346_
	);
	LUT3 #(
		.INIT('h0b)
	) name3597 (
		_w5326_,
		_w5345_,
		_w5346_,
		_w5347_
	);
	LUT2 #(
		.INIT('hb)
	) name3598 (
		_w5344_,
		_w5347_,
		_w5348_
	);
	LUT2 #(
		.INIT('h8)
	) name3599 (
		\u1_u2_rx_data_st_r_reg[6]/P0001 ,
		\u1_u2_rx_data_valid_r_reg/NET0131 ,
		_w5349_
	);
	LUT2 #(
		.INIT('h2)
	) name3600 (
		\u1_u2_dtmp_r_reg[14]/P0001 ,
		\u1_u2_dtmp_sel_r_reg/P0001 ,
		_w5350_
	);
	LUT4 #(
		.INIT('h4c5f)
	) name3601 (
		_w5325_,
		_w5326_,
		_w5349_,
		_w5350_,
		_w5351_
	);
	LUT2 #(
		.INIT('h8)
	) name3602 (
		\sram_data_i[14]_pad ,
		\u1_u2_dtmp_sel_r_reg/P0001 ,
		_w5352_
	);
	LUT2 #(
		.INIT('hd)
	) name3603 (
		_w5351_,
		_w5352_,
		_w5353_
	);
	LUT2 #(
		.INIT('h8)
	) name3604 (
		\u1_u2_rx_data_st_r_reg[7]/P0001 ,
		\u1_u2_rx_data_valid_r_reg/NET0131 ,
		_w5354_
	);
	LUT2 #(
		.INIT('h2)
	) name3605 (
		\u1_u2_dtmp_r_reg[15]/P0001 ,
		\u1_u2_dtmp_sel_r_reg/P0001 ,
		_w5355_
	);
	LUT4 #(
		.INIT('h4c5f)
	) name3606 (
		_w5325_,
		_w5326_,
		_w5354_,
		_w5355_,
		_w5356_
	);
	LUT2 #(
		.INIT('h8)
	) name3607 (
		\sram_data_i[15]_pad ,
		\u1_u2_dtmp_sel_r_reg/P0001 ,
		_w5357_
	);
	LUT2 #(
		.INIT('hd)
	) name3608 (
		_w5356_,
		_w5357_,
		_w5358_
	);
	LUT2 #(
		.INIT('h8)
	) name3609 (
		\u1_u2_rx_data_st_r_reg[0]/P0001 ,
		\u1_u2_rx_data_valid_r_reg/NET0131 ,
		_w5359_
	);
	LUT3 #(
		.INIT('h40)
	) name3610 (
		\u1_u2_dtmp_sel_r_reg/P0001 ,
		\u1_u2_rx_data_st_r_reg[0]/P0001 ,
		\u1_u2_rx_data_valid_r_reg/NET0131 ,
		_w5360_
	);
	LUT2 #(
		.INIT('h2)
	) name3611 (
		\u1_u2_dtmp_r_reg[16]/P0001 ,
		\u1_u2_dtmp_sel_r_reg/P0001 ,
		_w5361_
	);
	LUT4 #(
		.INIT('h083f)
	) name3612 (
		\u1_u2_rx_data_valid_r_reg/NET0131 ,
		_w3191_,
		_w5360_,
		_w5361_,
		_w5362_
	);
	LUT2 #(
		.INIT('h8)
	) name3613 (
		\sram_data_i[16]_pad ,
		\u1_u2_dtmp_sel_r_reg/P0001 ,
		_w5363_
	);
	LUT2 #(
		.INIT('hd)
	) name3614 (
		_w5362_,
		_w5363_,
		_w5364_
	);
	LUT2 #(
		.INIT('h8)
	) name3615 (
		\u1_u2_rx_data_st_r_reg[1]/P0001 ,
		\u1_u2_rx_data_valid_r_reg/NET0131 ,
		_w5365_
	);
	LUT3 #(
		.INIT('h40)
	) name3616 (
		\u1_u2_dtmp_sel_r_reg/P0001 ,
		\u1_u2_rx_data_st_r_reg[1]/P0001 ,
		\u1_u2_rx_data_valid_r_reg/NET0131 ,
		_w5366_
	);
	LUT2 #(
		.INIT('h2)
	) name3617 (
		\u1_u2_dtmp_r_reg[17]/P0001 ,
		\u1_u2_dtmp_sel_r_reg/P0001 ,
		_w5367_
	);
	LUT4 #(
		.INIT('h083f)
	) name3618 (
		\u1_u2_rx_data_valid_r_reg/NET0131 ,
		_w3191_,
		_w5366_,
		_w5367_,
		_w5368_
	);
	LUT2 #(
		.INIT('h8)
	) name3619 (
		\sram_data_i[17]_pad ,
		\u1_u2_dtmp_sel_r_reg/P0001 ,
		_w5369_
	);
	LUT2 #(
		.INIT('hd)
	) name3620 (
		_w5368_,
		_w5369_,
		_w5370_
	);
	LUT3 #(
		.INIT('h40)
	) name3621 (
		\u1_u2_dtmp_sel_r_reg/P0001 ,
		\u1_u2_rx_data_st_r_reg[2]/P0001 ,
		\u1_u2_rx_data_valid_r_reg/NET0131 ,
		_w5371_
	);
	LUT2 #(
		.INIT('h2)
	) name3622 (
		\u1_u2_dtmp_r_reg[18]/P0001 ,
		\u1_u2_dtmp_sel_r_reg/P0001 ,
		_w5372_
	);
	LUT4 #(
		.INIT('h083f)
	) name3623 (
		\u1_u2_rx_data_valid_r_reg/NET0131 ,
		_w3191_,
		_w5371_,
		_w5372_,
		_w5373_
	);
	LUT2 #(
		.INIT('h8)
	) name3624 (
		\sram_data_i[18]_pad ,
		\u1_u2_dtmp_sel_r_reg/P0001 ,
		_w5374_
	);
	LUT2 #(
		.INIT('hd)
	) name3625 (
		_w5373_,
		_w5374_,
		_w5375_
	);
	LUT3 #(
		.INIT('h40)
	) name3626 (
		\u1_u2_dtmp_sel_r_reg/P0001 ,
		\u1_u2_rx_data_st_r_reg[3]/P0001 ,
		\u1_u2_rx_data_valid_r_reg/NET0131 ,
		_w5376_
	);
	LUT2 #(
		.INIT('h2)
	) name3627 (
		\u1_u2_dtmp_r_reg[19]/P0001 ,
		\u1_u2_dtmp_sel_r_reg/P0001 ,
		_w5377_
	);
	LUT4 #(
		.INIT('h083f)
	) name3628 (
		\u1_u2_rx_data_valid_r_reg/NET0131 ,
		_w3191_,
		_w5376_,
		_w5377_,
		_w5378_
	);
	LUT2 #(
		.INIT('h8)
	) name3629 (
		\sram_data_i[19]_pad ,
		\u1_u2_dtmp_sel_r_reg/P0001 ,
		_w5379_
	);
	LUT2 #(
		.INIT('hd)
	) name3630 (
		_w5378_,
		_w5379_,
		_w5380_
	);
	LUT3 #(
		.INIT('h40)
	) name3631 (
		\u1_u2_dtmp_sel_r_reg/P0001 ,
		\u1_u2_rx_data_st_r_reg[4]/P0001 ,
		\u1_u2_rx_data_valid_r_reg/NET0131 ,
		_w5381_
	);
	LUT2 #(
		.INIT('h2)
	) name3632 (
		\u1_u2_dtmp_r_reg[20]/P0001 ,
		\u1_u2_dtmp_sel_r_reg/P0001 ,
		_w5382_
	);
	LUT4 #(
		.INIT('h083f)
	) name3633 (
		\u1_u2_rx_data_valid_r_reg/NET0131 ,
		_w3191_,
		_w5381_,
		_w5382_,
		_w5383_
	);
	LUT2 #(
		.INIT('h8)
	) name3634 (
		\sram_data_i[20]_pad ,
		\u1_u2_dtmp_sel_r_reg/P0001 ,
		_w5384_
	);
	LUT2 #(
		.INIT('hd)
	) name3635 (
		_w5383_,
		_w5384_,
		_w5385_
	);
	LUT3 #(
		.INIT('h40)
	) name3636 (
		\u1_u2_dtmp_sel_r_reg/P0001 ,
		\u1_u2_rx_data_st_r_reg[5]/P0001 ,
		\u1_u2_rx_data_valid_r_reg/NET0131 ,
		_w5386_
	);
	LUT2 #(
		.INIT('h2)
	) name3637 (
		\u1_u2_dtmp_r_reg[21]/P0001 ,
		\u1_u2_dtmp_sel_r_reg/P0001 ,
		_w5387_
	);
	LUT4 #(
		.INIT('h083f)
	) name3638 (
		\u1_u2_rx_data_valid_r_reg/NET0131 ,
		_w3191_,
		_w5386_,
		_w5387_,
		_w5388_
	);
	LUT2 #(
		.INIT('h8)
	) name3639 (
		\sram_data_i[21]_pad ,
		\u1_u2_dtmp_sel_r_reg/P0001 ,
		_w5389_
	);
	LUT2 #(
		.INIT('hd)
	) name3640 (
		_w5388_,
		_w5389_,
		_w5390_
	);
	LUT3 #(
		.INIT('h40)
	) name3641 (
		\u1_u2_dtmp_sel_r_reg/P0001 ,
		\u1_u2_rx_data_st_r_reg[6]/P0001 ,
		\u1_u2_rx_data_valid_r_reg/NET0131 ,
		_w5391_
	);
	LUT2 #(
		.INIT('h2)
	) name3642 (
		\u1_u2_dtmp_r_reg[22]/P0001 ,
		\u1_u2_dtmp_sel_r_reg/P0001 ,
		_w5392_
	);
	LUT4 #(
		.INIT('h083f)
	) name3643 (
		\u1_u2_rx_data_valid_r_reg/NET0131 ,
		_w3191_,
		_w5391_,
		_w5392_,
		_w5393_
	);
	LUT2 #(
		.INIT('h8)
	) name3644 (
		\sram_data_i[22]_pad ,
		\u1_u2_dtmp_sel_r_reg/P0001 ,
		_w5394_
	);
	LUT2 #(
		.INIT('hd)
	) name3645 (
		_w5393_,
		_w5394_,
		_w5395_
	);
	LUT3 #(
		.INIT('h40)
	) name3646 (
		\u1_u2_dtmp_sel_r_reg/P0001 ,
		\u1_u2_rx_data_st_r_reg[7]/P0001 ,
		\u1_u2_rx_data_valid_r_reg/NET0131 ,
		_w5396_
	);
	LUT2 #(
		.INIT('h2)
	) name3647 (
		\u1_u2_dtmp_r_reg[23]/P0001 ,
		\u1_u2_dtmp_sel_r_reg/P0001 ,
		_w5397_
	);
	LUT4 #(
		.INIT('h083f)
	) name3648 (
		\u1_u2_rx_data_valid_r_reg/NET0131 ,
		_w3191_,
		_w5396_,
		_w5397_,
		_w5398_
	);
	LUT2 #(
		.INIT('h8)
	) name3649 (
		\sram_data_i[23]_pad ,
		\u1_u2_dtmp_sel_r_reg/P0001 ,
		_w5399_
	);
	LUT2 #(
		.INIT('hd)
	) name3650 (
		_w5398_,
		_w5399_,
		_w5400_
	);
	LUT3 #(
		.INIT('h80)
	) name3651 (
		\u1_u2_adr_cb_reg[0]/NET0131 ,
		\u1_u2_adr_cb_reg[1]/NET0131 ,
		\u1_u2_rx_data_valid_r_reg/NET0131 ,
		_w5401_
	);
	LUT2 #(
		.INIT('h2)
	) name3652 (
		\u1_u2_dtmp_r_reg[24]/P0001 ,
		\u1_u2_dtmp_sel_r_reg/P0001 ,
		_w5402_
	);
	LUT4 #(
		.INIT('h083f)
	) name3653 (
		\u1_u2_rx_data_valid_r_reg/NET0131 ,
		_w3182_,
		_w5360_,
		_w5402_,
		_w5403_
	);
	LUT2 #(
		.INIT('h8)
	) name3654 (
		\sram_data_i[24]_pad ,
		\u1_u2_dtmp_sel_r_reg/P0001 ,
		_w5404_
	);
	LUT2 #(
		.INIT('hd)
	) name3655 (
		_w5403_,
		_w5404_,
		_w5405_
	);
	LUT2 #(
		.INIT('h8)
	) name3656 (
		_w3182_,
		_w5366_,
		_w5406_
	);
	LUT2 #(
		.INIT('h2)
	) name3657 (
		\u1_u2_dtmp_r_reg[25]/P0001 ,
		\u1_u2_dtmp_sel_r_reg/P0001 ,
		_w5407_
	);
	LUT2 #(
		.INIT('h8)
	) name3658 (
		\sram_data_i[25]_pad ,
		\u1_u2_dtmp_sel_r_reg/P0001 ,
		_w5408_
	);
	LUT3 #(
		.INIT('h0b)
	) name3659 (
		_w5401_,
		_w5407_,
		_w5408_,
		_w5409_
	);
	LUT2 #(
		.INIT('hb)
	) name3660 (
		_w5406_,
		_w5409_,
		_w5410_
	);
	LUT4 #(
		.INIT('h0800)
	) name3661 (
		\u1_u2_adr_cb_reg[0]/NET0131 ,
		\u1_u2_adr_cb_reg[1]/NET0131 ,
		\u1_u2_dtmp_sel_r_reg/P0001 ,
		\u1_u2_rx_data_valid_r_reg/NET0131 ,
		_w5411_
	);
	LUT2 #(
		.INIT('h8)
	) name3662 (
		\u1_u2_rx_data_st_r_reg[2]/P0001 ,
		_w5411_,
		_w5412_
	);
	LUT2 #(
		.INIT('h2)
	) name3663 (
		\u1_u2_dtmp_r_reg[26]/P0001 ,
		\u1_u2_dtmp_sel_r_reg/P0001 ,
		_w5413_
	);
	LUT2 #(
		.INIT('h8)
	) name3664 (
		\sram_data_i[26]_pad ,
		\u1_u2_dtmp_sel_r_reg/P0001 ,
		_w5414_
	);
	LUT3 #(
		.INIT('h0b)
	) name3665 (
		_w5401_,
		_w5413_,
		_w5414_,
		_w5415_
	);
	LUT2 #(
		.INIT('hb)
	) name3666 (
		_w5412_,
		_w5415_,
		_w5416_
	);
	LUT2 #(
		.INIT('h8)
	) name3667 (
		\u1_u2_rx_data_st_r_reg[3]/P0001 ,
		_w5411_,
		_w5417_
	);
	LUT2 #(
		.INIT('h2)
	) name3668 (
		\u1_u2_dtmp_r_reg[27]/P0001 ,
		\u1_u2_dtmp_sel_r_reg/P0001 ,
		_w5418_
	);
	LUT2 #(
		.INIT('h8)
	) name3669 (
		\sram_data_i[27]_pad ,
		\u1_u2_dtmp_sel_r_reg/P0001 ,
		_w5419_
	);
	LUT3 #(
		.INIT('h0b)
	) name3670 (
		_w5401_,
		_w5418_,
		_w5419_,
		_w5420_
	);
	LUT2 #(
		.INIT('hb)
	) name3671 (
		_w5417_,
		_w5420_,
		_w5421_
	);
	LUT2 #(
		.INIT('h8)
	) name3672 (
		\u1_u2_rx_data_st_r_reg[4]/P0001 ,
		_w5411_,
		_w5422_
	);
	LUT2 #(
		.INIT('h2)
	) name3673 (
		\u1_u2_dtmp_r_reg[28]/P0001 ,
		\u1_u2_dtmp_sel_r_reg/P0001 ,
		_w5423_
	);
	LUT2 #(
		.INIT('h8)
	) name3674 (
		\sram_data_i[28]_pad ,
		\u1_u2_dtmp_sel_r_reg/P0001 ,
		_w5424_
	);
	LUT3 #(
		.INIT('h0b)
	) name3675 (
		_w5401_,
		_w5423_,
		_w5424_,
		_w5425_
	);
	LUT2 #(
		.INIT('hb)
	) name3676 (
		_w5422_,
		_w5425_,
		_w5426_
	);
	LUT2 #(
		.INIT('h8)
	) name3677 (
		\u1_u2_rx_data_st_r_reg[5]/P0001 ,
		_w5411_,
		_w5427_
	);
	LUT2 #(
		.INIT('h2)
	) name3678 (
		\u1_u2_dtmp_r_reg[29]/P0001 ,
		\u1_u2_dtmp_sel_r_reg/P0001 ,
		_w5428_
	);
	LUT2 #(
		.INIT('h8)
	) name3679 (
		\sram_data_i[29]_pad ,
		\u1_u2_dtmp_sel_r_reg/P0001 ,
		_w5429_
	);
	LUT3 #(
		.INIT('h0b)
	) name3680 (
		_w5401_,
		_w5428_,
		_w5429_,
		_w5430_
	);
	LUT2 #(
		.INIT('hb)
	) name3681 (
		_w5427_,
		_w5430_,
		_w5431_
	);
	LUT2 #(
		.INIT('h8)
	) name3682 (
		\u1_u2_rx_data_st_r_reg[6]/P0001 ,
		_w5411_,
		_w5432_
	);
	LUT2 #(
		.INIT('h2)
	) name3683 (
		\u1_u2_dtmp_r_reg[30]/P0001 ,
		\u1_u2_dtmp_sel_r_reg/P0001 ,
		_w5433_
	);
	LUT2 #(
		.INIT('h8)
	) name3684 (
		\sram_data_i[30]_pad ,
		\u1_u2_dtmp_sel_r_reg/P0001 ,
		_w5434_
	);
	LUT3 #(
		.INIT('h0b)
	) name3685 (
		_w5401_,
		_w5433_,
		_w5434_,
		_w5435_
	);
	LUT2 #(
		.INIT('hb)
	) name3686 (
		_w5432_,
		_w5435_,
		_w5436_
	);
	LUT2 #(
		.INIT('h8)
	) name3687 (
		_w3182_,
		_w5396_,
		_w5437_
	);
	LUT2 #(
		.INIT('h2)
	) name3688 (
		\u1_u2_dtmp_r_reg[31]/P0001 ,
		\u1_u2_dtmp_sel_r_reg/P0001 ,
		_w5438_
	);
	LUT2 #(
		.INIT('h8)
	) name3689 (
		\sram_data_i[31]_pad ,
		\u1_u2_dtmp_sel_r_reg/P0001 ,
		_w5439_
	);
	LUT3 #(
		.INIT('h0b)
	) name3690 (
		_w5401_,
		_w5438_,
		_w5439_,
		_w5440_
	);
	LUT2 #(
		.INIT('hb)
	) name3691 (
		_w5437_,
		_w5440_,
		_w5441_
	);
	LUT2 #(
		.INIT('h2)
	) name3692 (
		\u1_u2_dtmp_r_reg[8]/P0001 ,
		\u1_u2_dtmp_sel_r_reg/P0001 ,
		_w5442_
	);
	LUT4 #(
		.INIT('h4c5f)
	) name3693 (
		_w5325_,
		_w5326_,
		_w5359_,
		_w5442_,
		_w5443_
	);
	LUT2 #(
		.INIT('h8)
	) name3694 (
		\sram_data_i[8]_pad ,
		\u1_u2_dtmp_sel_r_reg/P0001 ,
		_w5444_
	);
	LUT2 #(
		.INIT('hd)
	) name3695 (
		_w5443_,
		_w5444_,
		_w5445_
	);
	LUT2 #(
		.INIT('h2)
	) name3696 (
		\u1_u2_dtmp_r_reg[9]/P0001 ,
		\u1_u2_dtmp_sel_r_reg/P0001 ,
		_w5446_
	);
	LUT4 #(
		.INIT('h4c5f)
	) name3697 (
		_w5325_,
		_w5326_,
		_w5365_,
		_w5446_,
		_w5447_
	);
	LUT2 #(
		.INIT('h8)
	) name3698 (
		\sram_data_i[9]_pad ,
		\u1_u2_dtmp_sel_r_reg/P0001 ,
		_w5448_
	);
	LUT2 #(
		.INIT('hd)
	) name3699 (
		_w5447_,
		_w5448_,
		_w5449_
	);
	LUT2 #(
		.INIT('h1)
	) name3700 (
		\u1_u2_adr_cb_reg[0]/NET0131 ,
		\u1_u2_adr_cb_reg[1]/NET0131 ,
		_w5450_
	);
	LUT3 #(
		.INIT('h10)
	) name3701 (
		\u1_u2_adr_cb_reg[0]/NET0131 ,
		\u1_u2_adr_cb_reg[1]/NET0131 ,
		\u1_u2_rx_data_valid_r_reg/NET0131 ,
		_w5451_
	);
	LUT2 #(
		.INIT('h2)
	) name3702 (
		\u1_u2_dtmp_r_reg[0]/P0001 ,
		\u1_u2_dtmp_sel_r_reg/P0001 ,
		_w5452_
	);
	LUT4 #(
		.INIT('h203f)
	) name3703 (
		\u1_u2_rx_data_valid_r_reg/NET0131 ,
		_w5360_,
		_w5450_,
		_w5452_,
		_w5453_
	);
	LUT2 #(
		.INIT('h8)
	) name3704 (
		\sram_data_i[0]_pad ,
		\u1_u2_dtmp_sel_r_reg/P0001 ,
		_w5454_
	);
	LUT2 #(
		.INIT('hd)
	) name3705 (
		_w5453_,
		_w5454_,
		_w5455_
	);
	LUT2 #(
		.INIT('h2)
	) name3706 (
		\u1_u2_dtmp_r_reg[1]/P0001 ,
		\u1_u2_dtmp_sel_r_reg/P0001 ,
		_w5456_
	);
	LUT4 #(
		.INIT('h203f)
	) name3707 (
		\u1_u2_rx_data_valid_r_reg/NET0131 ,
		_w5366_,
		_w5450_,
		_w5456_,
		_w5457_
	);
	LUT2 #(
		.INIT('h8)
	) name3708 (
		\sram_data_i[1]_pad ,
		\u1_u2_dtmp_sel_r_reg/P0001 ,
		_w5458_
	);
	LUT2 #(
		.INIT('hd)
	) name3709 (
		_w5457_,
		_w5458_,
		_w5459_
	);
	LUT4 #(
		.INIT('h0100)
	) name3710 (
		\u1_u2_adr_cb_reg[0]/NET0131 ,
		\u1_u2_adr_cb_reg[1]/NET0131 ,
		\u1_u2_dtmp_sel_r_reg/P0001 ,
		\u1_u2_rx_data_valid_r_reg/NET0131 ,
		_w5460_
	);
	LUT2 #(
		.INIT('h2)
	) name3711 (
		\u1_u2_dtmp_r_reg[2]/P0001 ,
		\u1_u2_dtmp_sel_r_reg/P0001 ,
		_w5461_
	);
	LUT4 #(
		.INIT('h4c5f)
	) name3712 (
		\u1_u2_rx_data_st_r_reg[2]/P0001 ,
		_w5451_,
		_w5460_,
		_w5461_,
		_w5462_
	);
	LUT2 #(
		.INIT('h8)
	) name3713 (
		\sram_data_i[2]_pad ,
		\u1_u2_dtmp_sel_r_reg/P0001 ,
		_w5463_
	);
	LUT2 #(
		.INIT('hd)
	) name3714 (
		_w5462_,
		_w5463_,
		_w5464_
	);
	LUT2 #(
		.INIT('h2)
	) name3715 (
		\u1_u2_dtmp_r_reg[3]/P0001 ,
		\u1_u2_dtmp_sel_r_reg/P0001 ,
		_w5465_
	);
	LUT4 #(
		.INIT('h4c5f)
	) name3716 (
		\u1_u2_rx_data_st_r_reg[3]/P0001 ,
		_w5451_,
		_w5460_,
		_w5465_,
		_w5466_
	);
	LUT2 #(
		.INIT('h8)
	) name3717 (
		\sram_data_i[3]_pad ,
		\u1_u2_dtmp_sel_r_reg/P0001 ,
		_w5467_
	);
	LUT2 #(
		.INIT('hd)
	) name3718 (
		_w5466_,
		_w5467_,
		_w5468_
	);
	LUT2 #(
		.INIT('h2)
	) name3719 (
		\u1_u2_dtmp_r_reg[4]/P0001 ,
		\u1_u2_dtmp_sel_r_reg/P0001 ,
		_w5469_
	);
	LUT4 #(
		.INIT('h4c5f)
	) name3720 (
		\u1_u2_rx_data_st_r_reg[4]/P0001 ,
		_w5451_,
		_w5460_,
		_w5469_,
		_w5470_
	);
	LUT2 #(
		.INIT('h8)
	) name3721 (
		\sram_data_i[4]_pad ,
		\u1_u2_dtmp_sel_r_reg/P0001 ,
		_w5471_
	);
	LUT2 #(
		.INIT('hd)
	) name3722 (
		_w5470_,
		_w5471_,
		_w5472_
	);
	LUT2 #(
		.INIT('h8)
	) name3723 (
		\u1_u2_rx_data_st_r_reg[5]/P0001 ,
		_w5460_,
		_w5473_
	);
	LUT2 #(
		.INIT('h2)
	) name3724 (
		\u1_u2_dtmp_r_reg[5]/P0001 ,
		\u1_u2_dtmp_sel_r_reg/P0001 ,
		_w5474_
	);
	LUT2 #(
		.INIT('h8)
	) name3725 (
		\sram_data_i[5]_pad ,
		\u1_u2_dtmp_sel_r_reg/P0001 ,
		_w5475_
	);
	LUT3 #(
		.INIT('h0b)
	) name3726 (
		_w5451_,
		_w5474_,
		_w5475_,
		_w5476_
	);
	LUT2 #(
		.INIT('hb)
	) name3727 (
		_w5473_,
		_w5476_,
		_w5477_
	);
	LUT2 #(
		.INIT('h8)
	) name3728 (
		\u1_u2_rx_data_st_r_reg[6]/P0001 ,
		_w5460_,
		_w5478_
	);
	LUT2 #(
		.INIT('h2)
	) name3729 (
		\u1_u2_dtmp_r_reg[6]/P0001 ,
		\u1_u2_dtmp_sel_r_reg/P0001 ,
		_w5479_
	);
	LUT2 #(
		.INIT('h8)
	) name3730 (
		\sram_data_i[6]_pad ,
		\u1_u2_dtmp_sel_r_reg/P0001 ,
		_w5480_
	);
	LUT3 #(
		.INIT('h0b)
	) name3731 (
		_w5451_,
		_w5479_,
		_w5480_,
		_w5481_
	);
	LUT2 #(
		.INIT('hb)
	) name3732 (
		_w5478_,
		_w5481_,
		_w5482_
	);
	LUT2 #(
		.INIT('h8)
	) name3733 (
		\u1_u2_rx_data_st_r_reg[7]/P0001 ,
		_w5460_,
		_w5483_
	);
	LUT2 #(
		.INIT('h2)
	) name3734 (
		\u1_u2_dtmp_r_reg[7]/P0001 ,
		\u1_u2_dtmp_sel_r_reg/P0001 ,
		_w5484_
	);
	LUT2 #(
		.INIT('h8)
	) name3735 (
		\sram_data_i[7]_pad ,
		\u1_u2_dtmp_sel_r_reg/P0001 ,
		_w5485_
	);
	LUT3 #(
		.INIT('h0b)
	) name3736 (
		_w5451_,
		_w5484_,
		_w5485_,
		_w5486_
	);
	LUT2 #(
		.INIT('hb)
	) name3737 (
		_w5483_,
		_w5486_,
		_w5487_
	);
	LUT3 #(
		.INIT('h40)
	) name3738 (
		\u1_u3_abort_reg/P0001 ,
		_w3209_,
		_w3225_,
		_w5488_
	);
	LUT3 #(
		.INIT('h51)
	) name3739 (
		\u1_u2_mack_r_reg/P0001 ,
		_w3224_,
		_w5488_,
		_w5489_
	);
	LUT3 #(
		.INIT('h02)
	) name3740 (
		\u5_state_reg[0]/P0001 ,
		\u5_state_reg[1]/P0001 ,
		\u5_state_reg[2]/P0001 ,
		_w5490_
	);
	LUT2 #(
		.INIT('h8)
	) name3741 (
		\u5_wb_req_s1_reg/P0001 ,
		\wb_addr_i[17]_pad ,
		_w5491_
	);
	LUT3 #(
		.INIT('h80)
	) name3742 (
		_w2224_,
		_w5490_,
		_w5491_,
		_w5492_
	);
	LUT4 #(
		.INIT('h0001)
	) name3743 (
		\u5_state_reg[0]/P0001 ,
		\u5_state_reg[3]/P0001 ,
		\u5_state_reg[4]/P0001 ,
		\u5_state_reg[5]/NET0131 ,
		_w5493_
	);
	LUT2 #(
		.INIT('h6)
	) name3744 (
		\u5_state_reg[1]/P0001 ,
		\u5_state_reg[2]/P0001 ,
		_w5494_
	);
	LUT3 #(
		.INIT('h40)
	) name3745 (
		\u2_wack_r_reg/P0001 ,
		_w5493_,
		_w5494_,
		_w5495_
	);
	LUT3 #(
		.INIT('h54)
	) name3746 (
		\u1_u2_word_done_r_reg/P0001 ,
		_w5492_,
		_w5495_,
		_w5496_
	);
	LUT2 #(
		.INIT('h2)
	) name3747 (
		rst_i_pad,
		\u2_wack_r_reg/P0001 ,
		_w5497_
	);
	LUT3 #(
		.INIT('h40)
	) name3748 (
		_w5489_,
		_w5496_,
		_w5497_,
		_w5498_
	);
	LUT3 #(
		.INIT('ha6)
	) name3749 (
		\u1_u3_new_sizeb_reg[4]/P0001 ,
		_w2803_,
		_w2805_,
		_w5499_
	);
	LUT4 #(
		.INIT('h45ba)
	) name3750 (
		_w3439_,
		_w3441_,
		_w3443_,
		_w5499_,
		_w5500_
	);
	LUT4 #(
		.INIT('h008e)
	) name3751 (
		\u1_u3_new_sizeb_reg[3]/P0001 ,
		_w2813_,
		_w3438_,
		_w3453_,
		_w5501_
	);
	LUT3 #(
		.INIT('ha6)
	) name3752 (
		\u1_u3_new_sizeb_reg[5]/P0001 ,
		_w2820_,
		_w2822_,
		_w5502_
	);
	LUT2 #(
		.INIT('h1)
	) name3753 (
		_w3448_,
		_w5502_,
		_w5503_
	);
	LUT4 #(
		.INIT('h4f00)
	) name3754 (
		_w3441_,
		_w3443_,
		_w5501_,
		_w5503_,
		_w5504_
	);
	LUT2 #(
		.INIT('h8)
	) name3755 (
		_w3448_,
		_w5502_,
		_w5505_
	);
	LUT2 #(
		.INIT('h4)
	) name3756 (
		_w3453_,
		_w5502_,
		_w5506_
	);
	LUT4 #(
		.INIT('h4500)
	) name3757 (
		_w3439_,
		_w3441_,
		_w3443_,
		_w5506_,
		_w5507_
	);
	LUT3 #(
		.INIT('hfe)
	) name3758 (
		_w5504_,
		_w5505_,
		_w5507_,
		_w5508_
	);
	LUT3 #(
		.INIT('ha6)
	) name3759 (
		\u1_u3_new_sizeb_reg[6]/P0001 ,
		_w2860_,
		_w2862_,
		_w5509_
	);
	LUT3 #(
		.INIT('h10)
	) name3760 (
		_w3447_,
		_w3448_,
		_w5509_,
		_w5510_
	);
	LUT4 #(
		.INIT('hba00)
	) name3761 (
		_w3439_,
		_w3441_,
		_w3443_,
		_w5510_,
		_w5511_
	);
	LUT4 #(
		.INIT('h45ff)
	) name3762 (
		_w3439_,
		_w3441_,
		_w3443_,
		_w3449_,
		_w5512_
	);
	LUT4 #(
		.INIT('h090b)
	) name3763 (
		_w3454_,
		_w5509_,
		_w5511_,
		_w5512_,
		_w5513_
	);
	LUT4 #(
		.INIT('h0107)
	) name3764 (
		\u1_u3_new_sizeb_reg[5]/P0001 ,
		_w2823_,
		_w3445_,
		_w3448_,
		_w5514_
	);
	LUT3 #(
		.INIT('ha6)
	) name3765 (
		\u1_u3_new_sizeb_reg[7]/P0001 ,
		_w2830_,
		_w2832_,
		_w5515_
	);
	LUT4 #(
		.INIT('h45ba)
	) name3766 (
		_w3461_,
		_w3506_,
		_w5514_,
		_w5515_,
		_w5516_
	);
	LUT3 #(
		.INIT('h08)
	) name3767 (
		rst_i_pad,
		\u5_state_reg[2]/P0001 ,
		\u5_wb_req_s1_reg/P0001 ,
		_w5517_
	);
	LUT4 #(
		.INIT('h0080)
	) name3768 (
		rst_i_pad,
		\u5_wb_req_s1_reg/P0001 ,
		\wb_addr_i[17]_pad ,
		wb_we_i_pad,
		_w5518_
	);
	LUT4 #(
		.INIT('h8880)
	) name3769 (
		_w2224_,
		_w5490_,
		_w5517_,
		_w5518_,
		_w5519_
	);
	LUT2 #(
		.INIT('h4)
	) name3770 (
		\u1_u2_word_done_r_reg/P0001 ,
		\u2_wack_r_reg/P0001 ,
		_w5520_
	);
	LUT3 #(
		.INIT('h20)
	) name3771 (
		rst_i_pad,
		\u5_state_reg[1]/P0001 ,
		\u5_state_reg[2]/P0001 ,
		_w5521_
	);
	LUT3 #(
		.INIT('h20)
	) name3772 (
		_w5493_,
		_w5520_,
		_w5521_,
		_w5522_
	);
	LUT3 #(
		.INIT('h40)
	) name3773 (
		\u1_u2_mack_r_reg/P0001 ,
		_w5493_,
		_w5521_,
		_w5523_
	);
	LUT4 #(
		.INIT('h020f)
	) name3774 (
		_w3224_,
		_w5488_,
		_w5522_,
		_w5523_,
		_w5524_
	);
	LUT2 #(
		.INIT('hb)
	) name3775 (
		_w5519_,
		_w5524_,
		_w5525_
	);
	LUT2 #(
		.INIT('h9)
	) name3776 (
		\u4_u3_csr0_reg[9]/P0001 ,
		\u4_u3_dma_in_cnt_reg[7]/P0001 ,
		_w5526_
	);
	LUT4 #(
		.INIT('h31c4)
	) name3777 (
		\u4_u3_csr0_reg[8]/P0001 ,
		\u4_u3_csr0_reg[9]/P0001 ,
		\u4_u3_dma_in_cnt_reg[6]/P0001 ,
		\u4_u3_dma_in_cnt_reg[7]/P0001 ,
		_w5527_
	);
	LUT4 #(
		.INIT('h40f0)
	) name3778 (
		_w4390_,
		_w4393_,
		_w4569_,
		_w5527_,
		_w5528_
	);
	LUT4 #(
		.INIT('hd000)
	) name3779 (
		_w4387_,
		_w4391_,
		_w4392_,
		_w5526_,
		_w5529_
	);
	LUT4 #(
		.INIT('hb777)
	) name3780 (
		\u4_u3_dma_in_cnt_reg[7]/P0001 ,
		\u4_u3_r5_reg/NET0131 ,
		_w4398_,
		_w4399_,
		_w5530_
	);
	LUT4 #(
		.INIT('h0802)
	) name3781 (
		\u4_u3_csr0_reg[8]/P0001 ,
		\u4_u3_csr0_reg[9]/P0001 ,
		\u4_u3_dma_in_cnt_reg[6]/P0001 ,
		\u4_u3_dma_in_cnt_reg[7]/P0001 ,
		_w5531_
	);
	LUT4 #(
		.INIT('h00b0)
	) name3782 (
		_w4390_,
		_w5529_,
		_w5530_,
		_w5531_,
		_w5532_
	);
	LUT4 #(
		.INIT('h0001)
	) name3783 (
		\u1_u3_buf0_rl_reg/P0001 ,
		\u1_u3_buf0_set_reg/P0001 ,
		\u4_u3_dma_in_cnt_reg[7]/P0001 ,
		\u4_u3_set_r_reg/P0001 ,
		_w5533_
	);
	LUT3 #(
		.INIT('h0e)
	) name3784 (
		\u4_u3_dma_in_cnt_reg[7]/P0001 ,
		\u4_u3_ep_match_r_reg/P0001 ,
		\u4_u3_r5_reg/NET0131 ,
		_w5534_
	);
	LUT2 #(
		.INIT('h4)
	) name3785 (
		_w5533_,
		_w5534_,
		_w5535_
	);
	LUT3 #(
		.INIT('ha2)
	) name3786 (
		\u4_u3_csr1_reg[0]/P0001 ,
		_w5530_,
		_w5535_,
		_w5536_
	);
	LUT3 #(
		.INIT('h70)
	) name3787 (
		_w5528_,
		_w5532_,
		_w5536_,
		_w5537_
	);
	LUT2 #(
		.INIT('h9)
	) name3788 (
		\u4_u0_csr0_reg[9]/P0001 ,
		\u4_u0_dma_in_cnt_reg[7]/P0001 ,
		_w5538_
	);
	LUT4 #(
		.INIT('hd000)
	) name3789 (
		_w4419_,
		_w4423_,
		_w4424_,
		_w5538_,
		_w5539_
	);
	LUT4 #(
		.INIT('hb777)
	) name3790 (
		\u4_u0_dma_in_cnt_reg[7]/P0001 ,
		\u4_u0_r5_reg/NET0131 ,
		_w4430_,
		_w4431_,
		_w5540_
	);
	LUT4 #(
		.INIT('h0802)
	) name3791 (
		\u4_u0_csr0_reg[8]/P0001 ,
		\u4_u0_csr0_reg[9]/P0001 ,
		\u4_u0_dma_in_cnt_reg[6]/P0001 ,
		\u4_u0_dma_in_cnt_reg[7]/P0001 ,
		_w5541_
	);
	LUT4 #(
		.INIT('h00b0)
	) name3792 (
		_w4422_,
		_w5539_,
		_w5540_,
		_w5541_,
		_w5542_
	);
	LUT4 #(
		.INIT('h31c4)
	) name3793 (
		\u4_u0_csr0_reg[8]/P0001 ,
		\u4_u0_csr0_reg[9]/P0001 ,
		\u4_u0_dma_in_cnt_reg[6]/P0001 ,
		\u4_u0_dma_in_cnt_reg[7]/P0001 ,
		_w5543_
	);
	LUT4 #(
		.INIT('h40f0)
	) name3794 (
		_w4422_,
		_w4425_,
		_w4592_,
		_w5543_,
		_w5544_
	);
	LUT4 #(
		.INIT('h0001)
	) name3795 (
		\u1_u3_buf0_rl_reg/P0001 ,
		\u1_u3_buf0_set_reg/P0001 ,
		\u4_u0_dma_in_cnt_reg[7]/P0001 ,
		\u4_u0_set_r_reg/P0001 ,
		_w5545_
	);
	LUT3 #(
		.INIT('h0e)
	) name3796 (
		\u4_u0_dma_in_cnt_reg[7]/P0001 ,
		\u4_u0_ep_match_r_reg/P0001 ,
		\u4_u0_r5_reg/NET0131 ,
		_w5546_
	);
	LUT2 #(
		.INIT('h4)
	) name3797 (
		_w5545_,
		_w5546_,
		_w5547_
	);
	LUT3 #(
		.INIT('ha2)
	) name3798 (
		\u4_u0_csr1_reg[0]/P0001 ,
		_w5540_,
		_w5547_,
		_w5548_
	);
	LUT3 #(
		.INIT('h70)
	) name3799 (
		_w5542_,
		_w5544_,
		_w5548_,
		_w5549_
	);
	LUT4 #(
		.INIT('h8c23)
	) name3800 (
		\u4_u1_csr0_reg[8]/P0001 ,
		\u4_u1_csr0_reg[9]/P0001 ,
		\u4_u1_dma_in_cnt_reg[6]/P0001 ,
		\u4_u1_dma_in_cnt_reg[7]/P0001 ,
		_w5550_
	);
	LUT4 #(
		.INIT('h31c4)
	) name3801 (
		\u4_u1_csr0_reg[8]/P0001 ,
		\u4_u1_csr0_reg[9]/P0001 ,
		\u4_u1_dma_in_cnt_reg[6]/P0001 ,
		\u4_u1_dma_in_cnt_reg[7]/P0001 ,
		_w5551_
	);
	LUT2 #(
		.INIT('h4)
	) name3802 (
		_w4460_,
		_w5551_,
		_w5552_
	);
	LUT4 #(
		.INIT('hef00)
	) name3803 (
		_w4463_,
		_w4468_,
		_w4469_,
		_w5552_,
		_w5553_
	);
	LUT4 #(
		.INIT('h1040)
	) name3804 (
		\u4_u1_csr0_reg[8]/P0001 ,
		\u4_u1_csr0_reg[9]/P0001 ,
		\u4_u1_dma_in_cnt_reg[6]/P0001 ,
		\u4_u1_dma_in_cnt_reg[7]/P0001 ,
		_w5554_
	);
	LUT2 #(
		.INIT('h2)
	) name3805 (
		_w4454_,
		_w5554_,
		_w5555_
	);
	LUT4 #(
		.INIT('hb777)
	) name3806 (
		\u4_u1_dma_in_cnt_reg[7]/P0001 ,
		\u4_u1_r5_reg/NET0131 ,
		_w4447_,
		_w4448_,
		_w5556_
	);
	LUT2 #(
		.INIT('h8)
	) name3807 (
		_w5555_,
		_w5556_,
		_w5557_
	);
	LUT4 #(
		.INIT('h0b00)
	) name3808 (
		_w4605_,
		_w5550_,
		_w5553_,
		_w5557_,
		_w5558_
	);
	LUT4 #(
		.INIT('h0001)
	) name3809 (
		\u1_u3_buf0_rl_reg/P0001 ,
		\u1_u3_buf0_set_reg/P0001 ,
		\u4_u1_dma_in_cnt_reg[7]/P0001 ,
		\u4_u1_set_r_reg/P0001 ,
		_w5559_
	);
	LUT3 #(
		.INIT('h0e)
	) name3810 (
		\u4_u1_dma_in_cnt_reg[7]/P0001 ,
		\u4_u1_ep_match_r_reg/P0001 ,
		\u4_u1_r5_reg/NET0131 ,
		_w5560_
	);
	LUT2 #(
		.INIT('h4)
	) name3811 (
		_w5559_,
		_w5560_,
		_w5561_
	);
	LUT3 #(
		.INIT('ha2)
	) name3812 (
		\u4_u1_csr1_reg[0]/P0001 ,
		_w5556_,
		_w5561_,
		_w5562_
	);
	LUT2 #(
		.INIT('h4)
	) name3813 (
		_w5558_,
		_w5562_,
		_w5563_
	);
	LUT4 #(
		.INIT('hf531)
	) name3814 (
		\u4_u2_csr0_reg[7]/P0001 ,
		\u4_u2_csr0_reg[8]/P0001 ,
		\u4_u2_dma_in_cnt_reg[5]/P0001 ,
		\u4_u2_dma_in_cnt_reg[6]/P0001 ,
		_w5564_
	);
	LUT4 #(
		.INIT('hef00)
	) name3815 (
		_w4491_,
		_w4496_,
		_w4497_,
		_w5564_,
		_w5565_
	);
	LUT4 #(
		.INIT('h8c23)
	) name3816 (
		\u4_u2_csr0_reg[8]/P0001 ,
		\u4_u2_csr0_reg[9]/P0001 ,
		\u4_u2_dma_in_cnt_reg[6]/P0001 ,
		\u4_u2_dma_in_cnt_reg[7]/P0001 ,
		_w5566_
	);
	LUT4 #(
		.INIT('h31c4)
	) name3817 (
		\u4_u2_csr0_reg[8]/P0001 ,
		\u4_u2_csr0_reg[9]/P0001 ,
		\u4_u2_dma_in_cnt_reg[6]/P0001 ,
		\u4_u2_dma_in_cnt_reg[7]/P0001 ,
		_w5567_
	);
	LUT2 #(
		.INIT('h4)
	) name3818 (
		_w4488_,
		_w5567_,
		_w5568_
	);
	LUT4 #(
		.INIT('hef00)
	) name3819 (
		_w4491_,
		_w4496_,
		_w4497_,
		_w5568_,
		_w5569_
	);
	LUT4 #(
		.INIT('h1040)
	) name3820 (
		\u4_u2_csr0_reg[8]/P0001 ,
		\u4_u2_csr0_reg[9]/P0001 ,
		\u4_u2_dma_in_cnt_reg[6]/P0001 ,
		\u4_u2_dma_in_cnt_reg[7]/P0001 ,
		_w5570_
	);
	LUT2 #(
		.INIT('h2)
	) name3821 (
		_w4610_,
		_w5570_,
		_w5571_
	);
	LUT4 #(
		.INIT('hb777)
	) name3822 (
		\u4_u2_dma_in_cnt_reg[7]/P0001 ,
		\u4_u2_r5_reg/NET0131 ,
		_w4504_,
		_w4505_,
		_w5572_
	);
	LUT2 #(
		.INIT('h8)
	) name3823 (
		_w5571_,
		_w5572_,
		_w5573_
	);
	LUT4 #(
		.INIT('h0b00)
	) name3824 (
		_w5565_,
		_w5566_,
		_w5569_,
		_w5573_,
		_w5574_
	);
	LUT4 #(
		.INIT('h0001)
	) name3825 (
		\u1_u3_buf0_rl_reg/P0001 ,
		\u1_u3_buf0_set_reg/P0001 ,
		\u4_u2_dma_in_cnt_reg[7]/P0001 ,
		\u4_u2_set_r_reg/P0001 ,
		_w5575_
	);
	LUT3 #(
		.INIT('h0e)
	) name3826 (
		\u4_u2_dma_in_cnt_reg[7]/P0001 ,
		\u4_u2_ep_match_r_reg/P0001 ,
		\u4_u2_r5_reg/NET0131 ,
		_w5576_
	);
	LUT2 #(
		.INIT('h4)
	) name3827 (
		_w5575_,
		_w5576_,
		_w5577_
	);
	LUT3 #(
		.INIT('ha2)
	) name3828 (
		\u4_u2_csr1_reg[0]/P0001 ,
		_w5572_,
		_w5577_,
		_w5578_
	);
	LUT2 #(
		.INIT('h4)
	) name3829 (
		_w5574_,
		_w5578_,
		_w5579_
	);
	LUT3 #(
		.INIT('h20)
	) name3830 (
		\u4_u3_csr1_reg[0]/P0001 ,
		\u4_u3_dma_out_cnt_reg[7]/P0001 ,
		\u4_u3_r5_reg/NET0131 ,
		_w5580_
	);
	LUT3 #(
		.INIT('h80)
	) name3831 (
		\u4_u3_csr1_reg[0]/P0001 ,
		\u4_u3_dma_out_cnt_reg[7]/P0001 ,
		\u4_u3_r5_reg/NET0131 ,
		_w5581_
	);
	LUT4 #(
		.INIT('h087f)
	) name3832 (
		_w4650_,
		_w4652_,
		_w5580_,
		_w5581_,
		_w5582_
	);
	LUT4 #(
		.INIT('h135f)
	) name3833 (
		\u4_u3_csr0_reg[7]/P0001 ,
		\u4_u3_csr0_reg[8]/P0001 ,
		\u4_u3_dma_out_cnt_reg[5]/P0001 ,
		\u4_u3_dma_out_cnt_reg[6]/P0001 ,
		_w5583_
	);
	LUT4 #(
		.INIT('hef00)
	) name3834 (
		_w4667_,
		_w4672_,
		_w4674_,
		_w5583_,
		_w5584_
	);
	LUT4 #(
		.INIT('hc832)
	) name3835 (
		\u4_u3_csr0_reg[8]/P0001 ,
		\u4_u3_csr0_reg[9]/P0001 ,
		\u4_u3_dma_out_cnt_reg[6]/P0001 ,
		\u4_u3_dma_out_cnt_reg[7]/P0001 ,
		_w5585_
	);
	LUT2 #(
		.INIT('h4)
	) name3836 (
		_w5584_,
		_w5585_,
		_w5586_
	);
	LUT4 #(
		.INIT('h134c)
	) name3837 (
		\u4_u3_csr0_reg[8]/P0001 ,
		\u4_u3_csr0_reg[9]/P0001 ,
		\u4_u3_dma_out_cnt_reg[6]/P0001 ,
		\u4_u3_dma_out_cnt_reg[7]/P0001 ,
		_w5587_
	);
	LUT3 #(
		.INIT('h2a)
	) name3838 (
		_w4569_,
		_w4676_,
		_w5587_,
		_w5588_
	);
	LUT4 #(
		.INIT('h0001)
	) name3839 (
		\u1_u3_buf0_rl_reg/P0001 ,
		\u1_u3_buf0_set_reg/P0001 ,
		\u4_u3_dma_out_cnt_reg[7]/P0001 ,
		\u4_u3_set_r_reg/P0001 ,
		_w5589_
	);
	LUT3 #(
		.INIT('ha8)
	) name3840 (
		\u4_u3_csr1_reg[0]/P0001 ,
		\u4_u3_dma_out_cnt_reg[7]/P0001 ,
		\u4_u3_ep_match_r_reg/P0001 ,
		_w5590_
	);
	LUT3 #(
		.INIT('h10)
	) name3841 (
		\u4_u3_r5_reg/NET0131 ,
		_w5589_,
		_w5590_,
		_w5591_
	);
	LUT4 #(
		.INIT('hdf55)
	) name3842 (
		_w5582_,
		_w5586_,
		_w5588_,
		_w5591_,
		_w5592_
	);
	LUT3 #(
		.INIT('h20)
	) name3843 (
		\u4_u0_csr1_reg[0]/P0001 ,
		\u4_u0_dma_out_cnt_reg[7]/P0001 ,
		\u4_u0_r5_reg/NET0131 ,
		_w5593_
	);
	LUT3 #(
		.INIT('h80)
	) name3844 (
		\u4_u0_csr1_reg[0]/P0001 ,
		\u4_u0_dma_out_cnt_reg[7]/P0001 ,
		\u4_u0_r5_reg/NET0131 ,
		_w5594_
	);
	LUT4 #(
		.INIT('h087f)
	) name3845 (
		_w4681_,
		_w4683_,
		_w5593_,
		_w5594_,
		_w5595_
	);
	LUT4 #(
		.INIT('h134c)
	) name3846 (
		\u4_u0_csr0_reg[8]/P0001 ,
		\u4_u0_csr0_reg[9]/P0001 ,
		\u4_u0_dma_out_cnt_reg[6]/P0001 ,
		\u4_u0_dma_out_cnt_reg[7]/P0001 ,
		_w5596_
	);
	LUT4 #(
		.INIT('h135f)
	) name3847 (
		\u4_u0_csr0_reg[7]/P0001 ,
		\u4_u0_csr0_reg[8]/P0001 ,
		\u4_u0_dma_out_cnt_reg[5]/P0001 ,
		\u4_u0_dma_out_cnt_reg[6]/P0001 ,
		_w5597_
	);
	LUT4 #(
		.INIT('hef00)
	) name3848 (
		_w4697_,
		_w4702_,
		_w4704_,
		_w5597_,
		_w5598_
	);
	LUT4 #(
		.INIT('hc832)
	) name3849 (
		\u4_u0_csr0_reg[8]/P0001 ,
		\u4_u0_csr0_reg[9]/P0001 ,
		\u4_u0_dma_out_cnt_reg[6]/P0001 ,
		\u4_u0_dma_out_cnt_reg[7]/P0001 ,
		_w5599_
	);
	LUT4 #(
		.INIT('h7077)
	) name3850 (
		_w4706_,
		_w5596_,
		_w5598_,
		_w5599_,
		_w5600_
	);
	LUT4 #(
		.INIT('h0001)
	) name3851 (
		\u1_u3_buf0_rl_reg/P0001 ,
		\u1_u3_buf0_set_reg/P0001 ,
		\u4_u0_dma_out_cnt_reg[7]/P0001 ,
		\u4_u0_set_r_reg/P0001 ,
		_w5601_
	);
	LUT3 #(
		.INIT('ha8)
	) name3852 (
		\u4_u0_csr1_reg[0]/P0001 ,
		\u4_u0_dma_out_cnt_reg[7]/P0001 ,
		\u4_u0_ep_match_r_reg/P0001 ,
		_w5602_
	);
	LUT3 #(
		.INIT('h10)
	) name3853 (
		\u4_u0_r5_reg/NET0131 ,
		_w5601_,
		_w5602_,
		_w5603_
	);
	LUT4 #(
		.INIT('h7f33)
	) name3854 (
		_w4592_,
		_w5595_,
		_w5600_,
		_w5603_,
		_w5604_
	);
	LUT3 #(
		.INIT('h20)
	) name3855 (
		\u4_u1_csr1_reg[0]/P0001 ,
		\u4_u1_dma_out_cnt_reg[7]/P0001 ,
		\u4_u1_r5_reg/NET0131 ,
		_w5605_
	);
	LUT3 #(
		.INIT('h80)
	) name3856 (
		\u4_u1_csr1_reg[0]/P0001 ,
		\u4_u1_dma_out_cnt_reg[7]/P0001 ,
		\u4_u1_r5_reg/NET0131 ,
		_w5606_
	);
	LUT4 #(
		.INIT('h087f)
	) name3857 (
		_w4711_,
		_w4713_,
		_w5605_,
		_w5606_,
		_w5607_
	);
	LUT4 #(
		.INIT('h134c)
	) name3858 (
		\u4_u1_csr0_reg[8]/P0001 ,
		\u4_u1_csr0_reg[9]/P0001 ,
		\u4_u1_dma_out_cnt_reg[6]/P0001 ,
		\u4_u1_dma_out_cnt_reg[7]/P0001 ,
		_w5608_
	);
	LUT4 #(
		.INIT('h135f)
	) name3859 (
		\u4_u1_csr0_reg[7]/P0001 ,
		\u4_u1_csr0_reg[8]/P0001 ,
		\u4_u1_dma_out_cnt_reg[5]/P0001 ,
		\u4_u1_dma_out_cnt_reg[6]/P0001 ,
		_w5609_
	);
	LUT4 #(
		.INIT('hef00)
	) name3860 (
		_w4728_,
		_w4733_,
		_w4735_,
		_w5609_,
		_w5610_
	);
	LUT4 #(
		.INIT('hc832)
	) name3861 (
		\u4_u1_csr0_reg[8]/P0001 ,
		\u4_u1_csr0_reg[9]/P0001 ,
		\u4_u1_dma_out_cnt_reg[6]/P0001 ,
		\u4_u1_dma_out_cnt_reg[7]/P0001 ,
		_w5611_
	);
	LUT4 #(
		.INIT('h7077)
	) name3862 (
		_w4737_,
		_w5608_,
		_w5610_,
		_w5611_,
		_w5612_
	);
	LUT4 #(
		.INIT('h0001)
	) name3863 (
		\u1_u3_buf0_rl_reg/P0001 ,
		\u1_u3_buf0_set_reg/P0001 ,
		\u4_u1_dma_out_cnt_reg[7]/P0001 ,
		\u4_u1_set_r_reg/P0001 ,
		_w5613_
	);
	LUT3 #(
		.INIT('ha8)
	) name3864 (
		\u4_u1_csr1_reg[0]/P0001 ,
		\u4_u1_dma_out_cnt_reg[7]/P0001 ,
		\u4_u1_ep_match_r_reg/P0001 ,
		_w5614_
	);
	LUT3 #(
		.INIT('h10)
	) name3865 (
		\u4_u1_r5_reg/NET0131 ,
		_w5613_,
		_w5614_,
		_w5615_
	);
	LUT4 #(
		.INIT('h7f33)
	) name3866 (
		_w4454_,
		_w5607_,
		_w5612_,
		_w5615_,
		_w5616_
	);
	LUT3 #(
		.INIT('h20)
	) name3867 (
		\u4_u2_csr1_reg[0]/P0001 ,
		\u4_u2_dma_out_cnt_reg[7]/P0001 ,
		\u4_u2_r5_reg/NET0131 ,
		_w5617_
	);
	LUT3 #(
		.INIT('h80)
	) name3868 (
		\u4_u2_csr1_reg[0]/P0001 ,
		\u4_u2_dma_out_cnt_reg[7]/P0001 ,
		\u4_u2_r5_reg/NET0131 ,
		_w5618_
	);
	LUT4 #(
		.INIT('h087f)
	) name3869 (
		_w4742_,
		_w4744_,
		_w5617_,
		_w5618_,
		_w5619_
	);
	LUT4 #(
		.INIT('h135f)
	) name3870 (
		\u4_u2_csr0_reg[7]/P0001 ,
		\u4_u2_csr0_reg[8]/P0001 ,
		\u4_u2_dma_out_cnt_reg[5]/P0001 ,
		\u4_u2_dma_out_cnt_reg[6]/P0001 ,
		_w5620_
	);
	LUT4 #(
		.INIT('hef00)
	) name3871 (
		_w4758_,
		_w4763_,
		_w4765_,
		_w5620_,
		_w5621_
	);
	LUT4 #(
		.INIT('hc832)
	) name3872 (
		\u4_u2_csr0_reg[8]/P0001 ,
		\u4_u2_csr0_reg[9]/P0001 ,
		\u4_u2_dma_out_cnt_reg[6]/P0001 ,
		\u4_u2_dma_out_cnt_reg[7]/P0001 ,
		_w5622_
	);
	LUT2 #(
		.INIT('h4)
	) name3873 (
		_w5621_,
		_w5622_,
		_w5623_
	);
	LUT4 #(
		.INIT('h134c)
	) name3874 (
		\u4_u2_csr0_reg[8]/P0001 ,
		\u4_u2_csr0_reg[9]/P0001 ,
		\u4_u2_dma_out_cnt_reg[6]/P0001 ,
		\u4_u2_dma_out_cnt_reg[7]/P0001 ,
		_w5624_
	);
	LUT3 #(
		.INIT('h2a)
	) name3875 (
		_w4610_,
		_w4767_,
		_w5624_,
		_w5625_
	);
	LUT4 #(
		.INIT('h0001)
	) name3876 (
		\u1_u3_buf0_rl_reg/P0001 ,
		\u1_u3_buf0_set_reg/P0001 ,
		\u4_u2_dma_out_cnt_reg[7]/P0001 ,
		\u4_u2_set_r_reg/P0001 ,
		_w5626_
	);
	LUT3 #(
		.INIT('ha8)
	) name3877 (
		\u4_u2_csr1_reg[0]/P0001 ,
		\u4_u2_dma_out_cnt_reg[7]/P0001 ,
		\u4_u2_ep_match_r_reg/P0001 ,
		_w5627_
	);
	LUT3 #(
		.INIT('h10)
	) name3878 (
		\u4_u2_r5_reg/NET0131 ,
		_w5626_,
		_w5627_,
		_w5628_
	);
	LUT4 #(
		.INIT('hdf55)
	) name3879 (
		_w5619_,
		_w5623_,
		_w5625_,
		_w5628_,
		_w5629_
	);
	LUT4 #(
		.INIT('h5450)
	) name3880 (
		\u4_u3_r5_reg/NET0131 ,
		_w4676_,
		_w4951_,
		_w4952_,
		_w5630_
	);
	LUT2 #(
		.INIT('h2)
	) name3881 (
		\u4_u3_ep_match_r_reg/P0001 ,
		\u4_u3_r5_reg/NET0131 ,
		_w5631_
	);
	LUT2 #(
		.INIT('h4)
	) name3882 (
		_w4402_,
		_w5631_,
		_w5632_
	);
	LUT4 #(
		.INIT('h8000)
	) name3883 (
		\u4_u3_r5_reg/NET0131 ,
		_w4652_,
		_w4953_,
		_w4954_,
		_w5633_
	);
	LUT3 #(
		.INIT('ha8)
	) name3884 (
		\u4_u3_dma_out_cnt_reg[10]/P0001 ,
		_w5632_,
		_w5633_,
		_w5634_
	);
	LUT2 #(
		.INIT('h1)
	) name3885 (
		\u4_u3_dma_out_cnt_reg[10]/P0001 ,
		\u4_u3_r5_reg/NET0131 ,
		_w5635_
	);
	LUT4 #(
		.INIT('hec00)
	) name3886 (
		_w4676_,
		_w4951_,
		_w4952_,
		_w5635_,
		_w5636_
	);
	LUT3 #(
		.INIT('h45)
	) name3887 (
		\u4_u3_dma_out_cnt_reg[10]/P0001 ,
		_w4402_,
		_w5631_,
		_w5637_
	);
	LUT3 #(
		.INIT('h8a)
	) name3888 (
		\u4_u3_csr1_reg[0]/P0001 ,
		_w5633_,
		_w5637_,
		_w5638_
	);
	LUT4 #(
		.INIT('h0b00)
	) name3889 (
		_w5630_,
		_w5634_,
		_w5636_,
		_w5638_,
		_w5639_
	);
	LUT4 #(
		.INIT('h5450)
	) name3890 (
		\u4_u0_r5_reg/NET0131 ,
		_w4706_,
		_w4981_,
		_w4982_,
		_w5640_
	);
	LUT2 #(
		.INIT('h2)
	) name3891 (
		\u4_u0_ep_match_r_reg/P0001 ,
		\u4_u0_r5_reg/NET0131 ,
		_w5641_
	);
	LUT2 #(
		.INIT('h4)
	) name3892 (
		_w4434_,
		_w5641_,
		_w5642_
	);
	LUT4 #(
		.INIT('h8000)
	) name3893 (
		\u4_u0_r5_reg/NET0131 ,
		_w4683_,
		_w4983_,
		_w4984_,
		_w5643_
	);
	LUT3 #(
		.INIT('ha8)
	) name3894 (
		\u4_u0_dma_out_cnt_reg[10]/P0001 ,
		_w5642_,
		_w5643_,
		_w5644_
	);
	LUT2 #(
		.INIT('h1)
	) name3895 (
		\u4_u0_dma_out_cnt_reg[10]/P0001 ,
		\u4_u0_r5_reg/NET0131 ,
		_w5645_
	);
	LUT4 #(
		.INIT('hec00)
	) name3896 (
		_w4706_,
		_w4981_,
		_w4982_,
		_w5645_,
		_w5646_
	);
	LUT3 #(
		.INIT('h45)
	) name3897 (
		\u4_u0_dma_out_cnt_reg[10]/P0001 ,
		_w4434_,
		_w5641_,
		_w5647_
	);
	LUT3 #(
		.INIT('h8a)
	) name3898 (
		\u4_u0_csr1_reg[0]/P0001 ,
		_w5643_,
		_w5647_,
		_w5648_
	);
	LUT4 #(
		.INIT('h0b00)
	) name3899 (
		_w5640_,
		_w5644_,
		_w5646_,
		_w5648_,
		_w5649_
	);
	LUT4 #(
		.INIT('h5450)
	) name3900 (
		\u4_u1_r5_reg/NET0131 ,
		_w4737_,
		_w5015_,
		_w5016_,
		_w5650_
	);
	LUT2 #(
		.INIT('h2)
	) name3901 (
		\u4_u1_ep_match_r_reg/P0001 ,
		\u4_u1_r5_reg/NET0131 ,
		_w5651_
	);
	LUT2 #(
		.INIT('h4)
	) name3902 (
		_w4453_,
		_w5651_,
		_w5652_
	);
	LUT4 #(
		.INIT('h8000)
	) name3903 (
		\u4_u1_r5_reg/NET0131 ,
		_w4713_,
		_w5017_,
		_w5018_,
		_w5653_
	);
	LUT3 #(
		.INIT('ha8)
	) name3904 (
		\u4_u1_dma_out_cnt_reg[10]/P0001 ,
		_w5652_,
		_w5653_,
		_w5654_
	);
	LUT2 #(
		.INIT('h1)
	) name3905 (
		\u4_u1_dma_out_cnt_reg[10]/P0001 ,
		\u4_u1_r5_reg/NET0131 ,
		_w5655_
	);
	LUT4 #(
		.INIT('hec00)
	) name3906 (
		_w4737_,
		_w5015_,
		_w5016_,
		_w5655_,
		_w5656_
	);
	LUT3 #(
		.INIT('h45)
	) name3907 (
		\u4_u1_dma_out_cnt_reg[10]/P0001 ,
		_w4453_,
		_w5651_,
		_w5657_
	);
	LUT3 #(
		.INIT('h8a)
	) name3908 (
		\u4_u1_csr1_reg[0]/P0001 ,
		_w5653_,
		_w5657_,
		_w5658_
	);
	LUT4 #(
		.INIT('h0b00)
	) name3909 (
		_w5650_,
		_w5654_,
		_w5656_,
		_w5658_,
		_w5659_
	);
	LUT4 #(
		.INIT('h007f)
	) name3910 (
		\u4_u2_csr0_reg[10]/P0001 ,
		\u4_u2_dma_out_cnt_reg[8]/P0001 ,
		\u4_u2_dma_out_cnt_reg[9]/P0001 ,
		\u4_u2_r5_reg/NET0131 ,
		_w5660_
	);
	LUT4 #(
		.INIT('h8f00)
	) name3911 (
		_w4767_,
		_w4768_,
		_w5056_,
		_w5660_,
		_w5661_
	);
	LUT2 #(
		.INIT('h2)
	) name3912 (
		\u4_u2_ep_match_r_reg/P0001 ,
		\u4_u2_r5_reg/NET0131 ,
		_w5662_
	);
	LUT2 #(
		.INIT('h4)
	) name3913 (
		_w4482_,
		_w5662_,
		_w5663_
	);
	LUT4 #(
		.INIT('h8000)
	) name3914 (
		\u4_u2_r5_reg/NET0131 ,
		_w4744_,
		_w5047_,
		_w5048_,
		_w5664_
	);
	LUT3 #(
		.INIT('ha8)
	) name3915 (
		\u4_u2_dma_out_cnt_reg[10]/P0001 ,
		_w5663_,
		_w5664_,
		_w5665_
	);
	LUT2 #(
		.INIT('h1)
	) name3916 (
		\u4_u2_dma_out_cnt_reg[10]/P0001 ,
		\u4_u2_r5_reg/NET0131 ,
		_w5666_
	);
	LUT2 #(
		.INIT('h4)
	) name3917 (
		_w5057_,
		_w5666_,
		_w5667_
	);
	LUT4 #(
		.INIT('h8f00)
	) name3918 (
		_w4767_,
		_w4768_,
		_w5056_,
		_w5667_,
		_w5668_
	);
	LUT3 #(
		.INIT('h45)
	) name3919 (
		\u4_u2_dma_out_cnt_reg[10]/P0001 ,
		_w4482_,
		_w5662_,
		_w5669_
	);
	LUT3 #(
		.INIT('h8a)
	) name3920 (
		\u4_u2_csr1_reg[0]/P0001 ,
		_w5664_,
		_w5669_,
		_w5670_
	);
	LUT4 #(
		.INIT('h0b00)
	) name3921 (
		_w5661_,
		_w5665_,
		_w5668_,
		_w5670_,
		_w5671_
	);
	LUT3 #(
		.INIT('h01)
	) name3922 (
		\u5_state_reg[0]/P0001 ,
		\u5_state_reg[1]/P0001 ,
		\u5_state_reg[2]/P0001 ,
		_w5672_
	);
	LUT3 #(
		.INIT('h02)
	) name3923 (
		\u5_state_reg[3]/P0001 ,
		\u5_state_reg[4]/P0001 ,
		\u5_state_reg[5]/NET0131 ,
		_w5673_
	);
	LUT2 #(
		.INIT('h8)
	) name3924 (
		_w5672_,
		_w5673_,
		_w5674_
	);
	LUT4 #(
		.INIT('h0111)
	) name3925 (
		\u5_state_reg[4]/P0001 ,
		_w5520_,
		_w5672_,
		_w5673_,
		_w5675_
	);
	LUT4 #(
		.INIT('h0111)
	) name3926 (
		\u1_u2_mack_r_reg/P0001 ,
		\u5_state_reg[4]/P0001 ,
		_w5672_,
		_w5673_,
		_w5676_
	);
	LUT4 #(
		.INIT('h020f)
	) name3927 (
		_w3224_,
		_w5488_,
		_w5675_,
		_w5676_,
		_w5677_
	);
	LUT4 #(
		.INIT('h0777)
	) name3928 (
		_w5493_,
		_w5494_,
		_w5672_,
		_w5673_,
		_w5678_
	);
	LUT2 #(
		.INIT('h2)
	) name3929 (
		rst_i_pad,
		_w5678_,
		_w5679_
	);
	LUT2 #(
		.INIT('h8)
	) name3930 (
		_w5677_,
		_w5679_,
		_w5680_
	);
	LUT2 #(
		.INIT('h8)
	) name3931 (
		\u4_u3_dma_in_cnt_reg[4]/P0001 ,
		\u4_u3_dma_in_cnt_reg[5]/P0001 ,
		_w5681_
	);
	LUT3 #(
		.INIT('h2a)
	) name3932 (
		\u4_u3_r5_reg/NET0131 ,
		_w4399_,
		_w5681_,
		_w5682_
	);
	LUT2 #(
		.INIT('h8)
	) name3933 (
		\u4_u3_csr1_reg[0]/P0001 ,
		\u4_u3_dma_in_cnt_reg[5]/P0001 ,
		_w5683_
	);
	LUT2 #(
		.INIT('h8)
	) name3934 (
		\u4_u3_csr1_reg[0]/P0001 ,
		\u4_u3_dma_in_cnt_reg[4]/P0001 ,
		_w5684_
	);
	LUT3 #(
		.INIT('h13)
	) name3935 (
		_w4399_,
		_w5683_,
		_w5684_,
		_w5685_
	);
	LUT2 #(
		.INIT('h2)
	) name3936 (
		_w5682_,
		_w5685_,
		_w5686_
	);
	LUT4 #(
		.INIT('h7310)
	) name3937 (
		\u4_u3_csr0_reg[5]/P0001 ,
		\u4_u3_csr0_reg[6]/P0001 ,
		\u4_u3_dma_in_cnt_reg[3]/P0001 ,
		\u4_u3_dma_in_cnt_reg[4]/P0001 ,
		_w5687_
	);
	LUT4 #(
		.INIT('h0b00)
	) name3938 (
		_w4384_,
		_w4385_,
		_w4386_,
		_w4389_,
		_w5688_
	);
	LUT2 #(
		.INIT('h9)
	) name3939 (
		\u4_u3_csr0_reg[7]/P0001 ,
		\u4_u3_dma_in_cnt_reg[5]/P0001 ,
		_w5689_
	);
	LUT4 #(
		.INIT('h0001)
	) name3940 (
		\u1_u3_buf0_rl_reg/P0001 ,
		\u1_u3_buf0_set_reg/P0001 ,
		\u4_u3_dma_in_cnt_reg[5]/P0001 ,
		\u4_u3_set_r_reg/P0001 ,
		_w5690_
	);
	LUT3 #(
		.INIT('ha8)
	) name3941 (
		\u4_u3_csr1_reg[0]/P0001 ,
		\u4_u3_dma_in_cnt_reg[5]/P0001 ,
		\u4_u3_ep_match_r_reg/P0001 ,
		_w5691_
	);
	LUT4 #(
		.INIT('h0700)
	) name3942 (
		_w4569_,
		_w5689_,
		_w5690_,
		_w5691_,
		_w5692_
	);
	LUT4 #(
		.INIT('h0d00)
	) name3943 (
		_w4569_,
		_w5689_,
		_w5690_,
		_w5691_,
		_w5693_
	);
	LUT4 #(
		.INIT('h0e1f)
	) name3944 (
		_w5687_,
		_w5688_,
		_w5692_,
		_w5693_,
		_w5694_
	);
	LUT3 #(
		.INIT('hcd)
	) name3945 (
		\u4_u3_r5_reg/NET0131 ,
		_w5686_,
		_w5694_,
		_w5695_
	);
	LUT2 #(
		.INIT('h8)
	) name3946 (
		\u4_u0_dma_in_cnt_reg[4]/P0001 ,
		\u4_u0_dma_in_cnt_reg[5]/P0001 ,
		_w5696_
	);
	LUT3 #(
		.INIT('h2a)
	) name3947 (
		\u4_u0_r5_reg/NET0131 ,
		_w4431_,
		_w5696_,
		_w5697_
	);
	LUT2 #(
		.INIT('h8)
	) name3948 (
		\u4_u0_csr1_reg[0]/P0001 ,
		\u4_u0_dma_in_cnt_reg[5]/P0001 ,
		_w5698_
	);
	LUT2 #(
		.INIT('h8)
	) name3949 (
		\u4_u0_csr1_reg[0]/P0001 ,
		\u4_u0_dma_in_cnt_reg[4]/P0001 ,
		_w5699_
	);
	LUT3 #(
		.INIT('h13)
	) name3950 (
		_w4431_,
		_w5698_,
		_w5699_,
		_w5700_
	);
	LUT2 #(
		.INIT('h2)
	) name3951 (
		_w5697_,
		_w5700_,
		_w5701_
	);
	LUT4 #(
		.INIT('h7310)
	) name3952 (
		\u4_u0_csr0_reg[5]/P0001 ,
		\u4_u0_csr0_reg[6]/P0001 ,
		\u4_u0_dma_in_cnt_reg[3]/P0001 ,
		\u4_u0_dma_in_cnt_reg[4]/P0001 ,
		_w5702_
	);
	LUT4 #(
		.INIT('h0b00)
	) name3953 (
		_w4416_,
		_w4417_,
		_w4418_,
		_w4421_,
		_w5703_
	);
	LUT2 #(
		.INIT('h9)
	) name3954 (
		\u4_u0_csr0_reg[7]/P0001 ,
		\u4_u0_dma_in_cnt_reg[5]/P0001 ,
		_w5704_
	);
	LUT4 #(
		.INIT('h0001)
	) name3955 (
		\u1_u3_buf0_rl_reg/P0001 ,
		\u1_u3_buf0_set_reg/P0001 ,
		\u4_u0_dma_in_cnt_reg[5]/P0001 ,
		\u4_u0_set_r_reg/P0001 ,
		_w5705_
	);
	LUT3 #(
		.INIT('ha8)
	) name3956 (
		\u4_u0_csr1_reg[0]/P0001 ,
		\u4_u0_dma_in_cnt_reg[5]/P0001 ,
		\u4_u0_ep_match_r_reg/P0001 ,
		_w5706_
	);
	LUT4 #(
		.INIT('h0700)
	) name3957 (
		_w4592_,
		_w5704_,
		_w5705_,
		_w5706_,
		_w5707_
	);
	LUT4 #(
		.INIT('h0d00)
	) name3958 (
		_w4592_,
		_w5704_,
		_w5705_,
		_w5706_,
		_w5708_
	);
	LUT4 #(
		.INIT('h0e1f)
	) name3959 (
		_w5702_,
		_w5703_,
		_w5707_,
		_w5708_,
		_w5709_
	);
	LUT3 #(
		.INIT('hcd)
	) name3960 (
		\u4_u0_r5_reg/NET0131 ,
		_w5701_,
		_w5709_,
		_w5710_
	);
	LUT2 #(
		.INIT('h9)
	) name3961 (
		\u4_u1_csr0_reg[7]/P0001 ,
		\u4_u1_dma_in_cnt_reg[5]/P0001 ,
		_w5711_
	);
	LUT2 #(
		.INIT('h8)
	) name3962 (
		_w4454_,
		_w5711_,
		_w5712_
	);
	LUT3 #(
		.INIT('hb0)
	) name3963 (
		\u4_u1_csr0_reg[6]/P0001 ,
		\u4_u1_dma_in_cnt_reg[4]/P0001 ,
		\u4_u1_ep_match_r_reg/P0001 ,
		_w5713_
	);
	LUT2 #(
		.INIT('h4)
	) name3964 (
		_w4453_,
		_w5713_,
		_w5714_
	);
	LUT4 #(
		.INIT('h0e0f)
	) name3965 (
		_w4463_,
		_w4468_,
		_w5712_,
		_w5714_,
		_w5715_
	);
	LUT4 #(
		.INIT('h60c0)
	) name3966 (
		\u4_u1_dma_in_cnt_reg[4]/P0001 ,
		\u4_u1_dma_in_cnt_reg[5]/P0001 ,
		\u4_u1_r5_reg/NET0131 ,
		_w4448_,
		_w5716_
	);
	LUT4 #(
		.INIT('h8c23)
	) name3967 (
		\u4_u1_csr0_reg[6]/P0001 ,
		\u4_u1_csr0_reg[7]/P0001 ,
		\u4_u1_dma_in_cnt_reg[4]/P0001 ,
		\u4_u1_dma_in_cnt_reg[5]/P0001 ,
		_w5717_
	);
	LUT4 #(
		.INIT('h0e0f)
	) name3968 (
		_w4463_,
		_w4468_,
		_w5716_,
		_w5717_,
		_w5718_
	);
	LUT4 #(
		.INIT('h0001)
	) name3969 (
		\u1_u3_buf0_rl_reg/P0001 ,
		\u1_u3_buf0_set_reg/P0001 ,
		\u4_u1_dma_in_cnt_reg[5]/P0001 ,
		\u4_u1_set_r_reg/P0001 ,
		_w5719_
	);
	LUT3 #(
		.INIT('h0e)
	) name3970 (
		\u4_u1_dma_in_cnt_reg[5]/P0001 ,
		\u4_u1_ep_match_r_reg/P0001 ,
		\u4_u1_r5_reg/NET0131 ,
		_w5720_
	);
	LUT2 #(
		.INIT('h4)
	) name3971 (
		_w5719_,
		_w5720_,
		_w5721_
	);
	LUT3 #(
		.INIT('ha8)
	) name3972 (
		\u4_u1_csr1_reg[0]/P0001 ,
		_w5716_,
		_w5721_,
		_w5722_
	);
	LUT3 #(
		.INIT('hb0)
	) name3973 (
		_w5715_,
		_w5718_,
		_w5722_,
		_w5723_
	);
	LUT2 #(
		.INIT('h9)
	) name3974 (
		\u4_u2_csr0_reg[7]/P0001 ,
		\u4_u2_dma_in_cnt_reg[5]/P0001 ,
		_w5724_
	);
	LUT2 #(
		.INIT('h8)
	) name3975 (
		_w4610_,
		_w5724_,
		_w5725_
	);
	LUT3 #(
		.INIT('hb0)
	) name3976 (
		\u4_u2_csr0_reg[6]/P0001 ,
		\u4_u2_dma_in_cnt_reg[4]/P0001 ,
		\u4_u2_ep_match_r_reg/P0001 ,
		_w5726_
	);
	LUT2 #(
		.INIT('h4)
	) name3977 (
		_w4482_,
		_w5726_,
		_w5727_
	);
	LUT4 #(
		.INIT('h0e0f)
	) name3978 (
		_w4491_,
		_w4496_,
		_w5725_,
		_w5727_,
		_w5728_
	);
	LUT2 #(
		.INIT('h8)
	) name3979 (
		\u4_u2_dma_in_cnt_reg[4]/P0001 ,
		\u4_u2_dma_in_cnt_reg[5]/P0001 ,
		_w5729_
	);
	LUT4 #(
		.INIT('h60c0)
	) name3980 (
		\u4_u2_dma_in_cnt_reg[4]/P0001 ,
		\u4_u2_dma_in_cnt_reg[5]/P0001 ,
		\u4_u2_r5_reg/NET0131 ,
		_w4505_,
		_w5730_
	);
	LUT4 #(
		.INIT('h8c23)
	) name3981 (
		\u4_u2_csr0_reg[6]/P0001 ,
		\u4_u2_csr0_reg[7]/P0001 ,
		\u4_u2_dma_in_cnt_reg[4]/P0001 ,
		\u4_u2_dma_in_cnt_reg[5]/P0001 ,
		_w5731_
	);
	LUT4 #(
		.INIT('h0e0f)
	) name3982 (
		_w4491_,
		_w4496_,
		_w5730_,
		_w5731_,
		_w5732_
	);
	LUT4 #(
		.INIT('h0001)
	) name3983 (
		\u1_u3_buf0_rl_reg/P0001 ,
		\u1_u3_buf0_set_reg/P0001 ,
		\u4_u2_dma_in_cnt_reg[5]/P0001 ,
		\u4_u2_set_r_reg/P0001 ,
		_w5733_
	);
	LUT3 #(
		.INIT('h0e)
	) name3984 (
		\u4_u2_dma_in_cnt_reg[5]/P0001 ,
		\u4_u2_ep_match_r_reg/P0001 ,
		\u4_u2_r5_reg/NET0131 ,
		_w5734_
	);
	LUT2 #(
		.INIT('h4)
	) name3985 (
		_w5733_,
		_w5734_,
		_w5735_
	);
	LUT3 #(
		.INIT('ha8)
	) name3986 (
		\u4_u2_csr1_reg[0]/P0001 ,
		_w5730_,
		_w5735_,
		_w5736_
	);
	LUT3 #(
		.INIT('hb0)
	) name3987 (
		_w5728_,
		_w5732_,
		_w5736_,
		_w5737_
	);
	LUT3 #(
		.INIT('h08)
	) name3988 (
		rst_i_pad,
		\u5_state_reg[4]/P0001 ,
		\u5_state_reg[5]/NET0131 ,
		_w5738_
	);
	LUT4 #(
		.INIT('h0001)
	) name3989 (
		\u5_state_reg[0]/P0001 ,
		\u5_state_reg[1]/P0001 ,
		\u5_state_reg[2]/P0001 ,
		\u5_state_reg[3]/P0001 ,
		_w5739_
	);
	LUT2 #(
		.INIT('h8)
	) name3990 (
		_w5738_,
		_w5739_,
		_w5740_
	);
	LUT2 #(
		.INIT('h8)
	) name3991 (
		\u1_u2_rx_data_valid_r_reg/NET0131 ,
		\u1_u2_sizu_c_reg[0]/P0001 ,
		_w5741_
	);
	LUT4 #(
		.INIT('h007f)
	) name3992 (
		\u1_u2_rx_data_valid_r_reg/NET0131 ,
		\u1_u2_sizu_c_reg[0]/P0001 ,
		\u1_u2_sizu_c_reg[1]/P0001 ,
		\u1_u2_sizu_c_reg[2]/P0001 ,
		_w5742_
	);
	LUT3 #(
		.INIT('h04)
	) name3993 (
		_w4783_,
		_w4787_,
		_w5742_,
		_w5743_
	);
	LUT3 #(
		.INIT('h20)
	) name3994 (
		rst_i_pad,
		\u1_u2_rx_dma_en_r_reg/P0001 ,
		\u1_u2_sizu_c_reg[3]/P0001 ,
		_w5744_
	);
	LUT3 #(
		.INIT('h02)
	) name3995 (
		rst_i_pad,
		\u1_u2_rx_dma_en_r_reg/P0001 ,
		\u1_u2_sizu_c_reg[3]/P0001 ,
		_w5745_
	);
	LUT3 #(
		.INIT('he4)
	) name3996 (
		_w4783_,
		_w5744_,
		_w5745_,
		_w5746_
	);
	LUT2 #(
		.INIT('h8)
	) name3997 (
		\u1_u2_sizu_c_reg[3]/P0001 ,
		\u1_u2_sizu_c_reg[4]/P0001 ,
		_w5747_
	);
	LUT4 #(
		.INIT('h6c00)
	) name3998 (
		\u1_u2_sizu_c_reg[3]/P0001 ,
		\u1_u2_sizu_c_reg[4]/P0001 ,
		_w4783_,
		_w4787_,
		_w5748_
	);
	LUT3 #(
		.INIT('h15)
	) name3999 (
		\u1_u2_sizu_c_reg[5]/P0001 ,
		_w4783_,
		_w5747_,
		_w5749_
	);
	LUT3 #(
		.INIT('h70)
	) name4000 (
		_w4783_,
		_w4784_,
		_w4787_,
		_w5750_
	);
	LUT2 #(
		.INIT('h4)
	) name4001 (
		_w5749_,
		_w5750_,
		_w5751_
	);
	LUT4 #(
		.INIT('h6a00)
	) name4002 (
		\u1_u2_sizu_c_reg[6]/P0001 ,
		_w4783_,
		_w4784_,
		_w4787_,
		_w5752_
	);
	LUT4 #(
		.INIT('h8000)
	) name4003 (
		\u1_u2_sizu_c_reg[3]/P0001 ,
		\u1_u2_sizu_c_reg[4]/P0001 ,
		\u1_u2_sizu_c_reg[5]/P0001 ,
		\u1_u2_sizu_c_reg[6]/P0001 ,
		_w5753_
	);
	LUT3 #(
		.INIT('h15)
	) name4004 (
		\u1_u2_sizu_c_reg[7]/P0001 ,
		_w4783_,
		_w5753_,
		_w5754_
	);
	LUT4 #(
		.INIT('h7f00)
	) name4005 (
		_w4783_,
		_w4784_,
		_w4785_,
		_w4787_,
		_w5755_
	);
	LUT2 #(
		.INIT('h4)
	) name4006 (
		_w5754_,
		_w5755_,
		_w5756_
	);
	LUT4 #(
		.INIT('h7f00)
	) name4007 (
		_w4783_,
		_w4785_,
		_w4788_,
		_w5314_,
		_w5757_
	);
	LUT3 #(
		.INIT('h02)
	) name4008 (
		rst_i_pad,
		\u1_u2_rx_dma_en_r_reg/P0001 ,
		\u1_u2_sizu_c_reg[9]/P0001 ,
		_w5758_
	);
	LUT4 #(
		.INIT('h8000)
	) name4009 (
		_w4783_,
		_w4785_,
		_w4788_,
		_w5758_,
		_w5759_
	);
	LUT2 #(
		.INIT('he)
	) name4010 (
		_w5757_,
		_w5759_,
		_w5760_
	);
	LUT4 #(
		.INIT('h0010)
	) name4011 (
		\u0_u0_state_reg[10]/P0001 ,
		\u0_u0_state_reg[7]/NET0131 ,
		\u0_u0_state_reg[8]/NET0131 ,
		\u0_u0_state_reg[9]/P0001 ,
		_w5761_
	);
	LUT4 #(
		.INIT('h8000)
	) name4012 (
		_w4094_,
		_w4098_,
		_w4101_,
		_w5761_,
		_w5762_
	);
	LUT4 #(
		.INIT('h8000)
	) name4013 (
		_w4097_,
		_w4108_,
		_w4109_,
		_w4323_,
		_w5763_
	);
	LUT2 #(
		.INIT('h9)
	) name4014 (
		\u0_u0_state_reg[1]/P0001 ,
		\u0_u0_state_reg[2]/NET0131 ,
		_w5764_
	);
	LUT3 #(
		.INIT('ha2)
	) name4015 (
		_w5762_,
		_w5763_,
		_w5764_,
		_w5765_
	);
	LUT4 #(
		.INIT('h0020)
	) name4016 (
		\u0_u0_T1_gt_3_0_mS_reg/P0001 ,
		\u0_u0_mode_hs_reg/P0001 ,
		\u0_u0_state_reg[1]/P0001 ,
		\u0_u0_state_reg[2]/NET0131 ,
		_w5766_
	);
	LUT2 #(
		.INIT('h4)
	) name4017 (
		_w4316_,
		_w5766_,
		_w5767_
	);
	LUT4 #(
		.INIT('h2a3f)
	) name4018 (
		_w4316_,
		_w4345_,
		_w4355_,
		_w5766_,
		_w5768_
	);
	LUT2 #(
		.INIT('h2)
	) name4019 (
		_w5763_,
		_w5768_,
		_w5769_
	);
	LUT2 #(
		.INIT('h4)
	) name4020 (
		\u0_u0_idle_cnt1_clr_reg/P0001 ,
		\u0_u0_idle_long_reg/P0001 ,
		_w5770_
	);
	LUT3 #(
		.INIT('h23)
	) name4021 (
		\u0_u0_T1_gt_5_0_mS_reg/P0001 ,
		\u0_u0_idle_cnt1_reg[4]/P0001 ,
		\u0_u0_ps_cnt_clr_reg/P0001 ,
		_w5771_
	);
	LUT3 #(
		.INIT('h10)
	) name4022 (
		\u0_u0_T1_gt_5_0_mS_reg/P0001 ,
		\u0_u0_idle_cnt1_next_reg[4]/P0001 ,
		\u0_u0_ps_cnt_clr_reg/P0001 ,
		_w5772_
	);
	LUT3 #(
		.INIT('h02)
	) name4023 (
		_w5770_,
		_w5771_,
		_w5772_,
		_w5773_
	);
	LUT3 #(
		.INIT('hd0)
	) name4024 (
		_w5763_,
		_w5768_,
		_w5773_,
		_w5774_
	);
	LUT2 #(
		.INIT('h4)
	) name4025 (
		_w5765_,
		_w5774_,
		_w5775_
	);
	LUT2 #(
		.INIT('h2)
	) name4026 (
		\u4_u0_buf0_orig_reg[26]/P0001 ,
		\u4_u0_dma_in_cnt_reg[7]/P0001 ,
		_w5776_
	);
	LUT4 #(
		.INIT('hf531)
	) name4027 (
		\u4_u0_buf0_orig_reg[27]/P0001 ,
		\u4_u0_buf0_orig_reg[28]/P0001 ,
		\u4_u0_dma_in_cnt_reg[8]/P0001 ,
		\u4_u0_dma_in_cnt_reg[9]/P0001 ,
		_w5777_
	);
	LUT4 #(
		.INIT('h8caf)
	) name4028 (
		\u4_u0_buf0_orig_reg[25]/P0001 ,
		\u4_u0_buf0_orig_reg[26]/P0001 ,
		\u4_u0_dma_in_cnt_reg[6]/P0001 ,
		\u4_u0_dma_in_cnt_reg[7]/P0001 ,
		_w5778_
	);
	LUT3 #(
		.INIT('h04)
	) name4029 (
		_w5776_,
		_w5777_,
		_w5778_,
		_w5779_
	);
	LUT4 #(
		.INIT('h8caf)
	) name4030 (
		\u4_u0_buf0_orig_reg[23]/P0001 ,
		\u4_u0_buf0_orig_reg[24]/P0001 ,
		\u4_u0_dma_in_cnt_reg[4]/P0001 ,
		\u4_u0_dma_in_cnt_reg[5]/P0001 ,
		_w5780_
	);
	LUT4 #(
		.INIT('hf531)
	) name4031 (
		\u4_u0_buf0_orig_reg[22]/P0001 ,
		\u4_u0_buf0_orig_reg[23]/P0001 ,
		\u4_u0_dma_in_cnt_reg[3]/P0001 ,
		\u4_u0_dma_in_cnt_reg[4]/P0001 ,
		_w5781_
	);
	LUT2 #(
		.INIT('h2)
	) name4032 (
		_w5780_,
		_w5781_,
		_w5782_
	);
	LUT4 #(
		.INIT('h08cc)
	) name4033 (
		\u4_u0_buf0_orig_reg[19]/P0001 ,
		\u4_u0_buf0_orig_reg[20]/P0001 ,
		\u4_u0_dma_in_cnt_reg[0]/P0001 ,
		\u4_u0_dma_in_cnt_reg[1]/P0001 ,
		_w5783_
	);
	LUT2 #(
		.INIT('h2)
	) name4034 (
		\u4_u0_buf0_orig_reg[21]/P0001 ,
		\u4_u0_dma_in_cnt_reg[2]/P0001 ,
		_w5784_
	);
	LUT3 #(
		.INIT('h02)
	) name4035 (
		\u4_u0_buf0_orig_reg[19]/P0001 ,
		\u4_u0_dma_in_cnt_reg[0]/P0001 ,
		\u4_u0_dma_in_cnt_reg[1]/P0001 ,
		_w5785_
	);
	LUT3 #(
		.INIT('h01)
	) name4036 (
		_w5783_,
		_w5784_,
		_w5785_,
		_w5786_
	);
	LUT4 #(
		.INIT('h8caf)
	) name4037 (
		\u4_u0_buf0_orig_reg[21]/P0001 ,
		\u4_u0_buf0_orig_reg[22]/P0001 ,
		\u4_u0_dma_in_cnt_reg[2]/P0001 ,
		\u4_u0_dma_in_cnt_reg[3]/P0001 ,
		_w5787_
	);
	LUT2 #(
		.INIT('h8)
	) name4038 (
		_w5780_,
		_w5787_,
		_w5788_
	);
	LUT4 #(
		.INIT('hf531)
	) name4039 (
		\u4_u0_buf0_orig_reg[24]/P0001 ,
		\u4_u0_buf0_orig_reg[25]/P0001 ,
		\u4_u0_dma_in_cnt_reg[5]/P0001 ,
		\u4_u0_dma_in_cnt_reg[6]/P0001 ,
		_w5789_
	);
	LUT3 #(
		.INIT('h40)
	) name4040 (
		_w5776_,
		_w5777_,
		_w5789_,
		_w5790_
	);
	LUT4 #(
		.INIT('h4500)
	) name4041 (
		_w5782_,
		_w5786_,
		_w5788_,
		_w5790_,
		_w5791_
	);
	LUT2 #(
		.INIT('h2)
	) name4042 (
		\u4_u0_csr1_reg[11]/P0001 ,
		\u4_u0_csr1_reg[12]/P0001 ,
		_w5792_
	);
	LUT3 #(
		.INIT('h8c)
	) name4043 (
		\u4_u0_buf0_orig_reg[30]/NET0131 ,
		\u4_u0_csr1_reg[0]/P0001 ,
		\u4_u0_dma_in_cnt_reg[11]/P0001 ,
		_w5793_
	);
	LUT4 #(
		.INIT('h5010)
	) name4044 (
		\u4_u0_buf0_orig_reg[27]/P0001 ,
		\u4_u0_buf0_orig_reg[28]/P0001 ,
		\u4_u0_dma_in_cnt_reg[8]/P0001 ,
		\u4_u0_dma_in_cnt_reg[9]/P0001 ,
		_w5794_
	);
	LUT4 #(
		.INIT('h8acf)
	) name4045 (
		\u4_u0_buf0_orig_reg[28]/P0001 ,
		\u4_u0_buf0_orig_reg[29]/NET0131 ,
		\u4_u0_dma_in_cnt_reg[10]/P0001 ,
		\u4_u0_dma_in_cnt_reg[9]/P0001 ,
		_w5795_
	);
	LUT4 #(
		.INIT('h0800)
	) name4046 (
		_w5792_,
		_w5793_,
		_w5794_,
		_w5795_,
		_w5796_
	);
	LUT4 #(
		.INIT('hf531)
	) name4047 (
		\u4_u0_buf0_orig_reg[29]/NET0131 ,
		\u4_u0_buf0_orig_reg[30]/NET0131 ,
		\u4_u0_dma_in_cnt_reg[10]/P0001 ,
		\u4_u0_dma_in_cnt_reg[11]/P0001 ,
		_w5797_
	);
	LUT3 #(
		.INIT('h08)
	) name4048 (
		_w5792_,
		_w5793_,
		_w5797_,
		_w5798_
	);
	LUT2 #(
		.INIT('h1)
	) name4049 (
		\u4_u0_dma_out_cnt_reg[10]/P0001 ,
		\u4_u0_dma_out_cnt_reg[11]/P0001 ,
		_w5799_
	);
	LUT4 #(
		.INIT('h0001)
	) name4050 (
		\u4_u0_dma_out_cnt_reg[2]/P0001 ,
		\u4_u0_dma_out_cnt_reg[3]/P0001 ,
		\u4_u0_dma_out_cnt_reg[4]/P0001 ,
		\u4_u0_dma_out_cnt_reg[5]/P0001 ,
		_w5800_
	);
	LUT4 #(
		.INIT('h8000)
	) name4051 (
		_w4682_,
		_w4984_,
		_w5799_,
		_w5800_,
		_w5801_
	);
	LUT3 #(
		.INIT('h20)
	) name4052 (
		\u4_u0_csr1_reg[0]/P0001 ,
		\u4_u0_csr1_reg[11]/P0001 ,
		\u4_u0_csr1_reg[12]/P0001 ,
		_w5802_
	);
	LUT3 #(
		.INIT('h45)
	) name4053 (
		_w5798_,
		_w5801_,
		_w5802_,
		_w5803_
	);
	LUT4 #(
		.INIT('hef00)
	) name4054 (
		_w5779_,
		_w5791_,
		_w5796_,
		_w5803_,
		_w5804_
	);
	LUT3 #(
		.INIT('h01)
	) name4055 (
		\u4_u0_r2_reg/P0001 ,
		\u4_u0_r4_reg/P0001 ,
		\u4_u0_r5_reg/NET0131 ,
		_w5805_
	);
	LUT2 #(
		.INIT('h4)
	) name4056 (
		_w5804_,
		_w5805_,
		_w5806_
	);
	LUT4 #(
		.INIT('hf531)
	) name4057 (
		\u4_u1_buf0_orig_reg[26]/P0001 ,
		\u4_u1_buf0_orig_reg[27]/P0001 ,
		\u4_u1_dma_in_cnt_reg[7]/P0001 ,
		\u4_u1_dma_in_cnt_reg[8]/P0001 ,
		_w5807_
	);
	LUT4 #(
		.INIT('h8caf)
	) name4058 (
		\u4_u1_buf0_orig_reg[25]/P0001 ,
		\u4_u1_buf0_orig_reg[26]/P0001 ,
		\u4_u1_dma_in_cnt_reg[6]/P0001 ,
		\u4_u1_dma_in_cnt_reg[7]/P0001 ,
		_w5808_
	);
	LUT2 #(
		.INIT('h2)
	) name4059 (
		_w5807_,
		_w5808_,
		_w5809_
	);
	LUT4 #(
		.INIT('h8caf)
	) name4060 (
		\u4_u1_buf0_orig_reg[23]/P0001 ,
		\u4_u1_buf0_orig_reg[24]/P0001 ,
		\u4_u1_dma_in_cnt_reg[4]/P0001 ,
		\u4_u1_dma_in_cnt_reg[5]/P0001 ,
		_w5810_
	);
	LUT4 #(
		.INIT('hf531)
	) name4061 (
		\u4_u1_buf0_orig_reg[22]/P0001 ,
		\u4_u1_buf0_orig_reg[23]/P0001 ,
		\u4_u1_dma_in_cnt_reg[3]/P0001 ,
		\u4_u1_dma_in_cnt_reg[4]/P0001 ,
		_w5811_
	);
	LUT2 #(
		.INIT('h2)
	) name4062 (
		_w5810_,
		_w5811_,
		_w5812_
	);
	LUT4 #(
		.INIT('h080a)
	) name4063 (
		\u4_u1_buf0_orig_reg[19]/P0001 ,
		\u4_u1_buf0_orig_reg[20]/P0001 ,
		\u4_u1_dma_in_cnt_reg[0]/P0001 ,
		\u4_u1_dma_in_cnt_reg[1]/P0001 ,
		_w5813_
	);
	LUT4 #(
		.INIT('hf531)
	) name4064 (
		\u4_u1_buf0_orig_reg[20]/P0001 ,
		\u4_u1_buf0_orig_reg[21]/P0001 ,
		\u4_u1_dma_in_cnt_reg[1]/P0001 ,
		\u4_u1_dma_in_cnt_reg[2]/P0001 ,
		_w5814_
	);
	LUT4 #(
		.INIT('h8caf)
	) name4065 (
		\u4_u1_buf0_orig_reg[21]/P0001 ,
		\u4_u1_buf0_orig_reg[22]/P0001 ,
		\u4_u1_dma_in_cnt_reg[2]/P0001 ,
		\u4_u1_dma_in_cnt_reg[3]/P0001 ,
		_w5815_
	);
	LUT4 #(
		.INIT('h8a00)
	) name4066 (
		_w5810_,
		_w5813_,
		_w5814_,
		_w5815_,
		_w5816_
	);
	LUT4 #(
		.INIT('hf531)
	) name4067 (
		\u4_u1_buf0_orig_reg[24]/P0001 ,
		\u4_u1_buf0_orig_reg[25]/P0001 ,
		\u4_u1_dma_in_cnt_reg[5]/P0001 ,
		\u4_u1_dma_in_cnt_reg[6]/P0001 ,
		_w5817_
	);
	LUT2 #(
		.INIT('h8)
	) name4068 (
		_w5807_,
		_w5817_,
		_w5818_
	);
	LUT4 #(
		.INIT('h5455)
	) name4069 (
		_w5809_,
		_w5812_,
		_w5816_,
		_w5818_,
		_w5819_
	);
	LUT2 #(
		.INIT('h4)
	) name4070 (
		\u4_u1_buf0_orig_reg[30]/NET0131 ,
		\u4_u1_dma_in_cnt_reg[11]/P0001 ,
		_w5820_
	);
	LUT2 #(
		.INIT('h2)
	) name4071 (
		\u4_u1_csr1_reg[11]/P0001 ,
		\u4_u1_csr1_reg[12]/P0001 ,
		_w5821_
	);
	LUT3 #(
		.INIT('h08)
	) name4072 (
		\u4_u1_csr1_reg[0]/P0001 ,
		\u4_u1_csr1_reg[11]/P0001 ,
		\u4_u1_csr1_reg[12]/P0001 ,
		_w5822_
	);
	LUT4 #(
		.INIT('h5010)
	) name4073 (
		\u4_u1_buf0_orig_reg[29]/NET0131 ,
		\u4_u1_buf0_orig_reg[30]/NET0131 ,
		\u4_u1_dma_in_cnt_reg[10]/P0001 ,
		\u4_u1_dma_in_cnt_reg[11]/P0001 ,
		_w5823_
	);
	LUT4 #(
		.INIT('h8caf)
	) name4074 (
		\u4_u1_buf0_orig_reg[27]/P0001 ,
		\u4_u1_buf0_orig_reg[28]/P0001 ,
		\u4_u1_dma_in_cnt_reg[8]/P0001 ,
		\u4_u1_dma_in_cnt_reg[9]/P0001 ,
		_w5824_
	);
	LUT4 #(
		.INIT('h0400)
	) name4075 (
		_w5820_,
		_w5822_,
		_w5823_,
		_w5824_,
		_w5825_
	);
	LUT2 #(
		.INIT('h2)
	) name4076 (
		\u4_u1_buf0_orig_reg[28]/P0001 ,
		\u4_u1_dma_in_cnt_reg[9]/P0001 ,
		_w5826_
	);
	LUT4 #(
		.INIT('hf531)
	) name4077 (
		\u4_u1_buf0_orig_reg[29]/NET0131 ,
		\u4_u1_buf0_orig_reg[30]/NET0131 ,
		\u4_u1_dma_in_cnt_reg[10]/P0001 ,
		\u4_u1_dma_in_cnt_reg[11]/P0001 ,
		_w5827_
	);
	LUT4 #(
		.INIT('h4044)
	) name4078 (
		_w5820_,
		_w5822_,
		_w5826_,
		_w5827_,
		_w5828_
	);
	LUT2 #(
		.INIT('h1)
	) name4079 (
		\u4_u1_dma_out_cnt_reg[10]/P0001 ,
		\u4_u1_dma_out_cnt_reg[11]/P0001 ,
		_w5829_
	);
	LUT4 #(
		.INIT('h0001)
	) name4080 (
		\u4_u1_dma_out_cnt_reg[2]/P0001 ,
		\u4_u1_dma_out_cnt_reg[3]/P0001 ,
		\u4_u1_dma_out_cnt_reg[4]/P0001 ,
		\u4_u1_dma_out_cnt_reg[5]/P0001 ,
		_w5830_
	);
	LUT4 #(
		.INIT('h8000)
	) name4081 (
		_w4712_,
		_w5018_,
		_w5829_,
		_w5830_,
		_w5831_
	);
	LUT3 #(
		.INIT('h20)
	) name4082 (
		\u4_u1_csr1_reg[0]/P0001 ,
		\u4_u1_csr1_reg[11]/P0001 ,
		\u4_u1_csr1_reg[12]/P0001 ,
		_w5832_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name4083 (
		_w5823_,
		_w5828_,
		_w5831_,
		_w5832_,
		_w5833_
	);
	LUT3 #(
		.INIT('h01)
	) name4084 (
		\u4_u1_r2_reg/P0001 ,
		\u4_u1_r4_reg/P0001 ,
		\u4_u1_r5_reg/NET0131 ,
		_w5834_
	);
	LUT4 #(
		.INIT('h8f00)
	) name4085 (
		_w5819_,
		_w5825_,
		_w5833_,
		_w5834_,
		_w5835_
	);
	LUT2 #(
		.INIT('h8)
	) name4086 (
		_w3740_,
		_w4856_,
		_w5836_
	);
	LUT4 #(
		.INIT('h0208)
	) name4087 (
		rst_i_pad,
		\u1_u2_rx_data_valid_r_reg/NET0131 ,
		\u1_u2_rx_dma_en_r_reg/P0001 ,
		\u1_u2_sizu_c_reg[0]/P0001 ,
		_w5837_
	);
	LUT3 #(
		.INIT('h48)
	) name4088 (
		\u1_u2_sizu_c_reg[1]/P0001 ,
		_w4787_,
		_w5741_,
		_w5838_
	);
	LUT2 #(
		.INIT('h8)
	) name4089 (
		_w2240_,
		_w2241_,
		_w5839_
	);
	LUT2 #(
		.INIT('h1)
	) name4090 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w5840_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name4091 (
		\u4_u0_buf1_reg[0]/P0001 ,
		\u4_u0_csr0_reg[0]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w5841_
	);
	LUT4 #(
		.INIT('hf53f)
	) name4092 (
		\u4_u0_buf0_reg[0]/P0001 ,
		\u4_u0_int_stat_reg[0]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w5842_
	);
	LUT4 #(
		.INIT('h0888)
	) name4093 (
		_w2240_,
		_w2241_,
		_w5841_,
		_w5842_,
		_w5843_
	);
	LUT2 #(
		.INIT('h8)
	) name4094 (
		_w2228_,
		_w2240_,
		_w5844_
	);
	LUT4 #(
		.INIT('hf5f3)
	) name4095 (
		\u4_u2_buf0_reg[0]/P0001 ,
		\u4_u2_csr0_reg[0]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w5845_
	);
	LUT4 #(
		.INIT('h5f3f)
	) name4096 (
		\u4_u2_buf1_reg[0]/P0001 ,
		\u4_u2_int_stat_reg[0]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w5846_
	);
	LUT4 #(
		.INIT('h0888)
	) name4097 (
		_w2228_,
		_w2240_,
		_w5845_,
		_w5846_,
		_w5847_
	);
	LUT2 #(
		.INIT('h8)
	) name4098 (
		_w2227_,
		_w2228_,
		_w5848_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name4099 (
		\u4_u3_buf1_reg[0]/P0001 ,
		\u4_u3_csr0_reg[0]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w5849_
	);
	LUT4 #(
		.INIT('hf53f)
	) name4100 (
		\u4_u3_buf0_reg[0]/P0001 ,
		\u4_u3_int_stat_reg[0]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w5850_
	);
	LUT4 #(
		.INIT('h0888)
	) name4101 (
		_w2227_,
		_w2228_,
		_w5849_,
		_w5850_,
		_w5851_
	);
	LUT3 #(
		.INIT('h01)
	) name4102 (
		_w5843_,
		_w5847_,
		_w5851_,
		_w5852_
	);
	LUT4 #(
		.INIT('h0008)
	) name4103 (
		\u4_funct_adr_reg[0]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w5853_
	);
	LUT4 #(
		.INIT('h0002)
	) name4104 (
		\u0_u0_usb_suspend_reg/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w5854_
	);
	LUT4 #(
		.INIT('h0080)
	) name4105 (
		\u4_int_srca_reg[0]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w5855_
	);
	LUT3 #(
		.INIT('h01)
	) name4106 (
		_w5853_,
		_w5854_,
		_w5855_,
		_w5856_
	);
	LUT4 #(
		.INIT('h0020)
	) name4107 (
		\u4_inta_msk_reg[0]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w5857_
	);
	LUT4 #(
		.INIT('h0200)
	) name4108 (
		\u1_sof_time_reg[0]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w5858_
	);
	LUT4 #(
		.INIT('h0800)
	) name4109 (
		\u4_utmi_vend_stat_r_reg[0]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w5859_
	);
	LUT3 #(
		.INIT('h01)
	) name4110 (
		_w5857_,
		_w5858_,
		_w5859_,
		_w5860_
	);
	LUT4 #(
		.INIT('h0001)
	) name4111 (
		\wb_addr_i[5]_pad ,
		\wb_addr_i[6]_pad ,
		\wb_addr_i[7]_pad ,
		\wb_addr_i[8]_pad ,
		_w5861_
	);
	LUT2 #(
		.INIT('h8)
	) name4112 (
		_w2227_,
		_w2241_,
		_w5862_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name4113 (
		\u4_u1_buf1_reg[0]/P0001 ,
		\u4_u1_csr0_reg[0]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w5863_
	);
	LUT4 #(
		.INIT('hf53f)
	) name4114 (
		\u4_u1_buf0_reg[0]/P0001 ,
		\u4_u1_int_stat_reg[0]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w5864_
	);
	LUT4 #(
		.INIT('h0888)
	) name4115 (
		_w2227_,
		_w2241_,
		_w5863_,
		_w5864_,
		_w5865_
	);
	LUT4 #(
		.INIT('h008f)
	) name4116 (
		_w5856_,
		_w5860_,
		_w5861_,
		_w5865_,
		_w5866_
	);
	LUT2 #(
		.INIT('h7)
	) name4117 (
		_w5852_,
		_w5866_,
		_w5867_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name4118 (
		\u4_u0_buf1_reg[1]/P0001 ,
		\u4_u0_csr0_reg[1]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w5868_
	);
	LUT4 #(
		.INIT('hf53f)
	) name4119 (
		\u4_u0_buf0_reg[1]/P0001 ,
		\u4_u0_int_stat_reg[1]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w5869_
	);
	LUT4 #(
		.INIT('h0888)
	) name4120 (
		_w2240_,
		_w2241_,
		_w5868_,
		_w5869_,
		_w5870_
	);
	LUT4 #(
		.INIT('hf5f3)
	) name4121 (
		\u4_u3_buf0_reg[1]/P0001 ,
		\u4_u3_csr0_reg[1]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w5871_
	);
	LUT4 #(
		.INIT('h5f3f)
	) name4122 (
		\u4_u3_buf1_reg[1]/P0001 ,
		\u4_u3_int_stat_reg[1]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w5872_
	);
	LUT4 #(
		.INIT('h0888)
	) name4123 (
		_w2227_,
		_w2228_,
		_w5871_,
		_w5872_,
		_w5873_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name4124 (
		\u4_u2_buf1_reg[1]/P0001 ,
		\u4_u2_csr0_reg[1]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w5874_
	);
	LUT4 #(
		.INIT('hf53f)
	) name4125 (
		\u4_u2_buf0_reg[1]/P0001 ,
		\u4_u2_int_stat_reg[1]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w5875_
	);
	LUT4 #(
		.INIT('h0888)
	) name4126 (
		_w2228_,
		_w2240_,
		_w5874_,
		_w5875_,
		_w5876_
	);
	LUT3 #(
		.INIT('h01)
	) name4127 (
		_w5870_,
		_w5873_,
		_w5876_,
		_w5877_
	);
	LUT4 #(
		.INIT('h0008)
	) name4128 (
		\u4_funct_adr_reg[1]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w5878_
	);
	LUT4 #(
		.INIT('h0002)
	) name4129 (
		\u0_u0_mode_hs_reg/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w5879_
	);
	LUT4 #(
		.INIT('h0080)
	) name4130 (
		\u4_int_srca_reg[1]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w5880_
	);
	LUT3 #(
		.INIT('h01)
	) name4131 (
		_w5878_,
		_w5879_,
		_w5880_,
		_w5881_
	);
	LUT4 #(
		.INIT('h0020)
	) name4132 (
		\u4_inta_msk_reg[1]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w5882_
	);
	LUT4 #(
		.INIT('h0200)
	) name4133 (
		\u1_sof_time_reg[1]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w5883_
	);
	LUT4 #(
		.INIT('h0800)
	) name4134 (
		\u4_utmi_vend_stat_r_reg[1]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w5884_
	);
	LUT3 #(
		.INIT('h01)
	) name4135 (
		_w5882_,
		_w5883_,
		_w5884_,
		_w5885_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name4136 (
		\u4_u1_buf1_reg[1]/P0001 ,
		\u4_u1_csr0_reg[1]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w5886_
	);
	LUT4 #(
		.INIT('hf53f)
	) name4137 (
		\u4_u1_buf0_reg[1]/P0001 ,
		\u4_u1_int_stat_reg[1]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w5887_
	);
	LUT4 #(
		.INIT('h0888)
	) name4138 (
		_w2227_,
		_w2241_,
		_w5886_,
		_w5887_,
		_w5888_
	);
	LUT4 #(
		.INIT('h00d5)
	) name4139 (
		_w5861_,
		_w5881_,
		_w5885_,
		_w5888_,
		_w5889_
	);
	LUT2 #(
		.INIT('h7)
	) name4140 (
		_w5877_,
		_w5889_,
		_w5890_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name4141 (
		\u4_u0_buf1_reg[2]/P0001 ,
		\u4_u0_csr0_reg[2]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w5891_
	);
	LUT4 #(
		.INIT('hf53f)
	) name4142 (
		\u4_u0_buf0_reg[2]/P0001 ,
		\u4_u0_int_stat_reg[2]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w5892_
	);
	LUT4 #(
		.INIT('h0888)
	) name4143 (
		_w2240_,
		_w2241_,
		_w5891_,
		_w5892_,
		_w5893_
	);
	LUT4 #(
		.INIT('hf5f3)
	) name4144 (
		\u4_u3_buf0_reg[2]/P0001 ,
		\u4_u3_csr0_reg[2]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w5894_
	);
	LUT4 #(
		.INIT('h5f3f)
	) name4145 (
		\u4_u3_buf1_reg[2]/P0001 ,
		\u4_u3_int_stat_reg[2]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w5895_
	);
	LUT4 #(
		.INIT('h0888)
	) name4146 (
		_w2227_,
		_w2228_,
		_w5894_,
		_w5895_,
		_w5896_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name4147 (
		\u4_u2_buf1_reg[2]/P0001 ,
		\u4_u2_csr0_reg[2]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w5897_
	);
	LUT4 #(
		.INIT('hf53f)
	) name4148 (
		\u4_u2_buf0_reg[2]/P0001 ,
		\u4_u2_int_stat_reg[2]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w5898_
	);
	LUT4 #(
		.INIT('h0888)
	) name4149 (
		_w2228_,
		_w2240_,
		_w5897_,
		_w5898_,
		_w5899_
	);
	LUT3 #(
		.INIT('h01)
	) name4150 (
		_w5893_,
		_w5896_,
		_w5899_,
		_w5900_
	);
	LUT4 #(
		.INIT('h0008)
	) name4151 (
		\u4_funct_adr_reg[2]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w5901_
	);
	LUT4 #(
		.INIT('h0002)
	) name4152 (
		\u0_u0_usb_attached_reg/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w5902_
	);
	LUT4 #(
		.INIT('h0080)
	) name4153 (
		\u4_int_srca_reg[2]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w5903_
	);
	LUT3 #(
		.INIT('h01)
	) name4154 (
		_w5901_,
		_w5902_,
		_w5903_,
		_w5904_
	);
	LUT4 #(
		.INIT('h0020)
	) name4155 (
		\u4_inta_msk_reg[2]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w5905_
	);
	LUT4 #(
		.INIT('h0200)
	) name4156 (
		\u1_sof_time_reg[2]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w5906_
	);
	LUT4 #(
		.INIT('h0800)
	) name4157 (
		\u4_utmi_vend_stat_r_reg[2]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w5907_
	);
	LUT3 #(
		.INIT('h01)
	) name4158 (
		_w5905_,
		_w5906_,
		_w5907_,
		_w5908_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name4159 (
		\u4_u1_buf1_reg[2]/P0001 ,
		\u4_u1_csr0_reg[2]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w5909_
	);
	LUT4 #(
		.INIT('hf53f)
	) name4160 (
		\u4_u1_buf0_reg[2]/P0001 ,
		\u4_u1_int_stat_reg[2]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w5910_
	);
	LUT4 #(
		.INIT('h0888)
	) name4161 (
		_w2227_,
		_w2241_,
		_w5909_,
		_w5910_,
		_w5911_
	);
	LUT4 #(
		.INIT('h00d5)
	) name4162 (
		_w5861_,
		_w5904_,
		_w5908_,
		_w5911_,
		_w5912_
	);
	LUT2 #(
		.INIT('h7)
	) name4163 (
		_w5900_,
		_w5912_,
		_w5913_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name4164 (
		\u4_u0_buf1_reg[3]/P0001 ,
		\u4_u0_csr0_reg[3]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w5914_
	);
	LUT4 #(
		.INIT('hf53f)
	) name4165 (
		\u4_u0_buf0_reg[3]/P0001 ,
		\u4_u0_int_stat_reg[3]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w5915_
	);
	LUT4 #(
		.INIT('h0888)
	) name4166 (
		_w2240_,
		_w2241_,
		_w5914_,
		_w5915_,
		_w5916_
	);
	LUT4 #(
		.INIT('hf5f3)
	) name4167 (
		\u4_u3_buf0_reg[3]/P0001 ,
		\u4_u3_csr0_reg[3]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w5917_
	);
	LUT4 #(
		.INIT('h5f3f)
	) name4168 (
		\u4_u3_buf1_reg[3]/P0001 ,
		\u4_u3_int_stat_reg[3]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w5918_
	);
	LUT4 #(
		.INIT('h0888)
	) name4169 (
		_w2227_,
		_w2228_,
		_w5917_,
		_w5918_,
		_w5919_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name4170 (
		\u4_u2_buf1_reg[3]/P0001 ,
		\u4_u2_csr0_reg[3]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w5920_
	);
	LUT4 #(
		.INIT('hf53f)
	) name4171 (
		\u4_u2_buf0_reg[3]/P0001 ,
		\u4_u2_int_stat_reg[3]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w5921_
	);
	LUT4 #(
		.INIT('h0888)
	) name4172 (
		_w2228_,
		_w2240_,
		_w5920_,
		_w5921_,
		_w5922_
	);
	LUT3 #(
		.INIT('h01)
	) name4173 (
		_w5916_,
		_w5919_,
		_w5922_,
		_w5923_
	);
	LUT4 #(
		.INIT('h0008)
	) name4174 (
		\u4_funct_adr_reg[3]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w5924_
	);
	LUT4 #(
		.INIT('h0200)
	) name4175 (
		\u1_sof_time_reg[3]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w5925_
	);
	LUT4 #(
		.INIT('h0080)
	) name4176 (
		\u4_int_srca_reg[3]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w5926_
	);
	LUT3 #(
		.INIT('h01)
	) name4177 (
		_w5924_,
		_w5925_,
		_w5926_,
		_w5927_
	);
	LUT4 #(
		.INIT('h0020)
	) name4178 (
		\u4_inta_msk_reg[3]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w5928_
	);
	LUT4 #(
		.INIT('h0002)
	) name4179 (
		\LineState_r_reg[0]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w5929_
	);
	LUT4 #(
		.INIT('h0800)
	) name4180 (
		\u4_utmi_vend_stat_r_reg[3]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w5930_
	);
	LUT3 #(
		.INIT('h01)
	) name4181 (
		_w5928_,
		_w5929_,
		_w5930_,
		_w5931_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name4182 (
		\u4_u1_buf1_reg[3]/P0001 ,
		\u4_u1_csr0_reg[3]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w5932_
	);
	LUT4 #(
		.INIT('hf53f)
	) name4183 (
		\u4_u1_buf0_reg[3]/P0001 ,
		\u4_u1_int_stat_reg[3]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w5933_
	);
	LUT4 #(
		.INIT('h0888)
	) name4184 (
		_w2227_,
		_w2241_,
		_w5932_,
		_w5933_,
		_w5934_
	);
	LUT4 #(
		.INIT('h00d5)
	) name4185 (
		_w5861_,
		_w5927_,
		_w5931_,
		_w5934_,
		_w5935_
	);
	LUT2 #(
		.INIT('h7)
	) name4186 (
		_w5923_,
		_w5935_,
		_w5936_
	);
	LUT3 #(
		.INIT('h82)
	) name4187 (
		\u1_u0_pid_reg[0]/NET0131 ,
		\u1_u0_pid_reg[2]/NET0131 ,
		\u1_u3_this_dpid_reg[1]/P0001 ,
		_w5937_
	);
	LUT3 #(
		.INIT('h82)
	) name4188 (
		\u1_u0_pid_reg[1]/NET0131 ,
		\u1_u0_pid_reg[3]/NET0131 ,
		\u1_u3_this_dpid_reg[0]/P0001 ,
		_w5938_
	);
	LUT2 #(
		.INIT('h7)
	) name4189 (
		_w5937_,
		_w5938_,
		_w5939_
	);
	LUT3 #(
		.INIT('hac)
	) name4190 (
		\u1_u2_sizu_c_reg[1]/P0001 ,
		\u1_u3_new_size_reg[1]/P0001 ,
		\u1_u3_out_to_small_r_reg/P0001 ,
		_w5940_
	);
	LUT3 #(
		.INIT('h59)
	) name4191 (
		\u1_u3_adr_reg[2]/P0001 ,
		_w2795_,
		_w2797_,
		_w5941_
	);
	LUT4 #(
		.INIT('h4db2)
	) name4192 (
		\u1_u3_adr_reg[1]/P0001 ,
		_w2785_,
		_w4071_,
		_w5941_,
		_w5942_
	);
	LUT3 #(
		.INIT('h59)
	) name4193 (
		\u1_u3_adr_reg[3]/P0001 ,
		_w2810_,
		_w2812_,
		_w5943_
	);
	LUT3 #(
		.INIT('he1)
	) name4194 (
		_w4073_,
		_w4075_,
		_w5943_,
		_w5944_
	);
	LUT2 #(
		.INIT('h4)
	) name4195 (
		\u4_u3_buf0_orig_reg[28]/P0001 ,
		\u4_u3_dma_out_cnt_reg[9]/P0001 ,
		_w5945_
	);
	LUT2 #(
		.INIT('h4)
	) name4196 (
		\u4_u3_buf0_orig_reg[27]/P0001 ,
		\u4_u3_dma_out_cnt_reg[8]/P0001 ,
		_w5946_
	);
	LUT2 #(
		.INIT('h2)
	) name4197 (
		\u4_u3_buf0_orig_reg[26]/P0001 ,
		\u4_u3_dma_out_cnt_reg[7]/P0001 ,
		_w5947_
	);
	LUT4 #(
		.INIT('h08ce)
	) name4198 (
		\u4_u3_buf0_orig_reg[26]/P0001 ,
		\u4_u3_buf0_orig_reg[27]/P0001 ,
		\u4_u3_dma_out_cnt_reg[7]/P0001 ,
		\u4_u3_dma_out_cnt_reg[8]/P0001 ,
		_w5948_
	);
	LUT2 #(
		.INIT('h2)
	) name4199 (
		\u4_u3_buf0_orig_reg[25]/P0001 ,
		\u4_u3_dma_out_cnt_reg[6]/P0001 ,
		_w5949_
	);
	LUT4 #(
		.INIT('h5010)
	) name4200 (
		\u4_u3_buf0_orig_reg[24]/P0001 ,
		\u4_u3_buf0_orig_reg[25]/P0001 ,
		\u4_u3_dma_out_cnt_reg[5]/P0001 ,
		\u4_u3_dma_out_cnt_reg[6]/P0001 ,
		_w5950_
	);
	LUT4 #(
		.INIT('h8caf)
	) name4201 (
		\u4_u3_buf0_orig_reg[22]/P0001 ,
		\u4_u3_buf0_orig_reg[23]/P0001 ,
		\u4_u3_dma_out_cnt_reg[3]/P0001 ,
		\u4_u3_dma_out_cnt_reg[4]/P0001 ,
		_w5951_
	);
	LUT4 #(
		.INIT('h080a)
	) name4202 (
		\u4_u3_buf0_orig_reg[22]/P0001 ,
		\u4_u3_buf0_orig_reg[23]/P0001 ,
		\u4_u3_dma_out_cnt_reg[3]/P0001 ,
		\u4_u3_dma_out_cnt_reg[4]/P0001 ,
		_w5952_
	);
	LUT4 #(
		.INIT('h8caf)
	) name4203 (
		\u4_u3_buf0_orig_reg[19]/P0001 ,
		\u4_u3_buf0_orig_reg[20]/P0001 ,
		\u4_u3_dma_in_cnt_reg[0]/P0001 ,
		\u4_u3_dma_out_cnt_reg[1]/P0001 ,
		_w5953_
	);
	LUT4 #(
		.INIT('hf531)
	) name4204 (
		\u4_u3_buf0_orig_reg[20]/P0001 ,
		\u4_u3_buf0_orig_reg[21]/P0001 ,
		\u4_u3_dma_out_cnt_reg[1]/P0001 ,
		\u4_u3_dma_out_cnt_reg[2]/P0001 ,
		_w5954_
	);
	LUT2 #(
		.INIT('h4)
	) name4205 (
		\u4_u3_buf0_orig_reg[21]/P0001 ,
		\u4_u3_dma_out_cnt_reg[2]/P0001 ,
		_w5955_
	);
	LUT4 #(
		.INIT('h008a)
	) name4206 (
		_w5951_,
		_w5953_,
		_w5954_,
		_w5955_,
		_w5956_
	);
	LUT2 #(
		.INIT('h2)
	) name4207 (
		\u4_u3_buf0_orig_reg[23]/P0001 ,
		\u4_u3_dma_out_cnt_reg[4]/P0001 ,
		_w5957_
	);
	LUT4 #(
		.INIT('hf531)
	) name4208 (
		\u4_u3_buf0_orig_reg[23]/P0001 ,
		\u4_u3_buf0_orig_reg[24]/P0001 ,
		\u4_u3_dma_out_cnt_reg[4]/P0001 ,
		\u4_u3_dma_out_cnt_reg[5]/P0001 ,
		_w5958_
	);
	LUT2 #(
		.INIT('h4)
	) name4209 (
		_w5949_,
		_w5958_,
		_w5959_
	);
	LUT4 #(
		.INIT('h5455)
	) name4210 (
		_w5950_,
		_w5952_,
		_w5956_,
		_w5959_,
		_w5960_
	);
	LUT4 #(
		.INIT('h8caf)
	) name4211 (
		\u4_u3_buf0_orig_reg[25]/P0001 ,
		\u4_u3_buf0_orig_reg[26]/P0001 ,
		\u4_u3_dma_out_cnt_reg[6]/P0001 ,
		\u4_u3_dma_out_cnt_reg[7]/P0001 ,
		_w5961_
	);
	LUT2 #(
		.INIT('h4)
	) name4212 (
		_w5946_,
		_w5961_,
		_w5962_
	);
	LUT4 #(
		.INIT('h5444)
	) name4213 (
		_w5945_,
		_w5948_,
		_w5960_,
		_w5962_,
		_w5963_
	);
	LUT2 #(
		.INIT('h2)
	) name4214 (
		\u4_u3_buf0_orig_reg[29]/NET0131 ,
		\u4_u3_dma_out_cnt_reg[10]/P0001 ,
		_w5964_
	);
	LUT2 #(
		.INIT('h9)
	) name4215 (
		\u4_u3_buf0_orig_reg[29]/NET0131 ,
		\u4_u3_dma_out_cnt_reg[10]/P0001 ,
		_w5965_
	);
	LUT2 #(
		.INIT('h2)
	) name4216 (
		\u4_u3_buf0_orig_reg[28]/P0001 ,
		\u4_u3_dma_out_cnt_reg[9]/P0001 ,
		_w5966_
	);
	LUT4 #(
		.INIT('h283c)
	) name4217 (
		\u4_u3_buf0_orig_reg[28]/P0001 ,
		\u4_u3_buf0_orig_reg[29]/NET0131 ,
		\u4_u3_dma_out_cnt_reg[10]/P0001 ,
		\u4_u3_dma_out_cnt_reg[9]/P0001 ,
		_w5967_
	);
	LUT4 #(
		.INIT('hea00)
	) name4218 (
		_w5948_,
		_w5960_,
		_w5962_,
		_w5967_,
		_w5968_
	);
	LUT4 #(
		.INIT('hff34)
	) name4219 (
		_w5963_,
		_w5965_,
		_w5966_,
		_w5968_,
		_w5969_
	);
	LUT2 #(
		.INIT('h4)
	) name4220 (
		\u4_u0_buf0_orig_reg[28]/P0001 ,
		\u4_u0_dma_out_cnt_reg[9]/P0001 ,
		_w5970_
	);
	LUT2 #(
		.INIT('h4)
	) name4221 (
		\u4_u0_buf0_orig_reg[27]/P0001 ,
		\u4_u0_dma_out_cnt_reg[8]/P0001 ,
		_w5971_
	);
	LUT2 #(
		.INIT('h2)
	) name4222 (
		\u4_u0_buf0_orig_reg[26]/P0001 ,
		\u4_u0_dma_out_cnt_reg[7]/P0001 ,
		_w5972_
	);
	LUT4 #(
		.INIT('h08ce)
	) name4223 (
		\u4_u0_buf0_orig_reg[26]/P0001 ,
		\u4_u0_buf0_orig_reg[27]/P0001 ,
		\u4_u0_dma_out_cnt_reg[7]/P0001 ,
		\u4_u0_dma_out_cnt_reg[8]/P0001 ,
		_w5973_
	);
	LUT2 #(
		.INIT('h2)
	) name4224 (
		\u4_u0_buf0_orig_reg[25]/P0001 ,
		\u4_u0_dma_out_cnt_reg[6]/P0001 ,
		_w5974_
	);
	LUT4 #(
		.INIT('h5010)
	) name4225 (
		\u4_u0_buf0_orig_reg[24]/P0001 ,
		\u4_u0_buf0_orig_reg[25]/P0001 ,
		\u4_u0_dma_out_cnt_reg[5]/P0001 ,
		\u4_u0_dma_out_cnt_reg[6]/P0001 ,
		_w5975_
	);
	LUT4 #(
		.INIT('h8caf)
	) name4226 (
		\u4_u0_buf0_orig_reg[22]/P0001 ,
		\u4_u0_buf0_orig_reg[23]/P0001 ,
		\u4_u0_dma_out_cnt_reg[3]/P0001 ,
		\u4_u0_dma_out_cnt_reg[4]/P0001 ,
		_w5976_
	);
	LUT4 #(
		.INIT('h080a)
	) name4227 (
		\u4_u0_buf0_orig_reg[22]/P0001 ,
		\u4_u0_buf0_orig_reg[23]/P0001 ,
		\u4_u0_dma_out_cnt_reg[3]/P0001 ,
		\u4_u0_dma_out_cnt_reg[4]/P0001 ,
		_w5977_
	);
	LUT4 #(
		.INIT('h8caf)
	) name4228 (
		\u4_u0_buf0_orig_reg[19]/P0001 ,
		\u4_u0_buf0_orig_reg[20]/P0001 ,
		\u4_u0_dma_in_cnt_reg[0]/P0001 ,
		\u4_u0_dma_out_cnt_reg[1]/P0001 ,
		_w5978_
	);
	LUT4 #(
		.INIT('hf531)
	) name4229 (
		\u4_u0_buf0_orig_reg[20]/P0001 ,
		\u4_u0_buf0_orig_reg[21]/P0001 ,
		\u4_u0_dma_out_cnt_reg[1]/P0001 ,
		\u4_u0_dma_out_cnt_reg[2]/P0001 ,
		_w5979_
	);
	LUT2 #(
		.INIT('h4)
	) name4230 (
		\u4_u0_buf0_orig_reg[21]/P0001 ,
		\u4_u0_dma_out_cnt_reg[2]/P0001 ,
		_w5980_
	);
	LUT4 #(
		.INIT('h008a)
	) name4231 (
		_w5976_,
		_w5978_,
		_w5979_,
		_w5980_,
		_w5981_
	);
	LUT2 #(
		.INIT('h2)
	) name4232 (
		\u4_u0_buf0_orig_reg[23]/P0001 ,
		\u4_u0_dma_out_cnt_reg[4]/P0001 ,
		_w5982_
	);
	LUT4 #(
		.INIT('hf531)
	) name4233 (
		\u4_u0_buf0_orig_reg[23]/P0001 ,
		\u4_u0_buf0_orig_reg[24]/P0001 ,
		\u4_u0_dma_out_cnt_reg[4]/P0001 ,
		\u4_u0_dma_out_cnt_reg[5]/P0001 ,
		_w5983_
	);
	LUT2 #(
		.INIT('h4)
	) name4234 (
		_w5974_,
		_w5983_,
		_w5984_
	);
	LUT4 #(
		.INIT('h5455)
	) name4235 (
		_w5975_,
		_w5977_,
		_w5981_,
		_w5984_,
		_w5985_
	);
	LUT4 #(
		.INIT('h8caf)
	) name4236 (
		\u4_u0_buf0_orig_reg[25]/P0001 ,
		\u4_u0_buf0_orig_reg[26]/P0001 ,
		\u4_u0_dma_out_cnt_reg[6]/P0001 ,
		\u4_u0_dma_out_cnt_reg[7]/P0001 ,
		_w5986_
	);
	LUT2 #(
		.INIT('h4)
	) name4237 (
		_w5971_,
		_w5986_,
		_w5987_
	);
	LUT4 #(
		.INIT('h5444)
	) name4238 (
		_w5970_,
		_w5973_,
		_w5985_,
		_w5987_,
		_w5988_
	);
	LUT2 #(
		.INIT('h2)
	) name4239 (
		\u4_u0_buf0_orig_reg[29]/NET0131 ,
		\u4_u0_dma_out_cnt_reg[10]/P0001 ,
		_w5989_
	);
	LUT2 #(
		.INIT('h9)
	) name4240 (
		\u4_u0_buf0_orig_reg[29]/NET0131 ,
		\u4_u0_dma_out_cnt_reg[10]/P0001 ,
		_w5990_
	);
	LUT2 #(
		.INIT('h2)
	) name4241 (
		\u4_u0_buf0_orig_reg[28]/P0001 ,
		\u4_u0_dma_out_cnt_reg[9]/P0001 ,
		_w5991_
	);
	LUT4 #(
		.INIT('h283c)
	) name4242 (
		\u4_u0_buf0_orig_reg[28]/P0001 ,
		\u4_u0_buf0_orig_reg[29]/NET0131 ,
		\u4_u0_dma_out_cnt_reg[10]/P0001 ,
		\u4_u0_dma_out_cnt_reg[9]/P0001 ,
		_w5992_
	);
	LUT4 #(
		.INIT('hea00)
	) name4243 (
		_w5973_,
		_w5985_,
		_w5987_,
		_w5992_,
		_w5993_
	);
	LUT4 #(
		.INIT('hff34)
	) name4244 (
		_w5988_,
		_w5990_,
		_w5991_,
		_w5993_,
		_w5994_
	);
	LUT2 #(
		.INIT('h4)
	) name4245 (
		\u4_u1_buf0_orig_reg[28]/P0001 ,
		\u4_u1_dma_out_cnt_reg[9]/P0001 ,
		_w5995_
	);
	LUT2 #(
		.INIT('h4)
	) name4246 (
		\u4_u1_buf0_orig_reg[27]/P0001 ,
		\u4_u1_dma_out_cnt_reg[8]/P0001 ,
		_w5996_
	);
	LUT2 #(
		.INIT('h2)
	) name4247 (
		\u4_u1_buf0_orig_reg[26]/P0001 ,
		\u4_u1_dma_out_cnt_reg[7]/P0001 ,
		_w5997_
	);
	LUT4 #(
		.INIT('h08ce)
	) name4248 (
		\u4_u1_buf0_orig_reg[26]/P0001 ,
		\u4_u1_buf0_orig_reg[27]/P0001 ,
		\u4_u1_dma_out_cnt_reg[7]/P0001 ,
		\u4_u1_dma_out_cnt_reg[8]/P0001 ,
		_w5998_
	);
	LUT2 #(
		.INIT('h2)
	) name4249 (
		\u4_u1_buf0_orig_reg[25]/P0001 ,
		\u4_u1_dma_out_cnt_reg[6]/P0001 ,
		_w5999_
	);
	LUT4 #(
		.INIT('h5010)
	) name4250 (
		\u4_u1_buf0_orig_reg[24]/P0001 ,
		\u4_u1_buf0_orig_reg[25]/P0001 ,
		\u4_u1_dma_out_cnt_reg[5]/P0001 ,
		\u4_u1_dma_out_cnt_reg[6]/P0001 ,
		_w6000_
	);
	LUT4 #(
		.INIT('h8caf)
	) name4251 (
		\u4_u1_buf0_orig_reg[22]/P0001 ,
		\u4_u1_buf0_orig_reg[23]/P0001 ,
		\u4_u1_dma_out_cnt_reg[3]/P0001 ,
		\u4_u1_dma_out_cnt_reg[4]/P0001 ,
		_w6001_
	);
	LUT4 #(
		.INIT('h080a)
	) name4252 (
		\u4_u1_buf0_orig_reg[22]/P0001 ,
		\u4_u1_buf0_orig_reg[23]/P0001 ,
		\u4_u1_dma_out_cnt_reg[3]/P0001 ,
		\u4_u1_dma_out_cnt_reg[4]/P0001 ,
		_w6002_
	);
	LUT4 #(
		.INIT('h8caf)
	) name4253 (
		\u4_u1_buf0_orig_reg[19]/P0001 ,
		\u4_u1_buf0_orig_reg[20]/P0001 ,
		\u4_u1_dma_in_cnt_reg[0]/P0001 ,
		\u4_u1_dma_out_cnt_reg[1]/P0001 ,
		_w6003_
	);
	LUT4 #(
		.INIT('hf531)
	) name4254 (
		\u4_u1_buf0_orig_reg[20]/P0001 ,
		\u4_u1_buf0_orig_reg[21]/P0001 ,
		\u4_u1_dma_out_cnt_reg[1]/P0001 ,
		\u4_u1_dma_out_cnt_reg[2]/P0001 ,
		_w6004_
	);
	LUT2 #(
		.INIT('h4)
	) name4255 (
		\u4_u1_buf0_orig_reg[21]/P0001 ,
		\u4_u1_dma_out_cnt_reg[2]/P0001 ,
		_w6005_
	);
	LUT4 #(
		.INIT('h008a)
	) name4256 (
		_w6001_,
		_w6003_,
		_w6004_,
		_w6005_,
		_w6006_
	);
	LUT2 #(
		.INIT('h2)
	) name4257 (
		\u4_u1_buf0_orig_reg[23]/P0001 ,
		\u4_u1_dma_out_cnt_reg[4]/P0001 ,
		_w6007_
	);
	LUT4 #(
		.INIT('hf531)
	) name4258 (
		\u4_u1_buf0_orig_reg[23]/P0001 ,
		\u4_u1_buf0_orig_reg[24]/P0001 ,
		\u4_u1_dma_out_cnt_reg[4]/P0001 ,
		\u4_u1_dma_out_cnt_reg[5]/P0001 ,
		_w6008_
	);
	LUT2 #(
		.INIT('h4)
	) name4259 (
		_w5999_,
		_w6008_,
		_w6009_
	);
	LUT4 #(
		.INIT('h5455)
	) name4260 (
		_w6000_,
		_w6002_,
		_w6006_,
		_w6009_,
		_w6010_
	);
	LUT4 #(
		.INIT('h8caf)
	) name4261 (
		\u4_u1_buf0_orig_reg[25]/P0001 ,
		\u4_u1_buf0_orig_reg[26]/P0001 ,
		\u4_u1_dma_out_cnt_reg[6]/P0001 ,
		\u4_u1_dma_out_cnt_reg[7]/P0001 ,
		_w6011_
	);
	LUT2 #(
		.INIT('h4)
	) name4262 (
		_w5996_,
		_w6011_,
		_w6012_
	);
	LUT4 #(
		.INIT('h5444)
	) name4263 (
		_w5995_,
		_w5998_,
		_w6010_,
		_w6012_,
		_w6013_
	);
	LUT2 #(
		.INIT('h2)
	) name4264 (
		\u4_u1_buf0_orig_reg[29]/NET0131 ,
		\u4_u1_dma_out_cnt_reg[10]/P0001 ,
		_w6014_
	);
	LUT2 #(
		.INIT('h9)
	) name4265 (
		\u4_u1_buf0_orig_reg[29]/NET0131 ,
		\u4_u1_dma_out_cnt_reg[10]/P0001 ,
		_w6015_
	);
	LUT2 #(
		.INIT('h2)
	) name4266 (
		\u4_u1_buf0_orig_reg[28]/P0001 ,
		\u4_u1_dma_out_cnt_reg[9]/P0001 ,
		_w6016_
	);
	LUT4 #(
		.INIT('h283c)
	) name4267 (
		\u4_u1_buf0_orig_reg[28]/P0001 ,
		\u4_u1_buf0_orig_reg[29]/NET0131 ,
		\u4_u1_dma_out_cnt_reg[10]/P0001 ,
		\u4_u1_dma_out_cnt_reg[9]/P0001 ,
		_w6017_
	);
	LUT4 #(
		.INIT('hea00)
	) name4268 (
		_w5998_,
		_w6010_,
		_w6012_,
		_w6017_,
		_w6018_
	);
	LUT4 #(
		.INIT('hff34)
	) name4269 (
		_w6013_,
		_w6015_,
		_w6016_,
		_w6018_,
		_w6019_
	);
	LUT2 #(
		.INIT('h4)
	) name4270 (
		\u4_u2_buf0_orig_reg[28]/P0001 ,
		\u4_u2_dma_out_cnt_reg[9]/P0001 ,
		_w6020_
	);
	LUT2 #(
		.INIT('h4)
	) name4271 (
		\u4_u2_buf0_orig_reg[27]/P0001 ,
		\u4_u2_dma_out_cnt_reg[8]/P0001 ,
		_w6021_
	);
	LUT2 #(
		.INIT('h2)
	) name4272 (
		\u4_u2_buf0_orig_reg[26]/P0001 ,
		\u4_u2_dma_out_cnt_reg[7]/P0001 ,
		_w6022_
	);
	LUT4 #(
		.INIT('h08ce)
	) name4273 (
		\u4_u2_buf0_orig_reg[26]/P0001 ,
		\u4_u2_buf0_orig_reg[27]/P0001 ,
		\u4_u2_dma_out_cnt_reg[7]/P0001 ,
		\u4_u2_dma_out_cnt_reg[8]/P0001 ,
		_w6023_
	);
	LUT2 #(
		.INIT('h2)
	) name4274 (
		\u4_u2_buf0_orig_reg[25]/P0001 ,
		\u4_u2_dma_out_cnt_reg[6]/P0001 ,
		_w6024_
	);
	LUT4 #(
		.INIT('h5010)
	) name4275 (
		\u4_u2_buf0_orig_reg[24]/P0001 ,
		\u4_u2_buf0_orig_reg[25]/P0001 ,
		\u4_u2_dma_out_cnt_reg[5]/P0001 ,
		\u4_u2_dma_out_cnt_reg[6]/P0001 ,
		_w6025_
	);
	LUT4 #(
		.INIT('h8caf)
	) name4276 (
		\u4_u2_buf0_orig_reg[22]/P0001 ,
		\u4_u2_buf0_orig_reg[23]/P0001 ,
		\u4_u2_dma_out_cnt_reg[3]/P0001 ,
		\u4_u2_dma_out_cnt_reg[4]/P0001 ,
		_w6026_
	);
	LUT4 #(
		.INIT('h080a)
	) name4277 (
		\u4_u2_buf0_orig_reg[22]/P0001 ,
		\u4_u2_buf0_orig_reg[23]/P0001 ,
		\u4_u2_dma_out_cnt_reg[3]/P0001 ,
		\u4_u2_dma_out_cnt_reg[4]/P0001 ,
		_w6027_
	);
	LUT4 #(
		.INIT('h8caf)
	) name4278 (
		\u4_u2_buf0_orig_reg[19]/P0001 ,
		\u4_u2_buf0_orig_reg[20]/P0001 ,
		\u4_u2_dma_in_cnt_reg[0]/P0001 ,
		\u4_u2_dma_out_cnt_reg[1]/P0001 ,
		_w6028_
	);
	LUT4 #(
		.INIT('hf531)
	) name4279 (
		\u4_u2_buf0_orig_reg[20]/P0001 ,
		\u4_u2_buf0_orig_reg[21]/P0001 ,
		\u4_u2_dma_out_cnt_reg[1]/P0001 ,
		\u4_u2_dma_out_cnt_reg[2]/P0001 ,
		_w6029_
	);
	LUT2 #(
		.INIT('h4)
	) name4280 (
		\u4_u2_buf0_orig_reg[21]/P0001 ,
		\u4_u2_dma_out_cnt_reg[2]/P0001 ,
		_w6030_
	);
	LUT4 #(
		.INIT('h008a)
	) name4281 (
		_w6026_,
		_w6028_,
		_w6029_,
		_w6030_,
		_w6031_
	);
	LUT2 #(
		.INIT('h2)
	) name4282 (
		\u4_u2_buf0_orig_reg[23]/P0001 ,
		\u4_u2_dma_out_cnt_reg[4]/P0001 ,
		_w6032_
	);
	LUT4 #(
		.INIT('hf531)
	) name4283 (
		\u4_u2_buf0_orig_reg[23]/P0001 ,
		\u4_u2_buf0_orig_reg[24]/P0001 ,
		\u4_u2_dma_out_cnt_reg[4]/P0001 ,
		\u4_u2_dma_out_cnt_reg[5]/P0001 ,
		_w6033_
	);
	LUT2 #(
		.INIT('h4)
	) name4284 (
		_w6024_,
		_w6033_,
		_w6034_
	);
	LUT4 #(
		.INIT('h5455)
	) name4285 (
		_w6025_,
		_w6027_,
		_w6031_,
		_w6034_,
		_w6035_
	);
	LUT4 #(
		.INIT('h8caf)
	) name4286 (
		\u4_u2_buf0_orig_reg[25]/P0001 ,
		\u4_u2_buf0_orig_reg[26]/P0001 ,
		\u4_u2_dma_out_cnt_reg[6]/P0001 ,
		\u4_u2_dma_out_cnt_reg[7]/P0001 ,
		_w6036_
	);
	LUT2 #(
		.INIT('h4)
	) name4287 (
		_w6021_,
		_w6036_,
		_w6037_
	);
	LUT4 #(
		.INIT('h5444)
	) name4288 (
		_w6020_,
		_w6023_,
		_w6035_,
		_w6037_,
		_w6038_
	);
	LUT2 #(
		.INIT('h9)
	) name4289 (
		\u4_u2_buf0_orig_reg[29]/NET0131 ,
		\u4_u2_dma_out_cnt_reg[10]/P0001 ,
		_w6039_
	);
	LUT2 #(
		.INIT('h2)
	) name4290 (
		\u4_u2_buf0_orig_reg[28]/P0001 ,
		\u4_u2_dma_out_cnt_reg[9]/P0001 ,
		_w6040_
	);
	LUT4 #(
		.INIT('h283c)
	) name4291 (
		\u4_u2_buf0_orig_reg[28]/P0001 ,
		\u4_u2_buf0_orig_reg[29]/NET0131 ,
		\u4_u2_dma_out_cnt_reg[10]/P0001 ,
		\u4_u2_dma_out_cnt_reg[9]/P0001 ,
		_w6041_
	);
	LUT4 #(
		.INIT('hea00)
	) name4292 (
		_w6023_,
		_w6035_,
		_w6037_,
		_w6041_,
		_w6042_
	);
	LUT4 #(
		.INIT('hff34)
	) name4293 (
		_w6038_,
		_w6039_,
		_w6040_,
		_w6042_,
		_w6043_
	);
	LUT2 #(
		.INIT('h9)
	) name4294 (
		\u4_u3_csr0_reg[8]/P0001 ,
		\u4_u3_dma_in_cnt_reg[6]/P0001 ,
		_w6044_
	);
	LUT2 #(
		.INIT('h8)
	) name4295 (
		_w4569_,
		_w6044_,
		_w6045_
	);
	LUT2 #(
		.INIT('h4)
	) name4296 (
		_w4564_,
		_w4569_,
		_w6046_
	);
	LUT3 #(
		.INIT('h13)
	) name4297 (
		_w4561_,
		_w6045_,
		_w6046_,
		_w6047_
	);
	LUT3 #(
		.INIT('h15)
	) name4298 (
		\u4_u3_dma_in_cnt_reg[6]/P0001 ,
		_w4399_,
		_w5681_,
		_w6048_
	);
	LUT3 #(
		.INIT('h2a)
	) name4299 (
		\u4_u3_r5_reg/NET0131 ,
		_w4398_,
		_w4399_,
		_w6049_
	);
	LUT2 #(
		.INIT('h4)
	) name4300 (
		_w4564_,
		_w6044_,
		_w6050_
	);
	LUT4 #(
		.INIT('h45cf)
	) name4301 (
		_w4561_,
		_w6048_,
		_w6049_,
		_w6050_,
		_w6051_
	);
	LUT4 #(
		.INIT('h0001)
	) name4302 (
		\u1_u3_buf0_rl_reg/P0001 ,
		\u1_u3_buf0_set_reg/P0001 ,
		\u4_u3_dma_in_cnt_reg[6]/P0001 ,
		\u4_u3_set_r_reg/P0001 ,
		_w6052_
	);
	LUT3 #(
		.INIT('h0e)
	) name4303 (
		\u4_u3_dma_in_cnt_reg[6]/P0001 ,
		\u4_u3_ep_match_r_reg/P0001 ,
		\u4_u3_r5_reg/NET0131 ,
		_w6053_
	);
	LUT2 #(
		.INIT('h4)
	) name4304 (
		_w6052_,
		_w6053_,
		_w6054_
	);
	LUT4 #(
		.INIT('haa20)
	) name4305 (
		\u4_u3_csr1_reg[0]/P0001 ,
		_w6048_,
		_w6049_,
		_w6054_,
		_w6055_
	);
	LUT3 #(
		.INIT('hb0)
	) name4306 (
		_w6047_,
		_w6051_,
		_w6055_,
		_w6056_
	);
	LUT4 #(
		.INIT('h0100)
	) name4307 (
		\u4_u3_dma_out_cnt_reg[4]/P0001 ,
		\u4_u3_dma_out_cnt_reg[5]/P0001 ,
		\u4_u3_dma_out_cnt_reg[6]/P0001 ,
		\u4_u3_r5_reg/NET0131 ,
		_w6057_
	);
	LUT3 #(
		.INIT('h80)
	) name4308 (
		\u4_u3_csr1_reg[0]/P0001 ,
		_w4652_,
		_w6057_,
		_w6058_
	);
	LUT3 #(
		.INIT('h80)
	) name4309 (
		\u4_u3_csr1_reg[0]/P0001 ,
		\u4_u3_dma_out_cnt_reg[6]/P0001 ,
		\u4_u3_r5_reg/NET0131 ,
		_w6059_
	);
	LUT3 #(
		.INIT('h70)
	) name4310 (
		_w4652_,
		_w4953_,
		_w6059_,
		_w6060_
	);
	LUT2 #(
		.INIT('h1)
	) name4311 (
		_w6058_,
		_w6060_,
		_w6061_
	);
	LUT2 #(
		.INIT('h6)
	) name4312 (
		\u4_u3_csr0_reg[8]/P0001 ,
		\u4_u3_dma_out_cnt_reg[6]/P0001 ,
		_w6062_
	);
	LUT4 #(
		.INIT('h8020)
	) name4313 (
		\u4_u3_csr0_reg[7]/P0001 ,
		\u4_u3_csr0_reg[8]/P0001 ,
		\u4_u3_dma_out_cnt_reg[5]/P0001 ,
		\u4_u3_dma_out_cnt_reg[6]/P0001 ,
		_w6063_
	);
	LUT2 #(
		.INIT('h2)
	) name4314 (
		_w4674_,
		_w6062_,
		_w6064_
	);
	LUT4 #(
		.INIT('h0e0f)
	) name4315 (
		_w4667_,
		_w4672_,
		_w6063_,
		_w6064_,
		_w6065_
	);
	LUT4 #(
		.INIT('h134c)
	) name4316 (
		\u4_u3_csr0_reg[7]/P0001 ,
		\u4_u3_csr0_reg[8]/P0001 ,
		\u4_u3_dma_out_cnt_reg[5]/P0001 ,
		\u4_u3_dma_out_cnt_reg[6]/P0001 ,
		_w6066_
	);
	LUT4 #(
		.INIT('hef00)
	) name4317 (
		_w4667_,
		_w4672_,
		_w4674_,
		_w6066_,
		_w6067_
	);
	LUT4 #(
		.INIT('h0001)
	) name4318 (
		\u1_u3_buf0_rl_reg/P0001 ,
		\u1_u3_buf0_set_reg/P0001 ,
		\u4_u3_dma_out_cnt_reg[6]/P0001 ,
		\u4_u3_set_r_reg/P0001 ,
		_w6068_
	);
	LUT3 #(
		.INIT('ha8)
	) name4319 (
		\u4_u3_csr1_reg[0]/P0001 ,
		\u4_u3_dma_out_cnt_reg[6]/P0001 ,
		\u4_u3_ep_match_r_reg/P0001 ,
		_w6069_
	);
	LUT3 #(
		.INIT('h10)
	) name4320 (
		\u4_u3_r5_reg/NET0131 ,
		_w6068_,
		_w6069_,
		_w6070_
	);
	LUT4 #(
		.INIT('hf700)
	) name4321 (
		_w4569_,
		_w6065_,
		_w6067_,
		_w6070_,
		_w6071_
	);
	LUT2 #(
		.INIT('hd)
	) name4322 (
		_w6061_,
		_w6071_,
		_w6072_
	);
	LUT2 #(
		.INIT('h9)
	) name4323 (
		\u4_u0_csr0_reg[8]/P0001 ,
		\u4_u0_dma_in_cnt_reg[6]/P0001 ,
		_w6073_
	);
	LUT2 #(
		.INIT('h8)
	) name4324 (
		_w4592_,
		_w6073_,
		_w6074_
	);
	LUT2 #(
		.INIT('h4)
	) name4325 (
		_w4587_,
		_w4592_,
		_w6075_
	);
	LUT3 #(
		.INIT('h13)
	) name4326 (
		_w4584_,
		_w6074_,
		_w6075_,
		_w6076_
	);
	LUT3 #(
		.INIT('h15)
	) name4327 (
		\u4_u0_dma_in_cnt_reg[6]/P0001 ,
		_w4431_,
		_w5696_,
		_w6077_
	);
	LUT3 #(
		.INIT('h2a)
	) name4328 (
		\u4_u0_r5_reg/NET0131 ,
		_w4430_,
		_w4431_,
		_w6078_
	);
	LUT2 #(
		.INIT('h4)
	) name4329 (
		_w4587_,
		_w6073_,
		_w6079_
	);
	LUT4 #(
		.INIT('h45cf)
	) name4330 (
		_w4584_,
		_w6077_,
		_w6078_,
		_w6079_,
		_w6080_
	);
	LUT4 #(
		.INIT('h0001)
	) name4331 (
		\u1_u3_buf0_rl_reg/P0001 ,
		\u1_u3_buf0_set_reg/P0001 ,
		\u4_u0_dma_in_cnt_reg[6]/P0001 ,
		\u4_u0_set_r_reg/P0001 ,
		_w6081_
	);
	LUT3 #(
		.INIT('h0e)
	) name4332 (
		\u4_u0_dma_in_cnt_reg[6]/P0001 ,
		\u4_u0_ep_match_r_reg/P0001 ,
		\u4_u0_r5_reg/NET0131 ,
		_w6082_
	);
	LUT2 #(
		.INIT('h4)
	) name4333 (
		_w6081_,
		_w6082_,
		_w6083_
	);
	LUT4 #(
		.INIT('haa20)
	) name4334 (
		\u4_u0_csr1_reg[0]/P0001 ,
		_w6077_,
		_w6078_,
		_w6083_,
		_w6084_
	);
	LUT3 #(
		.INIT('hb0)
	) name4335 (
		_w6076_,
		_w6080_,
		_w6084_,
		_w6085_
	);
	LUT4 #(
		.INIT('hb777)
	) name4336 (
		\u4_u0_dma_out_cnt_reg[6]/P0001 ,
		\u4_u0_r5_reg/NET0131 ,
		_w4683_,
		_w4983_,
		_w6086_
	);
	LUT4 #(
		.INIT('h0001)
	) name4337 (
		\u1_u3_buf0_rl_reg/P0001 ,
		\u1_u3_buf0_set_reg/P0001 ,
		\u4_u0_dma_out_cnt_reg[6]/P0001 ,
		\u4_u0_set_r_reg/P0001 ,
		_w6087_
	);
	LUT3 #(
		.INIT('h0e)
	) name4338 (
		\u4_u0_dma_out_cnt_reg[6]/P0001 ,
		\u4_u0_ep_match_r_reg/P0001 ,
		\u4_u0_r5_reg/NET0131 ,
		_w6088_
	);
	LUT2 #(
		.INIT('h4)
	) name4339 (
		_w6087_,
		_w6088_,
		_w6089_
	);
	LUT2 #(
		.INIT('h2)
	) name4340 (
		_w6086_,
		_w6089_,
		_w6090_
	);
	LUT2 #(
		.INIT('h6)
	) name4341 (
		\u4_u0_csr0_reg[8]/P0001 ,
		\u4_u0_dma_out_cnt_reg[6]/P0001 ,
		_w6091_
	);
	LUT4 #(
		.INIT('h8020)
	) name4342 (
		\u4_u0_csr0_reg[7]/P0001 ,
		\u4_u0_csr0_reg[8]/P0001 ,
		\u4_u0_dma_out_cnt_reg[5]/P0001 ,
		\u4_u0_dma_out_cnt_reg[6]/P0001 ,
		_w6092_
	);
	LUT2 #(
		.INIT('h2)
	) name4343 (
		_w4704_,
		_w6091_,
		_w6093_
	);
	LUT4 #(
		.INIT('h0e0f)
	) name4344 (
		_w4697_,
		_w4702_,
		_w6092_,
		_w6093_,
		_w6094_
	);
	LUT4 #(
		.INIT('h134c)
	) name4345 (
		\u4_u0_csr0_reg[7]/P0001 ,
		\u4_u0_csr0_reg[8]/P0001 ,
		\u4_u0_dma_out_cnt_reg[5]/P0001 ,
		\u4_u0_dma_out_cnt_reg[6]/P0001 ,
		_w6095_
	);
	LUT4 #(
		.INIT('hef00)
	) name4346 (
		_w4697_,
		_w4702_,
		_w4704_,
		_w6095_,
		_w6096_
	);
	LUT2 #(
		.INIT('h8)
	) name4347 (
		_w4592_,
		_w6086_,
		_w6097_
	);
	LUT4 #(
		.INIT('h5155)
	) name4348 (
		_w6090_,
		_w6094_,
		_w6096_,
		_w6097_,
		_w6098_
	);
	LUT2 #(
		.INIT('h8)
	) name4349 (
		\u4_u0_csr1_reg[0]/P0001 ,
		_w6098_,
		_w6099_
	);
	LUT3 #(
		.INIT('h2a)
	) name4350 (
		\u4_u1_r5_reg/NET0131 ,
		_w4447_,
		_w4448_,
		_w6100_
	);
	LUT2 #(
		.INIT('h8)
	) name4351 (
		\u4_u1_csr1_reg[0]/P0001 ,
		\u4_u1_dma_in_cnt_reg[6]/P0001 ,
		_w6101_
	);
	LUT3 #(
		.INIT('h80)
	) name4352 (
		\u4_u1_csr1_reg[0]/P0001 ,
		\u4_u1_dma_in_cnt_reg[4]/P0001 ,
		\u4_u1_dma_in_cnt_reg[5]/P0001 ,
		_w6102_
	);
	LUT3 #(
		.INIT('h13)
	) name4353 (
		_w4448_,
		_w6101_,
		_w6102_,
		_w6103_
	);
	LUT2 #(
		.INIT('h2)
	) name4354 (
		_w6100_,
		_w6103_,
		_w6104_
	);
	LUT2 #(
		.INIT('h9)
	) name4355 (
		\u4_u1_csr0_reg[8]/P0001 ,
		\u4_u1_dma_in_cnt_reg[6]/P0001 ,
		_w6105_
	);
	LUT4 #(
		.INIT('h31c4)
	) name4356 (
		\u4_u1_csr0_reg[7]/P0001 ,
		\u4_u1_csr0_reg[8]/P0001 ,
		\u4_u1_dma_in_cnt_reg[5]/P0001 ,
		\u4_u1_dma_in_cnt_reg[6]/P0001 ,
		_w6106_
	);
	LUT4 #(
		.INIT('hef00)
	) name4357 (
		_w4463_,
		_w4468_,
		_w4469_,
		_w6106_,
		_w6107_
	);
	LUT4 #(
		.INIT('h0802)
	) name4358 (
		\u4_u1_csr0_reg[7]/P0001 ,
		\u4_u1_csr0_reg[8]/P0001 ,
		\u4_u1_dma_in_cnt_reg[5]/P0001 ,
		\u4_u1_dma_in_cnt_reg[6]/P0001 ,
		_w6108_
	);
	LUT2 #(
		.INIT('h8)
	) name4359 (
		_w4469_,
		_w6105_,
		_w6109_
	);
	LUT4 #(
		.INIT('h0e0f)
	) name4360 (
		_w4463_,
		_w4468_,
		_w6108_,
		_w6109_,
		_w6110_
	);
	LUT4 #(
		.INIT('h0001)
	) name4361 (
		\u1_u3_buf0_rl_reg/P0001 ,
		\u1_u3_buf0_set_reg/P0001 ,
		\u4_u1_dma_in_cnt_reg[6]/P0001 ,
		\u4_u1_set_r_reg/P0001 ,
		_w6111_
	);
	LUT3 #(
		.INIT('ha8)
	) name4362 (
		\u4_u1_csr1_reg[0]/P0001 ,
		\u4_u1_dma_in_cnt_reg[6]/P0001 ,
		\u4_u1_ep_match_r_reg/P0001 ,
		_w6112_
	);
	LUT3 #(
		.INIT('h10)
	) name4363 (
		\u4_u1_r5_reg/NET0131 ,
		_w6111_,
		_w6112_,
		_w6113_
	);
	LUT4 #(
		.INIT('hdf00)
	) name4364 (
		_w4454_,
		_w6107_,
		_w6110_,
		_w6113_,
		_w6114_
	);
	LUT2 #(
		.INIT('he)
	) name4365 (
		_w6104_,
		_w6114_,
		_w6115_
	);
	LUT4 #(
		.INIT('h0100)
	) name4366 (
		\u4_u1_dma_out_cnt_reg[4]/P0001 ,
		\u4_u1_dma_out_cnt_reg[5]/P0001 ,
		\u4_u1_dma_out_cnt_reg[6]/P0001 ,
		\u4_u1_r5_reg/NET0131 ,
		_w6116_
	);
	LUT3 #(
		.INIT('h80)
	) name4367 (
		\u4_u1_csr1_reg[0]/P0001 ,
		_w4713_,
		_w6116_,
		_w6117_
	);
	LUT3 #(
		.INIT('h80)
	) name4368 (
		\u4_u1_csr1_reg[0]/P0001 ,
		\u4_u1_dma_out_cnt_reg[6]/P0001 ,
		\u4_u1_r5_reg/NET0131 ,
		_w6118_
	);
	LUT3 #(
		.INIT('h70)
	) name4369 (
		_w4713_,
		_w5017_,
		_w6118_,
		_w6119_
	);
	LUT2 #(
		.INIT('h1)
	) name4370 (
		_w6117_,
		_w6119_,
		_w6120_
	);
	LUT2 #(
		.INIT('h6)
	) name4371 (
		\u4_u1_csr0_reg[8]/P0001 ,
		\u4_u1_dma_out_cnt_reg[6]/P0001 ,
		_w6121_
	);
	LUT4 #(
		.INIT('h8020)
	) name4372 (
		\u4_u1_csr0_reg[7]/P0001 ,
		\u4_u1_csr0_reg[8]/P0001 ,
		\u4_u1_dma_out_cnt_reg[5]/P0001 ,
		\u4_u1_dma_out_cnt_reg[6]/P0001 ,
		_w6122_
	);
	LUT2 #(
		.INIT('h2)
	) name4373 (
		_w4735_,
		_w6121_,
		_w6123_
	);
	LUT4 #(
		.INIT('h0e0f)
	) name4374 (
		_w4728_,
		_w4733_,
		_w6122_,
		_w6123_,
		_w6124_
	);
	LUT4 #(
		.INIT('h134c)
	) name4375 (
		\u4_u1_csr0_reg[7]/P0001 ,
		\u4_u1_csr0_reg[8]/P0001 ,
		\u4_u1_dma_out_cnt_reg[5]/P0001 ,
		\u4_u1_dma_out_cnt_reg[6]/P0001 ,
		_w6125_
	);
	LUT4 #(
		.INIT('hef00)
	) name4376 (
		_w4728_,
		_w4733_,
		_w4735_,
		_w6125_,
		_w6126_
	);
	LUT4 #(
		.INIT('h0001)
	) name4377 (
		\u1_u3_buf0_rl_reg/P0001 ,
		\u1_u3_buf0_set_reg/P0001 ,
		\u4_u1_dma_out_cnt_reg[6]/P0001 ,
		\u4_u1_set_r_reg/P0001 ,
		_w6127_
	);
	LUT3 #(
		.INIT('ha8)
	) name4378 (
		\u4_u1_csr1_reg[0]/P0001 ,
		\u4_u1_dma_out_cnt_reg[6]/P0001 ,
		\u4_u1_ep_match_r_reg/P0001 ,
		_w6128_
	);
	LUT3 #(
		.INIT('h10)
	) name4379 (
		\u4_u1_r5_reg/NET0131 ,
		_w6127_,
		_w6128_,
		_w6129_
	);
	LUT4 #(
		.INIT('hf700)
	) name4380 (
		_w4454_,
		_w6124_,
		_w6126_,
		_w6129_,
		_w6130_
	);
	LUT2 #(
		.INIT('hd)
	) name4381 (
		_w6120_,
		_w6130_,
		_w6131_
	);
	LUT3 #(
		.INIT('h15)
	) name4382 (
		\u4_u2_dma_in_cnt_reg[6]/P0001 ,
		_w4505_,
		_w5729_,
		_w6132_
	);
	LUT2 #(
		.INIT('h8)
	) name4383 (
		\u4_u2_csr1_reg[0]/P0001 ,
		\u4_u2_r5_reg/NET0131 ,
		_w6133_
	);
	LUT3 #(
		.INIT('h70)
	) name4384 (
		_w4504_,
		_w4505_,
		_w6133_,
		_w6134_
	);
	LUT4 #(
		.INIT('h0001)
	) name4385 (
		\u1_u3_buf0_rl_reg/P0001 ,
		\u1_u3_buf0_set_reg/P0001 ,
		\u4_u2_dma_in_cnt_reg[6]/P0001 ,
		\u4_u2_set_r_reg/P0001 ,
		_w6135_
	);
	LUT4 #(
		.INIT('h00a8)
	) name4386 (
		\u4_u2_csr1_reg[0]/P0001 ,
		\u4_u2_dma_in_cnt_reg[6]/P0001 ,
		\u4_u2_ep_match_r_reg/P0001 ,
		\u4_u2_r5_reg/NET0131 ,
		_w6136_
	);
	LUT2 #(
		.INIT('h4)
	) name4387 (
		_w6135_,
		_w6136_,
		_w6137_
	);
	LUT3 #(
		.INIT('h0b)
	) name4388 (
		_w6132_,
		_w6134_,
		_w6137_,
		_w6138_
	);
	LUT2 #(
		.INIT('h9)
	) name4389 (
		\u4_u2_csr0_reg[8]/P0001 ,
		\u4_u2_dma_in_cnt_reg[6]/P0001 ,
		_w6139_
	);
	LUT4 #(
		.INIT('h31c4)
	) name4390 (
		\u4_u2_csr0_reg[7]/P0001 ,
		\u4_u2_csr0_reg[8]/P0001 ,
		\u4_u2_dma_in_cnt_reg[5]/P0001 ,
		\u4_u2_dma_in_cnt_reg[6]/P0001 ,
		_w6140_
	);
	LUT4 #(
		.INIT('hef00)
	) name4391 (
		_w4491_,
		_w4496_,
		_w4497_,
		_w6140_,
		_w6141_
	);
	LUT4 #(
		.INIT('h0802)
	) name4392 (
		\u4_u2_csr0_reg[7]/P0001 ,
		\u4_u2_csr0_reg[8]/P0001 ,
		\u4_u2_dma_in_cnt_reg[5]/P0001 ,
		\u4_u2_dma_in_cnt_reg[6]/P0001 ,
		_w6142_
	);
	LUT2 #(
		.INIT('h8)
	) name4393 (
		_w4497_,
		_w6139_,
		_w6143_
	);
	LUT4 #(
		.INIT('h0e0f)
	) name4394 (
		_w4491_,
		_w4496_,
		_w6142_,
		_w6143_,
		_w6144_
	);
	LUT3 #(
		.INIT('h8a)
	) name4395 (
		_w4610_,
		_w6132_,
		_w6134_,
		_w6145_
	);
	LUT4 #(
		.INIT('h4555)
	) name4396 (
		_w6138_,
		_w6141_,
		_w6144_,
		_w6145_,
		_w6146_
	);
	LUT4 #(
		.INIT('h0100)
	) name4397 (
		\u4_u2_dma_out_cnt_reg[4]/P0001 ,
		\u4_u2_dma_out_cnt_reg[5]/P0001 ,
		\u4_u2_dma_out_cnt_reg[6]/P0001 ,
		\u4_u2_r5_reg/NET0131 ,
		_w6147_
	);
	LUT3 #(
		.INIT('h80)
	) name4398 (
		\u4_u2_csr1_reg[0]/P0001 ,
		_w4744_,
		_w6147_,
		_w6148_
	);
	LUT3 #(
		.INIT('h80)
	) name4399 (
		\u4_u2_csr1_reg[0]/P0001 ,
		\u4_u2_dma_out_cnt_reg[6]/P0001 ,
		\u4_u2_r5_reg/NET0131 ,
		_w6149_
	);
	LUT3 #(
		.INIT('h70)
	) name4400 (
		_w4744_,
		_w5047_,
		_w6149_,
		_w6150_
	);
	LUT2 #(
		.INIT('h1)
	) name4401 (
		_w6148_,
		_w6150_,
		_w6151_
	);
	LUT2 #(
		.INIT('h6)
	) name4402 (
		\u4_u2_csr0_reg[8]/P0001 ,
		\u4_u2_dma_out_cnt_reg[6]/P0001 ,
		_w6152_
	);
	LUT4 #(
		.INIT('h8020)
	) name4403 (
		\u4_u2_csr0_reg[7]/P0001 ,
		\u4_u2_csr0_reg[8]/P0001 ,
		\u4_u2_dma_out_cnt_reg[5]/P0001 ,
		\u4_u2_dma_out_cnt_reg[6]/P0001 ,
		_w6153_
	);
	LUT2 #(
		.INIT('h2)
	) name4404 (
		_w4765_,
		_w6152_,
		_w6154_
	);
	LUT4 #(
		.INIT('h0e0f)
	) name4405 (
		_w4758_,
		_w4763_,
		_w6153_,
		_w6154_,
		_w6155_
	);
	LUT4 #(
		.INIT('h134c)
	) name4406 (
		\u4_u2_csr0_reg[7]/P0001 ,
		\u4_u2_csr0_reg[8]/P0001 ,
		\u4_u2_dma_out_cnt_reg[5]/P0001 ,
		\u4_u2_dma_out_cnt_reg[6]/P0001 ,
		_w6156_
	);
	LUT4 #(
		.INIT('hef00)
	) name4407 (
		_w4758_,
		_w4763_,
		_w4765_,
		_w6156_,
		_w6157_
	);
	LUT4 #(
		.INIT('h0001)
	) name4408 (
		\u1_u3_buf0_rl_reg/P0001 ,
		\u1_u3_buf0_set_reg/P0001 ,
		\u4_u2_dma_out_cnt_reg[6]/P0001 ,
		\u4_u2_set_r_reg/P0001 ,
		_w6158_
	);
	LUT3 #(
		.INIT('ha8)
	) name4409 (
		\u4_u2_csr1_reg[0]/P0001 ,
		\u4_u2_dma_out_cnt_reg[6]/P0001 ,
		\u4_u2_ep_match_r_reg/P0001 ,
		_w6159_
	);
	LUT3 #(
		.INIT('h10)
	) name4410 (
		\u4_u2_r5_reg/NET0131 ,
		_w6158_,
		_w6159_,
		_w6160_
	);
	LUT4 #(
		.INIT('hf700)
	) name4411 (
		_w4610_,
		_w6155_,
		_w6157_,
		_w6160_,
		_w6161_
	);
	LUT2 #(
		.INIT('hd)
	) name4412 (
		_w6151_,
		_w6161_,
		_w6162_
	);
	LUT2 #(
		.INIT('h9)
	) name4413 (
		\u4_u3_csr0_reg[6]/P0001 ,
		\u4_u3_dma_in_cnt_reg[4]/P0001 ,
		_w6163_
	);
	LUT3 #(
		.INIT('h02)
	) name4414 (
		_w4389_,
		_w4560_,
		_w6163_,
		_w6164_
	);
	LUT3 #(
		.INIT('hc4)
	) name4415 (
		_w4559_,
		_w4569_,
		_w6163_,
		_w6165_
	);
	LUT3 #(
		.INIT('hb7)
	) name4416 (
		\u4_u3_dma_in_cnt_reg[4]/P0001 ,
		\u4_u3_r5_reg/NET0131 ,
		_w4399_,
		_w6166_
	);
	LUT4 #(
		.INIT('h3100)
	) name4417 (
		_w4389_,
		_w4559_,
		_w4560_,
		_w6163_,
		_w6167_
	);
	LUT4 #(
		.INIT('h0040)
	) name4418 (
		_w6164_,
		_w6165_,
		_w6166_,
		_w6167_,
		_w6168_
	);
	LUT4 #(
		.INIT('h0001)
	) name4419 (
		\u1_u3_buf0_rl_reg/P0001 ,
		\u1_u3_buf0_set_reg/P0001 ,
		\u4_u3_dma_in_cnt_reg[4]/P0001 ,
		\u4_u3_set_r_reg/P0001 ,
		_w6169_
	);
	LUT3 #(
		.INIT('h0e)
	) name4420 (
		\u4_u3_dma_in_cnt_reg[4]/P0001 ,
		\u4_u3_ep_match_r_reg/P0001 ,
		\u4_u3_r5_reg/NET0131 ,
		_w6170_
	);
	LUT2 #(
		.INIT('h4)
	) name4421 (
		_w6169_,
		_w6170_,
		_w6171_
	);
	LUT3 #(
		.INIT('ha2)
	) name4422 (
		\u4_u3_csr1_reg[0]/P0001 ,
		_w6166_,
		_w6171_,
		_w6172_
	);
	LUT2 #(
		.INIT('h4)
	) name4423 (
		_w6168_,
		_w6172_,
		_w6173_
	);
	LUT2 #(
		.INIT('h9)
	) name4424 (
		\u4_u0_csr0_reg[6]/P0001 ,
		\u4_u0_dma_in_cnt_reg[4]/P0001 ,
		_w6174_
	);
	LUT3 #(
		.INIT('hc4)
	) name4425 (
		_w4582_,
		_w4592_,
		_w6174_,
		_w6175_
	);
	LUT4 #(
		.INIT('h3100)
	) name4426 (
		_w4421_,
		_w4582_,
		_w4583_,
		_w6174_,
		_w6176_
	);
	LUT3 #(
		.INIT('h02)
	) name4427 (
		_w4421_,
		_w4583_,
		_w6174_,
		_w6177_
	);
	LUT3 #(
		.INIT('hb7)
	) name4428 (
		\u4_u0_dma_in_cnt_reg[4]/P0001 ,
		\u4_u0_r5_reg/NET0131 ,
		_w4431_,
		_w6178_
	);
	LUT4 #(
		.INIT('h0200)
	) name4429 (
		_w6175_,
		_w6176_,
		_w6177_,
		_w6178_,
		_w6179_
	);
	LUT4 #(
		.INIT('h0001)
	) name4430 (
		\u1_u3_buf0_rl_reg/P0001 ,
		\u1_u3_buf0_set_reg/P0001 ,
		\u4_u0_dma_in_cnt_reg[4]/P0001 ,
		\u4_u0_set_r_reg/P0001 ,
		_w6180_
	);
	LUT3 #(
		.INIT('h0e)
	) name4431 (
		\u4_u0_dma_in_cnt_reg[4]/P0001 ,
		\u4_u0_ep_match_r_reg/P0001 ,
		\u4_u0_r5_reg/NET0131 ,
		_w6181_
	);
	LUT2 #(
		.INIT('h4)
	) name4432 (
		_w6180_,
		_w6181_,
		_w6182_
	);
	LUT3 #(
		.INIT('ha2)
	) name4433 (
		\u4_u0_csr1_reg[0]/P0001 ,
		_w6178_,
		_w6182_,
		_w6183_
	);
	LUT2 #(
		.INIT('h4)
	) name4434 (
		_w6179_,
		_w6183_,
		_w6184_
	);
	LUT3 #(
		.INIT('hb7)
	) name4435 (
		\u4_u1_dma_in_cnt_reg[4]/P0001 ,
		\u4_u1_r5_reg/NET0131 ,
		_w4448_,
		_w6185_
	);
	LUT2 #(
		.INIT('h9)
	) name4436 (
		\u4_u1_csr0_reg[6]/P0001 ,
		\u4_u1_dma_in_cnt_reg[4]/P0001 ,
		_w6186_
	);
	LUT4 #(
		.INIT('hf531)
	) name4437 (
		\u4_u1_csr0_reg[4]/P0001 ,
		\u4_u1_csr0_reg[5]/P0001 ,
		\u4_u1_dma_in_cnt_reg[2]/P0001 ,
		\u4_u1_dma_in_cnt_reg[3]/P0001 ,
		_w6187_
	);
	LUT4 #(
		.INIT('h0b00)
	) name4438 (
		_w4465_,
		_w4466_,
		_w6186_,
		_w6187_,
		_w6188_
	);
	LUT4 #(
		.INIT('h1040)
	) name4439 (
		\u4_u1_csr0_reg[5]/P0001 ,
		\u4_u1_csr0_reg[6]/P0001 ,
		\u4_u1_dma_in_cnt_reg[3]/P0001 ,
		\u4_u1_dma_in_cnt_reg[4]/P0001 ,
		_w6189_
	);
	LUT2 #(
		.INIT('h2)
	) name4440 (
		_w4454_,
		_w6189_,
		_w6190_
	);
	LUT4 #(
		.INIT('h8c23)
	) name4441 (
		\u4_u1_csr0_reg[5]/P0001 ,
		\u4_u1_csr0_reg[6]/P0001 ,
		\u4_u1_dma_in_cnt_reg[3]/P0001 ,
		\u4_u1_dma_in_cnt_reg[4]/P0001 ,
		_w6191_
	);
	LUT4 #(
		.INIT('h4f00)
	) name4442 (
		_w4465_,
		_w4466_,
		_w6187_,
		_w6191_,
		_w6192_
	);
	LUT4 #(
		.INIT('h0020)
	) name4443 (
		_w6185_,
		_w6188_,
		_w6190_,
		_w6192_,
		_w6193_
	);
	LUT4 #(
		.INIT('h0001)
	) name4444 (
		\u1_u3_buf0_rl_reg/P0001 ,
		\u1_u3_buf0_set_reg/P0001 ,
		\u4_u1_dma_in_cnt_reg[4]/P0001 ,
		\u4_u1_set_r_reg/P0001 ,
		_w6194_
	);
	LUT3 #(
		.INIT('h0e)
	) name4445 (
		\u4_u1_dma_in_cnt_reg[4]/P0001 ,
		\u4_u1_ep_match_r_reg/P0001 ,
		\u4_u1_r5_reg/NET0131 ,
		_w6195_
	);
	LUT2 #(
		.INIT('h4)
	) name4446 (
		_w6194_,
		_w6195_,
		_w6196_
	);
	LUT3 #(
		.INIT('ha2)
	) name4447 (
		\u4_u1_csr1_reg[0]/P0001 ,
		_w6185_,
		_w6196_,
		_w6197_
	);
	LUT2 #(
		.INIT('h4)
	) name4448 (
		_w6193_,
		_w6197_,
		_w6198_
	);
	LUT3 #(
		.INIT('hb7)
	) name4449 (
		\u4_u2_dma_in_cnt_reg[4]/P0001 ,
		\u4_u2_r5_reg/NET0131 ,
		_w4505_,
		_w6199_
	);
	LUT2 #(
		.INIT('h9)
	) name4450 (
		\u4_u2_csr0_reg[6]/P0001 ,
		\u4_u2_dma_in_cnt_reg[4]/P0001 ,
		_w6200_
	);
	LUT4 #(
		.INIT('hf531)
	) name4451 (
		\u4_u2_csr0_reg[4]/P0001 ,
		\u4_u2_csr0_reg[5]/P0001 ,
		\u4_u2_dma_in_cnt_reg[2]/P0001 ,
		\u4_u2_dma_in_cnt_reg[3]/P0001 ,
		_w6201_
	);
	LUT4 #(
		.INIT('h0b00)
	) name4452 (
		_w4493_,
		_w4494_,
		_w6200_,
		_w6201_,
		_w6202_
	);
	LUT4 #(
		.INIT('h1040)
	) name4453 (
		\u4_u2_csr0_reg[5]/P0001 ,
		\u4_u2_csr0_reg[6]/P0001 ,
		\u4_u2_dma_in_cnt_reg[3]/P0001 ,
		\u4_u2_dma_in_cnt_reg[4]/P0001 ,
		_w6203_
	);
	LUT2 #(
		.INIT('h2)
	) name4454 (
		_w4610_,
		_w6203_,
		_w6204_
	);
	LUT4 #(
		.INIT('h8c23)
	) name4455 (
		\u4_u2_csr0_reg[5]/P0001 ,
		\u4_u2_csr0_reg[6]/P0001 ,
		\u4_u2_dma_in_cnt_reg[3]/P0001 ,
		\u4_u2_dma_in_cnt_reg[4]/P0001 ,
		_w6205_
	);
	LUT4 #(
		.INIT('h4f00)
	) name4456 (
		_w4493_,
		_w4494_,
		_w6201_,
		_w6205_,
		_w6206_
	);
	LUT4 #(
		.INIT('h0020)
	) name4457 (
		_w6199_,
		_w6202_,
		_w6204_,
		_w6206_,
		_w6207_
	);
	LUT4 #(
		.INIT('h0001)
	) name4458 (
		\u1_u3_buf0_rl_reg/P0001 ,
		\u1_u3_buf0_set_reg/P0001 ,
		\u4_u2_dma_in_cnt_reg[4]/P0001 ,
		\u4_u2_set_r_reg/P0001 ,
		_w6208_
	);
	LUT3 #(
		.INIT('h0e)
	) name4459 (
		\u4_u2_dma_in_cnt_reg[4]/P0001 ,
		\u4_u2_ep_match_r_reg/P0001 ,
		\u4_u2_r5_reg/NET0131 ,
		_w6209_
	);
	LUT2 #(
		.INIT('h4)
	) name4460 (
		_w6208_,
		_w6209_,
		_w6210_
	);
	LUT3 #(
		.INIT('ha2)
	) name4461 (
		\u4_u2_csr1_reg[0]/P0001 ,
		_w6199_,
		_w6210_,
		_w6211_
	);
	LUT2 #(
		.INIT('h4)
	) name4462 (
		_w6207_,
		_w6211_,
		_w6212_
	);
	LUT4 #(
		.INIT('h135f)
	) name4463 (
		\u4_u3_csr0_reg[4]/P0001 ,
		\u4_u3_csr0_reg[5]/P0001 ,
		\u4_u3_dma_out_cnt_reg[2]/P0001 ,
		\u4_u3_dma_out_cnt_reg[3]/P0001 ,
		_w6213_
	);
	LUT2 #(
		.INIT('h6)
	) name4464 (
		\u4_u3_csr0_reg[6]/P0001 ,
		\u4_u3_dma_out_cnt_reg[4]/P0001 ,
		_w6214_
	);
	LUT4 #(
		.INIT('hc832)
	) name4465 (
		\u4_u3_csr0_reg[5]/P0001 ,
		\u4_u3_csr0_reg[6]/P0001 ,
		\u4_u3_dma_out_cnt_reg[3]/P0001 ,
		\u4_u3_dma_out_cnt_reg[4]/P0001 ,
		_w6215_
	);
	LUT4 #(
		.INIT('h4f00)
	) name4466 (
		_w4669_,
		_w4670_,
		_w6213_,
		_w6215_,
		_w6216_
	);
	LUT4 #(
		.INIT('hb000)
	) name4467 (
		_w4669_,
		_w4670_,
		_w6213_,
		_w6214_,
		_w6217_
	);
	LUT3 #(
		.INIT('hb7)
	) name4468 (
		\u4_u3_dma_out_cnt_reg[4]/P0001 ,
		\u4_u3_r5_reg/NET0131 ,
		_w4652_,
		_w6218_
	);
	LUT4 #(
		.INIT('h0104)
	) name4469 (
		\u4_u3_csr0_reg[5]/P0001 ,
		\u4_u3_csr0_reg[6]/P0001 ,
		\u4_u3_dma_out_cnt_reg[3]/P0001 ,
		\u4_u3_dma_out_cnt_reg[4]/P0001 ,
		_w6219_
	);
	LUT4 #(
		.INIT('h00b7)
	) name4470 (
		\u4_u3_dma_out_cnt_reg[4]/P0001 ,
		\u4_u3_r5_reg/NET0131 ,
		_w4652_,
		_w6219_,
		_w6220_
	);
	LUT4 #(
		.INIT('h0200)
	) name4471 (
		_w4569_,
		_w6216_,
		_w6217_,
		_w6220_,
		_w6221_
	);
	LUT4 #(
		.INIT('h0001)
	) name4472 (
		\u1_u3_buf0_rl_reg/P0001 ,
		\u1_u3_buf0_set_reg/P0001 ,
		\u4_u3_dma_out_cnt_reg[4]/P0001 ,
		\u4_u3_set_r_reg/P0001 ,
		_w6222_
	);
	LUT3 #(
		.INIT('h0e)
	) name4473 (
		\u4_u3_dma_out_cnt_reg[4]/P0001 ,
		\u4_u3_ep_match_r_reg/P0001 ,
		\u4_u3_r5_reg/NET0131 ,
		_w6223_
	);
	LUT2 #(
		.INIT('h4)
	) name4474 (
		_w6222_,
		_w6223_,
		_w6224_
	);
	LUT3 #(
		.INIT('ha2)
	) name4475 (
		\u4_u3_csr1_reg[0]/P0001 ,
		_w6218_,
		_w6224_,
		_w6225_
	);
	LUT2 #(
		.INIT('h4)
	) name4476 (
		_w6221_,
		_w6225_,
		_w6226_
	);
	LUT4 #(
		.INIT('h135f)
	) name4477 (
		\u4_u0_csr0_reg[4]/P0001 ,
		\u4_u0_csr0_reg[5]/P0001 ,
		\u4_u0_dma_out_cnt_reg[2]/P0001 ,
		\u4_u0_dma_out_cnt_reg[3]/P0001 ,
		_w6227_
	);
	LUT2 #(
		.INIT('h6)
	) name4478 (
		\u4_u0_csr0_reg[6]/P0001 ,
		\u4_u0_dma_out_cnt_reg[4]/P0001 ,
		_w6228_
	);
	LUT4 #(
		.INIT('hc832)
	) name4479 (
		\u4_u0_csr0_reg[5]/P0001 ,
		\u4_u0_csr0_reg[6]/P0001 ,
		\u4_u0_dma_out_cnt_reg[3]/P0001 ,
		\u4_u0_dma_out_cnt_reg[4]/P0001 ,
		_w6229_
	);
	LUT4 #(
		.INIT('h4f00)
	) name4480 (
		_w4699_,
		_w4700_,
		_w6227_,
		_w6229_,
		_w6230_
	);
	LUT4 #(
		.INIT('hb000)
	) name4481 (
		_w4699_,
		_w4700_,
		_w6227_,
		_w6228_,
		_w6231_
	);
	LUT3 #(
		.INIT('hb7)
	) name4482 (
		\u4_u0_dma_out_cnt_reg[4]/P0001 ,
		\u4_u0_r5_reg/NET0131 ,
		_w4683_,
		_w6232_
	);
	LUT4 #(
		.INIT('h0104)
	) name4483 (
		\u4_u0_csr0_reg[5]/P0001 ,
		\u4_u0_csr0_reg[6]/P0001 ,
		\u4_u0_dma_out_cnt_reg[3]/P0001 ,
		\u4_u0_dma_out_cnt_reg[4]/P0001 ,
		_w6233_
	);
	LUT4 #(
		.INIT('h00b7)
	) name4484 (
		\u4_u0_dma_out_cnt_reg[4]/P0001 ,
		\u4_u0_r5_reg/NET0131 ,
		_w4683_,
		_w6233_,
		_w6234_
	);
	LUT4 #(
		.INIT('h0200)
	) name4485 (
		_w4592_,
		_w6230_,
		_w6231_,
		_w6234_,
		_w6235_
	);
	LUT4 #(
		.INIT('h0001)
	) name4486 (
		\u1_u3_buf0_rl_reg/P0001 ,
		\u1_u3_buf0_set_reg/P0001 ,
		\u4_u0_dma_out_cnt_reg[4]/P0001 ,
		\u4_u0_set_r_reg/P0001 ,
		_w6236_
	);
	LUT3 #(
		.INIT('h0e)
	) name4487 (
		\u4_u0_dma_out_cnt_reg[4]/P0001 ,
		\u4_u0_ep_match_r_reg/P0001 ,
		\u4_u0_r5_reg/NET0131 ,
		_w6237_
	);
	LUT2 #(
		.INIT('h4)
	) name4488 (
		_w6236_,
		_w6237_,
		_w6238_
	);
	LUT3 #(
		.INIT('ha2)
	) name4489 (
		\u4_u0_csr1_reg[0]/P0001 ,
		_w6232_,
		_w6238_,
		_w6239_
	);
	LUT2 #(
		.INIT('h4)
	) name4490 (
		_w6235_,
		_w6239_,
		_w6240_
	);
	LUT4 #(
		.INIT('h135f)
	) name4491 (
		\u4_u1_csr0_reg[4]/P0001 ,
		\u4_u1_csr0_reg[5]/P0001 ,
		\u4_u1_dma_out_cnt_reg[2]/P0001 ,
		\u4_u1_dma_out_cnt_reg[3]/P0001 ,
		_w6241_
	);
	LUT2 #(
		.INIT('h6)
	) name4492 (
		\u4_u1_csr0_reg[6]/P0001 ,
		\u4_u1_dma_out_cnt_reg[4]/P0001 ,
		_w6242_
	);
	LUT4 #(
		.INIT('hc832)
	) name4493 (
		\u4_u1_csr0_reg[5]/P0001 ,
		\u4_u1_csr0_reg[6]/P0001 ,
		\u4_u1_dma_out_cnt_reg[3]/P0001 ,
		\u4_u1_dma_out_cnt_reg[4]/P0001 ,
		_w6243_
	);
	LUT4 #(
		.INIT('h4f00)
	) name4494 (
		_w4730_,
		_w4731_,
		_w6241_,
		_w6243_,
		_w6244_
	);
	LUT4 #(
		.INIT('hb000)
	) name4495 (
		_w4730_,
		_w4731_,
		_w6241_,
		_w6242_,
		_w6245_
	);
	LUT3 #(
		.INIT('hb7)
	) name4496 (
		\u4_u1_dma_out_cnt_reg[4]/P0001 ,
		\u4_u1_r5_reg/NET0131 ,
		_w4713_,
		_w6246_
	);
	LUT4 #(
		.INIT('h0104)
	) name4497 (
		\u4_u1_csr0_reg[5]/P0001 ,
		\u4_u1_csr0_reg[6]/P0001 ,
		\u4_u1_dma_out_cnt_reg[3]/P0001 ,
		\u4_u1_dma_out_cnt_reg[4]/P0001 ,
		_w6247_
	);
	LUT4 #(
		.INIT('h00b7)
	) name4498 (
		\u4_u1_dma_out_cnt_reg[4]/P0001 ,
		\u4_u1_r5_reg/NET0131 ,
		_w4713_,
		_w6247_,
		_w6248_
	);
	LUT4 #(
		.INIT('h0200)
	) name4499 (
		_w4454_,
		_w6244_,
		_w6245_,
		_w6248_,
		_w6249_
	);
	LUT4 #(
		.INIT('h0001)
	) name4500 (
		\u1_u3_buf0_rl_reg/P0001 ,
		\u1_u3_buf0_set_reg/P0001 ,
		\u4_u1_dma_out_cnt_reg[4]/P0001 ,
		\u4_u1_set_r_reg/P0001 ,
		_w6250_
	);
	LUT3 #(
		.INIT('h0e)
	) name4501 (
		\u4_u1_dma_out_cnt_reg[4]/P0001 ,
		\u4_u1_ep_match_r_reg/P0001 ,
		\u4_u1_r5_reg/NET0131 ,
		_w6251_
	);
	LUT2 #(
		.INIT('h4)
	) name4502 (
		_w6250_,
		_w6251_,
		_w6252_
	);
	LUT3 #(
		.INIT('ha2)
	) name4503 (
		\u4_u1_csr1_reg[0]/P0001 ,
		_w6246_,
		_w6252_,
		_w6253_
	);
	LUT2 #(
		.INIT('h4)
	) name4504 (
		_w6249_,
		_w6253_,
		_w6254_
	);
	LUT4 #(
		.INIT('h135f)
	) name4505 (
		\u4_u2_csr0_reg[4]/P0001 ,
		\u4_u2_csr0_reg[5]/P0001 ,
		\u4_u2_dma_out_cnt_reg[2]/P0001 ,
		\u4_u2_dma_out_cnt_reg[3]/P0001 ,
		_w6255_
	);
	LUT2 #(
		.INIT('h6)
	) name4506 (
		\u4_u2_csr0_reg[6]/P0001 ,
		\u4_u2_dma_out_cnt_reg[4]/P0001 ,
		_w6256_
	);
	LUT4 #(
		.INIT('hc832)
	) name4507 (
		\u4_u2_csr0_reg[5]/P0001 ,
		\u4_u2_csr0_reg[6]/P0001 ,
		\u4_u2_dma_out_cnt_reg[3]/P0001 ,
		\u4_u2_dma_out_cnt_reg[4]/P0001 ,
		_w6257_
	);
	LUT4 #(
		.INIT('h4f00)
	) name4508 (
		_w4760_,
		_w4761_,
		_w6255_,
		_w6257_,
		_w6258_
	);
	LUT4 #(
		.INIT('hb000)
	) name4509 (
		_w4760_,
		_w4761_,
		_w6255_,
		_w6256_,
		_w6259_
	);
	LUT3 #(
		.INIT('hb7)
	) name4510 (
		\u4_u2_dma_out_cnt_reg[4]/P0001 ,
		\u4_u2_r5_reg/NET0131 ,
		_w4744_,
		_w6260_
	);
	LUT4 #(
		.INIT('h0104)
	) name4511 (
		\u4_u2_csr0_reg[5]/P0001 ,
		\u4_u2_csr0_reg[6]/P0001 ,
		\u4_u2_dma_out_cnt_reg[3]/P0001 ,
		\u4_u2_dma_out_cnt_reg[4]/P0001 ,
		_w6261_
	);
	LUT4 #(
		.INIT('h00b7)
	) name4512 (
		\u4_u2_dma_out_cnt_reg[4]/P0001 ,
		\u4_u2_r5_reg/NET0131 ,
		_w4744_,
		_w6261_,
		_w6262_
	);
	LUT4 #(
		.INIT('h0200)
	) name4513 (
		_w4610_,
		_w6258_,
		_w6259_,
		_w6262_,
		_w6263_
	);
	LUT4 #(
		.INIT('h0001)
	) name4514 (
		\u1_u3_buf0_rl_reg/P0001 ,
		\u1_u3_buf0_set_reg/P0001 ,
		\u4_u2_dma_out_cnt_reg[4]/P0001 ,
		\u4_u2_set_r_reg/P0001 ,
		_w6264_
	);
	LUT3 #(
		.INIT('h0e)
	) name4515 (
		\u4_u2_dma_out_cnt_reg[4]/P0001 ,
		\u4_u2_ep_match_r_reg/P0001 ,
		\u4_u2_r5_reg/NET0131 ,
		_w6265_
	);
	LUT2 #(
		.INIT('h4)
	) name4516 (
		_w6264_,
		_w6265_,
		_w6266_
	);
	LUT3 #(
		.INIT('ha2)
	) name4517 (
		\u4_u2_csr1_reg[0]/P0001 ,
		_w6260_,
		_w6266_,
		_w6267_
	);
	LUT2 #(
		.INIT('h4)
	) name4518 (
		_w6263_,
		_w6267_,
		_w6268_
	);
	LUT4 #(
		.INIT('h10f0)
	) name4519 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u3_buf1_reg[0]/P0001 ,
		\u4_u3_ep_match_r_reg/P0001 ,
		_w6269_
	);
	LUT4 #(
		.INIT('hc800)
	) name4520 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_idin_reg[0]/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u3_ep_match_r_reg/P0001 ,
		_w6270_
	);
	LUT2 #(
		.INIT('h1)
	) name4521 (
		_w6269_,
		_w6270_,
		_w6271_
	);
	LUT3 #(
		.INIT('h07)
	) name4522 (
		_w2231_,
		_w2320_,
		_w6271_,
		_w6272_
	);
	LUT3 #(
		.INIT('h80)
	) name4523 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_data_i[0]_pad ,
		_w6273_
	);
	LUT3 #(
		.INIT('h2a)
	) name4524 (
		rst_i_pad,
		_w2231_,
		_w6273_,
		_w6274_
	);
	LUT2 #(
		.INIT('hb)
	) name4525 (
		_w6272_,
		_w6274_,
		_w6275_
	);
	LUT4 #(
		.INIT('h10f0)
	) name4526 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u3_buf1_reg[12]/P0001 ,
		\u4_u3_ep_match_r_reg/P0001 ,
		_w6276_
	);
	LUT4 #(
		.INIT('hc800)
	) name4527 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_idin_reg[12]/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u3_ep_match_r_reg/P0001 ,
		_w6277_
	);
	LUT2 #(
		.INIT('h1)
	) name4528 (
		_w6276_,
		_w6277_,
		_w6278_
	);
	LUT3 #(
		.INIT('h07)
	) name4529 (
		_w2231_,
		_w2320_,
		_w6278_,
		_w6279_
	);
	LUT3 #(
		.INIT('h80)
	) name4530 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_data_i[12]_pad ,
		_w6280_
	);
	LUT3 #(
		.INIT('h2a)
	) name4531 (
		rst_i_pad,
		_w2231_,
		_w6280_,
		_w6281_
	);
	LUT2 #(
		.INIT('hb)
	) name4532 (
		_w6279_,
		_w6281_,
		_w6282_
	);
	LUT4 #(
		.INIT('h10f0)
	) name4533 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u3_buf1_reg[16]/P0001 ,
		\u4_u3_ep_match_r_reg/P0001 ,
		_w6283_
	);
	LUT4 #(
		.INIT('hc800)
	) name4534 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_idin_reg[16]/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u3_ep_match_r_reg/P0001 ,
		_w6284_
	);
	LUT2 #(
		.INIT('h1)
	) name4535 (
		_w6283_,
		_w6284_,
		_w6285_
	);
	LUT3 #(
		.INIT('h07)
	) name4536 (
		_w2231_,
		_w2320_,
		_w6285_,
		_w6286_
	);
	LUT3 #(
		.INIT('h80)
	) name4537 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_data_i[16]_pad ,
		_w6287_
	);
	LUT3 #(
		.INIT('h2a)
	) name4538 (
		rst_i_pad,
		_w2231_,
		_w6287_,
		_w6288_
	);
	LUT2 #(
		.INIT('hb)
	) name4539 (
		_w6286_,
		_w6288_,
		_w6289_
	);
	LUT4 #(
		.INIT('h10f0)
	) name4540 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u3_buf1_reg[17]/P0001 ,
		\u4_u3_ep_match_r_reg/P0001 ,
		_w6290_
	);
	LUT4 #(
		.INIT('hc800)
	) name4541 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_idin_reg[17]/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u3_ep_match_r_reg/P0001 ,
		_w6291_
	);
	LUT2 #(
		.INIT('h1)
	) name4542 (
		_w6290_,
		_w6291_,
		_w6292_
	);
	LUT3 #(
		.INIT('h07)
	) name4543 (
		_w2231_,
		_w2320_,
		_w6292_,
		_w6293_
	);
	LUT3 #(
		.INIT('h80)
	) name4544 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_data_i[17]_pad ,
		_w6294_
	);
	LUT3 #(
		.INIT('h2a)
	) name4545 (
		rst_i_pad,
		_w2231_,
		_w6294_,
		_w6295_
	);
	LUT2 #(
		.INIT('hb)
	) name4546 (
		_w6293_,
		_w6295_,
		_w6296_
	);
	LUT4 #(
		.INIT('h10f0)
	) name4547 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u3_buf1_reg[18]/P0001 ,
		\u4_u3_ep_match_r_reg/P0001 ,
		_w6297_
	);
	LUT4 #(
		.INIT('hc800)
	) name4548 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_idin_reg[18]/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u3_ep_match_r_reg/P0001 ,
		_w6298_
	);
	LUT2 #(
		.INIT('h1)
	) name4549 (
		_w6297_,
		_w6298_,
		_w6299_
	);
	LUT3 #(
		.INIT('h07)
	) name4550 (
		_w2231_,
		_w2320_,
		_w6299_,
		_w6300_
	);
	LUT3 #(
		.INIT('h80)
	) name4551 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_data_i[18]_pad ,
		_w6301_
	);
	LUT3 #(
		.INIT('h2a)
	) name4552 (
		rst_i_pad,
		_w2231_,
		_w6301_,
		_w6302_
	);
	LUT2 #(
		.INIT('hb)
	) name4553 (
		_w6300_,
		_w6302_,
		_w6303_
	);
	LUT4 #(
		.INIT('h10f0)
	) name4554 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u3_buf1_reg[19]/P0001 ,
		\u4_u3_ep_match_r_reg/P0001 ,
		_w6304_
	);
	LUT4 #(
		.INIT('hc800)
	) name4555 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_idin_reg[19]/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u3_ep_match_r_reg/P0001 ,
		_w6305_
	);
	LUT2 #(
		.INIT('h1)
	) name4556 (
		_w6304_,
		_w6305_,
		_w6306_
	);
	LUT3 #(
		.INIT('h07)
	) name4557 (
		_w2231_,
		_w2320_,
		_w6306_,
		_w6307_
	);
	LUT3 #(
		.INIT('h80)
	) name4558 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_data_i[19]_pad ,
		_w6308_
	);
	LUT3 #(
		.INIT('h2a)
	) name4559 (
		rst_i_pad,
		_w2231_,
		_w6308_,
		_w6309_
	);
	LUT2 #(
		.INIT('hb)
	) name4560 (
		_w6307_,
		_w6309_,
		_w6310_
	);
	LUT4 #(
		.INIT('h10f0)
	) name4561 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u3_buf1_reg[1]/P0001 ,
		\u4_u3_ep_match_r_reg/P0001 ,
		_w6311_
	);
	LUT4 #(
		.INIT('hc800)
	) name4562 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_idin_reg[1]/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u3_ep_match_r_reg/P0001 ,
		_w6312_
	);
	LUT2 #(
		.INIT('h1)
	) name4563 (
		_w6311_,
		_w6312_,
		_w6313_
	);
	LUT3 #(
		.INIT('h07)
	) name4564 (
		_w2231_,
		_w2320_,
		_w6313_,
		_w6314_
	);
	LUT3 #(
		.INIT('h80)
	) name4565 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_data_i[1]_pad ,
		_w6315_
	);
	LUT3 #(
		.INIT('h2a)
	) name4566 (
		rst_i_pad,
		_w2231_,
		_w6315_,
		_w6316_
	);
	LUT2 #(
		.INIT('hb)
	) name4567 (
		_w6314_,
		_w6316_,
		_w6317_
	);
	LUT4 #(
		.INIT('h10f0)
	) name4568 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u3_buf1_reg[20]/P0001 ,
		\u4_u3_ep_match_r_reg/P0001 ,
		_w6318_
	);
	LUT4 #(
		.INIT('hc800)
	) name4569 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_idin_reg[20]/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u3_ep_match_r_reg/P0001 ,
		_w6319_
	);
	LUT2 #(
		.INIT('h1)
	) name4570 (
		_w6318_,
		_w6319_,
		_w6320_
	);
	LUT3 #(
		.INIT('h07)
	) name4571 (
		_w2231_,
		_w2320_,
		_w6320_,
		_w6321_
	);
	LUT3 #(
		.INIT('h80)
	) name4572 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_data_i[20]_pad ,
		_w6322_
	);
	LUT3 #(
		.INIT('h2a)
	) name4573 (
		rst_i_pad,
		_w2231_,
		_w6322_,
		_w6323_
	);
	LUT2 #(
		.INIT('hb)
	) name4574 (
		_w6321_,
		_w6323_,
		_w6324_
	);
	LUT4 #(
		.INIT('h10f0)
	) name4575 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u3_buf1_reg[21]/P0001 ,
		\u4_u3_ep_match_r_reg/P0001 ,
		_w6325_
	);
	LUT4 #(
		.INIT('hc800)
	) name4576 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_idin_reg[21]/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u3_ep_match_r_reg/P0001 ,
		_w6326_
	);
	LUT2 #(
		.INIT('h1)
	) name4577 (
		_w6325_,
		_w6326_,
		_w6327_
	);
	LUT3 #(
		.INIT('h07)
	) name4578 (
		_w2231_,
		_w2320_,
		_w6327_,
		_w6328_
	);
	LUT3 #(
		.INIT('h80)
	) name4579 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_data_i[21]_pad ,
		_w6329_
	);
	LUT3 #(
		.INIT('h2a)
	) name4580 (
		rst_i_pad,
		_w2231_,
		_w6329_,
		_w6330_
	);
	LUT2 #(
		.INIT('hb)
	) name4581 (
		_w6328_,
		_w6330_,
		_w6331_
	);
	LUT4 #(
		.INIT('h10f0)
	) name4582 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u3_buf1_reg[22]/P0001 ,
		\u4_u3_ep_match_r_reg/P0001 ,
		_w6332_
	);
	LUT4 #(
		.INIT('hc800)
	) name4583 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_idin_reg[22]/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u3_ep_match_r_reg/P0001 ,
		_w6333_
	);
	LUT2 #(
		.INIT('h1)
	) name4584 (
		_w6332_,
		_w6333_,
		_w6334_
	);
	LUT3 #(
		.INIT('h07)
	) name4585 (
		_w2231_,
		_w2320_,
		_w6334_,
		_w6335_
	);
	LUT3 #(
		.INIT('h80)
	) name4586 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_data_i[22]_pad ,
		_w6336_
	);
	LUT3 #(
		.INIT('h2a)
	) name4587 (
		rst_i_pad,
		_w2231_,
		_w6336_,
		_w6337_
	);
	LUT2 #(
		.INIT('hb)
	) name4588 (
		_w6335_,
		_w6337_,
		_w6338_
	);
	LUT4 #(
		.INIT('h10f0)
	) name4589 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u3_buf1_reg[23]/P0001 ,
		\u4_u3_ep_match_r_reg/P0001 ,
		_w6339_
	);
	LUT4 #(
		.INIT('hc800)
	) name4590 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_idin_reg[23]/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u3_ep_match_r_reg/P0001 ,
		_w6340_
	);
	LUT2 #(
		.INIT('h1)
	) name4591 (
		_w6339_,
		_w6340_,
		_w6341_
	);
	LUT3 #(
		.INIT('h07)
	) name4592 (
		_w2231_,
		_w2320_,
		_w6341_,
		_w6342_
	);
	LUT3 #(
		.INIT('h80)
	) name4593 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_data_i[23]_pad ,
		_w6343_
	);
	LUT3 #(
		.INIT('h2a)
	) name4594 (
		rst_i_pad,
		_w2231_,
		_w6343_,
		_w6344_
	);
	LUT2 #(
		.INIT('hb)
	) name4595 (
		_w6342_,
		_w6344_,
		_w6345_
	);
	LUT4 #(
		.INIT('h10f0)
	) name4596 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u3_buf1_reg[24]/P0001 ,
		\u4_u3_ep_match_r_reg/P0001 ,
		_w6346_
	);
	LUT4 #(
		.INIT('hc800)
	) name4597 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_idin_reg[24]/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u3_ep_match_r_reg/P0001 ,
		_w6347_
	);
	LUT2 #(
		.INIT('h1)
	) name4598 (
		_w6346_,
		_w6347_,
		_w6348_
	);
	LUT3 #(
		.INIT('h07)
	) name4599 (
		_w2231_,
		_w2320_,
		_w6348_,
		_w6349_
	);
	LUT3 #(
		.INIT('h80)
	) name4600 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_data_i[24]_pad ,
		_w6350_
	);
	LUT3 #(
		.INIT('h2a)
	) name4601 (
		rst_i_pad,
		_w2231_,
		_w6350_,
		_w6351_
	);
	LUT2 #(
		.INIT('hb)
	) name4602 (
		_w6349_,
		_w6351_,
		_w6352_
	);
	LUT4 #(
		.INIT('h10f0)
	) name4603 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u3_buf1_reg[25]/P0001 ,
		\u4_u3_ep_match_r_reg/P0001 ,
		_w6353_
	);
	LUT4 #(
		.INIT('hc800)
	) name4604 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_idin_reg[25]/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u3_ep_match_r_reg/P0001 ,
		_w6354_
	);
	LUT2 #(
		.INIT('h1)
	) name4605 (
		_w6353_,
		_w6354_,
		_w6355_
	);
	LUT3 #(
		.INIT('h07)
	) name4606 (
		_w2231_,
		_w2320_,
		_w6355_,
		_w6356_
	);
	LUT3 #(
		.INIT('h80)
	) name4607 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_data_i[25]_pad ,
		_w6357_
	);
	LUT3 #(
		.INIT('h2a)
	) name4608 (
		rst_i_pad,
		_w2231_,
		_w6357_,
		_w6358_
	);
	LUT2 #(
		.INIT('hb)
	) name4609 (
		_w6356_,
		_w6358_,
		_w6359_
	);
	LUT4 #(
		.INIT('h10f0)
	) name4610 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u3_buf1_reg[26]/P0001 ,
		\u4_u3_ep_match_r_reg/P0001 ,
		_w6360_
	);
	LUT4 #(
		.INIT('hc800)
	) name4611 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_idin_reg[26]/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u3_ep_match_r_reg/P0001 ,
		_w6361_
	);
	LUT2 #(
		.INIT('h1)
	) name4612 (
		_w6360_,
		_w6361_,
		_w6362_
	);
	LUT3 #(
		.INIT('h07)
	) name4613 (
		_w2231_,
		_w2320_,
		_w6362_,
		_w6363_
	);
	LUT3 #(
		.INIT('h80)
	) name4614 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_data_i[26]_pad ,
		_w6364_
	);
	LUT3 #(
		.INIT('h2a)
	) name4615 (
		rst_i_pad,
		_w2231_,
		_w6364_,
		_w6365_
	);
	LUT2 #(
		.INIT('hb)
	) name4616 (
		_w6363_,
		_w6365_,
		_w6366_
	);
	LUT4 #(
		.INIT('h10f0)
	) name4617 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u3_buf1_reg[27]/P0001 ,
		\u4_u3_ep_match_r_reg/P0001 ,
		_w6367_
	);
	LUT4 #(
		.INIT('hc800)
	) name4618 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_idin_reg[27]/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u3_ep_match_r_reg/P0001 ,
		_w6368_
	);
	LUT2 #(
		.INIT('h1)
	) name4619 (
		_w6367_,
		_w6368_,
		_w6369_
	);
	LUT3 #(
		.INIT('h07)
	) name4620 (
		_w2231_,
		_w2320_,
		_w6369_,
		_w6370_
	);
	LUT3 #(
		.INIT('h80)
	) name4621 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_data_i[27]_pad ,
		_w6371_
	);
	LUT3 #(
		.INIT('h2a)
	) name4622 (
		rst_i_pad,
		_w2231_,
		_w6371_,
		_w6372_
	);
	LUT2 #(
		.INIT('hb)
	) name4623 (
		_w6370_,
		_w6372_,
		_w6373_
	);
	LUT4 #(
		.INIT('h10f0)
	) name4624 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u3_buf1_reg[28]/P0001 ,
		\u4_u3_ep_match_r_reg/P0001 ,
		_w6374_
	);
	LUT4 #(
		.INIT('hc800)
	) name4625 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_idin_reg[28]/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u3_ep_match_r_reg/P0001 ,
		_w6375_
	);
	LUT2 #(
		.INIT('h1)
	) name4626 (
		_w6374_,
		_w6375_,
		_w6376_
	);
	LUT3 #(
		.INIT('h07)
	) name4627 (
		_w2231_,
		_w2320_,
		_w6376_,
		_w6377_
	);
	LUT3 #(
		.INIT('h80)
	) name4628 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_data_i[28]_pad ,
		_w6378_
	);
	LUT3 #(
		.INIT('h2a)
	) name4629 (
		rst_i_pad,
		_w2231_,
		_w6378_,
		_w6379_
	);
	LUT2 #(
		.INIT('hb)
	) name4630 (
		_w6377_,
		_w6379_,
		_w6380_
	);
	LUT4 #(
		.INIT('h10f0)
	) name4631 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u3_buf1_reg[29]/P0001 ,
		\u4_u3_ep_match_r_reg/P0001 ,
		_w6381_
	);
	LUT4 #(
		.INIT('hc800)
	) name4632 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_idin_reg[29]/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u3_ep_match_r_reg/P0001 ,
		_w6382_
	);
	LUT2 #(
		.INIT('h1)
	) name4633 (
		_w6381_,
		_w6382_,
		_w6383_
	);
	LUT3 #(
		.INIT('h07)
	) name4634 (
		_w2231_,
		_w2320_,
		_w6383_,
		_w6384_
	);
	LUT3 #(
		.INIT('h80)
	) name4635 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_data_i[29]_pad ,
		_w6385_
	);
	LUT3 #(
		.INIT('h2a)
	) name4636 (
		rst_i_pad,
		_w2231_,
		_w6385_,
		_w6386_
	);
	LUT2 #(
		.INIT('hb)
	) name4637 (
		_w6384_,
		_w6386_,
		_w6387_
	);
	LUT4 #(
		.INIT('h10f0)
	) name4638 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u3_buf1_reg[2]/P0001 ,
		\u4_u3_ep_match_r_reg/P0001 ,
		_w6388_
	);
	LUT4 #(
		.INIT('hc800)
	) name4639 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_idin_reg[2]/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u3_ep_match_r_reg/P0001 ,
		_w6389_
	);
	LUT2 #(
		.INIT('h1)
	) name4640 (
		_w6388_,
		_w6389_,
		_w6390_
	);
	LUT3 #(
		.INIT('h07)
	) name4641 (
		_w2231_,
		_w2320_,
		_w6390_,
		_w6391_
	);
	LUT3 #(
		.INIT('h80)
	) name4642 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_data_i[2]_pad ,
		_w6392_
	);
	LUT3 #(
		.INIT('h2a)
	) name4643 (
		rst_i_pad,
		_w2231_,
		_w6392_,
		_w6393_
	);
	LUT2 #(
		.INIT('hb)
	) name4644 (
		_w6391_,
		_w6393_,
		_w6394_
	);
	LUT4 #(
		.INIT('h10f0)
	) name4645 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u3_buf1_reg[30]/P0001 ,
		\u4_u3_ep_match_r_reg/P0001 ,
		_w6395_
	);
	LUT4 #(
		.INIT('hc800)
	) name4646 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_idin_reg[30]/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u3_ep_match_r_reg/P0001 ,
		_w6396_
	);
	LUT2 #(
		.INIT('h1)
	) name4647 (
		_w6395_,
		_w6396_,
		_w6397_
	);
	LUT3 #(
		.INIT('h07)
	) name4648 (
		_w2231_,
		_w2320_,
		_w6397_,
		_w6398_
	);
	LUT3 #(
		.INIT('h80)
	) name4649 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_data_i[30]_pad ,
		_w6399_
	);
	LUT3 #(
		.INIT('h2a)
	) name4650 (
		rst_i_pad,
		_w2231_,
		_w6399_,
		_w6400_
	);
	LUT2 #(
		.INIT('hb)
	) name4651 (
		_w6398_,
		_w6400_,
		_w6401_
	);
	LUT4 #(
		.INIT('h10f0)
	) name4652 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u3_buf1_reg[31]/P0001 ,
		\u4_u3_ep_match_r_reg/P0001 ,
		_w6402_
	);
	LUT4 #(
		.INIT('hc800)
	) name4653 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_idin_reg[31]/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u3_ep_match_r_reg/P0001 ,
		_w6403_
	);
	LUT2 #(
		.INIT('h1)
	) name4654 (
		_w6402_,
		_w6403_,
		_w6404_
	);
	LUT3 #(
		.INIT('h07)
	) name4655 (
		_w2231_,
		_w2320_,
		_w6404_,
		_w6405_
	);
	LUT3 #(
		.INIT('h80)
	) name4656 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_data_i[31]_pad ,
		_w6406_
	);
	LUT3 #(
		.INIT('h2a)
	) name4657 (
		rst_i_pad,
		_w2231_,
		_w6406_,
		_w6407_
	);
	LUT2 #(
		.INIT('hb)
	) name4658 (
		_w6405_,
		_w6407_,
		_w6408_
	);
	LUT4 #(
		.INIT('h10f0)
	) name4659 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u3_buf1_reg[3]/P0001 ,
		\u4_u3_ep_match_r_reg/P0001 ,
		_w6409_
	);
	LUT4 #(
		.INIT('hc800)
	) name4660 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_idin_reg[3]/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u3_ep_match_r_reg/P0001 ,
		_w6410_
	);
	LUT2 #(
		.INIT('h1)
	) name4661 (
		_w6409_,
		_w6410_,
		_w6411_
	);
	LUT3 #(
		.INIT('h07)
	) name4662 (
		_w2231_,
		_w2320_,
		_w6411_,
		_w6412_
	);
	LUT3 #(
		.INIT('h80)
	) name4663 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_data_i[3]_pad ,
		_w6413_
	);
	LUT3 #(
		.INIT('h2a)
	) name4664 (
		rst_i_pad,
		_w2231_,
		_w6413_,
		_w6414_
	);
	LUT2 #(
		.INIT('hb)
	) name4665 (
		_w6412_,
		_w6414_,
		_w6415_
	);
	LUT4 #(
		.INIT('h10f0)
	) name4666 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u3_buf1_reg[8]/P0001 ,
		\u4_u3_ep_match_r_reg/P0001 ,
		_w6416_
	);
	LUT4 #(
		.INIT('hc800)
	) name4667 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_idin_reg[8]/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u3_ep_match_r_reg/P0001 ,
		_w6417_
	);
	LUT2 #(
		.INIT('h1)
	) name4668 (
		_w6416_,
		_w6417_,
		_w6418_
	);
	LUT3 #(
		.INIT('h07)
	) name4669 (
		_w2231_,
		_w2320_,
		_w6418_,
		_w6419_
	);
	LUT3 #(
		.INIT('h80)
	) name4670 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_data_i[8]_pad ,
		_w6420_
	);
	LUT3 #(
		.INIT('h2a)
	) name4671 (
		rst_i_pad,
		_w2231_,
		_w6420_,
		_w6421_
	);
	LUT2 #(
		.INIT('hb)
	) name4672 (
		_w6419_,
		_w6421_,
		_w6422_
	);
	LUT4 #(
		.INIT('h10f0)
	) name4673 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u3_buf1_reg[9]/P0001 ,
		\u4_u3_ep_match_r_reg/P0001 ,
		_w6423_
	);
	LUT4 #(
		.INIT('hc800)
	) name4674 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_idin_reg[9]/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u3_ep_match_r_reg/P0001 ,
		_w6424_
	);
	LUT2 #(
		.INIT('h1)
	) name4675 (
		_w6423_,
		_w6424_,
		_w6425_
	);
	LUT3 #(
		.INIT('h07)
	) name4676 (
		_w2231_,
		_w2320_,
		_w6425_,
		_w6426_
	);
	LUT3 #(
		.INIT('h80)
	) name4677 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_data_i[9]_pad ,
		_w6427_
	);
	LUT3 #(
		.INIT('h2a)
	) name4678 (
		rst_i_pad,
		_w2231_,
		_w6427_,
		_w6428_
	);
	LUT2 #(
		.INIT('hb)
	) name4679 (
		_w6426_,
		_w6428_,
		_w6429_
	);
	LUT3 #(
		.INIT('h80)
	) name4680 (
		\u5_wb_req_s1_reg/P0001 ,
		\wb_addr_i[17]_pad ,
		wb_we_i_pad,
		_w6430_
	);
	LUT4 #(
		.INIT('h1555)
	) name4681 (
		\u5_state_reg[1]/P0001 ,
		\u5_wb_req_s1_reg/P0001 ,
		\wb_addr_i[17]_pad ,
		wb_we_i_pad,
		_w6431_
	);
	LUT4 #(
		.INIT('h0080)
	) name4682 (
		rst_i_pad,
		_w2224_,
		_w5490_,
		_w6431_,
		_w6432_
	);
	LUT3 #(
		.INIT('hb0)
	) name4683 (
		\u1_u2_word_done_r_reg/P0001 ,
		\u2_wack_r_reg/P0001 ,
		\u5_state_reg[1]/P0001 ,
		_w6433_
	);
	LUT2 #(
		.INIT('h4)
	) name4684 (
		\u1_u2_mack_r_reg/P0001 ,
		\u5_state_reg[1]/P0001 ,
		_w6434_
	);
	LUT4 #(
		.INIT('h020f)
	) name4685 (
		_w3224_,
		_w5488_,
		_w6433_,
		_w6434_,
		_w6435_
	);
	LUT3 #(
		.INIT('h20)
	) name4686 (
		rst_i_pad,
		\u5_state_reg[2]/P0001 ,
		_w5493_,
		_w6436_
	);
	LUT3 #(
		.INIT('hba)
	) name4687 (
		_w6432_,
		_w6435_,
		_w6436_,
		_w6437_
	);
	LUT4 #(
		.INIT('hff80)
	) name4688 (
		\u1_u2_adr_cb_reg[0]/NET0131 ,
		\u1_u2_adr_cb_reg[1]/NET0131 ,
		\u1_u2_rx_data_valid_r_reg/NET0131 ,
		\u1_u2_wr_last_reg/P0001 ,
		_w6438_
	);
	LUT2 #(
		.INIT('h2)
	) name4689 (
		\u1_u2_rx_data_done_r2_reg/P0001 ,
		\u1_u3_abort_reg/P0001 ,
		_w6439_
	);
	LUT4 #(
		.INIT('h3038)
	) name4690 (
		\u1_u2_rx_data_done_r2_reg/P0001 ,
		\u1_u2_state_reg[2]/NET0131 ,
		\u1_u2_state_reg[3]/NET0131 ,
		\u1_u3_abort_reg/P0001 ,
		_w6440_
	);
	LUT3 #(
		.INIT('h0e)
	) name4691 (
		\u1_u2_adr_cb_reg[0]/NET0131 ,
		\u1_u2_adr_cb_reg[1]/NET0131 ,
		\u1_u2_rx_data_valid_r_reg/NET0131 ,
		_w6441_
	);
	LUT4 #(
		.INIT('h8000)
	) name4692 (
		_w3204_,
		_w3209_,
		_w6440_,
		_w6441_,
		_w6442_
	);
	LUT4 #(
		.INIT('h10f0)
	) name4693 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u0_buf1_reg[0]/P0001 ,
		\u4_u0_ep_match_r_reg/P0001 ,
		_w6443_
	);
	LUT4 #(
		.INIT('hc800)
	) name4694 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_idin_reg[0]/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u0_ep_match_r_reg/P0001 ,
		_w6444_
	);
	LUT2 #(
		.INIT('h1)
	) name4695 (
		_w6443_,
		_w6444_,
		_w6445_
	);
	LUT3 #(
		.INIT('h07)
	) name4696 (
		_w2243_,
		_w2320_,
		_w6445_,
		_w6446_
	);
	LUT3 #(
		.INIT('h2a)
	) name4697 (
		rst_i_pad,
		_w2243_,
		_w6273_,
		_w6447_
	);
	LUT2 #(
		.INIT('hb)
	) name4698 (
		_w6446_,
		_w6447_,
		_w6448_
	);
	LUT4 #(
		.INIT('h10f0)
	) name4699 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u0_buf1_reg[12]/P0001 ,
		\u4_u0_ep_match_r_reg/P0001 ,
		_w6449_
	);
	LUT4 #(
		.INIT('hc800)
	) name4700 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_idin_reg[12]/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u0_ep_match_r_reg/P0001 ,
		_w6450_
	);
	LUT2 #(
		.INIT('h1)
	) name4701 (
		_w6449_,
		_w6450_,
		_w6451_
	);
	LUT3 #(
		.INIT('h07)
	) name4702 (
		_w2243_,
		_w2320_,
		_w6451_,
		_w6452_
	);
	LUT3 #(
		.INIT('h2a)
	) name4703 (
		rst_i_pad,
		_w2243_,
		_w6280_,
		_w6453_
	);
	LUT2 #(
		.INIT('hb)
	) name4704 (
		_w6452_,
		_w6453_,
		_w6454_
	);
	LUT4 #(
		.INIT('h10f0)
	) name4705 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u0_buf1_reg[16]/P0001 ,
		\u4_u0_ep_match_r_reg/P0001 ,
		_w6455_
	);
	LUT4 #(
		.INIT('hc800)
	) name4706 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_idin_reg[16]/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u0_ep_match_r_reg/P0001 ,
		_w6456_
	);
	LUT2 #(
		.INIT('h1)
	) name4707 (
		_w6455_,
		_w6456_,
		_w6457_
	);
	LUT3 #(
		.INIT('h07)
	) name4708 (
		_w2243_,
		_w2320_,
		_w6457_,
		_w6458_
	);
	LUT3 #(
		.INIT('h2a)
	) name4709 (
		rst_i_pad,
		_w2243_,
		_w6287_,
		_w6459_
	);
	LUT2 #(
		.INIT('hb)
	) name4710 (
		_w6458_,
		_w6459_,
		_w6460_
	);
	LUT4 #(
		.INIT('h10f0)
	) name4711 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u0_buf1_reg[17]/P0001 ,
		\u4_u0_ep_match_r_reg/P0001 ,
		_w6461_
	);
	LUT4 #(
		.INIT('hc800)
	) name4712 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_idin_reg[17]/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u0_ep_match_r_reg/P0001 ,
		_w6462_
	);
	LUT2 #(
		.INIT('h1)
	) name4713 (
		_w6461_,
		_w6462_,
		_w6463_
	);
	LUT3 #(
		.INIT('h07)
	) name4714 (
		_w2243_,
		_w2320_,
		_w6463_,
		_w6464_
	);
	LUT3 #(
		.INIT('h2a)
	) name4715 (
		rst_i_pad,
		_w2243_,
		_w6294_,
		_w6465_
	);
	LUT2 #(
		.INIT('hb)
	) name4716 (
		_w6464_,
		_w6465_,
		_w6466_
	);
	LUT4 #(
		.INIT('h10f0)
	) name4717 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u0_buf1_reg[18]/P0001 ,
		\u4_u0_ep_match_r_reg/P0001 ,
		_w6467_
	);
	LUT4 #(
		.INIT('hc800)
	) name4718 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_idin_reg[18]/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u0_ep_match_r_reg/P0001 ,
		_w6468_
	);
	LUT2 #(
		.INIT('h1)
	) name4719 (
		_w6467_,
		_w6468_,
		_w6469_
	);
	LUT3 #(
		.INIT('h07)
	) name4720 (
		_w2243_,
		_w2320_,
		_w6469_,
		_w6470_
	);
	LUT3 #(
		.INIT('h2a)
	) name4721 (
		rst_i_pad,
		_w2243_,
		_w6301_,
		_w6471_
	);
	LUT2 #(
		.INIT('hb)
	) name4722 (
		_w6470_,
		_w6471_,
		_w6472_
	);
	LUT4 #(
		.INIT('h10f0)
	) name4723 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u0_buf1_reg[19]/P0001 ,
		\u4_u0_ep_match_r_reg/P0001 ,
		_w6473_
	);
	LUT4 #(
		.INIT('hc800)
	) name4724 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_idin_reg[19]/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u0_ep_match_r_reg/P0001 ,
		_w6474_
	);
	LUT2 #(
		.INIT('h1)
	) name4725 (
		_w6473_,
		_w6474_,
		_w6475_
	);
	LUT3 #(
		.INIT('h07)
	) name4726 (
		_w2243_,
		_w2320_,
		_w6475_,
		_w6476_
	);
	LUT3 #(
		.INIT('h2a)
	) name4727 (
		rst_i_pad,
		_w2243_,
		_w6308_,
		_w6477_
	);
	LUT2 #(
		.INIT('hb)
	) name4728 (
		_w6476_,
		_w6477_,
		_w6478_
	);
	LUT4 #(
		.INIT('h10f0)
	) name4729 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u0_buf1_reg[1]/P0001 ,
		\u4_u0_ep_match_r_reg/P0001 ,
		_w6479_
	);
	LUT4 #(
		.INIT('hc800)
	) name4730 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_idin_reg[1]/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u0_ep_match_r_reg/P0001 ,
		_w6480_
	);
	LUT2 #(
		.INIT('h1)
	) name4731 (
		_w6479_,
		_w6480_,
		_w6481_
	);
	LUT3 #(
		.INIT('h07)
	) name4732 (
		_w2243_,
		_w2320_,
		_w6481_,
		_w6482_
	);
	LUT3 #(
		.INIT('h2a)
	) name4733 (
		rst_i_pad,
		_w2243_,
		_w6315_,
		_w6483_
	);
	LUT2 #(
		.INIT('hb)
	) name4734 (
		_w6482_,
		_w6483_,
		_w6484_
	);
	LUT4 #(
		.INIT('h10f0)
	) name4735 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u0_buf1_reg[20]/P0001 ,
		\u4_u0_ep_match_r_reg/P0001 ,
		_w6485_
	);
	LUT4 #(
		.INIT('hc800)
	) name4736 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_idin_reg[20]/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u0_ep_match_r_reg/P0001 ,
		_w6486_
	);
	LUT2 #(
		.INIT('h1)
	) name4737 (
		_w6485_,
		_w6486_,
		_w6487_
	);
	LUT3 #(
		.INIT('h07)
	) name4738 (
		_w2243_,
		_w2320_,
		_w6487_,
		_w6488_
	);
	LUT3 #(
		.INIT('h2a)
	) name4739 (
		rst_i_pad,
		_w2243_,
		_w6322_,
		_w6489_
	);
	LUT2 #(
		.INIT('hb)
	) name4740 (
		_w6488_,
		_w6489_,
		_w6490_
	);
	LUT4 #(
		.INIT('h10f0)
	) name4741 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u0_buf1_reg[21]/P0001 ,
		\u4_u0_ep_match_r_reg/P0001 ,
		_w6491_
	);
	LUT4 #(
		.INIT('hc800)
	) name4742 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_idin_reg[21]/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u0_ep_match_r_reg/P0001 ,
		_w6492_
	);
	LUT2 #(
		.INIT('h1)
	) name4743 (
		_w6491_,
		_w6492_,
		_w6493_
	);
	LUT3 #(
		.INIT('h07)
	) name4744 (
		_w2243_,
		_w2320_,
		_w6493_,
		_w6494_
	);
	LUT3 #(
		.INIT('h2a)
	) name4745 (
		rst_i_pad,
		_w2243_,
		_w6329_,
		_w6495_
	);
	LUT2 #(
		.INIT('hb)
	) name4746 (
		_w6494_,
		_w6495_,
		_w6496_
	);
	LUT4 #(
		.INIT('h10f0)
	) name4747 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u0_buf1_reg[22]/P0001 ,
		\u4_u0_ep_match_r_reg/P0001 ,
		_w6497_
	);
	LUT4 #(
		.INIT('hc800)
	) name4748 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_idin_reg[22]/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u0_ep_match_r_reg/P0001 ,
		_w6498_
	);
	LUT2 #(
		.INIT('h1)
	) name4749 (
		_w6497_,
		_w6498_,
		_w6499_
	);
	LUT3 #(
		.INIT('h07)
	) name4750 (
		_w2243_,
		_w2320_,
		_w6499_,
		_w6500_
	);
	LUT3 #(
		.INIT('h2a)
	) name4751 (
		rst_i_pad,
		_w2243_,
		_w6336_,
		_w6501_
	);
	LUT2 #(
		.INIT('hb)
	) name4752 (
		_w6500_,
		_w6501_,
		_w6502_
	);
	LUT4 #(
		.INIT('h10f0)
	) name4753 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u0_buf1_reg[23]/P0001 ,
		\u4_u0_ep_match_r_reg/P0001 ,
		_w6503_
	);
	LUT4 #(
		.INIT('hc800)
	) name4754 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_idin_reg[23]/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u0_ep_match_r_reg/P0001 ,
		_w6504_
	);
	LUT2 #(
		.INIT('h1)
	) name4755 (
		_w6503_,
		_w6504_,
		_w6505_
	);
	LUT3 #(
		.INIT('h07)
	) name4756 (
		_w2243_,
		_w2320_,
		_w6505_,
		_w6506_
	);
	LUT3 #(
		.INIT('h2a)
	) name4757 (
		rst_i_pad,
		_w2243_,
		_w6343_,
		_w6507_
	);
	LUT2 #(
		.INIT('hb)
	) name4758 (
		_w6506_,
		_w6507_,
		_w6508_
	);
	LUT4 #(
		.INIT('h10f0)
	) name4759 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u0_buf1_reg[24]/P0001 ,
		\u4_u0_ep_match_r_reg/P0001 ,
		_w6509_
	);
	LUT4 #(
		.INIT('hc800)
	) name4760 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_idin_reg[24]/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u0_ep_match_r_reg/P0001 ,
		_w6510_
	);
	LUT2 #(
		.INIT('h1)
	) name4761 (
		_w6509_,
		_w6510_,
		_w6511_
	);
	LUT3 #(
		.INIT('h07)
	) name4762 (
		_w2243_,
		_w2320_,
		_w6511_,
		_w6512_
	);
	LUT3 #(
		.INIT('h2a)
	) name4763 (
		rst_i_pad,
		_w2243_,
		_w6350_,
		_w6513_
	);
	LUT2 #(
		.INIT('hb)
	) name4764 (
		_w6512_,
		_w6513_,
		_w6514_
	);
	LUT4 #(
		.INIT('h10f0)
	) name4765 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u0_buf1_reg[25]/P0001 ,
		\u4_u0_ep_match_r_reg/P0001 ,
		_w6515_
	);
	LUT4 #(
		.INIT('hc800)
	) name4766 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_idin_reg[25]/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u0_ep_match_r_reg/P0001 ,
		_w6516_
	);
	LUT2 #(
		.INIT('h1)
	) name4767 (
		_w6515_,
		_w6516_,
		_w6517_
	);
	LUT3 #(
		.INIT('h07)
	) name4768 (
		_w2243_,
		_w2320_,
		_w6517_,
		_w6518_
	);
	LUT3 #(
		.INIT('h2a)
	) name4769 (
		rst_i_pad,
		_w2243_,
		_w6357_,
		_w6519_
	);
	LUT2 #(
		.INIT('hb)
	) name4770 (
		_w6518_,
		_w6519_,
		_w6520_
	);
	LUT4 #(
		.INIT('h8acf)
	) name4771 (
		\u4_buf1_reg[26]/NET0131 ,
		\u4_buf1_reg[27]/P0001 ,
		\u4_csr_reg[10]/P0001 ,
		\u4_csr_reg[9]/NET0131 ,
		_w6521_
	);
	LUT2 #(
		.INIT('h1)
	) name4772 (
		\u4_buf1_reg[28]/P0001 ,
		\u4_buf1_reg[29]/P0001 ,
		_w6522_
	);
	LUT3 #(
		.INIT('h31)
	) name4773 (
		\u4_buf1_reg[27]/P0001 ,
		\u4_buf1_reg[30]/P0001 ,
		\u4_csr_reg[10]/P0001 ,
		_w6523_
	);
	LUT3 #(
		.INIT('h40)
	) name4774 (
		_w6521_,
		_w6522_,
		_w6523_,
		_w6524_
	);
	LUT4 #(
		.INIT('h8caf)
	) name4775 (
		\u4_buf1_reg[24]/NET0131 ,
		\u4_buf1_reg[25]/NET0131 ,
		\u4_csr_reg[7]/P0001 ,
		\u4_csr_reg[8]/P0001 ,
		_w6525_
	);
	LUT4 #(
		.INIT('hf531)
	) name4776 (
		\u4_buf1_reg[23]/NET0131 ,
		\u4_buf1_reg[24]/NET0131 ,
		\u4_csr_reg[6]/NET0131 ,
		\u4_csr_reg[7]/P0001 ,
		_w6526_
	);
	LUT2 #(
		.INIT('h2)
	) name4777 (
		_w6525_,
		_w6526_,
		_w6527_
	);
	LUT4 #(
		.INIT('hf531)
	) name4778 (
		\u4_buf1_reg[21]/NET0131 ,
		\u4_buf1_reg[22]/NET0131 ,
		\u4_csr_reg[4]/NET0131 ,
		\u4_csr_reg[5]/NET0131 ,
		_w6528_
	);
	LUT4 #(
		.INIT('h8caf)
	) name4779 (
		\u4_buf1_reg[20]/NET0131 ,
		\u4_buf1_reg[21]/NET0131 ,
		\u4_csr_reg[3]/P0001 ,
		\u4_csr_reg[4]/NET0131 ,
		_w6529_
	);
	LUT2 #(
		.INIT('h2)
	) name4780 (
		_w6528_,
		_w6529_,
		_w6530_
	);
	LUT4 #(
		.INIT('h5010)
	) name4781 (
		\u4_buf1_reg[17]/NET0131 ,
		\u4_buf1_reg[18]/P0001 ,
		\u4_csr_reg[0]/P0001 ,
		\u4_csr_reg[1]/P0001 ,
		_w6531_
	);
	LUT4 #(
		.INIT('h8caf)
	) name4782 (
		\u4_buf1_reg[18]/P0001 ,
		\u4_buf1_reg[19]/NET0131 ,
		\u4_csr_reg[1]/P0001 ,
		\u4_csr_reg[2]/NET0131 ,
		_w6532_
	);
	LUT4 #(
		.INIT('hf531)
	) name4783 (
		\u4_buf1_reg[19]/NET0131 ,
		\u4_buf1_reg[20]/NET0131 ,
		\u4_csr_reg[2]/NET0131 ,
		\u4_csr_reg[3]/P0001 ,
		_w6533_
	);
	LUT4 #(
		.INIT('h8a00)
	) name4784 (
		_w6528_,
		_w6531_,
		_w6532_,
		_w6533_,
		_w6534_
	);
	LUT4 #(
		.INIT('h8caf)
	) name4785 (
		\u4_buf1_reg[22]/NET0131 ,
		\u4_buf1_reg[23]/NET0131 ,
		\u4_csr_reg[5]/NET0131 ,
		\u4_csr_reg[6]/NET0131 ,
		_w6535_
	);
	LUT2 #(
		.INIT('h8)
	) name4786 (
		_w6525_,
		_w6535_,
		_w6536_
	);
	LUT4 #(
		.INIT('h5455)
	) name4787 (
		_w6527_,
		_w6530_,
		_w6534_,
		_w6536_,
		_w6537_
	);
	LUT4 #(
		.INIT('hf531)
	) name4788 (
		\u4_buf1_reg[25]/NET0131 ,
		\u4_buf1_reg[26]/NET0131 ,
		\u4_csr_reg[8]/P0001 ,
		\u4_csr_reg[9]/NET0131 ,
		_w6538_
	);
	LUT3 #(
		.INIT('h80)
	) name4789 (
		_w6522_,
		_w6523_,
		_w6538_,
		_w6539_
	);
	LUT3 #(
		.INIT('hea)
	) name4790 (
		_w6524_,
		_w6537_,
		_w6539_,
		_w6540_
	);
	LUT4 #(
		.INIT('h10f0)
	) name4791 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u0_buf1_reg[26]/P0001 ,
		\u4_u0_ep_match_r_reg/P0001 ,
		_w6541_
	);
	LUT4 #(
		.INIT('hc800)
	) name4792 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_idin_reg[26]/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u0_ep_match_r_reg/P0001 ,
		_w6542_
	);
	LUT2 #(
		.INIT('h1)
	) name4793 (
		_w6541_,
		_w6542_,
		_w6543_
	);
	LUT3 #(
		.INIT('h07)
	) name4794 (
		_w2243_,
		_w2320_,
		_w6543_,
		_w6544_
	);
	LUT3 #(
		.INIT('h2a)
	) name4795 (
		rst_i_pad,
		_w2243_,
		_w6364_,
		_w6545_
	);
	LUT2 #(
		.INIT('hb)
	) name4796 (
		_w6544_,
		_w6545_,
		_w6546_
	);
	LUT4 #(
		.INIT('h10f0)
	) name4797 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u0_buf1_reg[27]/P0001 ,
		\u4_u0_ep_match_r_reg/P0001 ,
		_w6547_
	);
	LUT4 #(
		.INIT('hc800)
	) name4798 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_idin_reg[27]/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u0_ep_match_r_reg/P0001 ,
		_w6548_
	);
	LUT2 #(
		.INIT('h1)
	) name4799 (
		_w6547_,
		_w6548_,
		_w6549_
	);
	LUT3 #(
		.INIT('h07)
	) name4800 (
		_w2243_,
		_w2320_,
		_w6549_,
		_w6550_
	);
	LUT3 #(
		.INIT('h2a)
	) name4801 (
		rst_i_pad,
		_w2243_,
		_w6371_,
		_w6551_
	);
	LUT2 #(
		.INIT('hb)
	) name4802 (
		_w6550_,
		_w6551_,
		_w6552_
	);
	LUT4 #(
		.INIT('h10f0)
	) name4803 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u0_buf1_reg[28]/P0001 ,
		\u4_u0_ep_match_r_reg/P0001 ,
		_w6553_
	);
	LUT4 #(
		.INIT('hc800)
	) name4804 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_idin_reg[28]/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u0_ep_match_r_reg/P0001 ,
		_w6554_
	);
	LUT2 #(
		.INIT('h1)
	) name4805 (
		_w6553_,
		_w6554_,
		_w6555_
	);
	LUT3 #(
		.INIT('h07)
	) name4806 (
		_w2243_,
		_w2320_,
		_w6555_,
		_w6556_
	);
	LUT3 #(
		.INIT('h2a)
	) name4807 (
		rst_i_pad,
		_w2243_,
		_w6378_,
		_w6557_
	);
	LUT2 #(
		.INIT('hb)
	) name4808 (
		_w6556_,
		_w6557_,
		_w6558_
	);
	LUT4 #(
		.INIT('h10f0)
	) name4809 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u0_buf1_reg[29]/P0001 ,
		\u4_u0_ep_match_r_reg/P0001 ,
		_w6559_
	);
	LUT4 #(
		.INIT('hc800)
	) name4810 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_idin_reg[29]/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u0_ep_match_r_reg/P0001 ,
		_w6560_
	);
	LUT2 #(
		.INIT('h1)
	) name4811 (
		_w6559_,
		_w6560_,
		_w6561_
	);
	LUT3 #(
		.INIT('h07)
	) name4812 (
		_w2243_,
		_w2320_,
		_w6561_,
		_w6562_
	);
	LUT3 #(
		.INIT('h2a)
	) name4813 (
		rst_i_pad,
		_w2243_,
		_w6385_,
		_w6563_
	);
	LUT2 #(
		.INIT('hb)
	) name4814 (
		_w6562_,
		_w6563_,
		_w6564_
	);
	LUT4 #(
		.INIT('h10f0)
	) name4815 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u0_buf1_reg[2]/P0001 ,
		\u4_u0_ep_match_r_reg/P0001 ,
		_w6565_
	);
	LUT4 #(
		.INIT('hc800)
	) name4816 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_idin_reg[2]/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u0_ep_match_r_reg/P0001 ,
		_w6566_
	);
	LUT2 #(
		.INIT('h1)
	) name4817 (
		_w6565_,
		_w6566_,
		_w6567_
	);
	LUT3 #(
		.INIT('h07)
	) name4818 (
		_w2243_,
		_w2320_,
		_w6567_,
		_w6568_
	);
	LUT3 #(
		.INIT('h2a)
	) name4819 (
		rst_i_pad,
		_w2243_,
		_w6392_,
		_w6569_
	);
	LUT2 #(
		.INIT('hb)
	) name4820 (
		_w6568_,
		_w6569_,
		_w6570_
	);
	LUT4 #(
		.INIT('h10f0)
	) name4821 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u0_buf1_reg[30]/P0001 ,
		\u4_u0_ep_match_r_reg/P0001 ,
		_w6571_
	);
	LUT4 #(
		.INIT('hc800)
	) name4822 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_idin_reg[30]/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u0_ep_match_r_reg/P0001 ,
		_w6572_
	);
	LUT2 #(
		.INIT('h1)
	) name4823 (
		_w6571_,
		_w6572_,
		_w6573_
	);
	LUT3 #(
		.INIT('h07)
	) name4824 (
		_w2243_,
		_w2320_,
		_w6573_,
		_w6574_
	);
	LUT3 #(
		.INIT('h2a)
	) name4825 (
		rst_i_pad,
		_w2243_,
		_w6399_,
		_w6575_
	);
	LUT2 #(
		.INIT('hb)
	) name4826 (
		_w6574_,
		_w6575_,
		_w6576_
	);
	LUT4 #(
		.INIT('h10f0)
	) name4827 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u0_buf1_reg[31]/P0001 ,
		\u4_u0_ep_match_r_reg/P0001 ,
		_w6577_
	);
	LUT4 #(
		.INIT('hc800)
	) name4828 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_idin_reg[31]/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u0_ep_match_r_reg/P0001 ,
		_w6578_
	);
	LUT2 #(
		.INIT('h1)
	) name4829 (
		_w6577_,
		_w6578_,
		_w6579_
	);
	LUT3 #(
		.INIT('h07)
	) name4830 (
		_w2243_,
		_w2320_,
		_w6579_,
		_w6580_
	);
	LUT3 #(
		.INIT('h2a)
	) name4831 (
		rst_i_pad,
		_w2243_,
		_w6406_,
		_w6581_
	);
	LUT2 #(
		.INIT('hb)
	) name4832 (
		_w6580_,
		_w6581_,
		_w6582_
	);
	LUT4 #(
		.INIT('h10f0)
	) name4833 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u0_buf1_reg[3]/P0001 ,
		\u4_u0_ep_match_r_reg/P0001 ,
		_w6583_
	);
	LUT4 #(
		.INIT('hc800)
	) name4834 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_idin_reg[3]/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u0_ep_match_r_reg/P0001 ,
		_w6584_
	);
	LUT2 #(
		.INIT('h1)
	) name4835 (
		_w6583_,
		_w6584_,
		_w6585_
	);
	LUT3 #(
		.INIT('h07)
	) name4836 (
		_w2243_,
		_w2320_,
		_w6585_,
		_w6586_
	);
	LUT3 #(
		.INIT('h2a)
	) name4837 (
		rst_i_pad,
		_w2243_,
		_w6413_,
		_w6587_
	);
	LUT2 #(
		.INIT('hb)
	) name4838 (
		_w6586_,
		_w6587_,
		_w6588_
	);
	LUT4 #(
		.INIT('h10f0)
	) name4839 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u0_buf1_reg[8]/P0001 ,
		\u4_u0_ep_match_r_reg/P0001 ,
		_w6589_
	);
	LUT4 #(
		.INIT('hc800)
	) name4840 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_idin_reg[8]/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u0_ep_match_r_reg/P0001 ,
		_w6590_
	);
	LUT2 #(
		.INIT('h1)
	) name4841 (
		_w6589_,
		_w6590_,
		_w6591_
	);
	LUT3 #(
		.INIT('h07)
	) name4842 (
		_w2243_,
		_w2320_,
		_w6591_,
		_w6592_
	);
	LUT3 #(
		.INIT('h2a)
	) name4843 (
		rst_i_pad,
		_w2243_,
		_w6420_,
		_w6593_
	);
	LUT2 #(
		.INIT('hb)
	) name4844 (
		_w6592_,
		_w6593_,
		_w6594_
	);
	LUT4 #(
		.INIT('h10f0)
	) name4845 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u0_buf1_reg[9]/P0001 ,
		\u4_u0_ep_match_r_reg/P0001 ,
		_w6595_
	);
	LUT4 #(
		.INIT('hc800)
	) name4846 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_idin_reg[9]/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u0_ep_match_r_reg/P0001 ,
		_w6596_
	);
	LUT2 #(
		.INIT('h1)
	) name4847 (
		_w6595_,
		_w6596_,
		_w6597_
	);
	LUT3 #(
		.INIT('h07)
	) name4848 (
		_w2243_,
		_w2320_,
		_w6597_,
		_w6598_
	);
	LUT3 #(
		.INIT('h2a)
	) name4849 (
		rst_i_pad,
		_w2243_,
		_w6427_,
		_w6599_
	);
	LUT2 #(
		.INIT('hb)
	) name4850 (
		_w6598_,
		_w6599_,
		_w6600_
	);
	LUT3 #(
		.INIT('h10)
	) name4851 (
		\u0_u0_T1_gt_5_0_mS_reg/P0001 ,
		\u0_u0_idle_cnt1_next_reg[7]/P0001 ,
		\u0_u0_ps_cnt_clr_reg/P0001 ,
		_w6601_
	);
	LUT3 #(
		.INIT('h23)
	) name4852 (
		\u0_u0_T1_gt_5_0_mS_reg/P0001 ,
		\u0_u0_idle_cnt1_reg[7]/P0001 ,
		\u0_u0_ps_cnt_clr_reg/P0001 ,
		_w6602_
	);
	LUT3 #(
		.INIT('h02)
	) name4853 (
		_w5770_,
		_w6601_,
		_w6602_,
		_w6603_
	);
	LUT3 #(
		.INIT('hd0)
	) name4854 (
		_w5763_,
		_w5768_,
		_w6603_,
		_w6604_
	);
	LUT2 #(
		.INIT('h4)
	) name4855 (
		_w5765_,
		_w6604_,
		_w6605_
	);
	LUT4 #(
		.INIT('h10f0)
	) name4856 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u1_buf1_reg[0]/P0001 ,
		\u4_u1_ep_match_r_reg/P0001 ,
		_w6606_
	);
	LUT4 #(
		.INIT('hc800)
	) name4857 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_idin_reg[0]/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u1_ep_match_r_reg/P0001 ,
		_w6607_
	);
	LUT2 #(
		.INIT('h1)
	) name4858 (
		_w6606_,
		_w6607_,
		_w6608_
	);
	LUT3 #(
		.INIT('h07)
	) name4859 (
		_w2260_,
		_w2320_,
		_w6608_,
		_w6609_
	);
	LUT3 #(
		.INIT('h2a)
	) name4860 (
		rst_i_pad,
		_w2260_,
		_w6273_,
		_w6610_
	);
	LUT2 #(
		.INIT('hb)
	) name4861 (
		_w6609_,
		_w6610_,
		_w6611_
	);
	LUT4 #(
		.INIT('h10f0)
	) name4862 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u1_buf1_reg[12]/P0001 ,
		\u4_u1_ep_match_r_reg/P0001 ,
		_w6612_
	);
	LUT4 #(
		.INIT('hc800)
	) name4863 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_idin_reg[12]/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u1_ep_match_r_reg/P0001 ,
		_w6613_
	);
	LUT2 #(
		.INIT('h1)
	) name4864 (
		_w6612_,
		_w6613_,
		_w6614_
	);
	LUT3 #(
		.INIT('h07)
	) name4865 (
		_w2260_,
		_w2320_,
		_w6614_,
		_w6615_
	);
	LUT3 #(
		.INIT('h2a)
	) name4866 (
		rst_i_pad,
		_w2260_,
		_w6280_,
		_w6616_
	);
	LUT2 #(
		.INIT('hb)
	) name4867 (
		_w6615_,
		_w6616_,
		_w6617_
	);
	LUT4 #(
		.INIT('h10f0)
	) name4868 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u1_buf1_reg[16]/P0001 ,
		\u4_u1_ep_match_r_reg/P0001 ,
		_w6618_
	);
	LUT4 #(
		.INIT('hc800)
	) name4869 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_idin_reg[16]/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u1_ep_match_r_reg/P0001 ,
		_w6619_
	);
	LUT2 #(
		.INIT('h1)
	) name4870 (
		_w6618_,
		_w6619_,
		_w6620_
	);
	LUT3 #(
		.INIT('h07)
	) name4871 (
		_w2260_,
		_w2320_,
		_w6620_,
		_w6621_
	);
	LUT3 #(
		.INIT('h2a)
	) name4872 (
		rst_i_pad,
		_w2260_,
		_w6287_,
		_w6622_
	);
	LUT2 #(
		.INIT('hb)
	) name4873 (
		_w6621_,
		_w6622_,
		_w6623_
	);
	LUT4 #(
		.INIT('h10f0)
	) name4874 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u1_buf1_reg[17]/P0001 ,
		\u4_u1_ep_match_r_reg/P0001 ,
		_w6624_
	);
	LUT4 #(
		.INIT('hc800)
	) name4875 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_idin_reg[17]/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u1_ep_match_r_reg/P0001 ,
		_w6625_
	);
	LUT2 #(
		.INIT('h1)
	) name4876 (
		_w6624_,
		_w6625_,
		_w6626_
	);
	LUT3 #(
		.INIT('h07)
	) name4877 (
		_w2260_,
		_w2320_,
		_w6626_,
		_w6627_
	);
	LUT3 #(
		.INIT('h2a)
	) name4878 (
		rst_i_pad,
		_w2260_,
		_w6294_,
		_w6628_
	);
	LUT2 #(
		.INIT('hb)
	) name4879 (
		_w6627_,
		_w6628_,
		_w6629_
	);
	LUT4 #(
		.INIT('h10f0)
	) name4880 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u1_buf1_reg[18]/P0001 ,
		\u4_u1_ep_match_r_reg/P0001 ,
		_w6630_
	);
	LUT4 #(
		.INIT('hc800)
	) name4881 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_idin_reg[18]/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u1_ep_match_r_reg/P0001 ,
		_w6631_
	);
	LUT2 #(
		.INIT('h1)
	) name4882 (
		_w6630_,
		_w6631_,
		_w6632_
	);
	LUT3 #(
		.INIT('h07)
	) name4883 (
		_w2260_,
		_w2320_,
		_w6632_,
		_w6633_
	);
	LUT3 #(
		.INIT('h2a)
	) name4884 (
		rst_i_pad,
		_w2260_,
		_w6301_,
		_w6634_
	);
	LUT2 #(
		.INIT('hb)
	) name4885 (
		_w6633_,
		_w6634_,
		_w6635_
	);
	LUT4 #(
		.INIT('h10f0)
	) name4886 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u1_buf1_reg[19]/P0001 ,
		\u4_u1_ep_match_r_reg/P0001 ,
		_w6636_
	);
	LUT4 #(
		.INIT('hc800)
	) name4887 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_idin_reg[19]/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u1_ep_match_r_reg/P0001 ,
		_w6637_
	);
	LUT2 #(
		.INIT('h1)
	) name4888 (
		_w6636_,
		_w6637_,
		_w6638_
	);
	LUT3 #(
		.INIT('h07)
	) name4889 (
		_w2260_,
		_w2320_,
		_w6638_,
		_w6639_
	);
	LUT3 #(
		.INIT('h2a)
	) name4890 (
		rst_i_pad,
		_w2260_,
		_w6308_,
		_w6640_
	);
	LUT2 #(
		.INIT('hb)
	) name4891 (
		_w6639_,
		_w6640_,
		_w6641_
	);
	LUT4 #(
		.INIT('h10f0)
	) name4892 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u1_buf1_reg[1]/P0001 ,
		\u4_u1_ep_match_r_reg/P0001 ,
		_w6642_
	);
	LUT4 #(
		.INIT('hc800)
	) name4893 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_idin_reg[1]/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u1_ep_match_r_reg/P0001 ,
		_w6643_
	);
	LUT2 #(
		.INIT('h1)
	) name4894 (
		_w6642_,
		_w6643_,
		_w6644_
	);
	LUT3 #(
		.INIT('h07)
	) name4895 (
		_w2260_,
		_w2320_,
		_w6644_,
		_w6645_
	);
	LUT3 #(
		.INIT('h2a)
	) name4896 (
		rst_i_pad,
		_w2260_,
		_w6315_,
		_w6646_
	);
	LUT2 #(
		.INIT('hb)
	) name4897 (
		_w6645_,
		_w6646_,
		_w6647_
	);
	LUT4 #(
		.INIT('h10f0)
	) name4898 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u1_buf1_reg[20]/P0001 ,
		\u4_u1_ep_match_r_reg/P0001 ,
		_w6648_
	);
	LUT4 #(
		.INIT('hc800)
	) name4899 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_idin_reg[20]/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u1_ep_match_r_reg/P0001 ,
		_w6649_
	);
	LUT2 #(
		.INIT('h1)
	) name4900 (
		_w6648_,
		_w6649_,
		_w6650_
	);
	LUT3 #(
		.INIT('h07)
	) name4901 (
		_w2260_,
		_w2320_,
		_w6650_,
		_w6651_
	);
	LUT3 #(
		.INIT('h2a)
	) name4902 (
		rst_i_pad,
		_w2260_,
		_w6322_,
		_w6652_
	);
	LUT2 #(
		.INIT('hb)
	) name4903 (
		_w6651_,
		_w6652_,
		_w6653_
	);
	LUT4 #(
		.INIT('h10f0)
	) name4904 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u1_buf1_reg[21]/P0001 ,
		\u4_u1_ep_match_r_reg/P0001 ,
		_w6654_
	);
	LUT4 #(
		.INIT('hc800)
	) name4905 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_idin_reg[21]/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u1_ep_match_r_reg/P0001 ,
		_w6655_
	);
	LUT2 #(
		.INIT('h1)
	) name4906 (
		_w6654_,
		_w6655_,
		_w6656_
	);
	LUT3 #(
		.INIT('h07)
	) name4907 (
		_w2260_,
		_w2320_,
		_w6656_,
		_w6657_
	);
	LUT3 #(
		.INIT('h2a)
	) name4908 (
		rst_i_pad,
		_w2260_,
		_w6329_,
		_w6658_
	);
	LUT2 #(
		.INIT('hb)
	) name4909 (
		_w6657_,
		_w6658_,
		_w6659_
	);
	LUT4 #(
		.INIT('h10f0)
	) name4910 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u1_buf1_reg[22]/P0001 ,
		\u4_u1_ep_match_r_reg/P0001 ,
		_w6660_
	);
	LUT4 #(
		.INIT('hc800)
	) name4911 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_idin_reg[22]/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u1_ep_match_r_reg/P0001 ,
		_w6661_
	);
	LUT2 #(
		.INIT('h1)
	) name4912 (
		_w6660_,
		_w6661_,
		_w6662_
	);
	LUT3 #(
		.INIT('h07)
	) name4913 (
		_w2260_,
		_w2320_,
		_w6662_,
		_w6663_
	);
	LUT3 #(
		.INIT('h2a)
	) name4914 (
		rst_i_pad,
		_w2260_,
		_w6336_,
		_w6664_
	);
	LUT2 #(
		.INIT('hb)
	) name4915 (
		_w6663_,
		_w6664_,
		_w6665_
	);
	LUT4 #(
		.INIT('h10f0)
	) name4916 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u1_buf1_reg[23]/P0001 ,
		\u4_u1_ep_match_r_reg/P0001 ,
		_w6666_
	);
	LUT4 #(
		.INIT('hc800)
	) name4917 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_idin_reg[23]/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u1_ep_match_r_reg/P0001 ,
		_w6667_
	);
	LUT2 #(
		.INIT('h1)
	) name4918 (
		_w6666_,
		_w6667_,
		_w6668_
	);
	LUT3 #(
		.INIT('h07)
	) name4919 (
		_w2260_,
		_w2320_,
		_w6668_,
		_w6669_
	);
	LUT3 #(
		.INIT('h2a)
	) name4920 (
		rst_i_pad,
		_w2260_,
		_w6343_,
		_w6670_
	);
	LUT2 #(
		.INIT('hb)
	) name4921 (
		_w6669_,
		_w6670_,
		_w6671_
	);
	LUT4 #(
		.INIT('h10f0)
	) name4922 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u1_buf1_reg[24]/P0001 ,
		\u4_u1_ep_match_r_reg/P0001 ,
		_w6672_
	);
	LUT4 #(
		.INIT('hc800)
	) name4923 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_idin_reg[24]/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u1_ep_match_r_reg/P0001 ,
		_w6673_
	);
	LUT2 #(
		.INIT('h1)
	) name4924 (
		_w6672_,
		_w6673_,
		_w6674_
	);
	LUT3 #(
		.INIT('h07)
	) name4925 (
		_w2260_,
		_w2320_,
		_w6674_,
		_w6675_
	);
	LUT3 #(
		.INIT('h2a)
	) name4926 (
		rst_i_pad,
		_w2260_,
		_w6350_,
		_w6676_
	);
	LUT2 #(
		.INIT('hb)
	) name4927 (
		_w6675_,
		_w6676_,
		_w6677_
	);
	LUT4 #(
		.INIT('h10f0)
	) name4928 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u1_buf1_reg[25]/P0001 ,
		\u4_u1_ep_match_r_reg/P0001 ,
		_w6678_
	);
	LUT4 #(
		.INIT('hc800)
	) name4929 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_idin_reg[25]/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u1_ep_match_r_reg/P0001 ,
		_w6679_
	);
	LUT2 #(
		.INIT('h1)
	) name4930 (
		_w6678_,
		_w6679_,
		_w6680_
	);
	LUT3 #(
		.INIT('h07)
	) name4931 (
		_w2260_,
		_w2320_,
		_w6680_,
		_w6681_
	);
	LUT3 #(
		.INIT('h2a)
	) name4932 (
		rst_i_pad,
		_w2260_,
		_w6357_,
		_w6682_
	);
	LUT2 #(
		.INIT('hb)
	) name4933 (
		_w6681_,
		_w6682_,
		_w6683_
	);
	LUT4 #(
		.INIT('h10f0)
	) name4934 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u1_buf1_reg[26]/P0001 ,
		\u4_u1_ep_match_r_reg/P0001 ,
		_w6684_
	);
	LUT4 #(
		.INIT('hc800)
	) name4935 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_idin_reg[26]/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u1_ep_match_r_reg/P0001 ,
		_w6685_
	);
	LUT2 #(
		.INIT('h1)
	) name4936 (
		_w6684_,
		_w6685_,
		_w6686_
	);
	LUT3 #(
		.INIT('h07)
	) name4937 (
		_w2260_,
		_w2320_,
		_w6686_,
		_w6687_
	);
	LUT3 #(
		.INIT('h2a)
	) name4938 (
		rst_i_pad,
		_w2260_,
		_w6364_,
		_w6688_
	);
	LUT2 #(
		.INIT('hb)
	) name4939 (
		_w6687_,
		_w6688_,
		_w6689_
	);
	LUT4 #(
		.INIT('h10f0)
	) name4940 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u1_buf1_reg[27]/P0001 ,
		\u4_u1_ep_match_r_reg/P0001 ,
		_w6690_
	);
	LUT4 #(
		.INIT('hc800)
	) name4941 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_idin_reg[27]/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u1_ep_match_r_reg/P0001 ,
		_w6691_
	);
	LUT2 #(
		.INIT('h1)
	) name4942 (
		_w6690_,
		_w6691_,
		_w6692_
	);
	LUT3 #(
		.INIT('h07)
	) name4943 (
		_w2260_,
		_w2320_,
		_w6692_,
		_w6693_
	);
	LUT3 #(
		.INIT('h2a)
	) name4944 (
		rst_i_pad,
		_w2260_,
		_w6371_,
		_w6694_
	);
	LUT2 #(
		.INIT('hb)
	) name4945 (
		_w6693_,
		_w6694_,
		_w6695_
	);
	LUT4 #(
		.INIT('h10f0)
	) name4946 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u1_buf1_reg[28]/P0001 ,
		\u4_u1_ep_match_r_reg/P0001 ,
		_w6696_
	);
	LUT4 #(
		.INIT('hc800)
	) name4947 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_idin_reg[28]/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u1_ep_match_r_reg/P0001 ,
		_w6697_
	);
	LUT2 #(
		.INIT('h1)
	) name4948 (
		_w6696_,
		_w6697_,
		_w6698_
	);
	LUT3 #(
		.INIT('h07)
	) name4949 (
		_w2260_,
		_w2320_,
		_w6698_,
		_w6699_
	);
	LUT3 #(
		.INIT('h2a)
	) name4950 (
		rst_i_pad,
		_w2260_,
		_w6378_,
		_w6700_
	);
	LUT2 #(
		.INIT('hb)
	) name4951 (
		_w6699_,
		_w6700_,
		_w6701_
	);
	LUT4 #(
		.INIT('h10f0)
	) name4952 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u1_buf1_reg[29]/P0001 ,
		\u4_u1_ep_match_r_reg/P0001 ,
		_w6702_
	);
	LUT4 #(
		.INIT('hc800)
	) name4953 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_idin_reg[29]/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u1_ep_match_r_reg/P0001 ,
		_w6703_
	);
	LUT2 #(
		.INIT('h1)
	) name4954 (
		_w6702_,
		_w6703_,
		_w6704_
	);
	LUT3 #(
		.INIT('h07)
	) name4955 (
		_w2260_,
		_w2320_,
		_w6704_,
		_w6705_
	);
	LUT3 #(
		.INIT('h2a)
	) name4956 (
		rst_i_pad,
		_w2260_,
		_w6385_,
		_w6706_
	);
	LUT2 #(
		.INIT('hb)
	) name4957 (
		_w6705_,
		_w6706_,
		_w6707_
	);
	LUT4 #(
		.INIT('h10f0)
	) name4958 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u1_buf1_reg[2]/P0001 ,
		\u4_u1_ep_match_r_reg/P0001 ,
		_w6708_
	);
	LUT4 #(
		.INIT('hc800)
	) name4959 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_idin_reg[2]/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u1_ep_match_r_reg/P0001 ,
		_w6709_
	);
	LUT2 #(
		.INIT('h1)
	) name4960 (
		_w6708_,
		_w6709_,
		_w6710_
	);
	LUT3 #(
		.INIT('h07)
	) name4961 (
		_w2260_,
		_w2320_,
		_w6710_,
		_w6711_
	);
	LUT3 #(
		.INIT('h2a)
	) name4962 (
		rst_i_pad,
		_w2260_,
		_w6392_,
		_w6712_
	);
	LUT2 #(
		.INIT('hb)
	) name4963 (
		_w6711_,
		_w6712_,
		_w6713_
	);
	LUT4 #(
		.INIT('h10f0)
	) name4964 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u1_buf1_reg[30]/P0001 ,
		\u4_u1_ep_match_r_reg/P0001 ,
		_w6714_
	);
	LUT4 #(
		.INIT('hc800)
	) name4965 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_idin_reg[30]/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u1_ep_match_r_reg/P0001 ,
		_w6715_
	);
	LUT2 #(
		.INIT('h1)
	) name4966 (
		_w6714_,
		_w6715_,
		_w6716_
	);
	LUT3 #(
		.INIT('h07)
	) name4967 (
		_w2260_,
		_w2320_,
		_w6716_,
		_w6717_
	);
	LUT3 #(
		.INIT('h2a)
	) name4968 (
		rst_i_pad,
		_w2260_,
		_w6399_,
		_w6718_
	);
	LUT2 #(
		.INIT('hb)
	) name4969 (
		_w6717_,
		_w6718_,
		_w6719_
	);
	LUT4 #(
		.INIT('h10f0)
	) name4970 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u1_buf1_reg[31]/P0001 ,
		\u4_u1_ep_match_r_reg/P0001 ,
		_w6720_
	);
	LUT4 #(
		.INIT('hc800)
	) name4971 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_idin_reg[31]/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u1_ep_match_r_reg/P0001 ,
		_w6721_
	);
	LUT2 #(
		.INIT('h1)
	) name4972 (
		_w6720_,
		_w6721_,
		_w6722_
	);
	LUT3 #(
		.INIT('h07)
	) name4973 (
		_w2260_,
		_w2320_,
		_w6722_,
		_w6723_
	);
	LUT3 #(
		.INIT('h2a)
	) name4974 (
		rst_i_pad,
		_w2260_,
		_w6406_,
		_w6724_
	);
	LUT2 #(
		.INIT('hb)
	) name4975 (
		_w6723_,
		_w6724_,
		_w6725_
	);
	LUT4 #(
		.INIT('h10f0)
	) name4976 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u1_buf1_reg[3]/P0001 ,
		\u4_u1_ep_match_r_reg/P0001 ,
		_w6726_
	);
	LUT4 #(
		.INIT('hc800)
	) name4977 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_idin_reg[3]/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u1_ep_match_r_reg/P0001 ,
		_w6727_
	);
	LUT2 #(
		.INIT('h1)
	) name4978 (
		_w6726_,
		_w6727_,
		_w6728_
	);
	LUT3 #(
		.INIT('h07)
	) name4979 (
		_w2260_,
		_w2320_,
		_w6728_,
		_w6729_
	);
	LUT3 #(
		.INIT('h2a)
	) name4980 (
		rst_i_pad,
		_w2260_,
		_w6413_,
		_w6730_
	);
	LUT2 #(
		.INIT('hb)
	) name4981 (
		_w6729_,
		_w6730_,
		_w6731_
	);
	LUT4 #(
		.INIT('h10f0)
	) name4982 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u1_buf1_reg[8]/P0001 ,
		\u4_u1_ep_match_r_reg/P0001 ,
		_w6732_
	);
	LUT4 #(
		.INIT('hc800)
	) name4983 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_idin_reg[8]/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u1_ep_match_r_reg/P0001 ,
		_w6733_
	);
	LUT2 #(
		.INIT('h1)
	) name4984 (
		_w6732_,
		_w6733_,
		_w6734_
	);
	LUT3 #(
		.INIT('h07)
	) name4985 (
		_w2260_,
		_w2320_,
		_w6734_,
		_w6735_
	);
	LUT3 #(
		.INIT('h2a)
	) name4986 (
		rst_i_pad,
		_w2260_,
		_w6420_,
		_w6736_
	);
	LUT2 #(
		.INIT('hb)
	) name4987 (
		_w6735_,
		_w6736_,
		_w6737_
	);
	LUT4 #(
		.INIT('h10f0)
	) name4988 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u1_buf1_reg[9]/P0001 ,
		\u4_u1_ep_match_r_reg/P0001 ,
		_w6738_
	);
	LUT4 #(
		.INIT('hc800)
	) name4989 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_idin_reg[9]/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u1_ep_match_r_reg/P0001 ,
		_w6739_
	);
	LUT2 #(
		.INIT('h1)
	) name4990 (
		_w6738_,
		_w6739_,
		_w6740_
	);
	LUT3 #(
		.INIT('h07)
	) name4991 (
		_w2260_,
		_w2320_,
		_w6740_,
		_w6741_
	);
	LUT3 #(
		.INIT('h2a)
	) name4992 (
		rst_i_pad,
		_w2260_,
		_w6427_,
		_w6742_
	);
	LUT2 #(
		.INIT('hb)
	) name4993 (
		_w6741_,
		_w6742_,
		_w6743_
	);
	LUT4 #(
		.INIT('h10f0)
	) name4994 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u2_buf1_reg[0]/P0001 ,
		\u4_u2_ep_match_r_reg/P0001 ,
		_w6744_
	);
	LUT4 #(
		.INIT('hc800)
	) name4995 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_idin_reg[0]/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u2_ep_match_r_reg/P0001 ,
		_w6745_
	);
	LUT2 #(
		.INIT('h1)
	) name4996 (
		_w6744_,
		_w6745_,
		_w6746_
	);
	LUT3 #(
		.INIT('h07)
	) name4997 (
		_w2267_,
		_w2320_,
		_w6746_,
		_w6747_
	);
	LUT3 #(
		.INIT('h2a)
	) name4998 (
		rst_i_pad,
		_w2267_,
		_w6273_,
		_w6748_
	);
	LUT2 #(
		.INIT('hb)
	) name4999 (
		_w6747_,
		_w6748_,
		_w6749_
	);
	LUT4 #(
		.INIT('h10f0)
	) name5000 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u2_buf1_reg[12]/P0001 ,
		\u4_u2_ep_match_r_reg/P0001 ,
		_w6750_
	);
	LUT4 #(
		.INIT('hc800)
	) name5001 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_idin_reg[12]/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u2_ep_match_r_reg/P0001 ,
		_w6751_
	);
	LUT2 #(
		.INIT('h1)
	) name5002 (
		_w6750_,
		_w6751_,
		_w6752_
	);
	LUT3 #(
		.INIT('h07)
	) name5003 (
		_w2267_,
		_w2320_,
		_w6752_,
		_w6753_
	);
	LUT3 #(
		.INIT('h2a)
	) name5004 (
		rst_i_pad,
		_w2267_,
		_w6280_,
		_w6754_
	);
	LUT2 #(
		.INIT('hb)
	) name5005 (
		_w6753_,
		_w6754_,
		_w6755_
	);
	LUT4 #(
		.INIT('h10f0)
	) name5006 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u2_buf1_reg[16]/P0001 ,
		\u4_u2_ep_match_r_reg/P0001 ,
		_w6756_
	);
	LUT4 #(
		.INIT('hc800)
	) name5007 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_idin_reg[16]/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u2_ep_match_r_reg/P0001 ,
		_w6757_
	);
	LUT2 #(
		.INIT('h1)
	) name5008 (
		_w6756_,
		_w6757_,
		_w6758_
	);
	LUT3 #(
		.INIT('h07)
	) name5009 (
		_w2267_,
		_w2320_,
		_w6758_,
		_w6759_
	);
	LUT3 #(
		.INIT('h2a)
	) name5010 (
		rst_i_pad,
		_w2267_,
		_w6287_,
		_w6760_
	);
	LUT2 #(
		.INIT('hb)
	) name5011 (
		_w6759_,
		_w6760_,
		_w6761_
	);
	LUT4 #(
		.INIT('h10f0)
	) name5012 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u2_buf1_reg[17]/P0001 ,
		\u4_u2_ep_match_r_reg/P0001 ,
		_w6762_
	);
	LUT4 #(
		.INIT('hc800)
	) name5013 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_idin_reg[17]/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u2_ep_match_r_reg/P0001 ,
		_w6763_
	);
	LUT2 #(
		.INIT('h1)
	) name5014 (
		_w6762_,
		_w6763_,
		_w6764_
	);
	LUT3 #(
		.INIT('h07)
	) name5015 (
		_w2267_,
		_w2320_,
		_w6764_,
		_w6765_
	);
	LUT3 #(
		.INIT('h2a)
	) name5016 (
		rst_i_pad,
		_w2267_,
		_w6294_,
		_w6766_
	);
	LUT2 #(
		.INIT('hb)
	) name5017 (
		_w6765_,
		_w6766_,
		_w6767_
	);
	LUT4 #(
		.INIT('h10f0)
	) name5018 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u2_buf1_reg[18]/P0001 ,
		\u4_u2_ep_match_r_reg/P0001 ,
		_w6768_
	);
	LUT4 #(
		.INIT('hc800)
	) name5019 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_idin_reg[18]/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u2_ep_match_r_reg/P0001 ,
		_w6769_
	);
	LUT2 #(
		.INIT('h1)
	) name5020 (
		_w6768_,
		_w6769_,
		_w6770_
	);
	LUT3 #(
		.INIT('h07)
	) name5021 (
		_w2267_,
		_w2320_,
		_w6770_,
		_w6771_
	);
	LUT3 #(
		.INIT('h2a)
	) name5022 (
		rst_i_pad,
		_w2267_,
		_w6301_,
		_w6772_
	);
	LUT2 #(
		.INIT('hb)
	) name5023 (
		_w6771_,
		_w6772_,
		_w6773_
	);
	LUT4 #(
		.INIT('h10f0)
	) name5024 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u2_buf1_reg[19]/P0001 ,
		\u4_u2_ep_match_r_reg/P0001 ,
		_w6774_
	);
	LUT4 #(
		.INIT('hc800)
	) name5025 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_idin_reg[19]/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u2_ep_match_r_reg/P0001 ,
		_w6775_
	);
	LUT2 #(
		.INIT('h1)
	) name5026 (
		_w6774_,
		_w6775_,
		_w6776_
	);
	LUT3 #(
		.INIT('h07)
	) name5027 (
		_w2267_,
		_w2320_,
		_w6776_,
		_w6777_
	);
	LUT3 #(
		.INIT('h2a)
	) name5028 (
		rst_i_pad,
		_w2267_,
		_w6308_,
		_w6778_
	);
	LUT2 #(
		.INIT('hb)
	) name5029 (
		_w6777_,
		_w6778_,
		_w6779_
	);
	LUT4 #(
		.INIT('h10f0)
	) name5030 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u2_buf1_reg[1]/P0001 ,
		\u4_u2_ep_match_r_reg/P0001 ,
		_w6780_
	);
	LUT4 #(
		.INIT('hc800)
	) name5031 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_idin_reg[1]/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u2_ep_match_r_reg/P0001 ,
		_w6781_
	);
	LUT2 #(
		.INIT('h1)
	) name5032 (
		_w6780_,
		_w6781_,
		_w6782_
	);
	LUT3 #(
		.INIT('h07)
	) name5033 (
		_w2267_,
		_w2320_,
		_w6782_,
		_w6783_
	);
	LUT3 #(
		.INIT('h2a)
	) name5034 (
		rst_i_pad,
		_w2267_,
		_w6315_,
		_w6784_
	);
	LUT2 #(
		.INIT('hb)
	) name5035 (
		_w6783_,
		_w6784_,
		_w6785_
	);
	LUT4 #(
		.INIT('h10f0)
	) name5036 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u2_buf1_reg[20]/P0001 ,
		\u4_u2_ep_match_r_reg/P0001 ,
		_w6786_
	);
	LUT4 #(
		.INIT('hc800)
	) name5037 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_idin_reg[20]/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u2_ep_match_r_reg/P0001 ,
		_w6787_
	);
	LUT2 #(
		.INIT('h1)
	) name5038 (
		_w6786_,
		_w6787_,
		_w6788_
	);
	LUT3 #(
		.INIT('h07)
	) name5039 (
		_w2267_,
		_w2320_,
		_w6788_,
		_w6789_
	);
	LUT3 #(
		.INIT('h2a)
	) name5040 (
		rst_i_pad,
		_w2267_,
		_w6322_,
		_w6790_
	);
	LUT2 #(
		.INIT('hb)
	) name5041 (
		_w6789_,
		_w6790_,
		_w6791_
	);
	LUT4 #(
		.INIT('h10f0)
	) name5042 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u2_buf1_reg[21]/P0001 ,
		\u4_u2_ep_match_r_reg/P0001 ,
		_w6792_
	);
	LUT4 #(
		.INIT('hc800)
	) name5043 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_idin_reg[21]/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u2_ep_match_r_reg/P0001 ,
		_w6793_
	);
	LUT2 #(
		.INIT('h1)
	) name5044 (
		_w6792_,
		_w6793_,
		_w6794_
	);
	LUT3 #(
		.INIT('h07)
	) name5045 (
		_w2267_,
		_w2320_,
		_w6794_,
		_w6795_
	);
	LUT3 #(
		.INIT('h2a)
	) name5046 (
		rst_i_pad,
		_w2267_,
		_w6329_,
		_w6796_
	);
	LUT2 #(
		.INIT('hb)
	) name5047 (
		_w6795_,
		_w6796_,
		_w6797_
	);
	LUT4 #(
		.INIT('h10f0)
	) name5048 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u2_buf1_reg[22]/P0001 ,
		\u4_u2_ep_match_r_reg/P0001 ,
		_w6798_
	);
	LUT4 #(
		.INIT('hc800)
	) name5049 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_idin_reg[22]/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u2_ep_match_r_reg/P0001 ,
		_w6799_
	);
	LUT2 #(
		.INIT('h1)
	) name5050 (
		_w6798_,
		_w6799_,
		_w6800_
	);
	LUT3 #(
		.INIT('h07)
	) name5051 (
		_w2267_,
		_w2320_,
		_w6800_,
		_w6801_
	);
	LUT3 #(
		.INIT('h2a)
	) name5052 (
		rst_i_pad,
		_w2267_,
		_w6336_,
		_w6802_
	);
	LUT2 #(
		.INIT('hb)
	) name5053 (
		_w6801_,
		_w6802_,
		_w6803_
	);
	LUT4 #(
		.INIT('h10f0)
	) name5054 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u2_buf1_reg[23]/P0001 ,
		\u4_u2_ep_match_r_reg/P0001 ,
		_w6804_
	);
	LUT4 #(
		.INIT('hc800)
	) name5055 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_idin_reg[23]/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u2_ep_match_r_reg/P0001 ,
		_w6805_
	);
	LUT2 #(
		.INIT('h1)
	) name5056 (
		_w6804_,
		_w6805_,
		_w6806_
	);
	LUT3 #(
		.INIT('h07)
	) name5057 (
		_w2267_,
		_w2320_,
		_w6806_,
		_w6807_
	);
	LUT3 #(
		.INIT('h2a)
	) name5058 (
		rst_i_pad,
		_w2267_,
		_w6343_,
		_w6808_
	);
	LUT2 #(
		.INIT('hb)
	) name5059 (
		_w6807_,
		_w6808_,
		_w6809_
	);
	LUT4 #(
		.INIT('h10f0)
	) name5060 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u2_buf1_reg[24]/P0001 ,
		\u4_u2_ep_match_r_reg/P0001 ,
		_w6810_
	);
	LUT4 #(
		.INIT('hc800)
	) name5061 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_idin_reg[24]/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u2_ep_match_r_reg/P0001 ,
		_w6811_
	);
	LUT2 #(
		.INIT('h1)
	) name5062 (
		_w6810_,
		_w6811_,
		_w6812_
	);
	LUT3 #(
		.INIT('h07)
	) name5063 (
		_w2267_,
		_w2320_,
		_w6812_,
		_w6813_
	);
	LUT3 #(
		.INIT('h2a)
	) name5064 (
		rst_i_pad,
		_w2267_,
		_w6350_,
		_w6814_
	);
	LUT2 #(
		.INIT('hb)
	) name5065 (
		_w6813_,
		_w6814_,
		_w6815_
	);
	LUT4 #(
		.INIT('h10f0)
	) name5066 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u2_buf1_reg[25]/P0001 ,
		\u4_u2_ep_match_r_reg/P0001 ,
		_w6816_
	);
	LUT4 #(
		.INIT('hc800)
	) name5067 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_idin_reg[25]/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u2_ep_match_r_reg/P0001 ,
		_w6817_
	);
	LUT2 #(
		.INIT('h1)
	) name5068 (
		_w6816_,
		_w6817_,
		_w6818_
	);
	LUT3 #(
		.INIT('h07)
	) name5069 (
		_w2267_,
		_w2320_,
		_w6818_,
		_w6819_
	);
	LUT3 #(
		.INIT('h2a)
	) name5070 (
		rst_i_pad,
		_w2267_,
		_w6357_,
		_w6820_
	);
	LUT2 #(
		.INIT('hb)
	) name5071 (
		_w6819_,
		_w6820_,
		_w6821_
	);
	LUT4 #(
		.INIT('h10f0)
	) name5072 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u2_buf1_reg[26]/P0001 ,
		\u4_u2_ep_match_r_reg/P0001 ,
		_w6822_
	);
	LUT4 #(
		.INIT('hc800)
	) name5073 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_idin_reg[26]/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u2_ep_match_r_reg/P0001 ,
		_w6823_
	);
	LUT2 #(
		.INIT('h1)
	) name5074 (
		_w6822_,
		_w6823_,
		_w6824_
	);
	LUT3 #(
		.INIT('h07)
	) name5075 (
		_w2267_,
		_w2320_,
		_w6824_,
		_w6825_
	);
	LUT3 #(
		.INIT('h2a)
	) name5076 (
		rst_i_pad,
		_w2267_,
		_w6364_,
		_w6826_
	);
	LUT2 #(
		.INIT('hb)
	) name5077 (
		_w6825_,
		_w6826_,
		_w6827_
	);
	LUT4 #(
		.INIT('h10f0)
	) name5078 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u2_buf1_reg[27]/P0001 ,
		\u4_u2_ep_match_r_reg/P0001 ,
		_w6828_
	);
	LUT4 #(
		.INIT('hc800)
	) name5079 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_idin_reg[27]/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u2_ep_match_r_reg/P0001 ,
		_w6829_
	);
	LUT2 #(
		.INIT('h1)
	) name5080 (
		_w6828_,
		_w6829_,
		_w6830_
	);
	LUT3 #(
		.INIT('h07)
	) name5081 (
		_w2267_,
		_w2320_,
		_w6830_,
		_w6831_
	);
	LUT3 #(
		.INIT('h2a)
	) name5082 (
		rst_i_pad,
		_w2267_,
		_w6371_,
		_w6832_
	);
	LUT2 #(
		.INIT('hb)
	) name5083 (
		_w6831_,
		_w6832_,
		_w6833_
	);
	LUT4 #(
		.INIT('h10f0)
	) name5084 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u2_buf1_reg[28]/P0001 ,
		\u4_u2_ep_match_r_reg/P0001 ,
		_w6834_
	);
	LUT4 #(
		.INIT('hc800)
	) name5085 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_idin_reg[28]/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u2_ep_match_r_reg/P0001 ,
		_w6835_
	);
	LUT2 #(
		.INIT('h1)
	) name5086 (
		_w6834_,
		_w6835_,
		_w6836_
	);
	LUT3 #(
		.INIT('h07)
	) name5087 (
		_w2267_,
		_w2320_,
		_w6836_,
		_w6837_
	);
	LUT3 #(
		.INIT('h2a)
	) name5088 (
		rst_i_pad,
		_w2267_,
		_w6378_,
		_w6838_
	);
	LUT2 #(
		.INIT('hb)
	) name5089 (
		_w6837_,
		_w6838_,
		_w6839_
	);
	LUT4 #(
		.INIT('h10f0)
	) name5090 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u2_buf1_reg[29]/P0001 ,
		\u4_u2_ep_match_r_reg/P0001 ,
		_w6840_
	);
	LUT4 #(
		.INIT('hc800)
	) name5091 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_idin_reg[29]/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u2_ep_match_r_reg/P0001 ,
		_w6841_
	);
	LUT2 #(
		.INIT('h1)
	) name5092 (
		_w6840_,
		_w6841_,
		_w6842_
	);
	LUT3 #(
		.INIT('h07)
	) name5093 (
		_w2267_,
		_w2320_,
		_w6842_,
		_w6843_
	);
	LUT3 #(
		.INIT('h2a)
	) name5094 (
		rst_i_pad,
		_w2267_,
		_w6385_,
		_w6844_
	);
	LUT2 #(
		.INIT('hb)
	) name5095 (
		_w6843_,
		_w6844_,
		_w6845_
	);
	LUT4 #(
		.INIT('h10f0)
	) name5096 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u2_buf1_reg[2]/P0001 ,
		\u4_u2_ep_match_r_reg/P0001 ,
		_w6846_
	);
	LUT4 #(
		.INIT('hc800)
	) name5097 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_idin_reg[2]/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u2_ep_match_r_reg/P0001 ,
		_w6847_
	);
	LUT2 #(
		.INIT('h1)
	) name5098 (
		_w6846_,
		_w6847_,
		_w6848_
	);
	LUT3 #(
		.INIT('h07)
	) name5099 (
		_w2267_,
		_w2320_,
		_w6848_,
		_w6849_
	);
	LUT3 #(
		.INIT('h2a)
	) name5100 (
		rst_i_pad,
		_w2267_,
		_w6392_,
		_w6850_
	);
	LUT2 #(
		.INIT('hb)
	) name5101 (
		_w6849_,
		_w6850_,
		_w6851_
	);
	LUT4 #(
		.INIT('h10f0)
	) name5102 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u2_buf1_reg[30]/P0001 ,
		\u4_u2_ep_match_r_reg/P0001 ,
		_w6852_
	);
	LUT4 #(
		.INIT('hc800)
	) name5103 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_idin_reg[30]/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u2_ep_match_r_reg/P0001 ,
		_w6853_
	);
	LUT2 #(
		.INIT('h1)
	) name5104 (
		_w6852_,
		_w6853_,
		_w6854_
	);
	LUT3 #(
		.INIT('h07)
	) name5105 (
		_w2267_,
		_w2320_,
		_w6854_,
		_w6855_
	);
	LUT3 #(
		.INIT('h2a)
	) name5106 (
		rst_i_pad,
		_w2267_,
		_w6399_,
		_w6856_
	);
	LUT2 #(
		.INIT('hb)
	) name5107 (
		_w6855_,
		_w6856_,
		_w6857_
	);
	LUT4 #(
		.INIT('h10f0)
	) name5108 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u2_buf1_reg[31]/P0001 ,
		\u4_u2_ep_match_r_reg/P0001 ,
		_w6858_
	);
	LUT4 #(
		.INIT('hc800)
	) name5109 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_idin_reg[31]/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u2_ep_match_r_reg/P0001 ,
		_w6859_
	);
	LUT2 #(
		.INIT('h1)
	) name5110 (
		_w6858_,
		_w6859_,
		_w6860_
	);
	LUT3 #(
		.INIT('h07)
	) name5111 (
		_w2267_,
		_w2320_,
		_w6860_,
		_w6861_
	);
	LUT3 #(
		.INIT('h2a)
	) name5112 (
		rst_i_pad,
		_w2267_,
		_w6406_,
		_w6862_
	);
	LUT2 #(
		.INIT('hb)
	) name5113 (
		_w6861_,
		_w6862_,
		_w6863_
	);
	LUT4 #(
		.INIT('h10f0)
	) name5114 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u2_buf1_reg[3]/P0001 ,
		\u4_u2_ep_match_r_reg/P0001 ,
		_w6864_
	);
	LUT4 #(
		.INIT('hc800)
	) name5115 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_idin_reg[3]/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u2_ep_match_r_reg/P0001 ,
		_w6865_
	);
	LUT2 #(
		.INIT('h1)
	) name5116 (
		_w6864_,
		_w6865_,
		_w6866_
	);
	LUT3 #(
		.INIT('h07)
	) name5117 (
		_w2267_,
		_w2320_,
		_w6866_,
		_w6867_
	);
	LUT3 #(
		.INIT('h2a)
	) name5118 (
		rst_i_pad,
		_w2267_,
		_w6413_,
		_w6868_
	);
	LUT2 #(
		.INIT('hb)
	) name5119 (
		_w6867_,
		_w6868_,
		_w6869_
	);
	LUT4 #(
		.INIT('h10f0)
	) name5120 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u2_buf1_reg[8]/P0001 ,
		\u4_u2_ep_match_r_reg/P0001 ,
		_w6870_
	);
	LUT4 #(
		.INIT('hc800)
	) name5121 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_idin_reg[8]/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u2_ep_match_r_reg/P0001 ,
		_w6871_
	);
	LUT2 #(
		.INIT('h1)
	) name5122 (
		_w6870_,
		_w6871_,
		_w6872_
	);
	LUT3 #(
		.INIT('h07)
	) name5123 (
		_w2267_,
		_w2320_,
		_w6872_,
		_w6873_
	);
	LUT3 #(
		.INIT('h2a)
	) name5124 (
		rst_i_pad,
		_w2267_,
		_w6420_,
		_w6874_
	);
	LUT2 #(
		.INIT('hb)
	) name5125 (
		_w6873_,
		_w6874_,
		_w6875_
	);
	LUT4 #(
		.INIT('h10f0)
	) name5126 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u2_buf1_reg[9]/P0001 ,
		\u4_u2_ep_match_r_reg/P0001 ,
		_w6876_
	);
	LUT4 #(
		.INIT('hc800)
	) name5127 (
		\u1_u3_buf1_set_reg/P0001 ,
		\u1_u3_idin_reg[9]/P0001 ,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u2_ep_match_r_reg/P0001 ,
		_w6877_
	);
	LUT2 #(
		.INIT('h1)
	) name5128 (
		_w6876_,
		_w6877_,
		_w6878_
	);
	LUT3 #(
		.INIT('h07)
	) name5129 (
		_w2267_,
		_w2320_,
		_w6878_,
		_w6879_
	);
	LUT3 #(
		.INIT('h2a)
	) name5130 (
		rst_i_pad,
		_w2267_,
		_w6427_,
		_w6880_
	);
	LUT2 #(
		.INIT('hb)
	) name5131 (
		_w6879_,
		_w6880_,
		_w6881_
	);
	LUT4 #(
		.INIT('h0008)
	) name5132 (
		\u0_rx_active_reg/P0001 ,
		\u0_rx_valid_reg/P0001 ,
		\u1_u0_state_reg[1]/P0001 ,
		\u1_u0_state_reg[3]/P0001 ,
		_w6882_
	);
	LUT3 #(
		.INIT('h08)
	) name5133 (
		rst_i_pad,
		\u1_u0_state_reg[0]/P0001 ,
		\u1_u0_state_reg[2]/P0001 ,
		_w6883_
	);
	LUT2 #(
		.INIT('h8)
	) name5134 (
		_w6882_,
		_w6883_,
		_w6884_
	);
	LUT3 #(
		.INIT('h04)
	) name5135 (
		_w3695_,
		_w4884_,
		_w4885_,
		_w6885_
	);
	LUT4 #(
		.INIT('h1000)
	) name5136 (
		\u0_rx_err_reg/P0001 ,
		_w3695_,
		_w4883_,
		_w5245_,
		_w6886_
	);
	LUT3 #(
		.INIT('h80)
	) name5137 (
		rst_i_pad,
		\u0_rx_active_reg/P0001 ,
		\u1_u0_state_reg[1]/P0001 ,
		_w6887_
	);
	LUT2 #(
		.INIT('h8)
	) name5138 (
		_w4881_,
		_w6887_,
		_w6888_
	);
	LUT4 #(
		.INIT('habaa)
	) name5139 (
		_w6884_,
		_w6885_,
		_w6886_,
		_w6888_,
		_w6889_
	);
	LUT2 #(
		.INIT('h9)
	) name5140 (
		\u0_rx_data_reg[6]/P0001 ,
		\u0_rx_data_reg[7]/P0001 ,
		_w6890_
	);
	LUT3 #(
		.INIT('h96)
	) name5141 (
		\u0_rx_data_reg[6]/P0001 ,
		\u0_rx_data_reg[7]/P0001 ,
		\u1_u0_crc16_sum_reg[8]/P0001 ,
		_w6891_
	);
	LUT2 #(
		.INIT('h9)
	) name5142 (
		\u0_rx_data_reg[0]/P0001 ,
		\u0_rx_data_reg[1]/P0001 ,
		_w6892_
	);
	LUT4 #(
		.INIT('h6996)
	) name5143 (
		\u0_rx_data_reg[0]/P0001 ,
		\u0_rx_data_reg[1]/P0001 ,
		\u0_rx_data_reg[2]/P0001 ,
		\u0_rx_data_reg[3]/P0001 ,
		_w6893_
	);
	LUT2 #(
		.INIT('h9)
	) name5144 (
		\u0_rx_data_reg[4]/P0001 ,
		\u0_rx_data_reg[5]/P0001 ,
		_w6894_
	);
	LUT2 #(
		.INIT('h6)
	) name5145 (
		\u1_u0_crc16_sum_reg[15]/P0001 ,
		\u1_u0_crc16_sum_reg[7]/P0001 ,
		_w6895_
	);
	LUT4 #(
		.INIT('h9669)
	) name5146 (
		_w6891_,
		_w6893_,
		_w6894_,
		_w6895_,
		_w6896_
	);
	LUT2 #(
		.INIT('h8)
	) name5147 (
		_w3671_,
		_w4884_,
		_w6897_
	);
	LUT4 #(
		.INIT('hb000)
	) name5148 (
		\u0_rx_err_reg/P0001 ,
		_w3695_,
		_w4881_,
		_w5245_,
		_w6898_
	);
	LUT2 #(
		.INIT('h8)
	) name5149 (
		_w4884_,
		_w4885_,
		_w6899_
	);
	LUT3 #(
		.INIT('h15)
	) name5150 (
		_w6897_,
		_w6898_,
		_w6899_,
		_w6900_
	);
	LUT3 #(
		.INIT('hea)
	) name5151 (
		_w6897_,
		_w6898_,
		_w6899_,
		_w6901_
	);
	LUT2 #(
		.INIT('h9)
	) name5152 (
		\u1_u0_crc16_sum_reg[11]/P0001 ,
		\u1_u0_crc16_sum_reg[12]/P0001 ,
		_w6902_
	);
	LUT4 #(
		.INIT('h6996)
	) name5153 (
		\u1_u0_crc16_sum_reg[10]/P0001 ,
		\u1_u0_crc16_sum_reg[13]/P0001 ,
		\u1_u0_crc16_sum_reg[14]/P0001 ,
		\u1_u0_crc16_sum_reg[9]/P0001 ,
		_w6903_
	);
	LUT2 #(
		.INIT('h6)
	) name5154 (
		_w6902_,
		_w6903_,
		_w6904_
	);
	LUT4 #(
		.INIT('h00ea)
	) name5155 (
		_w6897_,
		_w6898_,
		_w6899_,
		_w6904_,
		_w6905_
	);
	LUT2 #(
		.INIT('h4)
	) name5156 (
		_w6896_,
		_w6905_,
		_w6906_
	);
	LUT4 #(
		.INIT('hea00)
	) name5157 (
		_w6897_,
		_w6898_,
		_w6899_,
		_w6904_,
		_w6907_
	);
	LUT2 #(
		.INIT('h6)
	) name5158 (
		_w6893_,
		_w6894_,
		_w6908_
	);
	LUT3 #(
		.INIT('h69)
	) name5159 (
		\u1_u0_crc16_sum_reg[15]/P0001 ,
		\u1_u0_crc16_sum_reg[7]/P0001 ,
		\u1_u0_crc16_sum_reg[8]/P0001 ,
		_w6909_
	);
	LUT4 #(
		.INIT('h9669)
	) name5160 (
		_w6890_,
		_w6893_,
		_w6894_,
		_w6909_,
		_w6910_
	);
	LUT2 #(
		.INIT('h2)
	) name5161 (
		\u0_rx_active_reg/P0001 ,
		\u1_u0_rx_active_r_reg/P0001 ,
		_w6911_
	);
	LUT4 #(
		.INIT('hdf00)
	) name5162 (
		\u0_rx_active_reg/P0001 ,
		\u0_rx_err_reg/P0001 ,
		\u0_rx_valid_reg/P0001 ,
		\u1_u0_crc16_sum_reg[15]/P0001 ,
		_w6912_
	);
	LUT2 #(
		.INIT('h2)
	) name5163 (
		\u1_u0_crc16_sum_reg[15]/P0001 ,
		_w3671_,
		_w6913_
	);
	LUT4 #(
		.INIT('h040f)
	) name5164 (
		_w4886_,
		_w6898_,
		_w6912_,
		_w6913_,
		_w6914_
	);
	LUT4 #(
		.INIT('h0700)
	) name5165 (
		_w6907_,
		_w6910_,
		_w6911_,
		_w6914_,
		_w6915_
	);
	LUT2 #(
		.INIT('hb)
	) name5166 (
		_w6906_,
		_w6915_,
		_w6916_
	);
	LUT2 #(
		.INIT('h6)
	) name5167 (
		\u1_u0_crc16_sum_reg[12]/P0001 ,
		\u1_u0_crc16_sum_reg[13]/P0001 ,
		_w6917_
	);
	LUT2 #(
		.INIT('h9)
	) name5168 (
		\u1_u0_crc16_sum_reg[14]/P0001 ,
		\u1_u0_crc16_sum_reg[15]/P0001 ,
		_w6918_
	);
	LUT4 #(
		.INIT('h6996)
	) name5169 (
		\u1_u0_crc16_sum_reg[9]/P0001 ,
		_w6893_,
		_w6917_,
		_w6918_,
		_w6919_
	);
	LUT2 #(
		.INIT('h6)
	) name5170 (
		\u1_u0_crc16_sum_reg[10]/P0001 ,
		\u1_u0_crc16_sum_reg[11]/P0001 ,
		_w6920_
	);
	LUT4 #(
		.INIT('h9669)
	) name5171 (
		\u0_rx_data_reg[4]/P0001 ,
		\u0_rx_data_reg[5]/P0001 ,
		\u1_u0_crc16_sum_reg[10]/P0001 ,
		\u1_u0_crc16_sum_reg[11]/P0001 ,
		_w6921_
	);
	LUT2 #(
		.INIT('h6)
	) name5172 (
		\u0_rx_data_reg[6]/P0001 ,
		_w6921_,
		_w6922_
	);
	LUT4 #(
		.INIT('h9669)
	) name5173 (
		\u1_u0_crc16_sum_reg[12]/P0001 ,
		\u1_u0_crc16_sum_reg[13]/P0001 ,
		\u1_u0_crc16_sum_reg[14]/P0001 ,
		\u1_u0_crc16_sum_reg[15]/P0001 ,
		_w6923_
	);
	LUT3 #(
		.INIT('h96)
	) name5174 (
		\u1_u0_crc16_sum_reg[9]/P0001 ,
		_w6893_,
		_w6923_,
		_w6924_
	);
	LUT4 #(
		.INIT('heaef)
	) name5175 (
		_w6900_,
		_w6919_,
		_w6922_,
		_w6924_,
		_w6925_
	);
	LUT2 #(
		.INIT('h2)
	) name5176 (
		\u1_u0_crc16_sum_reg[1]/P0001 ,
		_w3671_,
		_w6926_
	);
	LUT4 #(
		.INIT('hdf00)
	) name5177 (
		\u0_rx_active_reg/P0001 ,
		\u0_rx_err_reg/P0001 ,
		\u0_rx_valid_reg/P0001 ,
		\u1_u0_crc16_sum_reg[1]/P0001 ,
		_w6927_
	);
	LUT2 #(
		.INIT('h1)
	) name5178 (
		_w6911_,
		_w6927_,
		_w6928_
	);
	LUT4 #(
		.INIT('h4f00)
	) name5179 (
		_w4886_,
		_w6898_,
		_w6926_,
		_w6928_,
		_w6929_
	);
	LUT2 #(
		.INIT('h7)
	) name5180 (
		_w6925_,
		_w6929_,
		_w6930_
	);
	LUT2 #(
		.INIT('h2)
	) name5181 (
		\u0_rx_active_reg/P0001 ,
		\u1_u0_state_reg[0]/P0001 ,
		_w6931_
	);
	LUT2 #(
		.INIT('h2)
	) name5182 (
		_w4881_,
		_w6931_,
		_w6932_
	);
	LUT3 #(
		.INIT('h10)
	) name5183 (
		_w6885_,
		_w6886_,
		_w6932_,
		_w6933_
	);
	LUT2 #(
		.INIT('h2)
	) name5184 (
		_w3671_,
		_w6931_,
		_w6934_
	);
	LUT2 #(
		.INIT('h8)
	) name5185 (
		_w4884_,
		_w4888_,
		_w6935_
	);
	LUT3 #(
		.INIT('h2a)
	) name5186 (
		rst_i_pad,
		_w4884_,
		_w4888_,
		_w6936_
	);
	LUT4 #(
		.INIT('h0013)
	) name5187 (
		\u1_u0_state_reg[0]/P0001 ,
		\u1_u0_state_reg[1]/P0001 ,
		\u1_u0_state_reg[2]/P0001 ,
		\u1_u0_state_reg[3]/P0001 ,
		_w6937_
	);
	LUT3 #(
		.INIT('hdc)
	) name5188 (
		\u0_rx_active_reg/P0001 ,
		\u1_u0_state_reg[0]/P0001 ,
		\u1_u0_state_reg[2]/P0001 ,
		_w6938_
	);
	LUT3 #(
		.INIT('h40)
	) name5189 (
		_w4883_,
		_w6937_,
		_w6938_,
		_w6939_
	);
	LUT3 #(
		.INIT('h04)
	) name5190 (
		_w6934_,
		_w6936_,
		_w6939_,
		_w6940_
	);
	LUT2 #(
		.INIT('hb)
	) name5191 (
		_w6933_,
		_w6940_,
		_w6941_
	);
	LUT4 #(
		.INIT('h0440)
	) name5192 (
		\u1_u2_word_done_r_reg/P0001 ,
		\u2_wack_r_reg/P0001 ,
		\u5_state_reg[1]/P0001 ,
		\u5_state_reg[2]/P0001 ,
		_w6942_
	);
	LUT4 #(
		.INIT('hae00)
	) name5193 (
		\u1_u2_mack_r_reg/P0001 ,
		_w3224_,
		_w5488_,
		_w6942_,
		_w6943_
	);
	LUT2 #(
		.INIT('he)
	) name5194 (
		_w5674_,
		_w6943_,
		_w6944_
	);
	LUT3 #(
		.INIT('ha6)
	) name5195 (
		\u1_u3_new_sizeb_reg[2]/P0001 ,
		_w2795_,
		_w2797_,
		_w6945_
	);
	LUT4 #(
		.INIT('he817)
	) name5196 (
		\u1_u3_new_sizeb_reg[1]/P0001 ,
		_w2785_,
		_w3440_,
		_w6945_,
		_w6946_
	);
	LUT4 #(
		.INIT('h0e08)
	) name5197 (
		\u1_u3_new_sizeb_reg[1]/P0001 ,
		_w2785_,
		_w3438_,
		_w3440_,
		_w6947_
	);
	LUT3 #(
		.INIT('ha6)
	) name5198 (
		\u1_u3_new_sizeb_reg[3]/P0001 ,
		_w2810_,
		_w2812_,
		_w6948_
	);
	LUT3 #(
		.INIT('he1)
	) name5199 (
		_w3442_,
		_w6947_,
		_w6948_,
		_w6949_
	);
	LUT4 #(
		.INIT('h135f)
	) name5200 (
		\u4_int_srcb_reg[4]/P0001 ,
		\u4_int_srcb_reg[6]/P0001 ,
		\u4_inta_msk_reg[4]/P0001 ,
		\u4_inta_msk_reg[6]/P0001 ,
		_w6950_
	);
	LUT4 #(
		.INIT('h135f)
	) name5201 (
		\u4_int_srcb_reg[5]/P0001 ,
		\u4_int_srcb_reg[7]/P0001 ,
		\u4_inta_msk_reg[5]/P0001 ,
		\u4_inta_msk_reg[7]/P0001 ,
		_w6951_
	);
	LUT4 #(
		.INIT('h0001)
	) name5202 (
		\u4_u0_inta_reg/P0001 ,
		\u4_u1_inta_reg/P0001 ,
		\u4_u2_inta_reg/P0001 ,
		\u4_u3_inta_reg/P0001 ,
		_w6952_
	);
	LUT4 #(
		.INIT('h135f)
	) name5203 (
		\u4_int_srcb_reg[0]/P0001 ,
		\u4_int_srcb_reg[3]/P0001 ,
		\u4_inta_msk_reg[0]/P0001 ,
		\u4_inta_msk_reg[3]/P0001 ,
		_w6953_
	);
	LUT4 #(
		.INIT('h8000)
	) name5204 (
		_w6950_,
		_w6951_,
		_w6952_,
		_w6953_,
		_w6954_
	);
	LUT4 #(
		.INIT('h135f)
	) name5205 (
		\u4_int_srcb_reg[2]/P0001 ,
		\u4_int_srcb_reg[8]/P0001 ,
		\u4_inta_msk_reg[2]/P0001 ,
		\u4_inta_msk_reg[8]/P0001 ,
		_w6955_
	);
	LUT2 #(
		.INIT('h8)
	) name5206 (
		\u4_int_srcb_reg[1]/P0001 ,
		\u4_inta_msk_reg[1]/P0001 ,
		_w6956_
	);
	LUT2 #(
		.INIT('h2)
	) name5207 (
		_w6955_,
		_w6956_,
		_w6957_
	);
	LUT2 #(
		.INIT('h7)
	) name5208 (
		_w6954_,
		_w6957_,
		_w6958_
	);
	LUT4 #(
		.INIT('h135f)
	) name5209 (
		\u4_int_srcb_reg[4]/P0001 ,
		\u4_int_srcb_reg[6]/P0001 ,
		\u4_intb_msk_reg[4]/P0001 ,
		\u4_intb_msk_reg[6]/P0001 ,
		_w6959_
	);
	LUT4 #(
		.INIT('h135f)
	) name5210 (
		\u4_int_srcb_reg[5]/P0001 ,
		\u4_int_srcb_reg[7]/P0001 ,
		\u4_intb_msk_reg[5]/P0001 ,
		\u4_intb_msk_reg[7]/P0001 ,
		_w6960_
	);
	LUT4 #(
		.INIT('h0001)
	) name5211 (
		\u4_u0_intb_reg/P0001 ,
		\u4_u1_intb_reg/P0001 ,
		\u4_u2_intb_reg/P0001 ,
		\u4_u3_intb_reg/P0001 ,
		_w6961_
	);
	LUT4 #(
		.INIT('h135f)
	) name5212 (
		\u4_int_srcb_reg[0]/P0001 ,
		\u4_int_srcb_reg[3]/P0001 ,
		\u4_intb_msk_reg[0]/P0001 ,
		\u4_intb_msk_reg[3]/P0001 ,
		_w6962_
	);
	LUT4 #(
		.INIT('h8000)
	) name5213 (
		_w6959_,
		_w6960_,
		_w6961_,
		_w6962_,
		_w6963_
	);
	LUT4 #(
		.INIT('h135f)
	) name5214 (
		\u4_int_srcb_reg[2]/P0001 ,
		\u4_int_srcb_reg[8]/P0001 ,
		\u4_intb_msk_reg[2]/P0001 ,
		\u4_intb_msk_reg[8]/P0001 ,
		_w6964_
	);
	LUT2 #(
		.INIT('h8)
	) name5215 (
		\u4_int_srcb_reg[1]/P0001 ,
		\u4_intb_msk_reg[1]/P0001 ,
		_w6965_
	);
	LUT2 #(
		.INIT('h2)
	) name5216 (
		_w6964_,
		_w6965_,
		_w6966_
	);
	LUT2 #(
		.INIT('h7)
	) name5217 (
		_w6963_,
		_w6966_,
		_w6967_
	);
	LUT4 #(
		.INIT('h0001)
	) name5218 (
		\u1_u3_buf0_rl_reg/P0001 ,
		\u1_u3_buf0_set_reg/P0001 ,
		\u4_u3_r5_reg/NET0131 ,
		\u4_u3_set_r_reg/P0001 ,
		_w6968_
	);
	LUT3 #(
		.INIT('h07)
	) name5219 (
		\u4_u3_csr0_reg[2]/P0001 ,
		\u4_u3_ep_match_r_reg/P0001 ,
		\u4_u3_r5_reg/NET0131 ,
		_w6969_
	);
	LUT4 #(
		.INIT('h8882)
	) name5220 (
		\u4_u3_csr1_reg[0]/P0001 ,
		\u4_u3_dma_in_cnt_reg[0]/P0001 ,
		_w6968_,
		_w6969_,
		_w6970_
	);
	LUT3 #(
		.INIT('h07)
	) name5221 (
		\u4_u0_csr0_reg[2]/P0001 ,
		\u4_u0_ep_match_r_reg/P0001 ,
		\u4_u0_r5_reg/NET0131 ,
		_w6971_
	);
	LUT4 #(
		.INIT('h8882)
	) name5222 (
		\u4_u0_csr1_reg[0]/P0001 ,
		\u4_u0_dma_in_cnt_reg[0]/P0001 ,
		_w6971_,
		_w5003_,
		_w6972_
	);
	LUT3 #(
		.INIT('h07)
	) name5223 (
		\u4_u1_csr0_reg[2]/P0001 ,
		\u4_u1_ep_match_r_reg/P0001 ,
		\u4_u1_r5_reg/NET0131 ,
		_w6973_
	);
	LUT4 #(
		.INIT('h8882)
	) name5224 (
		\u4_u1_csr1_reg[0]/P0001 ,
		\u4_u1_dma_in_cnt_reg[0]/P0001 ,
		_w6973_,
		_w5037_,
		_w6974_
	);
	LUT3 #(
		.INIT('h07)
	) name5225 (
		\u4_u2_csr0_reg[2]/P0001 ,
		\u4_u2_ep_match_r_reg/P0001 ,
		\u4_u2_r5_reg/NET0131 ,
		_w6975_
	);
	LUT4 #(
		.INIT('h0001)
	) name5226 (
		\u1_u3_buf0_rl_reg/P0001 ,
		\u1_u3_buf0_set_reg/P0001 ,
		\u4_u2_r5_reg/NET0131 ,
		\u4_u2_set_r_reg/P0001 ,
		_w6976_
	);
	LUT4 #(
		.INIT('h8882)
	) name5227 (
		\u4_u2_csr1_reg[0]/P0001 ,
		\u4_u2_dma_in_cnt_reg[0]/P0001 ,
		_w6975_,
		_w6976_,
		_w6977_
	);
	LUT2 #(
		.INIT('h6)
	) name5228 (
		\u4_u3_csr0_reg[3]/NET0131 ,
		\u4_u3_dma_out_cnt_reg[1]/P0001 ,
		_w6978_
	);
	LUT3 #(
		.INIT('h90)
	) name5229 (
		\u4_u3_dma_in_cnt_reg[0]/P0001 ,
		\u4_u3_dma_out_cnt_reg[1]/P0001 ,
		\u4_u3_r5_reg/NET0131 ,
		_w6979_
	);
	LUT4 #(
		.INIT('h0082)
	) name5230 (
		_w4569_,
		_w4668_,
		_w6978_,
		_w6979_,
		_w6980_
	);
	LUT4 #(
		.INIT('h0001)
	) name5231 (
		\u1_u3_buf0_rl_reg/P0001 ,
		\u1_u3_buf0_set_reg/P0001 ,
		\u4_u3_dma_out_cnt_reg[1]/P0001 ,
		\u4_u3_set_r_reg/P0001 ,
		_w6981_
	);
	LUT3 #(
		.INIT('h0e)
	) name5232 (
		\u4_u3_dma_out_cnt_reg[1]/P0001 ,
		\u4_u3_ep_match_r_reg/P0001 ,
		\u4_u3_r5_reg/NET0131 ,
		_w6982_
	);
	LUT4 #(
		.INIT('h8a88)
	) name5233 (
		\u4_u3_csr1_reg[0]/P0001 ,
		_w6979_,
		_w6981_,
		_w6982_,
		_w6983_
	);
	LUT2 #(
		.INIT('h4)
	) name5234 (
		_w6980_,
		_w6983_,
		_w6984_
	);
	LUT4 #(
		.INIT('hec80)
	) name5235 (
		\u4_u3_csr0_reg[2]/P0001 ,
		\u4_u3_csr0_reg[3]/NET0131 ,
		\u4_u3_dma_in_cnt_reg[0]/P0001 ,
		\u4_u3_dma_out_cnt_reg[1]/P0001 ,
		_w6985_
	);
	LUT2 #(
		.INIT('h6)
	) name5236 (
		\u4_u3_csr0_reg[4]/P0001 ,
		\u4_u3_dma_out_cnt_reg[2]/P0001 ,
		_w6986_
	);
	LUT4 #(
		.INIT('h1eff)
	) name5237 (
		\u4_u3_dma_in_cnt_reg[0]/P0001 ,
		\u4_u3_dma_out_cnt_reg[1]/P0001 ,
		\u4_u3_dma_out_cnt_reg[2]/P0001 ,
		\u4_u3_r5_reg/NET0131 ,
		_w6987_
	);
	LUT4 #(
		.INIT('h8200)
	) name5238 (
		_w4569_,
		_w6985_,
		_w6986_,
		_w6987_,
		_w6988_
	);
	LUT4 #(
		.INIT('h0001)
	) name5239 (
		\u1_u3_buf0_rl_reg/P0001 ,
		\u1_u3_buf0_set_reg/P0001 ,
		\u4_u3_dma_out_cnt_reg[2]/P0001 ,
		\u4_u3_set_r_reg/P0001 ,
		_w6989_
	);
	LUT3 #(
		.INIT('h0e)
	) name5240 (
		\u4_u3_dma_out_cnt_reg[2]/P0001 ,
		\u4_u3_ep_match_r_reg/P0001 ,
		\u4_u3_r5_reg/NET0131 ,
		_w6990_
	);
	LUT4 #(
		.INIT('h2a22)
	) name5241 (
		\u4_u3_csr1_reg[0]/P0001 ,
		_w6987_,
		_w6989_,
		_w6990_,
		_w6991_
	);
	LUT2 #(
		.INIT('h4)
	) name5242 (
		_w6988_,
		_w6991_,
		_w6992_
	);
	LUT4 #(
		.INIT('h6f3f)
	) name5243 (
		\u4_u3_dma_out_cnt_reg[2]/P0001 ,
		\u4_u3_dma_out_cnt_reg[3]/P0001 ,
		\u4_u3_r5_reg/NET0131 ,
		_w4651_,
		_w6993_
	);
	LUT2 #(
		.INIT('h2)
	) name5244 (
		\u4_u3_csr1_reg[0]/P0001 ,
		_w6993_,
		_w6994_
	);
	LUT2 #(
		.INIT('h6)
	) name5245 (
		\u4_u3_csr0_reg[5]/P0001 ,
		\u4_u3_dma_out_cnt_reg[3]/P0001 ,
		_w6995_
	);
	LUT4 #(
		.INIT('h00f4)
	) name5246 (
		_w4669_,
		_w4670_,
		_w4671_,
		_w6995_,
		_w6996_
	);
	LUT4 #(
		.INIT('h134c)
	) name5247 (
		\u4_u3_csr0_reg[4]/P0001 ,
		\u4_u3_csr0_reg[5]/P0001 ,
		\u4_u3_dma_out_cnt_reg[2]/P0001 ,
		\u4_u3_dma_out_cnt_reg[3]/P0001 ,
		_w6997_
	);
	LUT4 #(
		.INIT('h20aa)
	) name5248 (
		_w4569_,
		_w4669_,
		_w4670_,
		_w6997_,
		_w6998_
	);
	LUT4 #(
		.INIT('h0001)
	) name5249 (
		\u1_u3_buf0_rl_reg/P0001 ,
		\u1_u3_buf0_set_reg/P0001 ,
		\u4_u3_dma_out_cnt_reg[3]/P0001 ,
		\u4_u3_set_r_reg/P0001 ,
		_w6999_
	);
	LUT3 #(
		.INIT('ha8)
	) name5250 (
		\u4_u3_csr1_reg[0]/P0001 ,
		\u4_u3_dma_out_cnt_reg[3]/P0001 ,
		\u4_u3_ep_match_r_reg/P0001 ,
		_w7000_
	);
	LUT3 #(
		.INIT('h10)
	) name5251 (
		\u4_u3_r5_reg/NET0131 ,
		_w6999_,
		_w7000_,
		_w7001_
	);
	LUT3 #(
		.INIT('hb0)
	) name5252 (
		_w6996_,
		_w6998_,
		_w7001_,
		_w7002_
	);
	LUT2 #(
		.INIT('he)
	) name5253 (
		_w6994_,
		_w7002_,
		_w7003_
	);
	LUT4 #(
		.INIT('h4000)
	) name5254 (
		\u1_u2_mack_r_reg/P0001 ,
		\u1_u2_state_reg[4]/NET0131 ,
		_w3205_,
		_w3206_,
		_w7004_
	);
	LUT3 #(
		.INIT('h04)
	) name5255 (
		\u1_u2_mack_r_reg/P0001 ,
		\u1_u2_state_reg[4]/NET0131 ,
		\u1_u3_abort_reg/P0001 ,
		_w7005_
	);
	LUT4 #(
		.INIT('ha800)
	) name5256 (
		_w3205_,
		_w3222_,
		_w3223_,
		_w7005_,
		_w7006_
	);
	LUT4 #(
		.INIT('h00f2)
	) name5257 (
		\u1_u2_state_reg[4]/NET0131 ,
		\u1_u2_wr_done_reg/P0001 ,
		\u1_u2_wr_last_reg/P0001 ,
		\u1_u3_abort_reg/P0001 ,
		_w7007_
	);
	LUT3 #(
		.INIT('h80)
	) name5258 (
		_w3209_,
		_w3214_,
		_w7007_,
		_w7008_
	);
	LUT4 #(
		.INIT('haaa8)
	) name5259 (
		rst_i_pad,
		_w7004_,
		_w7006_,
		_w7008_,
		_w7009_
	);
	LUT2 #(
		.INIT('h6)
	) name5260 (
		\u4_u0_csr0_reg[3]/NET0131 ,
		\u4_u0_dma_out_cnt_reg[1]/P0001 ,
		_w7010_
	);
	LUT3 #(
		.INIT('h90)
	) name5261 (
		\u4_u0_dma_in_cnt_reg[0]/P0001 ,
		\u4_u0_dma_out_cnt_reg[1]/P0001 ,
		\u4_u0_r5_reg/NET0131 ,
		_w7011_
	);
	LUT4 #(
		.INIT('h0082)
	) name5262 (
		_w4592_,
		_w4698_,
		_w7010_,
		_w7011_,
		_w7012_
	);
	LUT4 #(
		.INIT('h0001)
	) name5263 (
		\u1_u3_buf0_rl_reg/P0001 ,
		\u1_u3_buf0_set_reg/P0001 ,
		\u4_u0_dma_out_cnt_reg[1]/P0001 ,
		\u4_u0_set_r_reg/P0001 ,
		_w7013_
	);
	LUT3 #(
		.INIT('h0e)
	) name5264 (
		\u4_u0_dma_out_cnt_reg[1]/P0001 ,
		\u4_u0_ep_match_r_reg/P0001 ,
		\u4_u0_r5_reg/NET0131 ,
		_w7014_
	);
	LUT4 #(
		.INIT('h8a88)
	) name5265 (
		\u4_u0_csr1_reg[0]/P0001 ,
		_w7011_,
		_w7013_,
		_w7014_,
		_w7015_
	);
	LUT2 #(
		.INIT('h4)
	) name5266 (
		_w7012_,
		_w7015_,
		_w7016_
	);
	LUT4 #(
		.INIT('hec80)
	) name5267 (
		\u4_u0_csr0_reg[2]/P0001 ,
		\u4_u0_csr0_reg[3]/NET0131 ,
		\u4_u0_dma_in_cnt_reg[0]/P0001 ,
		\u4_u0_dma_out_cnt_reg[1]/P0001 ,
		_w7017_
	);
	LUT2 #(
		.INIT('h6)
	) name5268 (
		\u4_u0_csr0_reg[4]/P0001 ,
		\u4_u0_dma_out_cnt_reg[2]/P0001 ,
		_w7018_
	);
	LUT4 #(
		.INIT('h1eff)
	) name5269 (
		\u4_u0_dma_in_cnt_reg[0]/P0001 ,
		\u4_u0_dma_out_cnt_reg[1]/P0001 ,
		\u4_u0_dma_out_cnt_reg[2]/P0001 ,
		\u4_u0_r5_reg/NET0131 ,
		_w7019_
	);
	LUT4 #(
		.INIT('h8200)
	) name5270 (
		_w4592_,
		_w7017_,
		_w7018_,
		_w7019_,
		_w7020_
	);
	LUT4 #(
		.INIT('h0001)
	) name5271 (
		\u1_u3_buf0_rl_reg/P0001 ,
		\u1_u3_buf0_set_reg/P0001 ,
		\u4_u0_dma_out_cnt_reg[2]/P0001 ,
		\u4_u0_set_r_reg/P0001 ,
		_w7021_
	);
	LUT3 #(
		.INIT('h0e)
	) name5272 (
		\u4_u0_dma_out_cnt_reg[2]/P0001 ,
		\u4_u0_ep_match_r_reg/P0001 ,
		\u4_u0_r5_reg/NET0131 ,
		_w7022_
	);
	LUT4 #(
		.INIT('h2a22)
	) name5273 (
		\u4_u0_csr1_reg[0]/P0001 ,
		_w7019_,
		_w7021_,
		_w7022_,
		_w7023_
	);
	LUT2 #(
		.INIT('h4)
	) name5274 (
		_w7020_,
		_w7023_,
		_w7024_
	);
	LUT4 #(
		.INIT('h6f3f)
	) name5275 (
		\u4_u0_dma_out_cnt_reg[2]/P0001 ,
		\u4_u0_dma_out_cnt_reg[3]/P0001 ,
		\u4_u0_r5_reg/NET0131 ,
		_w4682_,
		_w7025_
	);
	LUT2 #(
		.INIT('h2)
	) name5276 (
		\u4_u0_csr1_reg[0]/P0001 ,
		_w7025_,
		_w7026_
	);
	LUT2 #(
		.INIT('h6)
	) name5277 (
		\u4_u0_csr0_reg[5]/P0001 ,
		\u4_u0_dma_out_cnt_reg[3]/P0001 ,
		_w7027_
	);
	LUT4 #(
		.INIT('h00f4)
	) name5278 (
		_w4699_,
		_w4700_,
		_w4701_,
		_w7027_,
		_w7028_
	);
	LUT4 #(
		.INIT('h134c)
	) name5279 (
		\u4_u0_csr0_reg[4]/P0001 ,
		\u4_u0_csr0_reg[5]/P0001 ,
		\u4_u0_dma_out_cnt_reg[2]/P0001 ,
		\u4_u0_dma_out_cnt_reg[3]/P0001 ,
		_w7029_
	);
	LUT4 #(
		.INIT('h20aa)
	) name5280 (
		_w4592_,
		_w4699_,
		_w4700_,
		_w7029_,
		_w7030_
	);
	LUT4 #(
		.INIT('h0001)
	) name5281 (
		\u1_u3_buf0_rl_reg/P0001 ,
		\u1_u3_buf0_set_reg/P0001 ,
		\u4_u0_dma_out_cnt_reg[3]/P0001 ,
		\u4_u0_set_r_reg/P0001 ,
		_w7031_
	);
	LUT3 #(
		.INIT('h0e)
	) name5282 (
		\u4_u0_dma_out_cnt_reg[3]/P0001 ,
		\u4_u0_ep_match_r_reg/P0001 ,
		\u4_u0_r5_reg/NET0131 ,
		_w7032_
	);
	LUT3 #(
		.INIT('h20)
	) name5283 (
		\u4_u0_csr1_reg[0]/P0001 ,
		_w7031_,
		_w7032_,
		_w7033_
	);
	LUT3 #(
		.INIT('hb0)
	) name5284 (
		_w7028_,
		_w7030_,
		_w7033_,
		_w7034_
	);
	LUT2 #(
		.INIT('he)
	) name5285 (
		_w7026_,
		_w7034_,
		_w7035_
	);
	LUT2 #(
		.INIT('h6)
	) name5286 (
		\u4_u1_csr0_reg[3]/NET0131 ,
		\u4_u1_dma_out_cnt_reg[1]/P0001 ,
		_w7036_
	);
	LUT3 #(
		.INIT('h90)
	) name5287 (
		\u4_u1_dma_in_cnt_reg[0]/P0001 ,
		\u4_u1_dma_out_cnt_reg[1]/P0001 ,
		\u4_u1_r5_reg/NET0131 ,
		_w7037_
	);
	LUT4 #(
		.INIT('h0082)
	) name5288 (
		_w4454_,
		_w4729_,
		_w7036_,
		_w7037_,
		_w7038_
	);
	LUT4 #(
		.INIT('h0001)
	) name5289 (
		\u1_u3_buf0_rl_reg/P0001 ,
		\u1_u3_buf0_set_reg/P0001 ,
		\u4_u1_dma_out_cnt_reg[1]/P0001 ,
		\u4_u1_set_r_reg/P0001 ,
		_w7039_
	);
	LUT3 #(
		.INIT('h0e)
	) name5290 (
		\u4_u1_dma_out_cnt_reg[1]/P0001 ,
		\u4_u1_ep_match_r_reg/P0001 ,
		\u4_u1_r5_reg/NET0131 ,
		_w7040_
	);
	LUT4 #(
		.INIT('h8a88)
	) name5291 (
		\u4_u1_csr1_reg[0]/P0001 ,
		_w7037_,
		_w7039_,
		_w7040_,
		_w7041_
	);
	LUT2 #(
		.INIT('h4)
	) name5292 (
		_w7038_,
		_w7041_,
		_w7042_
	);
	LUT4 #(
		.INIT('hec80)
	) name5293 (
		\u4_u1_csr0_reg[2]/P0001 ,
		\u4_u1_csr0_reg[3]/NET0131 ,
		\u4_u1_dma_in_cnt_reg[0]/P0001 ,
		\u4_u1_dma_out_cnt_reg[1]/P0001 ,
		_w7043_
	);
	LUT2 #(
		.INIT('h6)
	) name5294 (
		\u4_u1_csr0_reg[4]/P0001 ,
		\u4_u1_dma_out_cnt_reg[2]/P0001 ,
		_w7044_
	);
	LUT4 #(
		.INIT('h1eff)
	) name5295 (
		\u4_u1_dma_in_cnt_reg[0]/P0001 ,
		\u4_u1_dma_out_cnt_reg[1]/P0001 ,
		\u4_u1_dma_out_cnt_reg[2]/P0001 ,
		\u4_u1_r5_reg/NET0131 ,
		_w7045_
	);
	LUT4 #(
		.INIT('h8200)
	) name5296 (
		_w4454_,
		_w7043_,
		_w7044_,
		_w7045_,
		_w7046_
	);
	LUT4 #(
		.INIT('h0001)
	) name5297 (
		\u1_u3_buf0_rl_reg/P0001 ,
		\u1_u3_buf0_set_reg/P0001 ,
		\u4_u1_dma_out_cnt_reg[2]/P0001 ,
		\u4_u1_set_r_reg/P0001 ,
		_w7047_
	);
	LUT3 #(
		.INIT('h0e)
	) name5298 (
		\u4_u1_dma_out_cnt_reg[2]/P0001 ,
		\u4_u1_ep_match_r_reg/P0001 ,
		\u4_u1_r5_reg/NET0131 ,
		_w7048_
	);
	LUT4 #(
		.INIT('h2a22)
	) name5299 (
		\u4_u1_csr1_reg[0]/P0001 ,
		_w7045_,
		_w7047_,
		_w7048_,
		_w7049_
	);
	LUT2 #(
		.INIT('h4)
	) name5300 (
		_w7046_,
		_w7049_,
		_w7050_
	);
	LUT4 #(
		.INIT('h6f3f)
	) name5301 (
		\u4_u1_dma_out_cnt_reg[2]/P0001 ,
		\u4_u1_dma_out_cnt_reg[3]/P0001 ,
		\u4_u1_r5_reg/NET0131 ,
		_w4712_,
		_w7051_
	);
	LUT2 #(
		.INIT('h2)
	) name5302 (
		\u4_u1_csr1_reg[0]/P0001 ,
		_w7051_,
		_w7052_
	);
	LUT2 #(
		.INIT('h6)
	) name5303 (
		\u4_u1_csr0_reg[5]/P0001 ,
		\u4_u1_dma_out_cnt_reg[3]/P0001 ,
		_w7053_
	);
	LUT4 #(
		.INIT('h00f4)
	) name5304 (
		_w4730_,
		_w4731_,
		_w4732_,
		_w7053_,
		_w7054_
	);
	LUT4 #(
		.INIT('h134c)
	) name5305 (
		\u4_u1_csr0_reg[4]/P0001 ,
		\u4_u1_csr0_reg[5]/P0001 ,
		\u4_u1_dma_out_cnt_reg[2]/P0001 ,
		\u4_u1_dma_out_cnt_reg[3]/P0001 ,
		_w7055_
	);
	LUT4 #(
		.INIT('h20aa)
	) name5306 (
		_w4454_,
		_w4730_,
		_w4731_,
		_w7055_,
		_w7056_
	);
	LUT4 #(
		.INIT('h0001)
	) name5307 (
		\u1_u3_buf0_rl_reg/P0001 ,
		\u1_u3_buf0_set_reg/P0001 ,
		\u4_u1_dma_out_cnt_reg[3]/P0001 ,
		\u4_u1_set_r_reg/P0001 ,
		_w7057_
	);
	LUT3 #(
		.INIT('h0e)
	) name5308 (
		\u4_u1_dma_out_cnt_reg[3]/P0001 ,
		\u4_u1_ep_match_r_reg/P0001 ,
		\u4_u1_r5_reg/NET0131 ,
		_w7058_
	);
	LUT3 #(
		.INIT('h20)
	) name5309 (
		\u4_u1_csr1_reg[0]/P0001 ,
		_w7057_,
		_w7058_,
		_w7059_
	);
	LUT3 #(
		.INIT('hb0)
	) name5310 (
		_w7054_,
		_w7056_,
		_w7059_,
		_w7060_
	);
	LUT2 #(
		.INIT('he)
	) name5311 (
		_w7052_,
		_w7060_,
		_w7061_
	);
	LUT2 #(
		.INIT('h6)
	) name5312 (
		\u4_u2_csr0_reg[3]/NET0131 ,
		\u4_u2_dma_out_cnt_reg[1]/P0001 ,
		_w7062_
	);
	LUT3 #(
		.INIT('h90)
	) name5313 (
		\u4_u2_dma_in_cnt_reg[0]/P0001 ,
		\u4_u2_dma_out_cnt_reg[1]/P0001 ,
		\u4_u2_r5_reg/NET0131 ,
		_w7063_
	);
	LUT4 #(
		.INIT('h0082)
	) name5314 (
		_w4610_,
		_w4759_,
		_w7062_,
		_w7063_,
		_w7064_
	);
	LUT4 #(
		.INIT('h0001)
	) name5315 (
		\u1_u3_buf0_rl_reg/P0001 ,
		\u1_u3_buf0_set_reg/P0001 ,
		\u4_u2_dma_out_cnt_reg[1]/P0001 ,
		\u4_u2_set_r_reg/P0001 ,
		_w7065_
	);
	LUT3 #(
		.INIT('h0e)
	) name5316 (
		\u4_u2_dma_out_cnt_reg[1]/P0001 ,
		\u4_u2_ep_match_r_reg/P0001 ,
		\u4_u2_r5_reg/NET0131 ,
		_w7066_
	);
	LUT4 #(
		.INIT('h8a88)
	) name5317 (
		\u4_u2_csr1_reg[0]/P0001 ,
		_w7063_,
		_w7065_,
		_w7066_,
		_w7067_
	);
	LUT2 #(
		.INIT('h4)
	) name5318 (
		_w7064_,
		_w7067_,
		_w7068_
	);
	LUT4 #(
		.INIT('hec80)
	) name5319 (
		\u4_u2_csr0_reg[2]/P0001 ,
		\u4_u2_csr0_reg[3]/NET0131 ,
		\u4_u2_dma_in_cnt_reg[0]/P0001 ,
		\u4_u2_dma_out_cnt_reg[1]/P0001 ,
		_w7069_
	);
	LUT2 #(
		.INIT('h6)
	) name5320 (
		\u4_u2_csr0_reg[4]/P0001 ,
		\u4_u2_dma_out_cnt_reg[2]/P0001 ,
		_w7070_
	);
	LUT4 #(
		.INIT('h1eff)
	) name5321 (
		\u4_u2_dma_in_cnt_reg[0]/P0001 ,
		\u4_u2_dma_out_cnt_reg[1]/P0001 ,
		\u4_u2_dma_out_cnt_reg[2]/P0001 ,
		\u4_u2_r5_reg/NET0131 ,
		_w7071_
	);
	LUT4 #(
		.INIT('h8200)
	) name5322 (
		_w4610_,
		_w7069_,
		_w7070_,
		_w7071_,
		_w7072_
	);
	LUT4 #(
		.INIT('h0001)
	) name5323 (
		\u1_u3_buf0_rl_reg/P0001 ,
		\u1_u3_buf0_set_reg/P0001 ,
		\u4_u2_dma_out_cnt_reg[2]/P0001 ,
		\u4_u2_set_r_reg/P0001 ,
		_w7073_
	);
	LUT3 #(
		.INIT('h0e)
	) name5324 (
		\u4_u2_dma_out_cnt_reg[2]/P0001 ,
		\u4_u2_ep_match_r_reg/P0001 ,
		\u4_u2_r5_reg/NET0131 ,
		_w7074_
	);
	LUT4 #(
		.INIT('h2a22)
	) name5325 (
		\u4_u2_csr1_reg[0]/P0001 ,
		_w7071_,
		_w7073_,
		_w7074_,
		_w7075_
	);
	LUT2 #(
		.INIT('h4)
	) name5326 (
		_w7072_,
		_w7075_,
		_w7076_
	);
	LUT4 #(
		.INIT('h6f3f)
	) name5327 (
		\u4_u2_dma_out_cnt_reg[2]/P0001 ,
		\u4_u2_dma_out_cnt_reg[3]/P0001 ,
		\u4_u2_r5_reg/NET0131 ,
		_w4743_,
		_w7077_
	);
	LUT2 #(
		.INIT('h2)
	) name5328 (
		\u4_u2_csr1_reg[0]/P0001 ,
		_w7077_,
		_w7078_
	);
	LUT2 #(
		.INIT('h6)
	) name5329 (
		\u4_u2_csr0_reg[5]/P0001 ,
		\u4_u2_dma_out_cnt_reg[3]/P0001 ,
		_w7079_
	);
	LUT4 #(
		.INIT('h00f4)
	) name5330 (
		_w4760_,
		_w4761_,
		_w4762_,
		_w7079_,
		_w7080_
	);
	LUT4 #(
		.INIT('h134c)
	) name5331 (
		\u4_u2_csr0_reg[4]/P0001 ,
		\u4_u2_csr0_reg[5]/P0001 ,
		\u4_u2_dma_out_cnt_reg[2]/P0001 ,
		\u4_u2_dma_out_cnt_reg[3]/P0001 ,
		_w7081_
	);
	LUT4 #(
		.INIT('h20aa)
	) name5332 (
		_w4610_,
		_w4760_,
		_w4761_,
		_w7081_,
		_w7082_
	);
	LUT4 #(
		.INIT('h0001)
	) name5333 (
		\u1_u3_buf0_rl_reg/P0001 ,
		\u1_u3_buf0_set_reg/P0001 ,
		\u4_u2_dma_out_cnt_reg[3]/P0001 ,
		\u4_u2_set_r_reg/P0001 ,
		_w7083_
	);
	LUT3 #(
		.INIT('ha8)
	) name5334 (
		\u4_u2_csr1_reg[0]/P0001 ,
		\u4_u2_dma_out_cnt_reg[3]/P0001 ,
		\u4_u2_ep_match_r_reg/P0001 ,
		_w7084_
	);
	LUT3 #(
		.INIT('h10)
	) name5335 (
		\u4_u2_r5_reg/NET0131 ,
		_w7083_,
		_w7084_,
		_w7085_
	);
	LUT3 #(
		.INIT('hb0)
	) name5336 (
		_w7080_,
		_w7082_,
		_w7085_,
		_w7086_
	);
	LUT2 #(
		.INIT('he)
	) name5337 (
		_w7078_,
		_w7086_,
		_w7087_
	);
	LUT2 #(
		.INIT('h9)
	) name5338 (
		\u4_u3_csr0_reg[4]/P0001 ,
		\u4_u3_dma_in_cnt_reg[2]/P0001 ,
		_w7088_
	);
	LUT3 #(
		.INIT('hc8)
	) name5339 (
		_w4560_,
		_w4569_,
		_w7088_,
		_w7089_
	);
	LUT4 #(
		.INIT('h87ff)
	) name5340 (
		\u4_u3_dma_in_cnt_reg[0]/P0001 ,
		\u4_u3_dma_in_cnt_reg[1]/P0001 ,
		\u4_u3_dma_in_cnt_reg[2]/P0001 ,
		\u4_u3_r5_reg/NET0131 ,
		_w7090_
	);
	LUT4 #(
		.INIT('hfb00)
	) name5341 (
		_w4384_,
		_w4385_,
		_w4388_,
		_w7090_,
		_w7091_
	);
	LUT4 #(
		.INIT('h0001)
	) name5342 (
		\u1_u3_buf0_rl_reg/P0001 ,
		\u1_u3_buf0_set_reg/P0001 ,
		\u4_u3_dma_in_cnt_reg[2]/P0001 ,
		\u4_u3_set_r_reg/P0001 ,
		_w7092_
	);
	LUT3 #(
		.INIT('h0e)
	) name5343 (
		\u4_u3_dma_in_cnt_reg[2]/P0001 ,
		\u4_u3_ep_match_r_reg/P0001 ,
		\u4_u3_r5_reg/NET0131 ,
		_w7093_
	);
	LUT4 #(
		.INIT('h2a22)
	) name5344 (
		\u4_u3_csr1_reg[0]/P0001 ,
		_w7090_,
		_w7092_,
		_w7093_,
		_w7094_
	);
	LUT3 #(
		.INIT('h70)
	) name5345 (
		_w7089_,
		_w7091_,
		_w7094_,
		_w7095_
	);
	LUT2 #(
		.INIT('h8)
	) name5346 (
		\u4_u3_csr1_reg[0]/P0001 ,
		\u4_u3_dma_in_cnt_reg[3]/P0001 ,
		_w7096_
	);
	LUT4 #(
		.INIT('h8000)
	) name5347 (
		\u4_u3_csr1_reg[0]/P0001 ,
		\u4_u3_dma_in_cnt_reg[0]/P0001 ,
		\u4_u3_dma_in_cnt_reg[1]/P0001 ,
		\u4_u3_dma_in_cnt_reg[2]/P0001 ,
		_w7097_
	);
	LUT4 #(
		.INIT('h2220)
	) name5348 (
		\u4_u3_r5_reg/NET0131 ,
		_w4399_,
		_w7096_,
		_w7097_,
		_w7098_
	);
	LUT2 #(
		.INIT('h9)
	) name5349 (
		\u4_u3_csr0_reg[5]/P0001 ,
		\u4_u3_dma_in_cnt_reg[3]/P0001 ,
		_w7099_
	);
	LUT4 #(
		.INIT('hf400)
	) name5350 (
		_w4384_,
		_w4385_,
		_w4388_,
		_w7099_,
		_w7100_
	);
	LUT4 #(
		.INIT('h31c4)
	) name5351 (
		\u4_u3_csr0_reg[4]/P0001 ,
		\u4_u3_csr0_reg[5]/P0001 ,
		\u4_u3_dma_in_cnt_reg[2]/P0001 ,
		\u4_u3_dma_in_cnt_reg[3]/P0001 ,
		_w7101_
	);
	LUT4 #(
		.INIT('h40f0)
	) name5352 (
		_w4384_,
		_w4385_,
		_w4569_,
		_w7101_,
		_w7102_
	);
	LUT4 #(
		.INIT('h0001)
	) name5353 (
		\u1_u3_buf0_rl_reg/P0001 ,
		\u1_u3_buf0_set_reg/P0001 ,
		\u4_u3_dma_in_cnt_reg[3]/P0001 ,
		\u4_u3_set_r_reg/P0001 ,
		_w7103_
	);
	LUT3 #(
		.INIT('ha8)
	) name5354 (
		\u4_u3_csr1_reg[0]/P0001 ,
		\u4_u3_dma_in_cnt_reg[3]/P0001 ,
		\u4_u3_ep_match_r_reg/P0001 ,
		_w7104_
	);
	LUT3 #(
		.INIT('h10)
	) name5355 (
		\u4_u3_r5_reg/NET0131 ,
		_w7103_,
		_w7104_,
		_w7105_
	);
	LUT4 #(
		.INIT('hefaa)
	) name5356 (
		_w7098_,
		_w7100_,
		_w7102_,
		_w7105_,
		_w7106_
	);
	LUT3 #(
		.INIT('h10)
	) name5357 (
		\u4_u3_dma_out_cnt_reg[4]/P0001 ,
		\u4_u3_dma_out_cnt_reg[5]/P0001 ,
		\u4_u3_r5_reg/NET0131 ,
		_w7107_
	);
	LUT3 #(
		.INIT('h80)
	) name5358 (
		\u4_u3_csr1_reg[0]/P0001 ,
		_w4652_,
		_w7107_,
		_w7108_
	);
	LUT3 #(
		.INIT('h80)
	) name5359 (
		\u4_u3_csr1_reg[0]/P0001 ,
		\u4_u3_dma_out_cnt_reg[5]/P0001 ,
		\u4_u3_r5_reg/NET0131 ,
		_w7109_
	);
	LUT3 #(
		.INIT('hb0)
	) name5360 (
		\u4_u3_dma_out_cnt_reg[4]/P0001 ,
		_w4652_,
		_w7109_,
		_w7110_
	);
	LUT2 #(
		.INIT('h1)
	) name5361 (
		_w7108_,
		_w7110_,
		_w7111_
	);
	LUT2 #(
		.INIT('h6)
	) name5362 (
		\u4_u3_csr0_reg[7]/P0001 ,
		\u4_u3_dma_out_cnt_reg[5]/P0001 ,
		_w7112_
	);
	LUT4 #(
		.INIT('hfe00)
	) name5363 (
		_w4667_,
		_w4672_,
		_w4673_,
		_w7112_,
		_w7113_
	);
	LUT4 #(
		.INIT('hc832)
	) name5364 (
		\u4_u3_csr0_reg[6]/P0001 ,
		\u4_u3_csr0_reg[7]/P0001 ,
		\u4_u3_dma_out_cnt_reg[4]/P0001 ,
		\u4_u3_dma_out_cnt_reg[5]/P0001 ,
		_w7114_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name5365 (
		_w4569_,
		_w4667_,
		_w4672_,
		_w7114_,
		_w7115_
	);
	LUT4 #(
		.INIT('h0001)
	) name5366 (
		\u1_u3_buf0_rl_reg/P0001 ,
		\u1_u3_buf0_set_reg/P0001 ,
		\u4_u3_dma_out_cnt_reg[5]/P0001 ,
		\u4_u3_set_r_reg/P0001 ,
		_w7116_
	);
	LUT3 #(
		.INIT('ha8)
	) name5367 (
		\u4_u3_csr1_reg[0]/P0001 ,
		\u4_u3_dma_out_cnt_reg[5]/P0001 ,
		\u4_u3_ep_match_r_reg/P0001 ,
		_w7117_
	);
	LUT3 #(
		.INIT('h10)
	) name5368 (
		\u4_u3_r5_reg/NET0131 ,
		_w7116_,
		_w7117_,
		_w7118_
	);
	LUT4 #(
		.INIT('hdf55)
	) name5369 (
		_w7111_,
		_w7113_,
		_w7115_,
		_w7118_,
		_w7119_
	);
	LUT2 #(
		.INIT('h9)
	) name5370 (
		\u4_u0_csr0_reg[4]/P0001 ,
		\u4_u0_dma_in_cnt_reg[2]/P0001 ,
		_w7120_
	);
	LUT3 #(
		.INIT('hc8)
	) name5371 (
		_w4583_,
		_w4592_,
		_w7120_,
		_w7121_
	);
	LUT4 #(
		.INIT('h87ff)
	) name5372 (
		\u4_u0_dma_in_cnt_reg[0]/P0001 ,
		\u4_u0_dma_in_cnt_reg[1]/P0001 ,
		\u4_u0_dma_in_cnt_reg[2]/P0001 ,
		\u4_u0_r5_reg/NET0131 ,
		_w7122_
	);
	LUT4 #(
		.INIT('hfb00)
	) name5373 (
		_w4416_,
		_w4417_,
		_w4420_,
		_w7122_,
		_w7123_
	);
	LUT4 #(
		.INIT('h0001)
	) name5374 (
		\u1_u3_buf0_rl_reg/P0001 ,
		\u1_u3_buf0_set_reg/P0001 ,
		\u4_u0_dma_in_cnt_reg[2]/P0001 ,
		\u4_u0_set_r_reg/P0001 ,
		_w7124_
	);
	LUT3 #(
		.INIT('h0e)
	) name5375 (
		\u4_u0_dma_in_cnt_reg[2]/P0001 ,
		\u4_u0_ep_match_r_reg/P0001 ,
		\u4_u0_r5_reg/NET0131 ,
		_w7125_
	);
	LUT4 #(
		.INIT('h2a22)
	) name5376 (
		\u4_u0_csr1_reg[0]/P0001 ,
		_w7122_,
		_w7124_,
		_w7125_,
		_w7126_
	);
	LUT3 #(
		.INIT('h70)
	) name5377 (
		_w7121_,
		_w7123_,
		_w7126_,
		_w7127_
	);
	LUT2 #(
		.INIT('h8)
	) name5378 (
		\u4_u0_csr1_reg[0]/P0001 ,
		\u4_u0_dma_in_cnt_reg[3]/P0001 ,
		_w7128_
	);
	LUT4 #(
		.INIT('h8000)
	) name5379 (
		\u4_u0_csr1_reg[0]/P0001 ,
		\u4_u0_dma_in_cnt_reg[0]/P0001 ,
		\u4_u0_dma_in_cnt_reg[1]/P0001 ,
		\u4_u0_dma_in_cnt_reg[2]/P0001 ,
		_w7129_
	);
	LUT4 #(
		.INIT('h2220)
	) name5380 (
		\u4_u0_r5_reg/NET0131 ,
		_w4431_,
		_w7128_,
		_w7129_,
		_w7130_
	);
	LUT2 #(
		.INIT('h9)
	) name5381 (
		\u4_u0_csr0_reg[5]/P0001 ,
		\u4_u0_dma_in_cnt_reg[3]/P0001 ,
		_w7131_
	);
	LUT4 #(
		.INIT('hf400)
	) name5382 (
		_w4416_,
		_w4417_,
		_w4420_,
		_w7131_,
		_w7132_
	);
	LUT4 #(
		.INIT('h31c4)
	) name5383 (
		\u4_u0_csr0_reg[4]/P0001 ,
		\u4_u0_csr0_reg[5]/P0001 ,
		\u4_u0_dma_in_cnt_reg[2]/P0001 ,
		\u4_u0_dma_in_cnt_reg[3]/P0001 ,
		_w7133_
	);
	LUT4 #(
		.INIT('h40f0)
	) name5384 (
		_w4416_,
		_w4417_,
		_w4592_,
		_w7133_,
		_w7134_
	);
	LUT4 #(
		.INIT('h0001)
	) name5385 (
		\u1_u3_buf0_rl_reg/P0001 ,
		\u1_u3_buf0_set_reg/P0001 ,
		\u4_u0_dma_in_cnt_reg[3]/P0001 ,
		\u4_u0_set_r_reg/P0001 ,
		_w7135_
	);
	LUT3 #(
		.INIT('ha8)
	) name5386 (
		\u4_u0_csr1_reg[0]/P0001 ,
		\u4_u0_dma_in_cnt_reg[3]/P0001 ,
		\u4_u0_ep_match_r_reg/P0001 ,
		_w7136_
	);
	LUT3 #(
		.INIT('h10)
	) name5387 (
		\u4_u0_r5_reg/NET0131 ,
		_w7135_,
		_w7136_,
		_w7137_
	);
	LUT4 #(
		.INIT('hefaa)
	) name5388 (
		_w7130_,
		_w7132_,
		_w7134_,
		_w7137_,
		_w7138_
	);
	LUT3 #(
		.INIT('h80)
	) name5389 (
		\u4_u0_csr1_reg[0]/P0001 ,
		_w4683_,
		_w4989_,
		_w7139_
	);
	LUT3 #(
		.INIT('h80)
	) name5390 (
		\u4_u0_csr1_reg[0]/P0001 ,
		\u4_u0_dma_out_cnt_reg[5]/P0001 ,
		\u4_u0_r5_reg/NET0131 ,
		_w7140_
	);
	LUT3 #(
		.INIT('hb0)
	) name5391 (
		\u4_u0_dma_out_cnt_reg[4]/P0001 ,
		_w4683_,
		_w7140_,
		_w7141_
	);
	LUT2 #(
		.INIT('h1)
	) name5392 (
		_w7139_,
		_w7141_,
		_w7142_
	);
	LUT2 #(
		.INIT('h6)
	) name5393 (
		\u4_u0_csr0_reg[7]/P0001 ,
		\u4_u0_dma_out_cnt_reg[5]/P0001 ,
		_w7143_
	);
	LUT4 #(
		.INIT('hfe00)
	) name5394 (
		_w4697_,
		_w4702_,
		_w4703_,
		_w7143_,
		_w7144_
	);
	LUT4 #(
		.INIT('hc832)
	) name5395 (
		\u4_u0_csr0_reg[6]/P0001 ,
		\u4_u0_csr0_reg[7]/P0001 ,
		\u4_u0_dma_out_cnt_reg[4]/P0001 ,
		\u4_u0_dma_out_cnt_reg[5]/P0001 ,
		_w7145_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name5396 (
		_w4592_,
		_w4697_,
		_w4702_,
		_w7145_,
		_w7146_
	);
	LUT4 #(
		.INIT('h0001)
	) name5397 (
		\u1_u3_buf0_rl_reg/P0001 ,
		\u1_u3_buf0_set_reg/P0001 ,
		\u4_u0_dma_out_cnt_reg[5]/P0001 ,
		\u4_u0_set_r_reg/P0001 ,
		_w7147_
	);
	LUT3 #(
		.INIT('ha8)
	) name5398 (
		\u4_u0_csr1_reg[0]/P0001 ,
		\u4_u0_dma_out_cnt_reg[5]/P0001 ,
		\u4_u0_ep_match_r_reg/P0001 ,
		_w7148_
	);
	LUT3 #(
		.INIT('h10)
	) name5399 (
		\u4_u0_r5_reg/NET0131 ,
		_w7147_,
		_w7148_,
		_w7149_
	);
	LUT4 #(
		.INIT('hdf55)
	) name5400 (
		_w7142_,
		_w7144_,
		_w7146_,
		_w7149_,
		_w7150_
	);
	LUT4 #(
		.INIT('h08ce)
	) name5401 (
		\u4_u1_csr0_reg[2]/P0001 ,
		\u4_u1_csr0_reg[3]/NET0131 ,
		\u4_u1_dma_in_cnt_reg[0]/P0001 ,
		\u4_u1_dma_in_cnt_reg[1]/P0001 ,
		_w7151_
	);
	LUT2 #(
		.INIT('h9)
	) name5402 (
		\u4_u1_csr0_reg[4]/P0001 ,
		\u4_u1_dma_in_cnt_reg[2]/P0001 ,
		_w7152_
	);
	LUT4 #(
		.INIT('h87ff)
	) name5403 (
		\u4_u1_dma_in_cnt_reg[0]/P0001 ,
		\u4_u1_dma_in_cnt_reg[1]/P0001 ,
		\u4_u1_dma_in_cnt_reg[2]/P0001 ,
		\u4_u1_r5_reg/NET0131 ,
		_w7153_
	);
	LUT4 #(
		.INIT('h2800)
	) name5404 (
		_w4454_,
		_w7151_,
		_w7152_,
		_w7153_,
		_w7154_
	);
	LUT4 #(
		.INIT('h0001)
	) name5405 (
		\u1_u3_buf0_rl_reg/P0001 ,
		\u1_u3_buf0_set_reg/P0001 ,
		\u4_u1_dma_in_cnt_reg[2]/P0001 ,
		\u4_u1_set_r_reg/P0001 ,
		_w7155_
	);
	LUT3 #(
		.INIT('h0e)
	) name5406 (
		\u4_u1_dma_in_cnt_reg[2]/P0001 ,
		\u4_u1_ep_match_r_reg/P0001 ,
		\u4_u1_r5_reg/NET0131 ,
		_w7156_
	);
	LUT4 #(
		.INIT('h2a22)
	) name5407 (
		\u4_u1_csr1_reg[0]/P0001 ,
		_w7153_,
		_w7155_,
		_w7156_,
		_w7157_
	);
	LUT2 #(
		.INIT('h4)
	) name5408 (
		_w7154_,
		_w7157_,
		_w7158_
	);
	LUT2 #(
		.INIT('h8)
	) name5409 (
		\u4_u1_csr1_reg[0]/P0001 ,
		\u4_u1_dma_in_cnt_reg[3]/P0001 ,
		_w7159_
	);
	LUT4 #(
		.INIT('h8000)
	) name5410 (
		\u4_u1_csr1_reg[0]/P0001 ,
		\u4_u1_dma_in_cnt_reg[0]/P0001 ,
		\u4_u1_dma_in_cnt_reg[1]/P0001 ,
		\u4_u1_dma_in_cnt_reg[2]/P0001 ,
		_w7160_
	);
	LUT4 #(
		.INIT('h2220)
	) name5411 (
		\u4_u1_r5_reg/NET0131 ,
		_w4448_,
		_w7159_,
		_w7160_,
		_w7161_
	);
	LUT2 #(
		.INIT('h9)
	) name5412 (
		\u4_u1_csr0_reg[5]/P0001 ,
		\u4_u1_dma_in_cnt_reg[3]/P0001 ,
		_w7162_
	);
	LUT4 #(
		.INIT('hf400)
	) name5413 (
		_w4465_,
		_w4466_,
		_w4467_,
		_w7162_,
		_w7163_
	);
	LUT4 #(
		.INIT('h31c4)
	) name5414 (
		\u4_u1_csr0_reg[4]/P0001 ,
		\u4_u1_csr0_reg[5]/P0001 ,
		\u4_u1_dma_in_cnt_reg[2]/P0001 ,
		\u4_u1_dma_in_cnt_reg[3]/P0001 ,
		_w7164_
	);
	LUT4 #(
		.INIT('h20aa)
	) name5415 (
		_w4454_,
		_w4465_,
		_w4466_,
		_w7164_,
		_w7165_
	);
	LUT4 #(
		.INIT('h0001)
	) name5416 (
		\u1_u3_buf0_rl_reg/P0001 ,
		\u1_u3_buf0_set_reg/P0001 ,
		\u4_u1_dma_in_cnt_reg[3]/P0001 ,
		\u4_u1_set_r_reg/P0001 ,
		_w7166_
	);
	LUT3 #(
		.INIT('ha8)
	) name5417 (
		\u4_u1_csr1_reg[0]/P0001 ,
		\u4_u1_dma_in_cnt_reg[3]/P0001 ,
		\u4_u1_ep_match_r_reg/P0001 ,
		_w7167_
	);
	LUT3 #(
		.INIT('h10)
	) name5418 (
		\u4_u1_r5_reg/NET0131 ,
		_w7166_,
		_w7167_,
		_w7168_
	);
	LUT4 #(
		.INIT('hefaa)
	) name5419 (
		_w7161_,
		_w7163_,
		_w7165_,
		_w7168_,
		_w7169_
	);
	LUT3 #(
		.INIT('h80)
	) name5420 (
		\u4_u1_csr1_reg[0]/P0001 ,
		_w4713_,
		_w5023_,
		_w7170_
	);
	LUT3 #(
		.INIT('h80)
	) name5421 (
		\u4_u1_csr1_reg[0]/P0001 ,
		\u4_u1_dma_out_cnt_reg[5]/P0001 ,
		\u4_u1_r5_reg/NET0131 ,
		_w7171_
	);
	LUT3 #(
		.INIT('hb0)
	) name5422 (
		\u4_u1_dma_out_cnt_reg[4]/P0001 ,
		_w4713_,
		_w7171_,
		_w7172_
	);
	LUT2 #(
		.INIT('h1)
	) name5423 (
		_w7170_,
		_w7172_,
		_w7173_
	);
	LUT2 #(
		.INIT('h6)
	) name5424 (
		\u4_u1_csr0_reg[7]/P0001 ,
		\u4_u1_dma_out_cnt_reg[5]/P0001 ,
		_w7174_
	);
	LUT4 #(
		.INIT('hfe00)
	) name5425 (
		_w4728_,
		_w4733_,
		_w4734_,
		_w7174_,
		_w7175_
	);
	LUT4 #(
		.INIT('hc832)
	) name5426 (
		\u4_u1_csr0_reg[6]/P0001 ,
		\u4_u1_csr0_reg[7]/P0001 ,
		\u4_u1_dma_out_cnt_reg[4]/P0001 ,
		\u4_u1_dma_out_cnt_reg[5]/P0001 ,
		_w7176_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name5427 (
		_w4454_,
		_w4728_,
		_w4733_,
		_w7176_,
		_w7177_
	);
	LUT4 #(
		.INIT('h0001)
	) name5428 (
		\u1_u3_buf0_rl_reg/P0001 ,
		\u1_u3_buf0_set_reg/P0001 ,
		\u4_u1_dma_out_cnt_reg[5]/P0001 ,
		\u4_u1_set_r_reg/P0001 ,
		_w7178_
	);
	LUT3 #(
		.INIT('ha8)
	) name5429 (
		\u4_u1_csr1_reg[0]/P0001 ,
		\u4_u1_dma_out_cnt_reg[5]/P0001 ,
		\u4_u1_ep_match_r_reg/P0001 ,
		_w7179_
	);
	LUT3 #(
		.INIT('h10)
	) name5430 (
		\u4_u1_r5_reg/NET0131 ,
		_w7178_,
		_w7179_,
		_w7180_
	);
	LUT4 #(
		.INIT('hdf55)
	) name5431 (
		_w7173_,
		_w7175_,
		_w7177_,
		_w7180_,
		_w7181_
	);
	LUT4 #(
		.INIT('h08ce)
	) name5432 (
		\u4_u2_csr0_reg[2]/P0001 ,
		\u4_u2_csr0_reg[3]/NET0131 ,
		\u4_u2_dma_in_cnt_reg[0]/P0001 ,
		\u4_u2_dma_in_cnt_reg[1]/P0001 ,
		_w7182_
	);
	LUT2 #(
		.INIT('h9)
	) name5433 (
		\u4_u2_csr0_reg[4]/P0001 ,
		\u4_u2_dma_in_cnt_reg[2]/P0001 ,
		_w7183_
	);
	LUT4 #(
		.INIT('h87ff)
	) name5434 (
		\u4_u2_dma_in_cnt_reg[0]/P0001 ,
		\u4_u2_dma_in_cnt_reg[1]/P0001 ,
		\u4_u2_dma_in_cnt_reg[2]/P0001 ,
		\u4_u2_r5_reg/NET0131 ,
		_w7184_
	);
	LUT4 #(
		.INIT('h2800)
	) name5435 (
		_w4610_,
		_w7182_,
		_w7183_,
		_w7184_,
		_w7185_
	);
	LUT4 #(
		.INIT('h0001)
	) name5436 (
		\u1_u3_buf0_rl_reg/P0001 ,
		\u1_u3_buf0_set_reg/P0001 ,
		\u4_u2_dma_in_cnt_reg[2]/P0001 ,
		\u4_u2_set_r_reg/P0001 ,
		_w7186_
	);
	LUT3 #(
		.INIT('h0e)
	) name5437 (
		\u4_u2_dma_in_cnt_reg[2]/P0001 ,
		\u4_u2_ep_match_r_reg/P0001 ,
		\u4_u2_r5_reg/NET0131 ,
		_w7187_
	);
	LUT4 #(
		.INIT('h2a22)
	) name5438 (
		\u4_u2_csr1_reg[0]/P0001 ,
		_w7184_,
		_w7186_,
		_w7187_,
		_w7188_
	);
	LUT2 #(
		.INIT('h4)
	) name5439 (
		_w7185_,
		_w7188_,
		_w7189_
	);
	LUT2 #(
		.INIT('h8)
	) name5440 (
		\u4_u2_csr1_reg[0]/P0001 ,
		\u4_u2_dma_in_cnt_reg[3]/P0001 ,
		_w7190_
	);
	LUT4 #(
		.INIT('h8000)
	) name5441 (
		\u4_u2_csr1_reg[0]/P0001 ,
		\u4_u2_dma_in_cnt_reg[0]/P0001 ,
		\u4_u2_dma_in_cnt_reg[1]/P0001 ,
		\u4_u2_dma_in_cnt_reg[2]/P0001 ,
		_w7191_
	);
	LUT4 #(
		.INIT('h2220)
	) name5442 (
		\u4_u2_r5_reg/NET0131 ,
		_w4505_,
		_w7190_,
		_w7191_,
		_w7192_
	);
	LUT2 #(
		.INIT('h9)
	) name5443 (
		\u4_u2_csr0_reg[5]/P0001 ,
		\u4_u2_dma_in_cnt_reg[3]/P0001 ,
		_w7193_
	);
	LUT4 #(
		.INIT('hf400)
	) name5444 (
		_w4493_,
		_w4494_,
		_w4495_,
		_w7193_,
		_w7194_
	);
	LUT4 #(
		.INIT('h31c4)
	) name5445 (
		\u4_u2_csr0_reg[4]/P0001 ,
		\u4_u2_csr0_reg[5]/P0001 ,
		\u4_u2_dma_in_cnt_reg[2]/P0001 ,
		\u4_u2_dma_in_cnt_reg[3]/P0001 ,
		_w7195_
	);
	LUT4 #(
		.INIT('h40f0)
	) name5446 (
		_w4493_,
		_w4494_,
		_w4610_,
		_w7195_,
		_w7196_
	);
	LUT4 #(
		.INIT('h0001)
	) name5447 (
		\u1_u3_buf0_rl_reg/P0001 ,
		\u1_u3_buf0_set_reg/P0001 ,
		\u4_u2_dma_in_cnt_reg[3]/P0001 ,
		\u4_u2_set_r_reg/P0001 ,
		_w7197_
	);
	LUT3 #(
		.INIT('ha8)
	) name5448 (
		\u4_u2_csr1_reg[0]/P0001 ,
		\u4_u2_dma_in_cnt_reg[3]/P0001 ,
		\u4_u2_ep_match_r_reg/P0001 ,
		_w7198_
	);
	LUT3 #(
		.INIT('h10)
	) name5449 (
		\u4_u2_r5_reg/NET0131 ,
		_w7197_,
		_w7198_,
		_w7199_
	);
	LUT4 #(
		.INIT('hefaa)
	) name5450 (
		_w7192_,
		_w7194_,
		_w7196_,
		_w7199_,
		_w7200_
	);
	LUT3 #(
		.INIT('h10)
	) name5451 (
		\u4_u2_dma_out_cnt_reg[4]/P0001 ,
		\u4_u2_dma_out_cnt_reg[5]/P0001 ,
		\u4_u2_r5_reg/NET0131 ,
		_w7201_
	);
	LUT3 #(
		.INIT('h80)
	) name5452 (
		\u4_u2_csr1_reg[0]/P0001 ,
		_w4744_,
		_w7201_,
		_w7202_
	);
	LUT3 #(
		.INIT('h80)
	) name5453 (
		\u4_u2_csr1_reg[0]/P0001 ,
		\u4_u2_dma_out_cnt_reg[5]/P0001 ,
		\u4_u2_r5_reg/NET0131 ,
		_w7203_
	);
	LUT3 #(
		.INIT('hb0)
	) name5454 (
		\u4_u2_dma_out_cnt_reg[4]/P0001 ,
		_w4744_,
		_w7203_,
		_w7204_
	);
	LUT2 #(
		.INIT('h1)
	) name5455 (
		_w7202_,
		_w7204_,
		_w7205_
	);
	LUT2 #(
		.INIT('h6)
	) name5456 (
		\u4_u2_csr0_reg[7]/P0001 ,
		\u4_u2_dma_out_cnt_reg[5]/P0001 ,
		_w7206_
	);
	LUT4 #(
		.INIT('hfe00)
	) name5457 (
		_w4758_,
		_w4763_,
		_w4764_,
		_w7206_,
		_w7207_
	);
	LUT4 #(
		.INIT('hc832)
	) name5458 (
		\u4_u2_csr0_reg[6]/P0001 ,
		\u4_u2_csr0_reg[7]/P0001 ,
		\u4_u2_dma_out_cnt_reg[4]/P0001 ,
		\u4_u2_dma_out_cnt_reg[5]/P0001 ,
		_w7208_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name5459 (
		_w4610_,
		_w4758_,
		_w4763_,
		_w7208_,
		_w7209_
	);
	LUT4 #(
		.INIT('h0001)
	) name5460 (
		\u1_u3_buf0_rl_reg/P0001 ,
		\u1_u3_buf0_set_reg/P0001 ,
		\u4_u2_dma_out_cnt_reg[5]/P0001 ,
		\u4_u2_set_r_reg/P0001 ,
		_w7210_
	);
	LUT3 #(
		.INIT('ha8)
	) name5461 (
		\u4_u2_csr1_reg[0]/P0001 ,
		\u4_u2_dma_out_cnt_reg[5]/P0001 ,
		\u4_u2_ep_match_r_reg/P0001 ,
		_w7211_
	);
	LUT3 #(
		.INIT('h10)
	) name5462 (
		\u4_u2_r5_reg/NET0131 ,
		_w7210_,
		_w7211_,
		_w7212_
	);
	LUT4 #(
		.INIT('hdf55)
	) name5463 (
		_w7205_,
		_w7207_,
		_w7209_,
		_w7212_,
		_w7213_
	);
	LUT4 #(
		.INIT('hf800)
	) name5464 (
		\u0_u0_idle_cnt1_reg[0]/P0001 ,
		\u0_u0_idle_cnt1_reg[1]/P0001 ,
		\u0_u0_idle_cnt1_reg[2]/P0001 ,
		\u0_u0_idle_cnt1_reg[3]/P0001 ,
		_w7214_
	);
	LUT2 #(
		.INIT('h1)
	) name5465 (
		\u0_u0_idle_cnt1_reg[6]/P0001 ,
		\u0_u0_idle_cnt1_reg[7]/P0001 ,
		_w7215_
	);
	LUT4 #(
		.INIT('h0001)
	) name5466 (
		\u0_u0_idle_cnt1_reg[4]/P0001 ,
		\u0_u0_idle_cnt1_reg[5]/P0001 ,
		\u0_u0_idle_cnt1_reg[6]/P0001 ,
		\u0_u0_idle_cnt1_reg[7]/P0001 ,
		_w7216_
	);
	LUT2 #(
		.INIT('h4)
	) name5467 (
		_w7214_,
		_w7216_,
		_w7217_
	);
	LUT3 #(
		.INIT('h0d)
	) name5468 (
		_w5763_,
		_w5768_,
		_w7217_,
		_w7218_
	);
	LUT2 #(
		.INIT('h4)
	) name5469 (
		_w5765_,
		_w7218_,
		_w7219_
	);
	LUT2 #(
		.INIT('h9)
	) name5470 (
		\u4_u3_csr0_reg[3]/NET0131 ,
		\u4_u3_dma_in_cnt_reg[1]/P0001 ,
		_w7220_
	);
	LUT3 #(
		.INIT('h60)
	) name5471 (
		\u4_u3_dma_in_cnt_reg[0]/P0001 ,
		\u4_u3_dma_in_cnt_reg[1]/P0001 ,
		\u4_u3_r5_reg/NET0131 ,
		_w7221_
	);
	LUT4 #(
		.INIT('h0048)
	) name5472 (
		_w4383_,
		_w4569_,
		_w7220_,
		_w7221_,
		_w7222_
	);
	LUT4 #(
		.INIT('h0001)
	) name5473 (
		\u1_u3_buf0_rl_reg/P0001 ,
		\u1_u3_buf0_set_reg/P0001 ,
		\u4_u3_dma_in_cnt_reg[1]/P0001 ,
		\u4_u3_set_r_reg/P0001 ,
		_w7223_
	);
	LUT3 #(
		.INIT('h0e)
	) name5474 (
		\u4_u3_dma_in_cnt_reg[1]/P0001 ,
		\u4_u3_ep_match_r_reg/P0001 ,
		\u4_u3_r5_reg/NET0131 ,
		_w7224_
	);
	LUT4 #(
		.INIT('h8a88)
	) name5475 (
		\u4_u3_csr1_reg[0]/P0001 ,
		_w7221_,
		_w7223_,
		_w7224_,
		_w7225_
	);
	LUT2 #(
		.INIT('h4)
	) name5476 (
		_w7222_,
		_w7225_,
		_w7226_
	);
	LUT2 #(
		.INIT('h9)
	) name5477 (
		\u4_u0_csr0_reg[3]/NET0131 ,
		\u4_u0_dma_in_cnt_reg[1]/P0001 ,
		_w7227_
	);
	LUT3 #(
		.INIT('h60)
	) name5478 (
		\u4_u0_dma_in_cnt_reg[0]/P0001 ,
		\u4_u0_dma_in_cnt_reg[1]/P0001 ,
		\u4_u0_r5_reg/NET0131 ,
		_w7228_
	);
	LUT4 #(
		.INIT('h0048)
	) name5479 (
		_w4415_,
		_w4592_,
		_w7227_,
		_w7228_,
		_w7229_
	);
	LUT4 #(
		.INIT('h0001)
	) name5480 (
		\u1_u3_buf0_rl_reg/P0001 ,
		\u1_u3_buf0_set_reg/P0001 ,
		\u4_u0_dma_in_cnt_reg[1]/P0001 ,
		\u4_u0_set_r_reg/P0001 ,
		_w7230_
	);
	LUT3 #(
		.INIT('h0e)
	) name5481 (
		\u4_u0_dma_in_cnt_reg[1]/P0001 ,
		\u4_u0_ep_match_r_reg/P0001 ,
		\u4_u0_r5_reg/NET0131 ,
		_w7231_
	);
	LUT4 #(
		.INIT('h8a88)
	) name5482 (
		\u4_u0_csr1_reg[0]/P0001 ,
		_w7228_,
		_w7230_,
		_w7231_,
		_w7232_
	);
	LUT2 #(
		.INIT('h4)
	) name5483 (
		_w7229_,
		_w7232_,
		_w7233_
	);
	LUT2 #(
		.INIT('h9)
	) name5484 (
		\u4_u1_csr0_reg[3]/NET0131 ,
		\u4_u1_dma_in_cnt_reg[1]/P0001 ,
		_w7234_
	);
	LUT3 #(
		.INIT('h60)
	) name5485 (
		\u4_u1_dma_in_cnt_reg[0]/P0001 ,
		\u4_u1_dma_in_cnt_reg[1]/P0001 ,
		\u4_u1_r5_reg/NET0131 ,
		_w7235_
	);
	LUT4 #(
		.INIT('h0028)
	) name5486 (
		_w4454_,
		_w4464_,
		_w7234_,
		_w7235_,
		_w7236_
	);
	LUT4 #(
		.INIT('h0001)
	) name5487 (
		\u1_u3_buf0_rl_reg/P0001 ,
		\u1_u3_buf0_set_reg/P0001 ,
		\u4_u1_dma_in_cnt_reg[1]/P0001 ,
		\u4_u1_set_r_reg/P0001 ,
		_w7237_
	);
	LUT3 #(
		.INIT('h0e)
	) name5488 (
		\u4_u1_dma_in_cnt_reg[1]/P0001 ,
		\u4_u1_ep_match_r_reg/P0001 ,
		\u4_u1_r5_reg/NET0131 ,
		_w7238_
	);
	LUT4 #(
		.INIT('h8a88)
	) name5489 (
		\u4_u1_csr1_reg[0]/P0001 ,
		_w7235_,
		_w7237_,
		_w7238_,
		_w7239_
	);
	LUT2 #(
		.INIT('h4)
	) name5490 (
		_w7236_,
		_w7239_,
		_w7240_
	);
	LUT2 #(
		.INIT('h9)
	) name5491 (
		\u4_u2_csr0_reg[3]/NET0131 ,
		\u4_u2_dma_in_cnt_reg[1]/P0001 ,
		_w7241_
	);
	LUT3 #(
		.INIT('h60)
	) name5492 (
		\u4_u2_dma_in_cnt_reg[0]/P0001 ,
		\u4_u2_dma_in_cnt_reg[1]/P0001 ,
		\u4_u2_r5_reg/NET0131 ,
		_w7242_
	);
	LUT4 #(
		.INIT('h0048)
	) name5493 (
		_w4492_,
		_w4610_,
		_w7241_,
		_w7242_,
		_w7243_
	);
	LUT4 #(
		.INIT('h0001)
	) name5494 (
		\u1_u3_buf0_rl_reg/P0001 ,
		\u1_u3_buf0_set_reg/P0001 ,
		\u4_u2_dma_in_cnt_reg[1]/P0001 ,
		\u4_u2_set_r_reg/P0001 ,
		_w7244_
	);
	LUT3 #(
		.INIT('h0e)
	) name5495 (
		\u4_u2_dma_in_cnt_reg[1]/P0001 ,
		\u4_u2_ep_match_r_reg/P0001 ,
		\u4_u2_r5_reg/NET0131 ,
		_w7245_
	);
	LUT4 #(
		.INIT('h8a88)
	) name5496 (
		\u4_u2_csr1_reg[0]/P0001 ,
		_w7242_,
		_w7244_,
		_w7245_,
		_w7246_
	);
	LUT2 #(
		.INIT('h4)
	) name5497 (
		_w7243_,
		_w7246_,
		_w7247_
	);
	LUT3 #(
		.INIT('h20)
	) name5498 (
		rst_i_pad,
		\u4_u2_int_re_reg/P0001 ,
		\u4_u2_int_stat_reg[0]/P0001 ,
		_w7248_
	);
	LUT3 #(
		.INIT('h08)
	) name5499 (
		\u1_u3_rx_ack_to_reg/P0001 ,
		\u1_u3_state_reg[3]/P0001 ,
		\u1_u3_state_reg[5]/P0001 ,
		_w7249_
	);
	LUT3 #(
		.INIT('h80)
	) name5500 (
		_w2127_,
		_w3699_,
		_w7249_,
		_w7250_
	);
	LUT2 #(
		.INIT('h4)
	) name5501 (
		\u1_u3_state_reg[2]/P0001 ,
		\u1_u3_tx_data_to_reg/P0001 ,
		_w7251_
	);
	LUT4 #(
		.INIT('h8000)
	) name5502 (
		\u1_u3_state_reg[4]/P0001 ,
		_w2127_,
		_w3676_,
		_w7251_,
		_w7252_
	);
	LUT3 #(
		.INIT('h08)
	) name5503 (
		rst_i_pad,
		\u4_u2_ep_match_r_reg/P0001 ,
		\u4_u2_int_re_reg/P0001 ,
		_w7253_
	);
	LUT4 #(
		.INIT('hfeaa)
	) name5504 (
		_w7248_,
		_w7250_,
		_w7252_,
		_w7253_,
		_w7254_
	);
	LUT3 #(
		.INIT('h40)
	) name5505 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_data_i[0]_pad ,
		_w7255_
	);
	LUT3 #(
		.INIT('h2a)
	) name5506 (
		rst_i_pad,
		_w2231_,
		_w7255_,
		_w7256_
	);
	LUT4 #(
		.INIT('hd8f0)
	) name5507 (
		\u1_u3_buf0_set_reg/P0001 ,
		\u1_u3_idin_reg[0]/P0001 ,
		\u4_u3_buf0_reg[0]/P0001 ,
		\u4_u3_ep_match_r_reg/P0001 ,
		_w7257_
	);
	LUT3 #(
		.INIT('hb8)
	) name5508 (
		\u4_u3_buf0_orig_reg[0]/P0001 ,
		_w2235_,
		_w7257_,
		_w7258_
	);
	LUT3 #(
		.INIT('h70)
	) name5509 (
		_w2231_,
		_w2232_,
		_w7258_,
		_w7259_
	);
	LUT2 #(
		.INIT('hd)
	) name5510 (
		_w7256_,
		_w7259_,
		_w7260_
	);
	LUT3 #(
		.INIT('h40)
	) name5511 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_data_i[12]_pad ,
		_w7261_
	);
	LUT3 #(
		.INIT('h2a)
	) name5512 (
		rst_i_pad,
		_w2231_,
		_w7261_,
		_w7262_
	);
	LUT4 #(
		.INIT('hd8f0)
	) name5513 (
		\u1_u3_buf0_set_reg/P0001 ,
		\u1_u3_idin_reg[12]/P0001 ,
		\u4_u3_buf0_reg[12]/P0001 ,
		\u4_u3_ep_match_r_reg/P0001 ,
		_w7263_
	);
	LUT3 #(
		.INIT('hb8)
	) name5514 (
		\u4_u3_buf0_orig_reg[12]/P0001 ,
		_w2235_,
		_w7263_,
		_w7264_
	);
	LUT3 #(
		.INIT('h70)
	) name5515 (
		_w2231_,
		_w2232_,
		_w7264_,
		_w7265_
	);
	LUT2 #(
		.INIT('hd)
	) name5516 (
		_w7262_,
		_w7265_,
		_w7266_
	);
	LUT3 #(
		.INIT('h40)
	) name5517 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_data_i[16]_pad ,
		_w7267_
	);
	LUT3 #(
		.INIT('h2a)
	) name5518 (
		rst_i_pad,
		_w2231_,
		_w7267_,
		_w7268_
	);
	LUT4 #(
		.INIT('hd8f0)
	) name5519 (
		\u1_u3_buf0_set_reg/P0001 ,
		\u1_u3_idin_reg[16]/P0001 ,
		\u4_u3_buf0_reg[16]/P0001 ,
		\u4_u3_ep_match_r_reg/P0001 ,
		_w7269_
	);
	LUT3 #(
		.INIT('hb8)
	) name5520 (
		\u4_u3_buf0_orig_reg[16]/P0001 ,
		_w2235_,
		_w7269_,
		_w7270_
	);
	LUT3 #(
		.INIT('h70)
	) name5521 (
		_w2231_,
		_w2232_,
		_w7270_,
		_w7271_
	);
	LUT2 #(
		.INIT('hd)
	) name5522 (
		_w7268_,
		_w7271_,
		_w7272_
	);
	LUT3 #(
		.INIT('h40)
	) name5523 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_data_i[17]_pad ,
		_w7273_
	);
	LUT3 #(
		.INIT('h2a)
	) name5524 (
		rst_i_pad,
		_w2231_,
		_w7273_,
		_w7274_
	);
	LUT4 #(
		.INIT('hd8f0)
	) name5525 (
		\u1_u3_buf0_set_reg/P0001 ,
		\u1_u3_idin_reg[17]/P0001 ,
		\u4_u3_buf0_reg[17]/P0001 ,
		\u4_u3_ep_match_r_reg/P0001 ,
		_w7275_
	);
	LUT3 #(
		.INIT('hb8)
	) name5526 (
		\u4_u3_buf0_orig_reg[17]/P0001 ,
		_w2235_,
		_w7275_,
		_w7276_
	);
	LUT3 #(
		.INIT('h70)
	) name5527 (
		_w2231_,
		_w2232_,
		_w7276_,
		_w7277_
	);
	LUT2 #(
		.INIT('hd)
	) name5528 (
		_w7274_,
		_w7277_,
		_w7278_
	);
	LUT3 #(
		.INIT('h40)
	) name5529 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_data_i[18]_pad ,
		_w7279_
	);
	LUT3 #(
		.INIT('h2a)
	) name5530 (
		rst_i_pad,
		_w2231_,
		_w7279_,
		_w7280_
	);
	LUT4 #(
		.INIT('hd8f0)
	) name5531 (
		\u1_u3_buf0_set_reg/P0001 ,
		\u1_u3_idin_reg[18]/P0001 ,
		\u4_u3_buf0_reg[18]/P0001 ,
		\u4_u3_ep_match_r_reg/P0001 ,
		_w7281_
	);
	LUT3 #(
		.INIT('hb8)
	) name5532 (
		\u4_u3_buf0_orig_reg[18]/P0001 ,
		_w2235_,
		_w7281_,
		_w7282_
	);
	LUT3 #(
		.INIT('h70)
	) name5533 (
		_w2231_,
		_w2232_,
		_w7282_,
		_w7283_
	);
	LUT2 #(
		.INIT('hd)
	) name5534 (
		_w7280_,
		_w7283_,
		_w7284_
	);
	LUT3 #(
		.INIT('h40)
	) name5535 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_data_i[19]_pad ,
		_w7285_
	);
	LUT3 #(
		.INIT('h2a)
	) name5536 (
		rst_i_pad,
		_w2231_,
		_w7285_,
		_w7286_
	);
	LUT4 #(
		.INIT('hd8f0)
	) name5537 (
		\u1_u3_buf0_set_reg/P0001 ,
		\u1_u3_idin_reg[19]/P0001 ,
		\u4_u3_buf0_reg[19]/P0001 ,
		\u4_u3_ep_match_r_reg/P0001 ,
		_w7287_
	);
	LUT3 #(
		.INIT('hb8)
	) name5538 (
		\u4_u3_buf0_orig_reg[19]/P0001 ,
		_w2235_,
		_w7287_,
		_w7288_
	);
	LUT3 #(
		.INIT('h70)
	) name5539 (
		_w2231_,
		_w2232_,
		_w7288_,
		_w7289_
	);
	LUT2 #(
		.INIT('hd)
	) name5540 (
		_w7286_,
		_w7289_,
		_w7290_
	);
	LUT3 #(
		.INIT('h40)
	) name5541 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_data_i[1]_pad ,
		_w7291_
	);
	LUT3 #(
		.INIT('h2a)
	) name5542 (
		rst_i_pad,
		_w2231_,
		_w7291_,
		_w7292_
	);
	LUT4 #(
		.INIT('hd8f0)
	) name5543 (
		\u1_u3_buf0_set_reg/P0001 ,
		\u1_u3_idin_reg[1]/P0001 ,
		\u4_u3_buf0_reg[1]/P0001 ,
		\u4_u3_ep_match_r_reg/P0001 ,
		_w7293_
	);
	LUT3 #(
		.INIT('hb8)
	) name5544 (
		\u4_u3_buf0_orig_reg[1]/P0001 ,
		_w2235_,
		_w7293_,
		_w7294_
	);
	LUT3 #(
		.INIT('h70)
	) name5545 (
		_w2231_,
		_w2232_,
		_w7294_,
		_w7295_
	);
	LUT2 #(
		.INIT('hd)
	) name5546 (
		_w7292_,
		_w7295_,
		_w7296_
	);
	LUT3 #(
		.INIT('h40)
	) name5547 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_data_i[20]_pad ,
		_w7297_
	);
	LUT3 #(
		.INIT('h2a)
	) name5548 (
		rst_i_pad,
		_w2231_,
		_w7297_,
		_w7298_
	);
	LUT4 #(
		.INIT('hd8f0)
	) name5549 (
		\u1_u3_buf0_set_reg/P0001 ,
		\u1_u3_idin_reg[20]/P0001 ,
		\u4_u3_buf0_reg[20]/P0001 ,
		\u4_u3_ep_match_r_reg/P0001 ,
		_w7299_
	);
	LUT3 #(
		.INIT('hb8)
	) name5550 (
		\u4_u3_buf0_orig_reg[20]/P0001 ,
		_w2235_,
		_w7299_,
		_w7300_
	);
	LUT3 #(
		.INIT('h70)
	) name5551 (
		_w2231_,
		_w2232_,
		_w7300_,
		_w7301_
	);
	LUT2 #(
		.INIT('hd)
	) name5552 (
		_w7298_,
		_w7301_,
		_w7302_
	);
	LUT3 #(
		.INIT('h40)
	) name5553 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_data_i[21]_pad ,
		_w7303_
	);
	LUT3 #(
		.INIT('h2a)
	) name5554 (
		rst_i_pad,
		_w2231_,
		_w7303_,
		_w7304_
	);
	LUT4 #(
		.INIT('hd8f0)
	) name5555 (
		\u1_u3_buf0_set_reg/P0001 ,
		\u1_u3_idin_reg[21]/P0001 ,
		\u4_u3_buf0_reg[21]/P0001 ,
		\u4_u3_ep_match_r_reg/P0001 ,
		_w7305_
	);
	LUT3 #(
		.INIT('hb8)
	) name5556 (
		\u4_u3_buf0_orig_reg[21]/P0001 ,
		_w2235_,
		_w7305_,
		_w7306_
	);
	LUT3 #(
		.INIT('h70)
	) name5557 (
		_w2231_,
		_w2232_,
		_w7306_,
		_w7307_
	);
	LUT2 #(
		.INIT('hd)
	) name5558 (
		_w7304_,
		_w7307_,
		_w7308_
	);
	LUT3 #(
		.INIT('h40)
	) name5559 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_data_i[22]_pad ,
		_w7309_
	);
	LUT3 #(
		.INIT('h2a)
	) name5560 (
		rst_i_pad,
		_w2231_,
		_w7309_,
		_w7310_
	);
	LUT4 #(
		.INIT('hd8f0)
	) name5561 (
		\u1_u3_buf0_set_reg/P0001 ,
		\u1_u3_idin_reg[22]/P0001 ,
		\u4_u3_buf0_reg[22]/P0001 ,
		\u4_u3_ep_match_r_reg/P0001 ,
		_w7311_
	);
	LUT3 #(
		.INIT('hb8)
	) name5562 (
		\u4_u3_buf0_orig_reg[22]/P0001 ,
		_w2235_,
		_w7311_,
		_w7312_
	);
	LUT3 #(
		.INIT('h70)
	) name5563 (
		_w2231_,
		_w2232_,
		_w7312_,
		_w7313_
	);
	LUT2 #(
		.INIT('hd)
	) name5564 (
		_w7310_,
		_w7313_,
		_w7314_
	);
	LUT3 #(
		.INIT('h40)
	) name5565 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_data_i[23]_pad ,
		_w7315_
	);
	LUT3 #(
		.INIT('h2a)
	) name5566 (
		rst_i_pad,
		_w2231_,
		_w7315_,
		_w7316_
	);
	LUT4 #(
		.INIT('hd8f0)
	) name5567 (
		\u1_u3_buf0_set_reg/P0001 ,
		\u1_u3_idin_reg[23]/P0001 ,
		\u4_u3_buf0_reg[23]/P0001 ,
		\u4_u3_ep_match_r_reg/P0001 ,
		_w7317_
	);
	LUT3 #(
		.INIT('hb8)
	) name5568 (
		\u4_u3_buf0_orig_reg[23]/P0001 ,
		_w2235_,
		_w7317_,
		_w7318_
	);
	LUT3 #(
		.INIT('h70)
	) name5569 (
		_w2231_,
		_w2232_,
		_w7318_,
		_w7319_
	);
	LUT2 #(
		.INIT('hd)
	) name5570 (
		_w7316_,
		_w7319_,
		_w7320_
	);
	LUT3 #(
		.INIT('h40)
	) name5571 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_data_i[24]_pad ,
		_w7321_
	);
	LUT3 #(
		.INIT('h2a)
	) name5572 (
		rst_i_pad,
		_w2231_,
		_w7321_,
		_w7322_
	);
	LUT4 #(
		.INIT('hd8f0)
	) name5573 (
		\u1_u3_buf0_set_reg/P0001 ,
		\u1_u3_idin_reg[24]/P0001 ,
		\u4_u3_buf0_reg[24]/P0001 ,
		\u4_u3_ep_match_r_reg/P0001 ,
		_w7323_
	);
	LUT3 #(
		.INIT('hb8)
	) name5574 (
		\u4_u3_buf0_orig_reg[24]/P0001 ,
		_w2235_,
		_w7323_,
		_w7324_
	);
	LUT3 #(
		.INIT('h70)
	) name5575 (
		_w2231_,
		_w2232_,
		_w7324_,
		_w7325_
	);
	LUT2 #(
		.INIT('hd)
	) name5576 (
		_w7322_,
		_w7325_,
		_w7326_
	);
	LUT3 #(
		.INIT('h40)
	) name5577 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_data_i[25]_pad ,
		_w7327_
	);
	LUT3 #(
		.INIT('h2a)
	) name5578 (
		rst_i_pad,
		_w2231_,
		_w7327_,
		_w7328_
	);
	LUT4 #(
		.INIT('hd8f0)
	) name5579 (
		\u1_u3_buf0_set_reg/P0001 ,
		\u1_u3_idin_reg[25]/P0001 ,
		\u4_u3_buf0_reg[25]/P0001 ,
		\u4_u3_ep_match_r_reg/P0001 ,
		_w7329_
	);
	LUT3 #(
		.INIT('hb8)
	) name5580 (
		\u4_u3_buf0_orig_reg[25]/P0001 ,
		_w2235_,
		_w7329_,
		_w7330_
	);
	LUT3 #(
		.INIT('h70)
	) name5581 (
		_w2231_,
		_w2232_,
		_w7330_,
		_w7331_
	);
	LUT2 #(
		.INIT('hd)
	) name5582 (
		_w7328_,
		_w7331_,
		_w7332_
	);
	LUT3 #(
		.INIT('h40)
	) name5583 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_data_i[26]_pad ,
		_w7333_
	);
	LUT3 #(
		.INIT('h2a)
	) name5584 (
		rst_i_pad,
		_w2231_,
		_w7333_,
		_w7334_
	);
	LUT4 #(
		.INIT('hd8f0)
	) name5585 (
		\u1_u3_buf0_set_reg/P0001 ,
		\u1_u3_idin_reg[26]/P0001 ,
		\u4_u3_buf0_reg[26]/P0001 ,
		\u4_u3_ep_match_r_reg/P0001 ,
		_w7335_
	);
	LUT3 #(
		.INIT('hb8)
	) name5586 (
		\u4_u3_buf0_orig_reg[26]/P0001 ,
		_w2235_,
		_w7335_,
		_w7336_
	);
	LUT3 #(
		.INIT('h70)
	) name5587 (
		_w2231_,
		_w2232_,
		_w7336_,
		_w7337_
	);
	LUT2 #(
		.INIT('hd)
	) name5588 (
		_w7334_,
		_w7337_,
		_w7338_
	);
	LUT3 #(
		.INIT('h40)
	) name5589 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_data_i[27]_pad ,
		_w7339_
	);
	LUT3 #(
		.INIT('h2a)
	) name5590 (
		rst_i_pad,
		_w2231_,
		_w7339_,
		_w7340_
	);
	LUT4 #(
		.INIT('hd8f0)
	) name5591 (
		\u1_u3_buf0_set_reg/P0001 ,
		\u1_u3_idin_reg[27]/P0001 ,
		\u4_u3_buf0_reg[27]/P0001 ,
		\u4_u3_ep_match_r_reg/P0001 ,
		_w7341_
	);
	LUT3 #(
		.INIT('hb8)
	) name5592 (
		\u4_u3_buf0_orig_reg[27]/P0001 ,
		_w2235_,
		_w7341_,
		_w7342_
	);
	LUT3 #(
		.INIT('h70)
	) name5593 (
		_w2231_,
		_w2232_,
		_w7342_,
		_w7343_
	);
	LUT2 #(
		.INIT('hd)
	) name5594 (
		_w7340_,
		_w7343_,
		_w7344_
	);
	LUT3 #(
		.INIT('h40)
	) name5595 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_data_i[28]_pad ,
		_w7345_
	);
	LUT3 #(
		.INIT('h2a)
	) name5596 (
		rst_i_pad,
		_w2231_,
		_w7345_,
		_w7346_
	);
	LUT4 #(
		.INIT('hd8f0)
	) name5597 (
		\u1_u3_buf0_set_reg/P0001 ,
		\u1_u3_idin_reg[28]/P0001 ,
		\u4_u3_buf0_reg[28]/P0001 ,
		\u4_u3_ep_match_r_reg/P0001 ,
		_w7347_
	);
	LUT3 #(
		.INIT('hb8)
	) name5598 (
		\u4_u3_buf0_orig_reg[28]/P0001 ,
		_w2235_,
		_w7347_,
		_w7348_
	);
	LUT3 #(
		.INIT('h70)
	) name5599 (
		_w2231_,
		_w2232_,
		_w7348_,
		_w7349_
	);
	LUT2 #(
		.INIT('hd)
	) name5600 (
		_w7346_,
		_w7349_,
		_w7350_
	);
	LUT3 #(
		.INIT('h40)
	) name5601 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_data_i[29]_pad ,
		_w7351_
	);
	LUT3 #(
		.INIT('h2a)
	) name5602 (
		rst_i_pad,
		_w2231_,
		_w7351_,
		_w7352_
	);
	LUT4 #(
		.INIT('hd8f0)
	) name5603 (
		\u1_u3_buf0_set_reg/P0001 ,
		\u1_u3_idin_reg[29]/P0001 ,
		\u4_u3_buf0_reg[29]/P0001 ,
		\u4_u3_ep_match_r_reg/P0001 ,
		_w7353_
	);
	LUT3 #(
		.INIT('hb8)
	) name5604 (
		\u4_u3_buf0_orig_reg[29]/NET0131 ,
		_w2235_,
		_w7353_,
		_w7354_
	);
	LUT3 #(
		.INIT('h70)
	) name5605 (
		_w2231_,
		_w2232_,
		_w7354_,
		_w7355_
	);
	LUT2 #(
		.INIT('hd)
	) name5606 (
		_w7352_,
		_w7355_,
		_w7356_
	);
	LUT3 #(
		.INIT('h40)
	) name5607 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_data_i[2]_pad ,
		_w7357_
	);
	LUT3 #(
		.INIT('h2a)
	) name5608 (
		rst_i_pad,
		_w2231_,
		_w7357_,
		_w7358_
	);
	LUT4 #(
		.INIT('hd8f0)
	) name5609 (
		\u1_u3_buf0_set_reg/P0001 ,
		\u1_u3_idin_reg[2]/P0001 ,
		\u4_u3_buf0_reg[2]/P0001 ,
		\u4_u3_ep_match_r_reg/P0001 ,
		_w7359_
	);
	LUT3 #(
		.INIT('hb8)
	) name5610 (
		\u4_u3_buf0_orig_reg[2]/P0001 ,
		_w2235_,
		_w7359_,
		_w7360_
	);
	LUT3 #(
		.INIT('h70)
	) name5611 (
		_w2231_,
		_w2232_,
		_w7360_,
		_w7361_
	);
	LUT2 #(
		.INIT('hd)
	) name5612 (
		_w7358_,
		_w7361_,
		_w7362_
	);
	LUT3 #(
		.INIT('h40)
	) name5613 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_data_i[30]_pad ,
		_w7363_
	);
	LUT3 #(
		.INIT('h2a)
	) name5614 (
		rst_i_pad,
		_w2231_,
		_w7363_,
		_w7364_
	);
	LUT4 #(
		.INIT('hd8f0)
	) name5615 (
		\u1_u3_buf0_set_reg/P0001 ,
		\u1_u3_idin_reg[30]/P0001 ,
		\u4_u3_buf0_reg[30]/P0001 ,
		\u4_u3_ep_match_r_reg/P0001 ,
		_w7365_
	);
	LUT3 #(
		.INIT('hb8)
	) name5616 (
		\u4_u3_buf0_orig_reg[30]/NET0131 ,
		_w2235_,
		_w7365_,
		_w7366_
	);
	LUT3 #(
		.INIT('h70)
	) name5617 (
		_w2231_,
		_w2232_,
		_w7366_,
		_w7367_
	);
	LUT2 #(
		.INIT('hd)
	) name5618 (
		_w7364_,
		_w7367_,
		_w7368_
	);
	LUT3 #(
		.INIT('h40)
	) name5619 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_data_i[31]_pad ,
		_w7369_
	);
	LUT3 #(
		.INIT('h2a)
	) name5620 (
		rst_i_pad,
		_w2231_,
		_w7369_,
		_w7370_
	);
	LUT4 #(
		.INIT('hd8f0)
	) name5621 (
		\u1_u3_buf0_set_reg/P0001 ,
		\u1_u3_idin_reg[31]/P0001 ,
		\u4_u3_buf0_reg[31]/P0001 ,
		\u4_u3_ep_match_r_reg/P0001 ,
		_w7371_
	);
	LUT3 #(
		.INIT('hb8)
	) name5622 (
		\u4_u3_buf0_orig_reg[31]/P0001 ,
		_w2235_,
		_w7371_,
		_w7372_
	);
	LUT3 #(
		.INIT('h70)
	) name5623 (
		_w2231_,
		_w2232_,
		_w7372_,
		_w7373_
	);
	LUT2 #(
		.INIT('hd)
	) name5624 (
		_w7370_,
		_w7373_,
		_w7374_
	);
	LUT3 #(
		.INIT('h40)
	) name5625 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_data_i[3]_pad ,
		_w7375_
	);
	LUT3 #(
		.INIT('h2a)
	) name5626 (
		rst_i_pad,
		_w2231_,
		_w7375_,
		_w7376_
	);
	LUT4 #(
		.INIT('hd8f0)
	) name5627 (
		\u1_u3_buf0_set_reg/P0001 ,
		\u1_u3_idin_reg[3]/P0001 ,
		\u4_u3_buf0_reg[3]/P0001 ,
		\u4_u3_ep_match_r_reg/P0001 ,
		_w7377_
	);
	LUT3 #(
		.INIT('hb8)
	) name5628 (
		\u4_u3_buf0_orig_reg[3]/P0001 ,
		_w2235_,
		_w7377_,
		_w7378_
	);
	LUT3 #(
		.INIT('h70)
	) name5629 (
		_w2231_,
		_w2232_,
		_w7378_,
		_w7379_
	);
	LUT2 #(
		.INIT('hd)
	) name5630 (
		_w7376_,
		_w7379_,
		_w7380_
	);
	LUT3 #(
		.INIT('h40)
	) name5631 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_data_i[8]_pad ,
		_w7381_
	);
	LUT3 #(
		.INIT('h2a)
	) name5632 (
		rst_i_pad,
		_w2231_,
		_w7381_,
		_w7382_
	);
	LUT4 #(
		.INIT('hd8f0)
	) name5633 (
		\u1_u3_buf0_set_reg/P0001 ,
		\u1_u3_idin_reg[8]/P0001 ,
		\u4_u3_buf0_reg[8]/P0001 ,
		\u4_u3_ep_match_r_reg/P0001 ,
		_w7383_
	);
	LUT3 #(
		.INIT('hb8)
	) name5634 (
		\u4_u3_buf0_orig_reg[8]/P0001 ,
		_w2235_,
		_w7383_,
		_w7384_
	);
	LUT3 #(
		.INIT('h70)
	) name5635 (
		_w2231_,
		_w2232_,
		_w7384_,
		_w7385_
	);
	LUT2 #(
		.INIT('hd)
	) name5636 (
		_w7382_,
		_w7385_,
		_w7386_
	);
	LUT3 #(
		.INIT('h40)
	) name5637 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_data_i[9]_pad ,
		_w7387_
	);
	LUT3 #(
		.INIT('h2a)
	) name5638 (
		rst_i_pad,
		_w2231_,
		_w7387_,
		_w7388_
	);
	LUT4 #(
		.INIT('hd8f0)
	) name5639 (
		\u1_u3_buf0_set_reg/P0001 ,
		\u1_u3_idin_reg[9]/P0001 ,
		\u4_u3_buf0_reg[9]/P0001 ,
		\u4_u3_ep_match_r_reg/P0001 ,
		_w7389_
	);
	LUT3 #(
		.INIT('hb8)
	) name5640 (
		\u4_u3_buf0_orig_reg[9]/P0001 ,
		_w2235_,
		_w7389_,
		_w7390_
	);
	LUT3 #(
		.INIT('h70)
	) name5641 (
		_w2231_,
		_w2232_,
		_w7390_,
		_w7391_
	);
	LUT2 #(
		.INIT('hd)
	) name5642 (
		_w7388_,
		_w7391_,
		_w7392_
	);
	LUT3 #(
		.INIT('h20)
	) name5643 (
		rst_i_pad,
		\u4_u3_int_re_reg/P0001 ,
		\u4_u3_int_stat_reg[0]/P0001 ,
		_w7393_
	);
	LUT3 #(
		.INIT('h08)
	) name5644 (
		rst_i_pad,
		\u4_u3_ep_match_r_reg/P0001 ,
		\u4_u3_int_re_reg/P0001 ,
		_w7394_
	);
	LUT4 #(
		.INIT('hfef0)
	) name5645 (
		_w7250_,
		_w7252_,
		_w7393_,
		_w7394_,
		_w7395_
	);
	LUT4 #(
		.INIT('h0010)
	) name5646 (
		\u1_u2_state_reg[0]/P0001 ,
		\u1_u2_state_reg[1]/NET0131 ,
		\u1_u2_state_reg[2]/NET0131 ,
		\u1_u2_state_reg[3]/NET0131 ,
		_w7396_
	);
	LUT3 #(
		.INIT('h80)
	) name5647 (
		_w3209_,
		_w6439_,
		_w7396_,
		_w7397_
	);
	LUT3 #(
		.INIT('h01)
	) name5648 (
		\u1_u2_wr_done_reg/P0001 ,
		\u1_u2_wr_last_reg/P0001 ,
		\u1_u3_abort_reg/P0001 ,
		_w7398_
	);
	LUT3 #(
		.INIT('h80)
	) name5649 (
		_w3209_,
		_w3214_,
		_w7398_,
		_w7399_
	);
	LUT3 #(
		.INIT('ha8)
	) name5650 (
		rst_i_pad,
		_w7397_,
		_w7399_,
		_w7400_
	);
	LUT3 #(
		.INIT('h2a)
	) name5651 (
		rst_i_pad,
		_w2243_,
		_w7255_,
		_w7401_
	);
	LUT4 #(
		.INIT('hd8f0)
	) name5652 (
		\u1_u3_buf0_set_reg/P0001 ,
		\u1_u3_idin_reg[0]/P0001 ,
		\u4_u0_buf0_reg[0]/P0001 ,
		\u4_u0_ep_match_r_reg/P0001 ,
		_w7402_
	);
	LUT3 #(
		.INIT('hb8)
	) name5653 (
		\u4_u0_buf0_orig_reg[0]/P0001 ,
		_w2245_,
		_w7402_,
		_w7403_
	);
	LUT3 #(
		.INIT('h70)
	) name5654 (
		_w2232_,
		_w2243_,
		_w7403_,
		_w7404_
	);
	LUT2 #(
		.INIT('hd)
	) name5655 (
		_w7401_,
		_w7404_,
		_w7405_
	);
	LUT3 #(
		.INIT('h2a)
	) name5656 (
		rst_i_pad,
		_w2243_,
		_w7261_,
		_w7406_
	);
	LUT4 #(
		.INIT('hd8f0)
	) name5657 (
		\u1_u3_buf0_set_reg/P0001 ,
		\u1_u3_idin_reg[12]/P0001 ,
		\u4_u0_buf0_reg[12]/P0001 ,
		\u4_u0_ep_match_r_reg/P0001 ,
		_w7407_
	);
	LUT3 #(
		.INIT('hb8)
	) name5658 (
		\u4_u0_buf0_orig_reg[12]/P0001 ,
		_w2245_,
		_w7407_,
		_w7408_
	);
	LUT3 #(
		.INIT('h70)
	) name5659 (
		_w2232_,
		_w2243_,
		_w7408_,
		_w7409_
	);
	LUT2 #(
		.INIT('hd)
	) name5660 (
		_w7406_,
		_w7409_,
		_w7410_
	);
	LUT3 #(
		.INIT('h2a)
	) name5661 (
		rst_i_pad,
		_w2243_,
		_w7267_,
		_w7411_
	);
	LUT4 #(
		.INIT('hd8f0)
	) name5662 (
		\u1_u3_buf0_set_reg/P0001 ,
		\u1_u3_idin_reg[16]/P0001 ,
		\u4_u0_buf0_reg[16]/P0001 ,
		\u4_u0_ep_match_r_reg/P0001 ,
		_w7412_
	);
	LUT3 #(
		.INIT('hb8)
	) name5663 (
		\u4_u0_buf0_orig_reg[16]/P0001 ,
		_w2245_,
		_w7412_,
		_w7413_
	);
	LUT3 #(
		.INIT('h70)
	) name5664 (
		_w2232_,
		_w2243_,
		_w7413_,
		_w7414_
	);
	LUT2 #(
		.INIT('hd)
	) name5665 (
		_w7411_,
		_w7414_,
		_w7415_
	);
	LUT3 #(
		.INIT('h2a)
	) name5666 (
		rst_i_pad,
		_w2243_,
		_w7273_,
		_w7416_
	);
	LUT4 #(
		.INIT('hd8f0)
	) name5667 (
		\u1_u3_buf0_set_reg/P0001 ,
		\u1_u3_idin_reg[17]/P0001 ,
		\u4_u0_buf0_reg[17]/P0001 ,
		\u4_u0_ep_match_r_reg/P0001 ,
		_w7417_
	);
	LUT3 #(
		.INIT('hb8)
	) name5668 (
		\u4_u0_buf0_orig_reg[17]/P0001 ,
		_w2245_,
		_w7417_,
		_w7418_
	);
	LUT3 #(
		.INIT('h70)
	) name5669 (
		_w2232_,
		_w2243_,
		_w7418_,
		_w7419_
	);
	LUT2 #(
		.INIT('hd)
	) name5670 (
		_w7416_,
		_w7419_,
		_w7420_
	);
	LUT3 #(
		.INIT('h2a)
	) name5671 (
		rst_i_pad,
		_w2243_,
		_w7279_,
		_w7421_
	);
	LUT4 #(
		.INIT('hd8f0)
	) name5672 (
		\u1_u3_buf0_set_reg/P0001 ,
		\u1_u3_idin_reg[18]/P0001 ,
		\u4_u0_buf0_reg[18]/P0001 ,
		\u4_u0_ep_match_r_reg/P0001 ,
		_w7422_
	);
	LUT3 #(
		.INIT('hb8)
	) name5673 (
		\u4_u0_buf0_orig_reg[18]/P0001 ,
		_w2245_,
		_w7422_,
		_w7423_
	);
	LUT3 #(
		.INIT('h70)
	) name5674 (
		_w2232_,
		_w2243_,
		_w7423_,
		_w7424_
	);
	LUT2 #(
		.INIT('hd)
	) name5675 (
		_w7421_,
		_w7424_,
		_w7425_
	);
	LUT3 #(
		.INIT('h2a)
	) name5676 (
		rst_i_pad,
		_w2243_,
		_w7285_,
		_w7426_
	);
	LUT4 #(
		.INIT('hd8f0)
	) name5677 (
		\u1_u3_buf0_set_reg/P0001 ,
		\u1_u3_idin_reg[19]/P0001 ,
		\u4_u0_buf0_reg[19]/P0001 ,
		\u4_u0_ep_match_r_reg/P0001 ,
		_w7427_
	);
	LUT3 #(
		.INIT('hb8)
	) name5678 (
		\u4_u0_buf0_orig_reg[19]/P0001 ,
		_w2245_,
		_w7427_,
		_w7428_
	);
	LUT3 #(
		.INIT('h70)
	) name5679 (
		_w2232_,
		_w2243_,
		_w7428_,
		_w7429_
	);
	LUT2 #(
		.INIT('hd)
	) name5680 (
		_w7426_,
		_w7429_,
		_w7430_
	);
	LUT3 #(
		.INIT('h2a)
	) name5681 (
		rst_i_pad,
		_w2243_,
		_w7291_,
		_w7431_
	);
	LUT4 #(
		.INIT('hd8f0)
	) name5682 (
		\u1_u3_buf0_set_reg/P0001 ,
		\u1_u3_idin_reg[1]/P0001 ,
		\u4_u0_buf0_reg[1]/P0001 ,
		\u4_u0_ep_match_r_reg/P0001 ,
		_w7432_
	);
	LUT3 #(
		.INIT('hb8)
	) name5683 (
		\u4_u0_buf0_orig_reg[1]/P0001 ,
		_w2245_,
		_w7432_,
		_w7433_
	);
	LUT3 #(
		.INIT('h70)
	) name5684 (
		_w2232_,
		_w2243_,
		_w7433_,
		_w7434_
	);
	LUT2 #(
		.INIT('hd)
	) name5685 (
		_w7431_,
		_w7434_,
		_w7435_
	);
	LUT3 #(
		.INIT('h2a)
	) name5686 (
		rst_i_pad,
		_w2243_,
		_w7297_,
		_w7436_
	);
	LUT4 #(
		.INIT('hd8f0)
	) name5687 (
		\u1_u3_buf0_set_reg/P0001 ,
		\u1_u3_idin_reg[20]/P0001 ,
		\u4_u0_buf0_reg[20]/P0001 ,
		\u4_u0_ep_match_r_reg/P0001 ,
		_w7437_
	);
	LUT3 #(
		.INIT('hb8)
	) name5688 (
		\u4_u0_buf0_orig_reg[20]/P0001 ,
		_w2245_,
		_w7437_,
		_w7438_
	);
	LUT3 #(
		.INIT('h70)
	) name5689 (
		_w2232_,
		_w2243_,
		_w7438_,
		_w7439_
	);
	LUT2 #(
		.INIT('hd)
	) name5690 (
		_w7436_,
		_w7439_,
		_w7440_
	);
	LUT3 #(
		.INIT('h2a)
	) name5691 (
		rst_i_pad,
		_w2243_,
		_w7303_,
		_w7441_
	);
	LUT4 #(
		.INIT('hd8f0)
	) name5692 (
		\u1_u3_buf0_set_reg/P0001 ,
		\u1_u3_idin_reg[21]/P0001 ,
		\u4_u0_buf0_reg[21]/P0001 ,
		\u4_u0_ep_match_r_reg/P0001 ,
		_w7442_
	);
	LUT3 #(
		.INIT('hb8)
	) name5693 (
		\u4_u0_buf0_orig_reg[21]/P0001 ,
		_w2245_,
		_w7442_,
		_w7443_
	);
	LUT3 #(
		.INIT('h70)
	) name5694 (
		_w2232_,
		_w2243_,
		_w7443_,
		_w7444_
	);
	LUT2 #(
		.INIT('hd)
	) name5695 (
		_w7441_,
		_w7444_,
		_w7445_
	);
	LUT3 #(
		.INIT('h2a)
	) name5696 (
		rst_i_pad,
		_w2243_,
		_w7309_,
		_w7446_
	);
	LUT4 #(
		.INIT('hd8f0)
	) name5697 (
		\u1_u3_buf0_set_reg/P0001 ,
		\u1_u3_idin_reg[22]/P0001 ,
		\u4_u0_buf0_reg[22]/P0001 ,
		\u4_u0_ep_match_r_reg/P0001 ,
		_w7447_
	);
	LUT3 #(
		.INIT('hb8)
	) name5698 (
		\u4_u0_buf0_orig_reg[22]/P0001 ,
		_w2245_,
		_w7447_,
		_w7448_
	);
	LUT3 #(
		.INIT('h70)
	) name5699 (
		_w2232_,
		_w2243_,
		_w7448_,
		_w7449_
	);
	LUT2 #(
		.INIT('hd)
	) name5700 (
		_w7446_,
		_w7449_,
		_w7450_
	);
	LUT3 #(
		.INIT('h2a)
	) name5701 (
		rst_i_pad,
		_w2243_,
		_w7315_,
		_w7451_
	);
	LUT4 #(
		.INIT('hd8f0)
	) name5702 (
		\u1_u3_buf0_set_reg/P0001 ,
		\u1_u3_idin_reg[23]/P0001 ,
		\u4_u0_buf0_reg[23]/P0001 ,
		\u4_u0_ep_match_r_reg/P0001 ,
		_w7452_
	);
	LUT3 #(
		.INIT('hb8)
	) name5703 (
		\u4_u0_buf0_orig_reg[23]/P0001 ,
		_w2245_,
		_w7452_,
		_w7453_
	);
	LUT3 #(
		.INIT('h70)
	) name5704 (
		_w2232_,
		_w2243_,
		_w7453_,
		_w7454_
	);
	LUT2 #(
		.INIT('hd)
	) name5705 (
		_w7451_,
		_w7454_,
		_w7455_
	);
	LUT3 #(
		.INIT('h2a)
	) name5706 (
		rst_i_pad,
		_w2243_,
		_w7321_,
		_w7456_
	);
	LUT4 #(
		.INIT('hd8f0)
	) name5707 (
		\u1_u3_buf0_set_reg/P0001 ,
		\u1_u3_idin_reg[24]/P0001 ,
		\u4_u0_buf0_reg[24]/P0001 ,
		\u4_u0_ep_match_r_reg/P0001 ,
		_w7457_
	);
	LUT3 #(
		.INIT('hb8)
	) name5708 (
		\u4_u0_buf0_orig_reg[24]/P0001 ,
		_w2245_,
		_w7457_,
		_w7458_
	);
	LUT3 #(
		.INIT('h70)
	) name5709 (
		_w2232_,
		_w2243_,
		_w7458_,
		_w7459_
	);
	LUT2 #(
		.INIT('hd)
	) name5710 (
		_w7456_,
		_w7459_,
		_w7460_
	);
	LUT3 #(
		.INIT('h2a)
	) name5711 (
		rst_i_pad,
		_w2243_,
		_w7327_,
		_w7461_
	);
	LUT4 #(
		.INIT('hd8f0)
	) name5712 (
		\u1_u3_buf0_set_reg/P0001 ,
		\u1_u3_idin_reg[25]/P0001 ,
		\u4_u0_buf0_reg[25]/P0001 ,
		\u4_u0_ep_match_r_reg/P0001 ,
		_w7462_
	);
	LUT3 #(
		.INIT('hb8)
	) name5713 (
		\u4_u0_buf0_orig_reg[25]/P0001 ,
		_w2245_,
		_w7462_,
		_w7463_
	);
	LUT3 #(
		.INIT('h70)
	) name5714 (
		_w2232_,
		_w2243_,
		_w7463_,
		_w7464_
	);
	LUT2 #(
		.INIT('hd)
	) name5715 (
		_w7461_,
		_w7464_,
		_w7465_
	);
	LUT3 #(
		.INIT('h2a)
	) name5716 (
		rst_i_pad,
		_w2243_,
		_w7333_,
		_w7466_
	);
	LUT4 #(
		.INIT('hd8f0)
	) name5717 (
		\u1_u3_buf0_set_reg/P0001 ,
		\u1_u3_idin_reg[26]/P0001 ,
		\u4_u0_buf0_reg[26]/P0001 ,
		\u4_u0_ep_match_r_reg/P0001 ,
		_w7467_
	);
	LUT3 #(
		.INIT('hb8)
	) name5718 (
		\u4_u0_buf0_orig_reg[26]/P0001 ,
		_w2245_,
		_w7467_,
		_w7468_
	);
	LUT3 #(
		.INIT('h70)
	) name5719 (
		_w2232_,
		_w2243_,
		_w7468_,
		_w7469_
	);
	LUT2 #(
		.INIT('hd)
	) name5720 (
		_w7466_,
		_w7469_,
		_w7470_
	);
	LUT3 #(
		.INIT('h2a)
	) name5721 (
		rst_i_pad,
		_w2243_,
		_w7339_,
		_w7471_
	);
	LUT4 #(
		.INIT('hd8f0)
	) name5722 (
		\u1_u3_buf0_set_reg/P0001 ,
		\u1_u3_idin_reg[27]/P0001 ,
		\u4_u0_buf0_reg[27]/P0001 ,
		\u4_u0_ep_match_r_reg/P0001 ,
		_w7472_
	);
	LUT3 #(
		.INIT('hb8)
	) name5723 (
		\u4_u0_buf0_orig_reg[27]/P0001 ,
		_w2245_,
		_w7472_,
		_w7473_
	);
	LUT3 #(
		.INIT('h70)
	) name5724 (
		_w2232_,
		_w2243_,
		_w7473_,
		_w7474_
	);
	LUT2 #(
		.INIT('hd)
	) name5725 (
		_w7471_,
		_w7474_,
		_w7475_
	);
	LUT3 #(
		.INIT('h2a)
	) name5726 (
		rst_i_pad,
		_w2243_,
		_w7345_,
		_w7476_
	);
	LUT4 #(
		.INIT('hd8f0)
	) name5727 (
		\u1_u3_buf0_set_reg/P0001 ,
		\u1_u3_idin_reg[28]/P0001 ,
		\u4_u0_buf0_reg[28]/P0001 ,
		\u4_u0_ep_match_r_reg/P0001 ,
		_w7477_
	);
	LUT3 #(
		.INIT('hb8)
	) name5728 (
		\u4_u0_buf0_orig_reg[28]/P0001 ,
		_w2245_,
		_w7477_,
		_w7478_
	);
	LUT3 #(
		.INIT('h70)
	) name5729 (
		_w2232_,
		_w2243_,
		_w7478_,
		_w7479_
	);
	LUT2 #(
		.INIT('hd)
	) name5730 (
		_w7476_,
		_w7479_,
		_w7480_
	);
	LUT3 #(
		.INIT('h2a)
	) name5731 (
		rst_i_pad,
		_w2243_,
		_w7351_,
		_w7481_
	);
	LUT4 #(
		.INIT('hd8f0)
	) name5732 (
		\u1_u3_buf0_set_reg/P0001 ,
		\u1_u3_idin_reg[29]/P0001 ,
		\u4_u0_buf0_reg[29]/P0001 ,
		\u4_u0_ep_match_r_reg/P0001 ,
		_w7482_
	);
	LUT3 #(
		.INIT('hb8)
	) name5733 (
		\u4_u0_buf0_orig_reg[29]/NET0131 ,
		_w2245_,
		_w7482_,
		_w7483_
	);
	LUT3 #(
		.INIT('h70)
	) name5734 (
		_w2232_,
		_w2243_,
		_w7483_,
		_w7484_
	);
	LUT2 #(
		.INIT('hd)
	) name5735 (
		_w7481_,
		_w7484_,
		_w7485_
	);
	LUT3 #(
		.INIT('h2a)
	) name5736 (
		rst_i_pad,
		_w2243_,
		_w7357_,
		_w7486_
	);
	LUT4 #(
		.INIT('hd8f0)
	) name5737 (
		\u1_u3_buf0_set_reg/P0001 ,
		\u1_u3_idin_reg[2]/P0001 ,
		\u4_u0_buf0_reg[2]/P0001 ,
		\u4_u0_ep_match_r_reg/P0001 ,
		_w7487_
	);
	LUT3 #(
		.INIT('hb8)
	) name5738 (
		\u4_u0_buf0_orig_reg[2]/P0001 ,
		_w2245_,
		_w7487_,
		_w7488_
	);
	LUT3 #(
		.INIT('h70)
	) name5739 (
		_w2232_,
		_w2243_,
		_w7488_,
		_w7489_
	);
	LUT2 #(
		.INIT('hd)
	) name5740 (
		_w7486_,
		_w7489_,
		_w7490_
	);
	LUT3 #(
		.INIT('h2a)
	) name5741 (
		rst_i_pad,
		_w2243_,
		_w7363_,
		_w7491_
	);
	LUT4 #(
		.INIT('hd8f0)
	) name5742 (
		\u1_u3_buf0_set_reg/P0001 ,
		\u1_u3_idin_reg[30]/P0001 ,
		\u4_u0_buf0_reg[30]/P0001 ,
		\u4_u0_ep_match_r_reg/P0001 ,
		_w7492_
	);
	LUT3 #(
		.INIT('hb8)
	) name5743 (
		\u4_u0_buf0_orig_reg[30]/NET0131 ,
		_w2245_,
		_w7492_,
		_w7493_
	);
	LUT3 #(
		.INIT('h70)
	) name5744 (
		_w2232_,
		_w2243_,
		_w7493_,
		_w7494_
	);
	LUT2 #(
		.INIT('hd)
	) name5745 (
		_w7491_,
		_w7494_,
		_w7495_
	);
	LUT3 #(
		.INIT('h2a)
	) name5746 (
		rst_i_pad,
		_w2243_,
		_w7369_,
		_w7496_
	);
	LUT4 #(
		.INIT('hd8f0)
	) name5747 (
		\u1_u3_buf0_set_reg/P0001 ,
		\u1_u3_idin_reg[31]/P0001 ,
		\u4_u0_buf0_reg[31]/P0001 ,
		\u4_u0_ep_match_r_reg/P0001 ,
		_w7497_
	);
	LUT3 #(
		.INIT('hb8)
	) name5748 (
		\u4_u0_buf0_orig_reg[31]/P0001 ,
		_w2245_,
		_w7497_,
		_w7498_
	);
	LUT3 #(
		.INIT('h70)
	) name5749 (
		_w2232_,
		_w2243_,
		_w7498_,
		_w7499_
	);
	LUT2 #(
		.INIT('hd)
	) name5750 (
		_w7496_,
		_w7499_,
		_w7500_
	);
	LUT3 #(
		.INIT('h2a)
	) name5751 (
		rst_i_pad,
		_w2243_,
		_w7375_,
		_w7501_
	);
	LUT4 #(
		.INIT('hd8f0)
	) name5752 (
		\u1_u3_buf0_set_reg/P0001 ,
		\u1_u3_idin_reg[3]/P0001 ,
		\u4_u0_buf0_reg[3]/P0001 ,
		\u4_u0_ep_match_r_reg/P0001 ,
		_w7502_
	);
	LUT3 #(
		.INIT('hb8)
	) name5753 (
		\u4_u0_buf0_orig_reg[3]/P0001 ,
		_w2245_,
		_w7502_,
		_w7503_
	);
	LUT3 #(
		.INIT('h70)
	) name5754 (
		_w2232_,
		_w2243_,
		_w7503_,
		_w7504_
	);
	LUT2 #(
		.INIT('hd)
	) name5755 (
		_w7501_,
		_w7504_,
		_w7505_
	);
	LUT3 #(
		.INIT('h2a)
	) name5756 (
		rst_i_pad,
		_w2243_,
		_w7381_,
		_w7506_
	);
	LUT4 #(
		.INIT('hd8f0)
	) name5757 (
		\u1_u3_buf0_set_reg/P0001 ,
		\u1_u3_idin_reg[8]/P0001 ,
		\u4_u0_buf0_reg[8]/P0001 ,
		\u4_u0_ep_match_r_reg/P0001 ,
		_w7507_
	);
	LUT3 #(
		.INIT('hb8)
	) name5758 (
		\u4_u0_buf0_orig_reg[8]/P0001 ,
		_w2245_,
		_w7507_,
		_w7508_
	);
	LUT3 #(
		.INIT('h70)
	) name5759 (
		_w2232_,
		_w2243_,
		_w7508_,
		_w7509_
	);
	LUT2 #(
		.INIT('hd)
	) name5760 (
		_w7506_,
		_w7509_,
		_w7510_
	);
	LUT3 #(
		.INIT('h2a)
	) name5761 (
		rst_i_pad,
		_w2243_,
		_w7387_,
		_w7511_
	);
	LUT4 #(
		.INIT('hd8f0)
	) name5762 (
		\u1_u3_buf0_set_reg/P0001 ,
		\u1_u3_idin_reg[9]/P0001 ,
		\u4_u0_buf0_reg[9]/P0001 ,
		\u4_u0_ep_match_r_reg/P0001 ,
		_w7512_
	);
	LUT3 #(
		.INIT('hb8)
	) name5763 (
		\u4_u0_buf0_orig_reg[9]/P0001 ,
		_w2245_,
		_w7512_,
		_w7513_
	);
	LUT3 #(
		.INIT('h70)
	) name5764 (
		_w2232_,
		_w2243_,
		_w7513_,
		_w7514_
	);
	LUT2 #(
		.INIT('hd)
	) name5765 (
		_w7511_,
		_w7514_,
		_w7515_
	);
	LUT3 #(
		.INIT('h10)
	) name5766 (
		\u0_u0_T1_gt_5_0_mS_reg/P0001 ,
		\u0_u0_idle_cnt1_next_reg[3]/P0001 ,
		\u0_u0_ps_cnt_clr_reg/P0001 ,
		_w7516_
	);
	LUT3 #(
		.INIT('h23)
	) name5767 (
		\u0_u0_T1_gt_5_0_mS_reg/P0001 ,
		\u0_u0_idle_cnt1_reg[3]/P0001 ,
		\u0_u0_ps_cnt_clr_reg/P0001 ,
		_w7517_
	);
	LUT3 #(
		.INIT('h02)
	) name5768 (
		_w5770_,
		_w7516_,
		_w7517_,
		_w7518_
	);
	LUT3 #(
		.INIT('hd0)
	) name5769 (
		_w5763_,
		_w5768_,
		_w7518_,
		_w7519_
	);
	LUT2 #(
		.INIT('h4)
	) name5770 (
		_w5765_,
		_w7519_,
		_w7520_
	);
	LUT3 #(
		.INIT('h20)
	) name5771 (
		rst_i_pad,
		\u4_u0_int_re_reg/P0001 ,
		\u4_u0_int_stat_reg[0]/P0001 ,
		_w7521_
	);
	LUT3 #(
		.INIT('h08)
	) name5772 (
		rst_i_pad,
		\u4_u0_ep_match_r_reg/P0001 ,
		\u4_u0_int_re_reg/P0001 ,
		_w7522_
	);
	LUT4 #(
		.INIT('hfef0)
	) name5773 (
		_w7250_,
		_w7252_,
		_w7521_,
		_w7522_,
		_w7523_
	);
	LUT3 #(
		.INIT('h2a)
	) name5774 (
		rst_i_pad,
		_w2260_,
		_w7255_,
		_w7524_
	);
	LUT4 #(
		.INIT('hd8f0)
	) name5775 (
		\u1_u3_buf0_set_reg/P0001 ,
		\u1_u3_idin_reg[0]/P0001 ,
		\u4_u1_buf0_reg[0]/P0001 ,
		\u4_u1_ep_match_r_reg/P0001 ,
		_w7525_
	);
	LUT3 #(
		.INIT('hb8)
	) name5776 (
		\u4_u1_buf0_orig_reg[0]/P0001 ,
		_w2262_,
		_w7525_,
		_w7526_
	);
	LUT3 #(
		.INIT('h70)
	) name5777 (
		_w2232_,
		_w2260_,
		_w7526_,
		_w7527_
	);
	LUT2 #(
		.INIT('hd)
	) name5778 (
		_w7524_,
		_w7527_,
		_w7528_
	);
	LUT3 #(
		.INIT('h2a)
	) name5779 (
		rst_i_pad,
		_w2260_,
		_w7261_,
		_w7529_
	);
	LUT4 #(
		.INIT('hd8f0)
	) name5780 (
		\u1_u3_buf0_set_reg/P0001 ,
		\u1_u3_idin_reg[12]/P0001 ,
		\u4_u1_buf0_reg[12]/P0001 ,
		\u4_u1_ep_match_r_reg/P0001 ,
		_w7530_
	);
	LUT3 #(
		.INIT('hb8)
	) name5781 (
		\u4_u1_buf0_orig_reg[12]/P0001 ,
		_w2262_,
		_w7530_,
		_w7531_
	);
	LUT3 #(
		.INIT('h70)
	) name5782 (
		_w2232_,
		_w2260_,
		_w7531_,
		_w7532_
	);
	LUT2 #(
		.INIT('hd)
	) name5783 (
		_w7529_,
		_w7532_,
		_w7533_
	);
	LUT3 #(
		.INIT('h2a)
	) name5784 (
		rst_i_pad,
		_w2260_,
		_w7267_,
		_w7534_
	);
	LUT4 #(
		.INIT('hd8f0)
	) name5785 (
		\u1_u3_buf0_set_reg/P0001 ,
		\u1_u3_idin_reg[16]/P0001 ,
		\u4_u1_buf0_reg[16]/P0001 ,
		\u4_u1_ep_match_r_reg/P0001 ,
		_w7535_
	);
	LUT3 #(
		.INIT('hb8)
	) name5786 (
		\u4_u1_buf0_orig_reg[16]/P0001 ,
		_w2262_,
		_w7535_,
		_w7536_
	);
	LUT3 #(
		.INIT('h70)
	) name5787 (
		_w2232_,
		_w2260_,
		_w7536_,
		_w7537_
	);
	LUT2 #(
		.INIT('hd)
	) name5788 (
		_w7534_,
		_w7537_,
		_w7538_
	);
	LUT3 #(
		.INIT('h2a)
	) name5789 (
		rst_i_pad,
		_w2260_,
		_w7273_,
		_w7539_
	);
	LUT4 #(
		.INIT('hd8f0)
	) name5790 (
		\u1_u3_buf0_set_reg/P0001 ,
		\u1_u3_idin_reg[17]/P0001 ,
		\u4_u1_buf0_reg[17]/P0001 ,
		\u4_u1_ep_match_r_reg/P0001 ,
		_w7540_
	);
	LUT3 #(
		.INIT('hb8)
	) name5791 (
		\u4_u1_buf0_orig_reg[17]/P0001 ,
		_w2262_,
		_w7540_,
		_w7541_
	);
	LUT3 #(
		.INIT('h70)
	) name5792 (
		_w2232_,
		_w2260_,
		_w7541_,
		_w7542_
	);
	LUT2 #(
		.INIT('hd)
	) name5793 (
		_w7539_,
		_w7542_,
		_w7543_
	);
	LUT3 #(
		.INIT('h2a)
	) name5794 (
		rst_i_pad,
		_w2260_,
		_w7279_,
		_w7544_
	);
	LUT4 #(
		.INIT('hd8f0)
	) name5795 (
		\u1_u3_buf0_set_reg/P0001 ,
		\u1_u3_idin_reg[18]/P0001 ,
		\u4_u1_buf0_reg[18]/P0001 ,
		\u4_u1_ep_match_r_reg/P0001 ,
		_w7545_
	);
	LUT3 #(
		.INIT('hb8)
	) name5796 (
		\u4_u1_buf0_orig_reg[18]/P0001 ,
		_w2262_,
		_w7545_,
		_w7546_
	);
	LUT3 #(
		.INIT('h70)
	) name5797 (
		_w2232_,
		_w2260_,
		_w7546_,
		_w7547_
	);
	LUT2 #(
		.INIT('hd)
	) name5798 (
		_w7544_,
		_w7547_,
		_w7548_
	);
	LUT3 #(
		.INIT('h2a)
	) name5799 (
		rst_i_pad,
		_w2260_,
		_w7285_,
		_w7549_
	);
	LUT4 #(
		.INIT('hd8f0)
	) name5800 (
		\u1_u3_buf0_set_reg/P0001 ,
		\u1_u3_idin_reg[19]/P0001 ,
		\u4_u1_buf0_reg[19]/P0001 ,
		\u4_u1_ep_match_r_reg/P0001 ,
		_w7550_
	);
	LUT3 #(
		.INIT('hb8)
	) name5801 (
		\u4_u1_buf0_orig_reg[19]/P0001 ,
		_w2262_,
		_w7550_,
		_w7551_
	);
	LUT3 #(
		.INIT('h70)
	) name5802 (
		_w2232_,
		_w2260_,
		_w7551_,
		_w7552_
	);
	LUT2 #(
		.INIT('hd)
	) name5803 (
		_w7549_,
		_w7552_,
		_w7553_
	);
	LUT3 #(
		.INIT('h2a)
	) name5804 (
		rst_i_pad,
		_w2260_,
		_w7291_,
		_w7554_
	);
	LUT4 #(
		.INIT('hd8f0)
	) name5805 (
		\u1_u3_buf0_set_reg/P0001 ,
		\u1_u3_idin_reg[1]/P0001 ,
		\u4_u1_buf0_reg[1]/P0001 ,
		\u4_u1_ep_match_r_reg/P0001 ,
		_w7555_
	);
	LUT3 #(
		.INIT('hb8)
	) name5806 (
		\u4_u1_buf0_orig_reg[1]/P0001 ,
		_w2262_,
		_w7555_,
		_w7556_
	);
	LUT3 #(
		.INIT('h70)
	) name5807 (
		_w2232_,
		_w2260_,
		_w7556_,
		_w7557_
	);
	LUT2 #(
		.INIT('hd)
	) name5808 (
		_w7554_,
		_w7557_,
		_w7558_
	);
	LUT3 #(
		.INIT('h2a)
	) name5809 (
		rst_i_pad,
		_w2260_,
		_w7297_,
		_w7559_
	);
	LUT4 #(
		.INIT('hd8f0)
	) name5810 (
		\u1_u3_buf0_set_reg/P0001 ,
		\u1_u3_idin_reg[20]/P0001 ,
		\u4_u1_buf0_reg[20]/P0001 ,
		\u4_u1_ep_match_r_reg/P0001 ,
		_w7560_
	);
	LUT3 #(
		.INIT('hb8)
	) name5811 (
		\u4_u1_buf0_orig_reg[20]/P0001 ,
		_w2262_,
		_w7560_,
		_w7561_
	);
	LUT3 #(
		.INIT('h70)
	) name5812 (
		_w2232_,
		_w2260_,
		_w7561_,
		_w7562_
	);
	LUT2 #(
		.INIT('hd)
	) name5813 (
		_w7559_,
		_w7562_,
		_w7563_
	);
	LUT3 #(
		.INIT('h2a)
	) name5814 (
		rst_i_pad,
		_w2260_,
		_w7303_,
		_w7564_
	);
	LUT4 #(
		.INIT('hd8f0)
	) name5815 (
		\u1_u3_buf0_set_reg/P0001 ,
		\u1_u3_idin_reg[21]/P0001 ,
		\u4_u1_buf0_reg[21]/P0001 ,
		\u4_u1_ep_match_r_reg/P0001 ,
		_w7565_
	);
	LUT3 #(
		.INIT('hb8)
	) name5816 (
		\u4_u1_buf0_orig_reg[21]/P0001 ,
		_w2262_,
		_w7565_,
		_w7566_
	);
	LUT3 #(
		.INIT('h70)
	) name5817 (
		_w2232_,
		_w2260_,
		_w7566_,
		_w7567_
	);
	LUT2 #(
		.INIT('hd)
	) name5818 (
		_w7564_,
		_w7567_,
		_w7568_
	);
	LUT3 #(
		.INIT('h2a)
	) name5819 (
		rst_i_pad,
		_w2260_,
		_w7309_,
		_w7569_
	);
	LUT4 #(
		.INIT('hd8f0)
	) name5820 (
		\u1_u3_buf0_set_reg/P0001 ,
		\u1_u3_idin_reg[22]/P0001 ,
		\u4_u1_buf0_reg[22]/P0001 ,
		\u4_u1_ep_match_r_reg/P0001 ,
		_w7570_
	);
	LUT3 #(
		.INIT('hb8)
	) name5821 (
		\u4_u1_buf0_orig_reg[22]/P0001 ,
		_w2262_,
		_w7570_,
		_w7571_
	);
	LUT3 #(
		.INIT('h70)
	) name5822 (
		_w2232_,
		_w2260_,
		_w7571_,
		_w7572_
	);
	LUT2 #(
		.INIT('hd)
	) name5823 (
		_w7569_,
		_w7572_,
		_w7573_
	);
	LUT3 #(
		.INIT('h2a)
	) name5824 (
		rst_i_pad,
		_w2260_,
		_w7315_,
		_w7574_
	);
	LUT4 #(
		.INIT('hd8f0)
	) name5825 (
		\u1_u3_buf0_set_reg/P0001 ,
		\u1_u3_idin_reg[23]/P0001 ,
		\u4_u1_buf0_reg[23]/P0001 ,
		\u4_u1_ep_match_r_reg/P0001 ,
		_w7575_
	);
	LUT3 #(
		.INIT('hb8)
	) name5826 (
		\u4_u1_buf0_orig_reg[23]/P0001 ,
		_w2262_,
		_w7575_,
		_w7576_
	);
	LUT3 #(
		.INIT('h70)
	) name5827 (
		_w2232_,
		_w2260_,
		_w7576_,
		_w7577_
	);
	LUT2 #(
		.INIT('hd)
	) name5828 (
		_w7574_,
		_w7577_,
		_w7578_
	);
	LUT3 #(
		.INIT('h2a)
	) name5829 (
		rst_i_pad,
		_w2260_,
		_w7321_,
		_w7579_
	);
	LUT4 #(
		.INIT('hd8f0)
	) name5830 (
		\u1_u3_buf0_set_reg/P0001 ,
		\u1_u3_idin_reg[24]/P0001 ,
		\u4_u1_buf0_reg[24]/P0001 ,
		\u4_u1_ep_match_r_reg/P0001 ,
		_w7580_
	);
	LUT3 #(
		.INIT('hb8)
	) name5831 (
		\u4_u1_buf0_orig_reg[24]/P0001 ,
		_w2262_,
		_w7580_,
		_w7581_
	);
	LUT3 #(
		.INIT('h70)
	) name5832 (
		_w2232_,
		_w2260_,
		_w7581_,
		_w7582_
	);
	LUT2 #(
		.INIT('hd)
	) name5833 (
		_w7579_,
		_w7582_,
		_w7583_
	);
	LUT3 #(
		.INIT('h2a)
	) name5834 (
		rst_i_pad,
		_w2260_,
		_w7327_,
		_w7584_
	);
	LUT4 #(
		.INIT('hd8f0)
	) name5835 (
		\u1_u3_buf0_set_reg/P0001 ,
		\u1_u3_idin_reg[25]/P0001 ,
		\u4_u1_buf0_reg[25]/P0001 ,
		\u4_u1_ep_match_r_reg/P0001 ,
		_w7585_
	);
	LUT3 #(
		.INIT('hb8)
	) name5836 (
		\u4_u1_buf0_orig_reg[25]/P0001 ,
		_w2262_,
		_w7585_,
		_w7586_
	);
	LUT3 #(
		.INIT('h70)
	) name5837 (
		_w2232_,
		_w2260_,
		_w7586_,
		_w7587_
	);
	LUT2 #(
		.INIT('hd)
	) name5838 (
		_w7584_,
		_w7587_,
		_w7588_
	);
	LUT3 #(
		.INIT('h2a)
	) name5839 (
		rst_i_pad,
		_w2260_,
		_w7333_,
		_w7589_
	);
	LUT4 #(
		.INIT('hd8f0)
	) name5840 (
		\u1_u3_buf0_set_reg/P0001 ,
		\u1_u3_idin_reg[26]/P0001 ,
		\u4_u1_buf0_reg[26]/P0001 ,
		\u4_u1_ep_match_r_reg/P0001 ,
		_w7590_
	);
	LUT3 #(
		.INIT('hb8)
	) name5841 (
		\u4_u1_buf0_orig_reg[26]/P0001 ,
		_w2262_,
		_w7590_,
		_w7591_
	);
	LUT3 #(
		.INIT('h70)
	) name5842 (
		_w2232_,
		_w2260_,
		_w7591_,
		_w7592_
	);
	LUT2 #(
		.INIT('hd)
	) name5843 (
		_w7589_,
		_w7592_,
		_w7593_
	);
	LUT3 #(
		.INIT('h2a)
	) name5844 (
		rst_i_pad,
		_w2260_,
		_w7339_,
		_w7594_
	);
	LUT4 #(
		.INIT('hd8f0)
	) name5845 (
		\u1_u3_buf0_set_reg/P0001 ,
		\u1_u3_idin_reg[27]/P0001 ,
		\u4_u1_buf0_reg[27]/P0001 ,
		\u4_u1_ep_match_r_reg/P0001 ,
		_w7595_
	);
	LUT3 #(
		.INIT('hb8)
	) name5846 (
		\u4_u1_buf0_orig_reg[27]/P0001 ,
		_w2262_,
		_w7595_,
		_w7596_
	);
	LUT3 #(
		.INIT('h70)
	) name5847 (
		_w2232_,
		_w2260_,
		_w7596_,
		_w7597_
	);
	LUT2 #(
		.INIT('hd)
	) name5848 (
		_w7594_,
		_w7597_,
		_w7598_
	);
	LUT3 #(
		.INIT('h2a)
	) name5849 (
		rst_i_pad,
		_w2260_,
		_w7345_,
		_w7599_
	);
	LUT4 #(
		.INIT('hd8f0)
	) name5850 (
		\u1_u3_buf0_set_reg/P0001 ,
		\u1_u3_idin_reg[28]/P0001 ,
		\u4_u1_buf0_reg[28]/P0001 ,
		\u4_u1_ep_match_r_reg/P0001 ,
		_w7600_
	);
	LUT3 #(
		.INIT('hb8)
	) name5851 (
		\u4_u1_buf0_orig_reg[28]/P0001 ,
		_w2262_,
		_w7600_,
		_w7601_
	);
	LUT3 #(
		.INIT('h70)
	) name5852 (
		_w2232_,
		_w2260_,
		_w7601_,
		_w7602_
	);
	LUT2 #(
		.INIT('hd)
	) name5853 (
		_w7599_,
		_w7602_,
		_w7603_
	);
	LUT3 #(
		.INIT('h2a)
	) name5854 (
		rst_i_pad,
		_w2260_,
		_w7351_,
		_w7604_
	);
	LUT4 #(
		.INIT('hd8f0)
	) name5855 (
		\u1_u3_buf0_set_reg/P0001 ,
		\u1_u3_idin_reg[29]/P0001 ,
		\u4_u1_buf0_reg[29]/P0001 ,
		\u4_u1_ep_match_r_reg/P0001 ,
		_w7605_
	);
	LUT3 #(
		.INIT('hb8)
	) name5856 (
		\u4_u1_buf0_orig_reg[29]/NET0131 ,
		_w2262_,
		_w7605_,
		_w7606_
	);
	LUT3 #(
		.INIT('h70)
	) name5857 (
		_w2232_,
		_w2260_,
		_w7606_,
		_w7607_
	);
	LUT2 #(
		.INIT('hd)
	) name5858 (
		_w7604_,
		_w7607_,
		_w7608_
	);
	LUT3 #(
		.INIT('h2a)
	) name5859 (
		rst_i_pad,
		_w2260_,
		_w7357_,
		_w7609_
	);
	LUT4 #(
		.INIT('hd8f0)
	) name5860 (
		\u1_u3_buf0_set_reg/P0001 ,
		\u1_u3_idin_reg[2]/P0001 ,
		\u4_u1_buf0_reg[2]/P0001 ,
		\u4_u1_ep_match_r_reg/P0001 ,
		_w7610_
	);
	LUT3 #(
		.INIT('hb8)
	) name5861 (
		\u4_u1_buf0_orig_reg[2]/P0001 ,
		_w2262_,
		_w7610_,
		_w7611_
	);
	LUT3 #(
		.INIT('h70)
	) name5862 (
		_w2232_,
		_w2260_,
		_w7611_,
		_w7612_
	);
	LUT2 #(
		.INIT('hd)
	) name5863 (
		_w7609_,
		_w7612_,
		_w7613_
	);
	LUT3 #(
		.INIT('h2a)
	) name5864 (
		rst_i_pad,
		_w2260_,
		_w7363_,
		_w7614_
	);
	LUT4 #(
		.INIT('hd8f0)
	) name5865 (
		\u1_u3_buf0_set_reg/P0001 ,
		\u1_u3_idin_reg[30]/P0001 ,
		\u4_u1_buf0_reg[30]/P0001 ,
		\u4_u1_ep_match_r_reg/P0001 ,
		_w7615_
	);
	LUT3 #(
		.INIT('hb8)
	) name5866 (
		\u4_u1_buf0_orig_reg[30]/NET0131 ,
		_w2262_,
		_w7615_,
		_w7616_
	);
	LUT3 #(
		.INIT('h70)
	) name5867 (
		_w2232_,
		_w2260_,
		_w7616_,
		_w7617_
	);
	LUT2 #(
		.INIT('hd)
	) name5868 (
		_w7614_,
		_w7617_,
		_w7618_
	);
	LUT3 #(
		.INIT('h2a)
	) name5869 (
		rst_i_pad,
		_w2260_,
		_w7369_,
		_w7619_
	);
	LUT4 #(
		.INIT('hd8f0)
	) name5870 (
		\u1_u3_buf0_set_reg/P0001 ,
		\u1_u3_idin_reg[31]/P0001 ,
		\u4_u1_buf0_reg[31]/P0001 ,
		\u4_u1_ep_match_r_reg/P0001 ,
		_w7620_
	);
	LUT3 #(
		.INIT('hb8)
	) name5871 (
		\u4_u1_buf0_orig_reg[31]/P0001 ,
		_w2262_,
		_w7620_,
		_w7621_
	);
	LUT3 #(
		.INIT('h70)
	) name5872 (
		_w2232_,
		_w2260_,
		_w7621_,
		_w7622_
	);
	LUT2 #(
		.INIT('hd)
	) name5873 (
		_w7619_,
		_w7622_,
		_w7623_
	);
	LUT3 #(
		.INIT('h2a)
	) name5874 (
		rst_i_pad,
		_w2260_,
		_w7375_,
		_w7624_
	);
	LUT4 #(
		.INIT('hd8f0)
	) name5875 (
		\u1_u3_buf0_set_reg/P0001 ,
		\u1_u3_idin_reg[3]/P0001 ,
		\u4_u1_buf0_reg[3]/P0001 ,
		\u4_u1_ep_match_r_reg/P0001 ,
		_w7625_
	);
	LUT3 #(
		.INIT('hb8)
	) name5876 (
		\u4_u1_buf0_orig_reg[3]/P0001 ,
		_w2262_,
		_w7625_,
		_w7626_
	);
	LUT3 #(
		.INIT('h70)
	) name5877 (
		_w2232_,
		_w2260_,
		_w7626_,
		_w7627_
	);
	LUT2 #(
		.INIT('hd)
	) name5878 (
		_w7624_,
		_w7627_,
		_w7628_
	);
	LUT3 #(
		.INIT('h2a)
	) name5879 (
		rst_i_pad,
		_w2260_,
		_w7381_,
		_w7629_
	);
	LUT4 #(
		.INIT('hd8f0)
	) name5880 (
		\u1_u3_buf0_set_reg/P0001 ,
		\u1_u3_idin_reg[8]/P0001 ,
		\u4_u1_buf0_reg[8]/P0001 ,
		\u4_u1_ep_match_r_reg/P0001 ,
		_w7630_
	);
	LUT3 #(
		.INIT('hb8)
	) name5881 (
		\u4_u1_buf0_orig_reg[8]/P0001 ,
		_w2262_,
		_w7630_,
		_w7631_
	);
	LUT3 #(
		.INIT('h70)
	) name5882 (
		_w2232_,
		_w2260_,
		_w7631_,
		_w7632_
	);
	LUT2 #(
		.INIT('hd)
	) name5883 (
		_w7629_,
		_w7632_,
		_w7633_
	);
	LUT3 #(
		.INIT('h2a)
	) name5884 (
		rst_i_pad,
		_w2260_,
		_w7387_,
		_w7634_
	);
	LUT4 #(
		.INIT('hd8f0)
	) name5885 (
		\u1_u3_buf0_set_reg/P0001 ,
		\u1_u3_idin_reg[9]/P0001 ,
		\u4_u1_buf0_reg[9]/P0001 ,
		\u4_u1_ep_match_r_reg/P0001 ,
		_w7635_
	);
	LUT3 #(
		.INIT('hb8)
	) name5886 (
		\u4_u1_buf0_orig_reg[9]/P0001 ,
		_w2262_,
		_w7635_,
		_w7636_
	);
	LUT3 #(
		.INIT('h70)
	) name5887 (
		_w2232_,
		_w2260_,
		_w7636_,
		_w7637_
	);
	LUT2 #(
		.INIT('hd)
	) name5888 (
		_w7634_,
		_w7637_,
		_w7638_
	);
	LUT3 #(
		.INIT('h20)
	) name5889 (
		rst_i_pad,
		\u4_u1_int_re_reg/P0001 ,
		\u4_u1_int_stat_reg[0]/P0001 ,
		_w7639_
	);
	LUT3 #(
		.INIT('h08)
	) name5890 (
		rst_i_pad,
		\u4_u1_ep_match_r_reg/P0001 ,
		\u4_u1_int_re_reg/P0001 ,
		_w7640_
	);
	LUT4 #(
		.INIT('hfef0)
	) name5891 (
		_w7250_,
		_w7252_,
		_w7639_,
		_w7640_,
		_w7641_
	);
	LUT3 #(
		.INIT('h2a)
	) name5892 (
		rst_i_pad,
		_w2267_,
		_w7255_,
		_w7642_
	);
	LUT4 #(
		.INIT('hd8f0)
	) name5893 (
		\u1_u3_buf0_set_reg/P0001 ,
		\u1_u3_idin_reg[0]/P0001 ,
		\u4_u2_buf0_reg[0]/P0001 ,
		\u4_u2_ep_match_r_reg/P0001 ,
		_w7643_
	);
	LUT3 #(
		.INIT('hb8)
	) name5894 (
		\u4_u2_buf0_orig_reg[0]/P0001 ,
		_w2269_,
		_w7643_,
		_w7644_
	);
	LUT3 #(
		.INIT('h70)
	) name5895 (
		_w2232_,
		_w2267_,
		_w7644_,
		_w7645_
	);
	LUT2 #(
		.INIT('hd)
	) name5896 (
		_w7642_,
		_w7645_,
		_w7646_
	);
	LUT3 #(
		.INIT('h2a)
	) name5897 (
		rst_i_pad,
		_w2267_,
		_w7261_,
		_w7647_
	);
	LUT4 #(
		.INIT('hd8f0)
	) name5898 (
		\u1_u3_buf0_set_reg/P0001 ,
		\u1_u3_idin_reg[12]/P0001 ,
		\u4_u2_buf0_reg[12]/P0001 ,
		\u4_u2_ep_match_r_reg/P0001 ,
		_w7648_
	);
	LUT3 #(
		.INIT('hb8)
	) name5899 (
		\u4_u2_buf0_orig_reg[12]/P0001 ,
		_w2269_,
		_w7648_,
		_w7649_
	);
	LUT3 #(
		.INIT('h70)
	) name5900 (
		_w2232_,
		_w2267_,
		_w7649_,
		_w7650_
	);
	LUT2 #(
		.INIT('hd)
	) name5901 (
		_w7647_,
		_w7650_,
		_w7651_
	);
	LUT3 #(
		.INIT('h2a)
	) name5902 (
		rst_i_pad,
		_w2267_,
		_w7267_,
		_w7652_
	);
	LUT4 #(
		.INIT('hd8f0)
	) name5903 (
		\u1_u3_buf0_set_reg/P0001 ,
		\u1_u3_idin_reg[16]/P0001 ,
		\u4_u2_buf0_reg[16]/P0001 ,
		\u4_u2_ep_match_r_reg/P0001 ,
		_w7653_
	);
	LUT3 #(
		.INIT('hb8)
	) name5904 (
		\u4_u2_buf0_orig_reg[16]/P0001 ,
		_w2269_,
		_w7653_,
		_w7654_
	);
	LUT3 #(
		.INIT('h70)
	) name5905 (
		_w2232_,
		_w2267_,
		_w7654_,
		_w7655_
	);
	LUT2 #(
		.INIT('hd)
	) name5906 (
		_w7652_,
		_w7655_,
		_w7656_
	);
	LUT3 #(
		.INIT('h2a)
	) name5907 (
		rst_i_pad,
		_w2267_,
		_w7273_,
		_w7657_
	);
	LUT4 #(
		.INIT('hd8f0)
	) name5908 (
		\u1_u3_buf0_set_reg/P0001 ,
		\u1_u3_idin_reg[17]/P0001 ,
		\u4_u2_buf0_reg[17]/P0001 ,
		\u4_u2_ep_match_r_reg/P0001 ,
		_w7658_
	);
	LUT3 #(
		.INIT('hb8)
	) name5909 (
		\u4_u2_buf0_orig_reg[17]/P0001 ,
		_w2269_,
		_w7658_,
		_w7659_
	);
	LUT3 #(
		.INIT('h70)
	) name5910 (
		_w2232_,
		_w2267_,
		_w7659_,
		_w7660_
	);
	LUT2 #(
		.INIT('hd)
	) name5911 (
		_w7657_,
		_w7660_,
		_w7661_
	);
	LUT3 #(
		.INIT('h2a)
	) name5912 (
		rst_i_pad,
		_w2267_,
		_w7279_,
		_w7662_
	);
	LUT4 #(
		.INIT('hd8f0)
	) name5913 (
		\u1_u3_buf0_set_reg/P0001 ,
		\u1_u3_idin_reg[18]/P0001 ,
		\u4_u2_buf0_reg[18]/P0001 ,
		\u4_u2_ep_match_r_reg/P0001 ,
		_w7663_
	);
	LUT3 #(
		.INIT('hb8)
	) name5914 (
		\u4_u2_buf0_orig_reg[18]/P0001 ,
		_w2269_,
		_w7663_,
		_w7664_
	);
	LUT3 #(
		.INIT('h70)
	) name5915 (
		_w2232_,
		_w2267_,
		_w7664_,
		_w7665_
	);
	LUT2 #(
		.INIT('hd)
	) name5916 (
		_w7662_,
		_w7665_,
		_w7666_
	);
	LUT3 #(
		.INIT('h2a)
	) name5917 (
		rst_i_pad,
		_w2267_,
		_w7285_,
		_w7667_
	);
	LUT4 #(
		.INIT('hd8f0)
	) name5918 (
		\u1_u3_buf0_set_reg/P0001 ,
		\u1_u3_idin_reg[19]/P0001 ,
		\u4_u2_buf0_reg[19]/P0001 ,
		\u4_u2_ep_match_r_reg/P0001 ,
		_w7668_
	);
	LUT3 #(
		.INIT('hb8)
	) name5919 (
		\u4_u2_buf0_orig_reg[19]/P0001 ,
		_w2269_,
		_w7668_,
		_w7669_
	);
	LUT3 #(
		.INIT('h70)
	) name5920 (
		_w2232_,
		_w2267_,
		_w7669_,
		_w7670_
	);
	LUT2 #(
		.INIT('hd)
	) name5921 (
		_w7667_,
		_w7670_,
		_w7671_
	);
	LUT3 #(
		.INIT('h2a)
	) name5922 (
		rst_i_pad,
		_w2267_,
		_w7291_,
		_w7672_
	);
	LUT4 #(
		.INIT('hd8f0)
	) name5923 (
		\u1_u3_buf0_set_reg/P0001 ,
		\u1_u3_idin_reg[1]/P0001 ,
		\u4_u2_buf0_reg[1]/P0001 ,
		\u4_u2_ep_match_r_reg/P0001 ,
		_w7673_
	);
	LUT3 #(
		.INIT('hb8)
	) name5924 (
		\u4_u2_buf0_orig_reg[1]/P0001 ,
		_w2269_,
		_w7673_,
		_w7674_
	);
	LUT3 #(
		.INIT('h70)
	) name5925 (
		_w2232_,
		_w2267_,
		_w7674_,
		_w7675_
	);
	LUT2 #(
		.INIT('hd)
	) name5926 (
		_w7672_,
		_w7675_,
		_w7676_
	);
	LUT3 #(
		.INIT('h2a)
	) name5927 (
		rst_i_pad,
		_w2267_,
		_w7297_,
		_w7677_
	);
	LUT4 #(
		.INIT('hd8f0)
	) name5928 (
		\u1_u3_buf0_set_reg/P0001 ,
		\u1_u3_idin_reg[20]/P0001 ,
		\u4_u2_buf0_reg[20]/P0001 ,
		\u4_u2_ep_match_r_reg/P0001 ,
		_w7678_
	);
	LUT3 #(
		.INIT('hb8)
	) name5929 (
		\u4_u2_buf0_orig_reg[20]/P0001 ,
		_w2269_,
		_w7678_,
		_w7679_
	);
	LUT3 #(
		.INIT('h70)
	) name5930 (
		_w2232_,
		_w2267_,
		_w7679_,
		_w7680_
	);
	LUT2 #(
		.INIT('hd)
	) name5931 (
		_w7677_,
		_w7680_,
		_w7681_
	);
	LUT3 #(
		.INIT('h2a)
	) name5932 (
		rst_i_pad,
		_w2267_,
		_w7303_,
		_w7682_
	);
	LUT4 #(
		.INIT('hd8f0)
	) name5933 (
		\u1_u3_buf0_set_reg/P0001 ,
		\u1_u3_idin_reg[21]/P0001 ,
		\u4_u2_buf0_reg[21]/P0001 ,
		\u4_u2_ep_match_r_reg/P0001 ,
		_w7683_
	);
	LUT3 #(
		.INIT('hb8)
	) name5934 (
		\u4_u2_buf0_orig_reg[21]/P0001 ,
		_w2269_,
		_w7683_,
		_w7684_
	);
	LUT3 #(
		.INIT('h70)
	) name5935 (
		_w2232_,
		_w2267_,
		_w7684_,
		_w7685_
	);
	LUT2 #(
		.INIT('hd)
	) name5936 (
		_w7682_,
		_w7685_,
		_w7686_
	);
	LUT3 #(
		.INIT('h2a)
	) name5937 (
		rst_i_pad,
		_w2267_,
		_w7309_,
		_w7687_
	);
	LUT4 #(
		.INIT('hd8f0)
	) name5938 (
		\u1_u3_buf0_set_reg/P0001 ,
		\u1_u3_idin_reg[22]/P0001 ,
		\u4_u2_buf0_reg[22]/P0001 ,
		\u4_u2_ep_match_r_reg/P0001 ,
		_w7688_
	);
	LUT3 #(
		.INIT('hb8)
	) name5939 (
		\u4_u2_buf0_orig_reg[22]/P0001 ,
		_w2269_,
		_w7688_,
		_w7689_
	);
	LUT3 #(
		.INIT('h70)
	) name5940 (
		_w2232_,
		_w2267_,
		_w7689_,
		_w7690_
	);
	LUT2 #(
		.INIT('hd)
	) name5941 (
		_w7687_,
		_w7690_,
		_w7691_
	);
	LUT3 #(
		.INIT('h2a)
	) name5942 (
		rst_i_pad,
		_w2267_,
		_w7315_,
		_w7692_
	);
	LUT4 #(
		.INIT('hd8f0)
	) name5943 (
		\u1_u3_buf0_set_reg/P0001 ,
		\u1_u3_idin_reg[23]/P0001 ,
		\u4_u2_buf0_reg[23]/P0001 ,
		\u4_u2_ep_match_r_reg/P0001 ,
		_w7693_
	);
	LUT3 #(
		.INIT('hb8)
	) name5944 (
		\u4_u2_buf0_orig_reg[23]/P0001 ,
		_w2269_,
		_w7693_,
		_w7694_
	);
	LUT3 #(
		.INIT('h70)
	) name5945 (
		_w2232_,
		_w2267_,
		_w7694_,
		_w7695_
	);
	LUT2 #(
		.INIT('hd)
	) name5946 (
		_w7692_,
		_w7695_,
		_w7696_
	);
	LUT3 #(
		.INIT('h2a)
	) name5947 (
		rst_i_pad,
		_w2267_,
		_w7321_,
		_w7697_
	);
	LUT4 #(
		.INIT('hd8f0)
	) name5948 (
		\u1_u3_buf0_set_reg/P0001 ,
		\u1_u3_idin_reg[24]/P0001 ,
		\u4_u2_buf0_reg[24]/P0001 ,
		\u4_u2_ep_match_r_reg/P0001 ,
		_w7698_
	);
	LUT3 #(
		.INIT('hb8)
	) name5949 (
		\u4_u2_buf0_orig_reg[24]/P0001 ,
		_w2269_,
		_w7698_,
		_w7699_
	);
	LUT3 #(
		.INIT('h70)
	) name5950 (
		_w2232_,
		_w2267_,
		_w7699_,
		_w7700_
	);
	LUT2 #(
		.INIT('hd)
	) name5951 (
		_w7697_,
		_w7700_,
		_w7701_
	);
	LUT3 #(
		.INIT('h2a)
	) name5952 (
		rst_i_pad,
		_w2267_,
		_w7327_,
		_w7702_
	);
	LUT4 #(
		.INIT('hd8f0)
	) name5953 (
		\u1_u3_buf0_set_reg/P0001 ,
		\u1_u3_idin_reg[25]/P0001 ,
		\u4_u2_buf0_reg[25]/P0001 ,
		\u4_u2_ep_match_r_reg/P0001 ,
		_w7703_
	);
	LUT3 #(
		.INIT('hb8)
	) name5954 (
		\u4_u2_buf0_orig_reg[25]/P0001 ,
		_w2269_,
		_w7703_,
		_w7704_
	);
	LUT3 #(
		.INIT('h70)
	) name5955 (
		_w2232_,
		_w2267_,
		_w7704_,
		_w7705_
	);
	LUT2 #(
		.INIT('hd)
	) name5956 (
		_w7702_,
		_w7705_,
		_w7706_
	);
	LUT3 #(
		.INIT('h2a)
	) name5957 (
		rst_i_pad,
		_w2267_,
		_w7333_,
		_w7707_
	);
	LUT4 #(
		.INIT('hd8f0)
	) name5958 (
		\u1_u3_buf0_set_reg/P0001 ,
		\u1_u3_idin_reg[26]/P0001 ,
		\u4_u2_buf0_reg[26]/P0001 ,
		\u4_u2_ep_match_r_reg/P0001 ,
		_w7708_
	);
	LUT3 #(
		.INIT('hb8)
	) name5959 (
		\u4_u2_buf0_orig_reg[26]/P0001 ,
		_w2269_,
		_w7708_,
		_w7709_
	);
	LUT3 #(
		.INIT('h70)
	) name5960 (
		_w2232_,
		_w2267_,
		_w7709_,
		_w7710_
	);
	LUT2 #(
		.INIT('hd)
	) name5961 (
		_w7707_,
		_w7710_,
		_w7711_
	);
	LUT3 #(
		.INIT('h2a)
	) name5962 (
		rst_i_pad,
		_w2267_,
		_w7339_,
		_w7712_
	);
	LUT4 #(
		.INIT('hd8f0)
	) name5963 (
		\u1_u3_buf0_set_reg/P0001 ,
		\u1_u3_idin_reg[27]/P0001 ,
		\u4_u2_buf0_reg[27]/P0001 ,
		\u4_u2_ep_match_r_reg/P0001 ,
		_w7713_
	);
	LUT3 #(
		.INIT('hb8)
	) name5964 (
		\u4_u2_buf0_orig_reg[27]/P0001 ,
		_w2269_,
		_w7713_,
		_w7714_
	);
	LUT3 #(
		.INIT('h70)
	) name5965 (
		_w2232_,
		_w2267_,
		_w7714_,
		_w7715_
	);
	LUT2 #(
		.INIT('hd)
	) name5966 (
		_w7712_,
		_w7715_,
		_w7716_
	);
	LUT3 #(
		.INIT('h2a)
	) name5967 (
		rst_i_pad,
		_w2267_,
		_w7345_,
		_w7717_
	);
	LUT4 #(
		.INIT('hd8f0)
	) name5968 (
		\u1_u3_buf0_set_reg/P0001 ,
		\u1_u3_idin_reg[28]/P0001 ,
		\u4_u2_buf0_reg[28]/P0001 ,
		\u4_u2_ep_match_r_reg/P0001 ,
		_w7718_
	);
	LUT3 #(
		.INIT('hb8)
	) name5969 (
		\u4_u2_buf0_orig_reg[28]/P0001 ,
		_w2269_,
		_w7718_,
		_w7719_
	);
	LUT3 #(
		.INIT('h70)
	) name5970 (
		_w2232_,
		_w2267_,
		_w7719_,
		_w7720_
	);
	LUT2 #(
		.INIT('hd)
	) name5971 (
		_w7717_,
		_w7720_,
		_w7721_
	);
	LUT3 #(
		.INIT('h2a)
	) name5972 (
		rst_i_pad,
		_w2267_,
		_w7351_,
		_w7722_
	);
	LUT4 #(
		.INIT('hd8f0)
	) name5973 (
		\u1_u3_buf0_set_reg/P0001 ,
		\u1_u3_idin_reg[29]/P0001 ,
		\u4_u2_buf0_reg[29]/P0001 ,
		\u4_u2_ep_match_r_reg/P0001 ,
		_w7723_
	);
	LUT3 #(
		.INIT('hb8)
	) name5974 (
		\u4_u2_buf0_orig_reg[29]/NET0131 ,
		_w2269_,
		_w7723_,
		_w7724_
	);
	LUT3 #(
		.INIT('h70)
	) name5975 (
		_w2232_,
		_w2267_,
		_w7724_,
		_w7725_
	);
	LUT2 #(
		.INIT('hd)
	) name5976 (
		_w7722_,
		_w7725_,
		_w7726_
	);
	LUT3 #(
		.INIT('h2a)
	) name5977 (
		rst_i_pad,
		_w2267_,
		_w7357_,
		_w7727_
	);
	LUT4 #(
		.INIT('hd8f0)
	) name5978 (
		\u1_u3_buf0_set_reg/P0001 ,
		\u1_u3_idin_reg[2]/P0001 ,
		\u4_u2_buf0_reg[2]/P0001 ,
		\u4_u2_ep_match_r_reg/P0001 ,
		_w7728_
	);
	LUT3 #(
		.INIT('hb8)
	) name5979 (
		\u4_u2_buf0_orig_reg[2]/P0001 ,
		_w2269_,
		_w7728_,
		_w7729_
	);
	LUT3 #(
		.INIT('h70)
	) name5980 (
		_w2232_,
		_w2267_,
		_w7729_,
		_w7730_
	);
	LUT2 #(
		.INIT('hd)
	) name5981 (
		_w7727_,
		_w7730_,
		_w7731_
	);
	LUT3 #(
		.INIT('h2a)
	) name5982 (
		rst_i_pad,
		_w2267_,
		_w7363_,
		_w7732_
	);
	LUT4 #(
		.INIT('hd8f0)
	) name5983 (
		\u1_u3_buf0_set_reg/P0001 ,
		\u1_u3_idin_reg[30]/P0001 ,
		\u4_u2_buf0_reg[30]/P0001 ,
		\u4_u2_ep_match_r_reg/P0001 ,
		_w7733_
	);
	LUT3 #(
		.INIT('hb8)
	) name5984 (
		\u4_u2_buf0_orig_reg[30]/NET0131 ,
		_w2269_,
		_w7733_,
		_w7734_
	);
	LUT3 #(
		.INIT('h70)
	) name5985 (
		_w2232_,
		_w2267_,
		_w7734_,
		_w7735_
	);
	LUT2 #(
		.INIT('hd)
	) name5986 (
		_w7732_,
		_w7735_,
		_w7736_
	);
	LUT3 #(
		.INIT('h2a)
	) name5987 (
		rst_i_pad,
		_w2267_,
		_w7369_,
		_w7737_
	);
	LUT4 #(
		.INIT('hd8f0)
	) name5988 (
		\u1_u3_buf0_set_reg/P0001 ,
		\u1_u3_idin_reg[31]/P0001 ,
		\u4_u2_buf0_reg[31]/P0001 ,
		\u4_u2_ep_match_r_reg/P0001 ,
		_w7738_
	);
	LUT3 #(
		.INIT('hb8)
	) name5989 (
		\u4_u2_buf0_orig_reg[31]/P0001 ,
		_w2269_,
		_w7738_,
		_w7739_
	);
	LUT3 #(
		.INIT('h70)
	) name5990 (
		_w2232_,
		_w2267_,
		_w7739_,
		_w7740_
	);
	LUT2 #(
		.INIT('hd)
	) name5991 (
		_w7737_,
		_w7740_,
		_w7741_
	);
	LUT3 #(
		.INIT('h2a)
	) name5992 (
		rst_i_pad,
		_w2267_,
		_w7375_,
		_w7742_
	);
	LUT4 #(
		.INIT('hd8f0)
	) name5993 (
		\u1_u3_buf0_set_reg/P0001 ,
		\u1_u3_idin_reg[3]/P0001 ,
		\u4_u2_buf0_reg[3]/P0001 ,
		\u4_u2_ep_match_r_reg/P0001 ,
		_w7743_
	);
	LUT3 #(
		.INIT('hb8)
	) name5994 (
		\u4_u2_buf0_orig_reg[3]/P0001 ,
		_w2269_,
		_w7743_,
		_w7744_
	);
	LUT3 #(
		.INIT('h70)
	) name5995 (
		_w2232_,
		_w2267_,
		_w7744_,
		_w7745_
	);
	LUT2 #(
		.INIT('hd)
	) name5996 (
		_w7742_,
		_w7745_,
		_w7746_
	);
	LUT3 #(
		.INIT('h2a)
	) name5997 (
		rst_i_pad,
		_w2267_,
		_w7381_,
		_w7747_
	);
	LUT4 #(
		.INIT('hd8f0)
	) name5998 (
		\u1_u3_buf0_set_reg/P0001 ,
		\u1_u3_idin_reg[8]/P0001 ,
		\u4_u2_buf0_reg[8]/P0001 ,
		\u4_u2_ep_match_r_reg/P0001 ,
		_w7748_
	);
	LUT3 #(
		.INIT('hb8)
	) name5999 (
		\u4_u2_buf0_orig_reg[8]/P0001 ,
		_w2269_,
		_w7748_,
		_w7749_
	);
	LUT3 #(
		.INIT('h70)
	) name6000 (
		_w2232_,
		_w2267_,
		_w7749_,
		_w7750_
	);
	LUT2 #(
		.INIT('hd)
	) name6001 (
		_w7747_,
		_w7750_,
		_w7751_
	);
	LUT3 #(
		.INIT('h2a)
	) name6002 (
		rst_i_pad,
		_w2267_,
		_w7387_,
		_w7752_
	);
	LUT4 #(
		.INIT('hd8f0)
	) name6003 (
		\u1_u3_buf0_set_reg/P0001 ,
		\u1_u3_idin_reg[9]/P0001 ,
		\u4_u2_buf0_reg[9]/P0001 ,
		\u4_u2_ep_match_r_reg/P0001 ,
		_w7753_
	);
	LUT3 #(
		.INIT('hb8)
	) name6004 (
		\u4_u2_buf0_orig_reg[9]/P0001 ,
		_w2269_,
		_w7753_,
		_w7754_
	);
	LUT3 #(
		.INIT('h70)
	) name6005 (
		_w2232_,
		_w2267_,
		_w7754_,
		_w7755_
	);
	LUT2 #(
		.INIT('hd)
	) name6006 (
		_w7752_,
		_w7755_,
		_w7756_
	);
	LUT3 #(
		.INIT('h0b)
	) name6007 (
		\u4_attach_r1_reg/P0001 ,
		\u4_attach_r_reg/P0001 ,
		\u4_int_srcb_reg[5]/P0001 ,
		_w7757_
	);
	LUT2 #(
		.INIT('h2)
	) name6008 (
		_w4041_,
		_w7757_,
		_w7758_
	);
	LUT3 #(
		.INIT('h0d)
	) name6009 (
		\u4_attach_r1_reg/P0001 ,
		\u4_attach_r_reg/P0001 ,
		\u4_int_srcb_reg[6]/P0001 ,
		_w7759_
	);
	LUT2 #(
		.INIT('h2)
	) name6010 (
		_w4041_,
		_w7759_,
		_w7760_
	);
	LUT3 #(
		.INIT('h80)
	) name6011 (
		\u0_u0_mode_hs_reg/P0001 ,
		\u4_csr_reg[11]/P0001 ,
		\u4_csr_reg[29]/P0001 ,
		_w7761_
	);
	LUT2 #(
		.INIT('h8)
	) name6012 (
		\u0_u0_mode_hs_reg/P0001 ,
		\u4_csr_reg[12]/P0001 ,
		_w7762_
	);
	LUT2 #(
		.INIT('h8)
	) name6013 (
		\u4_csr_reg[24]/P0001 ,
		\u4_csr_reg[27]/NET0131 ,
		_w7763_
	);
	LUT4 #(
		.INIT('h8000)
	) name6014 (
		\u0_u0_mode_hs_reg/P0001 ,
		\u4_csr_reg[12]/P0001 ,
		\u4_csr_reg[24]/P0001 ,
		\u4_csr_reg[27]/NET0131 ,
		_w7764_
	);
	LUT3 #(
		.INIT('h15)
	) name6015 (
		_w2118_,
		_w7761_,
		_w7764_,
		_w7765_
	);
	LUT3 #(
		.INIT('h08)
	) name6016 (
		\u0_u0_mode_hs_reg/P0001 ,
		\u4_csr_reg[11]/P0001 ,
		\u4_csr_reg[28]/P0001 ,
		_w7766_
	);
	LUT2 #(
		.INIT('h2)
	) name6017 (
		_w7764_,
		_w7766_,
		_w7767_
	);
	LUT4 #(
		.INIT('haaea)
	) name6018 (
		_w2118_,
		_w7761_,
		_w7764_,
		_w7766_,
		_w7768_
	);
	LUT2 #(
		.INIT('h4)
	) name6019 (
		\u1_u3_setup_token_reg/P0001 ,
		\u4_csr_reg[28]/P0001 ,
		_w7769_
	);
	LUT2 #(
		.INIT('h4)
	) name6020 (
		_w2503_,
		_w7769_,
		_w7770_
	);
	LUT2 #(
		.INIT('h2)
	) name6021 (
		_w7768_,
		_w7770_,
		_w7771_
	);
	LUT4 #(
		.INIT('h0080)
	) name6022 (
		\u0_u0_mode_hs_reg/P0001 ,
		\u4_csr_reg[11]/P0001 ,
		\u4_csr_reg[12]/P0001 ,
		\u4_csr_reg[29]/P0001 ,
		_w7772_
	);
	LUT2 #(
		.INIT('h8)
	) name6023 (
		_w7763_,
		_w7772_,
		_w7773_
	);
	LUT3 #(
		.INIT('h31)
	) name6024 (
		_w7765_,
		_w7767_,
		_w7773_,
		_w7774_
	);
	LUT4 #(
		.INIT('h8000)
	) name6025 (
		\u1_u0_pid_reg[0]/NET0131 ,
		\u1_u0_pid_reg[1]/NET0131 ,
		\u1_u0_pid_reg[2]/NET0131 ,
		\u1_u0_pid_reg[3]/NET0131 ,
		_w7775_
	);
	LUT4 #(
		.INIT('h1500)
	) name6026 (
		_w2118_,
		_w7763_,
		_w7772_,
		_w7775_,
		_w7776_
	);
	LUT4 #(
		.INIT('h1500)
	) name6027 (
		_w2118_,
		_w7761_,
		_w7764_,
		_w7775_,
		_w7777_
	);
	LUT2 #(
		.INIT('h1)
	) name6028 (
		_w7776_,
		_w7777_,
		_w7778_
	);
	LUT3 #(
		.INIT('h20)
	) name6029 (
		_w7764_,
		_w7766_,
		_w7775_,
		_w7779_
	);
	LUT3 #(
		.INIT('h08)
	) name6030 (
		\u0_u0_mode_hs_reg/P0001 ,
		\u4_csr_reg[12]/P0001 ,
		\u4_csr_reg[25]/P0001 ,
		_w7780_
	);
	LUT4 #(
		.INIT('h001f)
	) name6031 (
		\u4_csr_reg[24]/P0001 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		\u4_csr_reg[28]/P0001 ,
		_w7781_
	);
	LUT4 #(
		.INIT('h7500)
	) name6032 (
		\u4_csr_reg[24]/P0001 ,
		_w7761_,
		_w7780_,
		_w7781_,
		_w7782_
	);
	LUT4 #(
		.INIT('h2220)
	) name6033 (
		_w7765_,
		_w7773_,
		_w7779_,
		_w7782_,
		_w7783_
	);
	LUT4 #(
		.INIT('hffae)
	) name6034 (
		_w7771_,
		_w7774_,
		_w7778_,
		_w7783_,
		_w7784_
	);
	LUT2 #(
		.INIT('h9)
	) name6035 (
		\u4_u2_buf0_orig_reg[28]/P0001 ,
		\u4_u2_dma_out_cnt_reg[9]/P0001 ,
		_w7785_
	);
	LUT4 #(
		.INIT('h15ea)
	) name6036 (
		_w6023_,
		_w6035_,
		_w6037_,
		_w7785_,
		_w7786_
	);
	LUT2 #(
		.INIT('h9)
	) name6037 (
		\u4_u3_buf0_orig_reg[28]/P0001 ,
		\u4_u3_dma_out_cnt_reg[9]/P0001 ,
		_w7787_
	);
	LUT4 #(
		.INIT('h15ea)
	) name6038 (
		_w5948_,
		_w5960_,
		_w5962_,
		_w7787_,
		_w7788_
	);
	LUT3 #(
		.INIT('h01)
	) name6039 (
		\u0_u0_state_reg[6]/NET0131 ,
		\u0_u0_state_reg[7]/NET0131 ,
		\u0_u0_state_reg[8]/NET0131 ,
		_w7789_
	);
	LUT2 #(
		.INIT('h8)
	) name6040 (
		_w4096_,
		_w7789_,
		_w7790_
	);
	LUT4 #(
		.INIT('h0001)
	) name6041 (
		\u0_u0_state_reg[0]/NET0131 ,
		\u0_u0_state_reg[1]/P0001 ,
		\u0_u0_state_reg[2]/NET0131 ,
		\u0_u0_state_reg[3]/P0001 ,
		_w7791_
	);
	LUT3 #(
		.INIT('h80)
	) name6042 (
		_w4096_,
		_w7789_,
		_w7791_,
		_w7792_
	);
	LUT3 #(
		.INIT('h01)
	) name6043 (
		\u0_u0_state_reg[10]/P0001 ,
		\u0_u0_state_reg[11]/NET0131 ,
		\u0_u0_state_reg[12]/NET0131 ,
		_w7793_
	);
	LUT4 #(
		.INIT('h0002)
	) name6044 (
		\u0_u0_state_reg[13]/NET0131 ,
		\u0_u0_state_reg[14]/P0001 ,
		\u0_u0_state_reg[4]/NET0131 ,
		\u0_u0_state_reg[9]/P0001 ,
		_w7794_
	);
	LUT2 #(
		.INIT('h8)
	) name6045 (
		_w7793_,
		_w7794_,
		_w7795_
	);
	LUT3 #(
		.INIT('h20)
	) name6046 (
		\u0_u0_T2_wakeup_reg/P0001 ,
		\u0_u0_state_reg[1]/P0001 ,
		\u0_u0_state_reg[5]/P0001 ,
		_w7796_
	);
	LUT4 #(
		.INIT('h0080)
	) name6047 (
		\u0_u0_T1_gt_3_0_mS_reg/P0001 ,
		\u0_u0_mode_hs_reg/P0001 ,
		\u0_u0_state_reg[1]/P0001 ,
		\u0_u0_state_reg[5]/P0001 ,
		_w7797_
	);
	LUT4 #(
		.INIT('h1000)
	) name6048 (
		\LineState_r_reg[0]/P0001 ,
		\LineState_r_reg[1]/P0001 ,
		\u0_u0_mode_hs_reg/P0001 ,
		\u0_u0_state_reg[4]/NET0131 ,
		_w7798_
	);
	LUT4 #(
		.INIT('h00fe)
	) name6049 (
		TermSel_pad_o_pad,
		_w7796_,
		_w7797_,
		_w7798_,
		_w7799_
	);
	LUT3 #(
		.INIT('h70)
	) name6050 (
		_w7792_,
		_w7795_,
		_w7799_,
		_w7800_
	);
	LUT2 #(
		.INIT('h1)
	) name6051 (
		\u0_u0_state_reg[10]/P0001 ,
		\u0_u0_state_reg[13]/NET0131 ,
		_w7801_
	);
	LUT2 #(
		.INIT('h6)
	) name6052 (
		\u0_u0_state_reg[1]/P0001 ,
		\u0_u0_state_reg[5]/P0001 ,
		_w7802_
	);
	LUT4 #(
		.INIT('h0002)
	) name6053 (
		\u0_u0_state_reg[0]/NET0131 ,
		\u0_u0_state_reg[7]/NET0131 ,
		\u0_u0_state_reg[8]/NET0131 ,
		\u0_u0_state_reg[9]/P0001 ,
		_w7803_
	);
	LUT3 #(
		.INIT('h01)
	) name6054 (
		\u0_u0_state_reg[14]/P0001 ,
		\u0_u0_state_reg[1]/P0001 ,
		\u0_u0_state_reg[2]/NET0131 ,
		_w7804_
	);
	LUT4 #(
		.INIT('h2000)
	) name6055 (
		_w4098_,
		_w7802_,
		_w7803_,
		_w7804_,
		_w7805_
	);
	LUT3 #(
		.INIT('h01)
	) name6056 (
		\u0_u0_state_reg[0]/NET0131 ,
		\u0_u0_state_reg[2]/NET0131 ,
		\u0_u0_state_reg[3]/P0001 ,
		_w7806_
	);
	LUT4 #(
		.INIT('h0102)
	) name6057 (
		\u0_u0_state_reg[14]/P0001 ,
		\u0_u0_state_reg[1]/P0001 ,
		\u0_u0_state_reg[5]/P0001 ,
		\u0_u0_state_reg[9]/P0001 ,
		_w7807_
	);
	LUT2 #(
		.INIT('h8)
	) name6058 (
		_w7806_,
		_w7807_,
		_w7808_
	);
	LUT4 #(
		.INIT('h575f)
	) name6059 (
		_w4100_,
		_w7790_,
		_w7805_,
		_w7808_,
		_w7809_
	);
	LUT3 #(
		.INIT('hae)
	) name6060 (
		_w7800_,
		_w7801_,
		_w7809_,
		_w7810_
	);
	LUT2 #(
		.INIT('h9)
	) name6061 (
		\u4_u0_buf0_orig_reg[28]/P0001 ,
		\u4_u0_dma_out_cnt_reg[9]/P0001 ,
		_w7811_
	);
	LUT4 #(
		.INIT('h15ea)
	) name6062 (
		_w5973_,
		_w5985_,
		_w5987_,
		_w7811_,
		_w7812_
	);
	LUT2 #(
		.INIT('h9)
	) name6063 (
		\u4_u1_buf0_orig_reg[28]/P0001 ,
		\u4_u1_dma_out_cnt_reg[9]/P0001 ,
		_w7813_
	);
	LUT4 #(
		.INIT('h15ea)
	) name6064 (
		_w5998_,
		_w6010_,
		_w6012_,
		_w7813_,
		_w7814_
	);
	LUT3 #(
		.INIT('hac)
	) name6065 (
		\sram_data_i[22]_pad ,
		\u4_dout_reg[22]/P0001 ,
		\wb_addr_i[17]_pad ,
		_w7815_
	);
	LUT3 #(
		.INIT('hac)
	) name6066 (
		\sram_data_i[23]_pad ,
		\u4_dout_reg[23]/P0001 ,
		\wb_addr_i[17]_pad ,
		_w7816_
	);
	LUT3 #(
		.INIT('hac)
	) name6067 (
		\sram_data_i[4]_pad ,
		\u4_dout_reg[4]/P0001 ,
		\wb_addr_i[17]_pad ,
		_w7817_
	);
	LUT3 #(
		.INIT('hac)
	) name6068 (
		\sram_data_i[7]_pad ,
		\u4_dout_reg[7]/P0001 ,
		\wb_addr_i[17]_pad ,
		_w7818_
	);
	LUT3 #(
		.INIT('hac)
	) name6069 (
		\u1_u2_sizu_c_reg[0]/P0001 ,
		\u1_u3_new_size_reg[0]/P0001 ,
		\u1_u3_out_to_small_r_reg/P0001 ,
		_w7819_
	);
	LUT2 #(
		.INIT('h9)
	) name6070 (
		\u4_u2_buf0_orig_reg[27]/P0001 ,
		\u4_u2_dma_out_cnt_reg[8]/P0001 ,
		_w7820_
	);
	LUT4 #(
		.INIT('h15ea)
	) name6071 (
		_w6022_,
		_w6035_,
		_w6036_,
		_w7820_,
		_w7821_
	);
	LUT4 #(
		.INIT('h0007)
	) name6072 (
		\u4_u3_buf0_orig_reg[19]/P0001 ,
		\u4_u3_buf0_orig_reg[20]/P0001 ,
		\u4_u3_buf0_orig_reg[21]/P0001 ,
		\u4_u3_buf0_orig_reg[22]/P0001 ,
		_w7822_
	);
	LUT2 #(
		.INIT('h1)
	) name6073 (
		\u4_u3_buf0_orig_reg[23]/P0001 ,
		\u4_u3_buf0_orig_reg[24]/P0001 ,
		_w7823_
	);
	LUT4 #(
		.INIT('h0001)
	) name6074 (
		\u4_u3_buf0_orig_reg[23]/P0001 ,
		\u4_u3_buf0_orig_reg[24]/P0001 ,
		\u4_u3_buf0_orig_reg[25]/P0001 ,
		\u4_u3_buf0_orig_reg[26]/P0001 ,
		_w7824_
	);
	LUT2 #(
		.INIT('h1)
	) name6075 (
		\u4_u3_buf0_orig_reg[27]/P0001 ,
		\u4_u3_buf0_orig_reg[28]/P0001 ,
		_w7825_
	);
	LUT3 #(
		.INIT('h01)
	) name6076 (
		\u4_u3_buf0_orig_reg[27]/P0001 ,
		\u4_u3_buf0_orig_reg[28]/P0001 ,
		\u4_u3_buf0_orig_reg[29]/NET0131 ,
		_w7826_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name6077 (
		\u4_u3_buf0_orig_reg[30]/NET0131 ,
		_w7822_,
		_w7824_,
		_w7826_,
		_w7827_
	);
	LUT3 #(
		.INIT('h59)
	) name6078 (
		\u1_u3_adr_reg[1]/P0001 ,
		_w2782_,
		_w2784_,
		_w7828_
	);
	LUT2 #(
		.INIT('h6)
	) name6079 (
		_w4071_,
		_w7828_,
		_w7829_
	);
	LUT2 #(
		.INIT('h9)
	) name6080 (
		\u4_u3_buf0_orig_reg[27]/P0001 ,
		\u4_u3_dma_out_cnt_reg[8]/P0001 ,
		_w7830_
	);
	LUT4 #(
		.INIT('h15ea)
	) name6081 (
		_w5947_,
		_w5960_,
		_w5961_,
		_w7830_,
		_w7831_
	);
	LUT2 #(
		.INIT('h1)
	) name6082 (
		\u4_u0_buf0_orig_reg[23]/P0001 ,
		\u4_u0_buf0_orig_reg[24]/P0001 ,
		_w7832_
	);
	LUT4 #(
		.INIT('h0001)
	) name6083 (
		\u4_u0_buf0_orig_reg[23]/P0001 ,
		\u4_u0_buf0_orig_reg[24]/P0001 ,
		\u4_u0_buf0_orig_reg[25]/P0001 ,
		\u4_u0_buf0_orig_reg[26]/P0001 ,
		_w7833_
	);
	LUT2 #(
		.INIT('h1)
	) name6084 (
		\u4_u0_buf0_orig_reg[21]/P0001 ,
		\u4_u0_buf0_orig_reg[22]/P0001 ,
		_w7834_
	);
	LUT4 #(
		.INIT('h0007)
	) name6085 (
		\u4_u0_buf0_orig_reg[19]/P0001 ,
		\u4_u0_buf0_orig_reg[20]/P0001 ,
		\u4_u0_buf0_orig_reg[21]/P0001 ,
		\u4_u0_buf0_orig_reg[22]/P0001 ,
		_w7835_
	);
	LUT3 #(
		.INIT('h01)
	) name6086 (
		\u4_u0_buf0_orig_reg[27]/P0001 ,
		\u4_u0_buf0_orig_reg[28]/P0001 ,
		\u4_u0_buf0_orig_reg[29]/NET0131 ,
		_w7836_
	);
	LUT3 #(
		.INIT('h80)
	) name6087 (
		_w7833_,
		_w7835_,
		_w7836_,
		_w7837_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name6088 (
		\u4_u0_buf0_orig_reg[30]/NET0131 ,
		_w7833_,
		_w7835_,
		_w7836_,
		_w7838_
	);
	LUT2 #(
		.INIT('h1)
	) name6089 (
		\u4_u0_buf0_orig_reg[27]/P0001 ,
		\u4_u0_buf0_orig_reg[28]/P0001 ,
		_w7839_
	);
	LUT4 #(
		.INIT('h0001)
	) name6090 (
		\u4_u0_buf0_orig_reg[27]/P0001 ,
		\u4_u0_buf0_orig_reg[28]/P0001 ,
		\u4_u0_buf0_orig_reg[29]/NET0131 ,
		\u4_u0_buf0_orig_reg[30]/NET0131 ,
		_w7840_
	);
	LUT3 #(
		.INIT('h80)
	) name6091 (
		_w7833_,
		_w7835_,
		_w7840_,
		_w7841_
	);
	LUT2 #(
		.INIT('he)
	) name6092 (
		_w7838_,
		_w7841_,
		_w7842_
	);
	LUT2 #(
		.INIT('h9)
	) name6093 (
		\u4_u0_buf0_orig_reg[27]/P0001 ,
		\u4_u0_dma_out_cnt_reg[8]/P0001 ,
		_w7843_
	);
	LUT4 #(
		.INIT('h15ea)
	) name6094 (
		_w5972_,
		_w5985_,
		_w5986_,
		_w7843_,
		_w7844_
	);
	LUT4 #(
		.INIT('h0007)
	) name6095 (
		\u4_u1_buf0_orig_reg[19]/P0001 ,
		\u4_u1_buf0_orig_reg[20]/P0001 ,
		\u4_u1_buf0_orig_reg[21]/P0001 ,
		\u4_u1_buf0_orig_reg[22]/P0001 ,
		_w7845_
	);
	LUT2 #(
		.INIT('h1)
	) name6096 (
		\u4_u1_buf0_orig_reg[23]/P0001 ,
		\u4_u1_buf0_orig_reg[24]/P0001 ,
		_w7846_
	);
	LUT4 #(
		.INIT('h0001)
	) name6097 (
		\u4_u1_buf0_orig_reg[23]/P0001 ,
		\u4_u1_buf0_orig_reg[24]/P0001 ,
		\u4_u1_buf0_orig_reg[25]/P0001 ,
		\u4_u1_buf0_orig_reg[26]/P0001 ,
		_w7847_
	);
	LUT2 #(
		.INIT('h1)
	) name6098 (
		\u4_u1_buf0_orig_reg[27]/P0001 ,
		\u4_u1_buf0_orig_reg[28]/P0001 ,
		_w7848_
	);
	LUT3 #(
		.INIT('h01)
	) name6099 (
		\u4_u1_buf0_orig_reg[27]/P0001 ,
		\u4_u1_buf0_orig_reg[28]/P0001 ,
		\u4_u1_buf0_orig_reg[29]/NET0131 ,
		_w7849_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name6100 (
		\u4_u1_buf0_orig_reg[30]/NET0131 ,
		_w7845_,
		_w7847_,
		_w7849_,
		_w7850_
	);
	LUT2 #(
		.INIT('h9)
	) name6101 (
		\u4_u1_buf0_orig_reg[27]/P0001 ,
		\u4_u1_dma_out_cnt_reg[8]/P0001 ,
		_w7851_
	);
	LUT4 #(
		.INIT('h15ea)
	) name6102 (
		_w5997_,
		_w6010_,
		_w6011_,
		_w7851_,
		_w7852_
	);
	LUT4 #(
		.INIT('h0007)
	) name6103 (
		\u4_u2_buf0_orig_reg[19]/P0001 ,
		\u4_u2_buf0_orig_reg[20]/P0001 ,
		\u4_u2_buf0_orig_reg[21]/P0001 ,
		\u4_u2_buf0_orig_reg[22]/P0001 ,
		_w7853_
	);
	LUT2 #(
		.INIT('h1)
	) name6104 (
		\u4_u2_buf0_orig_reg[23]/P0001 ,
		\u4_u2_buf0_orig_reg[24]/P0001 ,
		_w7854_
	);
	LUT4 #(
		.INIT('h0001)
	) name6105 (
		\u4_u2_buf0_orig_reg[23]/P0001 ,
		\u4_u2_buf0_orig_reg[24]/P0001 ,
		\u4_u2_buf0_orig_reg[25]/P0001 ,
		\u4_u2_buf0_orig_reg[26]/P0001 ,
		_w7855_
	);
	LUT2 #(
		.INIT('h1)
	) name6106 (
		\u4_u2_buf0_orig_reg[27]/P0001 ,
		\u4_u2_buf0_orig_reg[28]/P0001 ,
		_w7856_
	);
	LUT3 #(
		.INIT('h01)
	) name6107 (
		\u4_u2_buf0_orig_reg[27]/P0001 ,
		\u4_u2_buf0_orig_reg[28]/P0001 ,
		\u4_u2_buf0_orig_reg[29]/NET0131 ,
		_w7857_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name6108 (
		\u4_u2_buf0_orig_reg[30]/NET0131 ,
		_w7853_,
		_w7855_,
		_w7857_,
		_w7858_
	);
	LUT4 #(
		.INIT('h2000)
	) name6109 (
		\u0_rx_active_reg/P0001 ,
		\u0_rx_err_reg/P0001 ,
		\u0_rx_valid_reg/P0001 ,
		\u1_u0_rxv1_reg/P0001 ,
		_w7859_
	);
	LUT4 #(
		.INIT('h005d)
	) name6110 (
		\u1_u0_rxv2_reg/P0001 ,
		_w3671_,
		_w3672_,
		_w7859_,
		_w7860_
	);
	LUT3 #(
		.INIT('h11)
	) name6111 (
		\u1_u0_rxv2_reg/P0001 ,
		_w3671_,
		_w3672_,
		_w7861_
	);
	LUT4 #(
		.INIT('h040f)
	) name6112 (
		_w4886_,
		_w6898_,
		_w7860_,
		_w7861_,
		_w7862_
	);
	LUT2 #(
		.INIT('h8)
	) name6113 (
		rst_i_pad,
		_w7862_,
		_w7863_
	);
	LUT2 #(
		.INIT('h8)
	) name6114 (
		\u1_u3_buffer_done_reg/P0001 ,
		\u1_u3_state_reg[8]/P0001 ,
		_w7864_
	);
	LUT4 #(
		.INIT('h4000)
	) name6115 (
		\u1_u3_buf0_not_aloc_reg/P0001 ,
		\u1_u3_buffer_done_reg/P0001 ,
		\u1_u3_state_reg[8]/P0001 ,
		\u4_u2_ep_match_r_reg/P0001 ,
		_w7865_
	);
	LUT2 #(
		.INIT('h1)
	) name6116 (
		\u4_u2_int_stat_reg[3]/P0001 ,
		_w7865_,
		_w7866_
	);
	LUT4 #(
		.INIT('h00fd)
	) name6117 (
		\u1_u3_in_token_reg/NET0131 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		\u4_u2_int_stat_reg[3]/P0001 ,
		_w7867_
	);
	LUT3 #(
		.INIT('hd0)
	) name6118 (
		_w2352_,
		_w2353_,
		_w7867_,
		_w7868_
	);
	LUT3 #(
		.INIT('h02)
	) name6119 (
		_w3890_,
		_w7866_,
		_w7868_,
		_w7869_
	);
	LUT4 #(
		.INIT('h4000)
	) name6120 (
		\u1_u3_buf0_not_aloc_reg/P0001 ,
		\u1_u3_buffer_done_reg/P0001 ,
		\u1_u3_state_reg[8]/P0001 ,
		\u4_u3_ep_match_r_reg/P0001 ,
		_w7870_
	);
	LUT2 #(
		.INIT('h1)
	) name6121 (
		\u4_u3_int_stat_reg[3]/P0001 ,
		_w7870_,
		_w7871_
	);
	LUT4 #(
		.INIT('h00fd)
	) name6122 (
		\u1_u3_in_token_reg/NET0131 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		\u4_u3_int_stat_reg[3]/P0001 ,
		_w7872_
	);
	LUT3 #(
		.INIT('hd0)
	) name6123 (
		_w2352_,
		_w2353_,
		_w7872_,
		_w7873_
	);
	LUT3 #(
		.INIT('h02)
	) name6124 (
		_w3893_,
		_w7871_,
		_w7873_,
		_w7874_
	);
	LUT4 #(
		.INIT('h0102)
	) name6125 (
		\u0_u0_state_reg[13]/NET0131 ,
		\u0_u0_state_reg[14]/P0001 ,
		\u0_u0_state_reg[4]/NET0131 ,
		\u0_u0_state_reg[9]/P0001 ,
		_w7875_
	);
	LUT2 #(
		.INIT('h8)
	) name6126 (
		_w7793_,
		_w7875_,
		_w7876_
	);
	LUT2 #(
		.INIT('h2)
	) name6127 (
		XcvSelect_pad_o_pad,
		_w7798_,
		_w7877_
	);
	LUT3 #(
		.INIT('h70)
	) name6128 (
		_w7792_,
		_w7876_,
		_w7877_,
		_w7878_
	);
	LUT2 #(
		.INIT('h4)
	) name6129 (
		\u0_u0_state_reg[13]/NET0131 ,
		\u0_u0_state_reg[14]/P0001 ,
		_w7879_
	);
	LUT4 #(
		.INIT('h0001)
	) name6130 (
		\u0_u0_state_reg[10]/P0001 ,
		\u0_u0_state_reg[11]/NET0131 ,
		\u0_u0_state_reg[12]/NET0131 ,
		\u0_u0_state_reg[9]/P0001 ,
		_w7880_
	);
	LUT4 #(
		.INIT('h8000)
	) name6131 (
		_w4096_,
		_w7789_,
		_w7791_,
		_w7880_,
		_w7881_
	);
	LUT3 #(
		.INIT('h80)
	) name6132 (
		\u0_u0_T1_gt_3_0_mS_reg/P0001 ,
		\u0_u0_mode_hs_reg/P0001 ,
		\u0_u0_state_reg[1]/P0001 ,
		_w7882_
	);
	LUT4 #(
		.INIT('h0015)
	) name6133 (
		_w4333_,
		_w7879_,
		_w7881_,
		_w7882_,
		_w7883_
	);
	LUT2 #(
		.INIT('hb)
	) name6134 (
		_w7878_,
		_w7883_,
		_w7884_
	);
	LUT3 #(
		.INIT('h31)
	) name6135 (
		susp_o_pad,
		\u4_int_srcb_reg[3]/P0001 ,
		\u4_suspend_r1_reg/P0001 ,
		_w7885_
	);
	LUT2 #(
		.INIT('h2)
	) name6136 (
		_w4041_,
		_w7885_,
		_w7886_
	);
	LUT3 #(
		.INIT('h23)
	) name6137 (
		susp_o_pad,
		\u4_int_srcb_reg[4]/P0001 ,
		\u4_suspend_r1_reg/P0001 ,
		_w7887_
	);
	LUT2 #(
		.INIT('h2)
	) name6138 (
		_w4041_,
		_w7887_,
		_w7888_
	);
	LUT3 #(
		.INIT('h10)
	) name6139 (
		\u0_u0_T1_gt_5_0_mS_reg/P0001 ,
		\u0_u0_idle_cnt1_next_reg[0]/P0001 ,
		\u0_u0_ps_cnt_clr_reg/P0001 ,
		_w7889_
	);
	LUT3 #(
		.INIT('h23)
	) name6140 (
		\u0_u0_T1_gt_5_0_mS_reg/P0001 ,
		\u0_u0_idle_cnt1_reg[0]/P0001 ,
		\u0_u0_ps_cnt_clr_reg/P0001 ,
		_w7890_
	);
	LUT3 #(
		.INIT('h02)
	) name6141 (
		_w5770_,
		_w7889_,
		_w7890_,
		_w7891_
	);
	LUT3 #(
		.INIT('hd0)
	) name6142 (
		_w5763_,
		_w5768_,
		_w7891_,
		_w7892_
	);
	LUT2 #(
		.INIT('h4)
	) name6143 (
		_w5765_,
		_w7892_,
		_w7893_
	);
	LUT3 #(
		.INIT('h10)
	) name6144 (
		\u0_u0_T1_gt_5_0_mS_reg/P0001 ,
		\u0_u0_idle_cnt1_next_reg[1]/P0001 ,
		\u0_u0_ps_cnt_clr_reg/P0001 ,
		_w7894_
	);
	LUT3 #(
		.INIT('h23)
	) name6145 (
		\u0_u0_T1_gt_5_0_mS_reg/P0001 ,
		\u0_u0_idle_cnt1_reg[1]/P0001 ,
		\u0_u0_ps_cnt_clr_reg/P0001 ,
		_w7895_
	);
	LUT3 #(
		.INIT('h02)
	) name6146 (
		_w5770_,
		_w7894_,
		_w7895_,
		_w7896_
	);
	LUT3 #(
		.INIT('hd0)
	) name6147 (
		_w5763_,
		_w5768_,
		_w7896_,
		_w7897_
	);
	LUT2 #(
		.INIT('h4)
	) name6148 (
		_w5765_,
		_w7897_,
		_w7898_
	);
	LUT3 #(
		.INIT('h10)
	) name6149 (
		\u0_u0_T1_gt_5_0_mS_reg/P0001 ,
		\u0_u0_idle_cnt1_next_reg[2]/P0001 ,
		\u0_u0_ps_cnt_clr_reg/P0001 ,
		_w7899_
	);
	LUT3 #(
		.INIT('h23)
	) name6150 (
		\u0_u0_T1_gt_5_0_mS_reg/P0001 ,
		\u0_u0_idle_cnt1_reg[2]/P0001 ,
		\u0_u0_ps_cnt_clr_reg/P0001 ,
		_w7900_
	);
	LUT3 #(
		.INIT('h02)
	) name6151 (
		_w5770_,
		_w7899_,
		_w7900_,
		_w7901_
	);
	LUT3 #(
		.INIT('hd0)
	) name6152 (
		_w5763_,
		_w5768_,
		_w7901_,
		_w7902_
	);
	LUT2 #(
		.INIT('h4)
	) name6153 (
		_w5765_,
		_w7902_,
		_w7903_
	);
	LUT3 #(
		.INIT('h10)
	) name6154 (
		\u0_u0_T1_gt_5_0_mS_reg/P0001 ,
		\u0_u0_idle_cnt1_next_reg[5]/P0001 ,
		\u0_u0_ps_cnt_clr_reg/P0001 ,
		_w7904_
	);
	LUT3 #(
		.INIT('h23)
	) name6155 (
		\u0_u0_T1_gt_5_0_mS_reg/P0001 ,
		\u0_u0_idle_cnt1_reg[5]/P0001 ,
		\u0_u0_ps_cnt_clr_reg/P0001 ,
		_w7905_
	);
	LUT3 #(
		.INIT('h02)
	) name6156 (
		_w5770_,
		_w7904_,
		_w7905_,
		_w7906_
	);
	LUT3 #(
		.INIT('hd0)
	) name6157 (
		_w5763_,
		_w5768_,
		_w7906_,
		_w7907_
	);
	LUT2 #(
		.INIT('h4)
	) name6158 (
		_w5765_,
		_w7907_,
		_w7908_
	);
	LUT3 #(
		.INIT('h10)
	) name6159 (
		\u0_u0_T1_gt_5_0_mS_reg/P0001 ,
		\u0_u0_idle_cnt1_next_reg[6]/P0001 ,
		\u0_u0_ps_cnt_clr_reg/P0001 ,
		_w7909_
	);
	LUT3 #(
		.INIT('h23)
	) name6160 (
		\u0_u0_T1_gt_5_0_mS_reg/P0001 ,
		\u0_u0_idle_cnt1_reg[6]/P0001 ,
		\u0_u0_ps_cnt_clr_reg/P0001 ,
		_w7910_
	);
	LUT3 #(
		.INIT('h02)
	) name6161 (
		_w5770_,
		_w7909_,
		_w7910_,
		_w7911_
	);
	LUT3 #(
		.INIT('hd0)
	) name6162 (
		_w5763_,
		_w5768_,
		_w7911_,
		_w7912_
	);
	LUT2 #(
		.INIT('h4)
	) name6163 (
		_w5765_,
		_w7912_,
		_w7913_
	);
	LUT4 #(
		.INIT('h0001)
	) name6164 (
		\u0_u0_idle_cnt1_reg[0]/P0001 ,
		\u0_u0_idle_cnt1_reg[1]/P0001 ,
		\u0_u0_idle_cnt1_reg[2]/P0001 ,
		\u0_u0_idle_cnt1_reg[3]/P0001 ,
		_w7914_
	);
	LUT2 #(
		.INIT('h8)
	) name6165 (
		\u0_u0_idle_cnt1_reg[4]/P0001 ,
		\u0_u0_idle_cnt1_reg[6]/P0001 ,
		_w7915_
	);
	LUT3 #(
		.INIT('h07)
	) name6166 (
		\u0_u0_idle_cnt1_reg[5]/P0001 ,
		\u0_u0_idle_cnt1_reg[6]/P0001 ,
		\u0_u0_idle_cnt1_reg[7]/P0001 ,
		_w7916_
	);
	LUT3 #(
		.INIT('hb0)
	) name6167 (
		_w7914_,
		_w7915_,
		_w7916_,
		_w7917_
	);
	LUT3 #(
		.INIT('h0d)
	) name6168 (
		_w5763_,
		_w5768_,
		_w7917_,
		_w7918_
	);
	LUT2 #(
		.INIT('h4)
	) name6169 (
		_w5765_,
		_w7918_,
		_w7919_
	);
	LUT4 #(
		.INIT('h4000)
	) name6170 (
		\u1_u3_buf0_not_aloc_reg/P0001 ,
		\u1_u3_buffer_done_reg/P0001 ,
		\u1_u3_state_reg[8]/P0001 ,
		\u4_u0_ep_match_r_reg/P0001 ,
		_w7920_
	);
	LUT2 #(
		.INIT('h1)
	) name6171 (
		\u4_u0_int_stat_reg[3]/P0001 ,
		_w7920_,
		_w7921_
	);
	LUT4 #(
		.INIT('h00fd)
	) name6172 (
		\u1_u3_in_token_reg/NET0131 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		\u4_u0_int_stat_reg[3]/P0001 ,
		_w7922_
	);
	LUT3 #(
		.INIT('hd0)
	) name6173 (
		_w2352_,
		_w2353_,
		_w7922_,
		_w7923_
	);
	LUT3 #(
		.INIT('h02)
	) name6174 (
		_w3896_,
		_w7921_,
		_w7923_,
		_w7924_
	);
	LUT3 #(
		.INIT('h04)
	) name6175 (
		_w7761_,
		_w7764_,
		_w7766_,
		_w7925_
	);
	LUT3 #(
		.INIT('h80)
	) name6176 (
		_w7763_,
		_w7772_,
		_w7775_,
		_w7926_
	);
	LUT2 #(
		.INIT('h8)
	) name6177 (
		_w7925_,
		_w7926_,
		_w7927_
	);
	LUT2 #(
		.INIT('h4)
	) name6178 (
		\u4_csr_reg[25]/P0001 ,
		\u4_csr_reg[28]/P0001 ,
		_w7928_
	);
	LUT4 #(
		.INIT('h0200)
	) name6179 (
		\u4_csr_reg[24]/P0001 ,
		\u4_csr_reg[25]/P0001 ,
		\u4_csr_reg[27]/NET0131 ,
		\u4_csr_reg[28]/P0001 ,
		_w7929_
	);
	LUT2 #(
		.INIT('h8)
	) name6180 (
		_w7772_,
		_w7929_,
		_w7930_
	);
	LUT3 #(
		.INIT('h20)
	) name6181 (
		_w7765_,
		_w7925_,
		_w7930_,
		_w7931_
	);
	LUT2 #(
		.INIT('h4)
	) name6182 (
		\u1_u3_setup_token_reg/P0001 ,
		\u4_csr_reg[29]/P0001 ,
		_w7932_
	);
	LUT2 #(
		.INIT('h8)
	) name6183 (
		_w2503_,
		_w7932_,
		_w7933_
	);
	LUT2 #(
		.INIT('h2)
	) name6184 (
		_w7768_,
		_w7933_,
		_w7934_
	);
	LUT3 #(
		.INIT('hfe)
	) name6185 (
		_w7927_,
		_w7931_,
		_w7934_,
		_w7935_
	);
	LUT2 #(
		.INIT('h2)
	) name6186 (
		\u0_u0_idle_long_reg/P0001 ,
		\u0_u0_ps_cnt_clr_reg/P0001 ,
		_w7936_
	);
	LUT3 #(
		.INIT('h02)
	) name6187 (
		\u0_u0_idle_long_reg/P0001 ,
		\u0_u0_ps_cnt_clr_reg/P0001 ,
		\u0_u0_ps_cnt_reg[0]/P0001 ,
		_w7937_
	);
	LUT3 #(
		.INIT('hd0)
	) name6188 (
		_w5763_,
		_w5768_,
		_w7937_,
		_w7938_
	);
	LUT2 #(
		.INIT('h4)
	) name6189 (
		_w5765_,
		_w7938_,
		_w7939_
	);
	LUT3 #(
		.INIT('hd0)
	) name6190 (
		_w5763_,
		_w5768_,
		_w7936_,
		_w7940_
	);
	LUT2 #(
		.INIT('h9)
	) name6191 (
		\u0_u0_ps_cnt_reg[0]/P0001 ,
		\u0_u0_ps_cnt_reg[1]/P0001 ,
		_w7941_
	);
	LUT4 #(
		.INIT('hffa2)
	) name6192 (
		_w5762_,
		_w5763_,
		_w5764_,
		_w7941_,
		_w7942_
	);
	LUT2 #(
		.INIT('h2)
	) name6193 (
		_w7940_,
		_w7942_,
		_w7943_
	);
	LUT3 #(
		.INIT('h78)
	) name6194 (
		\u0_u0_ps_cnt_reg[0]/P0001 ,
		\u0_u0_ps_cnt_reg[1]/P0001 ,
		\u0_u0_ps_cnt_reg[2]/P0001 ,
		_w7944_
	);
	LUT4 #(
		.INIT('ha2ff)
	) name6195 (
		_w5762_,
		_w5763_,
		_w5764_,
		_w7944_,
		_w7945_
	);
	LUT2 #(
		.INIT('h2)
	) name6196 (
		_w7940_,
		_w7945_,
		_w7946_
	);
	LUT4 #(
		.INIT('h7f80)
	) name6197 (
		\u0_u0_ps_cnt_reg[0]/P0001 ,
		\u0_u0_ps_cnt_reg[1]/P0001 ,
		\u0_u0_ps_cnt_reg[2]/P0001 ,
		\u0_u0_ps_cnt_reg[3]/P0001 ,
		_w7947_
	);
	LUT2 #(
		.INIT('h8)
	) name6198 (
		_w7936_,
		_w7947_,
		_w7948_
	);
	LUT3 #(
		.INIT('hd0)
	) name6199 (
		_w5763_,
		_w5768_,
		_w7948_,
		_w7949_
	);
	LUT2 #(
		.INIT('h4)
	) name6200 (
		_w5765_,
		_w7949_,
		_w7950_
	);
	LUT4 #(
		.INIT('h8000)
	) name6201 (
		\u1_u3_rx_ack_to_cnt_reg[0]/P0001 ,
		\u1_u3_rx_ack_to_cnt_reg[1]/P0001 ,
		\u1_u3_rx_ack_to_cnt_reg[2]/P0001 ,
		\u1_u3_rx_ack_to_cnt_reg[3]/P0001 ,
		_w7951_
	);
	LUT3 #(
		.INIT('h14)
	) name6202 (
		\u1_u3_rx_ack_to_clr_reg/P0001 ,
		\u1_u3_rx_ack_to_cnt_reg[4]/P0001 ,
		_w7951_,
		_w7952_
	);
	LUT2 #(
		.INIT('h4)
	) name6203 (
		_w4316_,
		_w4324_,
		_w7953_
	);
	LUT4 #(
		.INIT('h0004)
	) name6204 (
		\u0_u0_T1_gt_3_0_mS_reg/P0001 ,
		\u0_u0_state_reg[1]/P0001 ,
		\u0_u0_state_reg[3]/P0001 ,
		\u0_u0_state_reg[6]/NET0131 ,
		_w7954_
	);
	LUT4 #(
		.INIT('h8000)
	) name6205 (
		_w4108_,
		_w4109_,
		_w4323_,
		_w7954_,
		_w7955_
	);
	LUT4 #(
		.INIT('h0001)
	) name6206 (
		\u0_u0_state_reg[0]/NET0131 ,
		\u0_u0_state_reg[10]/P0001 ,
		\u0_u0_state_reg[7]/NET0131 ,
		\u0_u0_state_reg[8]/NET0131 ,
		_w7956_
	);
	LUT3 #(
		.INIT('h80)
	) name6207 (
		_w4098_,
		_w4101_,
		_w7956_,
		_w7957_
	);
	LUT3 #(
		.INIT('h06)
	) name6208 (
		\u0_u0_state_reg[13]/NET0131 ,
		\u0_u0_state_reg[14]/P0001 ,
		\u0_u0_state_reg[9]/P0001 ,
		_w7958_
	);
	LUT2 #(
		.INIT('h2)
	) name6209 (
		\u0_u0_state_reg[13]/NET0131 ,
		\u0_u0_state_reg[1]/P0001 ,
		_w7959_
	);
	LUT3 #(
		.INIT('h8c)
	) name6210 (
		_w4117_,
		_w7958_,
		_w7959_,
		_w7960_
	);
	LUT4 #(
		.INIT('h0777)
	) name6211 (
		_w7953_,
		_w7955_,
		_w7957_,
		_w7960_,
		_w7961_
	);
	LUT4 #(
		.INIT('h8000)
	) name6212 (
		_w4099_,
		_w4108_,
		_w4109_,
		_w4323_,
		_w7962_
	);
	LUT4 #(
		.INIT('h0e00)
	) name6213 (
		\u0_u0_T2_gt_100_uS_reg/P0001 ,
		\u0_u0_state_reg[1]/P0001 ,
		\u0_u0_state_reg[3]/P0001 ,
		\u0_u0_state_reg[6]/NET0131 ,
		_w7963_
	);
	LUT2 #(
		.INIT('h1)
	) name6214 (
		\u0_u0_me_cnt_100_ms_reg/P0001 ,
		\u0_u0_state_reg[1]/P0001 ,
		_w7964_
	);
	LUT4 #(
		.INIT('h3f15)
	) name6215 (
		_w5762_,
		_w7962_,
		_w7963_,
		_w7964_,
		_w7965_
	);
	LUT3 #(
		.INIT('h2a)
	) name6216 (
		_w4103_,
		_w7961_,
		_w7965_,
		_w7966_
	);
	LUT4 #(
		.INIT('h8000)
	) name6217 (
		\u1_u3_tx_data_to_cnt_reg[0]/P0001 ,
		\u1_u3_tx_data_to_cnt_reg[1]/P0001 ,
		\u1_u3_tx_data_to_cnt_reg[2]/P0001 ,
		\u1_u3_tx_data_to_cnt_reg[3]/P0001 ,
		_w7967_
	);
	LUT3 #(
		.INIT('h14)
	) name6218 (
		\u0_rx_active_reg/P0001 ,
		\u1_u3_tx_data_to_cnt_reg[4]/P0001 ,
		_w7967_,
		_w7968_
	);
	LUT4 #(
		.INIT('h4000)
	) name6219 (
		\u1_u3_buf0_not_aloc_reg/P0001 ,
		\u1_u3_buffer_done_reg/P0001 ,
		\u1_u3_state_reg[8]/P0001 ,
		\u4_u1_ep_match_r_reg/P0001 ,
		_w7969_
	);
	LUT2 #(
		.INIT('h1)
	) name6220 (
		\u4_u1_int_stat_reg[3]/P0001 ,
		_w7969_,
		_w7970_
	);
	LUT4 #(
		.INIT('h00fd)
	) name6221 (
		\u1_u3_in_token_reg/NET0131 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		\u4_u1_int_stat_reg[3]/P0001 ,
		_w7971_
	);
	LUT3 #(
		.INIT('hd0)
	) name6222 (
		_w2352_,
		_w2353_,
		_w7971_,
		_w7972_
	);
	LUT3 #(
		.INIT('h02)
	) name6223 (
		_w3899_,
		_w7970_,
		_w7972_,
		_w7973_
	);
	LUT4 #(
		.INIT('h6996)
	) name6224 (
		\u0_rx_data_reg[6]/P0001 ,
		\u0_rx_data_reg[7]/P0001 ,
		\u1_u0_crc16_sum_reg[8]/P0001 ,
		\u1_u0_crc16_sum_reg[9]/P0001 ,
		_w7974_
	);
	LUT3 #(
		.INIT('h96)
	) name6225 (
		_w6920_,
		_w6923_,
		_w7974_,
		_w7975_
	);
	LUT4 #(
		.INIT('hc888)
	) name6226 (
		_w3671_,
		_w4884_,
		_w4885_,
		_w6898_,
		_w7976_
	);
	LUT2 #(
		.INIT('h2)
	) name6227 (
		\u1_u0_crc16_sum_reg[0]/P0001 ,
		_w3671_,
		_w7977_
	);
	LUT4 #(
		.INIT('hdf00)
	) name6228 (
		\u0_rx_active_reg/P0001 ,
		\u0_rx_err_reg/P0001 ,
		\u0_rx_valid_reg/P0001 ,
		\u1_u0_crc16_sum_reg[0]/P0001 ,
		_w7978_
	);
	LUT2 #(
		.INIT('h1)
	) name6229 (
		_w6911_,
		_w7978_,
		_w7979_
	);
	LUT4 #(
		.INIT('h4f00)
	) name6230 (
		_w4886_,
		_w6898_,
		_w7977_,
		_w7979_,
		_w7980_
	);
	LUT4 #(
		.INIT('h60ff)
	) name6231 (
		_w6908_,
		_w7975_,
		_w7976_,
		_w7980_,
		_w7981_
	);
	LUT3 #(
		.INIT('h31)
	) name6232 (
		\u0_rx_active_reg/P0001 ,
		\u1_u0_crc16_sum_reg[10]/P0001 ,
		\u1_u0_rx_active_r_reg/P0001 ,
		_w7982_
	);
	LUT4 #(
		.INIT('h1500)
	) name6233 (
		_w6897_,
		_w6898_,
		_w6899_,
		_w7982_,
		_w7983_
	);
	LUT3 #(
		.INIT('h31)
	) name6234 (
		\u0_rx_active_reg/P0001 ,
		\u1_u0_crc16_sum_reg[2]/P0001 ,
		\u1_u0_rx_active_r_reg/P0001 ,
		_w7984_
	);
	LUT4 #(
		.INIT('hea00)
	) name6235 (
		_w6897_,
		_w6898_,
		_w6899_,
		_w7984_,
		_w7985_
	);
	LUT2 #(
		.INIT('h1)
	) name6236 (
		_w7983_,
		_w7985_,
		_w7986_
	);
	LUT3 #(
		.INIT('h31)
	) name6237 (
		\u0_rx_active_reg/P0001 ,
		\u1_u0_crc16_sum_reg[11]/P0001 ,
		\u1_u0_rx_active_r_reg/P0001 ,
		_w7987_
	);
	LUT4 #(
		.INIT('h1500)
	) name6238 (
		_w6897_,
		_w6898_,
		_w6899_,
		_w7987_,
		_w7988_
	);
	LUT3 #(
		.INIT('h31)
	) name6239 (
		\u0_rx_active_reg/P0001 ,
		\u1_u0_crc16_sum_reg[3]/P0001 ,
		\u1_u0_rx_active_r_reg/P0001 ,
		_w7989_
	);
	LUT4 #(
		.INIT('hea00)
	) name6240 (
		_w6897_,
		_w6898_,
		_w6899_,
		_w7989_,
		_w7990_
	);
	LUT2 #(
		.INIT('h1)
	) name6241 (
		_w7988_,
		_w7990_,
		_w7991_
	);
	LUT3 #(
		.INIT('h31)
	) name6242 (
		\u0_rx_active_reg/P0001 ,
		\u1_u0_crc16_sum_reg[12]/P0001 ,
		\u1_u0_rx_active_r_reg/P0001 ,
		_w7992_
	);
	LUT4 #(
		.INIT('h1500)
	) name6243 (
		_w6897_,
		_w6898_,
		_w6899_,
		_w7992_,
		_w7993_
	);
	LUT3 #(
		.INIT('h31)
	) name6244 (
		\u0_rx_active_reg/P0001 ,
		\u1_u0_crc16_sum_reg[4]/P0001 ,
		\u1_u0_rx_active_r_reg/P0001 ,
		_w7994_
	);
	LUT4 #(
		.INIT('hea00)
	) name6245 (
		_w6897_,
		_w6898_,
		_w6899_,
		_w7994_,
		_w7995_
	);
	LUT2 #(
		.INIT('h1)
	) name6246 (
		_w7993_,
		_w7995_,
		_w7996_
	);
	LUT3 #(
		.INIT('h31)
	) name6247 (
		\u0_rx_active_reg/P0001 ,
		\u1_u0_crc16_sum_reg[13]/P0001 ,
		\u1_u0_rx_active_r_reg/P0001 ,
		_w7997_
	);
	LUT4 #(
		.INIT('h1500)
	) name6248 (
		_w6897_,
		_w6898_,
		_w6899_,
		_w7997_,
		_w7998_
	);
	LUT3 #(
		.INIT('h31)
	) name6249 (
		\u0_rx_active_reg/P0001 ,
		\u1_u0_crc16_sum_reg[5]/P0001 ,
		\u1_u0_rx_active_r_reg/P0001 ,
		_w7999_
	);
	LUT4 #(
		.INIT('hea00)
	) name6250 (
		_w6897_,
		_w6898_,
		_w6899_,
		_w7999_,
		_w8000_
	);
	LUT2 #(
		.INIT('h1)
	) name6251 (
		_w7998_,
		_w8000_,
		_w8001_
	);
	LUT3 #(
		.INIT('h31)
	) name6252 (
		\u0_rx_active_reg/P0001 ,
		\u1_u0_crc16_sum_reg[14]/P0001 ,
		\u1_u0_rx_active_r_reg/P0001 ,
		_w8002_
	);
	LUT4 #(
		.INIT('h1500)
	) name6253 (
		_w6897_,
		_w6898_,
		_w6899_,
		_w8002_,
		_w8003_
	);
	LUT3 #(
		.INIT('h31)
	) name6254 (
		\u0_rx_active_reg/P0001 ,
		\u1_u0_crc16_sum_reg[6]/P0001 ,
		\u1_u0_rx_active_r_reg/P0001 ,
		_w8004_
	);
	LUT4 #(
		.INIT('hea00)
	) name6255 (
		_w6897_,
		_w6898_,
		_w6899_,
		_w8004_,
		_w8005_
	);
	LUT2 #(
		.INIT('h1)
	) name6256 (
		_w8003_,
		_w8005_,
		_w8006_
	);
	LUT4 #(
		.INIT('hea00)
	) name6257 (
		_w6897_,
		_w6898_,
		_w6899_,
		_w7974_,
		_w8007_
	);
	LUT2 #(
		.INIT('h2)
	) name6258 (
		\u1_u0_crc16_sum_reg[2]/P0001 ,
		_w3671_,
		_w8008_
	);
	LUT4 #(
		.INIT('hdf00)
	) name6259 (
		\u0_rx_active_reg/P0001 ,
		\u0_rx_err_reg/P0001 ,
		\u0_rx_valid_reg/P0001 ,
		\u1_u0_crc16_sum_reg[2]/P0001 ,
		_w8009_
	);
	LUT2 #(
		.INIT('h1)
	) name6260 (
		_w6911_,
		_w8009_,
		_w8010_
	);
	LUT4 #(
		.INIT('h4f00)
	) name6261 (
		_w4886_,
		_w6898_,
		_w8008_,
		_w8010_,
		_w8011_
	);
	LUT2 #(
		.INIT('hb)
	) name6262 (
		_w8007_,
		_w8011_,
		_w8012_
	);
	LUT4 #(
		.INIT('h6996)
	) name6263 (
		\u0_rx_data_reg[5]/P0001 ,
		\u0_rx_data_reg[6]/P0001 ,
		\u1_u0_crc16_sum_reg[10]/P0001 ,
		\u1_u0_crc16_sum_reg[9]/P0001 ,
		_w8013_
	);
	LUT2 #(
		.INIT('h1)
	) name6264 (
		_w6911_,
		_w8013_,
		_w8014_
	);
	LUT4 #(
		.INIT('hea00)
	) name6265 (
		_w6897_,
		_w6898_,
		_w6899_,
		_w8014_,
		_w8015_
	);
	LUT4 #(
		.INIT('h1500)
	) name6266 (
		_w6897_,
		_w6898_,
		_w6899_,
		_w7989_,
		_w8016_
	);
	LUT2 #(
		.INIT('h1)
	) name6267 (
		_w8015_,
		_w8016_,
		_w8017_
	);
	LUT4 #(
		.INIT('h00ea)
	) name6268 (
		_w6897_,
		_w6898_,
		_w6899_,
		_w6921_,
		_w8018_
	);
	LUT2 #(
		.INIT('h2)
	) name6269 (
		\u1_u0_crc16_sum_reg[4]/P0001 ,
		_w3671_,
		_w8019_
	);
	LUT4 #(
		.INIT('hdf00)
	) name6270 (
		\u0_rx_active_reg/P0001 ,
		\u0_rx_err_reg/P0001 ,
		\u0_rx_valid_reg/P0001 ,
		\u1_u0_crc16_sum_reg[4]/P0001 ,
		_w8020_
	);
	LUT2 #(
		.INIT('h1)
	) name6271 (
		_w6911_,
		_w8020_,
		_w8021_
	);
	LUT4 #(
		.INIT('h4f00)
	) name6272 (
		_w4886_,
		_w6898_,
		_w8019_,
		_w8021_,
		_w8022_
	);
	LUT2 #(
		.INIT('hb)
	) name6273 (
		_w8018_,
		_w8022_,
		_w8023_
	);
	LUT4 #(
		.INIT('h6996)
	) name6274 (
		\u0_rx_data_reg[3]/P0001 ,
		\u0_rx_data_reg[4]/P0001 ,
		\u1_u0_crc16_sum_reg[11]/P0001 ,
		\u1_u0_crc16_sum_reg[12]/P0001 ,
		_w8024_
	);
	LUT2 #(
		.INIT('h1)
	) name6275 (
		_w6911_,
		_w8024_,
		_w8025_
	);
	LUT4 #(
		.INIT('hea00)
	) name6276 (
		_w6897_,
		_w6898_,
		_w6899_,
		_w8025_,
		_w8026_
	);
	LUT4 #(
		.INIT('h1500)
	) name6277 (
		_w6897_,
		_w6898_,
		_w6899_,
		_w7999_,
		_w8027_
	);
	LUT2 #(
		.INIT('h1)
	) name6278 (
		_w8026_,
		_w8027_,
		_w8028_
	);
	LUT4 #(
		.INIT('h9669)
	) name6279 (
		\u0_rx_data_reg[2]/P0001 ,
		\u0_rx_data_reg[3]/P0001 ,
		\u1_u0_crc16_sum_reg[12]/P0001 ,
		\u1_u0_crc16_sum_reg[13]/P0001 ,
		_w8029_
	);
	LUT2 #(
		.INIT('h4)
	) name6280 (
		_w6911_,
		_w8029_,
		_w8030_
	);
	LUT4 #(
		.INIT('hea00)
	) name6281 (
		_w6897_,
		_w6898_,
		_w6899_,
		_w8030_,
		_w8031_
	);
	LUT4 #(
		.INIT('h1500)
	) name6282 (
		_w6897_,
		_w6898_,
		_w6899_,
		_w8004_,
		_w8032_
	);
	LUT2 #(
		.INIT('h1)
	) name6283 (
		_w8031_,
		_w8032_,
		_w8033_
	);
	LUT4 #(
		.INIT('h6996)
	) name6284 (
		\u0_rx_data_reg[1]/P0001 ,
		\u0_rx_data_reg[2]/P0001 ,
		\u1_u0_crc16_sum_reg[13]/P0001 ,
		\u1_u0_crc16_sum_reg[14]/P0001 ,
		_w8034_
	);
	LUT2 #(
		.INIT('h1)
	) name6285 (
		_w6911_,
		_w8034_,
		_w8035_
	);
	LUT4 #(
		.INIT('hea00)
	) name6286 (
		_w6897_,
		_w6898_,
		_w6899_,
		_w8035_,
		_w8036_
	);
	LUT3 #(
		.INIT('h31)
	) name6287 (
		\u0_rx_active_reg/P0001 ,
		\u1_u0_crc16_sum_reg[7]/P0001 ,
		\u1_u0_rx_active_r_reg/P0001 ,
		_w8037_
	);
	LUT4 #(
		.INIT('h1500)
	) name6288 (
		_w6897_,
		_w6898_,
		_w6899_,
		_w8037_,
		_w8038_
	);
	LUT2 #(
		.INIT('h1)
	) name6289 (
		_w8036_,
		_w8038_,
		_w8039_
	);
	LUT3 #(
		.INIT('h96)
	) name6290 (
		\u1_u0_crc16_sum_reg[0]/P0001 ,
		\u1_u0_crc16_sum_reg[14]/P0001 ,
		\u1_u0_crc16_sum_reg[15]/P0001 ,
		_w8040_
	);
	LUT2 #(
		.INIT('h9)
	) name6291 (
		_w6892_,
		_w8040_,
		_w8041_
	);
	LUT4 #(
		.INIT('hea00)
	) name6292 (
		_w6897_,
		_w6898_,
		_w6899_,
		_w8041_,
		_w8042_
	);
	LUT2 #(
		.INIT('h2)
	) name6293 (
		\u1_u0_crc16_sum_reg[8]/P0001 ,
		_w3671_,
		_w8043_
	);
	LUT4 #(
		.INIT('hdf00)
	) name6294 (
		\u0_rx_active_reg/P0001 ,
		\u0_rx_err_reg/P0001 ,
		\u0_rx_valid_reg/P0001 ,
		\u1_u0_crc16_sum_reg[8]/P0001 ,
		_w8044_
	);
	LUT2 #(
		.INIT('h1)
	) name6295 (
		_w6911_,
		_w8044_,
		_w8045_
	);
	LUT4 #(
		.INIT('h4f00)
	) name6296 (
		_w4886_,
		_w6898_,
		_w8043_,
		_w8045_,
		_w8046_
	);
	LUT2 #(
		.INIT('hb)
	) name6297 (
		_w8042_,
		_w8046_,
		_w8047_
	);
	LUT3 #(
		.INIT('h96)
	) name6298 (
		\u0_rx_data_reg[0]/P0001 ,
		\u1_u0_crc16_sum_reg[15]/P0001 ,
		\u1_u0_crc16_sum_reg[1]/P0001 ,
		_w8048_
	);
	LUT2 #(
		.INIT('h1)
	) name6299 (
		_w6911_,
		_w8048_,
		_w8049_
	);
	LUT4 #(
		.INIT('hea00)
	) name6300 (
		_w6897_,
		_w6898_,
		_w6899_,
		_w8049_,
		_w8050_
	);
	LUT3 #(
		.INIT('h31)
	) name6301 (
		\u0_rx_active_reg/P0001 ,
		\u1_u0_crc16_sum_reg[9]/P0001 ,
		\u1_u0_rx_active_r_reg/P0001 ,
		_w8051_
	);
	LUT4 #(
		.INIT('h1500)
	) name6302 (
		_w6897_,
		_w6898_,
		_w6899_,
		_w8051_,
		_w8052_
	);
	LUT2 #(
		.INIT('h1)
	) name6303 (
		_w8050_,
		_w8052_,
		_w8053_
	);
	LUT4 #(
		.INIT('h8acf)
	) name6304 (
		\u4_buf0_reg[26]/NET0131 ,
		\u4_buf0_reg[27]/P0001 ,
		\u4_csr_reg[10]/P0001 ,
		\u4_csr_reg[9]/NET0131 ,
		_w8054_
	);
	LUT2 #(
		.INIT('h1)
	) name6305 (
		\u4_buf0_reg[28]/P0001 ,
		\u4_buf0_reg[29]/P0001 ,
		_w8055_
	);
	LUT3 #(
		.INIT('h31)
	) name6306 (
		\u4_buf0_reg[27]/P0001 ,
		\u4_buf0_reg[30]/P0001 ,
		\u4_csr_reg[10]/P0001 ,
		_w8056_
	);
	LUT3 #(
		.INIT('h40)
	) name6307 (
		_w8054_,
		_w8055_,
		_w8056_,
		_w8057_
	);
	LUT4 #(
		.INIT('h8caf)
	) name6308 (
		\u4_buf0_reg[24]/NET0131 ,
		\u4_buf0_reg[25]/NET0131 ,
		\u4_csr_reg[7]/P0001 ,
		\u4_csr_reg[8]/P0001 ,
		_w8058_
	);
	LUT4 #(
		.INIT('hf531)
	) name6309 (
		\u4_buf0_reg[23]/NET0131 ,
		\u4_buf0_reg[24]/NET0131 ,
		\u4_csr_reg[6]/NET0131 ,
		\u4_csr_reg[7]/P0001 ,
		_w8059_
	);
	LUT2 #(
		.INIT('h2)
	) name6310 (
		_w8058_,
		_w8059_,
		_w8060_
	);
	LUT4 #(
		.INIT('hf531)
	) name6311 (
		\u4_buf0_reg[21]/NET0131 ,
		\u4_buf0_reg[22]/NET0131 ,
		\u4_csr_reg[4]/NET0131 ,
		\u4_csr_reg[5]/NET0131 ,
		_w8061_
	);
	LUT4 #(
		.INIT('h8caf)
	) name6312 (
		\u4_buf0_reg[20]/NET0131 ,
		\u4_buf0_reg[21]/NET0131 ,
		\u4_csr_reg[3]/P0001 ,
		\u4_csr_reg[4]/NET0131 ,
		_w8062_
	);
	LUT2 #(
		.INIT('h2)
	) name6313 (
		_w8061_,
		_w8062_,
		_w8063_
	);
	LUT4 #(
		.INIT('h5010)
	) name6314 (
		\u4_buf0_reg[17]/NET0131 ,
		\u4_buf0_reg[18]/P0001 ,
		\u4_csr_reg[0]/P0001 ,
		\u4_csr_reg[1]/P0001 ,
		_w8064_
	);
	LUT4 #(
		.INIT('h8caf)
	) name6315 (
		\u4_buf0_reg[18]/P0001 ,
		\u4_buf0_reg[19]/NET0131 ,
		\u4_csr_reg[1]/P0001 ,
		\u4_csr_reg[2]/NET0131 ,
		_w8065_
	);
	LUT4 #(
		.INIT('hf531)
	) name6316 (
		\u4_buf0_reg[19]/NET0131 ,
		\u4_buf0_reg[20]/NET0131 ,
		\u4_csr_reg[2]/NET0131 ,
		\u4_csr_reg[3]/P0001 ,
		_w8066_
	);
	LUT4 #(
		.INIT('h8a00)
	) name6317 (
		_w8061_,
		_w8064_,
		_w8065_,
		_w8066_,
		_w8067_
	);
	LUT4 #(
		.INIT('h8caf)
	) name6318 (
		\u4_buf0_reg[22]/NET0131 ,
		\u4_buf0_reg[23]/NET0131 ,
		\u4_csr_reg[5]/NET0131 ,
		\u4_csr_reg[6]/NET0131 ,
		_w8068_
	);
	LUT2 #(
		.INIT('h8)
	) name6319 (
		_w8058_,
		_w8068_,
		_w8069_
	);
	LUT4 #(
		.INIT('h5455)
	) name6320 (
		_w8060_,
		_w8063_,
		_w8067_,
		_w8069_,
		_w8070_
	);
	LUT4 #(
		.INIT('hf531)
	) name6321 (
		\u4_buf0_reg[25]/NET0131 ,
		\u4_buf0_reg[26]/NET0131 ,
		\u4_csr_reg[8]/P0001 ,
		\u4_csr_reg[9]/NET0131 ,
		_w8071_
	);
	LUT3 #(
		.INIT('h80)
	) name6322 (
		_w8055_,
		_w8056_,
		_w8071_,
		_w8072_
	);
	LUT3 #(
		.INIT('hea)
	) name6323 (
		_w8057_,
		_w8070_,
		_w8072_,
		_w8073_
	);
	LUT3 #(
		.INIT('h20)
	) name6324 (
		rst_i_pad,
		\u4_u2_int_re_reg/P0001 ,
		\u4_u2_int_stat_reg[4]/P0001 ,
		_w8074_
	);
	LUT3 #(
		.INIT('h40)
	) name6325 (
		\u1_u3_buf1_not_aloc_reg/P0001 ,
		\u1_u3_buffer_done_reg/P0001 ,
		\u1_u3_state_reg[8]/P0001 ,
		_w8075_
	);
	LUT4 #(
		.INIT('h0d00)
	) name6326 (
		_w2352_,
		_w2353_,
		_w2356_,
		_w8075_,
		_w8076_
	);
	LUT3 #(
		.INIT('hec)
	) name6327 (
		_w7253_,
		_w8074_,
		_w8076_,
		_w8077_
	);
	LUT4 #(
		.INIT('h0001)
	) name6328 (
		\u4_u3_csr0_reg[3]/NET0131 ,
		\u4_u3_csr0_reg[4]/P0001 ,
		\u4_u3_csr0_reg[5]/P0001 ,
		\u4_u3_csr0_reg[6]/P0001 ,
		_w8078_
	);
	LUT4 #(
		.INIT('h0001)
	) name6329 (
		\u4_u3_csr0_reg[0]/P0001 ,
		\u4_u3_csr0_reg[10]/P0001 ,
		\u4_u3_csr0_reg[1]/P0001 ,
		\u4_u3_csr0_reg[2]/P0001 ,
		_w8079_
	);
	LUT3 #(
		.INIT('h01)
	) name6330 (
		\u4_u3_csr0_reg[7]/P0001 ,
		\u4_u3_csr0_reg[8]/P0001 ,
		\u4_u3_csr0_reg[9]/P0001 ,
		_w8080_
	);
	LUT3 #(
		.INIT('h80)
	) name6331 (
		_w8078_,
		_w8079_,
		_w8080_,
		_w8081_
	);
	LUT2 #(
		.INIT('h2)
	) name6332 (
		_w4394_,
		_w4566_,
		_w8082_
	);
	LUT3 #(
		.INIT('h23)
	) name6333 (
		\u4_u3_csr0_reg[10]/P0001 ,
		\u4_u3_dma_in_cnt_reg[11]/P0001 ,
		\u4_u3_dma_in_cnt_reg[8]/P0001 ,
		_w8083_
	);
	LUT2 #(
		.INIT('h8)
	) name6334 (
		_w4896_,
		_w8083_,
		_w8084_
	);
	LUT4 #(
		.INIT('h8f00)
	) name6335 (
		_w4561_,
		_w4565_,
		_w8082_,
		_w8084_,
		_w8085_
	);
	LUT2 #(
		.INIT('h1)
	) name6336 (
		_w8081_,
		_w8085_,
		_w8086_
	);
	LUT3 #(
		.INIT('h20)
	) name6337 (
		rst_i_pad,
		\u4_u3_int_re_reg/P0001 ,
		\u4_u3_int_stat_reg[4]/P0001 ,
		_w8087_
	);
	LUT3 #(
		.INIT('hf8)
	) name6338 (
		_w7394_,
		_w8076_,
		_w8087_,
		_w8088_
	);
	LUT4 #(
		.INIT('h0001)
	) name6339 (
		\u4_u0_csr0_reg[3]/NET0131 ,
		\u4_u0_csr0_reg[4]/P0001 ,
		\u4_u0_csr0_reg[5]/P0001 ,
		\u4_u0_csr0_reg[6]/P0001 ,
		_w8089_
	);
	LUT4 #(
		.INIT('h0001)
	) name6340 (
		\u4_u0_csr0_reg[0]/P0001 ,
		\u4_u0_csr0_reg[10]/P0001 ,
		\u4_u0_csr0_reg[1]/P0001 ,
		\u4_u0_csr0_reg[2]/P0001 ,
		_w8090_
	);
	LUT3 #(
		.INIT('h01)
	) name6341 (
		\u4_u0_csr0_reg[7]/P0001 ,
		\u4_u0_csr0_reg[8]/P0001 ,
		\u4_u0_csr0_reg[9]/P0001 ,
		_w8091_
	);
	LUT3 #(
		.INIT('h80)
	) name6342 (
		_w8089_,
		_w8090_,
		_w8091_,
		_w8092_
	);
	LUT2 #(
		.INIT('h2)
	) name6343 (
		_w4426_,
		_w4589_,
		_w8093_
	);
	LUT3 #(
		.INIT('h23)
	) name6344 (
		\u4_u0_csr0_reg[10]/P0001 ,
		\u4_u0_dma_in_cnt_reg[11]/P0001 ,
		\u4_u0_dma_in_cnt_reg[8]/P0001 ,
		_w8094_
	);
	LUT2 #(
		.INIT('h8)
	) name6345 (
		_w4910_,
		_w8094_,
		_w8095_
	);
	LUT4 #(
		.INIT('h8f00)
	) name6346 (
		_w4584_,
		_w4588_,
		_w8093_,
		_w8095_,
		_w8096_
	);
	LUT2 #(
		.INIT('h1)
	) name6347 (
		_w8092_,
		_w8096_,
		_w8097_
	);
	LUT3 #(
		.INIT('h20)
	) name6348 (
		rst_i_pad,
		\u4_u0_int_re_reg/P0001 ,
		\u4_u0_int_stat_reg[4]/P0001 ,
		_w8098_
	);
	LUT3 #(
		.INIT('hf8)
	) name6349 (
		_w7522_,
		_w8076_,
		_w8098_,
		_w8099_
	);
	LUT4 #(
		.INIT('h0001)
	) name6350 (
		\u4_u1_csr0_reg[3]/NET0131 ,
		\u4_u1_csr0_reg[4]/P0001 ,
		\u4_u1_csr0_reg[5]/P0001 ,
		\u4_u1_csr0_reg[6]/P0001 ,
		_w8100_
	);
	LUT4 #(
		.INIT('h0001)
	) name6351 (
		\u4_u1_csr0_reg[0]/P0001 ,
		\u4_u1_csr0_reg[10]/P0001 ,
		\u4_u1_csr0_reg[1]/P0001 ,
		\u4_u1_csr0_reg[2]/P0001 ,
		_w8101_
	);
	LUT3 #(
		.INIT('h01)
	) name6352 (
		\u4_u1_csr0_reg[7]/P0001 ,
		\u4_u1_csr0_reg[8]/P0001 ,
		\u4_u1_csr0_reg[9]/P0001 ,
		_w8102_
	);
	LUT3 #(
		.INIT('h80)
	) name6353 (
		_w8100_,
		_w8101_,
		_w8102_,
		_w8103_
	);
	LUT3 #(
		.INIT('h40)
	) name6354 (
		_w4473_,
		_w4929_,
		_w5110_,
		_w8104_
	);
	LUT3 #(
		.INIT('h80)
	) name6355 (
		_w4606_,
		_w4929_,
		_w5110_,
		_w8105_
	);
	LUT4 #(
		.INIT('h0203)
	) name6356 (
		_w4605_,
		_w8103_,
		_w8104_,
		_w8105_,
		_w8106_
	);
	LUT3 #(
		.INIT('h20)
	) name6357 (
		rst_i_pad,
		\u4_u1_int_re_reg/P0001 ,
		\u4_u1_int_stat_reg[4]/P0001 ,
		_w8107_
	);
	LUT3 #(
		.INIT('hf8)
	) name6358 (
		_w7640_,
		_w8076_,
		_w8107_,
		_w8108_
	);
	LUT2 #(
		.INIT('h4)
	) name6359 (
		\u0_u0_T1_gt_3_0_mS_reg/P0001 ,
		\u0_u0_state_reg[9]/P0001 ,
		_w8109_
	);
	LUT3 #(
		.INIT('hc8)
	) name6360 (
		_w4316_,
		_w4324_,
		_w8109_,
		_w8110_
	);
	LUT4 #(
		.INIT('h0ddd)
	) name6361 (
		_w4347_,
		_w4357_,
		_w5763_,
		_w8110_,
		_w8111_
	);
	LUT2 #(
		.INIT('h8)
	) name6362 (
		\u0_u0_T1_gt_5_0_mS_reg/P0001 ,
		\u0_u0_resume_req_s_reg/P0001 ,
		_w8112_
	);
	LUT3 #(
		.INIT('h70)
	) name6363 (
		\u0_u0_T1_gt_5_0_mS_reg/P0001 ,
		\u0_u0_resume_req_s_reg/P0001 ,
		\u0_u0_state_reg[9]/P0001 ,
		_w8113_
	);
	LUT3 #(
		.INIT('h23)
	) name6364 (
		_w4119_,
		_w4354_,
		_w8113_,
		_w8114_
	);
	LUT4 #(
		.INIT('hbb0b)
	) name6365 (
		\u0_u0_T2_gt_1_0_mS_reg/P0001 ,
		_w4199_,
		_w4343_,
		_w8114_,
		_w8115_
	);
	LUT3 #(
		.INIT('h2a)
	) name6366 (
		_w4103_,
		_w8111_,
		_w8115_,
		_w8116_
	);
	LUT3 #(
		.INIT('h23)
	) name6367 (
		\u4_u2_csr0_reg[10]/P0001 ,
		\u4_u2_dma_in_cnt_reg[11]/P0001 ,
		\u4_u2_dma_in_cnt_reg[8]/P0001 ,
		_w8117_
	);
	LUT4 #(
		.INIT('h0023)
	) name6368 (
		\u4_u2_csr0_reg[9]/P0001 ,
		\u4_u2_dma_in_cnt_reg[10]/P0001 ,
		\u4_u2_dma_in_cnt_reg[7]/P0001 ,
		\u4_u2_dma_in_cnt_reg[9]/P0001 ,
		_w8118_
	);
	LUT2 #(
		.INIT('h8)
	) name6369 (
		_w8117_,
		_w8118_,
		_w8119_
	);
	LUT4 #(
		.INIT('h0001)
	) name6370 (
		\u4_u2_csr0_reg[3]/NET0131 ,
		\u4_u2_csr0_reg[4]/P0001 ,
		\u4_u2_csr0_reg[5]/P0001 ,
		\u4_u2_csr0_reg[6]/P0001 ,
		_w8120_
	);
	LUT4 #(
		.INIT('h0001)
	) name6371 (
		\u4_u2_csr0_reg[0]/P0001 ,
		\u4_u2_csr0_reg[10]/P0001 ,
		\u4_u2_csr0_reg[1]/P0001 ,
		\u4_u2_csr0_reg[2]/P0001 ,
		_w8121_
	);
	LUT3 #(
		.INIT('h01)
	) name6372 (
		\u4_u2_csr0_reg[7]/P0001 ,
		\u4_u2_csr0_reg[8]/P0001 ,
		\u4_u2_csr0_reg[9]/P0001 ,
		_w8122_
	);
	LUT3 #(
		.INIT('h80)
	) name6373 (
		_w8120_,
		_w8121_,
		_w8122_,
		_w8123_
	);
	LUT4 #(
		.INIT('h0002)
	) name6374 (
		\u4_u2_csr0_reg[10]/P0001 ,
		\u4_u2_dma_in_cnt_reg[10]/P0001 ,
		\u4_u2_dma_in_cnt_reg[8]/P0001 ,
		\u4_u2_dma_in_cnt_reg[9]/P0001 ,
		_w8124_
	);
	LUT2 #(
		.INIT('h8)
	) name6375 (
		_w8117_,
		_w8124_,
		_w8125_
	);
	LUT3 #(
		.INIT('h01)
	) name6376 (
		_w8119_,
		_w8123_,
		_w8125_,
		_w8126_
	);
	LUT3 #(
		.INIT('h02)
	) name6377 (
		_w4500_,
		_w8123_,
		_w8125_,
		_w8127_
	);
	LUT3 #(
		.INIT('hec)
	) name6378 (
		_w4499_,
		_w8126_,
		_w8127_,
		_w8128_
	);
	LUT4 #(
		.INIT('he0f0)
	) name6379 (
		\LineState_r_reg[0]/P0001 ,
		\LineState_r_reg[1]/P0001 ,
		\OpMode_pad_o[1]_pad ,
		\u0_u0_state_reg[4]/NET0131 ,
		_w8129_
	);
	LUT2 #(
		.INIT('h8)
	) name6380 (
		\u0_u0_T2_wakeup_reg/P0001 ,
		\u0_u0_state_reg[5]/P0001 ,
		_w8130_
	);
	LUT2 #(
		.INIT('h1)
	) name6381 (
		_w8129_,
		_w8130_,
		_w8131_
	);
	LUT4 #(
		.INIT('h143c)
	) name6382 (
		\u0_u0_T2_wakeup_reg/P0001 ,
		\u0_u0_state_reg[13]/NET0131 ,
		\u0_u0_state_reg[14]/P0001 ,
		\u0_u0_state_reg[5]/P0001 ,
		_w8132_
	);
	LUT4 #(
		.INIT('habaf)
	) name6383 (
		_w4199_,
		_w7881_,
		_w8131_,
		_w8132_,
		_w8133_
	);
	LUT2 #(
		.INIT('h4)
	) name6384 (
		\u4_csr_reg[24]/P0001 ,
		\u4_csr_reg[28]/P0001 ,
		_w8134_
	);
	LUT3 #(
		.INIT('h07)
	) name6385 (
		_w7772_,
		_w7928_,
		_w8134_,
		_w8135_
	);
	LUT3 #(
		.INIT('h08)
	) name6386 (
		\u0_u0_mode_hs_reg/P0001 ,
		\u4_csr_reg[12]/P0001 ,
		\u4_csr_reg[28]/P0001 ,
		_w8136_
	);
	LUT4 #(
		.INIT('h0070)
	) name6387 (
		\u0_u0_mode_hs_reg/P0001 ,
		\u4_csr_reg[11]/P0001 ,
		\u4_csr_reg[24]/P0001 ,
		\u4_csr_reg[25]/P0001 ,
		_w8137_
	);
	LUT3 #(
		.INIT('h2a)
	) name6388 (
		\u4_csr_reg[26]/NET0131 ,
		_w8136_,
		_w8137_,
		_w8138_
	);
	LUT3 #(
		.INIT('h23)
	) name6389 (
		\u1_u3_setup_token_reg/P0001 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[28]/P0001 ,
		_w8139_
	);
	LUT4 #(
		.INIT('h7770)
	) name6390 (
		_w2503_,
		_w7932_,
		_w8139_,
		_w2356_,
		_w8140_
	);
	LUT4 #(
		.INIT('h0015)
	) name6391 (
		\u4_csr_reg[27]/NET0131 ,
		_w8135_,
		_w8138_,
		_w8140_,
		_w8141_
	);
	LUT3 #(
		.INIT('h08)
	) name6392 (
		\u0_u0_mode_hs_reg/P0001 ,
		\u4_csr_reg[12]/P0001 ,
		\u4_csr_reg[29]/P0001 ,
		_w8142_
	);
	LUT4 #(
		.INIT('h8088)
	) name6393 (
		\u0_u0_mode_hs_reg/P0001 ,
		\u4_csr_reg[11]/P0001 ,
		\u4_csr_reg[24]/P0001 ,
		\u4_csr_reg[28]/P0001 ,
		_w8143_
	);
	LUT2 #(
		.INIT('h4)
	) name6394 (
		_w8142_,
		_w8143_,
		_w8144_
	);
	LUT4 #(
		.INIT('h7000)
	) name6395 (
		\u0_u0_mode_hs_reg/P0001 ,
		\u4_csr_reg[11]/P0001 ,
		\u4_csr_reg[24]/P0001 ,
		\u4_csr_reg[27]/NET0131 ,
		_w8145_
	);
	LUT3 #(
		.INIT('h8d)
	) name6396 (
		\u4_csr_reg[24]/P0001 ,
		\u4_csr_reg[25]/P0001 ,
		\u4_csr_reg[28]/P0001 ,
		_w8146_
	);
	LUT4 #(
		.INIT('h008a)
	) name6397 (
		_w2120_,
		_w7762_,
		_w8145_,
		_w8146_,
		_w8147_
	);
	LUT3 #(
		.INIT('h08)
	) name6398 (
		\u1_u0_pid_reg[0]/NET0131 ,
		\u1_u0_pid_reg[1]/NET0131 ,
		\u1_u0_pid_reg[3]/NET0131 ,
		_w8148_
	);
	LUT3 #(
		.INIT('h04)
	) name6399 (
		_w7762_,
		_w8145_,
		_w8148_,
		_w8149_
	);
	LUT3 #(
		.INIT('h0b)
	) name6400 (
		_w8144_,
		_w8147_,
		_w8149_,
		_w8150_
	);
	LUT2 #(
		.INIT('hb)
	) name6401 (
		_w8141_,
		_w8150_,
		_w8151_
	);
	LUT2 #(
		.INIT('h8)
	) name6402 (
		\u0_u0_idle_cnt1_reg[4]/P0001 ,
		\u0_u0_idle_cnt1_reg[5]/P0001 ,
		_w8152_
	);
	LUT3 #(
		.INIT('h8a)
	) name6403 (
		_w7215_,
		_w7914_,
		_w8152_,
		_w8153_
	);
	LUT3 #(
		.INIT('h0d)
	) name6404 (
		_w5763_,
		_w5768_,
		_w8153_,
		_w8154_
	);
	LUT2 #(
		.INIT('h4)
	) name6405 (
		_w5765_,
		_w8154_,
		_w8155_
	);
	LUT4 #(
		.INIT('h9ccc)
	) name6406 (
		\u4_u3_buf0_orig_reg[25]/P0001 ,
		\u4_u3_buf0_orig_reg[26]/P0001 ,
		_w7822_,
		_w7823_,
		_w8156_
	);
	LUT3 #(
		.INIT('hac)
	) name6407 (
		\sram_data_i[16]_pad ,
		\u4_dout_reg[16]/P0001 ,
		\wb_addr_i[17]_pad ,
		_w8157_
	);
	LUT3 #(
		.INIT('hac)
	) name6408 (
		\sram_data_i[17]_pad ,
		\u4_dout_reg[17]/P0001 ,
		\wb_addr_i[17]_pad ,
		_w8158_
	);
	LUT3 #(
		.INIT('hac)
	) name6409 (
		\sram_data_i[18]_pad ,
		\u4_dout_reg[18]/P0001 ,
		\wb_addr_i[17]_pad ,
		_w8159_
	);
	LUT3 #(
		.INIT('hac)
	) name6410 (
		\sram_data_i[19]_pad ,
		\u4_dout_reg[19]/P0001 ,
		\wb_addr_i[17]_pad ,
		_w8160_
	);
	LUT3 #(
		.INIT('hac)
	) name6411 (
		\sram_data_i[20]_pad ,
		\u4_dout_reg[20]/P0001 ,
		\wb_addr_i[17]_pad ,
		_w8161_
	);
	LUT3 #(
		.INIT('hac)
	) name6412 (
		\sram_data_i[21]_pad ,
		\u4_dout_reg[21]/P0001 ,
		\wb_addr_i[17]_pad ,
		_w8162_
	);
	LUT3 #(
		.INIT('hac)
	) name6413 (
		\sram_data_i[25]_pad ,
		\u4_dout_reg[25]/P0001 ,
		\wb_addr_i[17]_pad ,
		_w8163_
	);
	LUT3 #(
		.INIT('hac)
	) name6414 (
		\sram_data_i[26]_pad ,
		\u4_dout_reg[26]/P0001 ,
		\wb_addr_i[17]_pad ,
		_w8164_
	);
	LUT3 #(
		.INIT('hac)
	) name6415 (
		\sram_data_i[27]_pad ,
		\u4_dout_reg[27]/P0001 ,
		\wb_addr_i[17]_pad ,
		_w8165_
	);
	LUT3 #(
		.INIT('hac)
	) name6416 (
		\sram_data_i[28]_pad ,
		\u4_dout_reg[28]/P0001 ,
		\wb_addr_i[17]_pad ,
		_w8166_
	);
	LUT3 #(
		.INIT('hac)
	) name6417 (
		\sram_data_i[29]_pad ,
		\u4_dout_reg[29]/P0001 ,
		\wb_addr_i[17]_pad ,
		_w8167_
	);
	LUT3 #(
		.INIT('hac)
	) name6418 (
		\sram_data_i[30]_pad ,
		\u4_dout_reg[30]/P0001 ,
		\wb_addr_i[17]_pad ,
		_w8168_
	);
	LUT3 #(
		.INIT('hac)
	) name6419 (
		\sram_data_i[31]_pad ,
		\u4_dout_reg[31]/P0001 ,
		\wb_addr_i[17]_pad ,
		_w8169_
	);
	LUT3 #(
		.INIT('hac)
	) name6420 (
		\sram_data_i[5]_pad ,
		\u4_dout_reg[5]/P0001 ,
		\wb_addr_i[17]_pad ,
		_w8170_
	);
	LUT3 #(
		.INIT('hac)
	) name6421 (
		\sram_data_i[6]_pad ,
		\u4_dout_reg[6]/P0001 ,
		\wb_addr_i[17]_pad ,
		_w8171_
	);
	LUT3 #(
		.INIT('hac)
	) name6422 (
		\sram_data_i[8]_pad ,
		\u4_dout_reg[8]/P0001 ,
		\wb_addr_i[17]_pad ,
		_w8172_
	);
	LUT3 #(
		.INIT('h01)
	) name6423 (
		\u4_u0_buf0_orig_reg[23]/P0001 ,
		\u4_u0_buf0_orig_reg[24]/P0001 ,
		\u4_u0_buf0_orig_reg[25]/P0001 ,
		_w8173_
	);
	LUT4 #(
		.INIT('hcaea)
	) name6424 (
		\u4_u0_buf0_orig_reg[26]/P0001 ,
		_w7833_,
		_w7835_,
		_w8173_,
		_w8174_
	);
	LUT3 #(
		.INIT('hac)
	) name6425 (
		\sram_data_i[24]_pad ,
		\u4_dout_reg[24]/P0001 ,
		\wb_addr_i[17]_pad ,
		_w8175_
	);
	LUT4 #(
		.INIT('h9ccc)
	) name6426 (
		\u4_u1_buf0_orig_reg[25]/P0001 ,
		\u4_u1_buf0_orig_reg[26]/P0001 ,
		_w7845_,
		_w7846_,
		_w8176_
	);
	LUT4 #(
		.INIT('h9ccc)
	) name6427 (
		\u4_u2_buf0_orig_reg[25]/P0001 ,
		\u4_u2_buf0_orig_reg[26]/P0001 ,
		_w7853_,
		_w7854_,
		_w8177_
	);
	LUT3 #(
		.INIT('h6a)
	) name6428 (
		\u4_u3_buf0_orig_reg[27]/P0001 ,
		_w7822_,
		_w7824_,
		_w8178_
	);
	LUT3 #(
		.INIT('h6a)
	) name6429 (
		\u4_u0_buf0_orig_reg[27]/P0001 ,
		_w7833_,
		_w7835_,
		_w8179_
	);
	LUT3 #(
		.INIT('h6a)
	) name6430 (
		\u4_u1_buf0_orig_reg[27]/P0001 ,
		_w7845_,
		_w7847_,
		_w8180_
	);
	LUT3 #(
		.INIT('ha6)
	) name6431 (
		\u1_u3_new_sizeb_reg[1]/P0001 ,
		_w2782_,
		_w2784_,
		_w8181_
	);
	LUT2 #(
		.INIT('h9)
	) name6432 (
		_w8181_,
		_w3440_,
		_w8182_
	);
	LUT3 #(
		.INIT('h6a)
	) name6433 (
		\u4_u2_buf0_orig_reg[27]/P0001 ,
		_w7853_,
		_w7855_,
		_w8183_
	);
	LUT2 #(
		.INIT('h1)
	) name6434 (
		\u1_u0_rxv1_reg/P0001 ,
		_w3671_,
		_w8184_
	);
	LUT4 #(
		.INIT('h0800)
	) name6435 (
		rst_i_pad,
		\u0_rx_active_reg/P0001 ,
		\u0_rx_err_reg/P0001 ,
		\u0_rx_valid_reg/P0001 ,
		_w8185_
	);
	LUT2 #(
		.INIT('h8)
	) name6436 (
		rst_i_pad,
		\u1_u0_rxv1_reg/P0001 ,
		_w8186_
	);
	LUT4 #(
		.INIT('h020f)
	) name6437 (
		_w3671_,
		_w3672_,
		_w8185_,
		_w8186_,
		_w8187_
	);
	LUT4 #(
		.INIT('h004f)
	) name6438 (
		_w4886_,
		_w6898_,
		_w8184_,
		_w8187_,
		_w8188_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name6439 (
		\u0_u0_state_reg[11]/NET0131 ,
		\u0_u0_state_reg[12]/NET0131 ,
		_w4112_,
		_w4119_,
		_w8189_
	);
	LUT4 #(
		.INIT('h3323)
	) name6440 (
		\u0_u0_chirp_cnt_is_6_reg/P0001 ,
		\u0_u0_chirp_cnt_reg[0]/P0001 ,
		_w4110_,
		_w8189_,
		_w8190_
	);
	LUT2 #(
		.INIT('h4)
	) name6441 (
		\u0_u0_chirp_cnt_is_6_reg/P0001 ,
		\u0_u0_chirp_cnt_reg[0]/P0001 ,
		_w8191_
	);
	LUT4 #(
		.INIT('h5155)
	) name6442 (
		\u0_u0_state_reg[10]/P0001 ,
		_w4110_,
		_w8189_,
		_w8191_,
		_w8192_
	);
	LUT2 #(
		.INIT('h4)
	) name6443 (
		_w8190_,
		_w8192_,
		_w8193_
	);
	LUT3 #(
		.INIT('h80)
	) name6444 (
		\u4_u2_csr1_reg[0]/P0001 ,
		_w3762_,
		_w3763_,
		_w8194_
	);
	LUT2 #(
		.INIT('h8)
	) name6445 (
		_w3761_,
		_w8194_,
		_w8195_
	);
	LUT3 #(
		.INIT('h80)
	) name6446 (
		\u4_u0_csr1_reg[0]/P0001 ,
		_w3755_,
		_w3756_,
		_w8196_
	);
	LUT3 #(
		.INIT('h07)
	) name6447 (
		\u4_u1_csr1_reg[0]/P0001 ,
		_w3768_,
		_w8196_,
		_w8197_
	);
	LUT3 #(
		.INIT('h80)
	) name6448 (
		\u4_u3_csr1_reg[0]/P0001 ,
		_w3761_,
		_w3773_,
		_w8198_
	);
	LUT3 #(
		.INIT('h80)
	) name6449 (
		\u4_csr_reg[15]/NET0131 ,
		_w3761_,
		_w3775_,
		_w8199_
	);
	LUT4 #(
		.INIT('hfffb)
	) name6450 (
		_w8195_,
		_w8197_,
		_w8198_,
		_w8199_,
		_w8200_
	);
	LUT3 #(
		.INIT('h80)
	) name6451 (
		\u4_u2_csr1_reg[1]/P0001 ,
		_w3762_,
		_w3763_,
		_w8201_
	);
	LUT2 #(
		.INIT('h8)
	) name6452 (
		_w3761_,
		_w8201_,
		_w8202_
	);
	LUT3 #(
		.INIT('h80)
	) name6453 (
		\u4_u0_csr1_reg[1]/P0001 ,
		_w3755_,
		_w3756_,
		_w8203_
	);
	LUT3 #(
		.INIT('h07)
	) name6454 (
		\u4_u1_csr1_reg[1]/P0001 ,
		_w3768_,
		_w8203_,
		_w8204_
	);
	LUT3 #(
		.INIT('h80)
	) name6455 (
		\u4_u3_csr1_reg[1]/P0001 ,
		_w3761_,
		_w3773_,
		_w8205_
	);
	LUT3 #(
		.INIT('h80)
	) name6456 (
		\u4_csr_reg[16]/P0001 ,
		_w3761_,
		_w3775_,
		_w8206_
	);
	LUT4 #(
		.INIT('hfffb)
	) name6457 (
		_w8202_,
		_w8204_,
		_w8205_,
		_w8206_,
		_w8207_
	);
	LUT3 #(
		.INIT('h80)
	) name6458 (
		\u4_u2_buf1_reg[5]/P0001 ,
		_w3762_,
		_w3763_,
		_w8208_
	);
	LUT2 #(
		.INIT('h8)
	) name6459 (
		_w3761_,
		_w8208_,
		_w8209_
	);
	LUT3 #(
		.INIT('h80)
	) name6460 (
		\u4_u0_buf1_reg[5]/P0001 ,
		_w3755_,
		_w3756_,
		_w8210_
	);
	LUT3 #(
		.INIT('h07)
	) name6461 (
		\u4_u1_buf1_reg[5]/P0001 ,
		_w3768_,
		_w8210_,
		_w8211_
	);
	LUT3 #(
		.INIT('h80)
	) name6462 (
		\u4_u3_buf1_reg[5]/P0001 ,
		_w3761_,
		_w3773_,
		_w8212_
	);
	LUT3 #(
		.INIT('h80)
	) name6463 (
		\u4_buf1_reg[5]/P0001 ,
		_w3761_,
		_w3775_,
		_w8213_
	);
	LUT4 #(
		.INIT('hfffb)
	) name6464 (
		_w8209_,
		_w8211_,
		_w8212_,
		_w8213_,
		_w8214_
	);
	LUT3 #(
		.INIT('h80)
	) name6465 (
		\u4_u2_csr1_reg[2]/P0001 ,
		_w3762_,
		_w3763_,
		_w8215_
	);
	LUT2 #(
		.INIT('h8)
	) name6466 (
		_w3761_,
		_w8215_,
		_w8216_
	);
	LUT3 #(
		.INIT('h80)
	) name6467 (
		\u4_u0_csr1_reg[2]/P0001 ,
		_w3755_,
		_w3756_,
		_w8217_
	);
	LUT3 #(
		.INIT('h07)
	) name6468 (
		\u4_u1_csr1_reg[2]/P0001 ,
		_w3768_,
		_w8217_,
		_w8218_
	);
	LUT3 #(
		.INIT('h80)
	) name6469 (
		\u4_u3_csr1_reg[2]/P0001 ,
		_w3761_,
		_w3773_,
		_w8219_
	);
	LUT3 #(
		.INIT('h80)
	) name6470 (
		\u4_csr_reg[17]/P0001 ,
		_w3761_,
		_w3775_,
		_w8220_
	);
	LUT4 #(
		.INIT('hfffb)
	) name6471 (
		_w8216_,
		_w8218_,
		_w8219_,
		_w8220_,
		_w8221_
	);
	LUT3 #(
		.INIT('h80)
	) name6472 (
		\u4_u2_csr0_reg[1]/P0001 ,
		_w3762_,
		_w3763_,
		_w8222_
	);
	LUT2 #(
		.INIT('h8)
	) name6473 (
		_w3761_,
		_w8222_,
		_w8223_
	);
	LUT3 #(
		.INIT('h80)
	) name6474 (
		\u4_u0_csr0_reg[1]/P0001 ,
		_w3755_,
		_w3756_,
		_w8224_
	);
	LUT3 #(
		.INIT('h07)
	) name6475 (
		\u4_u1_csr0_reg[1]/P0001 ,
		_w3768_,
		_w8224_,
		_w8225_
	);
	LUT3 #(
		.INIT('h80)
	) name6476 (
		\u4_u3_csr0_reg[1]/P0001 ,
		_w3761_,
		_w3773_,
		_w8226_
	);
	LUT3 #(
		.INIT('h80)
	) name6477 (
		\u4_csr_reg[1]/P0001 ,
		_w3761_,
		_w3775_,
		_w8227_
	);
	LUT4 #(
		.INIT('hfffb)
	) name6478 (
		_w8223_,
		_w8225_,
		_w8226_,
		_w8227_,
		_w8228_
	);
	LUT3 #(
		.INIT('h80)
	) name6479 (
		\u4_u2_csr1_reg[7]/P0001 ,
		_w3762_,
		_w3763_,
		_w8229_
	);
	LUT2 #(
		.INIT('h8)
	) name6480 (
		_w3761_,
		_w8229_,
		_w8230_
	);
	LUT3 #(
		.INIT('h80)
	) name6481 (
		\u4_u0_csr1_reg[7]/P0001 ,
		_w3755_,
		_w3756_,
		_w8231_
	);
	LUT3 #(
		.INIT('h07)
	) name6482 (
		\u4_u1_csr1_reg[7]/P0001 ,
		_w3768_,
		_w8231_,
		_w8232_
	);
	LUT3 #(
		.INIT('h80)
	) name6483 (
		\u4_u3_csr1_reg[7]/P0001 ,
		_w3761_,
		_w3773_,
		_w8233_
	);
	LUT3 #(
		.INIT('h80)
	) name6484 (
		\u4_csr_reg[22]/P0001 ,
		_w3761_,
		_w3775_,
		_w8234_
	);
	LUT4 #(
		.INIT('hfffb)
	) name6485 (
		_w8230_,
		_w8232_,
		_w8233_,
		_w8234_,
		_w8235_
	);
	LUT3 #(
		.INIT('h80)
	) name6486 (
		\u4_u2_csr1_reg[8]/P0001 ,
		_w3762_,
		_w3763_,
		_w8236_
	);
	LUT2 #(
		.INIT('h8)
	) name6487 (
		_w3761_,
		_w8236_,
		_w8237_
	);
	LUT3 #(
		.INIT('h80)
	) name6488 (
		\u4_u0_csr1_reg[8]/P0001 ,
		_w3755_,
		_w3756_,
		_w8238_
	);
	LUT3 #(
		.INIT('h07)
	) name6489 (
		\u4_u1_csr1_reg[8]/P0001 ,
		_w3768_,
		_w8238_,
		_w8239_
	);
	LUT3 #(
		.INIT('h80)
	) name6490 (
		\u4_u3_csr1_reg[8]/P0001 ,
		_w3761_,
		_w3773_,
		_w8240_
	);
	LUT3 #(
		.INIT('h80)
	) name6491 (
		\u4_csr_reg[23]/P0001 ,
		_w3761_,
		_w3775_,
		_w8241_
	);
	LUT4 #(
		.INIT('hfffb)
	) name6492 (
		_w8237_,
		_w8239_,
		_w8240_,
		_w8241_,
		_w8242_
	);
	LUT3 #(
		.INIT('h80)
	) name6493 (
		\u4_u2_csr1_reg[9]/P0001 ,
		_w3762_,
		_w3763_,
		_w8243_
	);
	LUT2 #(
		.INIT('h8)
	) name6494 (
		_w3761_,
		_w8243_,
		_w8244_
	);
	LUT3 #(
		.INIT('h80)
	) name6495 (
		\u4_u0_csr1_reg[9]/P0001 ,
		_w3755_,
		_w3756_,
		_w8245_
	);
	LUT3 #(
		.INIT('h07)
	) name6496 (
		\u4_u1_csr1_reg[9]/P0001 ,
		_w3768_,
		_w8245_,
		_w8246_
	);
	LUT3 #(
		.INIT('h80)
	) name6497 (
		\u4_u3_csr1_reg[9]/P0001 ,
		_w3761_,
		_w3773_,
		_w8247_
	);
	LUT3 #(
		.INIT('h80)
	) name6498 (
		\u4_csr_reg[24]/P0001 ,
		_w3761_,
		_w3775_,
		_w8248_
	);
	LUT4 #(
		.INIT('hfffb)
	) name6499 (
		_w8244_,
		_w8246_,
		_w8247_,
		_w8248_,
		_w8249_
	);
	LUT3 #(
		.INIT('h80)
	) name6500 (
		\u4_u2_csr1_reg[10]/P0001 ,
		_w3762_,
		_w3763_,
		_w8250_
	);
	LUT2 #(
		.INIT('h8)
	) name6501 (
		_w3761_,
		_w8250_,
		_w8251_
	);
	LUT3 #(
		.INIT('h80)
	) name6502 (
		\u4_u0_csr1_reg[10]/P0001 ,
		_w3755_,
		_w3756_,
		_w8252_
	);
	LUT3 #(
		.INIT('h07)
	) name6503 (
		\u4_u1_csr1_reg[10]/P0001 ,
		_w3768_,
		_w8252_,
		_w8253_
	);
	LUT3 #(
		.INIT('h80)
	) name6504 (
		\u4_u3_csr1_reg[10]/P0001 ,
		_w3761_,
		_w3773_,
		_w8254_
	);
	LUT3 #(
		.INIT('h80)
	) name6505 (
		\u4_csr_reg[25]/P0001 ,
		_w3761_,
		_w3775_,
		_w8255_
	);
	LUT4 #(
		.INIT('hfffb)
	) name6506 (
		_w8251_,
		_w8253_,
		_w8254_,
		_w8255_,
		_w8256_
	);
	LUT3 #(
		.INIT('h80)
	) name6507 (
		\u4_u2_csr1_reg[11]/P0001 ,
		_w3762_,
		_w3763_,
		_w8257_
	);
	LUT2 #(
		.INIT('h8)
	) name6508 (
		_w3761_,
		_w8257_,
		_w8258_
	);
	LUT3 #(
		.INIT('h80)
	) name6509 (
		\u4_u0_csr1_reg[11]/P0001 ,
		_w3755_,
		_w3756_,
		_w8259_
	);
	LUT3 #(
		.INIT('h07)
	) name6510 (
		\u4_u1_csr1_reg[11]/P0001 ,
		_w3768_,
		_w8259_,
		_w8260_
	);
	LUT3 #(
		.INIT('h80)
	) name6511 (
		\u4_u3_csr1_reg[11]/P0001 ,
		_w3761_,
		_w3773_,
		_w8261_
	);
	LUT3 #(
		.INIT('h80)
	) name6512 (
		\u4_csr_reg[26]/NET0131 ,
		_w3761_,
		_w3775_,
		_w8262_
	);
	LUT4 #(
		.INIT('hfffb)
	) name6513 (
		_w8258_,
		_w8260_,
		_w8261_,
		_w8262_,
		_w8263_
	);
	LUT3 #(
		.INIT('h80)
	) name6514 (
		\u4_u2_csr1_reg[12]/P0001 ,
		_w3762_,
		_w3763_,
		_w8264_
	);
	LUT2 #(
		.INIT('h8)
	) name6515 (
		_w3761_,
		_w8264_,
		_w8265_
	);
	LUT3 #(
		.INIT('h80)
	) name6516 (
		\u4_u0_csr1_reg[12]/P0001 ,
		_w3755_,
		_w3756_,
		_w8266_
	);
	LUT3 #(
		.INIT('h07)
	) name6517 (
		\u4_u1_csr1_reg[12]/P0001 ,
		_w3768_,
		_w8266_,
		_w8267_
	);
	LUT3 #(
		.INIT('h80)
	) name6518 (
		\u4_u3_csr1_reg[12]/P0001 ,
		_w3761_,
		_w3773_,
		_w8268_
	);
	LUT3 #(
		.INIT('h80)
	) name6519 (
		\u4_csr_reg[27]/NET0131 ,
		_w3761_,
		_w3775_,
		_w8269_
	);
	LUT4 #(
		.INIT('hfffb)
	) name6520 (
		_w8265_,
		_w8267_,
		_w8268_,
		_w8269_,
		_w8270_
	);
	LUT3 #(
		.INIT('h80)
	) name6521 (
		\u4_u2_uc_dpd_reg[0]/P0001 ,
		_w3762_,
		_w3763_,
		_w8271_
	);
	LUT2 #(
		.INIT('h8)
	) name6522 (
		_w3761_,
		_w8271_,
		_w8272_
	);
	LUT3 #(
		.INIT('h80)
	) name6523 (
		\u4_u0_uc_dpd_reg[0]/P0001 ,
		_w3755_,
		_w3756_,
		_w8273_
	);
	LUT3 #(
		.INIT('h07)
	) name6524 (
		\u4_u1_uc_dpd_reg[0]/P0001 ,
		_w3768_,
		_w8273_,
		_w8274_
	);
	LUT3 #(
		.INIT('h80)
	) name6525 (
		\u4_u3_uc_dpd_reg[0]/P0001 ,
		_w3761_,
		_w3773_,
		_w8275_
	);
	LUT3 #(
		.INIT('h80)
	) name6526 (
		\u4_csr_reg[28]/P0001 ,
		_w3761_,
		_w3775_,
		_w8276_
	);
	LUT4 #(
		.INIT('hfffb)
	) name6527 (
		_w8272_,
		_w8274_,
		_w8275_,
		_w8276_,
		_w8277_
	);
	LUT3 #(
		.INIT('h80)
	) name6528 (
		\u4_u2_uc_dpd_reg[1]/P0001 ,
		_w3762_,
		_w3763_,
		_w8278_
	);
	LUT2 #(
		.INIT('h8)
	) name6529 (
		_w3761_,
		_w8278_,
		_w8279_
	);
	LUT3 #(
		.INIT('h80)
	) name6530 (
		\u4_u0_uc_dpd_reg[1]/P0001 ,
		_w3755_,
		_w3756_,
		_w8280_
	);
	LUT3 #(
		.INIT('h07)
	) name6531 (
		\u4_u1_uc_dpd_reg[1]/P0001 ,
		_w3768_,
		_w8280_,
		_w8281_
	);
	LUT3 #(
		.INIT('h80)
	) name6532 (
		\u4_u3_uc_dpd_reg[1]/P0001 ,
		_w3761_,
		_w3773_,
		_w8282_
	);
	LUT3 #(
		.INIT('h80)
	) name6533 (
		\u4_csr_reg[29]/P0001 ,
		_w3761_,
		_w3775_,
		_w8283_
	);
	LUT4 #(
		.INIT('hfffb)
	) name6534 (
		_w8279_,
		_w8281_,
		_w8282_,
		_w8283_,
		_w8284_
	);
	LUT3 #(
		.INIT('h80)
	) name6535 (
		\u4_u2_csr0_reg[2]/P0001 ,
		_w3762_,
		_w3763_,
		_w8285_
	);
	LUT2 #(
		.INIT('h8)
	) name6536 (
		_w3761_,
		_w8285_,
		_w8286_
	);
	LUT3 #(
		.INIT('h80)
	) name6537 (
		\u4_u0_csr0_reg[2]/P0001 ,
		_w3755_,
		_w3756_,
		_w8287_
	);
	LUT3 #(
		.INIT('h07)
	) name6538 (
		\u4_u1_csr0_reg[2]/P0001 ,
		_w3768_,
		_w8287_,
		_w8288_
	);
	LUT3 #(
		.INIT('h80)
	) name6539 (
		\u4_u3_csr0_reg[2]/P0001 ,
		_w3761_,
		_w3773_,
		_w8289_
	);
	LUT3 #(
		.INIT('h80)
	) name6540 (
		\u4_csr_reg[2]/NET0131 ,
		_w3761_,
		_w3775_,
		_w8290_
	);
	LUT4 #(
		.INIT('hfffb)
	) name6541 (
		_w8286_,
		_w8288_,
		_w8289_,
		_w8290_,
		_w8291_
	);
	LUT3 #(
		.INIT('h80)
	) name6542 (
		\u4_u2_uc_bsel_reg[0]/P0001 ,
		_w3762_,
		_w3763_,
		_w8292_
	);
	LUT2 #(
		.INIT('h8)
	) name6543 (
		_w3761_,
		_w8292_,
		_w8293_
	);
	LUT3 #(
		.INIT('h80)
	) name6544 (
		\u4_u0_uc_bsel_reg[0]/P0001 ,
		_w3755_,
		_w3756_,
		_w8294_
	);
	LUT3 #(
		.INIT('h07)
	) name6545 (
		\u4_u1_uc_bsel_reg[0]/P0001 ,
		_w3768_,
		_w8294_,
		_w8295_
	);
	LUT3 #(
		.INIT('h80)
	) name6546 (
		\u4_u3_uc_bsel_reg[0]/P0001 ,
		_w3761_,
		_w3773_,
		_w8296_
	);
	LUT3 #(
		.INIT('h80)
	) name6547 (
		\u4_csr_reg[30]/NET0131 ,
		_w3761_,
		_w3775_,
		_w8297_
	);
	LUT4 #(
		.INIT('hfffb)
	) name6548 (
		_w8293_,
		_w8295_,
		_w8296_,
		_w8297_,
		_w8298_
	);
	LUT3 #(
		.INIT('h80)
	) name6549 (
		\u4_u2_uc_bsel_reg[1]/P0001 ,
		_w3762_,
		_w3763_,
		_w8299_
	);
	LUT2 #(
		.INIT('h8)
	) name6550 (
		_w3761_,
		_w8299_,
		_w8300_
	);
	LUT3 #(
		.INIT('h80)
	) name6551 (
		\u4_u0_uc_bsel_reg[1]/P0001 ,
		_w3755_,
		_w3756_,
		_w8301_
	);
	LUT3 #(
		.INIT('h07)
	) name6552 (
		\u4_u1_uc_bsel_reg[1]/P0001 ,
		_w3768_,
		_w8301_,
		_w8302_
	);
	LUT3 #(
		.INIT('h80)
	) name6553 (
		\u4_u3_uc_bsel_reg[1]/P0001 ,
		_w3761_,
		_w3773_,
		_w8303_
	);
	LUT3 #(
		.INIT('h80)
	) name6554 (
		\u4_csr_reg[31]/P0001 ,
		_w3761_,
		_w3775_,
		_w8304_
	);
	LUT4 #(
		.INIT('hfffb)
	) name6555 (
		_w8300_,
		_w8302_,
		_w8303_,
		_w8304_,
		_w8305_
	);
	LUT3 #(
		.INIT('h80)
	) name6556 (
		\u4_u2_csr0_reg[3]/NET0131 ,
		_w3762_,
		_w3763_,
		_w8306_
	);
	LUT2 #(
		.INIT('h8)
	) name6557 (
		_w3761_,
		_w8306_,
		_w8307_
	);
	LUT3 #(
		.INIT('h80)
	) name6558 (
		\u4_u0_csr0_reg[3]/NET0131 ,
		_w3755_,
		_w3756_,
		_w8308_
	);
	LUT3 #(
		.INIT('h07)
	) name6559 (
		\u4_u1_csr0_reg[3]/NET0131 ,
		_w3768_,
		_w8308_,
		_w8309_
	);
	LUT3 #(
		.INIT('h80)
	) name6560 (
		\u4_u3_csr0_reg[3]/NET0131 ,
		_w3761_,
		_w3773_,
		_w8310_
	);
	LUT3 #(
		.INIT('h80)
	) name6561 (
		\u4_csr_reg[3]/P0001 ,
		_w3761_,
		_w3775_,
		_w8311_
	);
	LUT4 #(
		.INIT('hfffb)
	) name6562 (
		_w8307_,
		_w8309_,
		_w8310_,
		_w8311_,
		_w8312_
	);
	LUT3 #(
		.INIT('h80)
	) name6563 (
		\u4_u2_csr0_reg[4]/P0001 ,
		_w3762_,
		_w3763_,
		_w8313_
	);
	LUT2 #(
		.INIT('h8)
	) name6564 (
		_w3761_,
		_w8313_,
		_w8314_
	);
	LUT3 #(
		.INIT('h80)
	) name6565 (
		\u4_u0_csr0_reg[4]/P0001 ,
		_w3755_,
		_w3756_,
		_w8315_
	);
	LUT3 #(
		.INIT('h07)
	) name6566 (
		\u4_u1_csr0_reg[4]/P0001 ,
		_w3768_,
		_w8315_,
		_w8316_
	);
	LUT3 #(
		.INIT('h80)
	) name6567 (
		\u4_u3_csr0_reg[4]/P0001 ,
		_w3761_,
		_w3773_,
		_w8317_
	);
	LUT3 #(
		.INIT('h80)
	) name6568 (
		\u4_csr_reg[4]/NET0131 ,
		_w3761_,
		_w3775_,
		_w8318_
	);
	LUT4 #(
		.INIT('hfffb)
	) name6569 (
		_w8314_,
		_w8316_,
		_w8317_,
		_w8318_,
		_w8319_
	);
	LUT3 #(
		.INIT('h80)
	) name6570 (
		\u4_u2_csr0_reg[5]/P0001 ,
		_w3762_,
		_w3763_,
		_w8320_
	);
	LUT2 #(
		.INIT('h8)
	) name6571 (
		_w3761_,
		_w8320_,
		_w8321_
	);
	LUT3 #(
		.INIT('h80)
	) name6572 (
		\u4_u0_csr0_reg[5]/P0001 ,
		_w3755_,
		_w3756_,
		_w8322_
	);
	LUT3 #(
		.INIT('h07)
	) name6573 (
		\u4_u1_csr0_reg[5]/P0001 ,
		_w3768_,
		_w8322_,
		_w8323_
	);
	LUT3 #(
		.INIT('h80)
	) name6574 (
		\u4_u3_csr0_reg[5]/P0001 ,
		_w3761_,
		_w3773_,
		_w8324_
	);
	LUT3 #(
		.INIT('h80)
	) name6575 (
		\u4_csr_reg[5]/NET0131 ,
		_w3761_,
		_w3775_,
		_w8325_
	);
	LUT4 #(
		.INIT('hfffb)
	) name6576 (
		_w8321_,
		_w8323_,
		_w8324_,
		_w8325_,
		_w8326_
	);
	LUT3 #(
		.INIT('h80)
	) name6577 (
		\u4_u2_csr0_reg[6]/P0001 ,
		_w3762_,
		_w3763_,
		_w8327_
	);
	LUT2 #(
		.INIT('h8)
	) name6578 (
		_w3761_,
		_w8327_,
		_w8328_
	);
	LUT3 #(
		.INIT('h80)
	) name6579 (
		\u4_u0_csr0_reg[6]/P0001 ,
		_w3755_,
		_w3756_,
		_w8329_
	);
	LUT3 #(
		.INIT('h07)
	) name6580 (
		\u4_u1_csr0_reg[6]/P0001 ,
		_w3768_,
		_w8329_,
		_w8330_
	);
	LUT3 #(
		.INIT('h80)
	) name6581 (
		\u4_u3_csr0_reg[6]/P0001 ,
		_w3761_,
		_w3773_,
		_w8331_
	);
	LUT3 #(
		.INIT('h80)
	) name6582 (
		\u4_csr_reg[6]/NET0131 ,
		_w3761_,
		_w3775_,
		_w8332_
	);
	LUT4 #(
		.INIT('hfffb)
	) name6583 (
		_w8328_,
		_w8330_,
		_w8331_,
		_w8332_,
		_w8333_
	);
	LUT3 #(
		.INIT('h80)
	) name6584 (
		\u4_u2_csr0_reg[7]/P0001 ,
		_w3762_,
		_w3763_,
		_w8334_
	);
	LUT2 #(
		.INIT('h8)
	) name6585 (
		_w3761_,
		_w8334_,
		_w8335_
	);
	LUT3 #(
		.INIT('h80)
	) name6586 (
		\u4_u0_csr0_reg[7]/P0001 ,
		_w3755_,
		_w3756_,
		_w8336_
	);
	LUT3 #(
		.INIT('h07)
	) name6587 (
		\u4_u1_csr0_reg[7]/P0001 ,
		_w3768_,
		_w8336_,
		_w8337_
	);
	LUT3 #(
		.INIT('h80)
	) name6588 (
		\u4_u3_csr0_reg[7]/P0001 ,
		_w3761_,
		_w3773_,
		_w8338_
	);
	LUT3 #(
		.INIT('h80)
	) name6589 (
		\u4_csr_reg[7]/P0001 ,
		_w3761_,
		_w3775_,
		_w8339_
	);
	LUT4 #(
		.INIT('hfffb)
	) name6590 (
		_w8335_,
		_w8337_,
		_w8338_,
		_w8339_,
		_w8340_
	);
	LUT3 #(
		.INIT('h80)
	) name6591 (
		\u4_u2_csr0_reg[8]/P0001 ,
		_w3762_,
		_w3763_,
		_w8341_
	);
	LUT2 #(
		.INIT('h8)
	) name6592 (
		_w3761_,
		_w8341_,
		_w8342_
	);
	LUT3 #(
		.INIT('h80)
	) name6593 (
		\u4_u0_csr0_reg[8]/P0001 ,
		_w3755_,
		_w3756_,
		_w8343_
	);
	LUT3 #(
		.INIT('h07)
	) name6594 (
		\u4_u1_csr0_reg[8]/P0001 ,
		_w3768_,
		_w8343_,
		_w8344_
	);
	LUT3 #(
		.INIT('h80)
	) name6595 (
		\u4_u3_csr0_reg[8]/P0001 ,
		_w3761_,
		_w3773_,
		_w8345_
	);
	LUT3 #(
		.INIT('h80)
	) name6596 (
		\u4_csr_reg[8]/P0001 ,
		_w3761_,
		_w3775_,
		_w8346_
	);
	LUT4 #(
		.INIT('hfffb)
	) name6597 (
		_w8342_,
		_w8344_,
		_w8345_,
		_w8346_,
		_w8347_
	);
	LUT3 #(
		.INIT('h80)
	) name6598 (
		\u4_u2_csr0_reg[9]/P0001 ,
		_w3762_,
		_w3763_,
		_w8348_
	);
	LUT2 #(
		.INIT('h8)
	) name6599 (
		_w3761_,
		_w8348_,
		_w8349_
	);
	LUT3 #(
		.INIT('h80)
	) name6600 (
		\u4_u0_csr0_reg[9]/P0001 ,
		_w3755_,
		_w3756_,
		_w8350_
	);
	LUT3 #(
		.INIT('h07)
	) name6601 (
		\u4_u1_csr0_reg[9]/P0001 ,
		_w3768_,
		_w8350_,
		_w8351_
	);
	LUT3 #(
		.INIT('h80)
	) name6602 (
		\u4_u3_csr0_reg[9]/P0001 ,
		_w3761_,
		_w3773_,
		_w8352_
	);
	LUT3 #(
		.INIT('h80)
	) name6603 (
		\u4_csr_reg[9]/NET0131 ,
		_w3761_,
		_w3775_,
		_w8353_
	);
	LUT4 #(
		.INIT('hfffb)
	) name6604 (
		_w8349_,
		_w8351_,
		_w8352_,
		_w8353_,
		_w8354_
	);
	LUT3 #(
		.INIT('h80)
	) name6605 (
		\u4_u2_buf1_reg[24]/P0001 ,
		_w3762_,
		_w3763_,
		_w8355_
	);
	LUT2 #(
		.INIT('h8)
	) name6606 (
		_w3761_,
		_w8355_,
		_w8356_
	);
	LUT3 #(
		.INIT('h80)
	) name6607 (
		\u4_u0_buf1_reg[24]/P0001 ,
		_w3755_,
		_w3756_,
		_w8357_
	);
	LUT3 #(
		.INIT('h07)
	) name6608 (
		\u4_u1_buf1_reg[24]/P0001 ,
		_w3768_,
		_w8357_,
		_w8358_
	);
	LUT3 #(
		.INIT('h80)
	) name6609 (
		\u4_u3_buf1_reg[24]/P0001 ,
		_w3761_,
		_w3773_,
		_w8359_
	);
	LUT3 #(
		.INIT('h80)
	) name6610 (
		\u4_buf1_reg[24]/NET0131 ,
		_w3761_,
		_w3775_,
		_w8360_
	);
	LUT4 #(
		.INIT('hfffb)
	) name6611 (
		_w8356_,
		_w8358_,
		_w8359_,
		_w8360_,
		_w8361_
	);
	LUT3 #(
		.INIT('h80)
	) name6612 (
		\u4_u2_buf0_reg[0]/P0001 ,
		_w3762_,
		_w3763_,
		_w8362_
	);
	LUT2 #(
		.INIT('h8)
	) name6613 (
		_w3761_,
		_w8362_,
		_w8363_
	);
	LUT3 #(
		.INIT('h80)
	) name6614 (
		\u4_u0_buf0_reg[0]/P0001 ,
		_w3755_,
		_w3756_,
		_w8364_
	);
	LUT3 #(
		.INIT('h07)
	) name6615 (
		\u4_u1_buf0_reg[0]/P0001 ,
		_w3768_,
		_w8364_,
		_w8365_
	);
	LUT3 #(
		.INIT('h80)
	) name6616 (
		\u4_u3_buf0_reg[0]/P0001 ,
		_w3761_,
		_w3773_,
		_w8366_
	);
	LUT3 #(
		.INIT('h80)
	) name6617 (
		\u4_buf0_reg[0]/P0001 ,
		_w3761_,
		_w3775_,
		_w8367_
	);
	LUT4 #(
		.INIT('hfffb)
	) name6618 (
		_w8363_,
		_w8365_,
		_w8366_,
		_w8367_,
		_w8368_
	);
	LUT3 #(
		.INIT('h80)
	) name6619 (
		\u4_u2_buf0_reg[10]/P0001 ,
		_w3762_,
		_w3763_,
		_w8369_
	);
	LUT2 #(
		.INIT('h8)
	) name6620 (
		_w3761_,
		_w8369_,
		_w8370_
	);
	LUT3 #(
		.INIT('h80)
	) name6621 (
		\u4_u0_buf0_reg[10]/P0001 ,
		_w3755_,
		_w3756_,
		_w8371_
	);
	LUT3 #(
		.INIT('h07)
	) name6622 (
		\u4_u1_buf0_reg[10]/P0001 ,
		_w3768_,
		_w8371_,
		_w8372_
	);
	LUT3 #(
		.INIT('h80)
	) name6623 (
		\u4_u3_buf0_reg[10]/P0001 ,
		_w3761_,
		_w3773_,
		_w8373_
	);
	LUT3 #(
		.INIT('h80)
	) name6624 (
		\u4_buf0_reg[10]/P0001 ,
		_w3761_,
		_w3775_,
		_w8374_
	);
	LUT4 #(
		.INIT('hfffb)
	) name6625 (
		_w8370_,
		_w8372_,
		_w8373_,
		_w8374_,
		_w8375_
	);
	LUT3 #(
		.INIT('h80)
	) name6626 (
		\u4_u2_buf0_reg[11]/P0001 ,
		_w3762_,
		_w3763_,
		_w8376_
	);
	LUT2 #(
		.INIT('h8)
	) name6627 (
		_w3761_,
		_w8376_,
		_w8377_
	);
	LUT3 #(
		.INIT('h80)
	) name6628 (
		\u4_u0_buf0_reg[11]/P0001 ,
		_w3755_,
		_w3756_,
		_w8378_
	);
	LUT3 #(
		.INIT('h07)
	) name6629 (
		\u4_u1_buf0_reg[11]/P0001 ,
		_w3768_,
		_w8378_,
		_w8379_
	);
	LUT3 #(
		.INIT('h80)
	) name6630 (
		\u4_u3_buf0_reg[11]/P0001 ,
		_w3761_,
		_w3773_,
		_w8380_
	);
	LUT3 #(
		.INIT('h80)
	) name6631 (
		\u4_buf0_reg[11]/P0001 ,
		_w3761_,
		_w3775_,
		_w8381_
	);
	LUT4 #(
		.INIT('hfffb)
	) name6632 (
		_w8377_,
		_w8379_,
		_w8380_,
		_w8381_,
		_w8382_
	);
	LUT3 #(
		.INIT('h80)
	) name6633 (
		\u4_u2_buf0_reg[12]/P0001 ,
		_w3762_,
		_w3763_,
		_w8383_
	);
	LUT2 #(
		.INIT('h8)
	) name6634 (
		_w3761_,
		_w8383_,
		_w8384_
	);
	LUT3 #(
		.INIT('h80)
	) name6635 (
		\u4_u0_buf0_reg[12]/P0001 ,
		_w3755_,
		_w3756_,
		_w8385_
	);
	LUT3 #(
		.INIT('h07)
	) name6636 (
		\u4_u1_buf0_reg[12]/P0001 ,
		_w3768_,
		_w8385_,
		_w8386_
	);
	LUT3 #(
		.INIT('h80)
	) name6637 (
		\u4_u3_buf0_reg[12]/P0001 ,
		_w3761_,
		_w3773_,
		_w8387_
	);
	LUT3 #(
		.INIT('h80)
	) name6638 (
		\u4_buf0_reg[12]/P0001 ,
		_w3761_,
		_w3775_,
		_w8388_
	);
	LUT4 #(
		.INIT('hfffb)
	) name6639 (
		_w8384_,
		_w8386_,
		_w8387_,
		_w8388_,
		_w8389_
	);
	LUT3 #(
		.INIT('h80)
	) name6640 (
		\u4_u2_buf0_reg[13]/P0001 ,
		_w3762_,
		_w3763_,
		_w8390_
	);
	LUT2 #(
		.INIT('h8)
	) name6641 (
		_w3761_,
		_w8390_,
		_w8391_
	);
	LUT3 #(
		.INIT('h80)
	) name6642 (
		\u4_u0_buf0_reg[13]/P0001 ,
		_w3755_,
		_w3756_,
		_w8392_
	);
	LUT3 #(
		.INIT('h07)
	) name6643 (
		\u4_u1_buf0_reg[13]/P0001 ,
		_w3768_,
		_w8392_,
		_w8393_
	);
	LUT3 #(
		.INIT('h80)
	) name6644 (
		\u4_u3_buf0_reg[13]/P0001 ,
		_w3761_,
		_w3773_,
		_w8394_
	);
	LUT3 #(
		.INIT('h80)
	) name6645 (
		\u4_buf0_reg[13]/P0001 ,
		_w3761_,
		_w3775_,
		_w8395_
	);
	LUT4 #(
		.INIT('hfffb)
	) name6646 (
		_w8391_,
		_w8393_,
		_w8394_,
		_w8395_,
		_w8396_
	);
	LUT3 #(
		.INIT('h80)
	) name6647 (
		\u4_u2_buf0_reg[14]/P0001 ,
		_w3762_,
		_w3763_,
		_w8397_
	);
	LUT2 #(
		.INIT('h8)
	) name6648 (
		_w3761_,
		_w8397_,
		_w8398_
	);
	LUT3 #(
		.INIT('h80)
	) name6649 (
		\u4_u0_buf0_reg[14]/P0001 ,
		_w3755_,
		_w3756_,
		_w8399_
	);
	LUT3 #(
		.INIT('h07)
	) name6650 (
		\u4_u1_buf0_reg[14]/P0001 ,
		_w3768_,
		_w8399_,
		_w8400_
	);
	LUT3 #(
		.INIT('h80)
	) name6651 (
		\u4_u3_buf0_reg[14]/P0001 ,
		_w3761_,
		_w3773_,
		_w8401_
	);
	LUT3 #(
		.INIT('h80)
	) name6652 (
		\u4_buf0_reg[14]/P0001 ,
		_w3761_,
		_w3775_,
		_w8402_
	);
	LUT4 #(
		.INIT('hfffb)
	) name6653 (
		_w8398_,
		_w8400_,
		_w8401_,
		_w8402_,
		_w8403_
	);
	LUT3 #(
		.INIT('h80)
	) name6654 (
		\u4_u2_buf0_reg[15]/P0001 ,
		_w3762_,
		_w3763_,
		_w8404_
	);
	LUT2 #(
		.INIT('h8)
	) name6655 (
		_w3761_,
		_w8404_,
		_w8405_
	);
	LUT3 #(
		.INIT('h80)
	) name6656 (
		\u4_u0_buf0_reg[15]/P0001 ,
		_w3755_,
		_w3756_,
		_w8406_
	);
	LUT3 #(
		.INIT('h07)
	) name6657 (
		\u4_u1_buf0_reg[15]/P0001 ,
		_w3768_,
		_w8406_,
		_w8407_
	);
	LUT3 #(
		.INIT('h80)
	) name6658 (
		\u4_u3_buf0_reg[15]/P0001 ,
		_w3761_,
		_w3773_,
		_w8408_
	);
	LUT3 #(
		.INIT('h80)
	) name6659 (
		\u4_buf0_reg[15]/P0001 ,
		_w3761_,
		_w3775_,
		_w8409_
	);
	LUT4 #(
		.INIT('hfffb)
	) name6660 (
		_w8405_,
		_w8407_,
		_w8408_,
		_w8409_,
		_w8410_
	);
	LUT3 #(
		.INIT('h80)
	) name6661 (
		\u4_u2_buf0_reg[16]/P0001 ,
		_w3762_,
		_w3763_,
		_w8411_
	);
	LUT2 #(
		.INIT('h8)
	) name6662 (
		_w3761_,
		_w8411_,
		_w8412_
	);
	LUT3 #(
		.INIT('h80)
	) name6663 (
		\u4_u0_buf0_reg[16]/P0001 ,
		_w3755_,
		_w3756_,
		_w8413_
	);
	LUT3 #(
		.INIT('h07)
	) name6664 (
		\u4_u1_buf0_reg[16]/P0001 ,
		_w3768_,
		_w8413_,
		_w8414_
	);
	LUT3 #(
		.INIT('h80)
	) name6665 (
		\u4_u3_buf0_reg[16]/P0001 ,
		_w3761_,
		_w3773_,
		_w8415_
	);
	LUT3 #(
		.INIT('h80)
	) name6666 (
		\u4_buf0_reg[16]/P0001 ,
		_w3761_,
		_w3775_,
		_w8416_
	);
	LUT4 #(
		.INIT('hfffb)
	) name6667 (
		_w8412_,
		_w8414_,
		_w8415_,
		_w8416_,
		_w8417_
	);
	LUT3 #(
		.INIT('h80)
	) name6668 (
		\u4_u2_buf0_reg[17]/P0001 ,
		_w3762_,
		_w3763_,
		_w8418_
	);
	LUT2 #(
		.INIT('h8)
	) name6669 (
		_w3761_,
		_w8418_,
		_w8419_
	);
	LUT3 #(
		.INIT('h80)
	) name6670 (
		\u4_u0_buf0_reg[17]/P0001 ,
		_w3755_,
		_w3756_,
		_w8420_
	);
	LUT3 #(
		.INIT('h07)
	) name6671 (
		\u4_u1_buf0_reg[17]/P0001 ,
		_w3768_,
		_w8420_,
		_w8421_
	);
	LUT3 #(
		.INIT('h80)
	) name6672 (
		\u4_u3_buf0_reg[17]/P0001 ,
		_w3761_,
		_w3773_,
		_w8422_
	);
	LUT3 #(
		.INIT('h80)
	) name6673 (
		\u4_buf0_reg[17]/NET0131 ,
		_w3761_,
		_w3775_,
		_w8423_
	);
	LUT4 #(
		.INIT('hfffb)
	) name6674 (
		_w8419_,
		_w8421_,
		_w8422_,
		_w8423_,
		_w8424_
	);
	LUT3 #(
		.INIT('h80)
	) name6675 (
		\u4_u2_buf0_reg[18]/P0001 ,
		_w3762_,
		_w3763_,
		_w8425_
	);
	LUT2 #(
		.INIT('h8)
	) name6676 (
		_w3761_,
		_w8425_,
		_w8426_
	);
	LUT3 #(
		.INIT('h80)
	) name6677 (
		\u4_u0_buf0_reg[18]/P0001 ,
		_w3755_,
		_w3756_,
		_w8427_
	);
	LUT3 #(
		.INIT('h07)
	) name6678 (
		\u4_u1_buf0_reg[18]/P0001 ,
		_w3768_,
		_w8427_,
		_w8428_
	);
	LUT3 #(
		.INIT('h80)
	) name6679 (
		\u4_u3_buf0_reg[18]/P0001 ,
		_w3761_,
		_w3773_,
		_w8429_
	);
	LUT3 #(
		.INIT('h80)
	) name6680 (
		\u4_buf0_reg[18]/P0001 ,
		_w3761_,
		_w3775_,
		_w8430_
	);
	LUT4 #(
		.INIT('hfffb)
	) name6681 (
		_w8426_,
		_w8428_,
		_w8429_,
		_w8430_,
		_w8431_
	);
	LUT3 #(
		.INIT('h80)
	) name6682 (
		\u4_u2_buf0_reg[19]/P0001 ,
		_w3762_,
		_w3763_,
		_w8432_
	);
	LUT2 #(
		.INIT('h8)
	) name6683 (
		_w3761_,
		_w8432_,
		_w8433_
	);
	LUT3 #(
		.INIT('h80)
	) name6684 (
		\u4_u0_buf0_reg[19]/P0001 ,
		_w3755_,
		_w3756_,
		_w8434_
	);
	LUT3 #(
		.INIT('h07)
	) name6685 (
		\u4_u1_buf0_reg[19]/P0001 ,
		_w3768_,
		_w8434_,
		_w8435_
	);
	LUT3 #(
		.INIT('h80)
	) name6686 (
		\u4_u3_buf0_reg[19]/P0001 ,
		_w3761_,
		_w3773_,
		_w8436_
	);
	LUT3 #(
		.INIT('h80)
	) name6687 (
		\u4_buf0_reg[19]/NET0131 ,
		_w3761_,
		_w3775_,
		_w8437_
	);
	LUT4 #(
		.INIT('hfffb)
	) name6688 (
		_w8433_,
		_w8435_,
		_w8436_,
		_w8437_,
		_w8438_
	);
	LUT3 #(
		.INIT('h80)
	) name6689 (
		\u4_u2_buf1_reg[6]/P0001 ,
		_w3762_,
		_w3763_,
		_w8439_
	);
	LUT2 #(
		.INIT('h8)
	) name6690 (
		_w3761_,
		_w8439_,
		_w8440_
	);
	LUT3 #(
		.INIT('h80)
	) name6691 (
		\u4_u0_buf1_reg[6]/P0001 ,
		_w3755_,
		_w3756_,
		_w8441_
	);
	LUT3 #(
		.INIT('h07)
	) name6692 (
		\u4_u1_buf1_reg[6]/P0001 ,
		_w3768_,
		_w8441_,
		_w8442_
	);
	LUT3 #(
		.INIT('h80)
	) name6693 (
		\u4_u3_buf1_reg[6]/P0001 ,
		_w3761_,
		_w3773_,
		_w8443_
	);
	LUT3 #(
		.INIT('h80)
	) name6694 (
		\u4_buf1_reg[6]/P0001 ,
		_w3761_,
		_w3775_,
		_w8444_
	);
	LUT4 #(
		.INIT('hfffb)
	) name6695 (
		_w8440_,
		_w8442_,
		_w8443_,
		_w8444_,
		_w8445_
	);
	LUT3 #(
		.INIT('h80)
	) name6696 (
		\u4_u2_buf0_reg[1]/P0001 ,
		_w3762_,
		_w3763_,
		_w8446_
	);
	LUT2 #(
		.INIT('h8)
	) name6697 (
		_w3761_,
		_w8446_,
		_w8447_
	);
	LUT3 #(
		.INIT('h80)
	) name6698 (
		\u4_u0_buf0_reg[1]/P0001 ,
		_w3755_,
		_w3756_,
		_w8448_
	);
	LUT3 #(
		.INIT('h07)
	) name6699 (
		\u4_u1_buf0_reg[1]/P0001 ,
		_w3768_,
		_w8448_,
		_w8449_
	);
	LUT3 #(
		.INIT('h80)
	) name6700 (
		\u4_u3_buf0_reg[1]/P0001 ,
		_w3761_,
		_w3773_,
		_w8450_
	);
	LUT3 #(
		.INIT('h80)
	) name6701 (
		\u4_buf0_reg[1]/P0001 ,
		_w3761_,
		_w3775_,
		_w8451_
	);
	LUT4 #(
		.INIT('hfffb)
	) name6702 (
		_w8447_,
		_w8449_,
		_w8450_,
		_w8451_,
		_w8452_
	);
	LUT3 #(
		.INIT('h80)
	) name6703 (
		\u4_u2_buf0_reg[20]/P0001 ,
		_w3762_,
		_w3763_,
		_w8453_
	);
	LUT2 #(
		.INIT('h8)
	) name6704 (
		_w3761_,
		_w8453_,
		_w8454_
	);
	LUT3 #(
		.INIT('h80)
	) name6705 (
		\u4_u0_buf0_reg[20]/P0001 ,
		_w3755_,
		_w3756_,
		_w8455_
	);
	LUT3 #(
		.INIT('h07)
	) name6706 (
		\u4_u1_buf0_reg[20]/P0001 ,
		_w3768_,
		_w8455_,
		_w8456_
	);
	LUT3 #(
		.INIT('h80)
	) name6707 (
		\u4_u3_buf0_reg[20]/P0001 ,
		_w3761_,
		_w3773_,
		_w8457_
	);
	LUT3 #(
		.INIT('h80)
	) name6708 (
		\u4_buf0_reg[20]/NET0131 ,
		_w3761_,
		_w3775_,
		_w8458_
	);
	LUT4 #(
		.INIT('hfffb)
	) name6709 (
		_w8454_,
		_w8456_,
		_w8457_,
		_w8458_,
		_w8459_
	);
	LUT3 #(
		.INIT('h80)
	) name6710 (
		\u4_u2_buf0_reg[21]/P0001 ,
		_w3762_,
		_w3763_,
		_w8460_
	);
	LUT2 #(
		.INIT('h8)
	) name6711 (
		_w3761_,
		_w8460_,
		_w8461_
	);
	LUT3 #(
		.INIT('h80)
	) name6712 (
		\u4_u0_buf0_reg[21]/P0001 ,
		_w3755_,
		_w3756_,
		_w8462_
	);
	LUT3 #(
		.INIT('h07)
	) name6713 (
		\u4_u1_buf0_reg[21]/P0001 ,
		_w3768_,
		_w8462_,
		_w8463_
	);
	LUT3 #(
		.INIT('h80)
	) name6714 (
		\u4_u3_buf0_reg[21]/P0001 ,
		_w3761_,
		_w3773_,
		_w8464_
	);
	LUT3 #(
		.INIT('h80)
	) name6715 (
		\u4_buf0_reg[21]/NET0131 ,
		_w3761_,
		_w3775_,
		_w8465_
	);
	LUT4 #(
		.INIT('hfffb)
	) name6716 (
		_w8461_,
		_w8463_,
		_w8464_,
		_w8465_,
		_w8466_
	);
	LUT3 #(
		.INIT('h80)
	) name6717 (
		\u4_u2_buf0_reg[22]/P0001 ,
		_w3762_,
		_w3763_,
		_w8467_
	);
	LUT2 #(
		.INIT('h8)
	) name6718 (
		_w3761_,
		_w8467_,
		_w8468_
	);
	LUT3 #(
		.INIT('h80)
	) name6719 (
		\u4_u0_buf0_reg[22]/P0001 ,
		_w3755_,
		_w3756_,
		_w8469_
	);
	LUT3 #(
		.INIT('h07)
	) name6720 (
		\u4_u1_buf0_reg[22]/P0001 ,
		_w3768_,
		_w8469_,
		_w8470_
	);
	LUT3 #(
		.INIT('h80)
	) name6721 (
		\u4_u3_buf0_reg[22]/P0001 ,
		_w3761_,
		_w3773_,
		_w8471_
	);
	LUT3 #(
		.INIT('h80)
	) name6722 (
		\u4_buf0_reg[22]/NET0131 ,
		_w3761_,
		_w3775_,
		_w8472_
	);
	LUT4 #(
		.INIT('hfffb)
	) name6723 (
		_w8468_,
		_w8470_,
		_w8471_,
		_w8472_,
		_w8473_
	);
	LUT3 #(
		.INIT('h80)
	) name6724 (
		\u4_u2_buf0_reg[23]/P0001 ,
		_w3762_,
		_w3763_,
		_w8474_
	);
	LUT2 #(
		.INIT('h8)
	) name6725 (
		_w3761_,
		_w8474_,
		_w8475_
	);
	LUT3 #(
		.INIT('h80)
	) name6726 (
		\u4_u0_buf0_reg[23]/P0001 ,
		_w3755_,
		_w3756_,
		_w8476_
	);
	LUT3 #(
		.INIT('h07)
	) name6727 (
		\u4_u1_buf0_reg[23]/P0001 ,
		_w3768_,
		_w8476_,
		_w8477_
	);
	LUT3 #(
		.INIT('h80)
	) name6728 (
		\u4_u3_buf0_reg[23]/P0001 ,
		_w3761_,
		_w3773_,
		_w8478_
	);
	LUT3 #(
		.INIT('h80)
	) name6729 (
		\u4_buf0_reg[23]/NET0131 ,
		_w3761_,
		_w3775_,
		_w8479_
	);
	LUT4 #(
		.INIT('hfffb)
	) name6730 (
		_w8475_,
		_w8477_,
		_w8478_,
		_w8479_,
		_w8480_
	);
	LUT3 #(
		.INIT('h80)
	) name6731 (
		\u4_u2_buf0_reg[24]/P0001 ,
		_w3762_,
		_w3763_,
		_w8481_
	);
	LUT2 #(
		.INIT('h8)
	) name6732 (
		_w3761_,
		_w8481_,
		_w8482_
	);
	LUT3 #(
		.INIT('h80)
	) name6733 (
		\u4_u0_buf0_reg[24]/P0001 ,
		_w3755_,
		_w3756_,
		_w8483_
	);
	LUT3 #(
		.INIT('h07)
	) name6734 (
		\u4_u1_buf0_reg[24]/P0001 ,
		_w3768_,
		_w8483_,
		_w8484_
	);
	LUT3 #(
		.INIT('h80)
	) name6735 (
		\u4_u3_buf0_reg[24]/P0001 ,
		_w3761_,
		_w3773_,
		_w8485_
	);
	LUT3 #(
		.INIT('h80)
	) name6736 (
		\u4_buf0_reg[24]/NET0131 ,
		_w3761_,
		_w3775_,
		_w8486_
	);
	LUT4 #(
		.INIT('hfffb)
	) name6737 (
		_w8482_,
		_w8484_,
		_w8485_,
		_w8486_,
		_w8487_
	);
	LUT3 #(
		.INIT('h80)
	) name6738 (
		\u4_u2_buf0_reg[25]/P0001 ,
		_w3762_,
		_w3763_,
		_w8488_
	);
	LUT2 #(
		.INIT('h8)
	) name6739 (
		_w3761_,
		_w8488_,
		_w8489_
	);
	LUT3 #(
		.INIT('h80)
	) name6740 (
		\u4_u0_buf0_reg[25]/P0001 ,
		_w3755_,
		_w3756_,
		_w8490_
	);
	LUT3 #(
		.INIT('h07)
	) name6741 (
		\u4_u1_buf0_reg[25]/P0001 ,
		_w3768_,
		_w8490_,
		_w8491_
	);
	LUT3 #(
		.INIT('h80)
	) name6742 (
		\u4_u3_buf0_reg[25]/P0001 ,
		_w3761_,
		_w3773_,
		_w8492_
	);
	LUT3 #(
		.INIT('h80)
	) name6743 (
		\u4_buf0_reg[25]/NET0131 ,
		_w3761_,
		_w3775_,
		_w8493_
	);
	LUT4 #(
		.INIT('hfffb)
	) name6744 (
		_w8489_,
		_w8491_,
		_w8492_,
		_w8493_,
		_w8494_
	);
	LUT3 #(
		.INIT('h80)
	) name6745 (
		\u4_u2_buf0_reg[26]/P0001 ,
		_w3762_,
		_w3763_,
		_w8495_
	);
	LUT2 #(
		.INIT('h8)
	) name6746 (
		_w3761_,
		_w8495_,
		_w8496_
	);
	LUT3 #(
		.INIT('h80)
	) name6747 (
		\u4_u0_buf0_reg[26]/P0001 ,
		_w3755_,
		_w3756_,
		_w8497_
	);
	LUT3 #(
		.INIT('h07)
	) name6748 (
		\u4_u1_buf0_reg[26]/P0001 ,
		_w3768_,
		_w8497_,
		_w8498_
	);
	LUT3 #(
		.INIT('h80)
	) name6749 (
		\u4_u3_buf0_reg[26]/P0001 ,
		_w3761_,
		_w3773_,
		_w8499_
	);
	LUT3 #(
		.INIT('h80)
	) name6750 (
		\u4_buf0_reg[26]/NET0131 ,
		_w3761_,
		_w3775_,
		_w8500_
	);
	LUT4 #(
		.INIT('hfffb)
	) name6751 (
		_w8496_,
		_w8498_,
		_w8499_,
		_w8500_,
		_w8501_
	);
	LUT3 #(
		.INIT('h80)
	) name6752 (
		\u4_u2_buf0_reg[27]/P0001 ,
		_w3762_,
		_w3763_,
		_w8502_
	);
	LUT2 #(
		.INIT('h8)
	) name6753 (
		_w3761_,
		_w8502_,
		_w8503_
	);
	LUT3 #(
		.INIT('h80)
	) name6754 (
		\u4_u0_buf0_reg[27]/P0001 ,
		_w3755_,
		_w3756_,
		_w8504_
	);
	LUT3 #(
		.INIT('h07)
	) name6755 (
		\u4_u1_buf0_reg[27]/P0001 ,
		_w3768_,
		_w8504_,
		_w8505_
	);
	LUT3 #(
		.INIT('h80)
	) name6756 (
		\u4_u3_buf0_reg[27]/P0001 ,
		_w3761_,
		_w3773_,
		_w8506_
	);
	LUT3 #(
		.INIT('h80)
	) name6757 (
		\u4_buf0_reg[27]/P0001 ,
		_w3761_,
		_w3775_,
		_w8507_
	);
	LUT4 #(
		.INIT('hfffb)
	) name6758 (
		_w8503_,
		_w8505_,
		_w8506_,
		_w8507_,
		_w8508_
	);
	LUT3 #(
		.INIT('h80)
	) name6759 (
		\u4_u2_buf0_reg[28]/P0001 ,
		_w3762_,
		_w3763_,
		_w8509_
	);
	LUT2 #(
		.INIT('h8)
	) name6760 (
		_w3761_,
		_w8509_,
		_w8510_
	);
	LUT3 #(
		.INIT('h80)
	) name6761 (
		\u4_u0_buf0_reg[28]/P0001 ,
		_w3755_,
		_w3756_,
		_w8511_
	);
	LUT3 #(
		.INIT('h07)
	) name6762 (
		\u4_u1_buf0_reg[28]/P0001 ,
		_w3768_,
		_w8511_,
		_w8512_
	);
	LUT3 #(
		.INIT('h80)
	) name6763 (
		\u4_u3_buf0_reg[28]/P0001 ,
		_w3761_,
		_w3773_,
		_w8513_
	);
	LUT3 #(
		.INIT('h80)
	) name6764 (
		\u4_buf0_reg[28]/P0001 ,
		_w3761_,
		_w3775_,
		_w8514_
	);
	LUT4 #(
		.INIT('hfffb)
	) name6765 (
		_w8510_,
		_w8512_,
		_w8513_,
		_w8514_,
		_w8515_
	);
	LUT3 #(
		.INIT('h80)
	) name6766 (
		\u4_u2_buf0_reg[29]/P0001 ,
		_w3762_,
		_w3763_,
		_w8516_
	);
	LUT2 #(
		.INIT('h8)
	) name6767 (
		_w3761_,
		_w8516_,
		_w8517_
	);
	LUT3 #(
		.INIT('h80)
	) name6768 (
		\u4_u0_buf0_reg[29]/P0001 ,
		_w3755_,
		_w3756_,
		_w8518_
	);
	LUT3 #(
		.INIT('h07)
	) name6769 (
		\u4_u1_buf0_reg[29]/P0001 ,
		_w3768_,
		_w8518_,
		_w8519_
	);
	LUT3 #(
		.INIT('h80)
	) name6770 (
		\u4_u3_buf0_reg[29]/P0001 ,
		_w3761_,
		_w3773_,
		_w8520_
	);
	LUT3 #(
		.INIT('h80)
	) name6771 (
		\u4_buf0_reg[29]/P0001 ,
		_w3761_,
		_w3775_,
		_w8521_
	);
	LUT4 #(
		.INIT('hfffb)
	) name6772 (
		_w8517_,
		_w8519_,
		_w8520_,
		_w8521_,
		_w8522_
	);
	LUT3 #(
		.INIT('h80)
	) name6773 (
		\u4_u2_buf0_reg[2]/P0001 ,
		_w3762_,
		_w3763_,
		_w8523_
	);
	LUT2 #(
		.INIT('h8)
	) name6774 (
		_w3761_,
		_w8523_,
		_w8524_
	);
	LUT3 #(
		.INIT('h80)
	) name6775 (
		\u4_u0_buf0_reg[2]/P0001 ,
		_w3755_,
		_w3756_,
		_w8525_
	);
	LUT3 #(
		.INIT('h07)
	) name6776 (
		\u4_u1_buf0_reg[2]/P0001 ,
		_w3768_,
		_w8525_,
		_w8526_
	);
	LUT3 #(
		.INIT('h80)
	) name6777 (
		\u4_u3_buf0_reg[2]/P0001 ,
		_w3761_,
		_w3773_,
		_w8527_
	);
	LUT3 #(
		.INIT('h80)
	) name6778 (
		\u4_buf0_reg[2]/P0001 ,
		_w3761_,
		_w3775_,
		_w8528_
	);
	LUT4 #(
		.INIT('hfffb)
	) name6779 (
		_w8524_,
		_w8526_,
		_w8527_,
		_w8528_,
		_w8529_
	);
	LUT3 #(
		.INIT('h80)
	) name6780 (
		\u4_u2_buf0_reg[30]/P0001 ,
		_w3762_,
		_w3763_,
		_w8530_
	);
	LUT2 #(
		.INIT('h8)
	) name6781 (
		_w3761_,
		_w8530_,
		_w8531_
	);
	LUT3 #(
		.INIT('h80)
	) name6782 (
		\u4_u0_buf0_reg[30]/P0001 ,
		_w3755_,
		_w3756_,
		_w8532_
	);
	LUT3 #(
		.INIT('h07)
	) name6783 (
		\u4_u1_buf0_reg[30]/P0001 ,
		_w3768_,
		_w8532_,
		_w8533_
	);
	LUT3 #(
		.INIT('h80)
	) name6784 (
		\u4_u3_buf0_reg[30]/P0001 ,
		_w3761_,
		_w3773_,
		_w8534_
	);
	LUT3 #(
		.INIT('h80)
	) name6785 (
		\u4_buf0_reg[30]/P0001 ,
		_w3761_,
		_w3775_,
		_w8535_
	);
	LUT4 #(
		.INIT('hfffb)
	) name6786 (
		_w8531_,
		_w8533_,
		_w8534_,
		_w8535_,
		_w8536_
	);
	LUT3 #(
		.INIT('h80)
	) name6787 (
		\u4_u2_buf0_reg[31]/P0001 ,
		_w3762_,
		_w3763_,
		_w8537_
	);
	LUT2 #(
		.INIT('h8)
	) name6788 (
		_w3761_,
		_w8537_,
		_w8538_
	);
	LUT3 #(
		.INIT('h80)
	) name6789 (
		\u4_u0_buf0_reg[31]/P0001 ,
		_w3755_,
		_w3756_,
		_w8539_
	);
	LUT3 #(
		.INIT('h07)
	) name6790 (
		\u4_u1_buf0_reg[31]/P0001 ,
		_w3768_,
		_w8539_,
		_w8540_
	);
	LUT3 #(
		.INIT('h80)
	) name6791 (
		\u4_u3_buf0_reg[31]/P0001 ,
		_w3761_,
		_w3773_,
		_w8541_
	);
	LUT3 #(
		.INIT('h80)
	) name6792 (
		\u4_buf0_reg[31]/P0001 ,
		_w3761_,
		_w3775_,
		_w8542_
	);
	LUT4 #(
		.INIT('hfffb)
	) name6793 (
		_w8538_,
		_w8540_,
		_w8541_,
		_w8542_,
		_w8543_
	);
	LUT3 #(
		.INIT('h80)
	) name6794 (
		\u4_u2_buf0_reg[3]/P0001 ,
		_w3762_,
		_w3763_,
		_w8544_
	);
	LUT2 #(
		.INIT('h8)
	) name6795 (
		_w3761_,
		_w8544_,
		_w8545_
	);
	LUT3 #(
		.INIT('h80)
	) name6796 (
		\u4_u0_buf0_reg[3]/P0001 ,
		_w3755_,
		_w3756_,
		_w8546_
	);
	LUT3 #(
		.INIT('h07)
	) name6797 (
		\u4_u1_buf0_reg[3]/P0001 ,
		_w3768_,
		_w8546_,
		_w8547_
	);
	LUT3 #(
		.INIT('h80)
	) name6798 (
		\u4_u3_buf0_reg[3]/P0001 ,
		_w3761_,
		_w3773_,
		_w8548_
	);
	LUT3 #(
		.INIT('h80)
	) name6799 (
		\u4_buf0_reg[3]/P0001 ,
		_w3761_,
		_w3775_,
		_w8549_
	);
	LUT4 #(
		.INIT('hfffb)
	) name6800 (
		_w8545_,
		_w8547_,
		_w8548_,
		_w8549_,
		_w8550_
	);
	LUT3 #(
		.INIT('h80)
	) name6801 (
		\u4_u2_buf0_reg[4]/P0001 ,
		_w3762_,
		_w3763_,
		_w8551_
	);
	LUT2 #(
		.INIT('h8)
	) name6802 (
		_w3761_,
		_w8551_,
		_w8552_
	);
	LUT3 #(
		.INIT('h80)
	) name6803 (
		\u4_u0_buf0_reg[4]/P0001 ,
		_w3755_,
		_w3756_,
		_w8553_
	);
	LUT3 #(
		.INIT('h07)
	) name6804 (
		\u4_u1_buf0_reg[4]/P0001 ,
		_w3768_,
		_w8553_,
		_w8554_
	);
	LUT3 #(
		.INIT('h80)
	) name6805 (
		\u4_u3_buf0_reg[4]/P0001 ,
		_w3761_,
		_w3773_,
		_w8555_
	);
	LUT3 #(
		.INIT('h80)
	) name6806 (
		\u4_buf0_reg[4]/P0001 ,
		_w3761_,
		_w3775_,
		_w8556_
	);
	LUT4 #(
		.INIT('hfffb)
	) name6807 (
		_w8552_,
		_w8554_,
		_w8555_,
		_w8556_,
		_w8557_
	);
	LUT3 #(
		.INIT('h80)
	) name6808 (
		\u4_u2_buf0_reg[5]/P0001 ,
		_w3762_,
		_w3763_,
		_w8558_
	);
	LUT2 #(
		.INIT('h8)
	) name6809 (
		_w3761_,
		_w8558_,
		_w8559_
	);
	LUT3 #(
		.INIT('h80)
	) name6810 (
		\u4_u0_buf0_reg[5]/P0001 ,
		_w3755_,
		_w3756_,
		_w8560_
	);
	LUT3 #(
		.INIT('h07)
	) name6811 (
		\u4_u1_buf0_reg[5]/P0001 ,
		_w3768_,
		_w8560_,
		_w8561_
	);
	LUT3 #(
		.INIT('h80)
	) name6812 (
		\u4_u3_buf0_reg[5]/P0001 ,
		_w3761_,
		_w3773_,
		_w8562_
	);
	LUT3 #(
		.INIT('h80)
	) name6813 (
		\u4_buf0_reg[5]/P0001 ,
		_w3761_,
		_w3775_,
		_w8563_
	);
	LUT4 #(
		.INIT('hfffb)
	) name6814 (
		_w8559_,
		_w8561_,
		_w8562_,
		_w8563_,
		_w8564_
	);
	LUT3 #(
		.INIT('h80)
	) name6815 (
		\u4_u2_buf0_reg[6]/P0001 ,
		_w3762_,
		_w3763_,
		_w8565_
	);
	LUT2 #(
		.INIT('h8)
	) name6816 (
		_w3761_,
		_w8565_,
		_w8566_
	);
	LUT3 #(
		.INIT('h80)
	) name6817 (
		\u4_u0_buf0_reg[6]/P0001 ,
		_w3755_,
		_w3756_,
		_w8567_
	);
	LUT3 #(
		.INIT('h07)
	) name6818 (
		\u4_u1_buf0_reg[6]/P0001 ,
		_w3768_,
		_w8567_,
		_w8568_
	);
	LUT3 #(
		.INIT('h80)
	) name6819 (
		\u4_u3_buf0_reg[6]/P0001 ,
		_w3761_,
		_w3773_,
		_w8569_
	);
	LUT3 #(
		.INIT('h80)
	) name6820 (
		\u4_buf0_reg[6]/P0001 ,
		_w3761_,
		_w3775_,
		_w8570_
	);
	LUT4 #(
		.INIT('hfffb)
	) name6821 (
		_w8566_,
		_w8568_,
		_w8569_,
		_w8570_,
		_w8571_
	);
	LUT3 #(
		.INIT('h80)
	) name6822 (
		\u4_u2_buf0_reg[7]/P0001 ,
		_w3762_,
		_w3763_,
		_w8572_
	);
	LUT2 #(
		.INIT('h8)
	) name6823 (
		_w3761_,
		_w8572_,
		_w8573_
	);
	LUT3 #(
		.INIT('h80)
	) name6824 (
		\u4_u0_buf0_reg[7]/P0001 ,
		_w3755_,
		_w3756_,
		_w8574_
	);
	LUT3 #(
		.INIT('h07)
	) name6825 (
		\u4_u1_buf0_reg[7]/P0001 ,
		_w3768_,
		_w8574_,
		_w8575_
	);
	LUT3 #(
		.INIT('h80)
	) name6826 (
		\u4_u3_buf0_reg[7]/P0001 ,
		_w3761_,
		_w3773_,
		_w8576_
	);
	LUT3 #(
		.INIT('h80)
	) name6827 (
		\u4_buf0_reg[7]/P0001 ,
		_w3761_,
		_w3775_,
		_w8577_
	);
	LUT4 #(
		.INIT('hfffb)
	) name6828 (
		_w8573_,
		_w8575_,
		_w8576_,
		_w8577_,
		_w8578_
	);
	LUT3 #(
		.INIT('h80)
	) name6829 (
		\u4_u2_buf0_reg[8]/P0001 ,
		_w3762_,
		_w3763_,
		_w8579_
	);
	LUT2 #(
		.INIT('h8)
	) name6830 (
		_w3761_,
		_w8579_,
		_w8580_
	);
	LUT3 #(
		.INIT('h80)
	) name6831 (
		\u4_u0_buf0_reg[8]/P0001 ,
		_w3755_,
		_w3756_,
		_w8581_
	);
	LUT3 #(
		.INIT('h07)
	) name6832 (
		\u4_u1_buf0_reg[8]/P0001 ,
		_w3768_,
		_w8581_,
		_w8582_
	);
	LUT3 #(
		.INIT('h80)
	) name6833 (
		\u4_u3_buf0_reg[8]/P0001 ,
		_w3761_,
		_w3773_,
		_w8583_
	);
	LUT3 #(
		.INIT('h80)
	) name6834 (
		\u4_buf0_reg[8]/P0001 ,
		_w3761_,
		_w3775_,
		_w8584_
	);
	LUT4 #(
		.INIT('hfffb)
	) name6835 (
		_w8580_,
		_w8582_,
		_w8583_,
		_w8584_,
		_w8585_
	);
	LUT3 #(
		.INIT('h80)
	) name6836 (
		\u4_u2_buf0_reg[9]/P0001 ,
		_w3762_,
		_w3763_,
		_w8586_
	);
	LUT2 #(
		.INIT('h8)
	) name6837 (
		_w3761_,
		_w8586_,
		_w8587_
	);
	LUT3 #(
		.INIT('h80)
	) name6838 (
		\u4_u0_buf0_reg[9]/P0001 ,
		_w3755_,
		_w3756_,
		_w8588_
	);
	LUT3 #(
		.INIT('h07)
	) name6839 (
		\u4_u1_buf0_reg[9]/P0001 ,
		_w3768_,
		_w8588_,
		_w8589_
	);
	LUT3 #(
		.INIT('h80)
	) name6840 (
		\u4_u3_buf0_reg[9]/P0001 ,
		_w3761_,
		_w3773_,
		_w8590_
	);
	LUT3 #(
		.INIT('h80)
	) name6841 (
		\u4_buf0_reg[9]/P0001 ,
		_w3761_,
		_w3775_,
		_w8591_
	);
	LUT4 #(
		.INIT('hfffb)
	) name6842 (
		_w8587_,
		_w8589_,
		_w8590_,
		_w8591_,
		_w8592_
	);
	LUT3 #(
		.INIT('h80)
	) name6843 (
		\u4_u2_buf1_reg[0]/P0001 ,
		_w3762_,
		_w3763_,
		_w8593_
	);
	LUT2 #(
		.INIT('h8)
	) name6844 (
		_w3761_,
		_w8593_,
		_w8594_
	);
	LUT3 #(
		.INIT('h80)
	) name6845 (
		\u4_u0_buf1_reg[0]/P0001 ,
		_w3755_,
		_w3756_,
		_w8595_
	);
	LUT3 #(
		.INIT('h07)
	) name6846 (
		\u4_u1_buf1_reg[0]/P0001 ,
		_w3768_,
		_w8595_,
		_w8596_
	);
	LUT3 #(
		.INIT('h80)
	) name6847 (
		\u4_u3_buf1_reg[0]/P0001 ,
		_w3761_,
		_w3773_,
		_w8597_
	);
	LUT3 #(
		.INIT('h80)
	) name6848 (
		\u4_buf1_reg[0]/P0001 ,
		_w3761_,
		_w3775_,
		_w8598_
	);
	LUT4 #(
		.INIT('hfffb)
	) name6849 (
		_w8594_,
		_w8596_,
		_w8597_,
		_w8598_,
		_w8599_
	);
	LUT3 #(
		.INIT('h80)
	) name6850 (
		\u4_u2_buf1_reg[10]/P0001 ,
		_w3762_,
		_w3763_,
		_w8600_
	);
	LUT2 #(
		.INIT('h8)
	) name6851 (
		_w3761_,
		_w8600_,
		_w8601_
	);
	LUT3 #(
		.INIT('h80)
	) name6852 (
		\u4_u0_buf1_reg[10]/P0001 ,
		_w3755_,
		_w3756_,
		_w8602_
	);
	LUT3 #(
		.INIT('h07)
	) name6853 (
		\u4_u1_buf1_reg[10]/P0001 ,
		_w3768_,
		_w8602_,
		_w8603_
	);
	LUT3 #(
		.INIT('h80)
	) name6854 (
		\u4_u3_buf1_reg[10]/P0001 ,
		_w3761_,
		_w3773_,
		_w8604_
	);
	LUT3 #(
		.INIT('h80)
	) name6855 (
		\u4_buf1_reg[10]/P0001 ,
		_w3761_,
		_w3775_,
		_w8605_
	);
	LUT4 #(
		.INIT('hfffb)
	) name6856 (
		_w8601_,
		_w8603_,
		_w8604_,
		_w8605_,
		_w8606_
	);
	LUT3 #(
		.INIT('h80)
	) name6857 (
		\u4_u2_buf1_reg[11]/P0001 ,
		_w3762_,
		_w3763_,
		_w8607_
	);
	LUT2 #(
		.INIT('h8)
	) name6858 (
		_w3761_,
		_w8607_,
		_w8608_
	);
	LUT3 #(
		.INIT('h80)
	) name6859 (
		\u4_u0_buf1_reg[11]/P0001 ,
		_w3755_,
		_w3756_,
		_w8609_
	);
	LUT3 #(
		.INIT('h07)
	) name6860 (
		\u4_u1_buf1_reg[11]/P0001 ,
		_w3768_,
		_w8609_,
		_w8610_
	);
	LUT3 #(
		.INIT('h80)
	) name6861 (
		\u4_u3_buf1_reg[11]/P0001 ,
		_w3761_,
		_w3773_,
		_w8611_
	);
	LUT3 #(
		.INIT('h80)
	) name6862 (
		\u4_buf1_reg[11]/P0001 ,
		_w3761_,
		_w3775_,
		_w8612_
	);
	LUT4 #(
		.INIT('hfffb)
	) name6863 (
		_w8608_,
		_w8610_,
		_w8611_,
		_w8612_,
		_w8613_
	);
	LUT3 #(
		.INIT('h80)
	) name6864 (
		\u4_u2_buf1_reg[12]/P0001 ,
		_w3762_,
		_w3763_,
		_w8614_
	);
	LUT2 #(
		.INIT('h8)
	) name6865 (
		_w3761_,
		_w8614_,
		_w8615_
	);
	LUT3 #(
		.INIT('h80)
	) name6866 (
		\u4_u0_buf1_reg[12]/P0001 ,
		_w3755_,
		_w3756_,
		_w8616_
	);
	LUT3 #(
		.INIT('h07)
	) name6867 (
		\u4_u1_buf1_reg[12]/P0001 ,
		_w3768_,
		_w8616_,
		_w8617_
	);
	LUT3 #(
		.INIT('h80)
	) name6868 (
		\u4_u3_buf1_reg[12]/P0001 ,
		_w3761_,
		_w3773_,
		_w8618_
	);
	LUT3 #(
		.INIT('h80)
	) name6869 (
		\u4_buf1_reg[12]/P0001 ,
		_w3761_,
		_w3775_,
		_w8619_
	);
	LUT4 #(
		.INIT('hfffb)
	) name6870 (
		_w8615_,
		_w8617_,
		_w8618_,
		_w8619_,
		_w8620_
	);
	LUT3 #(
		.INIT('h80)
	) name6871 (
		\u4_u2_buf1_reg[13]/P0001 ,
		_w3762_,
		_w3763_,
		_w8621_
	);
	LUT2 #(
		.INIT('h8)
	) name6872 (
		_w3761_,
		_w8621_,
		_w8622_
	);
	LUT3 #(
		.INIT('h80)
	) name6873 (
		\u4_u0_buf1_reg[13]/P0001 ,
		_w3755_,
		_w3756_,
		_w8623_
	);
	LUT3 #(
		.INIT('h07)
	) name6874 (
		\u4_u1_buf1_reg[13]/P0001 ,
		_w3768_,
		_w8623_,
		_w8624_
	);
	LUT3 #(
		.INIT('h80)
	) name6875 (
		\u4_u3_buf1_reg[13]/P0001 ,
		_w3761_,
		_w3773_,
		_w8625_
	);
	LUT3 #(
		.INIT('h80)
	) name6876 (
		\u4_buf1_reg[13]/P0001 ,
		_w3761_,
		_w3775_,
		_w8626_
	);
	LUT4 #(
		.INIT('hfffb)
	) name6877 (
		_w8622_,
		_w8624_,
		_w8625_,
		_w8626_,
		_w8627_
	);
	LUT3 #(
		.INIT('h80)
	) name6878 (
		\u4_u2_buf1_reg[14]/P0001 ,
		_w3762_,
		_w3763_,
		_w8628_
	);
	LUT2 #(
		.INIT('h8)
	) name6879 (
		_w3761_,
		_w8628_,
		_w8629_
	);
	LUT3 #(
		.INIT('h80)
	) name6880 (
		\u4_u0_buf1_reg[14]/P0001 ,
		_w3755_,
		_w3756_,
		_w8630_
	);
	LUT3 #(
		.INIT('h07)
	) name6881 (
		\u4_u1_buf1_reg[14]/P0001 ,
		_w3768_,
		_w8630_,
		_w8631_
	);
	LUT3 #(
		.INIT('h80)
	) name6882 (
		\u4_u3_buf1_reg[14]/P0001 ,
		_w3761_,
		_w3773_,
		_w8632_
	);
	LUT3 #(
		.INIT('h80)
	) name6883 (
		\u4_buf1_reg[14]/P0001 ,
		_w3761_,
		_w3775_,
		_w8633_
	);
	LUT4 #(
		.INIT('hfffb)
	) name6884 (
		_w8629_,
		_w8631_,
		_w8632_,
		_w8633_,
		_w8634_
	);
	LUT3 #(
		.INIT('h80)
	) name6885 (
		\u4_u2_buf1_reg[15]/P0001 ,
		_w3762_,
		_w3763_,
		_w8635_
	);
	LUT2 #(
		.INIT('h8)
	) name6886 (
		_w3761_,
		_w8635_,
		_w8636_
	);
	LUT3 #(
		.INIT('h80)
	) name6887 (
		\u4_u0_buf1_reg[15]/P0001 ,
		_w3755_,
		_w3756_,
		_w8637_
	);
	LUT3 #(
		.INIT('h07)
	) name6888 (
		\u4_u1_buf1_reg[15]/P0001 ,
		_w3768_,
		_w8637_,
		_w8638_
	);
	LUT3 #(
		.INIT('h80)
	) name6889 (
		\u4_u3_buf1_reg[15]/P0001 ,
		_w3761_,
		_w3773_,
		_w8639_
	);
	LUT3 #(
		.INIT('h80)
	) name6890 (
		\u4_buf1_reg[15]/P0001 ,
		_w3761_,
		_w3775_,
		_w8640_
	);
	LUT4 #(
		.INIT('hfffb)
	) name6891 (
		_w8636_,
		_w8638_,
		_w8639_,
		_w8640_,
		_w8641_
	);
	LUT3 #(
		.INIT('h80)
	) name6892 (
		\u4_u2_buf1_reg[16]/P0001 ,
		_w3762_,
		_w3763_,
		_w8642_
	);
	LUT2 #(
		.INIT('h8)
	) name6893 (
		_w3761_,
		_w8642_,
		_w8643_
	);
	LUT3 #(
		.INIT('h80)
	) name6894 (
		\u4_u0_buf1_reg[16]/P0001 ,
		_w3755_,
		_w3756_,
		_w8644_
	);
	LUT3 #(
		.INIT('h07)
	) name6895 (
		\u4_u1_buf1_reg[16]/P0001 ,
		_w3768_,
		_w8644_,
		_w8645_
	);
	LUT3 #(
		.INIT('h80)
	) name6896 (
		\u4_u3_buf1_reg[16]/P0001 ,
		_w3761_,
		_w3773_,
		_w8646_
	);
	LUT3 #(
		.INIT('h80)
	) name6897 (
		\u4_buf1_reg[16]/P0001 ,
		_w3761_,
		_w3775_,
		_w8647_
	);
	LUT4 #(
		.INIT('hfffb)
	) name6898 (
		_w8643_,
		_w8645_,
		_w8646_,
		_w8647_,
		_w8648_
	);
	LUT3 #(
		.INIT('h80)
	) name6899 (
		\u4_u2_buf1_reg[17]/P0001 ,
		_w3762_,
		_w3763_,
		_w8649_
	);
	LUT2 #(
		.INIT('h8)
	) name6900 (
		_w3761_,
		_w8649_,
		_w8650_
	);
	LUT3 #(
		.INIT('h80)
	) name6901 (
		\u4_u0_buf1_reg[17]/P0001 ,
		_w3755_,
		_w3756_,
		_w8651_
	);
	LUT3 #(
		.INIT('h07)
	) name6902 (
		\u4_u1_buf1_reg[17]/P0001 ,
		_w3768_,
		_w8651_,
		_w8652_
	);
	LUT3 #(
		.INIT('h80)
	) name6903 (
		\u4_u3_buf1_reg[17]/P0001 ,
		_w3761_,
		_w3773_,
		_w8653_
	);
	LUT3 #(
		.INIT('h80)
	) name6904 (
		\u4_buf1_reg[17]/NET0131 ,
		_w3761_,
		_w3775_,
		_w8654_
	);
	LUT4 #(
		.INIT('hfffb)
	) name6905 (
		_w8650_,
		_w8652_,
		_w8653_,
		_w8654_,
		_w8655_
	);
	LUT3 #(
		.INIT('h80)
	) name6906 (
		\u4_u2_buf1_reg[18]/P0001 ,
		_w3762_,
		_w3763_,
		_w8656_
	);
	LUT2 #(
		.INIT('h8)
	) name6907 (
		_w3761_,
		_w8656_,
		_w8657_
	);
	LUT3 #(
		.INIT('h80)
	) name6908 (
		\u4_u0_buf1_reg[18]/P0001 ,
		_w3755_,
		_w3756_,
		_w8658_
	);
	LUT3 #(
		.INIT('h07)
	) name6909 (
		\u4_u1_buf1_reg[18]/P0001 ,
		_w3768_,
		_w8658_,
		_w8659_
	);
	LUT3 #(
		.INIT('h80)
	) name6910 (
		\u4_u3_buf1_reg[18]/P0001 ,
		_w3761_,
		_w3773_,
		_w8660_
	);
	LUT3 #(
		.INIT('h80)
	) name6911 (
		\u4_buf1_reg[18]/P0001 ,
		_w3761_,
		_w3775_,
		_w8661_
	);
	LUT4 #(
		.INIT('hfffb)
	) name6912 (
		_w8657_,
		_w8659_,
		_w8660_,
		_w8661_,
		_w8662_
	);
	LUT3 #(
		.INIT('h80)
	) name6913 (
		\u4_u2_buf1_reg[19]/P0001 ,
		_w3762_,
		_w3763_,
		_w8663_
	);
	LUT2 #(
		.INIT('h8)
	) name6914 (
		_w3761_,
		_w8663_,
		_w8664_
	);
	LUT3 #(
		.INIT('h80)
	) name6915 (
		\u4_u0_buf1_reg[19]/P0001 ,
		_w3755_,
		_w3756_,
		_w8665_
	);
	LUT3 #(
		.INIT('h07)
	) name6916 (
		\u4_u1_buf1_reg[19]/P0001 ,
		_w3768_,
		_w8665_,
		_w8666_
	);
	LUT3 #(
		.INIT('h80)
	) name6917 (
		\u4_u3_buf1_reg[19]/P0001 ,
		_w3761_,
		_w3773_,
		_w8667_
	);
	LUT3 #(
		.INIT('h80)
	) name6918 (
		\u4_buf1_reg[19]/NET0131 ,
		_w3761_,
		_w3775_,
		_w8668_
	);
	LUT4 #(
		.INIT('hfffb)
	) name6919 (
		_w8664_,
		_w8666_,
		_w8667_,
		_w8668_,
		_w8669_
	);
	LUT3 #(
		.INIT('h80)
	) name6920 (
		\u4_u2_buf1_reg[1]/P0001 ,
		_w3762_,
		_w3763_,
		_w8670_
	);
	LUT2 #(
		.INIT('h8)
	) name6921 (
		_w3761_,
		_w8670_,
		_w8671_
	);
	LUT3 #(
		.INIT('h80)
	) name6922 (
		\u4_u0_buf1_reg[1]/P0001 ,
		_w3755_,
		_w3756_,
		_w8672_
	);
	LUT3 #(
		.INIT('h07)
	) name6923 (
		\u4_u1_buf1_reg[1]/P0001 ,
		_w3768_,
		_w8672_,
		_w8673_
	);
	LUT3 #(
		.INIT('h80)
	) name6924 (
		\u4_u3_buf1_reg[1]/P0001 ,
		_w3761_,
		_w3773_,
		_w8674_
	);
	LUT3 #(
		.INIT('h80)
	) name6925 (
		\u4_buf1_reg[1]/P0001 ,
		_w3761_,
		_w3775_,
		_w8675_
	);
	LUT4 #(
		.INIT('hfffb)
	) name6926 (
		_w8671_,
		_w8673_,
		_w8674_,
		_w8675_,
		_w8676_
	);
	LUT3 #(
		.INIT('h80)
	) name6927 (
		\u4_u2_buf1_reg[20]/P0001 ,
		_w3762_,
		_w3763_,
		_w8677_
	);
	LUT2 #(
		.INIT('h8)
	) name6928 (
		_w3761_,
		_w8677_,
		_w8678_
	);
	LUT3 #(
		.INIT('h80)
	) name6929 (
		\u4_u0_buf1_reg[20]/P0001 ,
		_w3755_,
		_w3756_,
		_w8679_
	);
	LUT3 #(
		.INIT('h07)
	) name6930 (
		\u4_u1_buf1_reg[20]/P0001 ,
		_w3768_,
		_w8679_,
		_w8680_
	);
	LUT3 #(
		.INIT('h80)
	) name6931 (
		\u4_u3_buf1_reg[20]/P0001 ,
		_w3761_,
		_w3773_,
		_w8681_
	);
	LUT3 #(
		.INIT('h80)
	) name6932 (
		\u4_buf1_reg[20]/NET0131 ,
		_w3761_,
		_w3775_,
		_w8682_
	);
	LUT4 #(
		.INIT('hfffb)
	) name6933 (
		_w8678_,
		_w8680_,
		_w8681_,
		_w8682_,
		_w8683_
	);
	LUT3 #(
		.INIT('h80)
	) name6934 (
		\u4_u2_buf1_reg[21]/P0001 ,
		_w3762_,
		_w3763_,
		_w8684_
	);
	LUT2 #(
		.INIT('h8)
	) name6935 (
		_w3761_,
		_w8684_,
		_w8685_
	);
	LUT3 #(
		.INIT('h80)
	) name6936 (
		\u4_u0_buf1_reg[21]/P0001 ,
		_w3755_,
		_w3756_,
		_w8686_
	);
	LUT3 #(
		.INIT('h07)
	) name6937 (
		\u4_u1_buf1_reg[21]/P0001 ,
		_w3768_,
		_w8686_,
		_w8687_
	);
	LUT3 #(
		.INIT('h80)
	) name6938 (
		\u4_u3_buf1_reg[21]/P0001 ,
		_w3761_,
		_w3773_,
		_w8688_
	);
	LUT3 #(
		.INIT('h80)
	) name6939 (
		\u4_buf1_reg[21]/NET0131 ,
		_w3761_,
		_w3775_,
		_w8689_
	);
	LUT4 #(
		.INIT('hfffb)
	) name6940 (
		_w8685_,
		_w8687_,
		_w8688_,
		_w8689_,
		_w8690_
	);
	LUT3 #(
		.INIT('h80)
	) name6941 (
		\u4_u2_buf1_reg[22]/P0001 ,
		_w3762_,
		_w3763_,
		_w8691_
	);
	LUT2 #(
		.INIT('h8)
	) name6942 (
		_w3761_,
		_w8691_,
		_w8692_
	);
	LUT3 #(
		.INIT('h80)
	) name6943 (
		\u4_u0_buf1_reg[22]/P0001 ,
		_w3755_,
		_w3756_,
		_w8693_
	);
	LUT3 #(
		.INIT('h07)
	) name6944 (
		\u4_u1_buf1_reg[22]/P0001 ,
		_w3768_,
		_w8693_,
		_w8694_
	);
	LUT3 #(
		.INIT('h80)
	) name6945 (
		\u4_u3_buf1_reg[22]/P0001 ,
		_w3761_,
		_w3773_,
		_w8695_
	);
	LUT3 #(
		.INIT('h80)
	) name6946 (
		\u4_buf1_reg[22]/NET0131 ,
		_w3761_,
		_w3775_,
		_w8696_
	);
	LUT4 #(
		.INIT('hfffb)
	) name6947 (
		_w8692_,
		_w8694_,
		_w8695_,
		_w8696_,
		_w8697_
	);
	LUT3 #(
		.INIT('h80)
	) name6948 (
		\u4_u2_buf1_reg[23]/P0001 ,
		_w3762_,
		_w3763_,
		_w8698_
	);
	LUT2 #(
		.INIT('h8)
	) name6949 (
		_w3761_,
		_w8698_,
		_w8699_
	);
	LUT3 #(
		.INIT('h80)
	) name6950 (
		\u4_u0_buf1_reg[23]/P0001 ,
		_w3755_,
		_w3756_,
		_w8700_
	);
	LUT3 #(
		.INIT('h07)
	) name6951 (
		\u4_u1_buf1_reg[23]/P0001 ,
		_w3768_,
		_w8700_,
		_w8701_
	);
	LUT3 #(
		.INIT('h80)
	) name6952 (
		\u4_u3_buf1_reg[23]/P0001 ,
		_w3761_,
		_w3773_,
		_w8702_
	);
	LUT3 #(
		.INIT('h80)
	) name6953 (
		\u4_buf1_reg[23]/NET0131 ,
		_w3761_,
		_w3775_,
		_w8703_
	);
	LUT4 #(
		.INIT('hfffb)
	) name6954 (
		_w8699_,
		_w8701_,
		_w8702_,
		_w8703_,
		_w8704_
	);
	LUT3 #(
		.INIT('h80)
	) name6955 (
		\u4_u2_buf1_reg[25]/P0001 ,
		_w3762_,
		_w3763_,
		_w8705_
	);
	LUT2 #(
		.INIT('h8)
	) name6956 (
		_w3761_,
		_w8705_,
		_w8706_
	);
	LUT3 #(
		.INIT('h80)
	) name6957 (
		\u4_u0_buf1_reg[25]/P0001 ,
		_w3755_,
		_w3756_,
		_w8707_
	);
	LUT3 #(
		.INIT('h07)
	) name6958 (
		\u4_u1_buf1_reg[25]/P0001 ,
		_w3768_,
		_w8707_,
		_w8708_
	);
	LUT3 #(
		.INIT('h80)
	) name6959 (
		\u4_u3_buf1_reg[25]/P0001 ,
		_w3761_,
		_w3773_,
		_w8709_
	);
	LUT3 #(
		.INIT('h80)
	) name6960 (
		\u4_buf1_reg[25]/NET0131 ,
		_w3761_,
		_w3775_,
		_w8710_
	);
	LUT4 #(
		.INIT('hfffb)
	) name6961 (
		_w8706_,
		_w8708_,
		_w8709_,
		_w8710_,
		_w8711_
	);
	LUT3 #(
		.INIT('h80)
	) name6962 (
		\u4_u2_buf1_reg[3]/P0001 ,
		_w3762_,
		_w3763_,
		_w8712_
	);
	LUT2 #(
		.INIT('h8)
	) name6963 (
		_w3761_,
		_w8712_,
		_w8713_
	);
	LUT3 #(
		.INIT('h80)
	) name6964 (
		\u4_u0_buf1_reg[3]/P0001 ,
		_w3755_,
		_w3756_,
		_w8714_
	);
	LUT3 #(
		.INIT('h07)
	) name6965 (
		\u4_u1_buf1_reg[3]/P0001 ,
		_w3768_,
		_w8714_,
		_w8715_
	);
	LUT3 #(
		.INIT('h80)
	) name6966 (
		\u4_u3_buf1_reg[3]/P0001 ,
		_w3761_,
		_w3773_,
		_w8716_
	);
	LUT3 #(
		.INIT('h80)
	) name6967 (
		\u4_buf1_reg[3]/P0001 ,
		_w3761_,
		_w3775_,
		_w8717_
	);
	LUT4 #(
		.INIT('hfffb)
	) name6968 (
		_w8713_,
		_w8715_,
		_w8716_,
		_w8717_,
		_w8718_
	);
	LUT3 #(
		.INIT('h80)
	) name6969 (
		\u4_u2_buf1_reg[26]/P0001 ,
		_w3762_,
		_w3763_,
		_w8719_
	);
	LUT2 #(
		.INIT('h8)
	) name6970 (
		_w3761_,
		_w8719_,
		_w8720_
	);
	LUT3 #(
		.INIT('h80)
	) name6971 (
		\u4_u0_buf1_reg[26]/P0001 ,
		_w3755_,
		_w3756_,
		_w8721_
	);
	LUT3 #(
		.INIT('h07)
	) name6972 (
		\u4_u1_buf1_reg[26]/P0001 ,
		_w3768_,
		_w8721_,
		_w8722_
	);
	LUT3 #(
		.INIT('h80)
	) name6973 (
		\u4_u3_buf1_reg[26]/P0001 ,
		_w3761_,
		_w3773_,
		_w8723_
	);
	LUT3 #(
		.INIT('h80)
	) name6974 (
		\u4_buf1_reg[26]/NET0131 ,
		_w3761_,
		_w3775_,
		_w8724_
	);
	LUT4 #(
		.INIT('hfffb)
	) name6975 (
		_w8720_,
		_w8722_,
		_w8723_,
		_w8724_,
		_w8725_
	);
	LUT3 #(
		.INIT('h80)
	) name6976 (
		\u4_u2_buf1_reg[27]/P0001 ,
		_w3762_,
		_w3763_,
		_w8726_
	);
	LUT2 #(
		.INIT('h8)
	) name6977 (
		_w3761_,
		_w8726_,
		_w8727_
	);
	LUT3 #(
		.INIT('h80)
	) name6978 (
		\u4_u0_buf1_reg[27]/P0001 ,
		_w3755_,
		_w3756_,
		_w8728_
	);
	LUT3 #(
		.INIT('h07)
	) name6979 (
		\u4_u1_buf1_reg[27]/P0001 ,
		_w3768_,
		_w8728_,
		_w8729_
	);
	LUT3 #(
		.INIT('h80)
	) name6980 (
		\u4_u3_buf1_reg[27]/P0001 ,
		_w3761_,
		_w3773_,
		_w8730_
	);
	LUT3 #(
		.INIT('h80)
	) name6981 (
		\u4_buf1_reg[27]/P0001 ,
		_w3761_,
		_w3775_,
		_w8731_
	);
	LUT4 #(
		.INIT('hfffb)
	) name6982 (
		_w8727_,
		_w8729_,
		_w8730_,
		_w8731_,
		_w8732_
	);
	LUT3 #(
		.INIT('h80)
	) name6983 (
		\u4_u2_buf1_reg[28]/P0001 ,
		_w3762_,
		_w3763_,
		_w8733_
	);
	LUT2 #(
		.INIT('h8)
	) name6984 (
		_w3761_,
		_w8733_,
		_w8734_
	);
	LUT3 #(
		.INIT('h80)
	) name6985 (
		\u4_u0_buf1_reg[28]/P0001 ,
		_w3755_,
		_w3756_,
		_w8735_
	);
	LUT3 #(
		.INIT('h07)
	) name6986 (
		\u4_u1_buf1_reg[28]/P0001 ,
		_w3768_,
		_w8735_,
		_w8736_
	);
	LUT3 #(
		.INIT('h80)
	) name6987 (
		\u4_u3_buf1_reg[28]/P0001 ,
		_w3761_,
		_w3773_,
		_w8737_
	);
	LUT3 #(
		.INIT('h80)
	) name6988 (
		\u4_buf1_reg[28]/P0001 ,
		_w3761_,
		_w3775_,
		_w8738_
	);
	LUT4 #(
		.INIT('hfffb)
	) name6989 (
		_w8734_,
		_w8736_,
		_w8737_,
		_w8738_,
		_w8739_
	);
	LUT3 #(
		.INIT('h80)
	) name6990 (
		\u4_u2_buf1_reg[29]/P0001 ,
		_w3762_,
		_w3763_,
		_w8740_
	);
	LUT2 #(
		.INIT('h8)
	) name6991 (
		_w3761_,
		_w8740_,
		_w8741_
	);
	LUT3 #(
		.INIT('h80)
	) name6992 (
		\u4_u0_buf1_reg[29]/P0001 ,
		_w3755_,
		_w3756_,
		_w8742_
	);
	LUT3 #(
		.INIT('h07)
	) name6993 (
		\u4_u1_buf1_reg[29]/P0001 ,
		_w3768_,
		_w8742_,
		_w8743_
	);
	LUT3 #(
		.INIT('h80)
	) name6994 (
		\u4_u3_buf1_reg[29]/P0001 ,
		_w3761_,
		_w3773_,
		_w8744_
	);
	LUT3 #(
		.INIT('h80)
	) name6995 (
		\u4_buf1_reg[29]/P0001 ,
		_w3761_,
		_w3775_,
		_w8745_
	);
	LUT4 #(
		.INIT('hfffb)
	) name6996 (
		_w8741_,
		_w8743_,
		_w8744_,
		_w8745_,
		_w8746_
	);
	LUT3 #(
		.INIT('h80)
	) name6997 (
		\u4_u2_buf1_reg[2]/P0001 ,
		_w3762_,
		_w3763_,
		_w8747_
	);
	LUT2 #(
		.INIT('h8)
	) name6998 (
		_w3761_,
		_w8747_,
		_w8748_
	);
	LUT3 #(
		.INIT('h80)
	) name6999 (
		\u4_u0_buf1_reg[2]/P0001 ,
		_w3755_,
		_w3756_,
		_w8749_
	);
	LUT3 #(
		.INIT('h07)
	) name7000 (
		\u4_u1_buf1_reg[2]/P0001 ,
		_w3768_,
		_w8749_,
		_w8750_
	);
	LUT3 #(
		.INIT('h80)
	) name7001 (
		\u4_u3_buf1_reg[2]/P0001 ,
		_w3761_,
		_w3773_,
		_w8751_
	);
	LUT3 #(
		.INIT('h80)
	) name7002 (
		\u4_buf1_reg[2]/P0001 ,
		_w3761_,
		_w3775_,
		_w8752_
	);
	LUT4 #(
		.INIT('hfffb)
	) name7003 (
		_w8748_,
		_w8750_,
		_w8751_,
		_w8752_,
		_w8753_
	);
	LUT3 #(
		.INIT('h80)
	) name7004 (
		\u4_u2_buf1_reg[30]/P0001 ,
		_w3762_,
		_w3763_,
		_w8754_
	);
	LUT2 #(
		.INIT('h8)
	) name7005 (
		_w3761_,
		_w8754_,
		_w8755_
	);
	LUT3 #(
		.INIT('h80)
	) name7006 (
		\u4_u0_buf1_reg[30]/P0001 ,
		_w3755_,
		_w3756_,
		_w8756_
	);
	LUT3 #(
		.INIT('h07)
	) name7007 (
		\u4_u1_buf1_reg[30]/P0001 ,
		_w3768_,
		_w8756_,
		_w8757_
	);
	LUT3 #(
		.INIT('h80)
	) name7008 (
		\u4_u3_buf1_reg[30]/P0001 ,
		_w3761_,
		_w3773_,
		_w8758_
	);
	LUT3 #(
		.INIT('h80)
	) name7009 (
		\u4_buf1_reg[30]/P0001 ,
		_w3761_,
		_w3775_,
		_w8759_
	);
	LUT4 #(
		.INIT('hfffb)
	) name7010 (
		_w8755_,
		_w8757_,
		_w8758_,
		_w8759_,
		_w8760_
	);
	LUT3 #(
		.INIT('h80)
	) name7011 (
		\u4_u2_buf1_reg[31]/P0001 ,
		_w3762_,
		_w3763_,
		_w8761_
	);
	LUT2 #(
		.INIT('h8)
	) name7012 (
		_w3761_,
		_w8761_,
		_w8762_
	);
	LUT3 #(
		.INIT('h80)
	) name7013 (
		\u4_u0_buf1_reg[31]/P0001 ,
		_w3755_,
		_w3756_,
		_w8763_
	);
	LUT3 #(
		.INIT('h07)
	) name7014 (
		\u4_u1_buf1_reg[31]/P0001 ,
		_w3768_,
		_w8763_,
		_w8764_
	);
	LUT3 #(
		.INIT('h80)
	) name7015 (
		\u4_u3_buf1_reg[31]/P0001 ,
		_w3761_,
		_w3773_,
		_w8765_
	);
	LUT3 #(
		.INIT('h80)
	) name7016 (
		\u4_buf1_reg[31]/P0001 ,
		_w3761_,
		_w3775_,
		_w8766_
	);
	LUT4 #(
		.INIT('hfffb)
	) name7017 (
		_w8762_,
		_w8764_,
		_w8765_,
		_w8766_,
		_w8767_
	);
	LUT3 #(
		.INIT('h80)
	) name7018 (
		\u4_u2_buf1_reg[4]/P0001 ,
		_w3762_,
		_w3763_,
		_w8768_
	);
	LUT2 #(
		.INIT('h8)
	) name7019 (
		_w3761_,
		_w8768_,
		_w8769_
	);
	LUT3 #(
		.INIT('h80)
	) name7020 (
		\u4_u0_buf1_reg[4]/P0001 ,
		_w3755_,
		_w3756_,
		_w8770_
	);
	LUT3 #(
		.INIT('h07)
	) name7021 (
		\u4_u1_buf1_reg[4]/P0001 ,
		_w3768_,
		_w8770_,
		_w8771_
	);
	LUT3 #(
		.INIT('h80)
	) name7022 (
		\u4_u3_buf1_reg[4]/P0001 ,
		_w3761_,
		_w3773_,
		_w8772_
	);
	LUT3 #(
		.INIT('h80)
	) name7023 (
		\u4_buf1_reg[4]/P0001 ,
		_w3761_,
		_w3775_,
		_w8773_
	);
	LUT4 #(
		.INIT('hfffb)
	) name7024 (
		_w8769_,
		_w8771_,
		_w8772_,
		_w8773_,
		_w8774_
	);
	LUT3 #(
		.INIT('h80)
	) name7025 (
		\u4_u2_buf1_reg[7]/P0001 ,
		_w3762_,
		_w3763_,
		_w8775_
	);
	LUT2 #(
		.INIT('h8)
	) name7026 (
		_w3761_,
		_w8775_,
		_w8776_
	);
	LUT3 #(
		.INIT('h80)
	) name7027 (
		\u4_u0_buf1_reg[7]/P0001 ,
		_w3755_,
		_w3756_,
		_w8777_
	);
	LUT3 #(
		.INIT('h07)
	) name7028 (
		\u4_u1_buf1_reg[7]/P0001 ,
		_w3768_,
		_w8777_,
		_w8778_
	);
	LUT3 #(
		.INIT('h80)
	) name7029 (
		\u4_u3_buf1_reg[7]/P0001 ,
		_w3761_,
		_w3773_,
		_w8779_
	);
	LUT3 #(
		.INIT('h80)
	) name7030 (
		\u4_buf1_reg[7]/P0001 ,
		_w3761_,
		_w3775_,
		_w8780_
	);
	LUT4 #(
		.INIT('hfffb)
	) name7031 (
		_w8776_,
		_w8778_,
		_w8779_,
		_w8780_,
		_w8781_
	);
	LUT3 #(
		.INIT('h80)
	) name7032 (
		\u4_u2_buf1_reg[8]/P0001 ,
		_w3762_,
		_w3763_,
		_w8782_
	);
	LUT2 #(
		.INIT('h8)
	) name7033 (
		_w3761_,
		_w8782_,
		_w8783_
	);
	LUT3 #(
		.INIT('h80)
	) name7034 (
		\u4_u0_buf1_reg[8]/P0001 ,
		_w3755_,
		_w3756_,
		_w8784_
	);
	LUT3 #(
		.INIT('h07)
	) name7035 (
		\u4_u1_buf1_reg[8]/P0001 ,
		_w3768_,
		_w8784_,
		_w8785_
	);
	LUT3 #(
		.INIT('h80)
	) name7036 (
		\u4_u3_buf1_reg[8]/P0001 ,
		_w3761_,
		_w3773_,
		_w8786_
	);
	LUT3 #(
		.INIT('h80)
	) name7037 (
		\u4_buf1_reg[8]/P0001 ,
		_w3761_,
		_w3775_,
		_w8787_
	);
	LUT4 #(
		.INIT('hfffb)
	) name7038 (
		_w8783_,
		_w8785_,
		_w8786_,
		_w8787_,
		_w8788_
	);
	LUT3 #(
		.INIT('h80)
	) name7039 (
		\u4_u2_buf1_reg[9]/P0001 ,
		_w3762_,
		_w3763_,
		_w8789_
	);
	LUT2 #(
		.INIT('h8)
	) name7040 (
		_w3761_,
		_w8789_,
		_w8790_
	);
	LUT3 #(
		.INIT('h80)
	) name7041 (
		\u4_u0_buf1_reg[9]/P0001 ,
		_w3755_,
		_w3756_,
		_w8791_
	);
	LUT3 #(
		.INIT('h07)
	) name7042 (
		\u4_u1_buf1_reg[9]/P0001 ,
		_w3768_,
		_w8791_,
		_w8792_
	);
	LUT3 #(
		.INIT('h80)
	) name7043 (
		\u4_u3_buf1_reg[9]/P0001 ,
		_w3761_,
		_w3773_,
		_w8793_
	);
	LUT3 #(
		.INIT('h80)
	) name7044 (
		\u4_buf1_reg[9]/P0001 ,
		_w3761_,
		_w3775_,
		_w8794_
	);
	LUT4 #(
		.INIT('hfffb)
	) name7045 (
		_w8790_,
		_w8792_,
		_w8793_,
		_w8794_,
		_w8795_
	);
	LUT3 #(
		.INIT('h80)
	) name7046 (
		\u4_u2_csr0_reg[0]/P0001 ,
		_w3762_,
		_w3763_,
		_w8796_
	);
	LUT2 #(
		.INIT('h8)
	) name7047 (
		_w3761_,
		_w8796_,
		_w8797_
	);
	LUT3 #(
		.INIT('h80)
	) name7048 (
		\u4_u0_csr0_reg[0]/P0001 ,
		_w3755_,
		_w3756_,
		_w8798_
	);
	LUT3 #(
		.INIT('h07)
	) name7049 (
		\u4_u1_csr0_reg[0]/P0001 ,
		_w3768_,
		_w8798_,
		_w8799_
	);
	LUT3 #(
		.INIT('h80)
	) name7050 (
		\u4_u3_csr0_reg[0]/P0001 ,
		_w3761_,
		_w3773_,
		_w8800_
	);
	LUT3 #(
		.INIT('h80)
	) name7051 (
		\u4_csr_reg[0]/P0001 ,
		_w3761_,
		_w3775_,
		_w8801_
	);
	LUT4 #(
		.INIT('hfffb)
	) name7052 (
		_w8797_,
		_w8799_,
		_w8800_,
		_w8801_,
		_w8802_
	);
	LUT3 #(
		.INIT('h80)
	) name7053 (
		\u4_u2_csr0_reg[10]/P0001 ,
		_w3762_,
		_w3763_,
		_w8803_
	);
	LUT2 #(
		.INIT('h8)
	) name7054 (
		_w3761_,
		_w8803_,
		_w8804_
	);
	LUT3 #(
		.INIT('h80)
	) name7055 (
		\u4_u0_csr0_reg[10]/P0001 ,
		_w3755_,
		_w3756_,
		_w8805_
	);
	LUT3 #(
		.INIT('h07)
	) name7056 (
		\u4_u1_csr0_reg[10]/P0001 ,
		_w3768_,
		_w8805_,
		_w8806_
	);
	LUT3 #(
		.INIT('h80)
	) name7057 (
		\u4_u3_csr0_reg[10]/P0001 ,
		_w3761_,
		_w3773_,
		_w8807_
	);
	LUT3 #(
		.INIT('h80)
	) name7058 (
		\u4_csr_reg[10]/P0001 ,
		_w3761_,
		_w3775_,
		_w8808_
	);
	LUT4 #(
		.INIT('hfffb)
	) name7059 (
		_w8804_,
		_w8806_,
		_w8807_,
		_w8808_,
		_w8809_
	);
	LUT3 #(
		.INIT('h80)
	) name7060 (
		\u4_u2_csr0_reg[11]/P0001 ,
		_w3762_,
		_w3763_,
		_w8810_
	);
	LUT2 #(
		.INIT('h8)
	) name7061 (
		_w3761_,
		_w8810_,
		_w8811_
	);
	LUT3 #(
		.INIT('h80)
	) name7062 (
		\u4_u0_csr0_reg[11]/P0001 ,
		_w3755_,
		_w3756_,
		_w8812_
	);
	LUT3 #(
		.INIT('h07)
	) name7063 (
		\u4_u1_csr0_reg[11]/P0001 ,
		_w3768_,
		_w8812_,
		_w8813_
	);
	LUT3 #(
		.INIT('h80)
	) name7064 (
		\u4_u3_csr0_reg[11]/P0001 ,
		_w3761_,
		_w3773_,
		_w8814_
	);
	LUT3 #(
		.INIT('h80)
	) name7065 (
		\u4_csr_reg[11]/P0001 ,
		_w3761_,
		_w3775_,
		_w8815_
	);
	LUT4 #(
		.INIT('hfffb)
	) name7066 (
		_w8811_,
		_w8813_,
		_w8814_,
		_w8815_,
		_w8816_
	);
	LUT3 #(
		.INIT('h80)
	) name7067 (
		\u4_u2_csr0_reg[12]/P0001 ,
		_w3762_,
		_w3763_,
		_w8817_
	);
	LUT2 #(
		.INIT('h8)
	) name7068 (
		_w3761_,
		_w8817_,
		_w8818_
	);
	LUT3 #(
		.INIT('h80)
	) name7069 (
		\u4_u0_csr0_reg[12]/P0001 ,
		_w3755_,
		_w3756_,
		_w8819_
	);
	LUT3 #(
		.INIT('h07)
	) name7070 (
		\u4_u1_csr0_reg[12]/P0001 ,
		_w3768_,
		_w8819_,
		_w8820_
	);
	LUT3 #(
		.INIT('h80)
	) name7071 (
		\u4_u3_csr0_reg[12]/P0001 ,
		_w3761_,
		_w3773_,
		_w8821_
	);
	LUT3 #(
		.INIT('h80)
	) name7072 (
		\u4_csr_reg[12]/P0001 ,
		_w3761_,
		_w3775_,
		_w8822_
	);
	LUT4 #(
		.INIT('hfffb)
	) name7073 (
		_w8818_,
		_w8820_,
		_w8821_,
		_w8822_,
		_w8823_
	);
	LUT3 #(
		.INIT('h0e)
	) name7074 (
		\u1_u2_mack_r_reg/P0001 ,
		\u1_u2_state_reg[2]/NET0131 ,
		\u1_u3_abort_reg/P0001 ,
		_w8824_
	);
	LUT3 #(
		.INIT('h80)
	) name7075 (
		_w3209_,
		_w3225_,
		_w8824_,
		_w8825_
	);
	LUT3 #(
		.INIT('h04)
	) name7076 (
		\u1_u2_rx_data_done_r2_reg/P0001 ,
		\u1_u2_state_reg[2]/NET0131 ,
		\u1_u3_abort_reg/P0001 ,
		_w8826_
	);
	LUT3 #(
		.INIT('h80)
	) name7077 (
		_w3209_,
		_w7396_,
		_w8826_,
		_w8827_
	);
	LUT3 #(
		.INIT('ha8)
	) name7078 (
		rst_i_pad,
		_w8825_,
		_w8827_,
		_w8828_
	);
	LUT4 #(
		.INIT('h0007)
	) name7079 (
		\u0_u0_idle_cnt1_reg[4]/P0001 ,
		\u0_u0_idle_cnt1_reg[5]/P0001 ,
		\u0_u0_idle_cnt1_reg[6]/P0001 ,
		\u0_u0_idle_cnt1_reg[7]/P0001 ,
		_w8829_
	);
	LUT4 #(
		.INIT('ha2ff)
	) name7080 (
		_w5762_,
		_w5763_,
		_w5764_,
		_w8829_,
		_w8830_
	);
	LUT2 #(
		.INIT('h1)
	) name7081 (
		_w5769_,
		_w8830_,
		_w8831_
	);
	LUT4 #(
		.INIT('h5155)
	) name7082 (
		\u0_u0_chirp_cnt_reg[1]/P0001 ,
		_w4110_,
		_w8189_,
		_w8191_,
		_w8832_
	);
	LUT3 #(
		.INIT('h40)
	) name7083 (
		\u0_u0_chirp_cnt_is_6_reg/P0001 ,
		\u0_u0_chirp_cnt_reg[0]/P0001 ,
		\u0_u0_chirp_cnt_reg[1]/P0001 ,
		_w8833_
	);
	LUT4 #(
		.INIT('h5155)
	) name7084 (
		\u0_u0_state_reg[10]/P0001 ,
		_w4110_,
		_w8189_,
		_w8833_,
		_w8834_
	);
	LUT2 #(
		.INIT('h4)
	) name7085 (
		_w8832_,
		_w8834_,
		_w8835_
	);
	LUT2 #(
		.INIT('h2)
	) name7086 (
		\u0_u0_chirp_cnt_reg[2]/P0001 ,
		\u0_u0_state_reg[10]/P0001 ,
		_w8836_
	);
	LUT4 #(
		.INIT('hdf00)
	) name7087 (
		_w4110_,
		_w8189_,
		_w8833_,
		_w8836_,
		_w8837_
	);
	LUT2 #(
		.INIT('h1)
	) name7088 (
		\u0_u0_chirp_cnt_reg[2]/P0001 ,
		\u0_u0_state_reg[10]/P0001 ,
		_w8838_
	);
	LUT2 #(
		.INIT('h8)
	) name7089 (
		_w8833_,
		_w8838_,
		_w8839_
	);
	LUT3 #(
		.INIT('h20)
	) name7090 (
		_w4110_,
		_w8189_,
		_w8839_,
		_w8840_
	);
	LUT2 #(
		.INIT('he)
	) name7091 (
		_w8837_,
		_w8840_,
		_w8841_
	);
	LUT4 #(
		.INIT('h8000)
	) name7092 (
		_w2224_,
		_w2226_,
		_w2229_,
		_w5861_,
		_w8842_
	);
	LUT4 #(
		.INIT('h0002)
	) name7093 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		\wb_data_i[0]_pad ,
		_w8843_
	);
	LUT2 #(
		.INIT('h8)
	) name7094 (
		_w8842_,
		_w8843_,
		_w8844_
	);
	LUT2 #(
		.INIT('h8)
	) name7095 (
		rst_i_pad,
		\u4_funct_adr_reg[0]/P0001 ,
		_w8845_
	);
	LUT3 #(
		.INIT('h02)
	) name7096 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w8846_
	);
	LUT3 #(
		.INIT('h80)
	) name7097 (
		rst_i_pad,
		\u5_wb_req_s1_reg/P0001 ,
		wb_we_i_pad,
		_w8847_
	);
	LUT4 #(
		.INIT('h8000)
	) name7098 (
		_w2224_,
		_w2226_,
		_w5861_,
		_w8847_,
		_w8848_
	);
	LUT3 #(
		.INIT('h15)
	) name7099 (
		_w8845_,
		_w8846_,
		_w8848_,
		_w8849_
	);
	LUT2 #(
		.INIT('h1)
	) name7100 (
		_w8844_,
		_w8849_,
		_w8850_
	);
	LUT4 #(
		.INIT('h0002)
	) name7101 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		\wb_data_i[1]_pad ,
		_w8851_
	);
	LUT2 #(
		.INIT('h8)
	) name7102 (
		_w8842_,
		_w8851_,
		_w8852_
	);
	LUT2 #(
		.INIT('h8)
	) name7103 (
		rst_i_pad,
		\u4_funct_adr_reg[1]/P0001 ,
		_w8853_
	);
	LUT3 #(
		.INIT('h07)
	) name7104 (
		_w8846_,
		_w8848_,
		_w8853_,
		_w8854_
	);
	LUT2 #(
		.INIT('h1)
	) name7105 (
		_w8852_,
		_w8854_,
		_w8855_
	);
	LUT4 #(
		.INIT('h0002)
	) name7106 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		\wb_data_i[2]_pad ,
		_w8856_
	);
	LUT2 #(
		.INIT('h8)
	) name7107 (
		_w8842_,
		_w8856_,
		_w8857_
	);
	LUT2 #(
		.INIT('h8)
	) name7108 (
		rst_i_pad,
		\u4_funct_adr_reg[2]/P0001 ,
		_w8858_
	);
	LUT3 #(
		.INIT('h07)
	) name7109 (
		_w8846_,
		_w8848_,
		_w8858_,
		_w8859_
	);
	LUT2 #(
		.INIT('h1)
	) name7110 (
		_w8857_,
		_w8859_,
		_w8860_
	);
	LUT4 #(
		.INIT('h0002)
	) name7111 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		\wb_data_i[3]_pad ,
		_w8861_
	);
	LUT2 #(
		.INIT('h8)
	) name7112 (
		_w8842_,
		_w8861_,
		_w8862_
	);
	LUT2 #(
		.INIT('h8)
	) name7113 (
		rst_i_pad,
		\u4_funct_adr_reg[3]/P0001 ,
		_w8863_
	);
	LUT3 #(
		.INIT('h07)
	) name7114 (
		_w8846_,
		_w8848_,
		_w8863_,
		_w8864_
	);
	LUT2 #(
		.INIT('h1)
	) name7115 (
		_w8862_,
		_w8864_,
		_w8865_
	);
	LUT4 #(
		.INIT('h0002)
	) name7116 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		\wb_data_i[4]_pad ,
		_w8866_
	);
	LUT2 #(
		.INIT('h8)
	) name7117 (
		_w8842_,
		_w8866_,
		_w8867_
	);
	LUT2 #(
		.INIT('h8)
	) name7118 (
		rst_i_pad,
		\u4_funct_adr_reg[4]/P0001 ,
		_w8868_
	);
	LUT3 #(
		.INIT('h07)
	) name7119 (
		_w8846_,
		_w8848_,
		_w8868_,
		_w8869_
	);
	LUT2 #(
		.INIT('h1)
	) name7120 (
		_w8867_,
		_w8869_,
		_w8870_
	);
	LUT4 #(
		.INIT('h0002)
	) name7121 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		\wb_data_i[5]_pad ,
		_w8871_
	);
	LUT2 #(
		.INIT('h8)
	) name7122 (
		_w8842_,
		_w8871_,
		_w8872_
	);
	LUT2 #(
		.INIT('h8)
	) name7123 (
		rst_i_pad,
		\u4_funct_adr_reg[5]/P0001 ,
		_w8873_
	);
	LUT3 #(
		.INIT('h07)
	) name7124 (
		_w8846_,
		_w8848_,
		_w8873_,
		_w8874_
	);
	LUT2 #(
		.INIT('h1)
	) name7125 (
		_w8872_,
		_w8874_,
		_w8875_
	);
	LUT4 #(
		.INIT('h0002)
	) name7126 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		\wb_data_i[6]_pad ,
		_w8876_
	);
	LUT2 #(
		.INIT('h8)
	) name7127 (
		_w8842_,
		_w8876_,
		_w8877_
	);
	LUT2 #(
		.INIT('h8)
	) name7128 (
		rst_i_pad,
		\u4_funct_adr_reg[6]/P0001 ,
		_w8878_
	);
	LUT3 #(
		.INIT('h07)
	) name7129 (
		_w8846_,
		_w8848_,
		_w8878_,
		_w8879_
	);
	LUT2 #(
		.INIT('h1)
	) name7130 (
		_w8877_,
		_w8879_,
		_w8880_
	);
	LUT4 #(
		.INIT('h0004)
	) name7131 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		\wb_data_i[0]_pad ,
		_w8881_
	);
	LUT2 #(
		.INIT('h8)
	) name7132 (
		_w8842_,
		_w8881_,
		_w8882_
	);
	LUT2 #(
		.INIT('h8)
	) name7133 (
		rst_i_pad,
		\u4_inta_msk_reg[0]/P0001 ,
		_w8883_
	);
	LUT3 #(
		.INIT('h04)
	) name7134 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w8884_
	);
	LUT3 #(
		.INIT('h13)
	) name7135 (
		_w8848_,
		_w8883_,
		_w8884_,
		_w8885_
	);
	LUT2 #(
		.INIT('h1)
	) name7136 (
		_w8882_,
		_w8885_,
		_w8886_
	);
	LUT4 #(
		.INIT('h0004)
	) name7137 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		\wb_data_i[1]_pad ,
		_w8887_
	);
	LUT2 #(
		.INIT('h8)
	) name7138 (
		_w8842_,
		_w8887_,
		_w8888_
	);
	LUT2 #(
		.INIT('h8)
	) name7139 (
		rst_i_pad,
		\u4_inta_msk_reg[1]/P0001 ,
		_w8889_
	);
	LUT3 #(
		.INIT('h07)
	) name7140 (
		_w8848_,
		_w8884_,
		_w8889_,
		_w8890_
	);
	LUT2 #(
		.INIT('h1)
	) name7141 (
		_w8888_,
		_w8890_,
		_w8891_
	);
	LUT4 #(
		.INIT('h0004)
	) name7142 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		\wb_data_i[2]_pad ,
		_w8892_
	);
	LUT2 #(
		.INIT('h8)
	) name7143 (
		_w8842_,
		_w8892_,
		_w8893_
	);
	LUT2 #(
		.INIT('h8)
	) name7144 (
		rst_i_pad,
		\u4_inta_msk_reg[2]/P0001 ,
		_w8894_
	);
	LUT3 #(
		.INIT('h07)
	) name7145 (
		_w8848_,
		_w8884_,
		_w8894_,
		_w8895_
	);
	LUT2 #(
		.INIT('h1)
	) name7146 (
		_w8893_,
		_w8895_,
		_w8896_
	);
	LUT4 #(
		.INIT('h0004)
	) name7147 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		\wb_data_i[3]_pad ,
		_w8897_
	);
	LUT2 #(
		.INIT('h8)
	) name7148 (
		_w8842_,
		_w8897_,
		_w8898_
	);
	LUT2 #(
		.INIT('h8)
	) name7149 (
		rst_i_pad,
		\u4_inta_msk_reg[3]/P0001 ,
		_w8899_
	);
	LUT3 #(
		.INIT('h07)
	) name7150 (
		_w8848_,
		_w8884_,
		_w8899_,
		_w8900_
	);
	LUT2 #(
		.INIT('h1)
	) name7151 (
		_w8898_,
		_w8900_,
		_w8901_
	);
	LUT4 #(
		.INIT('h0004)
	) name7152 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		\wb_data_i[4]_pad ,
		_w8902_
	);
	LUT2 #(
		.INIT('h8)
	) name7153 (
		_w8842_,
		_w8902_,
		_w8903_
	);
	LUT2 #(
		.INIT('h8)
	) name7154 (
		rst_i_pad,
		\u4_inta_msk_reg[4]/P0001 ,
		_w8904_
	);
	LUT3 #(
		.INIT('h07)
	) name7155 (
		_w8848_,
		_w8884_,
		_w8904_,
		_w8905_
	);
	LUT2 #(
		.INIT('h1)
	) name7156 (
		_w8903_,
		_w8905_,
		_w8906_
	);
	LUT4 #(
		.INIT('h0004)
	) name7157 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		\wb_data_i[5]_pad ,
		_w8907_
	);
	LUT2 #(
		.INIT('h8)
	) name7158 (
		_w8842_,
		_w8907_,
		_w8908_
	);
	LUT2 #(
		.INIT('h8)
	) name7159 (
		rst_i_pad,
		\u4_inta_msk_reg[5]/P0001 ,
		_w8909_
	);
	LUT3 #(
		.INIT('h07)
	) name7160 (
		_w8848_,
		_w8884_,
		_w8909_,
		_w8910_
	);
	LUT2 #(
		.INIT('h1)
	) name7161 (
		_w8908_,
		_w8910_,
		_w8911_
	);
	LUT4 #(
		.INIT('h0004)
	) name7162 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		\wb_data_i[6]_pad ,
		_w8912_
	);
	LUT2 #(
		.INIT('h8)
	) name7163 (
		_w8842_,
		_w8912_,
		_w8913_
	);
	LUT2 #(
		.INIT('h8)
	) name7164 (
		rst_i_pad,
		\u4_inta_msk_reg[6]/P0001 ,
		_w8914_
	);
	LUT3 #(
		.INIT('h07)
	) name7165 (
		_w8848_,
		_w8884_,
		_w8914_,
		_w8915_
	);
	LUT2 #(
		.INIT('h1)
	) name7166 (
		_w8913_,
		_w8915_,
		_w8916_
	);
	LUT4 #(
		.INIT('h0004)
	) name7167 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		\wb_data_i[7]_pad ,
		_w8917_
	);
	LUT2 #(
		.INIT('h8)
	) name7168 (
		_w8842_,
		_w8917_,
		_w8918_
	);
	LUT2 #(
		.INIT('h8)
	) name7169 (
		rst_i_pad,
		\u4_inta_msk_reg[7]/P0001 ,
		_w8919_
	);
	LUT3 #(
		.INIT('h07)
	) name7170 (
		_w8848_,
		_w8884_,
		_w8919_,
		_w8920_
	);
	LUT2 #(
		.INIT('h1)
	) name7171 (
		_w8918_,
		_w8920_,
		_w8921_
	);
	LUT4 #(
		.INIT('h0004)
	) name7172 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		\wb_data_i[8]_pad ,
		_w8922_
	);
	LUT2 #(
		.INIT('h8)
	) name7173 (
		_w8842_,
		_w8922_,
		_w8923_
	);
	LUT2 #(
		.INIT('h8)
	) name7174 (
		rst_i_pad,
		\u4_inta_msk_reg[8]/P0001 ,
		_w8924_
	);
	LUT3 #(
		.INIT('h07)
	) name7175 (
		_w8848_,
		_w8884_,
		_w8924_,
		_w8925_
	);
	LUT2 #(
		.INIT('h1)
	) name7176 (
		_w8923_,
		_w8925_,
		_w8926_
	);
	LUT4 #(
		.INIT('h0004)
	) name7177 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		\wb_data_i[16]_pad ,
		_w8927_
	);
	LUT2 #(
		.INIT('h8)
	) name7178 (
		_w8842_,
		_w8927_,
		_w8928_
	);
	LUT2 #(
		.INIT('h8)
	) name7179 (
		rst_i_pad,
		\u4_intb_msk_reg[0]/P0001 ,
		_w8929_
	);
	LUT3 #(
		.INIT('h07)
	) name7180 (
		_w8848_,
		_w8884_,
		_w8929_,
		_w8930_
	);
	LUT2 #(
		.INIT('h1)
	) name7181 (
		_w8928_,
		_w8930_,
		_w8931_
	);
	LUT4 #(
		.INIT('h0004)
	) name7182 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		\wb_data_i[17]_pad ,
		_w8932_
	);
	LUT2 #(
		.INIT('h8)
	) name7183 (
		_w8842_,
		_w8932_,
		_w8933_
	);
	LUT2 #(
		.INIT('h8)
	) name7184 (
		rst_i_pad,
		\u4_intb_msk_reg[1]/P0001 ,
		_w8934_
	);
	LUT3 #(
		.INIT('h07)
	) name7185 (
		_w8848_,
		_w8884_,
		_w8934_,
		_w8935_
	);
	LUT2 #(
		.INIT('h1)
	) name7186 (
		_w8933_,
		_w8935_,
		_w8936_
	);
	LUT4 #(
		.INIT('h0004)
	) name7187 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		\wb_data_i[18]_pad ,
		_w8937_
	);
	LUT2 #(
		.INIT('h8)
	) name7188 (
		_w8842_,
		_w8937_,
		_w8938_
	);
	LUT2 #(
		.INIT('h8)
	) name7189 (
		rst_i_pad,
		\u4_intb_msk_reg[2]/P0001 ,
		_w8939_
	);
	LUT3 #(
		.INIT('h07)
	) name7190 (
		_w8848_,
		_w8884_,
		_w8939_,
		_w8940_
	);
	LUT2 #(
		.INIT('h1)
	) name7191 (
		_w8938_,
		_w8940_,
		_w8941_
	);
	LUT4 #(
		.INIT('h0004)
	) name7192 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		\wb_data_i[19]_pad ,
		_w8942_
	);
	LUT2 #(
		.INIT('h8)
	) name7193 (
		_w8842_,
		_w8942_,
		_w8943_
	);
	LUT2 #(
		.INIT('h8)
	) name7194 (
		rst_i_pad,
		\u4_intb_msk_reg[3]/P0001 ,
		_w8944_
	);
	LUT3 #(
		.INIT('h07)
	) name7195 (
		_w8848_,
		_w8884_,
		_w8944_,
		_w8945_
	);
	LUT2 #(
		.INIT('h1)
	) name7196 (
		_w8943_,
		_w8945_,
		_w8946_
	);
	LUT4 #(
		.INIT('h0004)
	) name7197 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		\wb_data_i[20]_pad ,
		_w8947_
	);
	LUT2 #(
		.INIT('h8)
	) name7198 (
		_w8842_,
		_w8947_,
		_w8948_
	);
	LUT2 #(
		.INIT('h8)
	) name7199 (
		rst_i_pad,
		\u4_intb_msk_reg[4]/P0001 ,
		_w8949_
	);
	LUT3 #(
		.INIT('h07)
	) name7200 (
		_w8848_,
		_w8884_,
		_w8949_,
		_w8950_
	);
	LUT2 #(
		.INIT('h1)
	) name7201 (
		_w8948_,
		_w8950_,
		_w8951_
	);
	LUT4 #(
		.INIT('h0004)
	) name7202 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		\wb_data_i[21]_pad ,
		_w8952_
	);
	LUT2 #(
		.INIT('h8)
	) name7203 (
		_w8842_,
		_w8952_,
		_w8953_
	);
	LUT2 #(
		.INIT('h8)
	) name7204 (
		rst_i_pad,
		\u4_intb_msk_reg[5]/P0001 ,
		_w8954_
	);
	LUT3 #(
		.INIT('h07)
	) name7205 (
		_w8848_,
		_w8884_,
		_w8954_,
		_w8955_
	);
	LUT2 #(
		.INIT('h1)
	) name7206 (
		_w8953_,
		_w8955_,
		_w8956_
	);
	LUT4 #(
		.INIT('h0004)
	) name7207 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		\wb_data_i[22]_pad ,
		_w8957_
	);
	LUT2 #(
		.INIT('h8)
	) name7208 (
		_w8842_,
		_w8957_,
		_w8958_
	);
	LUT2 #(
		.INIT('h8)
	) name7209 (
		rst_i_pad,
		\u4_intb_msk_reg[6]/P0001 ,
		_w8959_
	);
	LUT3 #(
		.INIT('h07)
	) name7210 (
		_w8848_,
		_w8884_,
		_w8959_,
		_w8960_
	);
	LUT2 #(
		.INIT('h1)
	) name7211 (
		_w8958_,
		_w8960_,
		_w8961_
	);
	LUT4 #(
		.INIT('h0004)
	) name7212 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		\wb_data_i[23]_pad ,
		_w8962_
	);
	LUT2 #(
		.INIT('h8)
	) name7213 (
		_w8842_,
		_w8962_,
		_w8963_
	);
	LUT2 #(
		.INIT('h8)
	) name7214 (
		rst_i_pad,
		\u4_intb_msk_reg[7]/P0001 ,
		_w8964_
	);
	LUT3 #(
		.INIT('h07)
	) name7215 (
		_w8848_,
		_w8884_,
		_w8964_,
		_w8965_
	);
	LUT2 #(
		.INIT('h1)
	) name7216 (
		_w8963_,
		_w8965_,
		_w8966_
	);
	LUT4 #(
		.INIT('h0004)
	) name7217 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		\wb_data_i[24]_pad ,
		_w8967_
	);
	LUT2 #(
		.INIT('h8)
	) name7218 (
		_w8842_,
		_w8967_,
		_w8968_
	);
	LUT2 #(
		.INIT('h8)
	) name7219 (
		rst_i_pad,
		\u4_intb_msk_reg[8]/P0001 ,
		_w8969_
	);
	LUT3 #(
		.INIT('h07)
	) name7220 (
		_w8848_,
		_w8884_,
		_w8969_,
		_w8970_
	);
	LUT2 #(
		.INIT('h1)
	) name7221 (
		_w8968_,
		_w8970_,
		_w8971_
	);
	LUT3 #(
		.INIT('h80)
	) name7222 (
		\u1_u3_rx_ack_to_cnt_reg[4]/P0001 ,
		\u1_u3_rx_ack_to_cnt_reg[5]/P0001 ,
		\u1_u3_rx_ack_to_cnt_reg[6]/P0001 ,
		_w8972_
	);
	LUT2 #(
		.INIT('h4)
	) name7223 (
		\u1_u3_rx_ack_to_clr_reg/P0001 ,
		\u1_u3_rx_ack_to_cnt_reg[7]/P0001 ,
		_w8973_
	);
	LUT3 #(
		.INIT('h70)
	) name7224 (
		_w7951_,
		_w8972_,
		_w8973_,
		_w8974_
	);
	LUT4 #(
		.INIT('h4000)
	) name7225 (
		\u1_u3_rx_ack_to_clr_reg/P0001 ,
		\u1_u3_rx_ack_to_cnt_reg[4]/P0001 ,
		\u1_u3_rx_ack_to_cnt_reg[5]/P0001 ,
		\u1_u3_rx_ack_to_cnt_reg[6]/P0001 ,
		_w8975_
	);
	LUT3 #(
		.INIT('h40)
	) name7226 (
		\u1_u3_rx_ack_to_cnt_reg[7]/P0001 ,
		_w7951_,
		_w8975_,
		_w8976_
	);
	LUT2 #(
		.INIT('he)
	) name7227 (
		_w8974_,
		_w8976_,
		_w8977_
	);
	LUT3 #(
		.INIT('h80)
	) name7228 (
		\u1_u3_tx_data_to_cnt_reg[4]/P0001 ,
		\u1_u3_tx_data_to_cnt_reg[5]/P0001 ,
		\u1_u3_tx_data_to_cnt_reg[6]/P0001 ,
		_w8978_
	);
	LUT4 #(
		.INIT('h1444)
	) name7229 (
		\u0_rx_active_reg/P0001 ,
		\u1_u3_tx_data_to_cnt_reg[7]/P0001 ,
		_w7967_,
		_w8978_,
		_w8979_
	);
	LUT4 #(
		.INIT('h2220)
	) name7230 (
		rst_i_pad,
		\u4_int_src_re_reg/P0001 ,
		\u4_int_srcb_reg[1]/P0001 ,
		\u4_pid_cs_err_r_reg/P0001 ,
		_w8980_
	);
	LUT4 #(
		.INIT('h2220)
	) name7231 (
		rst_i_pad,
		\u4_int_src_re_reg/P0001 ,
		\u4_int_srcb_reg[7]/P0001 ,
		\u4_rx_err_r_reg/P0001 ,
		_w8981_
	);
	LUT4 #(
		.INIT('h2220)
	) name7232 (
		rst_i_pad,
		\u4_int_src_re_reg/P0001 ,
		\u4_int_srcb_reg[8]/P0001 ,
		\u4_usb_reset_r_reg/P0001 ,
		_w8982_
	);
	LUT4 #(
		.INIT('h0004)
	) name7233 (
		\u0_u0_state_reg[11]/NET0131 ,
		\u0_u0_state_reg[12]/NET0131 ,
		\u0_u0_state_reg[1]/P0001 ,
		\u0_u0_state_reg[2]/NET0131 ,
		_w8983_
	);
	LUT4 #(
		.INIT('h8000)
	) name7234 (
		_w4098_,
		_w4108_,
		_w4109_,
		_w8983_,
		_w8984_
	);
	LUT4 #(
		.INIT('hef00)
	) name7235 (
		\LineState_r_reg[0]/P0001 ,
		\LineState_r_reg[1]/P0001 ,
		\u0_u0_ls_se0_r_reg/P0001 ,
		\u0_u0_state_reg[13]/NET0131 ,
		_w8985_
	);
	LUT3 #(
		.INIT('h45)
	) name7236 (
		\u0_u0_chirp_cnt_is_6_reg/P0001 ,
		_w4112_,
		_w8985_,
		_w8986_
	);
	LUT2 #(
		.INIT('h2)
	) name7237 (
		_w8984_,
		_w8986_,
		_w8987_
	);
	LUT3 #(
		.INIT('h02)
	) name7238 (
		\u0_u0_state_reg[13]/NET0131 ,
		\u0_u0_state_reg[14]/P0001 ,
		\u0_u0_state_reg[9]/P0001 ,
		_w8988_
	);
	LUT2 #(
		.INIT('h4)
	) name7239 (
		_w4117_,
		_w8988_,
		_w8989_
	);
	LUT4 #(
		.INIT('h0002)
	) name7240 (
		\u0_u0_state_reg[11]/NET0131 ,
		\u0_u0_state_reg[12]/NET0131 ,
		\u0_u0_state_reg[1]/P0001 ,
		\u0_u0_state_reg[2]/NET0131 ,
		_w8990_
	);
	LUT4 #(
		.INIT('h8000)
	) name7241 (
		_w4098_,
		_w4108_,
		_w4109_,
		_w8990_,
		_w8991_
	);
	LUT3 #(
		.INIT('h45)
	) name7242 (
		\u0_u0_chirp_cnt_is_6_reg/P0001 ,
		_w4119_,
		_w8985_,
		_w8992_
	);
	LUT4 #(
		.INIT('h7707)
	) name7243 (
		_w7957_,
		_w8989_,
		_w8991_,
		_w8992_,
		_w8993_
	);
	LUT3 #(
		.INIT('h8a)
	) name7244 (
		_w4103_,
		_w8987_,
		_w8993_,
		_w8994_
	);
	LUT4 #(
		.INIT('h0008)
	) name7245 (
		rst_i_pad,
		\u0_u0_state_reg[3]/P0001 ,
		\u0_u0_state_reg[6]/NET0131 ,
		usb_vbus_pad_i_pad,
		_w8995_
	);
	LUT4 #(
		.INIT('h0100)
	) name7246 (
		_w4119_,
		_w4354_,
		_w8112_,
		_w8995_,
		_w8996_
	);
	LUT2 #(
		.INIT('h8)
	) name7247 (
		_w7962_,
		_w8996_,
		_w8997_
	);
	LUT4 #(
		.INIT('h3f37)
	) name7248 (
		\u0_u0_state_reg[3]/P0001 ,
		_w4345_,
		_w4355_,
		_w4356_,
		_w8998_
	);
	LUT4 #(
		.INIT('h8088)
	) name7249 (
		_w4103_,
		_w5763_,
		_w5767_,
		_w8998_,
		_w8999_
	);
	LUT2 #(
		.INIT('he)
	) name7250 (
		_w8997_,
		_w8999_,
		_w9000_
	);
	LUT4 #(
		.INIT('h00e0)
	) name7251 (
		resume_req_i_pad,
		\resume_req_r_reg/P0001 ,
		rst_i_pad,
		\suspend_clr_wr_reg/P0001 ,
		_w9001_
	);
	LUT4 #(
		.INIT('h8acf)
	) name7252 (
		\u4_u0_buf0_orig_reg[28]/P0001 ,
		\u4_u0_buf0_orig_reg[29]/NET0131 ,
		\u4_u0_dma_out_cnt_reg[10]/P0001 ,
		\u4_u0_dma_out_cnt_reg[9]/P0001 ,
		_w9002_
	);
	LUT4 #(
		.INIT('hea00)
	) name7253 (
		_w5973_,
		_w5985_,
		_w5987_,
		_w9002_,
		_w9003_
	);
	LUT4 #(
		.INIT('h008a)
	) name7254 (
		\u4_u0_buf0_orig_reg[28]/P0001 ,
		\u4_u0_buf0_orig_reg[29]/NET0131 ,
		\u4_u0_dma_out_cnt_reg[10]/P0001 ,
		\u4_u0_dma_out_cnt_reg[9]/P0001 ,
		_w9004_
	);
	LUT2 #(
		.INIT('h9)
	) name7255 (
		\u4_u0_buf0_orig_reg[30]/NET0131 ,
		\u4_u0_dma_out_cnt_reg[11]/P0001 ,
		_w9005_
	);
	LUT4 #(
		.INIT('h01fe)
	) name7256 (
		_w5989_,
		_w9003_,
		_w9004_,
		_w9005_,
		_w9006_
	);
	LUT4 #(
		.INIT('h8acf)
	) name7257 (
		\u4_u3_buf0_orig_reg[28]/P0001 ,
		\u4_u3_buf0_orig_reg[29]/NET0131 ,
		\u4_u3_dma_out_cnt_reg[10]/P0001 ,
		\u4_u3_dma_out_cnt_reg[9]/P0001 ,
		_w9007_
	);
	LUT4 #(
		.INIT('hea00)
	) name7258 (
		_w5948_,
		_w5960_,
		_w5962_,
		_w9007_,
		_w9008_
	);
	LUT4 #(
		.INIT('h008a)
	) name7259 (
		\u4_u3_buf0_orig_reg[28]/P0001 ,
		\u4_u3_buf0_orig_reg[29]/NET0131 ,
		\u4_u3_dma_out_cnt_reg[10]/P0001 ,
		\u4_u3_dma_out_cnt_reg[9]/P0001 ,
		_w9009_
	);
	LUT2 #(
		.INIT('h9)
	) name7260 (
		\u4_u3_buf0_orig_reg[30]/NET0131 ,
		\u4_u3_dma_out_cnt_reg[11]/P0001 ,
		_w9010_
	);
	LUT4 #(
		.INIT('h01fe)
	) name7261 (
		_w5964_,
		_w9008_,
		_w9009_,
		_w9010_,
		_w9011_
	);
	LUT3 #(
		.INIT('hac)
	) name7262 (
		\sram_data_i[10]_pad ,
		\u4_dout_reg[10]/P0001 ,
		\wb_addr_i[17]_pad ,
		_w9012_
	);
	LUT3 #(
		.INIT('hac)
	) name7263 (
		\sram_data_i[11]_pad ,
		\u4_dout_reg[11]/P0001 ,
		\wb_addr_i[17]_pad ,
		_w9013_
	);
	LUT3 #(
		.INIT('hac)
	) name7264 (
		\sram_data_i[9]_pad ,
		\u4_dout_reg[9]/P0001 ,
		\wb_addr_i[17]_pad ,
		_w9014_
	);
	LUT4 #(
		.INIT('h8000)
	) name7265 (
		\u0_u0_idle_cnt1_reg[0]/P0001 ,
		\u0_u0_idle_cnt1_reg[1]/P0001 ,
		\u0_u0_idle_cnt1_reg[2]/P0001 ,
		\u0_u0_idle_cnt1_reg[3]/P0001 ,
		_w9015_
	);
	LUT2 #(
		.INIT('h6)
	) name7266 (
		\u0_u0_idle_cnt1_reg[4]/P0001 ,
		_w9015_,
		_w9016_
	);
	LUT4 #(
		.INIT('h8acf)
	) name7267 (
		\u4_u1_buf0_orig_reg[28]/P0001 ,
		\u4_u1_buf0_orig_reg[29]/NET0131 ,
		\u4_u1_dma_out_cnt_reg[10]/P0001 ,
		\u4_u1_dma_out_cnt_reg[9]/P0001 ,
		_w9017_
	);
	LUT4 #(
		.INIT('hea00)
	) name7268 (
		_w5998_,
		_w6010_,
		_w6012_,
		_w9017_,
		_w9018_
	);
	LUT4 #(
		.INIT('h008a)
	) name7269 (
		\u4_u1_buf0_orig_reg[28]/P0001 ,
		\u4_u1_buf0_orig_reg[29]/NET0131 ,
		\u4_u1_dma_out_cnt_reg[10]/P0001 ,
		\u4_u1_dma_out_cnt_reg[9]/P0001 ,
		_w9019_
	);
	LUT2 #(
		.INIT('h9)
	) name7270 (
		\u4_u1_buf0_orig_reg[30]/NET0131 ,
		\u4_u1_dma_out_cnt_reg[11]/P0001 ,
		_w9020_
	);
	LUT4 #(
		.INIT('h01fe)
	) name7271 (
		_w6014_,
		_w9018_,
		_w9019_,
		_w9020_,
		_w9021_
	);
	LUT4 #(
		.INIT('h8acf)
	) name7272 (
		\u4_u2_buf0_orig_reg[28]/P0001 ,
		\u4_u2_buf0_orig_reg[29]/NET0131 ,
		\u4_u2_dma_out_cnt_reg[10]/P0001 ,
		\u4_u2_dma_out_cnt_reg[9]/P0001 ,
		_w9022_
	);
	LUT2 #(
		.INIT('h9)
	) name7273 (
		\u4_u2_buf0_orig_reg[30]/NET0131 ,
		\u4_u2_dma_out_cnt_reg[11]/P0001 ,
		_w9023_
	);
	LUT4 #(
		.INIT('hc431)
	) name7274 (
		\u4_u2_buf0_orig_reg[29]/NET0131 ,
		\u4_u2_buf0_orig_reg[30]/NET0131 ,
		\u4_u2_dma_out_cnt_reg[10]/P0001 ,
		\u4_u2_dma_out_cnt_reg[11]/P0001 ,
		_w9024_
	);
	LUT2 #(
		.INIT('h4)
	) name7275 (
		_w9022_,
		_w9024_,
		_w9025_
	);
	LUT2 #(
		.INIT('h4)
	) name7276 (
		_w6040_,
		_w9024_,
		_w9026_
	);
	LUT4 #(
		.INIT('h1500)
	) name7277 (
		_w6023_,
		_w6035_,
		_w6037_,
		_w9026_,
		_w9027_
	);
	LUT2 #(
		.INIT('h1)
	) name7278 (
		_w9025_,
		_w9027_,
		_w9028_
	);
	LUT4 #(
		.INIT('h7130)
	) name7279 (
		\u4_u2_buf0_orig_reg[28]/P0001 ,
		\u4_u2_buf0_orig_reg[29]/NET0131 ,
		\u4_u2_dma_out_cnt_reg[10]/P0001 ,
		\u4_u2_dma_out_cnt_reg[9]/P0001 ,
		_w9029_
	);
	LUT4 #(
		.INIT('hf351)
	) name7280 (
		\u4_u2_buf0_orig_reg[28]/P0001 ,
		\u4_u2_buf0_orig_reg[29]/NET0131 ,
		\u4_u2_dma_out_cnt_reg[10]/P0001 ,
		\u4_u2_dma_out_cnt_reg[9]/P0001 ,
		_w9030_
	);
	LUT4 #(
		.INIT('h1500)
	) name7281 (
		_w6023_,
		_w6035_,
		_w6037_,
		_w9030_,
		_w9031_
	);
	LUT3 #(
		.INIT('h01)
	) name7282 (
		_w9023_,
		_w9029_,
		_w9031_,
		_w9032_
	);
	LUT2 #(
		.INIT('hd)
	) name7283 (
		_w9028_,
		_w9032_,
		_w9033_
	);
	LUT2 #(
		.INIT('h9)
	) name7284 (
		\u4_u2_buf0_orig_reg[25]/P0001 ,
		\u4_u2_dma_out_cnt_reg[6]/P0001 ,
		_w9034_
	);
	LUT4 #(
		.INIT('h1040)
	) name7285 (
		\u4_u2_buf0_orig_reg[24]/P0001 ,
		\u4_u2_buf0_orig_reg[25]/P0001 ,
		\u4_u2_dma_out_cnt_reg[5]/P0001 ,
		\u4_u2_dma_out_cnt_reg[6]/P0001 ,
		_w9035_
	);
	LUT2 #(
		.INIT('h2)
	) name7286 (
		_w6033_,
		_w9034_,
		_w9036_
	);
	LUT4 #(
		.INIT('h0e0f)
	) name7287 (
		_w6027_,
		_w6031_,
		_w9035_,
		_w9036_,
		_w9037_
	);
	LUT4 #(
		.INIT('h8c23)
	) name7288 (
		\u4_u2_buf0_orig_reg[24]/P0001 ,
		\u4_u2_buf0_orig_reg[25]/P0001 ,
		\u4_u2_dma_out_cnt_reg[5]/P0001 ,
		\u4_u2_dma_out_cnt_reg[6]/P0001 ,
		_w9038_
	);
	LUT4 #(
		.INIT('hef00)
	) name7289 (
		_w6027_,
		_w6031_,
		_w6033_,
		_w9038_,
		_w9039_
	);
	LUT2 #(
		.INIT('h2)
	) name7290 (
		_w9037_,
		_w9039_,
		_w9040_
	);
	LUT2 #(
		.INIT('h9)
	) name7291 (
		\u4_u3_buf0_orig_reg[25]/P0001 ,
		\u4_u3_dma_out_cnt_reg[6]/P0001 ,
		_w9041_
	);
	LUT4 #(
		.INIT('h1040)
	) name7292 (
		\u4_u3_buf0_orig_reg[24]/P0001 ,
		\u4_u3_buf0_orig_reg[25]/P0001 ,
		\u4_u3_dma_out_cnt_reg[5]/P0001 ,
		\u4_u3_dma_out_cnt_reg[6]/P0001 ,
		_w9042_
	);
	LUT2 #(
		.INIT('h2)
	) name7293 (
		_w5958_,
		_w9041_,
		_w9043_
	);
	LUT4 #(
		.INIT('h0e0f)
	) name7294 (
		_w5952_,
		_w5956_,
		_w9042_,
		_w9043_,
		_w9044_
	);
	LUT4 #(
		.INIT('h8c23)
	) name7295 (
		\u4_u3_buf0_orig_reg[24]/P0001 ,
		\u4_u3_buf0_orig_reg[25]/P0001 ,
		\u4_u3_dma_out_cnt_reg[5]/P0001 ,
		\u4_u3_dma_out_cnt_reg[6]/P0001 ,
		_w9045_
	);
	LUT4 #(
		.INIT('hef00)
	) name7296 (
		_w5952_,
		_w5956_,
		_w5958_,
		_w9045_,
		_w9046_
	);
	LUT2 #(
		.INIT('h2)
	) name7297 (
		_w9044_,
		_w9046_,
		_w9047_
	);
	LUT2 #(
		.INIT('h9)
	) name7298 (
		\u4_u0_buf0_orig_reg[25]/P0001 ,
		\u4_u0_dma_out_cnt_reg[6]/P0001 ,
		_w9048_
	);
	LUT4 #(
		.INIT('h1040)
	) name7299 (
		\u4_u0_buf0_orig_reg[24]/P0001 ,
		\u4_u0_buf0_orig_reg[25]/P0001 ,
		\u4_u0_dma_out_cnt_reg[5]/P0001 ,
		\u4_u0_dma_out_cnt_reg[6]/P0001 ,
		_w9049_
	);
	LUT2 #(
		.INIT('h2)
	) name7300 (
		_w5983_,
		_w9048_,
		_w9050_
	);
	LUT4 #(
		.INIT('h0e0f)
	) name7301 (
		_w5977_,
		_w5981_,
		_w9049_,
		_w9050_,
		_w9051_
	);
	LUT4 #(
		.INIT('h8c23)
	) name7302 (
		\u4_u0_buf0_orig_reg[24]/P0001 ,
		\u4_u0_buf0_orig_reg[25]/P0001 ,
		\u4_u0_dma_out_cnt_reg[5]/P0001 ,
		\u4_u0_dma_out_cnt_reg[6]/P0001 ,
		_w9052_
	);
	LUT4 #(
		.INIT('hef00)
	) name7303 (
		_w5977_,
		_w5981_,
		_w5983_,
		_w9052_,
		_w9053_
	);
	LUT2 #(
		.INIT('h2)
	) name7304 (
		_w9051_,
		_w9053_,
		_w9054_
	);
	LUT2 #(
		.INIT('h9)
	) name7305 (
		\u4_u1_buf0_orig_reg[25]/P0001 ,
		\u4_u1_dma_out_cnt_reg[6]/P0001 ,
		_w9055_
	);
	LUT4 #(
		.INIT('h1040)
	) name7306 (
		\u4_u1_buf0_orig_reg[24]/P0001 ,
		\u4_u1_buf0_orig_reg[25]/P0001 ,
		\u4_u1_dma_out_cnt_reg[5]/P0001 ,
		\u4_u1_dma_out_cnt_reg[6]/P0001 ,
		_w9056_
	);
	LUT2 #(
		.INIT('h2)
	) name7307 (
		_w6008_,
		_w9055_,
		_w9057_
	);
	LUT4 #(
		.INIT('h0e0f)
	) name7308 (
		_w6002_,
		_w6006_,
		_w9056_,
		_w9057_,
		_w9058_
	);
	LUT4 #(
		.INIT('h8c23)
	) name7309 (
		\u4_u1_buf0_orig_reg[24]/P0001 ,
		\u4_u1_buf0_orig_reg[25]/P0001 ,
		\u4_u1_dma_out_cnt_reg[5]/P0001 ,
		\u4_u1_dma_out_cnt_reg[6]/P0001 ,
		_w9059_
	);
	LUT4 #(
		.INIT('hef00)
	) name7310 (
		_w6002_,
		_w6006_,
		_w6008_,
		_w9059_,
		_w9060_
	);
	LUT2 #(
		.INIT('h2)
	) name7311 (
		_w9058_,
		_w9060_,
		_w9061_
	);
	LUT3 #(
		.INIT('h59)
	) name7312 (
		\u1_u3_adr_reg[0]/P0001 ,
		_w2788_,
		_w2790_,
		_w9062_
	);
	LUT2 #(
		.INIT('h6)
	) name7313 (
		\u4_u3_buf0_orig_reg[23]/P0001 ,
		_w7822_,
		_w9063_
	);
	LUT2 #(
		.INIT('h6)
	) name7314 (
		\u4_u0_buf0_orig_reg[23]/P0001 ,
		_w7835_,
		_w9064_
	);
	LUT2 #(
		.INIT('h6)
	) name7315 (
		\u4_u1_buf0_orig_reg[23]/P0001 ,
		_w7845_,
		_w9065_
	);
	LUT2 #(
		.INIT('h6)
	) name7316 (
		\u4_u2_buf0_orig_reg[23]/P0001 ,
		_w7853_,
		_w9066_
	);
	LUT3 #(
		.INIT('h02)
	) name7317 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_data_i[24]_pad ,
		_w9067_
	);
	LUT2 #(
		.INIT('h8)
	) name7318 (
		rst_i_pad,
		\u4_u2_iena_reg[0]/P0001 ,
		_w9068_
	);
	LUT3 #(
		.INIT('h08)
	) name7319 (
		rst_i_pad,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w9069_
	);
	LUT4 #(
		.INIT('h7270)
	) name7320 (
		_w2267_,
		_w9067_,
		_w9068_,
		_w9069_,
		_w9070_
	);
	LUT3 #(
		.INIT('h02)
	) name7321 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_data_i[25]_pad ,
		_w9071_
	);
	LUT2 #(
		.INIT('h8)
	) name7322 (
		rst_i_pad,
		\u4_u2_iena_reg[1]/P0001 ,
		_w9072_
	);
	LUT4 #(
		.INIT('h5f08)
	) name7323 (
		_w2267_,
		_w9069_,
		_w9071_,
		_w9072_,
		_w9073_
	);
	LUT3 #(
		.INIT('h02)
	) name7324 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_data_i[26]_pad ,
		_w9074_
	);
	LUT2 #(
		.INIT('h8)
	) name7325 (
		rst_i_pad,
		\u4_u2_iena_reg[2]/P0001 ,
		_w9075_
	);
	LUT4 #(
		.INIT('h5f08)
	) name7326 (
		_w2267_,
		_w9069_,
		_w9074_,
		_w9075_,
		_w9076_
	);
	LUT3 #(
		.INIT('h02)
	) name7327 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_data_i[27]_pad ,
		_w9077_
	);
	LUT2 #(
		.INIT('h8)
	) name7328 (
		rst_i_pad,
		\u4_u2_iena_reg[3]/P0001 ,
		_w9078_
	);
	LUT4 #(
		.INIT('h5f08)
	) name7329 (
		_w2267_,
		_w9069_,
		_w9077_,
		_w9078_,
		_w9079_
	);
	LUT3 #(
		.INIT('h02)
	) name7330 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_data_i[28]_pad ,
		_w9080_
	);
	LUT2 #(
		.INIT('h8)
	) name7331 (
		rst_i_pad,
		\u4_u2_iena_reg[4]/P0001 ,
		_w9081_
	);
	LUT4 #(
		.INIT('h5f08)
	) name7332 (
		_w2267_,
		_w9069_,
		_w9080_,
		_w9081_,
		_w9082_
	);
	LUT3 #(
		.INIT('h02)
	) name7333 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_data_i[29]_pad ,
		_w9083_
	);
	LUT2 #(
		.INIT('h8)
	) name7334 (
		rst_i_pad,
		\u4_u2_iena_reg[5]/P0001 ,
		_w9084_
	);
	LUT4 #(
		.INIT('h5f08)
	) name7335 (
		_w2267_,
		_w9069_,
		_w9083_,
		_w9084_,
		_w9085_
	);
	LUT3 #(
		.INIT('h02)
	) name7336 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_data_i[16]_pad ,
		_w9086_
	);
	LUT2 #(
		.INIT('h8)
	) name7337 (
		rst_i_pad,
		\u4_u2_ienb_reg[0]/P0001 ,
		_w9087_
	);
	LUT4 #(
		.INIT('h5f08)
	) name7338 (
		_w2267_,
		_w9069_,
		_w9086_,
		_w9087_,
		_w9088_
	);
	LUT3 #(
		.INIT('h02)
	) name7339 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_data_i[17]_pad ,
		_w9089_
	);
	LUT2 #(
		.INIT('h8)
	) name7340 (
		rst_i_pad,
		\u4_u2_ienb_reg[1]/P0001 ,
		_w9090_
	);
	LUT4 #(
		.INIT('h5f08)
	) name7341 (
		_w2267_,
		_w9069_,
		_w9089_,
		_w9090_,
		_w9091_
	);
	LUT3 #(
		.INIT('h02)
	) name7342 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_data_i[18]_pad ,
		_w9092_
	);
	LUT2 #(
		.INIT('h8)
	) name7343 (
		rst_i_pad,
		\u4_u2_ienb_reg[2]/P0001 ,
		_w9093_
	);
	LUT4 #(
		.INIT('h5f08)
	) name7344 (
		_w2267_,
		_w9069_,
		_w9092_,
		_w9093_,
		_w9094_
	);
	LUT3 #(
		.INIT('h02)
	) name7345 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_data_i[19]_pad ,
		_w9095_
	);
	LUT2 #(
		.INIT('h8)
	) name7346 (
		rst_i_pad,
		\u4_u2_ienb_reg[3]/P0001 ,
		_w9096_
	);
	LUT4 #(
		.INIT('h5f08)
	) name7347 (
		_w2267_,
		_w9069_,
		_w9095_,
		_w9096_,
		_w9097_
	);
	LUT3 #(
		.INIT('h02)
	) name7348 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_data_i[20]_pad ,
		_w9098_
	);
	LUT2 #(
		.INIT('h8)
	) name7349 (
		rst_i_pad,
		\u4_u2_ienb_reg[4]/P0001 ,
		_w9099_
	);
	LUT4 #(
		.INIT('h5f08)
	) name7350 (
		_w2267_,
		_w9069_,
		_w9098_,
		_w9099_,
		_w9100_
	);
	LUT3 #(
		.INIT('h02)
	) name7351 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_data_i[21]_pad ,
		_w9101_
	);
	LUT2 #(
		.INIT('h8)
	) name7352 (
		rst_i_pad,
		\u4_u2_ienb_reg[5]/P0001 ,
		_w9102_
	);
	LUT4 #(
		.INIT('h5f08)
	) name7353 (
		_w2267_,
		_w9069_,
		_w9101_,
		_w9102_,
		_w9103_
	);
	LUT3 #(
		.INIT('h20)
	) name7354 (
		rst_i_pad,
		\u4_u2_int_re_reg/P0001 ,
		\u4_u2_int_stat_reg[1]/P0001 ,
		_w9104_
	);
	LUT3 #(
		.INIT('hd0)
	) name7355 (
		\u0_rx_active_reg/P0001 ,
		\u0_rx_err_reg/P0001 ,
		\u4_u2_ep_match_r_reg/P0001 ,
		_w9105_
	);
	LUT3 #(
		.INIT('h80)
	) name7356 (
		_w3671_,
		_w3890_,
		_w9105_,
		_w9106_
	);
	LUT3 #(
		.INIT('hdc)
	) name7357 (
		_w3682_,
		_w9104_,
		_w9106_,
		_w9107_
	);
	LUT3 #(
		.INIT('h01)
	) name7358 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_data_i[13]_pad ,
		_w9108_
	);
	LUT2 #(
		.INIT('h8)
	) name7359 (
		rst_i_pad,
		\u4_u2_ots_stop_reg/P0001 ,
		_w9109_
	);
	LUT3 #(
		.INIT('h02)
	) name7360 (
		rst_i_pad,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w9110_
	);
	LUT4 #(
		.INIT('h7270)
	) name7361 (
		_w2267_,
		_w9108_,
		_w9109_,
		_w9110_,
		_w9111_
	);
	LUT3 #(
		.INIT('h2a)
	) name7362 (
		\u4_u3_buf0_orig_reg[9]/P0001 ,
		_w2231_,
		_w2232_,
		_w9112_
	);
	LUT2 #(
		.INIT('hd)
	) name7363 (
		_w7388_,
		_w9112_,
		_w9113_
	);
	LUT3 #(
		.INIT('h2a)
	) name7364 (
		\u4_u3_buf0_orig_reg[7]/P0001 ,
		_w2231_,
		_w2232_,
		_w9114_
	);
	LUT2 #(
		.INIT('hd)
	) name7365 (
		_w2519_,
		_w9114_,
		_w9115_
	);
	LUT3 #(
		.INIT('h2a)
	) name7366 (
		\u4_u3_buf0_orig_reg[0]/P0001 ,
		_w2231_,
		_w2232_,
		_w9116_
	);
	LUT2 #(
		.INIT('hd)
	) name7367 (
		_w7256_,
		_w9116_,
		_w9117_
	);
	LUT3 #(
		.INIT('h2a)
	) name7368 (
		\u4_u3_buf0_orig_reg[10]/P0001 ,
		_w2231_,
		_w2232_,
		_w9118_
	);
	LUT2 #(
		.INIT('hd)
	) name7369 (
		_w2275_,
		_w9118_,
		_w9119_
	);
	LUT3 #(
		.INIT('h2a)
	) name7370 (
		\u4_u3_buf0_orig_reg[11]/P0001 ,
		_w2231_,
		_w2232_,
		_w9120_
	);
	LUT2 #(
		.INIT('hd)
	) name7371 (
		_w2390_,
		_w9120_,
		_w9121_
	);
	LUT3 #(
		.INIT('h2a)
	) name7372 (
		\u4_u3_buf0_orig_reg[12]/P0001 ,
		_w2231_,
		_w2232_,
		_w9122_
	);
	LUT2 #(
		.INIT('hd)
	) name7373 (
		_w7262_,
		_w9122_,
		_w9123_
	);
	LUT3 #(
		.INIT('h2a)
	) name7374 (
		\u4_u3_buf0_orig_reg[14]/P0001 ,
		_w2231_,
		_w2232_,
		_w9124_
	);
	LUT2 #(
		.INIT('hd)
	) name7375 (
		_w2234_,
		_w9124_,
		_w9125_
	);
	LUT3 #(
		.INIT('h2a)
	) name7376 (
		\u4_u3_buf0_orig_reg[15]/P0001 ,
		_w2231_,
		_w2232_,
		_w9126_
	);
	LUT2 #(
		.INIT('hd)
	) name7377 (
		_w2396_,
		_w9126_,
		_w9127_
	);
	LUT3 #(
		.INIT('h2a)
	) name7378 (
		\u4_u3_buf0_orig_reg[16]/P0001 ,
		_w2231_,
		_w2232_,
		_w9128_
	);
	LUT2 #(
		.INIT('hd)
	) name7379 (
		_w7268_,
		_w9128_,
		_w9129_
	);
	LUT3 #(
		.INIT('h2a)
	) name7380 (
		\u4_u3_buf0_orig_reg[17]/P0001 ,
		_w2231_,
		_w2232_,
		_w9130_
	);
	LUT2 #(
		.INIT('hd)
	) name7381 (
		_w7274_,
		_w9130_,
		_w9131_
	);
	LUT3 #(
		.INIT('h2a)
	) name7382 (
		\u4_u3_buf0_orig_reg[18]/P0001 ,
		_w2231_,
		_w2232_,
		_w9132_
	);
	LUT2 #(
		.INIT('hd)
	) name7383 (
		_w7280_,
		_w9132_,
		_w9133_
	);
	LUT3 #(
		.INIT('h2a)
	) name7384 (
		\u4_u3_buf0_orig_reg[19]/P0001 ,
		_w2231_,
		_w2232_,
		_w9134_
	);
	LUT2 #(
		.INIT('hd)
	) name7385 (
		_w7286_,
		_w9134_,
		_w9135_
	);
	LUT3 #(
		.INIT('h2a)
	) name7386 (
		\u4_u3_buf0_orig_reg[1]/P0001 ,
		_w2231_,
		_w2232_,
		_w9136_
	);
	LUT2 #(
		.INIT('hd)
	) name7387 (
		_w7292_,
		_w9136_,
		_w9137_
	);
	LUT3 #(
		.INIT('h2a)
	) name7388 (
		\u4_u3_buf0_orig_reg[20]/P0001 ,
		_w2231_,
		_w2232_,
		_w9138_
	);
	LUT2 #(
		.INIT('hd)
	) name7389 (
		_w7298_,
		_w9138_,
		_w9139_
	);
	LUT3 #(
		.INIT('h2a)
	) name7390 (
		\u4_u3_buf0_orig_reg[22]/P0001 ,
		_w2231_,
		_w2232_,
		_w9140_
	);
	LUT2 #(
		.INIT('hd)
	) name7391 (
		_w7310_,
		_w9140_,
		_w9141_
	);
	LUT3 #(
		.INIT('h2a)
	) name7392 (
		\u4_u3_buf0_orig_reg[23]/P0001 ,
		_w2231_,
		_w2232_,
		_w9142_
	);
	LUT2 #(
		.INIT('hd)
	) name7393 (
		_w7316_,
		_w9142_,
		_w9143_
	);
	LUT3 #(
		.INIT('h2a)
	) name7394 (
		\u4_u3_buf0_orig_reg[24]/P0001 ,
		_w2231_,
		_w2232_,
		_w9144_
	);
	LUT2 #(
		.INIT('hd)
	) name7395 (
		_w7322_,
		_w9144_,
		_w9145_
	);
	LUT3 #(
		.INIT('h2a)
	) name7396 (
		\u4_u3_buf0_orig_reg[25]/P0001 ,
		_w2231_,
		_w2232_,
		_w9146_
	);
	LUT2 #(
		.INIT('hd)
	) name7397 (
		_w7328_,
		_w9146_,
		_w9147_
	);
	LUT3 #(
		.INIT('h2a)
	) name7398 (
		\u4_u3_buf0_orig_reg[26]/P0001 ,
		_w2231_,
		_w2232_,
		_w9148_
	);
	LUT2 #(
		.INIT('hd)
	) name7399 (
		_w7334_,
		_w9148_,
		_w9149_
	);
	LUT3 #(
		.INIT('h2a)
	) name7400 (
		\u4_u3_buf0_orig_reg[27]/P0001 ,
		_w2231_,
		_w2232_,
		_w9150_
	);
	LUT2 #(
		.INIT('hd)
	) name7401 (
		_w7340_,
		_w9150_,
		_w9151_
	);
	LUT3 #(
		.INIT('h2a)
	) name7402 (
		\u4_u3_buf0_orig_reg[28]/P0001 ,
		_w2231_,
		_w2232_,
		_w9152_
	);
	LUT2 #(
		.INIT('hd)
	) name7403 (
		_w7346_,
		_w9152_,
		_w9153_
	);
	LUT3 #(
		.INIT('h2a)
	) name7404 (
		\u4_u3_buf0_orig_reg[29]/NET0131 ,
		_w2231_,
		_w2232_,
		_w9154_
	);
	LUT2 #(
		.INIT('hd)
	) name7405 (
		_w7352_,
		_w9154_,
		_w9155_
	);
	LUT3 #(
		.INIT('h2a)
	) name7406 (
		\u4_u3_buf0_orig_reg[2]/P0001 ,
		_w2231_,
		_w2232_,
		_w9156_
	);
	LUT2 #(
		.INIT('hd)
	) name7407 (
		_w7358_,
		_w9156_,
		_w9157_
	);
	LUT3 #(
		.INIT('h2a)
	) name7408 (
		\u4_u3_buf0_orig_reg[30]/NET0131 ,
		_w2231_,
		_w2232_,
		_w9158_
	);
	LUT2 #(
		.INIT('hd)
	) name7409 (
		_w7364_,
		_w9158_,
		_w9159_
	);
	LUT3 #(
		.INIT('h2a)
	) name7410 (
		\u4_u3_buf0_orig_reg[31]/P0001 ,
		_w2231_,
		_w2232_,
		_w9160_
	);
	LUT2 #(
		.INIT('hd)
	) name7411 (
		_w7370_,
		_w9160_,
		_w9161_
	);
	LUT3 #(
		.INIT('h2a)
	) name7412 (
		\u4_u3_buf0_orig_reg[3]/P0001 ,
		_w2231_,
		_w2232_,
		_w9162_
	);
	LUT2 #(
		.INIT('hd)
	) name7413 (
		_w7376_,
		_w9162_,
		_w9163_
	);
	LUT3 #(
		.INIT('h2a)
	) name7414 (
		\u4_u3_buf0_orig_reg[4]/P0001 ,
		_w2231_,
		_w2232_,
		_w9164_
	);
	LUT2 #(
		.INIT('hd)
	) name7415 (
		_w2507_,
		_w9164_,
		_w9165_
	);
	LUT3 #(
		.INIT('h2a)
	) name7416 (
		\u4_u3_buf0_orig_reg[5]/P0001 ,
		_w2231_,
		_w2232_,
		_w9166_
	);
	LUT2 #(
		.INIT('hd)
	) name7417 (
		_w2513_,
		_w9166_,
		_w9167_
	);
	LUT3 #(
		.INIT('h2a)
	) name7418 (
		\u4_u3_buf0_orig_reg[6]/P0001 ,
		_w2231_,
		_w2232_,
		_w9168_
	);
	LUT2 #(
		.INIT('hd)
	) name7419 (
		_w2409_,
		_w9168_,
		_w9169_
	);
	LUT3 #(
		.INIT('h01)
	) name7420 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_data_i[15]_pad ,
		_w9170_
	);
	LUT2 #(
		.INIT('h8)
	) name7421 (
		rst_i_pad,
		\u4_u2_csr1_reg[0]/P0001 ,
		_w9171_
	);
	LUT4 #(
		.INIT('h5f08)
	) name7422 (
		_w2267_,
		_w9110_,
		_w9170_,
		_w9171_,
		_w9172_
	);
	LUT3 #(
		.INIT('h01)
	) name7423 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_data_i[0]_pad ,
		_w9173_
	);
	LUT2 #(
		.INIT('h8)
	) name7424 (
		rst_i_pad,
		\u4_u3_csr0_reg[0]/P0001 ,
		_w9174_
	);
	LUT4 #(
		.INIT('h5f08)
	) name7425 (
		_w2231_,
		_w9110_,
		_w9173_,
		_w9174_,
		_w9175_
	);
	LUT3 #(
		.INIT('h01)
	) name7426 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_data_i[10]_pad ,
		_w9176_
	);
	LUT2 #(
		.INIT('h8)
	) name7427 (
		rst_i_pad,
		\u4_u3_csr0_reg[10]/P0001 ,
		_w9177_
	);
	LUT4 #(
		.INIT('h5f08)
	) name7428 (
		_w2231_,
		_w9110_,
		_w9176_,
		_w9177_,
		_w9178_
	);
	LUT3 #(
		.INIT('h01)
	) name7429 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_data_i[11]_pad ,
		_w9179_
	);
	LUT2 #(
		.INIT('h8)
	) name7430 (
		rst_i_pad,
		\u4_u3_csr0_reg[11]/P0001 ,
		_w9180_
	);
	LUT4 #(
		.INIT('h5f08)
	) name7431 (
		_w2231_,
		_w9110_,
		_w9179_,
		_w9180_,
		_w9181_
	);
	LUT3 #(
		.INIT('h01)
	) name7432 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_data_i[12]_pad ,
		_w9182_
	);
	LUT2 #(
		.INIT('h8)
	) name7433 (
		rst_i_pad,
		\u4_u3_csr0_reg[12]/P0001 ,
		_w9183_
	);
	LUT4 #(
		.INIT('h5f08)
	) name7434 (
		_w2231_,
		_w9110_,
		_w9182_,
		_w9183_,
		_w9184_
	);
	LUT3 #(
		.INIT('h01)
	) name7435 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_data_i[1]_pad ,
		_w9185_
	);
	LUT2 #(
		.INIT('h8)
	) name7436 (
		rst_i_pad,
		\u4_u3_csr0_reg[1]/P0001 ,
		_w9186_
	);
	LUT4 #(
		.INIT('h5f08)
	) name7437 (
		_w2231_,
		_w9110_,
		_w9185_,
		_w9186_,
		_w9187_
	);
	LUT3 #(
		.INIT('h01)
	) name7438 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_data_i[2]_pad ,
		_w9188_
	);
	LUT2 #(
		.INIT('h8)
	) name7439 (
		rst_i_pad,
		\u4_u3_csr0_reg[2]/P0001 ,
		_w9189_
	);
	LUT4 #(
		.INIT('h5f08)
	) name7440 (
		_w2231_,
		_w9110_,
		_w9188_,
		_w9189_,
		_w9190_
	);
	LUT3 #(
		.INIT('h01)
	) name7441 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_data_i[3]_pad ,
		_w9191_
	);
	LUT2 #(
		.INIT('h8)
	) name7442 (
		rst_i_pad,
		\u4_u3_csr0_reg[3]/NET0131 ,
		_w9192_
	);
	LUT4 #(
		.INIT('h5f08)
	) name7443 (
		_w2231_,
		_w9110_,
		_w9191_,
		_w9192_,
		_w9193_
	);
	LUT3 #(
		.INIT('h01)
	) name7444 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_data_i[4]_pad ,
		_w9194_
	);
	LUT2 #(
		.INIT('h8)
	) name7445 (
		rst_i_pad,
		\u4_u3_csr0_reg[4]/P0001 ,
		_w9195_
	);
	LUT4 #(
		.INIT('h5f08)
	) name7446 (
		_w2231_,
		_w9110_,
		_w9194_,
		_w9195_,
		_w9196_
	);
	LUT3 #(
		.INIT('h01)
	) name7447 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_data_i[5]_pad ,
		_w9197_
	);
	LUT2 #(
		.INIT('h8)
	) name7448 (
		rst_i_pad,
		\u4_u3_csr0_reg[5]/P0001 ,
		_w9198_
	);
	LUT4 #(
		.INIT('h5f08)
	) name7449 (
		_w2231_,
		_w9110_,
		_w9197_,
		_w9198_,
		_w9199_
	);
	LUT3 #(
		.INIT('h01)
	) name7450 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_data_i[6]_pad ,
		_w9200_
	);
	LUT2 #(
		.INIT('h8)
	) name7451 (
		rst_i_pad,
		\u4_u3_csr0_reg[6]/P0001 ,
		_w9201_
	);
	LUT4 #(
		.INIT('h5f08)
	) name7452 (
		_w2231_,
		_w9110_,
		_w9200_,
		_w9201_,
		_w9202_
	);
	LUT3 #(
		.INIT('h01)
	) name7453 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_data_i[7]_pad ,
		_w9203_
	);
	LUT2 #(
		.INIT('h8)
	) name7454 (
		rst_i_pad,
		\u4_u3_csr0_reg[7]/P0001 ,
		_w9204_
	);
	LUT4 #(
		.INIT('h5f08)
	) name7455 (
		_w2231_,
		_w9110_,
		_w9203_,
		_w9204_,
		_w9205_
	);
	LUT3 #(
		.INIT('h01)
	) name7456 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_data_i[8]_pad ,
		_w9206_
	);
	LUT2 #(
		.INIT('h8)
	) name7457 (
		rst_i_pad,
		\u4_u3_csr0_reg[8]/P0001 ,
		_w9207_
	);
	LUT4 #(
		.INIT('h5f08)
	) name7458 (
		_w2231_,
		_w9110_,
		_w9206_,
		_w9207_,
		_w9208_
	);
	LUT3 #(
		.INIT('h01)
	) name7459 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_data_i[9]_pad ,
		_w9209_
	);
	LUT2 #(
		.INIT('h8)
	) name7460 (
		rst_i_pad,
		\u4_u3_csr0_reg[9]/P0001 ,
		_w9210_
	);
	LUT4 #(
		.INIT('h5f08)
	) name7461 (
		_w2231_,
		_w9110_,
		_w9209_,
		_w9210_,
		_w9211_
	);
	LUT2 #(
		.INIT('h8)
	) name7462 (
		rst_i_pad,
		\u4_u3_csr1_reg[0]/P0001 ,
		_w9212_
	);
	LUT4 #(
		.INIT('h5f08)
	) name7463 (
		_w2231_,
		_w9110_,
		_w9170_,
		_w9212_,
		_w9213_
	);
	LUT3 #(
		.INIT('h01)
	) name7464 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_data_i[25]_pad ,
		_w9214_
	);
	LUT2 #(
		.INIT('h8)
	) name7465 (
		rst_i_pad,
		\u4_u3_csr1_reg[10]/P0001 ,
		_w9215_
	);
	LUT4 #(
		.INIT('h5f08)
	) name7466 (
		_w2231_,
		_w9110_,
		_w9214_,
		_w9215_,
		_w9216_
	);
	LUT3 #(
		.INIT('h01)
	) name7467 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_data_i[26]_pad ,
		_w9217_
	);
	LUT2 #(
		.INIT('h8)
	) name7468 (
		rst_i_pad,
		\u4_u3_csr1_reg[11]/P0001 ,
		_w9218_
	);
	LUT4 #(
		.INIT('h5f08)
	) name7469 (
		_w2231_,
		_w9110_,
		_w9217_,
		_w9218_,
		_w9219_
	);
	LUT3 #(
		.INIT('h01)
	) name7470 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_data_i[27]_pad ,
		_w9220_
	);
	LUT2 #(
		.INIT('h8)
	) name7471 (
		rst_i_pad,
		\u4_u3_csr1_reg[12]/P0001 ,
		_w9221_
	);
	LUT4 #(
		.INIT('h5f08)
	) name7472 (
		_w2231_,
		_w9110_,
		_w9220_,
		_w9221_,
		_w9222_
	);
	LUT3 #(
		.INIT('h01)
	) name7473 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_data_i[16]_pad ,
		_w9223_
	);
	LUT2 #(
		.INIT('h8)
	) name7474 (
		rst_i_pad,
		\u4_u3_csr1_reg[1]/P0001 ,
		_w9224_
	);
	LUT4 #(
		.INIT('h5f08)
	) name7475 (
		_w2231_,
		_w9110_,
		_w9223_,
		_w9224_,
		_w9225_
	);
	LUT3 #(
		.INIT('h01)
	) name7476 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_data_i[17]_pad ,
		_w9226_
	);
	LUT2 #(
		.INIT('h8)
	) name7477 (
		rst_i_pad,
		\u4_u3_csr1_reg[2]/P0001 ,
		_w9227_
	);
	LUT4 #(
		.INIT('h5f08)
	) name7478 (
		_w2231_,
		_w9110_,
		_w9226_,
		_w9227_,
		_w9228_
	);
	LUT3 #(
		.INIT('h01)
	) name7479 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_data_i[18]_pad ,
		_w9229_
	);
	LUT2 #(
		.INIT('h8)
	) name7480 (
		rst_i_pad,
		\u4_u3_csr1_reg[3]/P0001 ,
		_w9230_
	);
	LUT4 #(
		.INIT('h5f08)
	) name7481 (
		_w2231_,
		_w9110_,
		_w9229_,
		_w9230_,
		_w9231_
	);
	LUT3 #(
		.INIT('h01)
	) name7482 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_data_i[19]_pad ,
		_w9232_
	);
	LUT2 #(
		.INIT('h8)
	) name7483 (
		rst_i_pad,
		\u4_u3_csr1_reg[4]/P0001 ,
		_w9233_
	);
	LUT4 #(
		.INIT('h5f08)
	) name7484 (
		_w2231_,
		_w9110_,
		_w9232_,
		_w9233_,
		_w9234_
	);
	LUT3 #(
		.INIT('h01)
	) name7485 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_data_i[20]_pad ,
		_w9235_
	);
	LUT2 #(
		.INIT('h8)
	) name7486 (
		rst_i_pad,
		\u4_u3_csr1_reg[5]/P0001 ,
		_w9236_
	);
	LUT4 #(
		.INIT('h5f08)
	) name7487 (
		_w2231_,
		_w9110_,
		_w9235_,
		_w9236_,
		_w9237_
	);
	LUT3 #(
		.INIT('h01)
	) name7488 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_data_i[21]_pad ,
		_w9238_
	);
	LUT2 #(
		.INIT('h8)
	) name7489 (
		rst_i_pad,
		\u4_u3_csr1_reg[6]/P0001 ,
		_w9239_
	);
	LUT4 #(
		.INIT('h5f08)
	) name7490 (
		_w2231_,
		_w9110_,
		_w9238_,
		_w9239_,
		_w9240_
	);
	LUT3 #(
		.INIT('h01)
	) name7491 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_data_i[24]_pad ,
		_w9241_
	);
	LUT2 #(
		.INIT('h8)
	) name7492 (
		rst_i_pad,
		\u4_u3_csr1_reg[9]/P0001 ,
		_w9242_
	);
	LUT4 #(
		.INIT('h5f08)
	) name7493 (
		_w2231_,
		_w9110_,
		_w9241_,
		_w9242_,
		_w9243_
	);
	LUT3 #(
		.INIT('h2a)
	) name7494 (
		\u4_u3_buf0_orig_reg[13]/P0001 ,
		_w2231_,
		_w2232_,
		_w9244_
	);
	LUT2 #(
		.INIT('hd)
	) name7495 (
		_w2315_,
		_w9244_,
		_w9245_
	);
	LUT3 #(
		.INIT('h02)
	) name7496 (
		\u4_u1_csr1_reg[7]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w9246_
	);
	LUT4 #(
		.INIT('h35ff)
	) name7497 (
		\u4_u1_buf0_reg[22]/P0001 ,
		\u4_u1_buf1_reg[22]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w9247_
	);
	LUT4 #(
		.INIT('h8088)
	) name7498 (
		_w2227_,
		_w2241_,
		_w9246_,
		_w9247_,
		_w9248_
	);
	LUT3 #(
		.INIT('h02)
	) name7499 (
		\u4_u3_csr1_reg[7]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w9249_
	);
	LUT4 #(
		.INIT('h35ff)
	) name7500 (
		\u4_u3_buf0_reg[22]/P0001 ,
		\u4_u3_buf1_reg[22]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w9250_
	);
	LUT4 #(
		.INIT('h8088)
	) name7501 (
		_w2227_,
		_w2228_,
		_w9249_,
		_w9250_,
		_w9251_
	);
	LUT3 #(
		.INIT('h02)
	) name7502 (
		\u4_u2_csr1_reg[7]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w9252_
	);
	LUT4 #(
		.INIT('h35ff)
	) name7503 (
		\u4_u2_buf0_reg[22]/P0001 ,
		\u4_u2_buf1_reg[22]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w9253_
	);
	LUT4 #(
		.INIT('h8088)
	) name7504 (
		_w2228_,
		_w2240_,
		_w9252_,
		_w9253_,
		_w9254_
	);
	LUT3 #(
		.INIT('h01)
	) name7505 (
		_w9248_,
		_w9251_,
		_w9254_,
		_w9255_
	);
	LUT4 #(
		.INIT('h0200)
	) name7506 (
		\u1_frame_no_r_reg[6]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w9256_
	);
	LUT4 #(
		.INIT('h0020)
	) name7507 (
		\u4_intb_msk_reg[6]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w9257_
	);
	LUT4 #(
		.INIT('h0080)
	) name7508 (
		\u4_int_srcb_reg[2]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w9258_
	);
	LUT4 #(
		.INIT('haaa8)
	) name7509 (
		_w5861_,
		_w9256_,
		_w9257_,
		_w9258_,
		_w9259_
	);
	LUT3 #(
		.INIT('h02)
	) name7510 (
		\u4_u0_csr1_reg[7]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w9260_
	);
	LUT4 #(
		.INIT('h35ff)
	) name7511 (
		\u4_u0_buf0_reg[22]/P0001 ,
		\u4_u0_buf1_reg[22]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w9261_
	);
	LUT4 #(
		.INIT('h8088)
	) name7512 (
		_w2240_,
		_w2241_,
		_w9260_,
		_w9261_,
		_w9262_
	);
	LUT2 #(
		.INIT('h1)
	) name7513 (
		_w9259_,
		_w9262_,
		_w9263_
	);
	LUT2 #(
		.INIT('h7)
	) name7514 (
		_w9255_,
		_w9263_,
		_w9264_
	);
	LUT3 #(
		.INIT('h2a)
	) name7515 (
		\u4_u3_buf0_orig_reg[8]/P0001 ,
		_w2231_,
		_w2232_,
		_w9265_
	);
	LUT2 #(
		.INIT('hd)
	) name7516 (
		_w7382_,
		_w9265_,
		_w9266_
	);
	LUT2 #(
		.INIT('h8)
	) name7517 (
		rst_i_pad,
		\u4_u3_iena_reg[0]/P0001 ,
		_w9267_
	);
	LUT4 #(
		.INIT('h7720)
	) name7518 (
		_w2231_,
		_w9067_,
		_w9069_,
		_w9267_,
		_w9268_
	);
	LUT2 #(
		.INIT('h8)
	) name7519 (
		rst_i_pad,
		\u4_u3_iena_reg[1]/P0001 ,
		_w9269_
	);
	LUT4 #(
		.INIT('h5f08)
	) name7520 (
		_w2231_,
		_w9069_,
		_w9071_,
		_w9269_,
		_w9270_
	);
	LUT2 #(
		.INIT('h8)
	) name7521 (
		rst_i_pad,
		\u4_u3_iena_reg[2]/P0001 ,
		_w9271_
	);
	LUT4 #(
		.INIT('h5f08)
	) name7522 (
		_w2231_,
		_w9069_,
		_w9074_,
		_w9271_,
		_w9272_
	);
	LUT2 #(
		.INIT('h8)
	) name7523 (
		rst_i_pad,
		\u4_u3_iena_reg[3]/P0001 ,
		_w9273_
	);
	LUT4 #(
		.INIT('h5f08)
	) name7524 (
		_w2231_,
		_w9069_,
		_w9077_,
		_w9273_,
		_w9274_
	);
	LUT2 #(
		.INIT('h8)
	) name7525 (
		rst_i_pad,
		\u4_u3_iena_reg[4]/P0001 ,
		_w9275_
	);
	LUT4 #(
		.INIT('h5f08)
	) name7526 (
		_w2231_,
		_w9069_,
		_w9080_,
		_w9275_,
		_w9276_
	);
	LUT2 #(
		.INIT('h8)
	) name7527 (
		rst_i_pad,
		\u4_u3_iena_reg[5]/P0001 ,
		_w9277_
	);
	LUT4 #(
		.INIT('h5f08)
	) name7528 (
		_w2231_,
		_w9069_,
		_w9083_,
		_w9277_,
		_w9278_
	);
	LUT2 #(
		.INIT('h8)
	) name7529 (
		rst_i_pad,
		\u4_u3_ienb_reg[0]/P0001 ,
		_w9279_
	);
	LUT4 #(
		.INIT('h5f08)
	) name7530 (
		_w2231_,
		_w9069_,
		_w9086_,
		_w9279_,
		_w9280_
	);
	LUT2 #(
		.INIT('h8)
	) name7531 (
		rst_i_pad,
		\u4_u3_ienb_reg[2]/P0001 ,
		_w9281_
	);
	LUT4 #(
		.INIT('h5f08)
	) name7532 (
		_w2231_,
		_w9069_,
		_w9092_,
		_w9281_,
		_w9282_
	);
	LUT2 #(
		.INIT('h8)
	) name7533 (
		rst_i_pad,
		\u4_u3_ienb_reg[3]/P0001 ,
		_w9283_
	);
	LUT4 #(
		.INIT('h5f08)
	) name7534 (
		_w2231_,
		_w9069_,
		_w9095_,
		_w9283_,
		_w9284_
	);
	LUT2 #(
		.INIT('h8)
	) name7535 (
		rst_i_pad,
		\u4_u3_ienb_reg[1]/P0001 ,
		_w9285_
	);
	LUT4 #(
		.INIT('h5f08)
	) name7536 (
		_w2231_,
		_w9069_,
		_w9089_,
		_w9285_,
		_w9286_
	);
	LUT2 #(
		.INIT('h8)
	) name7537 (
		rst_i_pad,
		\u4_u3_ienb_reg[4]/P0001 ,
		_w9287_
	);
	LUT4 #(
		.INIT('h5f08)
	) name7538 (
		_w2231_,
		_w9069_,
		_w9098_,
		_w9287_,
		_w9288_
	);
	LUT2 #(
		.INIT('h8)
	) name7539 (
		rst_i_pad,
		\u4_u3_ienb_reg[5]/P0001 ,
		_w9289_
	);
	LUT4 #(
		.INIT('h5f08)
	) name7540 (
		_w2231_,
		_w9069_,
		_w9101_,
		_w9289_,
		_w9290_
	);
	LUT3 #(
		.INIT('h20)
	) name7541 (
		rst_i_pad,
		\u4_u3_int_re_reg/P0001 ,
		\u4_u3_int_stat_reg[1]/P0001 ,
		_w9291_
	);
	LUT3 #(
		.INIT('hd0)
	) name7542 (
		\u0_rx_active_reg/P0001 ,
		\u0_rx_err_reg/P0001 ,
		\u4_u3_ep_match_r_reg/P0001 ,
		_w9292_
	);
	LUT3 #(
		.INIT('h80)
	) name7543 (
		_w3671_,
		_w3893_,
		_w9292_,
		_w9293_
	);
	LUT3 #(
		.INIT('hdc)
	) name7544 (
		_w3682_,
		_w9291_,
		_w9293_,
		_w9294_
	);
	LUT2 #(
		.INIT('h8)
	) name7545 (
		rst_i_pad,
		\u4_u3_ots_stop_reg/P0001 ,
		_w9295_
	);
	LUT4 #(
		.INIT('h7720)
	) name7546 (
		_w2231_,
		_w9108_,
		_w9110_,
		_w9295_,
		_w9296_
	);
	LUT3 #(
		.INIT('h02)
	) name7547 (
		\u4_u1_csr0_reg[7]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w9297_
	);
	LUT4 #(
		.INIT('h35ff)
	) name7548 (
		\u4_u1_buf0_reg[7]/P0001 ,
		\u4_u1_buf1_reg[7]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w9298_
	);
	LUT4 #(
		.INIT('h8088)
	) name7549 (
		_w2227_,
		_w2241_,
		_w9297_,
		_w9298_,
		_w9299_
	);
	LUT3 #(
		.INIT('h02)
	) name7550 (
		\u4_u3_csr0_reg[7]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w9300_
	);
	LUT4 #(
		.INIT('h35ff)
	) name7551 (
		\u4_u3_buf0_reg[7]/P0001 ,
		\u4_u3_buf1_reg[7]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w9301_
	);
	LUT4 #(
		.INIT('h8088)
	) name7552 (
		_w2227_,
		_w2228_,
		_w9300_,
		_w9301_,
		_w9302_
	);
	LUT3 #(
		.INIT('h02)
	) name7553 (
		\u4_u2_csr0_reg[7]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w9303_
	);
	LUT4 #(
		.INIT('h35ff)
	) name7554 (
		\u4_u2_buf0_reg[7]/P0001 ,
		\u4_u2_buf1_reg[7]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w9304_
	);
	LUT4 #(
		.INIT('h8088)
	) name7555 (
		_w2228_,
		_w2240_,
		_w9303_,
		_w9304_,
		_w9305_
	);
	LUT3 #(
		.INIT('h01)
	) name7556 (
		_w9299_,
		_w9302_,
		_w9305_,
		_w9306_
	);
	LUT4 #(
		.INIT('h0800)
	) name7557 (
		\u4_utmi_vend_stat_r_reg[7]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w9307_
	);
	LUT4 #(
		.INIT('h0020)
	) name7558 (
		\u4_inta_msk_reg[7]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w9308_
	);
	LUT4 #(
		.INIT('h0200)
	) name7559 (
		\u1_sof_time_reg[7]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w9309_
	);
	LUT4 #(
		.INIT('haaa8)
	) name7560 (
		_w5861_,
		_w9307_,
		_w9308_,
		_w9309_,
		_w9310_
	);
	LUT3 #(
		.INIT('h02)
	) name7561 (
		\u4_u0_csr0_reg[7]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w9311_
	);
	LUT4 #(
		.INIT('h35ff)
	) name7562 (
		\u4_u0_buf0_reg[7]/P0001 ,
		\u4_u0_buf1_reg[7]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w9312_
	);
	LUT4 #(
		.INIT('h8088)
	) name7563 (
		_w2240_,
		_w2241_,
		_w9311_,
		_w9312_,
		_w9313_
	);
	LUT2 #(
		.INIT('h1)
	) name7564 (
		_w9310_,
		_w9313_,
		_w9314_
	);
	LUT2 #(
		.INIT('h7)
	) name7565 (
		_w9306_,
		_w9314_,
		_w9315_
	);
	LUT3 #(
		.INIT('h2a)
	) name7566 (
		\u4_u0_buf0_orig_reg[0]/P0001 ,
		_w2232_,
		_w2243_,
		_w9316_
	);
	LUT2 #(
		.INIT('hd)
	) name7567 (
		_w7401_,
		_w9316_,
		_w9317_
	);
	LUT3 #(
		.INIT('h2a)
	) name7568 (
		\u4_u0_buf0_orig_reg[10]/P0001 ,
		_w2232_,
		_w2243_,
		_w9318_
	);
	LUT2 #(
		.INIT('hd)
	) name7569 (
		_w2280_,
		_w9318_,
		_w9319_
	);
	LUT3 #(
		.INIT('h2a)
	) name7570 (
		\u4_u0_buf0_orig_reg[11]/P0001 ,
		_w2232_,
		_w2243_,
		_w9320_
	);
	LUT2 #(
		.INIT('hd)
	) name7571 (
		_w2414_,
		_w9320_,
		_w9321_
	);
	LUT3 #(
		.INIT('h2a)
	) name7572 (
		\u4_u0_buf0_orig_reg[12]/P0001 ,
		_w2232_,
		_w2243_,
		_w9322_
	);
	LUT2 #(
		.INIT('hd)
	) name7573 (
		_w7406_,
		_w9322_,
		_w9323_
	);
	LUT3 #(
		.INIT('h2a)
	) name7574 (
		\u4_u0_buf0_orig_reg[13]/P0001 ,
		_w2232_,
		_w2243_,
		_w9324_
	);
	LUT2 #(
		.INIT('hd)
	) name7575 (
		_w2328_,
		_w9324_,
		_w9325_
	);
	LUT3 #(
		.INIT('h2a)
	) name7576 (
		\u4_u0_buf0_orig_reg[14]/P0001 ,
		_w2232_,
		_w2243_,
		_w9326_
	);
	LUT2 #(
		.INIT('hd)
	) name7577 (
		_w2244_,
		_w9326_,
		_w9327_
	);
	LUT3 #(
		.INIT('h2a)
	) name7578 (
		\u4_u0_buf0_orig_reg[15]/P0001 ,
		_w2232_,
		_w2243_,
		_w9328_
	);
	LUT2 #(
		.INIT('hd)
	) name7579 (
		_w2419_,
		_w9328_,
		_w9329_
	);
	LUT3 #(
		.INIT('h2a)
	) name7580 (
		\u4_u0_buf0_orig_reg[16]/P0001 ,
		_w2232_,
		_w2243_,
		_w9330_
	);
	LUT2 #(
		.INIT('hd)
	) name7581 (
		_w7411_,
		_w9330_,
		_w9331_
	);
	LUT3 #(
		.INIT('h2a)
	) name7582 (
		\u4_u0_buf0_orig_reg[17]/P0001 ,
		_w2232_,
		_w2243_,
		_w9332_
	);
	LUT2 #(
		.INIT('hd)
	) name7583 (
		_w7416_,
		_w9332_,
		_w9333_
	);
	LUT3 #(
		.INIT('h2a)
	) name7584 (
		\u4_u0_buf0_orig_reg[18]/P0001 ,
		_w2232_,
		_w2243_,
		_w9334_
	);
	LUT2 #(
		.INIT('hd)
	) name7585 (
		_w7421_,
		_w9334_,
		_w9335_
	);
	LUT3 #(
		.INIT('h2a)
	) name7586 (
		\u4_u0_buf0_orig_reg[19]/P0001 ,
		_w2232_,
		_w2243_,
		_w9336_
	);
	LUT2 #(
		.INIT('hd)
	) name7587 (
		_w7426_,
		_w9336_,
		_w9337_
	);
	LUT3 #(
		.INIT('h2a)
	) name7588 (
		\u4_u0_buf0_orig_reg[1]/P0001 ,
		_w2232_,
		_w2243_,
		_w9338_
	);
	LUT2 #(
		.INIT('hd)
	) name7589 (
		_w7431_,
		_w9338_,
		_w9339_
	);
	LUT3 #(
		.INIT('h2a)
	) name7590 (
		\u4_u0_buf0_orig_reg[20]/P0001 ,
		_w2232_,
		_w2243_,
		_w9340_
	);
	LUT2 #(
		.INIT('hd)
	) name7591 (
		_w7436_,
		_w9340_,
		_w9341_
	);
	LUT3 #(
		.INIT('h2a)
	) name7592 (
		\u4_u0_buf0_orig_reg[21]/P0001 ,
		_w2232_,
		_w2243_,
		_w9342_
	);
	LUT2 #(
		.INIT('hd)
	) name7593 (
		_w7441_,
		_w9342_,
		_w9343_
	);
	LUT3 #(
		.INIT('h2a)
	) name7594 (
		\u4_u0_buf0_orig_reg[22]/P0001 ,
		_w2232_,
		_w2243_,
		_w9344_
	);
	LUT2 #(
		.INIT('hd)
	) name7595 (
		_w7446_,
		_w9344_,
		_w9345_
	);
	LUT3 #(
		.INIT('h2a)
	) name7596 (
		\u4_u0_buf0_orig_reg[23]/P0001 ,
		_w2232_,
		_w2243_,
		_w9346_
	);
	LUT2 #(
		.INIT('hd)
	) name7597 (
		_w7451_,
		_w9346_,
		_w9347_
	);
	LUT3 #(
		.INIT('h2a)
	) name7598 (
		\u4_u0_buf0_orig_reg[24]/P0001 ,
		_w2232_,
		_w2243_,
		_w9348_
	);
	LUT2 #(
		.INIT('hd)
	) name7599 (
		_w7456_,
		_w9348_,
		_w9349_
	);
	LUT3 #(
		.INIT('h2a)
	) name7600 (
		\u4_u0_buf0_orig_reg[25]/P0001 ,
		_w2232_,
		_w2243_,
		_w9350_
	);
	LUT2 #(
		.INIT('hd)
	) name7601 (
		_w7461_,
		_w9350_,
		_w9351_
	);
	LUT3 #(
		.INIT('h2a)
	) name7602 (
		\u4_u0_buf0_orig_reg[26]/P0001 ,
		_w2232_,
		_w2243_,
		_w9352_
	);
	LUT2 #(
		.INIT('hd)
	) name7603 (
		_w7466_,
		_w9352_,
		_w9353_
	);
	LUT3 #(
		.INIT('h2a)
	) name7604 (
		\u4_u0_buf0_orig_reg[27]/P0001 ,
		_w2232_,
		_w2243_,
		_w9354_
	);
	LUT2 #(
		.INIT('hd)
	) name7605 (
		_w7471_,
		_w9354_,
		_w9355_
	);
	LUT3 #(
		.INIT('h2a)
	) name7606 (
		\u4_u0_buf0_orig_reg[28]/P0001 ,
		_w2232_,
		_w2243_,
		_w9356_
	);
	LUT2 #(
		.INIT('hd)
	) name7607 (
		_w7476_,
		_w9356_,
		_w9357_
	);
	LUT3 #(
		.INIT('h2a)
	) name7608 (
		\u4_u0_buf0_orig_reg[29]/NET0131 ,
		_w2232_,
		_w2243_,
		_w9358_
	);
	LUT2 #(
		.INIT('hd)
	) name7609 (
		_w7481_,
		_w9358_,
		_w9359_
	);
	LUT3 #(
		.INIT('h2a)
	) name7610 (
		\u4_u0_buf0_orig_reg[2]/P0001 ,
		_w2232_,
		_w2243_,
		_w9360_
	);
	LUT2 #(
		.INIT('hd)
	) name7611 (
		_w7486_,
		_w9360_,
		_w9361_
	);
	LUT3 #(
		.INIT('h2a)
	) name7612 (
		\u4_u0_buf0_orig_reg[30]/NET0131 ,
		_w2232_,
		_w2243_,
		_w9362_
	);
	LUT2 #(
		.INIT('hd)
	) name7613 (
		_w7491_,
		_w9362_,
		_w9363_
	);
	LUT3 #(
		.INIT('h2a)
	) name7614 (
		\u4_u0_buf0_orig_reg[31]/P0001 ,
		_w2232_,
		_w2243_,
		_w9364_
	);
	LUT2 #(
		.INIT('hd)
	) name7615 (
		_w7496_,
		_w9364_,
		_w9365_
	);
	LUT3 #(
		.INIT('h2a)
	) name7616 (
		\u4_u0_buf0_orig_reg[3]/P0001 ,
		_w2232_,
		_w2243_,
		_w9366_
	);
	LUT2 #(
		.INIT('hd)
	) name7617 (
		_w7501_,
		_w9366_,
		_w9367_
	);
	LUT3 #(
		.INIT('h2a)
	) name7618 (
		\u4_u0_buf0_orig_reg[4]/P0001 ,
		_w2232_,
		_w2243_,
		_w9368_
	);
	LUT2 #(
		.INIT('hd)
	) name7619 (
		_w2545_,
		_w9368_,
		_w9369_
	);
	LUT3 #(
		.INIT('h2a)
	) name7620 (
		\u4_u0_buf0_orig_reg[5]/P0001 ,
		_w2232_,
		_w2243_,
		_w9370_
	);
	LUT2 #(
		.INIT('hd)
	) name7621 (
		_w2550_,
		_w9370_,
		_w9371_
	);
	LUT3 #(
		.INIT('h2a)
	) name7622 (
		\u4_u0_buf0_orig_reg[6]/P0001 ,
		_w2232_,
		_w2243_,
		_w9372_
	);
	LUT2 #(
		.INIT('hd)
	) name7623 (
		_w2424_,
		_w9372_,
		_w9373_
	);
	LUT3 #(
		.INIT('h2a)
	) name7624 (
		\u4_u0_buf0_orig_reg[7]/P0001 ,
		_w2232_,
		_w2243_,
		_w9374_
	);
	LUT2 #(
		.INIT('hd)
	) name7625 (
		_w2555_,
		_w9374_,
		_w9375_
	);
	LUT3 #(
		.INIT('h2a)
	) name7626 (
		\u4_u0_buf0_orig_reg[8]/P0001 ,
		_w2232_,
		_w2243_,
		_w9376_
	);
	LUT2 #(
		.INIT('hd)
	) name7627 (
		_w7506_,
		_w9376_,
		_w9377_
	);
	LUT3 #(
		.INIT('h2a)
	) name7628 (
		\u4_u0_buf0_orig_reg[9]/P0001 ,
		_w2232_,
		_w2243_,
		_w9378_
	);
	LUT2 #(
		.INIT('hd)
	) name7629 (
		_w7511_,
		_w9378_,
		_w9379_
	);
	LUT3 #(
		.INIT('h02)
	) name7630 (
		\u4_u1_csr1_reg[8]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w9380_
	);
	LUT4 #(
		.INIT('h35ff)
	) name7631 (
		\u4_u1_buf0_reg[23]/P0001 ,
		\u4_u1_buf1_reg[23]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w9381_
	);
	LUT4 #(
		.INIT('h8088)
	) name7632 (
		_w2227_,
		_w2241_,
		_w9380_,
		_w9381_,
		_w9382_
	);
	LUT3 #(
		.INIT('h02)
	) name7633 (
		\u4_u2_csr1_reg[8]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w9383_
	);
	LUT4 #(
		.INIT('h35ff)
	) name7634 (
		\u4_u2_buf0_reg[23]/P0001 ,
		\u4_u2_buf1_reg[23]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w9384_
	);
	LUT4 #(
		.INIT('h8088)
	) name7635 (
		_w2228_,
		_w2240_,
		_w9383_,
		_w9384_,
		_w9385_
	);
	LUT3 #(
		.INIT('h02)
	) name7636 (
		\u4_u3_csr1_reg[8]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w9386_
	);
	LUT4 #(
		.INIT('h35ff)
	) name7637 (
		\u4_u3_buf0_reg[23]/P0001 ,
		\u4_u3_buf1_reg[23]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w9387_
	);
	LUT4 #(
		.INIT('h8088)
	) name7638 (
		_w2227_,
		_w2228_,
		_w9386_,
		_w9387_,
		_w9388_
	);
	LUT3 #(
		.INIT('h01)
	) name7639 (
		_w9382_,
		_w9385_,
		_w9388_,
		_w9389_
	);
	LUT4 #(
		.INIT('h0200)
	) name7640 (
		\u1_frame_no_r_reg[7]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w9390_
	);
	LUT4 #(
		.INIT('h0020)
	) name7641 (
		\u4_intb_msk_reg[7]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w9391_
	);
	LUT4 #(
		.INIT('h0080)
	) name7642 (
		\u4_int_srcb_reg[3]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w9392_
	);
	LUT4 #(
		.INIT('haaa8)
	) name7643 (
		_w5861_,
		_w9390_,
		_w9391_,
		_w9392_,
		_w9393_
	);
	LUT3 #(
		.INIT('h02)
	) name7644 (
		\u4_u0_csr1_reg[8]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w9394_
	);
	LUT4 #(
		.INIT('h35ff)
	) name7645 (
		\u4_u0_buf0_reg[23]/P0001 ,
		\u4_u0_buf1_reg[23]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w9395_
	);
	LUT4 #(
		.INIT('h8088)
	) name7646 (
		_w2240_,
		_w2241_,
		_w9394_,
		_w9395_,
		_w9396_
	);
	LUT2 #(
		.INIT('h1)
	) name7647 (
		_w9393_,
		_w9396_,
		_w9397_
	);
	LUT2 #(
		.INIT('h7)
	) name7648 (
		_w9389_,
		_w9397_,
		_w9398_
	);
	LUT4 #(
		.INIT('h2000)
	) name7649 (
		\u0_rx_active_reg/P0001 ,
		\u0_rx_err_reg/P0001 ,
		\u0_rx_valid_reg/P0001 ,
		\u1_u0_rxv2_reg/P0001 ,
		_w9399_
	);
	LUT4 #(
		.INIT('hba00)
	) name7650 (
		_w3671_,
		_w4886_,
		_w6898_,
		_w9399_,
		_w9400_
	);
	LUT2 #(
		.INIT('h8)
	) name7651 (
		rst_i_pad,
		\u4_u0_csr0_reg[0]/P0001 ,
		_w9401_
	);
	LUT4 #(
		.INIT('h5f08)
	) name7652 (
		_w2243_,
		_w9110_,
		_w9173_,
		_w9401_,
		_w9402_
	);
	LUT2 #(
		.INIT('h8)
	) name7653 (
		rst_i_pad,
		\u4_u0_csr0_reg[10]/P0001 ,
		_w9403_
	);
	LUT4 #(
		.INIT('h5f08)
	) name7654 (
		_w2243_,
		_w9110_,
		_w9176_,
		_w9403_,
		_w9404_
	);
	LUT2 #(
		.INIT('h8)
	) name7655 (
		rst_i_pad,
		\u4_u0_csr0_reg[11]/P0001 ,
		_w9405_
	);
	LUT4 #(
		.INIT('h5f08)
	) name7656 (
		_w2243_,
		_w9110_,
		_w9179_,
		_w9405_,
		_w9406_
	);
	LUT2 #(
		.INIT('h8)
	) name7657 (
		rst_i_pad,
		\u4_u0_csr0_reg[12]/P0001 ,
		_w9407_
	);
	LUT4 #(
		.INIT('h5f08)
	) name7658 (
		_w2243_,
		_w9110_,
		_w9182_,
		_w9407_,
		_w9408_
	);
	LUT2 #(
		.INIT('h8)
	) name7659 (
		rst_i_pad,
		\u4_u0_csr0_reg[1]/P0001 ,
		_w9409_
	);
	LUT4 #(
		.INIT('h5f08)
	) name7660 (
		_w2243_,
		_w9110_,
		_w9185_,
		_w9409_,
		_w9410_
	);
	LUT2 #(
		.INIT('h8)
	) name7661 (
		rst_i_pad,
		\u4_u0_csr0_reg[2]/P0001 ,
		_w9411_
	);
	LUT4 #(
		.INIT('h5f08)
	) name7662 (
		_w2243_,
		_w9110_,
		_w9188_,
		_w9411_,
		_w9412_
	);
	LUT2 #(
		.INIT('h8)
	) name7663 (
		rst_i_pad,
		\u4_u0_csr0_reg[3]/NET0131 ,
		_w9413_
	);
	LUT4 #(
		.INIT('h5f08)
	) name7664 (
		_w2243_,
		_w9110_,
		_w9191_,
		_w9413_,
		_w9414_
	);
	LUT2 #(
		.INIT('h8)
	) name7665 (
		rst_i_pad,
		\u4_u0_csr0_reg[4]/P0001 ,
		_w9415_
	);
	LUT4 #(
		.INIT('h5f08)
	) name7666 (
		_w2243_,
		_w9110_,
		_w9194_,
		_w9415_,
		_w9416_
	);
	LUT2 #(
		.INIT('h8)
	) name7667 (
		rst_i_pad,
		\u4_u0_csr0_reg[5]/P0001 ,
		_w9417_
	);
	LUT4 #(
		.INIT('h5f08)
	) name7668 (
		_w2243_,
		_w9110_,
		_w9197_,
		_w9417_,
		_w9418_
	);
	LUT2 #(
		.INIT('h8)
	) name7669 (
		rst_i_pad,
		\u4_u0_csr0_reg[6]/P0001 ,
		_w9419_
	);
	LUT4 #(
		.INIT('h5f08)
	) name7670 (
		_w2243_,
		_w9110_,
		_w9200_,
		_w9419_,
		_w9420_
	);
	LUT2 #(
		.INIT('h8)
	) name7671 (
		rst_i_pad,
		\u4_u0_csr0_reg[7]/P0001 ,
		_w9421_
	);
	LUT4 #(
		.INIT('h5f08)
	) name7672 (
		_w2243_,
		_w9110_,
		_w9203_,
		_w9421_,
		_w9422_
	);
	LUT2 #(
		.INIT('h8)
	) name7673 (
		rst_i_pad,
		\u4_u0_csr0_reg[8]/P0001 ,
		_w9423_
	);
	LUT4 #(
		.INIT('h5f08)
	) name7674 (
		_w2243_,
		_w9110_,
		_w9206_,
		_w9423_,
		_w9424_
	);
	LUT2 #(
		.INIT('h8)
	) name7675 (
		rst_i_pad,
		\u4_u0_csr0_reg[9]/P0001 ,
		_w9425_
	);
	LUT4 #(
		.INIT('h5f08)
	) name7676 (
		_w2243_,
		_w9110_,
		_w9209_,
		_w9425_,
		_w9426_
	);
	LUT2 #(
		.INIT('h8)
	) name7677 (
		rst_i_pad,
		\u4_u0_csr1_reg[0]/P0001 ,
		_w9427_
	);
	LUT4 #(
		.INIT('h5f08)
	) name7678 (
		_w2243_,
		_w9110_,
		_w9170_,
		_w9427_,
		_w9428_
	);
	LUT2 #(
		.INIT('h8)
	) name7679 (
		rst_i_pad,
		\u4_u0_csr1_reg[10]/P0001 ,
		_w9429_
	);
	LUT4 #(
		.INIT('h5f08)
	) name7680 (
		_w2243_,
		_w9110_,
		_w9214_,
		_w9429_,
		_w9430_
	);
	LUT2 #(
		.INIT('h8)
	) name7681 (
		rst_i_pad,
		\u4_u0_csr1_reg[11]/P0001 ,
		_w9431_
	);
	LUT4 #(
		.INIT('h5f08)
	) name7682 (
		_w2243_,
		_w9110_,
		_w9217_,
		_w9431_,
		_w9432_
	);
	LUT2 #(
		.INIT('h8)
	) name7683 (
		rst_i_pad,
		\u4_u0_csr1_reg[12]/P0001 ,
		_w9433_
	);
	LUT4 #(
		.INIT('h5f08)
	) name7684 (
		_w2243_,
		_w9110_,
		_w9220_,
		_w9433_,
		_w9434_
	);
	LUT2 #(
		.INIT('h8)
	) name7685 (
		rst_i_pad,
		\u4_u0_csr1_reg[1]/P0001 ,
		_w9435_
	);
	LUT4 #(
		.INIT('h5f08)
	) name7686 (
		_w2243_,
		_w9110_,
		_w9223_,
		_w9435_,
		_w9436_
	);
	LUT2 #(
		.INIT('h8)
	) name7687 (
		rst_i_pad,
		\u4_u0_csr1_reg[2]/P0001 ,
		_w9437_
	);
	LUT4 #(
		.INIT('h5f08)
	) name7688 (
		_w2243_,
		_w9110_,
		_w9226_,
		_w9437_,
		_w9438_
	);
	LUT2 #(
		.INIT('h8)
	) name7689 (
		rst_i_pad,
		\u4_u0_csr1_reg[3]/P0001 ,
		_w9439_
	);
	LUT4 #(
		.INIT('h5f08)
	) name7690 (
		_w2243_,
		_w9110_,
		_w9229_,
		_w9439_,
		_w9440_
	);
	LUT2 #(
		.INIT('h8)
	) name7691 (
		rst_i_pad,
		\u4_u0_csr1_reg[4]/P0001 ,
		_w9441_
	);
	LUT4 #(
		.INIT('h5f08)
	) name7692 (
		_w2243_,
		_w9110_,
		_w9232_,
		_w9441_,
		_w9442_
	);
	LUT2 #(
		.INIT('h8)
	) name7693 (
		rst_i_pad,
		\u4_u0_csr1_reg[5]/P0001 ,
		_w9443_
	);
	LUT4 #(
		.INIT('h5f08)
	) name7694 (
		_w2243_,
		_w9110_,
		_w9235_,
		_w9443_,
		_w9444_
	);
	LUT2 #(
		.INIT('h8)
	) name7695 (
		rst_i_pad,
		\u4_u0_csr1_reg[6]/P0001 ,
		_w9445_
	);
	LUT4 #(
		.INIT('h5f08)
	) name7696 (
		_w2243_,
		_w9110_,
		_w9238_,
		_w9445_,
		_w9446_
	);
	LUT2 #(
		.INIT('h8)
	) name7697 (
		rst_i_pad,
		\u4_u0_csr1_reg[9]/P0001 ,
		_w9447_
	);
	LUT4 #(
		.INIT('h5f08)
	) name7698 (
		_w2243_,
		_w9110_,
		_w9241_,
		_w9447_,
		_w9448_
	);
	LUT3 #(
		.INIT('h2a)
	) name7699 (
		\u4_u3_buf0_orig_reg[21]/P0001 ,
		_w2231_,
		_w2232_,
		_w9449_
	);
	LUT2 #(
		.INIT('hd)
	) name7700 (
		_w7304_,
		_w9449_,
		_w9450_
	);
	LUT2 #(
		.INIT('h8)
	) name7701 (
		rst_i_pad,
		\u4_u0_iena_reg[0]/P0001 ,
		_w9451_
	);
	LUT4 #(
		.INIT('h7720)
	) name7702 (
		_w2243_,
		_w9067_,
		_w9069_,
		_w9451_,
		_w9452_
	);
	LUT2 #(
		.INIT('h8)
	) name7703 (
		rst_i_pad,
		\u4_u0_iena_reg[1]/P0001 ,
		_w9453_
	);
	LUT4 #(
		.INIT('h5f08)
	) name7704 (
		_w2243_,
		_w9069_,
		_w9071_,
		_w9453_,
		_w9454_
	);
	LUT2 #(
		.INIT('h8)
	) name7705 (
		rst_i_pad,
		\u4_u0_iena_reg[2]/P0001 ,
		_w9455_
	);
	LUT4 #(
		.INIT('h5f08)
	) name7706 (
		_w2243_,
		_w9069_,
		_w9074_,
		_w9455_,
		_w9456_
	);
	LUT2 #(
		.INIT('h8)
	) name7707 (
		rst_i_pad,
		\u4_u0_iena_reg[3]/P0001 ,
		_w9457_
	);
	LUT4 #(
		.INIT('h5f08)
	) name7708 (
		_w2243_,
		_w9069_,
		_w9077_,
		_w9457_,
		_w9458_
	);
	LUT2 #(
		.INIT('h8)
	) name7709 (
		rst_i_pad,
		\u4_u0_iena_reg[4]/P0001 ,
		_w9459_
	);
	LUT4 #(
		.INIT('h5f08)
	) name7710 (
		_w2243_,
		_w9069_,
		_w9080_,
		_w9459_,
		_w9460_
	);
	LUT2 #(
		.INIT('h8)
	) name7711 (
		rst_i_pad,
		\u4_u0_iena_reg[5]/P0001 ,
		_w9461_
	);
	LUT4 #(
		.INIT('h5f08)
	) name7712 (
		_w2243_,
		_w9069_,
		_w9083_,
		_w9461_,
		_w9462_
	);
	LUT2 #(
		.INIT('h8)
	) name7713 (
		rst_i_pad,
		\u4_u0_ienb_reg[0]/P0001 ,
		_w9463_
	);
	LUT4 #(
		.INIT('h5f08)
	) name7714 (
		_w2243_,
		_w9069_,
		_w9086_,
		_w9463_,
		_w9464_
	);
	LUT2 #(
		.INIT('h8)
	) name7715 (
		rst_i_pad,
		\u4_u0_ienb_reg[1]/P0001 ,
		_w9465_
	);
	LUT4 #(
		.INIT('h5f08)
	) name7716 (
		_w2243_,
		_w9069_,
		_w9089_,
		_w9465_,
		_w9466_
	);
	LUT2 #(
		.INIT('h8)
	) name7717 (
		rst_i_pad,
		\u4_u0_ienb_reg[2]/P0001 ,
		_w9467_
	);
	LUT4 #(
		.INIT('h5f08)
	) name7718 (
		_w2243_,
		_w9069_,
		_w9092_,
		_w9467_,
		_w9468_
	);
	LUT2 #(
		.INIT('h8)
	) name7719 (
		rst_i_pad,
		\u4_u0_ienb_reg[3]/P0001 ,
		_w9469_
	);
	LUT4 #(
		.INIT('h5f08)
	) name7720 (
		_w2243_,
		_w9069_,
		_w9095_,
		_w9469_,
		_w9470_
	);
	LUT2 #(
		.INIT('h8)
	) name7721 (
		rst_i_pad,
		\u4_u0_ienb_reg[4]/P0001 ,
		_w9471_
	);
	LUT4 #(
		.INIT('h5f08)
	) name7722 (
		_w2243_,
		_w9069_,
		_w9098_,
		_w9471_,
		_w9472_
	);
	LUT2 #(
		.INIT('h8)
	) name7723 (
		rst_i_pad,
		\u4_u0_ienb_reg[5]/P0001 ,
		_w9473_
	);
	LUT4 #(
		.INIT('h5f08)
	) name7724 (
		_w2243_,
		_w9069_,
		_w9101_,
		_w9473_,
		_w9474_
	);
	LUT3 #(
		.INIT('h20)
	) name7725 (
		rst_i_pad,
		\u4_u0_int_re_reg/P0001 ,
		\u4_u0_int_stat_reg[1]/P0001 ,
		_w9475_
	);
	LUT3 #(
		.INIT('hd0)
	) name7726 (
		\u0_rx_active_reg/P0001 ,
		\u0_rx_err_reg/P0001 ,
		\u4_u0_ep_match_r_reg/P0001 ,
		_w9476_
	);
	LUT3 #(
		.INIT('h80)
	) name7727 (
		_w3671_,
		_w3896_,
		_w9476_,
		_w9477_
	);
	LUT3 #(
		.INIT('hdc)
	) name7728 (
		_w3682_,
		_w9475_,
		_w9477_,
		_w9478_
	);
	LUT2 #(
		.INIT('h8)
	) name7729 (
		rst_i_pad,
		\u4_u0_ots_stop_reg/P0001 ,
		_w9479_
	);
	LUT4 #(
		.INIT('h7720)
	) name7730 (
		_w2243_,
		_w9108_,
		_w9110_,
		_w9479_,
		_w9480_
	);
	LUT3 #(
		.INIT('h2a)
	) name7731 (
		\u4_u1_buf0_orig_reg[0]/P0001 ,
		_w2232_,
		_w2260_,
		_w9481_
	);
	LUT2 #(
		.INIT('hd)
	) name7732 (
		_w7524_,
		_w9481_,
		_w9482_
	);
	LUT3 #(
		.INIT('h2a)
	) name7733 (
		\u4_u1_buf0_orig_reg[10]/P0001 ,
		_w2232_,
		_w2260_,
		_w9483_
	);
	LUT2 #(
		.INIT('hd)
	) name7734 (
		_w2285_,
		_w9483_,
		_w9484_
	);
	LUT3 #(
		.INIT('h2a)
	) name7735 (
		\u4_u1_buf0_orig_reg[11]/P0001 ,
		_w2232_,
		_w2260_,
		_w9485_
	);
	LUT2 #(
		.INIT('hd)
	) name7736 (
		_w2435_,
		_w9485_,
		_w9486_
	);
	LUT3 #(
		.INIT('h2a)
	) name7737 (
		\u4_u1_buf0_orig_reg[12]/P0001 ,
		_w2232_,
		_w2260_,
		_w9487_
	);
	LUT2 #(
		.INIT('hd)
	) name7738 (
		_w7529_,
		_w9487_,
		_w9488_
	);
	LUT3 #(
		.INIT('h2a)
	) name7739 (
		\u4_u1_buf0_orig_reg[13]/P0001 ,
		_w2232_,
		_w2260_,
		_w9489_
	);
	LUT2 #(
		.INIT('hd)
	) name7740 (
		_w2339_,
		_w9489_,
		_w9490_
	);
	LUT3 #(
		.INIT('h2a)
	) name7741 (
		\u4_u1_buf0_orig_reg[14]/P0001 ,
		_w2232_,
		_w2260_,
		_w9491_
	);
	LUT2 #(
		.INIT('hd)
	) name7742 (
		_w2261_,
		_w9491_,
		_w9492_
	);
	LUT3 #(
		.INIT('h2a)
	) name7743 (
		\u4_u1_buf0_orig_reg[15]/P0001 ,
		_w2232_,
		_w2260_,
		_w9493_
	);
	LUT2 #(
		.INIT('hd)
	) name7744 (
		_w2440_,
		_w9493_,
		_w9494_
	);
	LUT3 #(
		.INIT('h2a)
	) name7745 (
		\u4_u1_buf0_orig_reg[16]/P0001 ,
		_w2232_,
		_w2260_,
		_w9495_
	);
	LUT2 #(
		.INIT('hd)
	) name7746 (
		_w7534_,
		_w9495_,
		_w9496_
	);
	LUT3 #(
		.INIT('h2a)
	) name7747 (
		\u4_u1_buf0_orig_reg[17]/P0001 ,
		_w2232_,
		_w2260_,
		_w9497_
	);
	LUT2 #(
		.INIT('hd)
	) name7748 (
		_w7539_,
		_w9497_,
		_w9498_
	);
	LUT3 #(
		.INIT('h2a)
	) name7749 (
		\u4_u1_buf0_orig_reg[18]/P0001 ,
		_w2232_,
		_w2260_,
		_w9499_
	);
	LUT2 #(
		.INIT('hd)
	) name7750 (
		_w7544_,
		_w9499_,
		_w9500_
	);
	LUT3 #(
		.INIT('h2a)
	) name7751 (
		\u4_u1_buf0_orig_reg[19]/P0001 ,
		_w2232_,
		_w2260_,
		_w9501_
	);
	LUT2 #(
		.INIT('hd)
	) name7752 (
		_w7549_,
		_w9501_,
		_w9502_
	);
	LUT3 #(
		.INIT('h2a)
	) name7753 (
		\u4_u1_buf0_orig_reg[1]/P0001 ,
		_w2232_,
		_w2260_,
		_w9503_
	);
	LUT2 #(
		.INIT('hd)
	) name7754 (
		_w7554_,
		_w9503_,
		_w9504_
	);
	LUT3 #(
		.INIT('h2a)
	) name7755 (
		\u4_u1_buf0_orig_reg[20]/P0001 ,
		_w2232_,
		_w2260_,
		_w9505_
	);
	LUT2 #(
		.INIT('hd)
	) name7756 (
		_w7559_,
		_w9505_,
		_w9506_
	);
	LUT3 #(
		.INIT('h2a)
	) name7757 (
		\u4_u1_buf0_orig_reg[21]/P0001 ,
		_w2232_,
		_w2260_,
		_w9507_
	);
	LUT2 #(
		.INIT('hd)
	) name7758 (
		_w7564_,
		_w9507_,
		_w9508_
	);
	LUT3 #(
		.INIT('h2a)
	) name7759 (
		\u4_u1_buf0_orig_reg[22]/P0001 ,
		_w2232_,
		_w2260_,
		_w9509_
	);
	LUT2 #(
		.INIT('hd)
	) name7760 (
		_w7569_,
		_w9509_,
		_w9510_
	);
	LUT3 #(
		.INIT('h2a)
	) name7761 (
		\u4_u1_buf0_orig_reg[23]/P0001 ,
		_w2232_,
		_w2260_,
		_w9511_
	);
	LUT2 #(
		.INIT('hd)
	) name7762 (
		_w7574_,
		_w9511_,
		_w9512_
	);
	LUT3 #(
		.INIT('h2a)
	) name7763 (
		\u4_u1_buf0_orig_reg[24]/P0001 ,
		_w2232_,
		_w2260_,
		_w9513_
	);
	LUT2 #(
		.INIT('hd)
	) name7764 (
		_w7579_,
		_w9513_,
		_w9514_
	);
	LUT3 #(
		.INIT('h2a)
	) name7765 (
		\u4_u1_buf0_orig_reg[25]/P0001 ,
		_w2232_,
		_w2260_,
		_w9515_
	);
	LUT2 #(
		.INIT('hd)
	) name7766 (
		_w7584_,
		_w9515_,
		_w9516_
	);
	LUT3 #(
		.INIT('h2a)
	) name7767 (
		\u4_u1_buf0_orig_reg[26]/P0001 ,
		_w2232_,
		_w2260_,
		_w9517_
	);
	LUT2 #(
		.INIT('hd)
	) name7768 (
		_w7589_,
		_w9517_,
		_w9518_
	);
	LUT3 #(
		.INIT('h2a)
	) name7769 (
		\u4_u1_buf0_orig_reg[27]/P0001 ,
		_w2232_,
		_w2260_,
		_w9519_
	);
	LUT2 #(
		.INIT('hd)
	) name7770 (
		_w7594_,
		_w9519_,
		_w9520_
	);
	LUT3 #(
		.INIT('h2a)
	) name7771 (
		\u4_u1_buf0_orig_reg[28]/P0001 ,
		_w2232_,
		_w2260_,
		_w9521_
	);
	LUT2 #(
		.INIT('hd)
	) name7772 (
		_w7599_,
		_w9521_,
		_w9522_
	);
	LUT3 #(
		.INIT('h2a)
	) name7773 (
		\u4_u1_buf0_orig_reg[29]/NET0131 ,
		_w2232_,
		_w2260_,
		_w9523_
	);
	LUT2 #(
		.INIT('hd)
	) name7774 (
		_w7604_,
		_w9523_,
		_w9524_
	);
	LUT3 #(
		.INIT('h2a)
	) name7775 (
		\u4_u1_buf0_orig_reg[2]/P0001 ,
		_w2232_,
		_w2260_,
		_w9525_
	);
	LUT2 #(
		.INIT('hd)
	) name7776 (
		_w7609_,
		_w9525_,
		_w9526_
	);
	LUT3 #(
		.INIT('h2a)
	) name7777 (
		\u4_u1_buf0_orig_reg[30]/NET0131 ,
		_w2232_,
		_w2260_,
		_w9527_
	);
	LUT2 #(
		.INIT('hd)
	) name7778 (
		_w7614_,
		_w9527_,
		_w9528_
	);
	LUT3 #(
		.INIT('h2a)
	) name7779 (
		\u4_u1_buf0_orig_reg[31]/P0001 ,
		_w2232_,
		_w2260_,
		_w9529_
	);
	LUT2 #(
		.INIT('hd)
	) name7780 (
		_w7619_,
		_w9529_,
		_w9530_
	);
	LUT3 #(
		.INIT('h2a)
	) name7781 (
		\u4_u1_buf0_orig_reg[3]/P0001 ,
		_w2232_,
		_w2260_,
		_w9531_
	);
	LUT2 #(
		.INIT('hd)
	) name7782 (
		_w7624_,
		_w9531_,
		_w9532_
	);
	LUT3 #(
		.INIT('h2a)
	) name7783 (
		\u4_u1_buf0_orig_reg[4]/P0001 ,
		_w2232_,
		_w2260_,
		_w9533_
	);
	LUT2 #(
		.INIT('hd)
	) name7784 (
		_w2578_,
		_w9533_,
		_w9534_
	);
	LUT3 #(
		.INIT('h2a)
	) name7785 (
		\u4_u1_buf0_orig_reg[5]/P0001 ,
		_w2232_,
		_w2260_,
		_w9535_
	);
	LUT2 #(
		.INIT('hd)
	) name7786 (
		_w2583_,
		_w9535_,
		_w9536_
	);
	LUT3 #(
		.INIT('h2a)
	) name7787 (
		\u4_u1_buf0_orig_reg[6]/P0001 ,
		_w2232_,
		_w2260_,
		_w9537_
	);
	LUT2 #(
		.INIT('hd)
	) name7788 (
		_w2451_,
		_w9537_,
		_w9538_
	);
	LUT3 #(
		.INIT('h2a)
	) name7789 (
		\u4_u1_buf0_orig_reg[7]/P0001 ,
		_w2232_,
		_w2260_,
		_w9539_
	);
	LUT2 #(
		.INIT('hd)
	) name7790 (
		_w2588_,
		_w9539_,
		_w9540_
	);
	LUT3 #(
		.INIT('h2a)
	) name7791 (
		\u4_u1_buf0_orig_reg[8]/P0001 ,
		_w2232_,
		_w2260_,
		_w9541_
	);
	LUT2 #(
		.INIT('hd)
	) name7792 (
		_w7629_,
		_w9541_,
		_w9542_
	);
	LUT3 #(
		.INIT('h2a)
	) name7793 (
		\u4_u1_buf0_orig_reg[9]/P0001 ,
		_w2232_,
		_w2260_,
		_w9543_
	);
	LUT2 #(
		.INIT('hd)
	) name7794 (
		_w7634_,
		_w9543_,
		_w9544_
	);
	LUT4 #(
		.INIT('hddcd)
	) name7795 (
		\u1_u2_mack_r_reg/P0001 ,
		\u1_u2_word_done_r_reg/P0001 ,
		_w3224_,
		_w5488_,
		_w9545_
	);
	LUT2 #(
		.INIT('h8)
	) name7796 (
		rst_i_pad,
		\u4_u1_csr0_reg[0]/P0001 ,
		_w9546_
	);
	LUT4 #(
		.INIT('h5f08)
	) name7797 (
		_w2260_,
		_w9110_,
		_w9173_,
		_w9546_,
		_w9547_
	);
	LUT2 #(
		.INIT('h8)
	) name7798 (
		rst_i_pad,
		\u4_u1_csr0_reg[10]/P0001 ,
		_w9548_
	);
	LUT4 #(
		.INIT('h5f08)
	) name7799 (
		_w2260_,
		_w9110_,
		_w9176_,
		_w9548_,
		_w9549_
	);
	LUT2 #(
		.INIT('h8)
	) name7800 (
		rst_i_pad,
		\u4_u1_csr0_reg[11]/P0001 ,
		_w9550_
	);
	LUT4 #(
		.INIT('h5f08)
	) name7801 (
		_w2260_,
		_w9110_,
		_w9179_,
		_w9550_,
		_w9551_
	);
	LUT2 #(
		.INIT('h8)
	) name7802 (
		rst_i_pad,
		\u4_u1_csr0_reg[12]/P0001 ,
		_w9552_
	);
	LUT4 #(
		.INIT('h5f08)
	) name7803 (
		_w2260_,
		_w9110_,
		_w9182_,
		_w9552_,
		_w9553_
	);
	LUT2 #(
		.INIT('h8)
	) name7804 (
		rst_i_pad,
		\u4_u1_csr0_reg[1]/P0001 ,
		_w9554_
	);
	LUT4 #(
		.INIT('h5f08)
	) name7805 (
		_w2260_,
		_w9110_,
		_w9185_,
		_w9554_,
		_w9555_
	);
	LUT2 #(
		.INIT('h8)
	) name7806 (
		rst_i_pad,
		\u4_u1_csr0_reg[2]/P0001 ,
		_w9556_
	);
	LUT4 #(
		.INIT('h5f08)
	) name7807 (
		_w2260_,
		_w9110_,
		_w9188_,
		_w9556_,
		_w9557_
	);
	LUT2 #(
		.INIT('h8)
	) name7808 (
		rst_i_pad,
		\u4_u1_csr0_reg[3]/NET0131 ,
		_w9558_
	);
	LUT4 #(
		.INIT('h5f08)
	) name7809 (
		_w2260_,
		_w9110_,
		_w9191_,
		_w9558_,
		_w9559_
	);
	LUT4 #(
		.INIT('h007f)
	) name7810 (
		\u1_u3_rx_ack_to_cnt_reg[0]/P0001 ,
		\u1_u3_rx_ack_to_cnt_reg[1]/P0001 ,
		\u1_u3_rx_ack_to_cnt_reg[2]/P0001 ,
		\u1_u3_rx_ack_to_cnt_reg[3]/P0001 ,
		_w9560_
	);
	LUT3 #(
		.INIT('h01)
	) name7811 (
		\u1_u3_rx_ack_to_clr_reg/P0001 ,
		_w7951_,
		_w9560_,
		_w9561_
	);
	LUT2 #(
		.INIT('h8)
	) name7812 (
		rst_i_pad,
		\u4_u1_csr0_reg[4]/P0001 ,
		_w9562_
	);
	LUT4 #(
		.INIT('h5f08)
	) name7813 (
		_w2260_,
		_w9110_,
		_w9194_,
		_w9562_,
		_w9563_
	);
	LUT2 #(
		.INIT('h8)
	) name7814 (
		rst_i_pad,
		\u4_u1_csr0_reg[5]/P0001 ,
		_w9564_
	);
	LUT4 #(
		.INIT('h5f08)
	) name7815 (
		_w2260_,
		_w9110_,
		_w9197_,
		_w9564_,
		_w9565_
	);
	LUT2 #(
		.INIT('h8)
	) name7816 (
		rst_i_pad,
		\u4_u1_csr0_reg[6]/P0001 ,
		_w9566_
	);
	LUT4 #(
		.INIT('h5f08)
	) name7817 (
		_w2260_,
		_w9110_,
		_w9200_,
		_w9566_,
		_w9567_
	);
	LUT2 #(
		.INIT('h8)
	) name7818 (
		rst_i_pad,
		\u4_u1_csr0_reg[7]/P0001 ,
		_w9568_
	);
	LUT4 #(
		.INIT('h5f08)
	) name7819 (
		_w2260_,
		_w9110_,
		_w9203_,
		_w9568_,
		_w9569_
	);
	LUT2 #(
		.INIT('h8)
	) name7820 (
		rst_i_pad,
		\u4_u1_csr0_reg[8]/P0001 ,
		_w9570_
	);
	LUT4 #(
		.INIT('h5f08)
	) name7821 (
		_w2260_,
		_w9110_,
		_w9206_,
		_w9570_,
		_w9571_
	);
	LUT2 #(
		.INIT('h8)
	) name7822 (
		rst_i_pad,
		\u4_u1_csr0_reg[9]/P0001 ,
		_w9572_
	);
	LUT4 #(
		.INIT('h5f08)
	) name7823 (
		_w2260_,
		_w9110_,
		_w9209_,
		_w9572_,
		_w9573_
	);
	LUT2 #(
		.INIT('h8)
	) name7824 (
		rst_i_pad,
		\u4_u1_csr1_reg[0]/P0001 ,
		_w9574_
	);
	LUT4 #(
		.INIT('h5f08)
	) name7825 (
		_w2260_,
		_w9110_,
		_w9170_,
		_w9574_,
		_w9575_
	);
	LUT2 #(
		.INIT('h8)
	) name7826 (
		rst_i_pad,
		\u4_u1_csr1_reg[10]/P0001 ,
		_w9576_
	);
	LUT4 #(
		.INIT('h5f08)
	) name7827 (
		_w2260_,
		_w9110_,
		_w9214_,
		_w9576_,
		_w9577_
	);
	LUT2 #(
		.INIT('h8)
	) name7828 (
		rst_i_pad,
		\u4_u1_csr1_reg[11]/P0001 ,
		_w9578_
	);
	LUT4 #(
		.INIT('h5f08)
	) name7829 (
		_w2260_,
		_w9110_,
		_w9217_,
		_w9578_,
		_w9579_
	);
	LUT2 #(
		.INIT('h8)
	) name7830 (
		rst_i_pad,
		\u4_u1_csr1_reg[12]/P0001 ,
		_w9580_
	);
	LUT4 #(
		.INIT('h5f08)
	) name7831 (
		_w2260_,
		_w9110_,
		_w9220_,
		_w9580_,
		_w9581_
	);
	LUT2 #(
		.INIT('h8)
	) name7832 (
		rst_i_pad,
		\u4_u1_csr1_reg[1]/P0001 ,
		_w9582_
	);
	LUT4 #(
		.INIT('h5f08)
	) name7833 (
		_w2260_,
		_w9110_,
		_w9223_,
		_w9582_,
		_w9583_
	);
	LUT2 #(
		.INIT('h8)
	) name7834 (
		rst_i_pad,
		\u4_u1_csr1_reg[2]/P0001 ,
		_w9584_
	);
	LUT4 #(
		.INIT('h5f08)
	) name7835 (
		_w2260_,
		_w9110_,
		_w9226_,
		_w9584_,
		_w9585_
	);
	LUT2 #(
		.INIT('h8)
	) name7836 (
		rst_i_pad,
		\u4_u1_csr1_reg[3]/P0001 ,
		_w9586_
	);
	LUT4 #(
		.INIT('h5f08)
	) name7837 (
		_w2260_,
		_w9110_,
		_w9229_,
		_w9586_,
		_w9587_
	);
	LUT2 #(
		.INIT('h8)
	) name7838 (
		rst_i_pad,
		\u4_u1_csr1_reg[4]/P0001 ,
		_w9588_
	);
	LUT4 #(
		.INIT('h5f08)
	) name7839 (
		_w2260_,
		_w9110_,
		_w9232_,
		_w9588_,
		_w9589_
	);
	LUT2 #(
		.INIT('h8)
	) name7840 (
		rst_i_pad,
		\u4_u1_csr1_reg[5]/P0001 ,
		_w9590_
	);
	LUT4 #(
		.INIT('h5f08)
	) name7841 (
		_w2260_,
		_w9110_,
		_w9235_,
		_w9590_,
		_w9591_
	);
	LUT2 #(
		.INIT('h8)
	) name7842 (
		rst_i_pad,
		\u4_u1_csr1_reg[6]/P0001 ,
		_w9592_
	);
	LUT4 #(
		.INIT('h5f08)
	) name7843 (
		_w2260_,
		_w9110_,
		_w9238_,
		_w9592_,
		_w9593_
	);
	LUT2 #(
		.INIT('h8)
	) name7844 (
		rst_i_pad,
		\u4_u1_csr1_reg[9]/P0001 ,
		_w9594_
	);
	LUT4 #(
		.INIT('h5f08)
	) name7845 (
		_w2260_,
		_w9110_,
		_w9241_,
		_w9594_,
		_w9595_
	);
	LUT4 #(
		.INIT('hcedf)
	) name7846 (
		\LineState_r_reg[0]/P0001 ,
		\LineState_r_reg[1]/P0001 ,
		\u0_u0_ls_j_r_reg/P0001 ,
		\u0_u0_ls_se0_r_reg/P0001 ,
		_w9596_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name7847 (
		\u0_u0_state_reg[11]/NET0131 ,
		\u0_u0_state_reg[12]/NET0131 ,
		_w4119_,
		_w9596_,
		_w9597_
	);
	LUT3 #(
		.INIT('h08)
	) name7848 (
		_w4110_,
		_w4122_,
		_w9597_,
		_w9598_
	);
	LUT4 #(
		.INIT('h007f)
	) name7849 (
		\u1_u3_tx_data_to_cnt_reg[0]/P0001 ,
		\u1_u3_tx_data_to_cnt_reg[1]/P0001 ,
		\u1_u3_tx_data_to_cnt_reg[2]/P0001 ,
		\u1_u3_tx_data_to_cnt_reg[3]/P0001 ,
		_w9599_
	);
	LUT3 #(
		.INIT('h01)
	) name7850 (
		\u0_rx_active_reg/P0001 ,
		_w7967_,
		_w9599_,
		_w9600_
	);
	LUT2 #(
		.INIT('h1)
	) name7851 (
		\u0_u0_T2_gt_1_0_mS_reg/P0001 ,
		\u0_u0_state_reg[4]/NET0131 ,
		_w9601_
	);
	LUT4 #(
		.INIT('h0004)
	) name7852 (
		\u0_u0_state_reg[10]/P0001 ,
		\u0_u0_state_reg[7]/NET0131 ,
		\u0_u0_state_reg[8]/NET0131 ,
		\u0_u0_state_reg[9]/P0001 ,
		_w9602_
	);
	LUT4 #(
		.INIT('h8000)
	) name7853 (
		_w4094_,
		_w4098_,
		_w4101_,
		_w9602_,
		_w9603_
	);
	LUT2 #(
		.INIT('h4)
	) name7854 (
		_w9601_,
		_w9603_,
		_w9604_
	);
	LUT3 #(
		.INIT('h70)
	) name7855 (
		\u0_u0_T1_gt_5_0_mS_reg/P0001 ,
		\u0_u0_resume_req_s_reg/P0001 ,
		\u0_u0_state_reg[4]/NET0131 ,
		_w9605_
	);
	LUT4 #(
		.INIT('h0c08)
	) name7856 (
		_w4119_,
		_w4341_,
		_w4354_,
		_w9605_,
		_w9606_
	);
	LUT4 #(
		.INIT('h00e0)
	) name7857 (
		\LineState_r_reg[0]/P0001 ,
		\LineState_r_reg[1]/P0001 ,
		\u0_u0_state_reg[4]/NET0131 ,
		\u0_u0_state_reg[5]/P0001 ,
		_w9607_
	);
	LUT4 #(
		.INIT('h153f)
	) name7858 (
		_w4319_,
		_w7962_,
		_w9606_,
		_w9607_,
		_w9608_
	);
	LUT3 #(
		.INIT('h8a)
	) name7859 (
		_w4103_,
		_w9604_,
		_w9608_,
		_w9609_
	);
	LUT2 #(
		.INIT('h8)
	) name7860 (
		rst_i_pad,
		\u4_u1_iena_reg[0]/P0001 ,
		_w9610_
	);
	LUT4 #(
		.INIT('h7720)
	) name7861 (
		_w2260_,
		_w9067_,
		_w9069_,
		_w9610_,
		_w9611_
	);
	LUT2 #(
		.INIT('h8)
	) name7862 (
		rst_i_pad,
		\u4_u1_iena_reg[1]/P0001 ,
		_w9612_
	);
	LUT4 #(
		.INIT('h5f08)
	) name7863 (
		_w2260_,
		_w9069_,
		_w9071_,
		_w9612_,
		_w9613_
	);
	LUT2 #(
		.INIT('h8)
	) name7864 (
		rst_i_pad,
		\u4_u1_iena_reg[2]/P0001 ,
		_w9614_
	);
	LUT4 #(
		.INIT('h5f08)
	) name7865 (
		_w2260_,
		_w9069_,
		_w9074_,
		_w9614_,
		_w9615_
	);
	LUT2 #(
		.INIT('h8)
	) name7866 (
		rst_i_pad,
		\u4_u1_iena_reg[3]/P0001 ,
		_w9616_
	);
	LUT4 #(
		.INIT('h5f08)
	) name7867 (
		_w2260_,
		_w9069_,
		_w9077_,
		_w9616_,
		_w9617_
	);
	LUT2 #(
		.INIT('h8)
	) name7868 (
		rst_i_pad,
		\u4_u1_iena_reg[4]/P0001 ,
		_w9618_
	);
	LUT4 #(
		.INIT('h5f08)
	) name7869 (
		_w2260_,
		_w9069_,
		_w9080_,
		_w9618_,
		_w9619_
	);
	LUT2 #(
		.INIT('h8)
	) name7870 (
		rst_i_pad,
		\u4_u1_iena_reg[5]/P0001 ,
		_w9620_
	);
	LUT4 #(
		.INIT('h5f08)
	) name7871 (
		_w2260_,
		_w9069_,
		_w9083_,
		_w9620_,
		_w9621_
	);
	LUT2 #(
		.INIT('h8)
	) name7872 (
		rst_i_pad,
		\u4_u1_ienb_reg[0]/P0001 ,
		_w9622_
	);
	LUT4 #(
		.INIT('h5f08)
	) name7873 (
		_w2260_,
		_w9069_,
		_w9086_,
		_w9622_,
		_w9623_
	);
	LUT2 #(
		.INIT('h8)
	) name7874 (
		rst_i_pad,
		\u4_u1_ienb_reg[1]/P0001 ,
		_w9624_
	);
	LUT4 #(
		.INIT('h5f08)
	) name7875 (
		_w2260_,
		_w9069_,
		_w9089_,
		_w9624_,
		_w9625_
	);
	LUT2 #(
		.INIT('h8)
	) name7876 (
		rst_i_pad,
		\u4_u1_ienb_reg[2]/P0001 ,
		_w9626_
	);
	LUT4 #(
		.INIT('h5f08)
	) name7877 (
		_w2260_,
		_w9069_,
		_w9092_,
		_w9626_,
		_w9627_
	);
	LUT2 #(
		.INIT('h8)
	) name7878 (
		rst_i_pad,
		\u4_u1_ienb_reg[3]/P0001 ,
		_w9628_
	);
	LUT4 #(
		.INIT('h5f08)
	) name7879 (
		_w2260_,
		_w9069_,
		_w9095_,
		_w9628_,
		_w9629_
	);
	LUT2 #(
		.INIT('h8)
	) name7880 (
		rst_i_pad,
		\u4_u1_ienb_reg[4]/P0001 ,
		_w9630_
	);
	LUT4 #(
		.INIT('h5f08)
	) name7881 (
		_w2260_,
		_w9069_,
		_w9098_,
		_w9630_,
		_w9631_
	);
	LUT2 #(
		.INIT('h8)
	) name7882 (
		rst_i_pad,
		\u4_u1_ienb_reg[5]/P0001 ,
		_w9632_
	);
	LUT4 #(
		.INIT('h5f08)
	) name7883 (
		_w2260_,
		_w9069_,
		_w9101_,
		_w9632_,
		_w9633_
	);
	LUT3 #(
		.INIT('h20)
	) name7884 (
		rst_i_pad,
		\u4_u1_int_re_reg/P0001 ,
		\u4_u1_int_stat_reg[1]/P0001 ,
		_w9634_
	);
	LUT3 #(
		.INIT('hd0)
	) name7885 (
		\u0_rx_active_reg/P0001 ,
		\u0_rx_err_reg/P0001 ,
		\u4_u1_ep_match_r_reg/P0001 ,
		_w9635_
	);
	LUT3 #(
		.INIT('h80)
	) name7886 (
		_w3671_,
		_w3899_,
		_w9635_,
		_w9636_
	);
	LUT3 #(
		.INIT('hdc)
	) name7887 (
		_w3682_,
		_w9634_,
		_w9636_,
		_w9637_
	);
	LUT2 #(
		.INIT('h8)
	) name7888 (
		rst_i_pad,
		\u4_u1_ots_stop_reg/P0001 ,
		_w9638_
	);
	LUT4 #(
		.INIT('h7720)
	) name7889 (
		_w2260_,
		_w9108_,
		_w9110_,
		_w9638_,
		_w9639_
	);
	LUT3 #(
		.INIT('h2a)
	) name7890 (
		\u4_u2_buf0_orig_reg[0]/P0001 ,
		_w2232_,
		_w2267_,
		_w9640_
	);
	LUT2 #(
		.INIT('hd)
	) name7891 (
		_w7642_,
		_w9640_,
		_w9641_
	);
	LUT3 #(
		.INIT('h2a)
	) name7892 (
		\u4_u2_buf0_orig_reg[10]/P0001 ,
		_w2232_,
		_w2267_,
		_w9642_
	);
	LUT2 #(
		.INIT('hd)
	) name7893 (
		_w2290_,
		_w9642_,
		_w9643_
	);
	LUT3 #(
		.INIT('h2a)
	) name7894 (
		\u4_u2_buf0_orig_reg[11]/P0001 ,
		_w2232_,
		_w2267_,
		_w9644_
	);
	LUT2 #(
		.INIT('hd)
	) name7895 (
		_w2456_,
		_w9644_,
		_w9645_
	);
	LUT3 #(
		.INIT('h2a)
	) name7896 (
		\u4_u2_buf0_orig_reg[12]/P0001 ,
		_w2232_,
		_w2267_,
		_w9646_
	);
	LUT2 #(
		.INIT('hd)
	) name7897 (
		_w7647_,
		_w9646_,
		_w9647_
	);
	LUT3 #(
		.INIT('h2a)
	) name7898 (
		\u4_u2_buf0_orig_reg[13]/P0001 ,
		_w2232_,
		_w2267_,
		_w9648_
	);
	LUT2 #(
		.INIT('hd)
	) name7899 (
		_w2361_,
		_w9648_,
		_w9649_
	);
	LUT3 #(
		.INIT('h2a)
	) name7900 (
		\u4_u2_buf0_orig_reg[14]/P0001 ,
		_w2232_,
		_w2267_,
		_w9650_
	);
	LUT2 #(
		.INIT('hd)
	) name7901 (
		_w2268_,
		_w9650_,
		_w9651_
	);
	LUT3 #(
		.INIT('h2a)
	) name7902 (
		\u4_u2_buf0_orig_reg[15]/P0001 ,
		_w2232_,
		_w2267_,
		_w9652_
	);
	LUT2 #(
		.INIT('hd)
	) name7903 (
		_w2461_,
		_w9652_,
		_w9653_
	);
	LUT3 #(
		.INIT('h2a)
	) name7904 (
		\u4_u2_buf0_orig_reg[16]/P0001 ,
		_w2232_,
		_w2267_,
		_w9654_
	);
	LUT2 #(
		.INIT('hd)
	) name7905 (
		_w7652_,
		_w9654_,
		_w9655_
	);
	LUT3 #(
		.INIT('h2a)
	) name7906 (
		\u4_u2_buf0_orig_reg[17]/P0001 ,
		_w2232_,
		_w2267_,
		_w9656_
	);
	LUT2 #(
		.INIT('hd)
	) name7907 (
		_w7657_,
		_w9656_,
		_w9657_
	);
	LUT3 #(
		.INIT('h2a)
	) name7908 (
		\u4_u2_buf0_orig_reg[18]/P0001 ,
		_w2232_,
		_w2267_,
		_w9658_
	);
	LUT2 #(
		.INIT('hd)
	) name7909 (
		_w7662_,
		_w9658_,
		_w9659_
	);
	LUT3 #(
		.INIT('h2a)
	) name7910 (
		\u4_u2_buf0_orig_reg[19]/P0001 ,
		_w2232_,
		_w2267_,
		_w9660_
	);
	LUT2 #(
		.INIT('hd)
	) name7911 (
		_w7667_,
		_w9660_,
		_w9661_
	);
	LUT3 #(
		.INIT('h2a)
	) name7912 (
		\u4_u2_buf0_orig_reg[1]/P0001 ,
		_w2232_,
		_w2267_,
		_w9662_
	);
	LUT2 #(
		.INIT('hd)
	) name7913 (
		_w7672_,
		_w9662_,
		_w9663_
	);
	LUT3 #(
		.INIT('h2a)
	) name7914 (
		\u4_u2_buf0_orig_reg[20]/P0001 ,
		_w2232_,
		_w2267_,
		_w9664_
	);
	LUT2 #(
		.INIT('hd)
	) name7915 (
		_w7677_,
		_w9664_,
		_w9665_
	);
	LUT3 #(
		.INIT('h2a)
	) name7916 (
		\u4_u2_buf0_orig_reg[21]/P0001 ,
		_w2232_,
		_w2267_,
		_w9666_
	);
	LUT2 #(
		.INIT('hd)
	) name7917 (
		_w7682_,
		_w9666_,
		_w9667_
	);
	LUT3 #(
		.INIT('h2a)
	) name7918 (
		\u4_u2_buf0_orig_reg[22]/P0001 ,
		_w2232_,
		_w2267_,
		_w9668_
	);
	LUT2 #(
		.INIT('hd)
	) name7919 (
		_w7687_,
		_w9668_,
		_w9669_
	);
	LUT3 #(
		.INIT('h2a)
	) name7920 (
		\u4_u2_buf0_orig_reg[23]/P0001 ,
		_w2232_,
		_w2267_,
		_w9670_
	);
	LUT2 #(
		.INIT('hd)
	) name7921 (
		_w7692_,
		_w9670_,
		_w9671_
	);
	LUT3 #(
		.INIT('h2a)
	) name7922 (
		\u4_u2_buf0_orig_reg[24]/P0001 ,
		_w2232_,
		_w2267_,
		_w9672_
	);
	LUT2 #(
		.INIT('hd)
	) name7923 (
		_w7697_,
		_w9672_,
		_w9673_
	);
	LUT3 #(
		.INIT('h2a)
	) name7924 (
		\u4_u2_buf0_orig_reg[25]/P0001 ,
		_w2232_,
		_w2267_,
		_w9674_
	);
	LUT2 #(
		.INIT('hd)
	) name7925 (
		_w7702_,
		_w9674_,
		_w9675_
	);
	LUT3 #(
		.INIT('h2a)
	) name7926 (
		\u4_u2_buf0_orig_reg[26]/P0001 ,
		_w2232_,
		_w2267_,
		_w9676_
	);
	LUT2 #(
		.INIT('hd)
	) name7927 (
		_w7707_,
		_w9676_,
		_w9677_
	);
	LUT3 #(
		.INIT('h2a)
	) name7928 (
		\u4_u2_buf0_orig_reg[27]/P0001 ,
		_w2232_,
		_w2267_,
		_w9678_
	);
	LUT2 #(
		.INIT('hd)
	) name7929 (
		_w7712_,
		_w9678_,
		_w9679_
	);
	LUT3 #(
		.INIT('h2a)
	) name7930 (
		\u4_u2_buf0_orig_reg[28]/P0001 ,
		_w2232_,
		_w2267_,
		_w9680_
	);
	LUT2 #(
		.INIT('hd)
	) name7931 (
		_w7717_,
		_w9680_,
		_w9681_
	);
	LUT3 #(
		.INIT('h2a)
	) name7932 (
		\u4_u2_buf0_orig_reg[29]/NET0131 ,
		_w2232_,
		_w2267_,
		_w9682_
	);
	LUT2 #(
		.INIT('hd)
	) name7933 (
		_w7722_,
		_w9682_,
		_w9683_
	);
	LUT3 #(
		.INIT('h2a)
	) name7934 (
		\u4_u2_buf0_orig_reg[2]/P0001 ,
		_w2232_,
		_w2267_,
		_w9684_
	);
	LUT2 #(
		.INIT('hd)
	) name7935 (
		_w7727_,
		_w9684_,
		_w9685_
	);
	LUT3 #(
		.INIT('h2a)
	) name7936 (
		\u4_u2_buf0_orig_reg[30]/NET0131 ,
		_w2232_,
		_w2267_,
		_w9686_
	);
	LUT2 #(
		.INIT('hd)
	) name7937 (
		_w7732_,
		_w9686_,
		_w9687_
	);
	LUT3 #(
		.INIT('h2a)
	) name7938 (
		\u4_u2_buf0_orig_reg[31]/P0001 ,
		_w2232_,
		_w2267_,
		_w9688_
	);
	LUT2 #(
		.INIT('hd)
	) name7939 (
		_w7737_,
		_w9688_,
		_w9689_
	);
	LUT3 #(
		.INIT('h2a)
	) name7940 (
		\u4_u2_buf0_orig_reg[3]/P0001 ,
		_w2232_,
		_w2267_,
		_w9690_
	);
	LUT2 #(
		.INIT('hd)
	) name7941 (
		_w7742_,
		_w9690_,
		_w9691_
	);
	LUT3 #(
		.INIT('h2a)
	) name7942 (
		\u4_u2_buf0_orig_reg[4]/P0001 ,
		_w2232_,
		_w2267_,
		_w9692_
	);
	LUT2 #(
		.INIT('hd)
	) name7943 (
		_w2611_,
		_w9692_,
		_w9693_
	);
	LUT3 #(
		.INIT('h2a)
	) name7944 (
		\u4_u2_buf0_orig_reg[5]/P0001 ,
		_w2232_,
		_w2267_,
		_w9694_
	);
	LUT2 #(
		.INIT('hd)
	) name7945 (
		_w2616_,
		_w9694_,
		_w9695_
	);
	LUT3 #(
		.INIT('h2a)
	) name7946 (
		\u4_u2_buf0_orig_reg[6]/P0001 ,
		_w2232_,
		_w2267_,
		_w9696_
	);
	LUT2 #(
		.INIT('hd)
	) name7947 (
		_w2472_,
		_w9696_,
		_w9697_
	);
	LUT3 #(
		.INIT('h2a)
	) name7948 (
		\u4_u2_buf0_orig_reg[7]/P0001 ,
		_w2232_,
		_w2267_,
		_w9698_
	);
	LUT2 #(
		.INIT('hd)
	) name7949 (
		_w2621_,
		_w9698_,
		_w9699_
	);
	LUT3 #(
		.INIT('h2a)
	) name7950 (
		\u4_u2_buf0_orig_reg[8]/P0001 ,
		_w2232_,
		_w2267_,
		_w9700_
	);
	LUT2 #(
		.INIT('hd)
	) name7951 (
		_w7747_,
		_w9700_,
		_w9701_
	);
	LUT3 #(
		.INIT('h2a)
	) name7952 (
		\u4_u2_buf0_orig_reg[9]/P0001 ,
		_w2232_,
		_w2267_,
		_w9702_
	);
	LUT2 #(
		.INIT('hd)
	) name7953 (
		_w7752_,
		_w9702_,
		_w9703_
	);
	LUT2 #(
		.INIT('h8)
	) name7954 (
		rst_i_pad,
		\u4_u2_csr0_reg[0]/P0001 ,
		_w9704_
	);
	LUT4 #(
		.INIT('h5f08)
	) name7955 (
		_w2267_,
		_w9110_,
		_w9173_,
		_w9704_,
		_w9705_
	);
	LUT2 #(
		.INIT('h8)
	) name7956 (
		rst_i_pad,
		\u4_u2_csr0_reg[10]/P0001 ,
		_w9706_
	);
	LUT4 #(
		.INIT('h5f08)
	) name7957 (
		_w2267_,
		_w9110_,
		_w9176_,
		_w9706_,
		_w9707_
	);
	LUT2 #(
		.INIT('h8)
	) name7958 (
		rst_i_pad,
		\u4_u2_csr0_reg[11]/P0001 ,
		_w9708_
	);
	LUT4 #(
		.INIT('h5f08)
	) name7959 (
		_w2267_,
		_w9110_,
		_w9179_,
		_w9708_,
		_w9709_
	);
	LUT2 #(
		.INIT('h8)
	) name7960 (
		rst_i_pad,
		\u4_u2_csr0_reg[12]/P0001 ,
		_w9710_
	);
	LUT4 #(
		.INIT('h5f08)
	) name7961 (
		_w2267_,
		_w9110_,
		_w9182_,
		_w9710_,
		_w9711_
	);
	LUT2 #(
		.INIT('h8)
	) name7962 (
		rst_i_pad,
		\u4_u2_csr0_reg[1]/P0001 ,
		_w9712_
	);
	LUT4 #(
		.INIT('h5f08)
	) name7963 (
		_w2267_,
		_w9110_,
		_w9185_,
		_w9712_,
		_w9713_
	);
	LUT2 #(
		.INIT('h8)
	) name7964 (
		rst_i_pad,
		\u4_u2_csr0_reg[2]/P0001 ,
		_w9714_
	);
	LUT4 #(
		.INIT('h5f08)
	) name7965 (
		_w2267_,
		_w9110_,
		_w9188_,
		_w9714_,
		_w9715_
	);
	LUT2 #(
		.INIT('h8)
	) name7966 (
		rst_i_pad,
		\u4_u2_csr0_reg[3]/NET0131 ,
		_w9716_
	);
	LUT4 #(
		.INIT('h5f08)
	) name7967 (
		_w2267_,
		_w9110_,
		_w9191_,
		_w9716_,
		_w9717_
	);
	LUT2 #(
		.INIT('h8)
	) name7968 (
		rst_i_pad,
		\u4_u2_csr0_reg[4]/P0001 ,
		_w9718_
	);
	LUT4 #(
		.INIT('h5f08)
	) name7969 (
		_w2267_,
		_w9110_,
		_w9194_,
		_w9718_,
		_w9719_
	);
	LUT2 #(
		.INIT('h8)
	) name7970 (
		rst_i_pad,
		\u4_u2_csr0_reg[5]/P0001 ,
		_w9720_
	);
	LUT4 #(
		.INIT('h5f08)
	) name7971 (
		_w2267_,
		_w9110_,
		_w9197_,
		_w9720_,
		_w9721_
	);
	LUT2 #(
		.INIT('h8)
	) name7972 (
		rst_i_pad,
		\u4_u2_csr0_reg[6]/P0001 ,
		_w9722_
	);
	LUT4 #(
		.INIT('h5f08)
	) name7973 (
		_w2267_,
		_w9110_,
		_w9200_,
		_w9722_,
		_w9723_
	);
	LUT2 #(
		.INIT('h8)
	) name7974 (
		rst_i_pad,
		\u4_u2_csr0_reg[7]/P0001 ,
		_w9724_
	);
	LUT4 #(
		.INIT('h5f08)
	) name7975 (
		_w2267_,
		_w9110_,
		_w9203_,
		_w9724_,
		_w9725_
	);
	LUT2 #(
		.INIT('h8)
	) name7976 (
		rst_i_pad,
		\u4_u2_csr0_reg[8]/P0001 ,
		_w9726_
	);
	LUT4 #(
		.INIT('h5f08)
	) name7977 (
		_w2267_,
		_w9110_,
		_w9206_,
		_w9726_,
		_w9727_
	);
	LUT2 #(
		.INIT('h8)
	) name7978 (
		rst_i_pad,
		\u4_u2_csr0_reg[9]/P0001 ,
		_w9728_
	);
	LUT4 #(
		.INIT('h5f08)
	) name7979 (
		_w2267_,
		_w9110_,
		_w9209_,
		_w9728_,
		_w9729_
	);
	LUT2 #(
		.INIT('h8)
	) name7980 (
		rst_i_pad,
		\u4_u2_csr1_reg[10]/P0001 ,
		_w9730_
	);
	LUT4 #(
		.INIT('h5f08)
	) name7981 (
		_w2267_,
		_w9110_,
		_w9214_,
		_w9730_,
		_w9731_
	);
	LUT2 #(
		.INIT('h8)
	) name7982 (
		rst_i_pad,
		\u4_u2_csr1_reg[11]/P0001 ,
		_w9732_
	);
	LUT4 #(
		.INIT('h5f08)
	) name7983 (
		_w2267_,
		_w9110_,
		_w9217_,
		_w9732_,
		_w9733_
	);
	LUT2 #(
		.INIT('h8)
	) name7984 (
		rst_i_pad,
		\u4_u2_csr1_reg[12]/P0001 ,
		_w9734_
	);
	LUT4 #(
		.INIT('h5f08)
	) name7985 (
		_w2267_,
		_w9110_,
		_w9220_,
		_w9734_,
		_w9735_
	);
	LUT2 #(
		.INIT('h8)
	) name7986 (
		rst_i_pad,
		\u4_u2_csr1_reg[1]/P0001 ,
		_w9736_
	);
	LUT4 #(
		.INIT('h5f08)
	) name7987 (
		_w2267_,
		_w9110_,
		_w9223_,
		_w9736_,
		_w9737_
	);
	LUT2 #(
		.INIT('h8)
	) name7988 (
		rst_i_pad,
		\u4_u2_csr1_reg[2]/P0001 ,
		_w9738_
	);
	LUT4 #(
		.INIT('h5f08)
	) name7989 (
		_w2267_,
		_w9110_,
		_w9226_,
		_w9738_,
		_w9739_
	);
	LUT2 #(
		.INIT('h8)
	) name7990 (
		rst_i_pad,
		\u4_u2_csr1_reg[3]/P0001 ,
		_w9740_
	);
	LUT4 #(
		.INIT('h5f08)
	) name7991 (
		_w2267_,
		_w9110_,
		_w9229_,
		_w9740_,
		_w9741_
	);
	LUT2 #(
		.INIT('h8)
	) name7992 (
		rst_i_pad,
		\u4_u2_csr1_reg[4]/P0001 ,
		_w9742_
	);
	LUT4 #(
		.INIT('h5f08)
	) name7993 (
		_w2267_,
		_w9110_,
		_w9232_,
		_w9742_,
		_w9743_
	);
	LUT2 #(
		.INIT('h8)
	) name7994 (
		rst_i_pad,
		\u4_u2_csr1_reg[5]/P0001 ,
		_w9744_
	);
	LUT4 #(
		.INIT('h5f08)
	) name7995 (
		_w2267_,
		_w9110_,
		_w9235_,
		_w9744_,
		_w9745_
	);
	LUT2 #(
		.INIT('h8)
	) name7996 (
		rst_i_pad,
		\u4_u2_csr1_reg[6]/P0001 ,
		_w9746_
	);
	LUT4 #(
		.INIT('h5f08)
	) name7997 (
		_w2267_,
		_w9110_,
		_w9238_,
		_w9746_,
		_w9747_
	);
	LUT2 #(
		.INIT('h8)
	) name7998 (
		rst_i_pad,
		\u4_u2_csr1_reg[9]/P0001 ,
		_w9748_
	);
	LUT4 #(
		.INIT('h5f08)
	) name7999 (
		_w2267_,
		_w9110_,
		_w9241_,
		_w9748_,
		_w9749_
	);
	LUT4 #(
		.INIT('h0080)
	) name8000 (
		_w5201_,
		_w5203_,
		_w5211_,
		_w5214_,
		_w9750_
	);
	LUT3 #(
		.INIT('h80)
	) name8001 (
		_w5197_,
		_w5206_,
		_w5215_,
		_w9751_
	);
	LUT4 #(
		.INIT('h8000)
	) name8002 (
		_w5237_,
		_w5239_,
		_w9750_,
		_w9751_,
		_w9752_
	);
	LUT4 #(
		.INIT('h0800)
	) name8003 (
		\u1_u3_state_reg[9]/P0001 ,
		\u4_csr_reg[15]/NET0131 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		_w9753_
	);
	LUT2 #(
		.INIT('h4)
	) name8004 (
		_w9752_,
		_w9753_,
		_w9754_
	);
	LUT4 #(
		.INIT('hdf00)
	) name8005 (
		\LineState_r_reg[0]/P0001 ,
		\LineState_r_reg[1]/P0001 ,
		\u0_u0_ls_j_r_reg/P0001 ,
		\u0_u0_state_reg[14]/P0001 ,
		_w9755_
	);
	LUT2 #(
		.INIT('h1)
	) name8006 (
		_w4117_,
		_w9755_,
		_w9756_
	);
	LUT4 #(
		.INIT('hbf00)
	) name8007 (
		\LineState_r_reg[0]/P0001 ,
		\LineState_r_reg[1]/P0001 ,
		\u0_u0_ls_k_r_reg/P0001 ,
		\u0_u0_state_reg[14]/P0001 ,
		_w9757_
	);
	LUT2 #(
		.INIT('h1)
	) name8008 (
		_w4117_,
		_w9757_,
		_w9758_
	);
	LUT4 #(
		.INIT('hf531)
	) name8009 (
		_w8984_,
		_w8991_,
		_w9756_,
		_w9758_,
		_w9759_
	);
	LUT2 #(
		.INIT('h2)
	) name8010 (
		_w4122_,
		_w9759_,
		_w9760_
	);
	LUT3 #(
		.INIT('h07)
	) name8011 (
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u2_ep_match_r_reg/P0001 ,
		\u4_u2_int_stat_reg[6]/P0001 ,
		_w9761_
	);
	LUT2 #(
		.INIT('h2)
	) name8012 (
		_w3890_,
		_w9761_,
		_w9762_
	);
	LUT3 #(
		.INIT('h07)
	) name8013 (
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u0_ep_match_r_reg/P0001 ,
		\u4_u0_int_stat_reg[6]/P0001 ,
		_w9763_
	);
	LUT2 #(
		.INIT('h2)
	) name8014 (
		_w3896_,
		_w9763_,
		_w9764_
	);
	LUT3 #(
		.INIT('h07)
	) name8015 (
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u1_ep_match_r_reg/P0001 ,
		\u4_u1_int_stat_reg[6]/P0001 ,
		_w9765_
	);
	LUT2 #(
		.INIT('h2)
	) name8016 (
		_w3899_,
		_w9765_,
		_w9766_
	);
	LUT4 #(
		.INIT('h20a0)
	) name8017 (
		rst_i_pad,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u0_csr1_reg[8]/P0001 ,
		\u4_u0_ots_stop_reg/P0001 ,
		_w9767_
	);
	LUT2 #(
		.INIT('h8)
	) name8018 (
		rst_i_pad,
		\wb_data_i[23]_pad ,
		_w9768_
	);
	LUT4 #(
		.INIT('hf870)
	) name8019 (
		_w2243_,
		_w5840_,
		_w9767_,
		_w9768_,
		_w9769_
	);
	LUT2 #(
		.INIT('h2)
	) name8020 (
		\u0_u0_state_reg[3]/P0001 ,
		_w4354_,
		_w9770_
	);
	LUT3 #(
		.INIT('hb0)
	) name8021 (
		\u0_u0_usb_suspend_reg/P0001 ,
		_w5768_,
		_w9770_,
		_w9771_
	);
	LUT4 #(
		.INIT('h0110)
	) name8022 (
		\u0_u0_state_reg[1]/P0001 ,
		\u0_u0_state_reg[2]/NET0131 ,
		\u0_u0_state_reg[4]/NET0131 ,
		\u0_u0_state_reg[5]/P0001 ,
		_w9772_
	);
	LUT4 #(
		.INIT('h8000)
	) name8023 (
		_w4109_,
		_w7789_,
		_w7793_,
		_w9772_,
		_w9773_
	);
	LUT2 #(
		.INIT('h1)
	) name8024 (
		\u0_u0_state_reg[3]/P0001 ,
		_w9773_,
		_w9774_
	);
	LUT3 #(
		.INIT('h23)
	) name8025 (
		\u0_u0_usb_suspend_reg/P0001 ,
		_w4333_,
		_w5768_,
		_w9775_
	);
	LUT3 #(
		.INIT('hea)
	) name8026 (
		_w9771_,
		_w9774_,
		_w9775_,
		_w9776_
	);
	LUT4 #(
		.INIT('h20a0)
	) name8027 (
		rst_i_pad,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u2_csr1_reg[8]/P0001 ,
		\u4_u2_ots_stop_reg/P0001 ,
		_w9777_
	);
	LUT4 #(
		.INIT('hf780)
	) name8028 (
		_w2267_,
		_w5840_,
		_w9768_,
		_w9777_,
		_w9778_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name8029 (
		\u4_u0_buf1_reg[4]/P0001 ,
		\u4_u0_csr0_reg[4]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w9779_
	);
	LUT4 #(
		.INIT('hf53f)
	) name8030 (
		\u4_u0_buf0_reg[4]/P0001 ,
		\u4_u0_int_stat_reg[4]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w9780_
	);
	LUT4 #(
		.INIT('h0888)
	) name8031 (
		_w2240_,
		_w2241_,
		_w9779_,
		_w9780_,
		_w9781_
	);
	LUT4 #(
		.INIT('hf5f3)
	) name8032 (
		\u4_u2_buf0_reg[4]/P0001 ,
		\u4_u2_csr0_reg[4]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w9782_
	);
	LUT4 #(
		.INIT('h5f3f)
	) name8033 (
		\u4_u2_buf1_reg[4]/P0001 ,
		\u4_u2_int_stat_reg[4]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w9783_
	);
	LUT4 #(
		.INIT('h0888)
	) name8034 (
		_w2228_,
		_w2240_,
		_w9782_,
		_w9783_,
		_w9784_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name8035 (
		\u4_u3_buf1_reg[4]/P0001 ,
		\u4_u3_csr0_reg[4]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w9785_
	);
	LUT4 #(
		.INIT('hf53f)
	) name8036 (
		\u4_u3_buf0_reg[4]/P0001 ,
		\u4_u3_int_stat_reg[4]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w9786_
	);
	LUT4 #(
		.INIT('h0888)
	) name8037 (
		_w2227_,
		_w2228_,
		_w9785_,
		_w9786_,
		_w9787_
	);
	LUT3 #(
		.INIT('h01)
	) name8038 (
		_w9781_,
		_w9784_,
		_w9787_,
		_w9788_
	);
	LUT4 #(
		.INIT('h0008)
	) name8039 (
		\u4_funct_adr_reg[4]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w9789_
	);
	LUT4 #(
		.INIT('h0020)
	) name8040 (
		\u4_inta_msk_reg[4]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w9790_
	);
	LUT2 #(
		.INIT('h1)
	) name8041 (
		_w9789_,
		_w9790_,
		_w9791_
	);
	LUT4 #(
		.INIT('h0002)
	) name8042 (
		\LineState_r_reg[1]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w9792_
	);
	LUT4 #(
		.INIT('h0800)
	) name8043 (
		\u4_utmi_vend_stat_r_reg[4]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w9793_
	);
	LUT4 #(
		.INIT('h0200)
	) name8044 (
		\u1_sof_time_reg[4]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w9794_
	);
	LUT3 #(
		.INIT('h01)
	) name8045 (
		_w9792_,
		_w9793_,
		_w9794_,
		_w9795_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name8046 (
		\u4_u1_buf1_reg[4]/P0001 ,
		\u4_u1_csr0_reg[4]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w9796_
	);
	LUT4 #(
		.INIT('hf53f)
	) name8047 (
		\u4_u1_buf0_reg[4]/P0001 ,
		\u4_u1_int_stat_reg[4]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w9797_
	);
	LUT4 #(
		.INIT('h0888)
	) name8048 (
		_w2227_,
		_w2241_,
		_w9796_,
		_w9797_,
		_w9798_
	);
	LUT4 #(
		.INIT('h00d5)
	) name8049 (
		_w5861_,
		_w9791_,
		_w9795_,
		_w9798_,
		_w9799_
	);
	LUT2 #(
		.INIT('h7)
	) name8050 (
		_w9788_,
		_w9799_,
		_w9800_
	);
	LUT4 #(
		.INIT('h20a0)
	) name8051 (
		rst_i_pad,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u3_csr1_reg[8]/P0001 ,
		\u4_u3_ots_stop_reg/P0001 ,
		_w9801_
	);
	LUT4 #(
		.INIT('hf780)
	) name8052 (
		_w2231_,
		_w5840_,
		_w9768_,
		_w9801_,
		_w9802_
	);
	LUT4 #(
		.INIT('h8000)
	) name8053 (
		\u0_u0_idle_cnt1_reg[4]/P0001 ,
		\u0_u0_idle_cnt1_reg[5]/P0001 ,
		\u0_u0_idle_cnt1_reg[6]/P0001 ,
		\u0_u0_idle_cnt1_reg[7]/P0001 ,
		_w9803_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name8054 (
		\u0_u0_idle_cnt1_reg[6]/P0001 ,
		\u0_u0_idle_cnt1_reg[7]/P0001 ,
		_w8152_,
		_w9015_,
		_w9804_
	);
	LUT4 #(
		.INIT('h20a0)
	) name8055 (
		rst_i_pad,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u1_csr1_reg[8]/P0001 ,
		\u4_u1_ots_stop_reg/P0001 ,
		_w9805_
	);
	LUT4 #(
		.INIT('hf780)
	) name8056 (
		_w2260_,
		_w5840_,
		_w9768_,
		_w9805_,
		_w9806_
	);
	LUT2 #(
		.INIT('h8)
	) name8057 (
		rst_i_pad,
		\wb_data_i[22]_pad ,
		_w9807_
	);
	LUT4 #(
		.INIT('ha8a0)
	) name8058 (
		rst_i_pad,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u3_csr1_reg[7]/P0001 ,
		\u4_u3_ots_stop_reg/P0001 ,
		_w9808_
	);
	LUT4 #(
		.INIT('hf780)
	) name8059 (
		_w2231_,
		_w5840_,
		_w9807_,
		_w9808_,
		_w9809_
	);
	LUT4 #(
		.INIT('ha8a0)
	) name8060 (
		rst_i_pad,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u0_csr1_reg[7]/P0001 ,
		\u4_u0_ots_stop_reg/P0001 ,
		_w9810_
	);
	LUT4 #(
		.INIT('hf780)
	) name8061 (
		_w2243_,
		_w5840_,
		_w9807_,
		_w9810_,
		_w9811_
	);
	LUT4 #(
		.INIT('ha8a0)
	) name8062 (
		rst_i_pad,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u1_csr1_reg[7]/P0001 ,
		\u4_u1_ots_stop_reg/P0001 ,
		_w9812_
	);
	LUT4 #(
		.INIT('hf780)
	) name8063 (
		_w2260_,
		_w5840_,
		_w9807_,
		_w9812_,
		_w9813_
	);
	LUT4 #(
		.INIT('ha8a0)
	) name8064 (
		rst_i_pad,
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u2_csr1_reg[7]/P0001 ,
		\u4_u2_ots_stop_reg/P0001 ,
		_w9814_
	);
	LUT4 #(
		.INIT('hf780)
	) name8065 (
		_w2267_,
		_w5840_,
		_w9807_,
		_w9814_,
		_w9815_
	);
	LUT3 #(
		.INIT('hac)
	) name8066 (
		\sram_data_i[12]_pad ,
		\u4_dout_reg[12]/P0001 ,
		\wb_addr_i[17]_pad ,
		_w9816_
	);
	LUT3 #(
		.INIT('hac)
	) name8067 (
		\sram_data_i[13]_pad ,
		\u4_dout_reg[13]/P0001 ,
		\wb_addr_i[17]_pad ,
		_w9817_
	);
	LUT3 #(
		.INIT('hac)
	) name8068 (
		\sram_data_i[15]_pad ,
		\u4_dout_reg[15]/P0001 ,
		\wb_addr_i[17]_pad ,
		_w9818_
	);
	LUT3 #(
		.INIT('h40)
	) name8069 (
		VControl_Load_pad_o_pad,
		rst_i_pad,
		\u4_utmi_vend_wr_r_reg/P0001 ,
		_w9819_
	);
	LUT4 #(
		.INIT('h0800)
	) name8070 (
		rst_i_pad,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w9820_
	);
	LUT3 #(
		.INIT('hec)
	) name8071 (
		_w8842_,
		_w9819_,
		_w9820_,
		_w9821_
	);
	LUT3 #(
		.INIT('hed)
	) name8072 (
		\LineState_r_reg[0]/P0001 ,
		\LineState_r_reg[1]/P0001 ,
		\u0_u0_mode_hs_reg/P0001 ,
		_w9822_
	);
	LUT3 #(
		.INIT('h12)
	) name8073 (
		\LineState_r_reg[0]/P0001 ,
		\LineState_r_reg[1]/P0001 ,
		\u0_u0_mode_hs_reg/P0001 ,
		_w9823_
	);
	LUT2 #(
		.INIT('h8)
	) name8074 (
		\u0_u0_idle_long_reg/P0001 ,
		\u0_u0_ls_idle_r_reg/P0001 ,
		_w9824_
	);
	LUT3 #(
		.INIT('ha8)
	) name8075 (
		rst_i_pad,
		\u0_u0_idle_long_reg/P0001 ,
		\u0_u0_ls_idle_r_reg/P0001 ,
		_w9825_
	);
	LUT3 #(
		.INIT('hd0)
	) name8076 (
		_w9822_,
		_w9824_,
		_w9825_,
		_w9826_
	);
	LUT3 #(
		.INIT('h02)
	) name8077 (
		\u4_u0_uc_bsel_reg[1]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w9827_
	);
	LUT4 #(
		.INIT('h35ff)
	) name8078 (
		\u4_u0_buf0_reg[31]/P0001 ,
		\u4_u0_buf1_reg[31]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w9828_
	);
	LUT4 #(
		.INIT('h8088)
	) name8079 (
		_w2240_,
		_w2241_,
		_w9827_,
		_w9828_,
		_w9829_
	);
	LUT3 #(
		.INIT('h02)
	) name8080 (
		\u4_u1_uc_bsel_reg[1]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w9830_
	);
	LUT4 #(
		.INIT('h35ff)
	) name8081 (
		\u4_u1_buf0_reg[31]/P0001 ,
		\u4_u1_buf1_reg[31]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w9831_
	);
	LUT4 #(
		.INIT('h8088)
	) name8082 (
		_w2227_,
		_w2241_,
		_w9830_,
		_w9831_,
		_w9832_
	);
	LUT2 #(
		.INIT('h1)
	) name8083 (
		_w9829_,
		_w9832_,
		_w9833_
	);
	LUT4 #(
		.INIT('h0200)
	) name8084 (
		\u1_mfm_cnt_reg[3]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w9834_
	);
	LUT2 #(
		.INIT('h8)
	) name8085 (
		_w5861_,
		_w9834_,
		_w9835_
	);
	LUT3 #(
		.INIT('h02)
	) name8086 (
		\u4_u3_uc_bsel_reg[1]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w9836_
	);
	LUT4 #(
		.INIT('h35ff)
	) name8087 (
		\u4_u3_buf0_reg[31]/P0001 ,
		\u4_u3_buf1_reg[31]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w9837_
	);
	LUT4 #(
		.INIT('h8088)
	) name8088 (
		_w2227_,
		_w2228_,
		_w9836_,
		_w9837_,
		_w9838_
	);
	LUT3 #(
		.INIT('h02)
	) name8089 (
		\u4_u2_uc_bsel_reg[1]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w9839_
	);
	LUT4 #(
		.INIT('h35ff)
	) name8090 (
		\u4_u2_buf0_reg[31]/P0001 ,
		\u4_u2_buf1_reg[31]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w9840_
	);
	LUT4 #(
		.INIT('h8088)
	) name8091 (
		_w2228_,
		_w2240_,
		_w9839_,
		_w9840_,
		_w9841_
	);
	LUT3 #(
		.INIT('h01)
	) name8092 (
		_w9835_,
		_w9838_,
		_w9841_,
		_w9842_
	);
	LUT2 #(
		.INIT('h7)
	) name8093 (
		_w9833_,
		_w9842_,
		_w9843_
	);
	LUT3 #(
		.INIT('h02)
	) name8094 (
		\u4_u0_uc_bsel_reg[0]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w9844_
	);
	LUT4 #(
		.INIT('h35ff)
	) name8095 (
		\u4_u0_buf0_reg[30]/P0001 ,
		\u4_u0_buf1_reg[30]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w9845_
	);
	LUT4 #(
		.INIT('h8088)
	) name8096 (
		_w2240_,
		_w2241_,
		_w9844_,
		_w9845_,
		_w9846_
	);
	LUT3 #(
		.INIT('h02)
	) name8097 (
		\u4_u1_uc_bsel_reg[0]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w9847_
	);
	LUT4 #(
		.INIT('h35ff)
	) name8098 (
		\u4_u1_buf0_reg[30]/P0001 ,
		\u4_u1_buf1_reg[30]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w9848_
	);
	LUT4 #(
		.INIT('h8088)
	) name8099 (
		_w2227_,
		_w2241_,
		_w9847_,
		_w9848_,
		_w9849_
	);
	LUT2 #(
		.INIT('h1)
	) name8100 (
		_w9846_,
		_w9849_,
		_w9850_
	);
	LUT4 #(
		.INIT('h0200)
	) name8101 (
		\u1_mfm_cnt_reg[2]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w9851_
	);
	LUT2 #(
		.INIT('h8)
	) name8102 (
		_w5861_,
		_w9851_,
		_w9852_
	);
	LUT3 #(
		.INIT('h02)
	) name8103 (
		\u4_u3_uc_bsel_reg[0]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w9853_
	);
	LUT4 #(
		.INIT('h35ff)
	) name8104 (
		\u4_u3_buf0_reg[30]/P0001 ,
		\u4_u3_buf1_reg[30]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w9854_
	);
	LUT4 #(
		.INIT('h8088)
	) name8105 (
		_w2227_,
		_w2228_,
		_w9853_,
		_w9854_,
		_w9855_
	);
	LUT3 #(
		.INIT('h02)
	) name8106 (
		\u4_u2_uc_bsel_reg[0]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w9856_
	);
	LUT4 #(
		.INIT('h35ff)
	) name8107 (
		\u4_u2_buf0_reg[30]/P0001 ,
		\u4_u2_buf1_reg[30]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w9857_
	);
	LUT4 #(
		.INIT('h8088)
	) name8108 (
		_w2228_,
		_w2240_,
		_w9856_,
		_w9857_,
		_w9858_
	);
	LUT3 #(
		.INIT('h01)
	) name8109 (
		_w9852_,
		_w9855_,
		_w9858_,
		_w9859_
	);
	LUT2 #(
		.INIT('h7)
	) name8110 (
		_w9850_,
		_w9859_,
		_w9860_
	);
	LUT4 #(
		.INIT('hf53f)
	) name8111 (
		\u4_u2_buf0_reg[29]/P0001 ,
		\u4_u2_iena_reg[5]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w9861_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name8112 (
		\u4_u2_buf1_reg[29]/P0001 ,
		\u4_u2_uc_dpd_reg[1]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w9862_
	);
	LUT4 #(
		.INIT('h0888)
	) name8113 (
		_w2228_,
		_w2240_,
		_w9861_,
		_w9862_,
		_w9863_
	);
	LUT4 #(
		.INIT('h5f3f)
	) name8114 (
		\u4_u0_buf1_reg[29]/P0001 ,
		\u4_u0_iena_reg[5]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w9864_
	);
	LUT4 #(
		.INIT('hf5f3)
	) name8115 (
		\u4_u0_buf0_reg[29]/P0001 ,
		\u4_u0_uc_dpd_reg[1]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w9865_
	);
	LUT4 #(
		.INIT('h0888)
	) name8116 (
		_w2240_,
		_w2241_,
		_w9864_,
		_w9865_,
		_w9866_
	);
	LUT2 #(
		.INIT('h1)
	) name8117 (
		_w9863_,
		_w9866_,
		_w9867_
	);
	LUT4 #(
		.INIT('h0200)
	) name8118 (
		\u1_mfm_cnt_reg[1]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w9868_
	);
	LUT2 #(
		.INIT('h8)
	) name8119 (
		_w5861_,
		_w9868_,
		_w9869_
	);
	LUT4 #(
		.INIT('hf5f3)
	) name8120 (
		\u4_u3_buf0_reg[29]/P0001 ,
		\u4_u3_uc_dpd_reg[1]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w9870_
	);
	LUT4 #(
		.INIT('h5f3f)
	) name8121 (
		\u4_u3_buf1_reg[29]/P0001 ,
		\u4_u3_iena_reg[5]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w9871_
	);
	LUT4 #(
		.INIT('h0888)
	) name8122 (
		_w2227_,
		_w2228_,
		_w9870_,
		_w9871_,
		_w9872_
	);
	LUT4 #(
		.INIT('h35ff)
	) name8123 (
		\u4_u1_buf0_reg[29]/P0001 ,
		\u4_u1_buf1_reg[29]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w9873_
	);
	LUT4 #(
		.INIT('hff53)
	) name8124 (
		\u4_u1_iena_reg[5]/P0001 ,
		\u4_u1_uc_dpd_reg[1]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w9874_
	);
	LUT4 #(
		.INIT('h0888)
	) name8125 (
		_w2227_,
		_w2241_,
		_w9873_,
		_w9874_,
		_w9875_
	);
	LUT3 #(
		.INIT('h01)
	) name8126 (
		_w9869_,
		_w9872_,
		_w9875_,
		_w9876_
	);
	LUT2 #(
		.INIT('h7)
	) name8127 (
		_w9867_,
		_w9876_,
		_w9877_
	);
	LUT4 #(
		.INIT('h2a00)
	) name8128 (
		rst_i_pad,
		\u1_u3_uc_bsel_set_reg/P0001 ,
		\u4_u2_ep_match_r_reg/P0001 ,
		\u4_u2_uc_bsel_reg[0]/P0001 ,
		_w9878_
	);
	LUT4 #(
		.INIT('h8000)
	) name8129 (
		rst_i_pad,
		\u1_u3_idin_reg[0]/P0001 ,
		\u1_u3_uc_bsel_set_reg/P0001 ,
		\u4_u2_ep_match_r_reg/P0001 ,
		_w9879_
	);
	LUT2 #(
		.INIT('he)
	) name8130 (
		_w9878_,
		_w9879_,
		_w9880_
	);
	LUT4 #(
		.INIT('h2a00)
	) name8131 (
		rst_i_pad,
		\u1_u3_uc_bsel_set_reg/P0001 ,
		\u4_u2_ep_match_r_reg/P0001 ,
		\u4_u2_uc_bsel_reg[1]/P0001 ,
		_w9881_
	);
	LUT4 #(
		.INIT('h8000)
	) name8132 (
		rst_i_pad,
		\u1_u3_idin_reg[1]/P0001 ,
		\u1_u3_uc_bsel_set_reg/P0001 ,
		\u4_u2_ep_match_r_reg/P0001 ,
		_w9882_
	);
	LUT2 #(
		.INIT('he)
	) name8133 (
		_w9881_,
		_w9882_,
		_w9883_
	);
	LUT4 #(
		.INIT('h2a00)
	) name8134 (
		rst_i_pad,
		\u1_u3_uc_bsel_set_reg/P0001 ,
		\u4_u2_ep_match_r_reg/P0001 ,
		\u4_u2_uc_dpd_reg[1]/P0001 ,
		_w9884_
	);
	LUT4 #(
		.INIT('h8000)
	) name8135 (
		rst_i_pad,
		\u1_u3_idin_reg[3]/P0001 ,
		\u1_u3_uc_bsel_set_reg/P0001 ,
		\u4_u2_ep_match_r_reg/P0001 ,
		_w9885_
	);
	LUT2 #(
		.INIT('he)
	) name8136 (
		_w9884_,
		_w9885_,
		_w9886_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name8137 (
		\u4_u3_buf1_reg[27]/P0001 ,
		\u4_u3_csr1_reg[12]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w9887_
	);
	LUT4 #(
		.INIT('hf53f)
	) name8138 (
		\u4_u3_buf0_reg[27]/P0001 ,
		\u4_u3_iena_reg[3]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w9888_
	);
	LUT4 #(
		.INIT('h0888)
	) name8139 (
		_w2227_,
		_w2228_,
		_w9887_,
		_w9888_,
		_w9889_
	);
	LUT4 #(
		.INIT('h5f3f)
	) name8140 (
		\u4_u2_buf1_reg[27]/P0001 ,
		\u4_u2_iena_reg[3]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w9890_
	);
	LUT4 #(
		.INIT('hf5f3)
	) name8141 (
		\u4_u2_buf0_reg[27]/P0001 ,
		\u4_u2_csr1_reg[12]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w9891_
	);
	LUT4 #(
		.INIT('h0888)
	) name8142 (
		_w2228_,
		_w2240_,
		_w9890_,
		_w9891_,
		_w9892_
	);
	LUT2 #(
		.INIT('h1)
	) name8143 (
		_w9889_,
		_w9892_,
		_w9893_
	);
	LUT4 #(
		.INIT('h0080)
	) name8144 (
		\u4_int_srcb_reg[7]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w9894_
	);
	LUT2 #(
		.INIT('h8)
	) name8145 (
		_w5861_,
		_w9894_,
		_w9895_
	);
	LUT4 #(
		.INIT('hf5f3)
	) name8146 (
		\u4_u1_buf0_reg[27]/P0001 ,
		\u4_u1_csr1_reg[12]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w9896_
	);
	LUT4 #(
		.INIT('h5f3f)
	) name8147 (
		\u4_u1_buf1_reg[27]/P0001 ,
		\u4_u1_iena_reg[3]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w9897_
	);
	LUT4 #(
		.INIT('h0888)
	) name8148 (
		_w2227_,
		_w2241_,
		_w9896_,
		_w9897_,
		_w9898_
	);
	LUT4 #(
		.INIT('h5f3f)
	) name8149 (
		\u4_u0_buf1_reg[27]/P0001 ,
		\u4_u0_iena_reg[3]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w9899_
	);
	LUT4 #(
		.INIT('hf5f3)
	) name8150 (
		\u4_u0_buf0_reg[27]/P0001 ,
		\u4_u0_csr1_reg[12]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w9900_
	);
	LUT4 #(
		.INIT('h0888)
	) name8151 (
		_w2240_,
		_w2241_,
		_w9899_,
		_w9900_,
		_w9901_
	);
	LUT3 #(
		.INIT('h01)
	) name8152 (
		_w9895_,
		_w9898_,
		_w9901_,
		_w9902_
	);
	LUT2 #(
		.INIT('h7)
	) name8153 (
		_w9893_,
		_w9902_,
		_w9903_
	);
	LUT4 #(
		.INIT('h2a00)
	) name8154 (
		rst_i_pad,
		\u1_u3_uc_bsel_set_reg/P0001 ,
		\u4_u3_ep_match_r_reg/P0001 ,
		\u4_u3_uc_bsel_reg[0]/P0001 ,
		_w9904_
	);
	LUT4 #(
		.INIT('h8000)
	) name8155 (
		rst_i_pad,
		\u1_u3_idin_reg[0]/P0001 ,
		\u1_u3_uc_bsel_set_reg/P0001 ,
		\u4_u3_ep_match_r_reg/P0001 ,
		_w9905_
	);
	LUT2 #(
		.INIT('he)
	) name8156 (
		_w9904_,
		_w9905_,
		_w9906_
	);
	LUT4 #(
		.INIT('h2a00)
	) name8157 (
		rst_i_pad,
		\u1_u3_uc_bsel_set_reg/P0001 ,
		\u4_u3_ep_match_r_reg/P0001 ,
		\u4_u3_uc_bsel_reg[1]/P0001 ,
		_w9907_
	);
	LUT4 #(
		.INIT('h8000)
	) name8158 (
		rst_i_pad,
		\u1_u3_idin_reg[1]/P0001 ,
		\u1_u3_uc_bsel_set_reg/P0001 ,
		\u4_u3_ep_match_r_reg/P0001 ,
		_w9908_
	);
	LUT2 #(
		.INIT('he)
	) name8159 (
		_w9907_,
		_w9908_,
		_w9909_
	);
	LUT4 #(
		.INIT('h2a00)
	) name8160 (
		rst_i_pad,
		\u1_u3_uc_bsel_set_reg/P0001 ,
		\u4_u3_ep_match_r_reg/P0001 ,
		\u4_u3_uc_dpd_reg[0]/P0001 ,
		_w9910_
	);
	LUT4 #(
		.INIT('h8000)
	) name8161 (
		rst_i_pad,
		\u1_u3_idin_reg[2]/P0001 ,
		\u1_u3_uc_bsel_set_reg/P0001 ,
		\u4_u3_ep_match_r_reg/P0001 ,
		_w9911_
	);
	LUT2 #(
		.INIT('he)
	) name8162 (
		_w9910_,
		_w9911_,
		_w9912_
	);
	LUT3 #(
		.INIT('h80)
	) name8163 (
		\u4_u1_buf1_reg[8]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w9913_
	);
	LUT4 #(
		.INIT('hf5f3)
	) name8164 (
		\u4_u1_buf0_reg[8]/P0001 ,
		\u4_u1_csr0_reg[8]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w9914_
	);
	LUT4 #(
		.INIT('h8088)
	) name8165 (
		_w2227_,
		_w2241_,
		_w9913_,
		_w9914_,
		_w9915_
	);
	LUT3 #(
		.INIT('h80)
	) name8166 (
		\u4_u2_buf1_reg[8]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w9916_
	);
	LUT4 #(
		.INIT('hf5f3)
	) name8167 (
		\u4_u2_buf0_reg[8]/P0001 ,
		\u4_u2_csr0_reg[8]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w9917_
	);
	LUT4 #(
		.INIT('h8088)
	) name8168 (
		_w2228_,
		_w2240_,
		_w9916_,
		_w9917_,
		_w9918_
	);
	LUT2 #(
		.INIT('h1)
	) name8169 (
		_w9915_,
		_w9918_,
		_w9919_
	);
	LUT3 #(
		.INIT('h80)
	) name8170 (
		\u4_u0_buf1_reg[8]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w9920_
	);
	LUT4 #(
		.INIT('hf5f3)
	) name8171 (
		\u4_u0_buf0_reg[8]/P0001 ,
		\u4_u0_csr0_reg[8]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w9921_
	);
	LUT4 #(
		.INIT('h8088)
	) name8172 (
		_w2240_,
		_w2241_,
		_w9920_,
		_w9921_,
		_w9922_
	);
	LUT3 #(
		.INIT('h80)
	) name8173 (
		\u4_u3_buf1_reg[8]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w9923_
	);
	LUT4 #(
		.INIT('hf5f3)
	) name8174 (
		\u4_u3_buf0_reg[8]/P0001 ,
		\u4_u3_csr0_reg[8]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w9924_
	);
	LUT4 #(
		.INIT('h8088)
	) name8175 (
		_w2227_,
		_w2228_,
		_w9923_,
		_w9924_,
		_w9925_
	);
	LUT4 #(
		.INIT('h0200)
	) name8176 (
		\u1_sof_time_reg[8]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w9926_
	);
	LUT4 #(
		.INIT('h0020)
	) name8177 (
		\u4_inta_msk_reg[8]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w9927_
	);
	LUT3 #(
		.INIT('ha8)
	) name8178 (
		_w5861_,
		_w9926_,
		_w9927_,
		_w9928_
	);
	LUT3 #(
		.INIT('h01)
	) name8179 (
		_w9922_,
		_w9925_,
		_w9928_,
		_w9929_
	);
	LUT2 #(
		.INIT('h7)
	) name8180 (
		_w9919_,
		_w9929_,
		_w9930_
	);
	LUT4 #(
		.INIT('h2a00)
	) name8181 (
		rst_i_pad,
		\u1_u3_uc_bsel_set_reg/P0001 ,
		\u4_u2_ep_match_r_reg/P0001 ,
		\u4_u2_uc_dpd_reg[0]/P0001 ,
		_w9931_
	);
	LUT4 #(
		.INIT('h8000)
	) name8182 (
		rst_i_pad,
		\u1_u3_idin_reg[2]/P0001 ,
		\u1_u3_uc_bsel_set_reg/P0001 ,
		\u4_u2_ep_match_r_reg/P0001 ,
		_w9932_
	);
	LUT2 #(
		.INIT('he)
	) name8183 (
		_w9931_,
		_w9932_,
		_w9933_
	);
	LUT4 #(
		.INIT('h2a00)
	) name8184 (
		rst_i_pad,
		\u1_u3_uc_bsel_set_reg/P0001 ,
		\u4_u3_ep_match_r_reg/P0001 ,
		\u4_u3_uc_dpd_reg[1]/P0001 ,
		_w9934_
	);
	LUT4 #(
		.INIT('h8000)
	) name8185 (
		rst_i_pad,
		\u1_u3_idin_reg[3]/P0001 ,
		\u1_u3_uc_bsel_set_reg/P0001 ,
		\u4_u3_ep_match_r_reg/P0001 ,
		_w9935_
	);
	LUT2 #(
		.INIT('he)
	) name8186 (
		_w9934_,
		_w9935_,
		_w9936_
	);
	LUT4 #(
		.INIT('h2a00)
	) name8187 (
		rst_i_pad,
		\u1_u3_uc_bsel_set_reg/P0001 ,
		\u4_u0_ep_match_r_reg/P0001 ,
		\u4_u0_uc_bsel_reg[0]/P0001 ,
		_w9937_
	);
	LUT4 #(
		.INIT('h8000)
	) name8188 (
		rst_i_pad,
		\u1_u3_idin_reg[0]/P0001 ,
		\u1_u3_uc_bsel_set_reg/P0001 ,
		\u4_u0_ep_match_r_reg/P0001 ,
		_w9938_
	);
	LUT2 #(
		.INIT('he)
	) name8189 (
		_w9937_,
		_w9938_,
		_w9939_
	);
	LUT4 #(
		.INIT('h2a00)
	) name8190 (
		rst_i_pad,
		\u1_u3_uc_bsel_set_reg/P0001 ,
		\u4_u0_ep_match_r_reg/P0001 ,
		\u4_u0_uc_bsel_reg[1]/P0001 ,
		_w9940_
	);
	LUT4 #(
		.INIT('h8000)
	) name8191 (
		rst_i_pad,
		\u1_u3_idin_reg[1]/P0001 ,
		\u1_u3_uc_bsel_set_reg/P0001 ,
		\u4_u0_ep_match_r_reg/P0001 ,
		_w9941_
	);
	LUT2 #(
		.INIT('he)
	) name8192 (
		_w9940_,
		_w9941_,
		_w9942_
	);
	LUT4 #(
		.INIT('h2a00)
	) name8193 (
		rst_i_pad,
		\u1_u3_uc_bsel_set_reg/P0001 ,
		\u4_u0_ep_match_r_reg/P0001 ,
		\u4_u0_uc_dpd_reg[0]/P0001 ,
		_w9943_
	);
	LUT4 #(
		.INIT('h8000)
	) name8194 (
		rst_i_pad,
		\u1_u3_idin_reg[2]/P0001 ,
		\u1_u3_uc_bsel_set_reg/P0001 ,
		\u4_u0_ep_match_r_reg/P0001 ,
		_w9944_
	);
	LUT2 #(
		.INIT('he)
	) name8195 (
		_w9943_,
		_w9944_,
		_w9945_
	);
	LUT4 #(
		.INIT('h2a00)
	) name8196 (
		rst_i_pad,
		\u1_u3_uc_bsel_set_reg/P0001 ,
		\u4_u0_ep_match_r_reg/P0001 ,
		\u4_u0_uc_dpd_reg[1]/P0001 ,
		_w9946_
	);
	LUT4 #(
		.INIT('h8000)
	) name8197 (
		rst_i_pad,
		\u1_u3_idin_reg[3]/P0001 ,
		\u1_u3_uc_bsel_set_reg/P0001 ,
		\u4_u0_ep_match_r_reg/P0001 ,
		_w9947_
	);
	LUT2 #(
		.INIT('he)
	) name8198 (
		_w9946_,
		_w9947_,
		_w9948_
	);
	LUT3 #(
		.INIT('h08)
	) name8199 (
		\u1_u0_pid_reg[0]/NET0131 ,
		\u1_u0_pid_reg[1]/NET0131 ,
		\u1_u0_pid_reg[2]/NET0131 ,
		_w9949_
	);
	LUT3 #(
		.INIT('h04)
	) name8200 (
		_w7762_,
		_w8145_,
		_w9949_,
		_w9950_
	);
	LUT3 #(
		.INIT('h02)
	) name8201 (
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		\u4_csr_reg[28]/P0001 ,
		_w9951_
	);
	LUT4 #(
		.INIT('h1357)
	) name8202 (
		_w2120_,
		_w7772_,
		_w8136_,
		_w9951_,
		_w9952_
	);
	LUT3 #(
		.INIT('h8a)
	) name8203 (
		_w3961_,
		_w7762_,
		_w8145_,
		_w9953_
	);
	LUT3 #(
		.INIT('hba)
	) name8204 (
		_w9950_,
		_w9952_,
		_w9953_,
		_w9954_
	);
	LUT4 #(
		.INIT('hc4c0)
	) name8205 (
		\u0_u0_me_cnt_100_ms_reg/P0001 ,
		_w4103_,
		_w4333_,
		_w5762_,
		_w9955_
	);
	LUT4 #(
		.INIT('h2a00)
	) name8206 (
		rst_i_pad,
		\u1_u3_uc_bsel_set_reg/P0001 ,
		\u4_u1_ep_match_r_reg/P0001 ,
		\u4_u1_uc_bsel_reg[0]/P0001 ,
		_w9956_
	);
	LUT4 #(
		.INIT('h8000)
	) name8207 (
		rst_i_pad,
		\u1_u3_idin_reg[0]/P0001 ,
		\u1_u3_uc_bsel_set_reg/P0001 ,
		\u4_u1_ep_match_r_reg/P0001 ,
		_w9957_
	);
	LUT2 #(
		.INIT('he)
	) name8208 (
		_w9956_,
		_w9957_,
		_w9958_
	);
	LUT4 #(
		.INIT('h2a00)
	) name8209 (
		rst_i_pad,
		\u1_u3_uc_bsel_set_reg/P0001 ,
		\u4_u1_ep_match_r_reg/P0001 ,
		\u4_u1_uc_bsel_reg[1]/P0001 ,
		_w9959_
	);
	LUT4 #(
		.INIT('h8000)
	) name8210 (
		rst_i_pad,
		\u1_u3_idin_reg[1]/P0001 ,
		\u1_u3_uc_bsel_set_reg/P0001 ,
		\u4_u1_ep_match_r_reg/P0001 ,
		_w9960_
	);
	LUT2 #(
		.INIT('he)
	) name8211 (
		_w9959_,
		_w9960_,
		_w9961_
	);
	LUT4 #(
		.INIT('h2a00)
	) name8212 (
		rst_i_pad,
		\u1_u3_uc_bsel_set_reg/P0001 ,
		\u4_u1_ep_match_r_reg/P0001 ,
		\u4_u1_uc_dpd_reg[0]/P0001 ,
		_w9962_
	);
	LUT4 #(
		.INIT('h8000)
	) name8213 (
		rst_i_pad,
		\u1_u3_idin_reg[2]/P0001 ,
		\u1_u3_uc_bsel_set_reg/P0001 ,
		\u4_u1_ep_match_r_reg/P0001 ,
		_w9963_
	);
	LUT2 #(
		.INIT('he)
	) name8214 (
		_w9962_,
		_w9963_,
		_w9964_
	);
	LUT4 #(
		.INIT('h2a00)
	) name8215 (
		rst_i_pad,
		\u1_u3_uc_bsel_set_reg/P0001 ,
		\u4_u1_ep_match_r_reg/P0001 ,
		\u4_u1_uc_dpd_reg[1]/P0001 ,
		_w9965_
	);
	LUT4 #(
		.INIT('h8000)
	) name8216 (
		rst_i_pad,
		\u1_u3_idin_reg[3]/P0001 ,
		\u1_u3_uc_bsel_set_reg/P0001 ,
		\u4_u1_ep_match_r_reg/P0001 ,
		_w9966_
	);
	LUT2 #(
		.INIT('he)
	) name8217 (
		_w9965_,
		_w9966_,
		_w9967_
	);
	LUT3 #(
		.INIT('h59)
	) name8218 (
		\u1_u3_new_sizeb_reg[0]/P0001 ,
		_w2788_,
		_w2790_,
		_w9968_
	);
	LUT3 #(
		.INIT('h10)
	) name8219 (
		\u0_u0_T2_wakeup_reg/P0001 ,
		\u0_u0_state_reg[4]/NET0131 ,
		\u0_u0_state_reg[5]/P0001 ,
		_w9969_
	);
	LUT3 #(
		.INIT('h07)
	) name8220 (
		\u0_u0_T1_gt_5_0_mS_reg/P0001 ,
		\u0_u0_resume_req_s_reg/P0001 ,
		\u0_u0_state_reg[5]/P0001 ,
		_w9970_
	);
	LUT4 #(
		.INIT('h0004)
	) name8221 (
		_w4119_,
		_w4341_,
		_w4354_,
		_w9970_,
		_w9971_
	);
	LUT4 #(
		.INIT('h135f)
	) name8222 (
		_w4319_,
		_w7962_,
		_w9969_,
		_w9971_,
		_w9972_
	);
	LUT2 #(
		.INIT('h2)
	) name8223 (
		_w4103_,
		_w9972_,
		_w9973_
	);
	LUT4 #(
		.INIT('h2a3f)
	) name8224 (
		\u0_u0_T2_gt_1_0_mS_reg/P0001 ,
		_w4320_,
		_w4338_,
		_w9603_,
		_w9974_
	);
	LUT2 #(
		.INIT('h2)
	) name8225 (
		_w4103_,
		_w9974_,
		_w9975_
	);
	LUT4 #(
		.INIT('h0020)
	) name8226 (
		\u4_intb_msk_reg[0]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w9976_
	);
	LUT4 #(
		.INIT('h0200)
	) name8227 (
		\u1_frame_no_r_reg[0]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w9977_
	);
	LUT3 #(
		.INIT('ha8)
	) name8228 (
		_w5861_,
		_w9976_,
		_w9977_,
		_w9978_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name8229 (
		\u4_u1_buf1_reg[16]/P0001 ,
		\u4_u1_csr1_reg[1]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w9979_
	);
	LUT4 #(
		.INIT('hf53f)
	) name8230 (
		\u4_u1_buf0_reg[16]/P0001 ,
		\u4_u1_ienb_reg[0]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w9980_
	);
	LUT4 #(
		.INIT('h0888)
	) name8231 (
		_w2227_,
		_w2241_,
		_w9979_,
		_w9980_,
		_w9981_
	);
	LUT2 #(
		.INIT('h1)
	) name8232 (
		_w9978_,
		_w9981_,
		_w9982_
	);
	LUT4 #(
		.INIT('hf5f3)
	) name8233 (
		\u4_u3_buf0_reg[16]/P0001 ,
		\u4_u3_csr1_reg[1]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w9983_
	);
	LUT4 #(
		.INIT('h5f3f)
	) name8234 (
		\u4_u3_buf1_reg[16]/P0001 ,
		\u4_u3_ienb_reg[0]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w9984_
	);
	LUT4 #(
		.INIT('h0888)
	) name8235 (
		_w2227_,
		_w2228_,
		_w9983_,
		_w9984_,
		_w9985_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name8236 (
		\u4_u0_buf1_reg[16]/P0001 ,
		\u4_u0_csr1_reg[1]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w9986_
	);
	LUT4 #(
		.INIT('hf53f)
	) name8237 (
		\u4_u0_buf0_reg[16]/P0001 ,
		\u4_u0_ienb_reg[0]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w9987_
	);
	LUT4 #(
		.INIT('h0888)
	) name8238 (
		_w2240_,
		_w2241_,
		_w9986_,
		_w9987_,
		_w9988_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name8239 (
		\u4_u2_buf1_reg[16]/P0001 ,
		\u4_u2_csr1_reg[1]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w9989_
	);
	LUT4 #(
		.INIT('hf53f)
	) name8240 (
		\u4_u2_buf0_reg[16]/P0001 ,
		\u4_u2_ienb_reg[0]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w9990_
	);
	LUT4 #(
		.INIT('h0888)
	) name8241 (
		_w2228_,
		_w2240_,
		_w9989_,
		_w9990_,
		_w9991_
	);
	LUT3 #(
		.INIT('h01)
	) name8242 (
		_w9985_,
		_w9988_,
		_w9991_,
		_w9992_
	);
	LUT2 #(
		.INIT('h7)
	) name8243 (
		_w9982_,
		_w9992_,
		_w9993_
	);
	LUT4 #(
		.INIT('h0020)
	) name8244 (
		\u4_intb_msk_reg[1]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w9994_
	);
	LUT4 #(
		.INIT('h0200)
	) name8245 (
		\u1_frame_no_r_reg[1]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w9995_
	);
	LUT3 #(
		.INIT('ha8)
	) name8246 (
		_w5861_,
		_w9994_,
		_w9995_,
		_w9996_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name8247 (
		\u4_u1_buf1_reg[17]/P0001 ,
		\u4_u1_csr1_reg[2]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w9997_
	);
	LUT4 #(
		.INIT('hf53f)
	) name8248 (
		\u4_u1_buf0_reg[17]/P0001 ,
		\u4_u1_ienb_reg[1]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w9998_
	);
	LUT4 #(
		.INIT('h0888)
	) name8249 (
		_w2227_,
		_w2241_,
		_w9997_,
		_w9998_,
		_w9999_
	);
	LUT2 #(
		.INIT('h1)
	) name8250 (
		_w9996_,
		_w9999_,
		_w10000_
	);
	LUT4 #(
		.INIT('hf5f3)
	) name8251 (
		\u4_u3_buf0_reg[17]/P0001 ,
		\u4_u3_csr1_reg[2]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w10001_
	);
	LUT4 #(
		.INIT('h5f3f)
	) name8252 (
		\u4_u3_buf1_reg[17]/P0001 ,
		\u4_u3_ienb_reg[1]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w10002_
	);
	LUT4 #(
		.INIT('h0888)
	) name8253 (
		_w2227_,
		_w2228_,
		_w10001_,
		_w10002_,
		_w10003_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name8254 (
		\u4_u0_buf1_reg[17]/P0001 ,
		\u4_u0_csr1_reg[2]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w10004_
	);
	LUT4 #(
		.INIT('hf53f)
	) name8255 (
		\u4_u0_buf0_reg[17]/P0001 ,
		\u4_u0_ienb_reg[1]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w10005_
	);
	LUT4 #(
		.INIT('h0888)
	) name8256 (
		_w2240_,
		_w2241_,
		_w10004_,
		_w10005_,
		_w10006_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name8257 (
		\u4_u2_buf1_reg[17]/P0001 ,
		\u4_u2_csr1_reg[2]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w10007_
	);
	LUT4 #(
		.INIT('hf53f)
	) name8258 (
		\u4_u2_buf0_reg[17]/P0001 ,
		\u4_u2_ienb_reg[1]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w10008_
	);
	LUT4 #(
		.INIT('h0888)
	) name8259 (
		_w2228_,
		_w2240_,
		_w10007_,
		_w10008_,
		_w10009_
	);
	LUT3 #(
		.INIT('h01)
	) name8260 (
		_w10003_,
		_w10006_,
		_w10009_,
		_w10010_
	);
	LUT2 #(
		.INIT('h7)
	) name8261 (
		_w10000_,
		_w10010_,
		_w10011_
	);
	LUT4 #(
		.INIT('h0020)
	) name8262 (
		\u4_intb_msk_reg[2]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w10012_
	);
	LUT4 #(
		.INIT('h0200)
	) name8263 (
		\u1_frame_no_r_reg[2]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w10013_
	);
	LUT3 #(
		.INIT('ha8)
	) name8264 (
		_w5861_,
		_w10012_,
		_w10013_,
		_w10014_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name8265 (
		\u4_u1_buf1_reg[18]/P0001 ,
		\u4_u1_csr1_reg[3]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w10015_
	);
	LUT4 #(
		.INIT('hf53f)
	) name8266 (
		\u4_u1_buf0_reg[18]/P0001 ,
		\u4_u1_ienb_reg[2]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w10016_
	);
	LUT4 #(
		.INIT('h0888)
	) name8267 (
		_w2227_,
		_w2241_,
		_w10015_,
		_w10016_,
		_w10017_
	);
	LUT2 #(
		.INIT('h1)
	) name8268 (
		_w10014_,
		_w10017_,
		_w10018_
	);
	LUT4 #(
		.INIT('hf5f3)
	) name8269 (
		\u4_u2_buf0_reg[18]/P0001 ,
		\u4_u2_csr1_reg[3]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w10019_
	);
	LUT4 #(
		.INIT('h5f3f)
	) name8270 (
		\u4_u2_buf1_reg[18]/P0001 ,
		\u4_u2_ienb_reg[2]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w10020_
	);
	LUT4 #(
		.INIT('h0888)
	) name8271 (
		_w2228_,
		_w2240_,
		_w10019_,
		_w10020_,
		_w10021_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name8272 (
		\u4_u0_buf1_reg[18]/P0001 ,
		\u4_u0_csr1_reg[3]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w10022_
	);
	LUT4 #(
		.INIT('hf53f)
	) name8273 (
		\u4_u0_buf0_reg[18]/P0001 ,
		\u4_u0_ienb_reg[2]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w10023_
	);
	LUT4 #(
		.INIT('h0888)
	) name8274 (
		_w2240_,
		_w2241_,
		_w10022_,
		_w10023_,
		_w10024_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name8275 (
		\u4_u3_buf1_reg[18]/P0001 ,
		\u4_u3_csr1_reg[3]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w10025_
	);
	LUT4 #(
		.INIT('hf53f)
	) name8276 (
		\u4_u3_buf0_reg[18]/P0001 ,
		\u4_u3_ienb_reg[2]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w10026_
	);
	LUT4 #(
		.INIT('h0888)
	) name8277 (
		_w2227_,
		_w2228_,
		_w10025_,
		_w10026_,
		_w10027_
	);
	LUT3 #(
		.INIT('h01)
	) name8278 (
		_w10021_,
		_w10024_,
		_w10027_,
		_w10028_
	);
	LUT2 #(
		.INIT('h7)
	) name8279 (
		_w10018_,
		_w10028_,
		_w10029_
	);
	LUT4 #(
		.INIT('h0020)
	) name8280 (
		\u4_intb_msk_reg[3]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w10030_
	);
	LUT4 #(
		.INIT('h0200)
	) name8281 (
		\u1_frame_no_r_reg[3]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w10031_
	);
	LUT3 #(
		.INIT('ha8)
	) name8282 (
		_w5861_,
		_w10030_,
		_w10031_,
		_w10032_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name8283 (
		\u4_u1_buf1_reg[19]/P0001 ,
		\u4_u1_csr1_reg[4]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w10033_
	);
	LUT4 #(
		.INIT('hf53f)
	) name8284 (
		\u4_u1_buf0_reg[19]/P0001 ,
		\u4_u1_ienb_reg[3]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w10034_
	);
	LUT4 #(
		.INIT('h0888)
	) name8285 (
		_w2227_,
		_w2241_,
		_w10033_,
		_w10034_,
		_w10035_
	);
	LUT2 #(
		.INIT('h1)
	) name8286 (
		_w10032_,
		_w10035_,
		_w10036_
	);
	LUT4 #(
		.INIT('hf5f3)
	) name8287 (
		\u4_u2_buf0_reg[19]/P0001 ,
		\u4_u2_csr1_reg[4]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w10037_
	);
	LUT4 #(
		.INIT('h5f3f)
	) name8288 (
		\u4_u2_buf1_reg[19]/P0001 ,
		\u4_u2_ienb_reg[3]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w10038_
	);
	LUT4 #(
		.INIT('h0888)
	) name8289 (
		_w2228_,
		_w2240_,
		_w10037_,
		_w10038_,
		_w10039_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name8290 (
		\u4_u0_buf1_reg[19]/P0001 ,
		\u4_u0_csr1_reg[4]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w10040_
	);
	LUT4 #(
		.INIT('hf53f)
	) name8291 (
		\u4_u0_buf0_reg[19]/P0001 ,
		\u4_u0_ienb_reg[3]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w10041_
	);
	LUT4 #(
		.INIT('h0888)
	) name8292 (
		_w2240_,
		_w2241_,
		_w10040_,
		_w10041_,
		_w10042_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name8293 (
		\u4_u3_buf1_reg[19]/P0001 ,
		\u4_u3_csr1_reg[4]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w10043_
	);
	LUT4 #(
		.INIT('hf53f)
	) name8294 (
		\u4_u3_buf0_reg[19]/P0001 ,
		\u4_u3_ienb_reg[3]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w10044_
	);
	LUT4 #(
		.INIT('h0888)
	) name8295 (
		_w2227_,
		_w2228_,
		_w10043_,
		_w10044_,
		_w10045_
	);
	LUT3 #(
		.INIT('h01)
	) name8296 (
		_w10039_,
		_w10042_,
		_w10045_,
		_w10046_
	);
	LUT2 #(
		.INIT('h7)
	) name8297 (
		_w10036_,
		_w10046_,
		_w10047_
	);
	LUT4 #(
		.INIT('h0080)
	) name8298 (
		\u4_int_srcb_reg[5]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w10048_
	);
	LUT4 #(
		.INIT('h0200)
	) name8299 (
		\u1_frame_no_r_reg[9]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w10049_
	);
	LUT3 #(
		.INIT('ha8)
	) name8300 (
		_w5861_,
		_w10048_,
		_w10049_,
		_w10050_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name8301 (
		\u4_u1_buf1_reg[25]/P0001 ,
		\u4_u1_csr1_reg[10]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w10051_
	);
	LUT4 #(
		.INIT('hf53f)
	) name8302 (
		\u4_u1_buf0_reg[25]/P0001 ,
		\u4_u1_iena_reg[1]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w10052_
	);
	LUT4 #(
		.INIT('h0888)
	) name8303 (
		_w2227_,
		_w2241_,
		_w10051_,
		_w10052_,
		_w10053_
	);
	LUT2 #(
		.INIT('h1)
	) name8304 (
		_w10050_,
		_w10053_,
		_w10054_
	);
	LUT4 #(
		.INIT('hf5f3)
	) name8305 (
		\u4_u3_buf0_reg[25]/P0001 ,
		\u4_u3_csr1_reg[10]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w10055_
	);
	LUT4 #(
		.INIT('h5f3f)
	) name8306 (
		\u4_u3_buf1_reg[25]/P0001 ,
		\u4_u3_iena_reg[1]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w10056_
	);
	LUT4 #(
		.INIT('h0888)
	) name8307 (
		_w2227_,
		_w2228_,
		_w10055_,
		_w10056_,
		_w10057_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name8308 (
		\u4_u0_buf1_reg[25]/P0001 ,
		\u4_u0_csr1_reg[10]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w10058_
	);
	LUT4 #(
		.INIT('hf53f)
	) name8309 (
		\u4_u0_buf0_reg[25]/P0001 ,
		\u4_u0_iena_reg[1]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w10059_
	);
	LUT4 #(
		.INIT('h0888)
	) name8310 (
		_w2240_,
		_w2241_,
		_w10058_,
		_w10059_,
		_w10060_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name8311 (
		\u4_u2_buf1_reg[25]/P0001 ,
		\u4_u2_csr1_reg[10]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w10061_
	);
	LUT4 #(
		.INIT('hf53f)
	) name8312 (
		\u4_u2_buf0_reg[25]/P0001 ,
		\u4_u2_iena_reg[1]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w10062_
	);
	LUT4 #(
		.INIT('h0888)
	) name8313 (
		_w2228_,
		_w2240_,
		_w10061_,
		_w10062_,
		_w10063_
	);
	LUT3 #(
		.INIT('h01)
	) name8314 (
		_w10057_,
		_w10060_,
		_w10063_,
		_w10064_
	);
	LUT2 #(
		.INIT('h7)
	) name8315 (
		_w10054_,
		_w10064_,
		_w10065_
	);
	LUT4 #(
		.INIT('h0080)
	) name8316 (
		\u4_int_srcb_reg[6]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w10066_
	);
	LUT4 #(
		.INIT('h0200)
	) name8317 (
		\u1_frame_no_r_reg[10]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w10067_
	);
	LUT3 #(
		.INIT('ha8)
	) name8318 (
		_w5861_,
		_w10066_,
		_w10067_,
		_w10068_
	);
	LUT4 #(
		.INIT('h5f3f)
	) name8319 (
		\u4_u1_buf1_reg[26]/P0001 ,
		\u4_u1_iena_reg[2]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w10069_
	);
	LUT4 #(
		.INIT('hf5f3)
	) name8320 (
		\u4_u1_buf0_reg[26]/P0001 ,
		\u4_u1_csr1_reg[11]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w10070_
	);
	LUT4 #(
		.INIT('h0888)
	) name8321 (
		_w2227_,
		_w2241_,
		_w10069_,
		_w10070_,
		_w10071_
	);
	LUT2 #(
		.INIT('h1)
	) name8322 (
		_w10068_,
		_w10071_,
		_w10072_
	);
	LUT4 #(
		.INIT('hf5f3)
	) name8323 (
		\u4_u3_buf0_reg[26]/P0001 ,
		\u4_u3_csr1_reg[11]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w10073_
	);
	LUT4 #(
		.INIT('h5f3f)
	) name8324 (
		\u4_u3_buf1_reg[26]/P0001 ,
		\u4_u3_iena_reg[2]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w10074_
	);
	LUT4 #(
		.INIT('h0888)
	) name8325 (
		_w2227_,
		_w2228_,
		_w10073_,
		_w10074_,
		_w10075_
	);
	LUT4 #(
		.INIT('h5f3f)
	) name8326 (
		\u4_u0_buf1_reg[26]/P0001 ,
		\u4_u0_iena_reg[2]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w10076_
	);
	LUT4 #(
		.INIT('hf5f3)
	) name8327 (
		\u4_u0_buf0_reg[26]/P0001 ,
		\u4_u0_csr1_reg[11]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w10077_
	);
	LUT4 #(
		.INIT('h0888)
	) name8328 (
		_w2240_,
		_w2241_,
		_w10076_,
		_w10077_,
		_w10078_
	);
	LUT4 #(
		.INIT('h5f3f)
	) name8329 (
		\u4_u2_buf1_reg[26]/P0001 ,
		\u4_u2_iena_reg[2]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w10079_
	);
	LUT4 #(
		.INIT('hf5f3)
	) name8330 (
		\u4_u2_buf0_reg[26]/P0001 ,
		\u4_u2_csr1_reg[11]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w10080_
	);
	LUT4 #(
		.INIT('h0888)
	) name8331 (
		_w2228_,
		_w2240_,
		_w10079_,
		_w10080_,
		_w10081_
	);
	LUT3 #(
		.INIT('h01)
	) name8332 (
		_w10075_,
		_w10078_,
		_w10081_,
		_w10082_
	);
	LUT2 #(
		.INIT('h7)
	) name8333 (
		_w10072_,
		_w10082_,
		_w10083_
	);
	LUT4 #(
		.INIT('h0080)
	) name8334 (
		\u4_int_srcb_reg[8]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w10084_
	);
	LUT4 #(
		.INIT('h0200)
	) name8335 (
		\u1_mfm_cnt_reg[0]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w10085_
	);
	LUT3 #(
		.INIT('ha8)
	) name8336 (
		_w5861_,
		_w10084_,
		_w10085_,
		_w10086_
	);
	LUT4 #(
		.INIT('h5f3f)
	) name8337 (
		\u4_u1_buf1_reg[28]/P0001 ,
		\u4_u1_iena_reg[4]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w10087_
	);
	LUT4 #(
		.INIT('hf5f3)
	) name8338 (
		\u4_u1_buf0_reg[28]/P0001 ,
		\u4_u1_uc_dpd_reg[0]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w10088_
	);
	LUT4 #(
		.INIT('h0888)
	) name8339 (
		_w2227_,
		_w2241_,
		_w10087_,
		_w10088_,
		_w10089_
	);
	LUT2 #(
		.INIT('h1)
	) name8340 (
		_w10086_,
		_w10089_,
		_w10090_
	);
	LUT4 #(
		.INIT('hf53f)
	) name8341 (
		\u4_u2_buf0_reg[28]/P0001 ,
		\u4_u2_iena_reg[4]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w10091_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name8342 (
		\u4_u2_buf1_reg[28]/P0001 ,
		\u4_u2_uc_dpd_reg[0]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w10092_
	);
	LUT4 #(
		.INIT('h0888)
	) name8343 (
		_w2228_,
		_w2240_,
		_w10091_,
		_w10092_,
		_w10093_
	);
	LUT4 #(
		.INIT('h5f3f)
	) name8344 (
		\u4_u0_buf1_reg[28]/P0001 ,
		\u4_u0_iena_reg[4]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w10094_
	);
	LUT4 #(
		.INIT('hf5f3)
	) name8345 (
		\u4_u0_buf0_reg[28]/P0001 ,
		\u4_u0_uc_dpd_reg[0]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w10095_
	);
	LUT4 #(
		.INIT('h0888)
	) name8346 (
		_w2240_,
		_w2241_,
		_w10094_,
		_w10095_,
		_w10096_
	);
	LUT4 #(
		.INIT('h5f3f)
	) name8347 (
		\u4_u3_buf1_reg[28]/P0001 ,
		\u4_u3_iena_reg[4]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w10097_
	);
	LUT4 #(
		.INIT('hf5f3)
	) name8348 (
		\u4_u3_buf0_reg[28]/P0001 ,
		\u4_u3_uc_dpd_reg[0]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w10098_
	);
	LUT4 #(
		.INIT('h0888)
	) name8349 (
		_w2227_,
		_w2228_,
		_w10097_,
		_w10098_,
		_w10099_
	);
	LUT3 #(
		.INIT('h01)
	) name8350 (
		_w10093_,
		_w10096_,
		_w10099_,
		_w10100_
	);
	LUT2 #(
		.INIT('h7)
	) name8351 (
		_w10090_,
		_w10100_,
		_w10101_
	);
	LUT4 #(
		.INIT('hf5f3)
	) name8352 (
		\u4_u2_buf0_reg[21]/P0001 ,
		\u4_u2_csr1_reg[6]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w10102_
	);
	LUT4 #(
		.INIT('h5f3f)
	) name8353 (
		\u4_u2_buf1_reg[21]/P0001 ,
		\u4_u2_ienb_reg[5]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w10103_
	);
	LUT4 #(
		.INIT('h0888)
	) name8354 (
		_w2228_,
		_w2240_,
		_w10102_,
		_w10103_,
		_w10104_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name8355 (
		\u4_u3_buf1_reg[21]/P0001 ,
		\u4_u3_csr1_reg[6]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w10105_
	);
	LUT4 #(
		.INIT('hf53f)
	) name8356 (
		\u4_u3_buf0_reg[21]/P0001 ,
		\u4_u3_ienb_reg[5]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w10106_
	);
	LUT4 #(
		.INIT('h0888)
	) name8357 (
		_w2227_,
		_w2228_,
		_w10105_,
		_w10106_,
		_w10107_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name8358 (
		\u4_u0_buf1_reg[21]/P0001 ,
		\u4_u0_csr1_reg[6]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w10108_
	);
	LUT4 #(
		.INIT('hf53f)
	) name8359 (
		\u4_u0_buf0_reg[21]/P0001 ,
		\u4_u0_ienb_reg[5]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w10109_
	);
	LUT4 #(
		.INIT('h0888)
	) name8360 (
		_w2240_,
		_w2241_,
		_w10108_,
		_w10109_,
		_w10110_
	);
	LUT3 #(
		.INIT('h01)
	) name8361 (
		_w10104_,
		_w10107_,
		_w10110_,
		_w10111_
	);
	LUT4 #(
		.INIT('h0200)
	) name8362 (
		\u1_frame_no_r_reg[5]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w10112_
	);
	LUT4 #(
		.INIT('h0020)
	) name8363 (
		\u4_intb_msk_reg[5]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w10113_
	);
	LUT4 #(
		.INIT('h0080)
	) name8364 (
		\u4_int_srcb_reg[1]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w10114_
	);
	LUT4 #(
		.INIT('haaa8)
	) name8365 (
		_w5861_,
		_w10112_,
		_w10113_,
		_w10114_,
		_w10115_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name8366 (
		\u4_u1_buf1_reg[21]/P0001 ,
		\u4_u1_csr1_reg[6]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w10116_
	);
	LUT4 #(
		.INIT('hf53f)
	) name8367 (
		\u4_u1_buf0_reg[21]/P0001 ,
		\u4_u1_ienb_reg[5]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w10117_
	);
	LUT4 #(
		.INIT('h0888)
	) name8368 (
		_w2227_,
		_w2241_,
		_w10116_,
		_w10117_,
		_w10118_
	);
	LUT2 #(
		.INIT('h1)
	) name8369 (
		_w10115_,
		_w10118_,
		_w10119_
	);
	LUT2 #(
		.INIT('h7)
	) name8370 (
		_w10111_,
		_w10119_,
		_w10120_
	);
	LUT4 #(
		.INIT('hf5f3)
	) name8371 (
		\u4_u3_buf0_reg[24]/P0001 ,
		\u4_u3_csr1_reg[9]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w10121_
	);
	LUT4 #(
		.INIT('h5f3f)
	) name8372 (
		\u4_u3_buf1_reg[24]/P0001 ,
		\u4_u3_iena_reg[0]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w10122_
	);
	LUT4 #(
		.INIT('h0888)
	) name8373 (
		_w2227_,
		_w2228_,
		_w10121_,
		_w10122_,
		_w10123_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name8374 (
		\u4_u2_buf1_reg[24]/P0001 ,
		\u4_u2_csr1_reg[9]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w10124_
	);
	LUT4 #(
		.INIT('hf53f)
	) name8375 (
		\u4_u2_buf0_reg[24]/P0001 ,
		\u4_u2_iena_reg[0]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w10125_
	);
	LUT4 #(
		.INIT('h0888)
	) name8376 (
		_w2228_,
		_w2240_,
		_w10124_,
		_w10125_,
		_w10126_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name8377 (
		\u4_u0_buf1_reg[24]/P0001 ,
		\u4_u0_csr1_reg[9]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w10127_
	);
	LUT4 #(
		.INIT('hf53f)
	) name8378 (
		\u4_u0_buf0_reg[24]/P0001 ,
		\u4_u0_iena_reg[0]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w10128_
	);
	LUT4 #(
		.INIT('h0888)
	) name8379 (
		_w2240_,
		_w2241_,
		_w10127_,
		_w10128_,
		_w10129_
	);
	LUT3 #(
		.INIT('h01)
	) name8380 (
		_w10123_,
		_w10126_,
		_w10129_,
		_w10130_
	);
	LUT4 #(
		.INIT('h0200)
	) name8381 (
		\u1_frame_no_r_reg[8]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w10131_
	);
	LUT4 #(
		.INIT('h0020)
	) name8382 (
		\u4_intb_msk_reg[8]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w10132_
	);
	LUT4 #(
		.INIT('h0080)
	) name8383 (
		\u4_int_srcb_reg[4]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w10133_
	);
	LUT4 #(
		.INIT('haaa8)
	) name8384 (
		_w5861_,
		_w10131_,
		_w10132_,
		_w10133_,
		_w10134_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name8385 (
		\u4_u1_buf1_reg[24]/P0001 ,
		\u4_u1_csr1_reg[9]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w10135_
	);
	LUT4 #(
		.INIT('hf53f)
	) name8386 (
		\u4_u1_buf0_reg[24]/P0001 ,
		\u4_u1_iena_reg[0]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w10136_
	);
	LUT4 #(
		.INIT('h0888)
	) name8387 (
		_w2227_,
		_w2241_,
		_w10135_,
		_w10136_,
		_w10137_
	);
	LUT2 #(
		.INIT('h1)
	) name8388 (
		_w10134_,
		_w10137_,
		_w10138_
	);
	LUT2 #(
		.INIT('h7)
	) name8389 (
		_w10130_,
		_w10138_,
		_w10139_
	);
	LUT4 #(
		.INIT('hf5f3)
	) name8390 (
		\u4_u3_buf0_reg[20]/P0001 ,
		\u4_u3_csr1_reg[5]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w10140_
	);
	LUT4 #(
		.INIT('h5f3f)
	) name8391 (
		\u4_u3_buf1_reg[20]/P0001 ,
		\u4_u3_ienb_reg[4]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w10141_
	);
	LUT4 #(
		.INIT('h0888)
	) name8392 (
		_w2227_,
		_w2228_,
		_w10140_,
		_w10141_,
		_w10142_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name8393 (
		\u4_u2_buf1_reg[20]/P0001 ,
		\u4_u2_csr1_reg[5]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w10143_
	);
	LUT4 #(
		.INIT('hf53f)
	) name8394 (
		\u4_u2_buf0_reg[20]/P0001 ,
		\u4_u2_ienb_reg[4]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w10144_
	);
	LUT4 #(
		.INIT('h0888)
	) name8395 (
		_w2228_,
		_w2240_,
		_w10143_,
		_w10144_,
		_w10145_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name8396 (
		\u4_u0_buf1_reg[20]/P0001 ,
		\u4_u0_csr1_reg[5]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w10146_
	);
	LUT4 #(
		.INIT('hf53f)
	) name8397 (
		\u4_u0_buf0_reg[20]/P0001 ,
		\u4_u0_ienb_reg[4]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w10147_
	);
	LUT4 #(
		.INIT('h0888)
	) name8398 (
		_w2240_,
		_w2241_,
		_w10146_,
		_w10147_,
		_w10148_
	);
	LUT3 #(
		.INIT('h01)
	) name8399 (
		_w10142_,
		_w10145_,
		_w10148_,
		_w10149_
	);
	LUT4 #(
		.INIT('h0200)
	) name8400 (
		\u1_frame_no_r_reg[4]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w10150_
	);
	LUT4 #(
		.INIT('h0020)
	) name8401 (
		\u4_intb_msk_reg[4]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w10151_
	);
	LUT4 #(
		.INIT('h0080)
	) name8402 (
		\u4_int_srcb_reg[0]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w10152_
	);
	LUT4 #(
		.INIT('haaa8)
	) name8403 (
		_w5861_,
		_w10150_,
		_w10151_,
		_w10152_,
		_w10153_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name8404 (
		\u4_u1_buf1_reg[20]/P0001 ,
		\u4_u1_csr1_reg[5]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w10154_
	);
	LUT4 #(
		.INIT('hf53f)
	) name8405 (
		\u4_u1_buf0_reg[20]/P0001 ,
		\u4_u1_ienb_reg[4]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w10155_
	);
	LUT4 #(
		.INIT('h0888)
	) name8406 (
		_w2227_,
		_w2241_,
		_w10154_,
		_w10155_,
		_w10156_
	);
	LUT2 #(
		.INIT('h1)
	) name8407 (
		_w10153_,
		_w10156_,
		_w10157_
	);
	LUT2 #(
		.INIT('h7)
	) name8408 (
		_w10149_,
		_w10157_,
		_w10158_
	);
	LUT3 #(
		.INIT('h07)
	) name8409 (
		\u1_u3_out_to_small_reg/P0001 ,
		\u4_u3_ep_match_r_reg/P0001 ,
		\u4_u3_int_stat_reg[6]/P0001 ,
		_w10159_
	);
	LUT2 #(
		.INIT('h2)
	) name8410 (
		_w3893_,
		_w10159_,
		_w10160_
	);
	LUT4 #(
		.INIT('h0020)
	) name8411 (
		rst_i_pad,
		\u0_u0_state_reg[1]/P0001 ,
		\u0_u0_state_reg[2]/NET0131 ,
		usb_vbus_pad_i_pad,
		_w10161_
	);
	LUT3 #(
		.INIT('h10)
	) name8412 (
		_w4355_,
		_w4356_,
		_w10161_,
		_w10162_
	);
	LUT2 #(
		.INIT('h8)
	) name8413 (
		_w5763_,
		_w10162_,
		_w10163_
	);
	LUT3 #(
		.INIT('hd0)
	) name8414 (
		\u0_u0_T1_gt_3_0_mS_reg/P0001 ,
		\u0_u0_mode_hs_reg/P0001 ,
		\u0_u0_state_reg[2]/NET0131 ,
		_w10164_
	);
	LUT3 #(
		.INIT('h45)
	) name8415 (
		_w4315_,
		_w4316_,
		_w10164_,
		_w10165_
	);
	LUT3 #(
		.INIT('h08)
	) name8416 (
		_w4103_,
		_w4326_,
		_w10165_,
		_w10166_
	);
	LUT2 #(
		.INIT('he)
	) name8417 (
		_w10163_,
		_w10166_,
		_w10167_
	);
	LUT4 #(
		.INIT('hf5f3)
	) name8418 (
		\u4_u3_buf0_reg[5]/P0001 ,
		\u4_u3_csr0_reg[5]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w10168_
	);
	LUT4 #(
		.INIT('h5f3f)
	) name8419 (
		\u4_u3_buf1_reg[5]/P0001 ,
		\u4_u3_int_stat_reg[5]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w10169_
	);
	LUT4 #(
		.INIT('h0888)
	) name8420 (
		_w2227_,
		_w2228_,
		_w10168_,
		_w10169_,
		_w10170_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name8421 (
		\u4_u2_buf1_reg[5]/P0001 ,
		\u4_u2_csr0_reg[5]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w10171_
	);
	LUT4 #(
		.INIT('hf53f)
	) name8422 (
		\u4_u2_buf0_reg[5]/P0001 ,
		\u4_u2_int_stat_reg[5]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w10172_
	);
	LUT4 #(
		.INIT('h0888)
	) name8423 (
		_w2228_,
		_w2240_,
		_w10171_,
		_w10172_,
		_w10173_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name8424 (
		\u4_u0_buf1_reg[5]/P0001 ,
		\u4_u0_csr0_reg[5]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w10174_
	);
	LUT4 #(
		.INIT('hf53f)
	) name8425 (
		\u4_u0_buf0_reg[5]/P0001 ,
		\u4_u0_int_stat_reg[5]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w10175_
	);
	LUT4 #(
		.INIT('h0888)
	) name8426 (
		_w2240_,
		_w2241_,
		_w10174_,
		_w10175_,
		_w10176_
	);
	LUT3 #(
		.INIT('h01)
	) name8427 (
		_w10170_,
		_w10173_,
		_w10176_,
		_w10177_
	);
	LUT4 #(
		.INIT('h0200)
	) name8428 (
		\u1_sof_time_reg[5]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w10178_
	);
	LUT4 #(
		.INIT('h0008)
	) name8429 (
		\u4_funct_adr_reg[5]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w10179_
	);
	LUT4 #(
		.INIT('h0800)
	) name8430 (
		\u4_utmi_vend_stat_r_reg[5]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w10180_
	);
	LUT4 #(
		.INIT('h0020)
	) name8431 (
		\u4_inta_msk_reg[5]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w10181_
	);
	LUT4 #(
		.INIT('h0001)
	) name8432 (
		_w10178_,
		_w10179_,
		_w10180_,
		_w10181_,
		_w10182_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name8433 (
		\u4_u1_buf1_reg[5]/P0001 ,
		\u4_u1_csr0_reg[5]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w10183_
	);
	LUT4 #(
		.INIT('hf53f)
	) name8434 (
		\u4_u1_buf0_reg[5]/P0001 ,
		\u4_u1_int_stat_reg[5]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w10184_
	);
	LUT4 #(
		.INIT('h0888)
	) name8435 (
		_w2227_,
		_w2241_,
		_w10183_,
		_w10184_,
		_w10185_
	);
	LUT3 #(
		.INIT('h0d)
	) name8436 (
		_w5861_,
		_w10182_,
		_w10185_,
		_w10186_
	);
	LUT2 #(
		.INIT('h7)
	) name8437 (
		_w10177_,
		_w10186_,
		_w10187_
	);
	LUT4 #(
		.INIT('hf5f3)
	) name8438 (
		\u4_u3_buf0_reg[6]/P0001 ,
		\u4_u3_csr0_reg[6]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w10188_
	);
	LUT4 #(
		.INIT('h5f3f)
	) name8439 (
		\u4_u3_buf1_reg[6]/P0001 ,
		\u4_u3_int_stat_reg[6]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w10189_
	);
	LUT4 #(
		.INIT('h0888)
	) name8440 (
		_w2227_,
		_w2228_,
		_w10188_,
		_w10189_,
		_w10190_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name8441 (
		\u4_u2_buf1_reg[6]/P0001 ,
		\u4_u2_csr0_reg[6]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w10191_
	);
	LUT4 #(
		.INIT('hf53f)
	) name8442 (
		\u4_u2_buf0_reg[6]/P0001 ,
		\u4_u2_int_stat_reg[6]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w10192_
	);
	LUT4 #(
		.INIT('h0888)
	) name8443 (
		_w2228_,
		_w2240_,
		_w10191_,
		_w10192_,
		_w10193_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name8444 (
		\u4_u0_buf1_reg[6]/P0001 ,
		\u4_u0_csr0_reg[6]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w10194_
	);
	LUT4 #(
		.INIT('hf53f)
	) name8445 (
		\u4_u0_buf0_reg[6]/P0001 ,
		\u4_u0_int_stat_reg[6]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w10195_
	);
	LUT4 #(
		.INIT('h0888)
	) name8446 (
		_w2240_,
		_w2241_,
		_w10194_,
		_w10195_,
		_w10196_
	);
	LUT3 #(
		.INIT('h01)
	) name8447 (
		_w10190_,
		_w10193_,
		_w10196_,
		_w10197_
	);
	LUT4 #(
		.INIT('h0008)
	) name8448 (
		\u4_funct_adr_reg[6]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w10198_
	);
	LUT4 #(
		.INIT('h0200)
	) name8449 (
		\u1_sof_time_reg[6]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w10199_
	);
	LUT4 #(
		.INIT('h0800)
	) name8450 (
		\u4_utmi_vend_stat_r_reg[6]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w10200_
	);
	LUT4 #(
		.INIT('h0020)
	) name8451 (
		\u4_inta_msk_reg[6]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w10201_
	);
	LUT4 #(
		.INIT('h0001)
	) name8452 (
		_w10198_,
		_w10199_,
		_w10200_,
		_w10201_,
		_w10202_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name8453 (
		\u4_u1_buf1_reg[6]/P0001 ,
		\u4_u1_csr0_reg[6]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w10203_
	);
	LUT4 #(
		.INIT('hf53f)
	) name8454 (
		\u4_u1_buf0_reg[6]/P0001 ,
		\u4_u1_int_stat_reg[6]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w10204_
	);
	LUT4 #(
		.INIT('h0888)
	) name8455 (
		_w2227_,
		_w2241_,
		_w10203_,
		_w10204_,
		_w10205_
	);
	LUT3 #(
		.INIT('h0d)
	) name8456 (
		_w5861_,
		_w10202_,
		_w10205_,
		_w10206_
	);
	LUT2 #(
		.INIT('h7)
	) name8457 (
		_w10197_,
		_w10206_,
		_w10207_
	);
	LUT4 #(
		.INIT('h08a8)
	) name8458 (
		rst_i_pad,
		\u5_state_reg[3]/P0001 ,
		\u5_wb_req_s1_reg/P0001 ,
		\wb_addr_i[17]_pad ,
		_w10208_
	);
	LUT3 #(
		.INIT('h80)
	) name8459 (
		_w2224_,
		_w5490_,
		_w10208_,
		_w10209_
	);
	LUT3 #(
		.INIT('hac)
	) name8460 (
		\sram_data_i[14]_pad ,
		\u4_dout_reg[14]/P0001 ,
		\wb_addr_i[17]_pad ,
		_w10210_
	);
	LUT4 #(
		.INIT('h8caf)
	) name8461 (
		\u4_u2_buf0_orig_reg[21]/P0001 ,
		\u4_u2_buf0_orig_reg[22]/P0001 ,
		\u4_u2_dma_out_cnt_reg[2]/P0001 ,
		\u4_u2_dma_out_cnt_reg[3]/P0001 ,
		_w10211_
	);
	LUT2 #(
		.INIT('h9)
	) name8462 (
		\u4_u2_buf0_orig_reg[23]/P0001 ,
		\u4_u2_dma_out_cnt_reg[4]/P0001 ,
		_w10212_
	);
	LUT4 #(
		.INIT('h31c4)
	) name8463 (
		\u4_u2_buf0_orig_reg[22]/P0001 ,
		\u4_u2_buf0_orig_reg[23]/P0001 ,
		\u4_u2_dma_out_cnt_reg[3]/P0001 ,
		\u4_u2_dma_out_cnt_reg[4]/P0001 ,
		_w10213_
	);
	LUT4 #(
		.INIT('h4f00)
	) name8464 (
		_w6028_,
		_w6029_,
		_w10211_,
		_w10213_,
		_w10214_
	);
	LUT4 #(
		.INIT('h0802)
	) name8465 (
		\u4_u2_buf0_orig_reg[22]/P0001 ,
		\u4_u2_buf0_orig_reg[23]/P0001 ,
		\u4_u2_dma_out_cnt_reg[3]/P0001 ,
		\u4_u2_dma_out_cnt_reg[4]/P0001 ,
		_w10215_
	);
	LUT4 #(
		.INIT('hb000)
	) name8466 (
		_w6028_,
		_w6029_,
		_w10211_,
		_w10212_,
		_w10216_
	);
	LUT3 #(
		.INIT('h01)
	) name8467 (
		_w10214_,
		_w10215_,
		_w10216_,
		_w10217_
	);
	LUT4 #(
		.INIT('h8caf)
	) name8468 (
		\u4_u2_buf0_orig_reg[24]/P0001 ,
		\u4_u2_buf0_orig_reg[25]/P0001 ,
		\u4_u2_dma_out_cnt_reg[5]/P0001 ,
		\u4_u2_dma_out_cnt_reg[6]/P0001 ,
		_w10218_
	);
	LUT4 #(
		.INIT('hef00)
	) name8469 (
		_w6027_,
		_w6031_,
		_w6033_,
		_w10218_,
		_w10219_
	);
	LUT2 #(
		.INIT('h9)
	) name8470 (
		\u4_u2_buf0_orig_reg[26]/P0001 ,
		\u4_u2_dma_out_cnt_reg[7]/P0001 ,
		_w10220_
	);
	LUT2 #(
		.INIT('h8)
	) name8471 (
		_w10218_,
		_w10220_,
		_w10221_
	);
	LUT4 #(
		.INIT('hef00)
	) name8472 (
		_w6027_,
		_w6031_,
		_w6033_,
		_w10221_,
		_w10222_
	);
	LUT4 #(
		.INIT('h005e)
	) name8473 (
		_w6024_,
		_w10219_,
		_w10220_,
		_w10222_,
		_w10223_
	);
	LUT4 #(
		.INIT('h8caf)
	) name8474 (
		\u4_u3_buf0_orig_reg[21]/P0001 ,
		\u4_u3_buf0_orig_reg[22]/P0001 ,
		\u4_u3_dma_out_cnt_reg[2]/P0001 ,
		\u4_u3_dma_out_cnt_reg[3]/P0001 ,
		_w10224_
	);
	LUT2 #(
		.INIT('h9)
	) name8475 (
		\u4_u3_buf0_orig_reg[23]/P0001 ,
		\u4_u3_dma_out_cnt_reg[4]/P0001 ,
		_w10225_
	);
	LUT4 #(
		.INIT('h31c4)
	) name8476 (
		\u4_u3_buf0_orig_reg[22]/P0001 ,
		\u4_u3_buf0_orig_reg[23]/P0001 ,
		\u4_u3_dma_out_cnt_reg[3]/P0001 ,
		\u4_u3_dma_out_cnt_reg[4]/P0001 ,
		_w10226_
	);
	LUT4 #(
		.INIT('h4f00)
	) name8477 (
		_w5953_,
		_w5954_,
		_w10224_,
		_w10226_,
		_w10227_
	);
	LUT4 #(
		.INIT('h0802)
	) name8478 (
		\u4_u3_buf0_orig_reg[22]/P0001 ,
		\u4_u3_buf0_orig_reg[23]/P0001 ,
		\u4_u3_dma_out_cnt_reg[3]/P0001 ,
		\u4_u3_dma_out_cnt_reg[4]/P0001 ,
		_w10228_
	);
	LUT4 #(
		.INIT('hb000)
	) name8479 (
		_w5953_,
		_w5954_,
		_w10224_,
		_w10225_,
		_w10229_
	);
	LUT3 #(
		.INIT('h01)
	) name8480 (
		_w10227_,
		_w10228_,
		_w10229_,
		_w10230_
	);
	LUT4 #(
		.INIT('h8caf)
	) name8481 (
		\u4_u3_buf0_orig_reg[24]/P0001 ,
		\u4_u3_buf0_orig_reg[25]/P0001 ,
		\u4_u3_dma_out_cnt_reg[5]/P0001 ,
		\u4_u3_dma_out_cnt_reg[6]/P0001 ,
		_w10231_
	);
	LUT4 #(
		.INIT('hef00)
	) name8482 (
		_w5952_,
		_w5956_,
		_w5958_,
		_w10231_,
		_w10232_
	);
	LUT2 #(
		.INIT('h9)
	) name8483 (
		\u4_u3_buf0_orig_reg[26]/P0001 ,
		\u4_u3_dma_out_cnt_reg[7]/P0001 ,
		_w10233_
	);
	LUT2 #(
		.INIT('h8)
	) name8484 (
		_w10231_,
		_w10233_,
		_w10234_
	);
	LUT4 #(
		.INIT('hef00)
	) name8485 (
		_w5952_,
		_w5956_,
		_w5958_,
		_w10234_,
		_w10235_
	);
	LUT4 #(
		.INIT('h005e)
	) name8486 (
		_w5949_,
		_w10232_,
		_w10233_,
		_w10235_,
		_w10236_
	);
	LUT4 #(
		.INIT('h8caf)
	) name8487 (
		\u4_u0_buf0_orig_reg[21]/P0001 ,
		\u4_u0_buf0_orig_reg[22]/P0001 ,
		\u4_u0_dma_out_cnt_reg[2]/P0001 ,
		\u4_u0_dma_out_cnt_reg[3]/P0001 ,
		_w10237_
	);
	LUT2 #(
		.INIT('h9)
	) name8488 (
		\u4_u0_buf0_orig_reg[23]/P0001 ,
		\u4_u0_dma_out_cnt_reg[4]/P0001 ,
		_w10238_
	);
	LUT4 #(
		.INIT('h31c4)
	) name8489 (
		\u4_u0_buf0_orig_reg[22]/P0001 ,
		\u4_u0_buf0_orig_reg[23]/P0001 ,
		\u4_u0_dma_out_cnt_reg[3]/P0001 ,
		\u4_u0_dma_out_cnt_reg[4]/P0001 ,
		_w10239_
	);
	LUT4 #(
		.INIT('h4f00)
	) name8490 (
		_w5978_,
		_w5979_,
		_w10237_,
		_w10239_,
		_w10240_
	);
	LUT4 #(
		.INIT('h0802)
	) name8491 (
		\u4_u0_buf0_orig_reg[22]/P0001 ,
		\u4_u0_buf0_orig_reg[23]/P0001 ,
		\u4_u0_dma_out_cnt_reg[3]/P0001 ,
		\u4_u0_dma_out_cnt_reg[4]/P0001 ,
		_w10241_
	);
	LUT4 #(
		.INIT('hb000)
	) name8492 (
		_w5978_,
		_w5979_,
		_w10237_,
		_w10238_,
		_w10242_
	);
	LUT3 #(
		.INIT('h01)
	) name8493 (
		_w10240_,
		_w10241_,
		_w10242_,
		_w10243_
	);
	LUT4 #(
		.INIT('h8caf)
	) name8494 (
		\u4_u0_buf0_orig_reg[24]/P0001 ,
		\u4_u0_buf0_orig_reg[25]/P0001 ,
		\u4_u0_dma_out_cnt_reg[5]/P0001 ,
		\u4_u0_dma_out_cnt_reg[6]/P0001 ,
		_w10244_
	);
	LUT4 #(
		.INIT('hef00)
	) name8495 (
		_w5977_,
		_w5981_,
		_w5983_,
		_w10244_,
		_w10245_
	);
	LUT4 #(
		.INIT('h31c4)
	) name8496 (
		\u4_u0_buf0_orig_reg[25]/P0001 ,
		\u4_u0_buf0_orig_reg[26]/P0001 ,
		\u4_u0_dma_out_cnt_reg[6]/P0001 ,
		\u4_u0_dma_out_cnt_reg[7]/P0001 ,
		_w10246_
	);
	LUT4 #(
		.INIT('h8c23)
	) name8497 (
		\u4_u0_buf0_orig_reg[25]/P0001 ,
		\u4_u0_buf0_orig_reg[26]/P0001 ,
		\u4_u0_dma_out_cnt_reg[6]/P0001 ,
		\u4_u0_dma_out_cnt_reg[7]/P0001 ,
		_w10247_
	);
	LUT4 #(
		.INIT('h45cf)
	) name8498 (
		_w5985_,
		_w10245_,
		_w10246_,
		_w10247_,
		_w10248_
	);
	LUT4 #(
		.INIT('h8caf)
	) name8499 (
		\u4_u1_buf0_orig_reg[21]/P0001 ,
		\u4_u1_buf0_orig_reg[22]/P0001 ,
		\u4_u1_dma_out_cnt_reg[2]/P0001 ,
		\u4_u1_dma_out_cnt_reg[3]/P0001 ,
		_w10249_
	);
	LUT2 #(
		.INIT('h9)
	) name8500 (
		\u4_u1_buf0_orig_reg[23]/P0001 ,
		\u4_u1_dma_out_cnt_reg[4]/P0001 ,
		_w10250_
	);
	LUT4 #(
		.INIT('h31c4)
	) name8501 (
		\u4_u1_buf0_orig_reg[22]/P0001 ,
		\u4_u1_buf0_orig_reg[23]/P0001 ,
		\u4_u1_dma_out_cnt_reg[3]/P0001 ,
		\u4_u1_dma_out_cnt_reg[4]/P0001 ,
		_w10251_
	);
	LUT4 #(
		.INIT('h4f00)
	) name8502 (
		_w6003_,
		_w6004_,
		_w10249_,
		_w10251_,
		_w10252_
	);
	LUT4 #(
		.INIT('h0802)
	) name8503 (
		\u4_u1_buf0_orig_reg[22]/P0001 ,
		\u4_u1_buf0_orig_reg[23]/P0001 ,
		\u4_u1_dma_out_cnt_reg[3]/P0001 ,
		\u4_u1_dma_out_cnt_reg[4]/P0001 ,
		_w10253_
	);
	LUT4 #(
		.INIT('hb000)
	) name8504 (
		_w6003_,
		_w6004_,
		_w10249_,
		_w10250_,
		_w10254_
	);
	LUT3 #(
		.INIT('h01)
	) name8505 (
		_w10252_,
		_w10253_,
		_w10254_,
		_w10255_
	);
	LUT4 #(
		.INIT('h8caf)
	) name8506 (
		\u4_u1_buf0_orig_reg[24]/P0001 ,
		\u4_u1_buf0_orig_reg[25]/P0001 ,
		\u4_u1_dma_out_cnt_reg[5]/P0001 ,
		\u4_u1_dma_out_cnt_reg[6]/P0001 ,
		_w10256_
	);
	LUT4 #(
		.INIT('hef00)
	) name8507 (
		_w6002_,
		_w6006_,
		_w6008_,
		_w10256_,
		_w10257_
	);
	LUT2 #(
		.INIT('h9)
	) name8508 (
		\u4_u1_buf0_orig_reg[26]/P0001 ,
		\u4_u1_dma_out_cnt_reg[7]/P0001 ,
		_w10258_
	);
	LUT2 #(
		.INIT('h8)
	) name8509 (
		_w10256_,
		_w10258_,
		_w10259_
	);
	LUT4 #(
		.INIT('hef00)
	) name8510 (
		_w6002_,
		_w6006_,
		_w6008_,
		_w10259_,
		_w10260_
	);
	LUT4 #(
		.INIT('h005e)
	) name8511 (
		_w5999_,
		_w10257_,
		_w10258_,
		_w10260_,
		_w10261_
	);
	LUT4 #(
		.INIT('h0080)
	) name8512 (
		rst_i_pad,
		\u0_tx_ready_reg/NET0131 ,
		\u1_u1_state_reg[2]/NET0131 ,
		\u1_u1_state_reg[4]/NET0131 ,
		_w10262_
	);
	LUT4 #(
		.INIT('h0002)
	) name8513 (
		rst_i_pad,
		\u0_tx_ready_reg/NET0131 ,
		\u1_u1_state_reg[0]/NET0131 ,
		\u1_u1_state_reg[1]/NET0131 ,
		_w10263_
	);
	LUT4 #(
		.INIT('heca0)
	) name8514 (
		_w1807_,
		_w1809_,
		_w10262_,
		_w10263_,
		_w10264_
	);
	LUT4 #(
		.INIT('h0f0e)
	) name8515 (
		\u0_u0_state_reg[3]/P0001 ,
		_w4333_,
		_w9770_,
		_w9773_,
		_w10265_
	);
	LUT3 #(
		.INIT('h02)
	) name8516 (
		\u4_u1_csr0_reg[10]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w10266_
	);
	LUT4 #(
		.INIT('h35ff)
	) name8517 (
		\u4_u1_buf0_reg[10]/P0001 ,
		\u4_u1_buf1_reg[10]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w10267_
	);
	LUT4 #(
		.INIT('h8088)
	) name8518 (
		_w2227_,
		_w2241_,
		_w10266_,
		_w10267_,
		_w10268_
	);
	LUT3 #(
		.INIT('h02)
	) name8519 (
		\u4_u3_csr0_reg[10]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w10269_
	);
	LUT4 #(
		.INIT('h35ff)
	) name8520 (
		\u4_u3_buf0_reg[10]/P0001 ,
		\u4_u3_buf1_reg[10]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w10270_
	);
	LUT4 #(
		.INIT('h8088)
	) name8521 (
		_w2227_,
		_w2228_,
		_w10269_,
		_w10270_,
		_w10271_
	);
	LUT2 #(
		.INIT('h1)
	) name8522 (
		_w10268_,
		_w10271_,
		_w10272_
	);
	LUT4 #(
		.INIT('h0200)
	) name8523 (
		\u1_sof_time_reg[10]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w10273_
	);
	LUT2 #(
		.INIT('h8)
	) name8524 (
		_w5861_,
		_w10273_,
		_w10274_
	);
	LUT3 #(
		.INIT('h02)
	) name8525 (
		\u4_u0_csr0_reg[10]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w10275_
	);
	LUT4 #(
		.INIT('h35ff)
	) name8526 (
		\u4_u0_buf0_reg[10]/P0001 ,
		\u4_u0_buf1_reg[10]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w10276_
	);
	LUT4 #(
		.INIT('h8088)
	) name8527 (
		_w2240_,
		_w2241_,
		_w10275_,
		_w10276_,
		_w10277_
	);
	LUT3 #(
		.INIT('h02)
	) name8528 (
		\u4_u2_csr0_reg[10]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w10278_
	);
	LUT4 #(
		.INIT('h35ff)
	) name8529 (
		\u4_u2_buf0_reg[10]/P0001 ,
		\u4_u2_buf1_reg[10]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w10279_
	);
	LUT4 #(
		.INIT('h8088)
	) name8530 (
		_w2228_,
		_w2240_,
		_w10278_,
		_w10279_,
		_w10280_
	);
	LUT3 #(
		.INIT('h01)
	) name8531 (
		_w10274_,
		_w10277_,
		_w10280_,
		_w10281_
	);
	LUT2 #(
		.INIT('h7)
	) name8532 (
		_w10272_,
		_w10281_,
		_w10282_
	);
	LUT3 #(
		.INIT('h02)
	) name8533 (
		\u4_u1_csr0_reg[11]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w10283_
	);
	LUT4 #(
		.INIT('h35ff)
	) name8534 (
		\u4_u1_buf0_reg[11]/P0001 ,
		\u4_u1_buf1_reg[11]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w10284_
	);
	LUT4 #(
		.INIT('h8088)
	) name8535 (
		_w2227_,
		_w2241_,
		_w10283_,
		_w10284_,
		_w10285_
	);
	LUT3 #(
		.INIT('h02)
	) name8536 (
		\u4_u3_csr0_reg[11]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w10286_
	);
	LUT4 #(
		.INIT('h35ff)
	) name8537 (
		\u4_u3_buf0_reg[11]/P0001 ,
		\u4_u3_buf1_reg[11]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w10287_
	);
	LUT4 #(
		.INIT('h8088)
	) name8538 (
		_w2227_,
		_w2228_,
		_w10286_,
		_w10287_,
		_w10288_
	);
	LUT2 #(
		.INIT('h1)
	) name8539 (
		_w10285_,
		_w10288_,
		_w10289_
	);
	LUT4 #(
		.INIT('h0200)
	) name8540 (
		\u1_sof_time_reg[11]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w10290_
	);
	LUT2 #(
		.INIT('h8)
	) name8541 (
		_w5861_,
		_w10290_,
		_w10291_
	);
	LUT3 #(
		.INIT('h02)
	) name8542 (
		\u4_u0_csr0_reg[11]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w10292_
	);
	LUT4 #(
		.INIT('h35ff)
	) name8543 (
		\u4_u0_buf0_reg[11]/P0001 ,
		\u4_u0_buf1_reg[11]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w10293_
	);
	LUT4 #(
		.INIT('h8088)
	) name8544 (
		_w2240_,
		_w2241_,
		_w10292_,
		_w10293_,
		_w10294_
	);
	LUT3 #(
		.INIT('h02)
	) name8545 (
		\u4_u2_csr0_reg[11]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w10295_
	);
	LUT4 #(
		.INIT('h35ff)
	) name8546 (
		\u4_u2_buf0_reg[11]/P0001 ,
		\u4_u2_buf1_reg[11]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w10296_
	);
	LUT4 #(
		.INIT('h8088)
	) name8547 (
		_w2228_,
		_w2240_,
		_w10295_,
		_w10296_,
		_w10297_
	);
	LUT3 #(
		.INIT('h01)
	) name8548 (
		_w10291_,
		_w10294_,
		_w10297_,
		_w10298_
	);
	LUT2 #(
		.INIT('h7)
	) name8549 (
		_w10289_,
		_w10298_,
		_w10299_
	);
	LUT3 #(
		.INIT('h02)
	) name8550 (
		\u4_u1_csr0_reg[9]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w10300_
	);
	LUT4 #(
		.INIT('h35ff)
	) name8551 (
		\u4_u1_buf0_reg[9]/P0001 ,
		\u4_u1_buf1_reg[9]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w10301_
	);
	LUT4 #(
		.INIT('h8088)
	) name8552 (
		_w2227_,
		_w2241_,
		_w10300_,
		_w10301_,
		_w10302_
	);
	LUT3 #(
		.INIT('h02)
	) name8553 (
		\u4_u3_csr0_reg[9]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w10303_
	);
	LUT4 #(
		.INIT('h35ff)
	) name8554 (
		\u4_u3_buf0_reg[9]/P0001 ,
		\u4_u3_buf1_reg[9]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w10304_
	);
	LUT4 #(
		.INIT('h8088)
	) name8555 (
		_w2227_,
		_w2228_,
		_w10303_,
		_w10304_,
		_w10305_
	);
	LUT2 #(
		.INIT('h1)
	) name8556 (
		_w10302_,
		_w10305_,
		_w10306_
	);
	LUT4 #(
		.INIT('h0200)
	) name8557 (
		\u1_sof_time_reg[9]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w10307_
	);
	LUT2 #(
		.INIT('h8)
	) name8558 (
		_w5861_,
		_w10307_,
		_w10308_
	);
	LUT3 #(
		.INIT('h02)
	) name8559 (
		\u4_u0_csr0_reg[9]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w10309_
	);
	LUT4 #(
		.INIT('h35ff)
	) name8560 (
		\u4_u0_buf0_reg[9]/P0001 ,
		\u4_u0_buf1_reg[9]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w10310_
	);
	LUT4 #(
		.INIT('h8088)
	) name8561 (
		_w2240_,
		_w2241_,
		_w10309_,
		_w10310_,
		_w10311_
	);
	LUT3 #(
		.INIT('h02)
	) name8562 (
		\u4_u2_csr0_reg[9]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w10312_
	);
	LUT4 #(
		.INIT('h35ff)
	) name8563 (
		\u4_u2_buf0_reg[9]/P0001 ,
		\u4_u2_buf1_reg[9]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w10313_
	);
	LUT4 #(
		.INIT('h8088)
	) name8564 (
		_w2228_,
		_w2240_,
		_w10312_,
		_w10313_,
		_w10314_
	);
	LUT3 #(
		.INIT('h01)
	) name8565 (
		_w10308_,
		_w10311_,
		_w10314_,
		_w10315_
	);
	LUT2 #(
		.INIT('h7)
	) name8566 (
		_w10306_,
		_w10315_,
		_w10316_
	);
	LUT2 #(
		.INIT('h8)
	) name8567 (
		\u1_u3_rx_ack_to_cnt_reg[4]/P0001 ,
		\u1_u3_rx_ack_to_cnt_reg[5]/P0001 ,
		_w10317_
	);
	LUT3 #(
		.INIT('h15)
	) name8568 (
		\u1_u3_rx_ack_to_cnt_reg[6]/P0001 ,
		_w7951_,
		_w10317_,
		_w10318_
	);
	LUT3 #(
		.INIT('h15)
	) name8569 (
		\u1_u3_rx_ack_to_clr_reg/P0001 ,
		_w7951_,
		_w8972_,
		_w10319_
	);
	LUT2 #(
		.INIT('h4)
	) name8570 (
		_w10318_,
		_w10319_,
		_w10320_
	);
	LUT2 #(
		.INIT('h8)
	) name8571 (
		\u1_u3_tx_data_to_cnt_reg[4]/P0001 ,
		\u1_u3_tx_data_to_cnt_reg[5]/P0001 ,
		_w10321_
	);
	LUT3 #(
		.INIT('h15)
	) name8572 (
		\u1_u3_tx_data_to_cnt_reg[6]/P0001 ,
		_w7967_,
		_w10321_,
		_w10322_
	);
	LUT3 #(
		.INIT('h15)
	) name8573 (
		\u0_rx_active_reg/P0001 ,
		_w7967_,
		_w8978_,
		_w10323_
	);
	LUT2 #(
		.INIT('h4)
	) name8574 (
		_w10322_,
		_w10323_,
		_w10324_
	);
	LUT3 #(
		.INIT('h0e)
	) name8575 (
		\LineState_r_reg[0]/P0001 ,
		\LineState_r_reg[1]/P0001 ,
		\u0_u0_state_reg[6]/NET0131 ,
		_w10325_
	);
	LUT2 #(
		.INIT('h2)
	) name8576 (
		_w4321_,
		_w10325_,
		_w10326_
	);
	LUT3 #(
		.INIT('h10)
	) name8577 (
		\u0_u0_T2_gt_100_uS_reg/P0001 ,
		\u0_u0_state_reg[3]/P0001 ,
		\u0_u0_state_reg[6]/NET0131 ,
		_w10327_
	);
	LUT4 #(
		.INIT('h135f)
	) name8578 (
		_w4319_,
		_w7962_,
		_w10326_,
		_w10327_,
		_w10328_
	);
	LUT2 #(
		.INIT('h2)
	) name8579 (
		_w4103_,
		_w10328_,
		_w10329_
	);
	LUT4 #(
		.INIT('hf807)
	) name8580 (
		\u4_u3_buf0_orig_reg[19]/P0001 ,
		\u4_u3_buf0_orig_reg[20]/P0001 ,
		\u4_u3_buf0_orig_reg[21]/P0001 ,
		\u4_u3_buf0_orig_reg[22]/P0001 ,
		_w10330_
	);
	LUT2 #(
		.INIT('h2)
	) name8581 (
		\u5_wb_req_s1_reg/P0001 ,
		wb_we_i_pad,
		_w10331_
	);
	LUT3 #(
		.INIT('h08)
	) name8582 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w10332_
	);
	LUT4 #(
		.INIT('h8000)
	) name8583 (
		_w2224_,
		_w2226_,
		_w5861_,
		_w10332_,
		_w10333_
	);
	LUT2 #(
		.INIT('h8)
	) name8584 (
		_w10331_,
		_w10333_,
		_w10334_
	);
	LUT4 #(
		.INIT('hf807)
	) name8585 (
		\u4_u0_buf0_orig_reg[19]/P0001 ,
		\u4_u0_buf0_orig_reg[20]/P0001 ,
		\u4_u0_buf0_orig_reg[21]/P0001 ,
		\u4_u0_buf0_orig_reg[22]/P0001 ,
		_w10335_
	);
	LUT4 #(
		.INIT('hf807)
	) name8586 (
		\u4_u1_buf0_orig_reg[19]/P0001 ,
		\u4_u1_buf0_orig_reg[20]/P0001 ,
		\u4_u1_buf0_orig_reg[21]/P0001 ,
		\u4_u1_buf0_orig_reg[22]/P0001 ,
		_w10336_
	);
	LUT4 #(
		.INIT('hf807)
	) name8587 (
		\u4_u2_buf0_orig_reg[19]/P0001 ,
		\u4_u2_buf0_orig_reg[20]/P0001 ,
		\u4_u2_buf0_orig_reg[21]/P0001 ,
		\u4_u2_buf0_orig_reg[22]/P0001 ,
		_w10337_
	);
	LUT4 #(
		.INIT('h7f80)
	) name8588 (
		\u0_u0_idle_cnt1_reg[0]/P0001 ,
		\u0_u0_idle_cnt1_reg[1]/P0001 ,
		\u0_u0_idle_cnt1_reg[2]/P0001 ,
		\u0_u0_idle_cnt1_reg[3]/P0001 ,
		_w10338_
	);
	LUT2 #(
		.INIT('h9)
	) name8589 (
		\u4_u1_buf0_orig_reg[24]/P0001 ,
		\u4_u1_dma_out_cnt_reg[5]/P0001 ,
		_w10339_
	);
	LUT4 #(
		.INIT('h01fe)
	) name8590 (
		_w6002_,
		_w6006_,
		_w6007_,
		_w10339_,
		_w10340_
	);
	LUT2 #(
		.INIT('h9)
	) name8591 (
		\u4_u3_buf0_orig_reg[24]/P0001 ,
		\u4_u3_dma_out_cnt_reg[5]/P0001 ,
		_w10341_
	);
	LUT4 #(
		.INIT('h01fe)
	) name8592 (
		_w5952_,
		_w5956_,
		_w5957_,
		_w10341_,
		_w10342_
	);
	LUT2 #(
		.INIT('h9)
	) name8593 (
		\u4_u0_buf0_orig_reg[24]/P0001 ,
		\u4_u0_dma_out_cnt_reg[5]/P0001 ,
		_w10343_
	);
	LUT4 #(
		.INIT('h01fe)
	) name8594 (
		_w5977_,
		_w5981_,
		_w5982_,
		_w10343_,
		_w10344_
	);
	LUT2 #(
		.INIT('h9)
	) name8595 (
		\u4_u2_buf0_orig_reg[24]/P0001 ,
		\u4_u2_dma_out_cnt_reg[5]/P0001 ,
		_w10345_
	);
	LUT4 #(
		.INIT('h01fe)
	) name8596 (
		_w6027_,
		_w6031_,
		_w6032_,
		_w10345_,
		_w10346_
	);
	LUT3 #(
		.INIT('h80)
	) name8597 (
		\u4_buf0_reg[11]/P0001 ,
		\u4_buf0_reg[13]/P0001 ,
		\u4_buf0_reg[14]/P0001 ,
		_w10347_
	);
	LUT3 #(
		.INIT('h80)
	) name8598 (
		\u4_buf0_reg[0]/P0001 ,
		\u4_buf0_reg[10]/P0001 ,
		\u4_buf0_reg[12]/P0001 ,
		_w10348_
	);
	LUT2 #(
		.INIT('h8)
	) name8599 (
		_w10347_,
		_w10348_,
		_w10349_
	);
	LUT4 #(
		.INIT('h8000)
	) name8600 (
		\u4_buf0_reg[3]/P0001 ,
		\u4_buf0_reg[4]/P0001 ,
		\u4_buf0_reg[5]/P0001 ,
		\u4_buf0_reg[6]/P0001 ,
		_w10350_
	);
	LUT4 #(
		.INIT('h8000)
	) name8601 (
		\u4_buf0_reg[15]/P0001 ,
		\u4_buf0_reg[16]/P0001 ,
		\u4_buf0_reg[1]/P0001 ,
		\u4_buf0_reg[2]/P0001 ,
		_w10351_
	);
	LUT3 #(
		.INIT('h80)
	) name8602 (
		\u4_buf0_reg[7]/P0001 ,
		\u4_buf0_reg[8]/P0001 ,
		\u4_buf0_reg[9]/P0001 ,
		_w10352_
	);
	LUT3 #(
		.INIT('h80)
	) name8603 (
		_w10350_,
		_w10351_,
		_w10352_,
		_w10353_
	);
	LUT2 #(
		.INIT('h8)
	) name8604 (
		_w10349_,
		_w10353_,
		_w10354_
	);
	LUT3 #(
		.INIT('hea)
	) name8605 (
		\u4_buf0_reg[31]/P0001 ,
		_w10349_,
		_w10353_,
		_w10355_
	);
	LUT3 #(
		.INIT('h80)
	) name8606 (
		\u4_buf1_reg[11]/P0001 ,
		\u4_buf1_reg[13]/P0001 ,
		\u4_buf1_reg[14]/P0001 ,
		_w10356_
	);
	LUT3 #(
		.INIT('h80)
	) name8607 (
		\u4_buf1_reg[0]/P0001 ,
		\u4_buf1_reg[10]/P0001 ,
		\u4_buf1_reg[12]/P0001 ,
		_w10357_
	);
	LUT2 #(
		.INIT('h8)
	) name8608 (
		_w10356_,
		_w10357_,
		_w10358_
	);
	LUT4 #(
		.INIT('h8000)
	) name8609 (
		\u4_buf1_reg[3]/P0001 ,
		\u4_buf1_reg[4]/P0001 ,
		\u4_buf1_reg[5]/P0001 ,
		\u4_buf1_reg[6]/P0001 ,
		_w10359_
	);
	LUT4 #(
		.INIT('h8000)
	) name8610 (
		\u4_buf1_reg[15]/P0001 ,
		\u4_buf1_reg[16]/P0001 ,
		\u4_buf1_reg[1]/P0001 ,
		\u4_buf1_reg[2]/P0001 ,
		_w10360_
	);
	LUT3 #(
		.INIT('h80)
	) name8611 (
		\u4_buf1_reg[7]/P0001 ,
		\u4_buf1_reg[8]/P0001 ,
		\u4_buf1_reg[9]/P0001 ,
		_w10361_
	);
	LUT3 #(
		.INIT('h80)
	) name8612 (
		_w10359_,
		_w10360_,
		_w10361_,
		_w10362_
	);
	LUT2 #(
		.INIT('h8)
	) name8613 (
		_w10358_,
		_w10362_,
		_w10363_
	);
	LUT3 #(
		.INIT('hea)
	) name8614 (
		\u4_buf1_reg[31]/P0001 ,
		_w10358_,
		_w10362_,
		_w10364_
	);
	LUT3 #(
		.INIT('h01)
	) name8615 (
		\u1_u0_state_reg[1]/P0001 ,
		\u1_u0_state_reg[2]/P0001 ,
		\u1_u0_state_reg[3]/P0001 ,
		_w10365_
	);
	LUT3 #(
		.INIT('h20)
	) name8616 (
		\u0_rx_active_reg/P0001 ,
		\u0_rx_data_reg[0]/P0001 ,
		\u0_rx_valid_reg/P0001 ,
		_w10366_
	);
	LUT2 #(
		.INIT('h8)
	) name8617 (
		rst_i_pad,
		\u1_u0_pid_reg[0]/NET0131 ,
		_w10367_
	);
	LUT3 #(
		.INIT('h80)
	) name8618 (
		rst_i_pad,
		\u0_rx_active_reg/P0001 ,
		\u0_rx_valid_reg/P0001 ,
		_w10368_
	);
	LUT4 #(
		.INIT('h7270)
	) name8619 (
		_w10365_,
		_w10366_,
		_w10367_,
		_w10368_,
		_w10369_
	);
	LUT3 #(
		.INIT('h20)
	) name8620 (
		\u0_rx_active_reg/P0001 ,
		\u0_rx_data_reg[1]/P0001 ,
		\u0_rx_valid_reg/P0001 ,
		_w10370_
	);
	LUT2 #(
		.INIT('h8)
	) name8621 (
		rst_i_pad,
		\u1_u0_pid_reg[1]/NET0131 ,
		_w10371_
	);
	LUT4 #(
		.INIT('h5f08)
	) name8622 (
		_w10365_,
		_w10368_,
		_w10370_,
		_w10371_,
		_w10372_
	);
	LUT3 #(
		.INIT('h20)
	) name8623 (
		\u0_rx_active_reg/P0001 ,
		\u0_rx_data_reg[2]/P0001 ,
		\u0_rx_valid_reg/P0001 ,
		_w10373_
	);
	LUT2 #(
		.INIT('h8)
	) name8624 (
		rst_i_pad,
		\u1_u0_pid_reg[2]/NET0131 ,
		_w10374_
	);
	LUT4 #(
		.INIT('h5f08)
	) name8625 (
		_w10365_,
		_w10368_,
		_w10373_,
		_w10374_,
		_w10375_
	);
	LUT3 #(
		.INIT('h20)
	) name8626 (
		\u0_rx_active_reg/P0001 ,
		\u0_rx_data_reg[3]/P0001 ,
		\u0_rx_valid_reg/P0001 ,
		_w10376_
	);
	LUT2 #(
		.INIT('h8)
	) name8627 (
		rst_i_pad,
		\u1_u0_pid_reg[3]/NET0131 ,
		_w10377_
	);
	LUT4 #(
		.INIT('h5f08)
	) name8628 (
		_w10365_,
		_w10368_,
		_w10376_,
		_w10377_,
		_w10378_
	);
	LUT3 #(
		.INIT('h02)
	) name8629 (
		\u4_u0_csr0_reg[12]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w10379_
	);
	LUT4 #(
		.INIT('h35ff)
	) name8630 (
		\u4_u0_buf0_reg[12]/P0001 ,
		\u4_u0_buf1_reg[12]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w10380_
	);
	LUT4 #(
		.INIT('h8088)
	) name8631 (
		_w2240_,
		_w2241_,
		_w10379_,
		_w10380_,
		_w10381_
	);
	LUT3 #(
		.INIT('h02)
	) name8632 (
		\u4_u3_csr0_reg[12]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w10382_
	);
	LUT4 #(
		.INIT('h35ff)
	) name8633 (
		\u4_u3_buf0_reg[12]/P0001 ,
		\u4_u3_buf1_reg[12]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w10383_
	);
	LUT4 #(
		.INIT('h8088)
	) name8634 (
		_w2227_,
		_w2228_,
		_w10382_,
		_w10383_,
		_w10384_
	);
	LUT3 #(
		.INIT('h02)
	) name8635 (
		\u4_u2_csr0_reg[12]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w10385_
	);
	LUT4 #(
		.INIT('h35ff)
	) name8636 (
		\u4_u2_buf0_reg[12]/P0001 ,
		\u4_u2_buf1_reg[12]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w10386_
	);
	LUT4 #(
		.INIT('h8088)
	) name8637 (
		_w2228_,
		_w2240_,
		_w10385_,
		_w10386_,
		_w10387_
	);
	LUT3 #(
		.INIT('h02)
	) name8638 (
		\u4_u1_csr0_reg[12]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w10388_
	);
	LUT4 #(
		.INIT('h35ff)
	) name8639 (
		\u4_u1_buf0_reg[12]/P0001 ,
		\u4_u1_buf1_reg[12]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w10389_
	);
	LUT4 #(
		.INIT('h8088)
	) name8640 (
		_w2227_,
		_w2241_,
		_w10388_,
		_w10389_,
		_w10390_
	);
	LUT4 #(
		.INIT('hfffe)
	) name8641 (
		_w10381_,
		_w10384_,
		_w10387_,
		_w10390_,
		_w10391_
	);
	LUT3 #(
		.INIT('h02)
	) name8642 (
		\u4_u2_ots_stop_reg/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w10392_
	);
	LUT4 #(
		.INIT('h35ff)
	) name8643 (
		\u4_u2_buf0_reg[13]/P0001 ,
		\u4_u2_buf1_reg[13]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w10393_
	);
	LUT4 #(
		.INIT('h8088)
	) name8644 (
		_w2228_,
		_w2240_,
		_w10392_,
		_w10393_,
		_w10394_
	);
	LUT3 #(
		.INIT('h02)
	) name8645 (
		\u4_u0_ots_stop_reg/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w10395_
	);
	LUT4 #(
		.INIT('h35ff)
	) name8646 (
		\u4_u0_buf0_reg[13]/P0001 ,
		\u4_u0_buf1_reg[13]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w10396_
	);
	LUT4 #(
		.INIT('h8088)
	) name8647 (
		_w2240_,
		_w2241_,
		_w10395_,
		_w10396_,
		_w10397_
	);
	LUT3 #(
		.INIT('h02)
	) name8648 (
		\u4_u3_ots_stop_reg/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w10398_
	);
	LUT4 #(
		.INIT('h35ff)
	) name8649 (
		\u4_u3_buf0_reg[13]/P0001 ,
		\u4_u3_buf1_reg[13]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w10399_
	);
	LUT4 #(
		.INIT('h8088)
	) name8650 (
		_w2227_,
		_w2228_,
		_w10398_,
		_w10399_,
		_w10400_
	);
	LUT3 #(
		.INIT('h02)
	) name8651 (
		\u4_u1_ots_stop_reg/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w10401_
	);
	LUT4 #(
		.INIT('h35ff)
	) name8652 (
		\u4_u1_buf0_reg[13]/P0001 ,
		\u4_u1_buf1_reg[13]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w10402_
	);
	LUT4 #(
		.INIT('h8088)
	) name8653 (
		_w2227_,
		_w2241_,
		_w10401_,
		_w10402_,
		_w10403_
	);
	LUT4 #(
		.INIT('hfffe)
	) name8654 (
		_w10394_,
		_w10397_,
		_w10400_,
		_w10403_,
		_w10404_
	);
	LUT3 #(
		.INIT('h02)
	) name8655 (
		\u4_u2_csr1_reg[0]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w10405_
	);
	LUT4 #(
		.INIT('h35ff)
	) name8656 (
		\u4_u2_buf0_reg[15]/P0001 ,
		\u4_u2_buf1_reg[15]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w10406_
	);
	LUT4 #(
		.INIT('h8088)
	) name8657 (
		_w2228_,
		_w2240_,
		_w10405_,
		_w10406_,
		_w10407_
	);
	LUT3 #(
		.INIT('h02)
	) name8658 (
		\u4_u0_csr1_reg[0]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w10408_
	);
	LUT4 #(
		.INIT('h35ff)
	) name8659 (
		\u4_u0_buf0_reg[15]/P0001 ,
		\u4_u0_buf1_reg[15]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w10409_
	);
	LUT4 #(
		.INIT('h8088)
	) name8660 (
		_w2240_,
		_w2241_,
		_w10408_,
		_w10409_,
		_w10410_
	);
	LUT3 #(
		.INIT('h02)
	) name8661 (
		\u4_u3_csr1_reg[0]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w10411_
	);
	LUT4 #(
		.INIT('h35ff)
	) name8662 (
		\u4_u3_buf0_reg[15]/P0001 ,
		\u4_u3_buf1_reg[15]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w10412_
	);
	LUT4 #(
		.INIT('h8088)
	) name8663 (
		_w2227_,
		_w2228_,
		_w10411_,
		_w10412_,
		_w10413_
	);
	LUT3 #(
		.INIT('h02)
	) name8664 (
		\u4_u1_csr1_reg[0]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w10414_
	);
	LUT4 #(
		.INIT('h35ff)
	) name8665 (
		\u4_u1_buf0_reg[15]/P0001 ,
		\u4_u1_buf1_reg[15]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w10415_
	);
	LUT4 #(
		.INIT('h8088)
	) name8666 (
		_w2227_,
		_w2241_,
		_w10414_,
		_w10415_,
		_w10416_
	);
	LUT4 #(
		.INIT('hfffe)
	) name8667 (
		_w10407_,
		_w10410_,
		_w10413_,
		_w10416_,
		_w10417_
	);
	LUT4 #(
		.INIT('h1450)
	) name8668 (
		\u1_u3_rx_ack_to_clr_reg/P0001 ,
		\u1_u3_rx_ack_to_cnt_reg[4]/P0001 ,
		\u1_u3_rx_ack_to_cnt_reg[5]/P0001 ,
		_w7951_,
		_w10418_
	);
	LUT3 #(
		.INIT('h2a)
	) name8669 (
		\u1_u0_pid_reg[4]/P0001 ,
		_w4883_,
		_w10365_,
		_w10419_
	);
	LUT3 #(
		.INIT('h80)
	) name8670 (
		\u0_rx_active_reg/P0001 ,
		\u0_rx_data_reg[4]/P0001 ,
		\u0_rx_valid_reg/P0001 ,
		_w10420_
	);
	LUT3 #(
		.INIT('h2a)
	) name8671 (
		rst_i_pad,
		_w10365_,
		_w10420_,
		_w10421_
	);
	LUT2 #(
		.INIT('hb)
	) name8672 (
		_w10419_,
		_w10421_,
		_w10422_
	);
	LUT3 #(
		.INIT('h2a)
	) name8673 (
		\u1_u0_pid_reg[5]/P0001 ,
		_w4883_,
		_w10365_,
		_w10423_
	);
	LUT3 #(
		.INIT('h80)
	) name8674 (
		\u0_rx_active_reg/P0001 ,
		\u0_rx_data_reg[5]/P0001 ,
		\u0_rx_valid_reg/P0001 ,
		_w10424_
	);
	LUT3 #(
		.INIT('h2a)
	) name8675 (
		rst_i_pad,
		_w10365_,
		_w10424_,
		_w10425_
	);
	LUT2 #(
		.INIT('hb)
	) name8676 (
		_w10423_,
		_w10425_,
		_w10426_
	);
	LUT3 #(
		.INIT('h2a)
	) name8677 (
		\u1_u0_pid_reg[6]/P0001 ,
		_w4883_,
		_w10365_,
		_w10427_
	);
	LUT3 #(
		.INIT('h80)
	) name8678 (
		\u0_rx_active_reg/P0001 ,
		\u0_rx_data_reg[6]/P0001 ,
		\u0_rx_valid_reg/P0001 ,
		_w10428_
	);
	LUT3 #(
		.INIT('h2a)
	) name8679 (
		rst_i_pad,
		_w10365_,
		_w10428_,
		_w10429_
	);
	LUT2 #(
		.INIT('hb)
	) name8680 (
		_w10427_,
		_w10429_,
		_w10430_
	);
	LUT3 #(
		.INIT('h2a)
	) name8681 (
		\u1_u0_pid_reg[7]/P0001 ,
		_w4883_,
		_w10365_,
		_w10431_
	);
	LUT3 #(
		.INIT('h80)
	) name8682 (
		\u0_rx_active_reg/P0001 ,
		\u0_rx_data_reg[7]/P0001 ,
		\u0_rx_valid_reg/P0001 ,
		_w10432_
	);
	LUT3 #(
		.INIT('h2a)
	) name8683 (
		rst_i_pad,
		_w10365_,
		_w10432_,
		_w10433_
	);
	LUT2 #(
		.INIT('hb)
	) name8684 (
		_w10431_,
		_w10433_,
		_w10434_
	);
	LUT4 #(
		.INIT('hdccc)
	) name8685 (
		\u0_rx_err_reg/P0001 ,
		\u1_u0_token_valid_r1_reg/P0001 ,
		_w3695_,
		_w4881_,
		_w10435_
	);
	LUT4 #(
		.INIT('h0008)
	) name8686 (
		\u5_wb_req_s1_reg/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		wb_we_i_pad,
		_w10436_
	);
	LUT3 #(
		.INIT('h80)
	) name8687 (
		_w2224_,
		_w2226_,
		_w10436_,
		_w10437_
	);
	LUT2 #(
		.INIT('h8)
	) name8688 (
		_w5839_,
		_w10437_,
		_w10438_
	);
	LUT4 #(
		.INIT('h1540)
	) name8689 (
		\u1_u3_rx_ack_to_clr_reg/P0001 ,
		\u1_u3_rx_ack_to_cnt_reg[0]/P0001 ,
		\u1_u3_rx_ack_to_cnt_reg[1]/P0001 ,
		\u1_u3_rx_ack_to_cnt_reg[2]/P0001 ,
		_w10439_
	);
	LUT4 #(
		.INIT('h1540)
	) name8690 (
		\u0_rx_active_reg/P0001 ,
		\u1_u3_tx_data_to_cnt_reg[0]/P0001 ,
		\u1_u3_tx_data_to_cnt_reg[1]/P0001 ,
		\u1_u3_tx_data_to_cnt_reg[2]/P0001 ,
		_w10440_
	);
	LUT4 #(
		.INIT('h1450)
	) name8691 (
		\u0_rx_active_reg/P0001 ,
		\u1_u3_tx_data_to_cnt_reg[4]/P0001 ,
		\u1_u3_tx_data_to_cnt_reg[5]/P0001 ,
		_w7967_,
		_w10441_
	);
	LUT2 #(
		.INIT('h8)
	) name8692 (
		_w5862_,
		_w10437_,
		_w10442_
	);
	LUT2 #(
		.INIT('he)
	) name8693 (
		\u4_u0_inta_reg/P0001 ,
		\u4_u0_intb_reg/P0001 ,
		_w10443_
	);
	LUT2 #(
		.INIT('he)
	) name8694 (
		\u4_u1_inta_reg/P0001 ,
		\u4_u1_intb_reg/P0001 ,
		_w10444_
	);
	LUT2 #(
		.INIT('he)
	) name8695 (
		\u4_u2_inta_reg/P0001 ,
		\u4_u2_intb_reg/P0001 ,
		_w10445_
	);
	LUT2 #(
		.INIT('he)
	) name8696 (
		\u4_u3_inta_reg/P0001 ,
		\u4_u3_intb_reg/P0001 ,
		_w10446_
	);
	LUT2 #(
		.INIT('h8)
	) name8697 (
		_w5844_,
		_w10437_,
		_w10447_
	);
	LUT2 #(
		.INIT('h4)
	) name8698 (
		\u0_u0_me_ps2_0_5_ms_reg/P0001 ,
		\u0_u0_me_ps2_reg[3]/P0001 ,
		_w10448_
	);
	LUT3 #(
		.INIT('h01)
	) name8699 (
		\u0_u0_me_ps2_reg[0]/P0001 ,
		\u0_u0_me_ps2_reg[1]/P0001 ,
		\u0_u0_me_ps2_reg[2]/P0001 ,
		_w10449_
	);
	LUT4 #(
		.INIT('h1000)
	) name8700 (
		\u0_u0_me_ps2_reg[4]/P0001 ,
		\u0_u0_me_ps2_reg[5]/P0001 ,
		\u0_u0_me_ps2_reg[6]/P0001 ,
		\u0_u0_me_ps2_reg[7]/P0001 ,
		_w10450_
	);
	LUT3 #(
		.INIT('h80)
	) name8701 (
		_w10448_,
		_w10449_,
		_w10450_,
		_w10451_
	);
	LUT4 #(
		.INIT('h9ccc)
	) name8702 (
		\u4_u3_buf0_orig_reg[27]/P0001 ,
		\u4_u3_buf0_orig_reg[28]/P0001 ,
		_w7822_,
		_w7824_,
		_w10452_
	);
	LUT4 #(
		.INIT('h9ccc)
	) name8703 (
		\u4_u1_buf0_orig_reg[27]/P0001 ,
		\u4_u1_buf0_orig_reg[28]/P0001 ,
		_w7845_,
		_w7847_,
		_w10453_
	);
	LUT4 #(
		.INIT('h9ccc)
	) name8704 (
		\u4_u0_buf0_orig_reg[27]/P0001 ,
		\u4_u0_buf0_orig_reg[28]/P0001 ,
		_w7833_,
		_w7835_,
		_w10454_
	);
	LUT3 #(
		.INIT('h6a)
	) name8705 (
		\u0_u0_idle_cnt1_reg[6]/P0001 ,
		_w8152_,
		_w9015_,
		_w10455_
	);
	LUT4 #(
		.INIT('h9ccc)
	) name8706 (
		\u4_u2_buf0_orig_reg[27]/P0001 ,
		\u4_u2_buf0_orig_reg[28]/P0001 ,
		_w7853_,
		_w7855_,
		_w10456_
	);
	LUT4 #(
		.INIT('h7310)
	) name8707 (
		\u4_u3_buf0_orig_reg[19]/P0001 ,
		\u4_u3_buf0_orig_reg[20]/P0001 ,
		\u4_u3_dma_in_cnt_reg[0]/P0001 ,
		\u4_u3_dma_out_cnt_reg[1]/P0001 ,
		_w10457_
	);
	LUT2 #(
		.INIT('h9)
	) name8708 (
		\u4_u3_buf0_orig_reg[21]/P0001 ,
		\u4_u3_dma_out_cnt_reg[2]/P0001 ,
		_w10458_
	);
	LUT2 #(
		.INIT('h9)
	) name8709 (
		_w10457_,
		_w10458_,
		_w10459_
	);
	LUT2 #(
		.INIT('h9)
	) name8710 (
		\u4_u3_buf0_orig_reg[22]/P0001 ,
		\u4_u3_dma_out_cnt_reg[3]/P0001 ,
		_w10460_
	);
	LUT4 #(
		.INIT('hf40b)
	) name8711 (
		_w5953_,
		_w5954_,
		_w5955_,
		_w10460_,
		_w10461_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name8712 (
		\u4_u2_buf0_orig_reg[29]/NET0131 ,
		_w7853_,
		_w7855_,
		_w7856_,
		_w10462_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name8713 (
		\u4_u0_buf0_orig_reg[29]/NET0131 ,
		_w7833_,
		_w7835_,
		_w7839_,
		_w10463_
	);
	LUT2 #(
		.INIT('he)
	) name8714 (
		_w7837_,
		_w10463_,
		_w10464_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name8715 (
		\u4_u3_buf0_orig_reg[29]/NET0131 ,
		_w7822_,
		_w7824_,
		_w7825_,
		_w10465_
	);
	LUT4 #(
		.INIT('h7310)
	) name8716 (
		\u4_u0_buf0_orig_reg[19]/P0001 ,
		\u4_u0_buf0_orig_reg[20]/P0001 ,
		\u4_u0_dma_in_cnt_reg[0]/P0001 ,
		\u4_u0_dma_out_cnt_reg[1]/P0001 ,
		_w10466_
	);
	LUT2 #(
		.INIT('h9)
	) name8717 (
		\u4_u0_buf0_orig_reg[21]/P0001 ,
		\u4_u0_dma_out_cnt_reg[2]/P0001 ,
		_w10467_
	);
	LUT2 #(
		.INIT('h9)
	) name8718 (
		_w10466_,
		_w10467_,
		_w10468_
	);
	LUT2 #(
		.INIT('h9)
	) name8719 (
		\u4_u0_buf0_orig_reg[22]/P0001 ,
		\u4_u0_dma_out_cnt_reg[3]/P0001 ,
		_w10469_
	);
	LUT4 #(
		.INIT('hf40b)
	) name8720 (
		_w5978_,
		_w5979_,
		_w5980_,
		_w10469_,
		_w10470_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name8721 (
		\u4_u1_buf0_orig_reg[29]/NET0131 ,
		_w7845_,
		_w7847_,
		_w7848_,
		_w10471_
	);
	LUT4 #(
		.INIT('h7310)
	) name8722 (
		\u4_u1_buf0_orig_reg[19]/P0001 ,
		\u4_u1_buf0_orig_reg[20]/P0001 ,
		\u4_u1_dma_in_cnt_reg[0]/P0001 ,
		\u4_u1_dma_out_cnt_reg[1]/P0001 ,
		_w10472_
	);
	LUT2 #(
		.INIT('h9)
	) name8723 (
		\u4_u1_buf0_orig_reg[21]/P0001 ,
		\u4_u1_dma_out_cnt_reg[2]/P0001 ,
		_w10473_
	);
	LUT2 #(
		.INIT('h9)
	) name8724 (
		_w10472_,
		_w10473_,
		_w10474_
	);
	LUT2 #(
		.INIT('h9)
	) name8725 (
		\u4_u1_buf0_orig_reg[22]/P0001 ,
		\u4_u1_dma_out_cnt_reg[3]/P0001 ,
		_w10475_
	);
	LUT4 #(
		.INIT('hf40b)
	) name8726 (
		_w6003_,
		_w6004_,
		_w6005_,
		_w10475_,
		_w10476_
	);
	LUT4 #(
		.INIT('h7310)
	) name8727 (
		\u4_u2_buf0_orig_reg[19]/P0001 ,
		\u4_u2_buf0_orig_reg[20]/P0001 ,
		\u4_u2_dma_in_cnt_reg[0]/P0001 ,
		\u4_u2_dma_out_cnt_reg[1]/P0001 ,
		_w10477_
	);
	LUT2 #(
		.INIT('h9)
	) name8728 (
		\u4_u2_buf0_orig_reg[21]/P0001 ,
		\u4_u2_dma_out_cnt_reg[2]/P0001 ,
		_w10478_
	);
	LUT2 #(
		.INIT('h9)
	) name8729 (
		_w10477_,
		_w10478_,
		_w10479_
	);
	LUT2 #(
		.INIT('h9)
	) name8730 (
		\u4_u2_buf0_orig_reg[22]/P0001 ,
		\u4_u2_dma_out_cnt_reg[3]/P0001 ,
		_w10480_
	);
	LUT4 #(
		.INIT('hf40b)
	) name8731 (
		_w6028_,
		_w6029_,
		_w6030_,
		_w10480_,
		_w10481_
	);
	LUT4 #(
		.INIT('h0008)
	) name8732 (
		\u1_u3_in_token_reg/NET0131 ,
		\u4_buf1_reg[0]/P0001 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		_w10482_
	);
	LUT3 #(
		.INIT('hc8)
	) name8733 (
		\u1_u3_buf0_na_reg/NET0131 ,
		\u4_buf1_reg[0]/P0001 ,
		\u4_csr_reg[30]/NET0131 ,
		_w10483_
	);
	LUT3 #(
		.INIT('h13)
	) name8734 (
		_w2352_,
		_w10482_,
		_w10483_,
		_w10484_
	);
	LUT4 #(
		.INIT('hccc4)
	) name8735 (
		\u1_u3_in_token_reg/NET0131 ,
		\u4_buf0_reg[0]/P0001 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		_w10485_
	);
	LUT3 #(
		.INIT('hd0)
	) name8736 (
		_w2352_,
		_w2353_,
		_w10485_,
		_w10486_
	);
	LUT2 #(
		.INIT('hd)
	) name8737 (
		_w10484_,
		_w10486_,
		_w10487_
	);
	LUT4 #(
		.INIT('h0008)
	) name8738 (
		\u1_u3_in_token_reg/NET0131 ,
		\u4_buf1_reg[10]/P0001 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		_w10488_
	);
	LUT3 #(
		.INIT('hc8)
	) name8739 (
		\u1_u3_buf0_na_reg/NET0131 ,
		\u4_buf1_reg[10]/P0001 ,
		\u4_csr_reg[30]/NET0131 ,
		_w10489_
	);
	LUT3 #(
		.INIT('h13)
	) name8740 (
		_w2352_,
		_w10488_,
		_w10489_,
		_w10490_
	);
	LUT4 #(
		.INIT('hccc4)
	) name8741 (
		\u1_u3_in_token_reg/NET0131 ,
		\u4_buf0_reg[10]/P0001 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		_w10491_
	);
	LUT3 #(
		.INIT('hd0)
	) name8742 (
		_w2352_,
		_w2353_,
		_w10491_,
		_w10492_
	);
	LUT2 #(
		.INIT('hd)
	) name8743 (
		_w10490_,
		_w10492_,
		_w10493_
	);
	LUT4 #(
		.INIT('h0008)
	) name8744 (
		\u1_u3_in_token_reg/NET0131 ,
		\u4_buf1_reg[11]/P0001 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		_w10494_
	);
	LUT3 #(
		.INIT('hc8)
	) name8745 (
		\u1_u3_buf0_na_reg/NET0131 ,
		\u4_buf1_reg[11]/P0001 ,
		\u4_csr_reg[30]/NET0131 ,
		_w10495_
	);
	LUT3 #(
		.INIT('h13)
	) name8746 (
		_w2352_,
		_w10494_,
		_w10495_,
		_w10496_
	);
	LUT4 #(
		.INIT('hccc4)
	) name8747 (
		\u1_u3_in_token_reg/NET0131 ,
		\u4_buf0_reg[11]/P0001 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		_w10497_
	);
	LUT3 #(
		.INIT('hd0)
	) name8748 (
		_w2352_,
		_w2353_,
		_w10497_,
		_w10498_
	);
	LUT2 #(
		.INIT('hd)
	) name8749 (
		_w10496_,
		_w10498_,
		_w10499_
	);
	LUT4 #(
		.INIT('h0008)
	) name8750 (
		\u1_u3_in_token_reg/NET0131 ,
		\u4_buf1_reg[12]/P0001 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		_w10500_
	);
	LUT3 #(
		.INIT('hc8)
	) name8751 (
		\u1_u3_buf0_na_reg/NET0131 ,
		\u4_buf1_reg[12]/P0001 ,
		\u4_csr_reg[30]/NET0131 ,
		_w10501_
	);
	LUT3 #(
		.INIT('h13)
	) name8752 (
		_w2352_,
		_w10500_,
		_w10501_,
		_w10502_
	);
	LUT4 #(
		.INIT('hccc4)
	) name8753 (
		\u1_u3_in_token_reg/NET0131 ,
		\u4_buf0_reg[12]/P0001 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		_w10503_
	);
	LUT3 #(
		.INIT('hd0)
	) name8754 (
		_w2352_,
		_w2353_,
		_w10503_,
		_w10504_
	);
	LUT2 #(
		.INIT('hd)
	) name8755 (
		_w10502_,
		_w10504_,
		_w10505_
	);
	LUT4 #(
		.INIT('h0008)
	) name8756 (
		\u1_u3_in_token_reg/NET0131 ,
		\u4_buf1_reg[13]/P0001 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		_w10506_
	);
	LUT3 #(
		.INIT('hc8)
	) name8757 (
		\u1_u3_buf0_na_reg/NET0131 ,
		\u4_buf1_reg[13]/P0001 ,
		\u4_csr_reg[30]/NET0131 ,
		_w10507_
	);
	LUT3 #(
		.INIT('h13)
	) name8758 (
		_w2352_,
		_w10506_,
		_w10507_,
		_w10508_
	);
	LUT4 #(
		.INIT('hccc4)
	) name8759 (
		\u1_u3_in_token_reg/NET0131 ,
		\u4_buf0_reg[13]/P0001 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		_w10509_
	);
	LUT3 #(
		.INIT('hd0)
	) name8760 (
		_w2352_,
		_w2353_,
		_w10509_,
		_w10510_
	);
	LUT2 #(
		.INIT('hd)
	) name8761 (
		_w10508_,
		_w10510_,
		_w10511_
	);
	LUT4 #(
		.INIT('h0008)
	) name8762 (
		\u1_u3_in_token_reg/NET0131 ,
		\u4_buf1_reg[14]/P0001 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		_w10512_
	);
	LUT3 #(
		.INIT('hc8)
	) name8763 (
		\u1_u3_buf0_na_reg/NET0131 ,
		\u4_buf1_reg[14]/P0001 ,
		\u4_csr_reg[30]/NET0131 ,
		_w10513_
	);
	LUT3 #(
		.INIT('h13)
	) name8764 (
		_w2352_,
		_w10512_,
		_w10513_,
		_w10514_
	);
	LUT4 #(
		.INIT('hccc4)
	) name8765 (
		\u1_u3_in_token_reg/NET0131 ,
		\u4_buf0_reg[14]/P0001 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		_w10515_
	);
	LUT3 #(
		.INIT('hd0)
	) name8766 (
		_w2352_,
		_w2353_,
		_w10515_,
		_w10516_
	);
	LUT2 #(
		.INIT('hd)
	) name8767 (
		_w10514_,
		_w10516_,
		_w10517_
	);
	LUT4 #(
		.INIT('h0008)
	) name8768 (
		\u1_u3_in_token_reg/NET0131 ,
		\u4_buf1_reg[16]/P0001 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		_w10518_
	);
	LUT3 #(
		.INIT('hc8)
	) name8769 (
		\u1_u3_buf0_na_reg/NET0131 ,
		\u4_buf1_reg[16]/P0001 ,
		\u4_csr_reg[30]/NET0131 ,
		_w10519_
	);
	LUT3 #(
		.INIT('h13)
	) name8770 (
		_w2352_,
		_w10518_,
		_w10519_,
		_w10520_
	);
	LUT4 #(
		.INIT('hccc4)
	) name8771 (
		\u1_u3_in_token_reg/NET0131 ,
		\u4_buf0_reg[16]/P0001 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		_w10521_
	);
	LUT3 #(
		.INIT('hd0)
	) name8772 (
		_w2352_,
		_w2353_,
		_w10521_,
		_w10522_
	);
	LUT2 #(
		.INIT('hd)
	) name8773 (
		_w10520_,
		_w10522_,
		_w10523_
	);
	LUT4 #(
		.INIT('h0008)
	) name8774 (
		\u1_u3_in_token_reg/NET0131 ,
		\u4_buf1_reg[1]/P0001 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		_w10524_
	);
	LUT3 #(
		.INIT('hc8)
	) name8775 (
		\u1_u3_buf0_na_reg/NET0131 ,
		\u4_buf1_reg[1]/P0001 ,
		\u4_csr_reg[30]/NET0131 ,
		_w10525_
	);
	LUT3 #(
		.INIT('h13)
	) name8776 (
		_w2352_,
		_w10524_,
		_w10525_,
		_w10526_
	);
	LUT4 #(
		.INIT('hccc4)
	) name8777 (
		\u1_u3_in_token_reg/NET0131 ,
		\u4_buf0_reg[1]/P0001 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		_w10527_
	);
	LUT3 #(
		.INIT('hd0)
	) name8778 (
		_w2352_,
		_w2353_,
		_w10527_,
		_w10528_
	);
	LUT2 #(
		.INIT('hd)
	) name8779 (
		_w10526_,
		_w10528_,
		_w10529_
	);
	LUT4 #(
		.INIT('h0008)
	) name8780 (
		\u1_u3_in_token_reg/NET0131 ,
		\u4_buf1_reg[2]/P0001 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		_w10530_
	);
	LUT3 #(
		.INIT('hc8)
	) name8781 (
		\u1_u3_buf0_na_reg/NET0131 ,
		\u4_buf1_reg[2]/P0001 ,
		\u4_csr_reg[30]/NET0131 ,
		_w10531_
	);
	LUT3 #(
		.INIT('h13)
	) name8782 (
		_w2352_,
		_w10530_,
		_w10531_,
		_w10532_
	);
	LUT4 #(
		.INIT('hccc4)
	) name8783 (
		\u1_u3_in_token_reg/NET0131 ,
		\u4_buf0_reg[2]/P0001 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		_w10533_
	);
	LUT3 #(
		.INIT('hd0)
	) name8784 (
		_w2352_,
		_w2353_,
		_w10533_,
		_w10534_
	);
	LUT2 #(
		.INIT('hd)
	) name8785 (
		_w10532_,
		_w10534_,
		_w10535_
	);
	LUT4 #(
		.INIT('h0008)
	) name8786 (
		\u1_u3_in_token_reg/NET0131 ,
		\u4_buf1_reg[3]/P0001 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		_w10536_
	);
	LUT3 #(
		.INIT('hc8)
	) name8787 (
		\u1_u3_buf0_na_reg/NET0131 ,
		\u4_buf1_reg[3]/P0001 ,
		\u4_csr_reg[30]/NET0131 ,
		_w10537_
	);
	LUT3 #(
		.INIT('h13)
	) name8788 (
		_w2352_,
		_w10536_,
		_w10537_,
		_w10538_
	);
	LUT4 #(
		.INIT('hccc4)
	) name8789 (
		\u1_u3_in_token_reg/NET0131 ,
		\u4_buf0_reg[3]/P0001 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		_w10539_
	);
	LUT3 #(
		.INIT('hd0)
	) name8790 (
		_w2352_,
		_w2353_,
		_w10539_,
		_w10540_
	);
	LUT2 #(
		.INIT('hd)
	) name8791 (
		_w10538_,
		_w10540_,
		_w10541_
	);
	LUT4 #(
		.INIT('h0008)
	) name8792 (
		\u1_u3_in_token_reg/NET0131 ,
		\u4_buf1_reg[4]/P0001 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		_w10542_
	);
	LUT3 #(
		.INIT('hc8)
	) name8793 (
		\u1_u3_buf0_na_reg/NET0131 ,
		\u4_buf1_reg[4]/P0001 ,
		\u4_csr_reg[30]/NET0131 ,
		_w10543_
	);
	LUT3 #(
		.INIT('h13)
	) name8794 (
		_w2352_,
		_w10542_,
		_w10543_,
		_w10544_
	);
	LUT4 #(
		.INIT('hccc4)
	) name8795 (
		\u1_u3_in_token_reg/NET0131 ,
		\u4_buf0_reg[4]/P0001 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		_w10545_
	);
	LUT3 #(
		.INIT('hd0)
	) name8796 (
		_w2352_,
		_w2353_,
		_w10545_,
		_w10546_
	);
	LUT2 #(
		.INIT('hd)
	) name8797 (
		_w10544_,
		_w10546_,
		_w10547_
	);
	LUT4 #(
		.INIT('h0008)
	) name8798 (
		\u1_u3_in_token_reg/NET0131 ,
		\u4_buf1_reg[5]/P0001 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		_w10548_
	);
	LUT3 #(
		.INIT('hc8)
	) name8799 (
		\u1_u3_buf0_na_reg/NET0131 ,
		\u4_buf1_reg[5]/P0001 ,
		\u4_csr_reg[30]/NET0131 ,
		_w10549_
	);
	LUT3 #(
		.INIT('h13)
	) name8800 (
		_w2352_,
		_w10548_,
		_w10549_,
		_w10550_
	);
	LUT4 #(
		.INIT('hccc4)
	) name8801 (
		\u1_u3_in_token_reg/NET0131 ,
		\u4_buf0_reg[5]/P0001 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		_w10551_
	);
	LUT3 #(
		.INIT('hd0)
	) name8802 (
		_w2352_,
		_w2353_,
		_w10551_,
		_w10552_
	);
	LUT2 #(
		.INIT('hd)
	) name8803 (
		_w10550_,
		_w10552_,
		_w10553_
	);
	LUT4 #(
		.INIT('h0008)
	) name8804 (
		\u1_u3_in_token_reg/NET0131 ,
		\u4_buf1_reg[6]/P0001 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		_w10554_
	);
	LUT3 #(
		.INIT('hc8)
	) name8805 (
		\u1_u3_buf0_na_reg/NET0131 ,
		\u4_buf1_reg[6]/P0001 ,
		\u4_csr_reg[30]/NET0131 ,
		_w10555_
	);
	LUT3 #(
		.INIT('h13)
	) name8806 (
		_w2352_,
		_w10554_,
		_w10555_,
		_w10556_
	);
	LUT4 #(
		.INIT('hccc4)
	) name8807 (
		\u1_u3_in_token_reg/NET0131 ,
		\u4_buf0_reg[6]/P0001 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		_w10557_
	);
	LUT3 #(
		.INIT('hd0)
	) name8808 (
		_w2352_,
		_w2353_,
		_w10557_,
		_w10558_
	);
	LUT2 #(
		.INIT('hd)
	) name8809 (
		_w10556_,
		_w10558_,
		_w10559_
	);
	LUT4 #(
		.INIT('h0008)
	) name8810 (
		\u1_u3_in_token_reg/NET0131 ,
		\u4_buf1_reg[7]/P0001 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		_w10560_
	);
	LUT3 #(
		.INIT('hc8)
	) name8811 (
		\u1_u3_buf0_na_reg/NET0131 ,
		\u4_buf1_reg[7]/P0001 ,
		\u4_csr_reg[30]/NET0131 ,
		_w10561_
	);
	LUT3 #(
		.INIT('h13)
	) name8812 (
		_w2352_,
		_w10560_,
		_w10561_,
		_w10562_
	);
	LUT4 #(
		.INIT('hccc4)
	) name8813 (
		\u1_u3_in_token_reg/NET0131 ,
		\u4_buf0_reg[7]/P0001 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		_w10563_
	);
	LUT3 #(
		.INIT('hd0)
	) name8814 (
		_w2352_,
		_w2353_,
		_w10563_,
		_w10564_
	);
	LUT2 #(
		.INIT('hd)
	) name8815 (
		_w10562_,
		_w10564_,
		_w10565_
	);
	LUT4 #(
		.INIT('h0008)
	) name8816 (
		\u1_u3_in_token_reg/NET0131 ,
		\u4_buf1_reg[8]/P0001 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		_w10566_
	);
	LUT3 #(
		.INIT('hc8)
	) name8817 (
		\u1_u3_buf0_na_reg/NET0131 ,
		\u4_buf1_reg[8]/P0001 ,
		\u4_csr_reg[30]/NET0131 ,
		_w10567_
	);
	LUT3 #(
		.INIT('h13)
	) name8818 (
		_w2352_,
		_w10566_,
		_w10567_,
		_w10568_
	);
	LUT4 #(
		.INIT('hccc4)
	) name8819 (
		\u1_u3_in_token_reg/NET0131 ,
		\u4_buf0_reg[8]/P0001 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		_w10569_
	);
	LUT3 #(
		.INIT('hd0)
	) name8820 (
		_w2352_,
		_w2353_,
		_w10569_,
		_w10570_
	);
	LUT2 #(
		.INIT('hd)
	) name8821 (
		_w10568_,
		_w10570_,
		_w10571_
	);
	LUT4 #(
		.INIT('h0008)
	) name8822 (
		\u1_u3_in_token_reg/NET0131 ,
		\u4_buf1_reg[9]/P0001 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		_w10572_
	);
	LUT3 #(
		.INIT('hc8)
	) name8823 (
		\u1_u3_buf0_na_reg/NET0131 ,
		\u4_buf1_reg[9]/P0001 ,
		\u4_csr_reg[30]/NET0131 ,
		_w10573_
	);
	LUT3 #(
		.INIT('h13)
	) name8824 (
		_w2352_,
		_w10572_,
		_w10573_,
		_w10574_
	);
	LUT4 #(
		.INIT('hccc4)
	) name8825 (
		\u1_u3_in_token_reg/NET0131 ,
		\u4_buf0_reg[9]/P0001 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		_w10575_
	);
	LUT3 #(
		.INIT('hd0)
	) name8826 (
		_w2352_,
		_w2353_,
		_w10575_,
		_w10576_
	);
	LUT2 #(
		.INIT('hd)
	) name8827 (
		_w10574_,
		_w10576_,
		_w10577_
	);
	LUT4 #(
		.INIT('h0008)
	) name8828 (
		\u1_u3_in_token_reg/NET0131 ,
		\u4_buf1_reg[15]/P0001 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		_w10578_
	);
	LUT3 #(
		.INIT('hc8)
	) name8829 (
		\u1_u3_buf0_na_reg/NET0131 ,
		\u4_buf1_reg[15]/P0001 ,
		\u4_csr_reg[30]/NET0131 ,
		_w10579_
	);
	LUT3 #(
		.INIT('h13)
	) name8830 (
		_w2352_,
		_w10578_,
		_w10579_,
		_w10580_
	);
	LUT4 #(
		.INIT('hccc4)
	) name8831 (
		\u1_u3_in_token_reg/NET0131 ,
		\u4_buf0_reg[15]/P0001 ,
		\u4_csr_reg[26]/NET0131 ,
		\u4_csr_reg[27]/NET0131 ,
		_w10581_
	);
	LUT3 #(
		.INIT('hd0)
	) name8832 (
		_w2352_,
		_w2353_,
		_w10581_,
		_w10582_
	);
	LUT2 #(
		.INIT('hd)
	) name8833 (
		_w10580_,
		_w10582_,
		_w10583_
	);
	LUT3 #(
		.INIT('h0d)
	) name8834 (
		\u1_u0_pid_reg[0]/NET0131 ,
		\u1_u0_pid_reg[1]/NET0131 ,
		\u1_u3_in_token_reg/NET0131 ,
		_w10584_
	);
	LUT3 #(
		.INIT('ha2)
	) name8835 (
		rst_i_pad,
		\u1_u0_pid_reg[2]/NET0131 ,
		\u1_u3_in_token_reg/NET0131 ,
		_w10585_
	);
	LUT4 #(
		.INIT('h0100)
	) name8836 (
		_w3721_,
		_w10584_,
		_w2116_,
		_w10585_,
		_w10586_
	);
	LUT4 #(
		.INIT('h8000)
	) name8837 (
		_w4093_,
		_w4098_,
		_w4101_,
		_w4331_,
		_w10587_
	);
	LUT3 #(
		.INIT('h07)
	) name8838 (
		\u0_u0_me_cnt_100_ms_reg/P0001 ,
		\u0_u0_state_reg[8]/NET0131 ,
		\u0_u0_usb_attached_reg/P0001 ,
		_w10588_
	);
	LUT2 #(
		.INIT('h1)
	) name8839 (
		_w10587_,
		_w10588_,
		_w10589_
	);
	LUT4 #(
		.INIT('hfe7f)
	) name8840 (
		\u0_u0_mode_hs_reg/P0001 ,
		\u1_u3_rx_ack_to_cnt_reg[1]/P0001 ,
		\u1_u3_rx_ack_to_cnt_reg[4]/P0001 ,
		\u1_u3_rx_ack_to_cnt_reg[5]/P0001 ,
		_w10590_
	);
	LUT4 #(
		.INIT('h0004)
	) name8841 (
		\u1_u3_rx_ack_to_cnt_reg[0]/P0001 ,
		\u1_u3_rx_ack_to_cnt_reg[2]/P0001 ,
		\u1_u3_rx_ack_to_cnt_reg[3]/P0001 ,
		\u1_u3_rx_ack_to_cnt_reg[6]/P0001 ,
		_w10591_
	);
	LUT3 #(
		.INIT('h10)
	) name8842 (
		\u1_u3_rx_ack_to_cnt_reg[7]/P0001 ,
		_w10590_,
		_w10591_,
		_w10592_
	);
	LUT4 #(
		.INIT('hfe7f)
	) name8843 (
		\u0_u0_mode_hs_reg/P0001 ,
		\u1_u3_tx_data_to_cnt_reg[1]/P0001 ,
		\u1_u3_tx_data_to_cnt_reg[4]/P0001 ,
		\u1_u3_tx_data_to_cnt_reg[5]/P0001 ,
		_w10593_
	);
	LUT4 #(
		.INIT('h0004)
	) name8844 (
		\u1_u3_tx_data_to_cnt_reg[0]/P0001 ,
		\u1_u3_tx_data_to_cnt_reg[2]/P0001 ,
		\u1_u3_tx_data_to_cnt_reg[3]/P0001 ,
		\u1_u3_tx_data_to_cnt_reg[6]/P0001 ,
		_w10594_
	);
	LUT3 #(
		.INIT('h10)
	) name8845 (
		\u1_u3_tx_data_to_cnt_reg[7]/P0001 ,
		_w10593_,
		_w10594_,
		_w10595_
	);
	LUT4 #(
		.INIT('h0200)
	) name8846 (
		\u0_u0_me_ps_reg[4]/P0001 ,
		\u0_u0_me_ps_reg[5]/P0001 ,
		\u0_u0_me_ps_reg[6]/P0001 ,
		\u0_u0_me_ps_reg[7]/P0001 ,
		_w10596_
	);
	LUT4 #(
		.INIT('h0010)
	) name8847 (
		\u0_u0_me_ps_reg[0]/P0001 ,
		\u0_u0_me_ps_reg[1]/P0001 ,
		\u0_u0_me_ps_reg[2]/P0001 ,
		\u0_u0_me_ps_reg[3]/P0001 ,
		_w10597_
	);
	LUT2 #(
		.INIT('h8)
	) name8848 (
		_w10596_,
		_w10597_,
		_w10598_
	);
	LUT2 #(
		.INIT('h8)
	) name8849 (
		_w2357_,
		_w3420_,
		_w10599_
	);
	LUT2 #(
		.INIT('h4)
	) name8850 (
		_w2357_,
		_w3420_,
		_w10600_
	);
	LUT3 #(
		.INIT('h02)
	) name8851 (
		\u1_u0_pid_reg[0]/NET0131 ,
		\u1_u0_pid_reg[1]/NET0131 ,
		\u1_u0_pid_reg[2]/NET0131 ,
		_w10601_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name8852 (
		rst_i_pad,
		\u1_u3_setup_token_reg/P0001 ,
		_w3721_,
		_w10601_,
		_w10602_
	);
	LUT4 #(
		.INIT('h35ff)
	) name8853 (
		\u4_u2_buf0_reg[14]/P0001 ,
		\u4_u2_buf1_reg[14]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w10603_
	);
	LUT3 #(
		.INIT('h08)
	) name8854 (
		_w2228_,
		_w2240_,
		_w10603_,
		_w10604_
	);
	LUT4 #(
		.INIT('h35ff)
	) name8855 (
		\u4_u3_buf0_reg[14]/P0001 ,
		\u4_u3_buf1_reg[14]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w10605_
	);
	LUT3 #(
		.INIT('h08)
	) name8856 (
		_w2227_,
		_w2228_,
		_w10605_,
		_w10606_
	);
	LUT4 #(
		.INIT('h35ff)
	) name8857 (
		\u4_u1_buf0_reg[14]/P0001 ,
		\u4_u1_buf1_reg[14]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w10607_
	);
	LUT3 #(
		.INIT('h08)
	) name8858 (
		_w2227_,
		_w2241_,
		_w10607_,
		_w10608_
	);
	LUT4 #(
		.INIT('h35ff)
	) name8859 (
		\u4_u0_buf0_reg[14]/P0001 ,
		\u4_u0_buf1_reg[14]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w10609_
	);
	LUT3 #(
		.INIT('h08)
	) name8860 (
		_w2240_,
		_w2241_,
		_w10609_,
		_w10610_
	);
	LUT4 #(
		.INIT('hfffe)
	) name8861 (
		_w10604_,
		_w10606_,
		_w10608_,
		_w10610_,
		_w10611_
	);
	LUT3 #(
		.INIT('h01)
	) name8862 (
		\u1_u2_sizd_c_reg[0]/P0001 ,
		\u1_u2_sizd_c_reg[10]/P0001 ,
		\u1_u2_sizd_c_reg[11]/P0001 ,
		_w10612_
	);
	LUT4 #(
		.INIT('h8000)
	) name8863 (
		_w2750_,
		_w2753_,
		_w2756_,
		_w10612_,
		_w10613_
	);
	LUT2 #(
		.INIT('he)
	) name8864 (
		\u1_u2_rx_data_done_r_reg/P0001 ,
		_w10613_,
		_w10614_
	);
	LUT2 #(
		.INIT('h8)
	) name8865 (
		_w5848_,
		_w10437_,
		_w10615_
	);
	LUT3 #(
		.INIT('h9c)
	) name8866 (
		\u4_u3_buf0_orig_reg[23]/P0001 ,
		\u4_u3_buf0_orig_reg[24]/P0001 ,
		_w7822_,
		_w10616_
	);
	LUT3 #(
		.INIT('h6a)
	) name8867 (
		\u4_u1_buf0_orig_reg[25]/P0001 ,
		_w7845_,
		_w7846_,
		_w10617_
	);
	LUT3 #(
		.INIT('h9c)
	) name8868 (
		\u4_u0_buf0_orig_reg[23]/P0001 ,
		\u4_u0_buf0_orig_reg[24]/P0001 ,
		_w7835_,
		_w10618_
	);
	LUT3 #(
		.INIT('h6a)
	) name8869 (
		\u4_u0_buf0_orig_reg[25]/P0001 ,
		_w7832_,
		_w7835_,
		_w10619_
	);
	LUT3 #(
		.INIT('h6a)
	) name8870 (
		\u4_u3_buf0_orig_reg[25]/P0001 ,
		_w7822_,
		_w7823_,
		_w10620_
	);
	LUT3 #(
		.INIT('h9c)
	) name8871 (
		\u4_u1_buf0_orig_reg[23]/P0001 ,
		\u4_u1_buf0_orig_reg[24]/P0001 ,
		_w7845_,
		_w10621_
	);
	LUT3 #(
		.INIT('h9c)
	) name8872 (
		\u4_u2_buf0_orig_reg[23]/P0001 ,
		\u4_u2_buf0_orig_reg[24]/P0001 ,
		_w7853_,
		_w10622_
	);
	LUT3 #(
		.INIT('h6a)
	) name8873 (
		\u4_u2_buf0_orig_reg[25]/P0001 ,
		_w7853_,
		_w7854_,
		_w10623_
	);
	LUT3 #(
		.INIT('h87)
	) name8874 (
		\u4_u0_buf0_orig_reg[19]/P0001 ,
		\u4_u0_buf0_orig_reg[20]/P0001 ,
		\u4_u0_buf0_orig_reg[21]/P0001 ,
		_w10624_
	);
	LUT3 #(
		.INIT('h87)
	) name8875 (
		\u4_u1_buf0_orig_reg[19]/P0001 ,
		\u4_u1_buf0_orig_reg[20]/P0001 ,
		\u4_u1_buf0_orig_reg[21]/P0001 ,
		_w10625_
	);
	LUT3 #(
		.INIT('h87)
	) name8876 (
		\u4_u2_buf0_orig_reg[19]/P0001 ,
		\u4_u2_buf0_orig_reg[20]/P0001 ,
		\u4_u2_buf0_orig_reg[21]/P0001 ,
		_w10626_
	);
	LUT3 #(
		.INIT('h87)
	) name8877 (
		\u4_u3_buf0_orig_reg[19]/P0001 ,
		\u4_u3_buf0_orig_reg[20]/P0001 ,
		\u4_u3_buf0_orig_reg[21]/P0001 ,
		_w10627_
	);
	LUT4 #(
		.INIT('h08aa)
	) name8878 (
		rst_i_pad,
		\u1_u3_out_token_reg/NET0131 ,
		_w2115_,
		_w3722_,
		_w10628_
	);
	LUT2 #(
		.INIT('h1)
	) name8879 (
		\u0_u0_mode_hs_reg/P0001 ,
		\u0_u0_state_reg[13]/NET0131 ,
		_w10629_
	);
	LUT4 #(
		.INIT('h0001)
	) name8880 (
		\u0_u0_state_reg[10]/P0001 ,
		\u0_u0_state_reg[13]/NET0131 ,
		\u0_u0_state_reg[7]/NET0131 ,
		\u0_u0_state_reg[8]/NET0131 ,
		_w10630_
	);
	LUT4 #(
		.INIT('h070f)
	) name8881 (
		_w4098_,
		_w4101_,
		_w10629_,
		_w10630_,
		_w10631_
	);
	LUT4 #(
		.INIT('h0400)
	) name8882 (
		\u0_u0_idle_cnt1_reg[0]/P0001 ,
		\u0_u0_idle_cnt1_reg[1]/P0001 ,
		\u0_u0_idle_cnt1_reg[2]/P0001 ,
		\u0_u0_idle_cnt1_reg[3]/P0001 ,
		_w10632_
	);
	LUT2 #(
		.INIT('h8)
	) name8883 (
		_w9803_,
		_w10632_,
		_w10633_
	);
	LUT2 #(
		.INIT('h8)
	) name8884 (
		\u4_u3_iena_reg[5]/P0001 ,
		\u4_u3_int_stat_reg[6]/P0001 ,
		_w10634_
	);
	LUT4 #(
		.INIT('h135f)
	) name8885 (
		\u4_u3_iena_reg[1]/P0001 ,
		\u4_u3_iena_reg[2]/P0001 ,
		\u4_u3_int_stat_reg[1]/P0001 ,
		\u4_u3_int_stat_reg[2]/P0001 ,
		_w10635_
	);
	LUT4 #(
		.INIT('h135f)
	) name8886 (
		\u4_u3_iena_reg[0]/P0001 ,
		\u4_u3_iena_reg[4]/P0001 ,
		\u4_u3_int_stat_reg[0]/P0001 ,
		\u4_u3_int_stat_reg[5]/P0001 ,
		_w10636_
	);
	LUT3 #(
		.INIT('ha8)
	) name8887 (
		\u4_u3_iena_reg[3]/P0001 ,
		\u4_u3_int_stat_reg[3]/P0001 ,
		\u4_u3_int_stat_reg[4]/P0001 ,
		_w10637_
	);
	LUT4 #(
		.INIT('hffbf)
	) name8888 (
		_w10634_,
		_w10635_,
		_w10636_,
		_w10637_,
		_w10638_
	);
	LUT2 #(
		.INIT('h8)
	) name8889 (
		\u4_u3_ienb_reg[1]/P0001 ,
		\u4_u3_int_stat_reg[1]/P0001 ,
		_w10639_
	);
	LUT4 #(
		.INIT('h135f)
	) name8890 (
		\u4_u3_ienb_reg[0]/P0001 ,
		\u4_u3_ienb_reg[2]/P0001 ,
		\u4_u3_int_stat_reg[0]/P0001 ,
		\u4_u3_int_stat_reg[2]/P0001 ,
		_w10640_
	);
	LUT3 #(
		.INIT('ha8)
	) name8891 (
		\u4_u3_ienb_reg[3]/P0001 ,
		\u4_u3_int_stat_reg[3]/P0001 ,
		\u4_u3_int_stat_reg[4]/P0001 ,
		_w10641_
	);
	LUT4 #(
		.INIT('h135f)
	) name8892 (
		\u4_u3_ienb_reg[4]/P0001 ,
		\u4_u3_ienb_reg[5]/P0001 ,
		\u4_u3_int_stat_reg[5]/P0001 ,
		\u4_u3_int_stat_reg[6]/P0001 ,
		_w10642_
	);
	LUT4 #(
		.INIT('hfbff)
	) name8893 (
		_w10639_,
		_w10640_,
		_w10641_,
		_w10642_,
		_w10643_
	);
	LUT2 #(
		.INIT('h8)
	) name8894 (
		\u4_u0_ienb_reg[5]/P0001 ,
		\u4_u0_int_stat_reg[6]/P0001 ,
		_w10644_
	);
	LUT4 #(
		.INIT('h135f)
	) name8895 (
		\u4_u0_ienb_reg[1]/P0001 ,
		\u4_u0_ienb_reg[4]/P0001 ,
		\u4_u0_int_stat_reg[1]/P0001 ,
		\u4_u0_int_stat_reg[5]/P0001 ,
		_w10645_
	);
	LUT4 #(
		.INIT('h135f)
	) name8896 (
		\u4_u0_ienb_reg[0]/P0001 ,
		\u4_u0_ienb_reg[2]/P0001 ,
		\u4_u0_int_stat_reg[0]/P0001 ,
		\u4_u0_int_stat_reg[2]/P0001 ,
		_w10646_
	);
	LUT3 #(
		.INIT('ha8)
	) name8897 (
		\u4_u0_ienb_reg[3]/P0001 ,
		\u4_u0_int_stat_reg[3]/P0001 ,
		\u4_u0_int_stat_reg[4]/P0001 ,
		_w10647_
	);
	LUT4 #(
		.INIT('hffbf)
	) name8898 (
		_w10644_,
		_w10645_,
		_w10646_,
		_w10647_,
		_w10648_
	);
	LUT2 #(
		.INIT('h8)
	) name8899 (
		\u4_u0_iena_reg[5]/P0001 ,
		\u4_u0_int_stat_reg[6]/P0001 ,
		_w10649_
	);
	LUT4 #(
		.INIT('h135f)
	) name8900 (
		\u4_u0_iena_reg[0]/P0001 ,
		\u4_u0_iena_reg[1]/P0001 ,
		\u4_u0_int_stat_reg[0]/P0001 ,
		\u4_u0_int_stat_reg[1]/P0001 ,
		_w10650_
	);
	LUT3 #(
		.INIT('ha8)
	) name8901 (
		\u4_u0_iena_reg[3]/P0001 ,
		\u4_u0_int_stat_reg[3]/P0001 ,
		\u4_u0_int_stat_reg[4]/P0001 ,
		_w10651_
	);
	LUT4 #(
		.INIT('h135f)
	) name8902 (
		\u4_u0_iena_reg[2]/P0001 ,
		\u4_u0_iena_reg[4]/P0001 ,
		\u4_u0_int_stat_reg[2]/P0001 ,
		\u4_u0_int_stat_reg[5]/P0001 ,
		_w10652_
	);
	LUT4 #(
		.INIT('hfbff)
	) name8903 (
		_w10649_,
		_w10650_,
		_w10651_,
		_w10652_,
		_w10653_
	);
	LUT2 #(
		.INIT('h8)
	) name8904 (
		\u4_u1_iena_reg[5]/P0001 ,
		\u4_u1_int_stat_reg[6]/P0001 ,
		_w10654_
	);
	LUT4 #(
		.INIT('h135f)
	) name8905 (
		\u4_u1_iena_reg[1]/P0001 ,
		\u4_u1_iena_reg[2]/P0001 ,
		\u4_u1_int_stat_reg[1]/P0001 ,
		\u4_u1_int_stat_reg[2]/P0001 ,
		_w10655_
	);
	LUT4 #(
		.INIT('h135f)
	) name8906 (
		\u4_u1_iena_reg[0]/P0001 ,
		\u4_u1_iena_reg[4]/P0001 ,
		\u4_u1_int_stat_reg[0]/P0001 ,
		\u4_u1_int_stat_reg[5]/P0001 ,
		_w10656_
	);
	LUT3 #(
		.INIT('ha8)
	) name8907 (
		\u4_u1_iena_reg[3]/P0001 ,
		\u4_u1_int_stat_reg[3]/P0001 ,
		\u4_u1_int_stat_reg[4]/P0001 ,
		_w10657_
	);
	LUT4 #(
		.INIT('hffbf)
	) name8908 (
		_w10654_,
		_w10655_,
		_w10656_,
		_w10657_,
		_w10658_
	);
	LUT2 #(
		.INIT('h8)
	) name8909 (
		\u4_u1_ienb_reg[5]/P0001 ,
		\u4_u1_int_stat_reg[6]/P0001 ,
		_w10659_
	);
	LUT4 #(
		.INIT('h135f)
	) name8910 (
		\u4_u1_ienb_reg[0]/P0001 ,
		\u4_u1_ienb_reg[1]/P0001 ,
		\u4_u1_int_stat_reg[0]/P0001 ,
		\u4_u1_int_stat_reg[1]/P0001 ,
		_w10660_
	);
	LUT3 #(
		.INIT('ha8)
	) name8911 (
		\u4_u1_ienb_reg[3]/P0001 ,
		\u4_u1_int_stat_reg[3]/P0001 ,
		\u4_u1_int_stat_reg[4]/P0001 ,
		_w10661_
	);
	LUT4 #(
		.INIT('h135f)
	) name8912 (
		\u4_u1_ienb_reg[2]/P0001 ,
		\u4_u1_ienb_reg[4]/P0001 ,
		\u4_u1_int_stat_reg[2]/P0001 ,
		\u4_u1_int_stat_reg[5]/P0001 ,
		_w10662_
	);
	LUT4 #(
		.INIT('hfbff)
	) name8913 (
		_w10659_,
		_w10660_,
		_w10661_,
		_w10662_,
		_w10663_
	);
	LUT2 #(
		.INIT('h8)
	) name8914 (
		\u4_u2_ienb_reg[1]/P0001 ,
		\u4_u2_int_stat_reg[1]/P0001 ,
		_w10664_
	);
	LUT4 #(
		.INIT('h135f)
	) name8915 (
		\u4_u2_ienb_reg[0]/P0001 ,
		\u4_u2_ienb_reg[2]/P0001 ,
		\u4_u2_int_stat_reg[0]/P0001 ,
		\u4_u2_int_stat_reg[2]/P0001 ,
		_w10665_
	);
	LUT4 #(
		.INIT('h135f)
	) name8916 (
		\u4_u2_ienb_reg[4]/P0001 ,
		\u4_u2_ienb_reg[5]/P0001 ,
		\u4_u2_int_stat_reg[5]/P0001 ,
		\u4_u2_int_stat_reg[6]/P0001 ,
		_w10666_
	);
	LUT3 #(
		.INIT('ha8)
	) name8917 (
		\u4_u2_ienb_reg[3]/P0001 ,
		\u4_u2_int_stat_reg[3]/P0001 ,
		\u4_u2_int_stat_reg[4]/P0001 ,
		_w10667_
	);
	LUT4 #(
		.INIT('hffbf)
	) name8918 (
		_w10664_,
		_w10665_,
		_w10666_,
		_w10667_,
		_w10668_
	);
	LUT2 #(
		.INIT('h8)
	) name8919 (
		\u4_u2_iena_reg[5]/P0001 ,
		\u4_u2_int_stat_reg[6]/P0001 ,
		_w10669_
	);
	LUT4 #(
		.INIT('h135f)
	) name8920 (
		\u4_u2_iena_reg[1]/P0001 ,
		\u4_u2_iena_reg[2]/P0001 ,
		\u4_u2_int_stat_reg[1]/P0001 ,
		\u4_u2_int_stat_reg[2]/P0001 ,
		_w10670_
	);
	LUT3 #(
		.INIT('ha8)
	) name8921 (
		\u4_u2_iena_reg[3]/P0001 ,
		\u4_u2_int_stat_reg[3]/P0001 ,
		\u4_u2_int_stat_reg[4]/P0001 ,
		_w10671_
	);
	LUT4 #(
		.INIT('h135f)
	) name8922 (
		\u4_u2_iena_reg[0]/P0001 ,
		\u4_u2_iena_reg[4]/P0001 ,
		\u4_u2_int_stat_reg[0]/P0001 ,
		\u4_u2_int_stat_reg[5]/P0001 ,
		_w10672_
	);
	LUT4 #(
		.INIT('hfbff)
	) name8923 (
		_w10669_,
		_w10670_,
		_w10671_,
		_w10672_,
		_w10673_
	);
	LUT4 #(
		.INIT('h0001)
	) name8924 (
		\u4_u2_buf0_orig_reg[23]/P0001 ,
		\u4_u2_buf0_orig_reg[24]/P0001 ,
		\u4_u2_buf0_orig_reg[27]/P0001 ,
		\u4_u2_buf0_orig_reg[28]/P0001 ,
		_w10674_
	);
	LUT2 #(
		.INIT('h1)
	) name8925 (
		\u4_u2_buf0_orig_reg[29]/NET0131 ,
		\u4_u2_buf0_orig_reg[30]/NET0131 ,
		_w10675_
	);
	LUT4 #(
		.INIT('h0001)
	) name8926 (
		\u4_u2_buf0_orig_reg[21]/P0001 ,
		\u4_u2_buf0_orig_reg[22]/P0001 ,
		\u4_u2_buf0_orig_reg[25]/P0001 ,
		\u4_u2_buf0_orig_reg[26]/P0001 ,
		_w10676_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name8927 (
		_w5264_,
		_w10674_,
		_w10675_,
		_w10676_,
		_w10677_
	);
	LUT4 #(
		.INIT('h0001)
	) name8928 (
		\u4_u1_buf0_orig_reg[23]/P0001 ,
		\u4_u1_buf0_orig_reg[24]/P0001 ,
		\u4_u1_buf0_orig_reg[27]/P0001 ,
		\u4_u1_buf0_orig_reg[28]/P0001 ,
		_w10678_
	);
	LUT2 #(
		.INIT('h1)
	) name8929 (
		\u4_u1_buf0_orig_reg[29]/NET0131 ,
		\u4_u1_buf0_orig_reg[30]/NET0131 ,
		_w10679_
	);
	LUT4 #(
		.INIT('h0001)
	) name8930 (
		\u4_u1_buf0_orig_reg[21]/P0001 ,
		\u4_u1_buf0_orig_reg[22]/P0001 ,
		\u4_u1_buf0_orig_reg[25]/P0001 ,
		\u4_u1_buf0_orig_reg[26]/P0001 ,
		_w10680_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name8931 (
		_w5821_,
		_w10678_,
		_w10679_,
		_w10680_,
		_w10681_
	);
	LUT4 #(
		.INIT('h0001)
	) name8932 (
		\u4_u3_buf0_orig_reg[23]/P0001 ,
		\u4_u3_buf0_orig_reg[24]/P0001 ,
		\u4_u3_buf0_orig_reg[27]/P0001 ,
		\u4_u3_buf0_orig_reg[28]/P0001 ,
		_w10682_
	);
	LUT2 #(
		.INIT('h1)
	) name8933 (
		\u4_u3_buf0_orig_reg[29]/NET0131 ,
		\u4_u3_buf0_orig_reg[30]/NET0131 ,
		_w10683_
	);
	LUT4 #(
		.INIT('h0001)
	) name8934 (
		\u4_u3_buf0_orig_reg[21]/P0001 ,
		\u4_u3_buf0_orig_reg[22]/P0001 ,
		\u4_u3_buf0_orig_reg[25]/P0001 ,
		\u4_u3_buf0_orig_reg[26]/P0001 ,
		_w10684_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name8935 (
		_w5297_,
		_w10682_,
		_w10683_,
		_w10684_,
		_w10685_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name8936 (
		_w5792_,
		_w7833_,
		_w7834_,
		_w7840_,
		_w10686_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name8937 (
		_w3395_,
		_w5048_,
		_w5272_,
		_w5273_,
		_w10687_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name8938 (
		_w3407_,
		_w4984_,
		_w5799_,
		_w5800_,
		_w10688_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name8939 (
		_w3401_,
		_w4954_,
		_w5303_,
		_w5304_,
		_w10689_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name8940 (
		_w3413_,
		_w5018_,
		_w5829_,
		_w5830_,
		_w10690_
	);
	LUT3 #(
		.INIT('h6c)
	) name8941 (
		\u0_u0_idle_cnt1_reg[4]/P0001 ,
		\u0_u0_idle_cnt1_reg[5]/P0001 ,
		_w9015_,
		_w10691_
	);
	LUT3 #(
		.INIT('h78)
	) name8942 (
		\u0_u0_idle_cnt1_reg[0]/P0001 ,
		\u0_u0_idle_cnt1_reg[1]/P0001 ,
		\u0_u0_idle_cnt1_reg[2]/P0001 ,
		_w10692_
	);
	LUT4 #(
		.INIT('h639c)
	) name8943 (
		\u4_u2_buf0_orig_reg[19]/P0001 ,
		\u4_u2_buf0_orig_reg[20]/P0001 ,
		\u4_u2_dma_in_cnt_reg[0]/P0001 ,
		\u4_u2_dma_out_cnt_reg[1]/P0001 ,
		_w10693_
	);
	LUT4 #(
		.INIT('h639c)
	) name8944 (
		\u4_u3_buf0_orig_reg[19]/P0001 ,
		\u4_u3_buf0_orig_reg[20]/P0001 ,
		\u4_u3_dma_in_cnt_reg[0]/P0001 ,
		\u4_u3_dma_out_cnt_reg[1]/P0001 ,
		_w10694_
	);
	LUT4 #(
		.INIT('h639c)
	) name8945 (
		\u4_u0_buf0_orig_reg[19]/P0001 ,
		\u4_u0_buf0_orig_reg[20]/P0001 ,
		\u4_u0_dma_in_cnt_reg[0]/P0001 ,
		\u4_u0_dma_out_cnt_reg[1]/P0001 ,
		_w10695_
	);
	LUT4 #(
		.INIT('h639c)
	) name8946 (
		\u4_u1_buf0_orig_reg[19]/P0001 ,
		\u4_u1_buf0_orig_reg[20]/P0001 ,
		\u4_u1_dma_in_cnt_reg[0]/P0001 ,
		\u4_u1_dma_out_cnt_reg[1]/P0001 ,
		_w10696_
	);
	LUT4 #(
		.INIT('h8c88)
	) name8947 (
		\dma_ack_i[3]_pad ,
		rst_i_pad,
		\u4_u3_dma_ack_clr1_reg/P0001 ,
		\u4_u3_dma_ack_wr1_reg/P0001 ,
		_w10697_
	);
	LUT4 #(
		.INIT('h8c88)
	) name8948 (
		\dma_ack_i[0]_pad ,
		rst_i_pad,
		\u4_u0_dma_ack_clr1_reg/P0001 ,
		\u4_u0_dma_ack_wr1_reg/P0001 ,
		_w10698_
	);
	LUT4 #(
		.INIT('h8c88)
	) name8949 (
		\dma_ack_i[1]_pad ,
		rst_i_pad,
		\u4_u1_dma_ack_clr1_reg/P0001 ,
		\u4_u1_dma_ack_wr1_reg/P0001 ,
		_w10699_
	);
	LUT4 #(
		.INIT('h8c88)
	) name8950 (
		\dma_ack_i[2]_pad ,
		rst_i_pad,
		\u4_u2_dma_ack_clr1_reg/P0001 ,
		\u4_u2_dma_ack_wr1_reg/P0001 ,
		_w10700_
	);
	LUT3 #(
		.INIT('h14)
	) name8951 (
		\u0_rx_active_reg/P0001 ,
		\u1_u3_tx_data_to_cnt_reg[0]/P0001 ,
		\u1_u3_tx_data_to_cnt_reg[1]/P0001 ,
		_w10701_
	);
	LUT3 #(
		.INIT('h14)
	) name8952 (
		\u1_u3_rx_ack_to_clr_reg/P0001 ,
		\u1_u3_rx_ack_to_cnt_reg[0]/P0001 ,
		\u1_u3_rx_ack_to_cnt_reg[1]/P0001 ,
		_w10702_
	);
	LUT2 #(
		.INIT('h1)
	) name8953 (
		\u1_u3_rx_ack_to_clr_reg/P0001 ,
		\u1_u3_rx_ack_to_cnt_reg[0]/P0001 ,
		_w10703_
	);
	LUT3 #(
		.INIT('h80)
	) name8954 (
		\u1_hms_cnt_reg[2]/P0001 ,
		\u1_hms_cnt_reg[3]/P0001 ,
		\u1_hms_cnt_reg[4]/P0001 ,
		_w10704_
	);
	LUT2 #(
		.INIT('h8)
	) name8955 (
		_w4516_,
		_w10704_,
		_w10705_
	);
	LUT4 #(
		.INIT('h2000)
	) name8956 (
		\u0_u0_ps_cnt_reg[0]/P0001 ,
		\u0_u0_ps_cnt_reg[1]/P0001 ,
		\u0_u0_ps_cnt_reg[2]/P0001 ,
		\u0_u0_ps_cnt_reg[3]/P0001 ,
		_w10706_
	);
	LUT4 #(
		.INIT('h1248)
	) name8957 (
		\u1_u0_pid_reg[2]/NET0131 ,
		\u1_u0_pid_reg[3]/NET0131 ,
		\u1_u0_pid_reg[6]/P0001 ,
		\u1_u0_pid_reg[7]/P0001 ,
		_w10707_
	);
	LUT4 #(
		.INIT('h1248)
	) name8958 (
		\u1_u0_pid_reg[0]/NET0131 ,
		\u1_u0_pid_reg[1]/NET0131 ,
		\u1_u0_pid_reg[4]/P0001 ,
		\u1_u0_pid_reg[5]/P0001 ,
		_w10708_
	);
	LUT2 #(
		.INIT('h7)
	) name8959 (
		_w10707_,
		_w10708_,
		_w10709_
	);
	LUT4 #(
		.INIT('h4f44)
	) name8960 (
		\LineState_pad_i[0]_pad ,
		\LineState_pad_i[1]_pad ,
		\u0_u0_resume_req_s_reg/P0001 ,
		\u0_u0_usb_suspend_reg/P0001 ,
		_w10710_
	);
	LUT4 #(
		.INIT('h88a8)
	) name8961 (
		rst_i_pad,
		\u4_u2_r1_reg/P0001 ,
		\u4_u2_r2_reg/P0001 ,
		\u4_u2_r4_reg/P0001 ,
		_w10711_
	);
	LUT4 #(
		.INIT('h88a8)
	) name8962 (
		rst_i_pad,
		\u4_u3_r1_reg/P0001 ,
		\u4_u3_r2_reg/P0001 ,
		\u4_u3_r4_reg/P0001 ,
		_w10712_
	);
	LUT4 #(
		.INIT('h88a8)
	) name8963 (
		rst_i_pad,
		\u4_u0_r1_reg/P0001 ,
		\u4_u0_r2_reg/P0001 ,
		\u4_u0_r4_reg/P0001 ,
		_w10713_
	);
	LUT4 #(
		.INIT('h88a8)
	) name8964 (
		rst_i_pad,
		\u4_u1_r1_reg/P0001 ,
		\u4_u1_r2_reg/P0001 ,
		\u4_u1_r4_reg/P0001 ,
		_w10714_
	);
	LUT2 #(
		.INIT('h8)
	) name8965 (
		_w2122_,
		_w7864_,
		_w10715_
	);
	LUT2 #(
		.INIT('h1)
	) name8966 (
		\u0_rx_active_reg/P0001 ,
		\u1_u3_tx_data_to_cnt_reg[0]/P0001 ,
		_w10716_
	);
	LUT2 #(
		.INIT('h6)
	) name8967 (
		\u4_u1_buf0_orig_reg[19]/P0001 ,
		\u4_u1_buf0_orig_reg[20]/P0001 ,
		_w10717_
	);
	LUT2 #(
		.INIT('h6)
	) name8968 (
		\u0_u0_idle_cnt1_reg[0]/P0001 ,
		\u0_u0_idle_cnt1_reg[1]/P0001 ,
		_w10718_
	);
	LUT3 #(
		.INIT('hfe)
	) name8969 (
		\u1_u2_state_reg[2]/NET0131 ,
		\u1_u2_state_reg[3]/NET0131 ,
		\u1_u2_state_reg[4]/NET0131 ,
		_w10719_
	);
	LUT3 #(
		.INIT('he0)
	) name8970 (
		\u1_u3_buf0_rl_reg/P0001 ,
		\u1_u3_buf0_set_reg/P0001 ,
		\u4_u3_r5_reg/NET0131 ,
		_w10720_
	);
	LUT3 #(
		.INIT('he0)
	) name8971 (
		\u1_u3_buf0_rl_reg/P0001 ,
		\u1_u3_buf0_set_reg/P0001 ,
		\u4_u0_r5_reg/NET0131 ,
		_w10721_
	);
	LUT3 #(
		.INIT('he0)
	) name8972 (
		\u1_u3_buf0_rl_reg/P0001 ,
		\u1_u3_buf0_set_reg/P0001 ,
		\u4_u2_r5_reg/NET0131 ,
		_w10722_
	);
	LUT3 #(
		.INIT('h04)
	) name8973 (
		\u1_u2_mack_r_reg/P0001 ,
		\u1_u2_state_reg[1]/NET0131 ,
		\u1_u3_abort_reg/P0001 ,
		_w10723_
	);
	LUT3 #(
		.INIT('hab)
	) name8974 (
		TxValid_pad_o_pad,
		\u1_u3_state_reg[2]/P0001 ,
		\u1_u3_state_reg[3]/P0001 ,
		_w10724_
	);
	LUT3 #(
		.INIT('h40)
	) name8975 (
		\u0_u0_chirp_cnt_reg[0]/P0001 ,
		\u0_u0_chirp_cnt_reg[1]/P0001 ,
		\u0_u0_chirp_cnt_reg[2]/P0001 ,
		_w10725_
	);
	LUT3 #(
		.INIT('he0)
	) name8976 (
		\u1_u3_buf0_rl_reg/P0001 ,
		\u1_u3_buf0_set_reg/P0001 ,
		\u4_u1_r5_reg/NET0131 ,
		_w10726_
	);
	LUT2 #(
		.INIT('h6)
	) name8977 (
		\u4_u0_buf0_orig_reg[19]/P0001 ,
		\u4_u0_dma_in_cnt_reg[0]/P0001 ,
		_w10727_
	);
	LUT2 #(
		.INIT('h6)
	) name8978 (
		\u4_u3_buf0_orig_reg[19]/P0001 ,
		\u4_u3_dma_in_cnt_reg[0]/P0001 ,
		_w10728_
	);
	LUT2 #(
		.INIT('h6)
	) name8979 (
		\u4_u2_buf0_orig_reg[19]/P0001 ,
		\u4_u2_dma_in_cnt_reg[0]/P0001 ,
		_w10729_
	);
	LUT2 #(
		.INIT('h6)
	) name8980 (
		\u4_u1_buf0_orig_reg[19]/P0001 ,
		\u4_u1_dma_in_cnt_reg[0]/P0001 ,
		_w10730_
	);
	LUT2 #(
		.INIT('h6)
	) name8981 (
		\u4_u3_buf0_orig_reg[19]/P0001 ,
		\u4_u3_buf0_orig_reg[20]/P0001 ,
		_w10731_
	);
	LUT2 #(
		.INIT('h6)
	) name8982 (
		\u4_u0_buf0_orig_reg[19]/P0001 ,
		\u4_u0_buf0_orig_reg[20]/P0001 ,
		_w10732_
	);
	LUT2 #(
		.INIT('h6)
	) name8983 (
		\u4_u2_buf0_orig_reg[19]/P0001 ,
		\u4_u2_buf0_orig_reg[20]/P0001 ,
		_w10733_
	);
	LUT2 #(
		.INIT('h2)
	) name8984 (
		\u1_u3_new_size_reg[11]/P0001 ,
		\u1_u3_out_to_small_r_reg/P0001 ,
		_w10734_
	);
	LUT2 #(
		.INIT('h2)
	) name8985 (
		\u1_u3_buffer_done_reg/P0001 ,
		\u1_u3_out_to_small_r_reg/P0001 ,
		_w10735_
	);
	LUT2 #(
		.INIT('h4)
	) name8986 (
		\u1_u2_adr_cw_reg[0]/NET0131 ,
		\u1_u2_mack_r_reg/P0001 ,
		_w10736_
	);
	LUT2 #(
		.INIT('h8)
	) name8987 (
		wb_cyc_i_pad,
		wb_stb_i_pad,
		_w10737_
	);
	LUT2 #(
		.INIT('h8)
	) name8988 (
		RxError_pad_i_pad,
		rst_i_pad,
		_w10738_
	);
	LUT2 #(
		.INIT('h8)
	) name8989 (
		RxActive_pad_i_pad,
		rst_i_pad,
		_w10739_
	);
	LUT2 #(
		.INIT('h8)
	) name8990 (
		RxValid_pad_i_pad,
		rst_i_pad,
		_w10740_
	);
	LUT2 #(
		.INIT('h8)
	) name8991 (
		\u1_u2_adr_cw_reg[0]/NET0131 ,
		\u1_u2_mack_r_reg/P0001 ,
		_w10741_
	);
	LUT4 #(
		.INIT('h9a99)
	) name8992 (
		\u1_u2_sizd_c_reg[1]/P0001 ,
		_w2748_,
		_w2757_,
		_w2758_,
		_w10742_
	);
	LUT4 #(
		.INIT('h0015)
	) name8993 (
		\u1_u2_tx_dma_en_r_reg/P0001 ,
		_w2766_,
		_w2773_,
		_w10742_,
		_w10743_
	);
	LUT2 #(
		.INIT('h2)
	) name8994 (
		rst_i_pad,
		_w10743_,
		_w10744_
	);
	LUT4 #(
		.INIT('h45ff)
	) name8995 (
		_w2779_,
		_w3916_,
		_w3922_,
		_w10744_,
		_w10745_
	);
	LUT4 #(
		.INIT('h20aa)
	) name8996 (
		\u4_csr_reg[2]/NET0131 ,
		_w2826_,
		_w2866_,
		_w2898_,
		_w10746_
	);
	LUT2 #(
		.INIT('he)
	) name8997 (
		_w2935_,
		_w10746_,
		_w10747_
	);
	LUT3 #(
		.INIT('h15)
	) name8998 (
		\u2_wack_r_reg/P0001 ,
		_w5493_,
		_w5494_,
		_w10748_
	);
	LUT3 #(
		.INIT('h45)
	) name8999 (
		\u1_u2_word_done_r_reg/P0001 ,
		_w5492_,
		_w10748_,
		_w10749_
	);
	LUT2 #(
		.INIT('h4)
	) name9000 (
		\u1_u2_word_done_r_reg/P0001 ,
		\wb_addr_i[2]_pad ,
		_w10750_
	);
	LUT3 #(
		.INIT('hb0)
	) name9001 (
		_w5492_,
		_w10748_,
		_w10750_,
		_w10751_
	);
	LUT4 #(
		.INIT('hbb8a)
	) name9002 (
		\u1_u2_adr_cw_reg[0]/NET0131 ,
		_w5489_,
		_w10749_,
		_w10751_,
		_w10752_
	);
	LUT2 #(
		.INIT('h4)
	) name9003 (
		\u1_u2_word_done_r_reg/P0001 ,
		\wb_addr_i[12]_pad ,
		_w10753_
	);
	LUT3 #(
		.INIT('hb0)
	) name9004 (
		_w5492_,
		_w10748_,
		_w10753_,
		_w10754_
	);
	LUT4 #(
		.INIT('hbb8a)
	) name9005 (
		\u1_u2_adr_cw_reg[10]/P0001 ,
		_w5489_,
		_w10749_,
		_w10754_,
		_w10755_
	);
	LUT2 #(
		.INIT('h4)
	) name9006 (
		\u1_u2_word_done_r_reg/P0001 ,
		\wb_addr_i[13]_pad ,
		_w10756_
	);
	LUT3 #(
		.INIT('hb0)
	) name9007 (
		_w5492_,
		_w10748_,
		_w10756_,
		_w10757_
	);
	LUT4 #(
		.INIT('hbb8a)
	) name9008 (
		\u1_u2_adr_cw_reg[11]/P0001 ,
		_w5489_,
		_w10749_,
		_w10757_,
		_w10758_
	);
	LUT2 #(
		.INIT('h4)
	) name9009 (
		\u1_u2_word_done_r_reg/P0001 ,
		\wb_addr_i[14]_pad ,
		_w10759_
	);
	LUT3 #(
		.INIT('hb0)
	) name9010 (
		_w5492_,
		_w10748_,
		_w10759_,
		_w10760_
	);
	LUT4 #(
		.INIT('hbb8a)
	) name9011 (
		\u1_u2_adr_cw_reg[12]/P0001 ,
		_w5489_,
		_w10749_,
		_w10760_,
		_w10761_
	);
	LUT2 #(
		.INIT('h4)
	) name9012 (
		\u1_u2_word_done_r_reg/P0001 ,
		\wb_addr_i[15]_pad ,
		_w10762_
	);
	LUT3 #(
		.INIT('hb0)
	) name9013 (
		_w5492_,
		_w10748_,
		_w10762_,
		_w10763_
	);
	LUT4 #(
		.INIT('hbb8a)
	) name9014 (
		\u1_u2_adr_cw_reg[13]/P0001 ,
		_w5489_,
		_w10749_,
		_w10763_,
		_w10764_
	);
	LUT2 #(
		.INIT('h4)
	) name9015 (
		\u1_u2_word_done_r_reg/P0001 ,
		\wb_addr_i[16]_pad ,
		_w10765_
	);
	LUT3 #(
		.INIT('hb0)
	) name9016 (
		_w5492_,
		_w10748_,
		_w10765_,
		_w10766_
	);
	LUT4 #(
		.INIT('hbb8a)
	) name9017 (
		\u1_u2_adr_cw_reg[14]/P0001 ,
		_w5489_,
		_w10749_,
		_w10766_,
		_w10767_
	);
	LUT2 #(
		.INIT('h4)
	) name9018 (
		\u1_u2_word_done_r_reg/P0001 ,
		\wb_addr_i[3]_pad ,
		_w10768_
	);
	LUT3 #(
		.INIT('hb0)
	) name9019 (
		_w5492_,
		_w10748_,
		_w10768_,
		_w10769_
	);
	LUT4 #(
		.INIT('hbb8a)
	) name9020 (
		\u1_u2_adr_cw_reg[1]/P0001 ,
		_w5489_,
		_w10749_,
		_w10769_,
		_w10770_
	);
	LUT2 #(
		.INIT('h4)
	) name9021 (
		\u1_u2_word_done_r_reg/P0001 ,
		\wb_addr_i[4]_pad ,
		_w10771_
	);
	LUT3 #(
		.INIT('hb0)
	) name9022 (
		_w5492_,
		_w10748_,
		_w10771_,
		_w10772_
	);
	LUT4 #(
		.INIT('hbb8a)
	) name9023 (
		\u1_u2_adr_cw_reg[2]/P0001 ,
		_w5489_,
		_w10749_,
		_w10772_,
		_w10773_
	);
	LUT2 #(
		.INIT('h4)
	) name9024 (
		\u1_u2_word_done_r_reg/P0001 ,
		\wb_addr_i[5]_pad ,
		_w10774_
	);
	LUT3 #(
		.INIT('hb0)
	) name9025 (
		_w5492_,
		_w10748_,
		_w10774_,
		_w10775_
	);
	LUT4 #(
		.INIT('hbb8a)
	) name9026 (
		\u1_u2_adr_cw_reg[3]/NET0131 ,
		_w5489_,
		_w10749_,
		_w10775_,
		_w10776_
	);
	LUT2 #(
		.INIT('h4)
	) name9027 (
		\u1_u2_word_done_r_reg/P0001 ,
		\wb_addr_i[6]_pad ,
		_w10777_
	);
	LUT3 #(
		.INIT('hb0)
	) name9028 (
		_w5492_,
		_w10748_,
		_w10777_,
		_w10778_
	);
	LUT4 #(
		.INIT('hbb8a)
	) name9029 (
		\u1_u2_adr_cw_reg[4]/P0001 ,
		_w5489_,
		_w10749_,
		_w10778_,
		_w10779_
	);
	LUT2 #(
		.INIT('h4)
	) name9030 (
		\u1_u2_word_done_r_reg/P0001 ,
		\wb_addr_i[7]_pad ,
		_w10780_
	);
	LUT3 #(
		.INIT('hb0)
	) name9031 (
		_w5492_,
		_w10748_,
		_w10780_,
		_w10781_
	);
	LUT4 #(
		.INIT('hbb8a)
	) name9032 (
		\u1_u2_adr_cw_reg[5]/NET0131 ,
		_w5489_,
		_w10749_,
		_w10781_,
		_w10782_
	);
	LUT2 #(
		.INIT('h4)
	) name9033 (
		\u1_u2_word_done_r_reg/P0001 ,
		\wb_addr_i[8]_pad ,
		_w10783_
	);
	LUT3 #(
		.INIT('hb0)
	) name9034 (
		_w5492_,
		_w10748_,
		_w10783_,
		_w10784_
	);
	LUT4 #(
		.INIT('hbb8a)
	) name9035 (
		\u1_u2_adr_cw_reg[6]/NET0131 ,
		_w5489_,
		_w10749_,
		_w10784_,
		_w10785_
	);
	LUT2 #(
		.INIT('h4)
	) name9036 (
		\u1_u2_word_done_r_reg/P0001 ,
		\wb_addr_i[9]_pad ,
		_w10786_
	);
	LUT3 #(
		.INIT('hb0)
	) name9037 (
		_w5492_,
		_w10748_,
		_w10786_,
		_w10787_
	);
	LUT4 #(
		.INIT('hbb8a)
	) name9038 (
		\u1_u2_adr_cw_reg[7]/NET0131 ,
		_w5489_,
		_w10749_,
		_w10787_,
		_w10788_
	);
	LUT2 #(
		.INIT('h4)
	) name9039 (
		\u1_u2_word_done_r_reg/P0001 ,
		\wb_addr_i[10]_pad ,
		_w10789_
	);
	LUT3 #(
		.INIT('hb0)
	) name9040 (
		_w5492_,
		_w10748_,
		_w10789_,
		_w10790_
	);
	LUT4 #(
		.INIT('hbb8a)
	) name9041 (
		\u1_u2_adr_cw_reg[8]/P0001 ,
		_w5489_,
		_w10749_,
		_w10790_,
		_w10791_
	);
	LUT2 #(
		.INIT('h4)
	) name9042 (
		\u1_u2_word_done_r_reg/P0001 ,
		\wb_addr_i[11]_pad ,
		_w10792_
	);
	LUT3 #(
		.INIT('hb0)
	) name9043 (
		_w5492_,
		_w10748_,
		_w10792_,
		_w10793_
	);
	LUT4 #(
		.INIT('hbb8a)
	) name9044 (
		\u1_u2_adr_cw_reg[9]/NET0131 ,
		_w5489_,
		_w10749_,
		_w10793_,
		_w10794_
	);
	LUT2 #(
		.INIT('h4)
	) name9045 (
		\u1_u2_word_done_r_reg/P0001 ,
		\wb_data_i[0]_pad ,
		_w10795_
	);
	LUT3 #(
		.INIT('hb0)
	) name9046 (
		_w5492_,
		_w10748_,
		_w10795_,
		_w10796_
	);
	LUT4 #(
		.INIT('hbb8a)
	) name9047 (
		\u1_u2_dout_r_reg[0]/P0001 ,
		_w5489_,
		_w10749_,
		_w10796_,
		_w10797_
	);
	LUT2 #(
		.INIT('h4)
	) name9048 (
		\u1_u2_word_done_r_reg/P0001 ,
		\wb_data_i[10]_pad ,
		_w10798_
	);
	LUT3 #(
		.INIT('hb0)
	) name9049 (
		_w5492_,
		_w10748_,
		_w10798_,
		_w10799_
	);
	LUT4 #(
		.INIT('hbb8a)
	) name9050 (
		\u1_u2_dout_r_reg[10]/P0001 ,
		_w5489_,
		_w10749_,
		_w10799_,
		_w10800_
	);
	LUT2 #(
		.INIT('h4)
	) name9051 (
		\u1_u2_word_done_r_reg/P0001 ,
		\wb_data_i[11]_pad ,
		_w10801_
	);
	LUT3 #(
		.INIT('hb0)
	) name9052 (
		_w5492_,
		_w10748_,
		_w10801_,
		_w10802_
	);
	LUT4 #(
		.INIT('hbb8a)
	) name9053 (
		\u1_u2_dout_r_reg[11]/P0001 ,
		_w5489_,
		_w10749_,
		_w10802_,
		_w10803_
	);
	LUT2 #(
		.INIT('h4)
	) name9054 (
		\u1_u2_word_done_r_reg/P0001 ,
		\wb_data_i[12]_pad ,
		_w10804_
	);
	LUT3 #(
		.INIT('hb0)
	) name9055 (
		_w5492_,
		_w10748_,
		_w10804_,
		_w10805_
	);
	LUT4 #(
		.INIT('hbb8a)
	) name9056 (
		\u1_u2_dout_r_reg[12]/P0001 ,
		_w5489_,
		_w10749_,
		_w10805_,
		_w10806_
	);
	LUT2 #(
		.INIT('h4)
	) name9057 (
		\u1_u2_word_done_r_reg/P0001 ,
		\wb_data_i[13]_pad ,
		_w10807_
	);
	LUT3 #(
		.INIT('hb0)
	) name9058 (
		_w5492_,
		_w10748_,
		_w10807_,
		_w10808_
	);
	LUT4 #(
		.INIT('hbb8a)
	) name9059 (
		\u1_u2_dout_r_reg[13]/P0001 ,
		_w5489_,
		_w10749_,
		_w10808_,
		_w10809_
	);
	LUT2 #(
		.INIT('h4)
	) name9060 (
		\u1_u2_word_done_r_reg/P0001 ,
		\wb_data_i[14]_pad ,
		_w10810_
	);
	LUT3 #(
		.INIT('hb0)
	) name9061 (
		_w5492_,
		_w10748_,
		_w10810_,
		_w10811_
	);
	LUT4 #(
		.INIT('hbb8a)
	) name9062 (
		\u1_u2_dout_r_reg[14]/P0001 ,
		_w5489_,
		_w10749_,
		_w10811_,
		_w10812_
	);
	LUT2 #(
		.INIT('h4)
	) name9063 (
		\u1_u2_word_done_r_reg/P0001 ,
		\wb_data_i[15]_pad ,
		_w10813_
	);
	LUT3 #(
		.INIT('hb0)
	) name9064 (
		_w5492_,
		_w10748_,
		_w10813_,
		_w10814_
	);
	LUT4 #(
		.INIT('hbb8a)
	) name9065 (
		\u1_u2_dout_r_reg[15]/P0001 ,
		_w5489_,
		_w10749_,
		_w10814_,
		_w10815_
	);
	LUT2 #(
		.INIT('h4)
	) name9066 (
		\u1_u2_word_done_r_reg/P0001 ,
		\wb_data_i[16]_pad ,
		_w10816_
	);
	LUT3 #(
		.INIT('hb0)
	) name9067 (
		_w5492_,
		_w10748_,
		_w10816_,
		_w10817_
	);
	LUT4 #(
		.INIT('hbb8a)
	) name9068 (
		\u1_u2_dout_r_reg[16]/P0001 ,
		_w5489_,
		_w10749_,
		_w10817_,
		_w10818_
	);
	LUT2 #(
		.INIT('h4)
	) name9069 (
		\u1_u2_word_done_r_reg/P0001 ,
		\wb_data_i[17]_pad ,
		_w10819_
	);
	LUT3 #(
		.INIT('hb0)
	) name9070 (
		_w5492_,
		_w10748_,
		_w10819_,
		_w10820_
	);
	LUT4 #(
		.INIT('hbb8a)
	) name9071 (
		\u1_u2_dout_r_reg[17]/P0001 ,
		_w5489_,
		_w10749_,
		_w10820_,
		_w10821_
	);
	LUT2 #(
		.INIT('h4)
	) name9072 (
		\u1_u2_word_done_r_reg/P0001 ,
		\wb_data_i[18]_pad ,
		_w10822_
	);
	LUT3 #(
		.INIT('hb0)
	) name9073 (
		_w5492_,
		_w10748_,
		_w10822_,
		_w10823_
	);
	LUT4 #(
		.INIT('hbb8a)
	) name9074 (
		\u1_u2_dout_r_reg[18]/P0001 ,
		_w5489_,
		_w10749_,
		_w10823_,
		_w10824_
	);
	LUT2 #(
		.INIT('h4)
	) name9075 (
		\u1_u2_word_done_r_reg/P0001 ,
		\wb_data_i[19]_pad ,
		_w10825_
	);
	LUT3 #(
		.INIT('hb0)
	) name9076 (
		_w5492_,
		_w10748_,
		_w10825_,
		_w10826_
	);
	LUT4 #(
		.INIT('hbb8a)
	) name9077 (
		\u1_u2_dout_r_reg[19]/P0001 ,
		_w5489_,
		_w10749_,
		_w10826_,
		_w10827_
	);
	LUT2 #(
		.INIT('h4)
	) name9078 (
		\u1_u2_word_done_r_reg/P0001 ,
		\wb_data_i[1]_pad ,
		_w10828_
	);
	LUT3 #(
		.INIT('hb0)
	) name9079 (
		_w5492_,
		_w10748_,
		_w10828_,
		_w10829_
	);
	LUT4 #(
		.INIT('hbb8a)
	) name9080 (
		\u1_u2_dout_r_reg[1]/P0001 ,
		_w5489_,
		_w10749_,
		_w10829_,
		_w10830_
	);
	LUT2 #(
		.INIT('h4)
	) name9081 (
		\u1_u2_word_done_r_reg/P0001 ,
		\wb_data_i[20]_pad ,
		_w10831_
	);
	LUT3 #(
		.INIT('hb0)
	) name9082 (
		_w5492_,
		_w10748_,
		_w10831_,
		_w10832_
	);
	LUT4 #(
		.INIT('hbb8a)
	) name9083 (
		\u1_u2_dout_r_reg[20]/P0001 ,
		_w5489_,
		_w10749_,
		_w10832_,
		_w10833_
	);
	LUT2 #(
		.INIT('h4)
	) name9084 (
		\u1_u2_word_done_r_reg/P0001 ,
		\wb_data_i[21]_pad ,
		_w10834_
	);
	LUT3 #(
		.INIT('hb0)
	) name9085 (
		_w5492_,
		_w10748_,
		_w10834_,
		_w10835_
	);
	LUT4 #(
		.INIT('hbb8a)
	) name9086 (
		\u1_u2_dout_r_reg[21]/P0001 ,
		_w5489_,
		_w10749_,
		_w10835_,
		_w10836_
	);
	LUT2 #(
		.INIT('h4)
	) name9087 (
		\u1_u2_word_done_r_reg/P0001 ,
		\wb_data_i[22]_pad ,
		_w10837_
	);
	LUT3 #(
		.INIT('hb0)
	) name9088 (
		_w5492_,
		_w10748_,
		_w10837_,
		_w10838_
	);
	LUT4 #(
		.INIT('hbb8a)
	) name9089 (
		\u1_u2_dout_r_reg[22]/P0001 ,
		_w5489_,
		_w10749_,
		_w10838_,
		_w10839_
	);
	LUT2 #(
		.INIT('h4)
	) name9090 (
		\u1_u2_word_done_r_reg/P0001 ,
		\wb_data_i[23]_pad ,
		_w10840_
	);
	LUT3 #(
		.INIT('hb0)
	) name9091 (
		_w5492_,
		_w10748_,
		_w10840_,
		_w10841_
	);
	LUT4 #(
		.INIT('hbb8a)
	) name9092 (
		\u1_u2_dout_r_reg[23]/P0001 ,
		_w5489_,
		_w10749_,
		_w10841_,
		_w10842_
	);
	LUT2 #(
		.INIT('h4)
	) name9093 (
		\u1_u2_word_done_r_reg/P0001 ,
		\wb_data_i[24]_pad ,
		_w10843_
	);
	LUT3 #(
		.INIT('hb0)
	) name9094 (
		_w5492_,
		_w10748_,
		_w10843_,
		_w10844_
	);
	LUT4 #(
		.INIT('hbb8a)
	) name9095 (
		\u1_u2_dout_r_reg[24]/P0001 ,
		_w5489_,
		_w10749_,
		_w10844_,
		_w10845_
	);
	LUT2 #(
		.INIT('h4)
	) name9096 (
		\u1_u2_word_done_r_reg/P0001 ,
		\wb_data_i[25]_pad ,
		_w10846_
	);
	LUT3 #(
		.INIT('hb0)
	) name9097 (
		_w5492_,
		_w10748_,
		_w10846_,
		_w10847_
	);
	LUT4 #(
		.INIT('hbb8a)
	) name9098 (
		\u1_u2_dout_r_reg[25]/P0001 ,
		_w5489_,
		_w10749_,
		_w10847_,
		_w10848_
	);
	LUT2 #(
		.INIT('h4)
	) name9099 (
		\u1_u2_word_done_r_reg/P0001 ,
		\wb_data_i[26]_pad ,
		_w10849_
	);
	LUT3 #(
		.INIT('hb0)
	) name9100 (
		_w5492_,
		_w10748_,
		_w10849_,
		_w10850_
	);
	LUT4 #(
		.INIT('hbb8a)
	) name9101 (
		\u1_u2_dout_r_reg[26]/P0001 ,
		_w5489_,
		_w10749_,
		_w10850_,
		_w10851_
	);
	LUT2 #(
		.INIT('h4)
	) name9102 (
		\u1_u2_word_done_r_reg/P0001 ,
		\wb_data_i[27]_pad ,
		_w10852_
	);
	LUT3 #(
		.INIT('hb0)
	) name9103 (
		_w5492_,
		_w10748_,
		_w10852_,
		_w10853_
	);
	LUT4 #(
		.INIT('hbb8a)
	) name9104 (
		\u1_u2_dout_r_reg[27]/P0001 ,
		_w5489_,
		_w10749_,
		_w10853_,
		_w10854_
	);
	LUT2 #(
		.INIT('h4)
	) name9105 (
		\u1_u2_word_done_r_reg/P0001 ,
		\wb_data_i[28]_pad ,
		_w10855_
	);
	LUT3 #(
		.INIT('hb0)
	) name9106 (
		_w5492_,
		_w10748_,
		_w10855_,
		_w10856_
	);
	LUT4 #(
		.INIT('hbb8a)
	) name9107 (
		\u1_u2_dout_r_reg[28]/P0001 ,
		_w5489_,
		_w10749_,
		_w10856_,
		_w10857_
	);
	LUT2 #(
		.INIT('h4)
	) name9108 (
		\u1_u2_word_done_r_reg/P0001 ,
		\wb_data_i[29]_pad ,
		_w10858_
	);
	LUT3 #(
		.INIT('hb0)
	) name9109 (
		_w5492_,
		_w10748_,
		_w10858_,
		_w10859_
	);
	LUT4 #(
		.INIT('hbb8a)
	) name9110 (
		\u1_u2_dout_r_reg[29]/P0001 ,
		_w5489_,
		_w10749_,
		_w10859_,
		_w10860_
	);
	LUT2 #(
		.INIT('h4)
	) name9111 (
		\u1_u2_word_done_r_reg/P0001 ,
		\wb_data_i[2]_pad ,
		_w10861_
	);
	LUT3 #(
		.INIT('hb0)
	) name9112 (
		_w5492_,
		_w10748_,
		_w10861_,
		_w10862_
	);
	LUT4 #(
		.INIT('hbb8a)
	) name9113 (
		\u1_u2_dout_r_reg[2]/P0001 ,
		_w5489_,
		_w10749_,
		_w10862_,
		_w10863_
	);
	LUT2 #(
		.INIT('h4)
	) name9114 (
		\u1_u2_word_done_r_reg/P0001 ,
		\wb_data_i[30]_pad ,
		_w10864_
	);
	LUT3 #(
		.INIT('hb0)
	) name9115 (
		_w5492_,
		_w10748_,
		_w10864_,
		_w10865_
	);
	LUT4 #(
		.INIT('hbb8a)
	) name9116 (
		\u1_u2_dout_r_reg[30]/P0001 ,
		_w5489_,
		_w10749_,
		_w10865_,
		_w10866_
	);
	LUT2 #(
		.INIT('h4)
	) name9117 (
		\u1_u2_word_done_r_reg/P0001 ,
		\wb_data_i[31]_pad ,
		_w10867_
	);
	LUT3 #(
		.INIT('hb0)
	) name9118 (
		_w5492_,
		_w10748_,
		_w10867_,
		_w10868_
	);
	LUT4 #(
		.INIT('hbb8a)
	) name9119 (
		\u1_u2_dout_r_reg[31]/P0001 ,
		_w5489_,
		_w10749_,
		_w10868_,
		_w10869_
	);
	LUT2 #(
		.INIT('h4)
	) name9120 (
		\u1_u2_word_done_r_reg/P0001 ,
		\wb_data_i[3]_pad ,
		_w10870_
	);
	LUT3 #(
		.INIT('hb0)
	) name9121 (
		_w5492_,
		_w10748_,
		_w10870_,
		_w10871_
	);
	LUT4 #(
		.INIT('hbb8a)
	) name9122 (
		\u1_u2_dout_r_reg[3]/P0001 ,
		_w5489_,
		_w10749_,
		_w10871_,
		_w10872_
	);
	LUT2 #(
		.INIT('h4)
	) name9123 (
		\u1_u2_word_done_r_reg/P0001 ,
		\wb_data_i[4]_pad ,
		_w10873_
	);
	LUT3 #(
		.INIT('hb0)
	) name9124 (
		_w5492_,
		_w10748_,
		_w10873_,
		_w10874_
	);
	LUT4 #(
		.INIT('hbb8a)
	) name9125 (
		\u1_u2_dout_r_reg[4]/P0001 ,
		_w5489_,
		_w10749_,
		_w10874_,
		_w10875_
	);
	LUT2 #(
		.INIT('h4)
	) name9126 (
		\u1_u2_word_done_r_reg/P0001 ,
		\wb_data_i[5]_pad ,
		_w10876_
	);
	LUT3 #(
		.INIT('hb0)
	) name9127 (
		_w5492_,
		_w10748_,
		_w10876_,
		_w10877_
	);
	LUT4 #(
		.INIT('hbb8a)
	) name9128 (
		\u1_u2_dout_r_reg[5]/P0001 ,
		_w5489_,
		_w10749_,
		_w10877_,
		_w10878_
	);
	LUT2 #(
		.INIT('h4)
	) name9129 (
		\u1_u2_word_done_r_reg/P0001 ,
		\wb_data_i[6]_pad ,
		_w10879_
	);
	LUT3 #(
		.INIT('hb0)
	) name9130 (
		_w5492_,
		_w10748_,
		_w10879_,
		_w10880_
	);
	LUT4 #(
		.INIT('hbb8a)
	) name9131 (
		\u1_u2_dout_r_reg[6]/P0001 ,
		_w5489_,
		_w10749_,
		_w10880_,
		_w10881_
	);
	LUT2 #(
		.INIT('h4)
	) name9132 (
		\u1_u2_word_done_r_reg/P0001 ,
		\wb_data_i[7]_pad ,
		_w10882_
	);
	LUT3 #(
		.INIT('hb0)
	) name9133 (
		_w5492_,
		_w10748_,
		_w10882_,
		_w10883_
	);
	LUT4 #(
		.INIT('hbb8a)
	) name9134 (
		\u1_u2_dout_r_reg[7]/P0001 ,
		_w5489_,
		_w10749_,
		_w10883_,
		_w10884_
	);
	LUT2 #(
		.INIT('h4)
	) name9135 (
		\u1_u2_word_done_r_reg/P0001 ,
		\wb_data_i[8]_pad ,
		_w10885_
	);
	LUT3 #(
		.INIT('hb0)
	) name9136 (
		_w5492_,
		_w10748_,
		_w10885_,
		_w10886_
	);
	LUT4 #(
		.INIT('hbb8a)
	) name9137 (
		\u1_u2_dout_r_reg[8]/P0001 ,
		_w5489_,
		_w10749_,
		_w10886_,
		_w10887_
	);
	LUT2 #(
		.INIT('h4)
	) name9138 (
		\u1_u2_word_done_r_reg/P0001 ,
		\wb_data_i[9]_pad ,
		_w10888_
	);
	LUT3 #(
		.INIT('hb0)
	) name9139 (
		_w5492_,
		_w10748_,
		_w10888_,
		_w10889_
	);
	LUT4 #(
		.INIT('hbb8a)
	) name9140 (
		\u1_u2_dout_r_reg[9]/P0001 ,
		_w5489_,
		_w10749_,
		_w10889_,
		_w10890_
	);
	LUT2 #(
		.INIT('h8)
	) name9141 (
		\u1_u2_mwe_reg/P0001 ,
		\u1_u2_word_done_r_reg/P0001 ,
		_w10891_
	);
	LUT2 #(
		.INIT('h4)
	) name9142 (
		\u1_u2_mack_r_reg/P0001 ,
		\u1_u2_mwe_reg/P0001 ,
		_w10892_
	);
	LUT4 #(
		.INIT('h020f)
	) name9143 (
		_w3224_,
		_w5488_,
		_w10891_,
		_w10892_,
		_w10893_
	);
	LUT3 #(
		.INIT('h80)
	) name9144 (
		_w2224_,
		_w2225_,
		_w6430_,
		_w10894_
	);
	LUT4 #(
		.INIT('h4404)
	) name9145 (
		_w5489_,
		_w5496_,
		_w6435_,
		_w10894_,
		_w10895_
	);
	LUT2 #(
		.INIT('hd)
	) name9146 (
		_w10893_,
		_w10895_,
		_w10896_
	);
	LUT3 #(
		.INIT('h20)
	) name9147 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w10897_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name9148 (
		\u4_utmi_vend_ctrl_r_reg[0]/P0001 ,
		\wb_data_i[0]_pad ,
		_w8842_,
		_w10897_,
		_w10898_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name9149 (
		\u4_utmi_vend_ctrl_r_reg[1]/P0001 ,
		\wb_data_i[1]_pad ,
		_w8842_,
		_w10897_,
		_w10899_
	);
	LUT4 #(
		.INIT('hcaaa)
	) name9150 (
		\u4_utmi_vend_ctrl_r_reg[2]/P0001 ,
		\wb_data_i[2]_pad ,
		_w8842_,
		_w10897_,
		_w10900_
	);
	LUT4 #(
		.INIT('h2000)
	) name9151 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		\wb_data_i[3]_pad ,
		_w10901_
	);
	LUT4 #(
		.INIT('hee2a)
	) name9152 (
		\u4_utmi_vend_ctrl_r_reg[3]/P0001 ,
		_w8842_,
		_w10897_,
		_w10901_,
		_w10902_
	);
	assign \dma_req_o[6]_pad  = 1'b0;
	assign \g37425/_0_  = _w1832_ ;
	assign \g37426/_0_  = _w1874_ ;
	assign \g37432/_0_  = _w1919_ ;
	assign \g37433/_0_  = _w1961_ ;
	assign \g37439/_0_  = _w2102_ ;
	assign \g37440/_0_  = _w2114_ ;
	assign \g37444/_00_  = _w2141_ ;
	assign \g37448/_0_  = _w2149_ ;
	assign \g37450/_0_  = _w2154_ ;
	assign \g37454/_0_  = _w2160_ ;
	assign \g37473/_0_  = _w2169_ ;
	assign \g37474/_0_  = _w2181_ ;
	assign \g37475/_0_  = _w2190_ ;
	assign \g37476/_0_  = _w2202_ ;
	assign \g37477/_0_  = _w2211_ ;
	assign \g37478/_0_  = _w2216_ ;
	assign \g37479/_0_  = _w2223_ ;
	assign \g37488/_0_  = _w2239_ ;
	assign \g37489/_0_  = _w2250_ ;
	assign \g37490/_0_  = _w2259_ ;
	assign \g37491/_0_  = _w2266_ ;
	assign \g37492/_0_  = _w2273_ ;
	assign \g37517/_0_  = _w2279_ ;
	assign \g37518/_0_  = _w2284_ ;
	assign \g37519/_0_  = _w2289_ ;
	assign \g37520/_0_  = _w2294_ ;
	assign \g37521/_0_  = _w2302_ ;
	assign \g37522/_0_  = _w2313_ ;
	assign \g37540/_0_  = _w2319_ ;
	assign \g37542/_0_  = _w2327_ ;
	assign \g37543/_0_  = _w2332_ ;
	assign \g37545/_0_  = _w2338_ ;
	assign \g37546/_0_  = _w2343_ ;
	assign \g37548/_0_  = _w2349_ ;
	assign \g37549/_0_  = _w2360_ ;
	assign \g37550/_0_  = _w2365_ ;
	assign \g37551/_0_  = _w2371_ ;
	assign \g37556/_0_  = _w2382_ ;
	assign \g37589/_0_  = _w2388_ ;
	assign \g37591/_0_  = _w2394_ ;
	assign \g37592/_0_  = _w2400_ ;
	assign \g37593/_0_  = _w2407_ ;
	assign \g37594/_0_  = _w2413_ ;
	assign \g37596/_0_  = _w2418_ ;
	assign \g37597/_0_  = _w2423_ ;
	assign \g37598/_0_  = _w2428_ ;
	assign \g37599/_0_  = _w2434_ ;
	assign \g37601/_0_  = _w2439_ ;
	assign \g37603/_0_  = _w2444_ ;
	assign \g37604/_0_  = _w2450_ ;
	assign \g37605/_0_  = _w2455_ ;
	assign \g37607/_0_  = _w2460_ ;
	assign \g37608/_0_  = _w2465_ ;
	assign \g37609/_0_  = _w2471_ ;
	assign \g37610/_0_  = _w2476_ ;
	assign \g37645/_0_  = _w2483_ ;
	assign \g37648/_0_  = _w2489_ ;
	assign \g37650/_0_  = _w2495_ ;
	assign \g37653/_0_  = _w2501_ ;
	assign \g37664/_3_  = _w2505_ ;
	assign \g37703/_0_  = _w2511_ ;
	assign \g37704/_0_  = _w2517_ ;
	assign \g37706/_0_  = _w2523_ ;
	assign \g37708/_0_  = _w2530_ ;
	assign \g37709/_0_  = _w2537_ ;
	assign \g37711/_0_  = _w2544_ ;
	assign \g37714/_0_  = _w2549_ ;
	assign \g37715/_0_  = _w2554_ ;
	assign \g37717/_0_  = _w2559_ ;
	assign \g37718/_0_  = _w2565_ ;
	assign \g37719/_0_  = _w2571_ ;
	assign \g37720/_0_  = _w2577_ ;
	assign \g37723/_0_  = _w2582_ ;
	assign \g37724/_0_  = _w2587_ ;
	assign \g37726/_0_  = _w2592_ ;
	assign \g37728/_0_  = _w2598_ ;
	assign \g37729/_0_  = _w2604_ ;
	assign \g37730/_0_  = _w2610_ ;
	assign \g37731/_0_  = _w2615_ ;
	assign \g37732/_0_  = _w2620_ ;
	assign \g37733/_0_  = _w2625_ ;
	assign \g37735/_0_  = _w2631_ ;
	assign \g37736/_0_  = _w2637_ ;
	assign \g37737/_0_  = _w2643_ ;
	assign \g37856/_0_  = _w2650_ ;
	assign \g37857/_0_  = _w2657_ ;
	assign \g37859/_0_  = _w2664_ ;
	assign \g37868/_0_  = _w2670_ ;
	assign \g37869/_0_  = _w2676_ ;
	assign \g37870/_0_  = _w2682_ ;
	assign \g37872/_0_  = _w2704_ ;
	assign \g37886/_0_  = _w2710_ ;
	assign \g37887/_0_  = _w2716_ ;
	assign \g37889/_0_  = _w2722_ ;
	assign \g37897/_0_  = _w2728_ ;
	assign \g37899/_0_  = _w2734_ ;
	assign \g37900/_0_  = _w2740_ ;
	assign \g37907/_0_  = _w2745_ ;
	assign \g37925/_0_  = _w2778_ ;
	assign \g37927/_0_  = _w2906_ ;
	assign \g37928/_0_  = _w2919_ ;
	assign \g37929/_0_  = _w2923_ ;
	assign \g37930/_0_  = _w2932_ ;
	assign \g37932/_0_  = _w2947_ ;
	assign \g37933/_0_  = _w2958_ ;
	assign \g37934/_0_  = _w2970_ ;
	assign \g37935/_0_  = _w2981_ ;
	assign \g37936/_0_  = _w2991_ ;
	assign \g37937/_0_  = _w3001_ ;
	assign \g37938/_0_  = _w3010_ ;
	assign \g37939/_0_  = _w3022_ ;
	assign \g37941/_0_  = _w3030_ ;
	assign \g37942/_0_  = _w3036_ ;
	assign \g37943/_0_  = _w3042_ ;
	assign \g37944/_0_  = _w3048_ ;
	assign \g37945/_0_  = _w3054_ ;
	assign \g38030/_3_  = _w3181_ ;
	assign \g38035/_0_  = _w3189_ ;
	assign \g38036/_0_  = _w3195_ ;
	assign \g38054/_0_  = _w3198_ ;
	assign \g38129/_0_  = _w3202_ ;
	assign \g38130/_0_  = _w3235_ ;
	assign \g38148/_3_  = _w3249_ ;
	assign \g38149/_3_  = _w3266_ ;
	assign \g38150/_3_  = _w3277_ ;
	assign \g38166/_0_  = _w3286_ ;
	assign \g38198/_0_  = _w3290_ ;
	assign \g38201/_0_  = _w3316_ ;
	assign \g38257/_0_  = _w3321_ ;
	assign \g38286/_0_  = _w3338_ ;
	assign \g38294/_3_  = _w3349_ ;
	assign \g38295/_3_  = _w3357_ ;
	assign \g38296/_3_  = _w3366_ ;
	assign \g38297/_3_  = _w3373_ ;
	assign \g38332/_0_  = _w3374_ ;
	assign \g38350/_0_  = _w3375_ ;
	assign \g38365/_3_  = _w3380_ ;
	assign \g38366/_3_  = _w3386_ ;
	assign \g38367/_3_  = _w3393_ ;
	assign \g38389/_0_  = _w3394_ ;
	assign \g38397/_0_  = _w3400_ ;
	assign \g38398/_0_  = _w3406_ ;
	assign \g38399/_0_  = _w3412_ ;
	assign \g38400/_0_  = _w3418_ ;
	assign \g38417/_3_  = _w3425_ ;
	assign \g38418/_3_  = _w3436_ ;
	assign \g38422/_0_  = _w3473_ ;
	assign \g38440/_0_  = _w3483_ ;
	assign \g38443/_0_  = _w3495_ ;
	assign \g38448/_3_  = _w3496_ ;
	assign \g38449/_0_  = _w3501_ ;
	assign \g38450/_0_  = _w3516_ ;
	assign \g38460/_0_  = _w3585_ ;
	assign \g38466/_0_  = _w3588_ ;
	assign \g38467/_0_  = _w3591_ ;
	assign \g38468/_0_  = _w3594_ ;
	assign \g38469/_0_  = _w3598_ ;
	assign \g38470/_0_  = _w3601_ ;
	assign \g38471/_0_  = _w3605_ ;
	assign \g38472/_0_  = _w3608_ ;
	assign \g38473/_0_  = _w3611_ ;
	assign \g38474/_0_  = _w3615_ ;
	assign \g38475/_0_  = _w3618_ ;
	assign \g38476/_0_  = _w3622_ ;
	assign \g38477/_0_  = _w3626_ ;
	assign \g38478/_0_  = _w3632_ ;
	assign \g38479/_0_  = _w3635_ ;
	assign \g38528/_0_  = _w3637_ ;
	assign \g38533/_0_  = _w3643_ ;
	assign \g38534/_0_  = _w3644_ ;
	assign \g38536/_0_  = _w3650_ ;
	assign \g38545/_0_  = _w3658_ ;
	assign \g38551/_0_  = _w3476_ ;
	assign \g38554/_0_  = _w3662_ ;
	assign \g38555/_0_  = _w3667_ ;
	assign \g38556/_0_  = _w3752_ ;
	assign \g38575/_0_  = _w3753_ ;
	assign \g38616/_0_  = _w3754_ ;
	assign \g38653/_0_  = _w3778_ ;
	assign \g38656/_0_  = _w3798_ ;
	assign \g38657/_0_  = _w3818_ ;
	assign \g38658/_0_  = _w3838_ ;
	assign \g38660/_0_  = _w3858_ ;
	assign \g38706/_0_  = _w3869_ ;
	assign \g38716/_0_  = _w3881_ ;
	assign \g38717/_0_  = _w3885_ ;
	assign \g38738/_1_  = _w1756_ ;
	assign \g38763/_0_  = _w3888_ ;
	assign \g38790/_0_  = _w3891_ ;
	assign \g38792/_0_  = _w3894_ ;
	assign \g38801/_0_  = _w3897_ ;
	assign \g38803/_0_  = _w3900_ ;
	assign \g38804/_0_  = _w3907_ ;
	assign \g38805/_0_  = _w3913_ ;
	assign \g38806/_0_  = _w3927_ ;
	assign \g38807/_0_  = _w3935_ ;
	assign \g38808/_0_  = _w3943_ ;
	assign \g38809/_0_  = _w3951_ ;
	assign \g38810/_0_  = _w3959_ ;
	assign \g38814/_0_  = _w3974_ ;
	assign \g38833/_0_  = _w3980_ ;
	assign \g38834/_0_  = _w3984_ ;
	assign \g38839/_0_  = _w3990_ ;
	assign \g38840/_0_  = _w3996_ ;
	assign \g38841/_0_  = _w4002_ ;
	assign \g38842/_0_  = _w4008_ ;
	assign \g38846/_0_  = _w4013_ ;
	assign \g38847/_0_  = _w4019_ ;
	assign \g38848/_0_  = _w4026_ ;
	assign \g38849/_0_  = _w4032_ ;
	assign \g38853/_0_  = _w4040_ ;
	assign \g38857/_0_  = _w4042_ ;
	assign \g38872/_0_  = _w4092_ ;
	assign \g38882/_0_  = _w4124_ ;
	assign \g38884/_0_  = _w4141_ ;
	assign \g38885/_0_  = _w4158_ ;
	assign \g38886/_0_  = _w4175_ ;
	assign \g38887/_0_  = _w4192_ ;
	assign \g38931/_0_  = _w4197_ ;
	assign \g38952/_0_  = _w4201_ ;
	assign \g38960/_0_  = _w4218_ ;
	assign \g38971/_0_  = _w4221_ ;
	assign \g38973/_0_  = _w4223_ ;
	assign \g38974/_0_  = _w4224_ ;
	assign \g38975/_0_  = _w4227_ ;
	assign \g38976/_0_  = _w4230_ ;
	assign \g38978/_0_  = _w4232_ ;
	assign \g38981/_0_  = _w4234_ ;
	assign \g38986/_0_  = _w4236_ ;
	assign \g38987/_0_  = _w4242_ ;
	assign \g39001/_3_  = _w4244_ ;
	assign \g39003/_3_  = _w4245_ ;
	assign \g39009/_3_  = _w4247_ ;
	assign \g39011/_3_  = _w4249_ ;
	assign \g39013/_3_  = _w4251_ ;
	assign \g39015/_2_  = _w4253_ ;
	assign \g39017/_2_  = _w4255_ ;
	assign \g39019/_2_  = _w4257_ ;
	assign \g39021/_2_  = _w4259_ ;
	assign \g39060/_0_  = _w4264_ ;
	assign \g39061/_3_  = _w4265_ ;
	assign \g39062/_0_  = _w4266_ ;
	assign \g39063/_0_  = _w4271_ ;
	assign \g39065/_0_  = _w4278_ ;
	assign \g39066/_0_  = _w4285_ ;
	assign \g39093/_0_  = _w4314_ ;
	assign \g39099/_2_  = _w4364_ ;
	assign \g39118/_0_  = _w4371_ ;
	assign \g39123/_0_  = _w4382_ ;
	assign \g39174/_0_  = _w4414_ ;
	assign \g39175/_0_  = _w4446_ ;
	assign \g39176/_0_  = _w4481_ ;
	assign \g39177/_0_  = _w4514_ ;
	assign \g39178/_0_  = _w4518_ ;
	assign \g39185/_0_  = _w4520_ ;
	assign \g39186/_0_  = _w4523_ ;
	assign \g39187/_0_  = _w4526_ ;
	assign \g39188/_0_  = _w4528_ ;
	assign \g39194/_0_  = _w4529_ ;
	assign \g39195/_0_  = _w4530_ ;
	assign \g39196/_0_  = _w4531_ ;
	assign \g39197/_0_  = _w4532_ ;
	assign \g39198/_0_  = _w4533_ ;
	assign \g39199/_0_  = _w4534_ ;
	assign \g39200/_0_  = _w4535_ ;
	assign \g39201/_0_  = _w4536_ ;
	assign \g39202/_0_  = _w4537_ ;
	assign \g39203/_0_  = _w4538_ ;
	assign \g39204/_0_  = _w4539_ ;
	assign \g39216/_3_  = _w4540_ ;
	assign \g39217/_3_  = _w4541_ ;
	assign \g39218/_0_  = _w4542_ ;
	assign \g39219/_0_  = _w4543_ ;
	assign \g39220/_0_  = _w4548_ ;
	assign \g39221/_0_  = _w4550_ ;
	assign \g39299/_0_  = _w4572_ ;
	assign \g39300/_0_  = _w4595_ ;
	assign \g39301/_0_  = _w4609_ ;
	assign \g39302/_0_  = _w4625_ ;
	assign \g39303/_0_  = _w4632_ ;
	assign \g39304/_0_  = _w4635_ ;
	assign \g39305/_0_  = _w4640_ ;
	assign \g39306/_0_  = _w4646_ ;
	assign \g39307/_0_  = _w4649_ ;
	assign \g39308/_0_  = _w4680_ ;
	assign \g39309/_0_  = _w4710_ ;
	assign \g39310/_0_  = _w4741_ ;
	assign \g39311/_0_  = _w4771_ ;
	assign \g39315/_0_  = _w4772_ ;
	assign \g39318/_0_  = _w4777_ ;
	assign \g39321/_0_  = _w4781_ ;
	assign \g39322/_0_  = _w4782_ ;
	assign \g39323/_0_  = _w4790_ ;
	assign \g39333/_0_  = _w4793_ ;
	assign \g39334/_0_  = _w4796_ ;
	assign \g39336/_0_  = _w4802_ ;
	assign \g39338/_0_  = _w4805_ ;
	assign \g39339/_0_  = _w4809_ ;
	assign \g39340/_0_  = _w4816_ ;
	assign \g39341/_0_  = _w4820_ ;
	assign \g39342/_0_  = _w4827_ ;
	assign \g39343/_0_  = _w4831_ ;
	assign \g39344/_0_  = _w4835_ ;
	assign \g39345/_0_  = _w4840_ ;
	assign \g39346/_0_  = _w4844_ ;
	assign \g39349/_0_  = _w4849_ ;
	assign \g39352/_3_  = _w4853_ ;
	assign \g39354/_3_  = _w4872_ ;
	assign \g39371/_3_  = _w4873_ ;
	assign \g39372/_3_  = _w4874_ ;
	assign \g39373/_3_  = _w4875_ ;
	assign \g39374/_3_  = _w4876_ ;
	assign \g39376/_0_  = _w4878_ ;
	assign \g39377/_0_  = _w4880_ ;
	assign \g39471/_0_  = _w4891_ ;
	assign \g39472/_0_  = _w4905_ ;
	assign \g39473/_0_  = _w4919_ ;
	assign \g39474/_0_  = _w4934_ ;
	assign \g39475/_0_  = _w4948_ ;
	assign \g39476/_0_  = _w4968_ ;
	assign \g39477/_0_  = _w4978_ ;
	assign \g39478/_0_  = _w4996_ ;
	assign \g39479/_0_  = _w5012_ ;
	assign \g39480/_0_  = _w5030_ ;
	assign \g39481/_0_  = _w5046_ ;
	assign \g39482/_0_  = _w5060_ ;
	assign \g39483/_0_  = _w5070_ ;
	assign \g39484/_0_  = _w5089_ ;
	assign \g39485/_0_  = _w5107_ ;
	assign \g39486/_0_  = _w5121_ ;
	assign \g39487/_0_  = _w5128_ ;
	assign \g39488/_0_  = _w5133_ ;
	assign \g39492/_0_  = _w5134_ ;
	assign \g39497/_0_  = _w5137_ ;
	assign \g39501/_0_  = _w5140_ ;
	assign \g39502/_0_  = _w5143_ ;
	assign \g39503/_0_  = _w5148_ ;
	assign \g39504/_0_  = _w5151_ ;
	assign \g39505/_0_  = _w5157_ ;
	assign \g39506/_0_  = _w5161_ ;
	assign \g39539/_0_  = _w5168_ ;
	assign \g39541/_0_  = _w5171_ ;
	assign \g39542/_0_  = _w5172_ ;
	assign \g39543/_0_  = _w5174_ ;
	assign \g39544/_0_  = _w5175_ ;
	assign \g39545/_0_  = _w5177_ ;
	assign \g39546/_0_  = _w5180_ ;
	assign \g39547/_0_  = _w5181_ ;
	assign \g39550/_0_  = _w5184_ ;
	assign \g39551/_0_  = _w5188_ ;
	assign \g39563/_0_  = _w5189_ ;
	assign \g39568/_00_  = _w5219_ ;
	assign \g39617/_0_  = _w5220_ ;
	assign \g39618/_0_  = _w5221_ ;
	assign \g39621/_0_  = _w5223_ ;
	assign \g39622/_0_  = _w5230_ ;
	assign \g39623/_0_  = _w5236_ ;
	assign \g39624/_00_  = _w5244_ ;
	assign \g39685/_0_  = _w5249_ ;
	assign \g39690/_0_  = _w5278_ ;
	assign \g39693/_0_  = _w5310_ ;
	assign \g39695/_0_  = _w5316_ ;
	assign \g39697/_0_  = _w5317_ ;
	assign \g39706/_0_  = _w5323_ ;
	assign \g39749/_0_  = _w5330_ ;
	assign \g39750/_0_  = _w5336_ ;
	assign \g39751/_0_  = _w5342_ ;
	assign \g39752/_0_  = _w5348_ ;
	assign \g39753/_0_  = _w5353_ ;
	assign \g39754/_0_  = _w5358_ ;
	assign \g39755/_0_  = _w5364_ ;
	assign \g39756/_0_  = _w5370_ ;
	assign \g39757/_0_  = _w5375_ ;
	assign \g39758/_0_  = _w5380_ ;
	assign \g39759/_0_  = _w5385_ ;
	assign \g39760/_0_  = _w5390_ ;
	assign \g39761/_0_  = _w5395_ ;
	assign \g39762/_0_  = _w5400_ ;
	assign \g39763/_0_  = _w5405_ ;
	assign \g39764/_0_  = _w5410_ ;
	assign \g39765/_0_  = _w5416_ ;
	assign \g39766/_0_  = _w5421_ ;
	assign \g39767/_0_  = _w5426_ ;
	assign \g39768/_0_  = _w5431_ ;
	assign \g39769/_0_  = _w5436_ ;
	assign \g39770/_0_  = _w5441_ ;
	assign \g39772/_0_  = _w5445_ ;
	assign \g39773/_0_  = _w5449_ ;
	assign \g39775/_3_  = _w5455_ ;
	assign \g39776/_3_  = _w5459_ ;
	assign \g39777/_3_  = _w5464_ ;
	assign \g39778/_3_  = _w5468_ ;
	assign \g39779/_3_  = _w5472_ ;
	assign \g39780/_3_  = _w5477_ ;
	assign \g39781/_3_  = _w5482_ ;
	assign \g39782/_3_  = _w5487_ ;
	assign \g39788/_3_  = _w5498_ ;
	assign \g39799/_0_  = _w5500_ ;
	assign \g39800/_0_  = _w5508_ ;
	assign \g39801/_0_  = _w5513_ ;
	assign \g39802/_0_  = _w5516_ ;
	assign \g39927/_0_  = _w5525_ ;
	assign \g39928/_0_  = _w5537_ ;
	assign \g39929/_0_  = _w5549_ ;
	assign \g39930/_0_  = _w5563_ ;
	assign \g39931/_0_  = _w5579_ ;
	assign \g39932/_0_  = _w5592_ ;
	assign \g39933/_0_  = _w5604_ ;
	assign \g39934/_0_  = _w5616_ ;
	assign \g39935/_0_  = _w5629_ ;
	assign \g39936/_0_  = _w5639_ ;
	assign \g39937/_0_  = _w5649_ ;
	assign \g39938/_0_  = _w5659_ ;
	assign \g39939/_0_  = _w5671_ ;
	assign \g39940/_0_  = _w5680_ ;
	assign \g39942/_0_  = _w5695_ ;
	assign \g39943/_0_  = _w5710_ ;
	assign \g39944/_0_  = _w5723_ ;
	assign \g39945/_0_  = _w5737_ ;
	assign \g39956/_0_  = _w5740_ ;
	assign \g39957/_0_  = _w5743_ ;
	assign \g39958/_0_  = _w5746_ ;
	assign \g39959/_0_  = _w5748_ ;
	assign \g39960/_0_  = _w5751_ ;
	assign \g39961/_0_  = _w5752_ ;
	assign \g39962/_0_  = _w5756_ ;
	assign \g39963/_0_  = _w5760_ ;
	assign \g39964/_0_  = _w5775_ ;
	assign \g39969/_0_  = _w5806_ ;
	assign \g39974/_0_  = _w5835_ ;
	assign \g39975/_0_  = _w5836_ ;
	assign \g39993/_0_  = _w5837_ ;
	assign \g39994/_0_  = _w5838_ ;
	assign \g40003/_0_  = _w5867_ ;
	assign \g40004/_0_  = _w5890_ ;
	assign \g40005/_0_  = _w5913_ ;
	assign \g40006/_0_  = _w5936_ ;
	assign \g40016/_0_  = _w5939_ ;
	assign \g40023/_3_  = _w5940_ ;
	assign \g40033/_0_  = _w5942_ ;
	assign \g40034/_0_  = _w5944_ ;
	assign \g40035/_0_  = _w5969_ ;
	assign \g40036/_0_  = _w5994_ ;
	assign \g40037/_0_  = _w6019_ ;
	assign \g40038/_0_  = _w6043_ ;
	assign \g40199/_0_  = _w6056_ ;
	assign \g40200/_0_  = _w6072_ ;
	assign \g40201/_0_  = _w6085_ ;
	assign \g40202/_0_  = _w6099_ ;
	assign \g40203/_0_  = _w6115_ ;
	assign \g40204/_0_  = _w6131_ ;
	assign \g40205/_0_  = _w6146_ ;
	assign \g40206/_0_  = _w6162_ ;
	assign \g40207/_0_  = _w6173_ ;
	assign \g40208/_0_  = _w6184_ ;
	assign \g40209/_0_  = _w6198_ ;
	assign \g40210/_0_  = _w6212_ ;
	assign \g40224/_0_  = _w6226_ ;
	assign \g40225/_0_  = _w6240_ ;
	assign \g40226/_0_  = _w6254_ ;
	assign \g40227/_0_  = _w6268_ ;
	assign \g40234/_0_  = _w6275_ ;
	assign \g40235/_0_  = _w6282_ ;
	assign \g40236/_0_  = _w6289_ ;
	assign \g40237/_0_  = _w6296_ ;
	assign \g40238/_0_  = _w6303_ ;
	assign \g40239/_0_  = _w6310_ ;
	assign \g40240/_0_  = _w6317_ ;
	assign \g40241/_0_  = _w6324_ ;
	assign \g40242/_0_  = _w6331_ ;
	assign \g40243/_0_  = _w6338_ ;
	assign \g40244/_0_  = _w6345_ ;
	assign \g40246/_0_  = _w6352_ ;
	assign \g40247/_0_  = _w6359_ ;
	assign \g40248/_0_  = _w6366_ ;
	assign \g40249/_0_  = _w6373_ ;
	assign \g40250/_0_  = _w6380_ ;
	assign \g40251/_0_  = _w6387_ ;
	assign \g40252/_0_  = _w6394_ ;
	assign \g40253/_0_  = _w6401_ ;
	assign \g40254/_0_  = _w6408_ ;
	assign \g40255/_0_  = _w6415_ ;
	assign \g40257/_0_  = _w6422_ ;
	assign \g40258/_0_  = _w6429_ ;
	assign \g40262/_0_  = _w6437_ ;
	assign \g40264/_0_  = _w6438_ ;
	assign \g40265/_0_  = _w6442_ ;
	assign \g40266/_0_  = _w6448_ ;
	assign \g40267/_0_  = _w6454_ ;
	assign \g40268/_0_  = _w6460_ ;
	assign \g40269/_0_  = _w6466_ ;
	assign \g40270/_0_  = _w6472_ ;
	assign \g40271/_0_  = _w6478_ ;
	assign \g40272/_0_  = _w6484_ ;
	assign \g40273/_0_  = _w6490_ ;
	assign \g40274/_0_  = _w6496_ ;
	assign \g40275/_0_  = _w6502_ ;
	assign \g40276/_0_  = _w6508_ ;
	assign \g40277/_0_  = _w6514_ ;
	assign \g40278/_0_  = _w6520_ ;
	assign \g40280/_2_  = _w6540_ ;
	assign \g40281/_0_  = _w6546_ ;
	assign \g40282/_0_  = _w6552_ ;
	assign \g40283/_0_  = _w6558_ ;
	assign \g40284/_0_  = _w6564_ ;
	assign \g40285/_0_  = _w6570_ ;
	assign \g40286/_0_  = _w6576_ ;
	assign \g40287/_0_  = _w6582_ ;
	assign \g40288/_0_  = _w6588_ ;
	assign \g40289/_0_  = _w6594_ ;
	assign \g40290/_0_  = _w6600_ ;
	assign \g40291/_0_  = _w6605_ ;
	assign \g40297/_0_  = _w6611_ ;
	assign \g40298/_0_  = _w6617_ ;
	assign \g40299/_0_  = _w6623_ ;
	assign \g40300/_0_  = _w6629_ ;
	assign \g40301/_0_  = _w6635_ ;
	assign \g40302/_0_  = _w6641_ ;
	assign \g40303/_0_  = _w6647_ ;
	assign \g40304/_0_  = _w6653_ ;
	assign \g40306/_0_  = _w6659_ ;
	assign \g40307/_0_  = _w6665_ ;
	assign \g40308/_0_  = _w6671_ ;
	assign \g40309/_0_  = _w6677_ ;
	assign \g40310/_0_  = _w6683_ ;
	assign \g40311/_0_  = _w6689_ ;
	assign \g40312/_0_  = _w6695_ ;
	assign \g40313/_0_  = _w6701_ ;
	assign \g40314/_0_  = _w6707_ ;
	assign \g40315/_0_  = _w6713_ ;
	assign \g40316/_0_  = _w6719_ ;
	assign \g40317/_0_  = _w6725_ ;
	assign \g40318/_0_  = _w6731_ ;
	assign \g40319/_0_  = _w6737_ ;
	assign \g40320/_0_  = _w6743_ ;
	assign \g40324/_0_  = _w4527_ ;
	assign \g40325/_0_  = _w6749_ ;
	assign \g40326/_0_  = _w6755_ ;
	assign \g40327/_0_  = _w6761_ ;
	assign \g40328/_0_  = _w6767_ ;
	assign \g40329/_0_  = _w6773_ ;
	assign \g40330/_0_  = _w6779_ ;
	assign \g40331/_0_  = _w6785_ ;
	assign \g40332/_0_  = _w6791_ ;
	assign \g40333/_0_  = _w6797_ ;
	assign \g40334/_0_  = _w6803_ ;
	assign \g40335/_0_  = _w6809_ ;
	assign \g40336/_0_  = _w6815_ ;
	assign \g40337/_0_  = _w6821_ ;
	assign \g40338/_0_  = _w6827_ ;
	assign \g40339/_0_  = _w6833_ ;
	assign \g40340/_0_  = _w6839_ ;
	assign \g40341/_0_  = _w6845_ ;
	assign \g40342/_0_  = _w6851_ ;
	assign \g40343/_0_  = _w6857_ ;
	assign \g40344/_0_  = _w6863_ ;
	assign \g40345/_0_  = _w6869_ ;
	assign \g40346/_0_  = _w6875_ ;
	assign \g40347/_0_  = _w6881_ ;
	assign \g40350/_0_  = _w6889_ ;
	assign \g40353/_0_  = _w6916_ ;
	assign \g40354/_0_  = _w6930_ ;
	assign \g40355/_0_  = _w6941_ ;
	assign \g40374/_0_  = _w6944_ ;
	assign \g40457/_0_  = _w6946_ ;
	assign \g40458/_0_  = _w6949_ ;
	assign \g40549/_0_  = _w6958_ ;
	assign \g40550/_0_  = _w6967_ ;
	assign \g40551/_0_  = _w6970_ ;
	assign \g40552/_0_  = _w6972_ ;
	assign \g40553/_0_  = _w6974_ ;
	assign \g40554/_0_  = _w6977_ ;
	assign \g40556/_0_  = _w6984_ ;
	assign \g40557/_0_  = _w6992_ ;
	assign \g40558/_0_  = _w7003_ ;
	assign \g40559/_0_  = _w7009_ ;
	assign \g40561/_0_  = _w7016_ ;
	assign \g40562/_0_  = _w7024_ ;
	assign \g40563/_0_  = _w7035_ ;
	assign \g40565/_0_  = _w7042_ ;
	assign \g40566/_0_  = _w7050_ ;
	assign \g40567/_0_  = _w7061_ ;
	assign \g40569/_0_  = _w7068_ ;
	assign \g40570/_0_  = _w7076_ ;
	assign \g40571/_0_  = _w7087_ ;
	assign \g40572/_0_  = _w7095_ ;
	assign \g40573/_0_  = _w7106_ ;
	assign \g40574/_0_  = _w7119_ ;
	assign \g40575/_0_  = _w7127_ ;
	assign \g40576/_0_  = _w7138_ ;
	assign \g40577/_0_  = _w7150_ ;
	assign \g40578/_0_  = _w7158_ ;
	assign \g40579/_0_  = _w7169_ ;
	assign \g40580/_0_  = _w7181_ ;
	assign \g40581/_0_  = _w7189_ ;
	assign \g40582/_0_  = _w7200_ ;
	assign \g40583/_0_  = _w7213_ ;
	assign \g40584/_0_  = _w7219_ ;
	assign \g40586/_0_  = _w7226_ ;
	assign \g40587/_0_  = _w7233_ ;
	assign \g40588/_0_  = _w7240_ ;
	assign \g40589/_0_  = _w7247_ ;
	assign \g40591/_0_  = _w7254_ ;
	assign \g40592/_0_  = _w7260_ ;
	assign \g40593/_0_  = _w7266_ ;
	assign \g40594/_0_  = _w7272_ ;
	assign \g40595/_0_  = _w7278_ ;
	assign \g40596/_0_  = _w7284_ ;
	assign \g40597/_0_  = _w7290_ ;
	assign \g40598/_0_  = _w7296_ ;
	assign \g40599/_0_  = _w7302_ ;
	assign \g40600/_0_  = _w7308_ ;
	assign \g40601/_0_  = _w7314_ ;
	assign \g40602/_0_  = _w7320_ ;
	assign \g40603/_0_  = _w7326_ ;
	assign \g40604/_0_  = _w7332_ ;
	assign \g40605/_0_  = _w7338_ ;
	assign \g40606/_0_  = _w7344_ ;
	assign \g40607/_0_  = _w7350_ ;
	assign \g40608/_0_  = _w7356_ ;
	assign \g40609/_0_  = _w7362_ ;
	assign \g40610/_0_  = _w7368_ ;
	assign \g40611/_0_  = _w7374_ ;
	assign \g40612/_0_  = _w7380_ ;
	assign \g40613/_0_  = _w7386_ ;
	assign \g40614/_0_  = _w7392_ ;
	assign \g40617/_0_  = _w7395_ ;
	assign \g40629/_0_  = _w7400_ ;
	assign \g40632/_0_  = _w7405_ ;
	assign \g40633/_0_  = _w7410_ ;
	assign \g40634/_0_  = _w7415_ ;
	assign \g40635/_0_  = _w7420_ ;
	assign \g40636/_0_  = _w7425_ ;
	assign \g40637/_0_  = _w7430_ ;
	assign \g40638/_0_  = _w7435_ ;
	assign \g40639/_0_  = _w7440_ ;
	assign \g40640/_0_  = _w7445_ ;
	assign \g40641/_0_  = _w7450_ ;
	assign \g40642/_0_  = _w7455_ ;
	assign \g40643/_0_  = _w7460_ ;
	assign \g40644/_0_  = _w7465_ ;
	assign \g40645/_0_  = _w7470_ ;
	assign \g40646/_0_  = _w7475_ ;
	assign \g40647/_0_  = _w7480_ ;
	assign \g40648/_0_  = _w7485_ ;
	assign \g40649/_0_  = _w7490_ ;
	assign \g40650/_0_  = _w7495_ ;
	assign \g40651/_0_  = _w7500_ ;
	assign \g40652/_0_  = _w7505_ ;
	assign \g40653/_0_  = _w7510_ ;
	assign \g40654/_0_  = _w7515_ ;
	assign \g40655/_0_  = _w7520_ ;
	assign \g40661/_0_  = _w7523_ ;
	assign \g40663/_0_  = _w7528_ ;
	assign \g40664/_0_  = _w7533_ ;
	assign \g40665/_0_  = _w7538_ ;
	assign \g40666/_0_  = _w7543_ ;
	assign \g40667/_0_  = _w7548_ ;
	assign \g40668/_0_  = _w7553_ ;
	assign \g40669/_0_  = _w7558_ ;
	assign \g40670/_0_  = _w7563_ ;
	assign \g40671/_0_  = _w7568_ ;
	assign \g40672/_0_  = _w7573_ ;
	assign \g40673/_0_  = _w7578_ ;
	assign \g40674/_0_  = _w7583_ ;
	assign \g40675/_0_  = _w7588_ ;
	assign \g40676/_0_  = _w7593_ ;
	assign \g40677/_0_  = _w7598_ ;
	assign \g40678/_0_  = _w7603_ ;
	assign \g40679/_0_  = _w7608_ ;
	assign \g40680/_0_  = _w7613_ ;
	assign \g40681/_0_  = _w7618_ ;
	assign \g40682/_0_  = _w7623_ ;
	assign \g40683/_0_  = _w7628_ ;
	assign \g40684/_0_  = _w7633_ ;
	assign \g40685/_0_  = _w7638_ ;
	assign \g40689/_0_  = _w7641_ ;
	assign \g40690/_0_  = _w7646_ ;
	assign \g40691/_0_  = _w7651_ ;
	assign \g40692/_0_  = _w7656_ ;
	assign \g40693/_0_  = _w7661_ ;
	assign \g40694/_0_  = _w7666_ ;
	assign \g40695/_0_  = _w7671_ ;
	assign \g40696/_0_  = _w7676_ ;
	assign \g40697/_0_  = _w7681_ ;
	assign \g40698/_0_  = _w7686_ ;
	assign \g40699/_0_  = _w7691_ ;
	assign \g40700/_0_  = _w7696_ ;
	assign \g40701/_0_  = _w7701_ ;
	assign \g40702/_0_  = _w7706_ ;
	assign \g40703/_0_  = _w7711_ ;
	assign \g40704/_0_  = _w7716_ ;
	assign \g40705/_0_  = _w7721_ ;
	assign \g40706/_0_  = _w7726_ ;
	assign \g40707/_0_  = _w7731_ ;
	assign \g40708/_0_  = _w7736_ ;
	assign \g40709/_0_  = _w7741_ ;
	assign \g40710/_0_  = _w7746_ ;
	assign \g40711/_0_  = _w7751_ ;
	assign \g40712/_0_  = _w7756_ ;
	assign \g40758/_00_  = _w7758_ ;
	assign \g40759/_0_  = _w7760_ ;
	assign \g40812/_0_  = _w7784_ ;
	assign \g40816/_0_  = _w7786_ ;
	assign \g40817/_0_  = _w7788_ ;
	assign \g40818/_0_  = _w7810_ ;
	assign \g40819/_0_  = _w7812_ ;
	assign \g40820/_0_  = _w7814_ ;
	assign \g40822/_3_  = _w7815_ ;
	assign \g40823/_3_  = _w7816_ ;
	assign \g40824/_3_  = _w7817_ ;
	assign \g40825/_3_  = _w7818_ ;
	assign \g40849/_3_  = _w7819_ ;
	assign \g40915/_0_  = _w7821_ ;
	assign \g40916/_0_  = _w7827_ ;
	assign \g40917/_0_  = _w7829_ ;
	assign \g40920/_0_  = _w7831_ ;
	assign \g40923/_0_  = _w7842_ ;
	assign \g40926/_0_  = _w7844_ ;
	assign \g40927/_0_  = _w7850_ ;
	assign \g40930/_0_  = _w7852_ ;
	assign \g40931/_0_  = _w7858_ ;
	assign \g41138/_0_  = _w7863_ ;
	assign \g41152/_0_  = _w7869_ ;
	assign \g41180/_0_  = _w7874_ ;
	assign \g41185/_0_  = _w7884_ ;
	assign \g41186/_0_  = _w7886_ ;
	assign \g41187/_0_  = _w7888_ ;
	assign \g41189/_0_  = _w7893_ ;
	assign \g41190/_0_  = _w7898_ ;
	assign \g41191/_0_  = _w7903_ ;
	assign \g41192/_0_  = _w7908_ ;
	assign \g41193/_0_  = _w7913_ ;
	assign \g41195/_0_  = _w7919_ ;
	assign \g41199/_0_  = _w7924_ ;
	assign \g41207/_0_  = _w7935_ ;
	assign \g41221/_0_  = _w7939_ ;
	assign \g41226/_0_  = _w7943_ ;
	assign \g41227/_0_  = _w7946_ ;
	assign \g41230/_0_  = _w7950_ ;
	assign \g41231/_0_  = _w7952_ ;
	assign \g41234/_0_  = _w7966_ ;
	assign \g41238/_0_  = _w7968_ ;
	assign \g41239/_0_  = _w7973_ ;
	assign \g41275/_0_  = _w7981_ ;
	assign \g41277/_0_  = _w7986_ ;
	assign \g41278/_0_  = _w7991_ ;
	assign \g41279/_0_  = _w7996_ ;
	assign \g41280/_0_  = _w8001_ ;
	assign \g41281/_0_  = _w8006_ ;
	assign \g41282/_0_  = _w8012_ ;
	assign \g41283/_0_  = _w8017_ ;
	assign \g41284/_0_  = _w8023_ ;
	assign \g41285/_0_  = _w8028_ ;
	assign \g41286/_0_  = _w8033_ ;
	assign \g41287/_0_  = _w8039_ ;
	assign \g41288/_0_  = _w8047_ ;
	assign \g41289/_0_  = _w8053_ ;
	assign \g41291/_3_  = _w8073_ ;
	assign \g41330/_0_  = _w8077_ ;
	assign \g41332/_0_  = _w8086_ ;
	assign \g41334/_0_  = _w8088_ ;
	assign \g41340/_0_  = _w8097_ ;
	assign \g41343/_0_  = _w8099_ ;
	assign \g41345/_0_  = _w8106_ ;
	assign \g41348/_0_  = _w8108_ ;
	assign \g41349/_0_  = _w8116_ ;
	assign \g41350/_0_  = _w8128_ ;
	assign \g41351/_0_  = _w8133_ ;
	assign \g41356/_0_  = _w8151_ ;
	assign \g41394/_0_  = _w8155_ ;
	assign \g41423/_0_  = _w8156_ ;
	assign \g41426/_3_  = _w8157_ ;
	assign \g41427/_3_  = _w8158_ ;
	assign \g41428/_3_  = _w8159_ ;
	assign \g41429/_3_  = _w8160_ ;
	assign \g41430/_3_  = _w8161_ ;
	assign \g41431/_3_  = _w8162_ ;
	assign \g41432/_3_  = _w8163_ ;
	assign \g41433/_3_  = _w8164_ ;
	assign \g41434/_3_  = _w8165_ ;
	assign \g41435/_3_  = _w8166_ ;
	assign \g41436/_3_  = _w8167_ ;
	assign \g41437/_3_  = _w8168_ ;
	assign \g41438/_3_  = _w8169_ ;
	assign \g41439/_3_  = _w8170_ ;
	assign \g41440/_3_  = _w8171_ ;
	assign \g41441/_3_  = _w8172_ ;
	assign \g41442/_0_  = _w8174_ ;
	assign \g41445/_3_  = _w8175_ ;
	assign \g41446/_0_  = _w8176_ ;
	assign \g41449/_0_  = _w8177_ ;
	assign \g41464/_0_  = _w8178_ ;
	assign \g41466/_0_  = _w8179_ ;
	assign \g41468/_0_  = _w8180_ ;
	assign \g41469/_0_  = _w8182_ ;
	assign \g41471/_0_  = _w8183_ ;
	assign \g41795/_0_  = _w8188_ ;
	assign \g41799/_0_  = _w8193_ ;
	assign \g41800/_0_  = _w8200_ ;
	assign \g41801/_0_  = _w8207_ ;
	assign \g41802/_0_  = _w8214_ ;
	assign \g41803/_0_  = _w8221_ ;
	assign \g41804/_0_  = _w8228_ ;
	assign \g41805/_0_  = _w8235_ ;
	assign \g41806/_0_  = _w8242_ ;
	assign \g41807/_0_  = _w8249_ ;
	assign \g41808/_0_  = _w8256_ ;
	assign \g41809/_0_  = _w8263_ ;
	assign \g41810/_0_  = _w8270_ ;
	assign \g41811/_0_  = _w8277_ ;
	assign \g41812/_0_  = _w8284_ ;
	assign \g41814/_0_  = _w8291_ ;
	assign \g41815/_0_  = _w8298_ ;
	assign \g41816/_0_  = _w8305_ ;
	assign \g41817/_0_  = _w8312_ ;
	assign \g41818/_0_  = _w8319_ ;
	assign \g41819/_0_  = _w8326_ ;
	assign \g41820/_0_  = _w8333_ ;
	assign \g41821/_0_  = _w8340_ ;
	assign \g41822/_0_  = _w8347_ ;
	assign \g41823/_0_  = _w8354_ ;
	assign \g41825/_0_  = _w8361_ ;
	assign \g41826/_0_  = _w8368_ ;
	assign \g41827/_0_  = _w8375_ ;
	assign \g41828/_0_  = _w8382_ ;
	assign \g41829/_0_  = _w8389_ ;
	assign \g41830/_0_  = _w8396_ ;
	assign \g41831/_0_  = _w8403_ ;
	assign \g41832/_0_  = _w8410_ ;
	assign \g41833/_0_  = _w8417_ ;
	assign \g41834/_0_  = _w8424_ ;
	assign \g41835/_0_  = _w8431_ ;
	assign \g41836/_0_  = _w8438_ ;
	assign \g41837/_0_  = _w8445_ ;
	assign \g41838/_0_  = _w8452_ ;
	assign \g41839/_0_  = _w8459_ ;
	assign \g41840/_0_  = _w8466_ ;
	assign \g41841/_0_  = _w8473_ ;
	assign \g41842/_0_  = _w8480_ ;
	assign \g41843/_0_  = _w8487_ ;
	assign \g41844/_0_  = _w8494_ ;
	assign \g41845/_0_  = _w8501_ ;
	assign \g41846/_0_  = _w8508_ ;
	assign \g41847/_0_  = _w8515_ ;
	assign \g41848/_0_  = _w8522_ ;
	assign \g41849/_0_  = _w8529_ ;
	assign \g41850/_0_  = _w8536_ ;
	assign \g41851/_0_  = _w8543_ ;
	assign \g41852/_0_  = _w8550_ ;
	assign \g41853/_0_  = _w8557_ ;
	assign \g41854/_0_  = _w8564_ ;
	assign \g41855/_0_  = _w8571_ ;
	assign \g41856/_0_  = _w8578_ ;
	assign \g41857/_0_  = _w8585_ ;
	assign \g41858/_0_  = _w8592_ ;
	assign \g41859/_0_  = _w8599_ ;
	assign \g41860/_0_  = _w8606_ ;
	assign \g41861/_0_  = _w8613_ ;
	assign \g41862/_0_  = _w8620_ ;
	assign \g41863/_0_  = _w8627_ ;
	assign \g41864/_0_  = _w8634_ ;
	assign \g41865/_0_  = _w8641_ ;
	assign \g41866/_0_  = _w8648_ ;
	assign \g41867/_0_  = _w8655_ ;
	assign \g41868/_0_  = _w8662_ ;
	assign \g41869/_0_  = _w8669_ ;
	assign \g41870/_0_  = _w8676_ ;
	assign \g41871/_0_  = _w8683_ ;
	assign \g41872/_0_  = _w8690_ ;
	assign \g41873/_0_  = _w8697_ ;
	assign \g41874/_0_  = _w8704_ ;
	assign \g41875/_0_  = _w8711_ ;
	assign \g41876/_0_  = _w8718_ ;
	assign \g41877/_0_  = _w8725_ ;
	assign \g41878/_0_  = _w8732_ ;
	assign \g41879/_0_  = _w8739_ ;
	assign \g41880/_0_  = _w8746_ ;
	assign \g41881/_0_  = _w8753_ ;
	assign \g41882/_0_  = _w8760_ ;
	assign \g41883/_0_  = _w8767_ ;
	assign \g41884/_0_  = _w8774_ ;
	assign \g41885/_0_  = _w8781_ ;
	assign \g41886/_0_  = _w8788_ ;
	assign \g41887/_0_  = _w8795_ ;
	assign \g41888/_0_  = _w8802_ ;
	assign \g41889/_0_  = _w8809_ ;
	assign \g41890/_0_  = _w8816_ ;
	assign \g41891/_0_  = _w8823_ ;
	assign \g41902/_0_  = _w8828_ ;
	assign \g41904/_0_  = _w8831_ ;
	assign \g41906/_0_  = _w8835_ ;
	assign \g41907/_0_  = _w8841_ ;
	assign \g41954/_0_  = _w8850_ ;
	assign \g41955/_0_  = _w8855_ ;
	assign \g41956/_0_  = _w8860_ ;
	assign \g41957/_0_  = _w8865_ ;
	assign \g41958/_0_  = _w8870_ ;
	assign \g41959/_0_  = _w8875_ ;
	assign \g41960/_0_  = _w8880_ ;
	assign \g41962/_0_  = _w8886_ ;
	assign \g41963/_0_  = _w8891_ ;
	assign \g41964/_0_  = _w8896_ ;
	assign \g41965/_0_  = _w8901_ ;
	assign \g41966/_0_  = _w8906_ ;
	assign \g41967/_0_  = _w8911_ ;
	assign \g41968/_0_  = _w8916_ ;
	assign \g41969/_0_  = _w8921_ ;
	assign \g41970/_0_  = _w8926_ ;
	assign \g41971/_0_  = _w8931_ ;
	assign \g41972/_0_  = _w8936_ ;
	assign \g41973/_0_  = _w8941_ ;
	assign \g41974/_0_  = _w8946_ ;
	assign \g41975/_0_  = _w8951_ ;
	assign \g41976/_0_  = _w8956_ ;
	assign \g41977/_0_  = _w8961_ ;
	assign \g41978/_0_  = _w8966_ ;
	assign \g41979/_0_  = _w8971_ ;
	assign \g42062/_0_  = _w8977_ ;
	assign \g42079/_0_  = _w8979_ ;
	assign \g42142/_0_  = _w8980_ ;
	assign \g42143/_0_  = _w8981_ ;
	assign \g42144/_0_  = _w8982_ ;
	assign \g42154/_0_  = _w8994_ ;
	assign \g42157/_0_  = _w9000_ ;
	assign \g42160/_0_  = _w9001_ ;
	assign \g42181/_0_  = _w9006_ ;
	assign \g42203/_0_  = _w9011_ ;
	assign \g42204/_3_  = _w9012_ ;
	assign \g42205/_3_  = _w9013_ ;
	assign \g42206/_3_  = _w9014_ ;
	assign \g42208/_0_  = _w9016_ ;
	assign \g42220/_0_  = _w9021_ ;
	assign \g42225/_0_  = _w9033_ ;
	assign \g42251/_0_  = _w9040_ ;
	assign \g42273/_0_  = _w9047_ ;
	assign \g42335/_0_  = _w9054_ ;
	assign \g42357/_0_  = _w9061_ ;
	assign \g42380/_0_  = _w9062_ ;
	assign \g42381/_0_  = _w9063_ ;
	assign \g42383/_0_  = _w9064_ ;
	assign \g42386/_0_  = _w9065_ ;
	assign \g42388/_0_  = _w9066_ ;
	assign \g42475/_0_  = _w9070_ ;
	assign \g42476/_0_  = _w9073_ ;
	assign \g42477/_0_  = _w9076_ ;
	assign \g42478/_0_  = _w9079_ ;
	assign \g42479/_0_  = _w9082_ ;
	assign \g42480/_0_  = _w9085_ ;
	assign \g42481/_0_  = _w9088_ ;
	assign \g42482/_0_  = _w9091_ ;
	assign \g42483/_0_  = _w9094_ ;
	assign \g42484/_0_  = _w9097_ ;
	assign \g42485/_0_  = _w9100_ ;
	assign \g42486/_0_  = _w9103_ ;
	assign \g42487/_0_  = _w9107_ ;
	assign \g42488/_0_  = _w9111_ ;
	assign \g42490/_0_  = _w9113_ ;
	assign \g42491/_0_  = _w9115_ ;
	assign \g42493/_0_  = _w9117_ ;
	assign \g42494/_0_  = _w9119_ ;
	assign \g42495/_0_  = _w9121_ ;
	assign \g42496/_0_  = _w9123_ ;
	assign \g42497/_0_  = _w9125_ ;
	assign \g42498/_0_  = _w9127_ ;
	assign \g42499/_0_  = _w9129_ ;
	assign \g42500/_0_  = _w9131_ ;
	assign \g42501/_0_  = _w9133_ ;
	assign \g42502/_0_  = _w9135_ ;
	assign \g42503/_0_  = _w9137_ ;
	assign \g42504/_0_  = _w9139_ ;
	assign \g42505/_0_  = _w9141_ ;
	assign \g42506/_0_  = _w9143_ ;
	assign \g42507/_0_  = _w9145_ ;
	assign \g42508/_0_  = _w9147_ ;
	assign \g42509/_0_  = _w9149_ ;
	assign \g42510/_0_  = _w9151_ ;
	assign \g42511/_0_  = _w9153_ ;
	assign \g42512/_0_  = _w9155_ ;
	assign \g42513/_0_  = _w9157_ ;
	assign \g42514/_0_  = _w9159_ ;
	assign \g42515/_0_  = _w9161_ ;
	assign \g42516/_0_  = _w9163_ ;
	assign \g42517/_0_  = _w9165_ ;
	assign \g42518/_0_  = _w9167_ ;
	assign \g42519/_0_  = _w9169_ ;
	assign \g42521/_0_  = _w9172_ ;
	assign \g42522/_0_  = _w9175_ ;
	assign \g42523/_0_  = _w9178_ ;
	assign \g42524/_0_  = _w9181_ ;
	assign \g42525/_0_  = _w9184_ ;
	assign \g42526/_0_  = _w9187_ ;
	assign \g42527/_0_  = _w9190_ ;
	assign \g42528/_0_  = _w9193_ ;
	assign \g42529/_0_  = _w9196_ ;
	assign \g42530/_0_  = _w9199_ ;
	assign \g42531/_0_  = _w9202_ ;
	assign \g42532/_0_  = _w9205_ ;
	assign \g42533/_0_  = _w9208_ ;
	assign \g42534/_0_  = _w9211_ ;
	assign \g42535/_0_  = _w9213_ ;
	assign \g42536/_0_  = _w9216_ ;
	assign \g42537/_0_  = _w9219_ ;
	assign \g42538/_0_  = _w9222_ ;
	assign \g42539/_0_  = _w9225_ ;
	assign \g42540/_0_  = _w9228_ ;
	assign \g42541/_0_  = _w9231_ ;
	assign \g42542/_0_  = _w9234_ ;
	assign \g42543/_0_  = _w9237_ ;
	assign \g42544/_0_  = _w9240_ ;
	assign \g42545/_0_  = _w9243_ ;
	assign \g42548/_0_  = _w9245_ ;
	assign \g42557/_0_  = _w9264_ ;
	assign \g42564/_0_  = _w9266_ ;
	assign \g42565/_0_  = _w9268_ ;
	assign \g42566/_0_  = _w9270_ ;
	assign \g42567/_0_  = _w9272_ ;
	assign \g42568/_0_  = _w9274_ ;
	assign \g42569/_0_  = _w9276_ ;
	assign \g42570/_0_  = _w9278_ ;
	assign \g42571/_0_  = _w9280_ ;
	assign \g42572/_0_  = _w9282_ ;
	assign \g42573/_0_  = _w9284_ ;
	assign \g42574/_0_  = _w9286_ ;
	assign \g42575/_0_  = _w9288_ ;
	assign \g42576/_0_  = _w9290_ ;
	assign \g42577/_0_  = _w9294_ ;
	assign \g42578/_0_  = _w9296_ ;
	assign \g42581/_0_  = _w9315_ ;
	assign \g42589/_0_  = _w9317_ ;
	assign \g42590/_0_  = _w9319_ ;
	assign \g42591/_0_  = _w9321_ ;
	assign \g42592/_0_  = _w9323_ ;
	assign \g42593/_0_  = _w9325_ ;
	assign \g42594/_0_  = _w9327_ ;
	assign \g42595/_0_  = _w9329_ ;
	assign \g42596/_0_  = _w9331_ ;
	assign \g42597/_0_  = _w9333_ ;
	assign \g42598/_0_  = _w9335_ ;
	assign \g42599/_0_  = _w9337_ ;
	assign \g42600/_0_  = _w9339_ ;
	assign \g42601/_0_  = _w9341_ ;
	assign \g42602/_0_  = _w9343_ ;
	assign \g42603/_0_  = _w9345_ ;
	assign \g42604/_0_  = _w9347_ ;
	assign \g42605/_0_  = _w9349_ ;
	assign \g42606/_0_  = _w9351_ ;
	assign \g42607/_0_  = _w9353_ ;
	assign \g42608/_0_  = _w9355_ ;
	assign \g42609/_0_  = _w9357_ ;
	assign \g42610/_0_  = _w9359_ ;
	assign \g42611/_0_  = _w9361_ ;
	assign \g42612/_0_  = _w9363_ ;
	assign \g42613/_0_  = _w9365_ ;
	assign \g42614/_0_  = _w9367_ ;
	assign \g42615/_0_  = _w9369_ ;
	assign \g42616/_0_  = _w9371_ ;
	assign \g42617/_0_  = _w9373_ ;
	assign \g42618/_0_  = _w9375_ ;
	assign \g42619/_0_  = _w9377_ ;
	assign \g42620/_0_  = _w9379_ ;
	assign \g42622/_0_  = _w9398_ ;
	assign \g42623/_0_  = _w9400_ ;
	assign \g42627/_0_  = _w9402_ ;
	assign \g42628/_0_  = _w9404_ ;
	assign \g42629/_0_  = _w9406_ ;
	assign \g42630/_0_  = _w9408_ ;
	assign \g42631/_0_  = _w9410_ ;
	assign \g42632/_0_  = _w9412_ ;
	assign \g42633/_0_  = _w9414_ ;
	assign \g42634/_0_  = _w9416_ ;
	assign \g42635/_0_  = _w9418_ ;
	assign \g42636/_0_  = _w9420_ ;
	assign \g42637/_0_  = _w9422_ ;
	assign \g42638/_0_  = _w9424_ ;
	assign \g42639/_0_  = _w9426_ ;
	assign \g42640/_0_  = _w9428_ ;
	assign \g42641/_0_  = _w9430_ ;
	assign \g42642/_0_  = _w9432_ ;
	assign \g42643/_0_  = _w9434_ ;
	assign \g42644/_0_  = _w9436_ ;
	assign \g42645/_0_  = _w9438_ ;
	assign \g42646/_0_  = _w9440_ ;
	assign \g42647/_0_  = _w9442_ ;
	assign \g42648/_0_  = _w9444_ ;
	assign \g42649/_0_  = _w9446_ ;
	assign \g42650/_0_  = _w9448_ ;
	assign \g42666/_0_  = _w9450_ ;
	assign \g42667/_0_  = _w9452_ ;
	assign \g42668/_0_  = _w9454_ ;
	assign \g42669/_0_  = _w9456_ ;
	assign \g42670/_0_  = _w9458_ ;
	assign \g42671/_0_  = _w9460_ ;
	assign \g42672/_0_  = _w9462_ ;
	assign \g42673/_0_  = _w9464_ ;
	assign \g42674/_0_  = _w9466_ ;
	assign \g42675/_0_  = _w9468_ ;
	assign \g42676/_0_  = _w9470_ ;
	assign \g42677/_0_  = _w9472_ ;
	assign \g42678/_0_  = _w9474_ ;
	assign \g42680/_0_  = _w9478_ ;
	assign \g42681/_0_  = _w9480_ ;
	assign \g42685/_0_  = _w9482_ ;
	assign \g42686/_0_  = _w9484_ ;
	assign \g42688/_0_  = _w9486_ ;
	assign \g42689/_0_  = _w9488_ ;
	assign \g42690/_0_  = _w9490_ ;
	assign \g42691/_0_  = _w9492_ ;
	assign \g42692/_0_  = _w9494_ ;
	assign \g42693/_0_  = _w9496_ ;
	assign \g42694/_0_  = _w9498_ ;
	assign \g42695/_0_  = _w9500_ ;
	assign \g42696/_0_  = _w9502_ ;
	assign \g42697/_0_  = _w9504_ ;
	assign \g42698/_0_  = _w9506_ ;
	assign \g42699/_0_  = _w9508_ ;
	assign \g42700/_0_  = _w9510_ ;
	assign \g42701/_0_  = _w9512_ ;
	assign \g42702/_0_  = _w9514_ ;
	assign \g42703/_0_  = _w9516_ ;
	assign \g42704/_0_  = _w9518_ ;
	assign \g42705/_0_  = _w9520_ ;
	assign \g42706/_0_  = _w9522_ ;
	assign \g42707/_0_  = _w9524_ ;
	assign \g42708/_0_  = _w9526_ ;
	assign \g42709/_0_  = _w9528_ ;
	assign \g42710/_0_  = _w9530_ ;
	assign \g42711/_0_  = _w9532_ ;
	assign \g42712/_0_  = _w9534_ ;
	assign \g42713/_0_  = _w9536_ ;
	assign \g42715/_0_  = _w9538_ ;
	assign \g42716/_0_  = _w9540_ ;
	assign \g42717/_0_  = _w9542_ ;
	assign \g42718/_0_  = _w9544_ ;
	assign \g42723/_1_  = _w9545_ ;
	assign \g42727/_0_  = _w9547_ ;
	assign \g42728/_0_  = _w9549_ ;
	assign \g42729/_0_  = _w9551_ ;
	assign \g42730/_0_  = _w9553_ ;
	assign \g42731/_0_  = _w9555_ ;
	assign \g42732/_0_  = _w9557_ ;
	assign \g42733/_0_  = _w9559_ ;
	assign \g42734/_0_  = _w9561_ ;
	assign \g42735/_0_  = _w9563_ ;
	assign \g42736/_0_  = _w9565_ ;
	assign \g42737/_0_  = _w9567_ ;
	assign \g42738/_0_  = _w9569_ ;
	assign \g42739/_0_  = _w9571_ ;
	assign \g42740/_0_  = _w9573_ ;
	assign \g42741/_0_  = _w9575_ ;
	assign \g42742/_0_  = _w9577_ ;
	assign \g42743/_0_  = _w9579_ ;
	assign \g42744/_0_  = _w9581_ ;
	assign \g42745/_0_  = _w9583_ ;
	assign \g42746/_0_  = _w9585_ ;
	assign \g42747/_0_  = _w9587_ ;
	assign \g42748/_0_  = _w9589_ ;
	assign \g42749/_0_  = _w9591_ ;
	assign \g42750/_0_  = _w9593_ ;
	assign \g42751/_0_  = _w9595_ ;
	assign \g42754/_0_  = _w9598_ ;
	assign \g42767/_0_  = _w9600_ ;
	assign \g42768/_0_  = _w9609_ ;
	assign \g42772/_0_  = _w9611_ ;
	assign \g42773/_0_  = _w9613_ ;
	assign \g42774/_0_  = _w9615_ ;
	assign \g42775/_0_  = _w9617_ ;
	assign \g42776/_0_  = _w9619_ ;
	assign \g42777/_0_  = _w9621_ ;
	assign \g42778/_0_  = _w9623_ ;
	assign \g42779/_0_  = _w9625_ ;
	assign \g42780/_0_  = _w9627_ ;
	assign \g42781/_0_  = _w9629_ ;
	assign \g42782/_0_  = _w9631_ ;
	assign \g42783/_0_  = _w9633_ ;
	assign \g42784/_0_  = _w9637_ ;
	assign \g42785/_0_  = _w9639_ ;
	assign \g42790/_0_  = _w9641_ ;
	assign \g42791/_0_  = _w9643_ ;
	assign \g42792/_0_  = _w9645_ ;
	assign \g42793/_0_  = _w9647_ ;
	assign \g42794/_0_  = _w9649_ ;
	assign \g42795/_0_  = _w9651_ ;
	assign \g42796/_0_  = _w9653_ ;
	assign \g42797/_0_  = _w9655_ ;
	assign \g42798/_0_  = _w9657_ ;
	assign \g42799/_0_  = _w9659_ ;
	assign \g42800/_0_  = _w9661_ ;
	assign \g42801/_0_  = _w9663_ ;
	assign \g42802/_0_  = _w9665_ ;
	assign \g42803/_0_  = _w9667_ ;
	assign \g42804/_0_  = _w9669_ ;
	assign \g42805/_0_  = _w9671_ ;
	assign \g42806/_0_  = _w9673_ ;
	assign \g42807/_0_  = _w9675_ ;
	assign \g42808/_0_  = _w9677_ ;
	assign \g42809/_0_  = _w9679_ ;
	assign \g42810/_0_  = _w9681_ ;
	assign \g42811/_0_  = _w9683_ ;
	assign \g42812/_0_  = _w9685_ ;
	assign \g42813/_0_  = _w9687_ ;
	assign \g42814/_0_  = _w9689_ ;
	assign \g42815/_0_  = _w9691_ ;
	assign \g42816/_0_  = _w9693_ ;
	assign \g42817/_0_  = _w9695_ ;
	assign \g42818/_0_  = _w9697_ ;
	assign \g42819/_0_  = _w9699_ ;
	assign \g42820/_0_  = _w9701_ ;
	assign \g42821/_0_  = _w9703_ ;
	assign \g42824/_0_  = _w9705_ ;
	assign \g42825/_0_  = _w9707_ ;
	assign \g42826/_0_  = _w9709_ ;
	assign \g42827/_0_  = _w9711_ ;
	assign \g42828/_0_  = _w9713_ ;
	assign \g42829/_0_  = _w9715_ ;
	assign \g42830/_0_  = _w9717_ ;
	assign \g42831/_0_  = _w9719_ ;
	assign \g42832/_0_  = _w9721_ ;
	assign \g42833/_0_  = _w9723_ ;
	assign \g42834/_0_  = _w9725_ ;
	assign \g42835/_0_  = _w9727_ ;
	assign \g42836/_0_  = _w9729_ ;
	assign \g42837/_0_  = _w9731_ ;
	assign \g42838/_0_  = _w9733_ ;
	assign \g42839/_0_  = _w9735_ ;
	assign \g42840/_0_  = _w9737_ ;
	assign \g42841/_0_  = _w9739_ ;
	assign \g42842/_0_  = _w9741_ ;
	assign \g42843/_0_  = _w9743_ ;
	assign \g42844/_0_  = _w9745_ ;
	assign \g42845/_0_  = _w9747_ ;
	assign \g42846/_0_  = _w9749_ ;
	assign \g42907/_0_  = _w9754_ ;
	assign \g42914/_0_  = _w9760_ ;
	assign \g42924/_0_  = _w9762_ ;
	assign \g42925/_0_  = _w9764_ ;
	assign \g42926/_0_  = _w9766_ ;
	assign \g42927/_0_  = _w9769_ ;
	assign \g42928/_0_  = _w9776_ ;
	assign \g42929/_0_  = _w9778_ ;
	assign \g42930/_0_  = _w9800_ ;
	assign \g42931/_0_  = _w9802_ ;
	assign \g42933/_0_  = _w9804_ ;
	assign \g42941/_0_  = _w9806_ ;
	assign \g42947/_0_  = _w9809_ ;
	assign \g42950/_0_  = _w9811_ ;
	assign \g42955/_0_  = _w9813_ ;
	assign \g42956/_0_  = _w9815_ ;
	assign \g42972/_3_  = _w9816_ ;
	assign \g42973/_3_  = _w9817_ ;
	assign \g42974/_3_  = _w9818_ ;
	assign \g43178/_0_  = _w9821_ ;
	assign \g43179/_0_  = _w9826_ ;
	assign \g43184/_0_  = _w9843_ ;
	assign \g43186/_0_  = _w9860_ ;
	assign \g43187/_0_  = _w9877_ ;
	assign \g43190/_0_  = _w9880_ ;
	assign \g43191/_0_  = _w9883_ ;
	assign \g43192/_0_  = _w9886_ ;
	assign \g43202/_0_  = _w9903_ ;
	assign \g43205/_0_  = _w9906_ ;
	assign \g43206/_0_  = _w9909_ ;
	assign \g43207/_0_  = _w9912_ ;
	assign \g43209/_2_  = _w9930_ ;
	assign \g43228/_0_  = _w9933_ ;
	assign \g43233/_0_  = _w9936_ ;
	assign \g43235/_0_  = _w9939_ ;
	assign \g43236/_0_  = _w9942_ ;
	assign \g43237/_0_  = _w9945_ ;
	assign \g43238/_0_  = _w9948_ ;
	assign \g43280/_0_  = _w9954_ ;
	assign \g43287/_0_  = _w9955_ ;
	assign \g43289/_0_  = _w9958_ ;
	assign \g43290/_0_  = _w9961_ ;
	assign \g43291/_0_  = _w9964_ ;
	assign \g43292/_0_  = _w9967_ ;
	assign \g43303/_0_  = _w9968_ ;
	assign \g43311/_0_  = _w9973_ ;
	assign \g43312/_0_  = _w9975_ ;
	assign \g43363/_0_  = _w9993_ ;
	assign \g43364/_0_  = _w10011_ ;
	assign \g43366/_0_  = _w10029_ ;
	assign \g43367/_0_  = _w10047_ ;
	assign \g43370/_0_  = _w10065_ ;
	assign \g43371/_0_  = _w10083_ ;
	assign \g43374/_0_  = _w10101_ ;
	assign \g43413/_0_  = _w10120_ ;
	assign \g43414/_0_  = _w10139_ ;
	assign \g43415/_0_  = _w10158_ ;
	assign \g43416/_0_  = _w10160_ ;
	assign \g43422/_0_  = _w10167_ ;
	assign \g43427/_0_  = _w10187_ ;
	assign \g43428/_0_  = _w10207_ ;
	assign \g43528/_1__syn_2  = _w6901_ ;
	assign \g43630/_0_  = _w10209_ ;
	assign \g43633/_3_  = _w10210_ ;
	assign \g43647/_0_  = _w10217_ ;
	assign \g43648/_0_  = _w10223_ ;
	assign \g43656/_0_  = _w10230_ ;
	assign \g43657/_0_  = _w10236_ ;
	assign \g43667/_0_  = _w10243_ ;
	assign \g43668/_0_  = _w10248_ ;
	assign \g43675/_0_  = _w10255_ ;
	assign \g43678/_0_  = _w10261_ ;
	assign \g43787/_0_  = _w10264_ ;
	assign \g44055/_0_  = _w10265_ ;
	assign \g44092/_0_  = _w10282_ ;
	assign \g44093/_0_  = _w10299_ ;
	assign \g44176/_0_  = _w10316_ ;
	assign \g44181/_0_  = _w10320_ ;
	assign \g44433/_0_  = _w10324_ ;
	assign \g44510/_0_  = _w10329_ ;
	assign \g44515/_2_  = _w10330_ ;
	assign \g44522/_0_  = _w10334_ ;
	assign \g44529/_2_  = _w10335_ ;
	assign \g44537/_2_  = _w10336_ ;
	assign \g44544/_2_  = _w10337_ ;
	assign \g44594/_0_  = _w10338_ ;
	assign \g44695/_0_  = _w10340_ ;
	assign \g44697/_0_  = _w10342_ ;
	assign \g44699/_0_  = _w10344_ ;
	assign \g44700/_0_  = _w10346_ ;
	assign \g44843/_0_  = _w10355_ ;
	assign \g44844/_0_  = _w10364_ ;
	assign \g44879/_0_  = _w10369_ ;
	assign \g44880/_0_  = _w10372_ ;
	assign \g44881/_0_  = _w10375_ ;
	assign \g44882/_0_  = _w10378_ ;
	assign \g44906/_2_  = _w10391_ ;
	assign \g44910/_0_  = _w10404_ ;
	assign \g44912/_0_  = _w10417_ ;
	assign \g44954/_0_  = _w10418_ ;
	assign \g45000/_0_  = _w10422_ ;
	assign \g45001/_0_  = _w10426_ ;
	assign \g45002/_0_  = _w10430_ ;
	assign \g45003/_0_  = _w10434_ ;
	assign \g45021/_1_  = _w4887_ ;
	assign \g45025/_0_  = _w10435_ ;
	assign \g45051/_0_  = _w10438_ ;
	assign \g45104/_0_  = _w10439_ ;
	assign \g45111/_0_  = _w10440_ ;
	assign \g45112/_0_  = _w10441_ ;
	assign \g45116/_0_  = _w10442_ ;
	assign \g45155/_0_  = _w3776_ ;
	assign \g45238/_0_  = _w10443_ ;
	assign \g45239/_0_  = _w10444_ ;
	assign \g45240/_0_  = _w10445_ ;
	assign \g45241/_0_  = _w10446_ ;
	assign \g45249/_0_  = _w10447_ ;
	assign \g45257/_0_  = _w10451_ ;
	assign \g45332/_0_  = _w10452_ ;
	assign \g45334/_0_  = _w10453_ ;
	assign \g45336/_0_  = _w10454_ ;
	assign \g45337/_0_  = _w10455_ ;
	assign \g45342/_0_  = _w10456_ ;
	assign \g45459/_0_  = _w10459_ ;
	assign \g45460/_0_  = _w10461_ ;
	assign \g45466/_0_  = _w10462_ ;
	assign \g45469/_0_  = _w10464_ ;
	assign \g45470/_0_  = _w10465_ ;
	assign \g45474/_0_  = _w10468_ ;
	assign \g45475/_0_  = _w10470_ ;
	assign \g45477/_0_  = _w10471_ ;
	assign \g45481/_0_  = _w10474_ ;
	assign \g45482/_0_  = _w10476_ ;
	assign \g45487/_0_  = _w10479_ ;
	assign \g45488/_0_  = _w10481_ ;
	assign \g45518/_3_  = _w10487_ ;
	assign \g45519/_3_  = _w10493_ ;
	assign \g45520/_3_  = _w10499_ ;
	assign \g45521/_3_  = _w10505_ ;
	assign \g45522/_3_  = _w10511_ ;
	assign \g45523/_3_  = _w10517_ ;
	assign \g45524/_3_  = _w10523_ ;
	assign \g45525/_3_  = _w10529_ ;
	assign \g45526/_3_  = _w10535_ ;
	assign \g45530/_3_  = _w10541_ ;
	assign \g45531/_3_  = _w10547_ ;
	assign \g45532/_3_  = _w10553_ ;
	assign \g45533/_3_  = _w10559_ ;
	assign \g45534/_3_  = _w10565_ ;
	assign \g45535/_3_  = _w10571_ ;
	assign \g45536/_3_  = _w10577_ ;
	assign \g45559/_3_  = _w10583_ ;
	assign \g45596/_0_  = _w10586_ ;
	assign \g45605/_0_  = _w10589_ ;
	assign \g45622/_0_  = _w10592_ ;
	assign \g45623/_0_  = _w10595_ ;
	assign \g45630/_0_  = _w10598_ ;
	assign \g45747/_0_  = _w10599_ ;
	assign \g45753/_0_  = _w10600_ ;
	assign \g45796/_0_  = _w10602_ ;
	assign \g45837/_0_  = _w10611_ ;
	assign \g45882/_0_  = _w10614_ ;
	assign \g45903/_0_  = _w10615_ ;
	assign \g45912/_0_  = _w10363_ ;
	assign \g45946/_0_  = _w10354_ ;
	assign \g45999/_0_  = _w10616_ ;
	assign \g46000/_0_  = _w10617_ ;
	assign \g46001/_0_  = _w10618_ ;
	assign \g46002/_0_  = _w10619_ ;
	assign \g46012/_0_  = _w10620_ ;
	assign \g46014/_0_  = _w10621_ ;
	assign \g46017/_0_  = _w10622_ ;
	assign \g46018/_0_  = _w10623_ ;
	assign \g46021/_0_  = _w10624_ ;
	assign \g46024/_0_  = _w10625_ ;
	assign \g46026/_0_  = _w10626_ ;
	assign \g46029/_0_  = _w10627_ ;
	assign \g46053/_0_  = _w10628_ ;
	assign \g46083/_0_  = _w10631_ ;
	assign \g46093/_0_  = _w10613_ ;
	assign \g46142/_0_  = _w10633_ ;
	assign \g46154/_1__syn_2  = _w6935_ ;
	assign \g46265/_0_  = _w10638_ ;
	assign \g46266/_0_  = _w10643_ ;
	assign \g46268/_0_  = _w10648_ ;
	assign \g46270/_0_  = _w10653_ ;
	assign \g46273/_0_  = _w10658_ ;
	assign \g46274/_0_  = _w10663_ ;
	assign \g46275/_0_  = _w10668_ ;
	assign \g46276/_0_  = _w10673_ ;
	assign \g46278/_0_  = _w10677_ ;
	assign \g46385/_0_  = _w10681_ ;
	assign \g46411/_0_  = _w10685_ ;
	assign \g46414/_0_  = _w10686_ ;
	assign \g46479/_0_  = _w10687_ ;
	assign \g46520/_0_  = _w10688_ ;
	assign \g46521/_0_  = _w10689_ ;
	assign \g46530/_0_  = _w10690_ ;
	assign \g46531/_0_  = _w10691_ ;
	assign \g46597/_0_  = _w10692_ ;
	assign \g46610/_0_  = _w10693_ ;
	assign \g46617/_0_  = _w10694_ ;
	assign \g46632/_0_  = _w10695_ ;
	assign \g46637/_0_  = _w10696_ ;
	assign \g46722/_0_  = _w10697_ ;
	assign \g46723/_0_  = _w10698_ ;
	assign \g46724/_0_  = _w10699_ ;
	assign \g46725/_0_  = _w10700_ ;
	assign \g46813/_0_  = _w3757_ ;
	assign \g46842/_0_  = _w3764_ ;
	assign \g46888/_0_  = _w3683_ ;
	assign \g46891/_0_  = _w10701_ ;
	assign \g46894/_0_  = _w9823_ ;
	assign \g46905/_0_  = _w10702_ ;
	assign \g46940/_0_  = _w10703_ ;
	assign \g46992/_0_  = _w3760_ ;
	assign \g46995/_0_  = _w3772_ ;
	assign \g47037/_3_  = _w10705_ ;
	assign \g47053/_0_  = _w10706_ ;
	assign \g47140/_0_  = _w10709_ ;
	assign \g47155/_3_  = _w10710_ ;
	assign \g47209/_0_  = _w10711_ ;
	assign \g47211/_0_  = _w10712_ ;
	assign \g47213/_0_  = _w10713_ ;
	assign \g47215/_0_  = _w10714_ ;
	assign \g47337/_0_  = _w10715_ ;
	assign \g47433/_0_  = _w10716_ ;
	assign \g47972/_0_  = _w10717_ ;
	assign \g47976/_0_  = _w10718_ ;
	assign \g48081/_0_  = _w10719_ ;
	assign \g48171/_0_  = _w10720_ ;
	assign \g48227/_0_  = _w10721_ ;
	assign \g48234/_1_  = _w2764_ ;
	assign \g48257/_1_  = _w3721_ ;
	assign \g48266/_0_  = _w2116_ ;
	assign \g48281/_0_  = _w10722_ ;
	assign \g48291/_1_  = _w10723_ ;
	assign \g48322/_0_  = _w10724_ ;
	assign \g48345/_0_  = _w10725_ ;
	assign \g48429/_0_  = _w10726_ ;
	assign \g48495/_1_  = _w4111_ ;
	assign \g48549/_0_  = _w4118_ ;
	assign \g48589/_0_  = _w2115_ ;
	assign \g48642/_0_  = _w4116_ ;
	assign \g48722/_0_  = _w10727_ ;
	assign \g48748/_0_  = _w10728_ ;
	assign \g48749/_0_  = _w10729_ ;
	assign \g48763/_0_  = _w10730_ ;
	assign \g48867/_0_  = _w10731_ ;
	assign \g48876/_0_  = _w10732_ ;
	assign \g48880/_0_  = _w10733_ ;
	assign \g49023/_0_  = _w4104_ ;
	assign \g49205/_0_  = _w10734_ ;
	assign \g49314/_0_  = _w10735_ ;
	assign \g49432/_0__syn_2  = _w10736_ ;
	assign \g49512/_0_  = _w10737_ ;
	assign \g49707/_0_  = _w10738_ ;
	assign \g49737/_0_  = _w10739_ ;
	assign \g49831/_0_  = _w10740_ ;
	assign \g49922/_1_  = _w10741_ ;
	assign \g50132/_0_  = _w4107_ ;
	assign \g51376/_0_  = _w1282_ ;
	assign \g51412/_0_  = _w862_ ;
	assign \g51822/_0_  = _w1492_ ;
	assign \g52114/_0_  = _w1072_ ;
	assign \g52156/_0_  = _w103_ ;
	assign \g54427/_0_  = _w2774_ ;
	assign \g54557/_0_  = _w10745_ ;
	assign \g54561/_3_  = _w3923_ ;
	assign \g55079/_0_  = _w10747_ ;
	assign \sram_adr_o[0]_pad  = _w10752_ ;
	assign \sram_adr_o[10]_pad  = _w10755_ ;
	assign \sram_adr_o[11]_pad  = _w10758_ ;
	assign \sram_adr_o[12]_pad  = _w10761_ ;
	assign \sram_adr_o[13]_pad  = _w10764_ ;
	assign \sram_adr_o[14]_pad  = _w10767_ ;
	assign \sram_adr_o[1]_pad  = _w10770_ ;
	assign \sram_adr_o[2]_pad  = _w10773_ ;
	assign \sram_adr_o[3]_pad  = _w10776_ ;
	assign \sram_adr_o[4]_pad  = _w10779_ ;
	assign \sram_adr_o[5]_pad  = _w10782_ ;
	assign \sram_adr_o[6]_pad  = _w10785_ ;
	assign \sram_adr_o[7]_pad  = _w10788_ ;
	assign \sram_adr_o[8]_pad  = _w10791_ ;
	assign \sram_adr_o[9]_pad  = _w10794_ ;
	assign \sram_data_o[0]_pad  = _w10797_ ;
	assign \sram_data_o[10]_pad  = _w10800_ ;
	assign \sram_data_o[11]_pad  = _w10803_ ;
	assign \sram_data_o[12]_pad  = _w10806_ ;
	assign \sram_data_o[13]_pad  = _w10809_ ;
	assign \sram_data_o[14]_pad  = _w10812_ ;
	assign \sram_data_o[15]_pad  = _w10815_ ;
	assign \sram_data_o[16]_pad  = _w10818_ ;
	assign \sram_data_o[17]_pad  = _w10821_ ;
	assign \sram_data_o[18]_pad  = _w10824_ ;
	assign \sram_data_o[19]_pad  = _w10827_ ;
	assign \sram_data_o[1]_pad  = _w10830_ ;
	assign \sram_data_o[20]_pad  = _w10833_ ;
	assign \sram_data_o[21]_pad  = _w10836_ ;
	assign \sram_data_o[22]_pad  = _w10839_ ;
	assign \sram_data_o[23]_pad  = _w10842_ ;
	assign \sram_data_o[24]_pad  = _w10845_ ;
	assign \sram_data_o[25]_pad  = _w10848_ ;
	assign \sram_data_o[26]_pad  = _w10851_ ;
	assign \sram_data_o[27]_pad  = _w10854_ ;
	assign \sram_data_o[28]_pad  = _w10857_ ;
	assign \sram_data_o[29]_pad  = _w10860_ ;
	assign \sram_data_o[2]_pad  = _w10863_ ;
	assign \sram_data_o[30]_pad  = _w10866_ ;
	assign \sram_data_o[31]_pad  = _w10869_ ;
	assign \sram_data_o[3]_pad  = _w10872_ ;
	assign \sram_data_o[4]_pad  = _w10875_ ;
	assign \sram_data_o[5]_pad  = _w10878_ ;
	assign \sram_data_o[6]_pad  = _w10881_ ;
	assign \sram_data_o[7]_pad  = _w10884_ ;
	assign \sram_data_o[8]_pad  = _w10887_ ;
	assign \sram_data_o[9]_pad  = _w10890_ ;
	assign sram_re_o_pad = 1'b1;
	assign sram_we_o_pad = _w10896_ ;
	assign \u4_utmi_vend_ctrl_r_reg[0]/P0001_reg_syn_3  = _w10898_ ;
	assign \u4_utmi_vend_ctrl_r_reg[1]/P0001_reg_syn_3  = _w10899_ ;
	assign \u4_utmi_vend_ctrl_r_reg[2]/P0001_reg_syn_3  = _w10900_ ;
	assign \u4_utmi_vend_ctrl_r_reg[3]/P0001_reg_syn_3  = _w10902_ ;
endmodule;