module top( \P1_BE_n_reg[0]/NET0131  , \P1_BE_n_reg[1]/NET0131  , \P1_BE_n_reg[2]/NET0131  , \P1_BE_n_reg[3]/NET0131  , \P1_ByteEnable_reg[0]/NET0131  , \P1_ByteEnable_reg[1]/NET0131  , \P1_ByteEnable_reg[2]/NET0131  , \P1_ByteEnable_reg[3]/NET0131  , \P1_CodeFetch_reg/NET0131  , \P1_D_C_n_reg/NET0131  , \P1_DataWidth_reg[0]/NET0131  , \P1_DataWidth_reg[1]/NET0131  , \P1_Datao_reg[0]/NET0131  , \P1_Datao_reg[10]/NET0131  , \P1_Datao_reg[11]/NET0131  , \P1_Datao_reg[12]/NET0131  , \P1_Datao_reg[13]/NET0131  , \P1_Datao_reg[14]/NET0131  , \P1_Datao_reg[15]/NET0131  , \P1_Datao_reg[16]/NET0131  , \P1_Datao_reg[17]/NET0131  , \P1_Datao_reg[18]/NET0131  , \P1_Datao_reg[19]/NET0131  , \P1_Datao_reg[1]/NET0131  , \P1_Datao_reg[20]/NET0131  , \P1_Datao_reg[21]/NET0131  , \P1_Datao_reg[22]/NET0131  , \P1_Datao_reg[23]/NET0131  , \P1_Datao_reg[24]/NET0131  , \P1_Datao_reg[25]/NET0131  , \P1_Datao_reg[26]/NET0131  , \P1_Datao_reg[27]/NET0131  , \P1_Datao_reg[28]/NET0131  , \P1_Datao_reg[29]/NET0131  , \P1_Datao_reg[2]/NET0131  , \P1_Datao_reg[30]/NET0131  , \P1_Datao_reg[3]/NET0131  , \P1_Datao_reg[4]/NET0131  , \P1_Datao_reg[5]/NET0131  , \P1_Datao_reg[6]/NET0131  , \P1_Datao_reg[7]/NET0131  , \P1_Datao_reg[8]/NET0131  , \P1_Datao_reg[9]/NET0131  , \P1_EAX_reg[0]/NET0131  , \P1_EAX_reg[10]/NET0131  , \P1_EAX_reg[11]/NET0131  , \P1_EAX_reg[12]/NET0131  , \P1_EAX_reg[13]/NET0131  , \P1_EAX_reg[14]/NET0131  , \P1_EAX_reg[15]/NET0131  , \P1_EAX_reg[16]/NET0131  , \P1_EAX_reg[17]/NET0131  , \P1_EAX_reg[18]/NET0131  , \P1_EAX_reg[19]/NET0131  , \P1_EAX_reg[1]/NET0131  , \P1_EAX_reg[20]/NET0131  , \P1_EAX_reg[21]/NET0131  , \P1_EAX_reg[22]/NET0131  , \P1_EAX_reg[23]/NET0131  , \P1_EAX_reg[24]/NET0131  , \P1_EAX_reg[25]/NET0131  , \P1_EAX_reg[26]/NET0131  , \P1_EAX_reg[27]/NET0131  , \P1_EAX_reg[28]/NET0131  , \P1_EAX_reg[29]/NET0131  , \P1_EAX_reg[2]/NET0131  , \P1_EAX_reg[30]/NET0131  , \P1_EAX_reg[31]/NET0131  , \P1_EAX_reg[3]/NET0131  , \P1_EAX_reg[4]/NET0131  , \P1_EAX_reg[5]/NET0131  , \P1_EAX_reg[6]/NET0131  , \P1_EAX_reg[7]/NET0131  , \P1_EAX_reg[8]/NET0131  , \P1_EAX_reg[9]/NET0131  , \P1_EBX_reg[0]/NET0131  , \P1_EBX_reg[10]/NET0131  , \P1_EBX_reg[11]/NET0131  , \P1_EBX_reg[12]/NET0131  , \P1_EBX_reg[13]/NET0131  , \P1_EBX_reg[14]/NET0131  , \P1_EBX_reg[15]/NET0131  , \P1_EBX_reg[16]/NET0131  , \P1_EBX_reg[17]/NET0131  , \P1_EBX_reg[18]/NET0131  , \P1_EBX_reg[19]/NET0131  , \P1_EBX_reg[1]/NET0131  , \P1_EBX_reg[20]/NET0131  , \P1_EBX_reg[21]/NET0131  , \P1_EBX_reg[22]/NET0131  , \P1_EBX_reg[23]/NET0131  , \P1_EBX_reg[24]/NET0131  , \P1_EBX_reg[25]/NET0131  , \P1_EBX_reg[26]/NET0131  , \P1_EBX_reg[27]/NET0131  , \P1_EBX_reg[28]/NET0131  , \P1_EBX_reg[29]/NET0131  , \P1_EBX_reg[2]/NET0131  , \P1_EBX_reg[30]/NET0131  , \P1_EBX_reg[31]/NET0131  , \P1_EBX_reg[3]/NET0131  , \P1_EBX_reg[4]/NET0131  , \P1_EBX_reg[5]/NET0131  , \P1_EBX_reg[6]/NET0131  , \P1_EBX_reg[7]/NET0131  , \P1_EBX_reg[8]/NET0131  , \P1_EBX_reg[9]/NET0131  , \P1_Flush_reg/NET0131  , \P1_InstAddrPointer_reg[0]/NET0131  , \P1_InstAddrPointer_reg[10]/NET0131  , \P1_InstAddrPointer_reg[11]/NET0131  , \P1_InstAddrPointer_reg[12]/NET0131  , \P1_InstAddrPointer_reg[13]/NET0131  , \P1_InstAddrPointer_reg[14]/NET0131  , \P1_InstAddrPointer_reg[15]/NET0131  , \P1_InstAddrPointer_reg[16]/NET0131  , \P1_InstAddrPointer_reg[17]/NET0131  , \P1_InstAddrPointer_reg[18]/NET0131  , \P1_InstAddrPointer_reg[19]/NET0131  , \P1_InstAddrPointer_reg[1]/NET0131  , \P1_InstAddrPointer_reg[20]/NET0131  , \P1_InstAddrPointer_reg[21]/NET0131  , \P1_InstAddrPointer_reg[22]/NET0131  , \P1_InstAddrPointer_reg[23]/NET0131  , \P1_InstAddrPointer_reg[24]/NET0131  , \P1_InstAddrPointer_reg[25]/NET0131  , \P1_InstAddrPointer_reg[26]/NET0131  , \P1_InstAddrPointer_reg[27]/NET0131  , \P1_InstAddrPointer_reg[28]/NET0131  , \P1_InstAddrPointer_reg[29]/NET0131  , \P1_InstAddrPointer_reg[2]/NET0131  , \P1_InstAddrPointer_reg[30]/NET0131  , \P1_InstAddrPointer_reg[31]/NET0131  , \P1_InstAddrPointer_reg[3]/NET0131  , \P1_InstAddrPointer_reg[4]/NET0131  , \P1_InstAddrPointer_reg[5]/NET0131  , \P1_InstAddrPointer_reg[6]/NET0131  , \P1_InstAddrPointer_reg[7]/NET0131  , \P1_InstAddrPointer_reg[8]/NET0131  , \P1_InstAddrPointer_reg[9]/NET0131  , \P1_InstQueueRd_Addr_reg[0]/NET0131  , \P1_InstQueueRd_Addr_reg[1]/NET0131  , \P1_InstQueueRd_Addr_reg[2]/NET0131  , \P1_InstQueueRd_Addr_reg[3]/NET0131  , \P1_InstQueueWr_Addr_reg[0]/NET0131  , \P1_InstQueueWr_Addr_reg[1]/NET0131  , \P1_InstQueueWr_Addr_reg[2]/NET0131  , \P1_InstQueueWr_Addr_reg[3]/NET0131  , \P1_InstQueue_reg[0][0]/NET0131  , \P1_InstQueue_reg[0][1]/NET0131  , \P1_InstQueue_reg[0][2]/NET0131  , \P1_InstQueue_reg[0][3]/NET0131  , \P1_InstQueue_reg[0][4]/NET0131  , \P1_InstQueue_reg[0][5]/NET0131  , \P1_InstQueue_reg[0][6]/NET0131  , \P1_InstQueue_reg[0][7]/NET0131  , \P1_InstQueue_reg[10][0]/NET0131  , \P1_InstQueue_reg[10][1]/NET0131  , \P1_InstQueue_reg[10][2]/NET0131  , \P1_InstQueue_reg[10][3]/NET0131  , \P1_InstQueue_reg[10][4]/NET0131  , \P1_InstQueue_reg[10][5]/NET0131  , \P1_InstQueue_reg[10][6]/NET0131  , \P1_InstQueue_reg[10][7]/NET0131  , \P1_InstQueue_reg[11][0]/NET0131  , \P1_InstQueue_reg[11][1]/NET0131  , \P1_InstQueue_reg[11][2]/NET0131  , \P1_InstQueue_reg[11][3]/NET0131  , \P1_InstQueue_reg[11][4]/NET0131  , \P1_InstQueue_reg[11][5]/NET0131  , \P1_InstQueue_reg[11][6]/NET0131  , \P1_InstQueue_reg[11][7]/NET0131  , \P1_InstQueue_reg[12][0]/NET0131  , \P1_InstQueue_reg[12][1]/NET0131  , \P1_InstQueue_reg[12][2]/NET0131  , \P1_InstQueue_reg[12][3]/NET0131  , \P1_InstQueue_reg[12][4]/NET0131  , \P1_InstQueue_reg[12][5]/NET0131  , \P1_InstQueue_reg[12][6]/NET0131  , \P1_InstQueue_reg[12][7]/NET0131  , \P1_InstQueue_reg[13][0]/NET0131  , \P1_InstQueue_reg[13][1]/NET0131  , \P1_InstQueue_reg[13][2]/NET0131  , \P1_InstQueue_reg[13][3]/NET0131  , \P1_InstQueue_reg[13][4]/NET0131  , \P1_InstQueue_reg[13][5]/NET0131  , \P1_InstQueue_reg[13][6]/NET0131  , \P1_InstQueue_reg[13][7]/NET0131  , \P1_InstQueue_reg[14][0]/NET0131  , \P1_InstQueue_reg[14][1]/NET0131  , \P1_InstQueue_reg[14][2]/NET0131  , \P1_InstQueue_reg[14][3]/NET0131  , \P1_InstQueue_reg[14][4]/NET0131  , \P1_InstQueue_reg[14][5]/NET0131  , \P1_InstQueue_reg[14][6]/NET0131  , \P1_InstQueue_reg[14][7]/NET0131  , \P1_InstQueue_reg[15][0]/NET0131  , \P1_InstQueue_reg[15][1]/NET0131  , \P1_InstQueue_reg[15][2]/NET0131  , \P1_InstQueue_reg[15][3]/NET0131  , \P1_InstQueue_reg[15][4]/NET0131  , \P1_InstQueue_reg[15][5]/NET0131  , \P1_InstQueue_reg[15][6]/NET0131  , \P1_InstQueue_reg[15][7]/NET0131  , \P1_InstQueue_reg[1][0]/NET0131  , \P1_InstQueue_reg[1][1]/NET0131  , \P1_InstQueue_reg[1][2]/NET0131  , \P1_InstQueue_reg[1][3]/NET0131  , \P1_InstQueue_reg[1][4]/NET0131  , \P1_InstQueue_reg[1][5]/NET0131  , \P1_InstQueue_reg[1][6]/NET0131  , \P1_InstQueue_reg[1][7]/NET0131  , \P1_InstQueue_reg[2][0]/NET0131  , \P1_InstQueue_reg[2][1]/NET0131  , \P1_InstQueue_reg[2][2]/NET0131  , \P1_InstQueue_reg[2][3]/NET0131  , \P1_InstQueue_reg[2][4]/NET0131  , \P1_InstQueue_reg[2][5]/NET0131  , \P1_InstQueue_reg[2][6]/NET0131  , \P1_InstQueue_reg[2][7]/NET0131  , \P1_InstQueue_reg[3][0]/NET0131  , \P1_InstQueue_reg[3][1]/NET0131  , \P1_InstQueue_reg[3][2]/NET0131  , \P1_InstQueue_reg[3][3]/NET0131  , \P1_InstQueue_reg[3][4]/NET0131  , \P1_InstQueue_reg[3][5]/NET0131  , \P1_InstQueue_reg[3][6]/NET0131  , \P1_InstQueue_reg[3][7]/NET0131  , \P1_InstQueue_reg[4][0]/NET0131  , \P1_InstQueue_reg[4][1]/NET0131  , \P1_InstQueue_reg[4][2]/NET0131  , \P1_InstQueue_reg[4][3]/NET0131  , \P1_InstQueue_reg[4][4]/NET0131  , \P1_InstQueue_reg[4][5]/NET0131  , \P1_InstQueue_reg[4][6]/NET0131  , \P1_InstQueue_reg[4][7]/NET0131  , \P1_InstQueue_reg[5][0]/NET0131  , \P1_InstQueue_reg[5][1]/NET0131  , \P1_InstQueue_reg[5][2]/NET0131  , \P1_InstQueue_reg[5][3]/NET0131  , \P1_InstQueue_reg[5][4]/NET0131  , \P1_InstQueue_reg[5][5]/NET0131  , \P1_InstQueue_reg[5][6]/NET0131  , \P1_InstQueue_reg[5][7]/NET0131  , \P1_InstQueue_reg[6][0]/NET0131  , \P1_InstQueue_reg[6][1]/NET0131  , \P1_InstQueue_reg[6][2]/NET0131  , \P1_InstQueue_reg[6][3]/NET0131  , \P1_InstQueue_reg[6][4]/NET0131  , \P1_InstQueue_reg[6][5]/NET0131  , \P1_InstQueue_reg[6][6]/NET0131  , \P1_InstQueue_reg[6][7]/NET0131  , \P1_InstQueue_reg[7][0]/NET0131  , \P1_InstQueue_reg[7][1]/NET0131  , \P1_InstQueue_reg[7][2]/NET0131  , \P1_InstQueue_reg[7][3]/NET0131  , \P1_InstQueue_reg[7][4]/NET0131  , \P1_InstQueue_reg[7][5]/NET0131  , \P1_InstQueue_reg[7][6]/NET0131  , \P1_InstQueue_reg[7][7]/NET0131  , \P1_InstQueue_reg[8][0]/NET0131  , \P1_InstQueue_reg[8][1]/NET0131  , \P1_InstQueue_reg[8][2]/NET0131  , \P1_InstQueue_reg[8][3]/NET0131  , \P1_InstQueue_reg[8][4]/NET0131  , \P1_InstQueue_reg[8][5]/NET0131  , \P1_InstQueue_reg[8][6]/NET0131  , \P1_InstQueue_reg[8][7]/NET0131  , \P1_InstQueue_reg[9][0]/NET0131  , \P1_InstQueue_reg[9][1]/NET0131  , \P1_InstQueue_reg[9][2]/NET0131  , \P1_InstQueue_reg[9][3]/NET0131  , \P1_InstQueue_reg[9][4]/NET0131  , \P1_InstQueue_reg[9][5]/NET0131  , \P1_InstQueue_reg[9][6]/NET0131  , \P1_InstQueue_reg[9][7]/NET0131  , \P1_M_IO_n_reg/NET0131  , \P1_MemoryFetch_reg/NET0131  , \P1_More_reg/NET0131  , \P1_PhyAddrPointer_reg[0]/NET0131  , \P1_PhyAddrPointer_reg[10]/NET0131  , \P1_PhyAddrPointer_reg[11]/NET0131  , \P1_PhyAddrPointer_reg[12]/NET0131  , \P1_PhyAddrPointer_reg[13]/NET0131  , \P1_PhyAddrPointer_reg[14]/NET0131  , \P1_PhyAddrPointer_reg[15]/NET0131  , \P1_PhyAddrPointer_reg[16]/NET0131  , \P1_PhyAddrPointer_reg[17]/NET0131  , \P1_PhyAddrPointer_reg[18]/NET0131  , \P1_PhyAddrPointer_reg[19]/NET0131  , \P1_PhyAddrPointer_reg[1]/NET0131  , \P1_PhyAddrPointer_reg[20]/NET0131  , \P1_PhyAddrPointer_reg[21]/NET0131  , \P1_PhyAddrPointer_reg[22]/NET0131  , \P1_PhyAddrPointer_reg[23]/NET0131  , \P1_PhyAddrPointer_reg[24]/NET0131  , \P1_PhyAddrPointer_reg[25]/NET0131  , \P1_PhyAddrPointer_reg[26]/NET0131  , \P1_PhyAddrPointer_reg[27]/NET0131  , \P1_PhyAddrPointer_reg[28]/NET0131  , \P1_PhyAddrPointer_reg[29]/NET0131  , \P1_PhyAddrPointer_reg[2]/NET0131  , \P1_PhyAddrPointer_reg[30]/NET0131  , \P1_PhyAddrPointer_reg[31]/NET0131  , \P1_PhyAddrPointer_reg[3]/NET0131  , \P1_PhyAddrPointer_reg[4]/NET0131  , \P1_PhyAddrPointer_reg[5]/NET0131  , \P1_PhyAddrPointer_reg[6]/NET0131  , \P1_PhyAddrPointer_reg[7]/NET0131  , \P1_PhyAddrPointer_reg[8]/NET0131  , \P1_PhyAddrPointer_reg[9]/NET0131  , \P1_ReadRequest_reg/NET0131  , \P1_RequestPending_reg/NET0131  , \P1_State2_reg[0]/NET0131  , \P1_State2_reg[1]/NET0131  , \P1_State2_reg[2]/NET0131  , \P1_State2_reg[3]/NET0131  , \P1_State_reg[0]/NET0131  , \P1_State_reg[1]/NET0131  , \P1_State_reg[2]/NET0131  , \P1_W_R_n_reg/NET0131  , \P1_lWord_reg[0]/NET0131  , \P1_lWord_reg[10]/NET0131  , \P1_lWord_reg[11]/NET0131  , \P1_lWord_reg[12]/NET0131  , \P1_lWord_reg[13]/NET0131  , \P1_lWord_reg[14]/NET0131  , \P1_lWord_reg[15]/NET0131  , \P1_lWord_reg[1]/NET0131  , \P1_lWord_reg[2]/NET0131  , \P1_lWord_reg[3]/NET0131  , \P1_lWord_reg[4]/NET0131  , \P1_lWord_reg[5]/NET0131  , \P1_lWord_reg[6]/NET0131  , \P1_lWord_reg[7]/NET0131  , \P1_lWord_reg[8]/NET0131  , \P1_lWord_reg[9]/NET0131  , \P1_rEIP_reg[0]/NET0131  , \P1_rEIP_reg[10]/NET0131  , \P1_rEIP_reg[11]/NET0131  , \P1_rEIP_reg[12]/NET0131  , \P1_rEIP_reg[13]/NET0131  , \P1_rEIP_reg[14]/NET0131  , \P1_rEIP_reg[15]/NET0131  , \P1_rEIP_reg[16]/NET0131  , \P1_rEIP_reg[17]/NET0131  , \P1_rEIP_reg[18]/NET0131  , \P1_rEIP_reg[19]/NET0131  , \P1_rEIP_reg[1]/NET0131  , \P1_rEIP_reg[20]/NET0131  , \P1_rEIP_reg[21]/NET0131  , \P1_rEIP_reg[22]/NET0131  , \P1_rEIP_reg[23]/NET0131  , \P1_rEIP_reg[24]/NET0131  , \P1_rEIP_reg[25]/NET0131  , \P1_rEIP_reg[26]/NET0131  , \P1_rEIP_reg[27]/NET0131  , \P1_rEIP_reg[28]/NET0131  , \P1_rEIP_reg[29]/NET0131  , \P1_rEIP_reg[2]/NET0131  , \P1_rEIP_reg[30]/NET0131  , \P1_rEIP_reg[31]/NET0131  , \P1_rEIP_reg[3]/NET0131  , \P1_rEIP_reg[4]/NET0131  , \P1_rEIP_reg[5]/NET0131  , \P1_rEIP_reg[6]/NET0131  , \P1_rEIP_reg[7]/NET0131  , \P1_rEIP_reg[8]/NET0131  , \P1_rEIP_reg[9]/NET0131  , \P1_uWord_reg[0]/NET0131  , \P1_uWord_reg[10]/NET0131  , \P1_uWord_reg[11]/NET0131  , \P1_uWord_reg[12]/NET0131  , \P1_uWord_reg[13]/NET0131  , \P1_uWord_reg[14]/NET0131  , \P1_uWord_reg[1]/NET0131  , \P1_uWord_reg[2]/NET0131  , \P1_uWord_reg[3]/NET0131  , \P1_uWord_reg[4]/NET0131  , \P1_uWord_reg[5]/NET0131  , \P1_uWord_reg[6]/NET0131  , \P1_uWord_reg[7]/NET0131  , \P1_uWord_reg[8]/NET0131  , \P1_uWord_reg[9]/NET0131  , \P2_ADS_n_reg/NET0131  , \P2_Address_reg[0]/NET0131  , \P2_Address_reg[10]/NET0131  , \P2_Address_reg[11]/NET0131  , \P2_Address_reg[12]/NET0131  , \P2_Address_reg[13]/NET0131  , \P2_Address_reg[14]/NET0131  , \P2_Address_reg[15]/NET0131  , \P2_Address_reg[16]/NET0131  , \P2_Address_reg[17]/NET0131  , \P2_Address_reg[18]/NET0131  , \P2_Address_reg[19]/NET0131  , \P2_Address_reg[1]/NET0131  , \P2_Address_reg[20]/NET0131  , \P2_Address_reg[21]/NET0131  , \P2_Address_reg[22]/NET0131  , \P2_Address_reg[23]/NET0131  , \P2_Address_reg[24]/NET0131  , \P2_Address_reg[25]/NET0131  , \P2_Address_reg[26]/NET0131  , \P2_Address_reg[27]/NET0131  , \P2_Address_reg[28]/NET0131  , \P2_Address_reg[29]/NET0131  , \P2_Address_reg[2]/NET0131  , \P2_Address_reg[3]/NET0131  , \P2_Address_reg[4]/NET0131  , \P2_Address_reg[5]/NET0131  , \P2_Address_reg[6]/NET0131  , \P2_Address_reg[7]/NET0131  , \P2_Address_reg[8]/NET0131  , \P2_Address_reg[9]/NET0131  , \P2_BE_n_reg[0]/NET0131  , \P2_BE_n_reg[1]/NET0131  , \P2_BE_n_reg[2]/NET0131  , \P2_BE_n_reg[3]/NET0131  , \P2_ByteEnable_reg[0]/NET0131  , \P2_ByteEnable_reg[1]/NET0131  , \P2_ByteEnable_reg[2]/NET0131  , \P2_ByteEnable_reg[3]/NET0131  , \P2_CodeFetch_reg/NET0131  , \P2_D_C_n_reg/NET0131  , \P2_DataWidth_reg[0]/NET0131  , \P2_DataWidth_reg[1]/NET0131  , \P2_Datao_reg[0]/NET0131  , \P2_Datao_reg[10]/NET0131  , \P2_Datao_reg[11]/NET0131  , \P2_Datao_reg[12]/NET0131  , \P2_Datao_reg[13]/NET0131  , \P2_Datao_reg[14]/NET0131  , \P2_Datao_reg[15]/NET0131  , \P2_Datao_reg[16]/NET0131  , \P2_Datao_reg[17]/NET0131  , \P2_Datao_reg[18]/NET0131  , \P2_Datao_reg[19]/NET0131  , \P2_Datao_reg[1]/NET0131  , \P2_Datao_reg[20]/NET0131  , \P2_Datao_reg[21]/NET0131  , \P2_Datao_reg[22]/NET0131  , \P2_Datao_reg[23]/NET0131  , \P2_Datao_reg[24]/NET0131  , \P2_Datao_reg[25]/NET0131  , \P2_Datao_reg[26]/NET0131  , \P2_Datao_reg[27]/NET0131  , \P2_Datao_reg[28]/NET0131  , \P2_Datao_reg[29]/NET0131  , \P2_Datao_reg[2]/NET0131  , \P2_Datao_reg[30]/NET0131  , \P2_Datao_reg[3]/NET0131  , \P2_Datao_reg[4]/NET0131  , \P2_Datao_reg[5]/NET0131  , \P2_Datao_reg[6]/NET0131  , \P2_Datao_reg[7]/NET0131  , \P2_Datao_reg[8]/NET0131  , \P2_Datao_reg[9]/NET0131  , \P2_EAX_reg[0]/NET0131  , \P2_EAX_reg[10]/NET0131  , \P2_EAX_reg[11]/NET0131  , \P2_EAX_reg[12]/NET0131  , \P2_EAX_reg[13]/NET0131  , \P2_EAX_reg[14]/NET0131  , \P2_EAX_reg[15]/NET0131  , \P2_EAX_reg[16]/NET0131  , \P2_EAX_reg[17]/NET0131  , \P2_EAX_reg[18]/NET0131  , \P2_EAX_reg[19]/NET0131  , \P2_EAX_reg[1]/NET0131  , \P2_EAX_reg[20]/NET0131  , \P2_EAX_reg[21]/NET0131  , \P2_EAX_reg[22]/NET0131  , \P2_EAX_reg[23]/NET0131  , \P2_EAX_reg[24]/NET0131  , \P2_EAX_reg[25]/NET0131  , \P2_EAX_reg[26]/NET0131  , \P2_EAX_reg[27]/NET0131  , \P2_EAX_reg[28]/NET0131  , \P2_EAX_reg[29]/NET0131  , \P2_EAX_reg[2]/NET0131  , \P2_EAX_reg[30]/NET0131  , \P2_EAX_reg[31]/NET0131  , \P2_EAX_reg[3]/NET0131  , \P2_EAX_reg[4]/NET0131  , \P2_EAX_reg[5]/NET0131  , \P2_EAX_reg[6]/NET0131  , \P2_EAX_reg[7]/NET0131  , \P2_EAX_reg[8]/NET0131  , \P2_EAX_reg[9]/NET0131  , \P2_EBX_reg[0]/NET0131  , \P2_EBX_reg[10]/NET0131  , \P2_EBX_reg[11]/NET0131  , \P2_EBX_reg[12]/NET0131  , \P2_EBX_reg[13]/NET0131  , \P2_EBX_reg[14]/NET0131  , \P2_EBX_reg[15]/NET0131  , \P2_EBX_reg[16]/NET0131  , \P2_EBX_reg[17]/NET0131  , \P2_EBX_reg[18]/NET0131  , \P2_EBX_reg[19]/NET0131  , \P2_EBX_reg[1]/NET0131  , \P2_EBX_reg[20]/NET0131  , \P2_EBX_reg[21]/NET0131  , \P2_EBX_reg[22]/NET0131  , \P2_EBX_reg[23]/NET0131  , \P2_EBX_reg[24]/NET0131  , \P2_EBX_reg[25]/NET0131  , \P2_EBX_reg[26]/NET0131  , \P2_EBX_reg[27]/NET0131  , \P2_EBX_reg[28]/NET0131  , \P2_EBX_reg[29]/NET0131  , \P2_EBX_reg[2]/NET0131  , \P2_EBX_reg[30]/NET0131  , \P2_EBX_reg[31]/NET0131  , \P2_EBX_reg[3]/NET0131  , \P2_EBX_reg[4]/NET0131  , \P2_EBX_reg[5]/NET0131  , \P2_EBX_reg[6]/NET0131  , \P2_EBX_reg[7]/NET0131  , \P2_EBX_reg[8]/NET0131  , \P2_EBX_reg[9]/NET0131  , \P2_Flush_reg/NET0131  , \P2_InstAddrPointer_reg[0]/NET0131  , \P2_InstAddrPointer_reg[10]/NET0131  , \P2_InstAddrPointer_reg[11]/NET0131  , \P2_InstAddrPointer_reg[12]/NET0131  , \P2_InstAddrPointer_reg[13]/NET0131  , \P2_InstAddrPointer_reg[14]/NET0131  , \P2_InstAddrPointer_reg[15]/NET0131  , \P2_InstAddrPointer_reg[16]/NET0131  , \P2_InstAddrPointer_reg[17]/NET0131  , \P2_InstAddrPointer_reg[18]/NET0131  , \P2_InstAddrPointer_reg[19]/NET0131  , \P2_InstAddrPointer_reg[1]/NET0131  , \P2_InstAddrPointer_reg[20]/NET0131  , \P2_InstAddrPointer_reg[21]/NET0131  , \P2_InstAddrPointer_reg[22]/NET0131  , \P2_InstAddrPointer_reg[23]/NET0131  , \P2_InstAddrPointer_reg[24]/NET0131  , \P2_InstAddrPointer_reg[25]/NET0131  , \P2_InstAddrPointer_reg[26]/NET0131  , \P2_InstAddrPointer_reg[27]/NET0131  , \P2_InstAddrPointer_reg[28]/NET0131  , \P2_InstAddrPointer_reg[29]/NET0131  , \P2_InstAddrPointer_reg[2]/NET0131  , \P2_InstAddrPointer_reg[30]/NET0131  , \P2_InstAddrPointer_reg[31]/NET0131  , \P2_InstAddrPointer_reg[3]/NET0131  , \P2_InstAddrPointer_reg[4]/NET0131  , \P2_InstAddrPointer_reg[5]/NET0131  , \P2_InstAddrPointer_reg[6]/NET0131  , \P2_InstAddrPointer_reg[7]/NET0131  , \P2_InstAddrPointer_reg[8]/NET0131  , \P2_InstAddrPointer_reg[9]/NET0131  , \P2_InstQueueRd_Addr_reg[0]/NET0131  , \P2_InstQueueRd_Addr_reg[1]/NET0131  , \P2_InstQueueRd_Addr_reg[2]/NET0131  , \P2_InstQueueRd_Addr_reg[3]/NET0131  , \P2_InstQueueWr_Addr_reg[0]/NET0131  , \P2_InstQueueWr_Addr_reg[1]/NET0131  , \P2_InstQueueWr_Addr_reg[2]/NET0131  , \P2_InstQueueWr_Addr_reg[3]/NET0131  , \P2_InstQueue_reg[0][0]/NET0131  , \P2_InstQueue_reg[0][1]/NET0131  , \P2_InstQueue_reg[0][2]/NET0131  , \P2_InstQueue_reg[0][3]/NET0131  , \P2_InstQueue_reg[0][4]/NET0131  , \P2_InstQueue_reg[0][5]/NET0131  , \P2_InstQueue_reg[0][6]/NET0131  , \P2_InstQueue_reg[0][7]/NET0131  , \P2_InstQueue_reg[10][0]/NET0131  , \P2_InstQueue_reg[10][1]/NET0131  , \P2_InstQueue_reg[10][2]/NET0131  , \P2_InstQueue_reg[10][3]/NET0131  , \P2_InstQueue_reg[10][4]/NET0131  , \P2_InstQueue_reg[10][5]/NET0131  , \P2_InstQueue_reg[10][6]/NET0131  , \P2_InstQueue_reg[10][7]/NET0131  , \P2_InstQueue_reg[11][0]/NET0131  , \P2_InstQueue_reg[11][1]/NET0131  , \P2_InstQueue_reg[11][2]/NET0131  , \P2_InstQueue_reg[11][3]/NET0131  , \P2_InstQueue_reg[11][4]/NET0131  , \P2_InstQueue_reg[11][5]/NET0131  , \P2_InstQueue_reg[11][6]/NET0131  , \P2_InstQueue_reg[11][7]/NET0131  , \P2_InstQueue_reg[12][0]/NET0131  , \P2_InstQueue_reg[12][1]/NET0131  , \P2_InstQueue_reg[12][2]/NET0131  , \P2_InstQueue_reg[12][3]/NET0131  , \P2_InstQueue_reg[12][4]/NET0131  , \P2_InstQueue_reg[12][5]/NET0131  , \P2_InstQueue_reg[12][6]/NET0131  , \P2_InstQueue_reg[12][7]/NET0131  , \P2_InstQueue_reg[13][0]/NET0131  , \P2_InstQueue_reg[13][1]/NET0131  , \P2_InstQueue_reg[13][2]/NET0131  , \P2_InstQueue_reg[13][3]/NET0131  , \P2_InstQueue_reg[13][4]/NET0131  , \P2_InstQueue_reg[13][5]/NET0131  , \P2_InstQueue_reg[13][6]/NET0131  , \P2_InstQueue_reg[13][7]/NET0131  , \P2_InstQueue_reg[14][0]/NET0131  , \P2_InstQueue_reg[14][1]/NET0131  , \P2_InstQueue_reg[14][2]/NET0131  , \P2_InstQueue_reg[14][3]/NET0131  , \P2_InstQueue_reg[14][4]/NET0131  , \P2_InstQueue_reg[14][5]/NET0131  , \P2_InstQueue_reg[14][6]/NET0131  , \P2_InstQueue_reg[14][7]/NET0131  , \P2_InstQueue_reg[15][0]/NET0131  , \P2_InstQueue_reg[15][1]/NET0131  , \P2_InstQueue_reg[15][2]/NET0131  , \P2_InstQueue_reg[15][3]/NET0131  , \P2_InstQueue_reg[15][4]/NET0131  , \P2_InstQueue_reg[15][5]/NET0131  , \P2_InstQueue_reg[15][6]/NET0131  , \P2_InstQueue_reg[15][7]/NET0131  , \P2_InstQueue_reg[1][0]/NET0131  , \P2_InstQueue_reg[1][1]/NET0131  , \P2_InstQueue_reg[1][2]/NET0131  , \P2_InstQueue_reg[1][3]/NET0131  , \P2_InstQueue_reg[1][4]/NET0131  , \P2_InstQueue_reg[1][5]/NET0131  , \P2_InstQueue_reg[1][6]/NET0131  , \P2_InstQueue_reg[1][7]/NET0131  , \P2_InstQueue_reg[2][0]/NET0131  , \P2_InstQueue_reg[2][1]/NET0131  , \P2_InstQueue_reg[2][2]/NET0131  , \P2_InstQueue_reg[2][3]/NET0131  , \P2_InstQueue_reg[2][4]/NET0131  , \P2_InstQueue_reg[2][5]/NET0131  , \P2_InstQueue_reg[2][6]/NET0131  , \P2_InstQueue_reg[2][7]/NET0131  , \P2_InstQueue_reg[3][0]/NET0131  , \P2_InstQueue_reg[3][1]/NET0131  , \P2_InstQueue_reg[3][2]/NET0131  , \P2_InstQueue_reg[3][3]/NET0131  , \P2_InstQueue_reg[3][4]/NET0131  , \P2_InstQueue_reg[3][5]/NET0131  , \P2_InstQueue_reg[3][6]/NET0131  , \P2_InstQueue_reg[3][7]/NET0131  , \P2_InstQueue_reg[4][0]/NET0131  , \P2_InstQueue_reg[4][1]/NET0131  , \P2_InstQueue_reg[4][2]/NET0131  , \P2_InstQueue_reg[4][3]/NET0131  , \P2_InstQueue_reg[4][4]/NET0131  , \P2_InstQueue_reg[4][5]/NET0131  , \P2_InstQueue_reg[4][6]/NET0131  , \P2_InstQueue_reg[4][7]/NET0131  , \P2_InstQueue_reg[5][0]/NET0131  , \P2_InstQueue_reg[5][1]/NET0131  , \P2_InstQueue_reg[5][2]/NET0131  , \P2_InstQueue_reg[5][3]/NET0131  , \P2_InstQueue_reg[5][4]/NET0131  , \P2_InstQueue_reg[5][5]/NET0131  , \P2_InstQueue_reg[5][6]/NET0131  , \P2_InstQueue_reg[5][7]/NET0131  , \P2_InstQueue_reg[6][0]/NET0131  , \P2_InstQueue_reg[6][1]/NET0131  , \P2_InstQueue_reg[6][2]/NET0131  , \P2_InstQueue_reg[6][3]/NET0131  , \P2_InstQueue_reg[6][4]/NET0131  , \P2_InstQueue_reg[6][5]/NET0131  , \P2_InstQueue_reg[6][6]/NET0131  , \P2_InstQueue_reg[6][7]/NET0131  , \P2_InstQueue_reg[7][0]/NET0131  , \P2_InstQueue_reg[7][1]/NET0131  , \P2_InstQueue_reg[7][2]/NET0131  , \P2_InstQueue_reg[7][3]/NET0131  , \P2_InstQueue_reg[7][4]/NET0131  , \P2_InstQueue_reg[7][5]/NET0131  , \P2_InstQueue_reg[7][6]/NET0131  , \P2_InstQueue_reg[7][7]/NET0131  , \P2_InstQueue_reg[8][0]/NET0131  , \P2_InstQueue_reg[8][1]/NET0131  , \P2_InstQueue_reg[8][2]/NET0131  , \P2_InstQueue_reg[8][3]/NET0131  , \P2_InstQueue_reg[8][4]/NET0131  , \P2_InstQueue_reg[8][5]/NET0131  , \P2_InstQueue_reg[8][6]/NET0131  , \P2_InstQueue_reg[8][7]/NET0131  , \P2_InstQueue_reg[9][0]/NET0131  , \P2_InstQueue_reg[9][1]/NET0131  , \P2_InstQueue_reg[9][2]/NET0131  , \P2_InstQueue_reg[9][3]/NET0131  , \P2_InstQueue_reg[9][4]/NET0131  , \P2_InstQueue_reg[9][5]/NET0131  , \P2_InstQueue_reg[9][6]/NET0131  , \P2_InstQueue_reg[9][7]/NET0131  , \P2_M_IO_n_reg/NET0131  , \P2_MemoryFetch_reg/NET0131  , \P2_More_reg/NET0131  , \P2_PhyAddrPointer_reg[0]/NET0131  , \P2_PhyAddrPointer_reg[10]/NET0131  , \P2_PhyAddrPointer_reg[11]/NET0131  , \P2_PhyAddrPointer_reg[12]/NET0131  , \P2_PhyAddrPointer_reg[13]/NET0131  , \P2_PhyAddrPointer_reg[14]/NET0131  , \P2_PhyAddrPointer_reg[15]/NET0131  , \P2_PhyAddrPointer_reg[16]/NET0131  , \P2_PhyAddrPointer_reg[17]/NET0131  , \P2_PhyAddrPointer_reg[18]/NET0131  , \P2_PhyAddrPointer_reg[19]/NET0131  , \P2_PhyAddrPointer_reg[1]/NET0131  , \P2_PhyAddrPointer_reg[20]/NET0131  , \P2_PhyAddrPointer_reg[21]/NET0131  , \P2_PhyAddrPointer_reg[22]/NET0131  , \P2_PhyAddrPointer_reg[23]/NET0131  , \P2_PhyAddrPointer_reg[24]/NET0131  , \P2_PhyAddrPointer_reg[25]/NET0131  , \P2_PhyAddrPointer_reg[26]/NET0131  , \P2_PhyAddrPointer_reg[27]/NET0131  , \P2_PhyAddrPointer_reg[28]/NET0131  , \P2_PhyAddrPointer_reg[29]/NET0131  , \P2_PhyAddrPointer_reg[2]/NET0131  , \P2_PhyAddrPointer_reg[30]/NET0131  , \P2_PhyAddrPointer_reg[31]/NET0131  , \P2_PhyAddrPointer_reg[3]/NET0131  , \P2_PhyAddrPointer_reg[4]/NET0131  , \P2_PhyAddrPointer_reg[5]/NET0131  , \P2_PhyAddrPointer_reg[6]/NET0131  , \P2_PhyAddrPointer_reg[7]/NET0131  , \P2_PhyAddrPointer_reg[8]/NET0131  , \P2_PhyAddrPointer_reg[9]/NET0131  , \P2_ReadRequest_reg/NET0131  , \P2_RequestPending_reg/NET0131  , \P2_State2_reg[0]/NET0131  , \P2_State2_reg[1]/NET0131  , \P2_State2_reg[2]/NET0131  , \P2_State2_reg[3]/NET0131  , \P2_State_reg[0]/NET0131  , \P2_State_reg[1]/NET0131  , \P2_State_reg[2]/NET0131  , \P2_W_R_n_reg/NET0131  , \P2_lWord_reg[0]/NET0131  , \P2_lWord_reg[10]/NET0131  , \P2_lWord_reg[11]/NET0131  , \P2_lWord_reg[12]/NET0131  , \P2_lWord_reg[13]/NET0131  , \P2_lWord_reg[14]/NET0131  , \P2_lWord_reg[15]/NET0131  , \P2_lWord_reg[1]/NET0131  , \P2_lWord_reg[2]/NET0131  , \P2_lWord_reg[3]/NET0131  , \P2_lWord_reg[4]/NET0131  , \P2_lWord_reg[5]/NET0131  , \P2_lWord_reg[6]/NET0131  , \P2_lWord_reg[7]/NET0131  , \P2_lWord_reg[8]/NET0131  , \P2_lWord_reg[9]/NET0131  , \P2_rEIP_reg[0]/NET0131  , \P2_rEIP_reg[10]/NET0131  , \P2_rEIP_reg[11]/NET0131  , \P2_rEIP_reg[12]/NET0131  , \P2_rEIP_reg[13]/NET0131  , \P2_rEIP_reg[14]/NET0131  , \P2_rEIP_reg[15]/NET0131  , \P2_rEIP_reg[16]/NET0131  , \P2_rEIP_reg[17]/NET0131  , \P2_rEIP_reg[18]/NET0131  , \P2_rEIP_reg[19]/NET0131  , \P2_rEIP_reg[1]/NET0131  , \P2_rEIP_reg[20]/NET0131  , \P2_rEIP_reg[21]/NET0131  , \P2_rEIP_reg[22]/NET0131  , \P2_rEIP_reg[23]/NET0131  , \P2_rEIP_reg[24]/NET0131  , \P2_rEIP_reg[25]/NET0131  , \P2_rEIP_reg[26]/NET0131  , \P2_rEIP_reg[27]/NET0131  , \P2_rEIP_reg[28]/NET0131  , \P2_rEIP_reg[29]/NET0131  , \P2_rEIP_reg[2]/NET0131  , \P2_rEIP_reg[30]/NET0131  , \P2_rEIP_reg[31]/NET0131  , \P2_rEIP_reg[3]/NET0131  , \P2_rEIP_reg[4]/NET0131  , \P2_rEIP_reg[5]/NET0131  , \P2_rEIP_reg[6]/NET0131  , \P2_rEIP_reg[7]/NET0131  , \P2_rEIP_reg[8]/NET0131  , \P2_rEIP_reg[9]/NET0131  , \P2_uWord_reg[0]/NET0131  , \P2_uWord_reg[10]/NET0131  , \P2_uWord_reg[11]/NET0131  , \P2_uWord_reg[12]/NET0131  , \P2_uWord_reg[13]/NET0131  , \P2_uWord_reg[14]/NET0131  , \P2_uWord_reg[1]/NET0131  , \P2_uWord_reg[2]/NET0131  , \P2_uWord_reg[3]/NET0131  , \P2_uWord_reg[4]/NET0131  , \P2_uWord_reg[5]/NET0131  , \P2_uWord_reg[6]/NET0131  , \P2_uWord_reg[7]/NET0131  , \P2_uWord_reg[8]/NET0131  , \P2_uWord_reg[9]/NET0131  , \P3_Address_reg[0]/NET0131  , \P3_Address_reg[10]/NET0131  , \P3_Address_reg[11]/NET0131  , \P3_Address_reg[12]/NET0131  , \P3_Address_reg[13]/NET0131  , \P3_Address_reg[14]/NET0131  , \P3_Address_reg[15]/NET0131  , \P3_Address_reg[16]/NET0131  , \P3_Address_reg[17]/NET0131  , \P3_Address_reg[18]/NET0131  , \P3_Address_reg[19]/NET0131  , \P3_Address_reg[1]/NET0131  , \P3_Address_reg[20]/NET0131  , \P3_Address_reg[21]/NET0131  , \P3_Address_reg[22]/NET0131  , \P3_Address_reg[23]/NET0131  , \P3_Address_reg[24]/NET0131  , \P3_Address_reg[25]/NET0131  , \P3_Address_reg[26]/NET0131  , \P3_Address_reg[27]/NET0131  , \P3_Address_reg[28]/NET0131  , \P3_Address_reg[29]/NET0131  , \P3_Address_reg[2]/NET0131  , \P3_Address_reg[3]/NET0131  , \P3_Address_reg[4]/NET0131  , \P3_Address_reg[5]/NET0131  , \P3_Address_reg[6]/NET0131  , \P3_Address_reg[7]/NET0131  , \P3_Address_reg[8]/NET0131  , \P3_Address_reg[9]/NET0131  , \P3_BE_n_reg[0]/NET0131  , \P3_BE_n_reg[1]/NET0131  , \P3_BE_n_reg[2]/NET0131  , \P3_BE_n_reg[3]/NET0131  , \P3_ByteEnable_reg[0]/NET0131  , \P3_ByteEnable_reg[1]/NET0131  , \P3_ByteEnable_reg[2]/NET0131  , \P3_ByteEnable_reg[3]/NET0131  , \P3_CodeFetch_reg/NET0131  , \P3_DataWidth_reg[0]/NET0131  , \P3_DataWidth_reg[1]/NET0131  , \P3_EAX_reg[0]/NET0131  , \P3_EAX_reg[10]/NET0131  , \P3_EAX_reg[11]/NET0131  , \P3_EAX_reg[12]/NET0131  , \P3_EAX_reg[13]/NET0131  , \P3_EAX_reg[14]/NET0131  , \P3_EAX_reg[15]/NET0131  , \P3_EAX_reg[16]/NET0131  , \P3_EAX_reg[17]/NET0131  , \P3_EAX_reg[18]/NET0131  , \P3_EAX_reg[19]/NET0131  , \P3_EAX_reg[1]/NET0131  , \P3_EAX_reg[20]/NET0131  , \P3_EAX_reg[21]/NET0131  , \P3_EAX_reg[22]/NET0131  , \P3_EAX_reg[23]/NET0131  , \P3_EAX_reg[24]/NET0131  , \P3_EAX_reg[25]/NET0131  , \P3_EAX_reg[26]/NET0131  , \P3_EAX_reg[27]/NET0131  , \P3_EAX_reg[28]/NET0131  , \P3_EAX_reg[29]/NET0131  , \P3_EAX_reg[2]/NET0131  , \P3_EAX_reg[30]/NET0131  , \P3_EAX_reg[31]/NET0131  , \P3_EAX_reg[3]/NET0131  , \P3_EAX_reg[4]/NET0131  , \P3_EAX_reg[5]/NET0131  , \P3_EAX_reg[6]/NET0131  , \P3_EAX_reg[7]/NET0131  , \P3_EAX_reg[8]/NET0131  , \P3_EAX_reg[9]/NET0131  , \P3_EBX_reg[0]/NET0131  , \P3_EBX_reg[10]/NET0131  , \P3_EBX_reg[11]/NET0131  , \P3_EBX_reg[12]/NET0131  , \P3_EBX_reg[13]/NET0131  , \P3_EBX_reg[14]/NET0131  , \P3_EBX_reg[15]/NET0131  , \P3_EBX_reg[16]/NET0131  , \P3_EBX_reg[17]/NET0131  , \P3_EBX_reg[18]/NET0131  , \P3_EBX_reg[19]/NET0131  , \P3_EBX_reg[1]/NET0131  , \P3_EBX_reg[20]/NET0131  , \P3_EBX_reg[21]/NET0131  , \P3_EBX_reg[22]/NET0131  , \P3_EBX_reg[23]/NET0131  , \P3_EBX_reg[24]/NET0131  , \P3_EBX_reg[25]/NET0131  , \P3_EBX_reg[26]/NET0131  , \P3_EBX_reg[27]/NET0131  , \P3_EBX_reg[28]/NET0131  , \P3_EBX_reg[29]/NET0131  , \P3_EBX_reg[2]/NET0131  , \P3_EBX_reg[30]/NET0131  , \P3_EBX_reg[31]/NET0131  , \P3_EBX_reg[3]/NET0131  , \P3_EBX_reg[4]/NET0131  , \P3_EBX_reg[5]/NET0131  , \P3_EBX_reg[6]/NET0131  , \P3_EBX_reg[7]/NET0131  , \P3_EBX_reg[8]/NET0131  , \P3_EBX_reg[9]/NET0131  , \P3_Flush_reg/NET0131  , \P3_InstAddrPointer_reg[0]/NET0131  , \P3_InstAddrPointer_reg[10]/NET0131  , \P3_InstAddrPointer_reg[11]/NET0131  , \P3_InstAddrPointer_reg[12]/NET0131  , \P3_InstAddrPointer_reg[13]/NET0131  , \P3_InstAddrPointer_reg[14]/NET0131  , \P3_InstAddrPointer_reg[15]/NET0131  , \P3_InstAddrPointer_reg[16]/NET0131  , \P3_InstAddrPointer_reg[17]/NET0131  , \P3_InstAddrPointer_reg[18]/NET0131  , \P3_InstAddrPointer_reg[19]/NET0131  , \P3_InstAddrPointer_reg[1]/NET0131  , \P3_InstAddrPointer_reg[20]/NET0131  , \P3_InstAddrPointer_reg[21]/NET0131  , \P3_InstAddrPointer_reg[22]/NET0131  , \P3_InstAddrPointer_reg[23]/NET0131  , \P3_InstAddrPointer_reg[24]/NET0131  , \P3_InstAddrPointer_reg[25]/NET0131  , \P3_InstAddrPointer_reg[26]/NET0131  , \P3_InstAddrPointer_reg[27]/NET0131  , \P3_InstAddrPointer_reg[28]/NET0131  , \P3_InstAddrPointer_reg[29]/NET0131  , \P3_InstAddrPointer_reg[2]/NET0131  , \P3_InstAddrPointer_reg[30]/NET0131  , \P3_InstAddrPointer_reg[31]/NET0131  , \P3_InstAddrPointer_reg[3]/NET0131  , \P3_InstAddrPointer_reg[4]/NET0131  , \P3_InstAddrPointer_reg[5]/NET0131  , \P3_InstAddrPointer_reg[6]/NET0131  , \P3_InstAddrPointer_reg[7]/NET0131  , \P3_InstAddrPointer_reg[8]/NET0131  , \P3_InstAddrPointer_reg[9]/NET0131  , \P3_InstQueueRd_Addr_reg[0]/NET0131  , \P3_InstQueueRd_Addr_reg[1]/NET0131  , \P3_InstQueueRd_Addr_reg[2]/NET0131  , \P3_InstQueueRd_Addr_reg[3]/NET0131  , \P3_InstQueueWr_Addr_reg[0]/NET0131  , \P3_InstQueueWr_Addr_reg[1]/NET0131  , \P3_InstQueueWr_Addr_reg[2]/NET0131  , \P3_InstQueueWr_Addr_reg[3]/NET0131  , \P3_InstQueue_reg[0][0]/NET0131  , \P3_InstQueue_reg[0][1]/NET0131  , \P3_InstQueue_reg[0][2]/NET0131  , \P3_InstQueue_reg[0][3]/NET0131  , \P3_InstQueue_reg[0][4]/NET0131  , \P3_InstQueue_reg[0][5]/NET0131  , \P3_InstQueue_reg[0][6]/NET0131  , \P3_InstQueue_reg[0][7]/NET0131  , \P3_InstQueue_reg[10][0]/NET0131  , \P3_InstQueue_reg[10][1]/NET0131  , \P3_InstQueue_reg[10][2]/NET0131  , \P3_InstQueue_reg[10][3]/NET0131  , \P3_InstQueue_reg[10][4]/NET0131  , \P3_InstQueue_reg[10][5]/NET0131  , \P3_InstQueue_reg[10][6]/NET0131  , \P3_InstQueue_reg[10][7]/NET0131  , \P3_InstQueue_reg[11][0]/NET0131  , \P3_InstQueue_reg[11][1]/NET0131  , \P3_InstQueue_reg[11][2]/NET0131  , \P3_InstQueue_reg[11][3]/NET0131  , \P3_InstQueue_reg[11][4]/NET0131  , \P3_InstQueue_reg[11][5]/NET0131  , \P3_InstQueue_reg[11][6]/NET0131  , \P3_InstQueue_reg[11][7]/NET0131  , \P3_InstQueue_reg[12][0]/NET0131  , \P3_InstQueue_reg[12][1]/NET0131  , \P3_InstQueue_reg[12][2]/NET0131  , \P3_InstQueue_reg[12][3]/NET0131  , \P3_InstQueue_reg[12][4]/NET0131  , \P3_InstQueue_reg[12][5]/NET0131  , \P3_InstQueue_reg[12][6]/NET0131  , \P3_InstQueue_reg[12][7]/NET0131  , \P3_InstQueue_reg[13][0]/NET0131  , \P3_InstQueue_reg[13][1]/NET0131  , \P3_InstQueue_reg[13][2]/NET0131  , \P3_InstQueue_reg[13][3]/NET0131  , \P3_InstQueue_reg[13][4]/NET0131  , \P3_InstQueue_reg[13][5]/NET0131  , \P3_InstQueue_reg[13][6]/NET0131  , \P3_InstQueue_reg[13][7]/NET0131  , \P3_InstQueue_reg[14][0]/NET0131  , \P3_InstQueue_reg[14][1]/NET0131  , \P3_InstQueue_reg[14][2]/NET0131  , \P3_InstQueue_reg[14][3]/NET0131  , \P3_InstQueue_reg[14][4]/NET0131  , \P3_InstQueue_reg[14][5]/NET0131  , \P3_InstQueue_reg[14][6]/NET0131  , \P3_InstQueue_reg[14][7]/NET0131  , \P3_InstQueue_reg[15][0]/NET0131  , \P3_InstQueue_reg[15][1]/NET0131  , \P3_InstQueue_reg[15][2]/NET0131  , \P3_InstQueue_reg[15][3]/NET0131  , \P3_InstQueue_reg[15][4]/NET0131  , \P3_InstQueue_reg[15][5]/NET0131  , \P3_InstQueue_reg[15][6]/NET0131  , \P3_InstQueue_reg[15][7]/NET0131  , \P3_InstQueue_reg[1][0]/NET0131  , \P3_InstQueue_reg[1][1]/NET0131  , \P3_InstQueue_reg[1][2]/NET0131  , \P3_InstQueue_reg[1][3]/NET0131  , \P3_InstQueue_reg[1][4]/NET0131  , \P3_InstQueue_reg[1][5]/NET0131  , \P3_InstQueue_reg[1][6]/NET0131  , \P3_InstQueue_reg[1][7]/NET0131  , \P3_InstQueue_reg[2][0]/NET0131  , \P3_InstQueue_reg[2][1]/NET0131  , \P3_InstQueue_reg[2][2]/NET0131  , \P3_InstQueue_reg[2][3]/NET0131  , \P3_InstQueue_reg[2][4]/NET0131  , \P3_InstQueue_reg[2][5]/NET0131  , \P3_InstQueue_reg[2][6]/NET0131  , \P3_InstQueue_reg[2][7]/NET0131  , \P3_InstQueue_reg[3][0]/NET0131  , \P3_InstQueue_reg[3][1]/NET0131  , \P3_InstQueue_reg[3][2]/NET0131  , \P3_InstQueue_reg[3][3]/NET0131  , \P3_InstQueue_reg[3][4]/NET0131  , \P3_InstQueue_reg[3][5]/NET0131  , \P3_InstQueue_reg[3][6]/NET0131  , \P3_InstQueue_reg[3][7]/NET0131  , \P3_InstQueue_reg[4][0]/NET0131  , \P3_InstQueue_reg[4][1]/NET0131  , \P3_InstQueue_reg[4][2]/NET0131  , \P3_InstQueue_reg[4][3]/NET0131  , \P3_InstQueue_reg[4][4]/NET0131  , \P3_InstQueue_reg[4][5]/NET0131  , \P3_InstQueue_reg[4][6]/NET0131  , \P3_InstQueue_reg[4][7]/NET0131  , \P3_InstQueue_reg[5][0]/NET0131  , \P3_InstQueue_reg[5][1]/NET0131  , \P3_InstQueue_reg[5][2]/NET0131  , \P3_InstQueue_reg[5][3]/NET0131  , \P3_InstQueue_reg[5][4]/NET0131  , \P3_InstQueue_reg[5][5]/NET0131  , \P3_InstQueue_reg[5][6]/NET0131  , \P3_InstQueue_reg[5][7]/NET0131  , \P3_InstQueue_reg[6][0]/NET0131  , \P3_InstQueue_reg[6][1]/NET0131  , \P3_InstQueue_reg[6][2]/NET0131  , \P3_InstQueue_reg[6][3]/NET0131  , \P3_InstQueue_reg[6][4]/NET0131  , \P3_InstQueue_reg[6][5]/NET0131  , \P3_InstQueue_reg[6][6]/NET0131  , \P3_InstQueue_reg[6][7]/NET0131  , \P3_InstQueue_reg[7][0]/NET0131  , \P3_InstQueue_reg[7][1]/NET0131  , \P3_InstQueue_reg[7][2]/NET0131  , \P3_InstQueue_reg[7][3]/NET0131  , \P3_InstQueue_reg[7][4]/NET0131  , \P3_InstQueue_reg[7][5]/NET0131  , \P3_InstQueue_reg[7][6]/NET0131  , \P3_InstQueue_reg[7][7]/NET0131  , \P3_InstQueue_reg[8][0]/NET0131  , \P3_InstQueue_reg[8][1]/NET0131  , \P3_InstQueue_reg[8][2]/NET0131  , \P3_InstQueue_reg[8][3]/NET0131  , \P3_InstQueue_reg[8][4]/NET0131  , \P3_InstQueue_reg[8][5]/NET0131  , \P3_InstQueue_reg[8][6]/NET0131  , \P3_InstQueue_reg[8][7]/NET0131  , \P3_InstQueue_reg[9][0]/NET0131  , \P3_InstQueue_reg[9][1]/NET0131  , \P3_InstQueue_reg[9][2]/NET0131  , \P3_InstQueue_reg[9][3]/NET0131  , \P3_InstQueue_reg[9][4]/NET0131  , \P3_InstQueue_reg[9][5]/NET0131  , \P3_InstQueue_reg[9][6]/NET0131  , \P3_InstQueue_reg[9][7]/NET0131  , \P3_MemoryFetch_reg/NET0131  , \P3_More_reg/NET0131  , \P3_PhyAddrPointer_reg[0]/NET0131  , \P3_PhyAddrPointer_reg[10]/NET0131  , \P3_PhyAddrPointer_reg[11]/NET0131  , \P3_PhyAddrPointer_reg[12]/NET0131  , \P3_PhyAddrPointer_reg[13]/NET0131  , \P3_PhyAddrPointer_reg[14]/NET0131  , \P3_PhyAddrPointer_reg[15]/NET0131  , \P3_PhyAddrPointer_reg[16]/NET0131  , \P3_PhyAddrPointer_reg[17]/NET0131  , \P3_PhyAddrPointer_reg[18]/NET0131  , \P3_PhyAddrPointer_reg[19]/NET0131  , \P3_PhyAddrPointer_reg[1]/NET0131  , \P3_PhyAddrPointer_reg[20]/NET0131  , \P3_PhyAddrPointer_reg[21]/NET0131  , \P3_PhyAddrPointer_reg[22]/NET0131  , \P3_PhyAddrPointer_reg[23]/NET0131  , \P3_PhyAddrPointer_reg[24]/NET0131  , \P3_PhyAddrPointer_reg[25]/NET0131  , \P3_PhyAddrPointer_reg[26]/NET0131  , \P3_PhyAddrPointer_reg[27]/NET0131  , \P3_PhyAddrPointer_reg[28]/NET0131  , \P3_PhyAddrPointer_reg[29]/NET0131  , \P3_PhyAddrPointer_reg[2]/NET0131  , \P3_PhyAddrPointer_reg[30]/NET0131  , \P3_PhyAddrPointer_reg[31]/NET0131  , \P3_PhyAddrPointer_reg[3]/NET0131  , \P3_PhyAddrPointer_reg[4]/NET0131  , \P3_PhyAddrPointer_reg[5]/NET0131  , \P3_PhyAddrPointer_reg[6]/NET0131  , \P3_PhyAddrPointer_reg[7]/NET0131  , \P3_PhyAddrPointer_reg[8]/NET0131  , \P3_PhyAddrPointer_reg[9]/NET0131  , \P3_ReadRequest_reg/NET0131  , \P3_RequestPending_reg/NET0131  , \P3_State2_reg[0]/NET0131  , \P3_State2_reg[1]/NET0131  , \P3_State2_reg[2]/NET0131  , \P3_State2_reg[3]/NET0131  , \P3_State_reg[0]/NET0131  , \P3_State_reg[1]/NET0131  , \P3_State_reg[2]/NET0131  , \P3_lWord_reg[0]/NET0131  , \P3_lWord_reg[10]/NET0131  , \P3_lWord_reg[11]/NET0131  , \P3_lWord_reg[12]/NET0131  , \P3_lWord_reg[13]/NET0131  , \P3_lWord_reg[14]/NET0131  , \P3_lWord_reg[15]/NET0131  , \P3_lWord_reg[1]/NET0131  , \P3_lWord_reg[2]/NET0131  , \P3_lWord_reg[3]/NET0131  , \P3_lWord_reg[4]/NET0131  , \P3_lWord_reg[5]/NET0131  , \P3_lWord_reg[6]/NET0131  , \P3_lWord_reg[7]/NET0131  , \P3_lWord_reg[8]/NET0131  , \P3_lWord_reg[9]/NET0131  , \P3_rEIP_reg[0]/NET0131  , \P3_rEIP_reg[10]/NET0131  , \P3_rEIP_reg[11]/NET0131  , \P3_rEIP_reg[12]/NET0131  , \P3_rEIP_reg[13]/NET0131  , \P3_rEIP_reg[14]/NET0131  , \P3_rEIP_reg[15]/NET0131  , \P3_rEIP_reg[16]/NET0131  , \P3_rEIP_reg[17]/NET0131  , \P3_rEIP_reg[18]/NET0131  , \P3_rEIP_reg[19]/NET0131  , \P3_rEIP_reg[1]/NET0131  , \P3_rEIP_reg[20]/NET0131  , \P3_rEIP_reg[21]/NET0131  , \P3_rEIP_reg[22]/NET0131  , \P3_rEIP_reg[23]/NET0131  , \P3_rEIP_reg[24]/NET0131  , \P3_rEIP_reg[25]/NET0131  , \P3_rEIP_reg[26]/NET0131  , \P3_rEIP_reg[27]/NET0131  , \P3_rEIP_reg[28]/NET0131  , \P3_rEIP_reg[29]/NET0131  , \P3_rEIP_reg[2]/NET0131  , \P3_rEIP_reg[30]/NET0131  , \P3_rEIP_reg[31]/NET0131  , \P3_rEIP_reg[3]/NET0131  , \P3_rEIP_reg[4]/NET0131  , \P3_rEIP_reg[5]/NET0131  , \P3_rEIP_reg[6]/NET0131  , \P3_rEIP_reg[7]/NET0131  , \P3_rEIP_reg[8]/NET0131  , \P3_rEIP_reg[9]/NET0131  , \P3_uWord_reg[0]/NET0131  , \P3_uWord_reg[10]/NET0131  , \P3_uWord_reg[11]/NET0131  , \P3_uWord_reg[12]/NET0131  , \P3_uWord_reg[13]/NET0131  , \P3_uWord_reg[14]/NET0131  , \P3_uWord_reg[1]/NET0131  , \P3_uWord_reg[2]/NET0131  , \P3_uWord_reg[3]/NET0131  , \P3_uWord_reg[4]/NET0131  , \P3_uWord_reg[5]/NET0131  , \P3_uWord_reg[6]/NET0131  , \P3_uWord_reg[7]/NET0131  , \P3_uWord_reg[8]/NET0131  , \P3_uWord_reg[9]/NET0131  , \address1[0]_pad  , \address1[10]_pad  , \address1[11]_pad  , \address1[12]_pad  , \address1[13]_pad  , \address1[14]_pad  , \address1[15]_pad  , \address1[16]_pad  , \address1[17]_pad  , \address1[18]_pad  , \address1[19]_pad  , \address1[1]_pad  , \address1[20]_pad  , \address1[21]_pad  , \address1[22]_pad  , \address1[23]_pad  , \address1[24]_pad  , \address1[25]_pad  , \address1[26]_pad  , \address1[27]_pad  , \address1[28]_pad  , \address1[29]_pad  , \address1[2]_pad  , \address1[3]_pad  , \address1[4]_pad  , \address1[5]_pad  , \address1[6]_pad  , \address1[7]_pad  , \address1[8]_pad  , \address1[9]_pad  , \ast1_pad  , \ast2_pad  , \bs16_pad  , \buf1_reg[0]/NET0131  , \buf1_reg[10]/NET0131  , \buf1_reg[11]/NET0131  , \buf1_reg[12]/NET0131  , \buf1_reg[13]/NET0131  , \buf1_reg[14]/NET0131  , \buf1_reg[15]/NET0131  , \buf1_reg[16]/NET0131  , \buf1_reg[17]/NET0131  , \buf1_reg[18]/NET0131  , \buf1_reg[19]/NET0131  , \buf1_reg[1]/NET0131  , \buf1_reg[20]/NET0131  , \buf1_reg[21]/NET0131  , \buf1_reg[22]/NET0131  , \buf1_reg[23]/NET0131  , \buf1_reg[24]/NET0131  , \buf1_reg[25]/NET0131  , \buf1_reg[26]/NET0131  , \buf1_reg[27]/NET0131  , \buf1_reg[28]/NET0131  , \buf1_reg[29]/NET0131  , \buf1_reg[2]/NET0131  , \buf1_reg[30]/NET0131  , \buf1_reg[3]/NET0131  , \buf1_reg[4]/NET0131  , \buf1_reg[5]/NET0131  , \buf1_reg[6]/NET0131  , \buf1_reg[7]/NET0131  , \buf1_reg[8]/NET0131  , \buf1_reg[9]/NET0131  , \buf2_reg[0]/NET0131  , \buf2_reg[10]/NET0131  , \buf2_reg[11]/NET0131  , \buf2_reg[12]/NET0131  , \buf2_reg[13]/NET0131  , \buf2_reg[14]/NET0131  , \buf2_reg[15]/NET0131  , \buf2_reg[16]/NET0131  , \buf2_reg[17]/NET0131  , \buf2_reg[18]/NET0131  , \buf2_reg[19]/NET0131  , \buf2_reg[1]/NET0131  , \buf2_reg[20]/NET0131  , \buf2_reg[21]/NET0131  , \buf2_reg[22]/NET0131  , \buf2_reg[23]/NET0131  , \buf2_reg[24]/NET0131  , \buf2_reg[25]/NET0131  , \buf2_reg[26]/NET0131  , \buf2_reg[27]/NET0131  , \buf2_reg[28]/NET0131  , \buf2_reg[29]/NET0131  , \buf2_reg[2]/NET0131  , \buf2_reg[30]/NET0131  , \buf2_reg[3]/NET0131  , \buf2_reg[4]/NET0131  , \buf2_reg[5]/NET0131  , \buf2_reg[6]/NET0131  , \buf2_reg[7]/NET0131  , \buf2_reg[8]/NET0131  , \buf2_reg[9]/NET0131  , \datai[0]_pad  , \datai[10]_pad  , \datai[11]_pad  , \datai[12]_pad  , \datai[13]_pad  , \datai[14]_pad  , \datai[15]_pad  , \datai[16]_pad  , \datai[17]_pad  , \datai[18]_pad  , \datai[19]_pad  , \datai[1]_pad  , \datai[20]_pad  , \datai[21]_pad  , \datai[22]_pad  , \datai[23]_pad  , \datai[24]_pad  , \datai[25]_pad  , \datai[26]_pad  , \datai[27]_pad  , \datai[28]_pad  , \datai[29]_pad  , \datai[2]_pad  , \datai[30]_pad  , \datai[31]_pad  , \datai[3]_pad  , \datai[4]_pad  , \datai[5]_pad  , \datai[6]_pad  , \datai[7]_pad  , \datai[8]_pad  , \datai[9]_pad  , \datao[0]_pad  , \datao[10]_pad  , \datao[11]_pad  , \datao[12]_pad  , \datao[13]_pad  , \datao[14]_pad  , \datao[15]_pad  , \datao[16]_pad  , \datao[17]_pad  , \datao[18]_pad  , \datao[19]_pad  , \datao[1]_pad  , \datao[20]_pad  , \datao[21]_pad  , \datao[22]_pad  , \datao[23]_pad  , \datao[24]_pad  , \datao[25]_pad  , \datao[26]_pad  , \datao[27]_pad  , \datao[28]_pad  , \datao[29]_pad  , \datao[2]_pad  , \datao[30]_pad  , \datao[3]_pad  , \datao[4]_pad  , \datao[5]_pad  , \datao[6]_pad  , \datao[7]_pad  , \datao[8]_pad  , \datao[9]_pad  , dc_pad , hold_pad , mio_pad , na_pad , \ready11_reg/NET0131  , \ready12_reg/NET0131  , \ready1_pad  , \ready21_reg/NET0131  , \ready22_reg/NET0131  , \ready2_pad  , wr_pad , \_al_n0  , \_al_n1  , \address2[0]_pad  , \address2[10]_pad  , \address2[11]_pad  , \address2[12]_pad  , \address2[13]_pad  , \address2[14]_pad  , \address2[15]_pad  , \address2[16]_pad  , \address2[17]_pad  , \address2[18]_pad  , \address2[19]_pad  , \address2[1]_pad  , \address2[20]_pad  , \address2[21]_pad  , \address2[22]_pad  , \address2[23]_pad  , \address2[24]_pad  , \address2[25]_pad  , \address2[26]_pad  , \address2[27]_pad  , \address2[28]_pad  , \address2[29]_pad  , \address2[2]_pad  , \address2[3]_pad  , \address2[4]_pad  , \address2[5]_pad  , \address2[6]_pad  , \address2[7]_pad  , \address2[8]_pad  , \address2[9]_pad  , \g133468/_2_  , \g133469/_2_  , \g133470/_2_  , \g133475/_0_  , \g133476/_2_  , \g133515/_0_  , \g133516/_0_  , \g133517/_0_  , \g133518/_0_  , \g133523/_0_  , \g133524/_0_  , \g133528/_0_  , \g133529/_0_  , \g133531/_0_  , \g133532/_0_  , \g133533/_0_  , \g133534/_0_  , \g133535/_0_  , \g133536/_0_  , \g133537/_0_  , \g133538/_0_  , \g133539/_0_  , \g133540/_0_  , \g133541/_0_  , \g133542/_0_  , \g133543/_0_  , \g133544/_0_  , \g133545/_0_  , \g133546/_0_  , \g133547/_0_  , \g133548/_0_  , \g133549/_0_  , \g133550/_0_  , \g133551/_0_  , \g133552/_0_  , \g133553/_0_  , \g133554/_0_  , \g133555/_0_  , \g133556/_0_  , \g133557/_0_  , \g133558/_0_  , \g133559/_0_  , \g133560/_0_  , \g133561/_0_  , \g133566/_0_  , \g133619/_0_  , \g133659/_0_  , \g133660/_0_  , \g133662/_0_  , \g133663/_0_  , \g133664/_0_  , \g133665/_0_  , \g133666/_0_  , \g133667/_0_  , \g133668/_0_  , \g133669/_0_  , \g133670/_0_  , \g133671/_0_  , \g133672/_0_  , \g133673/_0_  , \g133674/_0_  , \g133675/_0_  , \g133676/_0_  , \g133677/_0_  , \g133678/_0_  , \g133679/_0_  , \g133680/_0_  , \g133681/_0_  , \g133682/_0_  , \g133683/_0_  , \g133684/_0_  , \g133685/_0_  , \g133686/_0_  , \g133687/_0_  , \g133688/_0_  , \g133689/_0_  , \g133690/_0_  , \g133691/_0_  , \g133694/_0_  , \g133697/_0_  , \g133702/_0_  , \g133703/_0_  , \g133756/_0_  , \g133792/_0_  , \g133793/_0_  , \g133794/_0_  , \g133796/_0_  , \g133797/_0_  , \g133798/_0_  , \g133799/_0_  , \g133800/_0_  , \g133801/_0_  , \g133802/_0_  , \g133803/_0_  , \g133804/_0_  , \g133806/_0_  , \g133807/_0_  , \g133808/_0_  , \g133812/_0_  , \g133813/_0_  , \g133814/_0_  , \g133817/_0_  , \g133821/_0_  , \g133824/_0_  , \g133826/_0_  , \g133828/_0_  , \g133864/_0_  , \g133865/_0_  , \g133867/_0_  , \g133868/_0_  , \g133869/_0_  , \g133871/_0_  , \g133872/_0_  , \g133873/_0_  , \g133874/_0_  , \g133875/_0_  , \g133876/_0_  , \g133877/_0_  , \g133878/_0_  , \g133879/_0_  , \g133881/_0_  , \g133882/_0_  , \g133883/_0_  , \g133884/_0_  , \g133885/_0_  , \g133886/_0_  , \g133887/_0_  , \g133888/_0_  , \g133889/_0_  , \g133890/_0_  , \g133891/_0_  , \g133892/_0_  , \g133893/_0_  , \g133894/_0_  , \g133895/_0_  , \g133896/_0_  , \g133897/_0_  , \g133898/_0_  , \g133910/_0_  , \g133911/_0_  , \g133912/_0_  , \g133915/_0_  , \g133917/_0_  , \g133929/_0_  , \g134014/_0_  , \g134040/_0_  , \g134041/_0_  , \g134042/_0_  , \g134043/_0_  , \g134044/_0_  , \g134045/_0_  , \g134046/_0_  , \g134047/_0_  , \g134048/_0_  , \g134049/_0_  , \g134050/_0_  , \g134051/_0_  , \g134052/_0_  , \g134053/_0_  , \g134054/_0_  , \g134056/_0_  , \g134059/_0_  , \g134064/_0_  , \g134067/_0_  , \g134068/_0_  , \g134069/_0_  , \g134070/_0_  , \g134071/_0_  , \g134073/_0_  , \g134076/_0_  , \g134131/_0_  , \g134132/_0_  , \g134156/_0_  , \g134157/_0_  , \g134158/_0_  , \g134159/_0_  , \g134163/_0_  , \g134164/_0_  , \g134165/_0_  , \g134166/_0_  , \g134167/_0_  , \g134168/_0_  , \g134169/_0_  , \g134170/_0_  , \g134171/_0_  , \g134172/_0_  , \g134173/_0_  , \g134174/_0_  , \g134176/_0_  , \g134177/_0_  , \g134178/_0_  , \g134179/_0_  , \g134181/_0_  , \g134183/_0_  , \g134184/_0_  , \g134185/_0_  , \g134186/_0_  , \g134187/_0_  , \g134188/_0_  , \g134189/_0_  , \g134190/_0_  , \g134191/_0_  , \g134194/_0_  , \g134202/_0_  , \g134207/_0_  , \g134214/_0_  , \g134216/_0_  , \g134226/_0_  , \g134228/_0_  , \g134360/_0_  , \g134383/_0_  , \g134412/_0_  , \g134413/_0_  , \g134419/_0_  , \g134420/_0_  , \g134421/_0_  , \g134422/_0_  , \g134423/_0_  , \g134424/_0_  , \g134426/_0_  , \g134429/_0_  , \g134431/_0_  , \g134433/_0_  , \g134434/_0_  , \g134435/_0_  , \g134436/_0_  , \g134438/_0_  , \g134439/_0_  , \g134441/_0_  , \g134442/_0_  , \g134443/_0_  , \g134445/_0_  , \g134446/_0_  , \g134447/_0_  , \g134448/_0_  , \g134449/_0_  , \g134450/_0_  , \g134451/_0_  , \g134453/_0_  , \g134454/_0_  , \g134455/_0_  , \g134457/_0_  , \g134458/_0_  , \g134459/_0_  , \g134460/_0_  , \g134469/_0_  , \g134470/_0_  , \g134471/_0_  , \g134472/_0_  , \g134479/_0_  , \g134480/_0_  , \g134481/_0_  , \g134482/_0_  , \g134490/_0_  , \g134491/_0_  , \g134496/_0_  , \g134506/_0_  , \g134508/_0_  , \g134579/_0_  , \g134603/_0_  , \g134604/_0_  , \g134605/_0_  , \g134606/_0_  , \g134607/_0_  , \g134608/_0_  , \g134609/_0_  , \g134610/_0_  , \g134611/_0_  , \g134612/_0_  , \g134613/_0_  , \g134614/_0_  , \g134615/_0_  , \g134616/_0_  , \g134617/_0_  , \g134618/_0_  , \g134619/_0_  , \g134620/_0_  , \g134621/_0_  , \g134632/_0_  , \g134633/_0_  , \g134636/_0_  , \g134637/_0_  , \g134638/_0_  , \g134639/_0_  , \g134645/_0_  , \g134646/_0_  , \g134648/_0_  , \g134649/_0_  , \g134650/_0_  , \g134651/_0_  , \g134652/_0_  , \g134656/_0_  , \g134657/_0_  , \g134658/_0_  , \g134664/_0_  , \g134665/_0_  , \g134671/_0_  , \g134672/_0_  , \g134686/_0_  , \g134687/_0_  , \g134735/_0_  , \g134908/_0_  , \g134909/_0_  , \g134910/_0_  , \g134920/_0_  , \g134921/_0_  , \g134922/_0_  , \g134923/_0_  , \g134925/_0_  , \g134926/_0_  , \g134928/_0_  , \g134929/_0_  , \g134933/_0_  , \g134934/_0_  , \g134935/_0_  , \g134936/_0_  , \g134937/_0_  , \g134938/_0_  , \g134940/_0_  , \g134941/_0_  , \g134943/_0_  , \g134945/_0_  , \g134946/_0_  , \g134947/_0_  , \g134948/_0_  , \g134949/_0_  , \g134950/_0_  , \g134959/_0_  , \g134960/_0_  , \g134961/_0_  , \g134979/_0_  , \g134980/_0_  , \g135054/_0_  , \g135061/_0_  , \g135072/_0_  , \g135100/_0_  , \g135127/_0_  , \g135128/_0_  , \g135129/_0_  , \g135130/_0_  , \g135132/_0_  , \g135133/_0_  , \g135134/_0_  , \g135135/_0_  , \g135136/_0_  , \g135137/_0_  , \g135138/_0_  , \g135139/_0_  , \g135140/_0_  , \g135141/_0_  , \g135142/_0_  , \g135145/_0_  , \g135146/_0_  , \g135151/_0_  , \g135154/_0_  , \g135155/_0_  , \g135158/_0_  , \g135163/_0_  , \g135164/_0_  , \g135165/_0_  , \g135192/_0_  , \g135197/_0_  , \g135217/_0_  , \g135225/_0_  , \g135231/_0_  , \g135272/_0_  , \g135290/_0_  , \g135291/_0_  , \g135293/_0_  , \g135294/_0_  , \g135295/_0_  , \g135296/_0_  , \g135297/_0_  , \g135412/_0_  , \g135437/_0_  , \g135438/_0_  , \g135443/_0_  , \g135444/_0_  , \g135445/_0_  , \g135446/_0_  , \g135447/_0_  , \g135448/_0_  , \g135449/_0_  , \g135450/_0_  , \g135451/_0_  , \g135452/_0_  , \g135454/_0_  , \g135455/_0_  , \g135456/_0_  , \g135457/_0_  , \g135458/_0_  , \g135463/_0_  , \g135466/_0_  , \g135473/_0_  , \g135481/_0_  , \g135497/_0_  , \g135503/_0_  , \g135505/_0_  , \g135506/_0_  , \g135557/_0_  , \g135558/_0_  , \g135569/_0_  , \g135570/_0_  , \g135571/_0_  , \g135572/_0_  , \g135573/_0_  , \g135575/_0_  , \g135578/_0_  , \g135754/_0_  , \g135755/_0_  , \g135756/_0_  , \g135767/_0_  , \g135768/_0_  , \g135769/_0_  , \g135777/_0_  , \g135778/_0_  , \g135779/_0_  , \g135872/_0_  , \g135873/_0_  , \g135875/_0_  , \g135877/_0_  , \g135878/_0_  , \g135879/_0_  , \g135880/_0_  , \g136087/_0_  , \g136118/_0_  , \g136119/_0_  , \g136120/_0_  , \g136121/_0_  , \g136122/_0_  , \g136123/_0_  , \g136124/_0_  , \g136125/_0_  , \g136126/_0_  , \g136127/_0_  , \g136128/_0_  , \g136129/_0_  , \g136130/_0_  , \g136131/_0_  , \g136132/_0_  , \g136133/_0_  , \g136172/_0_  , \g136173/_0_  , \g136174/_0_  , \g136175/_0_  , \g136177/_0_  , \g136178/_0_  , \g136242/_0_  , \g136243/_0_  , \g136244/_0_  , \g136246/_0_  , \g136248/_0_  , \g136249/_0_  , \g136250/_0_  , \g136251/_0_  , \g136252/_0_  , \g136253/_0_  , \g136254/_0_  , \g136255/_0_  , \g136256/_0_  , \g136257/_0_  , \g136258/_0_  , \g136259/_0_  , \g136260/_0_  , \g136261/_0_  , \g136262/_0_  , \g136263/_0_  , \g136264/_0_  , \g136265/_0_  , \g136266/_0_  , \g136267/_0_  , \g136268/_0_  , \g136269/_0_  , \g136270/_0_  , \g136271/_0_  , \g136272/_0_  , \g136273/_0_  , \g136274/_0_  , \g136275/_0_  , \g136276/_0_  , \g136277/_0_  , \g136279/_0_  , \g136280/_0_  , \g136281/_0_  , \g136282/_0_  , \g136283/_0_  , \g136285/_0_  , \g136286/_0_  , \g136287/_0_  , \g136288/_0_  , \g136289/_0_  , \g136290/_0_  , \g136291/_0_  , \g136292/_0_  , \g136293/_0_  , \g136295/_0_  , \g136467/_0_  , \g136468/_0_  , \g136469/_0_  , \g136470/_0_  , \g136472/_0_  , \g136473/_0_  , \g136474/_0_  , \g136476/_0_  , \g136479/_0_  , \g136480/_0_  , \g136481/_0_  , \g136482/_0_  , \g136483/_0_  , \g136484/_0_  , \g136485/_0_  , \g136486/_0_  , \g136528/_0_  , \g136529/_0_  , \g136530/_0_  , \g136531/_0_  , \g136532/_0_  , \g136533/_0_  , \g136534/_0_  , \g136535/_0_  , \g136536/_0_  , \g136537/_0_  , \g136538/_0_  , \g136539/_0_  , \g136540/_0_  , \g136541/_0_  , \g136542/_0_  , \g136543/_0_  , \g136544/_0_  , \g136545/_0_  , \g136546/_0_  , \g136547/_0_  , \g136548/_0_  , \g136549/_0_  , \g136550/_0_  , \g136551/_0_  , \g136552/_0_  , \g136553/_0_  , \g136554/_0_  , \g136555/_0_  , \g136556/_0_  , \g136557/_0_  , \g136558/_0_  , \g136559/_0_  , \g136560/_0_  , \g136561/_0_  , \g136562/_0_  , \g136563/_0_  , \g136564/_0_  , \g136565/_0_  , \g136566/_0_  , \g136567/_0_  , \g136568/_0_  , \g136570/_0_  , \g136571/_0_  , \g136572/_0_  , \g136573/_0_  , \g136574/_0_  , \g136575/_0_  , \g136576/_0_  , \g136577/_0_  , \g136578/_0_  , \g136579/_0_  , \g136580/_0_  , \g136582/_0_  , \g136583/_0_  , \g136584/_0_  , \g136585/_0_  , \g136586/_0_  , \g136587/_0_  , \g136588/_0_  , \g136589/_0_  , \g136590/_0_  , \g136591/_0_  , \g136592/_0_  , \g136593/_0_  , \g136594/_0_  , \g136595/_0_  , \g136596/_0_  , \g136597/_0_  , \g136598/_0_  , \g136599/_0_  , \g136600/_0_  , \g136601/_0_  , \g136602/_0_  , \g136603/_0_  , \g136604/_0_  , \g136605/_0_  , \g136606/_0_  , \g136607/_0_  , \g136609/_0_  , \g136610/_0_  , \g136611/_0_  , \g136616/_0_  , \g136617/_0_  , \g136618/_0_  , \g136619/_0_  , \g136626/_0_  , \g136628/_0_  , \g136646/_0_  , \g136649/_0_  , \g136662/_0_  , \g136666/_0_  , \g136695/_0_  , \g136696/_0_  , \g136699/_0_  , \g136762/_0_  , \g136763/_0_  , \g136764/_0_  , \g136765/_0_  , \g136768/_0_  , \g136769/_0_  , \g137051/_0_  , \g137052/_0_  , \g137053/_0_  , \g137054/_0_  , \g137055/_0_  , \g137056/_0_  , \g137057/_0_  , \g137060/_0_  , \g137061/_0_  , \g137063/_0_  , \g137064/_0_  , \g137065/_0_  , \g137067/_0_  , \g137069/_0_  , \g137072/_0_  , \g137073/_0_  , \g137075/_0_  , \g137111/_0_  , \g137122/_0_  , \g137133/_0_  , \g137134/_0_  , \g137135/_0_  , \g137136/_0_  , \g137137/_0_  , \g137138/_0_  , \g137144/_0_  , \g137145/_0_  , \g137146/_0_  , \g137149/_0_  , \g137234/_0_  , \g137237/_0_  , \g137238/_0_  , \g137294/_0_  , \g137295/_0_  , \g137296/_0_  , \g137297/_0_  , \g137298/_0_  , \g137299/_0_  , \g137300/_0_  , \g137301/_0_  , \g137302/_0_  , \g137303/_0_  , \g137304/_0_  , \g137305/_0_  , \g137306/_0_  , \g137307/_0_  , \g137308/_0_  , \g137309/_0_  , \g137310/_0_  , \g137311/_0_  , \g137312/_0_  , \g137313/_0_  , \g137314/_0_  , \g137315/_0_  , \g137316/_0_  , \g137317/_0_  , \g137318/_0_  , \g137319/_0_  , \g137320/_0_  , \g137321/_0_  , \g137322/_0_  , \g137323/_0_  , \g137324/_0_  , \g137325/_0_  , \g137327/_0_  , \g137328/_0_  , \g137329/_0_  , \g137330/_0_  , \g137331/_0_  , \g137332/_0_  , \g137333/_0_  , \g137334/_0_  , \g137335/_0_  , \g137336/_0_  , \g137337/_0_  , \g137338/_0_  , \g137339/_0_  , \g137340/_0_  , \g137341/_0_  , \g137342/_0_  , \g137343/_0_  , \g137344/_0_  , \g137345/_0_  , \g137346/_0_  , \g137347/_0_  , \g137349/_0_  , \g137350/_0_  , \g137351/_0_  , \g137352/_0_  , \g137353/_0_  , \g137354/_0_  , \g137448/_0_  , \g137483/_0_  , \g137484/_0_  , \g137485/_0_  , \g137486/_0_  , \g137487/_0_  , \g137488/_0_  , \g137491/_0_  , \g137492/_0_  , \g137493/_0_  , \g137494/_0_  , \g137495/_0_  , \g137496/_0_  , \g137497/_0_  , \g137499/_0_  , \g137501/_0_  , \g137502/_0_  , \g137503/_0_  , \g137504/_0_  , \g137505/_0_  , \g137506/_0_  , \g137507/_0_  , \g137508/_0_  , \g137509/_0_  , \g137511/_0_  , \g137512/_0_  , \g137513/_0_  , \g137514/_0_  , \g137515/_0_  , \g137516/_0_  , \g137517/_0_  , \g137519/_0_  , \g137520/_0_  , \g137521/_0_  , \g137524/_0_  , \g137541/_0_  , \g137547/_0_  , \g137554/_0_  , \g137559/_0_  , \g137566/_0_  , \g137571/_0_  , \g137778/_0_  , \g137782/_0_  , \g137783/_0_  , \g137784/_0_  , \g137785/_0_  , \g137786/_0_  , \g137820/_0_  , \g137821/_0_  , \g137822/_0_  , \g137823/_0_  , \g137824/_0_  , \g137825/_0_  , \g137826/_0_  , \g137827/_0_  , \g137828/_0_  , \g137829/_0_  , \g137830/_0_  , \g137831/_0_  , \g137832/_0_  , \g137833/_0_  , \g137834/_0_  , \g137835/_0_  , \g137836/_0_  , \g137837/_0_  , \g137838/_0_  , \g137839/_0_  , \g137840/_0_  , \g137841/_0_  , \g137842/_0_  , \g137843/_0_  , \g137844/_0_  , \g137845/_0_  , \g137846/_0_  , \g137847/_0_  , \g137848/_0_  , \g137849/_0_  , \g137850/_0_  , \g137851/_0_  , \g137852/_0_  , \g137853/_0_  , \g137854/_0_  , \g137855/_0_  , \g137856/_0_  , \g137857/_0_  , \g137858/_0_  , \g137859/_0_  , \g137860/_0_  , \g137861/_0_  , \g137862/_0_  , \g137863/_0_  , \g137864/_0_  , \g137865/_0_  , \g137866/_0_  , \g137867/_0_  , \g137868/_0_  , \g137869/_0_  , \g137870/_0_  , \g137871/_0_  , \g137872/_0_  , \g137873/_0_  , \g137874/_0_  , \g137875/_0_  , \g137876/_0_  , \g137877/_0_  , \g137878/_0_  , \g137879/_0_  , \g137880/_0_  , \g137881/_0_  , \g137882/_0_  , \g137883/_0_  , \g137884/_0_  , \g137885/_0_  , \g137886/_0_  , \g137887/_0_  , \g137888/_0_  , \g137889/_0_  , \g137890/_0_  , \g137891/_0_  , \g137892/_0_  , \g137893/_0_  , \g137894/_0_  , \g137895/_0_  , \g137896/_0_  , \g137897/_0_  , \g137898/_0_  , \g137899/_0_  , \g137900/_0_  , \g137901/_0_  , \g137902/_0_  , \g137903/_0_  , \g138338/_0_  , \g138340/_0_  , \g138341/_0_  , \g138346/_0_  , \g138347/_0_  , \g138375/_0_  , \g138395/_0_  , \g138396/_0_  , \g138397/_0_  , \g138398/_0_  , \g138400/_0_  , \g138401/_0_  , \g138402/_0_  , \g138403/_0_  , \g138404/_0_  , \g138405/_0_  , \g138406/_0_  , \g138407/_0_  , \g138408/_0_  , \g138409/_0_  , \g138410/_0_  , \g138411/_0_  , \g138412/_0_  , \g138419/_0_  , \g138420/_0_  , \g138421/_0_  , \g138422/_0_  , \g138423/_0_  , \g138424/_0_  , \g138425/_0_  , \g138426/_0_  , \g138427/_0_  , \g138428/_0_  , \g138429/_0_  , \g138430/_0_  , \g138431/_0_  , \g138432/_0_  , \g138433/_0_  , \g138434/_0_  , \g138435/_0_  , \g138436/_0_  , \g138437/_0_  , \g138438/_0_  , \g138439/_0_  , \g138440/_0_  , \g138441/_0_  , \g138442/_0_  , \g138443/_0_  , \g138908/_0_  , \g138909/_0_  , \g138910/_0_  , \g138914/_0_  , \g138915/_0_  , \g138917/_0_  , \g138918/_0_  , \g138919/_0_  , \g138920/_0_  , \g138921/_0_  , \g138925/_0_  , \g138926/_0_  , \g138927/_0_  , \g138930/_0_  , \g138931/_0_  , \g138932/_0_  , \g138960/_0_  , \g138962/_0_  , \g139037/_0_  , \g139038/_0_  , \g139040/_0_  , \g139043/_0_  , \g139044/_0_  , \g139045/_0_  , \g139046/_0_  , \g139047/_0_  , \g139048/_0_  , \g139049/_0_  , \g139050/_0_  , \g139051/_0_  , \g139053/_0_  , \g139054/_0_  , \g139055/_0_  , \g139056/_0_  , \g139057/_0_  , \g139058/_0_  , \g139059/_0_  , \g139060/_0_  , \g139062/_0_  , \g139063/_0_  , \g139064/_0_  , \g139099/_0_  , \g139126/_0_  , \g139127/_0_  , \g139128/_0_  , \g139129/_0_  , \g139130/_0_  , \g139131/_0_  , \g139132/_0_  , \g139133/_0_  , \g139134/_0_  , \g139135/_0_  , \g139136/_0_  , \g139137/_0_  , \g139138/_0_  , \g139139/_0_  , \g139140/_0_  , \g139141/_0_  , \g139260/_0_  , \g139263/_0_  , \g139267/_0_  , \g139270/_0_  , \g139273/_0_  , \g139276/_0_  , \g139279/_0_  , \g139283/_0_  , \g139286/_0_  , \g139289/_0_  , \g139292/_0_  , \g139295/_0_  , \g139298/_0_  , \g139302/_0_  , \g139305/_0_  , \g139309/_0_  , \g139871/_0_  , \g139872/_0_  , \g139873/_0_  , \g139874/_0_  , \g139875/_0_  , \g139876/_0_  , \g139877/_0_  , \g139878/_0_  , \g139879/_0_  , \g139880/_0_  , \g139881/_0_  , \g139882/_0_  , \g139883/_0_  , \g139884/_0_  , \g139885/_0_  , \g139886/_0_  , \g139887/_0_  , \g139888/_0_  , \g139889/_0_  , \g139890/_0_  , \g139891/_0_  , \g139892/_0_  , \g139893/_0_  , \g139895/_0_  , \g139896/_0_  , \g139899/_0_  , \g139901/_0_  , \g139902/_0_  , \g139903/_0_  , \g139904/_0_  , \g140285/_0_  , \g140288/_0_  , \g140329/_0_  , \g140774/_0_  , \g140832/_0_  , \g140834/_0_  , \g140836/_0_  , \g140838/_0_  , \g140840/_0_  , \g140842/_0_  , \g140844/_0_  , \g140846/_0_  , \g140847/_0_  , \g140848/_0_  , \g140850/_0_  , \g140851/_0_  , \g140852/_0_  , \g140853/_0_  , \g140855/_0_  , \g140857/_0_  , \g140861/_0_  , \g140923/_0_  , \g141178/_0_  , \g141179/_0_  , \g141180/_0_  , \g141480/_0_  , \g141495/_0_  , \g141497/_0_  , \g141562/_0_  , \g141563/_0_  , \g141564/_0_  , \g141589/_0_  , \g141617/_0_  , \g141618/_0_  , \g141621/_0_  , \g141625/_0_  , \g141626/_0_  , \g141630/_0_  , \g141634/_0_  , \g141638/_0_  , \g141642/_0_  , \g141646/_0_  , \g141649/_0_  , \g141651/_0_  , \g141652/_0_  , \g141655/_0_  , \g141658/_0_  , \g141661/_0_  , \g141663/_0_  , \g141664/_0_  , \g141667/_0_  , \g141671/_0_  , \g141706/_0_  , \g141976/_0_  , \g141977/_0_  , \g141994/_0_  , \g142246/_0_  , \g142247/_0_  , \g142253/_0_  , \g142689/_0_  , \g142693/_0_  , \g142701/_0_  , \g142704/_0_  , \g142707/_0_  , \g142710/_0_  , \g142713/_0_  , \g142714/_0_  , \g142717/_0_  , \g142720/_0_  , \g142723/_0_  , \g142727/_0_  , \g142734/_0_  , \g143080/_0_  , \g143081/_0_  , \g143083/_0_  , \g143149/_0_  , \g143150/_0_  , \g143153/_0_  , \g143752/_0_  , \g143753/_0_  , \g143759/_0_  , \g144242/_0_  , \g144243/_0_  , \g144244/_0_  , \g144245/_0_  , \g144246/_0_  , \g144249/_0_  , \g145699/_0_  , \g145700/_0_  , \g145702/_0_  , \g145756/_0_  , \g145757/_0_  , \g145758/_0_  , \g146850/_0_  , \g146851/_0_  , \g146864/_0_  , \g147277/_0_  , \g147278/_0_  , \g147279/_0_  , \g147304/_0_  , \g147305/_0_  , \g147306/_0_  , \g147338/_3_  , \g147339/_3_  , \g147340/_3_  , \g147341/_3_  , \g147342/_3_  , \g147343/_3_  , \g147344/_3_  , \g147345/_3_  , \g147346/_3_  , \g147347/_3_  , \g147348/_3_  , \g147349/_3_  , \g147350/_3_  , \g147351/_3_  , \g147352/_3_  , \g147353/_3_  , \g147354/_3_  , \g147355/_3_  , \g147356/_3_  , \g147357/_3_  , \g147358/_3_  , \g147359/_3_  , \g147360/_3_  , \g147362/_3_  , \g147363/_3_  , \g147364/_3_  , \g147365/_3_  , \g147366/_3_  , \g147367/_3_  , \g147368/_3_  , \g147369/_3_  , \g148630/_0_  , \g148631/_0_  , \g148676/_0_  , \g148785/_0_  , \g148788/_0_  , \g148789/_0_  , \g148834/_0_  , \g148836/_0_  , \g148838/_0_  , \g149836/_0_  , \g149837/_0_  , \g149838/_0_  , \g150142/_0_  , \g152366/_0_  , \g152367/_0_  , \g152368/_0_  , \g152426/_0_  , \g152427/_0_  , \g152428/_0_  , \g152586/_0_  , \g152587/_0_  , \g152588/_0_  , \g153217/_0_  , \g154117/_0_  , \g154118/_0_  , \g154130/_0_  , \g154269/_0_  , \g154270/_0_  , \g154284/_0_  , \g154682/_0_  , \g155004/_0_  , \g155020/_0_  , \g155121/_0_  , \g155124/_0_  , \g155126/_0_  , \g155228/_0_  , \g155229/_0_  , \g155230/_0_  , \g155326/_0_  , \g155327/_0_  , \g155330/_0_  , \g155353/_0_  , \g155354/_0_  , \g155356/_0_  , \g155602/_0_  , \g155633/_0_  , \g155634/_0_  , \g155699/_0_  , \g155708/_0_  , \g155715/_0_  , \g156008/_0_  , \g156013/_0_  , \g156019/_0_  , \g156352/_0_  , \g156353/_0_  , \g156356/_0_  , \g156359/_0_  , \g156360/_0_  , \g156361/_0_  , \g156464/_0_  , \g156465/_0_  , \g156469/_0_  , \g156777/_0_  , \g156778/_0_  , \g156789/_0_  , \g158956/_0_  , \g158957/_0_  , \g158966/_0_  , \g159429/_1_  , \g159477/_1_  , \g159500/_1_  , \g159681/_0_  , \g159890/_0_  , \g159950/_0_  , \g160246/_0_  , \g160846/_0_  , \g160860/_0_  , \g160961/_0_  , \g160987/_0_  , \g161000/_0_  , \g161005/_0_  , \g161042/_0_  , \g161119/_0_  , \g161143/_0_  , \g161150/_0_  , \g161172/_0_  , \g161207/_0_  , \g161315/_0_  , \g161332/_0_  , \g161421/_0_  , \g161492/_0_  , \g161541/_0_  , \g161623/_0_  , \g161655/_0_  , \g161678/_0_  , \g161709/_0_  , \g161737/_0_  , \g161751/_0_  , \g161756/_0_  , \g162016/_0_  , \g162020/_0_  , \g162024/_0_  , \g163326/_0_  , \g163326/_3_  , \g174072/_1_  , \g174360/_1_  , \g174391/_0_  , \g180307/_0_  , \g180335/_0_  , \g180369/_0_  , \g180385/_0_  , \g180395/_0_  , \g180442/_0_  , \g180453/_0_  , \g180524/_0_  , \g180586/_0_  , \g180596/_0_  , \g180606/_0_  , \g180654/_0_  , \g180715/_0_  , \g180805/_0_  , \g180836/_0_  , \g180929/_0_  , \g180944/_0_  , \g180975/_0_  , \g181036/_0_  , \g181072/_0_  , \g181083/_0_  , \g181093/_0_  , \g181127/_0_  , \g181137/_0_  , \g181150/_0_  , \g181160/_0_  , \g181180/_0_  , \g181191/_0_  , \g181238/_0_  , \g181262/_0_  , \g181270/_0_  , \g181280/_0_  , \g181315/_0_  , \g181366/_0_  , \g181385/_0_  , \g181458/_0_  , \g181464/_0_  , \g181478/_0_  , \g181522/_0_  , \g181537/_0_  , \g181584/_0_  , \g181669/_0_  , \g181681/_0_  , \g181719/_0_  , \g181778/_0_  , \g181840/_0_  , \g181936/_0_  , \g181986/_0_  , \g182000/_0_  , \g182083/_0_  , \g182179/_0_  , \g182201/_0_  , \g182227/_0_  , \g182316/_0_  , \g182358/_0_  , \g182473/_0_  , \g182678/_0_  , \g53/_0_  );
  input \P1_BE_n_reg[0]/NET0131  ;
  input \P1_BE_n_reg[1]/NET0131  ;
  input \P1_BE_n_reg[2]/NET0131  ;
  input \P1_BE_n_reg[3]/NET0131  ;
  input \P1_ByteEnable_reg[0]/NET0131  ;
  input \P1_ByteEnable_reg[1]/NET0131  ;
  input \P1_ByteEnable_reg[2]/NET0131  ;
  input \P1_ByteEnable_reg[3]/NET0131  ;
  input \P1_CodeFetch_reg/NET0131  ;
  input \P1_D_C_n_reg/NET0131  ;
  input \P1_DataWidth_reg[0]/NET0131  ;
  input \P1_DataWidth_reg[1]/NET0131  ;
  input \P1_Datao_reg[0]/NET0131  ;
  input \P1_Datao_reg[10]/NET0131  ;
  input \P1_Datao_reg[11]/NET0131  ;
  input \P1_Datao_reg[12]/NET0131  ;
  input \P1_Datao_reg[13]/NET0131  ;
  input \P1_Datao_reg[14]/NET0131  ;
  input \P1_Datao_reg[15]/NET0131  ;
  input \P1_Datao_reg[16]/NET0131  ;
  input \P1_Datao_reg[17]/NET0131  ;
  input \P1_Datao_reg[18]/NET0131  ;
  input \P1_Datao_reg[19]/NET0131  ;
  input \P1_Datao_reg[1]/NET0131  ;
  input \P1_Datao_reg[20]/NET0131  ;
  input \P1_Datao_reg[21]/NET0131  ;
  input \P1_Datao_reg[22]/NET0131  ;
  input \P1_Datao_reg[23]/NET0131  ;
  input \P1_Datao_reg[24]/NET0131  ;
  input \P1_Datao_reg[25]/NET0131  ;
  input \P1_Datao_reg[26]/NET0131  ;
  input \P1_Datao_reg[27]/NET0131  ;
  input \P1_Datao_reg[28]/NET0131  ;
  input \P1_Datao_reg[29]/NET0131  ;
  input \P1_Datao_reg[2]/NET0131  ;
  input \P1_Datao_reg[30]/NET0131  ;
  input \P1_Datao_reg[3]/NET0131  ;
  input \P1_Datao_reg[4]/NET0131  ;
  input \P1_Datao_reg[5]/NET0131  ;
  input \P1_Datao_reg[6]/NET0131  ;
  input \P1_Datao_reg[7]/NET0131  ;
  input \P1_Datao_reg[8]/NET0131  ;
  input \P1_Datao_reg[9]/NET0131  ;
  input \P1_EAX_reg[0]/NET0131  ;
  input \P1_EAX_reg[10]/NET0131  ;
  input \P1_EAX_reg[11]/NET0131  ;
  input \P1_EAX_reg[12]/NET0131  ;
  input \P1_EAX_reg[13]/NET0131  ;
  input \P1_EAX_reg[14]/NET0131  ;
  input \P1_EAX_reg[15]/NET0131  ;
  input \P1_EAX_reg[16]/NET0131  ;
  input \P1_EAX_reg[17]/NET0131  ;
  input \P1_EAX_reg[18]/NET0131  ;
  input \P1_EAX_reg[19]/NET0131  ;
  input \P1_EAX_reg[1]/NET0131  ;
  input \P1_EAX_reg[20]/NET0131  ;
  input \P1_EAX_reg[21]/NET0131  ;
  input \P1_EAX_reg[22]/NET0131  ;
  input \P1_EAX_reg[23]/NET0131  ;
  input \P1_EAX_reg[24]/NET0131  ;
  input \P1_EAX_reg[25]/NET0131  ;
  input \P1_EAX_reg[26]/NET0131  ;
  input \P1_EAX_reg[27]/NET0131  ;
  input \P1_EAX_reg[28]/NET0131  ;
  input \P1_EAX_reg[29]/NET0131  ;
  input \P1_EAX_reg[2]/NET0131  ;
  input \P1_EAX_reg[30]/NET0131  ;
  input \P1_EAX_reg[31]/NET0131  ;
  input \P1_EAX_reg[3]/NET0131  ;
  input \P1_EAX_reg[4]/NET0131  ;
  input \P1_EAX_reg[5]/NET0131  ;
  input \P1_EAX_reg[6]/NET0131  ;
  input \P1_EAX_reg[7]/NET0131  ;
  input \P1_EAX_reg[8]/NET0131  ;
  input \P1_EAX_reg[9]/NET0131  ;
  input \P1_EBX_reg[0]/NET0131  ;
  input \P1_EBX_reg[10]/NET0131  ;
  input \P1_EBX_reg[11]/NET0131  ;
  input \P1_EBX_reg[12]/NET0131  ;
  input \P1_EBX_reg[13]/NET0131  ;
  input \P1_EBX_reg[14]/NET0131  ;
  input \P1_EBX_reg[15]/NET0131  ;
  input \P1_EBX_reg[16]/NET0131  ;
  input \P1_EBX_reg[17]/NET0131  ;
  input \P1_EBX_reg[18]/NET0131  ;
  input \P1_EBX_reg[19]/NET0131  ;
  input \P1_EBX_reg[1]/NET0131  ;
  input \P1_EBX_reg[20]/NET0131  ;
  input \P1_EBX_reg[21]/NET0131  ;
  input \P1_EBX_reg[22]/NET0131  ;
  input \P1_EBX_reg[23]/NET0131  ;
  input \P1_EBX_reg[24]/NET0131  ;
  input \P1_EBX_reg[25]/NET0131  ;
  input \P1_EBX_reg[26]/NET0131  ;
  input \P1_EBX_reg[27]/NET0131  ;
  input \P1_EBX_reg[28]/NET0131  ;
  input \P1_EBX_reg[29]/NET0131  ;
  input \P1_EBX_reg[2]/NET0131  ;
  input \P1_EBX_reg[30]/NET0131  ;
  input \P1_EBX_reg[31]/NET0131  ;
  input \P1_EBX_reg[3]/NET0131  ;
  input \P1_EBX_reg[4]/NET0131  ;
  input \P1_EBX_reg[5]/NET0131  ;
  input \P1_EBX_reg[6]/NET0131  ;
  input \P1_EBX_reg[7]/NET0131  ;
  input \P1_EBX_reg[8]/NET0131  ;
  input \P1_EBX_reg[9]/NET0131  ;
  input \P1_Flush_reg/NET0131  ;
  input \P1_InstAddrPointer_reg[0]/NET0131  ;
  input \P1_InstAddrPointer_reg[10]/NET0131  ;
  input \P1_InstAddrPointer_reg[11]/NET0131  ;
  input \P1_InstAddrPointer_reg[12]/NET0131  ;
  input \P1_InstAddrPointer_reg[13]/NET0131  ;
  input \P1_InstAddrPointer_reg[14]/NET0131  ;
  input \P1_InstAddrPointer_reg[15]/NET0131  ;
  input \P1_InstAddrPointer_reg[16]/NET0131  ;
  input \P1_InstAddrPointer_reg[17]/NET0131  ;
  input \P1_InstAddrPointer_reg[18]/NET0131  ;
  input \P1_InstAddrPointer_reg[19]/NET0131  ;
  input \P1_InstAddrPointer_reg[1]/NET0131  ;
  input \P1_InstAddrPointer_reg[20]/NET0131  ;
  input \P1_InstAddrPointer_reg[21]/NET0131  ;
  input \P1_InstAddrPointer_reg[22]/NET0131  ;
  input \P1_InstAddrPointer_reg[23]/NET0131  ;
  input \P1_InstAddrPointer_reg[24]/NET0131  ;
  input \P1_InstAddrPointer_reg[25]/NET0131  ;
  input \P1_InstAddrPointer_reg[26]/NET0131  ;
  input \P1_InstAddrPointer_reg[27]/NET0131  ;
  input \P1_InstAddrPointer_reg[28]/NET0131  ;
  input \P1_InstAddrPointer_reg[29]/NET0131  ;
  input \P1_InstAddrPointer_reg[2]/NET0131  ;
  input \P1_InstAddrPointer_reg[30]/NET0131  ;
  input \P1_InstAddrPointer_reg[31]/NET0131  ;
  input \P1_InstAddrPointer_reg[3]/NET0131  ;
  input \P1_InstAddrPointer_reg[4]/NET0131  ;
  input \P1_InstAddrPointer_reg[5]/NET0131  ;
  input \P1_InstAddrPointer_reg[6]/NET0131  ;
  input \P1_InstAddrPointer_reg[7]/NET0131  ;
  input \P1_InstAddrPointer_reg[8]/NET0131  ;
  input \P1_InstAddrPointer_reg[9]/NET0131  ;
  input \P1_InstQueueRd_Addr_reg[0]/NET0131  ;
  input \P1_InstQueueRd_Addr_reg[1]/NET0131  ;
  input \P1_InstQueueRd_Addr_reg[2]/NET0131  ;
  input \P1_InstQueueRd_Addr_reg[3]/NET0131  ;
  input \P1_InstQueueWr_Addr_reg[0]/NET0131  ;
  input \P1_InstQueueWr_Addr_reg[1]/NET0131  ;
  input \P1_InstQueueWr_Addr_reg[2]/NET0131  ;
  input \P1_InstQueueWr_Addr_reg[3]/NET0131  ;
  input \P1_InstQueue_reg[0][0]/NET0131  ;
  input \P1_InstQueue_reg[0][1]/NET0131  ;
  input \P1_InstQueue_reg[0][2]/NET0131  ;
  input \P1_InstQueue_reg[0][3]/NET0131  ;
  input \P1_InstQueue_reg[0][4]/NET0131  ;
  input \P1_InstQueue_reg[0][5]/NET0131  ;
  input \P1_InstQueue_reg[0][6]/NET0131  ;
  input \P1_InstQueue_reg[0][7]/NET0131  ;
  input \P1_InstQueue_reg[10][0]/NET0131  ;
  input \P1_InstQueue_reg[10][1]/NET0131  ;
  input \P1_InstQueue_reg[10][2]/NET0131  ;
  input \P1_InstQueue_reg[10][3]/NET0131  ;
  input \P1_InstQueue_reg[10][4]/NET0131  ;
  input \P1_InstQueue_reg[10][5]/NET0131  ;
  input \P1_InstQueue_reg[10][6]/NET0131  ;
  input \P1_InstQueue_reg[10][7]/NET0131  ;
  input \P1_InstQueue_reg[11][0]/NET0131  ;
  input \P1_InstQueue_reg[11][1]/NET0131  ;
  input \P1_InstQueue_reg[11][2]/NET0131  ;
  input \P1_InstQueue_reg[11][3]/NET0131  ;
  input \P1_InstQueue_reg[11][4]/NET0131  ;
  input \P1_InstQueue_reg[11][5]/NET0131  ;
  input \P1_InstQueue_reg[11][6]/NET0131  ;
  input \P1_InstQueue_reg[11][7]/NET0131  ;
  input \P1_InstQueue_reg[12][0]/NET0131  ;
  input \P1_InstQueue_reg[12][1]/NET0131  ;
  input \P1_InstQueue_reg[12][2]/NET0131  ;
  input \P1_InstQueue_reg[12][3]/NET0131  ;
  input \P1_InstQueue_reg[12][4]/NET0131  ;
  input \P1_InstQueue_reg[12][5]/NET0131  ;
  input \P1_InstQueue_reg[12][6]/NET0131  ;
  input \P1_InstQueue_reg[12][7]/NET0131  ;
  input \P1_InstQueue_reg[13][0]/NET0131  ;
  input \P1_InstQueue_reg[13][1]/NET0131  ;
  input \P1_InstQueue_reg[13][2]/NET0131  ;
  input \P1_InstQueue_reg[13][3]/NET0131  ;
  input \P1_InstQueue_reg[13][4]/NET0131  ;
  input \P1_InstQueue_reg[13][5]/NET0131  ;
  input \P1_InstQueue_reg[13][6]/NET0131  ;
  input \P1_InstQueue_reg[13][7]/NET0131  ;
  input \P1_InstQueue_reg[14][0]/NET0131  ;
  input \P1_InstQueue_reg[14][1]/NET0131  ;
  input \P1_InstQueue_reg[14][2]/NET0131  ;
  input \P1_InstQueue_reg[14][3]/NET0131  ;
  input \P1_InstQueue_reg[14][4]/NET0131  ;
  input \P1_InstQueue_reg[14][5]/NET0131  ;
  input \P1_InstQueue_reg[14][6]/NET0131  ;
  input \P1_InstQueue_reg[14][7]/NET0131  ;
  input \P1_InstQueue_reg[15][0]/NET0131  ;
  input \P1_InstQueue_reg[15][1]/NET0131  ;
  input \P1_InstQueue_reg[15][2]/NET0131  ;
  input \P1_InstQueue_reg[15][3]/NET0131  ;
  input \P1_InstQueue_reg[15][4]/NET0131  ;
  input \P1_InstQueue_reg[15][5]/NET0131  ;
  input \P1_InstQueue_reg[15][6]/NET0131  ;
  input \P1_InstQueue_reg[15][7]/NET0131  ;
  input \P1_InstQueue_reg[1][0]/NET0131  ;
  input \P1_InstQueue_reg[1][1]/NET0131  ;
  input \P1_InstQueue_reg[1][2]/NET0131  ;
  input \P1_InstQueue_reg[1][3]/NET0131  ;
  input \P1_InstQueue_reg[1][4]/NET0131  ;
  input \P1_InstQueue_reg[1][5]/NET0131  ;
  input \P1_InstQueue_reg[1][6]/NET0131  ;
  input \P1_InstQueue_reg[1][7]/NET0131  ;
  input \P1_InstQueue_reg[2][0]/NET0131  ;
  input \P1_InstQueue_reg[2][1]/NET0131  ;
  input \P1_InstQueue_reg[2][2]/NET0131  ;
  input \P1_InstQueue_reg[2][3]/NET0131  ;
  input \P1_InstQueue_reg[2][4]/NET0131  ;
  input \P1_InstQueue_reg[2][5]/NET0131  ;
  input \P1_InstQueue_reg[2][6]/NET0131  ;
  input \P1_InstQueue_reg[2][7]/NET0131  ;
  input \P1_InstQueue_reg[3][0]/NET0131  ;
  input \P1_InstQueue_reg[3][1]/NET0131  ;
  input \P1_InstQueue_reg[3][2]/NET0131  ;
  input \P1_InstQueue_reg[3][3]/NET0131  ;
  input \P1_InstQueue_reg[3][4]/NET0131  ;
  input \P1_InstQueue_reg[3][5]/NET0131  ;
  input \P1_InstQueue_reg[3][6]/NET0131  ;
  input \P1_InstQueue_reg[3][7]/NET0131  ;
  input \P1_InstQueue_reg[4][0]/NET0131  ;
  input \P1_InstQueue_reg[4][1]/NET0131  ;
  input \P1_InstQueue_reg[4][2]/NET0131  ;
  input \P1_InstQueue_reg[4][3]/NET0131  ;
  input \P1_InstQueue_reg[4][4]/NET0131  ;
  input \P1_InstQueue_reg[4][5]/NET0131  ;
  input \P1_InstQueue_reg[4][6]/NET0131  ;
  input \P1_InstQueue_reg[4][7]/NET0131  ;
  input \P1_InstQueue_reg[5][0]/NET0131  ;
  input \P1_InstQueue_reg[5][1]/NET0131  ;
  input \P1_InstQueue_reg[5][2]/NET0131  ;
  input \P1_InstQueue_reg[5][3]/NET0131  ;
  input \P1_InstQueue_reg[5][4]/NET0131  ;
  input \P1_InstQueue_reg[5][5]/NET0131  ;
  input \P1_InstQueue_reg[5][6]/NET0131  ;
  input \P1_InstQueue_reg[5][7]/NET0131  ;
  input \P1_InstQueue_reg[6][0]/NET0131  ;
  input \P1_InstQueue_reg[6][1]/NET0131  ;
  input \P1_InstQueue_reg[6][2]/NET0131  ;
  input \P1_InstQueue_reg[6][3]/NET0131  ;
  input \P1_InstQueue_reg[6][4]/NET0131  ;
  input \P1_InstQueue_reg[6][5]/NET0131  ;
  input \P1_InstQueue_reg[6][6]/NET0131  ;
  input \P1_InstQueue_reg[6][7]/NET0131  ;
  input \P1_InstQueue_reg[7][0]/NET0131  ;
  input \P1_InstQueue_reg[7][1]/NET0131  ;
  input \P1_InstQueue_reg[7][2]/NET0131  ;
  input \P1_InstQueue_reg[7][3]/NET0131  ;
  input \P1_InstQueue_reg[7][4]/NET0131  ;
  input \P1_InstQueue_reg[7][5]/NET0131  ;
  input \P1_InstQueue_reg[7][6]/NET0131  ;
  input \P1_InstQueue_reg[7][7]/NET0131  ;
  input \P1_InstQueue_reg[8][0]/NET0131  ;
  input \P1_InstQueue_reg[8][1]/NET0131  ;
  input \P1_InstQueue_reg[8][2]/NET0131  ;
  input \P1_InstQueue_reg[8][3]/NET0131  ;
  input \P1_InstQueue_reg[8][4]/NET0131  ;
  input \P1_InstQueue_reg[8][5]/NET0131  ;
  input \P1_InstQueue_reg[8][6]/NET0131  ;
  input \P1_InstQueue_reg[8][7]/NET0131  ;
  input \P1_InstQueue_reg[9][0]/NET0131  ;
  input \P1_InstQueue_reg[9][1]/NET0131  ;
  input \P1_InstQueue_reg[9][2]/NET0131  ;
  input \P1_InstQueue_reg[9][3]/NET0131  ;
  input \P1_InstQueue_reg[9][4]/NET0131  ;
  input \P1_InstQueue_reg[9][5]/NET0131  ;
  input \P1_InstQueue_reg[9][6]/NET0131  ;
  input \P1_InstQueue_reg[9][7]/NET0131  ;
  input \P1_M_IO_n_reg/NET0131  ;
  input \P1_MemoryFetch_reg/NET0131  ;
  input \P1_More_reg/NET0131  ;
  input \P1_PhyAddrPointer_reg[0]/NET0131  ;
  input \P1_PhyAddrPointer_reg[10]/NET0131  ;
  input \P1_PhyAddrPointer_reg[11]/NET0131  ;
  input \P1_PhyAddrPointer_reg[12]/NET0131  ;
  input \P1_PhyAddrPointer_reg[13]/NET0131  ;
  input \P1_PhyAddrPointer_reg[14]/NET0131  ;
  input \P1_PhyAddrPointer_reg[15]/NET0131  ;
  input \P1_PhyAddrPointer_reg[16]/NET0131  ;
  input \P1_PhyAddrPointer_reg[17]/NET0131  ;
  input \P1_PhyAddrPointer_reg[18]/NET0131  ;
  input \P1_PhyAddrPointer_reg[19]/NET0131  ;
  input \P1_PhyAddrPointer_reg[1]/NET0131  ;
  input \P1_PhyAddrPointer_reg[20]/NET0131  ;
  input \P1_PhyAddrPointer_reg[21]/NET0131  ;
  input \P1_PhyAddrPointer_reg[22]/NET0131  ;
  input \P1_PhyAddrPointer_reg[23]/NET0131  ;
  input \P1_PhyAddrPointer_reg[24]/NET0131  ;
  input \P1_PhyAddrPointer_reg[25]/NET0131  ;
  input \P1_PhyAddrPointer_reg[26]/NET0131  ;
  input \P1_PhyAddrPointer_reg[27]/NET0131  ;
  input \P1_PhyAddrPointer_reg[28]/NET0131  ;
  input \P1_PhyAddrPointer_reg[29]/NET0131  ;
  input \P1_PhyAddrPointer_reg[2]/NET0131  ;
  input \P1_PhyAddrPointer_reg[30]/NET0131  ;
  input \P1_PhyAddrPointer_reg[31]/NET0131  ;
  input \P1_PhyAddrPointer_reg[3]/NET0131  ;
  input \P1_PhyAddrPointer_reg[4]/NET0131  ;
  input \P1_PhyAddrPointer_reg[5]/NET0131  ;
  input \P1_PhyAddrPointer_reg[6]/NET0131  ;
  input \P1_PhyAddrPointer_reg[7]/NET0131  ;
  input \P1_PhyAddrPointer_reg[8]/NET0131  ;
  input \P1_PhyAddrPointer_reg[9]/NET0131  ;
  input \P1_ReadRequest_reg/NET0131  ;
  input \P1_RequestPending_reg/NET0131  ;
  input \P1_State2_reg[0]/NET0131  ;
  input \P1_State2_reg[1]/NET0131  ;
  input \P1_State2_reg[2]/NET0131  ;
  input \P1_State2_reg[3]/NET0131  ;
  input \P1_State_reg[0]/NET0131  ;
  input \P1_State_reg[1]/NET0131  ;
  input \P1_State_reg[2]/NET0131  ;
  input \P1_W_R_n_reg/NET0131  ;
  input \P1_lWord_reg[0]/NET0131  ;
  input \P1_lWord_reg[10]/NET0131  ;
  input \P1_lWord_reg[11]/NET0131  ;
  input \P1_lWord_reg[12]/NET0131  ;
  input \P1_lWord_reg[13]/NET0131  ;
  input \P1_lWord_reg[14]/NET0131  ;
  input \P1_lWord_reg[15]/NET0131  ;
  input \P1_lWord_reg[1]/NET0131  ;
  input \P1_lWord_reg[2]/NET0131  ;
  input \P1_lWord_reg[3]/NET0131  ;
  input \P1_lWord_reg[4]/NET0131  ;
  input \P1_lWord_reg[5]/NET0131  ;
  input \P1_lWord_reg[6]/NET0131  ;
  input \P1_lWord_reg[7]/NET0131  ;
  input \P1_lWord_reg[8]/NET0131  ;
  input \P1_lWord_reg[9]/NET0131  ;
  input \P1_rEIP_reg[0]/NET0131  ;
  input \P1_rEIP_reg[10]/NET0131  ;
  input \P1_rEIP_reg[11]/NET0131  ;
  input \P1_rEIP_reg[12]/NET0131  ;
  input \P1_rEIP_reg[13]/NET0131  ;
  input \P1_rEIP_reg[14]/NET0131  ;
  input \P1_rEIP_reg[15]/NET0131  ;
  input \P1_rEIP_reg[16]/NET0131  ;
  input \P1_rEIP_reg[17]/NET0131  ;
  input \P1_rEIP_reg[18]/NET0131  ;
  input \P1_rEIP_reg[19]/NET0131  ;
  input \P1_rEIP_reg[1]/NET0131  ;
  input \P1_rEIP_reg[20]/NET0131  ;
  input \P1_rEIP_reg[21]/NET0131  ;
  input \P1_rEIP_reg[22]/NET0131  ;
  input \P1_rEIP_reg[23]/NET0131  ;
  input \P1_rEIP_reg[24]/NET0131  ;
  input \P1_rEIP_reg[25]/NET0131  ;
  input \P1_rEIP_reg[26]/NET0131  ;
  input \P1_rEIP_reg[27]/NET0131  ;
  input \P1_rEIP_reg[28]/NET0131  ;
  input \P1_rEIP_reg[29]/NET0131  ;
  input \P1_rEIP_reg[2]/NET0131  ;
  input \P1_rEIP_reg[30]/NET0131  ;
  input \P1_rEIP_reg[31]/NET0131  ;
  input \P1_rEIP_reg[3]/NET0131  ;
  input \P1_rEIP_reg[4]/NET0131  ;
  input \P1_rEIP_reg[5]/NET0131  ;
  input \P1_rEIP_reg[6]/NET0131  ;
  input \P1_rEIP_reg[7]/NET0131  ;
  input \P1_rEIP_reg[8]/NET0131  ;
  input \P1_rEIP_reg[9]/NET0131  ;
  input \P1_uWord_reg[0]/NET0131  ;
  input \P1_uWord_reg[10]/NET0131  ;
  input \P1_uWord_reg[11]/NET0131  ;
  input \P1_uWord_reg[12]/NET0131  ;
  input \P1_uWord_reg[13]/NET0131  ;
  input \P1_uWord_reg[14]/NET0131  ;
  input \P1_uWord_reg[1]/NET0131  ;
  input \P1_uWord_reg[2]/NET0131  ;
  input \P1_uWord_reg[3]/NET0131  ;
  input \P1_uWord_reg[4]/NET0131  ;
  input \P1_uWord_reg[5]/NET0131  ;
  input \P1_uWord_reg[6]/NET0131  ;
  input \P1_uWord_reg[7]/NET0131  ;
  input \P1_uWord_reg[8]/NET0131  ;
  input \P1_uWord_reg[9]/NET0131  ;
  input \P2_ADS_n_reg/NET0131  ;
  input \P2_Address_reg[0]/NET0131  ;
  input \P2_Address_reg[10]/NET0131  ;
  input \P2_Address_reg[11]/NET0131  ;
  input \P2_Address_reg[12]/NET0131  ;
  input \P2_Address_reg[13]/NET0131  ;
  input \P2_Address_reg[14]/NET0131  ;
  input \P2_Address_reg[15]/NET0131  ;
  input \P2_Address_reg[16]/NET0131  ;
  input \P2_Address_reg[17]/NET0131  ;
  input \P2_Address_reg[18]/NET0131  ;
  input \P2_Address_reg[19]/NET0131  ;
  input \P2_Address_reg[1]/NET0131  ;
  input \P2_Address_reg[20]/NET0131  ;
  input \P2_Address_reg[21]/NET0131  ;
  input \P2_Address_reg[22]/NET0131  ;
  input \P2_Address_reg[23]/NET0131  ;
  input \P2_Address_reg[24]/NET0131  ;
  input \P2_Address_reg[25]/NET0131  ;
  input \P2_Address_reg[26]/NET0131  ;
  input \P2_Address_reg[27]/NET0131  ;
  input \P2_Address_reg[28]/NET0131  ;
  input \P2_Address_reg[29]/NET0131  ;
  input \P2_Address_reg[2]/NET0131  ;
  input \P2_Address_reg[3]/NET0131  ;
  input \P2_Address_reg[4]/NET0131  ;
  input \P2_Address_reg[5]/NET0131  ;
  input \P2_Address_reg[6]/NET0131  ;
  input \P2_Address_reg[7]/NET0131  ;
  input \P2_Address_reg[8]/NET0131  ;
  input \P2_Address_reg[9]/NET0131  ;
  input \P2_BE_n_reg[0]/NET0131  ;
  input \P2_BE_n_reg[1]/NET0131  ;
  input \P2_BE_n_reg[2]/NET0131  ;
  input \P2_BE_n_reg[3]/NET0131  ;
  input \P2_ByteEnable_reg[0]/NET0131  ;
  input \P2_ByteEnable_reg[1]/NET0131  ;
  input \P2_ByteEnable_reg[2]/NET0131  ;
  input \P2_ByteEnable_reg[3]/NET0131  ;
  input \P2_CodeFetch_reg/NET0131  ;
  input \P2_D_C_n_reg/NET0131  ;
  input \P2_DataWidth_reg[0]/NET0131  ;
  input \P2_DataWidth_reg[1]/NET0131  ;
  input \P2_Datao_reg[0]/NET0131  ;
  input \P2_Datao_reg[10]/NET0131  ;
  input \P2_Datao_reg[11]/NET0131  ;
  input \P2_Datao_reg[12]/NET0131  ;
  input \P2_Datao_reg[13]/NET0131  ;
  input \P2_Datao_reg[14]/NET0131  ;
  input \P2_Datao_reg[15]/NET0131  ;
  input \P2_Datao_reg[16]/NET0131  ;
  input \P2_Datao_reg[17]/NET0131  ;
  input \P2_Datao_reg[18]/NET0131  ;
  input \P2_Datao_reg[19]/NET0131  ;
  input \P2_Datao_reg[1]/NET0131  ;
  input \P2_Datao_reg[20]/NET0131  ;
  input \P2_Datao_reg[21]/NET0131  ;
  input \P2_Datao_reg[22]/NET0131  ;
  input \P2_Datao_reg[23]/NET0131  ;
  input \P2_Datao_reg[24]/NET0131  ;
  input \P2_Datao_reg[25]/NET0131  ;
  input \P2_Datao_reg[26]/NET0131  ;
  input \P2_Datao_reg[27]/NET0131  ;
  input \P2_Datao_reg[28]/NET0131  ;
  input \P2_Datao_reg[29]/NET0131  ;
  input \P2_Datao_reg[2]/NET0131  ;
  input \P2_Datao_reg[30]/NET0131  ;
  input \P2_Datao_reg[3]/NET0131  ;
  input \P2_Datao_reg[4]/NET0131  ;
  input \P2_Datao_reg[5]/NET0131  ;
  input \P2_Datao_reg[6]/NET0131  ;
  input \P2_Datao_reg[7]/NET0131  ;
  input \P2_Datao_reg[8]/NET0131  ;
  input \P2_Datao_reg[9]/NET0131  ;
  input \P2_EAX_reg[0]/NET0131  ;
  input \P2_EAX_reg[10]/NET0131  ;
  input \P2_EAX_reg[11]/NET0131  ;
  input \P2_EAX_reg[12]/NET0131  ;
  input \P2_EAX_reg[13]/NET0131  ;
  input \P2_EAX_reg[14]/NET0131  ;
  input \P2_EAX_reg[15]/NET0131  ;
  input \P2_EAX_reg[16]/NET0131  ;
  input \P2_EAX_reg[17]/NET0131  ;
  input \P2_EAX_reg[18]/NET0131  ;
  input \P2_EAX_reg[19]/NET0131  ;
  input \P2_EAX_reg[1]/NET0131  ;
  input \P2_EAX_reg[20]/NET0131  ;
  input \P2_EAX_reg[21]/NET0131  ;
  input \P2_EAX_reg[22]/NET0131  ;
  input \P2_EAX_reg[23]/NET0131  ;
  input \P2_EAX_reg[24]/NET0131  ;
  input \P2_EAX_reg[25]/NET0131  ;
  input \P2_EAX_reg[26]/NET0131  ;
  input \P2_EAX_reg[27]/NET0131  ;
  input \P2_EAX_reg[28]/NET0131  ;
  input \P2_EAX_reg[29]/NET0131  ;
  input \P2_EAX_reg[2]/NET0131  ;
  input \P2_EAX_reg[30]/NET0131  ;
  input \P2_EAX_reg[31]/NET0131  ;
  input \P2_EAX_reg[3]/NET0131  ;
  input \P2_EAX_reg[4]/NET0131  ;
  input \P2_EAX_reg[5]/NET0131  ;
  input \P2_EAX_reg[6]/NET0131  ;
  input \P2_EAX_reg[7]/NET0131  ;
  input \P2_EAX_reg[8]/NET0131  ;
  input \P2_EAX_reg[9]/NET0131  ;
  input \P2_EBX_reg[0]/NET0131  ;
  input \P2_EBX_reg[10]/NET0131  ;
  input \P2_EBX_reg[11]/NET0131  ;
  input \P2_EBX_reg[12]/NET0131  ;
  input \P2_EBX_reg[13]/NET0131  ;
  input \P2_EBX_reg[14]/NET0131  ;
  input \P2_EBX_reg[15]/NET0131  ;
  input \P2_EBX_reg[16]/NET0131  ;
  input \P2_EBX_reg[17]/NET0131  ;
  input \P2_EBX_reg[18]/NET0131  ;
  input \P2_EBX_reg[19]/NET0131  ;
  input \P2_EBX_reg[1]/NET0131  ;
  input \P2_EBX_reg[20]/NET0131  ;
  input \P2_EBX_reg[21]/NET0131  ;
  input \P2_EBX_reg[22]/NET0131  ;
  input \P2_EBX_reg[23]/NET0131  ;
  input \P2_EBX_reg[24]/NET0131  ;
  input \P2_EBX_reg[25]/NET0131  ;
  input \P2_EBX_reg[26]/NET0131  ;
  input \P2_EBX_reg[27]/NET0131  ;
  input \P2_EBX_reg[28]/NET0131  ;
  input \P2_EBX_reg[29]/NET0131  ;
  input \P2_EBX_reg[2]/NET0131  ;
  input \P2_EBX_reg[30]/NET0131  ;
  input \P2_EBX_reg[31]/NET0131  ;
  input \P2_EBX_reg[3]/NET0131  ;
  input \P2_EBX_reg[4]/NET0131  ;
  input \P2_EBX_reg[5]/NET0131  ;
  input \P2_EBX_reg[6]/NET0131  ;
  input \P2_EBX_reg[7]/NET0131  ;
  input \P2_EBX_reg[8]/NET0131  ;
  input \P2_EBX_reg[9]/NET0131  ;
  input \P2_Flush_reg/NET0131  ;
  input \P2_InstAddrPointer_reg[0]/NET0131  ;
  input \P2_InstAddrPointer_reg[10]/NET0131  ;
  input \P2_InstAddrPointer_reg[11]/NET0131  ;
  input \P2_InstAddrPointer_reg[12]/NET0131  ;
  input \P2_InstAddrPointer_reg[13]/NET0131  ;
  input \P2_InstAddrPointer_reg[14]/NET0131  ;
  input \P2_InstAddrPointer_reg[15]/NET0131  ;
  input \P2_InstAddrPointer_reg[16]/NET0131  ;
  input \P2_InstAddrPointer_reg[17]/NET0131  ;
  input \P2_InstAddrPointer_reg[18]/NET0131  ;
  input \P2_InstAddrPointer_reg[19]/NET0131  ;
  input \P2_InstAddrPointer_reg[1]/NET0131  ;
  input \P2_InstAddrPointer_reg[20]/NET0131  ;
  input \P2_InstAddrPointer_reg[21]/NET0131  ;
  input \P2_InstAddrPointer_reg[22]/NET0131  ;
  input \P2_InstAddrPointer_reg[23]/NET0131  ;
  input \P2_InstAddrPointer_reg[24]/NET0131  ;
  input \P2_InstAddrPointer_reg[25]/NET0131  ;
  input \P2_InstAddrPointer_reg[26]/NET0131  ;
  input \P2_InstAddrPointer_reg[27]/NET0131  ;
  input \P2_InstAddrPointer_reg[28]/NET0131  ;
  input \P2_InstAddrPointer_reg[29]/NET0131  ;
  input \P2_InstAddrPointer_reg[2]/NET0131  ;
  input \P2_InstAddrPointer_reg[30]/NET0131  ;
  input \P2_InstAddrPointer_reg[31]/NET0131  ;
  input \P2_InstAddrPointer_reg[3]/NET0131  ;
  input \P2_InstAddrPointer_reg[4]/NET0131  ;
  input \P2_InstAddrPointer_reg[5]/NET0131  ;
  input \P2_InstAddrPointer_reg[6]/NET0131  ;
  input \P2_InstAddrPointer_reg[7]/NET0131  ;
  input \P2_InstAddrPointer_reg[8]/NET0131  ;
  input \P2_InstAddrPointer_reg[9]/NET0131  ;
  input \P2_InstQueueRd_Addr_reg[0]/NET0131  ;
  input \P2_InstQueueRd_Addr_reg[1]/NET0131  ;
  input \P2_InstQueueRd_Addr_reg[2]/NET0131  ;
  input \P2_InstQueueRd_Addr_reg[3]/NET0131  ;
  input \P2_InstQueueWr_Addr_reg[0]/NET0131  ;
  input \P2_InstQueueWr_Addr_reg[1]/NET0131  ;
  input \P2_InstQueueWr_Addr_reg[2]/NET0131  ;
  input \P2_InstQueueWr_Addr_reg[3]/NET0131  ;
  input \P2_InstQueue_reg[0][0]/NET0131  ;
  input \P2_InstQueue_reg[0][1]/NET0131  ;
  input \P2_InstQueue_reg[0][2]/NET0131  ;
  input \P2_InstQueue_reg[0][3]/NET0131  ;
  input \P2_InstQueue_reg[0][4]/NET0131  ;
  input \P2_InstQueue_reg[0][5]/NET0131  ;
  input \P2_InstQueue_reg[0][6]/NET0131  ;
  input \P2_InstQueue_reg[0][7]/NET0131  ;
  input \P2_InstQueue_reg[10][0]/NET0131  ;
  input \P2_InstQueue_reg[10][1]/NET0131  ;
  input \P2_InstQueue_reg[10][2]/NET0131  ;
  input \P2_InstQueue_reg[10][3]/NET0131  ;
  input \P2_InstQueue_reg[10][4]/NET0131  ;
  input \P2_InstQueue_reg[10][5]/NET0131  ;
  input \P2_InstQueue_reg[10][6]/NET0131  ;
  input \P2_InstQueue_reg[10][7]/NET0131  ;
  input \P2_InstQueue_reg[11][0]/NET0131  ;
  input \P2_InstQueue_reg[11][1]/NET0131  ;
  input \P2_InstQueue_reg[11][2]/NET0131  ;
  input \P2_InstQueue_reg[11][3]/NET0131  ;
  input \P2_InstQueue_reg[11][4]/NET0131  ;
  input \P2_InstQueue_reg[11][5]/NET0131  ;
  input \P2_InstQueue_reg[11][6]/NET0131  ;
  input \P2_InstQueue_reg[11][7]/NET0131  ;
  input \P2_InstQueue_reg[12][0]/NET0131  ;
  input \P2_InstQueue_reg[12][1]/NET0131  ;
  input \P2_InstQueue_reg[12][2]/NET0131  ;
  input \P2_InstQueue_reg[12][3]/NET0131  ;
  input \P2_InstQueue_reg[12][4]/NET0131  ;
  input \P2_InstQueue_reg[12][5]/NET0131  ;
  input \P2_InstQueue_reg[12][6]/NET0131  ;
  input \P2_InstQueue_reg[12][7]/NET0131  ;
  input \P2_InstQueue_reg[13][0]/NET0131  ;
  input \P2_InstQueue_reg[13][1]/NET0131  ;
  input \P2_InstQueue_reg[13][2]/NET0131  ;
  input \P2_InstQueue_reg[13][3]/NET0131  ;
  input \P2_InstQueue_reg[13][4]/NET0131  ;
  input \P2_InstQueue_reg[13][5]/NET0131  ;
  input \P2_InstQueue_reg[13][6]/NET0131  ;
  input \P2_InstQueue_reg[13][7]/NET0131  ;
  input \P2_InstQueue_reg[14][0]/NET0131  ;
  input \P2_InstQueue_reg[14][1]/NET0131  ;
  input \P2_InstQueue_reg[14][2]/NET0131  ;
  input \P2_InstQueue_reg[14][3]/NET0131  ;
  input \P2_InstQueue_reg[14][4]/NET0131  ;
  input \P2_InstQueue_reg[14][5]/NET0131  ;
  input \P2_InstQueue_reg[14][6]/NET0131  ;
  input \P2_InstQueue_reg[14][7]/NET0131  ;
  input \P2_InstQueue_reg[15][0]/NET0131  ;
  input \P2_InstQueue_reg[15][1]/NET0131  ;
  input \P2_InstQueue_reg[15][2]/NET0131  ;
  input \P2_InstQueue_reg[15][3]/NET0131  ;
  input \P2_InstQueue_reg[15][4]/NET0131  ;
  input \P2_InstQueue_reg[15][5]/NET0131  ;
  input \P2_InstQueue_reg[15][6]/NET0131  ;
  input \P2_InstQueue_reg[15][7]/NET0131  ;
  input \P2_InstQueue_reg[1][0]/NET0131  ;
  input \P2_InstQueue_reg[1][1]/NET0131  ;
  input \P2_InstQueue_reg[1][2]/NET0131  ;
  input \P2_InstQueue_reg[1][3]/NET0131  ;
  input \P2_InstQueue_reg[1][4]/NET0131  ;
  input \P2_InstQueue_reg[1][5]/NET0131  ;
  input \P2_InstQueue_reg[1][6]/NET0131  ;
  input \P2_InstQueue_reg[1][7]/NET0131  ;
  input \P2_InstQueue_reg[2][0]/NET0131  ;
  input \P2_InstQueue_reg[2][1]/NET0131  ;
  input \P2_InstQueue_reg[2][2]/NET0131  ;
  input \P2_InstQueue_reg[2][3]/NET0131  ;
  input \P2_InstQueue_reg[2][4]/NET0131  ;
  input \P2_InstQueue_reg[2][5]/NET0131  ;
  input \P2_InstQueue_reg[2][6]/NET0131  ;
  input \P2_InstQueue_reg[2][7]/NET0131  ;
  input \P2_InstQueue_reg[3][0]/NET0131  ;
  input \P2_InstQueue_reg[3][1]/NET0131  ;
  input \P2_InstQueue_reg[3][2]/NET0131  ;
  input \P2_InstQueue_reg[3][3]/NET0131  ;
  input \P2_InstQueue_reg[3][4]/NET0131  ;
  input \P2_InstQueue_reg[3][5]/NET0131  ;
  input \P2_InstQueue_reg[3][6]/NET0131  ;
  input \P2_InstQueue_reg[3][7]/NET0131  ;
  input \P2_InstQueue_reg[4][0]/NET0131  ;
  input \P2_InstQueue_reg[4][1]/NET0131  ;
  input \P2_InstQueue_reg[4][2]/NET0131  ;
  input \P2_InstQueue_reg[4][3]/NET0131  ;
  input \P2_InstQueue_reg[4][4]/NET0131  ;
  input \P2_InstQueue_reg[4][5]/NET0131  ;
  input \P2_InstQueue_reg[4][6]/NET0131  ;
  input \P2_InstQueue_reg[4][7]/NET0131  ;
  input \P2_InstQueue_reg[5][0]/NET0131  ;
  input \P2_InstQueue_reg[5][1]/NET0131  ;
  input \P2_InstQueue_reg[5][2]/NET0131  ;
  input \P2_InstQueue_reg[5][3]/NET0131  ;
  input \P2_InstQueue_reg[5][4]/NET0131  ;
  input \P2_InstQueue_reg[5][5]/NET0131  ;
  input \P2_InstQueue_reg[5][6]/NET0131  ;
  input \P2_InstQueue_reg[5][7]/NET0131  ;
  input \P2_InstQueue_reg[6][0]/NET0131  ;
  input \P2_InstQueue_reg[6][1]/NET0131  ;
  input \P2_InstQueue_reg[6][2]/NET0131  ;
  input \P2_InstQueue_reg[6][3]/NET0131  ;
  input \P2_InstQueue_reg[6][4]/NET0131  ;
  input \P2_InstQueue_reg[6][5]/NET0131  ;
  input \P2_InstQueue_reg[6][6]/NET0131  ;
  input \P2_InstQueue_reg[6][7]/NET0131  ;
  input \P2_InstQueue_reg[7][0]/NET0131  ;
  input \P2_InstQueue_reg[7][1]/NET0131  ;
  input \P2_InstQueue_reg[7][2]/NET0131  ;
  input \P2_InstQueue_reg[7][3]/NET0131  ;
  input \P2_InstQueue_reg[7][4]/NET0131  ;
  input \P2_InstQueue_reg[7][5]/NET0131  ;
  input \P2_InstQueue_reg[7][6]/NET0131  ;
  input \P2_InstQueue_reg[7][7]/NET0131  ;
  input \P2_InstQueue_reg[8][0]/NET0131  ;
  input \P2_InstQueue_reg[8][1]/NET0131  ;
  input \P2_InstQueue_reg[8][2]/NET0131  ;
  input \P2_InstQueue_reg[8][3]/NET0131  ;
  input \P2_InstQueue_reg[8][4]/NET0131  ;
  input \P2_InstQueue_reg[8][5]/NET0131  ;
  input \P2_InstQueue_reg[8][6]/NET0131  ;
  input \P2_InstQueue_reg[8][7]/NET0131  ;
  input \P2_InstQueue_reg[9][0]/NET0131  ;
  input \P2_InstQueue_reg[9][1]/NET0131  ;
  input \P2_InstQueue_reg[9][2]/NET0131  ;
  input \P2_InstQueue_reg[9][3]/NET0131  ;
  input \P2_InstQueue_reg[9][4]/NET0131  ;
  input \P2_InstQueue_reg[9][5]/NET0131  ;
  input \P2_InstQueue_reg[9][6]/NET0131  ;
  input \P2_InstQueue_reg[9][7]/NET0131  ;
  input \P2_M_IO_n_reg/NET0131  ;
  input \P2_MemoryFetch_reg/NET0131  ;
  input \P2_More_reg/NET0131  ;
  input \P2_PhyAddrPointer_reg[0]/NET0131  ;
  input \P2_PhyAddrPointer_reg[10]/NET0131  ;
  input \P2_PhyAddrPointer_reg[11]/NET0131  ;
  input \P2_PhyAddrPointer_reg[12]/NET0131  ;
  input \P2_PhyAddrPointer_reg[13]/NET0131  ;
  input \P2_PhyAddrPointer_reg[14]/NET0131  ;
  input \P2_PhyAddrPointer_reg[15]/NET0131  ;
  input \P2_PhyAddrPointer_reg[16]/NET0131  ;
  input \P2_PhyAddrPointer_reg[17]/NET0131  ;
  input \P2_PhyAddrPointer_reg[18]/NET0131  ;
  input \P2_PhyAddrPointer_reg[19]/NET0131  ;
  input \P2_PhyAddrPointer_reg[1]/NET0131  ;
  input \P2_PhyAddrPointer_reg[20]/NET0131  ;
  input \P2_PhyAddrPointer_reg[21]/NET0131  ;
  input \P2_PhyAddrPointer_reg[22]/NET0131  ;
  input \P2_PhyAddrPointer_reg[23]/NET0131  ;
  input \P2_PhyAddrPointer_reg[24]/NET0131  ;
  input \P2_PhyAddrPointer_reg[25]/NET0131  ;
  input \P2_PhyAddrPointer_reg[26]/NET0131  ;
  input \P2_PhyAddrPointer_reg[27]/NET0131  ;
  input \P2_PhyAddrPointer_reg[28]/NET0131  ;
  input \P2_PhyAddrPointer_reg[29]/NET0131  ;
  input \P2_PhyAddrPointer_reg[2]/NET0131  ;
  input \P2_PhyAddrPointer_reg[30]/NET0131  ;
  input \P2_PhyAddrPointer_reg[31]/NET0131  ;
  input \P2_PhyAddrPointer_reg[3]/NET0131  ;
  input \P2_PhyAddrPointer_reg[4]/NET0131  ;
  input \P2_PhyAddrPointer_reg[5]/NET0131  ;
  input \P2_PhyAddrPointer_reg[6]/NET0131  ;
  input \P2_PhyAddrPointer_reg[7]/NET0131  ;
  input \P2_PhyAddrPointer_reg[8]/NET0131  ;
  input \P2_PhyAddrPointer_reg[9]/NET0131  ;
  input \P2_ReadRequest_reg/NET0131  ;
  input \P2_RequestPending_reg/NET0131  ;
  input \P2_State2_reg[0]/NET0131  ;
  input \P2_State2_reg[1]/NET0131  ;
  input \P2_State2_reg[2]/NET0131  ;
  input \P2_State2_reg[3]/NET0131  ;
  input \P2_State_reg[0]/NET0131  ;
  input \P2_State_reg[1]/NET0131  ;
  input \P2_State_reg[2]/NET0131  ;
  input \P2_W_R_n_reg/NET0131  ;
  input \P2_lWord_reg[0]/NET0131  ;
  input \P2_lWord_reg[10]/NET0131  ;
  input \P2_lWord_reg[11]/NET0131  ;
  input \P2_lWord_reg[12]/NET0131  ;
  input \P2_lWord_reg[13]/NET0131  ;
  input \P2_lWord_reg[14]/NET0131  ;
  input \P2_lWord_reg[15]/NET0131  ;
  input \P2_lWord_reg[1]/NET0131  ;
  input \P2_lWord_reg[2]/NET0131  ;
  input \P2_lWord_reg[3]/NET0131  ;
  input \P2_lWord_reg[4]/NET0131  ;
  input \P2_lWord_reg[5]/NET0131  ;
  input \P2_lWord_reg[6]/NET0131  ;
  input \P2_lWord_reg[7]/NET0131  ;
  input \P2_lWord_reg[8]/NET0131  ;
  input \P2_lWord_reg[9]/NET0131  ;
  input \P2_rEIP_reg[0]/NET0131  ;
  input \P2_rEIP_reg[10]/NET0131  ;
  input \P2_rEIP_reg[11]/NET0131  ;
  input \P2_rEIP_reg[12]/NET0131  ;
  input \P2_rEIP_reg[13]/NET0131  ;
  input \P2_rEIP_reg[14]/NET0131  ;
  input \P2_rEIP_reg[15]/NET0131  ;
  input \P2_rEIP_reg[16]/NET0131  ;
  input \P2_rEIP_reg[17]/NET0131  ;
  input \P2_rEIP_reg[18]/NET0131  ;
  input \P2_rEIP_reg[19]/NET0131  ;
  input \P2_rEIP_reg[1]/NET0131  ;
  input \P2_rEIP_reg[20]/NET0131  ;
  input \P2_rEIP_reg[21]/NET0131  ;
  input \P2_rEIP_reg[22]/NET0131  ;
  input \P2_rEIP_reg[23]/NET0131  ;
  input \P2_rEIP_reg[24]/NET0131  ;
  input \P2_rEIP_reg[25]/NET0131  ;
  input \P2_rEIP_reg[26]/NET0131  ;
  input \P2_rEIP_reg[27]/NET0131  ;
  input \P2_rEIP_reg[28]/NET0131  ;
  input \P2_rEIP_reg[29]/NET0131  ;
  input \P2_rEIP_reg[2]/NET0131  ;
  input \P2_rEIP_reg[30]/NET0131  ;
  input \P2_rEIP_reg[31]/NET0131  ;
  input \P2_rEIP_reg[3]/NET0131  ;
  input \P2_rEIP_reg[4]/NET0131  ;
  input \P2_rEIP_reg[5]/NET0131  ;
  input \P2_rEIP_reg[6]/NET0131  ;
  input \P2_rEIP_reg[7]/NET0131  ;
  input \P2_rEIP_reg[8]/NET0131  ;
  input \P2_rEIP_reg[9]/NET0131  ;
  input \P2_uWord_reg[0]/NET0131  ;
  input \P2_uWord_reg[10]/NET0131  ;
  input \P2_uWord_reg[11]/NET0131  ;
  input \P2_uWord_reg[12]/NET0131  ;
  input \P2_uWord_reg[13]/NET0131  ;
  input \P2_uWord_reg[14]/NET0131  ;
  input \P2_uWord_reg[1]/NET0131  ;
  input \P2_uWord_reg[2]/NET0131  ;
  input \P2_uWord_reg[3]/NET0131  ;
  input \P2_uWord_reg[4]/NET0131  ;
  input \P2_uWord_reg[5]/NET0131  ;
  input \P2_uWord_reg[6]/NET0131  ;
  input \P2_uWord_reg[7]/NET0131  ;
  input \P2_uWord_reg[8]/NET0131  ;
  input \P2_uWord_reg[9]/NET0131  ;
  input \P3_Address_reg[0]/NET0131  ;
  input \P3_Address_reg[10]/NET0131  ;
  input \P3_Address_reg[11]/NET0131  ;
  input \P3_Address_reg[12]/NET0131  ;
  input \P3_Address_reg[13]/NET0131  ;
  input \P3_Address_reg[14]/NET0131  ;
  input \P3_Address_reg[15]/NET0131  ;
  input \P3_Address_reg[16]/NET0131  ;
  input \P3_Address_reg[17]/NET0131  ;
  input \P3_Address_reg[18]/NET0131  ;
  input \P3_Address_reg[19]/NET0131  ;
  input \P3_Address_reg[1]/NET0131  ;
  input \P3_Address_reg[20]/NET0131  ;
  input \P3_Address_reg[21]/NET0131  ;
  input \P3_Address_reg[22]/NET0131  ;
  input \P3_Address_reg[23]/NET0131  ;
  input \P3_Address_reg[24]/NET0131  ;
  input \P3_Address_reg[25]/NET0131  ;
  input \P3_Address_reg[26]/NET0131  ;
  input \P3_Address_reg[27]/NET0131  ;
  input \P3_Address_reg[28]/NET0131  ;
  input \P3_Address_reg[29]/NET0131  ;
  input \P3_Address_reg[2]/NET0131  ;
  input \P3_Address_reg[3]/NET0131  ;
  input \P3_Address_reg[4]/NET0131  ;
  input \P3_Address_reg[5]/NET0131  ;
  input \P3_Address_reg[6]/NET0131  ;
  input \P3_Address_reg[7]/NET0131  ;
  input \P3_Address_reg[8]/NET0131  ;
  input \P3_Address_reg[9]/NET0131  ;
  input \P3_BE_n_reg[0]/NET0131  ;
  input \P3_BE_n_reg[1]/NET0131  ;
  input \P3_BE_n_reg[2]/NET0131  ;
  input \P3_BE_n_reg[3]/NET0131  ;
  input \P3_ByteEnable_reg[0]/NET0131  ;
  input \P3_ByteEnable_reg[1]/NET0131  ;
  input \P3_ByteEnable_reg[2]/NET0131  ;
  input \P3_ByteEnable_reg[3]/NET0131  ;
  input \P3_CodeFetch_reg/NET0131  ;
  input \P3_DataWidth_reg[0]/NET0131  ;
  input \P3_DataWidth_reg[1]/NET0131  ;
  input \P3_EAX_reg[0]/NET0131  ;
  input \P3_EAX_reg[10]/NET0131  ;
  input \P3_EAX_reg[11]/NET0131  ;
  input \P3_EAX_reg[12]/NET0131  ;
  input \P3_EAX_reg[13]/NET0131  ;
  input \P3_EAX_reg[14]/NET0131  ;
  input \P3_EAX_reg[15]/NET0131  ;
  input \P3_EAX_reg[16]/NET0131  ;
  input \P3_EAX_reg[17]/NET0131  ;
  input \P3_EAX_reg[18]/NET0131  ;
  input \P3_EAX_reg[19]/NET0131  ;
  input \P3_EAX_reg[1]/NET0131  ;
  input \P3_EAX_reg[20]/NET0131  ;
  input \P3_EAX_reg[21]/NET0131  ;
  input \P3_EAX_reg[22]/NET0131  ;
  input \P3_EAX_reg[23]/NET0131  ;
  input \P3_EAX_reg[24]/NET0131  ;
  input \P3_EAX_reg[25]/NET0131  ;
  input \P3_EAX_reg[26]/NET0131  ;
  input \P3_EAX_reg[27]/NET0131  ;
  input \P3_EAX_reg[28]/NET0131  ;
  input \P3_EAX_reg[29]/NET0131  ;
  input \P3_EAX_reg[2]/NET0131  ;
  input \P3_EAX_reg[30]/NET0131  ;
  input \P3_EAX_reg[31]/NET0131  ;
  input \P3_EAX_reg[3]/NET0131  ;
  input \P3_EAX_reg[4]/NET0131  ;
  input \P3_EAX_reg[5]/NET0131  ;
  input \P3_EAX_reg[6]/NET0131  ;
  input \P3_EAX_reg[7]/NET0131  ;
  input \P3_EAX_reg[8]/NET0131  ;
  input \P3_EAX_reg[9]/NET0131  ;
  input \P3_EBX_reg[0]/NET0131  ;
  input \P3_EBX_reg[10]/NET0131  ;
  input \P3_EBX_reg[11]/NET0131  ;
  input \P3_EBX_reg[12]/NET0131  ;
  input \P3_EBX_reg[13]/NET0131  ;
  input \P3_EBX_reg[14]/NET0131  ;
  input \P3_EBX_reg[15]/NET0131  ;
  input \P3_EBX_reg[16]/NET0131  ;
  input \P3_EBX_reg[17]/NET0131  ;
  input \P3_EBX_reg[18]/NET0131  ;
  input \P3_EBX_reg[19]/NET0131  ;
  input \P3_EBX_reg[1]/NET0131  ;
  input \P3_EBX_reg[20]/NET0131  ;
  input \P3_EBX_reg[21]/NET0131  ;
  input \P3_EBX_reg[22]/NET0131  ;
  input \P3_EBX_reg[23]/NET0131  ;
  input \P3_EBX_reg[24]/NET0131  ;
  input \P3_EBX_reg[25]/NET0131  ;
  input \P3_EBX_reg[26]/NET0131  ;
  input \P3_EBX_reg[27]/NET0131  ;
  input \P3_EBX_reg[28]/NET0131  ;
  input \P3_EBX_reg[29]/NET0131  ;
  input \P3_EBX_reg[2]/NET0131  ;
  input \P3_EBX_reg[30]/NET0131  ;
  input \P3_EBX_reg[31]/NET0131  ;
  input \P3_EBX_reg[3]/NET0131  ;
  input \P3_EBX_reg[4]/NET0131  ;
  input \P3_EBX_reg[5]/NET0131  ;
  input \P3_EBX_reg[6]/NET0131  ;
  input \P3_EBX_reg[7]/NET0131  ;
  input \P3_EBX_reg[8]/NET0131  ;
  input \P3_EBX_reg[9]/NET0131  ;
  input \P3_Flush_reg/NET0131  ;
  input \P3_InstAddrPointer_reg[0]/NET0131  ;
  input \P3_InstAddrPointer_reg[10]/NET0131  ;
  input \P3_InstAddrPointer_reg[11]/NET0131  ;
  input \P3_InstAddrPointer_reg[12]/NET0131  ;
  input \P3_InstAddrPointer_reg[13]/NET0131  ;
  input \P3_InstAddrPointer_reg[14]/NET0131  ;
  input \P3_InstAddrPointer_reg[15]/NET0131  ;
  input \P3_InstAddrPointer_reg[16]/NET0131  ;
  input \P3_InstAddrPointer_reg[17]/NET0131  ;
  input \P3_InstAddrPointer_reg[18]/NET0131  ;
  input \P3_InstAddrPointer_reg[19]/NET0131  ;
  input \P3_InstAddrPointer_reg[1]/NET0131  ;
  input \P3_InstAddrPointer_reg[20]/NET0131  ;
  input \P3_InstAddrPointer_reg[21]/NET0131  ;
  input \P3_InstAddrPointer_reg[22]/NET0131  ;
  input \P3_InstAddrPointer_reg[23]/NET0131  ;
  input \P3_InstAddrPointer_reg[24]/NET0131  ;
  input \P3_InstAddrPointer_reg[25]/NET0131  ;
  input \P3_InstAddrPointer_reg[26]/NET0131  ;
  input \P3_InstAddrPointer_reg[27]/NET0131  ;
  input \P3_InstAddrPointer_reg[28]/NET0131  ;
  input \P3_InstAddrPointer_reg[29]/NET0131  ;
  input \P3_InstAddrPointer_reg[2]/NET0131  ;
  input \P3_InstAddrPointer_reg[30]/NET0131  ;
  input \P3_InstAddrPointer_reg[31]/NET0131  ;
  input \P3_InstAddrPointer_reg[3]/NET0131  ;
  input \P3_InstAddrPointer_reg[4]/NET0131  ;
  input \P3_InstAddrPointer_reg[5]/NET0131  ;
  input \P3_InstAddrPointer_reg[6]/NET0131  ;
  input \P3_InstAddrPointer_reg[7]/NET0131  ;
  input \P3_InstAddrPointer_reg[8]/NET0131  ;
  input \P3_InstAddrPointer_reg[9]/NET0131  ;
  input \P3_InstQueueRd_Addr_reg[0]/NET0131  ;
  input \P3_InstQueueRd_Addr_reg[1]/NET0131  ;
  input \P3_InstQueueRd_Addr_reg[2]/NET0131  ;
  input \P3_InstQueueRd_Addr_reg[3]/NET0131  ;
  input \P3_InstQueueWr_Addr_reg[0]/NET0131  ;
  input \P3_InstQueueWr_Addr_reg[1]/NET0131  ;
  input \P3_InstQueueWr_Addr_reg[2]/NET0131  ;
  input \P3_InstQueueWr_Addr_reg[3]/NET0131  ;
  input \P3_InstQueue_reg[0][0]/NET0131  ;
  input \P3_InstQueue_reg[0][1]/NET0131  ;
  input \P3_InstQueue_reg[0][2]/NET0131  ;
  input \P3_InstQueue_reg[0][3]/NET0131  ;
  input \P3_InstQueue_reg[0][4]/NET0131  ;
  input \P3_InstQueue_reg[0][5]/NET0131  ;
  input \P3_InstQueue_reg[0][6]/NET0131  ;
  input \P3_InstQueue_reg[0][7]/NET0131  ;
  input \P3_InstQueue_reg[10][0]/NET0131  ;
  input \P3_InstQueue_reg[10][1]/NET0131  ;
  input \P3_InstQueue_reg[10][2]/NET0131  ;
  input \P3_InstQueue_reg[10][3]/NET0131  ;
  input \P3_InstQueue_reg[10][4]/NET0131  ;
  input \P3_InstQueue_reg[10][5]/NET0131  ;
  input \P3_InstQueue_reg[10][6]/NET0131  ;
  input \P3_InstQueue_reg[10][7]/NET0131  ;
  input \P3_InstQueue_reg[11][0]/NET0131  ;
  input \P3_InstQueue_reg[11][1]/NET0131  ;
  input \P3_InstQueue_reg[11][2]/NET0131  ;
  input \P3_InstQueue_reg[11][3]/NET0131  ;
  input \P3_InstQueue_reg[11][4]/NET0131  ;
  input \P3_InstQueue_reg[11][5]/NET0131  ;
  input \P3_InstQueue_reg[11][6]/NET0131  ;
  input \P3_InstQueue_reg[11][7]/NET0131  ;
  input \P3_InstQueue_reg[12][0]/NET0131  ;
  input \P3_InstQueue_reg[12][1]/NET0131  ;
  input \P3_InstQueue_reg[12][2]/NET0131  ;
  input \P3_InstQueue_reg[12][3]/NET0131  ;
  input \P3_InstQueue_reg[12][4]/NET0131  ;
  input \P3_InstQueue_reg[12][5]/NET0131  ;
  input \P3_InstQueue_reg[12][6]/NET0131  ;
  input \P3_InstQueue_reg[12][7]/NET0131  ;
  input \P3_InstQueue_reg[13][0]/NET0131  ;
  input \P3_InstQueue_reg[13][1]/NET0131  ;
  input \P3_InstQueue_reg[13][2]/NET0131  ;
  input \P3_InstQueue_reg[13][3]/NET0131  ;
  input \P3_InstQueue_reg[13][4]/NET0131  ;
  input \P3_InstQueue_reg[13][5]/NET0131  ;
  input \P3_InstQueue_reg[13][6]/NET0131  ;
  input \P3_InstQueue_reg[13][7]/NET0131  ;
  input \P3_InstQueue_reg[14][0]/NET0131  ;
  input \P3_InstQueue_reg[14][1]/NET0131  ;
  input \P3_InstQueue_reg[14][2]/NET0131  ;
  input \P3_InstQueue_reg[14][3]/NET0131  ;
  input \P3_InstQueue_reg[14][4]/NET0131  ;
  input \P3_InstQueue_reg[14][5]/NET0131  ;
  input \P3_InstQueue_reg[14][6]/NET0131  ;
  input \P3_InstQueue_reg[14][7]/NET0131  ;
  input \P3_InstQueue_reg[15][0]/NET0131  ;
  input \P3_InstQueue_reg[15][1]/NET0131  ;
  input \P3_InstQueue_reg[15][2]/NET0131  ;
  input \P3_InstQueue_reg[15][3]/NET0131  ;
  input \P3_InstQueue_reg[15][4]/NET0131  ;
  input \P3_InstQueue_reg[15][5]/NET0131  ;
  input \P3_InstQueue_reg[15][6]/NET0131  ;
  input \P3_InstQueue_reg[15][7]/NET0131  ;
  input \P3_InstQueue_reg[1][0]/NET0131  ;
  input \P3_InstQueue_reg[1][1]/NET0131  ;
  input \P3_InstQueue_reg[1][2]/NET0131  ;
  input \P3_InstQueue_reg[1][3]/NET0131  ;
  input \P3_InstQueue_reg[1][4]/NET0131  ;
  input \P3_InstQueue_reg[1][5]/NET0131  ;
  input \P3_InstQueue_reg[1][6]/NET0131  ;
  input \P3_InstQueue_reg[1][7]/NET0131  ;
  input \P3_InstQueue_reg[2][0]/NET0131  ;
  input \P3_InstQueue_reg[2][1]/NET0131  ;
  input \P3_InstQueue_reg[2][2]/NET0131  ;
  input \P3_InstQueue_reg[2][3]/NET0131  ;
  input \P3_InstQueue_reg[2][4]/NET0131  ;
  input \P3_InstQueue_reg[2][5]/NET0131  ;
  input \P3_InstQueue_reg[2][6]/NET0131  ;
  input \P3_InstQueue_reg[2][7]/NET0131  ;
  input \P3_InstQueue_reg[3][0]/NET0131  ;
  input \P3_InstQueue_reg[3][1]/NET0131  ;
  input \P3_InstQueue_reg[3][2]/NET0131  ;
  input \P3_InstQueue_reg[3][3]/NET0131  ;
  input \P3_InstQueue_reg[3][4]/NET0131  ;
  input \P3_InstQueue_reg[3][5]/NET0131  ;
  input \P3_InstQueue_reg[3][6]/NET0131  ;
  input \P3_InstQueue_reg[3][7]/NET0131  ;
  input \P3_InstQueue_reg[4][0]/NET0131  ;
  input \P3_InstQueue_reg[4][1]/NET0131  ;
  input \P3_InstQueue_reg[4][2]/NET0131  ;
  input \P3_InstQueue_reg[4][3]/NET0131  ;
  input \P3_InstQueue_reg[4][4]/NET0131  ;
  input \P3_InstQueue_reg[4][5]/NET0131  ;
  input \P3_InstQueue_reg[4][6]/NET0131  ;
  input \P3_InstQueue_reg[4][7]/NET0131  ;
  input \P3_InstQueue_reg[5][0]/NET0131  ;
  input \P3_InstQueue_reg[5][1]/NET0131  ;
  input \P3_InstQueue_reg[5][2]/NET0131  ;
  input \P3_InstQueue_reg[5][3]/NET0131  ;
  input \P3_InstQueue_reg[5][4]/NET0131  ;
  input \P3_InstQueue_reg[5][5]/NET0131  ;
  input \P3_InstQueue_reg[5][6]/NET0131  ;
  input \P3_InstQueue_reg[5][7]/NET0131  ;
  input \P3_InstQueue_reg[6][0]/NET0131  ;
  input \P3_InstQueue_reg[6][1]/NET0131  ;
  input \P3_InstQueue_reg[6][2]/NET0131  ;
  input \P3_InstQueue_reg[6][3]/NET0131  ;
  input \P3_InstQueue_reg[6][4]/NET0131  ;
  input \P3_InstQueue_reg[6][5]/NET0131  ;
  input \P3_InstQueue_reg[6][6]/NET0131  ;
  input \P3_InstQueue_reg[6][7]/NET0131  ;
  input \P3_InstQueue_reg[7][0]/NET0131  ;
  input \P3_InstQueue_reg[7][1]/NET0131  ;
  input \P3_InstQueue_reg[7][2]/NET0131  ;
  input \P3_InstQueue_reg[7][3]/NET0131  ;
  input \P3_InstQueue_reg[7][4]/NET0131  ;
  input \P3_InstQueue_reg[7][5]/NET0131  ;
  input \P3_InstQueue_reg[7][6]/NET0131  ;
  input \P3_InstQueue_reg[7][7]/NET0131  ;
  input \P3_InstQueue_reg[8][0]/NET0131  ;
  input \P3_InstQueue_reg[8][1]/NET0131  ;
  input \P3_InstQueue_reg[8][2]/NET0131  ;
  input \P3_InstQueue_reg[8][3]/NET0131  ;
  input \P3_InstQueue_reg[8][4]/NET0131  ;
  input \P3_InstQueue_reg[8][5]/NET0131  ;
  input \P3_InstQueue_reg[8][6]/NET0131  ;
  input \P3_InstQueue_reg[8][7]/NET0131  ;
  input \P3_InstQueue_reg[9][0]/NET0131  ;
  input \P3_InstQueue_reg[9][1]/NET0131  ;
  input \P3_InstQueue_reg[9][2]/NET0131  ;
  input \P3_InstQueue_reg[9][3]/NET0131  ;
  input \P3_InstQueue_reg[9][4]/NET0131  ;
  input \P3_InstQueue_reg[9][5]/NET0131  ;
  input \P3_InstQueue_reg[9][6]/NET0131  ;
  input \P3_InstQueue_reg[9][7]/NET0131  ;
  input \P3_MemoryFetch_reg/NET0131  ;
  input \P3_More_reg/NET0131  ;
  input \P3_PhyAddrPointer_reg[0]/NET0131  ;
  input \P3_PhyAddrPointer_reg[10]/NET0131  ;
  input \P3_PhyAddrPointer_reg[11]/NET0131  ;
  input \P3_PhyAddrPointer_reg[12]/NET0131  ;
  input \P3_PhyAddrPointer_reg[13]/NET0131  ;
  input \P3_PhyAddrPointer_reg[14]/NET0131  ;
  input \P3_PhyAddrPointer_reg[15]/NET0131  ;
  input \P3_PhyAddrPointer_reg[16]/NET0131  ;
  input \P3_PhyAddrPointer_reg[17]/NET0131  ;
  input \P3_PhyAddrPointer_reg[18]/NET0131  ;
  input \P3_PhyAddrPointer_reg[19]/NET0131  ;
  input \P3_PhyAddrPointer_reg[1]/NET0131  ;
  input \P3_PhyAddrPointer_reg[20]/NET0131  ;
  input \P3_PhyAddrPointer_reg[21]/NET0131  ;
  input \P3_PhyAddrPointer_reg[22]/NET0131  ;
  input \P3_PhyAddrPointer_reg[23]/NET0131  ;
  input \P3_PhyAddrPointer_reg[24]/NET0131  ;
  input \P3_PhyAddrPointer_reg[25]/NET0131  ;
  input \P3_PhyAddrPointer_reg[26]/NET0131  ;
  input \P3_PhyAddrPointer_reg[27]/NET0131  ;
  input \P3_PhyAddrPointer_reg[28]/NET0131  ;
  input \P3_PhyAddrPointer_reg[29]/NET0131  ;
  input \P3_PhyAddrPointer_reg[2]/NET0131  ;
  input \P3_PhyAddrPointer_reg[30]/NET0131  ;
  input \P3_PhyAddrPointer_reg[31]/NET0131  ;
  input \P3_PhyAddrPointer_reg[3]/NET0131  ;
  input \P3_PhyAddrPointer_reg[4]/NET0131  ;
  input \P3_PhyAddrPointer_reg[5]/NET0131  ;
  input \P3_PhyAddrPointer_reg[6]/NET0131  ;
  input \P3_PhyAddrPointer_reg[7]/NET0131  ;
  input \P3_PhyAddrPointer_reg[8]/NET0131  ;
  input \P3_PhyAddrPointer_reg[9]/NET0131  ;
  input \P3_ReadRequest_reg/NET0131  ;
  input \P3_RequestPending_reg/NET0131  ;
  input \P3_State2_reg[0]/NET0131  ;
  input \P3_State2_reg[1]/NET0131  ;
  input \P3_State2_reg[2]/NET0131  ;
  input \P3_State2_reg[3]/NET0131  ;
  input \P3_State_reg[0]/NET0131  ;
  input \P3_State_reg[1]/NET0131  ;
  input \P3_State_reg[2]/NET0131  ;
  input \P3_lWord_reg[0]/NET0131  ;
  input \P3_lWord_reg[10]/NET0131  ;
  input \P3_lWord_reg[11]/NET0131  ;
  input \P3_lWord_reg[12]/NET0131  ;
  input \P3_lWord_reg[13]/NET0131  ;
  input \P3_lWord_reg[14]/NET0131  ;
  input \P3_lWord_reg[15]/NET0131  ;
  input \P3_lWord_reg[1]/NET0131  ;
  input \P3_lWord_reg[2]/NET0131  ;
  input \P3_lWord_reg[3]/NET0131  ;
  input \P3_lWord_reg[4]/NET0131  ;
  input \P3_lWord_reg[5]/NET0131  ;
  input \P3_lWord_reg[6]/NET0131  ;
  input \P3_lWord_reg[7]/NET0131  ;
  input \P3_lWord_reg[8]/NET0131  ;
  input \P3_lWord_reg[9]/NET0131  ;
  input \P3_rEIP_reg[0]/NET0131  ;
  input \P3_rEIP_reg[10]/NET0131  ;
  input \P3_rEIP_reg[11]/NET0131  ;
  input \P3_rEIP_reg[12]/NET0131  ;
  input \P3_rEIP_reg[13]/NET0131  ;
  input \P3_rEIP_reg[14]/NET0131  ;
  input \P3_rEIP_reg[15]/NET0131  ;
  input \P3_rEIP_reg[16]/NET0131  ;
  input \P3_rEIP_reg[17]/NET0131  ;
  input \P3_rEIP_reg[18]/NET0131  ;
  input \P3_rEIP_reg[19]/NET0131  ;
  input \P3_rEIP_reg[1]/NET0131  ;
  input \P3_rEIP_reg[20]/NET0131  ;
  input \P3_rEIP_reg[21]/NET0131  ;
  input \P3_rEIP_reg[22]/NET0131  ;
  input \P3_rEIP_reg[23]/NET0131  ;
  input \P3_rEIP_reg[24]/NET0131  ;
  input \P3_rEIP_reg[25]/NET0131  ;
  input \P3_rEIP_reg[26]/NET0131  ;
  input \P3_rEIP_reg[27]/NET0131  ;
  input \P3_rEIP_reg[28]/NET0131  ;
  input \P3_rEIP_reg[29]/NET0131  ;
  input \P3_rEIP_reg[2]/NET0131  ;
  input \P3_rEIP_reg[30]/NET0131  ;
  input \P3_rEIP_reg[31]/NET0131  ;
  input \P3_rEIP_reg[3]/NET0131  ;
  input \P3_rEIP_reg[4]/NET0131  ;
  input \P3_rEIP_reg[5]/NET0131  ;
  input \P3_rEIP_reg[6]/NET0131  ;
  input \P3_rEIP_reg[7]/NET0131  ;
  input \P3_rEIP_reg[8]/NET0131  ;
  input \P3_rEIP_reg[9]/NET0131  ;
  input \P3_uWord_reg[0]/NET0131  ;
  input \P3_uWord_reg[10]/NET0131  ;
  input \P3_uWord_reg[11]/NET0131  ;
  input \P3_uWord_reg[12]/NET0131  ;
  input \P3_uWord_reg[13]/NET0131  ;
  input \P3_uWord_reg[14]/NET0131  ;
  input \P3_uWord_reg[1]/NET0131  ;
  input \P3_uWord_reg[2]/NET0131  ;
  input \P3_uWord_reg[3]/NET0131  ;
  input \P3_uWord_reg[4]/NET0131  ;
  input \P3_uWord_reg[5]/NET0131  ;
  input \P3_uWord_reg[6]/NET0131  ;
  input \P3_uWord_reg[7]/NET0131  ;
  input \P3_uWord_reg[8]/NET0131  ;
  input \P3_uWord_reg[9]/NET0131  ;
  input \address1[0]_pad  ;
  input \address1[10]_pad  ;
  input \address1[11]_pad  ;
  input \address1[12]_pad  ;
  input \address1[13]_pad  ;
  input \address1[14]_pad  ;
  input \address1[15]_pad  ;
  input \address1[16]_pad  ;
  input \address1[17]_pad  ;
  input \address1[18]_pad  ;
  input \address1[19]_pad  ;
  input \address1[1]_pad  ;
  input \address1[20]_pad  ;
  input \address1[21]_pad  ;
  input \address1[22]_pad  ;
  input \address1[23]_pad  ;
  input \address1[24]_pad  ;
  input \address1[25]_pad  ;
  input \address1[26]_pad  ;
  input \address1[27]_pad  ;
  input \address1[28]_pad  ;
  input \address1[29]_pad  ;
  input \address1[2]_pad  ;
  input \address1[3]_pad  ;
  input \address1[4]_pad  ;
  input \address1[5]_pad  ;
  input \address1[6]_pad  ;
  input \address1[7]_pad  ;
  input \address1[8]_pad  ;
  input \address1[9]_pad  ;
  input \ast1_pad  ;
  input \ast2_pad  ;
  input \bs16_pad  ;
  input \buf1_reg[0]/NET0131  ;
  input \buf1_reg[10]/NET0131  ;
  input \buf1_reg[11]/NET0131  ;
  input \buf1_reg[12]/NET0131  ;
  input \buf1_reg[13]/NET0131  ;
  input \buf1_reg[14]/NET0131  ;
  input \buf1_reg[15]/NET0131  ;
  input \buf1_reg[16]/NET0131  ;
  input \buf1_reg[17]/NET0131  ;
  input \buf1_reg[18]/NET0131  ;
  input \buf1_reg[19]/NET0131  ;
  input \buf1_reg[1]/NET0131  ;
  input \buf1_reg[20]/NET0131  ;
  input \buf1_reg[21]/NET0131  ;
  input \buf1_reg[22]/NET0131  ;
  input \buf1_reg[23]/NET0131  ;
  input \buf1_reg[24]/NET0131  ;
  input \buf1_reg[25]/NET0131  ;
  input \buf1_reg[26]/NET0131  ;
  input \buf1_reg[27]/NET0131  ;
  input \buf1_reg[28]/NET0131  ;
  input \buf1_reg[29]/NET0131  ;
  input \buf1_reg[2]/NET0131  ;
  input \buf1_reg[30]/NET0131  ;
  input \buf1_reg[3]/NET0131  ;
  input \buf1_reg[4]/NET0131  ;
  input \buf1_reg[5]/NET0131  ;
  input \buf1_reg[6]/NET0131  ;
  input \buf1_reg[7]/NET0131  ;
  input \buf1_reg[8]/NET0131  ;
  input \buf1_reg[9]/NET0131  ;
  input \buf2_reg[0]/NET0131  ;
  input \buf2_reg[10]/NET0131  ;
  input \buf2_reg[11]/NET0131  ;
  input \buf2_reg[12]/NET0131  ;
  input \buf2_reg[13]/NET0131  ;
  input \buf2_reg[14]/NET0131  ;
  input \buf2_reg[15]/NET0131  ;
  input \buf2_reg[16]/NET0131  ;
  input \buf2_reg[17]/NET0131  ;
  input \buf2_reg[18]/NET0131  ;
  input \buf2_reg[19]/NET0131  ;
  input \buf2_reg[1]/NET0131  ;
  input \buf2_reg[20]/NET0131  ;
  input \buf2_reg[21]/NET0131  ;
  input \buf2_reg[22]/NET0131  ;
  input \buf2_reg[23]/NET0131  ;
  input \buf2_reg[24]/NET0131  ;
  input \buf2_reg[25]/NET0131  ;
  input \buf2_reg[26]/NET0131  ;
  input \buf2_reg[27]/NET0131  ;
  input \buf2_reg[28]/NET0131  ;
  input \buf2_reg[29]/NET0131  ;
  input \buf2_reg[2]/NET0131  ;
  input \buf2_reg[30]/NET0131  ;
  input \buf2_reg[3]/NET0131  ;
  input \buf2_reg[4]/NET0131  ;
  input \buf2_reg[5]/NET0131  ;
  input \buf2_reg[6]/NET0131  ;
  input \buf2_reg[7]/NET0131  ;
  input \buf2_reg[8]/NET0131  ;
  input \buf2_reg[9]/NET0131  ;
  input \datai[0]_pad  ;
  input \datai[10]_pad  ;
  input \datai[11]_pad  ;
  input \datai[12]_pad  ;
  input \datai[13]_pad  ;
  input \datai[14]_pad  ;
  input \datai[15]_pad  ;
  input \datai[16]_pad  ;
  input \datai[17]_pad  ;
  input \datai[18]_pad  ;
  input \datai[19]_pad  ;
  input \datai[1]_pad  ;
  input \datai[20]_pad  ;
  input \datai[21]_pad  ;
  input \datai[22]_pad  ;
  input \datai[23]_pad  ;
  input \datai[24]_pad  ;
  input \datai[25]_pad  ;
  input \datai[26]_pad  ;
  input \datai[27]_pad  ;
  input \datai[28]_pad  ;
  input \datai[29]_pad  ;
  input \datai[2]_pad  ;
  input \datai[30]_pad  ;
  input \datai[31]_pad  ;
  input \datai[3]_pad  ;
  input \datai[4]_pad  ;
  input \datai[5]_pad  ;
  input \datai[6]_pad  ;
  input \datai[7]_pad  ;
  input \datai[8]_pad  ;
  input \datai[9]_pad  ;
  input \datao[0]_pad  ;
  input \datao[10]_pad  ;
  input \datao[11]_pad  ;
  input \datao[12]_pad  ;
  input \datao[13]_pad  ;
  input \datao[14]_pad  ;
  input \datao[15]_pad  ;
  input \datao[16]_pad  ;
  input \datao[17]_pad  ;
  input \datao[18]_pad  ;
  input \datao[19]_pad  ;
  input \datao[1]_pad  ;
  input \datao[20]_pad  ;
  input \datao[21]_pad  ;
  input \datao[22]_pad  ;
  input \datao[23]_pad  ;
  input \datao[24]_pad  ;
  input \datao[25]_pad  ;
  input \datao[26]_pad  ;
  input \datao[27]_pad  ;
  input \datao[28]_pad  ;
  input \datao[29]_pad  ;
  input \datao[2]_pad  ;
  input \datao[30]_pad  ;
  input \datao[3]_pad  ;
  input \datao[4]_pad  ;
  input \datao[5]_pad  ;
  input \datao[6]_pad  ;
  input \datao[7]_pad  ;
  input \datao[8]_pad  ;
  input \datao[9]_pad  ;
  input dc_pad ;
  input hold_pad ;
  input mio_pad ;
  input na_pad ;
  input \ready11_reg/NET0131  ;
  input \ready12_reg/NET0131  ;
  input \ready1_pad  ;
  input \ready21_reg/NET0131  ;
  input \ready22_reg/NET0131  ;
  input \ready2_pad  ;
  input wr_pad ;
  output \_al_n0  ;
  output \_al_n1  ;
  output \address2[0]_pad  ;
  output \address2[10]_pad  ;
  output \address2[11]_pad  ;
  output \address2[12]_pad  ;
  output \address2[13]_pad  ;
  output \address2[14]_pad  ;
  output \address2[15]_pad  ;
  output \address2[16]_pad  ;
  output \address2[17]_pad  ;
  output \address2[18]_pad  ;
  output \address2[19]_pad  ;
  output \address2[1]_pad  ;
  output \address2[20]_pad  ;
  output \address2[21]_pad  ;
  output \address2[22]_pad  ;
  output \address2[23]_pad  ;
  output \address2[24]_pad  ;
  output \address2[25]_pad  ;
  output \address2[26]_pad  ;
  output \address2[27]_pad  ;
  output \address2[28]_pad  ;
  output \address2[29]_pad  ;
  output \address2[2]_pad  ;
  output \address2[3]_pad  ;
  output \address2[4]_pad  ;
  output \address2[5]_pad  ;
  output \address2[6]_pad  ;
  output \address2[7]_pad  ;
  output \address2[8]_pad  ;
  output \address2[9]_pad  ;
  output \g133468/_2_  ;
  output \g133469/_2_  ;
  output \g133470/_2_  ;
  output \g133475/_0_  ;
  output \g133476/_2_  ;
  output \g133515/_0_  ;
  output \g133516/_0_  ;
  output \g133517/_0_  ;
  output \g133518/_0_  ;
  output \g133523/_0_  ;
  output \g133524/_0_  ;
  output \g133528/_0_  ;
  output \g133529/_0_  ;
  output \g133531/_0_  ;
  output \g133532/_0_  ;
  output \g133533/_0_  ;
  output \g133534/_0_  ;
  output \g133535/_0_  ;
  output \g133536/_0_  ;
  output \g133537/_0_  ;
  output \g133538/_0_  ;
  output \g133539/_0_  ;
  output \g133540/_0_  ;
  output \g133541/_0_  ;
  output \g133542/_0_  ;
  output \g133543/_0_  ;
  output \g133544/_0_  ;
  output \g133545/_0_  ;
  output \g133546/_0_  ;
  output \g133547/_0_  ;
  output \g133548/_0_  ;
  output \g133549/_0_  ;
  output \g133550/_0_  ;
  output \g133551/_0_  ;
  output \g133552/_0_  ;
  output \g133553/_0_  ;
  output \g133554/_0_  ;
  output \g133555/_0_  ;
  output \g133556/_0_  ;
  output \g133557/_0_  ;
  output \g133558/_0_  ;
  output \g133559/_0_  ;
  output \g133560/_0_  ;
  output \g133561/_0_  ;
  output \g133566/_0_  ;
  output \g133619/_0_  ;
  output \g133659/_0_  ;
  output \g133660/_0_  ;
  output \g133662/_0_  ;
  output \g133663/_0_  ;
  output \g133664/_0_  ;
  output \g133665/_0_  ;
  output \g133666/_0_  ;
  output \g133667/_0_  ;
  output \g133668/_0_  ;
  output \g133669/_0_  ;
  output \g133670/_0_  ;
  output \g133671/_0_  ;
  output \g133672/_0_  ;
  output \g133673/_0_  ;
  output \g133674/_0_  ;
  output \g133675/_0_  ;
  output \g133676/_0_  ;
  output \g133677/_0_  ;
  output \g133678/_0_  ;
  output \g133679/_0_  ;
  output \g133680/_0_  ;
  output \g133681/_0_  ;
  output \g133682/_0_  ;
  output \g133683/_0_  ;
  output \g133684/_0_  ;
  output \g133685/_0_  ;
  output \g133686/_0_  ;
  output \g133687/_0_  ;
  output \g133688/_0_  ;
  output \g133689/_0_  ;
  output \g133690/_0_  ;
  output \g133691/_0_  ;
  output \g133694/_0_  ;
  output \g133697/_0_  ;
  output \g133702/_0_  ;
  output \g133703/_0_  ;
  output \g133756/_0_  ;
  output \g133792/_0_  ;
  output \g133793/_0_  ;
  output \g133794/_0_  ;
  output \g133796/_0_  ;
  output \g133797/_0_  ;
  output \g133798/_0_  ;
  output \g133799/_0_  ;
  output \g133800/_0_  ;
  output \g133801/_0_  ;
  output \g133802/_0_  ;
  output \g133803/_0_  ;
  output \g133804/_0_  ;
  output \g133806/_0_  ;
  output \g133807/_0_  ;
  output \g133808/_0_  ;
  output \g133812/_0_  ;
  output \g133813/_0_  ;
  output \g133814/_0_  ;
  output \g133817/_0_  ;
  output \g133821/_0_  ;
  output \g133824/_0_  ;
  output \g133826/_0_  ;
  output \g133828/_0_  ;
  output \g133864/_0_  ;
  output \g133865/_0_  ;
  output \g133867/_0_  ;
  output \g133868/_0_  ;
  output \g133869/_0_  ;
  output \g133871/_0_  ;
  output \g133872/_0_  ;
  output \g133873/_0_  ;
  output \g133874/_0_  ;
  output \g133875/_0_  ;
  output \g133876/_0_  ;
  output \g133877/_0_  ;
  output \g133878/_0_  ;
  output \g133879/_0_  ;
  output \g133881/_0_  ;
  output \g133882/_0_  ;
  output \g133883/_0_  ;
  output \g133884/_0_  ;
  output \g133885/_0_  ;
  output \g133886/_0_  ;
  output \g133887/_0_  ;
  output \g133888/_0_  ;
  output \g133889/_0_  ;
  output \g133890/_0_  ;
  output \g133891/_0_  ;
  output \g133892/_0_  ;
  output \g133893/_0_  ;
  output \g133894/_0_  ;
  output \g133895/_0_  ;
  output \g133896/_0_  ;
  output \g133897/_0_  ;
  output \g133898/_0_  ;
  output \g133910/_0_  ;
  output \g133911/_0_  ;
  output \g133912/_0_  ;
  output \g133915/_0_  ;
  output \g133917/_0_  ;
  output \g133929/_0_  ;
  output \g134014/_0_  ;
  output \g134040/_0_  ;
  output \g134041/_0_  ;
  output \g134042/_0_  ;
  output \g134043/_0_  ;
  output \g134044/_0_  ;
  output \g134045/_0_  ;
  output \g134046/_0_  ;
  output \g134047/_0_  ;
  output \g134048/_0_  ;
  output \g134049/_0_  ;
  output \g134050/_0_  ;
  output \g134051/_0_  ;
  output \g134052/_0_  ;
  output \g134053/_0_  ;
  output \g134054/_0_  ;
  output \g134056/_0_  ;
  output \g134059/_0_  ;
  output \g134064/_0_  ;
  output \g134067/_0_  ;
  output \g134068/_0_  ;
  output \g134069/_0_  ;
  output \g134070/_0_  ;
  output \g134071/_0_  ;
  output \g134073/_0_  ;
  output \g134076/_0_  ;
  output \g134131/_0_  ;
  output \g134132/_0_  ;
  output \g134156/_0_  ;
  output \g134157/_0_  ;
  output \g134158/_0_  ;
  output \g134159/_0_  ;
  output \g134163/_0_  ;
  output \g134164/_0_  ;
  output \g134165/_0_  ;
  output \g134166/_0_  ;
  output \g134167/_0_  ;
  output \g134168/_0_  ;
  output \g134169/_0_  ;
  output \g134170/_0_  ;
  output \g134171/_0_  ;
  output \g134172/_0_  ;
  output \g134173/_0_  ;
  output \g134174/_0_  ;
  output \g134176/_0_  ;
  output \g134177/_0_  ;
  output \g134178/_0_  ;
  output \g134179/_0_  ;
  output \g134181/_0_  ;
  output \g134183/_0_  ;
  output \g134184/_0_  ;
  output \g134185/_0_  ;
  output \g134186/_0_  ;
  output \g134187/_0_  ;
  output \g134188/_0_  ;
  output \g134189/_0_  ;
  output \g134190/_0_  ;
  output \g134191/_0_  ;
  output \g134194/_0_  ;
  output \g134202/_0_  ;
  output \g134207/_0_  ;
  output \g134214/_0_  ;
  output \g134216/_0_  ;
  output \g134226/_0_  ;
  output \g134228/_0_  ;
  output \g134360/_0_  ;
  output \g134383/_0_  ;
  output \g134412/_0_  ;
  output \g134413/_0_  ;
  output \g134419/_0_  ;
  output \g134420/_0_  ;
  output \g134421/_0_  ;
  output \g134422/_0_  ;
  output \g134423/_0_  ;
  output \g134424/_0_  ;
  output \g134426/_0_  ;
  output \g134429/_0_  ;
  output \g134431/_0_  ;
  output \g134433/_0_  ;
  output \g134434/_0_  ;
  output \g134435/_0_  ;
  output \g134436/_0_  ;
  output \g134438/_0_  ;
  output \g134439/_0_  ;
  output \g134441/_0_  ;
  output \g134442/_0_  ;
  output \g134443/_0_  ;
  output \g134445/_0_  ;
  output \g134446/_0_  ;
  output \g134447/_0_  ;
  output \g134448/_0_  ;
  output \g134449/_0_  ;
  output \g134450/_0_  ;
  output \g134451/_0_  ;
  output \g134453/_0_  ;
  output \g134454/_0_  ;
  output \g134455/_0_  ;
  output \g134457/_0_  ;
  output \g134458/_0_  ;
  output \g134459/_0_  ;
  output \g134460/_0_  ;
  output \g134469/_0_  ;
  output \g134470/_0_  ;
  output \g134471/_0_  ;
  output \g134472/_0_  ;
  output \g134479/_0_  ;
  output \g134480/_0_  ;
  output \g134481/_0_  ;
  output \g134482/_0_  ;
  output \g134490/_0_  ;
  output \g134491/_0_  ;
  output \g134496/_0_  ;
  output \g134506/_0_  ;
  output \g134508/_0_  ;
  output \g134579/_0_  ;
  output \g134603/_0_  ;
  output \g134604/_0_  ;
  output \g134605/_0_  ;
  output \g134606/_0_  ;
  output \g134607/_0_  ;
  output \g134608/_0_  ;
  output \g134609/_0_  ;
  output \g134610/_0_  ;
  output \g134611/_0_  ;
  output \g134612/_0_  ;
  output \g134613/_0_  ;
  output \g134614/_0_  ;
  output \g134615/_0_  ;
  output \g134616/_0_  ;
  output \g134617/_0_  ;
  output \g134618/_0_  ;
  output \g134619/_0_  ;
  output \g134620/_0_  ;
  output \g134621/_0_  ;
  output \g134632/_0_  ;
  output \g134633/_0_  ;
  output \g134636/_0_  ;
  output \g134637/_0_  ;
  output \g134638/_0_  ;
  output \g134639/_0_  ;
  output \g134645/_0_  ;
  output \g134646/_0_  ;
  output \g134648/_0_  ;
  output \g134649/_0_  ;
  output \g134650/_0_  ;
  output \g134651/_0_  ;
  output \g134652/_0_  ;
  output \g134656/_0_  ;
  output \g134657/_0_  ;
  output \g134658/_0_  ;
  output \g134664/_0_  ;
  output \g134665/_0_  ;
  output \g134671/_0_  ;
  output \g134672/_0_  ;
  output \g134686/_0_  ;
  output \g134687/_0_  ;
  output \g134735/_0_  ;
  output \g134908/_0_  ;
  output \g134909/_0_  ;
  output \g134910/_0_  ;
  output \g134920/_0_  ;
  output \g134921/_0_  ;
  output \g134922/_0_  ;
  output \g134923/_0_  ;
  output \g134925/_0_  ;
  output \g134926/_0_  ;
  output \g134928/_0_  ;
  output \g134929/_0_  ;
  output \g134933/_0_  ;
  output \g134934/_0_  ;
  output \g134935/_0_  ;
  output \g134936/_0_  ;
  output \g134937/_0_  ;
  output \g134938/_0_  ;
  output \g134940/_0_  ;
  output \g134941/_0_  ;
  output \g134943/_0_  ;
  output \g134945/_0_  ;
  output \g134946/_0_  ;
  output \g134947/_0_  ;
  output \g134948/_0_  ;
  output \g134949/_0_  ;
  output \g134950/_0_  ;
  output \g134959/_0_  ;
  output \g134960/_0_  ;
  output \g134961/_0_  ;
  output \g134979/_0_  ;
  output \g134980/_0_  ;
  output \g135054/_0_  ;
  output \g135061/_0_  ;
  output \g135072/_0_  ;
  output \g135100/_0_  ;
  output \g135127/_0_  ;
  output \g135128/_0_  ;
  output \g135129/_0_  ;
  output \g135130/_0_  ;
  output \g135132/_0_  ;
  output \g135133/_0_  ;
  output \g135134/_0_  ;
  output \g135135/_0_  ;
  output \g135136/_0_  ;
  output \g135137/_0_  ;
  output \g135138/_0_  ;
  output \g135139/_0_  ;
  output \g135140/_0_  ;
  output \g135141/_0_  ;
  output \g135142/_0_  ;
  output \g135145/_0_  ;
  output \g135146/_0_  ;
  output \g135151/_0_  ;
  output \g135154/_0_  ;
  output \g135155/_0_  ;
  output \g135158/_0_  ;
  output \g135163/_0_  ;
  output \g135164/_0_  ;
  output \g135165/_0_  ;
  output \g135192/_0_  ;
  output \g135197/_0_  ;
  output \g135217/_0_  ;
  output \g135225/_0_  ;
  output \g135231/_0_  ;
  output \g135272/_0_  ;
  output \g135290/_0_  ;
  output \g135291/_0_  ;
  output \g135293/_0_  ;
  output \g135294/_0_  ;
  output \g135295/_0_  ;
  output \g135296/_0_  ;
  output \g135297/_0_  ;
  output \g135412/_0_  ;
  output \g135437/_0_  ;
  output \g135438/_0_  ;
  output \g135443/_0_  ;
  output \g135444/_0_  ;
  output \g135445/_0_  ;
  output \g135446/_0_  ;
  output \g135447/_0_  ;
  output \g135448/_0_  ;
  output \g135449/_0_  ;
  output \g135450/_0_  ;
  output \g135451/_0_  ;
  output \g135452/_0_  ;
  output \g135454/_0_  ;
  output \g135455/_0_  ;
  output \g135456/_0_  ;
  output \g135457/_0_  ;
  output \g135458/_0_  ;
  output \g135463/_0_  ;
  output \g135466/_0_  ;
  output \g135473/_0_  ;
  output \g135481/_0_  ;
  output \g135497/_0_  ;
  output \g135503/_0_  ;
  output \g135505/_0_  ;
  output \g135506/_0_  ;
  output \g135557/_0_  ;
  output \g135558/_0_  ;
  output \g135569/_0_  ;
  output \g135570/_0_  ;
  output \g135571/_0_  ;
  output \g135572/_0_  ;
  output \g135573/_0_  ;
  output \g135575/_0_  ;
  output \g135578/_0_  ;
  output \g135754/_0_  ;
  output \g135755/_0_  ;
  output \g135756/_0_  ;
  output \g135767/_0_  ;
  output \g135768/_0_  ;
  output \g135769/_0_  ;
  output \g135777/_0_  ;
  output \g135778/_0_  ;
  output \g135779/_0_  ;
  output \g135872/_0_  ;
  output \g135873/_0_  ;
  output \g135875/_0_  ;
  output \g135877/_0_  ;
  output \g135878/_0_  ;
  output \g135879/_0_  ;
  output \g135880/_0_  ;
  output \g136087/_0_  ;
  output \g136118/_0_  ;
  output \g136119/_0_  ;
  output \g136120/_0_  ;
  output \g136121/_0_  ;
  output \g136122/_0_  ;
  output \g136123/_0_  ;
  output \g136124/_0_  ;
  output \g136125/_0_  ;
  output \g136126/_0_  ;
  output \g136127/_0_  ;
  output \g136128/_0_  ;
  output \g136129/_0_  ;
  output \g136130/_0_  ;
  output \g136131/_0_  ;
  output \g136132/_0_  ;
  output \g136133/_0_  ;
  output \g136172/_0_  ;
  output \g136173/_0_  ;
  output \g136174/_0_  ;
  output \g136175/_0_  ;
  output \g136177/_0_  ;
  output \g136178/_0_  ;
  output \g136242/_0_  ;
  output \g136243/_0_  ;
  output \g136244/_0_  ;
  output \g136246/_0_  ;
  output \g136248/_0_  ;
  output \g136249/_0_  ;
  output \g136250/_0_  ;
  output \g136251/_0_  ;
  output \g136252/_0_  ;
  output \g136253/_0_  ;
  output \g136254/_0_  ;
  output \g136255/_0_  ;
  output \g136256/_0_  ;
  output \g136257/_0_  ;
  output \g136258/_0_  ;
  output \g136259/_0_  ;
  output \g136260/_0_  ;
  output \g136261/_0_  ;
  output \g136262/_0_  ;
  output \g136263/_0_  ;
  output \g136264/_0_  ;
  output \g136265/_0_  ;
  output \g136266/_0_  ;
  output \g136267/_0_  ;
  output \g136268/_0_  ;
  output \g136269/_0_  ;
  output \g136270/_0_  ;
  output \g136271/_0_  ;
  output \g136272/_0_  ;
  output \g136273/_0_  ;
  output \g136274/_0_  ;
  output \g136275/_0_  ;
  output \g136276/_0_  ;
  output \g136277/_0_  ;
  output \g136279/_0_  ;
  output \g136280/_0_  ;
  output \g136281/_0_  ;
  output \g136282/_0_  ;
  output \g136283/_0_  ;
  output \g136285/_0_  ;
  output \g136286/_0_  ;
  output \g136287/_0_  ;
  output \g136288/_0_  ;
  output \g136289/_0_  ;
  output \g136290/_0_  ;
  output \g136291/_0_  ;
  output \g136292/_0_  ;
  output \g136293/_0_  ;
  output \g136295/_0_  ;
  output \g136467/_0_  ;
  output \g136468/_0_  ;
  output \g136469/_0_  ;
  output \g136470/_0_  ;
  output \g136472/_0_  ;
  output \g136473/_0_  ;
  output \g136474/_0_  ;
  output \g136476/_0_  ;
  output \g136479/_0_  ;
  output \g136480/_0_  ;
  output \g136481/_0_  ;
  output \g136482/_0_  ;
  output \g136483/_0_  ;
  output \g136484/_0_  ;
  output \g136485/_0_  ;
  output \g136486/_0_  ;
  output \g136528/_0_  ;
  output \g136529/_0_  ;
  output \g136530/_0_  ;
  output \g136531/_0_  ;
  output \g136532/_0_  ;
  output \g136533/_0_  ;
  output \g136534/_0_  ;
  output \g136535/_0_  ;
  output \g136536/_0_  ;
  output \g136537/_0_  ;
  output \g136538/_0_  ;
  output \g136539/_0_  ;
  output \g136540/_0_  ;
  output \g136541/_0_  ;
  output \g136542/_0_  ;
  output \g136543/_0_  ;
  output \g136544/_0_  ;
  output \g136545/_0_  ;
  output \g136546/_0_  ;
  output \g136547/_0_  ;
  output \g136548/_0_  ;
  output \g136549/_0_  ;
  output \g136550/_0_  ;
  output \g136551/_0_  ;
  output \g136552/_0_  ;
  output \g136553/_0_  ;
  output \g136554/_0_  ;
  output \g136555/_0_  ;
  output \g136556/_0_  ;
  output \g136557/_0_  ;
  output \g136558/_0_  ;
  output \g136559/_0_  ;
  output \g136560/_0_  ;
  output \g136561/_0_  ;
  output \g136562/_0_  ;
  output \g136563/_0_  ;
  output \g136564/_0_  ;
  output \g136565/_0_  ;
  output \g136566/_0_  ;
  output \g136567/_0_  ;
  output \g136568/_0_  ;
  output \g136570/_0_  ;
  output \g136571/_0_  ;
  output \g136572/_0_  ;
  output \g136573/_0_  ;
  output \g136574/_0_  ;
  output \g136575/_0_  ;
  output \g136576/_0_  ;
  output \g136577/_0_  ;
  output \g136578/_0_  ;
  output \g136579/_0_  ;
  output \g136580/_0_  ;
  output \g136582/_0_  ;
  output \g136583/_0_  ;
  output \g136584/_0_  ;
  output \g136585/_0_  ;
  output \g136586/_0_  ;
  output \g136587/_0_  ;
  output \g136588/_0_  ;
  output \g136589/_0_  ;
  output \g136590/_0_  ;
  output \g136591/_0_  ;
  output \g136592/_0_  ;
  output \g136593/_0_  ;
  output \g136594/_0_  ;
  output \g136595/_0_  ;
  output \g136596/_0_  ;
  output \g136597/_0_  ;
  output \g136598/_0_  ;
  output \g136599/_0_  ;
  output \g136600/_0_  ;
  output \g136601/_0_  ;
  output \g136602/_0_  ;
  output \g136603/_0_  ;
  output \g136604/_0_  ;
  output \g136605/_0_  ;
  output \g136606/_0_  ;
  output \g136607/_0_  ;
  output \g136609/_0_  ;
  output \g136610/_0_  ;
  output \g136611/_0_  ;
  output \g136616/_0_  ;
  output \g136617/_0_  ;
  output \g136618/_0_  ;
  output \g136619/_0_  ;
  output \g136626/_0_  ;
  output \g136628/_0_  ;
  output \g136646/_0_  ;
  output \g136649/_0_  ;
  output \g136662/_0_  ;
  output \g136666/_0_  ;
  output \g136695/_0_  ;
  output \g136696/_0_  ;
  output \g136699/_0_  ;
  output \g136762/_0_  ;
  output \g136763/_0_  ;
  output \g136764/_0_  ;
  output \g136765/_0_  ;
  output \g136768/_0_  ;
  output \g136769/_0_  ;
  output \g137051/_0_  ;
  output \g137052/_0_  ;
  output \g137053/_0_  ;
  output \g137054/_0_  ;
  output \g137055/_0_  ;
  output \g137056/_0_  ;
  output \g137057/_0_  ;
  output \g137060/_0_  ;
  output \g137061/_0_  ;
  output \g137063/_0_  ;
  output \g137064/_0_  ;
  output \g137065/_0_  ;
  output \g137067/_0_  ;
  output \g137069/_0_  ;
  output \g137072/_0_  ;
  output \g137073/_0_  ;
  output \g137075/_0_  ;
  output \g137111/_0_  ;
  output \g137122/_0_  ;
  output \g137133/_0_  ;
  output \g137134/_0_  ;
  output \g137135/_0_  ;
  output \g137136/_0_  ;
  output \g137137/_0_  ;
  output \g137138/_0_  ;
  output \g137144/_0_  ;
  output \g137145/_0_  ;
  output \g137146/_0_  ;
  output \g137149/_0_  ;
  output \g137234/_0_  ;
  output \g137237/_0_  ;
  output \g137238/_0_  ;
  output \g137294/_0_  ;
  output \g137295/_0_  ;
  output \g137296/_0_  ;
  output \g137297/_0_  ;
  output \g137298/_0_  ;
  output \g137299/_0_  ;
  output \g137300/_0_  ;
  output \g137301/_0_  ;
  output \g137302/_0_  ;
  output \g137303/_0_  ;
  output \g137304/_0_  ;
  output \g137305/_0_  ;
  output \g137306/_0_  ;
  output \g137307/_0_  ;
  output \g137308/_0_  ;
  output \g137309/_0_  ;
  output \g137310/_0_  ;
  output \g137311/_0_  ;
  output \g137312/_0_  ;
  output \g137313/_0_  ;
  output \g137314/_0_  ;
  output \g137315/_0_  ;
  output \g137316/_0_  ;
  output \g137317/_0_  ;
  output \g137318/_0_  ;
  output \g137319/_0_  ;
  output \g137320/_0_  ;
  output \g137321/_0_  ;
  output \g137322/_0_  ;
  output \g137323/_0_  ;
  output \g137324/_0_  ;
  output \g137325/_0_  ;
  output \g137327/_0_  ;
  output \g137328/_0_  ;
  output \g137329/_0_  ;
  output \g137330/_0_  ;
  output \g137331/_0_  ;
  output \g137332/_0_  ;
  output \g137333/_0_  ;
  output \g137334/_0_  ;
  output \g137335/_0_  ;
  output \g137336/_0_  ;
  output \g137337/_0_  ;
  output \g137338/_0_  ;
  output \g137339/_0_  ;
  output \g137340/_0_  ;
  output \g137341/_0_  ;
  output \g137342/_0_  ;
  output \g137343/_0_  ;
  output \g137344/_0_  ;
  output \g137345/_0_  ;
  output \g137346/_0_  ;
  output \g137347/_0_  ;
  output \g137349/_0_  ;
  output \g137350/_0_  ;
  output \g137351/_0_  ;
  output \g137352/_0_  ;
  output \g137353/_0_  ;
  output \g137354/_0_  ;
  output \g137448/_0_  ;
  output \g137483/_0_  ;
  output \g137484/_0_  ;
  output \g137485/_0_  ;
  output \g137486/_0_  ;
  output \g137487/_0_  ;
  output \g137488/_0_  ;
  output \g137491/_0_  ;
  output \g137492/_0_  ;
  output \g137493/_0_  ;
  output \g137494/_0_  ;
  output \g137495/_0_  ;
  output \g137496/_0_  ;
  output \g137497/_0_  ;
  output \g137499/_0_  ;
  output \g137501/_0_  ;
  output \g137502/_0_  ;
  output \g137503/_0_  ;
  output \g137504/_0_  ;
  output \g137505/_0_  ;
  output \g137506/_0_  ;
  output \g137507/_0_  ;
  output \g137508/_0_  ;
  output \g137509/_0_  ;
  output \g137511/_0_  ;
  output \g137512/_0_  ;
  output \g137513/_0_  ;
  output \g137514/_0_  ;
  output \g137515/_0_  ;
  output \g137516/_0_  ;
  output \g137517/_0_  ;
  output \g137519/_0_  ;
  output \g137520/_0_  ;
  output \g137521/_0_  ;
  output \g137524/_0_  ;
  output \g137541/_0_  ;
  output \g137547/_0_  ;
  output \g137554/_0_  ;
  output \g137559/_0_  ;
  output \g137566/_0_  ;
  output \g137571/_0_  ;
  output \g137778/_0_  ;
  output \g137782/_0_  ;
  output \g137783/_0_  ;
  output \g137784/_0_  ;
  output \g137785/_0_  ;
  output \g137786/_0_  ;
  output \g137820/_0_  ;
  output \g137821/_0_  ;
  output \g137822/_0_  ;
  output \g137823/_0_  ;
  output \g137824/_0_  ;
  output \g137825/_0_  ;
  output \g137826/_0_  ;
  output \g137827/_0_  ;
  output \g137828/_0_  ;
  output \g137829/_0_  ;
  output \g137830/_0_  ;
  output \g137831/_0_  ;
  output \g137832/_0_  ;
  output \g137833/_0_  ;
  output \g137834/_0_  ;
  output \g137835/_0_  ;
  output \g137836/_0_  ;
  output \g137837/_0_  ;
  output \g137838/_0_  ;
  output \g137839/_0_  ;
  output \g137840/_0_  ;
  output \g137841/_0_  ;
  output \g137842/_0_  ;
  output \g137843/_0_  ;
  output \g137844/_0_  ;
  output \g137845/_0_  ;
  output \g137846/_0_  ;
  output \g137847/_0_  ;
  output \g137848/_0_  ;
  output \g137849/_0_  ;
  output \g137850/_0_  ;
  output \g137851/_0_  ;
  output \g137852/_0_  ;
  output \g137853/_0_  ;
  output \g137854/_0_  ;
  output \g137855/_0_  ;
  output \g137856/_0_  ;
  output \g137857/_0_  ;
  output \g137858/_0_  ;
  output \g137859/_0_  ;
  output \g137860/_0_  ;
  output \g137861/_0_  ;
  output \g137862/_0_  ;
  output \g137863/_0_  ;
  output \g137864/_0_  ;
  output \g137865/_0_  ;
  output \g137866/_0_  ;
  output \g137867/_0_  ;
  output \g137868/_0_  ;
  output \g137869/_0_  ;
  output \g137870/_0_  ;
  output \g137871/_0_  ;
  output \g137872/_0_  ;
  output \g137873/_0_  ;
  output \g137874/_0_  ;
  output \g137875/_0_  ;
  output \g137876/_0_  ;
  output \g137877/_0_  ;
  output \g137878/_0_  ;
  output \g137879/_0_  ;
  output \g137880/_0_  ;
  output \g137881/_0_  ;
  output \g137882/_0_  ;
  output \g137883/_0_  ;
  output \g137884/_0_  ;
  output \g137885/_0_  ;
  output \g137886/_0_  ;
  output \g137887/_0_  ;
  output \g137888/_0_  ;
  output \g137889/_0_  ;
  output \g137890/_0_  ;
  output \g137891/_0_  ;
  output \g137892/_0_  ;
  output \g137893/_0_  ;
  output \g137894/_0_  ;
  output \g137895/_0_  ;
  output \g137896/_0_  ;
  output \g137897/_0_  ;
  output \g137898/_0_  ;
  output \g137899/_0_  ;
  output \g137900/_0_  ;
  output \g137901/_0_  ;
  output \g137902/_0_  ;
  output \g137903/_0_  ;
  output \g138338/_0_  ;
  output \g138340/_0_  ;
  output \g138341/_0_  ;
  output \g138346/_0_  ;
  output \g138347/_0_  ;
  output \g138375/_0_  ;
  output \g138395/_0_  ;
  output \g138396/_0_  ;
  output \g138397/_0_  ;
  output \g138398/_0_  ;
  output \g138400/_0_  ;
  output \g138401/_0_  ;
  output \g138402/_0_  ;
  output \g138403/_0_  ;
  output \g138404/_0_  ;
  output \g138405/_0_  ;
  output \g138406/_0_  ;
  output \g138407/_0_  ;
  output \g138408/_0_  ;
  output \g138409/_0_  ;
  output \g138410/_0_  ;
  output \g138411/_0_  ;
  output \g138412/_0_  ;
  output \g138419/_0_  ;
  output \g138420/_0_  ;
  output \g138421/_0_  ;
  output \g138422/_0_  ;
  output \g138423/_0_  ;
  output \g138424/_0_  ;
  output \g138425/_0_  ;
  output \g138426/_0_  ;
  output \g138427/_0_  ;
  output \g138428/_0_  ;
  output \g138429/_0_  ;
  output \g138430/_0_  ;
  output \g138431/_0_  ;
  output \g138432/_0_  ;
  output \g138433/_0_  ;
  output \g138434/_0_  ;
  output \g138435/_0_  ;
  output \g138436/_0_  ;
  output \g138437/_0_  ;
  output \g138438/_0_  ;
  output \g138439/_0_  ;
  output \g138440/_0_  ;
  output \g138441/_0_  ;
  output \g138442/_0_  ;
  output \g138443/_0_  ;
  output \g138908/_0_  ;
  output \g138909/_0_  ;
  output \g138910/_0_  ;
  output \g138914/_0_  ;
  output \g138915/_0_  ;
  output \g138917/_0_  ;
  output \g138918/_0_  ;
  output \g138919/_0_  ;
  output \g138920/_0_  ;
  output \g138921/_0_  ;
  output \g138925/_0_  ;
  output \g138926/_0_  ;
  output \g138927/_0_  ;
  output \g138930/_0_  ;
  output \g138931/_0_  ;
  output \g138932/_0_  ;
  output \g138960/_0_  ;
  output \g138962/_0_  ;
  output \g139037/_0_  ;
  output \g139038/_0_  ;
  output \g139040/_0_  ;
  output \g139043/_0_  ;
  output \g139044/_0_  ;
  output \g139045/_0_  ;
  output \g139046/_0_  ;
  output \g139047/_0_  ;
  output \g139048/_0_  ;
  output \g139049/_0_  ;
  output \g139050/_0_  ;
  output \g139051/_0_  ;
  output \g139053/_0_  ;
  output \g139054/_0_  ;
  output \g139055/_0_  ;
  output \g139056/_0_  ;
  output \g139057/_0_  ;
  output \g139058/_0_  ;
  output \g139059/_0_  ;
  output \g139060/_0_  ;
  output \g139062/_0_  ;
  output \g139063/_0_  ;
  output \g139064/_0_  ;
  output \g139099/_0_  ;
  output \g139126/_0_  ;
  output \g139127/_0_  ;
  output \g139128/_0_  ;
  output \g139129/_0_  ;
  output \g139130/_0_  ;
  output \g139131/_0_  ;
  output \g139132/_0_  ;
  output \g139133/_0_  ;
  output \g139134/_0_  ;
  output \g139135/_0_  ;
  output \g139136/_0_  ;
  output \g139137/_0_  ;
  output \g139138/_0_  ;
  output \g139139/_0_  ;
  output \g139140/_0_  ;
  output \g139141/_0_  ;
  output \g139260/_0_  ;
  output \g139263/_0_  ;
  output \g139267/_0_  ;
  output \g139270/_0_  ;
  output \g139273/_0_  ;
  output \g139276/_0_  ;
  output \g139279/_0_  ;
  output \g139283/_0_  ;
  output \g139286/_0_  ;
  output \g139289/_0_  ;
  output \g139292/_0_  ;
  output \g139295/_0_  ;
  output \g139298/_0_  ;
  output \g139302/_0_  ;
  output \g139305/_0_  ;
  output \g139309/_0_  ;
  output \g139871/_0_  ;
  output \g139872/_0_  ;
  output \g139873/_0_  ;
  output \g139874/_0_  ;
  output \g139875/_0_  ;
  output \g139876/_0_  ;
  output \g139877/_0_  ;
  output \g139878/_0_  ;
  output \g139879/_0_  ;
  output \g139880/_0_  ;
  output \g139881/_0_  ;
  output \g139882/_0_  ;
  output \g139883/_0_  ;
  output \g139884/_0_  ;
  output \g139885/_0_  ;
  output \g139886/_0_  ;
  output \g139887/_0_  ;
  output \g139888/_0_  ;
  output \g139889/_0_  ;
  output \g139890/_0_  ;
  output \g139891/_0_  ;
  output \g139892/_0_  ;
  output \g139893/_0_  ;
  output \g139895/_0_  ;
  output \g139896/_0_  ;
  output \g139899/_0_  ;
  output \g139901/_0_  ;
  output \g139902/_0_  ;
  output \g139903/_0_  ;
  output \g139904/_0_  ;
  output \g140285/_0_  ;
  output \g140288/_0_  ;
  output \g140329/_0_  ;
  output \g140774/_0_  ;
  output \g140832/_0_  ;
  output \g140834/_0_  ;
  output \g140836/_0_  ;
  output \g140838/_0_  ;
  output \g140840/_0_  ;
  output \g140842/_0_  ;
  output \g140844/_0_  ;
  output \g140846/_0_  ;
  output \g140847/_0_  ;
  output \g140848/_0_  ;
  output \g140850/_0_  ;
  output \g140851/_0_  ;
  output \g140852/_0_  ;
  output \g140853/_0_  ;
  output \g140855/_0_  ;
  output \g140857/_0_  ;
  output \g140861/_0_  ;
  output \g140923/_0_  ;
  output \g141178/_0_  ;
  output \g141179/_0_  ;
  output \g141180/_0_  ;
  output \g141480/_0_  ;
  output \g141495/_0_  ;
  output \g141497/_0_  ;
  output \g141562/_0_  ;
  output \g141563/_0_  ;
  output \g141564/_0_  ;
  output \g141589/_0_  ;
  output \g141617/_0_  ;
  output \g141618/_0_  ;
  output \g141621/_0_  ;
  output \g141625/_0_  ;
  output \g141626/_0_  ;
  output \g141630/_0_  ;
  output \g141634/_0_  ;
  output \g141638/_0_  ;
  output \g141642/_0_  ;
  output \g141646/_0_  ;
  output \g141649/_0_  ;
  output \g141651/_0_  ;
  output \g141652/_0_  ;
  output \g141655/_0_  ;
  output \g141658/_0_  ;
  output \g141661/_0_  ;
  output \g141663/_0_  ;
  output \g141664/_0_  ;
  output \g141667/_0_  ;
  output \g141671/_0_  ;
  output \g141706/_0_  ;
  output \g141976/_0_  ;
  output \g141977/_0_  ;
  output \g141994/_0_  ;
  output \g142246/_0_  ;
  output \g142247/_0_  ;
  output \g142253/_0_  ;
  output \g142689/_0_  ;
  output \g142693/_0_  ;
  output \g142701/_0_  ;
  output \g142704/_0_  ;
  output \g142707/_0_  ;
  output \g142710/_0_  ;
  output \g142713/_0_  ;
  output \g142714/_0_  ;
  output \g142717/_0_  ;
  output \g142720/_0_  ;
  output \g142723/_0_  ;
  output \g142727/_0_  ;
  output \g142734/_0_  ;
  output \g143080/_0_  ;
  output \g143081/_0_  ;
  output \g143083/_0_  ;
  output \g143149/_0_  ;
  output \g143150/_0_  ;
  output \g143153/_0_  ;
  output \g143752/_0_  ;
  output \g143753/_0_  ;
  output \g143759/_0_  ;
  output \g144242/_0_  ;
  output \g144243/_0_  ;
  output \g144244/_0_  ;
  output \g144245/_0_  ;
  output \g144246/_0_  ;
  output \g144249/_0_  ;
  output \g145699/_0_  ;
  output \g145700/_0_  ;
  output \g145702/_0_  ;
  output \g145756/_0_  ;
  output \g145757/_0_  ;
  output \g145758/_0_  ;
  output \g146850/_0_  ;
  output \g146851/_0_  ;
  output \g146864/_0_  ;
  output \g147277/_0_  ;
  output \g147278/_0_  ;
  output \g147279/_0_  ;
  output \g147304/_0_  ;
  output \g147305/_0_  ;
  output \g147306/_0_  ;
  output \g147338/_3_  ;
  output \g147339/_3_  ;
  output \g147340/_3_  ;
  output \g147341/_3_  ;
  output \g147342/_3_  ;
  output \g147343/_3_  ;
  output \g147344/_3_  ;
  output \g147345/_3_  ;
  output \g147346/_3_  ;
  output \g147347/_3_  ;
  output \g147348/_3_  ;
  output \g147349/_3_  ;
  output \g147350/_3_  ;
  output \g147351/_3_  ;
  output \g147352/_3_  ;
  output \g147353/_3_  ;
  output \g147354/_3_  ;
  output \g147355/_3_  ;
  output \g147356/_3_  ;
  output \g147357/_3_  ;
  output \g147358/_3_  ;
  output \g147359/_3_  ;
  output \g147360/_3_  ;
  output \g147362/_3_  ;
  output \g147363/_3_  ;
  output \g147364/_3_  ;
  output \g147365/_3_  ;
  output \g147366/_3_  ;
  output \g147367/_3_  ;
  output \g147368/_3_  ;
  output \g147369/_3_  ;
  output \g148630/_0_  ;
  output \g148631/_0_  ;
  output \g148676/_0_  ;
  output \g148785/_0_  ;
  output \g148788/_0_  ;
  output \g148789/_0_  ;
  output \g148834/_0_  ;
  output \g148836/_0_  ;
  output \g148838/_0_  ;
  output \g149836/_0_  ;
  output \g149837/_0_  ;
  output \g149838/_0_  ;
  output \g150142/_0_  ;
  output \g152366/_0_  ;
  output \g152367/_0_  ;
  output \g152368/_0_  ;
  output \g152426/_0_  ;
  output \g152427/_0_  ;
  output \g152428/_0_  ;
  output \g152586/_0_  ;
  output \g152587/_0_  ;
  output \g152588/_0_  ;
  output \g153217/_0_  ;
  output \g154117/_0_  ;
  output \g154118/_0_  ;
  output \g154130/_0_  ;
  output \g154269/_0_  ;
  output \g154270/_0_  ;
  output \g154284/_0_  ;
  output \g154682/_0_  ;
  output \g155004/_0_  ;
  output \g155020/_0_  ;
  output \g155121/_0_  ;
  output \g155124/_0_  ;
  output \g155126/_0_  ;
  output \g155228/_0_  ;
  output \g155229/_0_  ;
  output \g155230/_0_  ;
  output \g155326/_0_  ;
  output \g155327/_0_  ;
  output \g155330/_0_  ;
  output \g155353/_0_  ;
  output \g155354/_0_  ;
  output \g155356/_0_  ;
  output \g155602/_0_  ;
  output \g155633/_0_  ;
  output \g155634/_0_  ;
  output \g155699/_0_  ;
  output \g155708/_0_  ;
  output \g155715/_0_  ;
  output \g156008/_0_  ;
  output \g156013/_0_  ;
  output \g156019/_0_  ;
  output \g156352/_0_  ;
  output \g156353/_0_  ;
  output \g156356/_0_  ;
  output \g156359/_0_  ;
  output \g156360/_0_  ;
  output \g156361/_0_  ;
  output \g156464/_0_  ;
  output \g156465/_0_  ;
  output \g156469/_0_  ;
  output \g156777/_0_  ;
  output \g156778/_0_  ;
  output \g156789/_0_  ;
  output \g158956/_0_  ;
  output \g158957/_0_  ;
  output \g158966/_0_  ;
  output \g159429/_1_  ;
  output \g159477/_1_  ;
  output \g159500/_1_  ;
  output \g159681/_0_  ;
  output \g159890/_0_  ;
  output \g159950/_0_  ;
  output \g160246/_0_  ;
  output \g160846/_0_  ;
  output \g160860/_0_  ;
  output \g160961/_0_  ;
  output \g160987/_0_  ;
  output \g161000/_0_  ;
  output \g161005/_0_  ;
  output \g161042/_0_  ;
  output \g161119/_0_  ;
  output \g161143/_0_  ;
  output \g161150/_0_  ;
  output \g161172/_0_  ;
  output \g161207/_0_  ;
  output \g161315/_0_  ;
  output \g161332/_0_  ;
  output \g161421/_0_  ;
  output \g161492/_0_  ;
  output \g161541/_0_  ;
  output \g161623/_0_  ;
  output \g161655/_0_  ;
  output \g161678/_0_  ;
  output \g161709/_0_  ;
  output \g161737/_0_  ;
  output \g161751/_0_  ;
  output \g161756/_0_  ;
  output \g162016/_0_  ;
  output \g162020/_0_  ;
  output \g162024/_0_  ;
  output \g163326/_0_  ;
  output \g163326/_3_  ;
  output \g174072/_1_  ;
  output \g174360/_1_  ;
  output \g174391/_0_  ;
  output \g180307/_0_  ;
  output \g180335/_0_  ;
  output \g180369/_0_  ;
  output \g180385/_0_  ;
  output \g180395/_0_  ;
  output \g180442/_0_  ;
  output \g180453/_0_  ;
  output \g180524/_0_  ;
  output \g180586/_0_  ;
  output \g180596/_0_  ;
  output \g180606/_0_  ;
  output \g180654/_0_  ;
  output \g180715/_0_  ;
  output \g180805/_0_  ;
  output \g180836/_0_  ;
  output \g180929/_0_  ;
  output \g180944/_0_  ;
  output \g180975/_0_  ;
  output \g181036/_0_  ;
  output \g181072/_0_  ;
  output \g181083/_0_  ;
  output \g181093/_0_  ;
  output \g181127/_0_  ;
  output \g181137/_0_  ;
  output \g181150/_0_  ;
  output \g181160/_0_  ;
  output \g181180/_0_  ;
  output \g181191/_0_  ;
  output \g181238/_0_  ;
  output \g181262/_0_  ;
  output \g181270/_0_  ;
  output \g181280/_0_  ;
  output \g181315/_0_  ;
  output \g181366/_0_  ;
  output \g181385/_0_  ;
  output \g181458/_0_  ;
  output \g181464/_0_  ;
  output \g181478/_0_  ;
  output \g181522/_0_  ;
  output \g181537/_0_  ;
  output \g181584/_0_  ;
  output \g181669/_0_  ;
  output \g181681/_0_  ;
  output \g181719/_0_  ;
  output \g181778/_0_  ;
  output \g181840/_0_  ;
  output \g181936/_0_  ;
  output \g181986/_0_  ;
  output \g182000/_0_  ;
  output \g182083/_0_  ;
  output \g182179/_0_  ;
  output \g182201/_0_  ;
  output \g182227/_0_  ;
  output \g182316/_0_  ;
  output \g182358/_0_  ;
  output \g182473/_0_  ;
  output \g182678/_0_  ;
  output \g53/_0_  ;
  wire n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , n6000 , n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , n6089 , n6090 , n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , n6170 , n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , n6230 , n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , n6240 , n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , n6250 , n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , n6259 , n6260 , n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , n6300 , n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , n6310 , n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , n6320 , n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , n6340 , n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , n6349 , n6350 , n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , n6359 , n6360 , n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , n6367 , n6368 , n6369 , n6370 , n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , n6380 , n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , n6390 , n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , n6400 , n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , n6409 , n6410 , n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , n6420 , n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , n6429 , n6430 , n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , n6439 , n6440 , n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , n6449 , n6450 , n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , n6460 , n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , n6470 , n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , n6480 , n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , n6490 , n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , n6499 , n6500 , n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , n6509 , n6510 , n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , n6519 , n6520 , n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , n6529 , n6530 , n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , n6539 , n6540 , n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , n6549 , n6550 , n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , n6559 , n6560 , n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , n6569 , n6570 , n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , n6579 , n6580 , n6581 , n6582 , n6583 , n6584 , n6585 , n6586 , n6587 , n6588 , n6589 , n6590 , n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , n6599 , n6600 , n6601 , n6602 , n6603 , n6604 , n6605 , n6606 , n6607 , n6608 , n6609 , n6610 , n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , n6617 , n6618 , n6619 , n6620 , n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , n6627 , n6628 , n6629 , n6630 , n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , n6639 , n6640 , n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , n6647 , n6648 , n6649 , n6650 , n6651 , n6652 , n6653 , n6654 , n6655 , n6656 , n6657 , n6658 , n6659 , n6660 , n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , n6667 , n6668 , n6669 , n6670 , n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , n6679 , n6680 , n6681 , n6682 , n6683 , n6684 , n6685 , n6686 , n6687 , n6688 , n6689 , n6690 , n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , n6697 , n6698 , n6699 , n6700 , n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , n6707 , n6708 , n6709 , n6710 , n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , n6717 , n6718 , n6719 , n6720 , n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , n6729 , n6730 , n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , n6739 , n6740 , n6741 , n6742 , n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , n6749 , n6750 , n6751 , n6752 , n6753 , n6754 , n6755 , n6756 , n6757 , n6758 , n6759 , n6760 , n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , n6770 , n6771 , n6772 , n6773 , n6774 , n6775 , n6776 , n6777 , n6778 , n6779 , n6780 , n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , n6789 , n6790 , n6791 , n6792 , n6793 , n6794 , n6795 , n6796 , n6797 , n6798 , n6799 , n6800 , n6801 , n6802 , n6803 , n6804 , n6805 , n6806 , n6807 , n6808 , n6809 , n6810 , n6811 , n6812 , n6813 , n6814 , n6815 , n6816 , n6817 , n6818 , n6819 , n6820 , n6821 , n6822 , n6823 , n6824 , n6825 , n6826 , n6827 , n6828 , n6829 , n6830 , n6831 , n6832 , n6833 , n6834 , n6835 , n6836 , n6837 , n6838 , n6839 , n6840 , n6841 , n6842 , n6843 , n6844 , n6845 , n6846 , n6847 , n6848 , n6849 , n6850 , n6851 , n6852 , n6853 , n6854 , n6855 , n6856 , n6857 , n6858 , n6859 , n6860 , n6861 , n6862 , n6863 , n6864 , n6865 , n6866 , n6867 , n6868 , n6869 , n6870 , n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , n6877 , n6878 , n6879 , n6880 , n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , n6887 , n6888 , n6889 , n6890 , n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , n6897 , n6898 , n6899 , n6900 , n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , n6907 , n6908 , n6909 , n6910 , n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , n6919 , n6920 , n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , n6927 , n6928 , n6929 , n6930 , n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , n6937 , n6938 , n6939 , n6940 , n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , n6949 , n6950 , n6951 , n6952 , n6953 , n6954 , n6955 , n6956 , n6957 , n6958 , n6959 , n6960 , n6961 , n6962 , n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , n6969 , n6970 , n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , n6979 , n6980 , n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , n6987 , n6988 , n6989 , n6990 , n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , n6997 , n6998 , n6999 , n7000 , n7001 , n7002 , n7003 , n7004 , n7005 , n7006 , n7007 , n7008 , n7009 , n7010 , n7011 , n7012 , n7013 , n7014 , n7015 , n7016 , n7017 , n7018 , n7019 , n7020 , n7021 , n7022 , n7023 , n7024 , n7025 , n7026 , n7027 , n7028 , n7029 , n7030 , n7031 , n7032 , n7033 , n7034 , n7035 , n7036 , n7037 , n7038 , n7039 , n7040 , n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , n7047 , n7048 , n7049 , n7050 , n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , n7057 , n7058 , n7059 , n7060 , n7061 , n7062 , n7063 , n7064 , n7065 , n7066 , n7067 , n7068 , n7069 , n7070 , n7071 , n7072 , n7073 , n7074 , n7075 , n7076 , n7077 , n7078 , n7079 , n7080 , n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , n7087 , n7088 , n7089 , n7090 , n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , n7097 , n7098 , n7099 , n7100 , n7101 , n7102 , n7103 , n7104 , n7105 , n7106 , n7107 , n7108 , n7109 , n7110 , n7111 , n7112 , n7113 , n7114 , n7115 , n7116 , n7117 , n7118 , n7119 , n7120 , n7121 , n7122 , n7123 , n7124 , n7125 , n7126 , n7127 , n7128 , n7129 , n7130 , n7131 , n7132 , n7133 , n7134 , n7135 , n7136 , n7137 , n7138 , n7139 , n7140 , n7141 , n7142 , n7143 , n7144 , n7145 , n7146 , n7147 , n7148 , n7149 , n7150 , n7151 , n7152 , n7153 , n7154 , n7155 , n7156 , n7157 , n7158 , n7159 , n7160 , n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , n7167 , n7168 , n7169 , n7170 , n7171 , n7172 , n7173 , n7174 , n7175 , n7176 , n7177 , n7178 , n7179 , n7180 , n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , n7187 , n7188 , n7189 , n7190 , n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , n7197 , n7198 , n7199 , n7200 , n7201 , n7202 , n7203 , n7204 , n7205 , n7206 , n7207 , n7208 , n7209 , n7210 , n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , n7217 , n7218 , n7219 , n7220 , n7221 , n7222 , n7223 , n7224 , n7225 , n7226 , n7227 , n7228 , n7229 , n7230 , n7231 , n7232 , n7233 , n7234 , n7235 , n7236 , n7237 , n7238 , n7239 , n7240 , n7241 , n7242 , n7243 , n7244 , n7245 , n7246 , n7247 , n7248 , n7249 , n7250 , n7251 , n7252 , n7253 , n7254 , n7255 , n7256 , n7257 , n7258 , n7259 , n7260 , n7261 , n7262 , n7263 , n7264 , n7265 , n7266 , n7267 , n7268 , n7269 , n7270 , n7271 , n7272 , n7273 , n7274 , n7275 , n7276 , n7277 , n7278 , n7279 , n7280 , n7281 , n7282 , n7283 , n7284 , n7285 , n7286 , n7287 , n7288 , n7289 , n7290 , n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , n7297 , n7298 , n7299 , n7300 , n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , n7307 , n7308 , n7309 , n7310 , n7311 , n7312 , n7313 , n7314 , n7315 , n7316 , n7317 , n7318 , n7319 , n7320 , n7321 , n7322 , n7323 , n7324 , n7325 , n7326 , n7327 , n7328 , n7329 , n7330 , n7331 , n7332 , n7333 , n7334 , n7335 , n7336 , n7337 , n7338 , n7339 , n7340 , n7341 , n7342 , n7343 , n7344 , n7345 , n7346 , n7347 , n7348 , n7349 , n7350 , n7351 , n7352 , n7353 , n7354 , n7355 , n7356 , n7357 , n7358 , n7359 , n7360 , n7361 , n7362 , n7363 , n7364 , n7365 , n7366 , n7367 , n7368 , n7369 , n7370 , n7371 , n7372 , n7373 , n7374 , n7375 , n7376 , n7377 , n7378 , n7379 , n7380 , n7381 , n7382 , n7383 , n7384 , n7385 , n7386 , n7387 , n7388 , n7389 , n7390 , n7391 , n7392 , n7393 , n7394 , n7395 , n7396 , n7397 , n7398 , n7399 , n7400 , n7401 , n7402 , n7403 , n7404 , n7405 , n7406 , n7407 , n7408 , n7409 , n7410 , n7411 , n7412 , n7413 , n7414 , n7415 , n7416 , n7417 , n7418 , n7419 , n7420 , n7421 , n7422 , n7423 , n7424 , n7425 , n7426 , n7427 , n7428 , n7429 , n7430 , n7431 , n7432 , n7433 , n7434 , n7435 , n7436 , n7437 , n7438 , n7439 , n7440 , n7441 , n7442 , n7443 , n7444 , n7445 , n7446 , n7447 , n7448 , n7449 , n7450 , n7451 , n7452 , n7453 , n7454 , n7455 , n7456 , n7457 , n7458 , n7459 , n7460 , n7461 , n7462 , n7463 , n7464 , n7465 , n7466 , n7467 , n7468 , n7469 , n7470 , n7471 , n7472 , n7473 , n7474 , n7475 , n7476 , n7477 , n7478 , n7479 , n7480 , n7481 , n7482 , n7483 , n7484 , n7485 , n7486 , n7487 , n7488 , n7489 , n7490 , n7491 , n7492 , n7493 , n7494 , n7495 , n7496 , n7497 , n7498 , n7499 , n7500 , n7501 , n7502 , n7503 , n7504 , n7505 , n7506 , n7507 , n7508 , n7509 , n7510 , n7511 , n7512 , n7513 , n7514 , n7515 , n7516 , n7517 , n7518 , n7519 , n7520 , n7521 , n7522 , n7523 , n7524 , n7525 , n7526 , n7527 , n7528 , n7529 , n7530 , n7531 , n7532 , n7533 , n7534 , n7535 , n7536 , n7537 , n7538 , n7539 , n7540 , n7541 , n7542 , n7543 , n7544 , n7545 , n7546 , n7547 , n7548 , n7549 , n7550 , n7551 , n7552 , n7553 , n7554 , n7555 , n7556 , n7557 , n7558 , n7559 , n7560 , n7561 , n7562 , n7563 , n7564 , n7565 , n7566 , n7567 , n7568 , n7569 , n7570 , n7571 , n7572 , n7573 , n7574 , n7575 , n7576 , n7577 , n7578 , n7579 , n7580 , n7581 , n7582 , n7583 , n7584 , n7585 , n7586 , n7587 , n7588 , n7589 , n7590 , n7591 , n7592 , n7593 , n7594 , n7595 , n7596 , n7597 , n7598 , n7599 , n7600 , n7601 , n7602 , n7603 , n7604 , n7605 , n7606 , n7607 , n7608 , n7609 , n7610 , n7611 , n7612 , n7613 , n7614 , n7615 , n7616 , n7617 , n7618 , n7619 , n7620 , n7621 , n7622 , n7623 , n7624 , n7625 , n7626 , n7627 , n7628 , n7629 , n7630 , n7631 , n7632 , n7633 , n7634 , n7635 , n7636 , n7637 , n7638 , n7639 , n7640 , n7641 , n7642 , n7643 , n7644 , n7645 , n7646 , n7647 , n7648 , n7649 , n7650 , n7651 , n7652 , n7653 , n7654 , n7655 , n7656 , n7657 , n7658 , n7659 , n7660 , n7661 , n7662 , n7663 , n7664 , n7665 , n7666 , n7667 , n7668 , n7669 , n7670 , n7671 , n7672 , n7673 , n7674 , n7675 , n7676 , n7677 , n7678 , n7679 , n7680 , n7681 , n7682 , n7683 , n7684 , n7685 , n7686 , n7687 , n7688 , n7689 , n7690 , n7691 , n7692 , n7693 , n7694 , n7695 , n7696 , n7697 , n7698 , n7699 , n7700 , n7701 , n7702 , n7703 , n7704 , n7705 , n7706 , n7707 , n7708 , n7709 , n7710 , n7711 , n7712 , n7713 , n7714 , n7715 , n7716 , n7717 , n7718 , n7719 , n7720 , n7721 , n7722 , n7723 , n7724 , n7725 , n7726 , n7727 , n7728 , n7729 , n7730 , n7731 , n7732 , n7733 , n7734 , n7735 , n7736 , n7737 , n7738 , n7739 , n7740 , n7741 , n7742 , n7743 , n7744 , n7745 , n7746 , n7747 , n7748 , n7749 , n7750 , n7751 , n7752 , n7753 , n7754 , n7755 , n7756 , n7757 , n7758 , n7759 , n7760 , n7761 , n7762 , n7763 , n7764 , n7765 , n7766 , n7767 , n7768 , n7769 , n7770 , n7771 , n7772 , n7773 , n7774 , n7775 , n7776 , n7777 , n7778 , n7779 , n7780 , n7781 , n7782 , n7783 , n7784 , n7785 , n7786 , n7787 , n7788 , n7789 , n7790 , n7791 , n7792 , n7793 , n7794 , n7795 , n7796 , n7797 , n7798 , n7799 , n7800 , n7801 , n7802 , n7803 , n7804 , n7805 , n7806 , n7807 , n7808 , n7809 , n7810 , n7811 , n7812 , n7813 , n7814 , n7815 , n7816 , n7817 , n7818 , n7819 , n7820 , n7821 , n7822 , n7823 , n7824 , n7825 , n7826 , n7827 , n7828 , n7829 , n7830 , n7831 , n7832 , n7833 , n7834 , n7835 , n7836 , n7837 , n7838 , n7839 , n7840 , n7841 , n7842 , n7843 , n7844 , n7845 , n7846 , n7847 , n7848 , n7849 , n7850 , n7851 , n7852 , n7853 , n7854 , n7855 , n7856 , n7857 , n7858 , n7859 , n7860 , n7861 , n7862 , n7863 , n7864 , n7865 , n7866 , n7867 , n7868 , n7869 , n7870 , n7871 , n7872 , n7873 , n7874 , n7875 , n7876 , n7877 , n7878 , n7879 , n7880 , n7881 , n7882 , n7883 , n7884 , n7885 , n7886 , n7887 , n7888 , n7889 , n7890 , n7891 , n7892 , n7893 , n7894 , n7895 , n7896 , n7897 , n7898 , n7899 , n7900 , n7901 , n7902 , n7903 , n7904 , n7905 , n7906 , n7907 , n7908 , n7909 , n7910 , n7911 , n7912 , n7913 , n7914 , n7915 , n7916 , n7917 , n7918 , n7919 , n7920 , n7921 , n7922 , n7923 , n7924 , n7925 , n7926 , n7927 , n7928 , n7929 , n7930 , n7931 , n7932 , n7933 , n7934 , n7935 , n7936 , n7937 , n7938 , n7939 , n7940 , n7941 , n7942 , n7943 , n7944 , n7945 , n7946 , n7947 , n7948 , n7949 , n7950 , n7951 , n7952 , n7953 , n7954 , n7955 , n7956 , n7957 , n7958 , n7959 , n7960 , n7961 , n7962 , n7963 , n7964 , n7965 , n7966 , n7967 , n7968 , n7969 , n7970 , n7971 , n7972 , n7973 , n7974 , n7975 , n7976 , n7977 , n7978 , n7979 , n7980 , n7981 , n7982 , n7983 , n7984 , n7985 , n7986 , n7987 , n7988 , n7989 , n7990 , n7991 , n7992 , n7993 , n7994 , n7995 , n7996 , n7997 , n7998 , n7999 , n8000 , n8001 , n8002 , n8003 , n8004 , n8005 , n8006 , n8007 , n8008 , n8009 , n8010 , n8011 , n8012 , n8013 , n8014 , n8015 , n8016 , n8017 , n8018 , n8019 , n8020 , n8021 , n8022 , n8023 , n8024 , n8025 , n8026 , n8027 , n8028 , n8029 , n8030 , n8031 , n8032 , n8033 , n8034 , n8035 , n8036 , n8037 , n8038 , n8039 , n8040 , n8041 , n8042 , n8043 , n8044 , n8045 , n8046 , n8047 , n8048 , n8049 , n8050 , n8051 , n8052 , n8053 , n8054 , n8055 , n8056 , n8057 , n8058 , n8059 , n8060 , n8061 , n8062 , n8063 , n8064 , n8065 , n8066 , n8067 , n8068 , n8069 , n8070 , n8071 , n8072 , n8073 , n8074 , n8075 , n8076 , n8077 , n8078 , n8079 , n8080 , n8081 , n8082 , n8083 , n8084 , n8085 , n8086 , n8087 , n8088 , n8089 , n8090 , n8091 , n8092 , n8093 , n8094 , n8095 , n8096 , n8097 , n8098 , n8099 , n8100 , n8101 , n8102 , n8103 , n8104 , n8105 , n8106 , n8107 , n8108 , n8109 , n8110 , n8111 , n8112 , n8113 , n8114 , n8115 , n8116 , n8117 , n8118 , n8119 , n8120 , n8121 , n8122 , n8123 , n8124 , n8125 , n8126 , n8127 , n8128 , n8129 , n8130 , n8131 , n8132 , n8133 , n8134 , n8135 , n8136 , n8137 , n8138 , n8139 , n8140 , n8141 , n8142 , n8143 , n8144 , n8145 , n8146 , n8147 , n8148 , n8149 , n8150 , n8151 , n8152 , n8153 , n8154 , n8155 , n8156 , n8157 , n8158 , n8159 , n8160 , n8161 , n8162 , n8163 , n8164 , n8165 , n8166 , n8167 , n8168 , n8169 , n8170 , n8171 , n8172 , n8173 , n8174 , n8175 , n8176 , n8177 , n8178 , n8179 , n8180 , n8181 , n8182 , n8183 , n8184 , n8185 , n8186 , n8187 , n8188 , n8189 , n8190 , n8191 , n8192 , n8193 , n8194 , n8195 , n8196 , n8197 , n8198 , n8199 , n8200 , n8201 , n8202 , n8203 , n8204 , n8205 , n8206 , n8207 , n8208 , n8209 , n8210 , n8211 , n8212 , n8213 , n8214 , n8215 , n8216 , n8217 , n8218 , n8219 , n8220 , n8221 , n8222 , n8223 , n8224 , n8225 , n8226 , n8227 , n8228 , n8229 , n8230 , n8231 , n8232 , n8233 , n8234 , n8235 , n8236 , n8237 , n8238 , n8239 , n8240 , n8241 , n8242 , n8243 , n8244 , n8245 , n8246 , n8247 , n8248 , n8249 , n8250 , n8251 , n8252 , n8253 , n8254 , n8255 , n8256 , n8257 , n8258 , n8259 , n8260 , n8261 , n8262 , n8263 , n8264 , n8265 , n8266 , n8267 , n8268 , n8269 , n8270 , n8271 , n8272 , n8273 , n8274 , n8275 , n8276 , n8277 , n8278 , n8279 , n8280 , n8281 , n8282 , n8283 , n8284 , n8285 , n8286 , n8287 , n8288 , n8289 , n8290 , n8291 , n8292 , n8293 , n8294 , n8295 , n8296 , n8297 , n8298 , n8299 , n8300 , n8301 , n8302 , n8303 , n8304 , n8305 , n8306 , n8307 , n8308 , n8309 , n8310 , n8311 , n8312 , n8313 , n8314 , n8315 , n8316 , n8317 , n8318 , n8319 , n8320 , n8321 , n8322 , n8323 , n8324 , n8325 , n8326 , n8327 , n8328 , n8329 , n8330 , n8331 , n8332 , n8333 , n8334 , n8335 , n8336 , n8337 , n8338 , n8339 , n8340 , n8341 , n8342 , n8343 , n8344 , n8345 , n8346 , n8347 , n8348 , n8349 , n8350 , n8351 , n8352 , n8353 , n8354 , n8355 , n8356 , n8357 , n8358 , n8359 , n8360 , n8361 , n8362 , n8363 , n8364 , n8365 , n8366 , n8367 , n8368 , n8369 , n8370 , n8371 , n8372 , n8373 , n8374 , n8375 , n8376 , n8377 , n8378 , n8379 , n8380 , n8381 , n8382 , n8383 , n8384 , n8385 , n8386 , n8387 , n8388 , n8389 , n8390 , n8391 , n8392 , n8393 , n8394 , n8395 , n8396 , n8397 , n8398 , n8399 , n8400 , n8401 , n8402 , n8403 , n8404 , n8405 , n8406 , n8407 , n8408 , n8409 , n8410 , n8411 , n8412 , n8413 , n8414 , n8415 , n8416 , n8417 , n8418 , n8419 , n8420 , n8421 , n8422 , n8423 , n8424 , n8425 , n8426 , n8427 , n8428 , n8429 , n8430 , n8431 , n8432 , n8433 , n8434 , n8435 , n8436 , n8437 , n8438 , n8439 , n8440 , n8441 , n8442 , n8443 , n8444 , n8445 , n8446 , n8447 , n8448 , n8449 , n8450 , n8451 , n8452 , n8453 , n8454 , n8455 , n8456 , n8457 , n8458 , n8459 , n8460 , n8461 , n8462 , n8463 , n8464 , n8465 , n8466 , n8467 , n8468 , n8469 , n8470 , n8471 , n8472 , n8473 , n8474 , n8475 , n8476 , n8477 , n8478 , n8479 , n8480 , n8481 , n8482 , n8483 , n8484 , n8485 , n8486 , n8487 , n8488 , n8489 , n8490 , n8491 , n8492 , n8493 , n8494 , n8495 , n8496 , n8497 , n8498 , n8499 , n8500 , n8501 , n8502 , n8503 , n8504 , n8505 , n8506 , n8507 , n8508 , n8509 , n8510 , n8511 , n8512 , n8513 , n8514 , n8515 , n8516 , n8517 , n8518 , n8519 , n8520 , n8521 , n8522 , n8523 , n8524 , n8525 , n8526 , n8527 , n8528 , n8529 , n8530 , n8531 , n8532 , n8533 , n8534 , n8535 , n8536 , n8537 , n8538 , n8539 , n8540 , n8541 , n8542 , n8543 , n8544 , n8545 , n8546 , n8547 , n8548 , n8549 , n8550 , n8551 , n8552 , n8553 , n8554 , n8555 , n8556 , n8557 , n8558 , n8559 , n8560 , n8561 , n8562 , n8563 , n8564 , n8565 , n8566 , n8567 , n8568 , n8569 , n8570 , n8571 , n8572 , n8573 , n8574 , n8575 , n8576 , n8577 , n8578 , n8579 , n8580 , n8581 , n8582 , n8583 , n8584 , n8585 , n8586 , n8587 , n8588 , n8589 , n8590 , n8591 , n8592 , n8593 , n8594 , n8595 , n8596 , n8597 , n8598 , n8599 , n8600 , n8601 , n8602 , n8603 , n8604 , n8605 , n8606 , n8607 , n8608 , n8609 , n8610 , n8611 , n8612 , n8613 , n8614 , n8615 , n8616 , n8617 , n8618 , n8619 , n8620 , n8621 , n8622 , n8623 , n8624 , n8625 , n8626 , n8627 , n8628 , n8629 , n8630 , n8631 , n8632 , n8633 , n8634 , n8635 , n8636 , n8637 , n8638 , n8639 , n8640 , n8641 , n8642 , n8643 , n8644 , n8645 , n8646 , n8647 , n8648 , n8649 , n8650 , n8651 , n8652 , n8653 , n8654 , n8655 , n8656 , n8657 , n8658 , n8659 , n8660 , n8661 , n8662 , n8663 , n8664 , n8665 , n8666 , n8667 , n8668 , n8669 , n8670 , n8671 , n8672 , n8673 , n8674 , n8675 , n8676 , n8677 , n8678 , n8679 , n8680 , n8681 , n8682 , n8683 , n8684 , n8685 , n8686 , n8687 , n8688 , n8689 , n8690 , n8691 , n8692 , n8693 , n8694 , n8695 , n8696 , n8697 , n8698 , n8699 , n8700 , n8701 , n8702 , n8703 , n8704 , n8705 , n8706 , n8707 , n8708 , n8709 , n8710 , n8711 , n8712 , n8713 , n8714 , n8715 , n8716 , n8717 , n8718 , n8719 , n8720 , n8721 , n8722 , n8723 , n8724 , n8725 , n8726 , n8727 , n8728 , n8729 , n8730 , n8731 , n8732 , n8733 , n8734 , n8735 , n8736 , n8737 , n8738 , n8739 , n8740 , n8741 , n8742 , n8743 , n8744 , n8745 , n8746 , n8747 , n8748 , n8749 , n8750 , n8751 , n8752 , n8753 , n8754 , n8755 , n8756 , n8757 , n8758 , n8759 , n8760 , n8761 , n8762 , n8763 , n8764 , n8765 , n8766 , n8767 , n8768 , n8769 , n8770 , n8771 , n8772 , n8773 , n8774 , n8775 , n8776 , n8777 , n8778 , n8779 , n8780 , n8781 , n8782 , n8783 , n8784 , n8785 , n8786 , n8787 , n8788 , n8789 , n8790 , n8791 , n8792 , n8793 , n8794 , n8795 , n8796 , n8797 , n8798 , n8799 , n8800 , n8801 , n8802 , n8803 , n8804 , n8805 , n8806 , n8807 , n8808 , n8809 , n8810 , n8811 , n8812 , n8813 , n8814 , n8815 , n8816 , n8817 , n8818 , n8819 , n8820 , n8821 , n8822 , n8823 , n8824 , n8825 , n8826 , n8827 , n8828 , n8829 , n8830 , n8831 , n8832 , n8833 , n8834 , n8835 , n8836 , n8837 , n8838 , n8839 , n8840 , n8841 , n8842 , n8843 , n8844 , n8845 , n8846 , n8847 , n8848 , n8849 , n8850 , n8851 , n8852 , n8853 , n8854 , n8855 , n8856 , n8857 , n8858 , n8859 , n8860 , n8861 , n8862 , n8863 , n8864 , n8865 , n8866 , n8867 , n8868 , n8869 , n8870 , n8871 , n8872 , n8873 , n8874 , n8875 , n8876 , n8877 , n8878 , n8879 , n8880 , n8881 , n8882 , n8883 , n8884 , n8885 , n8886 , n8887 , n8888 , n8889 , n8890 , n8891 , n8892 , n8893 , n8894 , n8895 , n8896 , n8897 , n8898 , n8899 , n8900 , n8901 , n8902 , n8903 , n8904 , n8905 , n8906 , n8907 , n8908 , n8909 , n8910 , n8911 , n8912 , n8913 , n8914 , n8915 , n8916 , n8917 , n8918 , n8919 , n8920 , n8921 , n8922 , n8923 , n8924 , n8925 , n8926 , n8927 , n8928 , n8929 , n8930 , n8931 , n8932 , n8933 , n8934 , n8935 , n8936 , n8937 , n8938 , n8939 , n8940 , n8941 , n8942 , n8943 , n8944 , n8945 , n8946 , n8947 , n8948 , n8949 , n8950 , n8951 , n8952 , n8953 , n8954 , n8955 , n8956 , n8957 , n8958 , n8959 , n8960 , n8961 , n8962 , n8963 , n8964 , n8965 , n8966 , n8967 , n8968 , n8969 , n8970 , n8971 , n8972 , n8973 , n8974 , n8975 , n8976 , n8977 , n8978 , n8979 , n8980 , n8981 , n8982 , n8983 , n8984 , n8985 , n8986 , n8987 , n8988 , n8989 , n8990 , n8991 , n8992 , n8993 , n8994 , n8995 , n8996 , n8997 , n8998 , n8999 , n9000 , n9001 , n9002 , n9003 , n9004 , n9005 , n9006 , n9007 , n9008 , n9009 , n9010 , n9011 , n9012 , n9013 , n9014 , n9015 , n9016 , n9017 , n9018 , n9019 , n9020 , n9021 , n9022 , n9023 , n9024 , n9025 , n9026 , n9027 , n9028 , n9029 , n9030 , n9031 , n9032 , n9033 , n9034 , n9035 , n9036 , n9037 , n9038 , n9039 , n9040 , n9041 , n9042 , n9043 , n9044 , n9045 , n9046 , n9047 , n9048 , n9049 , n9050 , n9051 , n9052 , n9053 , n9054 , n9055 , n9056 , n9057 , n9058 , n9059 , n9060 , n9061 , n9062 , n9063 , n9064 , n9065 , n9066 , n9067 , n9068 , n9069 , n9070 , n9071 , n9072 , n9073 , n9074 , n9075 , n9076 , n9077 , n9078 , n9079 , n9080 , n9081 , n9082 , n9083 , n9084 , n9085 , n9086 , n9087 , n9088 , n9089 , n9090 , n9091 , n9092 , n9093 , n9094 , n9095 , n9096 , n9097 , n9098 , n9099 , n9100 , n9101 , n9102 , n9103 , n9104 , n9105 , n9106 , n9107 , n9108 , n9109 , n9110 , n9111 , n9112 , n9113 , n9114 , n9115 , n9116 , n9117 , n9118 , n9119 , n9120 , n9121 , n9122 , n9123 , n9124 , n9125 , n9126 , n9127 , n9128 , n9129 , n9130 , n9131 , n9132 , n9133 , n9134 , n9135 , n9136 , n9137 , n9138 , n9139 , n9140 , n9141 , n9142 , n9143 , n9144 , n9145 , n9146 , n9147 , n9148 , n9149 , n9150 , n9151 , n9152 , n9153 , n9154 , n9155 , n9156 , n9157 , n9158 , n9159 , n9160 , n9161 , n9162 , n9163 , n9164 , n9165 , n9166 , n9167 , n9168 , n9169 , n9170 , n9171 , n9172 , n9173 , n9174 , n9175 , n9176 , n9177 , n9178 , n9179 , n9180 , n9181 , n9182 , n9183 , n9184 , n9185 , n9186 , n9187 , n9188 , n9189 , n9190 , n9191 , n9192 , n9193 , n9194 , n9195 , n9196 , n9197 , n9198 , n9199 , n9200 , n9201 , n9202 , n9203 , n9204 , n9205 , n9206 , n9207 , n9208 , n9209 , n9210 , n9211 , n9212 , n9213 , n9214 , n9215 , n9216 , n9217 , n9218 , n9219 , n9220 , n9221 , n9222 , n9223 , n9224 , n9225 , n9226 , n9227 , n9228 , n9229 , n9230 , n9231 , n9232 , n9233 , n9234 , n9235 , n9236 , n9237 , n9238 , n9239 , n9240 , n9241 , n9242 , n9243 , n9244 , n9245 , n9246 , n9247 , n9248 , n9249 , n9250 , n9251 , n9252 , n9253 , n9254 , n9255 , n9256 , n9257 , n9258 , n9259 , n9260 , n9261 , n9262 , n9263 , n9264 , n9265 , n9266 , n9267 , n9268 , n9269 , n9270 , n9271 , n9272 , n9273 , n9274 , n9275 , n9276 , n9277 , n9278 , n9279 , n9280 , n9281 , n9282 , n9283 , n9284 , n9285 , n9286 , n9287 , n9288 , n9289 , n9290 , n9291 , n9292 , n9293 , n9294 , n9295 , n9296 , n9297 , n9298 , n9299 , n9300 , n9301 , n9302 , n9303 , n9304 , n9305 , n9306 , n9307 , n9308 , n9309 , n9310 , n9311 , n9312 , n9313 , n9314 , n9315 , n9316 , n9317 , n9318 , n9319 , n9320 , n9321 , n9322 , n9323 , n9324 , n9325 , n9326 , n9327 , n9328 , n9329 , n9330 , n9331 , n9332 , n9333 , n9334 , n9335 , n9336 , n9337 , n9338 , n9339 , n9340 , n9341 , n9342 , n9343 , n9344 , n9345 , n9346 , n9347 , n9348 , n9349 , n9350 , n9351 , n9352 , n9353 , n9354 , n9355 , n9356 , n9357 , n9358 , n9359 , n9360 , n9361 , n9362 , n9363 , n9364 , n9365 , n9366 , n9367 , n9368 , n9369 , n9370 , n9371 , n9372 , n9373 , n9374 , n9375 , n9376 , n9377 , n9378 , n9379 , n9380 , n9381 , n9382 , n9383 , n9384 , n9385 , n9386 , n9387 , n9388 , n9389 , n9390 , n9391 , n9392 , n9393 , n9394 , n9395 , n9396 , n9397 , n9398 , n9399 , n9400 , n9401 , n9402 , n9403 , n9404 , n9405 , n9406 , n9407 , n9408 , n9409 , n9410 , n9411 , n9412 , n9413 , n9414 , n9415 , n9416 , n9417 , n9418 , n9419 , n9420 , n9421 , n9422 , n9423 , n9424 , n9425 , n9426 , n9427 , n9428 , n9429 , n9430 , n9431 , n9432 , n9433 , n9434 , n9435 , n9436 , n9437 , n9438 , n9439 , n9440 , n9441 , n9442 , n9443 , n9444 , n9445 , n9446 , n9447 , n9448 , n9449 , n9450 , n9451 , n9452 , n9453 , n9454 , n9455 , n9456 , n9457 , n9458 , n9459 , n9460 , n9461 , n9462 , n9463 , n9464 , n9465 , n9466 , n9467 , n9468 , n9469 , n9470 , n9471 , n9472 , n9473 , n9474 , n9475 , n9476 , n9477 , n9478 , n9479 , n9480 , n9481 , n9482 , n9483 , n9484 , n9485 , n9486 , n9487 , n9488 , n9489 , n9490 , n9491 , n9492 , n9493 , n9494 , n9495 , n9496 , n9497 , n9498 , n9499 , n9500 , n9501 , n9502 , n9503 , n9504 , n9505 , n9506 , n9507 , n9508 , n9509 , n9510 , n9511 , n9512 , n9513 , n9514 , n9515 , n9516 , n9517 , n9518 , n9519 , n9520 , n9521 , n9522 , n9523 , n9524 , n9525 , n9526 , n9527 , n9528 , n9529 , n9530 , n9531 , n9532 , n9533 , n9534 , n9535 , n9536 , n9537 , n9538 , n9539 , n9540 , n9541 , n9542 , n9543 , n9544 , n9545 , n9546 , n9547 , n9548 , n9549 , n9550 , n9551 , n9552 , n9553 , n9554 , n9555 , n9556 , n9557 , n9558 , n9559 , n9560 , n9561 , n9562 , n9563 , n9564 , n9565 , n9566 , n9567 , n9568 , n9569 , n9570 , n9571 , n9572 , n9573 , n9574 , n9575 , n9576 , n9577 , n9578 , n9579 , n9580 , n9581 , n9582 , n9583 , n9584 , n9585 , n9586 , n9587 , n9588 , n9589 , n9590 , n9591 , n9592 , n9593 , n9594 , n9595 , n9596 , n9597 , n9598 , n9599 , n9600 , n9601 , n9602 , n9603 , n9604 , n9605 , n9606 , n9607 , n9608 , n9609 , n9610 , n9611 , n9612 , n9613 , n9614 , n9615 , n9616 , n9617 , n9618 , n9619 , n9620 , n9621 , n9622 , n9623 , n9624 , n9625 , n9626 , n9627 , n9628 , n9629 , n9630 , n9631 , n9632 , n9633 , n9634 , n9635 , n9636 , n9637 , n9638 , n9639 , n9640 , n9641 , n9642 , n9643 , n9644 , n9645 , n9646 , n9647 , n9648 , n9649 , n9650 , n9651 , n9652 , n9653 , n9654 , n9655 , n9656 , n9657 , n9658 , n9659 , n9660 , n9661 , n9662 , n9663 , n9664 , n9665 , n9666 , n9667 , n9668 , n9669 , n9670 , n9671 , n9672 , n9673 , n9674 , n9675 , n9676 , n9677 , n9678 , n9679 , n9680 , n9681 , n9682 , n9683 , n9684 , n9685 , n9686 , n9687 , n9688 , n9689 , n9690 , n9691 , n9692 , n9693 , n9694 , n9695 , n9696 , n9697 , n9698 , n9699 , n9700 , n9701 , n9702 , n9703 , n9704 , n9705 , n9706 , n9707 , n9708 , n9709 , n9710 , n9711 , n9712 , n9713 , n9714 , n9715 , n9716 , n9717 , n9718 , n9719 , n9720 , n9721 , n9722 , n9723 , n9724 , n9725 , n9726 , n9727 , n9728 , n9729 , n9730 , n9731 , n9732 , n9733 , n9734 , n9735 , n9736 , n9737 , n9738 , n9739 , n9740 , n9741 , n9742 , n9743 , n9744 , n9745 , n9746 , n9747 , n9748 , n9749 , n9750 , n9751 , n9752 , n9753 , n9754 , n9755 , n9756 , n9757 , n9758 , n9759 , n9760 , n9761 , n9762 , n9763 , n9764 , n9765 , n9766 , n9767 , n9768 , n9769 , n9770 , n9771 , n9772 , n9773 , n9774 , n9775 , n9776 , n9777 , n9778 , n9779 , n9780 , n9781 , n9782 , n9783 , n9784 , n9785 , n9786 , n9787 , n9788 , n9789 , n9790 , n9791 , n9792 , n9793 , n9794 , n9795 , n9796 , n9797 , n9798 , n9799 , n9800 , n9801 , n9802 , n9803 , n9804 , n9805 , n9806 , n9807 , n9808 , n9809 , n9810 , n9811 , n9812 , n9813 , n9814 , n9815 , n9816 , n9817 , n9818 , n9819 , n9820 , n9821 , n9822 , n9823 , n9824 , n9825 , n9826 , n9827 , n9828 , n9829 , n9830 , n9831 , n9832 , n9833 , n9834 , n9835 , n9836 , n9837 , n9838 , n9839 , n9840 , n9841 , n9842 , n9843 , n9844 , n9845 , n9846 , n9847 , n9848 , n9849 , n9850 , n9851 , n9852 , n9853 , n9854 , n9855 , n9856 , n9857 , n9858 , n9859 , n9860 , n9861 , n9862 , n9863 , n9864 , n9865 , n9866 , n9867 , n9868 , n9869 , n9870 , n9871 , n9872 , n9873 , n9874 , n9875 , n9876 , n9877 , n9878 , n9879 , n9880 , n9881 , n9882 , n9883 , n9884 , n9885 , n9886 , n9887 , n9888 , n9889 , n9890 , n9891 , n9892 , n9893 , n9894 , n9895 , n9896 , n9897 , n9898 , n9899 , n9900 , n9901 , n9902 , n9903 , n9904 , n9905 , n9906 , n9907 , n9908 , n9909 , n9910 , n9911 , n9912 , n9913 , n9914 , n9915 , n9916 , n9917 , n9918 , n9919 , n9920 , n9921 , n9922 , n9923 , n9924 , n9925 , n9926 , n9927 , n9928 , n9929 , n9930 , n9931 , n9932 , n9933 , n9934 , n9935 , n9936 , n9937 , n9938 , n9939 , n9940 , n9941 , n9942 , n9943 , n9944 , n9945 , n9946 , n9947 , n9948 , n9949 , n9950 , n9951 , n9952 , n9953 , n9954 , n9955 , n9956 , n9957 , n9958 , n9959 , n9960 , n9961 , n9962 , n9963 , n9964 , n9965 , n9966 , n9967 , n9968 , n9969 , n9970 , n9971 , n9972 , n9973 , n9974 , n9975 , n9976 , n9977 , n9978 , n9979 , n9980 , n9981 , n9982 , n9983 , n9984 , n9985 , n9986 , n9987 , n9988 , n9989 , n9990 , n9991 , n9992 , n9993 , n9994 , n9995 , n9996 , n9997 , n9998 , n9999 , n10000 , n10001 , n10002 , n10003 , n10004 , n10005 , n10006 , n10007 , n10008 , n10009 , n10010 , n10011 , n10012 , n10013 , n10014 , n10015 , n10016 , n10017 , n10018 , n10019 , n10020 , n10021 , n10022 , n10023 , n10024 , n10025 , n10026 , n10027 , n10028 , n10029 , n10030 , n10031 , n10032 , n10033 , n10034 , n10035 , n10036 , n10037 , n10038 , n10039 , n10040 , n10041 , n10042 , n10043 , n10044 , n10045 , n10046 , n10047 , n10048 , n10049 , n10050 , n10051 , n10052 , n10053 , n10054 , n10055 , n10056 , n10057 , n10058 , n10059 , n10060 , n10061 , n10062 , n10063 , n10064 , n10065 , n10066 , n10067 , n10068 , n10069 , n10070 , n10071 , n10072 , n10073 , n10074 , n10075 , n10076 , n10077 , n10078 , n10079 , n10080 , n10081 , n10082 , n10083 , n10084 , n10085 , n10086 , n10087 , n10088 , n10089 , n10090 , n10091 , n10092 , n10093 , n10094 , n10095 , n10096 , n10097 , n10098 , n10099 , n10100 , n10101 , n10102 , n10103 , n10104 , n10105 , n10106 , n10107 , n10108 , n10109 , n10110 , n10111 , n10112 , n10113 , n10114 , n10115 , n10116 , n10117 , n10118 , n10119 , n10120 , n10121 , n10122 , n10123 , n10124 , n10125 , n10126 , n10127 , n10128 , n10129 , n10130 , n10131 , n10132 , n10133 , n10134 , n10135 , n10136 , n10137 , n10138 , n10139 , n10140 , n10141 , n10142 , n10143 , n10144 , n10145 , n10146 , n10147 , n10148 , n10149 , n10150 , n10151 , n10152 , n10153 , n10154 , n10155 , n10156 , n10157 , n10158 , n10159 , n10160 , n10161 , n10162 , n10163 , n10164 , n10165 , n10166 , n10167 , n10168 , n10169 , n10170 , n10171 , n10172 , n10173 , n10174 , n10175 , n10176 , n10177 , n10178 , n10179 , n10180 , n10181 , n10182 , n10183 , n10184 , n10185 , n10186 , n10187 , n10188 , n10189 , n10190 , n10191 , n10192 , n10193 , n10194 , n10195 , n10196 , n10197 , n10198 , n10199 , n10200 , n10201 , n10202 , n10203 , n10204 , n10205 , n10206 , n10207 , n10208 , n10209 , n10210 , n10211 , n10212 , n10213 , n10214 , n10215 , n10216 , n10217 , n10218 , n10219 , n10220 , n10221 , n10222 , n10223 , n10224 , n10225 , n10226 , n10227 , n10228 , n10229 , n10230 , n10231 , n10232 , n10233 , n10234 , n10235 , n10236 , n10237 , n10238 , n10239 , n10240 , n10241 , n10242 , n10243 , n10244 , n10245 , n10246 , n10247 , n10248 , n10249 , n10250 , n10251 , n10252 , n10253 , n10254 , n10255 , n10256 , n10257 , n10258 , n10259 , n10260 , n10261 , n10262 , n10263 , n10264 , n10265 , n10266 , n10267 , n10268 , n10269 , n10270 , n10271 , n10272 , n10273 , n10274 , n10275 , n10276 , n10277 , n10278 , n10279 , n10280 , n10281 , n10282 , n10283 , n10284 , n10285 , n10286 , n10287 , n10288 , n10289 , n10290 , n10291 , n10292 , n10293 , n10294 , n10295 , n10296 , n10297 , n10298 , n10299 , n10300 , n10301 , n10302 , n10303 , n10304 , n10305 , n10306 , n10307 , n10308 , n10309 , n10310 , n10311 , n10312 , n10313 , n10314 , n10315 , n10316 , n10317 , n10318 , n10319 , n10320 , n10321 , n10322 , n10323 , n10324 , n10325 , n10326 , n10327 , n10328 , n10329 , n10330 , n10331 , n10332 , n10333 , n10334 , n10335 , n10336 , n10337 , n10338 , n10339 , n10340 , n10341 , n10342 , n10343 , n10344 , n10345 , n10346 , n10347 , n10348 , n10349 , n10350 , n10351 , n10352 , n10353 , n10354 , n10355 , n10356 , n10357 , n10358 , n10359 , n10360 , n10361 , n10362 , n10363 , n10364 , n10365 , n10366 , n10367 , n10368 , n10369 , n10370 , n10371 , n10372 , n10373 , n10374 , n10375 , n10376 , n10377 , n10378 , n10379 , n10380 , n10381 , n10382 , n10383 , n10384 , n10385 , n10386 , n10387 , n10388 , n10389 , n10390 , n10391 , n10392 , n10393 , n10394 , n10395 , n10396 , n10397 , n10398 , n10399 , n10400 , n10401 , n10402 , n10403 , n10404 , n10405 , n10406 , n10407 , n10408 , n10409 , n10410 , n10411 , n10412 , n10413 , n10414 , n10415 , n10416 , n10417 , n10418 , n10419 , n10420 , n10421 , n10422 , n10423 , n10424 , n10425 , n10426 , n10427 , n10428 , n10429 , n10430 , n10431 , n10432 , n10433 , n10434 , n10435 , n10436 , n10437 , n10438 , n10439 , n10440 , n10441 , n10442 , n10443 , n10444 , n10445 , n10446 , n10447 , n10448 , n10449 , n10450 , n10451 , n10452 , n10453 , n10454 , n10455 , n10456 , n10457 , n10458 , n10459 , n10460 , n10461 , n10462 , n10463 , n10464 , n10465 , n10466 , n10467 , n10468 , n10469 , n10470 , n10471 , n10472 , n10473 , n10474 , n10475 , n10476 , n10477 , n10478 , n10479 , n10480 , n10481 , n10482 , n10483 , n10484 , n10485 , n10486 , n10487 , n10488 , n10489 , n10490 , n10491 , n10492 , n10493 , n10494 , n10495 , n10496 , n10497 , n10498 , n10499 , n10500 , n10501 , n10502 , n10503 , n10504 , n10505 , n10506 , n10507 , n10508 , n10509 , n10510 , n10511 , n10512 , n10513 , n10514 , n10515 , n10516 , n10517 , n10518 , n10519 , n10520 , n10521 , n10522 , n10523 , n10524 , n10525 , n10526 , n10527 , n10528 , n10529 , n10530 , n10531 , n10532 , n10533 , n10534 , n10535 , n10536 , n10537 , n10538 , n10539 , n10540 , n10541 , n10542 , n10543 , n10544 , n10545 , n10546 , n10547 , n10548 , n10549 , n10550 , n10551 , n10552 , n10553 , n10554 , n10555 , n10556 , n10557 , n10558 , n10559 , n10560 , n10561 , n10562 , n10563 , n10564 , n10565 , n10566 , n10567 , n10568 , n10569 , n10570 , n10571 , n10572 , n10573 , n10574 , n10575 , n10576 , n10577 , n10578 , n10579 , n10580 , n10581 , n10582 , n10583 , n10584 , n10585 , n10586 , n10587 , n10588 , n10589 , n10590 , n10591 , n10592 , n10593 , n10594 , n10595 , n10596 , n10597 , n10598 , n10599 , n10600 , n10601 , n10602 , n10603 , n10604 , n10605 , n10606 , n10607 , n10608 , n10609 , n10610 , n10611 , n10612 , n10613 , n10614 , n10615 , n10616 , n10617 , n10618 , n10619 , n10620 , n10621 , n10622 , n10623 , n10624 , n10625 , n10626 , n10627 , n10628 , n10629 , n10630 , n10631 , n10632 , n10633 , n10634 , n10635 , n10636 , n10637 , n10638 , n10639 , n10640 , n10641 , n10642 , n10643 , n10644 , n10645 , n10646 , n10647 , n10648 , n10649 , n10650 , n10651 , n10652 , n10653 , n10654 , n10655 , n10656 , n10657 , n10658 , n10659 , n10660 , n10661 , n10662 , n10663 , n10664 , n10665 , n10666 , n10667 , n10668 , n10669 , n10670 , n10671 , n10672 , n10673 , n10674 , n10675 , n10676 , n10677 , n10678 , n10679 , n10680 , n10681 , n10682 , n10683 , n10684 , n10685 , n10686 , n10687 , n10688 , n10689 , n10690 , n10691 , n10692 , n10693 , n10694 , n10695 , n10696 , n10697 , n10698 , n10699 , n10700 , n10701 , n10702 , n10703 , n10704 , n10705 , n10706 , n10707 , n10708 , n10709 , n10710 , n10711 , n10712 , n10713 , n10714 , n10715 , n10716 , n10717 , n10718 , n10719 , n10720 , n10721 , n10722 , n10723 , n10724 , n10725 , n10726 , n10727 , n10728 , n10729 , n10730 , n10731 , n10732 , n10733 , n10734 , n10735 , n10736 , n10737 , n10738 , n10739 , n10740 , n10741 , n10742 , n10743 , n10744 , n10745 , n10746 , n10747 , n10748 , n10749 , n10750 , n10751 , n10752 , n10753 , n10754 , n10755 , n10756 , n10757 , n10758 , n10759 , n10760 , n10761 , n10762 , n10763 , n10764 , n10765 , n10766 , n10767 , n10768 , n10769 , n10770 , n10771 , n10772 , n10773 , n10774 , n10775 , n10776 , n10777 , n10778 , n10779 , n10780 , n10781 , n10782 , n10783 , n10784 , n10785 , n10786 , n10787 , n10788 , n10789 , n10790 , n10791 , n10792 , n10793 , n10794 , n10795 , n10796 , n10797 , n10798 , n10799 , n10800 , n10801 , n10802 , n10803 , n10804 , n10805 , n10806 , n10807 , n10808 , n10809 , n10810 , n10811 , n10812 , n10813 , n10814 , n10815 , n10816 , n10817 , n10818 , n10819 , n10820 , n10821 , n10822 , n10823 , n10824 , n10825 , n10826 , n10827 , n10828 , n10829 , n10830 , n10831 , n10832 , n10833 , n10834 , n10835 , n10836 , n10837 , n10838 , n10839 , n10840 , n10841 , n10842 , n10843 , n10844 , n10845 , n10846 , n10847 , n10848 , n10849 , n10850 , n10851 , n10852 , n10853 , n10854 , n10855 , n10856 , n10857 , n10858 , n10859 , n10860 , n10861 , n10862 , n10863 , n10864 , n10865 , n10866 , n10867 , n10868 , n10869 , n10870 , n10871 , n10872 , n10873 , n10874 , n10875 , n10876 , n10877 , n10878 , n10879 , n10880 , n10881 , n10882 , n10883 , n10884 , n10885 , n10886 , n10887 , n10888 , n10889 , n10890 , n10891 , n10892 , n10893 , n10894 , n10895 , n10896 , n10897 , n10898 , n10899 , n10900 , n10901 , n10902 , n10903 , n10904 , n10905 , n10906 , n10907 , n10908 , n10909 , n10910 , n10911 , n10912 , n10913 , n10914 , n10915 , n10916 , n10917 , n10918 , n10919 , n10920 , n10921 , n10922 , n10923 , n10924 , n10925 , n10926 , n10927 , n10928 , n10929 , n10930 , n10931 , n10932 , n10933 , n10934 , n10935 , n10936 , n10937 , n10938 , n10939 , n10940 , n10941 , n10942 , n10943 , n10944 , n10945 , n10946 , n10947 , n10948 , n10949 , n10950 , n10951 , n10952 , n10953 , n10954 , n10955 , n10956 , n10957 , n10958 , n10959 , n10960 , n10961 , n10962 , n10963 , n10964 , n10965 , n10966 , n10967 , n10968 , n10969 , n10970 , n10971 , n10972 , n10973 , n10974 , n10975 , n10976 , n10977 , n10978 , n10979 , n10980 , n10981 , n10982 , n10983 , n10984 , n10985 , n10986 , n10987 , n10988 , n10989 , n10990 , n10991 , n10992 , n10993 , n10994 , n10995 , n10996 , n10997 , n10998 , n10999 , n11000 , n11001 , n11002 , n11003 , n11004 , n11005 , n11006 , n11007 , n11008 , n11009 , n11010 , n11011 , n11012 , n11013 , n11014 , n11015 , n11016 , n11017 , n11018 , n11019 , n11020 , n11021 , n11022 , n11023 , n11024 , n11025 , n11026 , n11027 , n11028 , n11029 , n11030 , n11031 , n11032 , n11033 , n11034 , n11035 , n11036 , n11037 , n11038 , n11039 , n11040 , n11041 , n11042 , n11043 , n11044 , n11045 , n11046 , n11047 , n11048 , n11049 , n11050 , n11051 , n11052 , n11053 , n11054 , n11055 , n11056 , n11057 , n11058 , n11059 , n11060 , n11061 , n11062 , n11063 , n11064 , n11065 , n11066 , n11067 , n11068 , n11069 , n11070 , n11071 , n11072 , n11073 , n11074 , n11075 , n11076 , n11077 , n11078 , n11079 , n11080 , n11081 , n11082 , n11083 , n11084 , n11085 , n11086 , n11087 , n11088 , n11089 , n11090 , n11091 , n11092 , n11093 , n11094 , n11095 , n11096 , n11097 , n11098 , n11099 , n11100 , n11101 , n11102 , n11103 , n11104 , n11105 , n11106 , n11107 , n11108 , n11109 , n11110 , n11111 , n11112 , n11113 , n11114 , n11115 , n11116 , n11117 , n11118 , n11119 , n11120 , n11121 , n11122 , n11123 , n11124 , n11125 , n11126 , n11127 , n11128 , n11129 , n11130 , n11131 , n11132 , n11133 , n11134 , n11135 , n11136 , n11137 , n11138 , n11139 , n11140 , n11141 , n11142 , n11143 , n11144 , n11145 , n11146 , n11147 , n11148 , n11149 , n11150 , n11151 , n11152 , n11153 , n11154 , n11155 , n11156 , n11157 , n11158 , n11159 , n11160 , n11161 , n11162 , n11163 , n11164 , n11165 , n11166 , n11167 , n11168 , n11169 , n11170 , n11171 , n11172 , n11173 , n11174 , n11175 , n11176 , n11177 , n11178 , n11179 , n11180 , n11181 , n11182 , n11183 , n11184 , n11185 , n11186 , n11187 , n11188 , n11189 , n11190 , n11191 , n11192 , n11193 , n11194 , n11195 , n11196 , n11197 , n11198 , n11199 , n11200 , n11201 , n11202 , n11203 , n11204 , n11205 , n11206 , n11207 , n11208 , n11209 , n11210 , n11211 , n11212 , n11213 , n11214 , n11215 , n11216 , n11217 , n11218 , n11219 , n11220 , n11221 , n11222 , n11223 , n11224 , n11225 , n11226 , n11227 , n11228 , n11229 , n11230 , n11231 , n11232 , n11233 , n11234 , n11235 , n11236 , n11237 , n11238 , n11239 , n11240 , n11241 , n11242 , n11243 , n11244 , n11245 , n11246 , n11247 , n11248 , n11249 , n11250 , n11251 , n11252 , n11253 , n11254 , n11255 , n11256 , n11257 , n11258 , n11259 , n11260 , n11261 , n11262 , n11263 , n11264 , n11265 , n11266 , n11267 , n11268 , n11269 , n11270 , n11271 , n11272 , n11273 , n11274 , n11275 , n11276 , n11277 , n11278 , n11279 , n11280 , n11281 , n11282 , n11283 , n11284 , n11285 , n11286 , n11287 , n11288 , n11289 , n11290 , n11291 , n11292 , n11293 , n11294 , n11295 , n11296 , n11297 , n11298 , n11299 , n11300 , n11301 , n11302 , n11303 , n11304 , n11305 , n11306 , n11307 , n11308 , n11309 , n11310 , n11311 , n11312 , n11313 , n11314 , n11315 , n11316 , n11317 , n11318 , n11319 , n11320 , n11321 , n11322 , n11323 , n11324 , n11325 , n11326 , n11327 , n11328 , n11329 , n11330 , n11331 , n11332 , n11333 , n11334 , n11335 , n11336 , n11337 , n11338 , n11339 , n11340 , n11341 , n11342 , n11343 , n11344 , n11345 , n11346 , n11347 , n11348 , n11349 , n11350 , n11351 , n11352 , n11353 , n11354 , n11355 , n11356 , n11357 , n11358 , n11359 , n11360 , n11361 , n11362 , n11363 , n11364 , n11365 , n11366 , n11367 , n11368 , n11369 , n11370 , n11371 , n11372 , n11373 , n11374 , n11375 , n11376 , n11377 , n11378 , n11379 , n11380 , n11381 , n11382 , n11383 , n11384 , n11385 , n11386 , n11387 , n11388 , n11389 , n11390 , n11391 , n11392 , n11393 , n11394 , n11395 , n11396 , n11397 , n11398 , n11399 , n11400 , n11401 , n11402 , n11403 , n11404 , n11405 , n11406 , n11407 , n11408 , n11409 , n11410 , n11411 , n11412 , n11413 , n11414 , n11415 , n11416 , n11417 , n11418 , n11419 , n11420 , n11421 , n11422 , n11423 , n11424 , n11425 , n11426 , n11427 , n11428 , n11429 , n11430 , n11431 , n11432 , n11433 , n11434 , n11435 , n11436 , n11437 , n11438 , n11439 , n11440 , n11441 , n11442 , n11443 , n11444 , n11445 , n11446 , n11447 , n11448 , n11449 , n11450 , n11451 , n11452 , n11453 , n11454 , n11455 , n11456 , n11457 , n11458 , n11459 , n11460 , n11461 , n11462 , n11463 , n11464 , n11465 , n11466 , n11467 , n11468 , n11469 , n11470 , n11471 , n11472 , n11473 , n11474 , n11475 , n11476 , n11477 , n11478 , n11479 , n11480 , n11481 , n11482 , n11483 , n11484 , n11485 , n11486 , n11487 , n11488 , n11489 , n11490 , n11491 , n11492 , n11493 , n11494 , n11495 , n11496 , n11497 , n11498 , n11499 , n11500 , n11501 , n11502 , n11503 , n11504 , n11505 , n11506 , n11507 , n11508 , n11509 , n11510 , n11511 , n11512 , n11513 , n11514 , n11515 , n11516 , n11517 , n11518 , n11519 , n11520 , n11521 , n11522 , n11523 , n11524 , n11525 , n11526 , n11527 , n11528 , n11529 , n11530 , n11531 , n11532 , n11533 , n11534 , n11535 , n11536 , n11537 , n11538 , n11539 , n11540 , n11541 , n11542 , n11543 , n11544 , n11545 , n11546 , n11547 , n11548 , n11549 , n11550 , n11551 , n11552 , n11553 , n11554 , n11555 , n11556 , n11557 , n11558 , n11559 , n11560 , n11561 , n11562 , n11563 , n11564 , n11565 , n11566 , n11567 , n11568 , n11569 , n11570 , n11571 , n11572 , n11573 , n11574 , n11575 , n11576 , n11577 , n11578 , n11579 , n11580 , n11581 , n11582 , n11583 , n11584 , n11585 , n11586 , n11587 , n11588 , n11589 , n11590 , n11591 , n11592 , n11593 , n11594 , n11595 , n11596 , n11597 , n11598 , n11599 , n11600 , n11601 , n11602 , n11603 , n11604 , n11605 , n11606 , n11607 , n11608 , n11609 , n11610 , n11611 , n11612 , n11613 , n11614 , n11615 , n11616 , n11617 , n11618 , n11619 , n11620 , n11621 , n11622 , n11623 , n11624 , n11625 , n11626 , n11627 , n11628 , n11629 , n11630 , n11631 , n11632 , n11633 , n11634 , n11635 , n11636 , n11637 , n11638 , n11639 , n11640 , n11641 , n11642 , n11643 , n11644 , n11645 , n11646 , n11647 , n11648 , n11649 , n11650 , n11651 , n11652 , n11653 , n11654 , n11655 , n11656 , n11657 , n11658 , n11659 , n11660 , n11661 , n11662 , n11663 , n11664 , n11665 , n11666 , n11667 , n11668 , n11669 , n11670 , n11671 , n11672 , n11673 , n11674 , n11675 , n11676 , n11677 , n11678 , n11679 , n11680 , n11681 , n11682 , n11683 , n11684 , n11685 , n11686 , n11687 , n11688 , n11689 , n11690 , n11691 , n11692 , n11693 , n11694 , n11695 , n11696 , n11697 , n11698 , n11699 , n11700 , n11701 , n11702 , n11703 , n11704 , n11705 , n11706 , n11707 , n11708 , n11709 , n11710 , n11711 , n11712 , n11713 , n11714 , n11715 , n11716 , n11717 , n11718 , n11719 , n11720 , n11721 , n11722 , n11723 , n11724 , n11725 , n11726 , n11727 , n11728 , n11729 , n11730 , n11731 , n11732 , n11733 , n11734 , n11735 , n11736 , n11737 , n11738 , n11739 , n11740 , n11741 , n11742 , n11743 , n11744 , n11745 , n11746 , n11747 , n11748 , n11749 , n11750 , n11751 , n11752 , n11753 , n11754 , n11755 , n11756 , n11757 , n11758 , n11759 , n11760 , n11761 , n11762 , n11763 , n11764 , n11765 , n11766 , n11767 , n11768 , n11769 , n11770 , n11771 , n11772 , n11773 , n11774 , n11775 , n11776 , n11777 , n11778 , n11779 , n11780 , n11781 , n11782 , n11783 , n11784 , n11785 , n11786 , n11787 , n11788 , n11789 , n11790 , n11791 , n11792 , n11793 , n11794 , n11795 , n11796 , n11797 , n11798 , n11799 , n11800 , n11801 , n11802 , n11803 , n11804 , n11805 , n11806 , n11807 , n11808 , n11809 , n11810 , n11811 , n11812 , n11813 , n11814 , n11815 , n11816 , n11817 , n11818 , n11819 , n11820 , n11821 , n11822 , n11823 , n11824 , n11825 , n11826 , n11827 , n11828 , n11829 , n11830 , n11831 , n11832 , n11833 , n11834 , n11835 , n11836 , n11837 , n11838 , n11839 , n11840 , n11841 , n11842 , n11843 , n11844 , n11845 , n11846 , n11847 , n11848 , n11849 , n11850 , n11851 , n11852 , n11853 , n11854 , n11855 , n11856 , n11857 , n11858 , n11859 , n11860 , n11861 , n11862 , n11863 , n11864 , n11865 , n11866 , n11867 , n11868 , n11869 , n11870 , n11871 , n11872 , n11873 , n11874 , n11875 , n11876 , n11877 , n11878 , n11879 , n11880 , n11881 , n11882 , n11883 , n11884 , n11885 , n11886 , n11887 , n11888 , n11889 , n11890 , n11891 , n11892 , n11893 , n11894 , n11895 , n11896 , n11897 , n11898 , n11899 , n11900 , n11901 , n11902 , n11903 , n11904 , n11905 , n11906 , n11907 , n11908 , n11909 , n11910 , n11911 , n11912 , n11913 , n11914 , n11915 , n11916 , n11917 , n11918 , n11919 , n11920 , n11921 , n11922 , n11923 , n11924 , n11925 , n11926 , n11927 , n11928 , n11929 , n11930 , n11931 , n11932 , n11933 , n11934 , n11935 , n11936 , n11937 , n11938 , n11939 , n11940 , n11941 , n11942 , n11943 , n11944 , n11945 , n11946 , n11947 , n11948 , n11949 , n11950 , n11951 , n11952 , n11953 , n11954 , n11955 , n11956 , n11957 , n11958 , n11959 , n11960 , n11961 , n11962 , n11963 , n11964 , n11965 , n11966 , n11967 , n11968 , n11969 , n11970 , n11971 , n11972 , n11973 , n11974 , n11975 , n11976 , n11977 , n11978 , n11979 , n11980 , n11981 , n11982 , n11983 , n11984 , n11985 , n11986 , n11987 , n11988 , n11989 , n11990 , n11991 , n11992 , n11993 , n11994 , n11995 , n11996 , n11997 , n11998 , n11999 , n12000 , n12001 , n12002 , n12003 , n12004 , n12005 , n12006 , n12007 , n12008 , n12009 , n12010 , n12011 , n12012 , n12013 , n12014 , n12015 , n12016 , n12017 , n12018 , n12019 , n12020 , n12021 , n12022 , n12023 , n12024 , n12025 , n12026 , n12027 , n12028 , n12029 , n12030 , n12031 , n12032 , n12033 , n12034 , n12035 , n12036 , n12037 , n12038 , n12039 , n12040 , n12041 , n12042 , n12043 , n12044 , n12045 , n12046 , n12047 , n12048 , n12049 , n12050 , n12051 , n12052 , n12053 , n12054 , n12055 , n12056 , n12057 , n12058 , n12059 , n12060 , n12061 , n12062 , n12063 , n12064 , n12065 , n12066 , n12067 , n12068 , n12069 , n12070 , n12071 , n12072 , n12073 , n12074 , n12075 , n12076 , n12077 , n12078 , n12079 , n12080 , n12081 , n12082 , n12083 , n12084 , n12085 , n12086 , n12087 , n12088 , n12089 , n12090 , n12091 , n12092 , n12093 , n12094 , n12095 , n12096 , n12097 , n12098 , n12099 , n12100 , n12101 , n12102 , n12103 , n12104 , n12105 , n12106 , n12107 , n12108 , n12109 , n12110 , n12111 , n12112 , n12113 , n12114 , n12115 , n12116 , n12117 , n12118 , n12119 , n12120 , n12121 , n12122 , n12123 , n12124 , n12125 , n12126 , n12127 , n12128 , n12129 , n12130 , n12131 , n12132 , n12133 , n12134 , n12135 , n12136 , n12137 , n12138 , n12139 , n12140 , n12141 , n12142 , n12143 , n12144 , n12145 , n12146 , n12147 , n12148 , n12149 , n12150 , n12151 , n12152 , n12153 , n12154 , n12155 , n12156 , n12157 , n12158 , n12159 , n12160 , n12161 , n12162 , n12163 , n12164 , n12165 , n12166 , n12167 , n12168 , n12169 , n12170 , n12171 , n12172 , n12173 , n12174 , n12175 , n12176 , n12177 , n12178 , n12179 , n12180 , n12181 , n12182 , n12183 , n12184 , n12185 , n12186 , n12187 , n12188 , n12189 , n12190 , n12191 , n12192 , n12193 , n12194 , n12195 , n12196 , n12197 , n12198 , n12199 , n12200 , n12201 , n12202 , n12203 , n12204 , n12205 , n12206 , n12207 , n12208 , n12209 , n12210 , n12211 , n12212 , n12213 , n12214 , n12215 , n12216 , n12217 , n12218 , n12219 , n12220 , n12221 , n12222 , n12223 , n12224 , n12225 , n12226 , n12227 , n12228 , n12229 , n12230 , n12231 , n12232 , n12233 , n12234 , n12235 , n12236 , n12237 , n12238 , n12239 , n12240 , n12241 , n12242 , n12243 , n12244 , n12245 , n12246 , n12247 , n12248 , n12249 , n12250 , n12251 , n12252 , n12253 , n12254 , n12255 , n12256 , n12257 , n12258 , n12259 , n12260 , n12261 , n12262 , n12263 , n12264 , n12265 , n12266 , n12267 , n12268 , n12269 , n12270 , n12271 , n12272 , n12273 , n12274 , n12275 , n12276 , n12277 , n12278 , n12279 , n12280 , n12281 , n12282 , n12283 , n12284 , n12285 , n12286 , n12287 , n12288 , n12289 , n12290 , n12291 , n12292 , n12293 , n12294 , n12295 , n12296 , n12297 , n12298 , n12299 , n12300 , n12301 , n12302 , n12303 , n12304 , n12305 , n12306 , n12307 , n12308 , n12309 , n12310 , n12311 , n12312 , n12313 , n12314 , n12315 , n12316 , n12317 , n12318 , n12319 , n12320 , n12321 , n12322 , n12323 , n12324 , n12325 , n12326 , n12327 , n12328 , n12329 , n12330 , n12331 , n12332 , n12333 , n12334 , n12335 , n12336 , n12337 , n12338 , n12339 , n12340 , n12341 , n12342 , n12343 , n12344 , n12345 , n12346 , n12347 , n12348 , n12349 , n12350 , n12351 , n12352 , n12353 , n12354 , n12355 , n12356 , n12357 , n12358 , n12359 , n12360 , n12361 , n12362 , n12363 , n12364 , n12365 , n12366 , n12367 , n12368 , n12369 , n12370 , n12371 , n12372 , n12373 , n12374 , n12375 , n12376 , n12377 , n12378 , n12379 , n12380 , n12381 , n12382 , n12383 , n12384 , n12385 , n12386 , n12387 , n12388 , n12389 , n12390 , n12391 , n12392 , n12393 , n12394 , n12395 , n12396 , n12397 , n12398 , n12399 , n12400 , n12401 , n12402 , n12403 , n12404 , n12405 , n12406 , n12407 , n12408 , n12409 , n12410 , n12411 , n12412 , n12413 , n12414 , n12415 , n12416 , n12417 , n12418 , n12419 , n12420 , n12421 , n12422 , n12423 , n12424 , n12425 , n12426 , n12427 , n12428 , n12429 , n12430 , n12431 , n12432 , n12433 , n12434 , n12435 , n12436 , n12437 , n12438 , n12439 , n12440 , n12441 , n12442 , n12443 , n12444 , n12445 , n12446 , n12447 , n12448 , n12449 , n12450 , n12451 , n12452 , n12453 , n12454 , n12455 , n12456 , n12457 , n12458 , n12459 , n12460 , n12461 , n12462 , n12463 , n12464 , n12465 , n12466 , n12467 , n12468 , n12469 , n12470 , n12471 , n12472 , n12473 , n12474 , n12475 , n12476 , n12477 , n12478 , n12479 , n12480 , n12481 , n12482 , n12483 , n12484 , n12485 , n12486 , n12487 , n12488 , n12489 , n12490 , n12491 , n12492 , n12493 , n12494 , n12495 , n12496 , n12497 , n12498 , n12499 , n12500 , n12501 , n12502 , n12503 , n12504 , n12505 , n12506 , n12507 , n12508 , n12509 , n12510 , n12511 , n12512 , n12513 , n12514 , n12515 , n12516 , n12517 , n12518 , n12519 , n12520 , n12521 , n12522 , n12523 , n12524 , n12525 , n12526 , n12527 , n12528 , n12529 , n12530 , n12531 , n12532 , n12533 , n12534 , n12535 , n12536 , n12537 , n12538 , n12539 , n12540 , n12541 , n12542 , n12543 , n12544 , n12545 , n12546 , n12547 , n12548 , n12549 , n12550 , n12551 , n12552 , n12553 , n12554 , n12555 , n12556 , n12557 , n12558 , n12559 , n12560 , n12561 , n12562 , n12563 , n12564 , n12565 , n12566 , n12567 , n12568 , n12569 , n12570 , n12571 , n12572 , n12573 , n12574 , n12575 , n12576 , n12577 , n12578 , n12579 , n12580 , n12581 , n12582 , n12583 , n12584 , n12585 , n12586 , n12587 , n12588 , n12589 , n12590 , n12591 , n12592 , n12593 , n12594 , n12595 , n12596 , n12597 , n12598 , n12599 , n12600 , n12601 , n12602 , n12603 , n12604 , n12605 , n12606 , n12607 , n12608 , n12609 , n12610 , n12611 , n12612 , n12613 , n12614 , n12615 , n12616 , n12617 , n12618 , n12619 , n12620 , n12621 , n12622 , n12623 , n12624 , n12625 , n12626 , n12627 , n12628 , n12629 , n12630 , n12631 , n12632 , n12633 , n12634 , n12635 , n12636 , n12637 , n12638 , n12639 , n12640 , n12641 , n12642 , n12643 , n12644 , n12645 , n12646 , n12647 , n12648 , n12649 , n12650 , n12651 , n12652 , n12653 , n12654 , n12655 , n12656 , n12657 , n12658 , n12659 , n12660 , n12661 , n12662 , n12663 , n12664 , n12665 , n12666 , n12667 , n12668 , n12669 , n12670 , n12671 , n12672 , n12673 , n12674 , n12675 , n12676 , n12677 , n12678 , n12679 , n12680 , n12681 , n12682 , n12683 , n12684 , n12685 , n12686 , n12687 , n12688 , n12689 , n12690 , n12691 , n12692 , n12693 , n12694 , n12695 , n12696 , n12697 , n12698 , n12699 , n12700 , n12701 , n12702 , n12703 , n12704 , n12705 , n12706 , n12707 , n12708 , n12709 , n12710 , n12711 , n12712 , n12713 , n12714 , n12715 , n12716 , n12717 , n12718 , n12719 , n12720 , n12721 , n12722 , n12723 , n12724 , n12725 , n12726 , n12727 , n12728 , n12729 , n12730 , n12731 , n12732 , n12733 , n12734 , n12735 , n12736 , n12737 , n12738 , n12739 , n12740 , n12741 , n12742 , n12743 , n12744 , n12745 , n12746 , n12747 , n12748 , n12749 , n12750 , n12751 , n12752 , n12753 , n12754 , n12755 , n12756 , n12757 , n12758 , n12759 , n12760 , n12761 , n12762 , n12763 , n12764 , n12765 , n12766 , n12767 , n12768 , n12769 , n12770 , n12771 , n12772 , n12773 , n12774 , n12775 , n12776 , n12777 , n12778 , n12779 , n12780 , n12781 , n12782 , n12783 , n12784 , n12785 , n12786 , n12787 , n12788 , n12789 , n12790 , n12791 , n12792 , n12793 , n12794 , n12795 , n12796 , n12797 , n12798 , n12799 , n12800 , n12801 , n12802 , n12803 , n12804 , n12805 , n12806 , n12807 , n12808 , n12809 , n12810 , n12811 , n12812 , n12813 , n12814 , n12815 , n12816 , n12817 , n12818 , n12819 , n12820 , n12821 , n12822 , n12823 , n12824 , n12825 , n12826 , n12827 , n12828 , n12829 , n12830 , n12831 , n12832 , n12833 , n12834 , n12835 , n12836 , n12837 , n12838 , n12839 , n12840 , n12841 , n12842 , n12843 , n12844 , n12845 , n12846 , n12847 , n12848 , n12849 , n12850 , n12851 , n12852 , n12853 , n12854 , n12855 , n12856 , n12857 , n12858 , n12859 , n12860 , n12861 , n12862 , n12863 , n12864 , n12865 , n12866 , n12867 , n12868 , n12869 , n12870 , n12871 , n12872 , n12873 , n12874 , n12875 , n12876 , n12877 , n12878 , n12879 , n12880 , n12881 , n12882 , n12883 , n12884 , n12885 , n12886 , n12887 , n12888 , n12889 , n12890 , n12891 , n12892 , n12893 , n12894 , n12895 , n12896 , n12897 , n12898 , n12899 , n12900 , n12901 , n12902 , n12903 , n12904 , n12905 , n12906 , n12907 , n12908 , n12909 , n12910 , n12911 , n12912 , n12913 , n12914 , n12915 , n12916 , n12917 , n12918 , n12919 , n12920 , n12921 , n12922 , n12923 , n12924 , n12925 , n12926 , n12927 , n12928 , n12929 , n12930 , n12931 , n12932 , n12933 , n12934 , n12935 , n12936 , n12937 , n12938 , n12939 , n12940 , n12941 , n12942 , n12943 , n12944 , n12945 , n12946 , n12947 , n12948 , n12949 , n12950 , n12951 , n12952 , n12953 , n12954 , n12955 , n12956 , n12957 , n12958 , n12959 , n12960 , n12961 , n12962 , n12963 , n12964 , n12965 , n12966 , n12967 , n12968 , n12969 , n12970 , n12971 , n12972 , n12973 , n12974 , n12975 , n12976 , n12977 , n12978 , n12979 , n12980 , n12981 , n12982 , n12983 , n12984 , n12985 , n12986 , n12987 , n12988 , n12989 , n12990 , n12991 , n12992 , n12993 , n12994 , n12995 , n12996 , n12997 , n12998 , n12999 , n13000 , n13001 , n13002 , n13003 , n13004 , n13005 , n13006 , n13007 , n13008 , n13009 , n13010 , n13011 , n13012 , n13013 , n13014 , n13015 , n13016 , n13017 , n13018 , n13019 , n13020 , n13021 , n13022 , n13023 , n13024 , n13025 , n13026 , n13027 , n13028 , n13029 , n13030 , n13031 , n13032 , n13033 , n13034 , n13035 , n13036 , n13037 , n13038 , n13039 , n13040 , n13041 , n13042 , n13043 , n13044 , n13045 , n13046 , n13047 , n13048 , n13049 , n13050 , n13051 , n13052 , n13053 , n13054 , n13055 , n13056 , n13057 , n13058 , n13059 , n13060 , n13061 , n13062 , n13063 , n13064 , n13065 , n13066 , n13067 , n13068 , n13069 , n13070 , n13071 , n13072 , n13073 , n13074 , n13075 , n13076 , n13077 , n13078 , n13079 , n13080 , n13081 , n13082 , n13083 , n13084 , n13085 , n13086 , n13087 , n13088 , n13089 , n13090 , n13091 , n13092 , n13093 , n13094 , n13095 , n13096 , n13097 , n13098 , n13099 , n13100 , n13101 , n13102 , n13103 , n13104 , n13105 , n13106 , n13107 , n13108 , n13109 , n13110 , n13111 , n13112 , n13113 , n13114 , n13115 , n13116 , n13117 , n13118 , n13119 , n13120 , n13121 , n13122 , n13123 , n13124 , n13125 , n13126 , n13127 , n13128 , n13129 , n13130 , n13131 , n13132 , n13133 , n13134 , n13135 , n13136 , n13137 , n13138 , n13139 , n13140 , n13141 , n13142 , n13143 , n13144 , n13145 , n13146 , n13147 , n13148 , n13149 , n13150 , n13151 , n13152 , n13153 , n13154 , n13155 , n13156 , n13157 , n13158 , n13159 , n13160 , n13161 , n13162 , n13163 , n13164 , n13165 , n13166 , n13167 , n13168 , n13169 , n13170 , n13171 , n13172 , n13173 , n13174 , n13175 , n13176 , n13177 , n13178 , n13179 , n13180 , n13181 , n13182 , n13183 , n13184 , n13185 , n13186 , n13187 , n13188 , n13189 , n13190 , n13191 , n13192 , n13193 , n13194 , n13195 , n13196 , n13197 , n13198 , n13199 , n13200 , n13201 , n13202 , n13203 , n13204 , n13205 , n13206 , n13207 , n13208 , n13209 , n13210 , n13211 , n13212 , n13213 , n13214 , n13215 , n13216 , n13217 , n13218 , n13219 , n13220 , n13221 , n13222 , n13223 , n13224 , n13225 , n13226 , n13227 , n13228 , n13229 , n13230 , n13231 , n13232 , n13233 , n13234 , n13235 , n13236 , n13237 , n13238 , n13239 , n13240 , n13241 , n13242 , n13243 , n13244 , n13245 , n13246 , n13247 , n13248 , n13249 , n13250 , n13251 , n13252 , n13253 , n13254 , n13255 , n13256 , n13257 , n13258 , n13259 , n13260 , n13261 , n13262 , n13263 , n13264 , n13265 , n13266 , n13267 , n13268 , n13269 , n13270 , n13271 , n13272 , n13273 , n13274 , n13275 , n13276 , n13277 , n13278 , n13279 , n13280 , n13281 , n13282 , n13283 , n13284 , n13285 , n13286 , n13287 , n13288 , n13289 , n13290 , n13291 , n13292 , n13293 , n13294 , n13295 , n13296 , n13297 , n13298 , n13299 , n13300 , n13301 , n13302 , n13303 , n13304 , n13305 , n13306 , n13307 , n13308 , n13309 , n13310 , n13311 , n13312 , n13313 , n13314 , n13315 , n13316 , n13317 , n13318 , n13319 , n13320 , n13321 , n13322 , n13323 , n13324 , n13325 , n13326 , n13327 , n13328 , n13329 , n13330 , n13331 , n13332 , n13333 , n13334 , n13335 , n13336 , n13337 , n13338 , n13339 , n13340 , n13341 , n13342 , n13343 , n13344 , n13345 , n13346 , n13347 , n13348 , n13349 , n13350 , n13351 , n13352 , n13353 , n13354 , n13355 , n13356 , n13357 , n13358 , n13359 , n13360 , n13361 , n13362 , n13363 , n13364 , n13365 , n13366 , n13367 , n13368 , n13369 , n13370 , n13371 , n13372 , n13373 , n13374 , n13375 , n13376 , n13377 , n13378 , n13379 , n13380 , n13381 , n13382 , n13383 , n13384 , n13385 , n13386 , n13387 , n13388 , n13389 , n13390 , n13391 , n13392 , n13393 , n13394 , n13395 , n13396 , n13397 , n13398 , n13399 , n13400 , n13401 , n13402 , n13403 , n13404 , n13405 , n13406 , n13407 , n13408 , n13409 , n13410 , n13411 , n13412 , n13413 , n13414 , n13415 , n13416 , n13417 , n13418 , n13419 , n13420 , n13421 , n13422 , n13423 , n13424 , n13425 , n13426 , n13427 , n13428 , n13429 , n13430 , n13431 , n13432 , n13433 , n13434 , n13435 , n13436 , n13437 , n13438 , n13439 , n13440 , n13441 , n13442 , n13443 , n13444 , n13445 , n13446 , n13447 , n13448 , n13449 , n13450 , n13451 , n13452 , n13453 , n13454 , n13455 , n13456 , n13457 , n13458 , n13459 , n13460 , n13461 , n13462 , n13463 , n13464 , n13465 , n13466 , n13467 , n13468 , n13469 , n13470 , n13471 , n13472 , n13473 , n13474 , n13475 , n13476 , n13477 , n13478 , n13479 , n13480 , n13481 , n13482 , n13483 , n13484 , n13485 , n13486 , n13487 , n13488 , n13489 , n13490 , n13491 , n13492 , n13493 , n13494 , n13495 , n13496 , n13497 , n13498 , n13499 , n13500 , n13501 , n13502 , n13503 , n13504 , n13505 , n13506 , n13507 , n13508 , n13509 , n13510 , n13511 , n13512 , n13513 , n13514 , n13515 , n13516 , n13517 , n13518 , n13519 , n13520 , n13521 , n13522 , n13523 , n13524 , n13525 , n13526 , n13527 , n13528 , n13529 , n13530 , n13531 , n13532 , n13533 , n13534 , n13535 , n13536 , n13537 , n13538 , n13539 , n13540 , n13541 , n13542 , n13543 , n13544 , n13545 , n13546 , n13547 , n13548 , n13549 , n13550 , n13551 , n13552 , n13553 , n13554 , n13555 , n13556 , n13557 , n13558 , n13559 , n13560 , n13561 , n13562 , n13563 , n13564 , n13565 , n13566 , n13567 , n13568 , n13569 , n13570 , n13571 , n13572 , n13573 , n13574 , n13575 , n13576 , n13577 , n13578 , n13579 , n13580 , n13581 , n13582 , n13583 , n13584 , n13585 , n13586 , n13587 , n13588 , n13589 , n13590 , n13591 , n13592 , n13593 , n13594 , n13595 , n13596 , n13597 , n13598 , n13599 , n13600 , n13601 , n13602 , n13603 , n13604 , n13605 , n13606 , n13607 , n13608 , n13609 , n13610 , n13611 , n13612 , n13613 , n13614 , n13615 , n13616 , n13617 , n13618 , n13619 , n13620 , n13621 , n13622 , n13623 , n13624 , n13625 , n13626 , n13627 , n13628 , n13629 , n13630 , n13631 , n13632 , n13633 , n13634 , n13635 , n13636 , n13637 , n13638 , n13639 , n13640 , n13641 , n13642 , n13643 , n13644 , n13645 , n13646 , n13647 , n13648 , n13649 , n13650 , n13651 , n13652 , n13653 , n13654 , n13655 , n13656 , n13657 , n13658 , n13659 , n13660 , n13661 , n13662 , n13663 , n13664 , n13665 , n13666 , n13667 , n13668 , n13669 , n13670 , n13671 , n13672 , n13673 , n13674 , n13675 , n13676 , n13677 , n13678 , n13679 , n13680 , n13681 , n13682 , n13683 , n13684 , n13685 , n13686 , n13687 , n13688 , n13689 , n13690 , n13691 , n13692 , n13693 , n13694 , n13695 , n13696 , n13697 , n13698 , n13699 , n13700 , n13701 , n13702 , n13703 , n13704 , n13705 , n13706 , n13707 , n13708 , n13709 , n13710 , n13711 , n13712 , n13713 , n13714 , n13715 , n13716 , n13717 , n13718 , n13719 , n13720 , n13721 , n13722 , n13723 , n13724 , n13725 , n13726 , n13727 , n13728 , n13729 , n13730 , n13731 , n13732 , n13733 , n13734 , n13735 , n13736 , n13737 , n13738 , n13739 , n13740 , n13741 , n13742 , n13743 , n13744 , n13745 , n13746 , n13747 , n13748 , n13749 , n13750 , n13751 , n13752 , n13753 , n13754 , n13755 , n13756 , n13757 , n13758 , n13759 , n13760 , n13761 , n13762 , n13763 , n13764 , n13765 , n13766 , n13767 , n13768 , n13769 , n13770 , n13771 , n13772 , n13773 , n13774 , n13775 , n13776 , n13777 , n13778 , n13779 , n13780 , n13781 , n13782 , n13783 , n13784 , n13785 , n13786 , n13787 , n13788 , n13789 , n13790 , n13791 , n13792 , n13793 , n13794 , n13795 , n13796 , n13797 , n13798 , n13799 , n13800 , n13801 , n13802 , n13803 , n13804 , n13805 , n13806 , n13807 , n13808 , n13809 , n13810 , n13811 , n13812 , n13813 , n13814 , n13815 , n13816 , n13817 , n13818 , n13819 , n13820 , n13821 , n13822 , n13823 , n13824 , n13825 , n13826 , n13827 , n13828 , n13829 , n13830 , n13831 , n13832 , n13833 , n13834 , n13835 , n13836 , n13837 , n13838 , n13839 , n13840 , n13841 , n13842 , n13843 , n13844 , n13845 , n13846 , n13847 , n13848 , n13849 , n13850 , n13851 , n13852 , n13853 , n13854 , n13855 , n13856 , n13857 , n13858 , n13859 , n13860 , n13861 , n13862 , n13863 , n13864 , n13865 , n13866 , n13867 , n13868 , n13869 , n13870 , n13871 , n13872 , n13873 , n13874 , n13875 , n13876 , n13877 , n13878 , n13879 , n13880 , n13881 , n13882 , n13883 , n13884 , n13885 , n13886 , n13887 , n13888 , n13889 , n13890 , n13891 , n13892 , n13893 , n13894 , n13895 , n13896 , n13897 , n13898 , n13899 , n13900 , n13901 , n13902 , n13903 , n13904 , n13905 , n13906 , n13907 , n13908 , n13909 , n13910 , n13911 , n13912 , n13913 , n13914 , n13915 , n13916 , n13917 , n13918 , n13919 , n13920 , n13921 , n13922 , n13923 , n13924 , n13925 , n13926 , n13927 , n13928 , n13929 , n13930 , n13931 , n13932 , n13933 , n13934 , n13935 , n13936 , n13937 , n13938 , n13939 , n13940 , n13941 , n13942 , n13943 , n13944 , n13945 , n13946 , n13947 , n13948 , n13949 , n13950 , n13951 , n13952 , n13953 , n13954 , n13955 , n13956 , n13957 , n13958 , n13959 , n13960 , n13961 , n13962 , n13963 , n13964 , n13965 , n13966 , n13967 , n13968 , n13969 , n13970 , n13971 , n13972 , n13973 , n13974 , n13975 , n13976 , n13977 , n13978 , n13979 , n13980 , n13981 , n13982 , n13983 , n13984 , n13985 , n13986 , n13987 , n13988 , n13989 , n13990 , n13991 , n13992 , n13993 , n13994 , n13995 , n13996 , n13997 , n13998 , n13999 , n14000 , n14001 , n14002 , n14003 , n14004 , n14005 , n14006 , n14007 , n14008 , n14009 , n14010 , n14011 , n14012 , n14013 , n14014 , n14015 , n14016 , n14017 , n14018 , n14019 , n14020 , n14021 , n14022 , n14023 , n14024 , n14025 , n14026 , n14027 , n14028 , n14029 , n14030 , n14031 , n14032 , n14033 , n14034 , n14035 , n14036 , n14037 , n14038 , n14039 , n14040 , n14041 , n14042 , n14043 , n14044 , n14045 , n14046 , n14047 , n14048 , n14049 , n14050 , n14051 , n14052 , n14053 , n14054 , n14055 , n14056 , n14057 , n14058 , n14059 , n14060 , n14061 , n14062 , n14063 , n14064 , n14065 , n14066 , n14067 , n14068 , n14069 , n14070 , n14071 , n14072 , n14073 , n14074 , n14075 , n14076 , n14077 , n14078 , n14079 , n14080 , n14081 , n14082 , n14083 , n14084 , n14085 , n14086 , n14087 , n14088 , n14089 , n14090 , n14091 , n14092 , n14093 , n14094 , n14095 , n14096 , n14097 , n14098 , n14099 , n14100 , n14101 , n14102 , n14103 , n14104 , n14105 , n14106 , n14107 , n14108 , n14109 , n14110 , n14111 , n14112 , n14113 , n14114 , n14115 , n14116 , n14117 , n14118 , n14119 , n14120 , n14121 , n14122 , n14123 , n14124 , n14125 , n14126 , n14127 , n14128 , n14129 , n14130 , n14131 , n14132 , n14133 , n14134 , n14135 , n14136 , n14137 , n14138 , n14139 , n14140 , n14141 , n14142 , n14143 , n14144 , n14145 , n14146 , n14147 , n14148 , n14149 , n14150 , n14151 , n14152 , n14153 , n14154 , n14155 , n14156 , n14157 , n14158 , n14159 , n14160 , n14161 , n14162 , n14163 , n14164 , n14165 , n14166 , n14167 , n14168 , n14169 , n14170 , n14171 , n14172 , n14173 , n14174 , n14175 , n14176 , n14177 , n14178 , n14179 , n14180 , n14181 , n14182 , n14183 , n14184 , n14185 , n14186 , n14187 , n14188 , n14189 , n14190 , n14191 , n14192 , n14193 , n14194 , n14195 , n14196 , n14197 , n14198 , n14199 , n14200 , n14201 , n14202 , n14203 , n14204 , n14205 , n14206 , n14207 , n14208 , n14209 , n14210 , n14211 , n14212 , n14213 , n14214 , n14215 , n14216 , n14217 , n14218 , n14219 , n14220 , n14221 , n14222 , n14223 , n14224 , n14225 , n14226 , n14227 , n14228 , n14229 , n14230 , n14231 , n14232 , n14233 , n14234 , n14235 , n14236 , n14237 , n14238 , n14239 , n14240 , n14241 , n14242 , n14243 , n14244 , n14245 , n14246 , n14247 , n14248 , n14249 , n14250 , n14251 , n14252 , n14253 , n14254 , n14255 , n14256 , n14257 , n14258 , n14259 , n14260 , n14261 , n14262 , n14263 , n14264 , n14265 , n14266 , n14267 , n14268 , n14269 , n14270 , n14271 , n14272 , n14273 , n14274 , n14275 , n14276 , n14277 , n14278 , n14279 , n14280 , n14281 , n14282 , n14283 , n14284 , n14285 , n14286 , n14287 , n14288 , n14289 , n14290 , n14291 , n14292 , n14293 , n14294 , n14295 , n14296 , n14297 , n14298 , n14299 , n14300 , n14301 , n14302 , n14303 , n14304 , n14305 , n14306 , n14307 , n14308 , n14309 , n14310 , n14311 , n14312 , n14313 , n14314 , n14315 , n14316 , n14317 , n14318 , n14319 , n14320 , n14321 , n14322 , n14323 , n14324 , n14325 , n14326 , n14327 , n14328 , n14329 , n14330 , n14331 , n14332 , n14333 , n14334 , n14335 , n14336 , n14337 , n14338 , n14339 , n14340 , n14341 , n14342 , n14343 , n14344 , n14345 , n14346 , n14347 , n14348 , n14349 , n14350 , n14351 , n14352 , n14353 , n14354 , n14355 , n14356 , n14357 , n14358 , n14359 , n14360 , n14361 , n14362 , n14363 , n14364 , n14365 , n14366 , n14367 , n14368 , n14369 , n14370 , n14371 , n14372 , n14373 , n14374 , n14375 , n14376 , n14377 , n14378 , n14379 , n14380 , n14381 , n14382 , n14383 , n14384 , n14385 , n14386 , n14387 , n14388 , n14389 , n14390 , n14391 , n14392 , n14393 , n14394 , n14395 , n14396 , n14397 , n14398 , n14399 , n14400 , n14401 , n14402 , n14403 , n14404 , n14405 , n14406 , n14407 , n14408 , n14409 , n14410 , n14411 , n14412 , n14413 , n14414 , n14415 , n14416 , n14417 , n14418 , n14419 , n14420 , n14421 , n14422 , n14423 , n14424 , n14425 , n14426 , n14427 , n14428 , n14429 , n14430 , n14431 , n14432 , n14433 , n14434 , n14435 , n14436 , n14437 , n14438 , n14439 , n14440 , n14441 , n14442 , n14443 , n14444 , n14445 , n14446 , n14447 , n14448 , n14449 , n14450 , n14451 , n14452 , n14453 , n14454 , n14455 , n14456 , n14457 , n14458 , n14459 , n14460 , n14461 , n14462 , n14463 , n14464 , n14465 , n14466 , n14467 , n14468 , n14469 , n14470 , n14471 , n14472 , n14473 , n14474 , n14475 , n14476 , n14477 , n14478 , n14479 , n14480 , n14481 , n14482 , n14483 , n14484 , n14485 , n14486 , n14487 , n14488 , n14489 , n14490 , n14491 , n14492 , n14493 , n14494 , n14495 , n14496 , n14497 , n14498 , n14499 , n14500 , n14501 , n14502 , n14503 , n14504 , n14505 , n14506 , n14507 , n14508 , n14509 , n14510 , n14511 , n14512 , n14513 , n14514 , n14515 , n14516 , n14517 , n14518 , n14519 , n14520 , n14521 , n14522 , n14523 , n14524 , n14525 , n14526 , n14527 , n14528 , n14529 , n14530 , n14531 , n14532 , n14533 , n14534 , n14535 , n14536 , n14537 , n14538 , n14539 , n14540 , n14541 , n14542 , n14543 , n14544 , n14545 , n14546 , n14547 , n14548 , n14549 , n14550 , n14551 , n14552 , n14553 , n14554 , n14555 , n14556 , n14557 , n14558 , n14559 , n14560 , n14561 , n14562 , n14563 , n14564 , n14565 , n14566 , n14567 , n14568 , n14569 , n14570 , n14571 , n14572 , n14573 , n14574 , n14575 , n14576 , n14577 , n14578 , n14579 , n14580 , n14581 , n14582 , n14583 , n14584 , n14585 , n14586 , n14587 , n14588 , n14589 , n14590 , n14591 , n14592 , n14593 , n14594 , n14595 , n14596 , n14597 , n14598 , n14599 , n14600 , n14601 , n14602 , n14603 , n14604 , n14605 , n14606 , n14607 , n14608 , n14609 , n14610 , n14611 , n14612 , n14613 , n14614 , n14615 , n14616 , n14617 , n14618 , n14619 , n14620 , n14621 , n14622 , n14623 , n14624 , n14625 , n14626 , n14627 , n14628 , n14629 , n14630 , n14631 , n14632 , n14633 , n14634 , n14635 , n14636 , n14637 , n14638 , n14639 , n14640 , n14641 , n14642 , n14643 , n14644 , n14645 , n14646 , n14647 , n14648 , n14649 , n14650 , n14651 , n14652 , n14653 , n14654 , n14655 , n14656 , n14657 , n14658 , n14659 , n14660 , n14661 , n14662 , n14663 , n14664 , n14665 , n14666 , n14667 , n14668 , n14669 , n14670 , n14671 , n14672 , n14673 , n14674 , n14675 , n14676 , n14677 , n14678 , n14679 , n14680 , n14681 , n14682 , n14683 , n14684 , n14685 , n14686 , n14687 , n14688 , n14689 , n14690 , n14691 , n14692 , n14693 , n14694 , n14695 , n14696 , n14697 , n14698 , n14699 , n14700 , n14701 , n14702 , n14703 , n14704 , n14705 , n14706 , n14707 , n14708 , n14709 , n14710 , n14711 , n14712 , n14713 , n14714 , n14715 , n14716 , n14717 , n14718 , n14719 , n14720 , n14721 , n14722 , n14723 , n14724 , n14725 , n14726 , n14727 , n14728 , n14729 , n14730 , n14731 , n14732 , n14733 , n14734 , n14735 , n14736 , n14737 , n14738 , n14739 , n14740 , n14741 , n14742 , n14743 , n14744 , n14745 , n14746 , n14747 , n14748 , n14749 , n14750 , n14751 , n14752 , n14753 , n14754 , n14755 , n14756 , n14757 , n14758 , n14759 , n14760 , n14761 , n14762 , n14763 , n14764 , n14765 , n14766 , n14767 , n14768 , n14769 , n14770 , n14771 , n14772 , n14773 , n14774 , n14775 , n14776 , n14777 , n14778 , n14779 , n14780 , n14781 , n14782 , n14783 , n14784 , n14785 , n14786 , n14787 , n14788 , n14789 , n14790 , n14791 , n14792 , n14793 , n14794 , n14795 , n14796 , n14797 , n14798 , n14799 , n14800 , n14801 , n14802 , n14803 , n14804 , n14805 , n14806 , n14807 , n14808 , n14809 , n14810 , n14811 , n14812 , n14813 , n14814 , n14815 , n14816 , n14817 , n14818 , n14819 , n14820 , n14821 , n14822 , n14823 , n14824 , n14825 , n14826 , n14827 , n14828 , n14829 , n14830 , n14831 , n14832 , n14833 , n14834 , n14835 , n14836 , n14837 , n14838 , n14839 , n14840 , n14841 , n14842 , n14843 , n14844 , n14845 , n14846 , n14847 , n14848 , n14849 , n14850 , n14851 , n14852 , n14853 , n14854 , n14855 , n14856 , n14857 , n14858 , n14859 , n14860 , n14861 , n14862 , n14863 , n14864 , n14865 , n14866 , n14867 , n14868 , n14869 , n14870 , n14871 , n14872 , n14873 , n14874 , n14875 , n14876 , n14877 , n14878 , n14879 , n14880 , n14881 , n14882 , n14883 , n14884 , n14885 , n14886 , n14887 , n14888 , n14889 , n14890 , n14891 , n14892 , n14893 , n14894 , n14895 , n14896 , n14897 , n14898 , n14899 , n14900 , n14901 , n14902 , n14903 , n14904 , n14905 , n14906 , n14907 , n14908 , n14909 , n14910 , n14911 , n14912 , n14913 , n14914 , n14915 , n14916 , n14917 , n14918 , n14919 , n14920 , n14921 , n14922 , n14923 , n14924 , n14925 , n14926 , n14927 , n14928 , n14929 , n14930 , n14931 , n14932 , n14933 , n14934 , n14935 , n14936 , n14937 , n14938 , n14939 , n14940 , n14941 , n14942 , n14943 , n14944 , n14945 , n14946 , n14947 , n14948 , n14949 , n14950 , n14951 , n14952 , n14953 , n14954 , n14955 , n14956 , n14957 , n14958 , n14959 , n14960 , n14961 , n14962 , n14963 , n14964 , n14965 , n14966 , n14967 , n14968 , n14969 , n14970 , n14971 , n14972 , n14973 , n14974 , n14975 , n14976 , n14977 , n14978 , n14979 , n14980 , n14981 , n14982 , n14983 , n14984 , n14985 , n14986 , n14987 , n14988 , n14989 , n14990 , n14991 , n14992 , n14993 , n14994 , n14995 , n14996 , n14997 , n14998 , n14999 , n15000 , n15001 , n15002 , n15003 , n15004 , n15005 , n15006 , n15007 , n15008 , n15009 , n15010 , n15011 , n15012 , n15013 , n15014 , n15015 , n15016 , n15017 , n15018 , n15019 , n15020 , n15021 , n15022 , n15023 , n15024 , n15025 , n15026 , n15027 , n15028 , n15029 , n15030 , n15031 , n15032 , n15033 , n15034 , n15035 , n15036 , n15037 , n15038 , n15039 , n15040 , n15041 , n15042 , n15043 , n15044 , n15045 , n15046 , n15047 , n15048 , n15049 , n15050 , n15051 , n15052 , n15053 , n15054 , n15055 , n15056 , n15057 , n15058 , n15059 , n15060 , n15061 , n15062 , n15063 , n15064 , n15065 , n15066 , n15067 , n15068 , n15069 , n15070 , n15071 , n15072 , n15073 , n15074 , n15075 , n15076 , n15077 , n15078 , n15079 , n15080 , n15081 , n15082 , n15083 , n15084 , n15085 , n15086 , n15087 , n15088 , n15089 , n15090 , n15091 , n15092 , n15093 , n15094 , n15095 , n15096 , n15097 , n15098 , n15099 , n15100 , n15101 , n15102 , n15103 , n15104 , n15105 , n15106 , n15107 , n15108 , n15109 , n15110 , n15111 , n15112 , n15113 , n15114 , n15115 , n15116 , n15117 , n15118 , n15119 , n15120 , n15121 , n15122 , n15123 , n15124 , n15125 , n15126 , n15127 , n15128 , n15129 , n15130 , n15131 , n15132 , n15133 , n15134 , n15135 , n15136 , n15137 , n15138 , n15139 , n15140 , n15141 , n15142 , n15143 , n15144 , n15145 , n15146 , n15147 , n15148 , n15149 , n15150 , n15151 , n15152 , n15153 , n15154 , n15155 , n15156 , n15157 , n15158 , n15159 , n15160 , n15161 , n15162 , n15163 , n15164 , n15165 , n15166 , n15167 , n15168 , n15169 , n15170 , n15171 , n15172 , n15173 , n15174 , n15175 , n15176 , n15177 , n15178 , n15179 , n15180 , n15181 , n15182 , n15183 , n15184 , n15185 , n15186 , n15187 , n15188 , n15189 , n15190 , n15191 , n15192 , n15193 , n15194 , n15195 , n15196 , n15197 , n15198 , n15199 , n15200 , n15201 , n15202 , n15203 , n15204 , n15205 , n15206 , n15207 , n15208 , n15209 , n15210 , n15211 , n15212 , n15213 , n15214 , n15215 , n15216 , n15217 , n15218 , n15219 , n15220 , n15221 , n15222 , n15223 , n15224 , n15225 , n15226 , n15227 , n15228 , n15229 , n15230 , n15231 , n15232 , n15233 , n15234 , n15235 , n15236 , n15237 , n15238 , n15239 , n15240 , n15241 , n15242 , n15243 , n15244 , n15245 , n15246 , n15247 , n15248 , n15249 , n15250 , n15251 , n15252 , n15253 , n15254 , n15255 , n15256 , n15257 , n15258 , n15259 , n15260 , n15261 , n15262 , n15263 , n15264 , n15265 , n15266 , n15267 , n15268 , n15269 , n15270 , n15271 , n15272 , n15273 , n15274 , n15275 , n15276 , n15277 , n15278 , n15279 , n15280 , n15281 , n15282 , n15283 , n15284 , n15285 , n15286 , n15287 , n15288 , n15289 , n15290 , n15291 , n15292 , n15293 , n15294 , n15295 , n15296 , n15297 , n15298 , n15299 , n15300 , n15301 , n15302 , n15303 , n15304 , n15305 , n15306 , n15307 , n15308 , n15309 , n15310 , n15311 , n15312 , n15313 , n15314 , n15315 , n15316 , n15317 , n15318 , n15319 , n15320 , n15321 , n15322 , n15323 , n15324 , n15325 , n15326 , n15327 , n15328 , n15329 , n15330 , n15331 , n15332 , n15333 , n15334 , n15335 , n15336 , n15337 , n15338 , n15339 , n15340 , n15341 , n15342 , n15343 , n15344 , n15345 , n15346 , n15347 , n15348 , n15349 , n15350 , n15351 , n15352 , n15353 , n15354 , n15355 , n15356 , n15357 , n15358 , n15359 , n15360 , n15361 , n15362 , n15363 , n15364 , n15365 , n15366 , n15367 , n15368 , n15369 , n15370 , n15371 , n15372 , n15373 , n15374 , n15375 , n15376 , n15377 , n15378 , n15379 , n15380 , n15381 , n15382 , n15383 , n15384 , n15385 , n15386 , n15387 , n15388 , n15389 , n15390 , n15391 , n15392 , n15393 , n15394 , n15395 , n15396 , n15397 , n15398 , n15399 , n15400 , n15401 , n15402 , n15403 , n15404 , n15405 , n15406 , n15407 , n15408 , n15409 , n15410 , n15411 , n15412 , n15413 , n15414 , n15415 , n15416 , n15417 , n15418 , n15419 , n15420 , n15421 , n15422 , n15423 , n15424 , n15425 , n15426 , n15427 , n15428 , n15429 , n15430 , n15431 , n15432 , n15433 , n15434 , n15435 , n15436 , n15437 , n15438 , n15439 , n15440 , n15441 , n15442 , n15443 , n15444 , n15445 , n15446 , n15447 , n15448 , n15449 , n15450 , n15451 , n15452 , n15453 , n15454 , n15455 , n15456 , n15457 , n15458 , n15459 , n15460 , n15461 , n15462 , n15463 , n15464 , n15465 , n15466 , n15467 , n15468 , n15469 , n15470 , n15471 , n15472 , n15473 , n15474 , n15475 , n15476 , n15477 , n15478 , n15479 , n15480 , n15481 , n15482 , n15483 , n15484 , n15485 , n15486 , n15487 , n15488 , n15489 , n15490 , n15491 , n15492 , n15493 , n15494 , n15495 , n15496 , n15497 , n15498 , n15499 , n15500 , n15501 , n15502 , n15503 , n15504 , n15505 , n15506 , n15507 , n15508 , n15509 , n15510 , n15511 , n15512 , n15513 , n15514 , n15515 , n15516 , n15517 , n15518 , n15519 , n15520 , n15521 , n15522 , n15523 , n15524 , n15525 , n15526 , n15527 , n15528 , n15529 , n15530 , n15531 , n15532 , n15533 , n15534 , n15535 , n15536 , n15537 , n15538 , n15539 , n15540 , n15541 , n15542 , n15543 , n15544 , n15545 , n15546 , n15547 , n15548 , n15549 , n15550 , n15551 , n15552 , n15553 , n15554 , n15555 , n15556 , n15557 , n15558 , n15559 , n15560 , n15561 , n15562 , n15563 , n15564 , n15565 , n15566 , n15567 , n15568 , n15569 , n15570 , n15571 , n15572 , n15573 , n15574 , n15575 , n15576 , n15577 , n15578 , n15579 , n15580 , n15581 , n15582 , n15583 , n15584 , n15585 , n15586 , n15587 , n15588 , n15589 , n15590 , n15591 , n15592 , n15593 , n15594 , n15595 , n15596 , n15597 , n15598 , n15599 , n15600 , n15601 , n15602 , n15603 , n15604 , n15605 , n15606 , n15607 , n15608 , n15609 , n15610 , n15611 , n15612 , n15613 , n15614 , n15615 , n15616 , n15617 , n15618 , n15619 , n15620 , n15621 , n15622 , n15623 , n15624 , n15625 , n15626 , n15627 , n15628 , n15629 , n15630 , n15631 , n15632 , n15633 , n15634 , n15635 , n15636 , n15637 , n15638 , n15639 , n15640 , n15641 , n15642 , n15643 , n15644 , n15645 , n15646 , n15647 , n15648 , n15649 , n15650 , n15651 , n15652 , n15653 , n15654 , n15655 , n15656 , n15657 , n15658 , n15659 , n15660 , n15661 , n15662 , n15663 , n15664 , n15665 , n15666 , n15667 , n15668 , n15669 , n15670 , n15671 , n15672 , n15673 , n15674 , n15675 , n15676 , n15677 , n15678 , n15679 , n15680 , n15681 , n15682 , n15683 , n15684 , n15685 , n15686 , n15687 , n15688 , n15689 , n15690 , n15691 , n15692 , n15693 , n15694 , n15695 , n15696 , n15697 , n15698 , n15699 , n15700 , n15701 , n15702 , n15703 , n15704 , n15705 , n15706 , n15707 , n15708 , n15709 , n15710 , n15711 , n15712 , n15713 , n15714 , n15715 , n15716 , n15717 , n15718 , n15719 , n15720 , n15721 , n15722 , n15723 , n15724 , n15725 , n15726 , n15727 , n15728 , n15729 , n15730 , n15731 , n15732 , n15733 , n15734 , n15735 , n15736 , n15737 , n15738 , n15739 , n15740 , n15741 , n15742 , n15743 , n15744 , n15745 , n15746 , n15747 , n15748 , n15749 , n15750 , n15751 , n15752 , n15753 , n15754 , n15755 , n15756 , n15757 , n15758 , n15759 , n15760 , n15761 , n15762 , n15763 , n15764 , n15765 , n15766 , n15767 , n15768 , n15769 , n15770 , n15771 , n15772 , n15773 , n15774 , n15775 , n15776 , n15777 , n15778 , n15779 , n15780 , n15781 , n15782 , n15783 , n15784 , n15785 , n15786 , n15787 , n15788 , n15789 , n15790 , n15791 , n15792 , n15793 , n15794 , n15795 , n15796 , n15797 , n15798 , n15799 , n15800 , n15801 , n15802 , n15803 , n15804 , n15805 , n15806 , n15807 , n15808 , n15809 , n15810 , n15811 , n15812 , n15813 , n15814 , n15815 , n15816 , n15817 , n15818 , n15819 , n15820 , n15821 , n15822 , n15823 , n15824 , n15825 , n15826 , n15827 , n15828 , n15829 , n15830 , n15831 , n15832 , n15833 , n15834 , n15835 , n15836 , n15837 , n15838 , n15839 , n15840 , n15841 , n15842 , n15843 , n15844 , n15845 , n15846 , n15847 , n15848 , n15849 , n15850 , n15851 , n15852 , n15853 , n15854 , n15855 , n15856 , n15857 , n15858 , n15859 , n15860 , n15861 , n15862 , n15863 , n15864 , n15865 , n15866 , n15867 , n15868 , n15869 , n15870 , n15871 , n15872 , n15873 , n15874 , n15875 , n15876 , n15877 , n15878 , n15879 , n15880 , n15881 , n15882 , n15883 , n15884 , n15885 , n15886 , n15887 , n15888 , n15889 , n15890 , n15891 , n15892 , n15893 , n15894 , n15895 , n15896 , n15897 , n15898 , n15899 , n15900 , n15901 , n15902 , n15903 , n15904 , n15905 , n15906 , n15907 , n15908 , n15909 , n15910 , n15911 , n15912 , n15913 , n15914 , n15915 , n15916 , n15917 , n15918 , n15919 , n15920 , n15921 , n15922 , n15923 , n15924 , n15925 , n15926 , n15927 , n15928 , n15929 , n15930 , n15931 , n15932 , n15933 , n15934 , n15935 , n15936 , n15937 , n15938 , n15939 , n15940 , n15941 , n15942 , n15943 , n15944 , n15945 , n15946 , n15947 , n15948 , n15949 , n15950 , n15951 , n15952 , n15953 , n15954 , n15955 , n15956 , n15957 , n15958 , n15959 , n15960 , n15961 , n15962 , n15963 , n15964 , n15965 , n15966 , n15967 , n15968 , n15969 , n15970 , n15971 , n15972 , n15973 , n15974 , n15975 , n15976 , n15977 , n15978 , n15979 , n15980 , n15981 , n15982 , n15983 , n15984 , n15985 , n15986 , n15987 , n15988 , n15989 , n15990 , n15991 , n15992 , n15993 , n15994 , n15995 , n15996 , n15997 , n15998 , n15999 , n16000 , n16001 , n16002 , n16003 , n16004 , n16005 , n16006 , n16007 , n16008 , n16009 , n16010 , n16011 , n16012 , n16013 , n16014 , n16015 , n16016 , n16017 , n16018 , n16019 , n16020 , n16021 , n16022 , n16023 , n16024 , n16025 , n16026 , n16027 , n16028 , n16029 , n16030 , n16031 , n16032 , n16033 , n16034 , n16035 , n16036 , n16037 , n16038 , n16039 , n16040 , n16041 , n16042 , n16043 , n16044 , n16045 , n16046 , n16047 , n16048 , n16049 , n16050 , n16051 , n16052 , n16053 , n16054 , n16055 , n16056 , n16057 , n16058 , n16059 , n16060 , n16061 , n16062 , n16063 , n16064 , n16065 , n16066 , n16067 , n16068 , n16069 , n16070 , n16071 , n16072 , n16073 , n16074 , n16075 , n16076 , n16077 , n16078 , n16079 , n16080 , n16081 , n16082 , n16083 , n16084 , n16085 , n16086 , n16087 , n16088 , n16089 , n16090 , n16091 , n16092 , n16093 , n16094 , n16095 , n16096 , n16097 , n16098 , n16099 , n16100 , n16101 , n16102 , n16103 , n16104 , n16105 , n16106 , n16107 , n16108 , n16109 , n16110 , n16111 , n16112 , n16113 , n16114 , n16115 , n16116 , n16117 , n16118 , n16119 , n16120 , n16121 , n16122 , n16123 , n16124 , n16125 , n16126 , n16127 , n16128 , n16129 , n16130 , n16131 , n16132 , n16133 , n16134 , n16135 , n16136 , n16137 , n16138 , n16139 , n16140 , n16141 , n16142 , n16143 , n16144 , n16145 , n16146 , n16147 , n16148 , n16149 , n16150 , n16151 , n16152 , n16153 , n16154 , n16155 , n16156 , n16157 , n16158 , n16159 , n16160 , n16161 , n16162 , n16163 , n16164 , n16165 , n16166 , n16167 , n16168 , n16169 , n16170 , n16171 , n16172 , n16173 , n16174 , n16175 , n16176 , n16177 , n16178 , n16179 , n16180 , n16181 , n16182 , n16183 , n16184 , n16185 , n16186 , n16187 , n16188 , n16189 , n16190 , n16191 , n16192 , n16193 , n16194 , n16195 , n16196 , n16197 , n16198 , n16199 , n16200 , n16201 , n16202 , n16203 , n16204 , n16205 , n16206 , n16207 , n16208 , n16209 , n16210 , n16211 , n16212 , n16213 , n16214 , n16215 , n16216 , n16217 , n16218 , n16219 , n16220 , n16221 , n16222 , n16223 , n16224 , n16225 , n16226 , n16227 , n16228 , n16229 , n16230 , n16231 , n16232 , n16233 , n16234 , n16235 , n16236 , n16237 , n16238 , n16239 , n16240 , n16241 , n16242 , n16243 , n16244 , n16245 , n16246 , n16247 , n16248 , n16249 , n16250 , n16251 , n16252 , n16253 , n16254 , n16255 , n16256 , n16257 , n16258 , n16259 , n16260 , n16261 , n16262 , n16263 , n16264 , n16265 , n16266 , n16267 , n16268 , n16269 , n16270 , n16271 , n16272 , n16273 , n16274 , n16275 , n16276 , n16277 , n16278 , n16279 , n16280 , n16281 , n16282 , n16283 , n16284 , n16285 , n16286 , n16287 , n16288 , n16289 , n16290 , n16291 , n16292 , n16293 , n16294 , n16295 , n16296 , n16297 , n16298 , n16299 , n16300 , n16301 , n16302 , n16303 , n16304 , n16305 , n16306 , n16307 , n16308 , n16309 , n16310 , n16311 , n16312 , n16313 , n16314 , n16315 , n16316 , n16317 , n16318 , n16319 , n16320 , n16321 , n16322 , n16323 , n16324 , n16325 , n16326 , n16327 , n16328 , n16329 , n16330 , n16331 , n16332 , n16333 , n16334 , n16335 , n16336 , n16337 , n16338 , n16339 , n16340 , n16341 , n16342 , n16343 , n16344 , n16345 , n16346 , n16347 , n16348 , n16349 , n16350 , n16351 , n16352 , n16353 , n16354 , n16355 , n16356 , n16357 , n16358 , n16359 , n16360 , n16361 , n16362 , n16363 , n16364 , n16365 , n16366 , n16367 , n16368 , n16369 , n16370 , n16371 , n16372 , n16373 , n16374 , n16375 , n16376 , n16377 , n16378 , n16379 , n16380 , n16381 , n16382 , n16383 , n16384 , n16385 , n16386 , n16387 , n16388 , n16389 , n16390 , n16391 , n16392 , n16393 , n16394 , n16395 , n16396 , n16397 , n16398 , n16399 , n16400 , n16401 , n16402 , n16403 , n16404 , n16405 , n16406 , n16407 , n16408 , n16409 , n16410 , n16411 , n16412 , n16413 , n16414 , n16415 , n16416 , n16417 , n16418 , n16419 , n16420 , n16421 , n16422 , n16423 , n16424 , n16425 , n16426 , n16427 , n16428 , n16429 , n16430 , n16431 , n16432 , n16433 , n16434 , n16435 , n16436 , n16437 , n16438 , n16439 , n16440 , n16441 , n16442 , n16443 , n16444 , n16445 , n16446 , n16447 , n16448 , n16449 , n16450 , n16451 , n16452 , n16453 , n16454 , n16455 , n16456 , n16457 , n16458 , n16459 , n16460 , n16461 , n16462 , n16463 , n16464 , n16465 , n16466 , n16467 , n16468 , n16469 , n16470 , n16471 , n16472 , n16473 , n16474 , n16475 , n16476 , n16477 , n16478 , n16479 , n16480 , n16481 , n16482 , n16483 , n16484 , n16485 , n16486 , n16487 , n16488 , n16489 , n16490 , n16491 , n16492 , n16493 , n16494 , n16495 , n16496 , n16497 , n16498 , n16499 , n16500 , n16501 , n16502 , n16503 , n16504 , n16505 , n16506 , n16507 , n16508 , n16509 , n16510 , n16511 , n16512 , n16513 , n16514 , n16515 , n16516 , n16517 , n16518 , n16519 , n16520 , n16521 , n16522 , n16523 , n16524 , n16525 , n16526 , n16527 , n16528 , n16529 , n16530 , n16531 , n16532 , n16533 , n16534 , n16535 , n16536 , n16537 , n16538 , n16539 , n16540 , n16541 , n16542 , n16543 , n16544 , n16545 , n16546 , n16547 , n16548 , n16549 , n16550 , n16551 , n16552 , n16553 , n16554 , n16555 , n16556 , n16557 , n16558 , n16559 , n16560 , n16561 , n16562 , n16563 , n16564 , n16565 , n16566 , n16567 , n16568 , n16569 , n16570 , n16571 , n16572 , n16573 , n16574 , n16575 , n16576 , n16577 , n16578 , n16579 , n16580 , n16581 , n16582 , n16583 , n16584 , n16585 , n16586 , n16587 , n16588 , n16589 , n16590 , n16591 , n16592 , n16593 , n16594 , n16595 , n16596 , n16597 , n16598 , n16599 , n16600 , n16601 , n16602 , n16603 , n16604 , n16605 , n16606 , n16607 , n16608 , n16609 , n16610 , n16611 , n16612 , n16613 , n16614 , n16615 , n16616 , n16617 , n16618 , n16619 , n16620 , n16621 , n16622 , n16623 , n16624 , n16625 , n16626 , n16627 , n16628 , n16629 , n16630 , n16631 , n16632 , n16633 , n16634 , n16635 , n16636 , n16637 , n16638 , n16639 , n16640 , n16641 , n16642 , n16643 , n16644 , n16645 , n16646 , n16647 , n16648 , n16649 , n16650 , n16651 , n16652 , n16653 , n16654 , n16655 , n16656 , n16657 , n16658 , n16659 , n16660 , n16661 , n16662 , n16663 , n16664 , n16665 , n16666 , n16667 , n16668 , n16669 , n16670 , n16671 , n16672 , n16673 , n16674 , n16675 , n16676 , n16677 , n16678 , n16679 , n16680 , n16681 , n16682 , n16683 , n16684 , n16685 , n16686 , n16687 , n16688 , n16689 , n16690 , n16691 , n16692 , n16693 , n16694 , n16695 , n16696 , n16697 , n16698 , n16699 , n16700 , n16701 , n16702 , n16703 , n16704 , n16705 , n16706 , n16707 , n16708 , n16709 , n16710 , n16711 , n16712 , n16713 , n16714 , n16715 , n16716 , n16717 , n16718 , n16719 , n16720 , n16721 , n16722 , n16723 , n16724 , n16725 , n16726 , n16727 , n16728 , n16729 , n16730 , n16731 , n16732 , n16733 , n16734 , n16735 , n16736 , n16737 , n16738 , n16739 , n16740 , n16741 , n16742 , n16743 , n16744 , n16745 , n16746 , n16747 , n16748 , n16749 , n16750 , n16751 , n16752 , n16753 , n16754 , n16755 , n16756 , n16757 , n16758 , n16759 , n16760 , n16761 , n16762 , n16763 , n16764 , n16765 , n16766 , n16767 , n16768 , n16769 , n16770 , n16771 , n16772 , n16773 , n16774 , n16775 , n16776 , n16777 , n16778 , n16779 , n16780 , n16781 , n16782 , n16783 , n16784 , n16785 , n16786 , n16787 , n16788 , n16789 , n16790 , n16791 , n16792 , n16793 , n16794 , n16795 , n16796 , n16797 , n16798 , n16799 , n16800 , n16801 , n16802 , n16803 , n16804 , n16805 , n16806 , n16807 , n16808 , n16809 , n16810 , n16811 , n16812 , n16813 , n16814 , n16815 , n16816 , n16817 , n16818 , n16819 , n16820 , n16821 , n16822 , n16823 , n16824 , n16825 , n16826 , n16827 , n16828 , n16829 , n16830 , n16831 , n16832 , n16833 , n16834 , n16835 , n16836 , n16837 , n16838 , n16839 , n16840 , n16841 , n16842 , n16843 , n16844 , n16845 , n16846 , n16847 , n16848 , n16849 , n16850 , n16851 , n16852 , n16853 , n16854 , n16855 , n16856 , n16857 , n16858 , n16859 , n16860 , n16861 , n16862 , n16863 , n16864 , n16865 , n16866 , n16867 , n16868 , n16869 , n16870 , n16871 , n16872 , n16873 , n16874 , n16875 , n16876 , n16877 , n16878 , n16879 , n16880 , n16881 , n16882 , n16883 , n16884 , n16885 , n16886 , n16887 , n16888 , n16889 , n16890 , n16891 , n16892 , n16893 , n16894 , n16895 , n16896 , n16897 , n16898 , n16899 , n16900 , n16901 , n16902 , n16903 , n16904 , n16905 , n16906 , n16907 , n16908 , n16909 , n16910 , n16911 , n16912 , n16913 , n16914 , n16915 , n16916 , n16917 , n16918 , n16919 , n16920 , n16921 , n16922 , n16923 , n16924 , n16925 , n16926 , n16927 , n16928 , n16929 , n16930 , n16931 , n16932 , n16933 , n16934 , n16935 , n16936 , n16937 , n16938 , n16939 , n16940 , n16941 , n16942 , n16943 , n16944 , n16945 , n16946 , n16947 , n16948 , n16949 , n16950 , n16951 , n16952 , n16953 , n16954 , n16955 , n16956 , n16957 , n16958 , n16959 , n16960 , n16961 , n16962 , n16963 , n16964 , n16965 , n16966 , n16967 , n16968 , n16969 , n16970 , n16971 , n16972 , n16973 , n16974 , n16975 , n16976 , n16977 , n16978 , n16979 , n16980 , n16981 , n16982 , n16983 , n16984 , n16985 , n16986 , n16987 , n16988 , n16989 , n16990 , n16991 , n16992 , n16993 , n16994 , n16995 , n16996 , n16997 , n16998 , n16999 , n17000 , n17001 , n17002 , n17003 , n17004 , n17005 , n17006 , n17007 , n17008 , n17009 , n17010 , n17011 , n17012 , n17013 , n17014 , n17015 , n17016 , n17017 , n17018 , n17019 , n17020 , n17021 , n17022 , n17023 , n17024 , n17025 , n17026 , n17027 , n17028 , n17029 , n17030 , n17031 , n17032 , n17033 , n17034 , n17035 , n17036 , n17037 , n17038 , n17039 , n17040 , n17041 , n17042 , n17043 , n17044 , n17045 , n17046 , n17047 , n17048 , n17049 , n17050 , n17051 , n17052 , n17053 , n17054 , n17055 , n17056 , n17057 , n17058 , n17059 , n17060 , n17061 , n17062 , n17063 , n17064 , n17065 , n17066 , n17067 , n17068 , n17069 , n17070 , n17071 , n17072 , n17073 , n17074 , n17075 , n17076 , n17077 , n17078 , n17079 , n17080 , n17081 , n17082 , n17083 , n17084 , n17085 , n17086 , n17087 , n17088 , n17089 , n17090 , n17091 , n17092 , n17093 , n17094 , n17095 , n17096 , n17097 , n17098 , n17099 , n17100 , n17101 , n17102 , n17103 , n17104 , n17105 , n17106 , n17107 , n17108 , n17109 , n17110 , n17111 , n17112 , n17113 , n17114 , n17115 , n17116 , n17117 , n17118 , n17119 , n17120 , n17121 , n17122 , n17123 , n17124 , n17125 , n17126 , n17127 , n17128 , n17129 , n17130 , n17131 , n17132 , n17133 , n17134 , n17135 , n17136 , n17137 , n17138 , n17139 , n17140 , n17141 , n17142 , n17143 , n17144 , n17145 , n17146 , n17147 , n17148 , n17149 , n17150 , n17151 , n17152 , n17153 , n17154 , n17155 , n17156 , n17157 , n17158 , n17159 , n17160 , n17161 , n17162 , n17163 , n17164 , n17165 , n17166 , n17167 , n17168 , n17169 , n17170 , n17171 , n17172 , n17173 , n17174 , n17175 , n17176 , n17177 , n17178 , n17179 , n17180 , n17181 , n17182 , n17183 , n17184 , n17185 , n17186 , n17187 , n17188 , n17189 , n17190 , n17191 , n17192 , n17193 , n17194 , n17195 , n17196 , n17197 , n17198 , n17199 , n17200 , n17201 , n17202 , n17203 , n17204 , n17205 , n17206 , n17207 , n17208 , n17209 , n17210 , n17211 , n17212 , n17213 , n17214 , n17215 , n17216 , n17217 , n17218 , n17219 , n17220 , n17221 , n17222 , n17223 , n17224 , n17225 , n17226 , n17227 , n17228 , n17229 , n17230 , n17231 , n17232 , n17233 , n17234 , n17235 , n17236 , n17237 , n17238 , n17239 , n17240 , n17241 , n17242 , n17243 , n17244 , n17245 , n17246 , n17247 , n17248 , n17249 , n17250 , n17251 , n17252 , n17253 , n17254 , n17255 , n17256 , n17257 , n17258 , n17259 , n17260 , n17261 , n17262 , n17263 , n17264 , n17265 , n17266 , n17267 , n17268 , n17269 , n17270 , n17271 , n17272 , n17273 , n17274 , n17275 , n17276 , n17277 , n17278 , n17279 , n17280 , n17281 , n17282 , n17283 , n17284 , n17285 , n17286 , n17287 , n17288 , n17289 , n17290 , n17291 , n17292 , n17293 , n17294 , n17295 , n17296 , n17297 , n17298 , n17299 , n17300 , n17301 , n17302 , n17303 , n17304 , n17305 , n17306 , n17307 , n17308 , n17309 , n17310 , n17311 , n17312 , n17313 , n17314 , n17315 , n17316 , n17317 , n17318 , n17319 , n17320 , n17321 , n17322 , n17323 , n17324 , n17325 , n17326 , n17327 , n17328 , n17329 , n17330 , n17331 , n17332 , n17333 , n17334 , n17335 , n17336 , n17337 , n17338 , n17339 , n17340 , n17341 , n17342 , n17343 , n17344 , n17345 , n17346 , n17347 , n17348 , n17349 , n17350 , n17351 , n17352 , n17353 , n17354 , n17355 , n17356 , n17357 , n17358 , n17359 , n17360 , n17361 , n17362 , n17363 , n17364 , n17365 , n17366 , n17367 , n17368 , n17369 , n17370 , n17371 , n17372 , n17373 , n17374 , n17375 , n17376 , n17377 , n17378 , n17379 , n17380 , n17381 , n17382 , n17383 , n17384 , n17385 , n17386 , n17387 , n17388 , n17389 , n17390 , n17391 , n17392 , n17393 , n17394 , n17395 , n17396 , n17397 , n17398 , n17399 , n17400 , n17401 , n17402 , n17403 , n17404 , n17405 , n17406 , n17407 , n17408 , n17409 , n17410 , n17411 , n17412 , n17413 , n17414 , n17415 , n17416 , n17417 , n17418 , n17419 , n17420 , n17421 , n17422 , n17423 , n17424 , n17425 , n17426 , n17427 , n17428 , n17429 , n17430 , n17431 , n17432 , n17433 , n17434 , n17435 , n17436 , n17437 , n17438 , n17439 , n17440 , n17441 , n17442 , n17443 , n17444 , n17445 , n17446 , n17447 , n17448 , n17449 , n17450 , n17451 , n17452 , n17453 , n17454 , n17455 , n17456 , n17457 , n17458 , n17459 , n17460 , n17461 , n17462 , n17463 , n17464 , n17465 , n17466 , n17467 , n17468 , n17469 , n17470 , n17471 , n17472 , n17473 , n17474 , n17475 , n17476 , n17477 , n17478 , n17479 , n17480 , n17481 , n17482 , n17483 , n17484 , n17485 , n17486 , n17487 , n17488 , n17489 , n17490 , n17491 , n17492 , n17493 , n17494 , n17495 , n17496 , n17497 , n17498 , n17499 , n17500 , n17501 , n17502 , n17503 , n17504 , n17505 , n17506 , n17507 , n17508 , n17509 , n17510 , n17511 , n17512 , n17513 , n17514 , n17515 , n17516 , n17517 , n17518 , n17519 , n17520 , n17521 , n17522 , n17523 , n17524 , n17525 , n17526 , n17527 , n17528 , n17529 , n17530 , n17531 , n17532 , n17533 , n17534 , n17535 , n17536 , n17537 , n17538 , n17539 , n17540 , n17541 , n17542 , n17543 , n17544 , n17545 , n17546 , n17547 , n17548 , n17549 , n17550 , n17551 , n17552 , n17553 , n17554 , n17555 , n17556 , n17557 , n17558 , n17559 , n17560 , n17561 , n17562 , n17563 , n17564 , n17565 , n17566 , n17567 , n17568 , n17569 , n17570 , n17571 , n17572 , n17573 , n17574 , n17575 , n17576 , n17577 , n17578 , n17579 , n17580 , n17581 , n17582 , n17583 , n17584 , n17585 , n17586 , n17587 , n17588 , n17589 , n17590 , n17591 , n17592 , n17593 , n17594 , n17595 , n17596 , n17597 , n17598 , n17599 , n17600 , n17601 , n17602 , n17603 , n17604 , n17605 , n17606 , n17607 , n17608 , n17609 , n17610 , n17611 , n17612 , n17613 , n17614 , n17615 , n17616 , n17617 , n17618 , n17619 , n17620 , n17621 , n17622 , n17623 , n17624 , n17625 , n17626 , n17627 , n17628 , n17629 , n17630 , n17631 , n17632 , n17633 , n17634 , n17635 , n17636 , n17637 , n17638 , n17639 , n17640 , n17641 , n17642 , n17643 , n17644 , n17645 , n17646 , n17647 , n17648 , n17649 , n17650 , n17651 , n17652 , n17653 , n17654 , n17655 , n17656 , n17657 , n17658 , n17659 , n17660 , n17661 , n17662 , n17663 , n17664 , n17665 , n17666 , n17667 , n17668 , n17669 , n17670 , n17671 , n17672 , n17673 , n17674 , n17675 , n17676 , n17677 , n17678 , n17679 , n17680 , n17681 , n17682 , n17683 , n17684 , n17685 , n17686 , n17687 , n17688 , n17689 , n17690 , n17691 , n17692 , n17693 , n17694 , n17695 , n17696 , n17697 , n17698 , n17699 , n17700 , n17701 , n17702 , n17703 , n17704 , n17705 , n17706 , n17707 , n17708 , n17709 , n17710 , n17711 , n17712 , n17713 , n17714 , n17715 , n17716 , n17717 , n17718 , n17719 , n17720 , n17721 , n17722 , n17723 , n17724 , n17725 , n17726 , n17727 , n17728 , n17729 , n17730 , n17731 , n17732 , n17733 , n17734 , n17735 , n17736 , n17737 , n17738 , n17739 , n17740 , n17741 , n17742 , n17743 , n17744 , n17745 , n17746 , n17747 , n17748 , n17749 , n17750 , n17751 , n17752 , n17753 , n17754 , n17755 , n17756 , n17757 , n17758 , n17759 , n17760 , n17761 , n17762 , n17763 , n17764 , n17765 , n17766 , n17767 , n17768 , n17769 , n17770 , n17771 , n17772 , n17773 , n17774 , n17775 , n17776 , n17777 , n17778 , n17779 , n17780 , n17781 , n17782 , n17783 , n17784 , n17785 , n17786 , n17787 , n17788 , n17789 , n17790 , n17791 , n17792 , n17793 , n17794 , n17795 , n17796 , n17797 , n17798 , n17799 , n17800 , n17801 , n17802 , n17803 , n17804 , n17805 , n17806 , n17807 , n17808 , n17809 , n17810 , n17811 , n17812 , n17813 , n17814 , n17815 , n17816 , n17817 , n17818 , n17819 , n17820 , n17821 , n17822 , n17823 , n17824 , n17825 , n17826 , n17827 , n17828 , n17829 , n17830 , n17831 , n17832 , n17833 , n17834 , n17835 , n17836 , n17837 , n17838 , n17839 , n17840 , n17841 , n17842 , n17843 , n17844 , n17845 , n17846 , n17847 , n17848 , n17849 , n17850 , n17851 , n17852 , n17853 , n17854 , n17855 , n17856 , n17857 , n17858 , n17859 , n17860 , n17861 , n17862 , n17863 , n17864 , n17865 , n17866 , n17867 , n17868 , n17869 , n17870 , n17871 , n17872 , n17873 , n17874 , n17875 , n17876 , n17877 , n17878 , n17879 , n17880 , n17881 , n17882 , n17883 , n17884 , n17885 , n17886 , n17887 , n17888 , n17889 , n17890 , n17891 , n17892 , n17893 , n17894 , n17895 , n17896 , n17897 , n17898 , n17899 , n17900 , n17901 , n17902 , n17903 , n17904 , n17905 , n17906 , n17907 , n17908 , n17909 , n17910 , n17911 , n17912 , n17913 , n17914 , n17915 , n17916 , n17917 , n17918 , n17919 , n17920 , n17921 , n17922 , n17923 , n17924 , n17925 , n17926 , n17927 , n17928 , n17929 , n17930 , n17931 , n17932 , n17933 , n17934 , n17935 , n17936 , n17937 , n17938 , n17939 , n17940 , n17941 , n17942 , n17943 , n17944 , n17945 , n17946 , n17947 , n17948 , n17949 , n17950 , n17951 , n17952 , n17953 , n17954 , n17955 , n17956 , n17957 , n17958 , n17959 , n17960 , n17961 , n17962 , n17963 , n17964 , n17965 , n17966 , n17967 , n17968 , n17969 , n17970 , n17971 , n17972 , n17973 , n17974 , n17975 , n17976 , n17977 , n17978 , n17979 , n17980 , n17981 , n17982 , n17983 , n17984 , n17985 , n17986 , n17987 , n17988 , n17989 , n17990 , n17991 , n17992 , n17993 , n17994 , n17995 , n17996 , n17997 , n17998 , n17999 , n18000 , n18001 , n18002 , n18003 , n18004 , n18005 , n18006 , n18007 , n18008 , n18009 , n18010 , n18011 , n18012 , n18013 , n18014 , n18015 , n18016 , n18017 , n18018 , n18019 , n18020 , n18021 , n18022 , n18023 , n18024 , n18025 , n18026 , n18027 , n18028 , n18029 , n18030 , n18031 , n18032 , n18033 , n18034 , n18035 , n18036 , n18037 , n18038 , n18039 , n18040 , n18041 , n18042 , n18043 , n18044 , n18045 , n18046 , n18047 , n18048 , n18049 , n18050 , n18051 , n18052 , n18053 , n18054 , n18055 , n18056 , n18057 , n18058 , n18059 , n18060 , n18061 , n18062 , n18063 , n18064 , n18065 , n18066 , n18067 , n18068 , n18069 , n18070 , n18071 , n18072 , n18073 , n18074 , n18075 , n18076 , n18077 , n18078 , n18079 , n18080 , n18081 , n18082 , n18083 , n18084 , n18085 , n18086 , n18087 , n18088 , n18089 , n18090 , n18091 , n18092 , n18093 , n18094 , n18095 , n18096 , n18097 , n18098 , n18099 , n18100 , n18101 , n18102 , n18103 , n18104 , n18105 , n18106 , n18107 , n18108 , n18109 , n18110 , n18111 , n18112 , n18113 , n18114 , n18115 , n18116 , n18117 , n18118 , n18119 , n18120 , n18121 , n18122 , n18123 , n18124 , n18125 , n18126 , n18127 , n18128 , n18129 , n18130 , n18131 , n18132 , n18133 , n18134 , n18135 , n18136 , n18137 , n18138 , n18139 , n18140 , n18141 , n18142 , n18143 , n18144 , n18145 , n18146 , n18147 , n18148 , n18149 , n18150 , n18151 , n18152 , n18153 , n18154 , n18155 , n18156 , n18157 , n18158 , n18159 , n18160 , n18161 , n18162 , n18163 , n18164 , n18165 , n18166 , n18167 , n18168 , n18169 , n18170 , n18171 , n18172 , n18173 , n18174 , n18175 , n18176 , n18177 , n18178 , n18179 , n18180 , n18181 , n18182 , n18183 , n18184 , n18185 , n18186 , n18187 , n18188 , n18189 , n18190 , n18191 , n18192 , n18193 , n18194 , n18195 , n18196 , n18197 , n18198 , n18199 , n18200 , n18201 , n18202 , n18203 , n18204 , n18205 , n18206 , n18207 , n18208 , n18209 , n18210 , n18211 , n18212 , n18213 , n18214 , n18215 , n18216 , n18217 , n18218 , n18219 , n18220 , n18221 , n18222 , n18223 , n18224 , n18225 , n18226 , n18227 , n18228 , n18229 , n18230 , n18231 , n18232 , n18233 , n18234 , n18235 , n18236 , n18237 , n18238 , n18239 , n18240 , n18241 , n18242 , n18243 , n18244 , n18245 , n18246 , n18247 , n18248 , n18249 , n18250 , n18251 , n18252 , n18253 , n18254 , n18255 , n18256 , n18257 , n18258 , n18259 , n18260 , n18261 , n18262 , n18263 , n18264 , n18265 , n18266 , n18267 , n18268 , n18269 , n18270 , n18271 , n18272 , n18273 , n18274 , n18275 , n18276 , n18277 , n18278 , n18279 , n18280 , n18281 , n18282 , n18283 , n18284 , n18285 , n18286 , n18287 , n18288 , n18289 , n18290 , n18291 , n18292 , n18293 , n18294 , n18295 , n18296 , n18297 , n18298 , n18299 , n18300 , n18301 , n18302 , n18303 , n18304 , n18305 , n18306 , n18307 , n18308 , n18309 , n18310 , n18311 , n18312 , n18313 , n18314 , n18315 , n18316 , n18317 , n18318 , n18319 , n18320 , n18321 , n18322 , n18323 , n18324 , n18325 , n18326 , n18327 , n18328 , n18329 , n18330 , n18331 , n18332 , n18333 , n18334 , n18335 , n18336 , n18337 , n18338 , n18339 , n18340 , n18341 , n18342 , n18343 , n18344 , n18345 , n18346 , n18347 , n18348 , n18349 , n18350 , n18351 , n18352 , n18353 , n18354 , n18355 , n18356 , n18357 , n18358 , n18359 , n18360 , n18361 , n18362 , n18363 , n18364 , n18365 , n18366 , n18367 , n18368 , n18369 , n18370 , n18371 , n18372 , n18373 , n18374 , n18375 , n18376 , n18377 , n18378 , n18379 , n18380 , n18381 , n18382 , n18383 , n18384 , n18385 , n18386 , n18387 , n18388 , n18389 , n18390 , n18391 , n18392 , n18393 , n18394 , n18395 , n18396 , n18397 , n18398 , n18399 , n18400 , n18401 , n18402 , n18403 , n18404 , n18405 , n18406 , n18407 , n18408 , n18409 , n18410 , n18411 , n18412 , n18413 , n18414 , n18415 , n18416 , n18417 , n18418 , n18419 , n18420 , n18421 , n18422 , n18423 , n18424 , n18425 , n18426 , n18427 , n18428 , n18429 , n18430 , n18431 , n18432 , n18433 , n18434 , n18435 , n18436 , n18437 , n18438 , n18439 , n18440 , n18441 , n18442 , n18443 , n18444 , n18445 , n18446 , n18447 , n18448 , n18449 , n18450 , n18451 , n18452 , n18453 , n18454 , n18455 , n18456 , n18457 , n18458 , n18459 , n18460 , n18461 , n18462 , n18463 , n18464 , n18465 , n18466 , n18467 , n18468 , n18469 , n18470 , n18471 , n18472 , n18473 , n18474 , n18475 , n18476 , n18477 , n18478 , n18479 , n18480 , n18481 , n18482 , n18483 , n18484 , n18485 , n18486 , n18487 , n18488 , n18489 , n18490 , n18491 , n18492 , n18493 , n18494 , n18495 , n18496 , n18497 , n18498 , n18499 , n18500 , n18501 , n18502 , n18503 , n18504 , n18505 , n18506 , n18507 , n18508 , n18509 , n18510 , n18511 , n18512 , n18513 , n18514 , n18515 , n18516 , n18517 , n18518 , n18519 , n18520 , n18521 , n18522 , n18523 , n18524 , n18525 , n18526 , n18527 , n18528 , n18529 , n18530 , n18531 , n18532 , n18533 , n18534 , n18535 , n18536 , n18537 , n18538 , n18539 , n18540 , n18541 , n18542 , n18543 , n18544 , n18545 , n18546 , n18547 , n18548 , n18549 , n18550 , n18551 , n18552 , n18553 , n18554 , n18555 , n18556 , n18557 , n18558 , n18559 , n18560 , n18561 , n18562 , n18563 , n18564 , n18565 , n18566 , n18567 , n18568 , n18569 , n18570 , n18571 , n18572 , n18573 , n18574 , n18575 , n18576 , n18577 , n18578 , n18579 , n18580 , n18581 , n18582 , n18583 , n18584 , n18585 , n18586 , n18587 , n18588 , n18589 , n18590 , n18591 , n18592 , n18593 , n18594 , n18595 , n18596 , n18597 , n18598 , n18599 , n18600 , n18601 , n18602 , n18603 , n18604 , n18605 , n18606 , n18607 , n18608 , n18609 , n18610 , n18611 , n18612 , n18613 , n18614 , n18615 , n18616 , n18617 , n18618 , n18619 , n18620 , n18621 , n18622 , n18623 , n18624 , n18625 , n18626 , n18627 , n18628 , n18629 , n18630 , n18631 , n18632 , n18633 , n18634 , n18635 , n18636 , n18637 , n18638 , n18639 , n18640 , n18641 , n18642 , n18643 , n18644 , n18645 , n18646 , n18647 , n18648 , n18649 , n18650 , n18651 , n18652 , n18653 , n18654 , n18655 , n18656 , n18657 , n18658 , n18659 , n18660 , n18661 , n18662 , n18663 , n18664 , n18665 , n18666 , n18667 , n18668 , n18669 , n18670 , n18671 , n18672 , n18673 , n18674 , n18675 , n18676 , n18677 , n18678 , n18679 , n18680 , n18681 , n18682 , n18683 , n18684 , n18685 , n18686 , n18687 , n18688 , n18689 , n18690 , n18691 , n18692 , n18693 , n18694 , n18695 , n18696 , n18697 , n18698 , n18699 , n18700 , n18701 , n18702 , n18703 , n18704 , n18705 , n18706 , n18707 , n18708 , n18709 , n18710 , n18711 , n18712 , n18713 , n18714 , n18715 , n18716 , n18717 , n18718 , n18719 , n18720 , n18721 , n18722 , n18723 , n18724 , n18725 , n18726 , n18727 , n18728 , n18729 , n18730 , n18731 , n18732 , n18733 , n18734 , n18735 , n18736 , n18737 , n18738 , n18739 , n18740 , n18741 , n18742 , n18743 , n18744 , n18745 , n18746 , n18747 , n18748 , n18749 , n18750 , n18751 , n18752 , n18753 , n18754 , n18755 , n18756 , n18757 , n18758 , n18759 , n18760 , n18761 , n18762 , n18763 , n18764 , n18765 , n18766 , n18767 , n18768 , n18769 , n18770 , n18771 , n18772 , n18773 , n18774 , n18775 , n18776 , n18777 , n18778 , n18779 , n18780 , n18781 , n18782 , n18783 , n18784 , n18785 , n18786 , n18787 , n18788 , n18789 , n18790 , n18791 , n18792 , n18793 , n18794 , n18795 , n18796 , n18797 , n18798 , n18799 , n18800 , n18801 , n18802 , n18803 , n18804 , n18805 , n18806 , n18807 , n18808 , n18809 , n18810 , n18811 , n18812 , n18813 , n18814 , n18815 , n18816 , n18817 , n18818 , n18819 , n18820 , n18821 , n18822 , n18823 , n18824 , n18825 , n18826 , n18827 , n18828 , n18829 , n18830 , n18831 , n18832 , n18833 , n18834 , n18835 , n18836 , n18837 , n18838 , n18839 , n18840 , n18841 , n18842 , n18843 , n18844 , n18845 , n18846 , n18847 , n18848 , n18849 , n18850 , n18851 , n18852 , n18853 , n18854 , n18855 , n18856 , n18857 , n18858 , n18859 , n18860 , n18861 , n18862 , n18863 , n18864 , n18865 , n18866 , n18867 , n18868 , n18869 , n18870 , n18871 , n18872 , n18873 , n18874 , n18875 , n18876 , n18877 , n18878 , n18879 , n18880 , n18881 , n18882 , n18883 , n18884 , n18885 , n18886 , n18887 , n18888 , n18889 , n18890 , n18891 , n18892 , n18893 , n18894 , n18895 , n18896 , n18897 , n18898 , n18899 , n18900 , n18901 , n18902 , n18903 , n18904 , n18905 , n18906 , n18907 , n18908 , n18909 , n18910 , n18911 , n18912 , n18913 , n18914 , n18915 , n18916 , n18917 , n18918 , n18919 , n18920 , n18921 , n18922 , n18923 , n18924 , n18925 , n18926 , n18927 , n18928 , n18929 , n18930 , n18931 , n18932 , n18933 , n18934 , n18935 , n18936 , n18937 , n18938 , n18939 , n18940 , n18941 , n18942 , n18943 , n18944 , n18945 , n18946 , n18947 , n18948 , n18949 , n18950 , n18951 , n18952 , n18953 , n18954 , n18955 , n18956 , n18957 , n18958 , n18959 , n18960 , n18961 , n18962 , n18963 , n18964 , n18965 , n18966 , n18967 , n18968 , n18969 , n18970 , n18971 , n18972 , n18973 , n18974 , n18975 , n18976 , n18977 , n18978 , n18979 , n18980 , n18981 , n18982 , n18983 , n18984 , n18985 , n18986 , n18987 , n18988 , n18989 , n18990 , n18991 , n18992 , n18993 , n18994 , n18995 , n18996 , n18997 , n18998 , n18999 , n19000 , n19001 , n19002 , n19003 , n19004 , n19005 , n19006 , n19007 , n19008 , n19009 , n19010 , n19011 , n19012 , n19013 , n19014 , n19015 , n19016 , n19017 , n19018 , n19019 , n19020 , n19021 , n19022 , n19023 , n19024 , n19025 , n19026 , n19027 , n19028 , n19029 , n19030 , n19031 , n19032 , n19033 , n19034 , n19035 , n19036 , n19037 , n19038 , n19039 , n19040 , n19041 , n19042 , n19043 , n19044 , n19045 , n19046 , n19047 , n19048 , n19049 , n19050 , n19051 , n19052 , n19053 , n19054 , n19055 , n19056 , n19057 , n19058 , n19059 , n19060 , n19061 , n19062 , n19063 , n19064 , n19065 , n19066 , n19067 , n19068 , n19069 , n19070 , n19071 , n19072 , n19073 , n19074 , n19075 , n19076 , n19077 , n19078 , n19079 , n19080 , n19081 , n19082 , n19083 , n19084 , n19085 , n19086 , n19087 , n19088 , n19089 , n19090 , n19091 , n19092 , n19093 , n19094 , n19095 , n19096 , n19097 , n19098 , n19099 , n19100 , n19101 , n19102 , n19103 , n19104 , n19105 , n19106 , n19107 , n19108 , n19109 , n19110 , n19111 , n19112 , n19113 , n19114 , n19115 , n19116 , n19117 , n19118 , n19119 , n19120 , n19121 , n19122 , n19123 , n19124 , n19125 , n19126 , n19127 , n19128 , n19129 , n19130 , n19131 , n19132 , n19133 , n19134 , n19135 , n19136 , n19137 , n19138 , n19139 , n19140 , n19141 , n19142 , n19143 , n19144 , n19145 , n19146 , n19147 , n19148 , n19149 , n19150 , n19151 , n19152 , n19153 , n19154 , n19155 , n19156 , n19157 , n19158 , n19159 , n19160 , n19161 , n19162 , n19163 , n19164 , n19165 , n19166 , n19167 , n19168 , n19169 , n19170 , n19171 , n19172 , n19173 , n19174 , n19175 , n19176 , n19177 , n19178 , n19179 , n19180 , n19181 , n19182 , n19183 , n19184 , n19185 , n19186 , n19187 , n19188 , n19189 , n19190 , n19191 , n19192 , n19193 , n19194 , n19195 , n19196 , n19197 , n19198 , n19199 , n19200 , n19201 , n19202 , n19203 , n19204 , n19205 , n19206 , n19207 , n19208 , n19209 , n19210 , n19211 , n19212 , n19213 , n19214 , n19215 , n19216 , n19217 , n19218 , n19219 , n19220 , n19221 , n19222 , n19223 , n19224 , n19225 , n19226 , n19227 , n19228 , n19229 , n19230 , n19231 , n19232 , n19233 , n19234 , n19235 , n19236 , n19237 , n19238 , n19239 , n19240 , n19241 , n19242 , n19243 , n19244 , n19245 , n19246 , n19247 , n19248 , n19249 , n19250 , n19251 , n19252 , n19253 , n19254 , n19255 , n19256 , n19257 , n19258 , n19259 , n19260 , n19261 , n19262 , n19263 , n19264 , n19265 , n19266 , n19267 , n19268 , n19269 , n19270 , n19271 , n19272 , n19273 , n19274 , n19275 , n19276 , n19277 , n19278 , n19279 , n19280 , n19281 , n19282 , n19283 , n19284 , n19285 , n19286 , n19287 , n19288 , n19289 , n19290 , n19291 , n19292 , n19293 , n19294 , n19295 , n19296 , n19297 , n19298 , n19299 , n19300 , n19301 , n19302 , n19303 , n19304 , n19305 , n19306 , n19307 , n19308 , n19309 , n19310 , n19311 , n19312 , n19313 , n19314 , n19315 , n19316 , n19317 , n19318 , n19319 , n19320 , n19321 , n19322 , n19323 , n19324 , n19325 , n19326 , n19327 , n19328 , n19329 , n19330 , n19331 , n19332 , n19333 , n19334 , n19335 , n19336 , n19337 , n19338 , n19339 , n19340 , n19341 , n19342 , n19343 , n19344 , n19345 , n19346 , n19347 , n19348 , n19349 , n19350 , n19351 , n19352 , n19353 , n19354 , n19355 , n19356 , n19357 , n19358 , n19359 , n19360 , n19361 , n19362 , n19363 , n19364 , n19365 , n19366 , n19367 , n19368 , n19369 , n19370 , n19371 , n19372 , n19373 , n19374 , n19375 , n19376 , n19377 , n19378 , n19379 , n19380 , n19381 , n19382 , n19383 , n19384 , n19385 , n19386 , n19387 , n19388 , n19389 , n19390 , n19391 , n19392 , n19393 , n19394 , n19395 , n19396 , n19397 , n19398 , n19399 , n19400 , n19401 , n19402 , n19403 , n19404 , n19405 , n19406 , n19407 , n19408 , n19409 , n19410 , n19411 , n19412 , n19413 , n19414 , n19415 , n19416 , n19417 , n19418 , n19419 , n19420 , n19421 , n19422 , n19423 , n19424 , n19425 , n19426 , n19427 , n19428 , n19429 , n19430 , n19431 , n19432 , n19433 , n19434 , n19435 , n19436 , n19437 , n19438 , n19439 , n19440 , n19441 , n19442 , n19443 , n19444 , n19445 , n19446 , n19447 , n19448 , n19449 , n19450 , n19451 , n19452 , n19453 , n19454 , n19455 , n19456 , n19457 , n19458 , n19459 , n19460 , n19461 , n19462 , n19463 , n19464 , n19465 , n19466 , n19467 , n19468 , n19469 , n19470 , n19471 , n19472 , n19473 , n19474 , n19475 , n19476 , n19477 , n19478 , n19479 , n19480 , n19481 , n19482 , n19483 , n19484 , n19485 , n19486 , n19487 , n19488 , n19489 , n19490 , n19491 , n19492 , n19493 , n19494 , n19495 , n19496 , n19497 , n19498 , n19499 , n19500 , n19501 , n19502 , n19503 , n19504 , n19505 , n19506 , n19507 , n19508 , n19509 , n19510 , n19511 , n19512 , n19513 , n19514 , n19515 , n19516 , n19517 , n19518 , n19519 , n19520 , n19521 , n19522 , n19523 , n19524 , n19525 , n19526 , n19527 , n19528 , n19529 , n19530 , n19531 , n19532 , n19533 , n19534 , n19535 , n19536 , n19537 , n19538 , n19539 , n19540 , n19541 , n19542 , n19543 , n19544 , n19545 , n19546 , n19547 , n19548 , n19549 , n19550 , n19551 , n19552 , n19553 , n19554 , n19555 , n19556 , n19557 , n19558 , n19559 , n19560 , n19561 , n19562 , n19563 , n19564 , n19565 , n19566 , n19567 , n19568 , n19569 , n19570 , n19571 , n19572 , n19573 , n19574 , n19575 , n19576 , n19577 , n19578 , n19579 , n19580 , n19581 , n19582 , n19583 , n19584 , n19585 , n19586 , n19587 , n19588 , n19589 , n19590 , n19591 , n19592 , n19593 , n19594 , n19595 , n19596 , n19597 , n19598 , n19599 , n19600 , n19601 , n19602 , n19603 , n19604 , n19605 , n19606 , n19607 , n19608 , n19609 , n19610 , n19611 , n19612 , n19613 , n19614 , n19615 , n19616 , n19617 , n19618 , n19619 , n19620 , n19621 , n19622 , n19623 , n19624 , n19625 , n19626 , n19627 , n19628 , n19629 , n19630 , n19631 , n19632 , n19633 , n19634 , n19635 , n19636 , n19637 , n19638 , n19639 , n19640 , n19641 , n19642 , n19643 , n19644 , n19645 , n19646 , n19647 , n19648 , n19649 , n19650 , n19651 , n19652 , n19653 , n19654 , n19655 , n19656 , n19657 , n19658 , n19659 , n19660 , n19661 , n19662 , n19663 , n19664 , n19665 , n19666 , n19667 , n19668 , n19669 , n19670 , n19671 , n19672 , n19673 , n19674 , n19675 , n19676 , n19677 , n19678 , n19679 , n19680 , n19681 , n19682 , n19683 , n19684 , n19685 , n19686 , n19687 , n19688 , n19689 , n19690 , n19691 , n19692 , n19693 , n19694 , n19695 , n19696 , n19697 , n19698 , n19699 , n19700 , n19701 , n19702 , n19703 , n19704 , n19705 , n19706 , n19707 , n19708 , n19709 , n19710 , n19711 , n19712 , n19713 , n19714 , n19715 , n19716 , n19717 , n19718 , n19719 , n19720 , n19721 , n19722 , n19723 , n19724 , n19725 , n19726 , n19727 , n19728 , n19729 , n19730 , n19731 , n19732 , n19733 , n19734 , n19735 , n19736 , n19737 , n19738 , n19739 , n19740 , n19741 , n19742 , n19743 , n19744 , n19745 , n19746 , n19747 , n19748 , n19749 , n19750 , n19751 , n19752 , n19753 , n19754 , n19755 , n19756 , n19757 , n19758 , n19759 , n19760 , n19761 , n19762 , n19763 , n19764 , n19765 , n19766 , n19767 , n19768 , n19769 , n19770 , n19771 , n19772 , n19773 , n19774 , n19775 , n19776 , n19777 , n19778 , n19779 , n19780 , n19781 , n19782 , n19783 , n19784 , n19785 , n19786 , n19787 , n19788 , n19789 , n19790 , n19791 , n19792 , n19793 , n19794 , n19795 , n19796 , n19797 , n19798 , n19799 , n19800 , n19801 , n19802 , n19803 , n19804 , n19805 , n19806 , n19807 , n19808 , n19809 , n19810 , n19811 , n19812 , n19813 , n19814 , n19815 , n19816 , n19817 , n19818 , n19819 , n19820 , n19821 , n19822 , n19823 , n19824 , n19825 , n19826 , n19827 , n19828 , n19829 , n19830 , n19831 , n19832 , n19833 , n19834 , n19835 , n19836 , n19837 , n19838 , n19839 , n19840 , n19841 , n19842 , n19843 , n19844 , n19845 , n19846 , n19847 , n19848 , n19849 , n19850 , n19851 , n19852 , n19853 , n19854 , n19855 , n19856 , n19857 , n19858 , n19859 , n19860 , n19861 , n19862 , n19863 , n19864 , n19865 , n19866 , n19867 , n19868 , n19869 , n19870 , n19871 , n19872 , n19873 , n19874 , n19875 , n19876 , n19877 , n19878 , n19879 , n19880 , n19881 , n19882 , n19883 , n19884 , n19885 , n19886 , n19887 , n19888 , n19889 , n19890 , n19891 , n19892 , n19893 , n19894 , n19895 , n19896 , n19897 , n19898 , n19899 , n19900 , n19901 , n19902 , n19903 , n19904 , n19905 , n19906 , n19907 , n19908 , n19909 , n19910 , n19911 , n19912 , n19913 , n19914 , n19915 , n19916 , n19917 , n19918 , n19919 , n19920 , n19921 , n19922 , n19923 , n19924 , n19925 , n19926 , n19927 , n19928 , n19929 , n19930 , n19931 , n19932 , n19933 , n19934 , n19935 , n19936 , n19937 , n19938 , n19939 , n19940 , n19941 , n19942 , n19943 , n19944 , n19945 , n19946 , n19947 , n19948 , n19949 , n19950 , n19951 , n19952 , n19953 , n19954 , n19955 , n19956 , n19957 , n19958 , n19959 , n19960 , n19961 , n19962 , n19963 , n19964 , n19965 , n19966 , n19967 , n19968 , n19969 , n19970 , n19971 , n19972 , n19973 , n19974 , n19975 , n19976 , n19977 , n19978 , n19979 , n19980 , n19981 , n19982 , n19983 , n19984 , n19985 , n19986 , n19987 , n19988 , n19989 , n19990 , n19991 , n19992 , n19993 , n19994 , n19995 , n19996 , n19997 , n19998 , n19999 , n20000 , n20001 , n20002 , n20003 , n20004 , n20005 , n20006 , n20007 , n20008 , n20009 , n20010 , n20011 , n20012 , n20013 , n20014 , n20015 , n20016 , n20017 , n20018 , n20019 , n20020 , n20021 , n20022 , n20023 , n20024 , n20025 , n20026 , n20027 , n20028 , n20029 , n20030 , n20031 , n20032 , n20033 , n20034 , n20035 , n20036 , n20037 , n20038 , n20039 , n20040 , n20041 , n20042 , n20043 , n20044 , n20045 , n20046 , n20047 , n20048 , n20049 , n20050 , n20051 , n20052 , n20053 , n20054 , n20055 , n20056 , n20057 , n20058 , n20059 , n20060 , n20061 , n20062 , n20063 , n20064 , n20065 , n20066 , n20067 , n20068 , n20069 , n20070 , n20071 , n20072 , n20073 , n20074 , n20075 , n20076 , n20077 , n20078 , n20079 , n20080 , n20081 , n20082 , n20083 , n20084 , n20085 , n20086 , n20087 , n20088 , n20089 , n20090 , n20091 , n20092 , n20093 , n20094 , n20095 , n20096 , n20097 , n20098 , n20099 , n20100 , n20101 , n20102 , n20103 , n20104 , n20105 , n20106 , n20107 , n20108 , n20109 , n20110 , n20111 , n20112 , n20113 , n20114 , n20115 , n20116 , n20117 , n20118 , n20119 , n20120 , n20121 , n20122 , n20123 , n20124 , n20125 , n20126 , n20127 , n20128 , n20129 , n20130 , n20131 , n20132 , n20133 , n20134 , n20135 , n20136 , n20137 , n20138 , n20139 , n20140 , n20141 , n20142 , n20143 , n20144 , n20145 , n20146 , n20147 , n20148 , n20149 , n20150 , n20151 , n20152 , n20153 , n20154 , n20155 , n20156 , n20157 , n20158 , n20159 , n20160 , n20161 , n20162 , n20163 , n20164 , n20165 , n20166 , n20167 , n20168 , n20169 , n20170 , n20171 , n20172 , n20173 , n20174 , n20175 , n20176 , n20177 , n20178 , n20179 , n20180 , n20181 , n20182 , n20183 , n20184 , n20185 , n20186 , n20187 , n20188 , n20189 , n20190 , n20191 , n20192 , n20193 , n20194 , n20195 , n20196 , n20197 , n20198 , n20199 , n20200 , n20201 , n20202 , n20203 , n20204 , n20205 , n20206 , n20207 , n20208 , n20209 , n20210 , n20211 , n20212 , n20213 , n20214 , n20215 , n20216 , n20217 , n20218 , n20219 , n20220 , n20221 , n20222 , n20223 , n20224 , n20225 , n20226 , n20227 , n20228 , n20229 , n20230 , n20231 , n20232 , n20233 , n20234 , n20235 , n20236 , n20237 , n20238 , n20239 , n20240 , n20241 , n20242 , n20243 , n20244 , n20245 , n20246 , n20247 , n20248 , n20249 , n20250 , n20251 , n20252 , n20253 , n20254 , n20255 , n20256 , n20257 , n20258 , n20259 , n20260 , n20261 , n20262 , n20263 , n20264 , n20265 , n20266 , n20267 , n20268 , n20269 , n20270 , n20271 , n20272 , n20273 , n20274 , n20275 , n20276 , n20277 , n20278 , n20279 , n20280 , n20281 , n20282 , n20283 , n20284 , n20285 , n20286 , n20287 , n20288 , n20289 , n20290 , n20291 , n20292 , n20293 , n20294 , n20295 , n20296 , n20297 , n20298 , n20299 , n20300 , n20301 , n20302 , n20303 , n20304 , n20305 , n20306 , n20307 , n20308 , n20309 , n20310 , n20311 , n20312 , n20313 , n20314 , n20315 , n20316 , n20317 , n20318 , n20319 , n20320 , n20321 , n20322 , n20323 , n20324 , n20325 , n20326 , n20327 , n20328 , n20329 , n20330 , n20331 , n20332 , n20333 , n20334 , n20335 , n20336 , n20337 , n20338 , n20339 , n20340 , n20341 , n20342 , n20343 , n20344 , n20345 , n20346 , n20347 , n20348 , n20349 , n20350 , n20351 , n20352 , n20353 , n20354 , n20355 , n20356 , n20357 , n20358 , n20359 , n20360 , n20361 , n20362 , n20363 , n20364 , n20365 , n20366 , n20367 , n20368 , n20369 , n20370 , n20371 , n20372 , n20373 , n20374 , n20375 , n20376 , n20377 , n20378 , n20379 , n20380 , n20381 , n20382 , n20383 , n20384 , n20385 , n20386 , n20387 , n20388 , n20389 , n20390 , n20391 , n20392 , n20393 , n20394 , n20395 , n20396 , n20397 , n20398 , n20399 , n20400 , n20401 , n20402 , n20403 , n20404 , n20405 , n20406 , n20407 , n20408 , n20409 , n20410 , n20411 , n20412 , n20413 , n20414 , n20415 , n20416 , n20417 , n20418 , n20419 , n20420 , n20421 , n20422 , n20423 , n20424 , n20425 , n20426 , n20427 , n20428 , n20429 , n20430 , n20431 , n20432 , n20433 , n20434 , n20435 , n20436 , n20437 , n20438 , n20439 , n20440 , n20441 , n20442 , n20443 , n20444 , n20445 , n20446 , n20447 , n20448 , n20449 , n20450 , n20451 , n20452 , n20453 , n20454 , n20455 , n20456 , n20457 , n20458 , n20459 , n20460 , n20461 , n20462 , n20463 , n20464 , n20465 , n20466 , n20467 , n20468 , n20469 , n20470 , n20471 , n20472 , n20473 , n20474 , n20475 , n20476 , n20477 , n20478 , n20479 , n20480 , n20481 , n20482 , n20483 , n20484 , n20485 , n20486 , n20487 , n20488 , n20489 , n20490 , n20491 , n20492 , n20493 , n20494 , n20495 , n20496 , n20497 , n20498 , n20499 , n20500 , n20501 , n20502 , n20503 , n20504 , n20505 , n20506 , n20507 , n20508 , n20509 , n20510 , n20511 , n20512 , n20513 , n20514 , n20515 , n20516 , n20517 , n20518 , n20519 , n20520 , n20521 , n20522 , n20523 , n20524 , n20525 , n20526 , n20527 , n20528 , n20529 , n20530 , n20531 , n20532 , n20533 , n20534 , n20535 , n20536 , n20537 , n20538 , n20539 , n20540 , n20541 , n20542 , n20543 , n20544 , n20545 , n20546 , n20547 , n20548 , n20549 , n20550 , n20551 , n20552 , n20553 , n20554 , n20555 , n20556 , n20557 , n20558 , n20559 , n20560 , n20561 , n20562 , n20563 , n20564 , n20565 , n20566 , n20567 , n20568 , n20569 , n20570 , n20571 , n20572 , n20573 , n20574 , n20575 , n20576 , n20577 , n20578 , n20579 , n20580 , n20581 , n20582 , n20583 , n20584 , n20585 , n20586 , n20587 , n20588 , n20589 , n20590 , n20591 , n20592 , n20593 , n20594 , n20595 , n20596 , n20597 , n20598 , n20599 , n20600 , n20601 , n20602 , n20603 , n20604 , n20605 , n20606 , n20607 , n20608 , n20609 , n20610 , n20611 , n20612 , n20613 , n20614 , n20615 , n20616 , n20617 , n20618 , n20619 , n20620 , n20621 , n20622 , n20623 , n20624 , n20625 , n20626 , n20627 , n20628 , n20629 , n20630 , n20631 , n20632 , n20633 , n20634 , n20635 , n20636 , n20637 , n20638 , n20639 , n20640 , n20641 , n20642 , n20643 , n20644 , n20645 , n20646 , n20647 , n20648 , n20649 , n20650 , n20651 , n20652 , n20653 , n20654 , n20655 , n20656 , n20657 , n20658 , n20659 , n20660 , n20661 , n20662 , n20663 , n20664 , n20665 , n20666 , n20667 , n20668 , n20669 , n20670 , n20671 , n20672 , n20673 , n20674 , n20675 , n20676 , n20677 , n20678 , n20679 , n20680 , n20681 , n20682 , n20683 , n20684 , n20685 , n20686 , n20687 , n20688 , n20689 , n20690 , n20691 , n20692 , n20693 , n20694 , n20695 , n20696 , n20697 , n20698 , n20699 , n20700 , n20701 , n20702 , n20703 , n20704 , n20705 , n20706 , n20707 , n20708 , n20709 , n20710 , n20711 , n20712 , n20713 , n20714 , n20715 , n20716 , n20717 , n20718 , n20719 , n20720 , n20721 , n20722 , n20723 , n20724 , n20725 , n20726 , n20727 , n20728 , n20729 , n20730 , n20731 , n20732 , n20733 , n20734 , n20735 , n20736 , n20737 , n20738 , n20739 , n20740 , n20741 , n20742 , n20743 , n20744 , n20745 , n20746 , n20747 , n20748 , n20749 , n20750 , n20751 , n20752 , n20753 , n20754 , n20755 , n20756 , n20757 , n20758 , n20759 , n20760 , n20761 , n20762 , n20763 , n20764 , n20765 , n20766 , n20767 , n20768 , n20769 , n20770 , n20771 , n20772 , n20773 , n20774 , n20775 , n20776 , n20777 , n20778 , n20779 , n20780 , n20781 , n20782 , n20783 , n20784 , n20785 , n20786 , n20787 , n20788 , n20789 , n20790 , n20791 , n20792 , n20793 , n20794 , n20795 , n20796 , n20797 , n20798 , n20799 , n20800 , n20801 , n20802 , n20803 , n20804 , n20805 , n20806 , n20807 , n20808 , n20809 , n20810 , n20811 , n20812 , n20813 , n20814 , n20815 , n20816 , n20817 , n20818 , n20819 , n20820 , n20821 , n20822 , n20823 , n20824 , n20825 , n20826 , n20827 , n20828 , n20829 , n20830 , n20831 , n20832 , n20833 , n20834 , n20835 , n20836 , n20837 , n20838 , n20839 , n20840 , n20841 , n20842 , n20843 , n20844 , n20845 , n20846 , n20847 , n20848 , n20849 , n20850 , n20851 , n20852 , n20853 , n20854 , n20855 , n20856 , n20857 , n20858 , n20859 , n20860 , n20861 , n20862 , n20863 , n20864 , n20865 , n20866 , n20867 , n20868 , n20869 , n20870 , n20871 , n20872 , n20873 , n20874 , n20875 , n20876 , n20877 , n20878 , n20879 , n20880 , n20881 , n20882 , n20883 , n20884 , n20885 , n20886 , n20887 , n20888 , n20889 , n20890 , n20891 , n20892 , n20893 , n20894 , n20895 , n20896 , n20897 , n20898 , n20899 , n20900 , n20901 , n20902 , n20903 , n20904 , n20905 , n20906 , n20907 , n20908 , n20909 , n20910 , n20911 , n20912 , n20913 , n20914 , n20915 , n20916 , n20917 , n20918 , n20919 , n20920 , n20921 , n20922 , n20923 , n20924 , n20925 , n20926 , n20927 , n20928 , n20929 , n20930 , n20931 , n20932 , n20933 , n20934 , n20935 , n20936 , n20937 , n20938 , n20939 , n20940 , n20941 , n20942 , n20943 , n20944 , n20945 , n20946 , n20947 , n20948 , n20949 , n20950 , n20951 , n20952 , n20953 , n20954 , n20955 , n20956 , n20957 , n20958 , n20959 , n20960 , n20961 , n20962 , n20963 , n20964 , n20965 , n20966 , n20967 , n20968 , n20969 , n20970 , n20971 , n20972 , n20973 , n20974 , n20975 , n20976 , n20977 , n20978 , n20979 , n20980 , n20981 , n20982 , n20983 , n20984 , n20985 , n20986 , n20987 , n20988 , n20989 , n20990 , n20991 , n20992 , n20993 , n20994 , n20995 , n20996 , n20997 , n20998 , n20999 , n21000 , n21001 , n21002 , n21003 , n21004 , n21005 , n21006 , n21007 , n21008 , n21009 , n21010 , n21011 , n21012 , n21013 , n21014 , n21015 , n21016 , n21017 , n21018 , n21019 , n21020 , n21021 , n21022 , n21023 , n21024 , n21025 , n21026 , n21027 , n21028 , n21029 , n21030 , n21031 , n21032 , n21033 , n21034 , n21035 , n21036 , n21037 , n21038 , n21039 , n21040 , n21041 , n21042 , n21043 , n21044 , n21045 , n21046 , n21047 , n21048 , n21049 , n21050 , n21051 , n21052 , n21053 , n21054 , n21055 , n21056 , n21057 , n21058 , n21059 , n21060 , n21061 , n21062 , n21063 , n21064 , n21065 , n21066 , n21067 , n21068 , n21069 , n21070 , n21071 , n21072 , n21073 , n21074 , n21075 , n21076 , n21077 , n21078 , n21079 , n21080 , n21081 , n21082 , n21083 , n21084 , n21085 , n21086 , n21087 , n21088 , n21089 , n21090 , n21091 , n21092 , n21093 , n21094 , n21095 , n21096 , n21097 , n21098 , n21099 , n21100 , n21101 , n21102 , n21103 , n21104 , n21105 , n21106 , n21107 , n21108 , n21109 , n21110 , n21111 , n21112 , n21113 , n21114 , n21115 , n21116 , n21117 , n21118 , n21119 , n21120 , n21121 , n21122 , n21123 , n21124 , n21125 , n21126 , n21127 , n21128 , n21129 , n21130 , n21131 , n21132 , n21133 , n21134 , n21135 , n21136 , n21137 , n21138 , n21139 , n21140 , n21141 , n21142 , n21143 , n21144 , n21145 , n21146 , n21147 , n21148 , n21149 , n21150 , n21151 , n21152 , n21153 , n21154 , n21155 , n21156 , n21157 , n21158 , n21159 , n21160 , n21161 , n21162 , n21163 , n21164 , n21165 , n21166 , n21167 , n21168 , n21169 , n21170 , n21171 , n21172 , n21173 , n21174 , n21175 , n21176 , n21177 , n21178 , n21179 , n21180 , n21181 , n21182 , n21183 , n21184 , n21185 , n21186 , n21187 , n21188 , n21189 , n21190 , n21191 , n21192 , n21193 , n21194 , n21195 , n21196 , n21197 , n21198 , n21199 , n21200 , n21201 , n21202 , n21203 , n21204 , n21205 , n21206 , n21207 , n21208 , n21209 , n21210 , n21211 , n21212 , n21213 , n21214 , n21215 , n21216 , n21217 , n21218 , n21219 , n21220 , n21221 , n21222 , n21223 , n21224 , n21225 , n21226 , n21227 , n21228 , n21229 , n21230 , n21231 , n21232 , n21233 , n21234 , n21235 , n21236 , n21237 , n21238 , n21239 , n21240 , n21241 , n21242 , n21243 , n21244 , n21245 , n21246 , n21247 , n21248 , n21249 , n21250 , n21251 , n21252 , n21253 , n21254 , n21255 , n21256 , n21257 , n21258 , n21259 , n21260 , n21261 , n21262 , n21263 , n21264 , n21265 , n21266 , n21267 , n21268 , n21269 , n21270 , n21271 , n21272 , n21273 , n21274 , n21275 , n21276 , n21277 , n21278 , n21279 , n21280 , n21281 , n21282 , n21283 , n21284 , n21285 , n21286 , n21287 , n21288 , n21289 , n21290 , n21291 , n21292 , n21293 , n21294 , n21295 , n21296 , n21297 , n21298 , n21299 , n21300 , n21301 , n21302 , n21303 , n21304 , n21305 , n21306 , n21307 , n21308 , n21309 , n21310 , n21311 , n21312 , n21313 , n21314 , n21315 , n21316 , n21317 , n21318 , n21319 , n21320 , n21321 , n21322 , n21323 , n21324 , n21325 , n21326 , n21327 , n21328 , n21329 , n21330 , n21331 , n21332 , n21333 , n21334 , n21335 , n21336 , n21337 , n21338 , n21339 , n21340 , n21341 , n21342 , n21343 , n21344 , n21345 , n21346 , n21347 , n21348 , n21349 , n21350 , n21351 , n21352 , n21353 , n21354 , n21355 , n21356 , n21357 , n21358 , n21359 , n21360 , n21361 , n21362 , n21363 , n21364 , n21365 , n21366 , n21367 , n21368 , n21369 , n21370 , n21371 , n21372 , n21373 , n21374 , n21375 , n21376 , n21377 , n21378 , n21379 , n21380 , n21381 , n21382 , n21383 , n21384 , n21385 , n21386 , n21387 , n21388 , n21389 , n21390 , n21391 , n21392 , n21393 , n21394 , n21395 , n21396 , n21397 , n21398 , n21399 , n21400 , n21401 , n21402 , n21403 , n21404 , n21405 , n21406 , n21407 , n21408 , n21409 , n21410 , n21411 , n21412 , n21413 , n21414 , n21415 , n21416 , n21417 , n21418 , n21419 , n21420 , n21421 , n21422 , n21423 , n21424 , n21425 , n21426 , n21427 , n21428 , n21429 , n21430 , n21431 , n21432 , n21433 , n21434 , n21435 , n21436 , n21437 , n21438 , n21439 , n21440 , n21441 , n21442 , n21443 , n21444 , n21445 , n21446 , n21447 , n21448 , n21449 , n21450 , n21451 , n21452 , n21453 , n21454 , n21455 , n21456 , n21457 , n21458 , n21459 , n21460 , n21461 , n21462 , n21463 , n21464 , n21465 , n21466 , n21467 , n21468 , n21469 , n21470 , n21471 , n21472 , n21473 , n21474 , n21475 , n21476 , n21477 , n21478 , n21479 , n21480 , n21481 , n21482 , n21483 , n21484 , n21485 , n21486 , n21487 , n21488 , n21489 , n21490 , n21491 , n21492 , n21493 , n21494 , n21495 , n21496 , n21497 , n21498 , n21499 , n21500 , n21501 , n21502 , n21503 , n21504 , n21505 , n21506 , n21507 , n21508 , n21509 , n21510 , n21511 , n21512 , n21513 , n21514 , n21515 , n21516 , n21517 , n21518 , n21519 , n21520 , n21521 , n21522 , n21523 , n21524 , n21525 , n21526 , n21527 , n21528 , n21529 , n21530 , n21531 , n21532 , n21533 , n21534 , n21535 , n21536 , n21537 , n21538 , n21539 , n21540 , n21541 , n21542 , n21543 , n21544 , n21545 , n21546 , n21547 , n21548 , n21549 , n21550 , n21551 , n21552 , n21553 , n21554 , n21555 , n21556 , n21557 , n21558 , n21559 , n21560 , n21561 , n21562 , n21563 , n21564 , n21565 , n21566 , n21567 , n21568 , n21569 , n21570 , n21571 , n21572 , n21573 , n21574 , n21575 , n21576 , n21577 , n21578 , n21579 , n21580 , n21581 , n21582 , n21583 , n21584 , n21585 , n21586 , n21587 , n21588 , n21589 , n21590 , n21591 , n21592 , n21593 , n21594 , n21595 , n21596 , n21597 , n21598 , n21599 , n21600 , n21601 , n21602 , n21603 , n21604 , n21605 , n21606 , n21607 , n21608 , n21609 , n21610 , n21611 , n21612 , n21613 , n21614 , n21615 , n21616 , n21617 , n21618 , n21619 , n21620 , n21621 , n21622 , n21623 , n21624 , n21625 , n21626 , n21627 , n21628 , n21629 , n21630 , n21631 , n21632 , n21633 , n21634 , n21635 , n21636 , n21637 , n21638 , n21639 , n21640 , n21641 , n21642 , n21643 , n21644 , n21645 , n21646 , n21647 , n21648 , n21649 , n21650 , n21651 , n21652 , n21653 , n21654 , n21655 , n21656 , n21657 , n21658 , n21659 , n21660 , n21661 , n21662 , n21663 , n21664 , n21665 , n21666 , n21667 , n21668 , n21669 , n21670 , n21671 , n21672 , n21673 , n21674 , n21675 , n21676 , n21677 , n21678 , n21679 , n21680 , n21681 , n21682 , n21683 , n21684 , n21685 , n21686 , n21687 , n21688 , n21689 , n21690 , n21691 , n21692 , n21693 , n21694 , n21695 , n21696 , n21697 , n21698 , n21699 , n21700 , n21701 , n21702 , n21703 , n21704 , n21705 , n21706 , n21707 , n21708 , n21709 , n21710 , n21711 , n21712 , n21713 , n21714 , n21715 , n21716 , n21717 , n21718 , n21719 , n21720 , n21721 , n21722 , n21723 , n21724 , n21725 , n21726 , n21727 , n21728 , n21729 , n21730 , n21731 , n21732 , n21733 , n21734 , n21735 , n21736 , n21737 , n21738 , n21739 , n21740 , n21741 , n21742 , n21743 , n21744 , n21745 , n21746 , n21747 , n21748 , n21749 , n21750 , n21751 , n21752 , n21753 , n21754 , n21755 , n21756 , n21757 , n21758 , n21759 , n21760 , n21761 , n21762 , n21763 , n21764 , n21765 , n21766 , n21767 , n21768 , n21769 , n21770 , n21771 , n21772 , n21773 , n21774 , n21775 , n21776 , n21777 , n21778 , n21779 , n21780 , n21781 , n21782 , n21783 , n21784 , n21785 , n21786 , n21787 , n21788 , n21789 , n21790 , n21791 , n21792 , n21793 , n21794 , n21795 , n21796 , n21797 , n21798 , n21799 , n21800 , n21801 , n21802 , n21803 , n21804 , n21805 , n21806 , n21807 , n21808 , n21809 , n21810 , n21811 , n21812 , n21813 , n21814 , n21815 , n21816 , n21817 , n21818 , n21819 , n21820 , n21821 , n21822 , n21823 , n21824 , n21825 , n21826 , n21827 , n21828 , n21829 , n21830 , n21831 , n21832 , n21833 , n21834 , n21835 , n21836 , n21837 , n21838 , n21839 , n21840 , n21841 , n21842 , n21843 , n21844 , n21845 , n21846 , n21847 , n21848 , n21849 , n21850 , n21851 , n21852 , n21853 , n21854 , n21855 , n21856 , n21857 , n21858 , n21859 , n21860 , n21861 , n21862 , n21863 , n21864 , n21865 , n21866 , n21867 , n21868 , n21869 , n21870 , n21871 , n21872 , n21873 , n21874 , n21875 , n21876 , n21877 , n21878 , n21879 , n21880 , n21881 , n21882 , n21883 , n21884 , n21885 , n21886 , n21887 , n21888 , n21889 , n21890 , n21891 , n21892 , n21893 , n21894 , n21895 , n21896 , n21897 , n21898 , n21899 , n21900 , n21901 , n21902 , n21903 , n21904 , n21905 , n21906 , n21907 , n21908 , n21909 , n21910 , n21911 , n21912 , n21913 , n21914 , n21915 , n21916 , n21917 , n21918 , n21919 , n21920 , n21921 , n21922 , n21923 , n21924 , n21925 , n21926 , n21927 , n21928 , n21929 , n21930 , n21931 , n21932 , n21933 , n21934 , n21935 , n21936 , n21937 , n21938 , n21939 , n21940 , n21941 , n21942 , n21943 , n21944 , n21945 , n21946 , n21947 , n21948 , n21949 , n21950 , n21951 , n21952 , n21953 , n21954 , n21955 , n21956 , n21957 , n21958 , n21959 , n21960 , n21961 , n21962 , n21963 , n21964 , n21965 , n21966 , n21967 , n21968 , n21969 , n21970 , n21971 , n21972 , n21973 , n21974 , n21975 , n21976 , n21977 , n21978 , n21979 , n21980 , n21981 , n21982 , n21983 , n21984 , n21985 , n21986 , n21987 , n21988 , n21989 , n21990 , n21991 , n21992 , n21993 , n21994 , n21995 , n21996 , n21997 , n21998 , n21999 , n22000 , n22001 , n22002 , n22003 , n22004 , n22005 , n22006 , n22007 , n22008 , n22009 , n22010 , n22011 , n22012 , n22013 , n22014 , n22015 , n22016 , n22017 , n22018 , n22019 , n22020 , n22021 , n22022 , n22023 , n22024 , n22025 , n22026 , n22027 , n22028 , n22029 , n22030 , n22031 , n22032 , n22033 , n22034 , n22035 , n22036 , n22037 , n22038 , n22039 , n22040 , n22041 , n22042 , n22043 , n22044 , n22045 , n22046 , n22047 , n22048 , n22049 , n22050 , n22051 , n22052 , n22053 , n22054 , n22055 , n22056 , n22057 , n22058 , n22059 , n22060 , n22061 , n22062 , n22063 , n22064 , n22065 , n22066 , n22067 , n22068 , n22069 , n22070 , n22071 , n22072 , n22073 , n22074 , n22075 , n22076 , n22077 , n22078 , n22079 , n22080 , n22081 , n22082 , n22083 , n22084 , n22085 , n22086 , n22087 , n22088 , n22089 , n22090 , n22091 , n22092 , n22093 , n22094 , n22095 , n22096 , n22097 , n22098 , n22099 , n22100 , n22101 , n22102 , n22103 , n22104 , n22105 , n22106 , n22107 , n22108 , n22109 , n22110 , n22111 , n22112 , n22113 , n22114 , n22115 , n22116 , n22117 , n22118 , n22119 , n22120 , n22121 , n22122 , n22123 , n22124 , n22125 , n22126 , n22127 , n22128 , n22129 , n22130 , n22131 , n22132 , n22133 , n22134 , n22135 , n22136 , n22137 , n22138 , n22139 , n22140 , n22141 , n22142 , n22143 , n22144 , n22145 , n22146 , n22147 , n22148 , n22149 , n22150 , n22151 , n22152 , n22153 , n22154 , n22155 , n22156 , n22157 , n22158 , n22159 , n22160 , n22161 , n22162 , n22163 , n22164 , n22165 , n22166 , n22167 , n22168 , n22169 , n22170 , n22171 , n22172 , n22173 , n22174 , n22175 , n22176 , n22177 , n22178 , n22179 , n22180 , n22181 , n22182 , n22183 , n22184 , n22185 , n22186 , n22187 , n22188 , n22189 , n22190 , n22191 , n22192 , n22193 , n22194 , n22195 , n22196 , n22197 , n22198 , n22199 , n22200 , n22201 , n22202 , n22203 , n22204 , n22205 , n22206 , n22207 , n22208 , n22209 , n22210 , n22211 , n22212 , n22213 , n22214 , n22215 , n22216 , n22217 , n22218 , n22219 , n22220 , n22221 , n22222 , n22223 , n22224 , n22225 , n22226 , n22227 , n22228 , n22229 , n22230 , n22231 , n22232 , n22233 , n22234 , n22235 , n22236 , n22237 , n22238 , n22239 , n22240 , n22241 , n22242 , n22243 , n22244 , n22245 , n22246 , n22247 , n22248 , n22249 , n22250 , n22251 , n22252 , n22253 , n22254 , n22255 , n22256 , n22257 , n22258 , n22259 , n22260 , n22261 , n22262 , n22263 , n22264 , n22265 , n22266 , n22267 , n22268 , n22269 , n22270 , n22271 , n22272 , n22273 , n22274 , n22275 , n22276 , n22277 , n22278 , n22279 , n22280 , n22281 , n22282 , n22283 , n22284 , n22285 , n22286 , n22287 , n22288 , n22289 , n22290 , n22291 , n22292 , n22293 , n22294 , n22295 , n22296 , n22297 , n22298 , n22299 , n22300 , n22301 , n22302 , n22303 , n22304 , n22305 , n22306 , n22307 , n22308 , n22309 , n22310 , n22311 , n22312 , n22313 , n22314 , n22315 , n22316 , n22317 , n22318 , n22319 , n22320 , n22321 , n22322 , n22323 , n22324 , n22325 , n22326 , n22327 , n22328 , n22329 , n22330 , n22331 , n22332 , n22333 , n22334 , n22335 , n22336 , n22337 , n22338 , n22339 , n22340 , n22341 , n22342 , n22343 , n22344 , n22345 , n22346 , n22347 , n22348 , n22349 , n22350 , n22351 , n22352 , n22353 , n22354 , n22355 , n22356 , n22357 , n22358 , n22359 , n22360 , n22361 , n22362 , n22363 , n22364 , n22365 , n22366 , n22367 , n22368 , n22369 , n22370 , n22371 , n22372 , n22373 , n22374 , n22375 , n22376 , n22377 , n22378 , n22379 , n22380 , n22381 , n22382 , n22383 , n22384 , n22385 , n22386 , n22387 , n22388 , n22389 , n22390 , n22391 , n22392 , n22393 , n22394 , n22395 , n22396 , n22397 , n22398 , n22399 , n22400 , n22401 , n22402 , n22403 , n22404 , n22405 , n22406 , n22407 , n22408 , n22409 , n22410 , n22411 , n22412 , n22413 , n22414 , n22415 , n22416 , n22417 , n22418 , n22419 , n22420 , n22421 , n22422 , n22423 , n22424 , n22425 , n22426 , n22427 , n22428 , n22429 , n22430 , n22431 , n22432 , n22433 , n22434 , n22435 , n22436 , n22437 , n22438 , n22439 , n22440 , n22441 , n22442 , n22443 , n22444 , n22445 , n22446 , n22447 , n22448 , n22449 , n22450 , n22451 , n22452 , n22453 , n22454 , n22455 , n22456 , n22457 , n22458 , n22459 , n22460 , n22461 , n22462 , n22463 , n22464 , n22465 , n22466 , n22467 , n22468 , n22469 , n22470 , n22471 , n22472 , n22473 , n22474 , n22475 , n22476 , n22477 , n22478 , n22479 , n22480 , n22481 , n22482 , n22483 , n22484 , n22485 , n22486 , n22487 , n22488 , n22489 , n22490 , n22491 , n22492 , n22493 , n22494 , n22495 , n22496 , n22497 , n22498 , n22499 , n22500 , n22501 , n22502 , n22503 , n22504 , n22505 , n22506 , n22507 , n22508 , n22509 , n22510 , n22511 , n22512 , n22513 , n22514 , n22515 , n22516 , n22517 , n22518 , n22519 , n22520 , n22521 , n22522 , n22523 , n22524 , n22525 , n22526 , n22527 , n22528 , n22529 , n22530 , n22531 , n22532 , n22533 , n22534 , n22535 , n22536 , n22537 , n22538 , n22539 , n22540 , n22541 , n22542 , n22543 , n22544 , n22545 , n22546 , n22547 , n22548 , n22549 , n22550 , n22551 , n22552 , n22553 , n22554 , n22555 , n22556 , n22557 , n22558 , n22559 , n22560 , n22561 , n22562 , n22563 , n22564 , n22565 , n22566 , n22567 , n22568 , n22569 , n22570 , n22571 , n22572 , n22573 , n22574 , n22575 , n22576 , n22577 , n22578 , n22579 , n22580 , n22581 , n22582 , n22583 , n22584 , n22585 , n22586 , n22587 , n22588 , n22589 , n22590 , n22591 , n22592 , n22593 , n22594 , n22595 , n22596 , n22597 , n22598 , n22599 , n22600 , n22601 , n22602 , n22603 , n22604 , n22605 , n22606 , n22607 , n22608 , n22609 , n22610 , n22611 , n22612 , n22613 , n22614 , n22615 , n22616 , n22617 , n22618 , n22619 , n22620 , n22621 , n22622 , n22623 , n22624 , n22625 , n22626 , n22627 , n22628 , n22629 , n22630 , n22631 , n22632 , n22633 , n22634 , n22635 , n22636 , n22637 , n22638 , n22639 , n22640 , n22641 , n22642 , n22643 , n22644 , n22645 , n22646 , n22647 , n22648 , n22649 , n22650 , n22651 , n22652 , n22653 , n22654 , n22655 , n22656 , n22657 , n22658 , n22659 , n22660 , n22661 , n22662 , n22663 , n22664 , n22665 , n22666 , n22667 , n22668 , n22669 , n22670 , n22671 , n22672 , n22673 , n22674 , n22675 , n22676 , n22677 , n22678 , n22679 , n22680 , n22681 , n22682 , n22683 , n22684 , n22685 , n22686 , n22687 , n22688 , n22689 , n22690 , n22691 , n22692 , n22693 , n22694 , n22695 , n22696 , n22697 , n22698 , n22699 , n22700 , n22701 , n22702 , n22703 , n22704 , n22705 , n22706 , n22707 , n22708 , n22709 , n22710 , n22711 , n22712 , n22713 , n22714 , n22715 , n22716 , n22717 , n22718 , n22719 , n22720 , n22721 , n22722 , n22723 , n22724 , n22725 , n22726 , n22727 , n22728 , n22729 , n22730 , n22731 , n22732 , n22733 , n22734 , n22735 , n22736 , n22737 , n22738 , n22739 , n22740 , n22741 , n22742 , n22743 , n22744 , n22745 , n22746 , n22747 , n22748 , n22749 , n22750 , n22751 , n22752 , n22753 , n22754 , n22755 , n22756 , n22757 , n22758 , n22759 , n22760 , n22761 , n22762 , n22763 , n22764 , n22765 , n22766 , n22767 , n22768 , n22769 , n22770 , n22771 , n22772 , n22773 , n22774 , n22775 , n22776 , n22777 , n22778 , n22779 , n22780 , n22781 , n22782 , n22783 , n22784 , n22785 , n22786 , n22787 , n22788 , n22789 , n22790 , n22791 , n22792 , n22793 , n22794 , n22795 , n22796 , n22797 , n22798 , n22799 , n22800 , n22801 , n22802 , n22803 , n22804 , n22805 , n22806 , n22807 , n22808 , n22809 , n22810 , n22811 , n22812 , n22813 , n22814 , n22815 , n22816 , n22817 , n22818 , n22819 , n22820 , n22821 , n22822 , n22823 , n22824 , n22825 , n22826 , n22827 , n22828 , n22829 , n22830 , n22831 , n22832 , n22833 , n22834 , n22835 , n22836 , n22837 , n22838 , n22839 , n22840 , n22841 , n22842 , n22843 , n22844 , n22845 , n22846 , n22847 , n22848 , n22849 , n22850 , n22851 , n22852 , n22853 , n22854 , n22855 , n22856 , n22857 , n22858 , n22859 , n22860 , n22861 , n22862 , n22863 , n22864 , n22865 , n22866 , n22867 , n22868 , n22869 , n22870 , n22871 , n22872 , n22873 , n22874 , n22875 , n22876 , n22877 , n22878 , n22879 , n22880 , n22881 , n22882 , n22883 , n22884 , n22885 , n22886 , n22887 , n22888 , n22889 , n22890 , n22891 , n22892 , n22893 , n22894 , n22895 , n22896 , n22897 , n22898 , n22899 , n22900 , n22901 , n22902 , n22903 , n22904 , n22905 , n22906 , n22907 , n22908 , n22909 , n22910 , n22911 , n22912 , n22913 , n22914 , n22915 , n22916 , n22917 , n22918 , n22919 , n22920 , n22921 , n22922 , n22923 , n22924 , n22925 , n22926 , n22927 , n22928 , n22929 , n22930 , n22931 , n22932 , n22933 , n22934 , n22935 , n22936 , n22937 , n22938 , n22939 , n22940 , n22941 , n22942 , n22943 , n22944 , n22945 , n22946 , n22947 , n22948 , n22949 , n22950 , n22951 , n22952 , n22953 , n22954 , n22955 , n22956 , n22957 , n22958 , n22959 , n22960 , n22961 , n22962 , n22963 , n22964 , n22965 , n22966 , n22967 , n22968 , n22969 , n22970 , n22971 , n22972 , n22973 , n22974 , n22975 , n22976 , n22977 , n22978 , n22979 , n22980 , n22981 , n22982 , n22983 , n22984 , n22985 , n22986 , n22987 , n22988 , n22989 , n22990 , n22991 , n22992 , n22993 , n22994 , n22995 , n22996 , n22997 , n22998 , n22999 , n23000 , n23001 , n23002 , n23003 , n23004 , n23005 , n23006 , n23007 , n23008 , n23009 , n23010 , n23011 , n23012 , n23013 , n23014 , n23015 , n23016 , n23017 , n23018 , n23019 , n23020 , n23021 , n23022 , n23023 , n23024 , n23025 , n23026 , n23027 , n23028 , n23029 , n23030 , n23031 , n23032 , n23033 , n23034 , n23035 , n23036 , n23037 , n23038 , n23039 , n23040 , n23041 , n23042 , n23043 , n23044 , n23045 , n23046 , n23047 , n23048 , n23049 , n23050 , n23051 , n23052 , n23053 , n23054 , n23055 , n23056 , n23057 , n23058 , n23059 , n23060 , n23061 , n23062 , n23063 , n23064 , n23065 , n23066 , n23067 , n23068 , n23069 , n23070 , n23071 , n23072 , n23073 , n23074 , n23075 , n23076 , n23077 , n23078 , n23079 , n23080 , n23081 , n23082 , n23083 , n23084 , n23085 , n23086 , n23087 , n23088 , n23089 , n23090 , n23091 , n23092 , n23093 , n23094 , n23095 , n23096 , n23097 , n23098 , n23099 , n23100 , n23101 , n23102 , n23103 , n23104 , n23105 , n23106 , n23107 , n23108 , n23109 , n23110 , n23111 , n23112 , n23113 , n23114 , n23115 , n23116 , n23117 , n23118 , n23119 , n23120 , n23121 , n23122 , n23123 , n23124 , n23125 , n23126 , n23127 , n23128 , n23129 , n23130 , n23131 , n23132 , n23133 , n23134 , n23135 , n23136 , n23137 , n23138 , n23139 , n23140 , n23141 , n23142 , n23143 , n23144 , n23145 , n23146 , n23147 , n23148 , n23149 , n23150 , n23151 , n23152 , n23153 , n23154 , n23155 , n23156 , n23157 , n23158 , n23159 , n23160 , n23161 , n23162 , n23163 , n23164 , n23165 , n23166 , n23167 , n23168 , n23169 , n23170 , n23171 , n23172 , n23173 , n23174 , n23175 , n23176 , n23177 , n23178 , n23179 , n23180 , n23181 , n23182 , n23183 , n23184 , n23185 , n23186 , n23187 , n23188 , n23189 , n23190 , n23191 , n23192 , n23193 , n23194 , n23195 , n23196 , n23197 , n23198 , n23199 , n23200 , n23201 , n23202 , n23203 , n23204 , n23205 , n23206 , n23207 , n23208 , n23209 , n23210 , n23211 , n23212 , n23213 , n23214 , n23215 , n23216 , n23217 , n23218 , n23219 , n23220 , n23221 , n23222 , n23223 , n23224 , n23225 , n23226 , n23227 , n23228 , n23229 , n23230 , n23231 , n23232 , n23233 , n23234 , n23235 , n23236 , n23237 , n23238 , n23239 , n23240 , n23241 , n23242 , n23243 , n23244 , n23245 , n23246 , n23247 , n23248 , n23249 , n23250 , n23251 , n23252 , n23253 , n23254 , n23255 , n23256 , n23257 , n23258 , n23259 , n23260 , n23261 , n23262 , n23263 , n23264 , n23265 , n23266 , n23267 , n23268 , n23269 , n23270 , n23271 , n23272 , n23273 , n23274 , n23275 , n23276 , n23277 , n23278 , n23279 , n23280 , n23281 , n23282 , n23283 , n23284 , n23285 , n23286 , n23287 , n23288 , n23289 , n23290 , n23291 , n23292 , n23293 , n23294 , n23295 , n23296 , n23297 , n23298 , n23299 , n23300 , n23301 , n23302 , n23303 , n23304 , n23305 , n23306 , n23307 , n23308 , n23309 , n23310 , n23311 , n23312 , n23313 , n23314 , n23315 , n23316 , n23317 , n23318 , n23319 , n23320 , n23321 , n23322 , n23323 , n23324 , n23325 , n23326 , n23327 , n23328 , n23329 , n23330 , n23331 , n23332 , n23333 , n23334 , n23335 , n23336 , n23337 , n23338 , n23339 , n23340 , n23341 , n23342 , n23343 , n23344 , n23345 , n23346 , n23347 , n23348 , n23349 , n23350 , n23351 , n23352 , n23353 , n23354 , n23355 , n23356 , n23357 , n23358 , n23359 , n23360 , n23361 , n23362 , n23363 , n23364 , n23365 , n23366 , n23367 , n23368 , n23369 , n23370 , n23371 , n23372 , n23373 , n23374 , n23375 , n23376 , n23377 , n23378 , n23379 , n23380 , n23381 , n23382 , n23383 , n23384 , n23385 , n23386 , n23387 , n23388 , n23389 , n23390 , n23391 , n23392 , n23393 , n23394 , n23395 , n23396 , n23397 , n23398 , n23399 , n23400 , n23401 , n23402 , n23403 , n23404 , n23405 , n23406 , n23407 , n23408 , n23409 , n23410 , n23411 , n23412 , n23413 , n23414 , n23415 , n23416 , n23417 , n23418 , n23419 , n23420 , n23421 , n23422 , n23423 , n23424 , n23425 , n23426 , n23427 , n23428 , n23429 , n23430 , n23431 , n23432 , n23433 , n23434 , n23435 , n23436 , n23437 , n23438 , n23439 , n23440 , n23441 , n23442 , n23443 , n23444 , n23445 , n23446 , n23447 , n23448 , n23449 , n23450 , n23451 , n23452 , n23453 , n23454 , n23455 , n23456 , n23457 , n23458 , n23459 , n23460 , n23461 , n23462 , n23463 , n23464 , n23465 , n23466 , n23467 , n23468 , n23469 , n23470 , n23471 , n23472 , n23473 , n23474 , n23475 , n23476 , n23477 , n23478 , n23479 , n23480 , n23481 , n23482 , n23483 , n23484 , n23485 , n23486 , n23487 , n23488 , n23489 , n23490 , n23491 , n23492 , n23493 , n23494 , n23495 , n23496 , n23497 , n23498 , n23499 , n23500 , n23501 , n23502 , n23503 , n23504 , n23505 , n23506 , n23507 , n23508 , n23509 , n23510 , n23511 , n23512 , n23513 , n23514 , n23515 , n23516 , n23517 , n23518 , n23519 , n23520 , n23521 , n23522 , n23523 , n23524 , n23525 , n23526 , n23527 , n23528 , n23529 , n23530 , n23531 , n23532 , n23533 , n23534 , n23535 , n23536 , n23537 , n23538 , n23539 , n23540 , n23541 , n23542 , n23543 , n23544 , n23545 , n23546 , n23547 , n23548 , n23549 , n23550 , n23551 , n23552 , n23553 , n23554 , n23555 , n23556 , n23557 , n23558 , n23559 , n23560 , n23561 , n23562 , n23563 , n23564 , n23565 , n23566 , n23567 , n23568 , n23569 , n23570 , n23571 , n23572 , n23573 , n23574 , n23575 , n23576 , n23577 , n23578 , n23579 , n23580 , n23581 , n23582 , n23583 , n23584 , n23585 , n23586 , n23587 , n23588 , n23589 , n23590 , n23591 , n23592 , n23593 , n23594 , n23595 , n23596 , n23597 , n23598 , n23599 , n23600 , n23601 , n23602 , n23603 , n23604 , n23605 , n23606 , n23607 , n23608 , n23609 , n23610 , n23611 , n23612 , n23613 , n23614 , n23615 , n23616 , n23617 , n23618 , n23619 , n23620 , n23621 , n23622 , n23623 , n23624 , n23625 , n23626 , n23627 , n23628 , n23629 , n23630 , n23631 , n23632 , n23633 , n23634 , n23635 , n23636 , n23637 , n23638 , n23639 , n23640 , n23641 , n23642 , n23643 , n23644 , n23645 , n23646 , n23647 , n23648 , n23649 , n23650 , n23651 , n23652 , n23653 , n23654 , n23655 , n23656 , n23657 , n23658 , n23659 , n23660 , n23661 , n23662 , n23663 , n23664 , n23665 , n23666 , n23667 , n23668 , n23669 , n23670 , n23671 , n23672 , n23673 , n23674 , n23675 , n23676 , n23677 , n23678 , n23679 , n23680 , n23681 , n23682 , n23683 , n23684 , n23685 , n23686 , n23687 , n23688 , n23689 , n23690 , n23691 , n23692 , n23693 , n23694 , n23695 , n23696 , n23697 , n23698 , n23699 , n23700 , n23701 , n23702 , n23703 , n23704 , n23705 , n23706 , n23707 , n23708 , n23709 , n23710 , n23711 , n23712 , n23713 , n23714 , n23715 , n23716 , n23717 , n23718 , n23719 , n23720 , n23721 , n23722 , n23723 , n23724 , n23725 , n23726 , n23727 , n23728 , n23729 , n23730 , n23731 , n23732 , n23733 , n23734 , n23735 , n23736 , n23737 , n23738 , n23739 , n23740 , n23741 , n23742 , n23743 , n23744 , n23745 , n23746 , n23747 , n23748 , n23749 , n23750 , n23751 , n23752 , n23753 , n23754 , n23755 , n23756 , n23757 , n23758 , n23759 , n23760 , n23761 , n23762 , n23763 , n23764 , n23765 , n23766 , n23767 , n23768 , n23769 , n23770 , n23771 , n23772 , n23773 , n23774 , n23775 , n23776 , n23777 , n23778 , n23779 , n23780 , n23781 , n23782 , n23783 , n23784 , n23785 , n23786 , n23787 , n23788 , n23789 , n23790 , n23791 , n23792 , n23793 , n23794 , n23795 , n23796 , n23797 , n23798 , n23799 , n23800 , n23801 , n23802 , n23803 , n23804 , n23805 , n23806 , n23807 , n23808 , n23809 , n23810 , n23811 , n23812 , n23813 , n23814 , n23815 , n23816 , n23817 , n23818 , n23819 , n23820 , n23821 , n23822 , n23823 , n23824 , n23825 , n23826 , n23827 , n23828 , n23829 , n23830 , n23831 , n23832 , n23833 , n23834 , n23835 , n23836 , n23837 , n23838 , n23839 , n23840 , n23841 , n23842 , n23843 , n23844 , n23845 , n23846 , n23847 , n23848 , n23849 , n23850 , n23851 , n23852 , n23853 , n23854 , n23855 , n23856 , n23857 , n23858 , n23859 , n23860 , n23861 , n23862 , n23863 , n23864 , n23865 , n23866 , n23867 , n23868 , n23869 , n23870 , n23871 , n23872 , n23873 , n23874 , n23875 , n23876 , n23877 , n23878 , n23879 , n23880 , n23881 , n23882 , n23883 , n23884 , n23885 , n23886 , n23887 , n23888 , n23889 , n23890 , n23891 , n23892 , n23893 , n23894 , n23895 , n23896 , n23897 , n23898 , n23899 , n23900 , n23901 , n23902 , n23903 , n23904 , n23905 , n23906 , n23907 , n23908 , n23909 , n23910 , n23911 , n23912 , n23913 , n23914 , n23915 , n23916 , n23917 , n23918 , n23919 , n23920 , n23921 , n23922 , n23923 , n23924 , n23925 , n23926 , n23927 , n23928 , n23929 , n23930 , n23931 , n23932 , n23933 , n23934 , n23935 , n23936 , n23937 , n23938 , n23939 , n23940 , n23941 , n23942 , n23943 , n23944 , n23945 , n23946 , n23947 , n23948 , n23949 , n23950 , n23951 , n23952 , n23953 , n23954 , n23955 , n23956 , n23957 , n23958 , n23959 , n23960 , n23961 , n23962 , n23963 , n23964 , n23965 , n23966 , n23967 , n23968 , n23969 , n23970 , n23971 , n23972 , n23973 , n23974 , n23975 , n23976 , n23977 , n23978 , n23979 , n23980 , n23981 , n23982 , n23983 , n23984 , n23985 , n23986 , n23987 , n23988 , n23989 , n23990 , n23991 , n23992 , n23993 , n23994 , n23995 , n23996 , n23997 , n23998 , n23999 , n24000 , n24001 , n24002 , n24003 , n24004 , n24005 , n24006 , n24007 , n24008 , n24009 , n24010 , n24011 , n24012 , n24013 , n24014 , n24015 , n24016 , n24017 , n24018 , n24019 , n24020 , n24021 , n24022 , n24023 , n24024 , n24025 , n24026 , n24027 , n24028 , n24029 , n24030 , n24031 , n24032 , n24033 , n24034 , n24035 , n24036 , n24037 , n24038 , n24039 , n24040 , n24041 , n24042 , n24043 , n24044 , n24045 , n24046 , n24047 , n24048 , n24049 , n24050 , n24051 , n24052 , n24053 , n24054 , n24055 , n24056 , n24057 , n24058 , n24059 , n24060 , n24061 , n24062 , n24063 , n24064 , n24065 , n24066 , n24067 , n24068 , n24069 , n24070 , n24071 , n24072 , n24073 , n24074 , n24075 , n24076 , n24077 , n24078 , n24079 , n24080 , n24081 , n24082 , n24083 , n24084 , n24085 , n24086 , n24087 , n24088 , n24089 , n24090 , n24091 , n24092 , n24093 , n24094 , n24095 , n24096 , n24097 , n24098 , n24099 , n24100 , n24101 , n24102 , n24103 , n24104 , n24105 , n24106 , n24107 , n24108 , n24109 , n24110 , n24111 , n24112 , n24113 , n24114 , n24115 , n24116 , n24117 , n24118 , n24119 , n24120 , n24121 , n24122 , n24123 , n24124 , n24125 , n24126 , n24127 , n24128 , n24129 , n24130 , n24131 , n24132 , n24133 , n24134 , n24135 , n24136 , n24137 , n24138 , n24139 , n24140 , n24141 , n24142 , n24143 , n24144 , n24145 , n24146 , n24147 , n24148 , n24149 , n24150 , n24151 , n24152 , n24153 , n24154 , n24155 , n24156 , n24157 , n24158 , n24159 , n24160 , n24161 , n24162 , n24163 , n24164 , n24165 , n24166 , n24167 , n24168 , n24169 , n24170 , n24171 , n24172 , n24173 , n24174 , n24175 , n24176 , n24177 , n24178 , n24179 , n24180 , n24181 , n24182 , n24183 , n24184 , n24185 , n24186 , n24187 , n24188 , n24189 , n24190 , n24191 , n24192 , n24193 , n24194 , n24195 , n24196 , n24197 , n24198 , n24199 , n24200 , n24201 , n24202 , n24203 , n24204 , n24205 , n24206 , n24207 , n24208 , n24209 , n24210 , n24211 , n24212 , n24213 , n24214 , n24215 , n24216 , n24217 , n24218 , n24219 , n24220 , n24221 , n24222 , n24223 , n24224 , n24225 , n24226 , n24227 , n24228 , n24229 , n24230 , n24231 , n24232 , n24233 , n24234 , n24235 , n24236 , n24237 , n24238 , n24239 , n24240 , n24241 , n24242 , n24243 , n24244 , n24245 , n24246 , n24247 , n24248 , n24249 , n24250 , n24251 , n24252 , n24253 , n24254 , n24255 , n24256 , n24257 , n24258 , n24259 , n24260 , n24261 , n24262 , n24263 , n24264 , n24265 , n24266 , n24267 , n24268 , n24269 , n24270 , n24271 , n24272 , n24273 , n24274 , n24275 , n24276 , n24277 , n24278 , n24279 , n24280 , n24281 , n24282 , n24283 , n24284 , n24285 , n24286 , n24287 , n24288 , n24289 , n24290 , n24291 , n24292 , n24293 , n24294 , n24295 , n24296 , n24297 , n24298 , n24299 , n24300 , n24301 , n24302 , n24303 , n24304 , n24305 , n24306 , n24307 , n24308 , n24309 , n24310 , n24311 , n24312 , n24313 , n24314 , n24315 , n24316 , n24317 , n24318 , n24319 , n24320 , n24321 , n24322 , n24323 , n24324 , n24325 , n24326 , n24327 , n24328 , n24329 , n24330 , n24331 , n24332 , n24333 , n24334 , n24335 , n24336 , n24337 , n24338 , n24339 , n24340 , n24341 , n24342 , n24343 , n24344 , n24345 , n24346 , n24347 , n24348 , n24349 , n24350 , n24351 , n24352 , n24353 , n24354 , n24355 , n24356 , n24357 , n24358 , n24359 , n24360 , n24361 , n24362 , n24363 , n24364 , n24365 , n24366 , n24367 , n24368 , n24369 , n24370 , n24371 , n24372 , n24373 , n24374 , n24375 , n24376 , n24377 , n24378 , n24379 , n24380 , n24381 , n24382 , n24383 , n24384 , n24385 , n24386 , n24387 , n24388 , n24389 , n24390 , n24391 , n24392 , n24393 , n24394 , n24395 , n24396 , n24397 , n24398 , n24399 , n24400 , n24401 , n24402 , n24403 , n24404 , n24405 , n24406 , n24407 , n24408 , n24409 , n24410 , n24411 , n24412 , n24413 , n24414 , n24415 , n24416 , n24417 , n24418 , n24419 , n24420 , n24421 , n24422 , n24423 , n24424 , n24425 , n24426 , n24427 , n24428 , n24429 , n24430 , n24431 , n24432 , n24433 , n24434 , n24435 , n24436 , n24437 , n24438 , n24439 , n24440 , n24441 , n24442 , n24443 , n24444 , n24445 , n24446 , n24447 , n24448 , n24449 , n24450 , n24451 , n24452 , n24453 , n24454 , n24455 , n24456 , n24457 , n24458 , n24459 , n24460 , n24461 , n24462 , n24463 , n24464 , n24465 , n24466 , n24467 , n24468 , n24469 , n24470 , n24471 , n24472 , n24473 , n24474 , n24475 , n24476 , n24477 , n24478 , n24479 , n24480 , n24481 , n24482 , n24483 , n24484 , n24485 , n24486 , n24487 , n24488 , n24489 , n24490 , n24491 , n24492 , n24493 , n24494 , n24495 , n24496 , n24497 , n24498 , n24499 , n24500 , n24501 , n24502 , n24503 , n24504 , n24505 , n24506 , n24507 , n24508 , n24509 , n24510 , n24511 , n24512 , n24513 , n24514 , n24515 , n24516 , n24517 , n24518 , n24519 , n24520 , n24521 , n24522 , n24523 , n24524 , n24525 , n24526 , n24527 , n24528 , n24529 , n24530 , n24531 , n24532 , n24533 , n24534 , n24535 , n24536 , n24537 , n24538 , n24539 , n24540 , n24541 , n24542 , n24543 , n24544 , n24545 , n24546 , n24547 , n24548 , n24549 , n24550 , n24551 , n24552 , n24553 , n24554 , n24555 , n24556 , n24557 , n24558 , n24559 , n24560 , n24561 , n24562 , n24563 , n24564 , n24565 , n24566 , n24567 , n24568 , n24569 , n24570 , n24571 , n24572 , n24573 , n24574 , n24575 , n24576 , n24577 , n24578 , n24579 , n24580 , n24581 , n24582 , n24583 , n24584 , n24585 , n24586 , n24587 , n24588 , n24589 , n24590 , n24591 , n24592 , n24593 , n24594 , n24595 , n24596 , n24597 , n24598 , n24599 , n24600 , n24601 , n24602 , n24603 , n24604 , n24605 , n24606 , n24607 , n24608 , n24609 , n24610 , n24611 , n24612 , n24613 , n24614 , n24615 , n24616 , n24617 , n24618 , n24619 , n24620 , n24621 , n24622 , n24623 , n24624 , n24625 , n24626 , n24627 , n24628 , n24629 , n24630 , n24631 , n24632 , n24633 , n24634 , n24635 , n24636 , n24637 , n24638 , n24639 , n24640 , n24641 , n24642 , n24643 , n24644 , n24645 , n24646 , n24647 , n24648 , n24649 , n24650 , n24651 , n24652 , n24653 , n24654 , n24655 , n24656 , n24657 , n24658 , n24659 , n24660 , n24661 , n24662 , n24663 , n24664 , n24665 , n24666 , n24667 , n24668 , n24669 , n24670 , n24671 , n24672 , n24673 , n24674 , n24675 , n24676 , n24677 , n24678 , n24679 , n24680 , n24681 , n24682 , n24683 , n24684 , n24685 , n24686 , n24687 , n24688 , n24689 , n24690 , n24691 , n24692 , n24693 , n24694 , n24695 , n24696 , n24697 , n24698 , n24699 , n24700 , n24701 , n24702 , n24703 , n24704 , n24705 , n24706 , n24707 , n24708 , n24709 , n24710 , n24711 , n24712 , n24713 , n24714 , n24715 , n24716 , n24717 , n24718 , n24719 , n24720 , n24721 , n24722 , n24723 , n24724 , n24725 , n24726 , n24727 , n24728 , n24729 , n24730 , n24731 , n24732 , n24733 , n24734 , n24735 , n24736 , n24737 , n24738 , n24739 , n24740 , n24741 , n24742 , n24743 , n24744 , n24745 , n24746 , n24747 , n24748 , n24749 , n24750 , n24751 , n24752 , n24753 , n24754 , n24755 , n24756 , n24757 , n24758 , n24759 , n24760 , n24761 , n24762 , n24763 , n24764 , n24765 , n24766 , n24767 , n24768 , n24769 , n24770 , n24771 , n24772 , n24773 , n24774 , n24775 , n24776 , n24777 , n24778 , n24779 , n24780 , n24781 , n24782 , n24783 , n24784 , n24785 , n24786 , n24787 , n24788 , n24789 , n24790 , n24791 , n24792 , n24793 , n24794 , n24795 , n24796 , n24797 , n24798 , n24799 , n24800 , n24801 , n24802 , n24803 , n24804 , n24805 , n24806 , n24807 , n24808 , n24809 , n24810 , n24811 , n24812 , n24813 , n24814 , n24815 , n24816 , n24817 , n24818 , n24819 , n24820 , n24821 , n24822 , n24823 , n24824 , n24825 , n24826 , n24827 , n24828 , n24829 , n24830 , n24831 , n24832 , n24833 , n24834 , n24835 , n24836 , n24837 , n24838 , n24839 , n24840 , n24841 , n24842 , n24843 , n24844 , n24845 , n24846 , n24847 , n24848 , n24849 , n24850 , n24851 , n24852 , n24853 , n24854 , n24855 , n24856 , n24857 , n24858 , n24859 , n24860 , n24861 , n24862 , n24863 , n24864 , n24865 , n24866 , n24867 , n24868 , n24869 , n24870 , n24871 , n24872 , n24873 , n24874 , n24875 , n24876 , n24877 , n24878 , n24879 , n24880 , n24881 , n24882 , n24883 , n24884 , n24885 , n24886 , n24887 , n24888 , n24889 , n24890 , n24891 , n24892 , n24893 , n24894 , n24895 , n24896 , n24897 , n24898 , n24899 , n24900 , n24901 , n24902 , n24903 , n24904 , n24905 , n24906 , n24907 , n24908 , n24909 , n24910 , n24911 , n24912 , n24913 , n24914 , n24915 , n24916 , n24917 , n24918 , n24919 , n24920 , n24921 , n24922 , n24923 , n24924 , n24925 , n24926 , n24927 , n24928 , n24929 , n24930 , n24931 , n24932 , n24933 , n24934 , n24935 , n24936 , n24937 , n24938 , n24939 , n24940 , n24941 , n24942 , n24943 , n24944 , n24945 , n24946 , n24947 , n24948 , n24949 , n24950 , n24951 , n24952 , n24953 , n24954 , n24955 , n24956 , n24957 , n24958 , n24959 , n24960 , n24961 , n24962 , n24963 , n24964 , n24965 , n24966 , n24967 , n24968 , n24969 , n24970 , n24971 , n24972 , n24973 , n24974 , n24975 , n24976 , n24977 , n24978 , n24979 , n24980 , n24981 , n24982 , n24983 , n24984 , n24985 , n24986 , n24987 , n24988 , n24989 , n24990 , n24991 , n24992 , n24993 , n24994 , n24995 , n24996 , n24997 , n24998 , n24999 , n25000 , n25001 , n25002 , n25003 , n25004 , n25005 , n25006 , n25007 , n25008 , n25009 , n25010 , n25011 , n25012 , n25013 , n25014 , n25015 , n25016 , n25017 , n25018 , n25019 , n25020 , n25021 , n25022 , n25023 , n25024 , n25025 , n25026 , n25027 , n25028 , n25029 , n25030 , n25031 , n25032 , n25033 , n25034 , n25035 , n25036 , n25037 , n25038 , n25039 , n25040 , n25041 , n25042 , n25043 , n25044 , n25045 , n25046 , n25047 , n25048 , n25049 , n25050 , n25051 , n25052 , n25053 , n25054 , n25055 , n25056 , n25057 , n25058 , n25059 , n25060 , n25061 , n25062 , n25063 , n25064 , n25065 , n25066 , n25067 , n25068 , n25069 , n25070 , n25071 , n25072 , n25073 , n25074 , n25075 , n25076 , n25077 , n25078 , n25079 , n25080 , n25081 , n25082 , n25083 , n25084 , n25085 , n25086 , n25087 , n25088 , n25089 , n25090 , n25091 , n25092 , n25093 , n25094 , n25095 , n25096 , n25097 , n25098 , n25099 , n25100 , n25101 , n25102 , n25103 , n25104 , n25105 , n25106 , n25107 , n25108 , n25109 , n25110 , n25111 , n25112 , n25113 , n25114 , n25115 , n25116 , n25117 , n25118 , n25119 , n25120 , n25121 , n25122 , n25123 , n25124 , n25125 , n25126 , n25127 , n25128 , n25129 , n25130 , n25131 , n25132 , n25133 , n25134 , n25135 , n25136 , n25137 , n25138 , n25139 , n25140 , n25141 , n25142 , n25143 , n25144 , n25145 , n25146 , n25147 , n25148 , n25149 , n25150 , n25151 , n25152 , n25153 , n25154 , n25155 , n25156 , n25157 , n25158 , n25159 , n25160 , n25161 , n25162 , n25163 , n25164 , n25165 , n25166 , n25167 , n25168 , n25169 , n25170 , n25171 , n25172 , n25173 , n25174 , n25175 , n25176 , n25177 , n25178 , n25179 , n25180 , n25181 , n25182 , n25183 , n25184 , n25185 , n25186 , n25187 , n25188 , n25189 , n25190 , n25191 , n25192 , n25193 , n25194 , n25195 , n25196 , n25197 , n25198 , n25199 , n25200 , n25201 , n25202 , n25203 , n25204 , n25205 , n25206 , n25207 , n25208 , n25209 , n25210 , n25211 , n25212 , n25213 , n25214 , n25215 , n25216 , n25217 , n25218 , n25219 , n25220 , n25221 , n25222 , n25223 , n25224 , n25225 , n25226 , n25227 , n25228 , n25229 , n25230 , n25231 , n25232 , n25233 , n25234 , n25235 , n25236 , n25237 , n25238 , n25239 , n25240 , n25241 , n25242 , n25243 , n25244 , n25245 , n25246 , n25247 , n25248 , n25249 , n25250 , n25251 , n25252 , n25253 , n25254 , n25255 , n25256 , n25257 , n25258 , n25259 , n25260 , n25261 , n25262 , n25263 , n25264 , n25265 , n25266 , n25267 , n25268 , n25269 , n25270 , n25271 , n25272 , n25273 , n25274 , n25275 , n25276 , n25277 , n25278 , n25279 , n25280 , n25281 , n25282 , n25283 , n25284 , n25285 , n25286 , n25287 , n25288 , n25289 , n25290 , n25291 , n25292 , n25293 , n25294 , n25295 , n25296 , n25297 , n25298 , n25299 , n25300 , n25301 , n25302 , n25303 , n25304 , n25305 , n25306 , n25307 , n25308 , n25309 , n25310 , n25311 , n25312 , n25313 , n25314 , n25315 , n25316 , n25317 , n25318 , n25319 , n25320 , n25321 , n25322 , n25323 , n25324 , n25325 , n25326 , n25327 , n25328 , n25329 , n25330 , n25331 , n25332 , n25333 , n25334 , n25335 , n25336 , n25337 , n25338 , n25339 , n25340 , n25341 , n25342 , n25343 , n25344 , n25345 , n25346 , n25347 , n25348 , n25349 , n25350 , n25351 , n25352 , n25353 , n25354 , n25355 , n25356 , n25357 , n25358 , n25359 , n25360 , n25361 , n25362 , n25363 , n25364 , n25365 , n25366 , n25367 , n25368 , n25369 , n25370 , n25371 , n25372 , n25373 , n25374 , n25375 , n25376 , n25377 , n25378 , n25379 , n25380 , n25381 , n25382 , n25383 , n25384 , n25385 , n25386 , n25387 , n25388 , n25389 , n25390 , n25391 , n25392 , n25393 , n25394 , n25395 , n25396 , n25397 , n25398 , n25399 , n25400 , n25401 , n25402 , n25403 , n25404 , n25405 , n25406 , n25407 , n25408 , n25409 , n25410 , n25411 , n25412 , n25413 , n25414 , n25415 , n25416 , n25417 , n25418 , n25419 , n25420 , n25421 , n25422 , n25423 , n25424 , n25425 , n25426 , n25427 , n25428 , n25429 , n25430 , n25431 , n25432 , n25433 , n25434 , n25435 , n25436 , n25437 , n25438 , n25439 , n25440 , n25441 , n25442 , n25443 , n25444 , n25445 , n25446 , n25447 , n25448 , n25449 , n25450 , n25451 , n25452 , n25453 , n25454 , n25455 , n25456 , n25457 , n25458 , n25459 , n25460 , n25461 , n25462 , n25463 , n25464 , n25465 , n25466 , n25467 , n25468 , n25469 , n25470 , n25471 , n25472 , n25473 , n25474 , n25475 , n25476 , n25477 , n25478 , n25479 , n25480 , n25481 , n25482 , n25483 , n25484 , n25485 , n25486 , n25487 , n25488 , n25489 , n25490 , n25491 , n25492 , n25493 , n25494 , n25495 , n25496 , n25497 , n25498 , n25499 , n25500 , n25501 , n25502 , n25503 , n25504 , n25505 , n25506 , n25507 , n25508 , n25509 , n25510 , n25511 , n25512 , n25513 , n25514 , n25515 , n25516 , n25517 , n25518 , n25519 , n25520 , n25521 , n25522 , n25523 , n25524 , n25525 , n25526 , n25527 , n25528 , n25529 , n25530 , n25531 , n25532 , n25533 , n25534 , n25535 , n25536 , n25537 , n25538 , n25539 , n25540 , n25541 , n25542 , n25543 , n25544 , n25545 , n25546 , n25547 , n25548 , n25549 , n25550 , n25551 , n25552 , n25553 , n25554 , n25555 , n25556 , n25557 , n25558 , n25559 , n25560 , n25561 , n25562 , n25563 , n25564 , n25565 , n25566 , n25567 , n25568 , n25569 , n25570 , n25571 , n25572 , n25573 , n25574 , n25575 , n25576 , n25577 , n25578 , n25579 , n25580 , n25581 , n25582 , n25583 , n25584 , n25585 , n25586 , n25587 , n25588 , n25589 , n25590 , n25591 , n25592 , n25593 , n25594 , n25595 , n25596 , n25597 , n25598 , n25599 , n25600 , n25601 , n25602 , n25603 , n25604 , n25605 , n25606 , n25607 , n25608 , n25609 , n25610 , n25611 , n25612 , n25613 , n25614 , n25615 , n25616 , n25617 , n25618 , n25619 , n25620 , n25621 , n25622 , n25623 , n25624 , n25625 , n25626 , n25627 , n25628 , n25629 , n25630 , n25631 , n25632 , n25633 , n25634 , n25635 , n25636 , n25637 , n25638 , n25639 , n25640 , n25641 , n25642 , n25643 , n25644 , n25645 , n25646 , n25647 , n25648 , n25649 , n25650 , n25651 , n25652 , n25653 , n25654 , n25655 , n25656 , n25657 , n25658 , n25659 , n25660 , n25661 , n25662 , n25663 , n25664 , n25665 , n25666 , n25667 , n25668 , n25669 , n25670 , n25671 , n25672 , n25673 , n25674 , n25675 , n25676 , n25677 , n25678 , n25679 , n25680 , n25681 , n25682 , n25683 , n25684 , n25685 , n25686 , n25687 , n25688 , n25689 , n25690 , n25691 , n25692 , n25693 , n25694 , n25695 , n25696 , n25697 , n25698 , n25699 , n25700 , n25701 , n25702 , n25703 , n25704 , n25705 , n25706 , n25707 , n25708 , n25709 , n25710 , n25711 , n25712 , n25713 , n25714 , n25715 , n25716 , n25717 , n25718 , n25719 , n25720 , n25721 , n25722 , n25723 , n25724 , n25725 , n25726 , n25727 , n25728 , n25729 , n25730 , n25731 , n25732 , n25733 , n25734 , n25735 , n25736 , n25737 , n25738 , n25739 , n25740 , n25741 , n25742 , n25743 , n25744 , n25745 , n25746 , n25747 , n25748 , n25749 , n25750 , n25751 , n25752 , n25753 , n25754 , n25755 , n25756 , n25757 , n25758 , n25759 , n25760 , n25761 , n25762 , n25763 , n25764 , n25765 , n25766 , n25767 , n25768 , n25769 , n25770 , n25771 , n25772 , n25773 , n25774 , n25775 , n25776 , n25777 , n25778 , n25779 , n25780 , n25781 , n25782 , n25783 , n25784 , n25785 , n25786 , n25787 , n25788 , n25789 , n25790 , n25791 , n25792 , n25793 , n25794 , n25795 , n25796 , n25797 , n25798 , n25799 , n25800 , n25801 , n25802 , n25803 , n25804 , n25805 , n25806 , n25807 , n25808 , n25809 , n25810 , n25811 , n25812 , n25813 , n25814 , n25815 , n25816 , n25817 , n25818 , n25819 , n25820 , n25821 , n25822 , n25823 , n25824 , n25825 , n25826 , n25827 , n25828 , n25829 , n25830 , n25831 , n25832 , n25833 , n25834 , n25835 , n25836 , n25837 , n25838 , n25839 , n25840 , n25841 , n25842 , n25843 , n25844 , n25845 , n25846 , n25847 , n25848 , n25849 , n25850 , n25851 , n25852 , n25853 , n25854 , n25855 , n25856 , n25857 , n25858 , n25859 , n25860 , n25861 , n25862 , n25863 , n25864 , n25865 , n25866 , n25867 , n25868 , n25869 , n25870 , n25871 , n25872 , n25873 , n25874 , n25875 , n25876 , n25877 , n25878 , n25879 , n25880 , n25881 , n25882 , n25883 , n25884 , n25885 , n25886 , n25887 , n25888 , n25889 , n25890 , n25891 , n25892 , n25893 , n25894 , n25895 , n25896 , n25897 , n25898 , n25899 , n25900 , n25901 , n25902 , n25903 , n25904 , n25905 , n25906 , n25907 , n25908 , n25909 , n25910 , n25911 , n25912 , n25913 , n25914 , n25915 , n25916 , n25917 , n25918 , n25919 , n25920 , n25921 , n25922 , n25923 , n25924 , n25925 , n25926 , n25927 , n25928 , n25929 , n25930 , n25931 , n25932 , n25933 , n25934 , n25935 , n25936 , n25937 , n25938 , n25939 , n25940 , n25941 , n25942 , n25943 , n25944 , n25945 , n25946 , n25947 , n25948 , n25949 , n25950 , n25951 , n25952 , n25953 , n25954 , n25955 , n25956 , n25957 , n25958 , n25959 , n25960 , n25961 , n25962 , n25963 , n25964 , n25965 , n25966 , n25967 , n25968 , n25969 , n25970 , n25971 , n25972 , n25973 , n25974 , n25975 , n25976 , n25977 , n25978 , n25979 , n25980 , n25981 , n25982 , n25983 , n25984 , n25985 , n25986 , n25987 , n25988 , n25989 , n25990 , n25991 , n25992 , n25993 , n25994 , n25995 , n25996 , n25997 , n25998 , n25999 , n26000 , n26001 , n26002 , n26003 , n26004 , n26005 , n26006 , n26007 , n26008 , n26009 , n26010 , n26011 , n26012 , n26013 , n26014 , n26015 , n26016 , n26017 , n26018 , n26019 , n26020 , n26021 , n26022 , n26023 , n26024 , n26025 , n26026 , n26027 , n26028 , n26029 , n26030 , n26031 , n26032 , n26033 , n26034 , n26035 , n26036 , n26037 , n26038 , n26039 , n26040 , n26041 , n26042 , n26043 , n26044 , n26045 , n26046 , n26047 , n26048 , n26049 , n26050 , n26051 , n26052 , n26053 , n26054 , n26055 , n26056 , n26057 , n26058 , n26059 , n26060 , n26061 , n26062 , n26063 , n26064 , n26065 , n26066 , n26067 , n26068 , n26069 , n26070 , n26071 , n26072 , n26073 , n26074 , n26075 , n26076 , n26077 , n26078 , n26079 , n26080 , n26081 , n26082 , n26083 , n26084 , n26085 , n26086 , n26087 , n26088 , n26089 , n26090 , n26091 , n26092 , n26093 , n26094 , n26095 , n26096 , n26097 , n26098 , n26099 , n26100 , n26101 , n26102 , n26103 , n26104 , n26105 , n26106 , n26107 , n26108 , n26109 , n26110 , n26111 , n26112 , n26113 , n26114 , n26115 , n26116 , n26117 , n26118 , n26119 , n26120 , n26121 , n26122 , n26123 , n26124 , n26125 , n26126 , n26127 , n26128 , n26129 , n26130 , n26131 , n26132 , n26133 , n26134 , n26135 , n26136 , n26137 , n26138 , n26139 , n26140 , n26141 , n26142 , n26143 , n26144 , n26145 , n26146 , n26147 , n26148 , n26149 , n26150 , n26151 , n26152 , n26153 , n26154 , n26155 , n26156 , n26157 , n26158 , n26159 , n26160 , n26161 , n26162 , n26163 , n26164 , n26165 , n26166 , n26167 , n26168 , n26169 , n26170 , n26171 , n26172 , n26173 , n26174 , n26175 , n26176 , n26177 , n26178 , n26179 , n26180 , n26181 , n26182 , n26183 , n26184 , n26185 , n26186 , n26187 , n26188 , n26189 , n26190 , n26191 , n26192 , n26193 , n26194 , n26195 , n26196 , n26197 , n26198 , n26199 , n26200 , n26201 , n26202 , n26203 , n26204 , n26205 , n26206 , n26207 , n26208 , n26209 , n26210 , n26211 , n26212 , n26213 , n26214 , n26215 , n26216 , n26217 , n26218 , n26219 , n26220 , n26221 , n26222 , n26223 , n26224 , n26225 , n26226 , n26227 , n26228 , n26229 , n26230 , n26231 , n26232 , n26233 , n26234 , n26235 , n26236 , n26237 , n26238 , n26239 , n26240 , n26241 , n26242 , n26243 , n26244 , n26245 , n26246 , n26247 , n26248 , n26249 , n26250 , n26251 , n26252 , n26253 , n26254 , n26255 , n26256 , n26257 , n26258 , n26259 , n26260 , n26261 , n26262 , n26263 , n26264 , n26265 , n26266 , n26267 , n26268 , n26269 , n26270 , n26271 , n26272 , n26273 , n26274 , n26275 , n26276 , n26277 , n26278 , n26279 , n26280 , n26281 , n26282 , n26283 , n26284 , n26285 , n26286 , n26287 , n26288 , n26289 , n26290 , n26291 , n26292 , n26293 , n26294 , n26295 , n26296 , n26297 , n26298 , n26299 , n26300 , n26301 , n26302 , n26303 , n26304 , n26305 , n26306 , n26307 , n26308 , n26309 , n26310 , n26311 , n26312 , n26313 , n26314 , n26315 , n26316 , n26317 , n26318 , n26319 , n26320 , n26321 , n26322 , n26323 , n26324 , n26325 , n26326 , n26327 , n26328 , n26329 , n26330 , n26331 , n26332 , n26333 , n26334 , n26335 , n26336 , n26337 , n26338 , n26339 , n26340 , n26341 , n26342 , n26343 , n26344 , n26345 , n26346 , n26347 , n26348 , n26349 , n26350 , n26351 , n26352 , n26353 , n26354 , n26355 , n26356 , n26357 , n26358 , n26359 , n26360 , n26361 , n26362 , n26363 , n26364 , n26365 , n26366 , n26367 , n26368 , n26369 , n26370 , n26371 , n26372 , n26373 , n26374 , n26375 , n26376 , n26377 , n26378 , n26379 , n26380 , n26381 , n26382 , n26383 , n26384 , n26385 , n26386 , n26387 , n26388 , n26389 , n26390 , n26391 , n26392 , n26393 , n26394 , n26395 , n26396 , n26397 , n26398 , n26399 , n26400 , n26401 , n26402 , n26403 , n26404 , n26405 , n26406 , n26407 , n26408 , n26409 , n26410 , n26411 , n26412 , n26413 , n26414 , n26415 , n26416 , n26417 , n26418 , n26419 , n26420 , n26421 , n26422 , n26423 , n26424 , n26425 , n26426 , n26427 , n26428 , n26429 , n26430 , n26431 , n26432 , n26433 , n26434 , n26435 , n26436 , n26437 , n26438 , n26439 , n26440 , n26441 , n26442 , n26443 , n26444 , n26445 , n26446 , n26447 , n26448 , n26449 , n26450 , n26451 , n26452 , n26453 , n26454 , n26455 , n26456 , n26457 , n26458 , n26459 , n26460 , n26461 , n26462 , n26463 , n26464 , n26465 , n26466 , n26467 , n26468 , n26469 , n26470 , n26471 , n26472 , n26473 , n26474 , n26475 , n26476 , n26477 , n26478 , n26479 , n26480 , n26481 , n26482 , n26483 , n26484 , n26485 , n26486 , n26487 , n26488 , n26489 , n26490 , n26491 , n26492 , n26493 , n26494 , n26495 , n26496 , n26497 , n26498 , n26499 , n26500 , n26501 , n26502 , n26503 , n26504 , n26505 , n26506 , n26507 , n26508 , n26509 , n26510 , n26511 , n26512 , n26513 , n26514 , n26515 , n26516 , n26517 , n26518 , n26519 , n26520 , n26521 , n26522 , n26523 , n26524 , n26525 , n26526 , n26527 , n26528 , n26529 , n26530 , n26531 , n26532 , n26533 , n26534 , n26535 , n26536 , n26537 , n26538 , n26539 , n26540 , n26541 , n26542 , n26543 , n26544 , n26545 , n26546 , n26547 , n26548 , n26549 , n26550 , n26551 , n26552 , n26553 , n26554 , n26555 , n26556 , n26557 , n26558 , n26559 , n26560 , n26561 , n26562 , n26563 , n26564 , n26565 , n26566 , n26567 , n26568 , n26569 , n26570 , n26571 , n26572 , n26573 , n26574 , n26575 , n26576 , n26577 , n26578 , n26579 , n26580 , n26581 , n26582 , n26583 , n26584 , n26585 , n26586 , n26587 , n26588 , n26589 , n26590 , n26591 , n26592 , n26593 , n26594 , n26595 , n26596 , n26597 , n26598 , n26599 , n26600 , n26601 , n26602 , n26603 , n26604 , n26605 , n26606 , n26607 , n26608 , n26609 , n26610 , n26611 , n26612 , n26613 , n26614 , n26615 , n26616 , n26617 , n26618 , n26619 , n26620 , n26621 , n26622 , n26623 , n26624 , n26625 , n26626 , n26627 , n26628 , n26629 , n26630 , n26631 , n26632 , n26633 , n26634 , n26635 , n26636 , n26637 , n26638 , n26639 , n26640 , n26641 , n26642 , n26643 , n26644 , n26645 , n26646 , n26647 , n26648 , n26649 , n26650 , n26651 , n26652 , n26653 , n26654 , n26655 , n26656 , n26657 , n26658 , n26659 , n26660 , n26661 , n26662 , n26663 , n26664 , n26665 , n26666 , n26667 , n26668 , n26669 , n26670 , n26671 , n26672 , n26673 , n26674 , n26675 , n26676 , n26677 , n26678 , n26679 , n26680 , n26681 , n26682 , n26683 , n26684 , n26685 , n26686 , n26687 , n26688 , n26689 , n26690 , n26691 , n26692 , n26693 , n26694 , n26695 , n26696 , n26697 , n26698 , n26699 , n26700 , n26701 , n26702 , n26703 , n26704 , n26705 , n26706 , n26707 , n26708 , n26709 , n26710 , n26711 , n26712 , n26713 , n26714 , n26715 , n26716 , n26717 , n26718 , n26719 , n26720 , n26721 , n26722 , n26723 , n26724 , n26725 , n26726 , n26727 , n26728 , n26729 , n26730 , n26731 , n26732 , n26733 , n26734 , n26735 , n26736 , n26737 , n26738 , n26739 , n26740 , n26741 , n26742 , n26743 , n26744 , n26745 , n26746 , n26747 , n26748 , n26749 , n26750 , n26751 , n26752 , n26753 , n26754 , n26755 , n26756 , n26757 , n26758 , n26759 , n26760 , n26761 , n26762 , n26763 , n26764 , n26765 , n26766 , n26767 , n26768 , n26769 , n26770 , n26771 , n26772 , n26773 , n26774 , n26775 , n26776 , n26777 , n26778 , n26779 , n26780 , n26781 , n26782 , n26783 , n26784 , n26785 , n26786 , n26787 , n26788 , n26789 , n26790 , n26791 , n26792 , n26793 , n26794 , n26795 , n26796 , n26797 , n26798 , n26799 , n26800 , n26801 , n26802 , n26803 , n26804 , n26805 , n26806 , n26807 , n26808 , n26809 , n26810 , n26811 , n26812 , n26813 , n26814 , n26815 , n26816 , n26817 , n26818 , n26819 , n26820 , n26821 , n26822 , n26823 , n26824 , n26825 , n26826 , n26827 , n26828 , n26829 , n26830 , n26831 , n26832 , n26833 , n26834 , n26835 , n26836 , n26837 , n26838 , n26839 , n26840 , n26841 , n26842 , n26843 , n26844 , n26845 , n26846 , n26847 , n26848 , n26849 , n26850 , n26851 , n26852 , n26853 , n26854 , n26855 , n26856 , n26857 , n26858 , n26859 , n26860 , n26861 , n26862 , n26863 , n26864 , n26865 , n26866 , n26867 , n26868 , n26869 , n26870 , n26871 , n26872 , n26873 , n26874 , n26875 , n26876 , n26877 , n26878 , n26879 , n26880 , n26881 , n26882 , n26883 , n26884 , n26885 , n26886 , n26887 , n26888 , n26889 , n26890 , n26891 , n26892 , n26893 , n26894 , n26895 , n26896 , n26897 , n26898 , n26899 , n26900 , n26901 , n26902 , n26903 , n26904 , n26905 , n26906 , n26907 , n26908 , n26909 , n26910 , n26911 , n26912 , n26913 , n26914 , n26915 , n26916 , n26917 , n26918 , n26919 , n26920 , n26921 , n26922 , n26923 , n26924 , n26925 , n26926 , n26927 , n26928 , n26929 , n26930 , n26931 , n26932 , n26933 , n26934 , n26935 , n26936 , n26937 , n26938 , n26939 , n26940 , n26941 , n26942 , n26943 , n26944 , n26945 , n26946 , n26947 , n26948 , n26949 , n26950 , n26951 , n26952 , n26953 , n26954 , n26955 , n26956 , n26957 , n26958 , n26959 , n26960 , n26961 , n26962 , n26963 , n26964 , n26965 , n26966 , n26967 , n26968 , n26969 , n26970 , n26971 , n26972 , n26973 , n26974 , n26975 , n26976 , n26977 , n26978 , n26979 , n26980 , n26981 , n26982 , n26983 , n26984 , n26985 , n26986 , n26987 , n26988 , n26989 , n26990 , n26991 , n26992 , n26993 , n26994 , n26995 , n26996 , n26997 , n26998 , n26999 , n27000 , n27001 , n27002 , n27003 , n27004 , n27005 , n27006 , n27007 , n27008 , n27009 , n27010 , n27011 , n27012 , n27013 , n27014 , n27015 , n27016 , n27017 , n27018 , n27019 , n27020 , n27021 , n27022 , n27023 , n27024 , n27025 , n27026 , n27027 , n27028 , n27029 , n27030 , n27031 , n27032 , n27033 , n27034 , n27035 , n27036 , n27037 , n27038 , n27039 , n27040 , n27041 , n27042 , n27043 , n27044 , n27045 , n27046 , n27047 , n27048 , n27049 , n27050 , n27051 , n27052 , n27053 , n27054 , n27055 , n27056 , n27057 , n27058 , n27059 , n27060 , n27061 , n27062 , n27063 , n27064 , n27065 , n27066 , n27067 , n27068 , n27069 , n27070 , n27071 , n27072 , n27073 , n27074 , n27075 , n27076 , n27077 , n27078 , n27079 , n27080 , n27081 , n27082 , n27083 , n27084 , n27085 , n27086 , n27087 , n27088 , n27089 , n27090 , n27091 , n27092 , n27093 , n27094 , n27095 , n27096 , n27097 , n27098 , n27099 , n27100 , n27101 , n27102 , n27103 , n27104 , n27105 , n27106 , n27107 , n27108 , n27109 , n27110 , n27111 , n27112 , n27113 , n27114 , n27115 , n27116 , n27117 , n27118 , n27119 , n27120 , n27121 , n27122 , n27123 , n27124 , n27125 , n27126 , n27127 , n27128 , n27129 , n27130 , n27131 , n27132 , n27133 , n27134 , n27135 , n27136 , n27137 , n27138 , n27139 , n27140 , n27141 , n27142 , n27143 , n27144 , n27145 , n27146 , n27147 , n27148 , n27149 , n27150 , n27151 , n27152 , n27153 , n27154 , n27155 , n27156 , n27157 , n27158 , n27159 , n27160 , n27161 , n27162 , n27163 , n27164 , n27165 , n27166 , n27167 , n27168 , n27169 , n27170 , n27171 , n27172 , n27173 , n27174 , n27175 , n27176 , n27177 , n27178 , n27179 , n27180 , n27181 , n27182 , n27183 , n27184 , n27185 , n27186 , n27187 , n27188 , n27189 , n27190 , n27191 , n27192 , n27193 , n27194 , n27195 , n27196 , n27197 , n27198 , n27199 , n27200 , n27201 , n27202 , n27203 , n27204 , n27205 , n27206 , n27207 , n27208 , n27209 , n27210 , n27211 , n27212 , n27213 , n27214 , n27215 , n27216 , n27217 , n27218 , n27219 , n27220 , n27221 , n27222 , n27223 , n27224 , n27225 , n27226 , n27227 , n27228 , n27229 , n27230 , n27231 , n27232 , n27233 , n27234 , n27235 , n27236 , n27237 , n27238 , n27239 , n27240 , n27241 , n27242 , n27243 , n27244 , n27245 , n27246 , n27247 , n27248 , n27249 , n27250 , n27251 , n27252 , n27253 , n27254 , n27255 , n27256 , n27257 , n27258 , n27259 , n27260 , n27261 , n27262 , n27263 , n27264 , n27265 , n27266 , n27267 , n27268 , n27269 , n27270 , n27271 , n27272 , n27273 , n27274 , n27275 , n27276 , n27277 , n27278 , n27279 , n27280 , n27281 , n27282 , n27283 , n27284 , n27285 , n27286 , n27287 , n27288 , n27289 , n27290 , n27291 , n27292 , n27293 , n27294 , n27295 , n27296 , n27297 , n27298 , n27299 , n27300 , n27301 , n27302 , n27303 , n27304 , n27305 , n27306 , n27307 , n27308 , n27309 , n27310 , n27311 , n27312 , n27313 , n27314 , n27315 , n27316 , n27317 , n27318 , n27319 , n27320 , n27321 , n27322 , n27323 , n27324 , n27325 , n27326 , n27327 , n27328 , n27329 , n27330 , n27331 , n27332 , n27333 , n27334 , n27335 , n27336 , n27337 , n27338 , n27339 , n27340 , n27341 , n27342 , n27343 , n27344 , n27345 , n27346 , n27347 , n27348 , n27349 , n27350 , n27351 , n27352 , n27353 , n27354 , n27355 , n27356 , n27357 , n27358 , n27359 , n27360 , n27361 , n27362 , n27363 , n27364 , n27365 , n27366 , n27367 , n27368 , n27369 , n27370 , n27371 , n27372 , n27373 , n27374 , n27375 , n27376 , n27377 , n27378 , n27379 , n27380 , n27381 , n27382 , n27383 , n27384 , n27385 , n27386 , n27387 , n27388 , n27389 , n27390 , n27391 , n27392 , n27393 , n27394 , n27395 , n27396 , n27397 , n27398 , n27399 , n27400 , n27401 , n27402 , n27403 , n27404 , n27405 , n27406 , n27407 , n27408 , n27409 , n27410 , n27411 , n27412 , n27413 , n27414 , n27415 , n27416 , n27417 , n27418 , n27419 , n27420 , n27421 , n27422 , n27423 , n27424 , n27425 , n27426 , n27427 , n27428 , n27429 , n27430 , n27431 , n27432 , n27433 , n27434 , n27435 , n27436 , n27437 , n27438 , n27439 , n27440 , n27441 , n27442 , n27443 , n27444 , n27445 , n27446 , n27447 , n27448 , n27449 , n27450 , n27451 , n27452 , n27453 , n27454 , n27455 , n27456 , n27457 , n27458 , n27459 , n27460 , n27461 , n27462 , n27463 , n27464 , n27465 , n27466 , n27467 , n27468 , n27469 , n27470 , n27471 , n27472 , n27473 , n27474 , n27475 , n27476 , n27477 , n27478 , n27479 , n27480 , n27481 , n27482 , n27483 , n27484 , n27485 , n27486 , n27487 , n27488 , n27489 , n27490 , n27491 , n27492 , n27493 , n27494 , n27495 , n27496 , n27497 , n27498 , n27499 , n27500 , n27501 , n27502 , n27503 , n27504 , n27505 , n27506 , n27507 , n27508 , n27509 , n27510 , n27511 , n27512 , n27513 , n27514 , n27515 , n27516 , n27517 , n27518 , n27519 , n27520 , n27521 , n27522 , n27523 , n27524 , n27525 , n27526 , n27527 , n27528 , n27529 , n27530 , n27531 , n27532 , n27533 , n27534 , n27535 , n27536 , n27537 , n27538 , n27539 , n27540 , n27541 , n27542 , n27543 , n27544 , n27545 , n27546 , n27547 , n27548 , n27549 , n27550 , n27551 , n27552 , n27553 , n27554 , n27555 , n27556 , n27557 , n27558 , n27559 , n27560 , n27561 , n27562 , n27563 , n27564 , n27565 , n27566 , n27567 , n27568 , n27569 , n27570 , n27571 , n27572 , n27573 , n27574 , n27575 , n27576 , n27577 , n27578 , n27579 , n27580 , n27581 , n27582 , n27583 , n27584 , n27585 , n27586 , n27587 , n27588 , n27589 , n27590 , n27591 , n27592 , n27593 , n27594 , n27595 , n27596 , n27597 , n27598 , n27599 , n27600 , n27601 , n27602 , n27603 , n27604 , n27605 , n27606 , n27607 , n27608 , n27609 , n27610 , n27611 , n27612 , n27613 , n27614 , n27615 , n27616 , n27617 , n27618 , n27619 , n27620 , n27621 , n27622 , n27623 , n27624 , n27625 , n27626 , n27627 , n27628 , n27629 , n27630 , n27631 , n27632 , n27633 , n27634 , n27635 , n27636 , n27637 , n27638 , n27639 , n27640 , n27641 , n27642 , n27643 , n27644 , n27645 , n27646 , n27647 , n27648 , n27649 , n27650 , n27651 , n27652 , n27653 , n27654 , n27655 , n27656 , n27657 , n27658 , n27659 , n27660 , n27661 , n27662 , n27663 , n27664 , n27665 , n27666 , n27667 , n27668 , n27669 , n27670 , n27671 , n27672 , n27673 , n27674 , n27675 , n27676 , n27677 , n27678 , n27679 , n27680 , n27681 , n27682 , n27683 , n27684 , n27685 , n27686 , n27687 , n27688 , n27689 , n27690 , n27691 , n27692 , n27693 , n27694 , n27695 , n27696 , n27697 , n27698 , n27699 , n27700 , n27701 , n27702 , n27703 , n27704 , n27705 , n27706 , n27707 , n27708 , n27709 , n27710 , n27711 , n27712 , n27713 , n27714 , n27715 , n27716 , n27717 , n27718 , n27719 , n27720 , n27721 , n27722 , n27723 , n27724 , n27725 , n27726 , n27727 , n27728 , n27729 , n27730 , n27731 , n27732 , n27733 , n27734 , n27735 , n27736 , n27737 , n27738 , n27739 , n27740 , n27741 , n27742 , n27743 , n27744 , n27745 , n27746 , n27747 , n27748 , n27749 , n27750 , n27751 , n27752 , n27753 , n27754 , n27755 , n27756 , n27757 , n27758 , n27759 , n27760 , n27761 , n27762 , n27763 , n27764 , n27765 , n27766 , n27767 , n27768 , n27769 , n27770 , n27771 , n27772 , n27773 , n27774 , n27775 , n27776 , n27777 , n27778 , n27779 , n27780 , n27781 , n27782 , n27783 , n27784 , n27785 , n27786 , n27787 , n27788 , n27789 , n27790 , n27791 , n27792 , n27793 , n27794 , n27795 , n27796 , n27797 , n27798 , n27799 , n27800 , n27801 , n27802 , n27803 , n27804 , n27805 , n27806 , n27807 , n27808 , n27809 , n27810 , n27811 , n27812 , n27813 , n27814 , n27815 , n27816 , n27817 , n27818 , n27819 , n27820 , n27821 , n27822 , n27823 , n27824 , n27825 , n27826 , n27827 , n27828 , n27829 , n27830 , n27831 , n27832 , n27833 , n27834 , n27835 , n27836 , n27837 , n27838 , n27839 , n27840 , n27841 , n27842 , n27843 , n27844 , n27845 , n27846 , n27847 , n27848 , n27849 , n27850 , n27851 , n27852 , n27853 , n27854 , n27855 , n27856 , n27857 , n27858 , n27859 , n27860 , n27861 , n27862 , n27863 , n27864 , n27865 , n27866 , n27867 , n27868 , n27869 , n27870 , n27871 , n27872 , n27873 , n27874 , n27875 , n27876 , n27877 , n27878 , n27879 , n27880 , n27881 , n27882 , n27883 , n27884 , n27885 , n27886 , n27887 , n27888 , n27889 , n27890 , n27891 , n27892 , n27893 , n27894 , n27895 , n27896 , n27897 , n27898 , n27899 , n27900 , n27901 , n27902 , n27903 , n27904 , n27905 , n27906 , n27907 , n27908 , n27909 , n27910 , n27911 , n27912 , n27913 , n27914 , n27915 , n27916 , n27917 , n27918 , n27919 , n27920 , n27921 , n27922 , n27923 , n27924 , n27925 , n27926 , n27927 , n27928 , n27929 , n27930 , n27931 , n27932 , n27933 , n27934 , n27935 , n27936 , n27937 , n27938 , n27939 , n27940 , n27941 , n27942 , n27943 , n27944 , n27945 , n27946 , n27947 , n27948 , n27949 , n27950 , n27951 , n27952 , n27953 , n27954 , n27955 , n27956 , n27957 , n27958 , n27959 , n27960 , n27961 , n27962 , n27963 , n27964 , n27965 , n27966 , n27967 , n27968 , n27969 , n27970 , n27971 , n27972 , n27973 , n27974 , n27975 , n27976 , n27977 , n27978 , n27979 , n27980 , n27981 , n27982 , n27983 , n27984 , n27985 , n27986 , n27987 , n27988 , n27989 , n27990 , n27991 , n27992 , n27993 , n27994 , n27995 , n27996 , n27997 , n27998 , n27999 , n28000 , n28001 , n28002 , n28003 , n28004 , n28005 , n28006 , n28007 , n28008 , n28009 , n28010 , n28011 , n28012 , n28013 , n28014 , n28015 , n28016 , n28017 , n28018 , n28019 , n28020 , n28021 , n28022 , n28023 , n28024 , n28025 , n28026 , n28027 , n28028 , n28029 , n28030 , n28031 , n28032 , n28033 , n28034 , n28035 , n28036 , n28037 , n28038 , n28039 , n28040 , n28041 , n28042 , n28043 , n28044 , n28045 , n28046 , n28047 , n28048 , n28049 , n28050 , n28051 , n28052 , n28053 , n28054 , n28055 , n28056 , n28057 , n28058 , n28059 , n28060 , n28061 , n28062 , n28063 , n28064 , n28065 , n28066 , n28067 , n28068 , n28069 , n28070 , n28071 , n28072 , n28073 , n28074 , n28075 , n28076 , n28077 , n28078 , n28079 , n28080 , n28081 , n28082 , n28083 , n28084 , n28085 , n28086 , n28087 , n28088 , n28089 , n28090 , n28091 , n28092 , n28093 , n28094 , n28095 , n28096 , n28097 , n28098 , n28099 , n28100 , n28101 , n28102 , n28103 , n28104 , n28105 , n28106 , n28107 , n28108 , n28109 , n28110 , n28111 , n28112 , n28113 , n28114 , n28115 , n28116 , n28117 , n28118 , n28119 , n28120 , n28121 , n28122 , n28123 , n28124 , n28125 , n28126 , n28127 , n28128 , n28129 , n28130 , n28131 , n28132 , n28133 , n28134 , n28135 , n28136 , n28137 , n28138 , n28139 , n28140 , n28141 , n28142 , n28143 , n28144 , n28145 , n28146 , n28147 , n28148 , n28149 , n28150 , n28151 , n28152 , n28153 , n28154 , n28155 , n28156 , n28157 , n28158 , n28159 , n28160 , n28161 , n28162 , n28163 , n28164 , n28165 , n28166 , n28167 , n28168 , n28169 , n28170 , n28171 , n28172 , n28173 , n28174 , n28175 , n28176 , n28177 , n28178 , n28179 , n28180 , n28181 , n28182 , n28183 , n28184 , n28185 , n28186 , n28187 , n28188 , n28189 , n28190 , n28191 , n28192 , n28193 , n28194 , n28195 , n28196 , n28197 , n28198 , n28199 , n28200 , n28201 , n28202 , n28203 , n28204 , n28205 , n28206 , n28207 , n28208 , n28209 , n28210 , n28211 , n28212 , n28213 , n28214 , n28215 , n28216 , n28217 , n28218 , n28219 , n28220 , n28221 , n28222 , n28223 , n28224 , n28225 , n28226 , n28227 , n28228 , n28229 , n28230 , n28231 , n28232 , n28233 , n28234 , n28235 , n28236 , n28237 , n28238 , n28239 , n28240 , n28241 , n28242 , n28243 , n28244 , n28245 , n28246 , n28247 , n28248 , n28249 , n28250 , n28251 , n28252 , n28253 , n28254 , n28255 , n28256 , n28257 , n28258 , n28259 , n28260 , n28261 , n28262 , n28263 , n28264 , n28265 , n28266 , n28267 , n28268 , n28269 , n28270 , n28271 , n28272 , n28273 , n28274 , n28275 , n28276 , n28277 , n28278 , n28279 , n28280 , n28281 , n28282 , n28283 , n28284 , n28285 , n28286 , n28287 , n28288 , n28289 , n28290 , n28291 , n28292 , n28293 , n28294 , n28295 , n28296 , n28297 , n28298 , n28299 , n28300 , n28301 , n28302 , n28303 , n28304 , n28305 , n28306 , n28307 , n28308 , n28309 , n28310 , n28311 , n28312 , n28313 , n28314 , n28315 , n28316 , n28317 , n28318 , n28319 , n28320 , n28321 , n28322 , n28323 , n28324 , n28325 , n28326 , n28327 , n28328 , n28329 , n28330 , n28331 , n28332 , n28333 , n28334 , n28335 , n28336 , n28337 , n28338 , n28339 , n28340 , n28341 , n28342 , n28343 , n28344 , n28345 , n28346 , n28347 , n28348 , n28349 , n28350 , n28351 , n28352 , n28353 , n28354 , n28355 , n28356 , n28357 , n28358 , n28359 , n28360 , n28361 , n28362 , n28363 , n28364 , n28365 , n28366 , n28367 , n28368 , n28369 , n28370 , n28371 , n28372 , n28373 , n28374 , n28375 , n28376 , n28377 , n28378 , n28379 , n28380 , n28381 , n28382 , n28383 , n28384 , n28385 , n28386 , n28387 , n28388 , n28389 , n28390 , n28391 , n28392 , n28393 , n28394 , n28395 , n28396 , n28397 , n28398 , n28399 , n28400 , n28401 , n28402 , n28403 , n28404 , n28405 , n28406 , n28407 , n28408 , n28409 , n28410 , n28411 , n28412 , n28413 , n28414 , n28415 , n28416 , n28417 , n28418 , n28419 , n28420 , n28421 , n28422 , n28423 , n28424 , n28425 , n28426 , n28427 , n28428 , n28429 , n28430 , n28431 , n28432 , n28433 , n28434 , n28435 , n28436 , n28437 , n28438 , n28439 , n28440 , n28441 , n28442 , n28443 , n28444 , n28445 , n28446 , n28447 , n28448 , n28449 , n28450 , n28451 , n28452 , n28453 , n28454 , n28455 , n28456 , n28457 , n28458 , n28459 , n28460 , n28461 , n28462 , n28463 , n28464 , n28465 , n28466 , n28467 , n28468 , n28469 , n28470 , n28471 , n28472 , n28473 , n28474 , n28475 , n28476 , n28477 , n28478 , n28479 , n28480 , n28481 , n28482 , n28483 , n28484 , n28485 , n28486 , n28487 , n28488 , n28489 , n28490 , n28491 , n28492 , n28493 , n28494 , n28495 , n28496 , n28497 , n28498 , n28499 , n28500 , n28501 , n28502 , n28503 , n28504 , n28505 , n28506 , n28507 , n28508 , n28509 , n28510 , n28511 , n28512 , n28513 , n28514 , n28515 , n28516 , n28517 , n28518 , n28519 , n28520 , n28521 , n28522 , n28523 , n28524 , n28525 , n28526 , n28527 , n28528 , n28529 , n28530 , n28531 , n28532 , n28533 , n28534 , n28535 , n28536 , n28537 , n28538 , n28539 , n28540 , n28541 , n28542 , n28543 , n28544 , n28545 , n28546 , n28547 , n28548 , n28549 , n28550 , n28551 , n28552 , n28553 , n28554 , n28555 , n28556 , n28557 , n28558 , n28559 , n28560 , n28561 , n28562 , n28563 , n28564 , n28565 , n28566 , n28567 , n28568 , n28569 , n28570 , n28571 , n28572 , n28573 , n28574 , n28575 , n28576 , n28577 , n28578 , n28579 , n28580 , n28581 , n28582 , n28583 , n28584 , n28585 , n28586 , n28587 , n28588 , n28589 , n28590 , n28591 , n28592 , n28593 , n28594 , n28595 , n28596 , n28597 , n28598 , n28599 , n28600 , n28601 , n28602 , n28603 , n28604 , n28605 , n28606 , n28607 , n28608 , n28609 , n28610 , n28611 , n28612 , n28613 , n28614 , n28615 , n28616 , n28617 , n28618 , n28619 , n28620 , n28621 , n28622 , n28623 , n28624 , n28625 , n28626 , n28627 , n28628 , n28629 , n28630 , n28631 , n28632 , n28633 , n28634 , n28635 , n28636 , n28637 , n28638 , n28639 , n28640 , n28641 , n28642 , n28643 , n28644 , n28645 , n28646 , n28647 , n28648 , n28649 , n28650 , n28651 , n28652 , n28653 , n28654 , n28655 , n28656 , n28657 , n28658 , n28659 , n28660 , n28661 , n28662 , n28663 , n28664 , n28665 , n28666 , n28667 , n28668 , n28669 , n28670 , n28671 , n28672 , n28673 , n28674 , n28675 , n28676 , n28677 , n28678 , n28679 , n28680 , n28681 , n28682 , n28683 , n28684 , n28685 , n28686 , n28687 , n28688 , n28689 , n28690 , n28691 , n28692 , n28693 , n28694 , n28695 , n28696 , n28697 , n28698 , n28699 , n28700 , n28701 , n28702 , n28703 , n28704 , n28705 , n28706 , n28707 , n28708 , n28709 , n28710 , n28711 , n28712 , n28713 , n28714 , n28715 , n28716 , n28717 , n28718 , n28719 , n28720 , n28721 , n28722 , n28723 , n28724 , n28725 , n28726 , n28727 , n28728 , n28729 , n28730 , n28731 , n28732 , n28733 , n28734 , n28735 , n28736 , n28737 , n28738 , n28739 , n28740 , n28741 , n28742 , n28743 , n28744 , n28745 , n28746 , n28747 , n28748 , n28749 , n28750 , n28751 , n28752 , n28753 , n28754 , n28755 , n28756 , n28757 , n28758 , n28759 , n28760 , n28761 , n28762 , n28763 , n28764 , n28765 , n28766 , n28767 , n28768 , n28769 , n28770 , n28771 , n28772 , n28773 , n28774 , n28775 , n28776 , n28777 , n28778 , n28779 , n28780 , n28781 , n28782 , n28783 , n28784 , n28785 , n28786 , n28787 , n28788 , n28789 , n28790 , n28791 , n28792 , n28793 , n28794 , n28795 , n28796 , n28797 , n28798 , n28799 , n28800 , n28801 , n28802 , n28803 , n28804 , n28805 , n28806 , n28807 , n28808 , n28809 , n28810 , n28811 , n28812 , n28813 , n28814 , n28815 , n28816 , n28817 , n28818 , n28819 , n28820 , n28821 , n28822 , n28823 , n28824 , n28825 , n28826 , n28827 , n28828 , n28829 , n28830 , n28831 , n28832 , n28833 , n28834 , n28835 , n28836 , n28837 , n28838 , n28839 , n28840 , n28841 , n28842 , n28843 , n28844 , n28845 , n28846 , n28847 , n28848 , n28849 , n28850 , n28851 , n28852 , n28853 , n28854 , n28855 , n28856 , n28857 , n28858 , n28859 , n28860 , n28861 , n28862 , n28863 , n28864 , n28865 , n28866 , n28867 , n28868 , n28869 , n28870 , n28871 , n28872 , n28873 , n28874 , n28875 , n28876 , n28877 , n28878 , n28879 , n28880 , n28881 , n28882 , n28883 , n28884 , n28885 , n28886 , n28887 , n28888 , n28889 , n28890 , n28891 , n28892 , n28893 , n28894 , n28895 , n28896 , n28897 , n28898 , n28899 , n28900 , n28901 , n28902 , n28903 , n28904 , n28905 , n28906 , n28907 , n28908 , n28909 , n28910 , n28911 , n28912 , n28913 , n28914 , n28915 , n28916 , n28917 , n28918 , n28919 , n28920 , n28921 , n28922 , n28923 , n28924 , n28925 , n28926 , n28927 , n28928 , n28929 , n28930 , n28931 , n28932 , n28933 , n28934 , n28935 , n28936 , n28937 , n28938 , n28939 , n28940 , n28941 , n28942 , n28943 , n28944 , n28945 , n28946 , n28947 , n28948 , n28949 , n28950 , n28951 , n28952 , n28953 , n28954 , n28955 , n28956 , n28957 , n28958 , n28959 , n28960 , n28961 , n28962 , n28963 , n28964 , n28965 , n28966 , n28967 , n28968 , n28969 , n28970 , n28971 , n28972 , n28973 , n28974 , n28975 , n28976 , n28977 , n28978 , n28979 , n28980 , n28981 , n28982 , n28983 , n28984 , n28985 , n28986 , n28987 , n28988 , n28989 , n28990 , n28991 , n28992 , n28993 , n28994 , n28995 , n28996 , n28997 , n28998 , n28999 , n29000 , n29001 , n29002 , n29003 , n29004 , n29005 , n29006 , n29007 , n29008 , n29009 , n29010 , n29011 , n29012 , n29013 , n29014 , n29015 , n29016 , n29017 , n29018 , n29019 , n29020 , n29021 , n29022 , n29023 , n29024 , n29025 , n29026 , n29027 , n29028 , n29029 , n29030 , n29031 , n29032 , n29033 , n29034 , n29035 , n29036 , n29037 , n29038 , n29039 , n29040 , n29041 , n29042 , n29043 , n29044 , n29045 , n29046 , n29047 , n29048 , n29049 , n29050 , n29051 , n29052 , n29053 , n29054 , n29055 , n29056 , n29057 , n29058 , n29059 , n29060 , n29061 , n29062 , n29063 , n29064 , n29065 , n29066 , n29067 , n29068 , n29069 , n29070 , n29071 , n29072 , n29073 , n29074 , n29075 , n29076 , n29077 , n29078 , n29079 , n29080 , n29081 , n29082 , n29083 , n29084 , n29085 , n29086 , n29087 , n29088 , n29089 , n29090 , n29091 , n29092 , n29093 , n29094 , n29095 , n29096 , n29097 , n29098 , n29099 , n29100 , n29101 , n29102 , n29103 , n29104 , n29105 , n29106 , n29107 , n29108 , n29109 , n29110 , n29111 , n29112 , n29113 , n29114 , n29115 , n29116 , n29117 , n29118 , n29119 , n29120 , n29121 , n29122 , n29123 , n29124 , n29125 , n29126 , n29127 , n29128 , n29129 , n29130 , n29131 , n29132 , n29133 , n29134 , n29135 , n29136 , n29137 , n29138 , n29139 , n29140 , n29141 , n29142 , n29143 , n29144 , n29145 , n29146 , n29147 , n29148 , n29149 , n29150 , n29151 , n29152 , n29153 , n29154 , n29155 , n29156 , n29157 , n29158 , n29159 , n29160 , n29161 , n29162 , n29163 , n29164 , n29165 , n29166 , n29167 , n29168 , n29169 , n29170 , n29171 , n29172 , n29173 , n29174 , n29175 , n29176 , n29177 , n29178 , n29179 , n29180 , n29181 , n29182 , n29183 , n29184 , n29185 , n29186 , n29187 , n29188 , n29189 , n29190 , n29191 , n29192 , n29193 , n29194 , n29195 , n29196 , n29197 , n29198 , n29199 , n29200 , n29201 , n29202 , n29203 , n29204 , n29205 , n29206 , n29207 , n29208 , n29209 , n29210 , n29211 , n29212 , n29213 , n29214 , n29215 , n29216 , n29217 , n29218 , n29219 , n29220 , n29221 , n29222 , n29223 , n29224 , n29225 , n29226 , n29227 , n29228 , n29229 , n29230 , n29231 , n29232 , n29233 , n29234 , n29235 , n29236 , n29237 , n29238 , n29239 , n29240 , n29241 , n29242 , n29243 , n29244 , n29245 , n29246 , n29247 , n29248 , n29249 , n29250 , n29251 , n29252 , n29253 , n29254 , n29255 , n29256 , n29257 , n29258 , n29259 , n29260 , n29261 , n29262 , n29263 , n29264 , n29265 , n29266 , n29267 , n29268 , n29269 , n29270 , n29271 , n29272 , n29273 , n29274 , n29275 , n29276 , n29277 , n29278 , n29279 , n29280 , n29281 , n29282 , n29283 , n29284 , n29285 , n29286 , n29287 , n29288 , n29289 , n29290 , n29291 , n29292 , n29293 , n29294 , n29295 , n29296 , n29297 , n29298 , n29299 , n29300 , n29301 , n29302 , n29303 , n29304 , n29305 , n29306 , n29307 , n29308 , n29309 , n29310 , n29311 , n29312 , n29313 , n29314 , n29315 , n29316 , n29317 , n29318 , n29319 , n29320 , n29321 , n29322 , n29323 , n29324 , n29325 , n29326 , n29327 , n29328 , n29329 , n29330 , n29331 , n29332 , n29333 , n29334 , n29335 , n29336 , n29337 , n29338 , n29339 , n29340 , n29341 , n29342 , n29343 , n29344 , n29345 , n29346 , n29347 , n29348 , n29349 , n29350 , n29351 , n29352 , n29353 , n29354 , n29355 , n29356 , n29357 , n29358 , n29359 , n29360 , n29361 , n29362 , n29363 , n29364 , n29365 , n29366 , n29367 , n29368 , n29369 , n29370 , n29371 , n29372 , n29373 , n29374 , n29375 , n29376 , n29377 , n29378 , n29379 , n29380 , n29381 , n29382 , n29383 , n29384 , n29385 , n29386 , n29387 , n29388 , n29389 , n29390 , n29391 , n29392 , n29393 , n29394 , n29395 , n29396 , n29397 , n29398 , n29399 , n29400 , n29401 , n29402 , n29403 , n29404 , n29405 , n29406 , n29407 , n29408 , n29409 , n29410 , n29411 , n29412 , n29413 , n29414 , n29415 , n29416 , n29417 , n29418 , n29419 , n29420 , n29421 , n29422 , n29423 , n29424 , n29425 , n29426 , n29427 , n29428 , n29429 , n29430 , n29431 , n29432 , n29433 , n29434 , n29435 , n29436 , n29437 , n29438 , n29439 , n29440 , n29441 , n29442 , n29443 , n29444 , n29445 , n29446 , n29447 , n29448 , n29449 , n29450 , n29451 , n29452 , n29453 , n29454 , n29455 , n29456 , n29457 , n29458 , n29459 , n29460 , n29461 , n29462 , n29463 , n29464 , n29465 , n29466 , n29467 , n29468 , n29469 , n29470 , n29471 , n29472 , n29473 , n29474 , n29475 , n29476 , n29477 , n29478 , n29479 , n29480 , n29481 , n29482 , n29483 , n29484 , n29485 , n29486 , n29487 , n29488 , n29489 , n29490 , n29491 , n29492 , n29493 , n29494 , n29495 , n29496 , n29497 , n29498 , n29499 , n29500 , n29501 , n29502 , n29503 , n29504 , n29505 , n29506 , n29507 , n29508 , n29509 , n29510 , n29511 , n29512 , n29513 , n29514 , n29515 , n29516 , n29517 , n29518 , n29519 , n29520 , n29521 , n29522 , n29523 , n29524 , n29525 , n29526 , n29527 , n29528 , n29529 , n29530 , n29531 , n29532 , n29533 , n29534 , n29535 , n29536 , n29537 , n29538 , n29539 , n29540 , n29541 , n29542 , n29543 , n29544 , n29545 , n29546 , n29547 , n29548 , n29549 , n29550 , n29551 , n29552 , n29553 , n29554 , n29555 , n29556 , n29557 , n29558 , n29559 , n29560 , n29561 , n29562 , n29563 , n29564 , n29565 , n29566 , n29567 , n29568 , n29569 , n29570 , n29571 , n29572 , n29573 , n29574 , n29575 , n29576 , n29577 , n29578 , n29579 , n29580 , n29581 , n29582 , n29583 , n29584 , n29585 , n29586 , n29587 , n29588 , n29589 , n29590 , n29591 , n29592 , n29593 , n29594 , n29595 , n29596 , n29597 , n29598 , n29599 , n29600 , n29601 , n29602 , n29603 , n29604 , n29605 , n29606 , n29607 , n29608 , n29609 , n29610 , n29611 , n29612 , n29613 , n29614 , n29615 , n29616 , n29617 , n29618 , n29619 , n29620 , n29621 , n29622 , n29623 , n29624 , n29625 , n29626 , n29627 , n29628 , n29629 , n29630 , n29631 , n29632 , n29633 , n29634 , n29635 , n29636 , n29637 , n29638 , n29639 , n29640 , n29641 , n29642 , n29643 , n29644 , n29645 , n29646 , n29647 , n29648 , n29649 , n29650 , n29651 , n29652 , n29653 , n29654 , n29655 , n29656 , n29657 , n29658 , n29659 , n29660 , n29661 , n29662 , n29663 , n29664 , n29665 , n29666 , n29667 , n29668 , n29669 , n29670 , n29671 , n29672 , n29673 , n29674 , n29675 , n29676 , n29677 , n29678 , n29679 , n29680 , n29681 , n29682 , n29683 , n29684 , n29685 , n29686 , n29687 , n29688 , n29689 , n29690 , n29691 , n29692 , n29693 , n29694 , n29695 , n29696 , n29697 , n29698 , n29699 , n29700 , n29701 , n29702 , n29703 , n29704 , n29705 , n29706 , n29707 , n29708 , n29709 , n29710 , n29711 , n29712 , n29713 , n29714 , n29715 , n29716 , n29717 , n29718 , n29719 , n29720 , n29721 , n29722 , n29723 , n29724 , n29725 , n29726 , n29727 , n29728 , n29729 , n29730 , n29731 , n29732 , n29733 , n29734 , n29735 , n29736 , n29737 , n29738 , n29739 , n29740 , n29741 , n29742 , n29743 , n29744 , n29745 , n29746 , n29747 , n29748 , n29749 , n29750 , n29751 , n29752 , n29753 , n29754 , n29755 , n29756 , n29757 , n29758 , n29759 , n29760 , n29761 , n29762 , n29763 , n29764 , n29765 , n29766 , n29767 , n29768 , n29769 , n29770 , n29771 , n29772 , n29773 , n29774 , n29775 , n29776 , n29777 , n29778 , n29779 , n29780 , n29781 , n29782 , n29783 , n29784 , n29785 , n29786 , n29787 , n29788 , n29789 , n29790 , n29791 , n29792 , n29793 , n29794 , n29795 , n29796 , n29797 , n29798 , n29799 , n29800 , n29801 , n29802 , n29803 , n29804 , n29805 , n29806 ;
  assign n1349 = ~\P1_Datao_reg[30]/NET0131  & ~\P2_Datao_reg[30]/NET0131  ;
  assign n1350 = ~\datao[30]_pad  & n1349 ;
  assign n1351 = \P2_Address_reg[0]/NET0131  & ~n1350 ;
  assign n1352 = \P3_Address_reg[0]/NET0131  & n1350 ;
  assign n1353 = ~n1351 & ~n1352 ;
  assign n1354 = \P2_Address_reg[10]/NET0131  & ~n1350 ;
  assign n1355 = \P3_Address_reg[10]/NET0131  & n1350 ;
  assign n1356 = ~n1354 & ~n1355 ;
  assign n1357 = \P2_Address_reg[11]/NET0131  & ~n1350 ;
  assign n1358 = \P3_Address_reg[11]/NET0131  & n1350 ;
  assign n1359 = ~n1357 & ~n1358 ;
  assign n1360 = \P2_Address_reg[12]/NET0131  & ~n1350 ;
  assign n1361 = \P3_Address_reg[12]/NET0131  & n1350 ;
  assign n1362 = ~n1360 & ~n1361 ;
  assign n1363 = \P2_Address_reg[13]/NET0131  & ~n1350 ;
  assign n1364 = \P3_Address_reg[13]/NET0131  & n1350 ;
  assign n1365 = ~n1363 & ~n1364 ;
  assign n1366 = \P2_Address_reg[14]/NET0131  & ~n1350 ;
  assign n1367 = \P3_Address_reg[14]/NET0131  & n1350 ;
  assign n1368 = ~n1366 & ~n1367 ;
  assign n1369 = \P2_Address_reg[15]/NET0131  & ~n1350 ;
  assign n1370 = \P3_Address_reg[15]/NET0131  & n1350 ;
  assign n1371 = ~n1369 & ~n1370 ;
  assign n1372 = \P2_Address_reg[16]/NET0131  & ~n1350 ;
  assign n1373 = \P3_Address_reg[16]/NET0131  & n1350 ;
  assign n1374 = ~n1372 & ~n1373 ;
  assign n1375 = \P2_Address_reg[17]/NET0131  & ~n1350 ;
  assign n1376 = \P3_Address_reg[17]/NET0131  & n1350 ;
  assign n1377 = ~n1375 & ~n1376 ;
  assign n1378 = \P2_Address_reg[18]/NET0131  & ~n1350 ;
  assign n1379 = \P3_Address_reg[18]/NET0131  & n1350 ;
  assign n1380 = ~n1378 & ~n1379 ;
  assign n1381 = \P2_Address_reg[19]/NET0131  & ~n1350 ;
  assign n1382 = \P3_Address_reg[19]/NET0131  & n1350 ;
  assign n1383 = ~n1381 & ~n1382 ;
  assign n1384 = \P2_Address_reg[1]/NET0131  & ~n1350 ;
  assign n1385 = \P3_Address_reg[1]/NET0131  & n1350 ;
  assign n1386 = ~n1384 & ~n1385 ;
  assign n1387 = \P2_Address_reg[20]/NET0131  & ~n1350 ;
  assign n1388 = \P3_Address_reg[20]/NET0131  & n1350 ;
  assign n1389 = ~n1387 & ~n1388 ;
  assign n1390 = \P2_Address_reg[21]/NET0131  & ~n1350 ;
  assign n1391 = \P3_Address_reg[21]/NET0131  & n1350 ;
  assign n1392 = ~n1390 & ~n1391 ;
  assign n1393 = \P2_Address_reg[22]/NET0131  & ~n1350 ;
  assign n1394 = \P3_Address_reg[22]/NET0131  & n1350 ;
  assign n1395 = ~n1393 & ~n1394 ;
  assign n1396 = \P2_Address_reg[23]/NET0131  & ~n1350 ;
  assign n1397 = \P3_Address_reg[23]/NET0131  & n1350 ;
  assign n1398 = ~n1396 & ~n1397 ;
  assign n1399 = \P2_Address_reg[24]/NET0131  & ~n1350 ;
  assign n1400 = \P3_Address_reg[24]/NET0131  & n1350 ;
  assign n1401 = ~n1399 & ~n1400 ;
  assign n1402 = \P2_Address_reg[25]/NET0131  & ~n1350 ;
  assign n1403 = \P3_Address_reg[25]/NET0131  & n1350 ;
  assign n1404 = ~n1402 & ~n1403 ;
  assign n1405 = \P2_Address_reg[26]/NET0131  & ~n1350 ;
  assign n1406 = \P3_Address_reg[26]/NET0131  & n1350 ;
  assign n1407 = ~n1405 & ~n1406 ;
  assign n1408 = \P2_Address_reg[27]/NET0131  & ~n1350 ;
  assign n1409 = \P3_Address_reg[27]/NET0131  & n1350 ;
  assign n1410 = ~n1408 & ~n1409 ;
  assign n1411 = \P2_Address_reg[28]/NET0131  & ~n1350 ;
  assign n1412 = \P3_Address_reg[28]/NET0131  & n1350 ;
  assign n1413 = ~n1411 & ~n1412 ;
  assign n1414 = \P2_Address_reg[29]/NET0131  & ~n1350 ;
  assign n1415 = \P3_Address_reg[29]/NET0131  & n1350 ;
  assign n1416 = ~n1414 & ~n1415 ;
  assign n1417 = \P2_Address_reg[2]/NET0131  & ~n1350 ;
  assign n1418 = \P3_Address_reg[2]/NET0131  & n1350 ;
  assign n1419 = ~n1417 & ~n1418 ;
  assign n1420 = \P2_Address_reg[3]/NET0131  & ~n1350 ;
  assign n1421 = \P3_Address_reg[3]/NET0131  & n1350 ;
  assign n1422 = ~n1420 & ~n1421 ;
  assign n1423 = \P2_Address_reg[4]/NET0131  & ~n1350 ;
  assign n1424 = \P3_Address_reg[4]/NET0131  & n1350 ;
  assign n1425 = ~n1423 & ~n1424 ;
  assign n1426 = \P2_Address_reg[5]/NET0131  & ~n1350 ;
  assign n1427 = \P3_Address_reg[5]/NET0131  & n1350 ;
  assign n1428 = ~n1426 & ~n1427 ;
  assign n1429 = \P2_Address_reg[6]/NET0131  & ~n1350 ;
  assign n1430 = \P3_Address_reg[6]/NET0131  & n1350 ;
  assign n1431 = ~n1429 & ~n1430 ;
  assign n1432 = \P2_Address_reg[7]/NET0131  & ~n1350 ;
  assign n1433 = \P3_Address_reg[7]/NET0131  & n1350 ;
  assign n1434 = ~n1432 & ~n1433 ;
  assign n1435 = \P2_Address_reg[8]/NET0131  & ~n1350 ;
  assign n1436 = \P3_Address_reg[8]/NET0131  & n1350 ;
  assign n1437 = ~n1435 & ~n1436 ;
  assign n1438 = \P2_Address_reg[9]/NET0131  & ~n1350 ;
  assign n1439 = \P3_Address_reg[9]/NET0131  & n1350 ;
  assign n1440 = ~n1438 & ~n1439 ;
  assign n1441 = \P2_InstQueueRd_Addr_reg[0]/NET0131  & \P2_InstQueueRd_Addr_reg[1]/NET0131  ;
  assign n1442 = \P2_InstQueueRd_Addr_reg[2]/NET0131  & n1441 ;
  assign n1443 = ~\P2_InstQueueRd_Addr_reg[2]/NET0131  & ~n1441 ;
  assign n1444 = ~n1442 & ~n1443 ;
  assign n1452 = ~\P2_InstQueueRd_Addr_reg[2]/NET0131  & \P2_InstQueueRd_Addr_reg[3]/NET0131  ;
  assign n1458 = ~\P2_InstQueueRd_Addr_reg[0]/NET0131  & \P2_InstQueueRd_Addr_reg[1]/NET0131  ;
  assign n1459 = n1452 & n1458 ;
  assign n1460 = \P2_InstQueue_reg[10][0]/NET0131  & n1459 ;
  assign n1446 = \P2_InstQueueRd_Addr_reg[2]/NET0131  & ~\P2_InstQueueRd_Addr_reg[3]/NET0131  ;
  assign n1461 = n1441 & n1446 ;
  assign n1462 = \P2_InstQueue_reg[7][0]/NET0131  & n1461 ;
  assign n1486 = ~n1460 & ~n1462 ;
  assign n1449 = ~\P2_InstQueueRd_Addr_reg[2]/NET0131  & ~\P2_InstQueueRd_Addr_reg[3]/NET0131  ;
  assign n1463 = ~\P2_InstQueueRd_Addr_reg[0]/NET0131  & ~\P2_InstQueueRd_Addr_reg[1]/NET0131  ;
  assign n1464 = n1449 & n1463 ;
  assign n1465 = \P2_InstQueue_reg[0][0]/NET0131  & n1464 ;
  assign n1455 = \P2_InstQueueRd_Addr_reg[2]/NET0131  & \P2_InstQueueRd_Addr_reg[3]/NET0131  ;
  assign n1466 = n1455 & n1463 ;
  assign n1467 = \P2_InstQueue_reg[12][0]/NET0131  & n1466 ;
  assign n1487 = ~n1465 & ~n1467 ;
  assign n1494 = n1486 & n1487 ;
  assign n1445 = \P2_InstQueueRd_Addr_reg[0]/NET0131  & ~\P2_InstQueueRd_Addr_reg[1]/NET0131  ;
  assign n1447 = n1445 & n1446 ;
  assign n1448 = \P2_InstQueue_reg[5][0]/NET0131  & n1447 ;
  assign n1450 = n1441 & n1449 ;
  assign n1451 = \P2_InstQueue_reg[3][0]/NET0131  & n1450 ;
  assign n1484 = ~n1448 & ~n1451 ;
  assign n1453 = n1445 & n1452 ;
  assign n1454 = \P2_InstQueue_reg[9][0]/NET0131  & n1453 ;
  assign n1456 = n1441 & n1455 ;
  assign n1457 = \P2_InstQueue_reg[15][0]/NET0131  & n1456 ;
  assign n1485 = ~n1454 & ~n1457 ;
  assign n1495 = n1484 & n1485 ;
  assign n1496 = n1494 & n1495 ;
  assign n1476 = n1446 & n1458 ;
  assign n1477 = \P2_InstQueue_reg[6][0]/NET0131  & n1476 ;
  assign n1478 = n1455 & n1458 ;
  assign n1479 = \P2_InstQueue_reg[14][0]/NET0131  & n1478 ;
  assign n1490 = ~n1477 & ~n1479 ;
  assign n1480 = n1441 & n1452 ;
  assign n1481 = \P2_InstQueue_reg[11][0]/NET0131  & n1480 ;
  assign n1482 = n1445 & n1455 ;
  assign n1483 = \P2_InstQueue_reg[13][0]/NET0131  & n1482 ;
  assign n1491 = ~n1481 & ~n1483 ;
  assign n1492 = n1490 & n1491 ;
  assign n1468 = n1445 & n1449 ;
  assign n1469 = \P2_InstQueue_reg[1][0]/NET0131  & n1468 ;
  assign n1470 = n1449 & n1458 ;
  assign n1471 = \P2_InstQueue_reg[2][0]/NET0131  & n1470 ;
  assign n1488 = ~n1469 & ~n1471 ;
  assign n1472 = n1452 & n1463 ;
  assign n1473 = \P2_InstQueue_reg[8][0]/NET0131  & n1472 ;
  assign n1474 = n1446 & n1463 ;
  assign n1475 = \P2_InstQueue_reg[4][0]/NET0131  & n1474 ;
  assign n1489 = ~n1473 & ~n1475 ;
  assign n1493 = n1488 & n1489 ;
  assign n1497 = n1492 & n1493 ;
  assign n1498 = n1496 & n1497 ;
  assign n1503 = \P2_InstQueue_reg[9][3]/NET0131  & n1453 ;
  assign n1504 = \P2_InstQueue_reg[7][3]/NET0131  & n1461 ;
  assign n1517 = ~n1503 & ~n1504 ;
  assign n1505 = \P2_InstQueue_reg[13][3]/NET0131  & n1482 ;
  assign n1506 = \P2_InstQueue_reg[4][3]/NET0131  & n1474 ;
  assign n1518 = ~n1505 & ~n1506 ;
  assign n1525 = n1517 & n1518 ;
  assign n1499 = \P2_InstQueue_reg[10][3]/NET0131  & n1459 ;
  assign n1500 = \P2_InstQueue_reg[3][3]/NET0131  & n1450 ;
  assign n1515 = ~n1499 & ~n1500 ;
  assign n1501 = \P2_InstQueue_reg[6][3]/NET0131  & n1476 ;
  assign n1502 = \P2_InstQueue_reg[12][3]/NET0131  & n1466 ;
  assign n1516 = ~n1501 & ~n1502 ;
  assign n1526 = n1515 & n1516 ;
  assign n1527 = n1525 & n1526 ;
  assign n1511 = \P2_InstQueue_reg[2][3]/NET0131  & n1470 ;
  assign n1512 = \P2_InstQueue_reg[0][3]/NET0131  & n1464 ;
  assign n1521 = ~n1511 & ~n1512 ;
  assign n1513 = \P2_InstQueue_reg[15][3]/NET0131  & n1456 ;
  assign n1514 = \P2_InstQueue_reg[14][3]/NET0131  & n1478 ;
  assign n1522 = ~n1513 & ~n1514 ;
  assign n1523 = n1521 & n1522 ;
  assign n1507 = \P2_InstQueue_reg[1][3]/NET0131  & n1468 ;
  assign n1508 = \P2_InstQueue_reg[11][3]/NET0131  & n1480 ;
  assign n1519 = ~n1507 & ~n1508 ;
  assign n1509 = \P2_InstQueue_reg[5][3]/NET0131  & n1447 ;
  assign n1510 = \P2_InstQueue_reg[8][3]/NET0131  & n1472 ;
  assign n1520 = ~n1509 & ~n1510 ;
  assign n1524 = n1519 & n1520 ;
  assign n1528 = n1523 & n1524 ;
  assign n1529 = n1527 & n1528 ;
  assign n1530 = ~n1498 & ~n1529 ;
  assign n1535 = \P2_InstQueue_reg[3][2]/NET0131  & n1450 ;
  assign n1536 = \P2_InstQueue_reg[14][2]/NET0131  & n1478 ;
  assign n1549 = ~n1535 & ~n1536 ;
  assign n1537 = \P2_InstQueue_reg[13][2]/NET0131  & n1482 ;
  assign n1538 = \P2_InstQueue_reg[4][2]/NET0131  & n1474 ;
  assign n1550 = ~n1537 & ~n1538 ;
  assign n1557 = n1549 & n1550 ;
  assign n1531 = \P2_InstQueue_reg[6][2]/NET0131  & n1476 ;
  assign n1532 = \P2_InstQueue_reg[11][2]/NET0131  & n1480 ;
  assign n1547 = ~n1531 & ~n1532 ;
  assign n1533 = \P2_InstQueue_reg[10][2]/NET0131  & n1459 ;
  assign n1534 = \P2_InstQueue_reg[8][2]/NET0131  & n1472 ;
  assign n1548 = ~n1533 & ~n1534 ;
  assign n1558 = n1547 & n1548 ;
  assign n1559 = n1557 & n1558 ;
  assign n1543 = \P2_InstQueue_reg[15][2]/NET0131  & n1456 ;
  assign n1544 = \P2_InstQueue_reg[2][2]/NET0131  & n1470 ;
  assign n1553 = ~n1543 & ~n1544 ;
  assign n1545 = \P2_InstQueue_reg[12][2]/NET0131  & n1466 ;
  assign n1546 = \P2_InstQueue_reg[0][2]/NET0131  & n1464 ;
  assign n1554 = ~n1545 & ~n1546 ;
  assign n1555 = n1553 & n1554 ;
  assign n1539 = \P2_InstQueue_reg[9][2]/NET0131  & n1453 ;
  assign n1540 = \P2_InstQueue_reg[7][2]/NET0131  & n1461 ;
  assign n1551 = ~n1539 & ~n1540 ;
  assign n1541 = \P2_InstQueue_reg[1][2]/NET0131  & n1468 ;
  assign n1542 = \P2_InstQueue_reg[5][2]/NET0131  & n1447 ;
  assign n1552 = ~n1541 & ~n1542 ;
  assign n1556 = n1551 & n1552 ;
  assign n1560 = n1555 & n1556 ;
  assign n1561 = n1559 & n1560 ;
  assign n1566 = \P2_InstQueue_reg[7][1]/NET0131  & n1461 ;
  assign n1567 = \P2_InstQueue_reg[11][1]/NET0131  & n1480 ;
  assign n1580 = ~n1566 & ~n1567 ;
  assign n1568 = \P2_InstQueue_reg[0][1]/NET0131  & n1464 ;
  assign n1569 = \P2_InstQueue_reg[10][1]/NET0131  & n1459 ;
  assign n1581 = ~n1568 & ~n1569 ;
  assign n1588 = n1580 & n1581 ;
  assign n1562 = \P2_InstQueue_reg[15][1]/NET0131  & n1456 ;
  assign n1563 = \P2_InstQueue_reg[5][1]/NET0131  & n1447 ;
  assign n1578 = ~n1562 & ~n1563 ;
  assign n1564 = \P2_InstQueue_reg[13][1]/NET0131  & n1482 ;
  assign n1565 = \P2_InstQueue_reg[12][1]/NET0131  & n1466 ;
  assign n1579 = ~n1564 & ~n1565 ;
  assign n1589 = n1578 & n1579 ;
  assign n1590 = n1588 & n1589 ;
  assign n1574 = \P2_InstQueue_reg[6][1]/NET0131  & n1476 ;
  assign n1575 = \P2_InstQueue_reg[4][1]/NET0131  & n1474 ;
  assign n1584 = ~n1574 & ~n1575 ;
  assign n1576 = \P2_InstQueue_reg[8][1]/NET0131  & n1472 ;
  assign n1577 = \P2_InstQueue_reg[14][1]/NET0131  & n1478 ;
  assign n1585 = ~n1576 & ~n1577 ;
  assign n1586 = n1584 & n1585 ;
  assign n1570 = \P2_InstQueue_reg[9][1]/NET0131  & n1453 ;
  assign n1571 = \P2_InstQueue_reg[3][1]/NET0131  & n1450 ;
  assign n1582 = ~n1570 & ~n1571 ;
  assign n1572 = \P2_InstQueue_reg[1][1]/NET0131  & n1468 ;
  assign n1573 = \P2_InstQueue_reg[2][1]/NET0131  & n1470 ;
  assign n1583 = ~n1572 & ~n1573 ;
  assign n1587 = n1582 & n1583 ;
  assign n1591 = n1586 & n1587 ;
  assign n1592 = n1590 & n1591 ;
  assign n1593 = n1561 & ~n1592 ;
  assign n1594 = n1530 & n1593 ;
  assign n1599 = \P2_InstQueue_reg[4][6]/NET0131  & n1474 ;
  assign n1600 = \P2_InstQueue_reg[2][6]/NET0131  & n1470 ;
  assign n1613 = ~n1599 & ~n1600 ;
  assign n1601 = \P2_InstQueue_reg[15][6]/NET0131  & n1456 ;
  assign n1602 = \P2_InstQueue_reg[1][6]/NET0131  & n1468 ;
  assign n1614 = ~n1601 & ~n1602 ;
  assign n1621 = n1613 & n1614 ;
  assign n1595 = \P2_InstQueue_reg[0][6]/NET0131  & n1464 ;
  assign n1596 = \P2_InstQueue_reg[11][6]/NET0131  & n1480 ;
  assign n1611 = ~n1595 & ~n1596 ;
  assign n1597 = \P2_InstQueue_reg[7][6]/NET0131  & n1461 ;
  assign n1598 = \P2_InstQueue_reg[10][6]/NET0131  & n1459 ;
  assign n1612 = ~n1597 & ~n1598 ;
  assign n1622 = n1611 & n1612 ;
  assign n1623 = n1621 & n1622 ;
  assign n1607 = \P2_InstQueue_reg[6][6]/NET0131  & n1476 ;
  assign n1608 = \P2_InstQueue_reg[9][6]/NET0131  & n1453 ;
  assign n1617 = ~n1607 & ~n1608 ;
  assign n1609 = \P2_InstQueue_reg[13][6]/NET0131  & n1482 ;
  assign n1610 = \P2_InstQueue_reg[12][6]/NET0131  & n1466 ;
  assign n1618 = ~n1609 & ~n1610 ;
  assign n1619 = n1617 & n1618 ;
  assign n1603 = \P2_InstQueue_reg[14][6]/NET0131  & n1478 ;
  assign n1604 = \P2_InstQueue_reg[8][6]/NET0131  & n1472 ;
  assign n1615 = ~n1603 & ~n1604 ;
  assign n1605 = \P2_InstQueue_reg[3][6]/NET0131  & n1450 ;
  assign n1606 = \P2_InstQueue_reg[5][6]/NET0131  & n1447 ;
  assign n1616 = ~n1605 & ~n1606 ;
  assign n1620 = n1615 & n1616 ;
  assign n1624 = n1619 & n1620 ;
  assign n1625 = n1623 & n1624 ;
  assign n1630 = \P2_InstQueue_reg[15][7]/NET0131  & n1456 ;
  assign n1631 = \P2_InstQueue_reg[2][7]/NET0131  & n1470 ;
  assign n1644 = ~n1630 & ~n1631 ;
  assign n1632 = \P2_InstQueue_reg[10][7]/NET0131  & n1459 ;
  assign n1633 = \P2_InstQueue_reg[9][7]/NET0131  & n1453 ;
  assign n1645 = ~n1632 & ~n1633 ;
  assign n1652 = n1644 & n1645 ;
  assign n1626 = \P2_InstQueue_reg[0][7]/NET0131  & n1464 ;
  assign n1627 = \P2_InstQueue_reg[11][7]/NET0131  & n1480 ;
  assign n1642 = ~n1626 & ~n1627 ;
  assign n1628 = \P2_InstQueue_reg[3][7]/NET0131  & n1450 ;
  assign n1629 = \P2_InstQueue_reg[12][7]/NET0131  & n1466 ;
  assign n1643 = ~n1628 & ~n1629 ;
  assign n1653 = n1642 & n1643 ;
  assign n1654 = n1652 & n1653 ;
  assign n1638 = \P2_InstQueue_reg[6][7]/NET0131  & n1476 ;
  assign n1639 = \P2_InstQueue_reg[1][7]/NET0131  & n1468 ;
  assign n1648 = ~n1638 & ~n1639 ;
  assign n1640 = \P2_InstQueue_reg[13][7]/NET0131  & n1482 ;
  assign n1641 = \P2_InstQueue_reg[4][7]/NET0131  & n1474 ;
  assign n1649 = ~n1640 & ~n1641 ;
  assign n1650 = n1648 & n1649 ;
  assign n1634 = \P2_InstQueue_reg[14][7]/NET0131  & n1478 ;
  assign n1635 = \P2_InstQueue_reg[8][7]/NET0131  & n1472 ;
  assign n1646 = ~n1634 & ~n1635 ;
  assign n1636 = \P2_InstQueue_reg[7][7]/NET0131  & n1461 ;
  assign n1637 = \P2_InstQueue_reg[5][7]/NET0131  & n1447 ;
  assign n1647 = ~n1636 & ~n1637 ;
  assign n1651 = n1646 & n1647 ;
  assign n1655 = n1650 & n1651 ;
  assign n1656 = n1654 & n1655 ;
  assign n1657 = n1625 & ~n1656 ;
  assign n1662 = \P2_InstQueue_reg[5][4]/NET0131  & n1447 ;
  assign n1663 = \P2_InstQueue_reg[9][4]/NET0131  & n1453 ;
  assign n1676 = ~n1662 & ~n1663 ;
  assign n1664 = \P2_InstQueue_reg[0][4]/NET0131  & n1464 ;
  assign n1665 = \P2_InstQueue_reg[10][4]/NET0131  & n1459 ;
  assign n1677 = ~n1664 & ~n1665 ;
  assign n1684 = n1676 & n1677 ;
  assign n1658 = \P2_InstQueue_reg[2][4]/NET0131  & n1470 ;
  assign n1659 = \P2_InstQueue_reg[13][4]/NET0131  & n1482 ;
  assign n1674 = ~n1658 & ~n1659 ;
  assign n1660 = \P2_InstQueue_reg[7][4]/NET0131  & n1461 ;
  assign n1661 = \P2_InstQueue_reg[14][4]/NET0131  & n1478 ;
  assign n1675 = ~n1660 & ~n1661 ;
  assign n1685 = n1674 & n1675 ;
  assign n1686 = n1684 & n1685 ;
  assign n1670 = \P2_InstQueue_reg[4][4]/NET0131  & n1474 ;
  assign n1671 = \P2_InstQueue_reg[12][4]/NET0131  & n1466 ;
  assign n1680 = ~n1670 & ~n1671 ;
  assign n1672 = \P2_InstQueue_reg[8][4]/NET0131  & n1472 ;
  assign n1673 = \P2_InstQueue_reg[6][4]/NET0131  & n1476 ;
  assign n1681 = ~n1672 & ~n1673 ;
  assign n1682 = n1680 & n1681 ;
  assign n1666 = \P2_InstQueue_reg[1][4]/NET0131  & n1468 ;
  assign n1667 = \P2_InstQueue_reg[3][4]/NET0131  & n1450 ;
  assign n1678 = ~n1666 & ~n1667 ;
  assign n1668 = \P2_InstQueue_reg[11][4]/NET0131  & n1480 ;
  assign n1669 = \P2_InstQueue_reg[15][4]/NET0131  & n1456 ;
  assign n1679 = ~n1668 & ~n1669 ;
  assign n1683 = n1678 & n1679 ;
  assign n1687 = n1682 & n1683 ;
  assign n1688 = n1686 & n1687 ;
  assign n1689 = n1657 & ~n1688 ;
  assign n1694 = \P2_InstQueue_reg[4][5]/NET0131  & n1474 ;
  assign n1695 = \P2_InstQueue_reg[1][5]/NET0131  & n1468 ;
  assign n1708 = ~n1694 & ~n1695 ;
  assign n1696 = \P2_InstQueue_reg[2][5]/NET0131  & n1470 ;
  assign n1697 = \P2_InstQueue_reg[8][5]/NET0131  & n1472 ;
  assign n1709 = ~n1696 & ~n1697 ;
  assign n1716 = n1708 & n1709 ;
  assign n1690 = \P2_InstQueue_reg[12][5]/NET0131  & n1466 ;
  assign n1691 = \P2_InstQueue_reg[5][5]/NET0131  & n1447 ;
  assign n1706 = ~n1690 & ~n1691 ;
  assign n1692 = \P2_InstQueue_reg[3][5]/NET0131  & n1450 ;
  assign n1693 = \P2_InstQueue_reg[0][5]/NET0131  & n1464 ;
  assign n1707 = ~n1692 & ~n1693 ;
  assign n1717 = n1706 & n1707 ;
  assign n1718 = n1716 & n1717 ;
  assign n1702 = \P2_InstQueue_reg[14][5]/NET0131  & n1478 ;
  assign n1703 = \P2_InstQueue_reg[11][5]/NET0131  & n1480 ;
  assign n1712 = ~n1702 & ~n1703 ;
  assign n1704 = \P2_InstQueue_reg[6][5]/NET0131  & n1476 ;
  assign n1705 = \P2_InstQueue_reg[13][5]/NET0131  & n1482 ;
  assign n1713 = ~n1704 & ~n1705 ;
  assign n1714 = n1712 & n1713 ;
  assign n1698 = \P2_InstQueue_reg[9][5]/NET0131  & n1453 ;
  assign n1699 = \P2_InstQueue_reg[7][5]/NET0131  & n1461 ;
  assign n1710 = ~n1698 & ~n1699 ;
  assign n1700 = \P2_InstQueue_reg[15][5]/NET0131  & n1456 ;
  assign n1701 = \P2_InstQueue_reg[10][5]/NET0131  & n1459 ;
  assign n1711 = ~n1700 & ~n1701 ;
  assign n1715 = n1710 & n1711 ;
  assign n1719 = n1714 & n1715 ;
  assign n1720 = n1718 & n1719 ;
  assign n1721 = n1689 & ~n1720 ;
  assign n1722 = n1594 & n1721 ;
  assign n1723 = n1498 & ~n1529 ;
  assign n1724 = n1561 & n1592 ;
  assign n1725 = n1723 & n1724 ;
  assign n1726 = n1721 & n1725 ;
  assign n1727 = ~n1722 & ~n1726 ;
  assign n1728 = ~n1625 & ~n1656 ;
  assign n1729 = n1688 & ~n1720 ;
  assign n1730 = n1728 & n1729 ;
  assign n1731 = n1530 & n1724 ;
  assign n1732 = n1730 & n1731 ;
  assign n1733 = n1593 & n1730 ;
  assign n1734 = n1530 & n1733 ;
  assign n1735 = ~n1732 & ~n1734 ;
  assign n1736 = n1498 & n1529 ;
  assign n1737 = n1724 & n1736 ;
  assign n1738 = n1720 & n1728 ;
  assign n1739 = n1737 & n1738 ;
  assign n1740 = n1688 & n1720 ;
  assign n1741 = n1657 & n1740 ;
  assign n1742 = n1594 & n1741 ;
  assign n1743 = n1731 & n1741 ;
  assign n1744 = ~n1561 & n1736 ;
  assign n1745 = n1730 & n1744 ;
  assign n1746 = ~n1743 & ~n1745 ;
  assign n1747 = ~n1742 & n1746 ;
  assign n1748 = ~n1739 & n1747 ;
  assign n1749 = n1735 & n1748 ;
  assign n1750 = n1727 & n1749 ;
  assign n1751 = ~n1625 & n1656 ;
  assign n1752 = ~n1592 & n1729 ;
  assign n1753 = n1751 & n1752 ;
  assign n1754 = n1744 & n1753 ;
  assign n1759 = n1592 & n1625 ;
  assign n1760 = n1656 & n1759 ;
  assign n1758 = n1529 & ~n1561 ;
  assign n1761 = n1740 & n1758 ;
  assign n1762 = n1760 & n1761 ;
  assign n1755 = n1740 & n1751 ;
  assign n1764 = ~n1498 & n1529 ;
  assign n1765 = n1593 & n1764 ;
  assign n1766 = n1755 & n1765 ;
  assign n1767 = ~n1762 & ~n1766 ;
  assign n1768 = ~n1754 & n1767 ;
  assign n1756 = ~n1689 & ~n1755 ;
  assign n1757 = n1737 & ~n1756 ;
  assign n1763 = n1723 & n1733 ;
  assign n1769 = ~n1757 & ~n1763 ;
  assign n1770 = n1768 & n1769 ;
  assign n1771 = ~n1750 & n1770 ;
  assign n1772 = n1444 & ~n1771 ;
  assign n1773 = ~\P2_InstQueueRd_Addr_reg[3]/NET0131  & \P2_InstQueueWr_Addr_reg[3]/NET0131  ;
  assign n1774 = ~\P2_InstQueueRd_Addr_reg[2]/NET0131  & \P2_InstQueueWr_Addr_reg[2]/NET0131  ;
  assign n1775 = \P2_InstQueueRd_Addr_reg[2]/NET0131  & ~\P2_InstQueueWr_Addr_reg[2]/NET0131  ;
  assign n1776 = ~\P2_InstQueueRd_Addr_reg[1]/NET0131  & \P2_InstQueueWr_Addr_reg[1]/NET0131  ;
  assign n1777 = \P2_InstQueueRd_Addr_reg[1]/NET0131  & ~\P2_InstQueueWr_Addr_reg[1]/NET0131  ;
  assign n1778 = \P2_InstQueueRd_Addr_reg[0]/NET0131  & ~\P2_InstQueueWr_Addr_reg[0]/NET0131  ;
  assign n1779 = ~n1777 & ~n1778 ;
  assign n1780 = ~n1776 & ~n1779 ;
  assign n1781 = ~n1775 & ~n1780 ;
  assign n1782 = ~n1774 & ~n1781 ;
  assign n1783 = n1773 & ~n1782 ;
  assign n1784 = \P2_InstQueueRd_Addr_reg[3]/NET0131  & ~\P2_InstQueueWr_Addr_reg[3]/NET0131  ;
  assign n1785 = ~n1782 & ~n1784 ;
  assign n1786 = ~n1773 & ~n1785 ;
  assign n1787 = ~n1774 & ~n1775 ;
  assign n1788 = n1780 & ~n1787 ;
  assign n1789 = ~n1780 & n1787 ;
  assign n1790 = ~n1788 & ~n1789 ;
  assign n1791 = ~n1786 & n1790 ;
  assign n1792 = ~n1783 & ~n1791 ;
  assign n1793 = ~n1776 & ~n1777 ;
  assign n1794 = ~\P2_InstQueueRd_Addr_reg[0]/NET0131  & \P2_InstQueueWr_Addr_reg[0]/NET0131  ;
  assign n1795 = ~n1778 & ~n1794 ;
  assign n1796 = n1793 & n1795 ;
  assign n1797 = ~n1783 & n1796 ;
  assign n1798 = ~n1792 & ~n1797 ;
  assign n1799 = ~\P2_InstQueueRd_Addr_reg[2]/NET0131  & ~n1798 ;
  assign n1800 = n1444 & n1798 ;
  assign n1801 = ~n1799 & ~n1800 ;
  assign n1802 = ~n1727 & n1801 ;
  assign n1835 = ~n1772 & ~n1802 ;
  assign n1806 = ~n1778 & ~n1793 ;
  assign n1807 = n1778 & n1793 ;
  assign n1808 = ~n1806 & ~n1807 ;
  assign n1809 = ~n1786 & ~n1808 ;
  assign n1810 = n1792 & ~n1809 ;
  assign n1813 = ~n1592 & n1745 ;
  assign n1814 = ~n1743 & ~n1813 ;
  assign n1822 = n1810 & ~n1814 ;
  assign n1803 = n1592 & n1745 ;
  assign n1804 = ~n1742 & ~n1803 ;
  assign n1805 = \ready12_reg/NET0131  & \ready21_reg/NET0131  ;
  assign n1811 = ~n1805 & ~n1810 ;
  assign n1812 = ~n1804 & ~n1811 ;
  assign n1815 = ~\P2_State_reg[0]/NET0131  & \P2_State_reg[1]/NET0131  ;
  assign n1816 = ~\P2_State_reg[2]/NET0131  & n1815 ;
  assign n1817 = ~\P2_State_reg[0]/NET0131  & ~\P2_State_reg[1]/NET0131  ;
  assign n1818 = \P2_State_reg[2]/NET0131  & n1817 ;
  assign n1819 = ~n1816 & ~n1818 ;
  assign n1820 = ~n1805 & ~n1819 ;
  assign n1821 = ~n1814 & ~n1820 ;
  assign n1823 = ~n1812 & ~n1821 ;
  assign n1824 = ~n1822 & n1823 ;
  assign n1825 = n1735 & n1824 ;
  assign n1826 = \P2_InstQueueRd_Addr_reg[2]/NET0131  & ~n1825 ;
  assign n1828 = ~n1814 & ~n1819 ;
  assign n1829 = n1804 & ~n1828 ;
  assign n1830 = n1811 & ~n1829 ;
  assign n1831 = ~n1739 & ~n1830 ;
  assign n1827 = \P2_InstQueueRd_Addr_reg[1]/NET0131  & \P2_InstQueueRd_Addr_reg[2]/NET0131  ;
  assign n1832 = ~\P2_InstQueueRd_Addr_reg[1]/NET0131  & ~\P2_InstQueueRd_Addr_reg[2]/NET0131  ;
  assign n1833 = ~n1827 & ~n1832 ;
  assign n1834 = ~n1831 & n1833 ;
  assign n1836 = ~n1826 & ~n1834 ;
  assign n1837 = n1835 & n1836 ;
  assign n1838 = \P2_InstQueueWr_Addr_reg[2]/NET0131  & n1837 ;
  assign n1860 = ~\P2_InstQueueRd_Addr_reg[3]/NET0131  & ~n1442 ;
  assign n1861 = ~n1456 & ~n1860 ;
  assign n1862 = ~n1771 & n1861 ;
  assign n1852 = ~n1814 & n1819 ;
  assign n1853 = ~n1747 & n1810 ;
  assign n1854 = ~n1852 & ~n1853 ;
  assign n1839 = ~\P2_InstQueueRd_Addr_reg[3]/NET0131  & ~n1827 ;
  assign n1840 = \P2_InstQueueRd_Addr_reg[3]/NET0131  & n1827 ;
  assign n1841 = ~n1839 & ~n1840 ;
  assign n1842 = ~n1805 & n1841 ;
  assign n1843 = \P2_InstQueueRd_Addr_reg[3]/NET0131  & n1805 ;
  assign n1844 = ~n1842 & ~n1843 ;
  assign n1855 = ~n1814 & ~n1844 ;
  assign n1856 = n1735 & ~n1855 ;
  assign n1857 = n1854 & n1856 ;
  assign n1858 = \P2_InstQueueRd_Addr_reg[3]/NET0131  & ~n1857 ;
  assign n1845 = ~n1810 & ~n1829 ;
  assign n1846 = ~n1844 & n1845 ;
  assign n1847 = ~n1443 & n1798 ;
  assign n1849 = \P2_InstQueueRd_Addr_reg[3]/NET0131  & n1847 ;
  assign n1848 = ~\P2_InstQueueRd_Addr_reg[3]/NET0131  & ~n1847 ;
  assign n1850 = ~n1727 & ~n1848 ;
  assign n1851 = ~n1849 & n1850 ;
  assign n1859 = n1739 & n1841 ;
  assign n1863 = ~n1851 & ~n1859 ;
  assign n1864 = ~n1846 & n1863 ;
  assign n1865 = ~n1858 & n1864 ;
  assign n1866 = ~n1862 & n1865 ;
  assign n1867 = \P2_InstQueueWr_Addr_reg[3]/NET0131  & n1866 ;
  assign n1868 = ~n1838 & ~n1867 ;
  assign n1870 = ~n1727 & n1798 ;
  assign n1871 = n1771 & ~n1870 ;
  assign n1908 = ~\P2_InstQueueRd_Addr_reg[0]/NET0131  & n1871 ;
  assign n1876 = n1726 & ~n1798 ;
  assign n1877 = n1722 & ~n1798 ;
  assign n1878 = ~n1876 & ~n1877 ;
  assign n1909 = \P2_InstQueueRd_Addr_reg[0]/NET0131  & n1878 ;
  assign n1910 = n1749 & n1909 ;
  assign n1911 = ~n1908 & ~n1910 ;
  assign n1912 = \P2_InstQueueWr_Addr_reg[0]/NET0131  & ~n1911 ;
  assign n1872 = ~n1445 & ~n1458 ;
  assign n1873 = ~n1871 & ~n1872 ;
  assign n1869 = ~\P2_InstQueueRd_Addr_reg[1]/NET0131  & ~n1831 ;
  assign n1874 = n1811 & ~n1852 ;
  assign n1875 = ~n1747 & ~n1874 ;
  assign n1879 = n1735 & n1878 ;
  assign n1880 = ~n1875 & n1879 ;
  assign n1881 = \P2_InstQueueRd_Addr_reg[1]/NET0131  & ~n1880 ;
  assign n1882 = ~n1869 & ~n1881 ;
  assign n1883 = ~n1873 & n1882 ;
  assign n1913 = \P2_InstQueueWr_Addr_reg[1]/NET0131  & n1883 ;
  assign n1914 = ~n1912 & ~n1913 ;
  assign n1915 = n1868 & n1914 ;
  assign n1884 = ~\P2_InstQueueWr_Addr_reg[1]/NET0131  & ~n1883 ;
  assign n1885 = ~\P2_InstQueueWr_Addr_reg[2]/NET0131  & ~n1837 ;
  assign n1886 = ~n1884 & ~n1885 ;
  assign n1887 = n1868 & ~n1886 ;
  assign n1888 = \P2_InstQueueWr_Addr_reg[3]/NET0131  & n1837 ;
  assign n1889 = ~n1866 & ~n1888 ;
  assign n1891 = ~n1804 & ~n1810 ;
  assign n1892 = n1805 & n1891 ;
  assign n1893 = ~n1810 & n1821 ;
  assign n1894 = ~n1892 & ~n1893 ;
  assign n1895 = \P2_Flush_reg/NET0131  & ~n1894 ;
  assign n1890 = n1732 & n1798 ;
  assign n1896 = ~n1795 & n1809 ;
  assign n1897 = n1792 & ~n1896 ;
  assign n1898 = n1734 & ~n1897 ;
  assign n1899 = ~n1890 & ~n1898 ;
  assign n1900 = ~n1895 & n1899 ;
  assign n1904 = ~\P2_More_reg/NET0131  & ~n1810 ;
  assign n1905 = ~n1824 & ~n1904 ;
  assign n1901 = n1734 & n1897 ;
  assign n1902 = n1732 & ~n1798 ;
  assign n1903 = n1878 & ~n1902 ;
  assign n1906 = ~n1901 & n1903 ;
  assign n1907 = ~n1905 & n1906 ;
  assign n1916 = n1900 & n1907 ;
  assign n1917 = ~n1889 & n1916 ;
  assign n1918 = ~n1887 & n1917 ;
  assign n1919 = ~n1915 & n1918 ;
  assign n1920 = ~\P2_DataWidth_reg[1]/NET0131  & ~n1805 ;
  assign n1921 = ~n1810 & ~n1819 ;
  assign n1922 = n1743 & n1921 ;
  assign n1923 = n1920 & n1922 ;
  assign n1924 = n1919 & ~n1923 ;
  assign n1925 = \P2_State2_reg[0]/NET0131  & ~\P2_State2_reg[3]/NET0131  ;
  assign n1926 = ~\P2_State2_reg[1]/NET0131  & \P2_State2_reg[2]/NET0131  ;
  assign n1927 = n1925 & n1926 ;
  assign n1928 = ~n1924 & n1927 ;
  assign n1929 = \P2_State2_reg[1]/NET0131  & ~\P2_State2_reg[2]/NET0131  ;
  assign n1930 = ~\P2_State2_reg[3]/NET0131  & n1929 ;
  assign n1931 = ~\P2_State2_reg[0]/NET0131  & n1930 ;
  assign n1932 = ~\P2_DataWidth_reg[1]/NET0131  & n1931 ;
  assign n1933 = ~\P2_State2_reg[2]/NET0131  & n1925 ;
  assign n1934 = ~\P2_State2_reg[1]/NET0131  & n1933 ;
  assign n1935 = ~\P2_State2_reg[0]/NET0131  & ~\P2_State2_reg[3]/NET0131  ;
  assign n1936 = \P2_State2_reg[2]/NET0131  & n1935 ;
  assign n1937 = ~n1933 & ~n1936 ;
  assign n1938 = n1805 & ~n1937 ;
  assign n1939 = ~n1934 & ~n1938 ;
  assign n1940 = ~\P2_State2_reg[1]/NET0131  & n1805 ;
  assign n1941 = ~n1939 & ~n1940 ;
  assign n1942 = ~n1932 & ~n1941 ;
  assign n1943 = ~n1928 & n1942 ;
  assign n1951 = ~\P1_InstQueueRd_Addr_reg[0]/NET0131  & ~\P1_InstQueueRd_Addr_reg[1]/NET0131  ;
  assign n1957 = ~\P1_InstQueueRd_Addr_reg[2]/NET0131  & ~\P1_InstQueueRd_Addr_reg[3]/NET0131  ;
  assign n1958 = n1951 & n1957 ;
  assign n1959 = \P1_InstQueue_reg[0][2]/NET0131  & n1958 ;
  assign n1960 = \P1_InstQueueRd_Addr_reg[2]/NET0131  & ~\P1_InstQueueRd_Addr_reg[3]/NET0131  ;
  assign n1961 = n1951 & n1960 ;
  assign n1962 = \P1_InstQueue_reg[4][2]/NET0131  & n1961 ;
  assign n1986 = ~n1959 & ~n1962 ;
  assign n1963 = \P1_InstQueueRd_Addr_reg[0]/NET0131  & ~\P1_InstQueueRd_Addr_reg[1]/NET0131  ;
  assign n1964 = n1960 & n1963 ;
  assign n1965 = \P1_InstQueue_reg[5][2]/NET0131  & n1964 ;
  assign n1966 = n1957 & n1963 ;
  assign n1967 = \P1_InstQueue_reg[1][2]/NET0131  & n1966 ;
  assign n1987 = ~n1965 & ~n1967 ;
  assign n1994 = n1986 & n1987 ;
  assign n1944 = ~\P1_InstQueueRd_Addr_reg[0]/NET0131  & \P1_InstQueueRd_Addr_reg[1]/NET0131  ;
  assign n1945 = ~\P1_InstQueueRd_Addr_reg[2]/NET0131  & \P1_InstQueueRd_Addr_reg[3]/NET0131  ;
  assign n1946 = n1944 & n1945 ;
  assign n1947 = \P1_InstQueue_reg[10][2]/NET0131  & n1946 ;
  assign n1948 = \P1_InstQueueRd_Addr_reg[0]/NET0131  & \P1_InstQueueRd_Addr_reg[1]/NET0131  ;
  assign n1949 = n1945 & n1948 ;
  assign n1950 = \P1_InstQueue_reg[11][2]/NET0131  & n1949 ;
  assign n1984 = ~n1947 & ~n1950 ;
  assign n1952 = \P1_InstQueueRd_Addr_reg[2]/NET0131  & \P1_InstQueueRd_Addr_reg[3]/NET0131  ;
  assign n1953 = n1951 & n1952 ;
  assign n1954 = \P1_InstQueue_reg[12][2]/NET0131  & n1953 ;
  assign n1955 = n1944 & n1952 ;
  assign n1956 = \P1_InstQueue_reg[14][2]/NET0131  & n1955 ;
  assign n1985 = ~n1954 & ~n1956 ;
  assign n1995 = n1984 & n1985 ;
  assign n1996 = n1994 & n1995 ;
  assign n1976 = n1948 & n1957 ;
  assign n1977 = \P1_InstQueue_reg[3][2]/NET0131  & n1976 ;
  assign n1978 = n1945 & n1963 ;
  assign n1979 = \P1_InstQueue_reg[9][2]/NET0131  & n1978 ;
  assign n1990 = ~n1977 & ~n1979 ;
  assign n1980 = n1952 & n1963 ;
  assign n1981 = \P1_InstQueue_reg[13][2]/NET0131  & n1980 ;
  assign n1982 = n1948 & n1952 ;
  assign n1983 = \P1_InstQueue_reg[15][2]/NET0131  & n1982 ;
  assign n1991 = ~n1981 & ~n1983 ;
  assign n1992 = n1990 & n1991 ;
  assign n1968 = n1948 & n1960 ;
  assign n1969 = \P1_InstQueue_reg[7][2]/NET0131  & n1968 ;
  assign n1970 = n1944 & n1957 ;
  assign n1971 = \P1_InstQueue_reg[2][2]/NET0131  & n1970 ;
  assign n1988 = ~n1969 & ~n1971 ;
  assign n1972 = n1944 & n1960 ;
  assign n1973 = \P1_InstQueue_reg[6][2]/NET0131  & n1972 ;
  assign n1974 = n1945 & n1951 ;
  assign n1975 = \P1_InstQueue_reg[8][2]/NET0131  & n1974 ;
  assign n1989 = ~n1973 & ~n1975 ;
  assign n1993 = n1988 & n1989 ;
  assign n1997 = n1992 & n1993 ;
  assign n1998 = n1996 & n1997 ;
  assign n2003 = \P1_InstQueue_reg[11][1]/NET0131  & n1949 ;
  assign n2004 = \P1_InstQueue_reg[9][1]/NET0131  & n1978 ;
  assign n2017 = ~n2003 & ~n2004 ;
  assign n2005 = \P1_InstQueue_reg[15][1]/NET0131  & n1982 ;
  assign n2006 = \P1_InstQueue_reg[3][1]/NET0131  & n1976 ;
  assign n2018 = ~n2005 & ~n2006 ;
  assign n2025 = n2017 & n2018 ;
  assign n1999 = \P1_InstQueue_reg[14][1]/NET0131  & n1955 ;
  assign n2000 = \P1_InstQueue_reg[0][1]/NET0131  & n1958 ;
  assign n2015 = ~n1999 & ~n2000 ;
  assign n2001 = \P1_InstQueue_reg[6][1]/NET0131  & n1972 ;
  assign n2002 = \P1_InstQueue_reg[12][1]/NET0131  & n1953 ;
  assign n2016 = ~n2001 & ~n2002 ;
  assign n2026 = n2015 & n2016 ;
  assign n2027 = n2025 & n2026 ;
  assign n2011 = \P1_InstQueue_reg[1][1]/NET0131  & n1966 ;
  assign n2012 = \P1_InstQueue_reg[2][1]/NET0131  & n1970 ;
  assign n2021 = ~n2011 & ~n2012 ;
  assign n2013 = \P1_InstQueue_reg[8][1]/NET0131  & n1974 ;
  assign n2014 = \P1_InstQueue_reg[7][1]/NET0131  & n1968 ;
  assign n2022 = ~n2013 & ~n2014 ;
  assign n2023 = n2021 & n2022 ;
  assign n2007 = \P1_InstQueue_reg[10][1]/NET0131  & n1946 ;
  assign n2008 = \P1_InstQueue_reg[5][1]/NET0131  & n1964 ;
  assign n2019 = ~n2007 & ~n2008 ;
  assign n2009 = \P1_InstQueue_reg[13][1]/NET0131  & n1980 ;
  assign n2010 = \P1_InstQueue_reg[4][1]/NET0131  & n1961 ;
  assign n2020 = ~n2009 & ~n2010 ;
  assign n2024 = n2019 & n2020 ;
  assign n2028 = n2023 & n2024 ;
  assign n2029 = n2027 & n2028 ;
  assign n2030 = n1998 & ~n2029 ;
  assign n2035 = \P1_InstQueue_reg[5][3]/NET0131  & n1964 ;
  assign n2036 = \P1_InstQueue_reg[4][3]/NET0131  & n1961 ;
  assign n2049 = ~n2035 & ~n2036 ;
  assign n2037 = \P1_InstQueue_reg[15][3]/NET0131  & n1982 ;
  assign n2038 = \P1_InstQueue_reg[13][3]/NET0131  & n1980 ;
  assign n2050 = ~n2037 & ~n2038 ;
  assign n2057 = n2049 & n2050 ;
  assign n2031 = \P1_InstQueue_reg[14][3]/NET0131  & n1955 ;
  assign n2032 = \P1_InstQueue_reg[7][3]/NET0131  & n1968 ;
  assign n2047 = ~n2031 & ~n2032 ;
  assign n2033 = \P1_InstQueue_reg[9][3]/NET0131  & n1978 ;
  assign n2034 = \P1_InstQueue_reg[8][3]/NET0131  & n1974 ;
  assign n2048 = ~n2033 & ~n2034 ;
  assign n2058 = n2047 & n2048 ;
  assign n2059 = n2057 & n2058 ;
  assign n2043 = \P1_InstQueue_reg[0][3]/NET0131  & n1958 ;
  assign n2044 = \P1_InstQueue_reg[11][3]/NET0131  & n1949 ;
  assign n2053 = ~n2043 & ~n2044 ;
  assign n2045 = \P1_InstQueue_reg[2][3]/NET0131  & n1970 ;
  assign n2046 = \P1_InstQueue_reg[12][3]/NET0131  & n1953 ;
  assign n2054 = ~n2045 & ~n2046 ;
  assign n2055 = n2053 & n2054 ;
  assign n2039 = \P1_InstQueue_reg[10][3]/NET0131  & n1946 ;
  assign n2040 = \P1_InstQueue_reg[3][3]/NET0131  & n1976 ;
  assign n2051 = ~n2039 & ~n2040 ;
  assign n2041 = \P1_InstQueue_reg[6][3]/NET0131  & n1972 ;
  assign n2042 = \P1_InstQueue_reg[1][3]/NET0131  & n1966 ;
  assign n2052 = ~n2041 & ~n2042 ;
  assign n2056 = n2051 & n2052 ;
  assign n2060 = n2055 & n2056 ;
  assign n2061 = n2059 & n2060 ;
  assign n2066 = \P1_InstQueue_reg[9][0]/NET0131  & n1978 ;
  assign n2067 = \P1_InstQueue_reg[7][0]/NET0131  & n1968 ;
  assign n2080 = ~n2066 & ~n2067 ;
  assign n2068 = \P1_InstQueue_reg[14][0]/NET0131  & n1955 ;
  assign n2069 = \P1_InstQueue_reg[4][0]/NET0131  & n1961 ;
  assign n2081 = ~n2068 & ~n2069 ;
  assign n2088 = n2080 & n2081 ;
  assign n2062 = \P1_InstQueue_reg[10][0]/NET0131  & n1946 ;
  assign n2063 = \P1_InstQueue_reg[5][0]/NET0131  & n1964 ;
  assign n2078 = ~n2062 & ~n2063 ;
  assign n2064 = \P1_InstQueue_reg[11][0]/NET0131  & n1949 ;
  assign n2065 = \P1_InstQueue_reg[2][0]/NET0131  & n1970 ;
  assign n2079 = ~n2064 & ~n2065 ;
  assign n2089 = n2078 & n2079 ;
  assign n2090 = n2088 & n2089 ;
  assign n2074 = \P1_InstQueue_reg[12][0]/NET0131  & n1953 ;
  assign n2075 = \P1_InstQueue_reg[1][0]/NET0131  & n1966 ;
  assign n2084 = ~n2074 & ~n2075 ;
  assign n2076 = \P1_InstQueue_reg[13][0]/NET0131  & n1980 ;
  assign n2077 = \P1_InstQueue_reg[0][0]/NET0131  & n1958 ;
  assign n2085 = ~n2076 & ~n2077 ;
  assign n2086 = n2084 & n2085 ;
  assign n2070 = \P1_InstQueue_reg[8][0]/NET0131  & n1974 ;
  assign n2071 = \P1_InstQueue_reg[6][0]/NET0131  & n1972 ;
  assign n2082 = ~n2070 & ~n2071 ;
  assign n2072 = \P1_InstQueue_reg[15][0]/NET0131  & n1982 ;
  assign n2073 = \P1_InstQueue_reg[3][0]/NET0131  & n1976 ;
  assign n2083 = ~n2072 & ~n2073 ;
  assign n2087 = n2082 & n2083 ;
  assign n2091 = n2086 & n2087 ;
  assign n2092 = n2090 & n2091 ;
  assign n2093 = ~n2061 & ~n2092 ;
  assign n2094 = n2030 & n2093 ;
  assign n2099 = \P1_InstQueue_reg[0][6]/NET0131  & n1958 ;
  assign n2100 = \P1_InstQueue_reg[4][6]/NET0131  & n1961 ;
  assign n2113 = ~n2099 & ~n2100 ;
  assign n2101 = \P1_InstQueue_reg[5][6]/NET0131  & n1964 ;
  assign n2102 = \P1_InstQueue_reg[1][6]/NET0131  & n1966 ;
  assign n2114 = ~n2101 & ~n2102 ;
  assign n2121 = n2113 & n2114 ;
  assign n2095 = \P1_InstQueue_reg[10][6]/NET0131  & n1946 ;
  assign n2096 = \P1_InstQueue_reg[11][6]/NET0131  & n1949 ;
  assign n2111 = ~n2095 & ~n2096 ;
  assign n2097 = \P1_InstQueue_reg[12][6]/NET0131  & n1953 ;
  assign n2098 = \P1_InstQueue_reg[14][6]/NET0131  & n1955 ;
  assign n2112 = ~n2097 & ~n2098 ;
  assign n2122 = n2111 & n2112 ;
  assign n2123 = n2121 & n2122 ;
  assign n2107 = \P1_InstQueue_reg[3][6]/NET0131  & n1976 ;
  assign n2108 = \P1_InstQueue_reg[9][6]/NET0131  & n1978 ;
  assign n2117 = ~n2107 & ~n2108 ;
  assign n2109 = \P1_InstQueue_reg[13][6]/NET0131  & n1980 ;
  assign n2110 = \P1_InstQueue_reg[15][6]/NET0131  & n1982 ;
  assign n2118 = ~n2109 & ~n2110 ;
  assign n2119 = n2117 & n2118 ;
  assign n2103 = \P1_InstQueue_reg[7][6]/NET0131  & n1968 ;
  assign n2104 = \P1_InstQueue_reg[2][6]/NET0131  & n1970 ;
  assign n2115 = ~n2103 & ~n2104 ;
  assign n2105 = \P1_InstQueue_reg[6][6]/NET0131  & n1972 ;
  assign n2106 = \P1_InstQueue_reg[8][6]/NET0131  & n1974 ;
  assign n2116 = ~n2105 & ~n2106 ;
  assign n2120 = n2115 & n2116 ;
  assign n2124 = n2119 & n2120 ;
  assign n2125 = n2123 & n2124 ;
  assign n2130 = \P1_InstQueue_reg[0][7]/NET0131  & n1958 ;
  assign n2131 = \P1_InstQueue_reg[4][7]/NET0131  & n1961 ;
  assign n2144 = ~n2130 & ~n2131 ;
  assign n2132 = \P1_InstQueue_reg[5][7]/NET0131  & n1964 ;
  assign n2133 = \P1_InstQueue_reg[1][7]/NET0131  & n1966 ;
  assign n2145 = ~n2132 & ~n2133 ;
  assign n2152 = n2144 & n2145 ;
  assign n2126 = \P1_InstQueue_reg[10][7]/NET0131  & n1946 ;
  assign n2127 = \P1_InstQueue_reg[11][7]/NET0131  & n1949 ;
  assign n2142 = ~n2126 & ~n2127 ;
  assign n2128 = \P1_InstQueue_reg[12][7]/NET0131  & n1953 ;
  assign n2129 = \P1_InstQueue_reg[14][7]/NET0131  & n1955 ;
  assign n2143 = ~n2128 & ~n2129 ;
  assign n2153 = n2142 & n2143 ;
  assign n2154 = n2152 & n2153 ;
  assign n2138 = \P1_InstQueue_reg[3][7]/NET0131  & n1976 ;
  assign n2139 = \P1_InstQueue_reg[9][7]/NET0131  & n1978 ;
  assign n2148 = ~n2138 & ~n2139 ;
  assign n2140 = \P1_InstQueue_reg[13][7]/NET0131  & n1980 ;
  assign n2141 = \P1_InstQueue_reg[15][7]/NET0131  & n1982 ;
  assign n2149 = ~n2140 & ~n2141 ;
  assign n2150 = n2148 & n2149 ;
  assign n2134 = \P1_InstQueue_reg[7][7]/NET0131  & n1968 ;
  assign n2135 = \P1_InstQueue_reg[2][7]/NET0131  & n1970 ;
  assign n2146 = ~n2134 & ~n2135 ;
  assign n2136 = \P1_InstQueue_reg[6][7]/NET0131  & n1972 ;
  assign n2137 = \P1_InstQueue_reg[8][7]/NET0131  & n1974 ;
  assign n2147 = ~n2136 & ~n2137 ;
  assign n2151 = n2146 & n2147 ;
  assign n2155 = n2150 & n2151 ;
  assign n2156 = n2154 & n2155 ;
  assign n2157 = n2125 & ~n2156 ;
  assign n2162 = \P1_InstQueue_reg[7][4]/NET0131  & n1968 ;
  assign n2163 = \P1_InstQueue_reg[0][4]/NET0131  & n1958 ;
  assign n2176 = ~n2162 & ~n2163 ;
  assign n2164 = \P1_InstQueue_reg[14][4]/NET0131  & n1955 ;
  assign n2165 = \P1_InstQueue_reg[1][4]/NET0131  & n1966 ;
  assign n2177 = ~n2164 & ~n2165 ;
  assign n2184 = n2176 & n2177 ;
  assign n2158 = \P1_InstQueue_reg[10][4]/NET0131  & n1946 ;
  assign n2159 = \P1_InstQueue_reg[5][4]/NET0131  & n1964 ;
  assign n2174 = ~n2158 & ~n2159 ;
  assign n2160 = \P1_InstQueue_reg[11][4]/NET0131  & n1949 ;
  assign n2161 = \P1_InstQueue_reg[12][4]/NET0131  & n1953 ;
  assign n2175 = ~n2160 & ~n2161 ;
  assign n2185 = n2174 & n2175 ;
  assign n2186 = n2184 & n2185 ;
  assign n2170 = \P1_InstQueue_reg[3][4]/NET0131  & n1976 ;
  assign n2171 = \P1_InstQueue_reg[4][4]/NET0131  & n1961 ;
  assign n2180 = ~n2170 & ~n2171 ;
  assign n2172 = \P1_InstQueue_reg[13][4]/NET0131  & n1980 ;
  assign n2173 = \P1_InstQueue_reg[9][4]/NET0131  & n1978 ;
  assign n2181 = ~n2172 & ~n2173 ;
  assign n2182 = n2180 & n2181 ;
  assign n2166 = \P1_InstQueue_reg[15][4]/NET0131  & n1982 ;
  assign n2167 = \P1_InstQueue_reg[6][4]/NET0131  & n1972 ;
  assign n2178 = ~n2166 & ~n2167 ;
  assign n2168 = \P1_InstQueue_reg[2][4]/NET0131  & n1970 ;
  assign n2169 = \P1_InstQueue_reg[8][4]/NET0131  & n1974 ;
  assign n2179 = ~n2168 & ~n2169 ;
  assign n2183 = n2178 & n2179 ;
  assign n2187 = n2182 & n2183 ;
  assign n2188 = n2186 & n2187 ;
  assign n2193 = \P1_InstQueue_reg[7][5]/NET0131  & n1968 ;
  assign n2194 = \P1_InstQueue_reg[0][5]/NET0131  & n1958 ;
  assign n2207 = ~n2193 & ~n2194 ;
  assign n2195 = \P1_InstQueue_reg[14][5]/NET0131  & n1955 ;
  assign n2196 = \P1_InstQueue_reg[1][5]/NET0131  & n1966 ;
  assign n2208 = ~n2195 & ~n2196 ;
  assign n2215 = n2207 & n2208 ;
  assign n2189 = \P1_InstQueue_reg[10][5]/NET0131  & n1946 ;
  assign n2190 = \P1_InstQueue_reg[5][5]/NET0131  & n1964 ;
  assign n2205 = ~n2189 & ~n2190 ;
  assign n2191 = \P1_InstQueue_reg[11][5]/NET0131  & n1949 ;
  assign n2192 = \P1_InstQueue_reg[12][5]/NET0131  & n1953 ;
  assign n2206 = ~n2191 & ~n2192 ;
  assign n2216 = n2205 & n2206 ;
  assign n2217 = n2215 & n2216 ;
  assign n2201 = \P1_InstQueue_reg[3][5]/NET0131  & n1976 ;
  assign n2202 = \P1_InstQueue_reg[9][5]/NET0131  & n1978 ;
  assign n2211 = ~n2201 & ~n2202 ;
  assign n2203 = \P1_InstQueue_reg[13][5]/NET0131  & n1980 ;
  assign n2204 = \P1_InstQueue_reg[4][5]/NET0131  & n1961 ;
  assign n2212 = ~n2203 & ~n2204 ;
  assign n2213 = n2211 & n2212 ;
  assign n2197 = \P1_InstQueue_reg[15][5]/NET0131  & n1982 ;
  assign n2198 = \P1_InstQueue_reg[6][5]/NET0131  & n1972 ;
  assign n2209 = ~n2197 & ~n2198 ;
  assign n2199 = \P1_InstQueue_reg[2][5]/NET0131  & n1970 ;
  assign n2200 = \P1_InstQueue_reg[8][5]/NET0131  & n1974 ;
  assign n2210 = ~n2199 & ~n2200 ;
  assign n2214 = n2209 & n2210 ;
  assign n2218 = n2213 & n2214 ;
  assign n2219 = n2217 & n2218 ;
  assign n2220 = n2188 & n2219 ;
  assign n2221 = n2157 & n2220 ;
  assign n2222 = n2094 & n2221 ;
  assign n2223 = n1998 & n2029 ;
  assign n2224 = n2093 & n2223 ;
  assign n2225 = n2221 & n2224 ;
  assign n2226 = ~n2125 & ~n2156 ;
  assign n2227 = n2188 & ~n2219 ;
  assign n2228 = n2226 & n2227 ;
  assign n2229 = ~n1998 & n2061 ;
  assign n2230 = n2092 & n2229 ;
  assign n2231 = n2228 & n2230 ;
  assign n2232 = ~n2225 & ~n2231 ;
  assign n2233 = ~n2222 & n2232 ;
  assign n2234 = n2092 & n2223 ;
  assign n2235 = n2061 & n2234 ;
  assign n2236 = n2219 & n2226 ;
  assign n2237 = n2235 & n2236 ;
  assign n2238 = n2233 & ~n2237 ;
  assign n2243 = n2224 & n2228 ;
  assign n2244 = n2094 & n2228 ;
  assign n2245 = ~n2243 & ~n2244 ;
  assign n2239 = n2157 & ~n2188 ;
  assign n2240 = ~n2219 & n2239 ;
  assign n2241 = n2234 & n2240 ;
  assign n2242 = n2094 & n2240 ;
  assign n2246 = ~n2241 & ~n2242 ;
  assign n2247 = n2245 & n2246 ;
  assign n2248 = n2238 & n2247 ;
  assign n2252 = n2235 & n2239 ;
  assign n2249 = ~n2061 & n2092 ;
  assign n2250 = n2030 & n2249 ;
  assign n2251 = n2228 & n2250 ;
  assign n2253 = n2061 & n2220 ;
  assign n2254 = ~n1998 & n2029 ;
  assign n2255 = n2125 & n2156 ;
  assign n2256 = n2254 & n2255 ;
  assign n2257 = n2253 & n2256 ;
  assign n2266 = ~n2251 & ~n2257 ;
  assign n2267 = ~n2252 & n2266 ;
  assign n2258 = ~n2125 & n2156 ;
  assign n2263 = ~n2029 & n2227 ;
  assign n2264 = n2258 & n2263 ;
  assign n2265 = n2230 & n2264 ;
  assign n2259 = n2253 & n2258 ;
  assign n2260 = n2234 & n2259 ;
  assign n2261 = n2030 & ~n2092 ;
  assign n2262 = n2259 & n2261 ;
  assign n2268 = ~n2260 & ~n2262 ;
  assign n2269 = ~n2265 & n2268 ;
  assign n2270 = n2267 & n2269 ;
  assign n2271 = ~n2248 & n2270 ;
  assign n2331 = ~n2061 & n2241 ;
  assign n2332 = ~n2242 & ~n2331 ;
  assign n2276 = ~\P1_InstQueueRd_Addr_reg[3]/NET0131  & \P1_InstQueueWr_Addr_reg[3]/NET0131  ;
  assign n2277 = ~\P1_InstQueueRd_Addr_reg[2]/NET0131  & \P1_InstQueueWr_Addr_reg[2]/NET0131  ;
  assign n2278 = \P1_InstQueueRd_Addr_reg[2]/NET0131  & ~\P1_InstQueueWr_Addr_reg[2]/NET0131  ;
  assign n2279 = ~\P1_InstQueueRd_Addr_reg[1]/NET0131  & \P1_InstQueueWr_Addr_reg[1]/NET0131  ;
  assign n2280 = \P1_InstQueueRd_Addr_reg[1]/NET0131  & ~\P1_InstQueueWr_Addr_reg[1]/NET0131  ;
  assign n2281 = \P1_InstQueueRd_Addr_reg[0]/NET0131  & ~\P1_InstQueueWr_Addr_reg[0]/NET0131  ;
  assign n2282 = ~n2280 & ~n2281 ;
  assign n2283 = ~n2279 & ~n2282 ;
  assign n2284 = ~n2278 & ~n2283 ;
  assign n2285 = ~n2277 & ~n2284 ;
  assign n2286 = n2276 & ~n2285 ;
  assign n2287 = \P1_InstQueueRd_Addr_reg[3]/NET0131  & ~\P1_InstQueueWr_Addr_reg[3]/NET0131  ;
  assign n2288 = ~n2285 & ~n2287 ;
  assign n2289 = ~n2276 & ~n2288 ;
  assign n2290 = ~n2277 & ~n2278 ;
  assign n2291 = n2283 & ~n2290 ;
  assign n2292 = ~n2283 & n2290 ;
  assign n2293 = ~n2291 & ~n2292 ;
  assign n2294 = ~n2289 & n2293 ;
  assign n2295 = ~n2286 & ~n2294 ;
  assign n2296 = ~n2279 & ~n2280 ;
  assign n2333 = ~\P1_InstQueueRd_Addr_reg[0]/NET0131  & \P1_InstQueueWr_Addr_reg[0]/NET0131  ;
  assign n2334 = ~n2281 & ~n2333 ;
  assign n2335 = n2296 & n2334 ;
  assign n2336 = ~n2286 & n2335 ;
  assign n2337 = ~n2295 & ~n2336 ;
  assign n2397 = ~n2332 & n2337 ;
  assign n2398 = n2271 & ~n2397 ;
  assign n2399 = ~n1944 & ~n1963 ;
  assign n2400 = ~n2398 & ~n2399 ;
  assign n2297 = ~n2281 & ~n2296 ;
  assign n2298 = n2281 & n2296 ;
  assign n2299 = ~n2297 & ~n2298 ;
  assign n2300 = ~n2289 & ~n2299 ;
  assign n2301 = n2295 & ~n2300 ;
  assign n2302 = n2029 & n2231 ;
  assign n2303 = ~n2222 & ~n2302 ;
  assign n2304 = ~n2301 & ~n2303 ;
  assign n2305 = ~n2029 & n2231 ;
  assign n2306 = ~n2225 & ~n2305 ;
  assign n2307 = ~\P1_State_reg[0]/NET0131  & \P1_State_reg[1]/NET0131  ;
  assign n2308 = ~\P1_State_reg[2]/NET0131  & n2307 ;
  assign n2309 = ~\P1_State_reg[0]/NET0131  & ~\P1_State_reg[1]/NET0131  ;
  assign n2310 = \P1_State_reg[2]/NET0131  & n2309 ;
  assign n2311 = ~n2308 & ~n2310 ;
  assign n2312 = ~n2301 & ~n2311 ;
  assign n2313 = ~n2306 & n2312 ;
  assign n2314 = ~n2304 & ~n2313 ;
  assign n2317 = \ready11_reg/NET0131  & \ready1_pad  ;
  assign n2401 = ~n2314 & ~n2317 ;
  assign n2402 = ~n2237 & ~n2401 ;
  assign n2403 = ~\P1_InstQueueRd_Addr_reg[1]/NET0131  & n2402 ;
  assign n2370 = n2242 & ~n2337 ;
  assign n2371 = n2331 & ~n2337 ;
  assign n2372 = ~n2370 & ~n2371 ;
  assign n2404 = n2245 & n2372 ;
  assign n2326 = ~n2306 & n2311 ;
  assign n2377 = ~n2301 & ~n2317 ;
  assign n2378 = ~n2326 & n2377 ;
  assign n2379 = ~n2233 & ~n2378 ;
  assign n2405 = \P1_InstQueueRd_Addr_reg[1]/NET0131  & ~n2379 ;
  assign n2406 = n2404 & n2405 ;
  assign n2407 = ~n2403 & ~n2406 ;
  assign n2408 = ~n2400 & ~n2407 ;
  assign n2410 = ~\P1_InstQueueWr_Addr_reg[1]/NET0131  & ~n2408 ;
  assign n2411 = ~\P1_InstQueueRd_Addr_reg[0]/NET0131  & n2398 ;
  assign n2412 = \P1_InstQueueRd_Addr_reg[0]/NET0131  & n2238 ;
  assign n2413 = n2404 & n2412 ;
  assign n2414 = ~n2411 & ~n2413 ;
  assign n2415 = \P1_InstQueueWr_Addr_reg[0]/NET0131  & ~n2414 ;
  assign n2416 = ~n2410 & n2415 ;
  assign n2409 = \P1_InstQueueWr_Addr_reg[1]/NET0131  & n2408 ;
  assign n2325 = ~n2233 & n2301 ;
  assign n2327 = n2245 & ~n2325 ;
  assign n2328 = ~n2326 & n2327 ;
  assign n2272 = ~\P1_InstQueueRd_Addr_reg[2]/NET0131  & ~n1948 ;
  assign n2350 = ~n2272 & n2337 ;
  assign n2351 = ~n2332 & ~n2350 ;
  assign n2352 = n2328 & ~n2351 ;
  assign n2353 = \P1_InstQueueRd_Addr_reg[3]/NET0131  & ~n2352 ;
  assign n2273 = \P1_InstQueueRd_Addr_reg[2]/NET0131  & n1948 ;
  assign n2347 = \P1_InstQueueRd_Addr_reg[3]/NET0131  & ~n2273 ;
  assign n2348 = ~n1968 & ~n2347 ;
  assign n2349 = ~n2271 & ~n2348 ;
  assign n2318 = \P1_InstQueueRd_Addr_reg[1]/NET0131  & \P1_InstQueueRd_Addr_reg[2]/NET0131  ;
  assign n2354 = ~\P1_InstQueueRd_Addr_reg[3]/NET0131  & ~n2318 ;
  assign n2355 = \P1_InstQueueRd_Addr_reg[3]/NET0131  & n2318 ;
  assign n2356 = ~n2354 & ~n2355 ;
  assign n2360 = ~n2317 & ~n2356 ;
  assign n2361 = ~\P1_InstQueueRd_Addr_reg[3]/NET0131  & n2317 ;
  assign n2362 = ~n2360 & ~n2361 ;
  assign n2363 = ~n2314 & n2362 ;
  assign n2357 = n2237 & n2356 ;
  assign n2358 = ~\P1_InstQueueRd_Addr_reg[3]/NET0131  & n2350 ;
  assign n2359 = ~n2332 & n2358 ;
  assign n2364 = ~n2357 & ~n2359 ;
  assign n2365 = ~n2363 & n2364 ;
  assign n2366 = ~n2349 & n2365 ;
  assign n2367 = ~n2353 & n2366 ;
  assign n2394 = \P1_InstQueueWr_Addr_reg[3]/NET0131  & n2367 ;
  assign n2274 = ~n2272 & ~n2273 ;
  assign n2275 = ~n2271 & n2274 ;
  assign n2319 = ~\P1_InstQueueRd_Addr_reg[1]/NET0131  & ~\P1_InstQueueRd_Addr_reg[2]/NET0131  ;
  assign n2320 = ~n2318 & ~n2319 ;
  assign n2330 = n2237 & n2320 ;
  assign n2338 = ~\P1_InstQueueRd_Addr_reg[2]/NET0131  & ~n2337 ;
  assign n2339 = n2274 & n2337 ;
  assign n2340 = ~n2338 & ~n2339 ;
  assign n2341 = ~n2332 & n2340 ;
  assign n2342 = ~n2330 & ~n2341 ;
  assign n2343 = ~n2275 & n2342 ;
  assign n2315 = \P1_InstQueueRd_Addr_reg[2]/NET0131  & ~n2232 ;
  assign n2316 = n2314 & ~n2315 ;
  assign n2321 = ~n2317 & ~n2320 ;
  assign n2322 = ~\P1_InstQueueRd_Addr_reg[2]/NET0131  & n2317 ;
  assign n2323 = ~n2321 & ~n2322 ;
  assign n2324 = ~n2316 & n2323 ;
  assign n2329 = \P1_InstQueueRd_Addr_reg[2]/NET0131  & ~n2328 ;
  assign n2344 = ~n2324 & ~n2329 ;
  assign n2345 = n2343 & n2344 ;
  assign n2417 = \P1_InstQueueWr_Addr_reg[2]/NET0131  & n2345 ;
  assign n2418 = ~n2394 & ~n2417 ;
  assign n2419 = ~n2409 & n2418 ;
  assign n2420 = ~n2416 & n2419 ;
  assign n2395 = ~\P1_InstQueueWr_Addr_reg[2]/NET0131  & ~n2345 ;
  assign n2396 = ~n2394 & n2395 ;
  assign n2346 = \P1_InstQueueWr_Addr_reg[3]/NET0131  & n2345 ;
  assign n2368 = ~n2346 & ~n2367 ;
  assign n2380 = ~\P1_More_reg/NET0131  & ~n2301 ;
  assign n2381 = n2379 & ~n2380 ;
  assign n2369 = n2243 & ~n2337 ;
  assign n2373 = ~n2369 & n2372 ;
  assign n2374 = n2300 & ~n2334 ;
  assign n2375 = n2295 & ~n2374 ;
  assign n2376 = n2244 & n2375 ;
  assign n2382 = n2373 & ~n2376 ;
  assign n2383 = ~n2381 & n2382 ;
  assign n2386 = n2304 & n2317 ;
  assign n2387 = ~n2311 & ~n2317 ;
  assign n2388 = ~n2306 & ~n2387 ;
  assign n2389 = ~n2301 & n2388 ;
  assign n2390 = ~n2386 & ~n2389 ;
  assign n2391 = \P1_Flush_reg/NET0131  & ~n2390 ;
  assign n2384 = n2244 & ~n2375 ;
  assign n2385 = n2243 & n2337 ;
  assign n2392 = ~n2384 & ~n2385 ;
  assign n2393 = ~n2391 & n2392 ;
  assign n2421 = n2383 & n2393 ;
  assign n2422 = ~n2368 & n2421 ;
  assign n2423 = ~n2396 & n2422 ;
  assign n2424 = ~n2420 & n2423 ;
  assign n2425 = ~\P1_DataWidth_reg[1]/NET0131  & ~n2317 ;
  assign n2426 = n2225 & n2312 ;
  assign n2427 = n2425 & n2426 ;
  assign n2428 = ~\P1_State2_reg[1]/NET0131  & ~n2427 ;
  assign n2429 = n2424 & n2428 ;
  assign n2430 = ~\P1_State2_reg[1]/NET0131  & \P1_State2_reg[2]/NET0131  ;
  assign n2431 = ~\P1_State2_reg[3]/NET0131  & n2430 ;
  assign n2432 = \P1_State2_reg[0]/NET0131  & n2431 ;
  assign n2433 = ~n2429 & n2432 ;
  assign n2438 = \P1_State2_reg[1]/NET0131  & \P1_State2_reg[2]/NET0131  ;
  assign n2439 = ~\P1_State2_reg[3]/NET0131  & n2438 ;
  assign n2440 = ~\P1_State2_reg[0]/NET0131  & n2439 ;
  assign n2434 = \P1_State2_reg[1]/NET0131  & ~\P1_State2_reg[2]/NET0131  ;
  assign n2435 = ~\P1_State2_reg[3]/NET0131  & n2434 ;
  assign n2441 = \P1_State2_reg[0]/NET0131  & n2435 ;
  assign n2442 = ~n2440 & ~n2441 ;
  assign n2443 = n2317 & ~n2442 ;
  assign n2436 = ~\P1_State2_reg[0]/NET0131  & n2435 ;
  assign n2437 = ~\P1_DataWidth_reg[1]/NET0131  & n2436 ;
  assign n2444 = \P1_State2_reg[0]/NET0131  & ~\P1_State2_reg[3]/NET0131  ;
  assign n2445 = ~\P1_State2_reg[2]/NET0131  & n2444 ;
  assign n2446 = ~\P1_State2_reg[1]/NET0131  & n2445 ;
  assign n2447 = ~n2317 & n2446 ;
  assign n2448 = ~n2437 & ~n2447 ;
  assign n2449 = ~n2443 & n2448 ;
  assign n2450 = ~n2433 & n2449 ;
  assign n2451 = \P3_State2_reg[0]/NET0131  & ~\P3_State2_reg[3]/NET0131  ;
  assign n2452 = ~\P3_State2_reg[1]/NET0131  & \P3_State2_reg[2]/NET0131  ;
  assign n2453 = n2451 & n2452 ;
  assign n2458 = \P3_InstQueueRd_Addr_reg[2]/NET0131  & ~\P3_InstQueueRd_Addr_reg[3]/NET0131  ;
  assign n2468 = ~\P3_InstQueueRd_Addr_reg[0]/NET0131  & ~\P3_InstQueueRd_Addr_reg[1]/NET0131  ;
  assign n2469 = n2458 & n2468 ;
  assign n2470 = \P3_InstQueue_reg[4][6]/NET0131  & n2469 ;
  assign n2471 = \P3_InstQueueRd_Addr_reg[2]/NET0131  & \P3_InstQueueRd_Addr_reg[3]/NET0131  ;
  assign n2472 = n2468 & n2471 ;
  assign n2473 = \P3_InstQueue_reg[12][6]/NET0131  & n2472 ;
  assign n2496 = ~n2470 & ~n2473 ;
  assign n2462 = ~\P3_InstQueueRd_Addr_reg[0]/NET0131  & \P3_InstQueueRd_Addr_reg[1]/NET0131  ;
  assign n2474 = n2458 & n2462 ;
  assign n2475 = \P3_InstQueue_reg[6][6]/NET0131  & n2474 ;
  assign n2463 = ~\P3_InstQueueRd_Addr_reg[2]/NET0131  & \P3_InstQueueRd_Addr_reg[3]/NET0131  ;
  assign n2476 = n2463 & n2468 ;
  assign n2477 = \P3_InstQueue_reg[8][6]/NET0131  & n2476 ;
  assign n2497 = ~n2475 & ~n2477 ;
  assign n2504 = n2496 & n2497 ;
  assign n2454 = ~\P3_InstQueueRd_Addr_reg[2]/NET0131  & ~\P3_InstQueueRd_Addr_reg[3]/NET0131  ;
  assign n2455 = \P3_InstQueueRd_Addr_reg[0]/NET0131  & ~\P3_InstQueueRd_Addr_reg[1]/NET0131  ;
  assign n2456 = n2454 & n2455 ;
  assign n2457 = \P3_InstQueue_reg[1][6]/NET0131  & n2456 ;
  assign n2459 = \P3_InstQueueRd_Addr_reg[0]/NET0131  & \P3_InstQueueRd_Addr_reg[1]/NET0131  ;
  assign n2460 = n2458 & n2459 ;
  assign n2461 = \P3_InstQueue_reg[7][6]/NET0131  & n2460 ;
  assign n2494 = ~n2457 & ~n2461 ;
  assign n2464 = n2462 & n2463 ;
  assign n2465 = \P3_InstQueue_reg[10][6]/NET0131  & n2464 ;
  assign n2466 = n2454 & n2462 ;
  assign n2467 = \P3_InstQueue_reg[2][6]/NET0131  & n2466 ;
  assign n2495 = ~n2465 & ~n2467 ;
  assign n2505 = n2494 & n2495 ;
  assign n2506 = n2504 & n2505 ;
  assign n2486 = n2459 & n2463 ;
  assign n2487 = \P3_InstQueue_reg[11][6]/NET0131  & n2486 ;
  assign n2488 = n2462 & n2471 ;
  assign n2489 = \P3_InstQueue_reg[14][6]/NET0131  & n2488 ;
  assign n2500 = ~n2487 & ~n2489 ;
  assign n2490 = n2455 & n2463 ;
  assign n2491 = \P3_InstQueue_reg[9][6]/NET0131  & n2490 ;
  assign n2492 = n2455 & n2458 ;
  assign n2493 = \P3_InstQueue_reg[5][6]/NET0131  & n2492 ;
  assign n2501 = ~n2491 & ~n2493 ;
  assign n2502 = n2500 & n2501 ;
  assign n2478 = n2455 & n2471 ;
  assign n2479 = \P3_InstQueue_reg[13][6]/NET0131  & n2478 ;
  assign n2480 = n2454 & n2459 ;
  assign n2481 = \P3_InstQueue_reg[3][6]/NET0131  & n2480 ;
  assign n2498 = ~n2479 & ~n2481 ;
  assign n2482 = n2454 & n2468 ;
  assign n2483 = \P3_InstQueue_reg[0][6]/NET0131  & n2482 ;
  assign n2484 = n2459 & n2471 ;
  assign n2485 = \P3_InstQueue_reg[15][6]/NET0131  & n2484 ;
  assign n2499 = ~n2483 & ~n2485 ;
  assign n2503 = n2498 & n2499 ;
  assign n2507 = n2502 & n2503 ;
  assign n2508 = n2506 & n2507 ;
  assign n2513 = \P3_InstQueue_reg[10][7]/NET0131  & n2464 ;
  assign n2514 = \P3_InstQueue_reg[13][7]/NET0131  & n2478 ;
  assign n2527 = ~n2513 & ~n2514 ;
  assign n2515 = \P3_InstQueue_reg[8][7]/NET0131  & n2476 ;
  assign n2516 = \P3_InstQueue_reg[4][7]/NET0131  & n2469 ;
  assign n2528 = ~n2515 & ~n2516 ;
  assign n2535 = n2527 & n2528 ;
  assign n2509 = \P3_InstQueue_reg[1][7]/NET0131  & n2456 ;
  assign n2510 = \P3_InstQueue_reg[11][7]/NET0131  & n2486 ;
  assign n2525 = ~n2509 & ~n2510 ;
  assign n2511 = \P3_InstQueue_reg[6][7]/NET0131  & n2474 ;
  assign n2512 = \P3_InstQueue_reg[15][7]/NET0131  & n2484 ;
  assign n2526 = ~n2511 & ~n2512 ;
  assign n2536 = n2525 & n2526 ;
  assign n2537 = n2535 & n2536 ;
  assign n2521 = \P3_InstQueue_reg[9][7]/NET0131  & n2490 ;
  assign n2522 = \P3_InstQueue_reg[3][7]/NET0131  & n2480 ;
  assign n2531 = ~n2521 & ~n2522 ;
  assign n2523 = \P3_InstQueue_reg[5][7]/NET0131  & n2492 ;
  assign n2524 = \P3_InstQueue_reg[7][7]/NET0131  & n2460 ;
  assign n2532 = ~n2523 & ~n2524 ;
  assign n2533 = n2531 & n2532 ;
  assign n2517 = \P3_InstQueue_reg[2][7]/NET0131  & n2466 ;
  assign n2518 = \P3_InstQueue_reg[14][7]/NET0131  & n2488 ;
  assign n2529 = ~n2517 & ~n2518 ;
  assign n2519 = \P3_InstQueue_reg[12][7]/NET0131  & n2472 ;
  assign n2520 = \P3_InstQueue_reg[0][7]/NET0131  & n2482 ;
  assign n2530 = ~n2519 & ~n2520 ;
  assign n2534 = n2529 & n2530 ;
  assign n2538 = n2533 & n2534 ;
  assign n2539 = n2537 & n2538 ;
  assign n2753 = ~n2508 & ~n2539 ;
  assign n2545 = \P3_InstQueue_reg[0][4]/NET0131  & n2482 ;
  assign n2546 = \P3_InstQueue_reg[11][4]/NET0131  & n2486 ;
  assign n2559 = ~n2545 & ~n2546 ;
  assign n2547 = \P3_InstQueue_reg[1][4]/NET0131  & n2456 ;
  assign n2548 = \P3_InstQueue_reg[2][4]/NET0131  & n2466 ;
  assign n2560 = ~n2547 & ~n2548 ;
  assign n2567 = n2559 & n2560 ;
  assign n2541 = \P3_InstQueue_reg[7][4]/NET0131  & n2460 ;
  assign n2542 = \P3_InstQueue_reg[13][4]/NET0131  & n2478 ;
  assign n2557 = ~n2541 & ~n2542 ;
  assign n2543 = \P3_InstQueue_reg[5][4]/NET0131  & n2492 ;
  assign n2544 = \P3_InstQueue_reg[15][4]/NET0131  & n2484 ;
  assign n2558 = ~n2543 & ~n2544 ;
  assign n2568 = n2557 & n2558 ;
  assign n2569 = n2567 & n2568 ;
  assign n2553 = \P3_InstQueue_reg[14][4]/NET0131  & n2488 ;
  assign n2554 = \P3_InstQueue_reg[6][4]/NET0131  & n2474 ;
  assign n2563 = ~n2553 & ~n2554 ;
  assign n2555 = \P3_InstQueue_reg[10][4]/NET0131  & n2464 ;
  assign n2556 = \P3_InstQueue_reg[8][4]/NET0131  & n2476 ;
  assign n2564 = ~n2555 & ~n2556 ;
  assign n2565 = n2563 & n2564 ;
  assign n2549 = \P3_InstQueue_reg[3][4]/NET0131  & n2480 ;
  assign n2550 = \P3_InstQueue_reg[12][4]/NET0131  & n2472 ;
  assign n2561 = ~n2549 & ~n2550 ;
  assign n2551 = \P3_InstQueue_reg[4][4]/NET0131  & n2469 ;
  assign n2552 = \P3_InstQueue_reg[9][4]/NET0131  & n2490 ;
  assign n2562 = ~n2551 & ~n2552 ;
  assign n2566 = n2561 & n2562 ;
  assign n2570 = n2565 & n2566 ;
  assign n2571 = n2569 & n2570 ;
  assign n2577 = \P3_InstQueue_reg[8][5]/NET0131  & n2476 ;
  assign n2578 = \P3_InstQueue_reg[0][5]/NET0131  & n2482 ;
  assign n2591 = ~n2577 & ~n2578 ;
  assign n2579 = \P3_InstQueue_reg[1][5]/NET0131  & n2456 ;
  assign n2580 = \P3_InstQueue_reg[13][5]/NET0131  & n2478 ;
  assign n2592 = ~n2579 & ~n2580 ;
  assign n2599 = n2591 & n2592 ;
  assign n2573 = \P3_InstQueue_reg[11][5]/NET0131  & n2486 ;
  assign n2574 = \P3_InstQueue_reg[5][5]/NET0131  & n2492 ;
  assign n2589 = ~n2573 & ~n2574 ;
  assign n2575 = \P3_InstQueue_reg[9][5]/NET0131  & n2490 ;
  assign n2576 = \P3_InstQueue_reg[10][5]/NET0131  & n2464 ;
  assign n2590 = ~n2575 & ~n2576 ;
  assign n2600 = n2589 & n2590 ;
  assign n2601 = n2599 & n2600 ;
  assign n2585 = \P3_InstQueue_reg[3][5]/NET0131  & n2480 ;
  assign n2586 = \P3_InstQueue_reg[7][5]/NET0131  & n2460 ;
  assign n2595 = ~n2585 & ~n2586 ;
  assign n2587 = \P3_InstQueue_reg[2][5]/NET0131  & n2466 ;
  assign n2588 = \P3_InstQueue_reg[6][5]/NET0131  & n2474 ;
  assign n2596 = ~n2587 & ~n2588 ;
  assign n2597 = n2595 & n2596 ;
  assign n2581 = \P3_InstQueue_reg[14][5]/NET0131  & n2488 ;
  assign n2582 = \P3_InstQueue_reg[4][5]/NET0131  & n2469 ;
  assign n2593 = ~n2581 & ~n2582 ;
  assign n2583 = \P3_InstQueue_reg[12][5]/NET0131  & n2472 ;
  assign n2584 = \P3_InstQueue_reg[15][5]/NET0131  & n2484 ;
  assign n2594 = ~n2583 & ~n2584 ;
  assign n2598 = n2593 & n2594 ;
  assign n2602 = n2597 & n2598 ;
  assign n2603 = n2601 & n2602 ;
  assign n2754 = n2571 & ~n2603 ;
  assign n2755 = n2753 & n2754 ;
  assign n2609 = \P3_InstQueue_reg[7][2]/NET0131  & n2460 ;
  assign n2610 = \P3_InstQueue_reg[4][2]/NET0131  & n2469 ;
  assign n2623 = ~n2609 & ~n2610 ;
  assign n2611 = \P3_InstQueue_reg[3][2]/NET0131  & n2480 ;
  assign n2612 = \P3_InstQueue_reg[0][2]/NET0131  & n2482 ;
  assign n2624 = ~n2611 & ~n2612 ;
  assign n2631 = n2623 & n2624 ;
  assign n2605 = \P3_InstQueue_reg[10][2]/NET0131  & n2464 ;
  assign n2606 = \P3_InstQueue_reg[1][2]/NET0131  & n2456 ;
  assign n2621 = ~n2605 & ~n2606 ;
  assign n2607 = \P3_InstQueue_reg[6][2]/NET0131  & n2474 ;
  assign n2608 = \P3_InstQueue_reg[11][2]/NET0131  & n2486 ;
  assign n2622 = ~n2607 & ~n2608 ;
  assign n2632 = n2621 & n2622 ;
  assign n2633 = n2631 & n2632 ;
  assign n2617 = \P3_InstQueue_reg[2][2]/NET0131  & n2466 ;
  assign n2618 = \P3_InstQueue_reg[5][2]/NET0131  & n2492 ;
  assign n2627 = ~n2617 & ~n2618 ;
  assign n2619 = \P3_InstQueue_reg[13][2]/NET0131  & n2478 ;
  assign n2620 = \P3_InstQueue_reg[9][2]/NET0131  & n2490 ;
  assign n2628 = ~n2619 & ~n2620 ;
  assign n2629 = n2627 & n2628 ;
  assign n2613 = \P3_InstQueue_reg[14][2]/NET0131  & n2488 ;
  assign n2614 = \P3_InstQueue_reg[12][2]/NET0131  & n2472 ;
  assign n2625 = ~n2613 & ~n2614 ;
  assign n2615 = \P3_InstQueue_reg[8][2]/NET0131  & n2476 ;
  assign n2616 = \P3_InstQueue_reg[15][2]/NET0131  & n2484 ;
  assign n2626 = ~n2615 & ~n2616 ;
  assign n2630 = n2625 & n2626 ;
  assign n2634 = n2629 & n2630 ;
  assign n2635 = n2633 & n2634 ;
  assign n2640 = \P3_InstQueue_reg[12][0]/NET0131  & n2472 ;
  assign n2641 = \P3_InstQueue_reg[4][0]/NET0131  & n2469 ;
  assign n2654 = ~n2640 & ~n2641 ;
  assign n2642 = \P3_InstQueue_reg[3][0]/NET0131  & n2480 ;
  assign n2643 = \P3_InstQueue_reg[0][0]/NET0131  & n2482 ;
  assign n2655 = ~n2642 & ~n2643 ;
  assign n2662 = n2654 & n2655 ;
  assign n2636 = \P3_InstQueue_reg[1][0]/NET0131  & n2456 ;
  assign n2637 = \P3_InstQueue_reg[15][0]/NET0131  & n2484 ;
  assign n2652 = ~n2636 & ~n2637 ;
  assign n2638 = \P3_InstQueue_reg[7][0]/NET0131  & n2460 ;
  assign n2639 = \P3_InstQueue_reg[9][0]/NET0131  & n2490 ;
  assign n2653 = ~n2638 & ~n2639 ;
  assign n2663 = n2652 & n2653 ;
  assign n2664 = n2662 & n2663 ;
  assign n2648 = \P3_InstQueue_reg[2][0]/NET0131  & n2466 ;
  assign n2649 = \P3_InstQueue_reg[13][0]/NET0131  & n2478 ;
  assign n2658 = ~n2648 & ~n2649 ;
  assign n2650 = \P3_InstQueue_reg[10][0]/NET0131  & n2464 ;
  assign n2651 = \P3_InstQueue_reg[11][0]/NET0131  & n2486 ;
  assign n2659 = ~n2650 & ~n2651 ;
  assign n2660 = n2658 & n2659 ;
  assign n2644 = \P3_InstQueue_reg[5][0]/NET0131  & n2492 ;
  assign n2645 = \P3_InstQueue_reg[8][0]/NET0131  & n2476 ;
  assign n2656 = ~n2644 & ~n2645 ;
  assign n2646 = \P3_InstQueue_reg[6][0]/NET0131  & n2474 ;
  assign n2647 = \P3_InstQueue_reg[14][0]/NET0131  & n2488 ;
  assign n2657 = ~n2646 & ~n2647 ;
  assign n2661 = n2656 & n2657 ;
  assign n2665 = n2660 & n2661 ;
  assign n2666 = n2664 & n2665 ;
  assign n2711 = \P3_InstQueue_reg[11][3]/NET0131  & n2486 ;
  assign n2712 = \P3_InstQueue_reg[5][3]/NET0131  & n2492 ;
  assign n2725 = ~n2711 & ~n2712 ;
  assign n2713 = \P3_InstQueue_reg[7][3]/NET0131  & n2460 ;
  assign n2714 = \P3_InstQueue_reg[14][3]/NET0131  & n2488 ;
  assign n2726 = ~n2713 & ~n2714 ;
  assign n2733 = n2725 & n2726 ;
  assign n2707 = \P3_InstQueue_reg[4][3]/NET0131  & n2469 ;
  assign n2708 = \P3_InstQueue_reg[13][3]/NET0131  & n2478 ;
  assign n2723 = ~n2707 & ~n2708 ;
  assign n2709 = \P3_InstQueue_reg[12][3]/NET0131  & n2472 ;
  assign n2710 = \P3_InstQueue_reg[6][3]/NET0131  & n2474 ;
  assign n2724 = ~n2709 & ~n2710 ;
  assign n2734 = n2723 & n2724 ;
  assign n2735 = n2733 & n2734 ;
  assign n2719 = \P3_InstQueue_reg[0][3]/NET0131  & n2482 ;
  assign n2720 = \P3_InstQueue_reg[9][3]/NET0131  & n2490 ;
  assign n2729 = ~n2719 & ~n2720 ;
  assign n2721 = \P3_InstQueue_reg[15][3]/NET0131  & n2484 ;
  assign n2722 = \P3_InstQueue_reg[10][3]/NET0131  & n2464 ;
  assign n2730 = ~n2721 & ~n2722 ;
  assign n2731 = n2729 & n2730 ;
  assign n2715 = \P3_InstQueue_reg[8][3]/NET0131  & n2476 ;
  assign n2716 = \P3_InstQueue_reg[2][3]/NET0131  & n2466 ;
  assign n2727 = ~n2715 & ~n2716 ;
  assign n2717 = \P3_InstQueue_reg[1][3]/NET0131  & n2456 ;
  assign n2718 = \P3_InstQueue_reg[3][3]/NET0131  & n2480 ;
  assign n2728 = ~n2717 & ~n2718 ;
  assign n2732 = n2727 & n2728 ;
  assign n2736 = n2731 & n2732 ;
  assign n2737 = n2735 & n2736 ;
  assign n2760 = ~n2666 & ~n2737 ;
  assign n2761 = n2635 & n2760 ;
  assign n2762 = n2755 & n2761 ;
  assign n2749 = ~n2635 & n2666 ;
  assign n2750 = n2737 & n2749 ;
  assign n2763 = n2750 & n2755 ;
  assign n2540 = n2508 & ~n2539 ;
  assign n2701 = n2571 & n2603 ;
  assign n2764 = n2540 & n2701 ;
  assign n2765 = n2761 & n2764 ;
  assign n2766 = ~n2763 & ~n2765 ;
  assign n2667 = n2635 & n2666 ;
  assign n2672 = \P3_InstQueue_reg[10][1]/NET0131  & n2464 ;
  assign n2673 = \P3_InstQueue_reg[3][1]/NET0131  & n2480 ;
  assign n2686 = ~n2672 & ~n2673 ;
  assign n2674 = \P3_InstQueue_reg[8][1]/NET0131  & n2476 ;
  assign n2675 = \P3_InstQueue_reg[12][1]/NET0131  & n2472 ;
  assign n2687 = ~n2674 & ~n2675 ;
  assign n2694 = n2686 & n2687 ;
  assign n2668 = \P3_InstQueue_reg[1][1]/NET0131  & n2456 ;
  assign n2669 = \P3_InstQueue_reg[11][1]/NET0131  & n2486 ;
  assign n2684 = ~n2668 & ~n2669 ;
  assign n2670 = \P3_InstQueue_reg[4][1]/NET0131  & n2469 ;
  assign n2671 = \P3_InstQueue_reg[14][1]/NET0131  & n2488 ;
  assign n2685 = ~n2670 & ~n2671 ;
  assign n2695 = n2684 & n2685 ;
  assign n2696 = n2694 & n2695 ;
  assign n2680 = \P3_InstQueue_reg[6][1]/NET0131  & n2474 ;
  assign n2681 = \P3_InstQueue_reg[5][1]/NET0131  & n2492 ;
  assign n2690 = ~n2680 & ~n2681 ;
  assign n2682 = \P3_InstQueue_reg[13][1]/NET0131  & n2478 ;
  assign n2683 = \P3_InstQueue_reg[15][1]/NET0131  & n2484 ;
  assign n2691 = ~n2682 & ~n2683 ;
  assign n2692 = n2690 & n2691 ;
  assign n2676 = \P3_InstQueue_reg[2][1]/NET0131  & n2466 ;
  assign n2677 = \P3_InstQueue_reg[9][1]/NET0131  & n2490 ;
  assign n2688 = ~n2676 & ~n2677 ;
  assign n2678 = \P3_InstQueue_reg[0][1]/NET0131  & n2482 ;
  assign n2679 = \P3_InstQueue_reg[7][1]/NET0131  & n2460 ;
  assign n2689 = ~n2678 & ~n2679 ;
  assign n2693 = n2688 & n2689 ;
  assign n2697 = n2692 & n2693 ;
  assign n2698 = n2696 & n2697 ;
  assign n2699 = n2667 & n2698 ;
  assign n2739 = n2603 & n2737 ;
  assign n2740 = n2699 & n2739 ;
  assign n2767 = n2740 & n2753 ;
  assign n2768 = n2766 & ~n2767 ;
  assign n2769 = ~n2762 & n2768 ;
  assign n2572 = n2540 & ~n2571 ;
  assign n2604 = n2572 & ~n2603 ;
  assign n2700 = n2604 & n2699 ;
  assign n2745 = n2635 & ~n2698 ;
  assign n2770 = n2604 & n2760 ;
  assign n2771 = n2745 & n2770 ;
  assign n2772 = ~n2700 & ~n2771 ;
  assign n2773 = n2769 & n2772 ;
  assign n2741 = ~n2508 & n2539 ;
  assign n2742 = n2571 & n2741 ;
  assign n2751 = ~n2603 & n2742 ;
  assign n2752 = n2750 & n2751 ;
  assign n2756 = n2667 & ~n2737 ;
  assign n2757 = n2755 & n2756 ;
  assign n2758 = ~n2752 & ~n2757 ;
  assign n2759 = ~n2698 & ~n2758 ;
  assign n2702 = n2508 & n2539 ;
  assign n2703 = ~n2635 & n2698 ;
  assign n2704 = n2702 & n2703 ;
  assign n2705 = n2701 & n2704 ;
  assign n2706 = ~n2700 & ~n2705 ;
  assign n2738 = ~n2706 & n2737 ;
  assign n2743 = ~n2572 & ~n2742 ;
  assign n2744 = n2740 & ~n2743 ;
  assign n2746 = ~n2666 & n2739 ;
  assign n2747 = n2745 & n2746 ;
  assign n2748 = n2742 & n2747 ;
  assign n2774 = ~n2744 & ~n2748 ;
  assign n2775 = ~n2738 & n2774 ;
  assign n2776 = ~n2759 & n2775 ;
  assign n2777 = ~n2773 & n2776 ;
  assign n2840 = n2700 & ~n2737 ;
  assign n2841 = ~n2771 & ~n2840 ;
  assign n2787 = ~\P3_InstQueueRd_Addr_reg[3]/NET0131  & \P3_InstQueueWr_Addr_reg[3]/NET0131  ;
  assign n2788 = \P3_InstQueueRd_Addr_reg[3]/NET0131  & ~\P3_InstQueueWr_Addr_reg[3]/NET0131  ;
  assign n2790 = ~\P3_InstQueueRd_Addr_reg[2]/NET0131  & \P3_InstQueueWr_Addr_reg[2]/NET0131  ;
  assign n2791 = \P3_InstQueueRd_Addr_reg[2]/NET0131  & ~\P3_InstQueueWr_Addr_reg[2]/NET0131  ;
  assign n2792 = ~\P3_InstQueueRd_Addr_reg[1]/NET0131  & \P3_InstQueueWr_Addr_reg[1]/NET0131  ;
  assign n2793 = \P3_InstQueueRd_Addr_reg[1]/NET0131  & ~\P3_InstQueueWr_Addr_reg[1]/NET0131  ;
  assign n2794 = \P3_InstQueueRd_Addr_reg[0]/NET0131  & ~\P3_InstQueueWr_Addr_reg[0]/NET0131  ;
  assign n2795 = ~n2793 & ~n2794 ;
  assign n2796 = ~n2792 & ~n2795 ;
  assign n2797 = ~n2791 & ~n2796 ;
  assign n2798 = ~n2790 & ~n2797 ;
  assign n2807 = ~n2788 & ~n2798 ;
  assign n2808 = ~n2787 & ~n2807 ;
  assign n2789 = ~n2787 & ~n2788 ;
  assign n2799 = n2789 & n2798 ;
  assign n2800 = ~n2789 & ~n2798 ;
  assign n2801 = ~n2799 & ~n2800 ;
  assign n2802 = ~n2790 & ~n2791 ;
  assign n2803 = n2796 & ~n2802 ;
  assign n2804 = ~n2796 & n2802 ;
  assign n2805 = ~n2803 & ~n2804 ;
  assign n2810 = ~n2792 & ~n2793 ;
  assign n2842 = ~\P3_InstQueueRd_Addr_reg[0]/NET0131  & \P3_InstQueueWr_Addr_reg[0]/NET0131  ;
  assign n2843 = ~n2794 & ~n2842 ;
  assign n2844 = n2810 & n2843 ;
  assign n2845 = n2805 & ~n2844 ;
  assign n2846 = n2801 & ~n2845 ;
  assign n2847 = ~n2808 & ~n2846 ;
  assign n2918 = ~n2841 & n2847 ;
  assign n2919 = n2777 & ~n2918 ;
  assign n2920 = ~n2459 & ~n2468 ;
  assign n2921 = ~n2919 & n2920 ;
  assign n2806 = n2801 & ~n2805 ;
  assign n2809 = ~n2806 & ~n2808 ;
  assign n2811 = n2794 & ~n2810 ;
  assign n2812 = ~n2794 & n2810 ;
  assign n2813 = ~n2811 & ~n2812 ;
  assign n2814 = ~n2808 & n2813 ;
  assign n2815 = ~n2809 & ~n2814 ;
  assign n2820 = n2698 & n2763 ;
  assign n2821 = ~n2698 & n2765 ;
  assign n2822 = ~n2820 & ~n2821 ;
  assign n2832 = ~n2815 & ~n2822 ;
  assign n2782 = ~\P3_State_reg[0]/NET0131  & \P3_State_reg[1]/NET0131  ;
  assign n2783 = ~\P3_State_reg[2]/NET0131  & n2782 ;
  assign n2784 = ~\P3_State_reg[0]/NET0131  & ~\P3_State_reg[1]/NET0131  ;
  assign n2785 = \P3_State_reg[2]/NET0131  & n2784 ;
  assign n2786 = ~n2783 & ~n2785 ;
  assign n2816 = ~n2786 & ~n2815 ;
  assign n2817 = ~n2698 & n2763 ;
  assign n2818 = n2698 & n2765 ;
  assign n2819 = ~n2817 & ~n2818 ;
  assign n2833 = n2816 & ~n2819 ;
  assign n2834 = ~n2832 & ~n2833 ;
  assign n2835 = \ready22_reg/NET0131  & \ready2_pad  ;
  assign n2922 = ~n2834 & ~n2835 ;
  assign n2923 = ~n2767 & ~n2922 ;
  assign n2924 = ~\P3_InstQueueRd_Addr_reg[1]/NET0131  & n2923 ;
  assign n2862 = ~n2815 & ~n2835 ;
  assign n2863 = n2821 & ~n2862 ;
  assign n2864 = n2820 & ~n2862 ;
  assign n2865 = ~n2863 & ~n2864 ;
  assign n2874 = ~n2786 & ~n2835 ;
  assign n2875 = ~n2815 & n2874 ;
  assign n2890 = ~n2819 & ~n2875 ;
  assign n2891 = n2865 & ~n2890 ;
  assign n2898 = ~n2841 & ~n2847 ;
  assign n2925 = n2891 & ~n2898 ;
  assign n2926 = \P3_InstQueueRd_Addr_reg[1]/NET0131  & ~n2762 ;
  assign n2927 = n2925 & n2926 ;
  assign n2928 = ~n2924 & ~n2927 ;
  assign n2929 = ~n2921 & ~n2928 ;
  assign n2931 = ~\P3_InstQueueWr_Addr_reg[1]/NET0131  & ~n2929 ;
  assign n2932 = ~\P3_InstQueueRd_Addr_reg[0]/NET0131  & n2919 ;
  assign n2933 = \P3_InstQueueRd_Addr_reg[0]/NET0131  & n2769 ;
  assign n2934 = ~n2898 & n2933 ;
  assign n2935 = ~n2932 & ~n2934 ;
  assign n2936 = \P3_InstQueueWr_Addr_reg[0]/NET0131  & ~n2935 ;
  assign n2937 = ~n2931 & n2936 ;
  assign n2823 = n2815 & ~n2822 ;
  assign n2824 = n2819 & ~n2823 ;
  assign n2825 = ~n2816 & ~n2824 ;
  assign n2826 = ~n2762 & ~n2825 ;
  assign n2827 = \P3_InstQueueRd_Addr_reg[2]/NET0131  & ~n2826 ;
  assign n2778 = \P3_InstQueueRd_Addr_reg[2]/NET0131  & n2459 ;
  assign n2779 = ~\P3_InstQueueRd_Addr_reg[2]/NET0131  & ~n2459 ;
  assign n2780 = ~n2778 & ~n2779 ;
  assign n2781 = ~n2777 & n2780 ;
  assign n2828 = \P3_InstQueueRd_Addr_reg[1]/NET0131  & \P3_InstQueueRd_Addr_reg[2]/NET0131  ;
  assign n2829 = ~\P3_InstQueueRd_Addr_reg[1]/NET0131  & ~\P3_InstQueueRd_Addr_reg[2]/NET0131  ;
  assign n2830 = ~n2828 & ~n2829 ;
  assign n2836 = ~n2830 & ~n2835 ;
  assign n2837 = ~\P3_InstQueueRd_Addr_reg[2]/NET0131  & n2835 ;
  assign n2838 = ~n2836 & ~n2837 ;
  assign n2839 = ~n2834 & n2838 ;
  assign n2831 = n2767 & n2830 ;
  assign n2848 = ~\P3_InstQueueRd_Addr_reg[2]/NET0131  & ~n2847 ;
  assign n2849 = n2780 & n2847 ;
  assign n2850 = ~n2848 & ~n2849 ;
  assign n2851 = ~n2841 & n2850 ;
  assign n2852 = ~n2831 & ~n2851 ;
  assign n2853 = ~n2839 & n2852 ;
  assign n2854 = ~n2781 & n2853 ;
  assign n2855 = ~n2827 & n2854 ;
  assign n2938 = \P3_InstQueueWr_Addr_reg[2]/NET0131  & n2855 ;
  assign n2857 = n2832 & ~n2835 ;
  assign n2858 = ~n2767 & ~n2857 ;
  assign n2859 = n2828 & ~n2858 ;
  assign n2860 = ~\P3_InstQueueRd_Addr_reg[3]/NET0131  & ~n2859 ;
  assign n2861 = ~n2767 & n2822 ;
  assign n2866 = \P3_InstQueueRd_Addr_reg[1]/NET0131  & n2471 ;
  assign n2867 = n2865 & n2866 ;
  assign n2868 = ~n2861 & ~n2867 ;
  assign n2869 = ~n2762 & ~n2868 ;
  assign n2870 = ~n2860 & ~n2869 ;
  assign n2871 = \P3_InstQueueRd_Addr_reg[3]/NET0131  & ~n2778 ;
  assign n2872 = ~n2460 & ~n2871 ;
  assign n2873 = ~n2777 & ~n2872 ;
  assign n2876 = n2828 & n2875 ;
  assign n2877 = \P3_InstQueueRd_Addr_reg[3]/NET0131  & ~n2876 ;
  assign n2878 = ~\P3_InstQueueRd_Addr_reg[3]/NET0131  & n2876 ;
  assign n2879 = ~n2877 & ~n2878 ;
  assign n2880 = ~n2819 & ~n2879 ;
  assign n2881 = ~n2779 & n2847 ;
  assign n2882 = \P3_InstQueueRd_Addr_reg[3]/NET0131  & n2881 ;
  assign n2883 = ~\P3_InstQueueRd_Addr_reg[3]/NET0131  & ~n2881 ;
  assign n2884 = ~n2882 & ~n2883 ;
  assign n2885 = ~n2841 & n2884 ;
  assign n2886 = ~n2880 & ~n2885 ;
  assign n2887 = ~n2873 & n2886 ;
  assign n2888 = ~n2870 & n2887 ;
  assign n2915 = \P3_InstQueueWr_Addr_reg[3]/NET0131  & n2888 ;
  assign n2930 = \P3_InstQueueWr_Addr_reg[1]/NET0131  & n2929 ;
  assign n2939 = ~n2915 & ~n2930 ;
  assign n2940 = ~n2938 & n2939 ;
  assign n2941 = ~n2937 & n2940 ;
  assign n2916 = ~\P3_InstQueueWr_Addr_reg[2]/NET0131  & ~n2855 ;
  assign n2917 = ~n2915 & n2916 ;
  assign n2856 = \P3_InstQueueWr_Addr_reg[3]/NET0131  & n2855 ;
  assign n2889 = ~n2856 & ~n2888 ;
  assign n2892 = ~\P3_More_reg/NET0131  & ~n2815 ;
  assign n2893 = ~n2891 & ~n2892 ;
  assign n2894 = ~n2698 & n2762 ;
  assign n2895 = n2814 & ~n2843 ;
  assign n2896 = ~n2809 & ~n2895 ;
  assign n2897 = n2894 & n2896 ;
  assign n2899 = n2698 & n2762 ;
  assign n2900 = ~n2847 & n2899 ;
  assign n2901 = ~n2898 & ~n2900 ;
  assign n2902 = ~n2897 & n2901 ;
  assign n2903 = ~n2893 & n2902 ;
  assign n2906 = n2786 & ~n2819 ;
  assign n2907 = ~n2835 & ~n2906 ;
  assign n2908 = n2765 & ~n2815 ;
  assign n2909 = n2763 & ~n2815 ;
  assign n2910 = ~n2908 & ~n2909 ;
  assign n2911 = \P3_Flush_reg/NET0131  & ~n2910 ;
  assign n2912 = ~n2907 & n2911 ;
  assign n2904 = n2894 & ~n2896 ;
  assign n2905 = n2847 & n2899 ;
  assign n2913 = ~n2904 & ~n2905 ;
  assign n2914 = ~n2912 & n2913 ;
  assign n2942 = n2903 & n2914 ;
  assign n2943 = ~n2889 & n2942 ;
  assign n2944 = ~n2917 & n2943 ;
  assign n2945 = ~n2941 & n2944 ;
  assign n2946 = ~\P3_DataWidth_reg[1]/NET0131  & ~n2835 ;
  assign n2947 = n2816 & n2946 ;
  assign n2948 = n2818 & n2947 ;
  assign n2949 = n2945 & ~n2948 ;
  assign n2950 = n2453 & ~n2949 ;
  assign n2951 = ~\P3_State2_reg[0]/NET0131  & ~\P3_State2_reg[3]/NET0131  ;
  assign n2952 = \P3_State2_reg[2]/NET0131  & n2951 ;
  assign n2953 = ~\P3_State2_reg[2]/NET0131  & n2451 ;
  assign n2954 = ~n2952 & ~n2953 ;
  assign n2955 = \P3_State2_reg[1]/NET0131  & ~n2954 ;
  assign n2956 = n2835 & n2955 ;
  assign n2957 = \P3_State2_reg[1]/NET0131  & ~\P3_State2_reg[2]/NET0131  ;
  assign n2958 = ~\P3_State2_reg[3]/NET0131  & n2957 ;
  assign n2959 = ~\P3_State2_reg[0]/NET0131  & n2958 ;
  assign n2960 = ~\P3_DataWidth_reg[1]/NET0131  & n2959 ;
  assign n2961 = ~\P3_State2_reg[1]/NET0131  & ~\P3_State2_reg[2]/NET0131  ;
  assign n2962 = \P3_State2_reg[0]/NET0131  & n2961 ;
  assign n2963 = ~\P3_State2_reg[3]/NET0131  & n2962 ;
  assign n2964 = ~n2835 & n2963 ;
  assign n2965 = ~n2960 & ~n2964 ;
  assign n2966 = ~n2956 & n2965 ;
  assign n2967 = ~n2950 & n2966 ;
  assign n2970 = \P3_DataWidth_reg[1]/NET0131  & n2959 ;
  assign n2968 = \P3_State2_reg[0]/NET0131  & n2958 ;
  assign n2969 = ~n2835 & n2968 ;
  assign n2971 = ~n2453 & ~n2952 ;
  assign n2972 = ~n2969 & n2971 ;
  assign n2973 = ~n2970 & n2972 ;
  assign n2974 = n1919 & n1923 ;
  assign n2975 = n1927 & ~n2974 ;
  assign n2976 = \P2_State2_reg[1]/NET0131  & \P2_State2_reg[2]/NET0131  ;
  assign n2979 = ~\P2_State2_reg[3]/NET0131  & n2976 ;
  assign n2980 = \P2_State2_reg[0]/NET0131  & n2979 ;
  assign n2981 = ~\P2_Flush_reg/NET0131  & \P2_InstQueueRd_Addr_reg[2]/NET0131  ;
  assign n2982 = \P2_InstQueueRd_Addr_reg[3]/NET0131  & ~n1463 ;
  assign n2983 = n2981 & n2982 ;
  assign n2984 = n2980 & ~n2983 ;
  assign n2988 = n1805 & n1933 ;
  assign n2977 = n1805 & n2976 ;
  assign n2978 = n1935 & ~n2977 ;
  assign n2985 = ~\P2_State2_reg[1]/NET0131  & ~\P2_State2_reg[2]/NET0131  ;
  assign n2986 = \P2_State2_reg[3]/NET0131  & n2985 ;
  assign n2987 = \P2_State2_reg[0]/NET0131  & n2986 ;
  assign n2989 = ~n2978 & ~n2987 ;
  assign n2990 = ~n2988 & n2989 ;
  assign n2991 = ~n2984 & n2990 ;
  assign n2992 = ~n2975 & n2991 ;
  assign n2993 = \P3_State2_reg[3]/NET0131  & n2961 ;
  assign n2994 = ~\P3_State2_reg[0]/NET0131  & n2993 ;
  assign n2995 = \P3_State2_reg[1]/NET0131  & \P3_State2_reg[2]/NET0131  ;
  assign n2996 = ~\P3_State2_reg[3]/NET0131  & n2995 ;
  assign n2997 = \P3_State2_reg[0]/NET0131  & n2996 ;
  assign n2998 = ~n2994 & ~n2997 ;
  assign n2999 = \P3_State2_reg[0]/NET0131  & ~n2947 ;
  assign n3000 = n2818 & ~n2999 ;
  assign n3001 = n2945 & n3000 ;
  assign n3002 = n2453 & ~n3001 ;
  assign n3007 = ~\P3_Flush_reg/NET0131  & \P3_InstQueueRd_Addr_reg[2]/NET0131  ;
  assign n3008 = \P3_InstQueueRd_Addr_reg[3]/NET0131  & ~n2468 ;
  assign n3009 = n3007 & n3008 ;
  assign n3010 = n2997 & ~n3009 ;
  assign n3005 = n2835 & n2995 ;
  assign n3006 = n2951 & ~n3005 ;
  assign n3003 = n2835 & n2953 ;
  assign n3004 = \P3_State2_reg[0]/NET0131  & n2993 ;
  assign n3011 = ~n3003 & ~n3004 ;
  assign n3012 = ~n3006 & n3011 ;
  assign n3013 = ~n3010 & n3012 ;
  assign n3014 = ~n3002 & n3013 ;
  assign n3025 = ~n2424 & n2432 ;
  assign n3016 = ~n2427 & n2432 ;
  assign n3020 = \P1_State2_reg[0]/NET0131  & n2439 ;
  assign n3021 = ~\P1_Flush_reg/NET0131  & \P1_InstQueueRd_Addr_reg[2]/NET0131  ;
  assign n3022 = \P1_InstQueueRd_Addr_reg[3]/NET0131  & ~n1951 ;
  assign n3023 = n3021 & n3022 ;
  assign n3024 = n3020 & ~n3023 ;
  assign n3026 = ~\P1_State2_reg[1]/NET0131  & ~\P1_State2_reg[2]/NET0131  ;
  assign n3027 = \P1_State2_reg[3]/NET0131  & n3026 ;
  assign n3028 = \P1_State2_reg[0]/NET0131  & n3027 ;
  assign n3015 = n2317 & n2445 ;
  assign n3017 = ~\P1_State2_reg[0]/NET0131  & ~\P1_State2_reg[3]/NET0131  ;
  assign n3018 = n2317 & n2438 ;
  assign n3019 = n3017 & ~n3018 ;
  assign n3029 = ~n3015 & ~n3019 ;
  assign n3030 = ~n3028 & n3029 ;
  assign n3031 = ~n3024 & n3030 ;
  assign n3032 = ~n3016 & n3031 ;
  assign n3033 = ~n3025 & n3032 ;
  assign n3035 = \P2_State2_reg[0]/NET0131  & n1930 ;
  assign n3036 = ~n1805 & n3035 ;
  assign n3034 = \P2_DataWidth_reg[1]/NET0131  & n1931 ;
  assign n3037 = ~n1927 & ~n1936 ;
  assign n3038 = ~n3034 & n3037 ;
  assign n3039 = ~n3036 & n3038 ;
  assign n3040 = ~\P2_State2_reg[0]/NET0131  & n2986 ;
  assign n3041 = ~n2980 & ~n3040 ;
  assign n3042 = ~\P1_State2_reg[0]/NET0131  & n3027 ;
  assign n3043 = ~n3020 & ~n3042 ;
  assign n3089 = ~\P2_InstQueueWr_Addr_reg[0]/NET0131  & ~\P2_InstQueueWr_Addr_reg[1]/NET0131  ;
  assign n3090 = ~\P2_InstQueueWr_Addr_reg[2]/NET0131  & n3089 ;
  assign n3091 = \P2_InstQueueWr_Addr_reg[3]/NET0131  & n3090 ;
  assign n3060 = ~\P2_Address_reg[26]/NET0131  & ~\P2_Address_reg[27]/NET0131  ;
  assign n3061 = ~\P2_Address_reg[28]/NET0131  & ~\P2_Address_reg[2]/NET0131  ;
  assign n3067 = n3060 & n3061 ;
  assign n3058 = ~\P2_Address_reg[22]/NET0131  & ~\P2_Address_reg[23]/NET0131  ;
  assign n3059 = ~\P2_Address_reg[24]/NET0131  & ~\P2_Address_reg[25]/NET0131  ;
  assign n3068 = n3058 & n3059 ;
  assign n3074 = n3067 & n3068 ;
  assign n3064 = ~\P2_Address_reg[7]/NET0131  & ~\P2_Address_reg[8]/NET0131  ;
  assign n3065 = ~\P2_Address_reg[9]/NET0131  & n3064 ;
  assign n3062 = ~\P2_Address_reg[3]/NET0131  & ~\P2_Address_reg[4]/NET0131  ;
  assign n3063 = ~\P2_Address_reg[5]/NET0131  & ~\P2_Address_reg[6]/NET0131  ;
  assign n3066 = n3062 & n3063 ;
  assign n3075 = n3065 & n3066 ;
  assign n3076 = n3074 & n3075 ;
  assign n3051 = ~\P2_Address_reg[0]/NET0131  & ~\P2_Address_reg[10]/NET0131  ;
  assign n3052 = ~\P2_Address_reg[11]/NET0131  & ~\P2_Address_reg[12]/NET0131  ;
  assign n3053 = ~\P2_Address_reg[13]/NET0131  & ~\P2_Address_reg[14]/NET0131  ;
  assign n3071 = n3052 & n3053 ;
  assign n3072 = n3051 & n3071 ;
  assign n3056 = ~\P2_Address_reg[19]/NET0131  & ~\P2_Address_reg[1]/NET0131  ;
  assign n3057 = ~\P2_Address_reg[20]/NET0131  & ~\P2_Address_reg[21]/NET0131  ;
  assign n3069 = n3056 & n3057 ;
  assign n3054 = ~\P2_Address_reg[15]/NET0131  & ~\P2_Address_reg[16]/NET0131  ;
  assign n3055 = ~\P2_Address_reg[17]/NET0131  & ~\P2_Address_reg[18]/NET0131  ;
  assign n3070 = n3054 & n3055 ;
  assign n3073 = n3069 & n3070 ;
  assign n3077 = n3072 & n3073 ;
  assign n3078 = n3076 & n3077 ;
  assign n3079 = \P2_Address_reg[29]/NET0131  & ~n3078 ;
  assign n3092 = \buf2_reg[28]/NET0131  & ~n3079 ;
  assign n3093 = \buf1_reg[28]/NET0131  & n3079 ;
  assign n3094 = ~n3092 & ~n3093 ;
  assign n3095 = n3091 & ~n3094 ;
  assign n3096 = \P2_InstQueueWr_Addr_reg[0]/NET0131  & ~\P2_InstQueueWr_Addr_reg[1]/NET0131  ;
  assign n3097 = ~\P2_InstQueueWr_Addr_reg[2]/NET0131  & n3096 ;
  assign n3098 = \P2_InstQueueWr_Addr_reg[3]/NET0131  & n3097 ;
  assign n3099 = \buf2_reg[20]/NET0131  & ~n3079 ;
  assign n3100 = \buf1_reg[20]/NET0131  & n3079 ;
  assign n3101 = ~n3099 & ~n3100 ;
  assign n3102 = n3098 & ~n3101 ;
  assign n3103 = ~n3095 & ~n3102 ;
  assign n3104 = \P2_DataWidth_reg[1]/NET0131  & ~n3103 ;
  assign n3044 = ~\P2_InstQueueWr_Addr_reg[0]/NET0131  & \P2_InstQueueWr_Addr_reg[1]/NET0131  ;
  assign n3045 = ~\P2_InstQueueWr_Addr_reg[2]/NET0131  & n3044 ;
  assign n3046 = \P2_InstQueueWr_Addr_reg[3]/NET0131  & n3045 ;
  assign n3047 = \P2_InstQueueWr_Addr_reg[0]/NET0131  & \P2_InstQueueWr_Addr_reg[1]/NET0131  ;
  assign n3048 = ~\P2_InstQueueWr_Addr_reg[2]/NET0131  & n3047 ;
  assign n3049 = \P2_InstQueueWr_Addr_reg[3]/NET0131  & n3048 ;
  assign n3050 = ~n3046 & ~n3049 ;
  assign n3080 = \buf2_reg[4]/NET0131  & ~n3079 ;
  assign n3081 = \buf1_reg[4]/NET0131  & n3079 ;
  assign n3082 = ~n3080 & ~n3081 ;
  assign n3083 = ~n3050 & ~n3082 ;
  assign n3084 = \P2_InstQueue_reg[11][4]/NET0131  & ~n3049 ;
  assign n3085 = ~n3046 & n3084 ;
  assign n3086 = ~n3083 & ~n3085 ;
  assign n3105 = ~n3091 & ~n3098 ;
  assign n3106 = \P2_DataWidth_reg[1]/NET0131  & ~n3105 ;
  assign n3107 = ~n3086 & ~n3106 ;
  assign n3108 = ~n3104 & ~n3107 ;
  assign n3109 = n1931 & ~n3108 ;
  assign n3087 = n1926 & n1935 ;
  assign n3088 = ~n3086 & n3087 ;
  assign n3110 = ~n1688 & n3049 ;
  assign n3111 = ~n3084 & ~n3110 ;
  assign n3112 = n3040 & ~n3111 ;
  assign n3113 = n1935 & n2985 ;
  assign n3114 = ~n1934 & ~n3113 ;
  assign n3115 = ~n2987 & n3114 ;
  assign n3116 = ~n1927 & ~n2979 ;
  assign n3117 = ~n3035 & n3116 ;
  assign n3118 = n3115 & n3117 ;
  assign n3119 = \P2_InstQueue_reg[11][4]/NET0131  & ~n3118 ;
  assign n3120 = ~n3112 & ~n3119 ;
  assign n3121 = ~n3088 & n3120 ;
  assign n3122 = ~n3109 & n3121 ;
  assign n3126 = \buf2_reg[7]/NET0131  & ~n3079 ;
  assign n3127 = \buf1_reg[7]/NET0131  & n3079 ;
  assign n3128 = ~n3126 & ~n3127 ;
  assign n3129 = ~n3050 & ~n3128 ;
  assign n3130 = \P2_InstQueue_reg[11][7]/NET0131  & ~n3049 ;
  assign n3131 = ~n3046 & n3130 ;
  assign n3132 = ~n3129 & ~n3131 ;
  assign n3124 = ~n3087 & n3106 ;
  assign n3125 = ~n1931 & ~n3087 ;
  assign n3133 = ~n3124 & ~n3125 ;
  assign n3134 = ~n3132 & n3133 ;
  assign n3135 = ~n1656 & n3049 ;
  assign n3136 = ~n3130 & ~n3135 ;
  assign n3137 = n3040 & ~n3136 ;
  assign n3123 = \P2_InstQueue_reg[11][7]/NET0131  & ~n3118 ;
  assign n3138 = \buf2_reg[23]/NET0131  & ~n3079 ;
  assign n3139 = \buf1_reg[23]/NET0131  & n3079 ;
  assign n3140 = ~n3138 & ~n3139 ;
  assign n3141 = n3034 & n3098 ;
  assign n3142 = ~n3140 & n3141 ;
  assign n3143 = ~n3123 & ~n3142 ;
  assign n3144 = ~n3137 & n3143 ;
  assign n3145 = ~n3134 & n3144 ;
  assign n3148 = \P1_DataWidth_reg[1]/NET0131  & n2436 ;
  assign n3146 = ~n2431 & ~n2440 ;
  assign n3147 = ~n2317 & n2441 ;
  assign n3149 = n3146 & ~n3147 ;
  assign n3150 = ~n3148 & n3149 ;
  assign n3151 = ~n3025 & n3150 ;
  assign n3161 = \P2_InstQueueWr_Addr_reg[2]/NET0131  & n3096 ;
  assign n3162 = \P2_InstQueueWr_Addr_reg[3]/NET0131  & n3161 ;
  assign n3163 = ~n3094 & n3162 ;
  assign n3164 = \P2_InstQueueWr_Addr_reg[2]/NET0131  & n3044 ;
  assign n3165 = \P2_InstQueueWr_Addr_reg[3]/NET0131  & n3164 ;
  assign n3166 = ~n3101 & n3165 ;
  assign n3167 = ~n3163 & ~n3166 ;
  assign n3168 = \P2_DataWidth_reg[1]/NET0131  & ~n3167 ;
  assign n3152 = ~\P2_InstQueueWr_Addr_reg[3]/NET0131  & n3090 ;
  assign n3153 = \P2_InstQueueWr_Addr_reg[2]/NET0131  & n3047 ;
  assign n3154 = \P2_InstQueueWr_Addr_reg[3]/NET0131  & n3153 ;
  assign n3155 = ~n3152 & ~n3154 ;
  assign n3156 = ~n3082 & ~n3155 ;
  assign n3157 = \P2_InstQueue_reg[0][4]/NET0131  & ~n3152 ;
  assign n3158 = ~n3154 & n3157 ;
  assign n3159 = ~n3156 & ~n3158 ;
  assign n3169 = ~n3162 & ~n3165 ;
  assign n3170 = \P2_DataWidth_reg[1]/NET0131  & ~n3169 ;
  assign n3171 = ~n3159 & ~n3170 ;
  assign n3172 = ~n3168 & ~n3171 ;
  assign n3173 = n1931 & ~n3172 ;
  assign n3160 = n3087 & ~n3159 ;
  assign n3174 = ~n1688 & n3152 ;
  assign n3175 = ~n3157 & ~n3174 ;
  assign n3176 = n3040 & ~n3175 ;
  assign n3177 = \P2_InstQueue_reg[0][4]/NET0131  & ~n3118 ;
  assign n3178 = ~n3176 & ~n3177 ;
  assign n3179 = ~n3160 & n3178 ;
  assign n3180 = ~n3173 & n3179 ;
  assign n3183 = ~n3128 & ~n3155 ;
  assign n3184 = \P2_InstQueue_reg[0][7]/NET0131  & ~n3152 ;
  assign n3185 = ~n3154 & n3184 ;
  assign n3186 = ~n3183 & ~n3185 ;
  assign n3182 = ~n3087 & n3170 ;
  assign n3187 = ~n3125 & ~n3182 ;
  assign n3188 = ~n3186 & n3187 ;
  assign n3189 = ~n1656 & n3152 ;
  assign n3190 = ~n3184 & ~n3189 ;
  assign n3191 = n3040 & ~n3190 ;
  assign n3181 = \P2_InstQueue_reg[0][7]/NET0131  & ~n3118 ;
  assign n3192 = n3034 & n3165 ;
  assign n3193 = ~n3140 & n3192 ;
  assign n3194 = ~n3181 & ~n3193 ;
  assign n3195 = ~n3191 & n3194 ;
  assign n3196 = ~n3188 & n3195 ;
  assign n3202 = ~n3046 & ~n3098 ;
  assign n3203 = ~n3128 & ~n3202 ;
  assign n3204 = \P2_InstQueue_reg[10][7]/NET0131  & ~n3046 ;
  assign n3205 = ~n3098 & n3204 ;
  assign n3206 = ~n3203 & ~n3205 ;
  assign n3198 = ~\P2_InstQueueWr_Addr_reg[3]/NET0131  & n3153 ;
  assign n3199 = ~n3091 & ~n3198 ;
  assign n3200 = \P2_DataWidth_reg[1]/NET0131  & ~n3199 ;
  assign n3201 = ~n3087 & n3200 ;
  assign n3207 = ~n3125 & ~n3201 ;
  assign n3208 = ~n3206 & n3207 ;
  assign n3209 = ~n1656 & n3046 ;
  assign n3210 = ~n3204 & ~n3209 ;
  assign n3211 = n3040 & ~n3210 ;
  assign n3197 = \P2_InstQueue_reg[10][7]/NET0131  & ~n3118 ;
  assign n3212 = n3034 & n3091 ;
  assign n3213 = ~n3140 & n3212 ;
  assign n3214 = ~n3197 & ~n3213 ;
  assign n3215 = ~n3211 & n3214 ;
  assign n3216 = ~n3208 & n3215 ;
  assign n3222 = n3091 & ~n3101 ;
  assign n3223 = ~n3094 & n3198 ;
  assign n3224 = ~n3222 & ~n3223 ;
  assign n3225 = \P2_DataWidth_reg[1]/NET0131  & ~n3224 ;
  assign n3217 = ~n3082 & ~n3202 ;
  assign n3218 = \P2_InstQueue_reg[10][4]/NET0131  & ~n3046 ;
  assign n3219 = ~n3098 & n3218 ;
  assign n3220 = ~n3217 & ~n3219 ;
  assign n3226 = ~n3200 & ~n3220 ;
  assign n3227 = ~n3225 & ~n3226 ;
  assign n3228 = n1931 & ~n3227 ;
  assign n3221 = n3087 & ~n3220 ;
  assign n3229 = ~n1688 & n3046 ;
  assign n3230 = ~n3218 & ~n3229 ;
  assign n3231 = n3040 & ~n3230 ;
  assign n3232 = \P2_InstQueue_reg[10][4]/NET0131  & ~n3118 ;
  assign n3233 = ~n3231 & ~n3232 ;
  assign n3234 = ~n3221 & n3233 ;
  assign n3235 = ~n3228 & n3234 ;
  assign n3244 = ~n3094 & n3098 ;
  assign n3245 = n3046 & ~n3101 ;
  assign n3246 = ~n3244 & ~n3245 ;
  assign n3247 = \P2_DataWidth_reg[1]/NET0131  & ~n3246 ;
  assign n3236 = \P2_InstQueueWr_Addr_reg[2]/NET0131  & n3089 ;
  assign n3237 = \P2_InstQueueWr_Addr_reg[3]/NET0131  & n3236 ;
  assign n3238 = ~n3049 & ~n3237 ;
  assign n3239 = ~n3082 & ~n3238 ;
  assign n3240 = \P2_InstQueue_reg[12][4]/NET0131  & ~n3237 ;
  assign n3241 = ~n3049 & n3240 ;
  assign n3242 = ~n3239 & ~n3241 ;
  assign n3248 = \P2_DataWidth_reg[1]/NET0131  & ~n3202 ;
  assign n3249 = ~n3242 & ~n3248 ;
  assign n3250 = ~n3247 & ~n3249 ;
  assign n3251 = n1931 & ~n3250 ;
  assign n3243 = n3087 & ~n3242 ;
  assign n3252 = ~n1688 & n3237 ;
  assign n3253 = ~n3240 & ~n3252 ;
  assign n3254 = n3040 & ~n3253 ;
  assign n3255 = \P2_InstQueue_reg[12][4]/NET0131  & ~n3118 ;
  assign n3256 = ~n3254 & ~n3255 ;
  assign n3257 = ~n3243 & n3256 ;
  assign n3258 = ~n3251 & n3257 ;
  assign n3261 = ~n3128 & ~n3238 ;
  assign n3262 = \P2_InstQueue_reg[12][7]/NET0131  & ~n3237 ;
  assign n3263 = ~n3049 & n3262 ;
  assign n3264 = ~n3261 & ~n3263 ;
  assign n3260 = ~n3087 & n3248 ;
  assign n3265 = ~n3125 & ~n3260 ;
  assign n3266 = ~n3264 & n3265 ;
  assign n3267 = ~n1656 & n3237 ;
  assign n3268 = ~n3262 & ~n3267 ;
  assign n3269 = n3040 & ~n3268 ;
  assign n3259 = \P2_InstQueue_reg[12][7]/NET0131  & ~n3118 ;
  assign n3270 = n3034 & n3046 ;
  assign n3271 = ~n3140 & n3270 ;
  assign n3272 = ~n3259 & ~n3271 ;
  assign n3273 = ~n3269 & n3272 ;
  assign n3274 = ~n3266 & n3273 ;
  assign n3281 = n3046 & ~n3094 ;
  assign n3282 = n3049 & ~n3101 ;
  assign n3283 = ~n3281 & ~n3282 ;
  assign n3284 = \P2_DataWidth_reg[1]/NET0131  & ~n3283 ;
  assign n3275 = ~n3162 & ~n3237 ;
  assign n3276 = ~n3082 & ~n3275 ;
  assign n3277 = \P2_InstQueue_reg[13][4]/NET0131  & ~n3162 ;
  assign n3278 = ~n3237 & n3277 ;
  assign n3279 = ~n3276 & ~n3278 ;
  assign n3285 = \P2_DataWidth_reg[1]/NET0131  & ~n3050 ;
  assign n3286 = ~n3279 & ~n3285 ;
  assign n3287 = ~n3284 & ~n3286 ;
  assign n3288 = n1931 & ~n3287 ;
  assign n3280 = n3087 & ~n3279 ;
  assign n3289 = ~n1688 & n3162 ;
  assign n3290 = ~n3277 & ~n3289 ;
  assign n3291 = n3040 & ~n3290 ;
  assign n3292 = \P2_InstQueue_reg[13][4]/NET0131  & ~n3118 ;
  assign n3293 = ~n3291 & ~n3292 ;
  assign n3294 = ~n3280 & n3293 ;
  assign n3295 = ~n3288 & n3294 ;
  assign n3298 = ~n3128 & ~n3275 ;
  assign n3299 = \P2_InstQueue_reg[13][7]/NET0131  & ~n3162 ;
  assign n3300 = ~n3237 & n3299 ;
  assign n3301 = ~n3298 & ~n3300 ;
  assign n3297 = ~n3087 & n3285 ;
  assign n3302 = ~n3125 & ~n3297 ;
  assign n3303 = ~n3301 & n3302 ;
  assign n3304 = ~n1656 & n3162 ;
  assign n3305 = ~n3299 & ~n3304 ;
  assign n3306 = n3040 & ~n3305 ;
  assign n3296 = \P2_InstQueue_reg[13][7]/NET0131  & ~n3118 ;
  assign n3307 = n3034 & n3049 ;
  assign n3308 = ~n3140 & n3307 ;
  assign n3309 = ~n3296 & ~n3308 ;
  assign n3310 = ~n3306 & n3309 ;
  assign n3311 = ~n3303 & n3310 ;
  assign n3317 = n3049 & ~n3094 ;
  assign n3318 = ~n3101 & n3237 ;
  assign n3319 = ~n3317 & ~n3318 ;
  assign n3320 = \P2_DataWidth_reg[1]/NET0131  & ~n3319 ;
  assign n3312 = ~n3082 & ~n3169 ;
  assign n3313 = \P2_InstQueue_reg[14][4]/NET0131  & ~n3165 ;
  assign n3314 = ~n3162 & n3313 ;
  assign n3315 = ~n3312 & ~n3314 ;
  assign n3321 = \P2_DataWidth_reg[1]/NET0131  & ~n3238 ;
  assign n3322 = ~n3315 & ~n3321 ;
  assign n3323 = ~n3320 & ~n3322 ;
  assign n3324 = n1931 & ~n3323 ;
  assign n3316 = n3087 & ~n3315 ;
  assign n3325 = ~n1688 & n3165 ;
  assign n3326 = ~n3313 & ~n3325 ;
  assign n3327 = n3040 & ~n3326 ;
  assign n3328 = \P2_InstQueue_reg[14][4]/NET0131  & ~n3118 ;
  assign n3329 = ~n3327 & ~n3328 ;
  assign n3330 = ~n3316 & n3329 ;
  assign n3331 = ~n3324 & n3330 ;
  assign n3334 = ~n3128 & ~n3169 ;
  assign n3335 = \P2_InstQueue_reg[14][7]/NET0131  & ~n3165 ;
  assign n3336 = ~n3162 & n3335 ;
  assign n3337 = ~n3334 & ~n3336 ;
  assign n3333 = ~n3087 & n3321 ;
  assign n3338 = ~n3125 & ~n3333 ;
  assign n3339 = ~n3337 & n3338 ;
  assign n3340 = ~n1656 & n3165 ;
  assign n3341 = ~n3335 & ~n3340 ;
  assign n3342 = n3040 & ~n3341 ;
  assign n3332 = \P2_InstQueue_reg[14][7]/NET0131  & ~n3118 ;
  assign n3343 = n3034 & n3237 ;
  assign n3344 = ~n3140 & n3343 ;
  assign n3345 = ~n3332 & ~n3344 ;
  assign n3346 = ~n3342 & n3345 ;
  assign n3347 = ~n3339 & n3346 ;
  assign n3354 = ~n3094 & n3237 ;
  assign n3355 = ~n3101 & n3162 ;
  assign n3356 = ~n3354 & ~n3355 ;
  assign n3357 = \P2_DataWidth_reg[1]/NET0131  & ~n3356 ;
  assign n3348 = ~n3154 & ~n3165 ;
  assign n3349 = ~n3082 & ~n3348 ;
  assign n3350 = \P2_InstQueue_reg[15][4]/NET0131  & ~n3154 ;
  assign n3351 = ~n3165 & n3350 ;
  assign n3352 = ~n3349 & ~n3351 ;
  assign n3358 = \P2_DataWidth_reg[1]/NET0131  & ~n3275 ;
  assign n3359 = ~n3352 & ~n3358 ;
  assign n3360 = ~n3357 & ~n3359 ;
  assign n3361 = n1931 & ~n3360 ;
  assign n3353 = n3087 & ~n3352 ;
  assign n3362 = ~n1688 & n3154 ;
  assign n3363 = ~n3350 & ~n3362 ;
  assign n3364 = n3040 & ~n3363 ;
  assign n3365 = \P2_InstQueue_reg[15][4]/NET0131  & ~n3118 ;
  assign n3366 = ~n3364 & ~n3365 ;
  assign n3367 = ~n3353 & n3366 ;
  assign n3368 = ~n3361 & n3367 ;
  assign n3371 = ~n3128 & ~n3348 ;
  assign n3372 = \P2_InstQueue_reg[15][7]/NET0131  & ~n3154 ;
  assign n3373 = ~n3165 & n3372 ;
  assign n3374 = ~n3371 & ~n3373 ;
  assign n3370 = ~n3087 & n3358 ;
  assign n3375 = ~n3125 & ~n3370 ;
  assign n3376 = ~n3374 & n3375 ;
  assign n3377 = ~n1656 & n3154 ;
  assign n3378 = ~n3372 & ~n3377 ;
  assign n3379 = n3040 & ~n3378 ;
  assign n3369 = \P2_InstQueue_reg[15][7]/NET0131  & ~n3118 ;
  assign n3380 = n3034 & n3162 ;
  assign n3381 = ~n3140 & n3380 ;
  assign n3382 = ~n3369 & ~n3381 ;
  assign n3383 = ~n3379 & n3382 ;
  assign n3384 = ~n3376 & n3383 ;
  assign n3388 = ~\P2_InstQueueWr_Addr_reg[3]/NET0131  & n3097 ;
  assign n3389 = ~n3152 & ~n3388 ;
  assign n3390 = ~n3128 & ~n3389 ;
  assign n3391 = \P2_InstQueue_reg[1][7]/NET0131  & ~n3388 ;
  assign n3392 = ~n3152 & n3391 ;
  assign n3393 = ~n3390 & ~n3392 ;
  assign n3386 = \P2_DataWidth_reg[1]/NET0131  & ~n3348 ;
  assign n3387 = ~n3087 & n3386 ;
  assign n3394 = ~n3125 & ~n3387 ;
  assign n3395 = ~n3393 & n3394 ;
  assign n3396 = ~n1656 & n3388 ;
  assign n3397 = ~n3391 & ~n3396 ;
  assign n3398 = n3040 & ~n3397 ;
  assign n3385 = \P2_InstQueue_reg[1][7]/NET0131  & ~n3118 ;
  assign n3399 = n3034 & n3154 ;
  assign n3400 = ~n3140 & n3399 ;
  assign n3401 = ~n3385 & ~n3400 ;
  assign n3402 = ~n3398 & n3401 ;
  assign n3403 = ~n3395 & n3402 ;
  assign n3409 = ~n3094 & n3165 ;
  assign n3410 = ~n3101 & n3154 ;
  assign n3411 = ~n3409 & ~n3410 ;
  assign n3412 = \P2_DataWidth_reg[1]/NET0131  & ~n3411 ;
  assign n3404 = ~n3082 & ~n3389 ;
  assign n3405 = \P2_InstQueue_reg[1][4]/NET0131  & ~n3388 ;
  assign n3406 = ~n3152 & n3405 ;
  assign n3407 = ~n3404 & ~n3406 ;
  assign n3413 = ~n3386 & ~n3407 ;
  assign n3414 = ~n3412 & ~n3413 ;
  assign n3415 = n1931 & ~n3414 ;
  assign n3408 = n3087 & ~n3407 ;
  assign n3416 = ~n1688 & n3388 ;
  assign n3417 = ~n3405 & ~n3416 ;
  assign n3418 = n3040 & ~n3417 ;
  assign n3419 = \P2_InstQueue_reg[1][4]/NET0131  & ~n3118 ;
  assign n3420 = ~n3418 & ~n3419 ;
  assign n3421 = ~n3408 & n3420 ;
  assign n3422 = ~n3415 & n3421 ;
  assign n3430 = ~n3101 & n3152 ;
  assign n3431 = ~n3094 & n3154 ;
  assign n3432 = ~n3430 & ~n3431 ;
  assign n3433 = \P2_DataWidth_reg[1]/NET0131  & ~n3432 ;
  assign n3423 = ~\P2_InstQueueWr_Addr_reg[3]/NET0131  & n3045 ;
  assign n3424 = ~n3388 & ~n3423 ;
  assign n3425 = ~n3082 & ~n3424 ;
  assign n3426 = \P2_InstQueue_reg[2][4]/NET0131  & ~n3423 ;
  assign n3427 = ~n3388 & n3426 ;
  assign n3428 = ~n3425 & ~n3427 ;
  assign n3434 = \P2_DataWidth_reg[1]/NET0131  & ~n3155 ;
  assign n3435 = ~n3428 & ~n3434 ;
  assign n3436 = ~n3433 & ~n3435 ;
  assign n3437 = n1931 & ~n3436 ;
  assign n3429 = n3087 & ~n3428 ;
  assign n3438 = ~n1688 & n3423 ;
  assign n3439 = ~n3426 & ~n3438 ;
  assign n3440 = n3040 & ~n3439 ;
  assign n3441 = \P2_InstQueue_reg[2][4]/NET0131  & ~n3118 ;
  assign n3442 = ~n3440 & ~n3441 ;
  assign n3443 = ~n3429 & n3442 ;
  assign n3444 = ~n3437 & n3443 ;
  assign n3447 = ~n3128 & ~n3424 ;
  assign n3448 = \P2_InstQueue_reg[2][7]/NET0131  & ~n3423 ;
  assign n3449 = ~n3388 & n3448 ;
  assign n3450 = ~n3447 & ~n3449 ;
  assign n3446 = ~n3087 & n3434 ;
  assign n3451 = ~n3125 & ~n3446 ;
  assign n3452 = ~n3450 & n3451 ;
  assign n3453 = ~n1656 & n3423 ;
  assign n3454 = ~n3448 & ~n3453 ;
  assign n3455 = n3040 & ~n3454 ;
  assign n3445 = \P2_InstQueue_reg[2][7]/NET0131  & ~n3118 ;
  assign n3456 = n3034 & n3152 ;
  assign n3457 = ~n3140 & n3456 ;
  assign n3458 = ~n3445 & ~n3457 ;
  assign n3459 = ~n3455 & n3458 ;
  assign n3460 = ~n3452 & n3459 ;
  assign n3468 = ~n3094 & n3152 ;
  assign n3469 = ~n3101 & n3388 ;
  assign n3470 = ~n3468 & ~n3469 ;
  assign n3471 = \P2_DataWidth_reg[1]/NET0131  & ~n3470 ;
  assign n3461 = ~\P2_InstQueueWr_Addr_reg[3]/NET0131  & n3048 ;
  assign n3462 = ~n3423 & ~n3461 ;
  assign n3463 = ~n3082 & ~n3462 ;
  assign n3464 = \P2_InstQueue_reg[3][4]/NET0131  & ~n3461 ;
  assign n3465 = ~n3423 & n3464 ;
  assign n3466 = ~n3463 & ~n3465 ;
  assign n3472 = \P2_DataWidth_reg[1]/NET0131  & ~n3389 ;
  assign n3473 = ~n3466 & ~n3472 ;
  assign n3474 = ~n3471 & ~n3473 ;
  assign n3475 = n1931 & ~n3474 ;
  assign n3467 = n3087 & ~n3466 ;
  assign n3476 = ~n1688 & n3461 ;
  assign n3477 = ~n3464 & ~n3476 ;
  assign n3478 = n3040 & ~n3477 ;
  assign n3479 = \P2_InstQueue_reg[3][4]/NET0131  & ~n3118 ;
  assign n3480 = ~n3478 & ~n3479 ;
  assign n3481 = ~n3467 & n3480 ;
  assign n3482 = ~n3475 & n3481 ;
  assign n3485 = ~n3128 & ~n3462 ;
  assign n3486 = \P2_InstQueue_reg[3][7]/NET0131  & ~n3461 ;
  assign n3487 = ~n3423 & n3486 ;
  assign n3488 = ~n3485 & ~n3487 ;
  assign n3484 = ~n3087 & n3472 ;
  assign n3489 = ~n3125 & ~n3484 ;
  assign n3490 = ~n3488 & n3489 ;
  assign n3491 = ~n1656 & n3461 ;
  assign n3492 = ~n3486 & ~n3491 ;
  assign n3493 = n3040 & ~n3492 ;
  assign n3483 = \P2_InstQueue_reg[3][7]/NET0131  & ~n3118 ;
  assign n3494 = n3034 & n3388 ;
  assign n3495 = ~n3140 & n3494 ;
  assign n3496 = ~n3483 & ~n3495 ;
  assign n3497 = ~n3493 & n3496 ;
  assign n3498 = ~n3490 & n3497 ;
  assign n3506 = ~n3094 & n3388 ;
  assign n3507 = ~n3101 & n3423 ;
  assign n3508 = ~n3506 & ~n3507 ;
  assign n3509 = \P2_DataWidth_reg[1]/NET0131  & ~n3508 ;
  assign n3499 = ~\P2_InstQueueWr_Addr_reg[3]/NET0131  & n3236 ;
  assign n3500 = ~n3461 & ~n3499 ;
  assign n3501 = ~n3082 & ~n3500 ;
  assign n3502 = \P2_InstQueue_reg[4][4]/NET0131  & ~n3499 ;
  assign n3503 = ~n3461 & n3502 ;
  assign n3504 = ~n3501 & ~n3503 ;
  assign n3510 = \P2_DataWidth_reg[1]/NET0131  & ~n3424 ;
  assign n3511 = ~n3504 & ~n3510 ;
  assign n3512 = ~n3509 & ~n3511 ;
  assign n3513 = n1931 & ~n3512 ;
  assign n3505 = n3087 & ~n3504 ;
  assign n3514 = ~n1688 & n3499 ;
  assign n3515 = ~n3502 & ~n3514 ;
  assign n3516 = n3040 & ~n3515 ;
  assign n3517 = \P2_InstQueue_reg[4][4]/NET0131  & ~n3118 ;
  assign n3518 = ~n3516 & ~n3517 ;
  assign n3519 = ~n3505 & n3518 ;
  assign n3520 = ~n3513 & n3519 ;
  assign n3523 = ~n3128 & ~n3500 ;
  assign n3524 = \P2_InstQueue_reg[4][7]/NET0131  & ~n3499 ;
  assign n3525 = ~n3461 & n3524 ;
  assign n3526 = ~n3523 & ~n3525 ;
  assign n3522 = ~n3087 & n3510 ;
  assign n3527 = ~n3125 & ~n3522 ;
  assign n3528 = ~n3526 & n3527 ;
  assign n3529 = ~n1656 & n3499 ;
  assign n3530 = ~n3524 & ~n3529 ;
  assign n3531 = n3040 & ~n3530 ;
  assign n3521 = \P2_InstQueue_reg[4][7]/NET0131  & ~n3118 ;
  assign n3532 = n3034 & n3423 ;
  assign n3533 = ~n3140 & n3532 ;
  assign n3534 = ~n3521 & ~n3533 ;
  assign n3535 = ~n3531 & n3534 ;
  assign n3536 = ~n3528 & n3535 ;
  assign n3544 = ~n3094 & n3423 ;
  assign n3545 = ~n3101 & n3461 ;
  assign n3546 = ~n3544 & ~n3545 ;
  assign n3547 = \P2_DataWidth_reg[1]/NET0131  & ~n3546 ;
  assign n3537 = ~\P2_InstQueueWr_Addr_reg[3]/NET0131  & n3161 ;
  assign n3538 = ~n3499 & ~n3537 ;
  assign n3539 = ~n3082 & ~n3538 ;
  assign n3540 = \P2_InstQueue_reg[5][4]/NET0131  & ~n3537 ;
  assign n3541 = ~n3499 & n3540 ;
  assign n3542 = ~n3539 & ~n3541 ;
  assign n3548 = \P2_DataWidth_reg[1]/NET0131  & ~n3462 ;
  assign n3549 = ~n3542 & ~n3548 ;
  assign n3550 = ~n3547 & ~n3549 ;
  assign n3551 = n1931 & ~n3550 ;
  assign n3543 = n3087 & ~n3542 ;
  assign n3552 = ~n1688 & n3537 ;
  assign n3553 = ~n3540 & ~n3552 ;
  assign n3554 = n3040 & ~n3553 ;
  assign n3555 = \P2_InstQueue_reg[5][4]/NET0131  & ~n3118 ;
  assign n3556 = ~n3554 & ~n3555 ;
  assign n3557 = ~n3543 & n3556 ;
  assign n3558 = ~n3551 & n3557 ;
  assign n3561 = ~n3128 & ~n3538 ;
  assign n3562 = \P2_InstQueue_reg[5][7]/NET0131  & ~n3537 ;
  assign n3563 = ~n3499 & n3562 ;
  assign n3564 = ~n3561 & ~n3563 ;
  assign n3560 = ~n3087 & n3548 ;
  assign n3565 = ~n3125 & ~n3560 ;
  assign n3566 = ~n3564 & n3565 ;
  assign n3567 = ~n1656 & n3537 ;
  assign n3568 = ~n3562 & ~n3567 ;
  assign n3569 = n3040 & ~n3568 ;
  assign n3559 = \P2_InstQueue_reg[5][7]/NET0131  & ~n3118 ;
  assign n3570 = n3034 & n3461 ;
  assign n3571 = ~n3140 & n3570 ;
  assign n3572 = ~n3559 & ~n3571 ;
  assign n3573 = ~n3569 & n3572 ;
  assign n3574 = ~n3566 & n3573 ;
  assign n3582 = ~n3094 & n3461 ;
  assign n3583 = ~n3101 & n3499 ;
  assign n3584 = ~n3582 & ~n3583 ;
  assign n3585 = \P2_DataWidth_reg[1]/NET0131  & ~n3584 ;
  assign n3575 = ~\P2_InstQueueWr_Addr_reg[3]/NET0131  & n3164 ;
  assign n3576 = ~n3537 & ~n3575 ;
  assign n3577 = ~n3082 & ~n3576 ;
  assign n3578 = \P2_InstQueue_reg[6][4]/NET0131  & ~n3575 ;
  assign n3579 = ~n3537 & n3578 ;
  assign n3580 = ~n3577 & ~n3579 ;
  assign n3586 = \P2_DataWidth_reg[1]/NET0131  & ~n3500 ;
  assign n3587 = ~n3580 & ~n3586 ;
  assign n3588 = ~n3585 & ~n3587 ;
  assign n3589 = n1931 & ~n3588 ;
  assign n3581 = n3087 & ~n3580 ;
  assign n3590 = ~n1688 & n3575 ;
  assign n3591 = ~n3578 & ~n3590 ;
  assign n3592 = n3040 & ~n3591 ;
  assign n3593 = \P2_InstQueue_reg[6][4]/NET0131  & ~n3118 ;
  assign n3594 = ~n3592 & ~n3593 ;
  assign n3595 = ~n3581 & n3594 ;
  assign n3596 = ~n3589 & n3595 ;
  assign n3599 = ~n3128 & ~n3576 ;
  assign n3600 = \P2_InstQueue_reg[6][7]/NET0131  & ~n3575 ;
  assign n3601 = ~n3537 & n3600 ;
  assign n3602 = ~n3599 & ~n3601 ;
  assign n3598 = ~n3087 & n3586 ;
  assign n3603 = ~n3125 & ~n3598 ;
  assign n3604 = ~n3602 & n3603 ;
  assign n3605 = ~n1656 & n3575 ;
  assign n3606 = ~n3600 & ~n3605 ;
  assign n3607 = n3040 & ~n3606 ;
  assign n3597 = \P2_InstQueue_reg[6][7]/NET0131  & ~n3118 ;
  assign n3608 = n3034 & n3499 ;
  assign n3609 = ~n3140 & n3608 ;
  assign n3610 = ~n3597 & ~n3609 ;
  assign n3611 = ~n3607 & n3610 ;
  assign n3612 = ~n3604 & n3611 ;
  assign n3619 = ~n3094 & n3499 ;
  assign n3620 = ~n3101 & n3537 ;
  assign n3621 = ~n3619 & ~n3620 ;
  assign n3622 = \P2_DataWidth_reg[1]/NET0131  & ~n3621 ;
  assign n3613 = ~n3198 & ~n3575 ;
  assign n3614 = ~n3082 & ~n3613 ;
  assign n3615 = \P2_InstQueue_reg[7][4]/NET0131  & ~n3198 ;
  assign n3616 = ~n3575 & n3615 ;
  assign n3617 = ~n3614 & ~n3616 ;
  assign n3623 = \P2_DataWidth_reg[1]/NET0131  & ~n3538 ;
  assign n3624 = ~n3617 & ~n3623 ;
  assign n3625 = ~n3622 & ~n3624 ;
  assign n3626 = n1931 & ~n3625 ;
  assign n3618 = n3087 & ~n3617 ;
  assign n3627 = ~n1688 & n3198 ;
  assign n3628 = ~n3615 & ~n3627 ;
  assign n3629 = n3040 & ~n3628 ;
  assign n3630 = \P2_InstQueue_reg[7][4]/NET0131  & ~n3118 ;
  assign n3631 = ~n3629 & ~n3630 ;
  assign n3632 = ~n3618 & n3631 ;
  assign n3633 = ~n3626 & n3632 ;
  assign n3636 = ~n3128 & ~n3613 ;
  assign n3637 = \P2_InstQueue_reg[7][7]/NET0131  & ~n3198 ;
  assign n3638 = ~n3575 & n3637 ;
  assign n3639 = ~n3636 & ~n3638 ;
  assign n3635 = ~n3087 & n3623 ;
  assign n3640 = ~n3125 & ~n3635 ;
  assign n3641 = ~n3639 & n3640 ;
  assign n3642 = ~n1656 & n3198 ;
  assign n3643 = ~n3637 & ~n3642 ;
  assign n3644 = n3040 & ~n3643 ;
  assign n3634 = \P2_InstQueue_reg[7][7]/NET0131  & ~n3118 ;
  assign n3645 = n3034 & n3537 ;
  assign n3646 = ~n3140 & n3645 ;
  assign n3647 = ~n3634 & ~n3646 ;
  assign n3648 = ~n3644 & n3647 ;
  assign n3649 = ~n3641 & n3648 ;
  assign n3655 = ~n3094 & n3537 ;
  assign n3656 = ~n3101 & n3575 ;
  assign n3657 = ~n3655 & ~n3656 ;
  assign n3658 = \P2_DataWidth_reg[1]/NET0131  & ~n3657 ;
  assign n3650 = ~n3082 & ~n3199 ;
  assign n3651 = \P2_InstQueue_reg[8][4]/NET0131  & ~n3091 ;
  assign n3652 = ~n3198 & n3651 ;
  assign n3653 = ~n3650 & ~n3652 ;
  assign n3659 = \P2_DataWidth_reg[1]/NET0131  & ~n3576 ;
  assign n3660 = ~n3653 & ~n3659 ;
  assign n3661 = ~n3658 & ~n3660 ;
  assign n3662 = n1931 & ~n3661 ;
  assign n3654 = n3087 & ~n3653 ;
  assign n3663 = ~n1688 & n3091 ;
  assign n3664 = ~n3651 & ~n3663 ;
  assign n3665 = n3040 & ~n3664 ;
  assign n3666 = \P2_InstQueue_reg[8][4]/NET0131  & ~n3118 ;
  assign n3667 = ~n3665 & ~n3666 ;
  assign n3668 = ~n3654 & n3667 ;
  assign n3669 = ~n3662 & n3668 ;
  assign n3672 = ~n3128 & ~n3199 ;
  assign n3673 = \P2_InstQueue_reg[8][7]/NET0131  & ~n3091 ;
  assign n3674 = ~n3198 & n3673 ;
  assign n3675 = ~n3672 & ~n3674 ;
  assign n3671 = ~n3087 & n3659 ;
  assign n3676 = ~n3125 & ~n3671 ;
  assign n3677 = ~n3675 & n3676 ;
  assign n3678 = ~n1656 & n3091 ;
  assign n3679 = ~n3673 & ~n3678 ;
  assign n3680 = n3040 & ~n3679 ;
  assign n3670 = \P2_InstQueue_reg[8][7]/NET0131  & ~n3118 ;
  assign n3681 = n3034 & n3575 ;
  assign n3682 = ~n3140 & n3681 ;
  assign n3683 = ~n3670 & ~n3682 ;
  assign n3684 = ~n3680 & n3683 ;
  assign n3685 = ~n3677 & n3684 ;
  assign n3691 = ~n3094 & n3575 ;
  assign n3692 = ~n3101 & n3198 ;
  assign n3693 = ~n3691 & ~n3692 ;
  assign n3694 = \P2_DataWidth_reg[1]/NET0131  & ~n3693 ;
  assign n3686 = ~n3082 & ~n3105 ;
  assign n3687 = \P2_InstQueue_reg[9][4]/NET0131  & ~n3098 ;
  assign n3688 = ~n3091 & n3687 ;
  assign n3689 = ~n3686 & ~n3688 ;
  assign n3695 = \P2_DataWidth_reg[1]/NET0131  & ~n3613 ;
  assign n3696 = ~n3689 & ~n3695 ;
  assign n3697 = ~n3694 & ~n3696 ;
  assign n3698 = n1931 & ~n3697 ;
  assign n3690 = n3087 & ~n3689 ;
  assign n3699 = ~n1688 & n3098 ;
  assign n3700 = ~n3687 & ~n3699 ;
  assign n3701 = n3040 & ~n3700 ;
  assign n3702 = \P2_InstQueue_reg[9][4]/NET0131  & ~n3118 ;
  assign n3703 = ~n3701 & ~n3702 ;
  assign n3704 = ~n3690 & n3703 ;
  assign n3705 = ~n3698 & n3704 ;
  assign n3708 = ~n3105 & ~n3128 ;
  assign n3709 = \P2_InstQueue_reg[9][7]/NET0131  & ~n3098 ;
  assign n3710 = ~n3091 & n3709 ;
  assign n3711 = ~n3708 & ~n3710 ;
  assign n3707 = ~n3087 & n3695 ;
  assign n3712 = ~n3125 & ~n3707 ;
  assign n3713 = ~n3711 & n3712 ;
  assign n3714 = ~n1656 & n3098 ;
  assign n3715 = ~n3709 & ~n3714 ;
  assign n3716 = n3040 & ~n3715 ;
  assign n3706 = \P2_InstQueue_reg[9][7]/NET0131  & ~n3118 ;
  assign n3717 = n3034 & n3198 ;
  assign n3718 = ~n3140 & n3717 ;
  assign n3719 = ~n3706 & ~n3718 ;
  assign n3720 = ~n3716 & n3719 ;
  assign n3721 = ~n3713 & n3720 ;
  assign n3722 = \P3_InstAddrPointer_reg[31]/NET0131  & n2896 ;
  assign n4115 = \P3_InstAddrPointer_reg[27]/NET0131  & \P3_InstAddrPointer_reg[28]/NET0131  ;
  assign n4116 = \P3_InstAddrPointer_reg[29]/NET0131  & n4115 ;
  assign n4123 = \P3_InstAddrPointer_reg[30]/NET0131  & n4116 ;
  assign n3756 = \P3_InstAddrPointer_reg[15]/NET0131  & \P3_InstAddrPointer_reg[16]/NET0131  ;
  assign n3757 = \P3_InstAddrPointer_reg[17]/NET0131  & n3756 ;
  assign n3754 = \P3_InstAddrPointer_reg[18]/NET0131  & \P3_InstAddrPointer_reg[19]/NET0131  ;
  assign n3755 = \P3_InstAddrPointer_reg[20]/NET0131  & n3754 ;
  assign n3758 = \P3_InstAddrPointer_reg[14]/NET0131  & \P3_InstAddrPointer_reg[21]/NET0131  ;
  assign n3759 = n3755 & n3758 ;
  assign n3760 = n3757 & n3759 ;
  assign n4094 = \P3_InstAddrPointer_reg[22]/NET0131  & n3760 ;
  assign n3761 = \P3_InstAddrPointer_reg[1]/NET0131  & \P3_InstAddrPointer_reg[2]/NET0131  ;
  assign n3762 = \P3_InstAddrPointer_reg[3]/NET0131  & n3761 ;
  assign n3763 = \P3_InstAddrPointer_reg[4]/NET0131  & n3762 ;
  assign n3764 = \P3_InstAddrPointer_reg[5]/NET0131  & n3763 ;
  assign n3765 = \P3_InstAddrPointer_reg[6]/NET0131  & n3764 ;
  assign n3766 = \P3_InstAddrPointer_reg[7]/NET0131  & n3765 ;
  assign n3777 = \P3_InstAddrPointer_reg[8]/NET0131  & \P3_InstAddrPointer_reg[9]/NET0131  ;
  assign n3778 = n3766 & n3777 ;
  assign n3779 = \P3_InstAddrPointer_reg[10]/NET0131  & \P3_InstAddrPointer_reg[11]/NET0131  ;
  assign n3780 = n3778 & n3779 ;
  assign n3781 = \P3_InstAddrPointer_reg[12]/NET0131  & \P3_InstAddrPointer_reg[13]/NET0131  ;
  assign n4095 = n3780 & n3781 ;
  assign n4096 = n4094 & n4095 ;
  assign n4088 = \P3_InstAddrPointer_reg[23]/NET0131  & \P3_InstAddrPointer_reg[24]/NET0131  ;
  assign n4089 = \P3_InstAddrPointer_reg[25]/NET0131  & n4088 ;
  assign n4108 = \P3_InstAddrPointer_reg[26]/NET0131  & n4089 ;
  assign n4109 = n4096 & n4108 ;
  assign n4132 = \P3_InstAddrPointer_reg[0]/NET0131  & n4109 ;
  assign n4133 = n4123 & n4132 ;
  assign n4134 = \P3_InstAddrPointer_reg[31]/NET0131  & ~n4133 ;
  assign n4124 = n4109 & n4123 ;
  assign n4126 = ~\P3_InstAddrPointer_reg[31]/NET0131  & n4124 ;
  assign n4135 = \P3_InstAddrPointer_reg[0]/NET0131  & n4126 ;
  assign n4136 = ~n4134 & ~n4135 ;
  assign n4137 = ~\P3_InstAddrPointer_reg[27]/NET0131  & ~n4132 ;
  assign n4138 = \P3_InstAddrPointer_reg[27]/NET0131  & n4132 ;
  assign n4139 = ~n4137 & ~n4138 ;
  assign n4140 = ~\P3_InstAddrPointer_reg[28]/NET0131  & ~n4138 ;
  assign n4141 = n4115 & n4132 ;
  assign n4142 = ~n4140 & ~n4141 ;
  assign n4143 = ~n4139 & ~n4142 ;
  assign n4144 = ~\P3_InstAddrPointer_reg[29]/NET0131  & ~n4141 ;
  assign n4145 = n4116 & n4132 ;
  assign n4146 = ~n4144 & ~n4145 ;
  assign n4147 = n4143 & ~n4146 ;
  assign n3767 = \P3_InstAddrPointer_reg[8]/NET0131  & n3766 ;
  assign n3768 = \P3_InstAddrPointer_reg[11]/NET0131  & \P3_InstAddrPointer_reg[12]/NET0131  ;
  assign n3769 = \P3_InstAddrPointer_reg[9]/NET0131  & n3768 ;
  assign n3770 = \P3_InstAddrPointer_reg[10]/NET0131  & n3769 ;
  assign n3771 = \P3_InstAddrPointer_reg[13]/NET0131  & n3770 ;
  assign n3772 = n3767 & n3771 ;
  assign n3773 = n3760 & n3772 ;
  assign n3775 = \P3_InstAddrPointer_reg[22]/NET0131  & n3773 ;
  assign n4090 = n3775 & n4089 ;
  assign n4148 = \P3_InstAddrPointer_reg[0]/NET0131  & n4090 ;
  assign n4149 = \P3_InstAddrPointer_reg[26]/NET0131  & n4148 ;
  assign n4150 = n4123 & n4149 ;
  assign n4091 = \P3_InstAddrPointer_reg[26]/NET0131  & n4090 ;
  assign n4117 = n4091 & n4116 ;
  assign n4151 = \P3_InstAddrPointer_reg[0]/NET0131  & n4117 ;
  assign n4152 = ~\P3_InstAddrPointer_reg[30]/NET0131  & ~n4151 ;
  assign n4153 = ~n4150 & ~n4152 ;
  assign n4154 = n4147 & ~n4153 ;
  assign n3727 = \P3_InstQueue_reg[14][7]/NET0131  & n2478 ;
  assign n3728 = \P3_InstQueue_reg[0][7]/NET0131  & n2484 ;
  assign n3741 = ~n3727 & ~n3728 ;
  assign n3729 = \P3_InstQueue_reg[5][7]/NET0131  & n2469 ;
  assign n3730 = \P3_InstQueue_reg[3][7]/NET0131  & n2466 ;
  assign n3742 = ~n3729 & ~n3730 ;
  assign n3749 = n3741 & n3742 ;
  assign n3723 = \P3_InstQueue_reg[8][7]/NET0131  & n2460 ;
  assign n3724 = \P3_InstQueue_reg[12][7]/NET0131  & n2486 ;
  assign n3739 = ~n3723 & ~n3724 ;
  assign n3725 = \P3_InstQueue_reg[2][7]/NET0131  & n2456 ;
  assign n3726 = \P3_InstQueue_reg[1][7]/NET0131  & n2482 ;
  assign n3740 = ~n3725 & ~n3726 ;
  assign n3750 = n3739 & n3740 ;
  assign n3751 = n3749 & n3750 ;
  assign n3735 = \P3_InstQueue_reg[7][7]/NET0131  & n2474 ;
  assign n3736 = \P3_InstQueue_reg[4][7]/NET0131  & n2480 ;
  assign n3745 = ~n3735 & ~n3736 ;
  assign n3737 = \P3_InstQueue_reg[13][7]/NET0131  & n2472 ;
  assign n3738 = \P3_InstQueue_reg[6][7]/NET0131  & n2492 ;
  assign n3746 = ~n3737 & ~n3738 ;
  assign n3747 = n3745 & n3746 ;
  assign n3731 = \P3_InstQueue_reg[9][7]/NET0131  & n2476 ;
  assign n3732 = \P3_InstQueue_reg[11][7]/NET0131  & n2464 ;
  assign n3743 = ~n3731 & ~n3732 ;
  assign n3733 = \P3_InstQueue_reg[10][7]/NET0131  & n2490 ;
  assign n3734 = \P3_InstQueue_reg[15][7]/NET0131  & n2488 ;
  assign n3744 = ~n3733 & ~n3734 ;
  assign n3748 = n3743 & n3744 ;
  assign n3752 = n3747 & n3748 ;
  assign n3753 = n3751 & n3752 ;
  assign n4159 = \P3_InstAddrPointer_reg[0]/NET0131  & n3763 ;
  assign n4160 = \P3_InstAddrPointer_reg[5]/NET0131  & n4159 ;
  assign n4161 = \P3_InstAddrPointer_reg[6]/NET0131  & n4160 ;
  assign n4162 = \P3_InstAddrPointer_reg[7]/NET0131  & n4161 ;
  assign n4177 = ~\P3_InstAddrPointer_reg[7]/NET0131  & ~n4161 ;
  assign n4178 = ~n4162 & ~n4177 ;
  assign n4179 = n3753 & ~n4178 ;
  assign n3870 = \P3_InstQueue_reg[8][2]/NET0131  & n2460 ;
  assign n3871 = \P3_InstQueue_reg[11][2]/NET0131  & n2464 ;
  assign n3884 = ~n3870 & ~n3871 ;
  assign n3872 = \P3_InstQueue_reg[10][2]/NET0131  & n2490 ;
  assign n3873 = \P3_InstQueue_reg[5][2]/NET0131  & n2469 ;
  assign n3885 = ~n3872 & ~n3873 ;
  assign n3892 = n3884 & n3885 ;
  assign n3866 = \P3_InstQueue_reg[14][2]/NET0131  & n2478 ;
  assign n3867 = \P3_InstQueue_reg[15][2]/NET0131  & n2488 ;
  assign n3882 = ~n3866 & ~n3867 ;
  assign n3868 = \P3_InstQueue_reg[3][2]/NET0131  & n2466 ;
  assign n3869 = \P3_InstQueue_reg[9][2]/NET0131  & n2476 ;
  assign n3883 = ~n3868 & ~n3869 ;
  assign n3893 = n3882 & n3883 ;
  assign n3894 = n3892 & n3893 ;
  assign n3878 = \P3_InstQueue_reg[7][2]/NET0131  & n2474 ;
  assign n3879 = \P3_InstQueue_reg[1][2]/NET0131  & n2482 ;
  assign n3888 = ~n3878 & ~n3879 ;
  assign n3880 = \P3_InstQueue_reg[6][2]/NET0131  & n2492 ;
  assign n3881 = \P3_InstQueue_reg[12][2]/NET0131  & n2486 ;
  assign n3889 = ~n3880 & ~n3881 ;
  assign n3890 = n3888 & n3889 ;
  assign n3874 = \P3_InstQueue_reg[4][2]/NET0131  & n2480 ;
  assign n3875 = \P3_InstQueue_reg[13][2]/NET0131  & n2472 ;
  assign n3886 = ~n3874 & ~n3875 ;
  assign n3876 = \P3_InstQueue_reg[2][2]/NET0131  & n2456 ;
  assign n3877 = \P3_InstQueue_reg[0][2]/NET0131  & n2484 ;
  assign n3887 = ~n3876 & ~n3877 ;
  assign n3891 = n3886 & n3887 ;
  assign n3895 = n3890 & n3891 ;
  assign n3896 = n3894 & n3895 ;
  assign n4186 = \P3_InstAddrPointer_reg[0]/NET0131  & \P3_InstAddrPointer_reg[1]/NET0131  ;
  assign n4187 = \P3_InstAddrPointer_reg[2]/NET0131  & n4186 ;
  assign n4188 = ~\P3_InstAddrPointer_reg[2]/NET0131  & ~n4186 ;
  assign n4189 = ~n4187 & ~n4188 ;
  assign n4190 = ~n3896 & n4189 ;
  assign n3904 = \P3_InstQueue_reg[10][1]/NET0131  & n2490 ;
  assign n3905 = \P3_InstQueue_reg[3][1]/NET0131  & n2466 ;
  assign n3918 = ~n3904 & ~n3905 ;
  assign n3906 = \P3_InstQueue_reg[8][1]/NET0131  & n2460 ;
  assign n3907 = \P3_InstQueue_reg[12][1]/NET0131  & n2486 ;
  assign n3919 = ~n3906 & ~n3907 ;
  assign n3926 = n3918 & n3919 ;
  assign n3900 = \P3_InstQueue_reg[6][1]/NET0131  & n2492 ;
  assign n3901 = \P3_InstQueue_reg[7][1]/NET0131  & n2474 ;
  assign n3916 = ~n3900 & ~n3901 ;
  assign n3902 = \P3_InstQueue_reg[9][1]/NET0131  & n2476 ;
  assign n3903 = \P3_InstQueue_reg[2][1]/NET0131  & n2456 ;
  assign n3917 = ~n3902 & ~n3903 ;
  assign n3927 = n3916 & n3917 ;
  assign n3928 = n3926 & n3927 ;
  assign n3912 = \P3_InstQueue_reg[0][1]/NET0131  & n2484 ;
  assign n3913 = \P3_InstQueue_reg[5][1]/NET0131  & n2469 ;
  assign n3922 = ~n3912 & ~n3913 ;
  assign n3914 = \P3_InstQueue_reg[11][1]/NET0131  & n2464 ;
  assign n3915 = \P3_InstQueue_reg[1][1]/NET0131  & n2482 ;
  assign n3923 = ~n3914 & ~n3915 ;
  assign n3924 = n3922 & n3923 ;
  assign n3908 = \P3_InstQueue_reg[13][1]/NET0131  & n2472 ;
  assign n3909 = \P3_InstQueue_reg[4][1]/NET0131  & n2480 ;
  assign n3920 = ~n3908 & ~n3909 ;
  assign n3910 = \P3_InstQueue_reg[14][1]/NET0131  & n2478 ;
  assign n3911 = \P3_InstQueue_reg[15][1]/NET0131  & n2488 ;
  assign n3921 = ~n3910 & ~n3911 ;
  assign n3925 = n3920 & n3921 ;
  assign n3929 = n3924 & n3925 ;
  assign n3930 = n3928 & n3929 ;
  assign n3931 = ~\P3_InstAddrPointer_reg[1]/NET0131  & ~n3930 ;
  assign n3932 = \P3_InstAddrPointer_reg[1]/NET0131  & n3930 ;
  assign n3937 = \P3_InstQueue_reg[7][0]/NET0131  & n2474 ;
  assign n3938 = \P3_InstQueue_reg[2][0]/NET0131  & n2456 ;
  assign n3951 = ~n3937 & ~n3938 ;
  assign n3939 = \P3_InstQueue_reg[1][0]/NET0131  & n2482 ;
  assign n3940 = \P3_InstQueue_reg[0][0]/NET0131  & n2484 ;
  assign n3952 = ~n3939 & ~n3940 ;
  assign n3959 = n3951 & n3952 ;
  assign n3933 = \P3_InstQueue_reg[8][0]/NET0131  & n2460 ;
  assign n3934 = \P3_InstQueue_reg[14][0]/NET0131  & n2478 ;
  assign n3949 = ~n3933 & ~n3934 ;
  assign n3935 = \P3_InstQueue_reg[3][0]/NET0131  & n2466 ;
  assign n3936 = \P3_InstQueue_reg[5][0]/NET0131  & n2469 ;
  assign n3950 = ~n3935 & ~n3936 ;
  assign n3960 = n3949 & n3950 ;
  assign n3961 = n3959 & n3960 ;
  assign n3945 = \P3_InstQueue_reg[13][0]/NET0131  & n2472 ;
  assign n3946 = \P3_InstQueue_reg[11][0]/NET0131  & n2464 ;
  assign n3955 = ~n3945 & ~n3946 ;
  assign n3947 = \P3_InstQueue_reg[6][0]/NET0131  & n2492 ;
  assign n3948 = \P3_InstQueue_reg[9][0]/NET0131  & n2476 ;
  assign n3956 = ~n3947 & ~n3948 ;
  assign n3957 = n3955 & n3956 ;
  assign n3941 = \P3_InstQueue_reg[12][0]/NET0131  & n2486 ;
  assign n3942 = \P3_InstQueue_reg[4][0]/NET0131  & n2480 ;
  assign n3953 = ~n3941 & ~n3942 ;
  assign n3943 = \P3_InstQueue_reg[10][0]/NET0131  & n2490 ;
  assign n3944 = \P3_InstQueue_reg[15][0]/NET0131  & n2488 ;
  assign n3954 = ~n3943 & ~n3944 ;
  assign n3958 = n3953 & n3954 ;
  assign n3962 = n3957 & n3958 ;
  assign n3963 = n3961 & n3962 ;
  assign n3964 = \P3_InstAddrPointer_reg[0]/NET0131  & ~n3963 ;
  assign n3965 = ~n3932 & n3964 ;
  assign n3966 = ~n3931 & ~n3965 ;
  assign n4191 = ~\P3_InstAddrPointer_reg[0]/NET0131  & \P3_InstAddrPointer_reg[1]/NET0131  ;
  assign n4192 = n3966 & ~n4191 ;
  assign n4193 = ~n4190 & n4192 ;
  assign n4194 = n3896 & ~n4189 ;
  assign n4006 = \P3_InstQueue_reg[11][3]/NET0131  & n2464 ;
  assign n4007 = \P3_InstQueue_reg[13][3]/NET0131  & n2472 ;
  assign n4020 = ~n4006 & ~n4007 ;
  assign n4008 = \P3_InstQueue_reg[1][3]/NET0131  & n2482 ;
  assign n4009 = \P3_InstQueue_reg[12][3]/NET0131  & n2486 ;
  assign n4021 = ~n4008 & ~n4009 ;
  assign n4028 = n4020 & n4021 ;
  assign n4002 = \P3_InstQueue_reg[5][3]/NET0131  & n2469 ;
  assign n4003 = \P3_InstQueue_reg[15][3]/NET0131  & n2488 ;
  assign n4018 = ~n4002 & ~n4003 ;
  assign n4004 = \P3_InstQueue_reg[10][3]/NET0131  & n2490 ;
  assign n4005 = \P3_InstQueue_reg[6][3]/NET0131  & n2492 ;
  assign n4019 = ~n4004 & ~n4005 ;
  assign n4029 = n4018 & n4019 ;
  assign n4030 = n4028 & n4029 ;
  assign n4014 = \P3_InstQueue_reg[8][3]/NET0131  & n2460 ;
  assign n4015 = \P3_InstQueue_reg[9][3]/NET0131  & n2476 ;
  assign n4024 = ~n4014 & ~n4015 ;
  assign n4016 = \P3_InstQueue_reg[14][3]/NET0131  & n2478 ;
  assign n4017 = \P3_InstQueue_reg[7][3]/NET0131  & n2474 ;
  assign n4025 = ~n4016 & ~n4017 ;
  assign n4026 = n4024 & n4025 ;
  assign n4010 = \P3_InstQueue_reg[4][3]/NET0131  & n2480 ;
  assign n4011 = \P3_InstQueue_reg[2][3]/NET0131  & n2456 ;
  assign n4022 = ~n4010 & ~n4011 ;
  assign n4012 = \P3_InstQueue_reg[0][3]/NET0131  & n2484 ;
  assign n4013 = \P3_InstQueue_reg[3][3]/NET0131  & n2466 ;
  assign n4023 = ~n4012 & ~n4013 ;
  assign n4027 = n4022 & n4023 ;
  assign n4031 = n4026 & n4027 ;
  assign n4032 = n4030 & n4031 ;
  assign n4195 = ~\P3_InstAddrPointer_reg[3]/NET0131  & ~n4187 ;
  assign n4196 = \P3_InstAddrPointer_reg[3]/NET0131  & n4187 ;
  assign n4197 = ~n4195 & ~n4196 ;
  assign n4198 = n4032 & ~n4197 ;
  assign n4199 = ~n4194 & ~n4198 ;
  assign n3974 = \P3_InstQueue_reg[6][4]/NET0131  & n2492 ;
  assign n3975 = \P3_InstQueue_reg[11][4]/NET0131  & n2464 ;
  assign n3988 = ~n3974 & ~n3975 ;
  assign n3976 = \P3_InstQueue_reg[9][4]/NET0131  & n2476 ;
  assign n3977 = \P3_InstQueue_reg[2][4]/NET0131  & n2456 ;
  assign n3989 = ~n3976 & ~n3977 ;
  assign n3996 = n3988 & n3989 ;
  assign n3970 = \P3_InstQueue_reg[10][4]/NET0131  & n2490 ;
  assign n3971 = \P3_InstQueue_reg[13][4]/NET0131  & n2472 ;
  assign n3986 = ~n3970 & ~n3971 ;
  assign n3972 = \P3_InstQueue_reg[15][4]/NET0131  & n2488 ;
  assign n3973 = \P3_InstQueue_reg[7][4]/NET0131  & n2474 ;
  assign n3987 = ~n3972 & ~n3973 ;
  assign n3997 = n3986 & n3987 ;
  assign n3998 = n3996 & n3997 ;
  assign n3982 = \P3_InstQueue_reg[5][4]/NET0131  & n2469 ;
  assign n3983 = \P3_InstQueue_reg[3][4]/NET0131  & n2466 ;
  assign n3992 = ~n3982 & ~n3983 ;
  assign n3984 = \P3_InstQueue_reg[8][4]/NET0131  & n2460 ;
  assign n3985 = \P3_InstQueue_reg[4][4]/NET0131  & n2480 ;
  assign n3993 = ~n3984 & ~n3985 ;
  assign n3994 = n3992 & n3993 ;
  assign n3978 = \P3_InstQueue_reg[0][4]/NET0131  & n2484 ;
  assign n3979 = \P3_InstQueue_reg[12][4]/NET0131  & n2486 ;
  assign n3990 = ~n3978 & ~n3979 ;
  assign n3980 = \P3_InstQueue_reg[1][4]/NET0131  & n2482 ;
  assign n3981 = \P3_InstQueue_reg[14][4]/NET0131  & n2478 ;
  assign n3991 = ~n3980 & ~n3981 ;
  assign n3995 = n3990 & n3991 ;
  assign n3999 = n3994 & n3995 ;
  assign n4000 = n3998 & n3999 ;
  assign n4200 = ~\P3_InstAddrPointer_reg[4]/NET0131  & ~n4196 ;
  assign n4201 = ~n4159 & ~n4200 ;
  assign n4202 = n4000 & ~n4201 ;
  assign n4203 = n4199 & ~n4202 ;
  assign n4204 = ~n4193 & n4203 ;
  assign n4205 = ~n4000 & n4201 ;
  assign n4206 = ~n4032 & n4197 ;
  assign n4207 = ~n4205 & ~n4206 ;
  assign n4208 = ~n4202 & ~n4207 ;
  assign n4209 = ~n4204 & ~n4208 ;
  assign n3838 = \P3_InstQueue_reg[4][6]/NET0131  & n2480 ;
  assign n3839 = \P3_InstQueue_reg[7][6]/NET0131  & n2474 ;
  assign n3852 = ~n3838 & ~n3839 ;
  assign n3840 = \P3_InstQueue_reg[11][6]/NET0131  & n2464 ;
  assign n3841 = \P3_InstQueue_reg[12][6]/NET0131  & n2486 ;
  assign n3853 = ~n3840 & ~n3841 ;
  assign n3860 = n3852 & n3853 ;
  assign n3834 = \P3_InstQueue_reg[2][6]/NET0131  & n2456 ;
  assign n3835 = \P3_InstQueue_reg[9][6]/NET0131  & n2476 ;
  assign n3850 = ~n3834 & ~n3835 ;
  assign n3836 = \P3_InstQueue_reg[15][6]/NET0131  & n2488 ;
  assign n3837 = \P3_InstQueue_reg[3][6]/NET0131  & n2466 ;
  assign n3851 = ~n3836 & ~n3837 ;
  assign n3861 = n3850 & n3851 ;
  assign n3862 = n3860 & n3861 ;
  assign n3846 = \P3_InstQueue_reg[5][6]/NET0131  & n2469 ;
  assign n3847 = \P3_InstQueue_reg[0][6]/NET0131  & n2484 ;
  assign n3856 = ~n3846 & ~n3847 ;
  assign n3848 = \P3_InstQueue_reg[10][6]/NET0131  & n2490 ;
  assign n3849 = \P3_InstQueue_reg[14][6]/NET0131  & n2478 ;
  assign n3857 = ~n3848 & ~n3849 ;
  assign n3858 = n3856 & n3857 ;
  assign n3842 = \P3_InstQueue_reg[1][6]/NET0131  & n2482 ;
  assign n3843 = \P3_InstQueue_reg[8][6]/NET0131  & n2460 ;
  assign n3854 = ~n3842 & ~n3843 ;
  assign n3844 = \P3_InstQueue_reg[13][6]/NET0131  & n2472 ;
  assign n3845 = \P3_InstQueue_reg[6][6]/NET0131  & n2492 ;
  assign n3855 = ~n3844 & ~n3845 ;
  assign n3859 = n3854 & n3855 ;
  assign n3863 = n3858 & n3859 ;
  assign n3864 = n3862 & n3863 ;
  assign n4180 = ~\P3_InstAddrPointer_reg[6]/NET0131  & ~n4160 ;
  assign n4181 = ~n4161 & ~n4180 ;
  assign n4182 = n3864 & ~n4181 ;
  assign n3804 = \P3_InstQueue_reg[4][5]/NET0131  & n2480 ;
  assign n3805 = \P3_InstQueue_reg[6][5]/NET0131  & n2492 ;
  assign n3818 = ~n3804 & ~n3805 ;
  assign n3806 = \P3_InstQueue_reg[11][5]/NET0131  & n2464 ;
  assign n3807 = \P3_InstQueue_reg[12][5]/NET0131  & n2486 ;
  assign n3819 = ~n3806 & ~n3807 ;
  assign n3826 = n3818 & n3819 ;
  assign n3800 = \P3_InstQueue_reg[2][5]/NET0131  & n2456 ;
  assign n3801 = \P3_InstQueue_reg[3][5]/NET0131  & n2466 ;
  assign n3816 = ~n3800 & ~n3801 ;
  assign n3802 = \P3_InstQueue_reg[15][5]/NET0131  & n2488 ;
  assign n3803 = \P3_InstQueue_reg[1][5]/NET0131  & n2482 ;
  assign n3817 = ~n3802 & ~n3803 ;
  assign n3827 = n3816 & n3817 ;
  assign n3828 = n3826 & n3827 ;
  assign n3812 = \P3_InstQueue_reg[5][5]/NET0131  & n2469 ;
  assign n3813 = \P3_InstQueue_reg[0][5]/NET0131  & n2484 ;
  assign n3822 = ~n3812 & ~n3813 ;
  assign n3814 = \P3_InstQueue_reg[13][5]/NET0131  & n2472 ;
  assign n3815 = \P3_InstQueue_reg[14][5]/NET0131  & n2478 ;
  assign n3823 = ~n3814 & ~n3815 ;
  assign n3824 = n3822 & n3823 ;
  assign n3808 = \P3_InstQueue_reg[10][5]/NET0131  & n2490 ;
  assign n3809 = \P3_InstQueue_reg[8][5]/NET0131  & n2460 ;
  assign n3820 = ~n3808 & ~n3809 ;
  assign n3810 = \P3_InstQueue_reg[9][5]/NET0131  & n2476 ;
  assign n3811 = \P3_InstQueue_reg[7][5]/NET0131  & n2474 ;
  assign n3821 = ~n3810 & ~n3811 ;
  assign n3825 = n3820 & n3821 ;
  assign n3829 = n3824 & n3825 ;
  assign n3830 = n3828 & n3829 ;
  assign n4183 = ~\P3_InstAddrPointer_reg[5]/NET0131  & ~n4159 ;
  assign n4184 = ~n4160 & ~n4183 ;
  assign n4185 = n3830 & ~n4184 ;
  assign n4210 = ~n4182 & ~n4185 ;
  assign n4211 = ~n4209 & n4210 ;
  assign n4212 = ~n4179 & n4211 ;
  assign n4221 = ~n4179 & ~n4182 ;
  assign n4222 = ~n3864 & n4181 ;
  assign n4223 = ~n3830 & n4184 ;
  assign n4224 = ~n4222 & ~n4223 ;
  assign n4225 = n4221 & ~n4224 ;
  assign n4218 = ~n3753 & n4178 ;
  assign n4163 = \P3_InstAddrPointer_reg[8]/NET0131  & n4162 ;
  assign n4219 = ~\P3_InstAddrPointer_reg[8]/NET0131  & ~n4162 ;
  assign n4220 = ~n4163 & ~n4219 ;
  assign n4226 = ~n4218 & ~n4220 ;
  assign n4227 = ~n4225 & n4226 ;
  assign n4067 = \P3_InstAddrPointer_reg[10]/NET0131  & n3778 ;
  assign n4155 = \P3_InstAddrPointer_reg[0]/NET0131  & n4067 ;
  assign n4213 = \P3_InstAddrPointer_reg[0]/NET0131  & n3778 ;
  assign n4214 = ~\P3_InstAddrPointer_reg[10]/NET0131  & ~n4213 ;
  assign n4215 = ~n4155 & ~n4214 ;
  assign n4216 = ~\P3_InstAddrPointer_reg[9]/NET0131  & ~n4163 ;
  assign n4217 = ~n4213 & ~n4216 ;
  assign n4228 = ~n4215 & ~n4217 ;
  assign n4229 = n4227 & n4228 ;
  assign n4230 = ~n4212 & n4229 ;
  assign n4156 = ~\P3_InstAddrPointer_reg[11]/NET0131  & ~n4155 ;
  assign n4157 = \P3_InstAddrPointer_reg[0]/NET0131  & n3780 ;
  assign n4158 = ~n4156 & ~n4157 ;
  assign n4164 = n3770 & n4163 ;
  assign n4165 = ~\P3_InstAddrPointer_reg[12]/NET0131  & ~n4157 ;
  assign n4166 = ~n4164 & ~n4165 ;
  assign n4167 = ~n4158 & ~n4166 ;
  assign n4168 = \P3_InstAddrPointer_reg[0]/NET0131  & n3772 ;
  assign n4169 = ~\P3_InstAddrPointer_reg[14]/NET0131  & ~n4168 ;
  assign n4064 = \P3_InstAddrPointer_reg[14]/NET0131  & n3772 ;
  assign n4170 = \P3_InstAddrPointer_reg[0]/NET0131  & n4064 ;
  assign n4171 = ~n4169 & ~n4170 ;
  assign n4057 = \P3_InstAddrPointer_reg[12]/NET0131  & n3780 ;
  assign n4173 = ~\P3_InstAddrPointer_reg[13]/NET0131  & ~n4057 ;
  assign n4172 = ~\P3_InstAddrPointer_reg[0]/NET0131  & ~\P3_InstAddrPointer_reg[13]/NET0131  ;
  assign n4174 = ~n4168 & ~n4172 ;
  assign n4175 = ~n4173 & n4174 ;
  assign n4176 = ~n4171 & ~n4175 ;
  assign n4231 = n4167 & n4176 ;
  assign n4232 = n4230 & n4231 ;
  assign n3782 = \P3_InstAddrPointer_reg[14]/NET0131  & n3781 ;
  assign n4233 = n3782 & n4157 ;
  assign n4234 = \P3_InstAddrPointer_reg[15]/NET0131  & n4233 ;
  assign n4235 = ~\P3_InstAddrPointer_reg[16]/NET0131  & ~n4234 ;
  assign n4236 = n3756 & n4233 ;
  assign n4237 = ~n4235 & ~n4236 ;
  assign n4238 = ~\P3_InstAddrPointer_reg[17]/NET0131  & ~n4236 ;
  assign n4239 = n3757 & n4170 ;
  assign n4240 = ~n4238 & ~n4239 ;
  assign n4241 = ~n4237 & ~n4240 ;
  assign n4242 = ~\P3_InstAddrPointer_reg[15]/NET0131  & ~n4233 ;
  assign n4243 = ~n4234 & ~n4242 ;
  assign n4244 = n4241 & ~n4243 ;
  assign n3783 = n3780 & n3782 ;
  assign n3784 = n3757 & n3783 ;
  assign n4245 = \P3_InstAddrPointer_reg[0]/NET0131  & n3784 ;
  assign n4246 = ~\P3_InstAddrPointer_reg[18]/NET0131  & ~n4245 ;
  assign n3794 = \P3_InstAddrPointer_reg[18]/NET0131  & n3784 ;
  assign n4247 = \P3_InstAddrPointer_reg[0]/NET0131  & n3794 ;
  assign n4248 = ~n4246 & ~n4247 ;
  assign n4249 = n4244 & ~n4248 ;
  assign n4250 = n4232 & n4249 ;
  assign n3785 = n3754 & n3784 ;
  assign n4251 = \P3_InstAddrPointer_reg[0]/NET0131  & n3785 ;
  assign n4252 = ~\P3_InstAddrPointer_reg[20]/NET0131  & ~n4251 ;
  assign n4253 = \P3_InstAddrPointer_reg[20]/NET0131  & n4251 ;
  assign n4254 = ~n4252 & ~n4253 ;
  assign n4255 = ~\P3_InstAddrPointer_reg[21]/NET0131  & ~n4253 ;
  assign n4256 = \P3_InstAddrPointer_reg[21]/NET0131  & n4253 ;
  assign n4257 = ~n4255 & ~n4256 ;
  assign n4258 = ~n4254 & ~n4257 ;
  assign n4102 = \P3_InstAddrPointer_reg[23]/NET0131  & n4096 ;
  assign n4259 = \P3_InstAddrPointer_reg[0]/NET0131  & n4102 ;
  assign n4260 = ~\P3_InstAddrPointer_reg[24]/NET0131  & ~n4259 ;
  assign n4261 = \P3_InstAddrPointer_reg[0]/NET0131  & n4096 ;
  assign n4262 = n4088 & n4261 ;
  assign n4263 = ~n4260 & ~n4262 ;
  assign n4264 = ~\P3_InstAddrPointer_reg[23]/NET0131  & ~n4261 ;
  assign n4265 = ~n4259 & ~n4264 ;
  assign n4266 = n4094 & n4168 ;
  assign n4267 = \P3_InstAddrPointer_reg[0]/NET0131  & n3773 ;
  assign n4268 = ~\P3_InstAddrPointer_reg[22]/NET0131  & ~n4267 ;
  assign n4269 = ~n4266 & ~n4268 ;
  assign n4270 = ~n4265 & ~n4269 ;
  assign n4271 = ~n4263 & n4270 ;
  assign n4272 = \P3_InstAddrPointer_reg[25]/NET0131  & ~n4262 ;
  assign n4273 = ~\P3_InstAddrPointer_reg[25]/NET0131  & n4262 ;
  assign n4274 = ~n4272 & ~n4273 ;
  assign n4275 = n4271 & n4274 ;
  assign n4276 = ~\P3_InstAddrPointer_reg[26]/NET0131  & ~n4148 ;
  assign n4277 = ~n4149 & ~n4276 ;
  assign n4278 = n4275 & ~n4277 ;
  assign n4279 = n4258 & n4278 ;
  assign n4280 = ~\P3_InstAddrPointer_reg[19]/NET0131  & ~n4247 ;
  assign n4281 = ~n4251 & ~n4280 ;
  assign n4282 = n4279 & ~n4281 ;
  assign n4283 = n4250 & n4282 ;
  assign n4284 = n4154 & n4283 ;
  assign n4286 = n4136 & n4284 ;
  assign n4285 = ~n4136 & ~n4284 ;
  assign n4287 = ~n3753 & ~n4285 ;
  assign n4288 = ~n4286 & n4287 ;
  assign n3897 = ~\P3_InstAddrPointer_reg[1]/NET0131  & ~\P3_InstAddrPointer_reg[2]/NET0131  ;
  assign n3898 = ~n3761 & ~n3897 ;
  assign n3899 = ~n3896 & n3898 ;
  assign n3967 = ~n3899 & n3966 ;
  assign n3968 = ~\P3_InstAddrPointer_reg[4]/NET0131  & ~n3762 ;
  assign n3969 = ~n3763 & ~n3968 ;
  assign n4001 = ~n3969 & n4000 ;
  assign n4033 = ~\P3_InstAddrPointer_reg[3]/NET0131  & ~n3761 ;
  assign n4034 = ~n3762 & ~n4033 ;
  assign n4035 = n4032 & ~n4034 ;
  assign n4036 = n3896 & ~n3898 ;
  assign n4037 = ~n4035 & ~n4036 ;
  assign n4038 = ~n4001 & n4037 ;
  assign n4039 = ~n3967 & n4038 ;
  assign n4040 = n3969 & ~n4000 ;
  assign n4041 = ~n4032 & n4034 ;
  assign n4042 = ~n4001 & n4041 ;
  assign n4043 = ~n4040 & ~n4042 ;
  assign n4044 = ~n4039 & n4043 ;
  assign n3798 = ~\P3_InstAddrPointer_reg[5]/NET0131  & ~n3763 ;
  assign n3799 = ~n3764 & ~n3798 ;
  assign n3831 = ~n3799 & n3830 ;
  assign n3832 = ~\P3_InstAddrPointer_reg[6]/NET0131  & ~n3764 ;
  assign n3833 = ~n3765 & ~n3832 ;
  assign n3865 = ~n3833 & n3864 ;
  assign n4045 = ~n3831 & ~n3865 ;
  assign n4046 = ~n4044 & n4045 ;
  assign n4047 = ~\P3_InstAddrPointer_reg[7]/NET0131  & ~n3765 ;
  assign n4048 = ~n3766 & ~n4047 ;
  assign n4049 = ~n3753 & n4048 ;
  assign n4050 = n3833 & ~n3864 ;
  assign n4051 = n3799 & ~n3830 ;
  assign n4052 = ~n3865 & n4051 ;
  assign n4053 = ~n4050 & ~n4052 ;
  assign n4054 = ~n4049 & n4053 ;
  assign n4055 = ~n4046 & n4054 ;
  assign n4056 = ~\P3_InstAddrPointer_reg[12]/NET0131  & ~n3780 ;
  assign n4058 = ~n4056 & ~n4057 ;
  assign n4059 = \P3_InstAddrPointer_reg[13]/NET0131  & n4058 ;
  assign n4060 = ~\P3_InstAddrPointer_reg[8]/NET0131  & ~n3766 ;
  assign n4061 = ~n3767 & ~n4060 ;
  assign n4062 = \P3_InstAddrPointer_reg[9]/NET0131  & n4061 ;
  assign n4063 = \P3_InstAddrPointer_reg[10]/NET0131  & n4062 ;
  assign n4070 = n3753 & ~n4048 ;
  assign n4071 = n4063 & ~n4070 ;
  assign n4065 = ~\P3_InstAddrPointer_reg[14]/NET0131  & ~n3772 ;
  assign n4066 = ~n4064 & ~n4065 ;
  assign n4068 = ~\P3_InstAddrPointer_reg[11]/NET0131  & ~n4067 ;
  assign n4069 = ~n3780 & ~n4068 ;
  assign n4072 = n4066 & n4069 ;
  assign n4073 = n4071 & n4072 ;
  assign n4074 = n4059 & n4073 ;
  assign n4075 = ~n4055 & n4074 ;
  assign n4076 = n3756 & n3783 ;
  assign n4077 = \P3_InstAddrPointer_reg[15]/NET0131  & n3783 ;
  assign n4078 = ~\P3_InstAddrPointer_reg[16]/NET0131  & ~n4077 ;
  assign n4079 = ~n4076 & ~n4078 ;
  assign n4080 = \P3_InstAddrPointer_reg[17]/NET0131  & n4079 ;
  assign n4081 = ~\P3_InstAddrPointer_reg[15]/NET0131  & ~n3783 ;
  assign n4082 = ~n4077 & ~n4081 ;
  assign n4083 = \P3_InstAddrPointer_reg[18]/NET0131  & n4082 ;
  assign n4084 = n4080 & n4083 ;
  assign n4085 = n4075 & n4084 ;
  assign n3774 = ~\P3_InstAddrPointer_reg[22]/NET0131  & ~n3773 ;
  assign n3776 = ~n3774 & ~n3775 ;
  assign n3786 = \P3_InstAddrPointer_reg[20]/NET0131  & n3785 ;
  assign n3787 = ~\P3_InstAddrPointer_reg[21]/NET0131  & ~n3786 ;
  assign n3788 = \P3_InstAddrPointer_reg[21]/NET0131  & n3786 ;
  assign n3789 = ~n3787 & ~n3788 ;
  assign n3790 = n3776 & n3789 ;
  assign n3791 = ~\P3_InstAddrPointer_reg[20]/NET0131  & ~n3785 ;
  assign n3792 = ~n3786 & ~n3791 ;
  assign n3793 = n3790 & n3792 ;
  assign n3795 = ~\P3_InstAddrPointer_reg[19]/NET0131  & n3794 ;
  assign n3796 = \P3_InstAddrPointer_reg[19]/NET0131  & ~n3794 ;
  assign n3797 = ~n3795 & ~n3796 ;
  assign n4086 = n3793 & ~n3797 ;
  assign n4087 = n4085 & n4086 ;
  assign n4092 = ~\P3_InstAddrPointer_reg[26]/NET0131  & ~n4090 ;
  assign n4093 = ~n4091 & ~n4092 ;
  assign n4097 = n4088 & n4096 ;
  assign n4098 = ~\P3_InstAddrPointer_reg[25]/NET0131  & ~n4097 ;
  assign n4099 = n4089 & n4096 ;
  assign n4100 = ~n4098 & ~n4099 ;
  assign n4101 = n4093 & n4100 ;
  assign n4103 = ~\P3_InstAddrPointer_reg[23]/NET0131  & ~n4096 ;
  assign n4104 = ~n4102 & ~n4103 ;
  assign n4105 = \P3_InstAddrPointer_reg[24]/NET0131  & n4104 ;
  assign n4106 = n4101 & n4105 ;
  assign n4107 = n4087 & n4106 ;
  assign n4110 = \P3_InstAddrPointer_reg[27]/NET0131  & n4109 ;
  assign n4111 = ~\P3_InstAddrPointer_reg[27]/NET0131  & ~n4109 ;
  assign n4112 = ~n4110 & ~n4111 ;
  assign n4113 = \P3_InstAddrPointer_reg[28]/NET0131  & n4112 ;
  assign n4114 = \P3_InstAddrPointer_reg[29]/NET0131  & n4113 ;
  assign n4118 = \P3_InstAddrPointer_reg[30]/NET0131  & ~n4117 ;
  assign n4119 = ~\P3_InstAddrPointer_reg[30]/NET0131  & n4117 ;
  assign n4120 = ~n4118 & ~n4119 ;
  assign n4121 = n4114 & ~n4120 ;
  assign n4122 = n4107 & n4121 ;
  assign n4125 = \P3_InstAddrPointer_reg[31]/NET0131  & ~n4124 ;
  assign n4127 = ~n4125 & ~n4126 ;
  assign n4129 = n4122 & n4127 ;
  assign n4128 = ~n4122 & ~n4127 ;
  assign n4130 = n3753 & ~n4128 ;
  assign n4131 = ~n4129 & n4130 ;
  assign n4289 = ~n2896 & ~n4131 ;
  assign n4290 = ~n4288 & n4289 ;
  assign n4291 = ~n3722 & ~n4290 ;
  assign n4292 = n2894 & ~n4291 ;
  assign n4293 = \P3_InstAddrPointer_reg[3]/NET0131  & ~n4188 ;
  assign n4294 = \P3_InstAddrPointer_reg[4]/NET0131  & n4293 ;
  assign n4295 = \P3_InstAddrPointer_reg[5]/NET0131  & n4294 ;
  assign n4296 = \P3_InstAddrPointer_reg[6]/NET0131  & n4295 ;
  assign n4297 = \P3_InstAddrPointer_reg[7]/NET0131  & n4296 ;
  assign n4298 = n3777 & n4297 ;
  assign n4299 = \P3_InstAddrPointer_reg[10]/NET0131  & n4298 ;
  assign n4300 = ~\P3_InstAddrPointer_reg[10]/NET0131  & ~n4298 ;
  assign n4301 = ~n4299 & ~n4300 ;
  assign n4302 = \P3_InstAddrPointer_reg[8]/NET0131  & n4297 ;
  assign n4303 = ~\P3_InstAddrPointer_reg[8]/NET0131  & ~n4297 ;
  assign n4304 = ~n4302 & ~n4303 ;
  assign n4305 = n3769 & n4304 ;
  assign n4306 = n4301 & n4305 ;
  assign n4307 = \P3_InstAddrPointer_reg[13]/NET0131  & n4306 ;
  assign n4308 = ~\P3_InstAddrPointer_reg[7]/NET0131  & ~n4296 ;
  assign n4309 = ~n4297 & ~n4308 ;
  assign n4310 = ~n3753 & n4309 ;
  assign n4311 = ~\P3_InstAddrPointer_reg[6]/NET0131  & ~n4295 ;
  assign n4312 = ~n4296 & ~n4311 ;
  assign n4313 = n3864 & ~n4312 ;
  assign n4314 = ~\P3_InstAddrPointer_reg[4]/NET0131  & ~n4293 ;
  assign n4315 = ~n4294 & ~n4314 ;
  assign n4316 = n4000 & ~n4315 ;
  assign n4317 = ~\P3_InstAddrPointer_reg[5]/NET0131  & ~n4294 ;
  assign n4318 = ~n4295 & ~n4317 ;
  assign n4319 = n3830 & ~n4318 ;
  assign n4320 = ~n4316 & ~n4319 ;
  assign n4321 = ~n3896 & ~n4189 ;
  assign n4322 = \P3_InstAddrPointer_reg[0]/NET0131  & ~\P3_InstAddrPointer_reg[1]/NET0131  ;
  assign n4323 = ~n4191 & ~n4322 ;
  assign n4324 = ~n3930 & ~n4323 ;
  assign n4325 = n3930 & n4323 ;
  assign n4326 = ~\P3_InstAddrPointer_reg[0]/NET0131  & ~n3963 ;
  assign n4327 = ~n4325 & n4326 ;
  assign n4328 = ~n4324 & ~n4327 ;
  assign n4329 = ~n4321 & n4328 ;
  assign n4330 = n3896 & n4189 ;
  assign n4331 = ~\P3_InstAddrPointer_reg[3]/NET0131  & n4188 ;
  assign n4332 = ~n4293 & ~n4331 ;
  assign n4333 = n4032 & ~n4332 ;
  assign n4334 = ~n4330 & ~n4333 ;
  assign n4335 = ~n4329 & n4334 ;
  assign n4336 = ~n4032 & n4332 ;
  assign n4337 = ~n4000 & n4315 ;
  assign n4338 = ~n4336 & ~n4337 ;
  assign n4339 = ~n4335 & n4338 ;
  assign n4340 = n4320 & ~n4339 ;
  assign n4341 = ~n3864 & n4312 ;
  assign n4342 = ~n3830 & n4318 ;
  assign n4343 = ~n4341 & ~n4342 ;
  assign n4344 = ~n4340 & n4343 ;
  assign n4345 = ~n4313 & ~n4344 ;
  assign n4346 = n3753 & ~n4309 ;
  assign n4347 = n4345 & ~n4346 ;
  assign n4348 = ~n4310 & ~n4347 ;
  assign n4349 = n4307 & ~n4348 ;
  assign n4350 = n3768 & n4299 ;
  assign n4351 = \P3_InstAddrPointer_reg[13]/NET0131  & n4350 ;
  assign n4352 = ~\P3_InstAddrPointer_reg[14]/NET0131  & ~n4351 ;
  assign n4353 = \P3_InstAddrPointer_reg[14]/NET0131  & n4351 ;
  assign n4354 = ~n4352 & ~n4353 ;
  assign n4355 = n3756 & n4354 ;
  assign n4356 = n4349 & n4355 ;
  assign n4357 = n3756 & n4353 ;
  assign n4358 = ~\P3_InstAddrPointer_reg[17]/NET0131  & ~n4357 ;
  assign n4359 = \P3_InstAddrPointer_reg[17]/NET0131  & n4357 ;
  assign n4360 = ~n4358 & ~n4359 ;
  assign n4361 = n3755 & n4360 ;
  assign n4362 = n4356 & n4361 ;
  assign n4363 = \P3_InstAddrPointer_reg[18]/NET0131  & n4359 ;
  assign n4364 = \P3_InstAddrPointer_reg[19]/NET0131  & n4363 ;
  assign n4365 = \P3_InstAddrPointer_reg[20]/NET0131  & n4364 ;
  assign n4366 = ~\P3_InstAddrPointer_reg[21]/NET0131  & ~n4365 ;
  assign n4367 = n3760 & n4351 ;
  assign n4368 = ~n4366 & ~n4367 ;
  assign n4369 = ~\P3_InstAddrPointer_reg[22]/NET0131  & ~n4367 ;
  assign n4370 = n4094 & n4351 ;
  assign n4371 = ~n4369 & ~n4370 ;
  assign n4372 = n4088 & n4371 ;
  assign n4373 = n4368 & n4372 ;
  assign n4374 = n4362 & n4373 ;
  assign n4375 = \P3_InstAddrPointer_reg[23]/NET0131  & n4370 ;
  assign n4376 = \P3_InstAddrPointer_reg[24]/NET0131  & n4375 ;
  assign n4377 = ~\P3_InstAddrPointer_reg[25]/NET0131  & ~n4376 ;
  assign n4378 = \P3_InstAddrPointer_reg[25]/NET0131  & n4376 ;
  assign n4379 = ~n4377 & ~n4378 ;
  assign n4380 = \P3_InstAddrPointer_reg[26]/NET0131  & n4379 ;
  assign n4381 = \P3_InstAddrPointer_reg[26]/NET0131  & n4378 ;
  assign n4382 = n4116 & n4381 ;
  assign n4383 = ~\P3_InstAddrPointer_reg[30]/NET0131  & ~n4382 ;
  assign n4384 = n4123 & n4381 ;
  assign n4385 = ~n4383 & ~n4384 ;
  assign n4386 = \P3_InstAddrPointer_reg[27]/NET0131  & n4381 ;
  assign n4387 = ~\P3_InstAddrPointer_reg[27]/NET0131  & ~n4381 ;
  assign n4388 = ~n4386 & ~n4387 ;
  assign n4389 = \P3_InstAddrPointer_reg[28]/NET0131  & n4388 ;
  assign n4390 = \P3_InstAddrPointer_reg[29]/NET0131  & n4389 ;
  assign n4391 = n4385 & n4390 ;
  assign n4392 = n4380 & n4391 ;
  assign n4393 = n4374 & n4392 ;
  assign n4394 = ~\P3_InstAddrPointer_reg[31]/NET0131  & ~n4384 ;
  assign n4395 = \P3_InstAddrPointer_reg[31]/NET0131  & n4384 ;
  assign n4396 = ~n4394 & ~n4395 ;
  assign n4398 = ~n4393 & ~n4396 ;
  assign n4397 = n4393 & n4396 ;
  assign n4399 = n2905 & ~n4397 ;
  assign n4400 = ~n4398 & n4399 ;
  assign n4405 = n2918 & n4396 ;
  assign n4404 = ~n2923 & ~n4127 ;
  assign n4401 = ~n2777 & ~n4136 ;
  assign n4402 = ~n2900 & n2925 ;
  assign n4403 = \P3_InstAddrPointer_reg[31]/NET0131  & ~n4402 ;
  assign n4406 = ~n4401 & ~n4403 ;
  assign n4407 = ~n4404 & n4406 ;
  assign n4408 = ~n4405 & n4407 ;
  assign n4409 = ~n4400 & n4408 ;
  assign n4410 = ~n4292 & n4409 ;
  assign n4411 = n2453 & ~n4410 ;
  assign n4412 = n2951 & n2961 ;
  assign n4413 = \P3_rEIP_reg[31]/NET0131  & n4412 ;
  assign n4414 = ~n2951 & n2961 ;
  assign n4415 = n2452 & n2951 ;
  assign n4416 = ~n2958 & ~n4415 ;
  assign n4417 = ~n2996 & n4416 ;
  assign n4418 = ~n4414 & n4417 ;
  assign n4419 = \P3_InstAddrPointer_reg[31]/NET0131  & ~n4418 ;
  assign n4420 = ~n4413 & ~n4419 ;
  assign n4421 = ~n4411 & n4420 ;
  assign n4422 = \P1_InstAddrPointer_reg[30]/NET0131  & n2375 ;
  assign n4454 = \P1_InstAddrPointer_reg[12]/NET0131  & \P1_InstAddrPointer_reg[13]/NET0131  ;
  assign n4455 = \P1_InstAddrPointer_reg[1]/NET0131  & \P1_InstAddrPointer_reg[2]/NET0131  ;
  assign n4456 = \P1_InstAddrPointer_reg[3]/NET0131  & n4455 ;
  assign n4457 = \P1_InstAddrPointer_reg[4]/NET0131  & n4456 ;
  assign n4458 = \P1_InstAddrPointer_reg[5]/NET0131  & n4457 ;
  assign n4459 = \P1_InstAddrPointer_reg[6]/NET0131  & n4458 ;
  assign n4461 = \P1_InstAddrPointer_reg[7]/NET0131  & \P1_InstAddrPointer_reg[8]/NET0131  ;
  assign n4460 = \P1_InstAddrPointer_reg[10]/NET0131  & \P1_InstAddrPointer_reg[9]/NET0131  ;
  assign n4462 = \P1_InstAddrPointer_reg[11]/NET0131  & n4460 ;
  assign n4463 = n4461 & n4462 ;
  assign n4464 = n4459 & n4463 ;
  assign n4465 = n4454 & n4464 ;
  assign n4466 = \P1_InstAddrPointer_reg[14]/NET0131  & \P1_InstAddrPointer_reg[15]/NET0131  ;
  assign n4467 = \P1_InstAddrPointer_reg[16]/NET0131  & n4466 ;
  assign n4468 = n4465 & n4467 ;
  assign n4469 = \P1_InstAddrPointer_reg[17]/NET0131  & \P1_InstAddrPointer_reg[18]/NET0131  ;
  assign n4470 = \P1_InstAddrPointer_reg[19]/NET0131  & n4469 ;
  assign n4471 = n4468 & n4470 ;
  assign n4472 = \P1_InstAddrPointer_reg[20]/NET0131  & \P1_InstAddrPointer_reg[21]/NET0131  ;
  assign n4477 = \P1_InstAddrPointer_reg[22]/NET0131  & \P1_InstAddrPointer_reg[23]/NET0131  ;
  assign n4478 = n4472 & n4477 ;
  assign n4479 = n4471 & n4478 ;
  assign n4483 = \P1_InstAddrPointer_reg[24]/NET0131  & n4479 ;
  assign n4484 = \P1_InstAddrPointer_reg[25]/NET0131  & n4483 ;
  assign n4489 = \P1_InstAddrPointer_reg[26]/NET0131  & n4484 ;
  assign n4490 = \P1_InstAddrPointer_reg[27]/NET0131  & n4489 ;
  assign n4807 = \P1_InstAddrPointer_reg[0]/NET0131  & n4490 ;
  assign n4808 = \P1_InstAddrPointer_reg[28]/NET0131  & n4807 ;
  assign n4809 = \P1_InstAddrPointer_reg[29]/NET0131  & n4808 ;
  assign n4810 = ~\P1_InstAddrPointer_reg[30]/NET0131  & ~n4809 ;
  assign n4811 = \P1_InstAddrPointer_reg[30]/NET0131  & n4809 ;
  assign n4812 = ~n4810 & ~n4811 ;
  assign n4813 = \P1_InstAddrPointer_reg[0]/NET0131  & \P1_InstAddrPointer_reg[1]/NET0131  ;
  assign n4814 = \P1_InstAddrPointer_reg[2]/NET0131  & n4813 ;
  assign n4815 = \P1_InstAddrPointer_reg[3]/NET0131  & n4814 ;
  assign n4816 = \P1_InstAddrPointer_reg[4]/NET0131  & n4815 ;
  assign n4817 = \P1_InstAddrPointer_reg[5]/NET0131  & n4816 ;
  assign n4818 = \P1_InstAddrPointer_reg[6]/NET0131  & n4817 ;
  assign n4819 = \P1_InstAddrPointer_reg[7]/NET0131  & n4818 ;
  assign n4820 = \P1_InstAddrPointer_reg[8]/NET0131  & n4819 ;
  assign n4821 = \P1_InstAddrPointer_reg[9]/NET0131  & n4820 ;
  assign n4822 = ~\P1_InstAddrPointer_reg[10]/NET0131  & ~n4821 ;
  assign n4496 = n4459 & n4461 ;
  assign n4497 = \P1_InstAddrPointer_reg[9]/NET0131  & n4496 ;
  assign n4771 = \P1_InstAddrPointer_reg[10]/NET0131  & n4497 ;
  assign n4823 = \P1_InstAddrPointer_reg[0]/NET0131  & n4771 ;
  assign n4824 = ~n4822 & ~n4823 ;
  assign n4427 = \P1_InstQueue_reg[7][7]/NET0131  & n1972 ;
  assign n4428 = \P1_InstQueue_reg[11][7]/NET0131  & n1946 ;
  assign n4441 = ~n4427 & ~n4428 ;
  assign n4429 = \P1_InstQueue_reg[10][7]/NET0131  & n1978 ;
  assign n4430 = \P1_InstQueue_reg[14][7]/NET0131  & n1980 ;
  assign n4442 = ~n4429 & ~n4430 ;
  assign n4449 = n4441 & n4442 ;
  assign n4423 = \P1_InstQueue_reg[8][7]/NET0131  & n1968 ;
  assign n4424 = \P1_InstQueue_reg[1][7]/NET0131  & n1958 ;
  assign n4439 = ~n4423 & ~n4424 ;
  assign n4425 = \P1_InstQueue_reg[12][7]/NET0131  & n1949 ;
  assign n4426 = \P1_InstQueue_reg[13][7]/NET0131  & n1953 ;
  assign n4440 = ~n4425 & ~n4426 ;
  assign n4450 = n4439 & n4440 ;
  assign n4451 = n4449 & n4450 ;
  assign n4435 = \P1_InstQueue_reg[2][7]/NET0131  & n1966 ;
  assign n4436 = \P1_InstQueue_reg[0][7]/NET0131  & n1982 ;
  assign n4445 = ~n4435 & ~n4436 ;
  assign n4437 = \P1_InstQueue_reg[3][7]/NET0131  & n1970 ;
  assign n4438 = \P1_InstQueue_reg[4][7]/NET0131  & n1976 ;
  assign n4446 = ~n4437 & ~n4438 ;
  assign n4447 = n4445 & n4446 ;
  assign n4431 = \P1_InstQueue_reg[9][7]/NET0131  & n1974 ;
  assign n4432 = \P1_InstQueue_reg[6][7]/NET0131  & n1964 ;
  assign n4443 = ~n4431 & ~n4432 ;
  assign n4433 = \P1_InstQueue_reg[5][7]/NET0131  & n1961 ;
  assign n4434 = \P1_InstQueue_reg[15][7]/NET0131  & n1955 ;
  assign n4444 = ~n4433 & ~n4434 ;
  assign n4448 = n4443 & n4444 ;
  assign n4452 = n4447 & n4448 ;
  assign n4453 = n4451 & n4452 ;
  assign n4825 = ~\P1_InstAddrPointer_reg[7]/NET0131  & ~n4818 ;
  assign n4826 = ~n4819 & ~n4825 ;
  assign n4827 = n4453 & ~n4826 ;
  assign n4547 = \P1_InstQueue_reg[4][5]/NET0131  & n1976 ;
  assign n4548 = \P1_InstQueue_reg[13][5]/NET0131  & n1953 ;
  assign n4561 = ~n4547 & ~n4548 ;
  assign n4549 = \P1_InstQueue_reg[12][5]/NET0131  & n1949 ;
  assign n4550 = \P1_InstQueue_reg[9][5]/NET0131  & n1974 ;
  assign n4562 = ~n4549 & ~n4550 ;
  assign n4569 = n4561 & n4562 ;
  assign n4543 = \P1_InstQueue_reg[1][5]/NET0131  & n1958 ;
  assign n4544 = \P1_InstQueue_reg[14][5]/NET0131  & n1980 ;
  assign n4559 = ~n4543 & ~n4544 ;
  assign n4545 = \P1_InstQueue_reg[3][5]/NET0131  & n1970 ;
  assign n4546 = \P1_InstQueue_reg[10][5]/NET0131  & n1978 ;
  assign n4560 = ~n4545 & ~n4546 ;
  assign n4570 = n4559 & n4560 ;
  assign n4571 = n4569 & n4570 ;
  assign n4555 = \P1_InstQueue_reg[15][5]/NET0131  & n1955 ;
  assign n4556 = \P1_InstQueue_reg[6][5]/NET0131  & n1964 ;
  assign n4565 = ~n4555 & ~n4556 ;
  assign n4557 = \P1_InstQueue_reg[5][5]/NET0131  & n1961 ;
  assign n4558 = \P1_InstQueue_reg[7][5]/NET0131  & n1972 ;
  assign n4566 = ~n4557 & ~n4558 ;
  assign n4567 = n4565 & n4566 ;
  assign n4551 = \P1_InstQueue_reg[0][5]/NET0131  & n1982 ;
  assign n4552 = \P1_InstQueue_reg[8][5]/NET0131  & n1968 ;
  assign n4563 = ~n4551 & ~n4552 ;
  assign n4553 = \P1_InstQueue_reg[2][5]/NET0131  & n1966 ;
  assign n4554 = \P1_InstQueue_reg[11][5]/NET0131  & n1946 ;
  assign n4564 = ~n4553 & ~n4554 ;
  assign n4568 = n4563 & n4564 ;
  assign n4572 = n4567 & n4568 ;
  assign n4573 = n4571 & n4572 ;
  assign n4828 = ~\P1_InstAddrPointer_reg[5]/NET0131  & ~n4816 ;
  assign n4829 = ~n4817 & ~n4828 ;
  assign n4830 = n4573 & ~n4829 ;
  assign n4513 = \P1_InstQueue_reg[15][6]/NET0131  & n1955 ;
  assign n4514 = \P1_InstQueue_reg[14][6]/NET0131  & n1980 ;
  assign n4527 = ~n4513 & ~n4514 ;
  assign n4515 = \P1_InstQueue_reg[8][6]/NET0131  & n1968 ;
  assign n4516 = \P1_InstQueue_reg[1][6]/NET0131  & n1958 ;
  assign n4528 = ~n4515 & ~n4516 ;
  assign n4535 = n4527 & n4528 ;
  assign n4509 = \P1_InstQueue_reg[3][6]/NET0131  & n1970 ;
  assign n4510 = \P1_InstQueue_reg[2][6]/NET0131  & n1966 ;
  assign n4525 = ~n4509 & ~n4510 ;
  assign n4511 = \P1_InstQueue_reg[7][6]/NET0131  & n1972 ;
  assign n4512 = \P1_InstQueue_reg[5][6]/NET0131  & n1961 ;
  assign n4526 = ~n4511 & ~n4512 ;
  assign n4536 = n4525 & n4526 ;
  assign n4537 = n4535 & n4536 ;
  assign n4521 = \P1_InstQueue_reg[6][6]/NET0131  & n1964 ;
  assign n4522 = \P1_InstQueue_reg[9][6]/NET0131  & n1974 ;
  assign n4531 = ~n4521 & ~n4522 ;
  assign n4523 = \P1_InstQueue_reg[4][6]/NET0131  & n1976 ;
  assign n4524 = \P1_InstQueue_reg[0][6]/NET0131  & n1982 ;
  assign n4532 = ~n4523 & ~n4524 ;
  assign n4533 = n4531 & n4532 ;
  assign n4517 = \P1_InstQueue_reg[12][6]/NET0131  & n1949 ;
  assign n4518 = \P1_InstQueue_reg[11][6]/NET0131  & n1946 ;
  assign n4529 = ~n4517 & ~n4518 ;
  assign n4519 = \P1_InstQueue_reg[10][6]/NET0131  & n1978 ;
  assign n4520 = \P1_InstQueue_reg[13][6]/NET0131  & n1953 ;
  assign n4530 = ~n4519 & ~n4520 ;
  assign n4534 = n4529 & n4530 ;
  assign n4538 = n4533 & n4534 ;
  assign n4539 = n4537 & n4538 ;
  assign n4831 = ~\P1_InstAddrPointer_reg[6]/NET0131  & ~n4817 ;
  assign n4832 = ~n4818 & ~n4831 ;
  assign n4833 = n4539 & ~n4832 ;
  assign n4834 = ~n4830 & ~n4833 ;
  assign n4835 = ~n4827 & n4834 ;
  assign n4581 = \P1_InstQueue_reg[2][4]/NET0131  & n1966 ;
  assign n4582 = \P1_InstQueue_reg[11][4]/NET0131  & n1946 ;
  assign n4595 = ~n4581 & ~n4582 ;
  assign n4583 = \P1_InstQueue_reg[14][4]/NET0131  & n1980 ;
  assign n4584 = \P1_InstQueue_reg[9][4]/NET0131  & n1974 ;
  assign n4596 = ~n4583 & ~n4584 ;
  assign n4603 = n4595 & n4596 ;
  assign n4577 = \P1_InstQueue_reg[0][4]/NET0131  & n1982 ;
  assign n4578 = \P1_InstQueue_reg[13][4]/NET0131  & n1953 ;
  assign n4593 = ~n4577 & ~n4578 ;
  assign n4579 = \P1_InstQueue_reg[10][4]/NET0131  & n1978 ;
  assign n4580 = \P1_InstQueue_reg[1][4]/NET0131  & n1958 ;
  assign n4594 = ~n4579 & ~n4580 ;
  assign n4604 = n4593 & n4594 ;
  assign n4605 = n4603 & n4604 ;
  assign n4589 = \P1_InstQueue_reg[4][4]/NET0131  & n1976 ;
  assign n4590 = \P1_InstQueue_reg[8][4]/NET0131  & n1968 ;
  assign n4599 = ~n4589 & ~n4590 ;
  assign n4591 = \P1_InstQueue_reg[3][4]/NET0131  & n1970 ;
  assign n4592 = \P1_InstQueue_reg[7][4]/NET0131  & n1972 ;
  assign n4600 = ~n4591 & ~n4592 ;
  assign n4601 = n4599 & n4600 ;
  assign n4585 = \P1_InstQueue_reg[12][4]/NET0131  & n1949 ;
  assign n4586 = \P1_InstQueue_reg[6][4]/NET0131  & n1964 ;
  assign n4597 = ~n4585 & ~n4586 ;
  assign n4587 = \P1_InstQueue_reg[5][4]/NET0131  & n1961 ;
  assign n4588 = \P1_InstQueue_reg[15][4]/NET0131  & n1955 ;
  assign n4598 = ~n4587 & ~n4588 ;
  assign n4602 = n4597 & n4598 ;
  assign n4606 = n4601 & n4602 ;
  assign n4607 = n4605 & n4606 ;
  assign n4836 = ~\P1_InstAddrPointer_reg[4]/NET0131  & ~n4815 ;
  assign n4837 = ~n4816 & ~n4836 ;
  assign n4838 = n4607 & ~n4837 ;
  assign n4684 = \P1_InstQueue_reg[12][1]/NET0131  & n1949 ;
  assign n4685 = \P1_InstQueue_reg[1][1]/NET0131  & n1958 ;
  assign n4698 = ~n4684 & ~n4685 ;
  assign n4686 = \P1_InstQueue_reg[5][1]/NET0131  & n1961 ;
  assign n4687 = \P1_InstQueue_reg[3][1]/NET0131  & n1970 ;
  assign n4699 = ~n4686 & ~n4687 ;
  assign n4706 = n4698 & n4699 ;
  assign n4680 = \P1_InstQueue_reg[14][1]/NET0131  & n1980 ;
  assign n4681 = \P1_InstQueue_reg[6][1]/NET0131  & n1964 ;
  assign n4696 = ~n4680 & ~n4681 ;
  assign n4682 = \P1_InstQueue_reg[4][1]/NET0131  & n1976 ;
  assign n4683 = \P1_InstQueue_reg[8][1]/NET0131  & n1968 ;
  assign n4697 = ~n4682 & ~n4683 ;
  assign n4707 = n4696 & n4697 ;
  assign n4708 = n4706 & n4707 ;
  assign n4692 = \P1_InstQueue_reg[10][1]/NET0131  & n1978 ;
  assign n4693 = \P1_InstQueue_reg[11][1]/NET0131  & n1946 ;
  assign n4702 = ~n4692 & ~n4693 ;
  assign n4694 = \P1_InstQueue_reg[9][1]/NET0131  & n1974 ;
  assign n4695 = \P1_InstQueue_reg[2][1]/NET0131  & n1966 ;
  assign n4703 = ~n4694 & ~n4695 ;
  assign n4704 = n4702 & n4703 ;
  assign n4688 = \P1_InstQueue_reg[13][1]/NET0131  & n1953 ;
  assign n4689 = \P1_InstQueue_reg[0][1]/NET0131  & n1982 ;
  assign n4700 = ~n4688 & ~n4689 ;
  assign n4690 = \P1_InstQueue_reg[7][1]/NET0131  & n1972 ;
  assign n4691 = \P1_InstQueue_reg[15][1]/NET0131  & n1955 ;
  assign n4701 = ~n4690 & ~n4691 ;
  assign n4705 = n4700 & n4701 ;
  assign n4709 = n4704 & n4705 ;
  assign n4710 = n4708 & n4709 ;
  assign n4839 = ~\P1_InstAddrPointer_reg[0]/NET0131  & ~\P1_InstAddrPointer_reg[1]/NET0131  ;
  assign n4840 = ~n4813 & ~n4839 ;
  assign n4841 = n4710 & ~n4840 ;
  assign n4711 = ~\P1_InstAddrPointer_reg[1]/NET0131  & ~n4710 ;
  assign n4717 = \P1_InstQueue_reg[8][0]/NET0131  & n1968 ;
  assign n4718 = \P1_InstQueue_reg[7][0]/NET0131  & n1972 ;
  assign n4731 = ~n4717 & ~n4718 ;
  assign n4719 = \P1_InstQueue_reg[12][0]/NET0131  & n1949 ;
  assign n4720 = \P1_InstQueue_reg[9][0]/NET0131  & n1974 ;
  assign n4732 = ~n4719 & ~n4720 ;
  assign n4739 = n4731 & n4732 ;
  assign n4713 = \P1_InstQueue_reg[13][0]/NET0131  & n1953 ;
  assign n4714 = \P1_InstQueue_reg[1][0]/NET0131  & n1958 ;
  assign n4729 = ~n4713 & ~n4714 ;
  assign n4715 = \P1_InstQueue_reg[14][0]/NET0131  & n1980 ;
  assign n4716 = \P1_InstQueue_reg[3][0]/NET0131  & n1970 ;
  assign n4730 = ~n4715 & ~n4716 ;
  assign n4740 = n4729 & n4730 ;
  assign n4741 = n4739 & n4740 ;
  assign n4725 = \P1_InstQueue_reg[11][0]/NET0131  & n1946 ;
  assign n4726 = \P1_InstQueue_reg[2][0]/NET0131  & n1966 ;
  assign n4735 = ~n4725 & ~n4726 ;
  assign n4727 = \P1_InstQueue_reg[6][0]/NET0131  & n1964 ;
  assign n4728 = \P1_InstQueue_reg[10][0]/NET0131  & n1978 ;
  assign n4736 = ~n4727 & ~n4728 ;
  assign n4737 = n4735 & n4736 ;
  assign n4721 = \P1_InstQueue_reg[5][0]/NET0131  & n1961 ;
  assign n4722 = \P1_InstQueue_reg[0][0]/NET0131  & n1982 ;
  assign n4733 = ~n4721 & ~n4722 ;
  assign n4723 = \P1_InstQueue_reg[4][0]/NET0131  & n1976 ;
  assign n4724 = \P1_InstQueue_reg[15][0]/NET0131  & n1955 ;
  assign n4734 = ~n4723 & ~n4724 ;
  assign n4738 = n4733 & n4734 ;
  assign n4742 = n4737 & n4738 ;
  assign n4743 = n4741 & n4742 ;
  assign n4842 = \P1_InstAddrPointer_reg[0]/NET0131  & n4743 ;
  assign n4843 = ~n4711 & n4842 ;
  assign n4844 = ~n4841 & ~n4843 ;
  assign n4613 = \P1_InstQueue_reg[2][3]/NET0131  & n1966 ;
  assign n4614 = \P1_InstQueue_reg[6][3]/NET0131  & n1964 ;
  assign n4627 = ~n4613 & ~n4614 ;
  assign n4615 = \P1_InstQueue_reg[9][3]/NET0131  & n1974 ;
  assign n4616 = \P1_InstQueue_reg[8][3]/NET0131  & n1968 ;
  assign n4628 = ~n4615 & ~n4616 ;
  assign n4635 = n4627 & n4628 ;
  assign n4609 = \P1_InstQueue_reg[7][3]/NET0131  & n1972 ;
  assign n4610 = \P1_InstQueue_reg[0][3]/NET0131  & n1982 ;
  assign n4625 = ~n4609 & ~n4610 ;
  assign n4611 = \P1_InstQueue_reg[14][3]/NET0131  & n1980 ;
  assign n4612 = \P1_InstQueue_reg[12][3]/NET0131  & n1949 ;
  assign n4626 = ~n4611 & ~n4612 ;
  assign n4636 = n4625 & n4626 ;
  assign n4637 = n4635 & n4636 ;
  assign n4621 = \P1_InstQueue_reg[5][3]/NET0131  & n1961 ;
  assign n4622 = \P1_InstQueue_reg[13][3]/NET0131  & n1953 ;
  assign n4631 = ~n4621 & ~n4622 ;
  assign n4623 = \P1_InstQueue_reg[3][3]/NET0131  & n1970 ;
  assign n4624 = \P1_InstQueue_reg[11][3]/NET0131  & n1946 ;
  assign n4632 = ~n4623 & ~n4624 ;
  assign n4633 = n4631 & n4632 ;
  assign n4617 = \P1_InstQueue_reg[15][3]/NET0131  & n1955 ;
  assign n4618 = \P1_InstQueue_reg[10][3]/NET0131  & n1978 ;
  assign n4629 = ~n4617 & ~n4618 ;
  assign n4619 = \P1_InstQueue_reg[1][3]/NET0131  & n1958 ;
  assign n4620 = \P1_InstQueue_reg[4][3]/NET0131  & n1976 ;
  assign n4630 = ~n4619 & ~n4620 ;
  assign n4634 = n4629 & n4630 ;
  assign n4638 = n4633 & n4634 ;
  assign n4639 = n4637 & n4638 ;
  assign n4845 = ~\P1_InstAddrPointer_reg[3]/NET0131  & ~n4814 ;
  assign n4846 = ~n4815 & ~n4845 ;
  assign n4847 = n4639 & ~n4846 ;
  assign n4647 = \P1_InstQueue_reg[10][2]/NET0131  & n1978 ;
  assign n4648 = \P1_InstQueue_reg[6][2]/NET0131  & n1964 ;
  assign n4663 = ~n4647 & ~n4648 ;
  assign n4649 = \P1_InstQueue_reg[5][2]/NET0131  & n1961 ;
  assign n4650 = \P1_InstQueue_reg[13][2]/NET0131  & n1953 ;
  assign n4664 = ~n4649 & ~n4650 ;
  assign n4670 = n4663 & n4664 ;
  assign n4643 = \P1_InstQueue_reg[3][2]/NET0131  & n1970 ;
  assign n4644 = \P1_InstQueue_reg[11][2]/NET0131  & n1946 ;
  assign n4661 = ~n4643 & ~n4644 ;
  assign n4645 = \P1_InstQueue_reg[8][2]/NET0131  & n1968 ;
  assign n4646 = \P1_InstQueue_reg[14][2]/NET0131  & n1980 ;
  assign n4662 = ~n4645 & ~n4646 ;
  assign n4671 = n4661 & n4662 ;
  assign n4672 = n4670 & n4671 ;
  assign n4658 = ~\P1_InstQueueRd_Addr_reg[2]/NET0131  & \P1_InstQueue_reg[2][2]/NET0131  ;
  assign n4659 = n1963 & n4658 ;
  assign n4660 = n2348 & n4659 ;
  assign n4657 = \P1_InstQueue_reg[4][2]/NET0131  & n1976 ;
  assign n4655 = \P1_InstQueue_reg[1][2]/NET0131  & n1958 ;
  assign n4656 = \P1_InstQueue_reg[7][2]/NET0131  & n1972 ;
  assign n4667 = ~n4655 & ~n4656 ;
  assign n4668 = ~n4657 & n4667 ;
  assign n4651 = \P1_InstQueue_reg[12][2]/NET0131  & n1949 ;
  assign n4652 = \P1_InstQueue_reg[0][2]/NET0131  & n1982 ;
  assign n4665 = ~n4651 & ~n4652 ;
  assign n4653 = \P1_InstQueue_reg[9][2]/NET0131  & n1974 ;
  assign n4654 = \P1_InstQueue_reg[15][2]/NET0131  & n1955 ;
  assign n4666 = ~n4653 & ~n4654 ;
  assign n4669 = n4665 & n4666 ;
  assign n4673 = n4668 & n4669 ;
  assign n4674 = ~n4660 & n4673 ;
  assign n4675 = n4672 & n4674 ;
  assign n4848 = ~\P1_InstAddrPointer_reg[2]/NET0131  & ~n4813 ;
  assign n4849 = ~n4814 & ~n4848 ;
  assign n4850 = n4675 & ~n4849 ;
  assign n4851 = ~n4847 & ~n4850 ;
  assign n4852 = n4844 & n4851 ;
  assign n4853 = ~n4639 & n4846 ;
  assign n4854 = ~n4675 & n4849 ;
  assign n4855 = ~n4847 & n4854 ;
  assign n4856 = ~n4853 & ~n4855 ;
  assign n4857 = ~n4852 & n4856 ;
  assign n4858 = ~n4838 & ~n4857 ;
  assign n4859 = ~n4607 & n4837 ;
  assign n4860 = ~n4573 & n4829 ;
  assign n4861 = ~n4859 & ~n4860 ;
  assign n4862 = ~n4858 & n4861 ;
  assign n4863 = n4835 & ~n4862 ;
  assign n4864 = ~n4453 & n4826 ;
  assign n4865 = ~n4539 & n4832 ;
  assign n4866 = ~n4864 & ~n4865 ;
  assign n4867 = ~n4827 & ~n4866 ;
  assign n4868 = ~\P1_InstAddrPointer_reg[8]/NET0131  & ~n4819 ;
  assign n4869 = ~n4820 & ~n4868 ;
  assign n4870 = ~\P1_InstAddrPointer_reg[9]/NET0131  & ~n4820 ;
  assign n4871 = ~n4821 & ~n4870 ;
  assign n4872 = ~n4869 & ~n4871 ;
  assign n4873 = ~n4867 & n4872 ;
  assign n4874 = ~n4863 & n4873 ;
  assign n4875 = ~n4824 & n4874 ;
  assign n4876 = ~\P1_InstAddrPointer_reg[11]/NET0131  & ~n4823 ;
  assign n4877 = n4463 & n4818 ;
  assign n4878 = ~n4876 & ~n4877 ;
  assign n4786 = \P1_InstAddrPointer_reg[12]/NET0131  & n4464 ;
  assign n4879 = \P1_InstAddrPointer_reg[0]/NET0131  & n4786 ;
  assign n4880 = ~\P1_InstAddrPointer_reg[13]/NET0131  & ~n4879 ;
  assign n4881 = n4454 & n4877 ;
  assign n4882 = ~n4880 & ~n4881 ;
  assign n4883 = ~\P1_InstAddrPointer_reg[12]/NET0131  & ~n4877 ;
  assign n4884 = ~n4879 & ~n4883 ;
  assign n4885 = ~n4882 & ~n4884 ;
  assign n4886 = ~n4878 & n4885 ;
  assign n4887 = n4875 & n4886 ;
  assign n4888 = n4467 & n4881 ;
  assign n4889 = n4470 & n4888 ;
  assign n4890 = n4478 & n4889 ;
  assign n4891 = ~\P1_InstAddrPointer_reg[24]/NET0131  & ~n4890 ;
  assign n4892 = \P1_InstAddrPointer_reg[0]/NET0131  & n4483 ;
  assign n4893 = ~n4891 & ~n4892 ;
  assign n4473 = n4471 & n4472 ;
  assign n4475 = \P1_InstAddrPointer_reg[22]/NET0131  & n4473 ;
  assign n4894 = \P1_InstAddrPointer_reg[0]/NET0131  & n4475 ;
  assign n4895 = ~\P1_InstAddrPointer_reg[23]/NET0131  & ~n4894 ;
  assign n4896 = ~n4890 & ~n4895 ;
  assign n4767 = \P1_InstAddrPointer_reg[20]/NET0131  & n4471 ;
  assign n4897 = \P1_InstAddrPointer_reg[0]/NET0131  & n4767 ;
  assign n4898 = ~\P1_InstAddrPointer_reg[21]/NET0131  & ~n4897 ;
  assign n4899 = n4472 & n4889 ;
  assign n4900 = ~n4898 & ~n4899 ;
  assign n4901 = ~\P1_InstAddrPointer_reg[22]/NET0131  & ~n4899 ;
  assign n4902 = ~n4894 & ~n4901 ;
  assign n4903 = ~n4900 & ~n4902 ;
  assign n4904 = ~n4896 & n4903 ;
  assign n4905 = ~n4893 & n4904 ;
  assign n4906 = ~\P1_InstAddrPointer_reg[25]/NET0131  & ~n4892 ;
  assign n4907 = \P1_InstAddrPointer_reg[25]/NET0131  & n4892 ;
  assign n4908 = ~n4906 & ~n4907 ;
  assign n4909 = n4905 & ~n4908 ;
  assign n4782 = n4465 & n4466 ;
  assign n4910 = \P1_InstAddrPointer_reg[0]/NET0131  & n4782 ;
  assign n4911 = \P1_InstAddrPointer_reg[14]/NET0131  & n4881 ;
  assign n4912 = ~\P1_InstAddrPointer_reg[15]/NET0131  & ~n4911 ;
  assign n4913 = ~n4910 & ~n4912 ;
  assign n4773 = \P1_InstAddrPointer_reg[17]/NET0131  & n4468 ;
  assign n4914 = \P1_InstAddrPointer_reg[0]/NET0131  & n4773 ;
  assign n4919 = ~\P1_InstAddrPointer_reg[18]/NET0131  & ~n4914 ;
  assign n4775 = n4468 & n4469 ;
  assign n4920 = \P1_InstAddrPointer_reg[0]/NET0131  & n4775 ;
  assign n4921 = ~n4919 & ~n4920 ;
  assign n4915 = ~\P1_InstAddrPointer_reg[17]/NET0131  & ~n4888 ;
  assign n4916 = ~n4914 & ~n4915 ;
  assign n4917 = ~\P1_InstAddrPointer_reg[16]/NET0131  & ~n4910 ;
  assign n4918 = ~n4888 & ~n4917 ;
  assign n4922 = ~n4916 & ~n4918 ;
  assign n4923 = ~n4921 & n4922 ;
  assign n4924 = ~n4913 & n4923 ;
  assign n4925 = ~\P1_InstAddrPointer_reg[19]/NET0131  & ~n4920 ;
  assign n4926 = ~n4889 & ~n4925 ;
  assign n4927 = ~\P1_InstAddrPointer_reg[20]/NET0131  & ~n4889 ;
  assign n4928 = ~n4897 & ~n4927 ;
  assign n4929 = ~n4926 & ~n4928 ;
  assign n4930 = ~\P1_InstAddrPointer_reg[14]/NET0131  & ~n4881 ;
  assign n4931 = ~n4911 & ~n4930 ;
  assign n4932 = n4929 & ~n4931 ;
  assign n4933 = n4924 & n4932 ;
  assign n4934 = n4909 & n4933 ;
  assign n4935 = n4887 & n4934 ;
  assign n4936 = ~\P1_InstAddrPointer_reg[28]/NET0131  & ~n4807 ;
  assign n4937 = ~n4808 & ~n4936 ;
  assign n4938 = ~\P1_InstAddrPointer_reg[26]/NET0131  & ~n4907 ;
  assign n4939 = \P1_InstAddrPointer_reg[0]/NET0131  & n4489 ;
  assign n4940 = ~n4938 & ~n4939 ;
  assign n4941 = ~\P1_InstAddrPointer_reg[27]/NET0131  & ~n4939 ;
  assign n4942 = ~n4807 & ~n4941 ;
  assign n4943 = ~n4940 & ~n4942 ;
  assign n4944 = ~n4937 & n4943 ;
  assign n4945 = ~\P1_InstAddrPointer_reg[29]/NET0131  & ~n4808 ;
  assign n4946 = ~n4809 & ~n4945 ;
  assign n4947 = n4944 & ~n4946 ;
  assign n4948 = n4935 & n4947 ;
  assign n4950 = ~n4812 & n4948 ;
  assign n4949 = n4812 & ~n4948 ;
  assign n4951 = ~n4453 & ~n4949 ;
  assign n4952 = ~n4950 & n4951 ;
  assign n4498 = ~\P1_InstAddrPointer_reg[9]/NET0131  & ~n4496 ;
  assign n4499 = ~n4497 & ~n4498 ;
  assign n4500 = \P1_InstAddrPointer_reg[7]/NET0131  & n4459 ;
  assign n4501 = ~\P1_InstAddrPointer_reg[8]/NET0131  & ~n4500 ;
  assign n4502 = ~n4496 & ~n4501 ;
  assign n4503 = ~\P1_InstAddrPointer_reg[7]/NET0131  & ~n4459 ;
  assign n4504 = ~n4500 & ~n4503 ;
  assign n4505 = n4453 & ~n4504 ;
  assign n4506 = n4502 & ~n4505 ;
  assign n4676 = ~\P1_InstAddrPointer_reg[1]/NET0131  & ~\P1_InstAddrPointer_reg[2]/NET0131  ;
  assign n4677 = ~n4455 & ~n4676 ;
  assign n4678 = ~n4675 & n4677 ;
  assign n4679 = n4675 & ~n4677 ;
  assign n4712 = \P1_InstAddrPointer_reg[1]/NET0131  & n4710 ;
  assign n4744 = \P1_InstAddrPointer_reg[0]/NET0131  & ~n4743 ;
  assign n4745 = ~n4712 & n4744 ;
  assign n4746 = ~n4711 & ~n4745 ;
  assign n4747 = ~n4679 & ~n4746 ;
  assign n4748 = ~n4678 & ~n4747 ;
  assign n4575 = ~\P1_InstAddrPointer_reg[4]/NET0131  & ~n4456 ;
  assign n4576 = ~n4457 & ~n4575 ;
  assign n4608 = ~n4576 & n4607 ;
  assign n4640 = ~\P1_InstAddrPointer_reg[3]/NET0131  & ~n4455 ;
  assign n4641 = ~n4456 & ~n4640 ;
  assign n4642 = n4639 & ~n4641 ;
  assign n4749 = ~n4608 & ~n4642 ;
  assign n4750 = ~n4748 & n4749 ;
  assign n4751 = n4576 & ~n4607 ;
  assign n4752 = ~n4639 & n4641 ;
  assign n4753 = ~n4608 & n4752 ;
  assign n4754 = ~n4751 & ~n4753 ;
  assign n4755 = ~n4750 & n4754 ;
  assign n4507 = ~\P1_InstAddrPointer_reg[6]/NET0131  & ~n4458 ;
  assign n4508 = ~n4459 & ~n4507 ;
  assign n4540 = ~n4508 & n4539 ;
  assign n4541 = ~\P1_InstAddrPointer_reg[5]/NET0131  & ~n4457 ;
  assign n4542 = ~n4458 & ~n4541 ;
  assign n4574 = ~n4542 & n4573 ;
  assign n4756 = ~n4540 & ~n4574 ;
  assign n4757 = ~n4755 & n4756 ;
  assign n4758 = ~n4453 & n4504 ;
  assign n4759 = n4508 & ~n4539 ;
  assign n4760 = n4542 & ~n4573 ;
  assign n4761 = ~n4540 & n4760 ;
  assign n4762 = ~n4759 & ~n4761 ;
  assign n4763 = ~n4758 & n4762 ;
  assign n4764 = ~n4757 & n4763 ;
  assign n4765 = n4506 & ~n4764 ;
  assign n4766 = n4499 & n4765 ;
  assign n4783 = ~\P1_InstAddrPointer_reg[16]/NET0131  & ~n4782 ;
  assign n4784 = ~n4468 & ~n4783 ;
  assign n4785 = \P1_InstAddrPointer_reg[17]/NET0131  & n4784 ;
  assign n4779 = ~\P1_InstAddrPointer_reg[11]/NET0131  & ~n4771 ;
  assign n4780 = ~n4464 & ~n4779 ;
  assign n4781 = \P1_InstAddrPointer_reg[12]/NET0131  & n4780 ;
  assign n4787 = ~\P1_InstAddrPointer_reg[13]/NET0131  & ~n4786 ;
  assign n4788 = ~n4465 & ~n4787 ;
  assign n4789 = n4466 & n4788 ;
  assign n4790 = n4781 & n4789 ;
  assign n4791 = n4785 & n4790 ;
  assign n4774 = ~\P1_InstAddrPointer_reg[18]/NET0131  & ~n4773 ;
  assign n4776 = ~n4774 & ~n4775 ;
  assign n4777 = \P1_InstAddrPointer_reg[19]/NET0131  & n4776 ;
  assign n4778 = \P1_InstAddrPointer_reg[20]/NET0131  & n4777 ;
  assign n4768 = ~\P1_InstAddrPointer_reg[21]/NET0131  & ~n4767 ;
  assign n4769 = ~n4473 & ~n4768 ;
  assign n4770 = ~\P1_InstAddrPointer_reg[10]/NET0131  & ~n4497 ;
  assign n4772 = ~n4770 & ~n4771 ;
  assign n4792 = n4769 & n4772 ;
  assign n4793 = n4778 & n4792 ;
  assign n4794 = n4791 & n4793 ;
  assign n4795 = n4766 & n4794 ;
  assign n4474 = ~\P1_InstAddrPointer_reg[22]/NET0131  & ~n4473 ;
  assign n4476 = ~n4474 & ~n4475 ;
  assign n4491 = ~\P1_InstAddrPointer_reg[27]/NET0131  & ~n4489 ;
  assign n4492 = ~n4490 & ~n4491 ;
  assign n4480 = ~\P1_InstAddrPointer_reg[23]/NET0131  & ~n4475 ;
  assign n4481 = ~n4479 & ~n4480 ;
  assign n4482 = \P1_InstAddrPointer_reg[24]/NET0131  & n4481 ;
  assign n4485 = ~\P1_InstAddrPointer_reg[25]/NET0131  & ~n4483 ;
  assign n4486 = ~n4484 & ~n4485 ;
  assign n4487 = \P1_InstAddrPointer_reg[26]/NET0131  & n4486 ;
  assign n4488 = n4482 & n4487 ;
  assign n4493 = \P1_InstAddrPointer_reg[28]/NET0131  & n4488 ;
  assign n4494 = n4492 & n4493 ;
  assign n4495 = \P1_InstAddrPointer_reg[29]/NET0131  & n4494 ;
  assign n4796 = n4476 & n4495 ;
  assign n4797 = n4795 & n4796 ;
  assign n4798 = \P1_InstAddrPointer_reg[28]/NET0131  & \P1_InstAddrPointer_reg[29]/NET0131  ;
  assign n4799 = n4490 & n4798 ;
  assign n4800 = \P1_InstAddrPointer_reg[30]/NET0131  & n4799 ;
  assign n4801 = ~\P1_InstAddrPointer_reg[30]/NET0131  & ~n4799 ;
  assign n4802 = ~n4800 & ~n4801 ;
  assign n4804 = n4797 & ~n4802 ;
  assign n4803 = ~n4797 & n4802 ;
  assign n4805 = n4453 & ~n4803 ;
  assign n4806 = ~n4804 & n4805 ;
  assign n4953 = ~n2375 & ~n4806 ;
  assign n4954 = ~n4952 & n4953 ;
  assign n4955 = ~n4422 & ~n4954 ;
  assign n4956 = n2244 & ~n4955 ;
  assign n4957 = \P1_InstAddrPointer_reg[3]/NET0131  & ~n4848 ;
  assign n4958 = \P1_InstAddrPointer_reg[4]/NET0131  & n4957 ;
  assign n4959 = \P1_InstAddrPointer_reg[5]/NET0131  & n4958 ;
  assign n4984 = ~\P1_InstAddrPointer_reg[5]/NET0131  & ~n4958 ;
  assign n4985 = ~n4959 & ~n4984 ;
  assign n4986 = n4573 & ~n4985 ;
  assign n4987 = ~\P1_InstAddrPointer_reg[4]/NET0131  & ~n4957 ;
  assign n4988 = ~n4958 & ~n4987 ;
  assign n4989 = n4607 & ~n4988 ;
  assign n4990 = ~n4986 & ~n4989 ;
  assign n4991 = ~\P1_InstAddrPointer_reg[3]/NET0131  & n4848 ;
  assign n4992 = ~n4957 & ~n4991 ;
  assign n4993 = n4639 & ~n4992 ;
  assign n4994 = n4675 & n4849 ;
  assign n4995 = ~n4993 & ~n4994 ;
  assign n4996 = ~n4710 & n4840 ;
  assign n4997 = ~\P1_InstAddrPointer_reg[0]/NET0131  & ~n4743 ;
  assign n4998 = ~n4996 & ~n4997 ;
  assign n4999 = ~n4841 & ~n4998 ;
  assign n5000 = n4995 & n4999 ;
  assign n5001 = ~n4639 & n4992 ;
  assign n5002 = ~n4675 & ~n4849 ;
  assign n5003 = ~n4993 & n5002 ;
  assign n5004 = ~n5001 & ~n5003 ;
  assign n5005 = ~n5000 & n5004 ;
  assign n5006 = n4990 & ~n5005 ;
  assign n5007 = ~n4573 & n4985 ;
  assign n5008 = ~n4607 & n4988 ;
  assign n5009 = ~n4986 & n5008 ;
  assign n5010 = ~n5007 & ~n5009 ;
  assign n5011 = ~n5006 & n5010 ;
  assign n4960 = \P1_InstAddrPointer_reg[6]/NET0131  & n4959 ;
  assign n4975 = \P1_InstAddrPointer_reg[7]/NET0131  & n4960 ;
  assign n4978 = ~\P1_InstAddrPointer_reg[7]/NET0131  & ~n4960 ;
  assign n4979 = ~n4975 & ~n4978 ;
  assign n4980 = n4453 & ~n4979 ;
  assign n4981 = ~\P1_InstAddrPointer_reg[6]/NET0131  & ~n4959 ;
  assign n4982 = ~n4960 & ~n4981 ;
  assign n4983 = n4539 & ~n4982 ;
  assign n5012 = ~n4980 & ~n4983 ;
  assign n5013 = ~n5011 & n5012 ;
  assign n5014 = ~n4453 & n4979 ;
  assign n5015 = ~n4539 & n4982 ;
  assign n5016 = ~n4980 & n5015 ;
  assign n5017 = ~n5014 & ~n5016 ;
  assign n5018 = ~n5013 & n5017 ;
  assign n4961 = n4461 & n4960 ;
  assign n4976 = ~\P1_InstAddrPointer_reg[8]/NET0131  & ~n4975 ;
  assign n4977 = ~n4961 & ~n4976 ;
  assign n5019 = \P1_InstAddrPointer_reg[9]/NET0131  & n4977 ;
  assign n5020 = ~n5018 & n5019 ;
  assign n4962 = n4460 & n4961 ;
  assign n5021 = \P1_InstAddrPointer_reg[9]/NET0131  & n4961 ;
  assign n5022 = ~\P1_InstAddrPointer_reg[10]/NET0131  & ~n5021 ;
  assign n5023 = ~n4962 & ~n5022 ;
  assign n5024 = n5020 & n5023 ;
  assign n4963 = \P1_InstAddrPointer_reg[11]/NET0131  & n4962 ;
  assign n5025 = ~\P1_InstAddrPointer_reg[11]/NET0131  & ~n4962 ;
  assign n5026 = ~n4963 & ~n5025 ;
  assign n5027 = n4454 & n5026 ;
  assign n5028 = n5024 & n5027 ;
  assign n4964 = \P1_InstAddrPointer_reg[12]/NET0131  & n4963 ;
  assign n4965 = \P1_InstAddrPointer_reg[13]/NET0131  & n4964 ;
  assign n4966 = n4467 & n4965 ;
  assign n5029 = \P1_InstAddrPointer_reg[14]/NET0131  & n4965 ;
  assign n5030 = \P1_InstAddrPointer_reg[15]/NET0131  & n5029 ;
  assign n5031 = ~\P1_InstAddrPointer_reg[16]/NET0131  & ~n5030 ;
  assign n5032 = ~n4966 & ~n5031 ;
  assign n5033 = ~\P1_InstAddrPointer_reg[14]/NET0131  & ~n4965 ;
  assign n5034 = ~n5029 & ~n5033 ;
  assign n5035 = \P1_InstAddrPointer_reg[15]/NET0131  & \P1_InstAddrPointer_reg[17]/NET0131  ;
  assign n5036 = n5034 & n5035 ;
  assign n5037 = n5032 & n5036 ;
  assign n5038 = n5028 & n5037 ;
  assign n4967 = \P1_InstAddrPointer_reg[17]/NET0131  & n4966 ;
  assign n4968 = ~\P1_InstAddrPointer_reg[18]/NET0131  & ~n4967 ;
  assign n4969 = n4469 & n4966 ;
  assign n4970 = ~n4968 & ~n4969 ;
  assign n4971 = ~\P1_InstAddrPointer_reg[19]/NET0131  & ~n4969 ;
  assign n4972 = n4470 & n4966 ;
  assign n4973 = ~n4971 & ~n4972 ;
  assign n4974 = n4472 & n4973 ;
  assign n5039 = n4970 & n4974 ;
  assign n5040 = n5038 & n5039 ;
  assign n5041 = n4478 & n4972 ;
  assign n5042 = \P1_InstAddrPointer_reg[24]/NET0131  & n5041 ;
  assign n5043 = ~\P1_InstAddrPointer_reg[25]/NET0131  & ~n5042 ;
  assign n5044 = \P1_InstAddrPointer_reg[25]/NET0131  & n5042 ;
  assign n5045 = ~n5043 & ~n5044 ;
  assign n5046 = n4472 & n4972 ;
  assign n5047 = ~\P1_InstAddrPointer_reg[22]/NET0131  & ~n5046 ;
  assign n5048 = \P1_InstAddrPointer_reg[22]/NET0131  & n5046 ;
  assign n5049 = ~n5047 & ~n5048 ;
  assign n5050 = \P1_InstAddrPointer_reg[23]/NET0131  & n5049 ;
  assign n5051 = \P1_InstAddrPointer_reg[24]/NET0131  & n5050 ;
  assign n5052 = n5045 & n5051 ;
  assign n5053 = n5040 & n5052 ;
  assign n5054 = ~\P1_InstAddrPointer_reg[26]/NET0131  & ~n5044 ;
  assign n5055 = \P1_InstAddrPointer_reg[26]/NET0131  & n5044 ;
  assign n5056 = ~n5054 & ~n5055 ;
  assign n5057 = n5053 & n5056 ;
  assign n5058 = \P1_InstAddrPointer_reg[27]/NET0131  & n5055 ;
  assign n5059 = ~\P1_InstAddrPointer_reg[27]/NET0131  & ~n5055 ;
  assign n5060 = ~n5058 & ~n5059 ;
  assign n5061 = n4798 & n5060 ;
  assign n5062 = n5057 & n5061 ;
  assign n5063 = n4798 & n5058 ;
  assign n5064 = ~\P1_InstAddrPointer_reg[30]/NET0131  & ~n5063 ;
  assign n5065 = \P1_InstAddrPointer_reg[30]/NET0131  & n5063 ;
  assign n5066 = ~n5064 & ~n5065 ;
  assign n5067 = ~n5062 & ~n5066 ;
  assign n5068 = \P1_InstAddrPointer_reg[30]/NET0131  & n5061 ;
  assign n5069 = n5057 & n5068 ;
  assign n5070 = n2385 & ~n5069 ;
  assign n5071 = ~n5067 & n5070 ;
  assign n5074 = n2337 & ~n5066 ;
  assign n5073 = ~\P1_InstAddrPointer_reg[30]/NET0131  & ~n2337 ;
  assign n5075 = ~n2332 & ~n5073 ;
  assign n5076 = ~n5074 & n5075 ;
  assign n5078 = n2377 & ~n4802 ;
  assign n5079 = ~n2222 & n2306 ;
  assign n5080 = n2301 & ~n5079 ;
  assign n5081 = ~n2302 & ~n5080 ;
  assign n5082 = ~n5078 & ~n5081 ;
  assign n5083 = ~n2369 & n2390 ;
  assign n5084 = ~n5082 & n5083 ;
  assign n5085 = \P1_InstAddrPointer_reg[30]/NET0131  & ~n5084 ;
  assign n5072 = ~n2271 & n4812 ;
  assign n5077 = ~n2402 & n4802 ;
  assign n5086 = ~n5072 & ~n5077 ;
  assign n5087 = ~n5085 & n5086 ;
  assign n5088 = ~n5076 & n5087 ;
  assign n5089 = ~n5071 & n5088 ;
  assign n5090 = ~n4956 & n5089 ;
  assign n5091 = n2432 & ~n5090 ;
  assign n5092 = n3017 & n3026 ;
  assign n5093 = \P1_rEIP_reg[30]/NET0131  & n5092 ;
  assign n5094 = ~n3017 & n3026 ;
  assign n5095 = ~\P1_State2_reg[0]/NET0131  & n2431 ;
  assign n5096 = ~n2435 & ~n2439 ;
  assign n5097 = ~n5095 & n5096 ;
  assign n5098 = ~n5094 & n5097 ;
  assign n5099 = \P1_InstAddrPointer_reg[30]/NET0131  & ~n5098 ;
  assign n5100 = ~n5093 & ~n5099 ;
  assign n5101 = ~n5091 & n5100 ;
  assign n5146 = ~\P1_InstQueueWr_Addr_reg[0]/NET0131  & ~\P1_InstQueueWr_Addr_reg[1]/NET0131  ;
  assign n5147 = ~\P1_InstQueueWr_Addr_reg[2]/NET0131  & n5146 ;
  assign n5148 = \P1_InstQueueWr_Addr_reg[3]/NET0131  & n5147 ;
  assign n5149 = \P1_InstQueueWr_Addr_reg[0]/NET0131  & ~\P1_InstQueueWr_Addr_reg[1]/NET0131  ;
  assign n5150 = ~\P1_InstQueueWr_Addr_reg[2]/NET0131  & n5149 ;
  assign n5151 = \P1_InstQueueWr_Addr_reg[3]/NET0131  & n5150 ;
  assign n5152 = ~n5148 & ~n5151 ;
  assign n5153 = \P1_DataWidth_reg[1]/NET0131  & ~n5152 ;
  assign n5118 = ~\address1[26]_pad  & ~\address1[27]_pad  ;
  assign n5119 = ~\address1[28]_pad  & ~\address1[2]_pad  ;
  assign n5125 = n5118 & n5119 ;
  assign n5116 = ~\address1[22]_pad  & ~\address1[23]_pad  ;
  assign n5117 = ~\address1[24]_pad  & ~\address1[25]_pad  ;
  assign n5126 = n5116 & n5117 ;
  assign n5132 = n5125 & n5126 ;
  assign n5122 = ~\address1[7]_pad  & ~\address1[8]_pad  ;
  assign n5123 = ~\address1[9]_pad  & n5122 ;
  assign n5120 = ~\address1[3]_pad  & ~\address1[4]_pad  ;
  assign n5121 = ~\address1[5]_pad  & ~\address1[6]_pad  ;
  assign n5124 = n5120 & n5121 ;
  assign n5133 = n5123 & n5124 ;
  assign n5134 = n5132 & n5133 ;
  assign n5109 = ~\address1[0]_pad  & ~\address1[10]_pad  ;
  assign n5110 = ~\address1[11]_pad  & ~\address1[12]_pad  ;
  assign n5111 = ~\address1[13]_pad  & ~\address1[14]_pad  ;
  assign n5129 = n5110 & n5111 ;
  assign n5130 = n5109 & n5129 ;
  assign n5114 = ~\address1[19]_pad  & ~\address1[1]_pad  ;
  assign n5115 = ~\address1[20]_pad  & ~\address1[21]_pad  ;
  assign n5127 = n5114 & n5115 ;
  assign n5112 = ~\address1[15]_pad  & ~\address1[16]_pad  ;
  assign n5113 = ~\address1[17]_pad  & ~\address1[18]_pad  ;
  assign n5128 = n5112 & n5113 ;
  assign n5131 = n5127 & n5128 ;
  assign n5135 = n5130 & n5131 ;
  assign n5136 = n5134 & n5135 ;
  assign n5137 = \address1[29]_pad  & ~n5136 ;
  assign n5155 = \datai[31]_pad  & ~n5137 ;
  assign n5165 = \datai[3]_pad  & ~n5137 ;
  assign n5166 = \buf1_reg[3]/NET0131  & n5137 ;
  assign n5167 = ~n5165 & ~n5166 ;
  assign n5168 = \datai[11]_pad  & ~n5137 ;
  assign n5169 = \buf1_reg[11]/NET0131  & n5137 ;
  assign n5170 = ~n5168 & ~n5169 ;
  assign n5203 = n5167 & n5170 ;
  assign n5171 = \datai[8]_pad  & ~n5137 ;
  assign n5172 = \buf1_reg[8]/NET0131  & n5137 ;
  assign n5173 = ~n5171 & ~n5172 ;
  assign n5174 = \datai[7]_pad  & ~n5137 ;
  assign n5175 = \buf1_reg[7]/NET0131  & n5137 ;
  assign n5176 = ~n5174 & ~n5175 ;
  assign n5204 = n5173 & n5176 ;
  assign n5211 = n5203 & n5204 ;
  assign n5138 = \datai[4]_pad  & ~n5137 ;
  assign n5139 = \buf1_reg[4]/NET0131  & n5137 ;
  assign n5140 = ~n5138 & ~n5139 ;
  assign n5156 = \datai[9]_pad  & ~n5137 ;
  assign n5157 = \buf1_reg[9]/NET0131  & n5137 ;
  assign n5158 = ~n5156 & ~n5157 ;
  assign n5201 = n5140 & n5158 ;
  assign n5159 = \datai[10]_pad  & ~n5137 ;
  assign n5160 = \buf1_reg[10]/NET0131  & n5137 ;
  assign n5161 = ~n5159 & ~n5160 ;
  assign n5162 = \datai[5]_pad  & ~n5137 ;
  assign n5163 = \buf1_reg[5]/NET0131  & n5137 ;
  assign n5164 = ~n5162 & ~n5163 ;
  assign n5202 = n5161 & n5164 ;
  assign n5212 = n5201 & n5202 ;
  assign n5213 = n5211 & n5212 ;
  assign n5189 = \datai[14]_pad  & ~n5137 ;
  assign n5190 = \buf1_reg[14]/NET0131  & n5137 ;
  assign n5191 = ~n5189 & ~n5190 ;
  assign n5192 = \datai[15]_pad  & ~n5137 ;
  assign n5193 = \buf1_reg[15]/NET0131  & n5137 ;
  assign n5194 = ~n5192 & ~n5193 ;
  assign n5207 = n5191 & n5194 ;
  assign n5195 = \datai[12]_pad  & ~n5137 ;
  assign n5196 = \buf1_reg[12]/NET0131  & n5137 ;
  assign n5197 = ~n5195 & ~n5196 ;
  assign n5198 = \datai[13]_pad  & ~n5137 ;
  assign n5199 = \buf1_reg[13]/NET0131  & n5137 ;
  assign n5200 = ~n5198 & ~n5199 ;
  assign n5208 = n5197 & n5200 ;
  assign n5209 = n5207 & n5208 ;
  assign n5177 = \datai[0]_pad  & ~n5137 ;
  assign n5178 = \buf1_reg[0]/NET0131  & n5137 ;
  assign n5179 = ~n5177 & ~n5178 ;
  assign n5180 = \datai[6]_pad  & ~n5137 ;
  assign n5181 = \buf1_reg[6]/NET0131  & n5137 ;
  assign n5182 = ~n5180 & ~n5181 ;
  assign n5205 = n5179 & n5182 ;
  assign n5183 = \datai[1]_pad  & ~n5137 ;
  assign n5184 = \buf1_reg[1]/NET0131  & n5137 ;
  assign n5185 = ~n5183 & ~n5184 ;
  assign n5186 = \datai[2]_pad  & ~n5137 ;
  assign n5187 = \buf1_reg[2]/NET0131  & n5137 ;
  assign n5188 = ~n5186 & ~n5187 ;
  assign n5206 = n5185 & n5188 ;
  assign n5210 = n5205 & n5206 ;
  assign n5214 = n5209 & n5210 ;
  assign n5215 = n5213 & n5214 ;
  assign n5228 = \datai[19]_pad  & ~n5137 ;
  assign n5229 = \buf1_reg[19]/NET0131  & n5137 ;
  assign n5230 = ~n5228 & ~n5229 ;
  assign n5231 = \datai[18]_pad  & ~n5137 ;
  assign n5232 = \buf1_reg[18]/NET0131  & n5137 ;
  assign n5233 = ~n5231 & ~n5232 ;
  assign n5242 = n5230 & n5233 ;
  assign n5234 = \datai[17]_pad  & ~n5137 ;
  assign n5235 = \buf1_reg[17]/NET0131  & n5137 ;
  assign n5236 = ~n5234 & ~n5235 ;
  assign n5237 = \datai[20]_pad  & ~n5137 ;
  assign n5238 = \buf1_reg[20]/NET0131  & n5137 ;
  assign n5239 = ~n5237 & ~n5238 ;
  assign n5243 = n5236 & n5239 ;
  assign n5244 = n5242 & n5243 ;
  assign n5216 = \datai[16]_pad  & ~n5137 ;
  assign n5217 = \buf1_reg[16]/NET0131  & n5137 ;
  assign n5218 = ~n5216 & ~n5217 ;
  assign n5219 = \datai[22]_pad  & ~n5137 ;
  assign n5220 = \buf1_reg[22]/NET0131  & n5137 ;
  assign n5221 = ~n5219 & ~n5220 ;
  assign n5240 = n5218 & n5221 ;
  assign n5222 = \datai[23]_pad  & ~n5137 ;
  assign n5223 = \buf1_reg[23]/NET0131  & n5137 ;
  assign n5224 = ~n5222 & ~n5223 ;
  assign n5225 = \datai[21]_pad  & ~n5137 ;
  assign n5226 = \buf1_reg[21]/NET0131  & n5137 ;
  assign n5227 = ~n5225 & ~n5226 ;
  assign n5241 = n5224 & n5227 ;
  assign n5245 = n5240 & n5241 ;
  assign n5246 = n5244 & n5245 ;
  assign n5247 = n5215 & n5246 ;
  assign n5248 = n5155 & ~n5247 ;
  assign n5249 = \datai[24]_pad  & ~n5137 ;
  assign n5250 = \buf1_reg[24]/NET0131  & n5137 ;
  assign n5251 = ~n5249 & ~n5250 ;
  assign n5252 = n5248 & ~n5251 ;
  assign n5253 = \datai[25]_pad  & ~n5137 ;
  assign n5254 = \buf1_reg[25]/NET0131  & n5137 ;
  assign n5255 = ~n5253 & ~n5254 ;
  assign n5256 = n5252 & ~n5255 ;
  assign n5257 = \datai[26]_pad  & ~n5137 ;
  assign n5258 = \buf1_reg[26]/NET0131  & n5137 ;
  assign n5259 = ~n5257 & ~n5258 ;
  assign n5260 = n5256 & ~n5259 ;
  assign n5261 = \datai[27]_pad  & ~n5137 ;
  assign n5262 = \buf1_reg[27]/NET0131  & n5137 ;
  assign n5263 = ~n5261 & ~n5262 ;
  assign n5264 = n5260 & ~n5263 ;
  assign n5265 = \datai[28]_pad  & ~n5137 ;
  assign n5266 = \buf1_reg[28]/NET0131  & n5137 ;
  assign n5267 = ~n5265 & ~n5266 ;
  assign n5268 = ~n5264 & n5267 ;
  assign n5269 = n5264 & ~n5267 ;
  assign n5270 = ~n5268 & ~n5269 ;
  assign n5271 = n5148 & ~n5270 ;
  assign n5272 = n5155 & ~n5215 ;
  assign n5273 = ~n5218 & n5272 ;
  assign n5274 = ~n5236 & n5273 ;
  assign n5275 = ~n5233 & n5274 ;
  assign n5276 = ~n5230 & n5275 ;
  assign n5277 = ~n5239 & n5276 ;
  assign n5278 = n5239 & ~n5276 ;
  assign n5279 = ~n5277 & ~n5278 ;
  assign n5280 = ~n5148 & ~n5279 ;
  assign n5281 = ~n5271 & ~n5280 ;
  assign n5282 = n5153 & ~n5281 ;
  assign n5102 = \P1_InstQueueWr_Addr_reg[0]/NET0131  & \P1_InstQueueWr_Addr_reg[1]/NET0131  ;
  assign n5103 = ~\P1_InstQueueWr_Addr_reg[2]/NET0131  & n5102 ;
  assign n5104 = \P1_InstQueueWr_Addr_reg[3]/NET0131  & n5103 ;
  assign n5105 = ~\P1_InstQueueWr_Addr_reg[0]/NET0131  & \P1_InstQueueWr_Addr_reg[1]/NET0131  ;
  assign n5106 = ~\P1_InstQueueWr_Addr_reg[2]/NET0131  & n5105 ;
  assign n5107 = \P1_InstQueueWr_Addr_reg[3]/NET0131  & n5106 ;
  assign n5108 = ~n5104 & ~n5107 ;
  assign n5141 = ~n5108 & ~n5140 ;
  assign n5142 = \P1_InstQueue_reg[11][4]/NET0131  & ~n5104 ;
  assign n5143 = ~n5107 & n5142 ;
  assign n5144 = ~n5141 & ~n5143 ;
  assign n5154 = n5144 & ~n5153 ;
  assign n5283 = n2436 & ~n5154 ;
  assign n5284 = ~n5282 & n5283 ;
  assign n5145 = n5095 & ~n5144 ;
  assign n5285 = ~n2188 & n5104 ;
  assign n5286 = ~n5142 & ~n5285 ;
  assign n5287 = n3042 & ~n5286 ;
  assign n5289 = ~n2432 & ~n2439 ;
  assign n5288 = ~n2445 & ~n5092 ;
  assign n5290 = ~n3028 & n5288 ;
  assign n5291 = n5289 & n5290 ;
  assign n5292 = \P1_InstQueue_reg[11][4]/NET0131  & ~n5291 ;
  assign n5293 = ~n5287 & ~n5292 ;
  assign n5294 = ~n5145 & n5293 ;
  assign n5295 = ~n5284 & n5294 ;
  assign n5304 = \buf2_reg[27]/NET0131  & ~n3079 ;
  assign n5305 = \buf1_reg[27]/NET0131  & n3079 ;
  assign n5306 = ~n5304 & ~n5305 ;
  assign n5307 = n3091 & ~n5306 ;
  assign n5308 = \buf2_reg[19]/NET0131  & ~n3079 ;
  assign n5309 = \buf1_reg[19]/NET0131  & n3079 ;
  assign n5310 = ~n5308 & ~n5309 ;
  assign n5311 = n3098 & ~n5310 ;
  assign n5312 = ~n5307 & ~n5311 ;
  assign n5313 = \P2_DataWidth_reg[1]/NET0131  & ~n5312 ;
  assign n5296 = \buf2_reg[3]/NET0131  & ~n3079 ;
  assign n5297 = \buf1_reg[3]/NET0131  & n3079 ;
  assign n5298 = ~n5296 & ~n5297 ;
  assign n5299 = ~n3050 & ~n5298 ;
  assign n5300 = \P2_InstQueue_reg[11][3]/NET0131  & ~n3049 ;
  assign n5301 = ~n3046 & n5300 ;
  assign n5302 = ~n5299 & ~n5301 ;
  assign n5314 = ~n3106 & ~n5302 ;
  assign n5315 = ~n5313 & ~n5314 ;
  assign n5316 = n1931 & ~n5315 ;
  assign n5303 = n3087 & ~n5302 ;
  assign n5317 = ~n1529 & n3049 ;
  assign n5318 = ~n5300 & ~n5317 ;
  assign n5319 = n3040 & ~n5318 ;
  assign n5320 = \P2_InstQueue_reg[11][3]/NET0131  & ~n3118 ;
  assign n5321 = ~n5319 & ~n5320 ;
  assign n5322 = ~n5303 & n5321 ;
  assign n5323 = ~n5316 & n5322 ;
  assign n5333 = \P1_InstQueueWr_Addr_reg[2]/NET0131  & n5149 ;
  assign n5334 = \P1_InstQueueWr_Addr_reg[3]/NET0131  & n5333 ;
  assign n5335 = \P1_InstQueueWr_Addr_reg[2]/NET0131  & n5105 ;
  assign n5336 = \P1_InstQueueWr_Addr_reg[3]/NET0131  & n5335 ;
  assign n5337 = ~n5334 & ~n5336 ;
  assign n5338 = \P1_DataWidth_reg[1]/NET0131  & ~n5337 ;
  assign n5340 = ~n5270 & n5334 ;
  assign n5341 = ~n5279 & ~n5334 ;
  assign n5342 = ~n5340 & ~n5341 ;
  assign n5343 = n5338 & ~n5342 ;
  assign n5324 = ~\P1_InstQueueWr_Addr_reg[3]/NET0131  & n5147 ;
  assign n5325 = \P1_InstQueueWr_Addr_reg[2]/NET0131  & n5102 ;
  assign n5326 = \P1_InstQueueWr_Addr_reg[3]/NET0131  & n5325 ;
  assign n5327 = ~n5324 & ~n5326 ;
  assign n5328 = ~n5140 & ~n5327 ;
  assign n5329 = \P1_InstQueue_reg[0][4]/NET0131  & ~n5324 ;
  assign n5330 = ~n5326 & n5329 ;
  assign n5331 = ~n5328 & ~n5330 ;
  assign n5339 = n5331 & ~n5338 ;
  assign n5344 = n2436 & ~n5339 ;
  assign n5345 = ~n5343 & n5344 ;
  assign n5332 = n5095 & ~n5331 ;
  assign n5346 = ~n2188 & n5324 ;
  assign n5347 = ~n5329 & ~n5346 ;
  assign n5348 = n3042 & ~n5347 ;
  assign n5349 = \P1_InstQueue_reg[0][4]/NET0131  & ~n5291 ;
  assign n5350 = ~n5348 & ~n5349 ;
  assign n5351 = ~n5332 & n5350 ;
  assign n5352 = ~n5345 & n5351 ;
  assign n5359 = ~\P1_InstQueueWr_Addr_reg[3]/NET0131  & n5325 ;
  assign n5360 = ~n5148 & ~n5359 ;
  assign n5361 = \P1_DataWidth_reg[1]/NET0131  & ~n5360 ;
  assign n5363 = ~n5270 & n5359 ;
  assign n5364 = ~n5279 & ~n5359 ;
  assign n5365 = ~n5363 & ~n5364 ;
  assign n5366 = n5361 & ~n5365 ;
  assign n5353 = ~n5107 & ~n5151 ;
  assign n5354 = ~n5140 & ~n5353 ;
  assign n5355 = \P1_InstQueue_reg[10][4]/NET0131  & ~n5107 ;
  assign n5356 = ~n5151 & n5355 ;
  assign n5357 = ~n5354 & ~n5356 ;
  assign n5362 = n5357 & ~n5361 ;
  assign n5367 = n2436 & ~n5362 ;
  assign n5368 = ~n5366 & n5367 ;
  assign n5358 = n5095 & ~n5357 ;
  assign n5369 = ~n2188 & n5107 ;
  assign n5370 = ~n5355 & ~n5369 ;
  assign n5371 = n3042 & ~n5370 ;
  assign n5372 = \P1_InstQueue_reg[10][4]/NET0131  & ~n5291 ;
  assign n5373 = ~n5371 & ~n5372 ;
  assign n5374 = ~n5358 & n5373 ;
  assign n5375 = ~n5368 & n5374 ;
  assign n5384 = \P1_DataWidth_reg[1]/NET0131  & ~n5353 ;
  assign n5386 = n5151 & ~n5270 ;
  assign n5387 = ~n5151 & ~n5279 ;
  assign n5388 = ~n5386 & ~n5387 ;
  assign n5389 = n5384 & ~n5388 ;
  assign n5376 = \P1_InstQueueWr_Addr_reg[2]/NET0131  & n5146 ;
  assign n5377 = \P1_InstQueueWr_Addr_reg[3]/NET0131  & n5376 ;
  assign n5378 = ~n5104 & ~n5377 ;
  assign n5379 = ~n5140 & ~n5378 ;
  assign n5380 = \P1_InstQueue_reg[12][4]/NET0131  & ~n5377 ;
  assign n5381 = ~n5104 & n5380 ;
  assign n5382 = ~n5379 & ~n5381 ;
  assign n5385 = n5382 & ~n5384 ;
  assign n5390 = n2436 & ~n5385 ;
  assign n5391 = ~n5389 & n5390 ;
  assign n5383 = n5095 & ~n5382 ;
  assign n5392 = ~n2188 & n5377 ;
  assign n5393 = ~n5380 & ~n5392 ;
  assign n5394 = n3042 & ~n5393 ;
  assign n5395 = \P1_InstQueue_reg[12][4]/NET0131  & ~n5291 ;
  assign n5396 = ~n5394 & ~n5395 ;
  assign n5397 = ~n5383 & n5396 ;
  assign n5398 = ~n5391 & n5397 ;
  assign n5405 = \P1_DataWidth_reg[1]/NET0131  & ~n5108 ;
  assign n5407 = n5107 & ~n5270 ;
  assign n5408 = ~n5107 & ~n5279 ;
  assign n5409 = ~n5407 & ~n5408 ;
  assign n5410 = n5405 & ~n5409 ;
  assign n5399 = ~n5334 & ~n5377 ;
  assign n5400 = ~n5140 & ~n5399 ;
  assign n5401 = \P1_InstQueue_reg[13][4]/NET0131  & ~n5334 ;
  assign n5402 = ~n5377 & n5401 ;
  assign n5403 = ~n5400 & ~n5402 ;
  assign n5406 = n5403 & ~n5405 ;
  assign n5411 = n2436 & ~n5406 ;
  assign n5412 = ~n5410 & n5411 ;
  assign n5404 = n5095 & ~n5403 ;
  assign n5413 = ~n2188 & n5334 ;
  assign n5414 = ~n5401 & ~n5413 ;
  assign n5415 = n3042 & ~n5414 ;
  assign n5416 = \P1_InstQueue_reg[13][4]/NET0131  & ~n5291 ;
  assign n5417 = ~n5415 & ~n5416 ;
  assign n5418 = ~n5404 & n5417 ;
  assign n5419 = ~n5412 & n5418 ;
  assign n5425 = \P1_DataWidth_reg[1]/NET0131  & ~n5378 ;
  assign n5427 = n5104 & ~n5270 ;
  assign n5428 = ~n5104 & ~n5279 ;
  assign n5429 = ~n5427 & ~n5428 ;
  assign n5430 = n5425 & ~n5429 ;
  assign n5420 = ~n5140 & ~n5337 ;
  assign n5421 = \P1_InstQueue_reg[14][4]/NET0131  & ~n5336 ;
  assign n5422 = ~n5334 & n5421 ;
  assign n5423 = ~n5420 & ~n5422 ;
  assign n5426 = n5423 & ~n5425 ;
  assign n5431 = n2436 & ~n5426 ;
  assign n5432 = ~n5430 & n5431 ;
  assign n5424 = n5095 & ~n5423 ;
  assign n5433 = ~n2188 & n5336 ;
  assign n5434 = ~n5421 & ~n5433 ;
  assign n5435 = n3042 & ~n5434 ;
  assign n5436 = \P1_InstQueue_reg[14][4]/NET0131  & ~n5291 ;
  assign n5437 = ~n5435 & ~n5436 ;
  assign n5438 = ~n5424 & n5437 ;
  assign n5439 = ~n5432 & n5438 ;
  assign n5446 = \P1_DataWidth_reg[1]/NET0131  & ~n5399 ;
  assign n5448 = ~n5270 & n5377 ;
  assign n5449 = ~n5279 & ~n5377 ;
  assign n5450 = ~n5448 & ~n5449 ;
  assign n5451 = n5446 & ~n5450 ;
  assign n5440 = ~n5326 & ~n5336 ;
  assign n5441 = ~n5140 & ~n5440 ;
  assign n5442 = \P1_InstQueue_reg[15][4]/NET0131  & ~n5326 ;
  assign n5443 = ~n5336 & n5442 ;
  assign n5444 = ~n5441 & ~n5443 ;
  assign n5447 = n5444 & ~n5446 ;
  assign n5452 = n2436 & ~n5447 ;
  assign n5453 = ~n5451 & n5452 ;
  assign n5445 = n5095 & ~n5444 ;
  assign n5454 = ~n2188 & n5326 ;
  assign n5455 = ~n5442 & ~n5454 ;
  assign n5456 = n3042 & ~n5455 ;
  assign n5457 = \P1_InstQueue_reg[15][4]/NET0131  & ~n5291 ;
  assign n5458 = ~n5456 & ~n5457 ;
  assign n5459 = ~n5445 & n5458 ;
  assign n5460 = ~n5453 & n5459 ;
  assign n5468 = \P1_DataWidth_reg[1]/NET0131  & ~n5440 ;
  assign n5470 = ~n5270 & n5336 ;
  assign n5471 = ~n5279 & ~n5336 ;
  assign n5472 = ~n5470 & ~n5471 ;
  assign n5473 = n5468 & ~n5472 ;
  assign n5461 = ~\P1_InstQueueWr_Addr_reg[3]/NET0131  & n5150 ;
  assign n5462 = ~n5324 & ~n5461 ;
  assign n5463 = ~n5140 & ~n5462 ;
  assign n5464 = \P1_InstQueue_reg[1][4]/NET0131  & ~n5461 ;
  assign n5465 = ~n5324 & n5464 ;
  assign n5466 = ~n5463 & ~n5465 ;
  assign n5469 = n5466 & ~n5468 ;
  assign n5474 = n2436 & ~n5469 ;
  assign n5475 = ~n5473 & n5474 ;
  assign n5467 = n5095 & ~n5466 ;
  assign n5476 = ~n2188 & n5461 ;
  assign n5477 = ~n5464 & ~n5476 ;
  assign n5478 = n3042 & ~n5477 ;
  assign n5479 = \P1_InstQueue_reg[1][4]/NET0131  & ~n5291 ;
  assign n5480 = ~n5478 & ~n5479 ;
  assign n5481 = ~n5467 & n5480 ;
  assign n5482 = ~n5475 & n5481 ;
  assign n5491 = \P1_DataWidth_reg[1]/NET0131  & ~n5462 ;
  assign n5493 = ~n5270 & n5324 ;
  assign n5494 = ~n5279 & ~n5324 ;
  assign n5495 = ~n5493 & ~n5494 ;
  assign n5496 = n5491 & ~n5495 ;
  assign n5483 = ~\P1_InstQueueWr_Addr_reg[3]/NET0131  & n5103 ;
  assign n5484 = ~\P1_InstQueueWr_Addr_reg[3]/NET0131  & n5106 ;
  assign n5485 = ~n5483 & ~n5484 ;
  assign n5486 = ~n5140 & ~n5485 ;
  assign n5487 = \P1_InstQueue_reg[3][4]/NET0131  & ~n5483 ;
  assign n5488 = ~n5484 & n5487 ;
  assign n5489 = ~n5486 & ~n5488 ;
  assign n5492 = n5489 & ~n5491 ;
  assign n5497 = n2436 & ~n5492 ;
  assign n5498 = ~n5496 & n5497 ;
  assign n5490 = n5095 & ~n5489 ;
  assign n5499 = ~n2188 & n5483 ;
  assign n5500 = ~n5487 & ~n5499 ;
  assign n5501 = n3042 & ~n5500 ;
  assign n5502 = \P1_InstQueue_reg[3][4]/NET0131  & ~n5291 ;
  assign n5503 = ~n5501 & ~n5502 ;
  assign n5504 = ~n5490 & n5503 ;
  assign n5505 = ~n5498 & n5504 ;
  assign n5512 = \P1_DataWidth_reg[1]/NET0131  & ~n5327 ;
  assign n5514 = ~n5270 & n5326 ;
  assign n5515 = ~n5279 & ~n5326 ;
  assign n5516 = ~n5514 & ~n5515 ;
  assign n5517 = n5512 & ~n5516 ;
  assign n5506 = ~n5461 & ~n5484 ;
  assign n5507 = ~n5140 & ~n5506 ;
  assign n5508 = \P1_InstQueue_reg[2][4]/NET0131  & ~n5484 ;
  assign n5509 = ~n5461 & n5508 ;
  assign n5510 = ~n5507 & ~n5509 ;
  assign n5513 = n5510 & ~n5512 ;
  assign n5518 = n2436 & ~n5513 ;
  assign n5519 = ~n5517 & n5518 ;
  assign n5511 = n5095 & ~n5510 ;
  assign n5520 = ~n2188 & n5484 ;
  assign n5521 = ~n5508 & ~n5520 ;
  assign n5522 = n3042 & ~n5521 ;
  assign n5523 = \P1_InstQueue_reg[2][4]/NET0131  & ~n5291 ;
  assign n5524 = ~n5522 & ~n5523 ;
  assign n5525 = ~n5511 & n5524 ;
  assign n5526 = ~n5519 & n5525 ;
  assign n5534 = \P1_DataWidth_reg[1]/NET0131  & ~n5506 ;
  assign n5536 = ~n5270 & n5461 ;
  assign n5537 = ~n5279 & ~n5461 ;
  assign n5538 = ~n5536 & ~n5537 ;
  assign n5539 = n5534 & ~n5538 ;
  assign n5527 = ~\P1_InstQueueWr_Addr_reg[3]/NET0131  & n5376 ;
  assign n5528 = ~n5483 & ~n5527 ;
  assign n5529 = ~n5140 & ~n5528 ;
  assign n5530 = \P1_InstQueue_reg[4][4]/NET0131  & ~n5527 ;
  assign n5531 = ~n5483 & n5530 ;
  assign n5532 = ~n5529 & ~n5531 ;
  assign n5535 = n5532 & ~n5534 ;
  assign n5540 = n2436 & ~n5535 ;
  assign n5541 = ~n5539 & n5540 ;
  assign n5533 = n5095 & ~n5532 ;
  assign n5542 = ~n2188 & n5527 ;
  assign n5543 = ~n5530 & ~n5542 ;
  assign n5544 = n3042 & ~n5543 ;
  assign n5545 = \P1_InstQueue_reg[4][4]/NET0131  & ~n5291 ;
  assign n5546 = ~n5544 & ~n5545 ;
  assign n5547 = ~n5533 & n5546 ;
  assign n5548 = ~n5541 & n5547 ;
  assign n5556 = \P1_DataWidth_reg[1]/NET0131  & ~n5485 ;
  assign n5558 = ~n5270 & n5484 ;
  assign n5559 = ~n5279 & ~n5484 ;
  assign n5560 = ~n5558 & ~n5559 ;
  assign n5561 = n5556 & ~n5560 ;
  assign n5549 = ~\P1_InstQueueWr_Addr_reg[3]/NET0131  & n5333 ;
  assign n5550 = ~n5527 & ~n5549 ;
  assign n5551 = ~n5140 & ~n5550 ;
  assign n5552 = \P1_InstQueue_reg[5][4]/NET0131  & ~n5549 ;
  assign n5553 = ~n5527 & n5552 ;
  assign n5554 = ~n5551 & ~n5553 ;
  assign n5557 = n5554 & ~n5556 ;
  assign n5562 = n2436 & ~n5557 ;
  assign n5563 = ~n5561 & n5562 ;
  assign n5555 = n5095 & ~n5554 ;
  assign n5564 = ~n2188 & n5549 ;
  assign n5565 = ~n5552 & ~n5564 ;
  assign n5566 = n3042 & ~n5565 ;
  assign n5567 = \P1_InstQueue_reg[5][4]/NET0131  & ~n5291 ;
  assign n5568 = ~n5566 & ~n5567 ;
  assign n5569 = ~n5555 & n5568 ;
  assign n5570 = ~n5563 & n5569 ;
  assign n5578 = \P1_DataWidth_reg[1]/NET0131  & ~n5528 ;
  assign n5580 = ~n5270 & n5483 ;
  assign n5581 = ~n5279 & ~n5483 ;
  assign n5582 = ~n5580 & ~n5581 ;
  assign n5583 = n5578 & ~n5582 ;
  assign n5571 = ~\P1_InstQueueWr_Addr_reg[3]/NET0131  & n5335 ;
  assign n5572 = ~n5549 & ~n5571 ;
  assign n5573 = ~n5140 & ~n5572 ;
  assign n5574 = \P1_InstQueue_reg[6][4]/NET0131  & ~n5571 ;
  assign n5575 = ~n5549 & n5574 ;
  assign n5576 = ~n5573 & ~n5575 ;
  assign n5579 = n5576 & ~n5578 ;
  assign n5584 = n2436 & ~n5579 ;
  assign n5585 = ~n5583 & n5584 ;
  assign n5577 = n5095 & ~n5576 ;
  assign n5586 = ~n2188 & n5571 ;
  assign n5587 = ~n5574 & ~n5586 ;
  assign n5588 = n3042 & ~n5587 ;
  assign n5589 = \P1_InstQueue_reg[6][4]/NET0131  & ~n5291 ;
  assign n5590 = ~n5588 & ~n5589 ;
  assign n5591 = ~n5577 & n5590 ;
  assign n5592 = ~n5585 & n5591 ;
  assign n5599 = \P1_DataWidth_reg[1]/NET0131  & ~n5550 ;
  assign n5601 = ~n5270 & n5527 ;
  assign n5602 = ~n5279 & ~n5527 ;
  assign n5603 = ~n5601 & ~n5602 ;
  assign n5604 = n5599 & ~n5603 ;
  assign n5593 = ~n5359 & ~n5571 ;
  assign n5594 = ~n5140 & ~n5593 ;
  assign n5595 = \P1_InstQueue_reg[7][4]/NET0131  & ~n5359 ;
  assign n5596 = ~n5571 & n5595 ;
  assign n5597 = ~n5594 & ~n5596 ;
  assign n5600 = n5597 & ~n5599 ;
  assign n5605 = n2436 & ~n5600 ;
  assign n5606 = ~n5604 & n5605 ;
  assign n5598 = n5095 & ~n5597 ;
  assign n5607 = ~n2188 & n5359 ;
  assign n5608 = ~n5595 & ~n5607 ;
  assign n5609 = n3042 & ~n5608 ;
  assign n5610 = \P1_InstQueue_reg[7][4]/NET0131  & ~n5291 ;
  assign n5611 = ~n5609 & ~n5610 ;
  assign n5612 = ~n5598 & n5611 ;
  assign n5613 = ~n5606 & n5612 ;
  assign n5619 = \P1_DataWidth_reg[1]/NET0131  & ~n5572 ;
  assign n5621 = ~n5270 & n5549 ;
  assign n5622 = ~n5279 & ~n5549 ;
  assign n5623 = ~n5621 & ~n5622 ;
  assign n5624 = n5619 & ~n5623 ;
  assign n5614 = ~n5140 & ~n5360 ;
  assign n5615 = \P1_InstQueue_reg[8][4]/NET0131  & ~n5148 ;
  assign n5616 = ~n5359 & n5615 ;
  assign n5617 = ~n5614 & ~n5616 ;
  assign n5620 = n5617 & ~n5619 ;
  assign n5625 = n2436 & ~n5620 ;
  assign n5626 = ~n5624 & n5625 ;
  assign n5618 = n5095 & ~n5617 ;
  assign n5627 = ~n2188 & n5148 ;
  assign n5628 = ~n5615 & ~n5627 ;
  assign n5629 = n3042 & ~n5628 ;
  assign n5630 = \P1_InstQueue_reg[8][4]/NET0131  & ~n5291 ;
  assign n5631 = ~n5629 & ~n5630 ;
  assign n5632 = ~n5618 & n5631 ;
  assign n5633 = ~n5626 & n5632 ;
  assign n5639 = \P1_DataWidth_reg[1]/NET0131  & ~n5593 ;
  assign n5641 = ~n5270 & n5571 ;
  assign n5642 = ~n5279 & ~n5571 ;
  assign n5643 = ~n5641 & ~n5642 ;
  assign n5644 = n5639 & ~n5643 ;
  assign n5634 = ~n5140 & ~n5152 ;
  assign n5635 = \P1_InstQueue_reg[9][4]/NET0131  & ~n5151 ;
  assign n5636 = ~n5148 & n5635 ;
  assign n5637 = ~n5634 & ~n5636 ;
  assign n5640 = n5637 & ~n5639 ;
  assign n5645 = n2436 & ~n5640 ;
  assign n5646 = ~n5644 & n5645 ;
  assign n5638 = n5095 & ~n5637 ;
  assign n5647 = ~n2188 & n5151 ;
  assign n5648 = ~n5635 & ~n5647 ;
  assign n5649 = n3042 & ~n5648 ;
  assign n5650 = \P1_InstQueue_reg[9][4]/NET0131  & ~n5291 ;
  assign n5651 = ~n5649 & ~n5650 ;
  assign n5652 = ~n5638 & n5651 ;
  assign n5653 = ~n5646 & n5652 ;
  assign n5659 = n3162 & ~n5306 ;
  assign n5660 = n3165 & ~n5310 ;
  assign n5661 = ~n5659 & ~n5660 ;
  assign n5662 = \P2_DataWidth_reg[1]/NET0131  & ~n5661 ;
  assign n5654 = ~n3155 & ~n5298 ;
  assign n5655 = \P2_InstQueue_reg[0][3]/NET0131  & ~n3152 ;
  assign n5656 = ~n3154 & n5655 ;
  assign n5657 = ~n5654 & ~n5656 ;
  assign n5663 = ~n3170 & ~n5657 ;
  assign n5664 = ~n5662 & ~n5663 ;
  assign n5665 = n1931 & ~n5664 ;
  assign n5658 = n3087 & ~n5657 ;
  assign n5666 = ~n1529 & n3152 ;
  assign n5667 = ~n5655 & ~n5666 ;
  assign n5668 = n3040 & ~n5667 ;
  assign n5669 = \P2_InstQueue_reg[0][3]/NET0131  & ~n3118 ;
  assign n5670 = ~n5668 & ~n5669 ;
  assign n5671 = ~n5658 & n5670 ;
  assign n5672 = ~n5665 & n5671 ;
  assign n5678 = n3091 & ~n5310 ;
  assign n5679 = n3198 & ~n5306 ;
  assign n5680 = ~n5678 & ~n5679 ;
  assign n5681 = \P2_DataWidth_reg[1]/NET0131  & ~n5680 ;
  assign n5673 = ~n3202 & ~n5298 ;
  assign n5674 = \P2_InstQueue_reg[10][3]/NET0131  & ~n3046 ;
  assign n5675 = ~n3098 & n5674 ;
  assign n5676 = ~n5673 & ~n5675 ;
  assign n5682 = ~n3200 & ~n5676 ;
  assign n5683 = ~n5681 & ~n5682 ;
  assign n5684 = n1931 & ~n5683 ;
  assign n5677 = n3087 & ~n5676 ;
  assign n5685 = ~n1529 & n3046 ;
  assign n5686 = ~n5674 & ~n5685 ;
  assign n5687 = n3040 & ~n5686 ;
  assign n5688 = \P2_InstQueue_reg[10][3]/NET0131  & ~n3118 ;
  assign n5689 = ~n5687 & ~n5688 ;
  assign n5690 = ~n5677 & n5689 ;
  assign n5691 = ~n5684 & n5690 ;
  assign n5697 = n3098 & ~n5306 ;
  assign n5698 = n3046 & ~n5310 ;
  assign n5699 = ~n5697 & ~n5698 ;
  assign n5700 = \P2_DataWidth_reg[1]/NET0131  & ~n5699 ;
  assign n5692 = ~n3238 & ~n5298 ;
  assign n5693 = \P2_InstQueue_reg[12][3]/NET0131  & ~n3237 ;
  assign n5694 = ~n3049 & n5693 ;
  assign n5695 = ~n5692 & ~n5694 ;
  assign n5701 = ~n3248 & ~n5695 ;
  assign n5702 = ~n5700 & ~n5701 ;
  assign n5703 = n1931 & ~n5702 ;
  assign n5696 = n3087 & ~n5695 ;
  assign n5704 = ~n1529 & n3237 ;
  assign n5705 = ~n5693 & ~n5704 ;
  assign n5706 = n3040 & ~n5705 ;
  assign n5707 = \P2_InstQueue_reg[12][3]/NET0131  & ~n3118 ;
  assign n5708 = ~n5706 & ~n5707 ;
  assign n5709 = ~n5696 & n5708 ;
  assign n5710 = ~n5703 & n5709 ;
  assign n5716 = n3046 & ~n5306 ;
  assign n5717 = n3049 & ~n5310 ;
  assign n5718 = ~n5716 & ~n5717 ;
  assign n5719 = \P2_DataWidth_reg[1]/NET0131  & ~n5718 ;
  assign n5711 = ~n3275 & ~n5298 ;
  assign n5712 = \P2_InstQueue_reg[13][3]/NET0131  & ~n3162 ;
  assign n5713 = ~n3237 & n5712 ;
  assign n5714 = ~n5711 & ~n5713 ;
  assign n5720 = ~n3285 & ~n5714 ;
  assign n5721 = ~n5719 & ~n5720 ;
  assign n5722 = n1931 & ~n5721 ;
  assign n5715 = n3087 & ~n5714 ;
  assign n5723 = ~n1529 & n3162 ;
  assign n5724 = ~n5712 & ~n5723 ;
  assign n5725 = n3040 & ~n5724 ;
  assign n5726 = \P2_InstQueue_reg[13][3]/NET0131  & ~n3118 ;
  assign n5727 = ~n5725 & ~n5726 ;
  assign n5728 = ~n5715 & n5727 ;
  assign n5729 = ~n5722 & n5728 ;
  assign n5735 = n3049 & ~n5306 ;
  assign n5736 = n3237 & ~n5310 ;
  assign n5737 = ~n5735 & ~n5736 ;
  assign n5738 = \P2_DataWidth_reg[1]/NET0131  & ~n5737 ;
  assign n5730 = ~n3169 & ~n5298 ;
  assign n5731 = \P2_InstQueue_reg[14][3]/NET0131  & ~n3165 ;
  assign n5732 = ~n3162 & n5731 ;
  assign n5733 = ~n5730 & ~n5732 ;
  assign n5739 = ~n3321 & ~n5733 ;
  assign n5740 = ~n5738 & ~n5739 ;
  assign n5741 = n1931 & ~n5740 ;
  assign n5734 = n3087 & ~n5733 ;
  assign n5742 = ~n1529 & n3165 ;
  assign n5743 = ~n5731 & ~n5742 ;
  assign n5744 = n3040 & ~n5743 ;
  assign n5745 = \P2_InstQueue_reg[14][3]/NET0131  & ~n3118 ;
  assign n5746 = ~n5744 & ~n5745 ;
  assign n5747 = ~n5734 & n5746 ;
  assign n5748 = ~n5741 & n5747 ;
  assign n5754 = n3237 & ~n5306 ;
  assign n5755 = n3162 & ~n5310 ;
  assign n5756 = ~n5754 & ~n5755 ;
  assign n5757 = \P2_DataWidth_reg[1]/NET0131  & ~n5756 ;
  assign n5749 = ~n3348 & ~n5298 ;
  assign n5750 = \P2_InstQueue_reg[15][3]/NET0131  & ~n3154 ;
  assign n5751 = ~n3165 & n5750 ;
  assign n5752 = ~n5749 & ~n5751 ;
  assign n5758 = ~n3358 & ~n5752 ;
  assign n5759 = ~n5757 & ~n5758 ;
  assign n5760 = n1931 & ~n5759 ;
  assign n5753 = n3087 & ~n5752 ;
  assign n5761 = ~n1529 & n3154 ;
  assign n5762 = ~n5750 & ~n5761 ;
  assign n5763 = n3040 & ~n5762 ;
  assign n5764 = \P2_InstQueue_reg[15][3]/NET0131  & ~n3118 ;
  assign n5765 = ~n5763 & ~n5764 ;
  assign n5766 = ~n5753 & n5765 ;
  assign n5767 = ~n5760 & n5766 ;
  assign n5773 = n3165 & ~n5306 ;
  assign n5774 = n3154 & ~n5310 ;
  assign n5775 = ~n5773 & ~n5774 ;
  assign n5776 = \P2_DataWidth_reg[1]/NET0131  & ~n5775 ;
  assign n5768 = ~n3389 & ~n5298 ;
  assign n5769 = \P2_InstQueue_reg[1][3]/NET0131  & ~n3388 ;
  assign n5770 = ~n3152 & n5769 ;
  assign n5771 = ~n5768 & ~n5770 ;
  assign n5777 = ~n3386 & ~n5771 ;
  assign n5778 = ~n5776 & ~n5777 ;
  assign n5779 = n1931 & ~n5778 ;
  assign n5772 = n3087 & ~n5771 ;
  assign n5780 = ~n1529 & n3388 ;
  assign n5781 = ~n5769 & ~n5780 ;
  assign n5782 = n3040 & ~n5781 ;
  assign n5783 = \P2_InstQueue_reg[1][3]/NET0131  & ~n3118 ;
  assign n5784 = ~n5782 & ~n5783 ;
  assign n5785 = ~n5772 & n5784 ;
  assign n5786 = ~n5779 & n5785 ;
  assign n5792 = n3152 & ~n5310 ;
  assign n5793 = n3154 & ~n5306 ;
  assign n5794 = ~n5792 & ~n5793 ;
  assign n5795 = \P2_DataWidth_reg[1]/NET0131  & ~n5794 ;
  assign n5787 = ~n3424 & ~n5298 ;
  assign n5788 = \P2_InstQueue_reg[2][3]/NET0131  & ~n3423 ;
  assign n5789 = ~n3388 & n5788 ;
  assign n5790 = ~n5787 & ~n5789 ;
  assign n5796 = ~n3434 & ~n5790 ;
  assign n5797 = ~n5795 & ~n5796 ;
  assign n5798 = n1931 & ~n5797 ;
  assign n5791 = n3087 & ~n5790 ;
  assign n5799 = ~n1529 & n3423 ;
  assign n5800 = ~n5788 & ~n5799 ;
  assign n5801 = n3040 & ~n5800 ;
  assign n5802 = \P2_InstQueue_reg[2][3]/NET0131  & ~n3118 ;
  assign n5803 = ~n5801 & ~n5802 ;
  assign n5804 = ~n5791 & n5803 ;
  assign n5805 = ~n5798 & n5804 ;
  assign n5811 = n3152 & ~n5306 ;
  assign n5812 = n3388 & ~n5310 ;
  assign n5813 = ~n5811 & ~n5812 ;
  assign n5814 = \P2_DataWidth_reg[1]/NET0131  & ~n5813 ;
  assign n5806 = ~n3462 & ~n5298 ;
  assign n5807 = \P2_InstQueue_reg[3][3]/NET0131  & ~n3461 ;
  assign n5808 = ~n3423 & n5807 ;
  assign n5809 = ~n5806 & ~n5808 ;
  assign n5815 = ~n3472 & ~n5809 ;
  assign n5816 = ~n5814 & ~n5815 ;
  assign n5817 = n1931 & ~n5816 ;
  assign n5810 = n3087 & ~n5809 ;
  assign n5818 = ~n1529 & n3461 ;
  assign n5819 = ~n5807 & ~n5818 ;
  assign n5820 = n3040 & ~n5819 ;
  assign n5821 = \P2_InstQueue_reg[3][3]/NET0131  & ~n3118 ;
  assign n5822 = ~n5820 & ~n5821 ;
  assign n5823 = ~n5810 & n5822 ;
  assign n5824 = ~n5817 & n5823 ;
  assign n5830 = n3388 & ~n5306 ;
  assign n5831 = n3423 & ~n5310 ;
  assign n5832 = ~n5830 & ~n5831 ;
  assign n5833 = \P2_DataWidth_reg[1]/NET0131  & ~n5832 ;
  assign n5825 = ~n3500 & ~n5298 ;
  assign n5826 = \P2_InstQueue_reg[4][3]/NET0131  & ~n3499 ;
  assign n5827 = ~n3461 & n5826 ;
  assign n5828 = ~n5825 & ~n5827 ;
  assign n5834 = ~n3510 & ~n5828 ;
  assign n5835 = ~n5833 & ~n5834 ;
  assign n5836 = n1931 & ~n5835 ;
  assign n5829 = n3087 & ~n5828 ;
  assign n5837 = ~n1529 & n3499 ;
  assign n5838 = ~n5826 & ~n5837 ;
  assign n5839 = n3040 & ~n5838 ;
  assign n5840 = \P2_InstQueue_reg[4][3]/NET0131  & ~n3118 ;
  assign n5841 = ~n5839 & ~n5840 ;
  assign n5842 = ~n5829 & n5841 ;
  assign n5843 = ~n5836 & n5842 ;
  assign n5849 = n3423 & ~n5306 ;
  assign n5850 = n3461 & ~n5310 ;
  assign n5851 = ~n5849 & ~n5850 ;
  assign n5852 = \P2_DataWidth_reg[1]/NET0131  & ~n5851 ;
  assign n5844 = ~n3538 & ~n5298 ;
  assign n5845 = \P2_InstQueue_reg[5][3]/NET0131  & ~n3537 ;
  assign n5846 = ~n3499 & n5845 ;
  assign n5847 = ~n5844 & ~n5846 ;
  assign n5853 = ~n3548 & ~n5847 ;
  assign n5854 = ~n5852 & ~n5853 ;
  assign n5855 = n1931 & ~n5854 ;
  assign n5848 = n3087 & ~n5847 ;
  assign n5856 = ~n1529 & n3537 ;
  assign n5857 = ~n5845 & ~n5856 ;
  assign n5858 = n3040 & ~n5857 ;
  assign n5859 = \P2_InstQueue_reg[5][3]/NET0131  & ~n3118 ;
  assign n5860 = ~n5858 & ~n5859 ;
  assign n5861 = ~n5848 & n5860 ;
  assign n5862 = ~n5855 & n5861 ;
  assign n5868 = n3461 & ~n5306 ;
  assign n5869 = n3499 & ~n5310 ;
  assign n5870 = ~n5868 & ~n5869 ;
  assign n5871 = \P2_DataWidth_reg[1]/NET0131  & ~n5870 ;
  assign n5863 = ~n3576 & ~n5298 ;
  assign n5864 = \P2_InstQueue_reg[6][3]/NET0131  & ~n3575 ;
  assign n5865 = ~n3537 & n5864 ;
  assign n5866 = ~n5863 & ~n5865 ;
  assign n5872 = ~n3586 & ~n5866 ;
  assign n5873 = ~n5871 & ~n5872 ;
  assign n5874 = n1931 & ~n5873 ;
  assign n5867 = n3087 & ~n5866 ;
  assign n5875 = ~n1529 & n3575 ;
  assign n5876 = ~n5864 & ~n5875 ;
  assign n5877 = n3040 & ~n5876 ;
  assign n5878 = \P2_InstQueue_reg[6][3]/NET0131  & ~n3118 ;
  assign n5879 = ~n5877 & ~n5878 ;
  assign n5880 = ~n5867 & n5879 ;
  assign n5881 = ~n5874 & n5880 ;
  assign n5887 = n3499 & ~n5306 ;
  assign n5888 = n3537 & ~n5310 ;
  assign n5889 = ~n5887 & ~n5888 ;
  assign n5890 = \P2_DataWidth_reg[1]/NET0131  & ~n5889 ;
  assign n5882 = ~n3613 & ~n5298 ;
  assign n5883 = \P2_InstQueue_reg[7][3]/NET0131  & ~n3198 ;
  assign n5884 = ~n3575 & n5883 ;
  assign n5885 = ~n5882 & ~n5884 ;
  assign n5891 = ~n3623 & ~n5885 ;
  assign n5892 = ~n5890 & ~n5891 ;
  assign n5893 = n1931 & ~n5892 ;
  assign n5886 = n3087 & ~n5885 ;
  assign n5894 = ~n1529 & n3198 ;
  assign n5895 = ~n5883 & ~n5894 ;
  assign n5896 = n3040 & ~n5895 ;
  assign n5897 = \P2_InstQueue_reg[7][3]/NET0131  & ~n3118 ;
  assign n5898 = ~n5896 & ~n5897 ;
  assign n5899 = ~n5886 & n5898 ;
  assign n5900 = ~n5893 & n5899 ;
  assign n5906 = n3537 & ~n5306 ;
  assign n5907 = n3575 & ~n5310 ;
  assign n5908 = ~n5906 & ~n5907 ;
  assign n5909 = \P2_DataWidth_reg[1]/NET0131  & ~n5908 ;
  assign n5901 = ~n3199 & ~n5298 ;
  assign n5902 = \P2_InstQueue_reg[8][3]/NET0131  & ~n3091 ;
  assign n5903 = ~n3198 & n5902 ;
  assign n5904 = ~n5901 & ~n5903 ;
  assign n5910 = ~n3659 & ~n5904 ;
  assign n5911 = ~n5909 & ~n5910 ;
  assign n5912 = n1931 & ~n5911 ;
  assign n5905 = n3087 & ~n5904 ;
  assign n5913 = ~n1529 & n3091 ;
  assign n5914 = ~n5902 & ~n5913 ;
  assign n5915 = n3040 & ~n5914 ;
  assign n5916 = \P2_InstQueue_reg[8][3]/NET0131  & ~n3118 ;
  assign n5917 = ~n5915 & ~n5916 ;
  assign n5918 = ~n5905 & n5917 ;
  assign n5919 = ~n5912 & n5918 ;
  assign n5925 = n3575 & ~n5306 ;
  assign n5926 = n3198 & ~n5310 ;
  assign n5927 = ~n5925 & ~n5926 ;
  assign n5928 = \P2_DataWidth_reg[1]/NET0131  & ~n5927 ;
  assign n5920 = ~n3105 & ~n5298 ;
  assign n5921 = \P2_InstQueue_reg[9][3]/NET0131  & ~n3098 ;
  assign n5922 = ~n3091 & n5921 ;
  assign n5923 = ~n5920 & ~n5922 ;
  assign n5929 = ~n3695 & ~n5923 ;
  assign n5930 = ~n5928 & ~n5929 ;
  assign n5931 = n1931 & ~n5930 ;
  assign n5924 = n3087 & ~n5923 ;
  assign n5932 = ~n1529 & n3098 ;
  assign n5933 = ~n5921 & ~n5932 ;
  assign n5934 = n3040 & ~n5933 ;
  assign n5935 = \P2_InstQueue_reg[9][3]/NET0131  & ~n3118 ;
  assign n5936 = ~n5934 & ~n5935 ;
  assign n5937 = ~n5924 & n5936 ;
  assign n5938 = ~n5931 & n5937 ;
  assign n5939 = \P1_InstAddrPointer_reg[29]/NET0131  & n2375 ;
  assign n5964 = \P1_InstAddrPointer_reg[28]/NET0131  & n4490 ;
  assign n5965 = ~\P1_InstAddrPointer_reg[29]/NET0131  & ~n5964 ;
  assign n5966 = ~n4799 & ~n5965 ;
  assign n5967 = ~\P1_InstAddrPointer_reg[17]/NET0131  & ~n4468 ;
  assign n5968 = ~n4773 & ~n5967 ;
  assign n5969 = \P1_InstAddrPointer_reg[10]/NET0131  & n4499 ;
  assign n5970 = n4781 & n5969 ;
  assign n5971 = n4467 & n4788 ;
  assign n5972 = n5970 & n5971 ;
  assign n5973 = n4765 & n5972 ;
  assign n5974 = n5968 & n5973 ;
  assign n5975 = n4778 & n5974 ;
  assign n5976 = \P1_InstAddrPointer_reg[22]/NET0131  & n4769 ;
  assign n5977 = n4494 & n5976 ;
  assign n5978 = n5975 & n5977 ;
  assign n5980 = ~n5966 & n5978 ;
  assign n5979 = n5966 & ~n5978 ;
  assign n5981 = n4453 & ~n5979 ;
  assign n5982 = ~n5980 & n5981 ;
  assign n5946 = ~n4844 & ~n4854 ;
  assign n5947 = ~n4838 & n4851 ;
  assign n5948 = ~n5946 & n5947 ;
  assign n5949 = ~n4838 & n4853 ;
  assign n5950 = ~n4859 & ~n5949 ;
  assign n5951 = ~n5948 & n5950 ;
  assign n5952 = n4835 & ~n5951 ;
  assign n5942 = ~n4864 & ~n4869 ;
  assign n5943 = ~n4833 & n4860 ;
  assign n5944 = ~n4865 & ~n5943 ;
  assign n5945 = ~n4827 & ~n5944 ;
  assign n5953 = n5942 & ~n5945 ;
  assign n5954 = ~n5952 & n5953 ;
  assign n5940 = ~n4824 & ~n4871 ;
  assign n5941 = ~n4878 & n5940 ;
  assign n5955 = ~n4884 & n5941 ;
  assign n5956 = n5954 & n5955 ;
  assign n5957 = ~n4882 & n5956 ;
  assign n5958 = n4934 & n5957 ;
  assign n5959 = n4944 & n5958 ;
  assign n5961 = n4946 & ~n5959 ;
  assign n5960 = ~n4946 & n5959 ;
  assign n5962 = ~n4453 & ~n5960 ;
  assign n5963 = ~n5961 & n5962 ;
  assign n5983 = ~n2375 & ~n5963 ;
  assign n5984 = ~n5982 & n5983 ;
  assign n5985 = ~n5939 & ~n5984 ;
  assign n5986 = n2244 & ~n5985 ;
  assign n5987 = \P1_InstAddrPointer_reg[28]/NET0131  & n5058 ;
  assign n5988 = ~\P1_InstAddrPointer_reg[29]/NET0131  & ~n5987 ;
  assign n5989 = ~n5063 & ~n5988 ;
  assign n5990 = \P1_InstAddrPointer_reg[20]/NET0131  & n4972 ;
  assign n5991 = ~\P1_InstAddrPointer_reg[20]/NET0131  & ~n4972 ;
  assign n5992 = ~n5990 & ~n5991 ;
  assign n5993 = \P1_InstAddrPointer_reg[21]/NET0131  & n5992 ;
  assign n5994 = ~n4999 & ~n5002 ;
  assign n5995 = n4995 & ~n5994 ;
  assign n5996 = ~n5001 & ~n5008 ;
  assign n5997 = ~n5995 & n5996 ;
  assign n5998 = n4990 & ~n5997 ;
  assign n5999 = ~n5007 & ~n5015 ;
  assign n6000 = ~n5998 & n5999 ;
  assign n6001 = ~n4983 & ~n6000 ;
  assign n6002 = ~n5014 & ~n6001 ;
  assign n6003 = n4977 & ~n4980 ;
  assign n6004 = n4460 & n6003 ;
  assign n6005 = ~n6002 & n6004 ;
  assign n6006 = ~\P1_InstAddrPointer_reg[15]/NET0131  & ~n5029 ;
  assign n6007 = ~n5030 & ~n6006 ;
  assign n6008 = \P1_InstAddrPointer_reg[14]/NET0131  & n5027 ;
  assign n6009 = n6007 & n6008 ;
  assign n6010 = n6005 & n6009 ;
  assign n6011 = n4470 & n5032 ;
  assign n6012 = n6010 & n6011 ;
  assign n6013 = n5993 & n6012 ;
  assign n6014 = n5051 & n6013 ;
  assign n6015 = \P1_InstAddrPointer_reg[26]/NET0131  & n5045 ;
  assign n6016 = \P1_InstAddrPointer_reg[27]/NET0131  & n6015 ;
  assign n6017 = ~\P1_InstAddrPointer_reg[28]/NET0131  & ~n5058 ;
  assign n6018 = ~n5987 & ~n6017 ;
  assign n6019 = n6016 & n6018 ;
  assign n6020 = n6014 & n6019 ;
  assign n6022 = n5989 & n6020 ;
  assign n6021 = ~n5989 & ~n6020 ;
  assign n6023 = n2385 & ~n6021 ;
  assign n6024 = ~n6022 & n6023 ;
  assign n6030 = n2397 & n5989 ;
  assign n6025 = ~n2271 & n4946 ;
  assign n6026 = ~n2325 & n2373 ;
  assign n6027 = n2390 & n6026 ;
  assign n6028 = \P1_InstAddrPointer_reg[29]/NET0131  & ~n6027 ;
  assign n6029 = ~n2402 & n5966 ;
  assign n6031 = ~n6028 & ~n6029 ;
  assign n6032 = ~n6025 & n6031 ;
  assign n6033 = ~n6030 & n6032 ;
  assign n6034 = ~n6024 & n6033 ;
  assign n6035 = ~n5986 & n6034 ;
  assign n6036 = n2432 & ~n6035 ;
  assign n6037 = \P1_rEIP_reg[29]/NET0131  & n5092 ;
  assign n6038 = \P1_InstAddrPointer_reg[29]/NET0131  & ~n5098 ;
  assign n6039 = ~n6037 & ~n6038 ;
  assign n6040 = ~n6036 & n6039 ;
  assign n6041 = \P3_InstAddrPointer_reg[28]/NET0131  & n2896 ;
  assign n6073 = ~n3966 & n4037 ;
  assign n6074 = ~n3899 & ~n4041 ;
  assign n6075 = ~n4035 & ~n6074 ;
  assign n6076 = ~n6073 & ~n6075 ;
  assign n6077 = ~n3831 & ~n4001 ;
  assign n6078 = ~n6076 & n6077 ;
  assign n6079 = ~n3831 & n4040 ;
  assign n6080 = ~n4051 & ~n6079 ;
  assign n6081 = ~n6078 & n6080 ;
  assign n6082 = ~n3865 & ~n4070 ;
  assign n6083 = ~n6081 & n6082 ;
  assign n6084 = ~n4049 & ~n4050 ;
  assign n6085 = ~n4070 & ~n6084 ;
  assign n6086 = ~n6083 & ~n6085 ;
  assign n6070 = ~\P3_InstAddrPointer_reg[10]/NET0131  & ~n3778 ;
  assign n6071 = ~n4067 & ~n6070 ;
  assign n6072 = \P3_InstAddrPointer_reg[11]/NET0131  & n6071 ;
  assign n6087 = n4062 & n6072 ;
  assign n6088 = ~n6086 & n6087 ;
  assign n6089 = n4066 & n4082 ;
  assign n6090 = n4059 & n6089 ;
  assign n6091 = n3754 & n4080 ;
  assign n6092 = n6090 & n6091 ;
  assign n6093 = n6088 & n6092 ;
  assign n6094 = n3793 & n4104 ;
  assign n6095 = n6093 & n6094 ;
  assign n6096 = ~\P3_InstAddrPointer_reg[24]/NET0131  & ~n4102 ;
  assign n6097 = ~n4097 & ~n6096 ;
  assign n6098 = n6095 & n6097 ;
  assign n6099 = n4101 & n4112 ;
  assign n6100 = n6098 & n6099 ;
  assign n6101 = ~\P3_InstAddrPointer_reg[28]/NET0131  & ~n4110 ;
  assign n6102 = n4109 & n4115 ;
  assign n6103 = ~n6101 & ~n6102 ;
  assign n6105 = ~n6100 & n6103 ;
  assign n6104 = n6100 & ~n6103 ;
  assign n6106 = n3753 & ~n6104 ;
  assign n6107 = ~n6105 & n6106 ;
  assign n6042 = n4176 & ~n4243 ;
  assign n6043 = ~n4217 & ~n4220 ;
  assign n6044 = ~n4215 & n6043 ;
  assign n6045 = n4167 & n6044 ;
  assign n6046 = ~n4192 & n4199 ;
  assign n6047 = n4190 & ~n4198 ;
  assign n6048 = ~n4206 & ~n6047 ;
  assign n6049 = ~n6046 & n6048 ;
  assign n6050 = ~n4185 & ~n4202 ;
  assign n6051 = ~n6049 & n6050 ;
  assign n6052 = ~n4185 & n4205 ;
  assign n6053 = ~n4223 & ~n6052 ;
  assign n6054 = ~n6051 & n6053 ;
  assign n6055 = n4221 & ~n6054 ;
  assign n6056 = ~n4179 & n4222 ;
  assign n6057 = ~n4218 & ~n6056 ;
  assign n6058 = ~n6055 & n6057 ;
  assign n6059 = n6045 & n6058 ;
  assign n6060 = n6042 & n6059 ;
  assign n6061 = ~n4248 & ~n4281 ;
  assign n6062 = n4241 & n6061 ;
  assign n6063 = ~n4139 & n6062 ;
  assign n6064 = n4279 & n6063 ;
  assign n6065 = n6060 & n6064 ;
  assign n6067 = ~n4142 & n6065 ;
  assign n6066 = n4142 & ~n6065 ;
  assign n6068 = ~n3753 & ~n6066 ;
  assign n6069 = ~n6067 & n6068 ;
  assign n6108 = ~n2896 & ~n6069 ;
  assign n6109 = ~n6107 & n6108 ;
  assign n6110 = ~n6041 & ~n6109 ;
  assign n6111 = n2894 & ~n6110 ;
  assign n6112 = ~\P3_InstAddrPointer_reg[28]/NET0131  & ~n4386 ;
  assign n6113 = n4115 & n4381 ;
  assign n6114 = ~n6112 & ~n6113 ;
  assign n6115 = ~n4335 & ~n4336 ;
  assign n6116 = n4320 & ~n6115 ;
  assign n6117 = ~n4319 & n4337 ;
  assign n6118 = ~n4342 & ~n6117 ;
  assign n6119 = ~n6116 & n6118 ;
  assign n6120 = ~n4313 & ~n4346 ;
  assign n6121 = ~n6119 & n6120 ;
  assign n6122 = n4341 & ~n4346 ;
  assign n6123 = ~n4310 & ~n6122 ;
  assign n6124 = ~n6121 & n6123 ;
  assign n6125 = n4307 & ~n6124 ;
  assign n6126 = n4355 & n6125 ;
  assign n6127 = n4361 & n6126 ;
  assign n6128 = n4373 & n6127 ;
  assign n6129 = n4379 & n6128 ;
  assign n6130 = \P3_InstAddrPointer_reg[26]/NET0131  & n6129 ;
  assign n6131 = n4388 & n6130 ;
  assign n6132 = ~n6114 & ~n6131 ;
  assign n6133 = n4389 & n6130 ;
  assign n6134 = n2905 & ~n6133 ;
  assign n6135 = ~n6132 & n6134 ;
  assign n6137 = ~\P3_InstAddrPointer_reg[28]/NET0131  & ~n2847 ;
  assign n6138 = ~n2841 & ~n6137 ;
  assign n6139 = n6114 & n6138 ;
  assign n6141 = ~n2766 & ~n2862 ;
  assign n6142 = ~n2906 & ~n6141 ;
  assign n6143 = n2901 & n6142 ;
  assign n6144 = \P3_InstAddrPointer_reg[28]/NET0131  & ~n6143 ;
  assign n6136 = ~n2777 & n4142 ;
  assign n6140 = ~n2923 & n6103 ;
  assign n6145 = ~n6136 & ~n6140 ;
  assign n6146 = ~n6144 & n6145 ;
  assign n6147 = ~n6139 & n6146 ;
  assign n6148 = ~n6135 & n6147 ;
  assign n6149 = ~n6111 & n6148 ;
  assign n6150 = n2453 & ~n6149 ;
  assign n6151 = \P3_rEIP_reg[28]/NET0131  & n4412 ;
  assign n6152 = \P3_InstAddrPointer_reg[28]/NET0131  & ~n4418 ;
  assign n6153 = ~n6151 & ~n6152 ;
  assign n6154 = ~n6150 & n6153 ;
  assign n6155 = \P2_InstAddrPointer_reg[29]/NET0131  & n1897 ;
  assign n6273 = \P2_InstQueue_reg[15][2]/NET0131  & n1478 ;
  assign n6274 = \P2_InstQueue_reg[5][2]/NET0131  & n1474 ;
  assign n6287 = ~n6273 & ~n6274 ;
  assign n6275 = \P2_InstQueue_reg[2][2]/NET0131  & n1468 ;
  assign n6276 = \P2_InstQueue_reg[13][2]/NET0131  & n1466 ;
  assign n6288 = ~n6275 & ~n6276 ;
  assign n6295 = n6287 & n6288 ;
  assign n6269 = \P2_InstQueue_reg[0][2]/NET0131  & n1456 ;
  assign n6270 = \P2_InstQueue_reg[4][2]/NET0131  & n1450 ;
  assign n6285 = ~n6269 & ~n6270 ;
  assign n6271 = \P2_InstQueue_reg[9][2]/NET0131  & n1472 ;
  assign n6272 = \P2_InstQueue_reg[1][2]/NET0131  & n1464 ;
  assign n6286 = ~n6271 & ~n6272 ;
  assign n6296 = n6285 & n6286 ;
  assign n6297 = n6295 & n6296 ;
  assign n6281 = \P2_InstQueue_reg[3][2]/NET0131  & n1470 ;
  assign n6282 = \P2_InstQueue_reg[10][2]/NET0131  & n1453 ;
  assign n6291 = ~n6281 & ~n6282 ;
  assign n6283 = \P2_InstQueue_reg[11][2]/NET0131  & n1459 ;
  assign n6284 = \P2_InstQueue_reg[7][2]/NET0131  & n1476 ;
  assign n6292 = ~n6283 & ~n6284 ;
  assign n6293 = n6291 & n6292 ;
  assign n6277 = \P2_InstQueue_reg[8][2]/NET0131  & n1461 ;
  assign n6278 = \P2_InstQueue_reg[6][2]/NET0131  & n1447 ;
  assign n6289 = ~n6277 & ~n6278 ;
  assign n6279 = \P2_InstQueue_reg[14][2]/NET0131  & n1482 ;
  assign n6280 = \P2_InstQueue_reg[12][2]/NET0131  & n1480 ;
  assign n6290 = ~n6279 & ~n6280 ;
  assign n6294 = n6289 & n6290 ;
  assign n6298 = n6293 & n6294 ;
  assign n6299 = n6297 & n6298 ;
  assign n6464 = \P2_InstAddrPointer_reg[1]/NET0131  & \P2_InstAddrPointer_reg[2]/NET0131  ;
  assign n6610 = ~\P2_InstAddrPointer_reg[1]/NET0131  & ~\P2_InstAddrPointer_reg[2]/NET0131  ;
  assign n6611 = ~n6464 & ~n6610 ;
  assign n6612 = ~n6299 & n6611 ;
  assign n6307 = \P2_InstQueue_reg[5][1]/NET0131  & n1474 ;
  assign n6308 = \P2_InstQueue_reg[1][1]/NET0131  & n1464 ;
  assign n6321 = ~n6307 & ~n6308 ;
  assign n6309 = \P2_InstQueue_reg[3][1]/NET0131  & n1470 ;
  assign n6310 = \P2_InstQueue_reg[10][1]/NET0131  & n1453 ;
  assign n6322 = ~n6309 & ~n6310 ;
  assign n6329 = n6321 & n6322 ;
  assign n6303 = \P2_InstQueue_reg[15][1]/NET0131  & n1478 ;
  assign n6304 = \P2_InstQueue_reg[9][1]/NET0131  & n1472 ;
  assign n6319 = ~n6303 & ~n6304 ;
  assign n6305 = \P2_InstQueue_reg[0][1]/NET0131  & n1456 ;
  assign n6306 = \P2_InstQueue_reg[7][1]/NET0131  & n1476 ;
  assign n6320 = ~n6305 & ~n6306 ;
  assign n6330 = n6319 & n6320 ;
  assign n6331 = n6329 & n6330 ;
  assign n6315 = \P2_InstQueue_reg[2][1]/NET0131  & n1468 ;
  assign n6316 = \P2_InstQueue_reg[12][1]/NET0131  & n1480 ;
  assign n6325 = ~n6315 & ~n6316 ;
  assign n6317 = \P2_InstQueue_reg[14][1]/NET0131  & n1482 ;
  assign n6318 = \P2_InstQueue_reg[11][1]/NET0131  & n1459 ;
  assign n6326 = ~n6317 & ~n6318 ;
  assign n6327 = n6325 & n6326 ;
  assign n6311 = \P2_InstQueue_reg[13][1]/NET0131  & n1466 ;
  assign n6312 = \P2_InstQueue_reg[4][1]/NET0131  & n1450 ;
  assign n6323 = ~n6311 & ~n6312 ;
  assign n6313 = \P2_InstQueue_reg[6][1]/NET0131  & n1447 ;
  assign n6314 = \P2_InstQueue_reg[8][1]/NET0131  & n1461 ;
  assign n6324 = ~n6313 & ~n6314 ;
  assign n6328 = n6323 & n6324 ;
  assign n6332 = n6327 & n6328 ;
  assign n6333 = n6331 & n6332 ;
  assign n6337 = ~\P2_InstAddrPointer_reg[1]/NET0131  & ~n6333 ;
  assign n6613 = \P2_InstAddrPointer_reg[1]/NET0131  & n6333 ;
  assign n6342 = \P2_InstQueue_reg[14][0]/NET0131  & n1482 ;
  assign n6343 = \P2_InstQueue_reg[1][0]/NET0131  & n1464 ;
  assign n6356 = ~n6342 & ~n6343 ;
  assign n6344 = \P2_InstQueue_reg[12][0]/NET0131  & n1480 ;
  assign n6345 = \P2_InstQueue_reg[2][0]/NET0131  & n1468 ;
  assign n6357 = ~n6344 & ~n6345 ;
  assign n6364 = n6356 & n6357 ;
  assign n6338 = \P2_InstQueue_reg[6][0]/NET0131  & n1447 ;
  assign n6339 = \P2_InstQueue_reg[5][0]/NET0131  & n1474 ;
  assign n6354 = ~n6338 & ~n6339 ;
  assign n6340 = \P2_InstQueue_reg[11][0]/NET0131  & n1459 ;
  assign n6341 = \P2_InstQueue_reg[3][0]/NET0131  & n1470 ;
  assign n6355 = ~n6340 & ~n6341 ;
  assign n6365 = n6354 & n6355 ;
  assign n6366 = n6364 & n6365 ;
  assign n6350 = \P2_InstQueue_reg[7][0]/NET0131  & n1476 ;
  assign n6351 = \P2_InstQueue_reg[13][0]/NET0131  & n1466 ;
  assign n6360 = ~n6350 & ~n6351 ;
  assign n6352 = \P2_InstQueue_reg[9][0]/NET0131  & n1472 ;
  assign n6353 = \P2_InstQueue_reg[15][0]/NET0131  & n1478 ;
  assign n6361 = ~n6352 & ~n6353 ;
  assign n6362 = n6360 & n6361 ;
  assign n6346 = \P2_InstQueue_reg[0][0]/NET0131  & n1456 ;
  assign n6347 = \P2_InstQueue_reg[8][0]/NET0131  & n1461 ;
  assign n6358 = ~n6346 & ~n6347 ;
  assign n6348 = \P2_InstQueue_reg[10][0]/NET0131  & n1453 ;
  assign n6349 = \P2_InstQueue_reg[4][0]/NET0131  & n1450 ;
  assign n6359 = ~n6348 & ~n6349 ;
  assign n6363 = n6358 & n6359 ;
  assign n6367 = n6362 & n6363 ;
  assign n6368 = n6366 & n6367 ;
  assign n6614 = \P2_InstAddrPointer_reg[0]/NET0131  & ~n6368 ;
  assign n6615 = ~n6613 & n6614 ;
  assign n6616 = ~n6337 & ~n6615 ;
  assign n6617 = ~n6612 & n6616 ;
  assign n6379 = \P2_InstQueue_reg[13][4]/NET0131  & n1466 ;
  assign n6380 = \P2_InstQueue_reg[11][4]/NET0131  & n1459 ;
  assign n6393 = ~n6379 & ~n6380 ;
  assign n6381 = \P2_InstQueue_reg[2][4]/NET0131  & n1468 ;
  assign n6382 = \P2_InstQueue_reg[9][4]/NET0131  & n1472 ;
  assign n6394 = ~n6381 & ~n6382 ;
  assign n6401 = n6393 & n6394 ;
  assign n6375 = \P2_InstQueue_reg[5][4]/NET0131  & n1474 ;
  assign n6376 = \P2_InstQueue_reg[6][4]/NET0131  & n1447 ;
  assign n6391 = ~n6375 & ~n6376 ;
  assign n6377 = \P2_InstQueue_reg[12][4]/NET0131  & n1480 ;
  assign n6378 = \P2_InstQueue_reg[0][4]/NET0131  & n1456 ;
  assign n6392 = ~n6377 & ~n6378 ;
  assign n6402 = n6391 & n6392 ;
  assign n6403 = n6401 & n6402 ;
  assign n6387 = \P2_InstQueue_reg[7][4]/NET0131  & n1476 ;
  assign n6388 = \P2_InstQueue_reg[3][4]/NET0131  & n1470 ;
  assign n6397 = ~n6387 & ~n6388 ;
  assign n6389 = \P2_InstQueue_reg[10][4]/NET0131  & n1453 ;
  assign n6390 = \P2_InstQueue_reg[1][4]/NET0131  & n1464 ;
  assign n6398 = ~n6389 & ~n6390 ;
  assign n6399 = n6397 & n6398 ;
  assign n6383 = \P2_InstQueue_reg[4][4]/NET0131  & n1450 ;
  assign n6384 = \P2_InstQueue_reg[14][4]/NET0131  & n1482 ;
  assign n6395 = ~n6383 & ~n6384 ;
  assign n6385 = \P2_InstQueue_reg[15][4]/NET0131  & n1478 ;
  assign n6386 = \P2_InstQueue_reg[8][4]/NET0131  & n1461 ;
  assign n6396 = ~n6385 & ~n6386 ;
  assign n6400 = n6395 & n6396 ;
  assign n6404 = n6399 & n6400 ;
  assign n6405 = n6403 & n6404 ;
  assign n6465 = \P2_InstAddrPointer_reg[3]/NET0131  & n6464 ;
  assign n6466 = \P2_InstAddrPointer_reg[4]/NET0131  & n6465 ;
  assign n6618 = ~\P2_InstAddrPointer_reg[4]/NET0131  & ~n6465 ;
  assign n6619 = ~n6466 & ~n6618 ;
  assign n6620 = n6405 & ~n6619 ;
  assign n6411 = \P2_InstQueue_reg[10][3]/NET0131  & n1453 ;
  assign n6412 = \P2_InstQueue_reg[12][3]/NET0131  & n1480 ;
  assign n6425 = ~n6411 & ~n6412 ;
  assign n6413 = \P2_InstQueue_reg[13][3]/NET0131  & n1466 ;
  assign n6414 = \P2_InstQueue_reg[11][3]/NET0131  & n1459 ;
  assign n6426 = ~n6413 & ~n6414 ;
  assign n6433 = n6425 & n6426 ;
  assign n6407 = \P2_InstQueue_reg[9][3]/NET0131  & n1472 ;
  assign n6408 = \P2_InstQueue_reg[4][3]/NET0131  & n1450 ;
  assign n6423 = ~n6407 & ~n6408 ;
  assign n6409 = \P2_InstQueue_reg[3][3]/NET0131  & n1470 ;
  assign n6410 = \P2_InstQueue_reg[14][3]/NET0131  & n1482 ;
  assign n6424 = ~n6409 & ~n6410 ;
  assign n6434 = n6423 & n6424 ;
  assign n6435 = n6433 & n6434 ;
  assign n6419 = \P2_InstQueue_reg[15][3]/NET0131  & n1478 ;
  assign n6420 = \P2_InstQueue_reg[6][3]/NET0131  & n1447 ;
  assign n6429 = ~n6419 & ~n6420 ;
  assign n6421 = \P2_InstQueue_reg[5][3]/NET0131  & n1474 ;
  assign n6422 = \P2_InstQueue_reg[7][3]/NET0131  & n1476 ;
  assign n6430 = ~n6421 & ~n6422 ;
  assign n6431 = n6429 & n6430 ;
  assign n6415 = \P2_InstQueue_reg[8][3]/NET0131  & n1461 ;
  assign n6416 = \P2_InstQueue_reg[0][3]/NET0131  & n1456 ;
  assign n6427 = ~n6415 & ~n6416 ;
  assign n6417 = \P2_InstQueue_reg[2][3]/NET0131  & n1468 ;
  assign n6418 = \P2_InstQueue_reg[1][3]/NET0131  & n1464 ;
  assign n6428 = ~n6417 & ~n6418 ;
  assign n6432 = n6427 & n6428 ;
  assign n6436 = n6431 & n6432 ;
  assign n6437 = n6435 & n6436 ;
  assign n6621 = ~\P2_InstAddrPointer_reg[3]/NET0131  & ~n6464 ;
  assign n6622 = ~n6465 & ~n6621 ;
  assign n6623 = n6437 & ~n6622 ;
  assign n6624 = n6299 & ~n6611 ;
  assign n6625 = ~n6623 & ~n6624 ;
  assign n6626 = ~n6620 & n6625 ;
  assign n6627 = ~n6617 & n6626 ;
  assign n6628 = ~n6405 & n6619 ;
  assign n6629 = ~n6437 & n6622 ;
  assign n6630 = ~n6620 & n6629 ;
  assign n6631 = ~n6628 & ~n6630 ;
  assign n6632 = ~n6627 & n6631 ;
  assign n6205 = \P2_InstQueue_reg[12][6]/NET0131  & n1480 ;
  assign n6206 = \P2_InstQueue_reg[6][6]/NET0131  & n1447 ;
  assign n6219 = ~n6205 & ~n6206 ;
  assign n6207 = \P2_InstQueue_reg[2][6]/NET0131  & n1468 ;
  assign n6208 = \P2_InstQueue_reg[7][6]/NET0131  & n1476 ;
  assign n6220 = ~n6207 & ~n6208 ;
  assign n6227 = n6219 & n6220 ;
  assign n6201 = \P2_InstQueue_reg[5][6]/NET0131  & n1474 ;
  assign n6202 = \P2_InstQueue_reg[0][6]/NET0131  & n1456 ;
  assign n6217 = ~n6201 & ~n6202 ;
  assign n6203 = \P2_InstQueue_reg[9][6]/NET0131  & n1472 ;
  assign n6204 = \P2_InstQueue_reg[11][6]/NET0131  & n1459 ;
  assign n6218 = ~n6203 & ~n6204 ;
  assign n6228 = n6217 & n6218 ;
  assign n6229 = n6227 & n6228 ;
  assign n6213 = \P2_InstQueue_reg[15][6]/NET0131  & n1478 ;
  assign n6214 = \P2_InstQueue_reg[14][6]/NET0131  & n1482 ;
  assign n6223 = ~n6213 & ~n6214 ;
  assign n6215 = \P2_InstQueue_reg[10][6]/NET0131  & n1453 ;
  assign n6216 = \P2_InstQueue_reg[3][6]/NET0131  & n1470 ;
  assign n6224 = ~n6215 & ~n6216 ;
  assign n6225 = n6223 & n6224 ;
  assign n6209 = \P2_InstQueue_reg[4][6]/NET0131  & n1450 ;
  assign n6210 = \P2_InstQueue_reg[1][6]/NET0131  & n1464 ;
  assign n6221 = ~n6209 & ~n6210 ;
  assign n6211 = \P2_InstQueue_reg[13][6]/NET0131  & n1466 ;
  assign n6212 = \P2_InstQueue_reg[8][6]/NET0131  & n1461 ;
  assign n6222 = ~n6211 & ~n6212 ;
  assign n6226 = n6221 & n6222 ;
  assign n6230 = n6225 & n6226 ;
  assign n6231 = n6229 & n6230 ;
  assign n6467 = \P2_InstAddrPointer_reg[5]/NET0131  & n6466 ;
  assign n6468 = \P2_InstAddrPointer_reg[6]/NET0131  & n6467 ;
  assign n6604 = ~\P2_InstAddrPointer_reg[6]/NET0131  & ~n6467 ;
  assign n6605 = ~n6468 & ~n6604 ;
  assign n6606 = n6231 & ~n6605 ;
  assign n6239 = \P2_InstQueue_reg[13][5]/NET0131  & n1466 ;
  assign n6240 = \P2_InstQueue_reg[3][5]/NET0131  & n1470 ;
  assign n6253 = ~n6239 & ~n6240 ;
  assign n6241 = \P2_InstQueue_reg[1][5]/NET0131  & n1464 ;
  assign n6242 = \P2_InstQueue_reg[0][5]/NET0131  & n1456 ;
  assign n6254 = ~n6241 & ~n6242 ;
  assign n6261 = n6253 & n6254 ;
  assign n6235 = \P2_InstQueue_reg[7][5]/NET0131  & n1476 ;
  assign n6236 = \P2_InstQueue_reg[11][5]/NET0131  & n1459 ;
  assign n6251 = ~n6235 & ~n6236 ;
  assign n6237 = \P2_InstQueue_reg[9][5]/NET0131  & n1472 ;
  assign n6238 = \P2_InstQueue_reg[12][5]/NET0131  & n1480 ;
  assign n6252 = ~n6237 & ~n6238 ;
  assign n6262 = n6251 & n6252 ;
  assign n6263 = n6261 & n6262 ;
  assign n6247 = \P2_InstQueue_reg[10][5]/NET0131  & n1453 ;
  assign n6248 = \P2_InstQueue_reg[15][5]/NET0131  & n1478 ;
  assign n6257 = ~n6247 & ~n6248 ;
  assign n6249 = \P2_InstQueue_reg[5][5]/NET0131  & n1474 ;
  assign n6250 = \P2_InstQueue_reg[14][5]/NET0131  & n1482 ;
  assign n6258 = ~n6249 & ~n6250 ;
  assign n6259 = n6257 & n6258 ;
  assign n6243 = \P2_InstQueue_reg[8][5]/NET0131  & n1461 ;
  assign n6244 = \P2_InstQueue_reg[6][5]/NET0131  & n1447 ;
  assign n6255 = ~n6243 & ~n6244 ;
  assign n6245 = \P2_InstQueue_reg[2][5]/NET0131  & n1468 ;
  assign n6246 = \P2_InstQueue_reg[4][5]/NET0131  & n1450 ;
  assign n6256 = ~n6245 & ~n6246 ;
  assign n6260 = n6255 & n6256 ;
  assign n6264 = n6259 & n6260 ;
  assign n6265 = n6263 & n6264 ;
  assign n6607 = ~\P2_InstAddrPointer_reg[5]/NET0131  & ~n6466 ;
  assign n6608 = ~n6467 & ~n6607 ;
  assign n6609 = n6265 & ~n6608 ;
  assign n6633 = ~n6606 & ~n6609 ;
  assign n6634 = ~n6632 & n6633 ;
  assign n6163 = \P2_InstQueue_reg[12][7]/NET0131  & n1480 ;
  assign n6164 = \P2_InstQueue_reg[2][7]/NET0131  & n1468 ;
  assign n6176 = ~n6163 & ~n6164 ;
  assign n6165 = \P2_InstQueue_reg[6][7]/NET0131  & n1447 ;
  assign n6166 = \P2_InstQueue_reg[7][7]/NET0131  & n1476 ;
  assign n6177 = ~n6165 & ~n6166 ;
  assign n6183 = n6176 & n6177 ;
  assign n6156 = \P2_InstQueue_reg[14][7]/NET0131  & n1482 ;
  assign n6157 = \P2_InstQueue_reg[9][7]/NET0131  & n1472 ;
  assign n6174 = ~n6156 & ~n6157 ;
  assign n6161 = \P2_InstQueue_reg[0][7]/NET0131  & n1456 ;
  assign n6162 = \P2_InstQueue_reg[10][7]/NET0131  & n1453 ;
  assign n6175 = ~n6161 & ~n6162 ;
  assign n6184 = n6174 & n6175 ;
  assign n6185 = n6183 & n6184 ;
  assign n6158 = \P2_InstQueue_reg[5][7]/NET0131  & n1463 ;
  assign n6159 = n1444 & n6158 ;
  assign n6160 = n1860 & n6159 ;
  assign n6173 = \P2_InstQueue_reg[4][7]/NET0131  & n1450 ;
  assign n6171 = \P2_InstQueue_reg[13][7]/NET0131  & n1466 ;
  assign n6172 = \P2_InstQueue_reg[1][7]/NET0131  & n1464 ;
  assign n6180 = ~n6171 & ~n6172 ;
  assign n6181 = ~n6173 & n6180 ;
  assign n6167 = \P2_InstQueue_reg[8][7]/NET0131  & n1461 ;
  assign n6168 = \P2_InstQueue_reg[11][7]/NET0131  & n1459 ;
  assign n6178 = ~n6167 & ~n6168 ;
  assign n6169 = \P2_InstQueue_reg[15][7]/NET0131  & n1478 ;
  assign n6170 = \P2_InstQueue_reg[3][7]/NET0131  & n1470 ;
  assign n6179 = ~n6169 & ~n6170 ;
  assign n6182 = n6178 & n6179 ;
  assign n6186 = n6181 & n6182 ;
  assign n6187 = ~n6160 & n6186 ;
  assign n6188 = n6185 & n6187 ;
  assign n6469 = \P2_InstAddrPointer_reg[7]/NET0131  & n6468 ;
  assign n6599 = ~\P2_InstAddrPointer_reg[7]/NET0131  & ~n6468 ;
  assign n6600 = ~n6469 & ~n6599 ;
  assign n6635 = ~n6188 & n6600 ;
  assign n6636 = ~n6231 & n6605 ;
  assign n6637 = ~n6265 & n6608 ;
  assign n6638 = ~n6606 & n6637 ;
  assign n6639 = ~n6636 & ~n6638 ;
  assign n6640 = ~n6635 & n6639 ;
  assign n6641 = ~n6634 & n6640 ;
  assign n6601 = n6188 & ~n6600 ;
  assign n6470 = \P2_InstAddrPointer_reg[8]/NET0131  & n6469 ;
  assign n6602 = ~\P2_InstAddrPointer_reg[8]/NET0131  & ~n6469 ;
  assign n6603 = ~n6470 & ~n6602 ;
  assign n6642 = ~n6601 & n6603 ;
  assign n6643 = ~n6641 & n6642 ;
  assign n6493 = \P2_InstAddrPointer_reg[10]/NET0131  & \P2_InstAddrPointer_reg[11]/NET0131  ;
  assign n6494 = \P2_InstAddrPointer_reg[7]/NET0131  & \P2_InstAddrPointer_reg[8]/NET0131  ;
  assign n6495 = \P2_InstAddrPointer_reg[9]/NET0131  & n6494 ;
  assign n6496 = n6468 & n6495 ;
  assign n6644 = ~\P2_InstAddrPointer_reg[9]/NET0131  & ~n6470 ;
  assign n6645 = ~n6496 & ~n6644 ;
  assign n6646 = n6493 & n6645 ;
  assign n6647 = \P2_InstAddrPointer_reg[12]/NET0131  & n6646 ;
  assign n6648 = n6643 & n6647 ;
  assign n6497 = n6493 & n6496 ;
  assign n6498 = \P2_InstAddrPointer_reg[12]/NET0131  & \P2_InstAddrPointer_reg[13]/NET0131  ;
  assign n6499 = \P2_InstAddrPointer_reg[14]/NET0131  & n6498 ;
  assign n6500 = n6497 & n6499 ;
  assign n6463 = \P2_InstAddrPointer_reg[10]/NET0131  & \P2_InstAddrPointer_reg[9]/NET0131  ;
  assign n6471 = n6463 & n6470 ;
  assign n6475 = \P2_InstAddrPointer_reg[11]/NET0131  & \P2_InstAddrPointer_reg[12]/NET0131  ;
  assign n6489 = n6471 & n6475 ;
  assign n6490 = \P2_InstAddrPointer_reg[13]/NET0131  & n6489 ;
  assign n6649 = ~\P2_InstAddrPointer_reg[14]/NET0131  & ~n6490 ;
  assign n6650 = ~n6500 & ~n6649 ;
  assign n6651 = \P2_InstAddrPointer_reg[15]/NET0131  & n6650 ;
  assign n6652 = ~\P2_InstAddrPointer_reg[13]/NET0131  & ~n6489 ;
  assign n6653 = ~n6490 & ~n6652 ;
  assign n6654 = \P2_InstAddrPointer_reg[16]/NET0131  & n6653 ;
  assign n6655 = n6651 & n6654 ;
  assign n6656 = n6648 & n6655 ;
  assign n6510 = \P2_InstAddrPointer_reg[15]/NET0131  & \P2_InstAddrPointer_reg[16]/NET0131  ;
  assign n6511 = n6499 & n6510 ;
  assign n6657 = n6497 & n6511 ;
  assign n6659 = \P2_InstAddrPointer_reg[17]/NET0131  & n6657 ;
  assign n6661 = \P2_InstAddrPointer_reg[18]/NET0131  & n6659 ;
  assign n6662 = ~\P2_InstAddrPointer_reg[18]/NET0131  & ~n6659 ;
  assign n6663 = ~n6661 & ~n6662 ;
  assign n6664 = \P2_InstAddrPointer_reg[19]/NET0131  & n6663 ;
  assign n6658 = ~\P2_InstAddrPointer_reg[17]/NET0131  & ~n6657 ;
  assign n6660 = ~n6658 & ~n6659 ;
  assign n6529 = \P2_InstAddrPointer_reg[17]/NET0131  & n6510 ;
  assign n6530 = \P2_InstAddrPointer_reg[18]/NET0131  & \P2_InstAddrPointer_reg[19]/NET0131  ;
  assign n6531 = n6529 & n6530 ;
  assign n6532 = n6500 & n6531 ;
  assign n6535 = \P2_InstAddrPointer_reg[20]/NET0131  & n6532 ;
  assign n6665 = ~\P2_InstAddrPointer_reg[20]/NET0131  & ~n6532 ;
  assign n6666 = ~n6535 & ~n6665 ;
  assign n6667 = n6660 & n6666 ;
  assign n6668 = n6664 & n6667 ;
  assign n6669 = n6656 & n6668 ;
  assign n6593 = ~\P2_InstAddrPointer_reg[21]/NET0131  & ~n6535 ;
  assign n6544 = \P2_InstAddrPointer_reg[20]/NET0131  & \P2_InstAddrPointer_reg[21]/NET0131  ;
  assign n6594 = n6532 & n6544 ;
  assign n6595 = ~n6593 & ~n6594 ;
  assign n6557 = \P2_InstAddrPointer_reg[23]/NET0131  & \P2_InstAddrPointer_reg[24]/NET0131  ;
  assign n6548 = \P2_InstAddrPointer_reg[22]/NET0131  & n6544 ;
  assign n6556 = n6532 & n6548 ;
  assign n6596 = ~\P2_InstAddrPointer_reg[22]/NET0131  & ~n6594 ;
  assign n6597 = ~n6556 & ~n6596 ;
  assign n6598 = n6557 & n6597 ;
  assign n6670 = n6595 & n6598 ;
  assign n6671 = n6669 & n6670 ;
  assign n6558 = n6556 & n6557 ;
  assign n6564 = \P2_InstAddrPointer_reg[25]/NET0131  & n6558 ;
  assign n6672 = ~\P2_InstAddrPointer_reg[25]/NET0131  & ~n6558 ;
  assign n6673 = ~n6564 & ~n6672 ;
  assign n6674 = \P2_InstAddrPointer_reg[26]/NET0131  & n6673 ;
  assign n6574 = \P2_InstAddrPointer_reg[26]/NET0131  & \P2_InstAddrPointer_reg[27]/NET0131  ;
  assign n6584 = n6564 & n6574 ;
  assign n6567 = \P2_InstAddrPointer_reg[26]/NET0131  & n6564 ;
  assign n6675 = ~\P2_InstAddrPointer_reg[27]/NET0131  & ~n6567 ;
  assign n6676 = ~n6584 & ~n6675 ;
  assign n6677 = \P2_InstAddrPointer_reg[28]/NET0131  & n6676 ;
  assign n6678 = n6674 & n6677 ;
  assign n6679 = n6671 & n6678 ;
  assign n6585 = \P2_InstAddrPointer_reg[28]/NET0131  & n6584 ;
  assign n6586 = \P2_InstAddrPointer_reg[29]/NET0131  & n6585 ;
  assign n6680 = ~\P2_InstAddrPointer_reg[29]/NET0131  & ~n6585 ;
  assign n6681 = ~n6586 & ~n6680 ;
  assign n6683 = ~n6679 & n6681 ;
  assign n6682 = n6679 & ~n6681 ;
  assign n6684 = n6188 & ~n6682 ;
  assign n6685 = ~n6683 & n6684 ;
  assign n6189 = \P2_InstAddrPointer_reg[0]/NET0131  & \P2_InstAddrPointer_reg[1]/NET0131  ;
  assign n6190 = \P2_InstAddrPointer_reg[2]/NET0131  & n6189 ;
  assign n6191 = \P2_InstAddrPointer_reg[3]/NET0131  & n6190 ;
  assign n6192 = \P2_InstAddrPointer_reg[4]/NET0131  & n6191 ;
  assign n6193 = \P2_InstAddrPointer_reg[5]/NET0131  & n6192 ;
  assign n6194 = \P2_InstAddrPointer_reg[6]/NET0131  & n6193 ;
  assign n6195 = ~\P2_InstAddrPointer_reg[7]/NET0131  & ~n6194 ;
  assign n6196 = \P2_InstAddrPointer_reg[7]/NET0131  & n6194 ;
  assign n6197 = ~n6195 & ~n6196 ;
  assign n6198 = n6188 & ~n6197 ;
  assign n6199 = ~\P2_InstAddrPointer_reg[6]/NET0131  & ~n6193 ;
  assign n6200 = ~n6194 & ~n6199 ;
  assign n6232 = ~n6200 & n6231 ;
  assign n6233 = ~\P2_InstAddrPointer_reg[5]/NET0131  & ~n6192 ;
  assign n6234 = ~n6193 & ~n6233 ;
  assign n6266 = ~n6234 & n6265 ;
  assign n6267 = ~n6232 & ~n6266 ;
  assign n6268 = ~n6198 & n6267 ;
  assign n6300 = ~\P2_InstAddrPointer_reg[2]/NET0131  & ~n6189 ;
  assign n6301 = ~n6190 & ~n6300 ;
  assign n6302 = ~n6299 & n6301 ;
  assign n6334 = ~\P2_InstAddrPointer_reg[0]/NET0131  & ~\P2_InstAddrPointer_reg[1]/NET0131  ;
  assign n6335 = ~n6189 & ~n6334 ;
  assign n6336 = n6333 & ~n6335 ;
  assign n6369 = \P2_InstAddrPointer_reg[0]/NET0131  & n6368 ;
  assign n6370 = ~n6337 & n6369 ;
  assign n6371 = ~n6336 & ~n6370 ;
  assign n6372 = ~n6302 & ~n6371 ;
  assign n6373 = ~\P2_InstAddrPointer_reg[4]/NET0131  & ~n6191 ;
  assign n6374 = ~n6192 & ~n6373 ;
  assign n6406 = ~n6374 & n6405 ;
  assign n6438 = ~\P2_InstAddrPointer_reg[3]/NET0131  & ~n6190 ;
  assign n6439 = ~n6191 & ~n6438 ;
  assign n6440 = n6437 & ~n6439 ;
  assign n6441 = n6299 & ~n6301 ;
  assign n6442 = ~n6440 & ~n6441 ;
  assign n6443 = ~n6406 & n6442 ;
  assign n6444 = ~n6372 & n6443 ;
  assign n6445 = n6374 & ~n6405 ;
  assign n6446 = ~n6437 & n6439 ;
  assign n6447 = ~n6406 & n6446 ;
  assign n6448 = ~n6445 & ~n6447 ;
  assign n6449 = ~n6444 & n6448 ;
  assign n6450 = n6268 & ~n6449 ;
  assign n6451 = n6200 & ~n6231 ;
  assign n6452 = n6234 & ~n6265 ;
  assign n6453 = ~n6232 & n6452 ;
  assign n6454 = ~n6451 & ~n6453 ;
  assign n6455 = ~n6198 & ~n6454 ;
  assign n6456 = ~n6188 & n6197 ;
  assign n6457 = ~\P2_InstAddrPointer_reg[8]/NET0131  & ~n6196 ;
  assign n6458 = \P2_InstAddrPointer_reg[8]/NET0131  & n6196 ;
  assign n6459 = ~n6457 & ~n6458 ;
  assign n6460 = ~n6456 & ~n6459 ;
  assign n6461 = ~n6455 & n6460 ;
  assign n6462 = ~n6450 & n6461 ;
  assign n6472 = \P2_InstAddrPointer_reg[0]/NET0131  & n6471 ;
  assign n6473 = \P2_InstAddrPointer_reg[11]/NET0131  & n6472 ;
  assign n6474 = ~\P2_InstAddrPointer_reg[12]/NET0131  & ~n6473 ;
  assign n6476 = n6472 & n6475 ;
  assign n6477 = ~n6474 & ~n6476 ;
  assign n6478 = ~\P2_InstAddrPointer_reg[9]/NET0131  & ~n6458 ;
  assign n6479 = \P2_InstAddrPointer_reg[9]/NET0131  & n6458 ;
  assign n6480 = ~n6478 & ~n6479 ;
  assign n6481 = ~\P2_InstAddrPointer_reg[10]/NET0131  & ~n6479 ;
  assign n6482 = ~n6472 & ~n6481 ;
  assign n6483 = ~n6480 & ~n6482 ;
  assign n6484 = ~\P2_InstAddrPointer_reg[11]/NET0131  & ~n6472 ;
  assign n6485 = ~n6473 & ~n6484 ;
  assign n6486 = n6483 & ~n6485 ;
  assign n6487 = ~n6477 & n6486 ;
  assign n6488 = n6462 & n6487 ;
  assign n6491 = \P2_InstAddrPointer_reg[0]/NET0131  & n6490 ;
  assign n6492 = ~\P2_InstAddrPointer_reg[14]/NET0131  & ~n6491 ;
  assign n6501 = \P2_InstAddrPointer_reg[0]/NET0131  & n6500 ;
  assign n6502 = ~n6492 & ~n6501 ;
  assign n6503 = ~\P2_InstAddrPointer_reg[15]/NET0131  & ~n6501 ;
  assign n6504 = \P2_InstAddrPointer_reg[15]/NET0131  & n6499 ;
  assign n6505 = n6473 & n6504 ;
  assign n6506 = ~n6503 & ~n6505 ;
  assign n6507 = ~n6502 & ~n6506 ;
  assign n6508 = ~\P2_InstAddrPointer_reg[16]/NET0131  & ~n6473 ;
  assign n6509 = ~\P2_InstAddrPointer_reg[16]/NET0131  & ~n6504 ;
  assign n6512 = ~n6509 & ~n6511 ;
  assign n6513 = \P2_InstAddrPointer_reg[0]/NET0131  & ~n6512 ;
  assign n6514 = n6497 & n6513 ;
  assign n6515 = ~n6508 & ~n6514 ;
  assign n6516 = n6507 & ~n6515 ;
  assign n6517 = ~\P2_InstAddrPointer_reg[13]/NET0131  & ~n6476 ;
  assign n6518 = ~n6491 & ~n6517 ;
  assign n6519 = n6516 & ~n6518 ;
  assign n6520 = n6488 & n6519 ;
  assign n6521 = n6501 & n6510 ;
  assign n6522 = ~\P2_InstAddrPointer_reg[17]/NET0131  & ~n6521 ;
  assign n6523 = \P2_InstAddrPointer_reg[17]/NET0131  & n6521 ;
  assign n6524 = ~n6522 & ~n6523 ;
  assign n6525 = ~\P2_InstAddrPointer_reg[18]/NET0131  & ~n6523 ;
  assign n6526 = \P2_InstAddrPointer_reg[18]/NET0131  & n6523 ;
  assign n6527 = ~n6525 & ~n6526 ;
  assign n6528 = ~n6524 & ~n6527 ;
  assign n6533 = \P2_InstAddrPointer_reg[0]/NET0131  & n6532 ;
  assign n6534 = ~\P2_InstAddrPointer_reg[20]/NET0131  & ~n6533 ;
  assign n6536 = \P2_InstAddrPointer_reg[0]/NET0131  & n6535 ;
  assign n6537 = ~n6534 & ~n6536 ;
  assign n6538 = ~\P2_InstAddrPointer_reg[19]/NET0131  & ~n6526 ;
  assign n6539 = ~n6533 & ~n6538 ;
  assign n6540 = ~n6537 & ~n6539 ;
  assign n6541 = n6528 & n6540 ;
  assign n6542 = n6520 & n6541 ;
  assign n6543 = ~\P2_InstAddrPointer_reg[21]/NET0131  & ~n6536 ;
  assign n6545 = n6533 & n6544 ;
  assign n6546 = ~n6543 & ~n6545 ;
  assign n6547 = ~\P2_InstAddrPointer_reg[22]/NET0131  & ~n6545 ;
  assign n6549 = n6533 & n6548 ;
  assign n6550 = ~n6547 & ~n6549 ;
  assign n6551 = ~n6546 & ~n6550 ;
  assign n6552 = ~\P2_InstAddrPointer_reg[23]/NET0131  & ~n6549 ;
  assign n6553 = \P2_InstAddrPointer_reg[23]/NET0131  & n6549 ;
  assign n6554 = ~n6552 & ~n6553 ;
  assign n6555 = ~\P2_InstAddrPointer_reg[24]/NET0131  & ~n6553 ;
  assign n6559 = \P2_InstAddrPointer_reg[0]/NET0131  & n6558 ;
  assign n6560 = ~n6555 & ~n6559 ;
  assign n6561 = ~n6554 & ~n6560 ;
  assign n6562 = n6551 & n6561 ;
  assign n6563 = n6542 & n6562 ;
  assign n6565 = \P2_InstAddrPointer_reg[0]/NET0131  & n6564 ;
  assign n6566 = ~\P2_InstAddrPointer_reg[26]/NET0131  & ~n6565 ;
  assign n6568 = \P2_InstAddrPointer_reg[0]/NET0131  & n6567 ;
  assign n6569 = ~n6566 & ~n6568 ;
  assign n6570 = ~\P2_InstAddrPointer_reg[25]/NET0131  & ~n6559 ;
  assign n6571 = ~n6565 & ~n6570 ;
  assign n6572 = ~n6569 & ~n6571 ;
  assign n6573 = ~\P2_InstAddrPointer_reg[27]/NET0131  & ~n6568 ;
  assign n6575 = n6565 & n6574 ;
  assign n6576 = ~n6573 & ~n6575 ;
  assign n6577 = ~\P2_InstAddrPointer_reg[28]/NET0131  & ~n6575 ;
  assign n6578 = \P2_InstAddrPointer_reg[28]/NET0131  & n6575 ;
  assign n6579 = ~n6577 & ~n6578 ;
  assign n6580 = ~n6576 & ~n6579 ;
  assign n6581 = n6572 & n6580 ;
  assign n6582 = n6563 & n6581 ;
  assign n6583 = ~\P2_InstAddrPointer_reg[29]/NET0131  & ~n6578 ;
  assign n6587 = \P2_InstAddrPointer_reg[0]/NET0131  & n6586 ;
  assign n6588 = ~n6583 & ~n6587 ;
  assign n6590 = n6582 & ~n6588 ;
  assign n6589 = ~n6582 & n6588 ;
  assign n6591 = ~n6188 & ~n6589 ;
  assign n6592 = ~n6590 & n6591 ;
  assign n6686 = ~n1897 & ~n6592 ;
  assign n6687 = ~n6685 & n6686 ;
  assign n6688 = ~n6155 & ~n6687 ;
  assign n6689 = n1734 & ~n6688 ;
  assign n6690 = \P2_InstAddrPointer_reg[3]/NET0131  & ~n6300 ;
  assign n6691 = \P2_InstAddrPointer_reg[4]/NET0131  & n6690 ;
  assign n6692 = \P2_InstAddrPointer_reg[5]/NET0131  & n6691 ;
  assign n6693 = \P2_InstAddrPointer_reg[6]/NET0131  & n6692 ;
  assign n6694 = \P2_InstAddrPointer_reg[7]/NET0131  & n6693 ;
  assign n6695 = ~\P2_InstAddrPointer_reg[7]/NET0131  & ~n6693 ;
  assign n6696 = ~n6694 & ~n6695 ;
  assign n6697 = ~n6188 & n6696 ;
  assign n6698 = ~\P2_InstAddrPointer_reg[6]/NET0131  & ~n6692 ;
  assign n6699 = ~n6693 & ~n6698 ;
  assign n6700 = n6231 & ~n6699 ;
  assign n6701 = ~\P2_InstAddrPointer_reg[5]/NET0131  & ~n6691 ;
  assign n6702 = ~n6692 & ~n6701 ;
  assign n6703 = n6265 & ~n6702 ;
  assign n6704 = ~n6700 & ~n6703 ;
  assign n6705 = ~\P2_InstAddrPointer_reg[4]/NET0131  & ~n6690 ;
  assign n6706 = ~n6691 & ~n6705 ;
  assign n6707 = n6405 & ~n6706 ;
  assign n6708 = ~\P2_InstAddrPointer_reg[3]/NET0131  & n6300 ;
  assign n6709 = ~n6690 & ~n6708 ;
  assign n6710 = n6437 & ~n6709 ;
  assign n6711 = ~n6707 & ~n6710 ;
  assign n6712 = n6299 & n6301 ;
  assign n6713 = ~n6299 & ~n6301 ;
  assign n6714 = ~n6333 & n6335 ;
  assign n6715 = ~\P2_InstAddrPointer_reg[0]/NET0131  & ~n6368 ;
  assign n6716 = ~n6714 & ~n6715 ;
  assign n6717 = ~n6336 & ~n6716 ;
  assign n6718 = ~n6713 & ~n6717 ;
  assign n6719 = ~n6712 & ~n6718 ;
  assign n6720 = n6711 & n6719 ;
  assign n6721 = ~n6405 & n6706 ;
  assign n6722 = ~n6437 & n6709 ;
  assign n6723 = ~n6707 & n6722 ;
  assign n6724 = ~n6721 & ~n6723 ;
  assign n6725 = ~n6720 & n6724 ;
  assign n6726 = n6704 & ~n6725 ;
  assign n6727 = ~n6231 & n6699 ;
  assign n6728 = ~n6265 & n6702 ;
  assign n6729 = ~n6700 & n6728 ;
  assign n6730 = ~n6727 & ~n6729 ;
  assign n6731 = ~n6726 & n6730 ;
  assign n6732 = ~n6697 & n6731 ;
  assign n6733 = n6188 & ~n6696 ;
  assign n6734 = ~\P2_InstAddrPointer_reg[8]/NET0131  & ~n6694 ;
  assign n6735 = \P2_InstAddrPointer_reg[8]/NET0131  & n6694 ;
  assign n6736 = ~n6734 & ~n6735 ;
  assign n6737 = ~n6733 & n6736 ;
  assign n6738 = \P2_InstAddrPointer_reg[9]/NET0131  & n6737 ;
  assign n6739 = ~n6732 & n6738 ;
  assign n6740 = \P2_InstAddrPointer_reg[9]/NET0131  & n6735 ;
  assign n6741 = ~\P2_InstAddrPointer_reg[10]/NET0131  & ~n6740 ;
  assign n6742 = n6463 & n6735 ;
  assign n6743 = ~n6741 & ~n6742 ;
  assign n6744 = n6475 & n6743 ;
  assign n6745 = \P2_InstAddrPointer_reg[13]/NET0131  & n6744 ;
  assign n6746 = n6739 & n6745 ;
  assign n6747 = n6475 & n6742 ;
  assign n6748 = \P2_InstAddrPointer_reg[13]/NET0131  & n6747 ;
  assign n6749 = ~\P2_InstAddrPointer_reg[14]/NET0131  & ~n6748 ;
  assign n6750 = \P2_InstAddrPointer_reg[14]/NET0131  & n6748 ;
  assign n6751 = ~n6749 & ~n6750 ;
  assign n6752 = n6510 & n6751 ;
  assign n6753 = \P2_InstAddrPointer_reg[15]/NET0131  & n6750 ;
  assign n6754 = \P2_InstAddrPointer_reg[16]/NET0131  & n6753 ;
  assign n6755 = ~\P2_InstAddrPointer_reg[17]/NET0131  & ~n6754 ;
  assign n6756 = n6529 & n6750 ;
  assign n6757 = ~n6755 & ~n6756 ;
  assign n6758 = n6530 & n6757 ;
  assign n6759 = \P2_InstAddrPointer_reg[20]/NET0131  & n6758 ;
  assign n6760 = n6752 & n6759 ;
  assign n6761 = n6746 & n6760 ;
  assign n6762 = n6531 & n6750 ;
  assign n6763 = \P2_InstAddrPointer_reg[20]/NET0131  & n6762 ;
  assign n6764 = ~\P2_InstAddrPointer_reg[21]/NET0131  & ~n6763 ;
  assign n6765 = n6544 & n6762 ;
  assign n6766 = ~n6764 & ~n6765 ;
  assign n6767 = n6761 & n6766 ;
  assign n6768 = ~\P2_InstAddrPointer_reg[22]/NET0131  & ~n6765 ;
  assign n6769 = \P2_InstAddrPointer_reg[22]/NET0131  & n6765 ;
  assign n6770 = ~n6768 & ~n6769 ;
  assign n6771 = n6557 & n6770 ;
  assign n6772 = n6767 & n6771 ;
  assign n6773 = n6557 & n6769 ;
  assign n6774 = \P2_InstAddrPointer_reg[25]/NET0131  & n6773 ;
  assign n6775 = \P2_InstAddrPointer_reg[26]/NET0131  & n6774 ;
  assign n6776 = ~\P2_InstAddrPointer_reg[27]/NET0131  & ~n6775 ;
  assign n6777 = n6574 & n6774 ;
  assign n6778 = ~n6776 & ~n6777 ;
  assign n6779 = \P2_InstAddrPointer_reg[28]/NET0131  & n6778 ;
  assign n6780 = ~\P2_InstAddrPointer_reg[25]/NET0131  & ~n6773 ;
  assign n6781 = ~n6774 & ~n6780 ;
  assign n6782 = \P2_InstAddrPointer_reg[26]/NET0131  & n6781 ;
  assign n6783 = n6779 & n6782 ;
  assign n6784 = n6772 & n6783 ;
  assign n6785 = \P2_InstAddrPointer_reg[28]/NET0131  & n6777 ;
  assign n6786 = \P2_InstAddrPointer_reg[29]/NET0131  & n6785 ;
  assign n6787 = ~\P2_InstAddrPointer_reg[29]/NET0131  & ~n6785 ;
  assign n6788 = ~n6786 & ~n6787 ;
  assign n6790 = ~n6784 & ~n6788 ;
  assign n6789 = n6784 & n6788 ;
  assign n6791 = n1890 & ~n6789 ;
  assign n6792 = ~n6790 & n6791 ;
  assign n6793 = n1870 & n6788 ;
  assign n6798 = ~n1771 & n6588 ;
  assign n6794 = n1805 & n1845 ;
  assign n6795 = n1854 & n1903 ;
  assign n6796 = ~n6794 & n6795 ;
  assign n6797 = \P2_InstAddrPointer_reg[29]/NET0131  & ~n6796 ;
  assign n6799 = ~n1831 & n6681 ;
  assign n6800 = ~n6797 & ~n6799 ;
  assign n6801 = ~n6798 & n6800 ;
  assign n6802 = ~n6793 & n6801 ;
  assign n6803 = ~n6792 & n6802 ;
  assign n6804 = ~n6689 & n6803 ;
  assign n6805 = n1927 & ~n6804 ;
  assign n6806 = \P2_rEIP_reg[29]/NET0131  & n3113 ;
  assign n6807 = ~n1935 & n2985 ;
  assign n6808 = ~n1930 & ~n2979 ;
  assign n6809 = ~n3087 & n6808 ;
  assign n6810 = ~n6807 & n6809 ;
  assign n6811 = \P2_InstAddrPointer_reg[29]/NET0131  & ~n6810 ;
  assign n6812 = ~n6806 & ~n6811 ;
  assign n6813 = ~n6805 & n6812 ;
  assign n6826 = n4460 & n4502 ;
  assign n6840 = n4758 & n6826 ;
  assign n6841 = ~n4757 & n4762 ;
  assign n6842 = n4506 & n5969 ;
  assign n6843 = ~n6841 & n6842 ;
  assign n6844 = ~n6840 & ~n6843 ;
  assign n6835 = ~\P1_InstAddrPointer_reg[20]/NET0131  & ~n4471 ;
  assign n6836 = ~n4767 & ~n6835 ;
  assign n6837 = n5976 & n6836 ;
  assign n6845 = ~\P1_InstAddrPointer_reg[19]/NET0131  & ~n4775 ;
  assign n6846 = ~n4471 & ~n6845 ;
  assign n6847 = n6837 & n6846 ;
  assign n6848 = n4776 & n4791 ;
  assign n6849 = n6847 & n6848 ;
  assign n6850 = ~n6844 & n6849 ;
  assign n6851 = ~n4481 & ~n6850 ;
  assign n6816 = n4748 & ~n4752 ;
  assign n6817 = ~n4642 & ~n6816 ;
  assign n6814 = ~n4574 & ~n4608 ;
  assign n6815 = ~n4505 & ~n4540 ;
  assign n6818 = n6814 & n6815 ;
  assign n6819 = n6817 & n6818 ;
  assign n6820 = ~n4574 & n4751 ;
  assign n6821 = ~n4760 & ~n6820 ;
  assign n6822 = ~n4759 & n6821 ;
  assign n6823 = n6815 & ~n6822 ;
  assign n6824 = ~n4758 & ~n6823 ;
  assign n6825 = ~n6819 & n6824 ;
  assign n6827 = \P1_InstAddrPointer_reg[11]/NET0131  & n6826 ;
  assign n6828 = ~n6825 & n6827 ;
  assign n6829 = ~\P1_InstAddrPointer_reg[12]/NET0131  & ~n4464 ;
  assign n6830 = ~n4786 & ~n6829 ;
  assign n6831 = n4789 & n6830 ;
  assign n6832 = n6828 & n6831 ;
  assign n6833 = n4777 & n4785 ;
  assign n6834 = n6832 & n6833 ;
  assign n6838 = n4481 & n6837 ;
  assign n6839 = n6834 & n6838 ;
  assign n6852 = n4453 & ~n6839 ;
  assign n6853 = ~n6851 & n6852 ;
  assign n6854 = n4834 & ~n5951 ;
  assign n6855 = n5944 & ~n6854 ;
  assign n6856 = ~n4827 & ~n6855 ;
  assign n6857 = n5940 & n5942 ;
  assign n6858 = ~n6856 & n6857 ;
  assign n6859 = n4886 & ~n4931 ;
  assign n6860 = n6858 & n6859 ;
  assign n6861 = n4924 & n6860 ;
  assign n6862 = ~n4900 & n4929 ;
  assign n6863 = ~n4902 & n6862 ;
  assign n6864 = n6861 & n6863 ;
  assign n6866 = n4896 & n6864 ;
  assign n6865 = ~n4896 & ~n6864 ;
  assign n6867 = ~n4453 & ~n6865 ;
  assign n6868 = ~n6866 & n6867 ;
  assign n6869 = ~n6853 & ~n6868 ;
  assign n6870 = ~n2375 & ~n6869 ;
  assign n6871 = \P1_InstAddrPointer_reg[23]/NET0131  & n2375 ;
  assign n6872 = ~n6870 & ~n6871 ;
  assign n6873 = n2244 & ~n6872 ;
  assign n6876 = ~\P1_InstAddrPointer_reg[23]/NET0131  & ~n5048 ;
  assign n6877 = ~n5041 & ~n6876 ;
  assign n6878 = n4469 & n5032 ;
  assign n6879 = n4974 & n6878 ;
  assign n6880 = n5049 & n6879 ;
  assign n6881 = n6010 & n6880 ;
  assign n6883 = n6877 & n6881 ;
  assign n6882 = ~n6877 & ~n6881 ;
  assign n6884 = n2385 & ~n6882 ;
  assign n6885 = ~n6883 & n6884 ;
  assign n6893 = n2337 & ~n6877 ;
  assign n6892 = ~\P1_InstAddrPointer_reg[23]/NET0131  & ~n2337 ;
  assign n6894 = ~n2332 & ~n6892 ;
  assign n6895 = ~n6893 & n6894 ;
  assign n6886 = n2401 & n4475 ;
  assign n6887 = ~\P1_InstAddrPointer_reg[23]/NET0131  & ~n6886 ;
  assign n6888 = ~n2233 & n4481 ;
  assign n6889 = ~n2369 & ~n6888 ;
  assign n6890 = ~n2379 & n6889 ;
  assign n6891 = ~n6887 & ~n6890 ;
  assign n6874 = n2237 & n4481 ;
  assign n6875 = ~n2271 & n4896 ;
  assign n6896 = ~n6874 & ~n6875 ;
  assign n6897 = ~n6891 & n6896 ;
  assign n6898 = ~n6895 & n6897 ;
  assign n6899 = ~n6885 & n6898 ;
  assign n6900 = ~n6873 & n6899 ;
  assign n6901 = n2432 & ~n6900 ;
  assign n6902 = \P1_rEIP_reg[23]/NET0131  & n5092 ;
  assign n6903 = \P1_InstAddrPointer_reg[23]/NET0131  & ~n5098 ;
  assign n6904 = ~n6902 & ~n6903 ;
  assign n6905 = ~n6901 & n6904 ;
  assign n6906 = \datai[29]_pad  & ~n5137 ;
  assign n6907 = \buf1_reg[29]/NET0131  & n5137 ;
  assign n6908 = ~n6906 & ~n6907 ;
  assign n6909 = n5269 & ~n6908 ;
  assign n6910 = \datai[30]_pad  & ~n5137 ;
  assign n6911 = \buf1_reg[30]/NET0131  & n5137 ;
  assign n6912 = ~n6910 & ~n6911 ;
  assign n6913 = n6909 & ~n6912 ;
  assign n6914 = n5155 & ~n6913 ;
  assign n6915 = ~n5155 & n6913 ;
  assign n6916 = ~n6914 & ~n6915 ;
  assign n6917 = n5148 & ~n6916 ;
  assign n6918 = ~n5227 & n5277 ;
  assign n6919 = ~n5221 & n6918 ;
  assign n6920 = n5224 & ~n6919 ;
  assign n6921 = ~n5224 & n6919 ;
  assign n6922 = ~n6920 & ~n6921 ;
  assign n6923 = n5151 & n6922 ;
  assign n6924 = ~n6917 & ~n6923 ;
  assign n6925 = \P1_DataWidth_reg[1]/NET0131  & ~n6924 ;
  assign n6926 = ~n5108 & ~n5176 ;
  assign n6927 = \P1_InstQueue_reg[11][7]/NET0131  & ~n5104 ;
  assign n6928 = ~n5107 & n6927 ;
  assign n6929 = ~n6926 & ~n6928 ;
  assign n6930 = ~n5153 & ~n6929 ;
  assign n6931 = ~n6925 & ~n6930 ;
  assign n6932 = n2436 & ~n6931 ;
  assign n6933 = n5095 & ~n6929 ;
  assign n6934 = ~n2156 & n5104 ;
  assign n6935 = ~n6927 & ~n6934 ;
  assign n6936 = n3042 & ~n6935 ;
  assign n6937 = \P1_InstQueue_reg[11][7]/NET0131  & ~n5291 ;
  assign n6938 = ~n6936 & ~n6937 ;
  assign n6939 = ~n6933 & n6938 ;
  assign n6940 = ~n6932 & n6939 ;
  assign n6941 = n5334 & ~n6916 ;
  assign n6942 = n5336 & n6922 ;
  assign n6943 = ~n6941 & ~n6942 ;
  assign n6944 = \P1_DataWidth_reg[1]/NET0131  & ~n6943 ;
  assign n6945 = ~n5176 & ~n5327 ;
  assign n6946 = \P1_InstQueue_reg[0][7]/NET0131  & ~n5324 ;
  assign n6947 = ~n5326 & n6946 ;
  assign n6948 = ~n6945 & ~n6947 ;
  assign n6949 = ~n5338 & ~n6948 ;
  assign n6950 = ~n6944 & ~n6949 ;
  assign n6951 = n2436 & ~n6950 ;
  assign n6952 = n5095 & ~n6948 ;
  assign n6953 = ~n2156 & n5324 ;
  assign n6954 = ~n6946 & ~n6953 ;
  assign n6955 = n3042 & ~n6954 ;
  assign n6956 = \P1_InstQueue_reg[0][7]/NET0131  & ~n5291 ;
  assign n6957 = ~n6955 & ~n6956 ;
  assign n6958 = ~n6952 & n6957 ;
  assign n6959 = ~n6951 & n6958 ;
  assign n6960 = n5359 & ~n6916 ;
  assign n6961 = n5148 & n6922 ;
  assign n6962 = ~n6960 & ~n6961 ;
  assign n6963 = \P1_DataWidth_reg[1]/NET0131  & ~n6962 ;
  assign n6964 = ~n5176 & ~n5353 ;
  assign n6965 = \P1_InstQueue_reg[10][7]/NET0131  & ~n5107 ;
  assign n6966 = ~n5151 & n6965 ;
  assign n6967 = ~n6964 & ~n6966 ;
  assign n6968 = ~n5361 & ~n6967 ;
  assign n6969 = ~n6963 & ~n6968 ;
  assign n6970 = n2436 & ~n6969 ;
  assign n6971 = n5095 & ~n6967 ;
  assign n6972 = ~n2156 & n5107 ;
  assign n6973 = ~n6965 & ~n6972 ;
  assign n6974 = n3042 & ~n6973 ;
  assign n6975 = \P1_InstQueue_reg[10][7]/NET0131  & ~n5291 ;
  assign n6976 = ~n6974 & ~n6975 ;
  assign n6977 = ~n6971 & n6976 ;
  assign n6978 = ~n6970 & n6977 ;
  assign n6979 = n5151 & ~n6916 ;
  assign n6980 = n5107 & n6922 ;
  assign n6981 = ~n6979 & ~n6980 ;
  assign n6982 = \P1_DataWidth_reg[1]/NET0131  & ~n6981 ;
  assign n6983 = ~n5176 & ~n5378 ;
  assign n6984 = \P1_InstQueue_reg[12][7]/NET0131  & ~n5377 ;
  assign n6985 = ~n5104 & n6984 ;
  assign n6986 = ~n6983 & ~n6985 ;
  assign n6987 = ~n5384 & ~n6986 ;
  assign n6988 = ~n6982 & ~n6987 ;
  assign n6989 = n2436 & ~n6988 ;
  assign n6990 = n5095 & ~n6986 ;
  assign n6991 = ~n2156 & n5377 ;
  assign n6992 = ~n6984 & ~n6991 ;
  assign n6993 = n3042 & ~n6992 ;
  assign n6994 = \P1_InstQueue_reg[12][7]/NET0131  & ~n5291 ;
  assign n6995 = ~n6993 & ~n6994 ;
  assign n6996 = ~n6990 & n6995 ;
  assign n6997 = ~n6989 & n6996 ;
  assign n6998 = n5107 & ~n6916 ;
  assign n6999 = n5104 & n6922 ;
  assign n7000 = ~n6998 & ~n6999 ;
  assign n7001 = \P1_DataWidth_reg[1]/NET0131  & ~n7000 ;
  assign n7002 = ~n5176 & ~n5399 ;
  assign n7003 = \P1_InstQueue_reg[13][7]/NET0131  & ~n5334 ;
  assign n7004 = ~n5377 & n7003 ;
  assign n7005 = ~n7002 & ~n7004 ;
  assign n7006 = ~n5405 & ~n7005 ;
  assign n7007 = ~n7001 & ~n7006 ;
  assign n7008 = n2436 & ~n7007 ;
  assign n7009 = n5095 & ~n7005 ;
  assign n7010 = ~n2156 & n5334 ;
  assign n7011 = ~n7003 & ~n7010 ;
  assign n7012 = n3042 & ~n7011 ;
  assign n7013 = \P1_InstQueue_reg[13][7]/NET0131  & ~n5291 ;
  assign n7014 = ~n7012 & ~n7013 ;
  assign n7015 = ~n7009 & n7014 ;
  assign n7016 = ~n7008 & n7015 ;
  assign n7017 = n5104 & ~n6916 ;
  assign n7018 = n5377 & n6922 ;
  assign n7019 = ~n7017 & ~n7018 ;
  assign n7020 = \P1_DataWidth_reg[1]/NET0131  & ~n7019 ;
  assign n7021 = ~n5176 & ~n5337 ;
  assign n7022 = \P1_InstQueue_reg[14][7]/NET0131  & ~n5336 ;
  assign n7023 = ~n5334 & n7022 ;
  assign n7024 = ~n7021 & ~n7023 ;
  assign n7025 = ~n5425 & ~n7024 ;
  assign n7026 = ~n7020 & ~n7025 ;
  assign n7027 = n2436 & ~n7026 ;
  assign n7028 = n5095 & ~n7024 ;
  assign n7029 = ~n2156 & n5336 ;
  assign n7030 = ~n7022 & ~n7029 ;
  assign n7031 = n3042 & ~n7030 ;
  assign n7032 = \P1_InstQueue_reg[14][7]/NET0131  & ~n5291 ;
  assign n7033 = ~n7031 & ~n7032 ;
  assign n7034 = ~n7028 & n7033 ;
  assign n7035 = ~n7027 & n7034 ;
  assign n7036 = n5377 & ~n6916 ;
  assign n7037 = n5334 & n6922 ;
  assign n7038 = ~n7036 & ~n7037 ;
  assign n7039 = \P1_DataWidth_reg[1]/NET0131  & ~n7038 ;
  assign n7040 = ~n5176 & ~n5440 ;
  assign n7041 = \P1_InstQueue_reg[15][7]/NET0131  & ~n5326 ;
  assign n7042 = ~n5336 & n7041 ;
  assign n7043 = ~n7040 & ~n7042 ;
  assign n7044 = ~n5446 & ~n7043 ;
  assign n7045 = ~n7039 & ~n7044 ;
  assign n7046 = n2436 & ~n7045 ;
  assign n7047 = n5095 & ~n7043 ;
  assign n7048 = ~n2156 & n5326 ;
  assign n7049 = ~n7041 & ~n7048 ;
  assign n7050 = n3042 & ~n7049 ;
  assign n7051 = \P1_InstQueue_reg[15][7]/NET0131  & ~n5291 ;
  assign n7052 = ~n7050 & ~n7051 ;
  assign n7053 = ~n7047 & n7052 ;
  assign n7054 = ~n7046 & n7053 ;
  assign n7055 = n5336 & ~n6916 ;
  assign n7056 = n5326 & n6922 ;
  assign n7057 = ~n7055 & ~n7056 ;
  assign n7058 = \P1_DataWidth_reg[1]/NET0131  & ~n7057 ;
  assign n7059 = ~n5176 & ~n5462 ;
  assign n7060 = \P1_InstQueue_reg[1][7]/NET0131  & ~n5461 ;
  assign n7061 = ~n5324 & n7060 ;
  assign n7062 = ~n7059 & ~n7061 ;
  assign n7063 = ~n5468 & ~n7062 ;
  assign n7064 = ~n7058 & ~n7063 ;
  assign n7065 = n2436 & ~n7064 ;
  assign n7066 = n5095 & ~n7062 ;
  assign n7067 = ~n2156 & n5461 ;
  assign n7068 = ~n7060 & ~n7067 ;
  assign n7069 = n3042 & ~n7068 ;
  assign n7070 = \P1_InstQueue_reg[1][7]/NET0131  & ~n5291 ;
  assign n7071 = ~n7069 & ~n7070 ;
  assign n7072 = ~n7066 & n7071 ;
  assign n7073 = ~n7065 & n7072 ;
  assign n7074 = n5326 & ~n6916 ;
  assign n7075 = n5324 & n6922 ;
  assign n7076 = ~n7074 & ~n7075 ;
  assign n7077 = \P1_DataWidth_reg[1]/NET0131  & ~n7076 ;
  assign n7078 = ~n5176 & ~n5506 ;
  assign n7079 = \P1_InstQueue_reg[2][7]/NET0131  & ~n5484 ;
  assign n7080 = ~n5461 & n7079 ;
  assign n7081 = ~n7078 & ~n7080 ;
  assign n7082 = ~n5512 & ~n7081 ;
  assign n7083 = ~n7077 & ~n7082 ;
  assign n7084 = n2436 & ~n7083 ;
  assign n7085 = n5095 & ~n7081 ;
  assign n7086 = ~n2156 & n5484 ;
  assign n7087 = ~n7079 & ~n7086 ;
  assign n7088 = n3042 & ~n7087 ;
  assign n7089 = \P1_InstQueue_reg[2][7]/NET0131  & ~n5291 ;
  assign n7090 = ~n7088 & ~n7089 ;
  assign n7091 = ~n7085 & n7090 ;
  assign n7092 = ~n7084 & n7091 ;
  assign n7093 = n5324 & ~n6916 ;
  assign n7094 = n5461 & n6922 ;
  assign n7095 = ~n7093 & ~n7094 ;
  assign n7096 = \P1_DataWidth_reg[1]/NET0131  & ~n7095 ;
  assign n7097 = ~n5176 & ~n5485 ;
  assign n7098 = \P1_InstQueue_reg[3][7]/NET0131  & ~n5483 ;
  assign n7099 = ~n5484 & n7098 ;
  assign n7100 = ~n7097 & ~n7099 ;
  assign n7101 = ~n5491 & ~n7100 ;
  assign n7102 = ~n7096 & ~n7101 ;
  assign n7103 = n2436 & ~n7102 ;
  assign n7104 = n5095 & ~n7100 ;
  assign n7105 = ~n2156 & n5483 ;
  assign n7106 = ~n7098 & ~n7105 ;
  assign n7107 = n3042 & ~n7106 ;
  assign n7108 = \P1_InstQueue_reg[3][7]/NET0131  & ~n5291 ;
  assign n7109 = ~n7107 & ~n7108 ;
  assign n7110 = ~n7104 & n7109 ;
  assign n7111 = ~n7103 & n7110 ;
  assign n7112 = n5461 & ~n6916 ;
  assign n7113 = n5484 & n6922 ;
  assign n7114 = ~n7112 & ~n7113 ;
  assign n7115 = \P1_DataWidth_reg[1]/NET0131  & ~n7114 ;
  assign n7116 = ~n5176 & ~n5528 ;
  assign n7117 = \P1_InstQueue_reg[4][7]/NET0131  & ~n5527 ;
  assign n7118 = ~n5483 & n7117 ;
  assign n7119 = ~n7116 & ~n7118 ;
  assign n7120 = ~n5534 & ~n7119 ;
  assign n7121 = ~n7115 & ~n7120 ;
  assign n7122 = n2436 & ~n7121 ;
  assign n7123 = n5095 & ~n7119 ;
  assign n7124 = ~n2156 & n5527 ;
  assign n7125 = ~n7117 & ~n7124 ;
  assign n7126 = n3042 & ~n7125 ;
  assign n7127 = \P1_InstQueue_reg[4][7]/NET0131  & ~n5291 ;
  assign n7128 = ~n7126 & ~n7127 ;
  assign n7129 = ~n7123 & n7128 ;
  assign n7130 = ~n7122 & n7129 ;
  assign n7131 = n5484 & ~n6916 ;
  assign n7132 = n5483 & n6922 ;
  assign n7133 = ~n7131 & ~n7132 ;
  assign n7134 = \P1_DataWidth_reg[1]/NET0131  & ~n7133 ;
  assign n7135 = ~n5176 & ~n5550 ;
  assign n7136 = \P1_InstQueue_reg[5][7]/NET0131  & ~n5549 ;
  assign n7137 = ~n5527 & n7136 ;
  assign n7138 = ~n7135 & ~n7137 ;
  assign n7139 = ~n5556 & ~n7138 ;
  assign n7140 = ~n7134 & ~n7139 ;
  assign n7141 = n2436 & ~n7140 ;
  assign n7142 = n5095 & ~n7138 ;
  assign n7143 = ~n2156 & n5549 ;
  assign n7144 = ~n7136 & ~n7143 ;
  assign n7145 = n3042 & ~n7144 ;
  assign n7146 = \P1_InstQueue_reg[5][7]/NET0131  & ~n5291 ;
  assign n7147 = ~n7145 & ~n7146 ;
  assign n7148 = ~n7142 & n7147 ;
  assign n7149 = ~n7141 & n7148 ;
  assign n7150 = n5483 & ~n6916 ;
  assign n7151 = n5527 & n6922 ;
  assign n7152 = ~n7150 & ~n7151 ;
  assign n7153 = \P1_DataWidth_reg[1]/NET0131  & ~n7152 ;
  assign n7154 = ~n5176 & ~n5572 ;
  assign n7155 = \P1_InstQueue_reg[6][7]/NET0131  & ~n5571 ;
  assign n7156 = ~n5549 & n7155 ;
  assign n7157 = ~n7154 & ~n7156 ;
  assign n7158 = ~n5578 & ~n7157 ;
  assign n7159 = ~n7153 & ~n7158 ;
  assign n7160 = n2436 & ~n7159 ;
  assign n7161 = n5095 & ~n7157 ;
  assign n7162 = ~n2156 & n5571 ;
  assign n7163 = ~n7155 & ~n7162 ;
  assign n7164 = n3042 & ~n7163 ;
  assign n7165 = \P1_InstQueue_reg[6][7]/NET0131  & ~n5291 ;
  assign n7166 = ~n7164 & ~n7165 ;
  assign n7167 = ~n7161 & n7166 ;
  assign n7168 = ~n7160 & n7167 ;
  assign n7169 = n5527 & ~n6916 ;
  assign n7170 = n5549 & n6922 ;
  assign n7171 = ~n7169 & ~n7170 ;
  assign n7172 = \P1_DataWidth_reg[1]/NET0131  & ~n7171 ;
  assign n7173 = ~n5176 & ~n5593 ;
  assign n7174 = \P1_InstQueue_reg[7][7]/NET0131  & ~n5359 ;
  assign n7175 = ~n5571 & n7174 ;
  assign n7176 = ~n7173 & ~n7175 ;
  assign n7177 = ~n5599 & ~n7176 ;
  assign n7178 = ~n7172 & ~n7177 ;
  assign n7179 = n2436 & ~n7178 ;
  assign n7180 = n5095 & ~n7176 ;
  assign n7181 = ~n2156 & n5359 ;
  assign n7182 = ~n7174 & ~n7181 ;
  assign n7183 = n3042 & ~n7182 ;
  assign n7184 = \P1_InstQueue_reg[7][7]/NET0131  & ~n5291 ;
  assign n7185 = ~n7183 & ~n7184 ;
  assign n7186 = ~n7180 & n7185 ;
  assign n7187 = ~n7179 & n7186 ;
  assign n7188 = n5549 & ~n6916 ;
  assign n7189 = n5571 & n6922 ;
  assign n7190 = ~n7188 & ~n7189 ;
  assign n7191 = \P1_DataWidth_reg[1]/NET0131  & ~n7190 ;
  assign n7192 = ~n5176 & ~n5360 ;
  assign n7193 = \P1_InstQueue_reg[8][7]/NET0131  & ~n5148 ;
  assign n7194 = ~n5359 & n7193 ;
  assign n7195 = ~n7192 & ~n7194 ;
  assign n7196 = ~n5619 & ~n7195 ;
  assign n7197 = ~n7191 & ~n7196 ;
  assign n7198 = n2436 & ~n7197 ;
  assign n7199 = n5095 & ~n7195 ;
  assign n7200 = ~n2156 & n5148 ;
  assign n7201 = ~n7193 & ~n7200 ;
  assign n7202 = n3042 & ~n7201 ;
  assign n7203 = \P1_InstQueue_reg[8][7]/NET0131  & ~n5291 ;
  assign n7204 = ~n7202 & ~n7203 ;
  assign n7205 = ~n7199 & n7204 ;
  assign n7206 = ~n7198 & n7205 ;
  assign n7207 = n5571 & ~n6916 ;
  assign n7208 = n5359 & n6922 ;
  assign n7209 = ~n7207 & ~n7208 ;
  assign n7210 = \P1_DataWidth_reg[1]/NET0131  & ~n7209 ;
  assign n7211 = ~n5152 & ~n5176 ;
  assign n7212 = \P1_InstQueue_reg[9][7]/NET0131  & ~n5151 ;
  assign n7213 = ~n5148 & n7212 ;
  assign n7214 = ~n7211 & ~n7213 ;
  assign n7215 = ~n5639 & ~n7214 ;
  assign n7216 = ~n7210 & ~n7215 ;
  assign n7217 = n2436 & ~n7216 ;
  assign n7218 = n5095 & ~n7214 ;
  assign n7219 = ~n2156 & n5151 ;
  assign n7220 = ~n7212 & ~n7219 ;
  assign n7221 = n3042 & ~n7220 ;
  assign n7222 = \P1_InstQueue_reg[9][7]/NET0131  & ~n5291 ;
  assign n7223 = ~n7221 & ~n7222 ;
  assign n7224 = ~n7218 & n7223 ;
  assign n7225 = ~n7217 & n7224 ;
  assign n7228 = \P1_InstAddrPointer_reg[26]/NET0131  & n2375 ;
  assign n7233 = ~\P1_InstAddrPointer_reg[26]/NET0131  & ~n4484 ;
  assign n7234 = ~n4489 & ~n7233 ;
  assign n7235 = n4482 & n5976 ;
  assign n7236 = n4486 & n7235 ;
  assign n7237 = n5975 & n7236 ;
  assign n7239 = ~n7234 & n7237 ;
  assign n7238 = n7234 & ~n7237 ;
  assign n7240 = n4453 & ~n7238 ;
  assign n7241 = ~n7239 & n7240 ;
  assign n7230 = n4935 & ~n4940 ;
  assign n7229 = ~n4935 & n4940 ;
  assign n7231 = ~n4453 & ~n7229 ;
  assign n7232 = ~n7230 & n7231 ;
  assign n7242 = ~n2375 & ~n7232 ;
  assign n7243 = ~n7241 & n7242 ;
  assign n7244 = ~n7228 & ~n7243 ;
  assign n7245 = n2244 & ~n7244 ;
  assign n7252 = ~n5053 & ~n5056 ;
  assign n7253 = n2385 & ~n5057 ;
  assign n7254 = ~n7252 & n7253 ;
  assign n7257 = ~n2337 & n5044 ;
  assign n7258 = ~n2332 & ~n7257 ;
  assign n7259 = n5056 & n7258 ;
  assign n7246 = n2222 & ~n2301 ;
  assign n7247 = ~n2302 & ~n7246 ;
  assign n7248 = n2317 & ~n7247 ;
  assign n7249 = ~n2389 & ~n7248 ;
  assign n7250 = n6026 & n7249 ;
  assign n7251 = \P1_InstAddrPointer_reg[26]/NET0131  & ~n7250 ;
  assign n7255 = ~n2271 & n4940 ;
  assign n7256 = ~n2402 & n7234 ;
  assign n7260 = ~n7255 & ~n7256 ;
  assign n7261 = ~n7251 & n7260 ;
  assign n7262 = ~n7259 & n7261 ;
  assign n7263 = ~n7254 & n7262 ;
  assign n7264 = ~n7245 & n7263 ;
  assign n7265 = n2432 & ~n7264 ;
  assign n7226 = \P1_rEIP_reg[26]/NET0131  & n5092 ;
  assign n7227 = \P1_InstAddrPointer_reg[26]/NET0131  & ~n5098 ;
  assign n7266 = ~n7226 & ~n7227 ;
  assign n7267 = ~n7265 & n7266 ;
  assign n7270 = \P1_InstAddrPointer_reg[24]/NET0131  & n2375 ;
  assign n7286 = n5975 & n7235 ;
  assign n7287 = ~\P1_InstAddrPointer_reg[24]/NET0131  & ~n4479 ;
  assign n7288 = ~n4483 & ~n7287 ;
  assign n7289 = ~n6839 & ~n7288 ;
  assign n7290 = ~n7286 & ~n7289 ;
  assign n7291 = n4453 & ~n7290 ;
  assign n7271 = ~n4863 & ~n4867 ;
  assign n7272 = ~n4869 & n5941 ;
  assign n7273 = n7271 & n7272 ;
  assign n7274 = ~n4913 & ~n4931 ;
  assign n7275 = n4885 & n7274 ;
  assign n7276 = n7273 & n7275 ;
  assign n7277 = n4923 & ~n4926 ;
  assign n7278 = n7276 & n7277 ;
  assign n7279 = ~n4928 & n7278 ;
  assign n7280 = n4904 & n7279 ;
  assign n7281 = n4893 & ~n7280 ;
  assign n7282 = n4933 & n5957 ;
  assign n7283 = n4905 & n7282 ;
  assign n7284 = ~n4453 & ~n7283 ;
  assign n7285 = ~n7281 & n7284 ;
  assign n7292 = ~n2375 & ~n7285 ;
  assign n7293 = ~n7291 & n7292 ;
  assign n7294 = ~n7270 & ~n7293 ;
  assign n7295 = n2244 & ~n7294 ;
  assign n7297 = ~\P1_InstAddrPointer_reg[24]/NET0131  & ~n5041 ;
  assign n7298 = ~n5042 & ~n7297 ;
  assign n7299 = \P1_InstAddrPointer_reg[10]/NET0131  & n5020 ;
  assign n7300 = n6009 & n7299 ;
  assign n7301 = n6011 & n7300 ;
  assign n7302 = n5050 & n5993 ;
  assign n7303 = n7301 & n7302 ;
  assign n7305 = n7298 & n7303 ;
  assign n7304 = ~n7298 & ~n7303 ;
  assign n7306 = n2385 & ~n7304 ;
  assign n7307 = ~n7305 & n7306 ;
  assign n7308 = ~n2301 & ~n2306 ;
  assign n7309 = \P1_InstAddrPointer_reg[24]/NET0131  & n7308 ;
  assign n7310 = n2314 & ~n7309 ;
  assign n7314 = n2317 & ~n7310 ;
  assign n7315 = n2311 & n7308 ;
  assign n7316 = n6026 & ~n7315 ;
  assign n7317 = ~n7314 & n7316 ;
  assign n7318 = \P1_InstAddrPointer_reg[24]/NET0131  & ~n7317 ;
  assign n7311 = ~n2317 & ~n7310 ;
  assign n7312 = ~n2237 & ~n7311 ;
  assign n7313 = n7288 & ~n7312 ;
  assign n7296 = ~n2271 & n4893 ;
  assign n7319 = n2397 & n7298 ;
  assign n7320 = ~n7296 & ~n7319 ;
  assign n7321 = ~n7313 & n7320 ;
  assign n7322 = ~n7318 & n7321 ;
  assign n7323 = ~n7307 & n7322 ;
  assign n7324 = ~n7295 & n7323 ;
  assign n7325 = n2432 & ~n7324 ;
  assign n7268 = \P1_rEIP_reg[24]/NET0131  & n5092 ;
  assign n7269 = \P1_InstAddrPointer_reg[24]/NET0131  & ~n5098 ;
  assign n7326 = ~n7268 & ~n7269 ;
  assign n7327 = ~n7325 & n7326 ;
  assign n7331 = \P3_InstAddrPointer_reg[15]/NET0131  & n2896 ;
  assign n7337 = n4232 & ~n4243 ;
  assign n7336 = ~n4232 & n4243 ;
  assign n7338 = ~n3753 & ~n7336 ;
  assign n7339 = ~n7337 & n7338 ;
  assign n7332 = ~n4075 & ~n4082 ;
  assign n7333 = n6088 & n6090 ;
  assign n7334 = ~n7332 & ~n7333 ;
  assign n7335 = n3753 & ~n7334 ;
  assign n7340 = ~n2896 & ~n7335 ;
  assign n7341 = ~n7339 & n7340 ;
  assign n7342 = ~n7331 & ~n7341 ;
  assign n7343 = n2894 & ~n7342 ;
  assign n7345 = \P3_InstAddrPointer_reg[15]/NET0131  & n4353 ;
  assign n7346 = ~\P3_InstAddrPointer_reg[15]/NET0131  & ~n4353 ;
  assign n7347 = ~n7345 & ~n7346 ;
  assign n7351 = n4349 & n4354 ;
  assign n7353 = ~n7347 & ~n7351 ;
  assign n7352 = \P3_InstAddrPointer_reg[15]/NET0131  & n7351 ;
  assign n7354 = n2905 & ~n7352 ;
  assign n7355 = ~n7353 & n7354 ;
  assign n7356 = ~n2923 & n3783 ;
  assign n7357 = ~\P3_InstAddrPointer_reg[15]/NET0131  & ~n7356 ;
  assign n7358 = n2891 & n4077 ;
  assign n7359 = ~n2768 & ~n7358 ;
  assign n7360 = ~n7357 & n7359 ;
  assign n7330 = ~n2777 & n4243 ;
  assign n7344 = ~\P3_InstAddrPointer_reg[15]/NET0131  & ~n2847 ;
  assign n7348 = ~n2841 & n7347 ;
  assign n7349 = n2901 & ~n7348 ;
  assign n7350 = ~n7344 & ~n7349 ;
  assign n7361 = ~n7330 & ~n7350 ;
  assign n7362 = ~n7360 & n7361 ;
  assign n7363 = ~n7355 & n7362 ;
  assign n7364 = ~n7343 & n7363 ;
  assign n7365 = n2453 & ~n7364 ;
  assign n7328 = \P3_rEIP_reg[15]/NET0131  & n4412 ;
  assign n7329 = \P3_InstAddrPointer_reg[15]/NET0131  & ~n4418 ;
  assign n7366 = ~n7328 & ~n7329 ;
  assign n7367 = ~n7365 & n7366 ;
  assign n7368 = \P3_InstAddrPointer_reg[22]/NET0131  & n2896 ;
  assign n7382 = n4080 & n7333 ;
  assign n7379 = ~\P3_InstAddrPointer_reg[18]/NET0131  & ~n3784 ;
  assign n7380 = n3796 & ~n7379 ;
  assign n7381 = n3792 & n7380 ;
  assign n7383 = n3789 & n7381 ;
  assign n7384 = n7382 & n7383 ;
  assign n7386 = ~n3776 & n7384 ;
  assign n7385 = n3776 & ~n7384 ;
  assign n7387 = n3753 & ~n7385 ;
  assign n7388 = ~n7386 & n7387 ;
  assign n7369 = ~n4171 & n4244 ;
  assign n7370 = ~n4175 & n6045 ;
  assign n7371 = n6058 & n7370 ;
  assign n7372 = n7369 & n7371 ;
  assign n7373 = n4258 & n6061 ;
  assign n7374 = n7372 & n7373 ;
  assign n7376 = ~n4269 & n7374 ;
  assign n7375 = n4269 & ~n7374 ;
  assign n7377 = ~n3753 & ~n7375 ;
  assign n7378 = ~n7376 & n7377 ;
  assign n7389 = ~n2896 & ~n7378 ;
  assign n7390 = ~n7388 & n7389 ;
  assign n7391 = ~n7368 & ~n7390 ;
  assign n7392 = n2894 & ~n7391 ;
  assign n7394 = n4368 & n6127 ;
  assign n7396 = ~n4371 & ~n7394 ;
  assign n7395 = \P3_InstAddrPointer_reg[22]/NET0131  & n7394 ;
  assign n7397 = n2905 & ~n7395 ;
  assign n7398 = ~n7396 & n7397 ;
  assign n7401 = ~n2834 & n2835 ;
  assign n7402 = ~n2825 & ~n2900 ;
  assign n7403 = ~n7401 & n7402 ;
  assign n7404 = ~n2898 & n7403 ;
  assign n7405 = \P3_InstAddrPointer_reg[22]/NET0131  & ~n7404 ;
  assign n7400 = ~n2923 & n3776 ;
  assign n7393 = ~n2777 & n4269 ;
  assign n7399 = n2918 & n4371 ;
  assign n7406 = ~n7393 & ~n7399 ;
  assign n7407 = ~n7400 & n7406 ;
  assign n7408 = ~n7405 & n7407 ;
  assign n7409 = ~n7398 & n7408 ;
  assign n7410 = ~n7392 & n7409 ;
  assign n7411 = n2453 & ~n7410 ;
  assign n7412 = \P3_rEIP_reg[22]/NET0131  & n4412 ;
  assign n7413 = \P3_InstAddrPointer_reg[22]/NET0131  & ~n4418 ;
  assign n7414 = ~n7412 & ~n7413 ;
  assign n7415 = ~n7411 & n7414 ;
  assign n7418 = \P2_InstAddrPointer_reg[15]/NET0131  & n1897 ;
  assign n7459 = ~\P2_InstAddrPointer_reg[15]/NET0131  & ~n6500 ;
  assign n7460 = \P2_InstAddrPointer_reg[15]/NET0131  & n6500 ;
  assign n7461 = ~n7459 & ~n7460 ;
  assign n7462 = n6463 & n6643 ;
  assign n7438 = ~\P2_InstAddrPointer_reg[11]/NET0131  & ~n6471 ;
  assign n7439 = ~n6497 & ~n7438 ;
  assign n7463 = n6499 & n7439 ;
  assign n7464 = n7462 & n7463 ;
  assign n7465 = ~n7461 & ~n7464 ;
  assign n7442 = ~n6616 & n6625 ;
  assign n7443 = n6612 & ~n6623 ;
  assign n7444 = ~n6629 & ~n7443 ;
  assign n7445 = ~n7442 & n7444 ;
  assign n7446 = ~n6609 & ~n6620 ;
  assign n7447 = ~n7445 & n7446 ;
  assign n7448 = ~n6609 & n6628 ;
  assign n7449 = ~n6637 & ~n7448 ;
  assign n7450 = ~n7447 & n7449 ;
  assign n7451 = ~n6601 & ~n6606 ;
  assign n7452 = ~n7450 & n7451 ;
  assign n7453 = ~n6635 & ~n6636 ;
  assign n7454 = ~n6601 & ~n7453 ;
  assign n7455 = ~n7452 & ~n7454 ;
  assign n7440 = n6498 & n7439 ;
  assign n7441 = n6463 & n6603 ;
  assign n7456 = n7440 & n7441 ;
  assign n7457 = ~n7455 & n7456 ;
  assign n7458 = n6651 & n7457 ;
  assign n7466 = n6188 & ~n7458 ;
  assign n7467 = ~n7465 & n7466 ;
  assign n7419 = n6371 & n6442 ;
  assign n7420 = n6302 & ~n6440 ;
  assign n7421 = ~n6446 & ~n7420 ;
  assign n7422 = ~n7419 & n7421 ;
  assign n7423 = ~n6406 & ~n7422 ;
  assign n7424 = ~n6445 & ~n6452 ;
  assign n7425 = ~n7423 & n7424 ;
  assign n7426 = n6268 & ~n7425 ;
  assign n7427 = ~n6198 & n6451 ;
  assign n7428 = ~n6456 & ~n7427 ;
  assign n7429 = ~n7426 & n7428 ;
  assign n7430 = ~n6459 & n7429 ;
  assign n7431 = n6483 & n7430 ;
  assign n7432 = ~n6477 & ~n6518 ;
  assign n7433 = ~n6485 & ~n6502 ;
  assign n7434 = n7432 & n7433 ;
  assign n7435 = ~n6188 & n7434 ;
  assign n7436 = n7431 & n7435 ;
  assign n7437 = ~n6506 & n7436 ;
  assign n7468 = n6267 & ~n6449 ;
  assign n7469 = n6454 & ~n7468 ;
  assign n7470 = ~n6198 & ~n7469 ;
  assign n7471 = n6460 & n6483 ;
  assign n7472 = ~n7470 & n7471 ;
  assign n7473 = n7434 & n7472 ;
  assign n7474 = ~n6188 & n6506 ;
  assign n7475 = ~n7473 & n7474 ;
  assign n7476 = ~n7437 & ~n7475 ;
  assign n7477 = ~n7467 & n7476 ;
  assign n7478 = ~n1897 & ~n7477 ;
  assign n7479 = ~n7418 & ~n7478 ;
  assign n7480 = n1734 & ~n7479 ;
  assign n7482 = ~\P2_InstAddrPointer_reg[15]/NET0131  & ~n6750 ;
  assign n7483 = ~n6753 & ~n7482 ;
  assign n7484 = n6463 & n6737 ;
  assign n7485 = ~n6732 & n7484 ;
  assign n7486 = ~\P2_InstAddrPointer_reg[13]/NET0131  & ~n6747 ;
  assign n7487 = ~n6748 & ~n7486 ;
  assign n7488 = \P2_InstAddrPointer_reg[14]/NET0131  & n7487 ;
  assign n7489 = ~\P2_InstAddrPointer_reg[11]/NET0131  & ~n6742 ;
  assign n7490 = \P2_InstAddrPointer_reg[11]/NET0131  & n6742 ;
  assign n7491 = ~n7489 & ~n7490 ;
  assign n7492 = \P2_InstAddrPointer_reg[12]/NET0131  & n7491 ;
  assign n7493 = n7488 & n7492 ;
  assign n7494 = n7485 & n7493 ;
  assign n7496 = n7483 & n7494 ;
  assign n7495 = ~n7483 & ~n7494 ;
  assign n7497 = n1890 & ~n7495 ;
  assign n7498 = ~n7496 & n7497 ;
  assign n7499 = ~n1727 & ~n6750 ;
  assign n7500 = ~n1853 & n1903 ;
  assign n7501 = n1894 & n7500 ;
  assign n7502 = ~n7499 & n7501 ;
  assign n7503 = \P2_InstAddrPointer_reg[15]/NET0131  & ~n7502 ;
  assign n7504 = ~n1771 & n6506 ;
  assign n7481 = ~n1831 & n7461 ;
  assign n7505 = n1870 & n7483 ;
  assign n7506 = ~n7481 & ~n7505 ;
  assign n7507 = ~n7504 & n7506 ;
  assign n7508 = ~n7503 & n7507 ;
  assign n7509 = ~n7498 & n7508 ;
  assign n7510 = ~n7480 & n7509 ;
  assign n7511 = n1927 & ~n7510 ;
  assign n7416 = \P2_rEIP_reg[15]/NET0131  & n3113 ;
  assign n7417 = \P2_InstAddrPointer_reg[15]/NET0131  & ~n6810 ;
  assign n7512 = ~n7416 & ~n7417 ;
  assign n7513 = ~n7511 & n7512 ;
  assign n7514 = \P2_InstAddrPointer_reg[22]/NET0131  & n1897 ;
  assign n7515 = n6487 & n7430 ;
  assign n7516 = n6519 & n7515 ;
  assign n7517 = n6541 & n7516 ;
  assign n7519 = ~n6546 & n7517 ;
  assign n7520 = n6550 & ~n7519 ;
  assign n7518 = n6551 & n7517 ;
  assign n7521 = ~n6188 & ~n7518 ;
  assign n7522 = ~n7520 & n7521 ;
  assign n7523 = n6529 & n6650 ;
  assign n7524 = n6664 & n7523 ;
  assign n7525 = n7457 & n7524 ;
  assign n7526 = \P2_InstAddrPointer_reg[21]/NET0131  & n6666 ;
  assign n7527 = n7525 & n7526 ;
  assign n7529 = n6597 & ~n7527 ;
  assign n7528 = ~n6597 & n7527 ;
  assign n7530 = n6188 & ~n7528 ;
  assign n7531 = ~n7529 & n7530 ;
  assign n7532 = ~n1897 & ~n7531 ;
  assign n7533 = ~n7522 & n7532 ;
  assign n7534 = ~n7514 & ~n7533 ;
  assign n7535 = n1734 & ~n7534 ;
  assign n7536 = ~\P2_InstAddrPointer_reg[18]/NET0131  & ~n6756 ;
  assign n7537 = \P2_InstAddrPointer_reg[18]/NET0131  & n6756 ;
  assign n7538 = ~n7536 & ~n7537 ;
  assign n7539 = ~n6719 & ~n6722 ;
  assign n7540 = n6711 & ~n7539 ;
  assign n7541 = ~n6721 & ~n6728 ;
  assign n7542 = ~n7540 & n7541 ;
  assign n7543 = n6704 & ~n7542 ;
  assign n7544 = ~n6697 & ~n6727 ;
  assign n7545 = ~n7543 & n7544 ;
  assign n7546 = n6738 & ~n7545 ;
  assign n7547 = n6745 & n7546 ;
  assign n7548 = \P2_InstAddrPointer_reg[17]/NET0131  & n6752 ;
  assign n7549 = n7547 & n7548 ;
  assign n7550 = n7538 & n7549 ;
  assign n7551 = ~\P2_InstAddrPointer_reg[19]/NET0131  & ~n7537 ;
  assign n7552 = ~n6762 & ~n7551 ;
  assign n7555 = n6544 & n7552 ;
  assign n7556 = n7550 & n7555 ;
  assign n7557 = ~n6770 & ~n7556 ;
  assign n7553 = n6548 & n7552 ;
  assign n7554 = n7550 & n7553 ;
  assign n7558 = n1890 & ~n7554 ;
  assign n7559 = ~n7557 & n7558 ;
  assign n7561 = \P2_InstAddrPointer_reg[22]/NET0131  & n1805 ;
  assign n7562 = ~n1805 & n6597 ;
  assign n7563 = ~n7561 & ~n7562 ;
  assign n7564 = ~n1804 & ~n7563 ;
  assign n7565 = \P2_InstAddrPointer_reg[22]/NET0131  & ~n1820 ;
  assign n7566 = ~n1819 & n7562 ;
  assign n7567 = ~n7565 & ~n7566 ;
  assign n7568 = ~n1814 & ~n7567 ;
  assign n7569 = ~n7564 & ~n7568 ;
  assign n7570 = ~n1810 & ~n7569 ;
  assign n7571 = n1870 & n6770 ;
  assign n7560 = ~n1771 & n6550 ;
  assign n7572 = \P2_InstAddrPointer_reg[22]/NET0131  & ~n7500 ;
  assign n7573 = n1739 & n6597 ;
  assign n7574 = ~n7572 & ~n7573 ;
  assign n7575 = ~n7560 & n7574 ;
  assign n7576 = ~n7571 & n7575 ;
  assign n7577 = ~n7570 & n7576 ;
  assign n7578 = ~n7559 & n7577 ;
  assign n7579 = ~n7535 & n7578 ;
  assign n7580 = n1927 & ~n7579 ;
  assign n7581 = \P2_rEIP_reg[22]/NET0131  & n3113 ;
  assign n7582 = \P2_InstAddrPointer_reg[22]/NET0131  & ~n6810 ;
  assign n7583 = ~n7581 & ~n7582 ;
  assign n7584 = ~n7580 & n7583 ;
  assign n7585 = \P2_InstAddrPointer_reg[26]/NET0131  & n1897 ;
  assign n7586 = ~\P2_InstAddrPointer_reg[26]/NET0131  & ~n6564 ;
  assign n7587 = ~n6567 & ~n7586 ;
  assign n7588 = n6671 & n6673 ;
  assign n7589 = ~n7587 & ~n7588 ;
  assign n7590 = n6663 & n7440 ;
  assign n7591 = n7523 & n7590 ;
  assign n7592 = n7462 & n7591 ;
  assign n7593 = ~\P2_InstAddrPointer_reg[19]/NET0131  & ~n6661 ;
  assign n7594 = ~n6532 & ~n7593 ;
  assign n7595 = n6544 & n7594 ;
  assign n7596 = n6598 & n7595 ;
  assign n7597 = n6674 & n7596 ;
  assign n7598 = n7592 & n7597 ;
  assign n7599 = n6188 & ~n7598 ;
  assign n7600 = ~n7589 & n7599 ;
  assign n7601 = ~n6459 & n6486 ;
  assign n7602 = n7429 & n7601 ;
  assign n7603 = n7432 & n7602 ;
  assign n7604 = n6516 & ~n6571 ;
  assign n7605 = n6541 & n7604 ;
  assign n7606 = n6562 & n7605 ;
  assign n7607 = n7603 & n7606 ;
  assign n7608 = ~n6569 & n7607 ;
  assign n7609 = n6569 & ~n7607 ;
  assign n7610 = ~n7608 & ~n7609 ;
  assign n7611 = ~n6188 & ~n7610 ;
  assign n7612 = ~n7600 & ~n7611 ;
  assign n7613 = ~n1897 & ~n7612 ;
  assign n7614 = ~n7585 & ~n7613 ;
  assign n7615 = n1734 & ~n7614 ;
  assign n7616 = ~\P2_InstAddrPointer_reg[26]/NET0131  & ~n6774 ;
  assign n7617 = ~n6775 & ~n7616 ;
  assign n7618 = \P2_InstAddrPointer_reg[25]/NET0131  & n6771 ;
  assign n7619 = n7556 & n7618 ;
  assign n7620 = ~n7617 & ~n7619 ;
  assign n7621 = \P2_InstAddrPointer_reg[23]/NET0131  & n6769 ;
  assign n7622 = ~\P2_InstAddrPointer_reg[23]/NET0131  & ~n6769 ;
  assign n7623 = ~n7621 & ~n7622 ;
  assign n7624 = ~\P2_InstAddrPointer_reg[24]/NET0131  & ~n7621 ;
  assign n7625 = ~n6773 & ~n7624 ;
  assign n7626 = n6782 & n7625 ;
  assign n7627 = n7623 & n7626 ;
  assign n7628 = n7554 & n7627 ;
  assign n7629 = n1890 & ~n7628 ;
  assign n7630 = ~n7620 & n7629 ;
  assign n7633 = n1798 & ~n7617 ;
  assign n7632 = ~\P2_InstAddrPointer_reg[26]/NET0131  & ~n1798 ;
  assign n7634 = ~n1727 & ~n7632 ;
  assign n7635 = ~n7633 & n7634 ;
  assign n7644 = ~n1805 & ~n7587 ;
  assign n7643 = ~\P2_InstAddrPointer_reg[26]/NET0131  & n1805 ;
  assign n7645 = n1845 & ~n7643 ;
  assign n7646 = ~n7644 & n7645 ;
  assign n7631 = ~n1771 & n6569 ;
  assign n7636 = ~n1853 & ~n1902 ;
  assign n7637 = ~n1893 & n7636 ;
  assign n7638 = \P2_InstAddrPointer_reg[26]/NET0131  & ~n7637 ;
  assign n7639 = ~n1810 & ~n1814 ;
  assign n7640 = ~n6564 & n7639 ;
  assign n7641 = ~n1739 & ~n7640 ;
  assign n7642 = n7587 & ~n7641 ;
  assign n7647 = ~n7638 & ~n7642 ;
  assign n7648 = ~n7631 & n7647 ;
  assign n7649 = ~n7646 & n7648 ;
  assign n7650 = ~n7635 & n7649 ;
  assign n7651 = ~n7630 & n7650 ;
  assign n7652 = ~n7615 & n7651 ;
  assign n7653 = n1927 & ~n7652 ;
  assign n7654 = \P2_rEIP_reg[26]/NET0131  & n3113 ;
  assign n7655 = \P2_InstAddrPointer_reg[26]/NET0131  & ~n6810 ;
  assign n7656 = ~n7654 & ~n7655 ;
  assign n7657 = ~n7653 & n7656 ;
  assign n7661 = \P1_InstAddrPointer_reg[20]/NET0131  & n2375 ;
  assign n7665 = n4928 & ~n7278 ;
  assign n7666 = ~n4453 & ~n7279 ;
  assign n7667 = ~n7665 & n7666 ;
  assign n7662 = ~n6834 & ~n6836 ;
  assign n7663 = ~n5975 & ~n7662 ;
  assign n7664 = n4453 & ~n7663 ;
  assign n7668 = ~n2375 & ~n7664 ;
  assign n7669 = ~n7667 & n7668 ;
  assign n7670 = ~n7661 & ~n7669 ;
  assign n7671 = n2244 & ~n7670 ;
  assign n7673 = n5992 & n7301 ;
  assign n7672 = ~n5992 & ~n7301 ;
  assign n7674 = n2385 & ~n7672 ;
  assign n7675 = ~n7673 & n7674 ;
  assign n7676 = n2387 & ~n6836 ;
  assign n7677 = n7308 & ~n7676 ;
  assign n7678 = n6026 & ~n7677 ;
  assign n7679 = \P1_InstAddrPointer_reg[20]/NET0131  & ~n7678 ;
  assign n7685 = ~n2337 & n4972 ;
  assign n7686 = ~n2332 & ~n7685 ;
  assign n7687 = n5992 & n7686 ;
  assign n7660 = ~n2271 & n4928 ;
  assign n7680 = n2237 & n6836 ;
  assign n7681 = ~\P1_InstAddrPointer_reg[20]/NET0131  & n2317 ;
  assign n7682 = ~n2317 & ~n6836 ;
  assign n7683 = ~n7681 & ~n7682 ;
  assign n7684 = ~n2314 & n7683 ;
  assign n7688 = ~n7680 & ~n7684 ;
  assign n7689 = ~n7660 & n7688 ;
  assign n7690 = ~n7687 & n7689 ;
  assign n7691 = ~n7679 & n7690 ;
  assign n7692 = ~n7675 & n7691 ;
  assign n7693 = ~n7671 & n7692 ;
  assign n7694 = n2432 & ~n7693 ;
  assign n7658 = \P1_rEIP_reg[20]/NET0131  & n5092 ;
  assign n7659 = \P1_InstAddrPointer_reg[20]/NET0131  & ~n5098 ;
  assign n7695 = ~n7658 & ~n7659 ;
  assign n7696 = ~n7694 & n7695 ;
  assign n7697 = ~n2436 & ~n5095 ;
  assign n7698 = ~n5108 & ~n5167 ;
  assign n7699 = \P1_InstQueue_reg[11][3]/NET0131  & ~n5104 ;
  assign n7700 = ~n5107 & n7699 ;
  assign n7701 = ~n7698 & ~n7700 ;
  assign n7702 = ~n7697 & ~n7701 ;
  assign n7703 = n2436 & n5153 ;
  assign n7704 = ~n7702 & ~n7703 ;
  assign n7709 = ~n5260 & n5263 ;
  assign n7710 = ~n5264 & ~n7709 ;
  assign n7711 = n5148 & n7710 ;
  assign n7705 = n5230 & ~n5275 ;
  assign n7706 = ~n5276 & ~n7705 ;
  assign n7707 = ~n5148 & n7706 ;
  assign n7708 = n5095 & ~n7701 ;
  assign n7712 = n5153 & ~n7708 ;
  assign n7713 = ~n7707 & n7712 ;
  assign n7714 = ~n7711 & n7713 ;
  assign n7715 = ~n7704 & ~n7714 ;
  assign n7716 = \P1_InstQueue_reg[11][3]/NET0131  & ~n5291 ;
  assign n7717 = ~n2061 & n5104 ;
  assign n7718 = ~n7699 & ~n7717 ;
  assign n7719 = n3042 & ~n7718 ;
  assign n7720 = ~n7716 & ~n7719 ;
  assign n7721 = ~n7715 & n7720 ;
  assign n7730 = \buf2_reg[30]/NET0131  & ~n3079 ;
  assign n7731 = \buf1_reg[30]/NET0131  & n3079 ;
  assign n7732 = ~n7730 & ~n7731 ;
  assign n7733 = n3091 & ~n7732 ;
  assign n7734 = \buf2_reg[22]/NET0131  & ~n3079 ;
  assign n7735 = \buf1_reg[22]/NET0131  & n3079 ;
  assign n7736 = ~n7734 & ~n7735 ;
  assign n7737 = n3098 & ~n7736 ;
  assign n7738 = ~n7733 & ~n7737 ;
  assign n7739 = \P2_DataWidth_reg[1]/NET0131  & ~n7738 ;
  assign n7722 = \buf2_reg[6]/NET0131  & ~n3079 ;
  assign n7723 = \buf1_reg[6]/NET0131  & n3079 ;
  assign n7724 = ~n7722 & ~n7723 ;
  assign n7725 = ~n3050 & ~n7724 ;
  assign n7726 = \P2_InstQueue_reg[11][6]/NET0131  & ~n3049 ;
  assign n7727 = ~n3046 & n7726 ;
  assign n7728 = ~n7725 & ~n7727 ;
  assign n7740 = ~n3106 & ~n7728 ;
  assign n7741 = ~n7739 & ~n7740 ;
  assign n7742 = n1931 & ~n7741 ;
  assign n7729 = n3087 & ~n7728 ;
  assign n7743 = ~n1625 & n3049 ;
  assign n7744 = ~n7726 & ~n7743 ;
  assign n7745 = n3040 & ~n7744 ;
  assign n7746 = \P2_InstQueue_reg[11][6]/NET0131  & ~n3118 ;
  assign n7747 = ~n7745 & ~n7746 ;
  assign n7748 = ~n7729 & n7747 ;
  assign n7749 = ~n7742 & n7748 ;
  assign n7750 = ~n5167 & ~n5327 ;
  assign n7751 = \P1_InstQueue_reg[0][3]/NET0131  & ~n5324 ;
  assign n7752 = ~n5326 & n7751 ;
  assign n7753 = ~n7750 & ~n7752 ;
  assign n7754 = ~n7697 & ~n7753 ;
  assign n7755 = n2436 & n5338 ;
  assign n7756 = ~n7754 & ~n7755 ;
  assign n7759 = n5334 & n7710 ;
  assign n7757 = ~n5334 & n7706 ;
  assign n7758 = n5095 & ~n7753 ;
  assign n7760 = n5338 & ~n7758 ;
  assign n7761 = ~n7757 & n7760 ;
  assign n7762 = ~n7759 & n7761 ;
  assign n7763 = ~n7756 & ~n7762 ;
  assign n7764 = \P1_InstQueue_reg[0][3]/NET0131  & ~n5291 ;
  assign n7765 = ~n2061 & n5324 ;
  assign n7766 = ~n7751 & ~n7765 ;
  assign n7767 = n3042 & ~n7766 ;
  assign n7768 = ~n7764 & ~n7767 ;
  assign n7769 = ~n7763 & n7768 ;
  assign n7770 = ~n5167 & ~n5353 ;
  assign n7771 = \P1_InstQueue_reg[10][3]/NET0131  & ~n5107 ;
  assign n7772 = ~n5151 & n7771 ;
  assign n7773 = ~n7770 & ~n7772 ;
  assign n7774 = ~n7697 & ~n7773 ;
  assign n7775 = n2436 & n5361 ;
  assign n7776 = ~n7774 & ~n7775 ;
  assign n7779 = n5359 & n7710 ;
  assign n7777 = ~n5359 & n7706 ;
  assign n7778 = n5095 & ~n7773 ;
  assign n7780 = n5361 & ~n7778 ;
  assign n7781 = ~n7777 & n7780 ;
  assign n7782 = ~n7779 & n7781 ;
  assign n7783 = ~n7776 & ~n7782 ;
  assign n7784 = \P1_InstQueue_reg[10][3]/NET0131  & ~n5291 ;
  assign n7785 = ~n2061 & n5107 ;
  assign n7786 = ~n7771 & ~n7785 ;
  assign n7787 = n3042 & ~n7786 ;
  assign n7788 = ~n7784 & ~n7787 ;
  assign n7789 = ~n7783 & n7788 ;
  assign n7790 = ~n5167 & ~n5378 ;
  assign n7791 = \P1_InstQueue_reg[12][3]/NET0131  & ~n5377 ;
  assign n7792 = ~n5104 & n7791 ;
  assign n7793 = ~n7790 & ~n7792 ;
  assign n7794 = ~n7697 & ~n7793 ;
  assign n7795 = n2436 & n5384 ;
  assign n7796 = ~n7794 & ~n7795 ;
  assign n7799 = n5151 & n7710 ;
  assign n7797 = ~n5151 & n7706 ;
  assign n7798 = n5095 & ~n7793 ;
  assign n7800 = n5384 & ~n7798 ;
  assign n7801 = ~n7797 & n7800 ;
  assign n7802 = ~n7799 & n7801 ;
  assign n7803 = ~n7796 & ~n7802 ;
  assign n7804 = \P1_InstQueue_reg[12][3]/NET0131  & ~n5291 ;
  assign n7805 = ~n2061 & n5377 ;
  assign n7806 = ~n7791 & ~n7805 ;
  assign n7807 = n3042 & ~n7806 ;
  assign n7808 = ~n7804 & ~n7807 ;
  assign n7809 = ~n7803 & n7808 ;
  assign n7810 = ~n5167 & ~n5399 ;
  assign n7811 = \P1_InstQueue_reg[13][3]/NET0131  & ~n5334 ;
  assign n7812 = ~n5377 & n7811 ;
  assign n7813 = ~n7810 & ~n7812 ;
  assign n7814 = ~n7697 & ~n7813 ;
  assign n7815 = n2436 & n5405 ;
  assign n7816 = ~n7814 & ~n7815 ;
  assign n7819 = n5107 & n7710 ;
  assign n7817 = ~n5107 & n7706 ;
  assign n7818 = n5095 & ~n7813 ;
  assign n7820 = n5405 & ~n7818 ;
  assign n7821 = ~n7817 & n7820 ;
  assign n7822 = ~n7819 & n7821 ;
  assign n7823 = ~n7816 & ~n7822 ;
  assign n7824 = \P1_InstQueue_reg[13][3]/NET0131  & ~n5291 ;
  assign n7825 = ~n2061 & n5334 ;
  assign n7826 = ~n7811 & ~n7825 ;
  assign n7827 = n3042 & ~n7826 ;
  assign n7828 = ~n7824 & ~n7827 ;
  assign n7829 = ~n7823 & n7828 ;
  assign n7830 = ~n5167 & ~n5337 ;
  assign n7831 = \P1_InstQueue_reg[14][3]/NET0131  & ~n5336 ;
  assign n7832 = ~n5334 & n7831 ;
  assign n7833 = ~n7830 & ~n7832 ;
  assign n7834 = ~n7697 & ~n7833 ;
  assign n7835 = n2436 & n5425 ;
  assign n7836 = ~n7834 & ~n7835 ;
  assign n7839 = n5104 & n7710 ;
  assign n7837 = ~n5104 & n7706 ;
  assign n7838 = n5095 & ~n7833 ;
  assign n7840 = n5425 & ~n7838 ;
  assign n7841 = ~n7837 & n7840 ;
  assign n7842 = ~n7839 & n7841 ;
  assign n7843 = ~n7836 & ~n7842 ;
  assign n7844 = \P1_InstQueue_reg[14][3]/NET0131  & ~n5291 ;
  assign n7845 = ~n2061 & n5336 ;
  assign n7846 = ~n7831 & ~n7845 ;
  assign n7847 = n3042 & ~n7846 ;
  assign n7848 = ~n7844 & ~n7847 ;
  assign n7849 = ~n7843 & n7848 ;
  assign n7850 = ~n5167 & ~n5440 ;
  assign n7851 = \P1_InstQueue_reg[15][3]/NET0131  & ~n5326 ;
  assign n7852 = ~n5336 & n7851 ;
  assign n7853 = ~n7850 & ~n7852 ;
  assign n7854 = ~n7697 & ~n7853 ;
  assign n7855 = n2436 & n5446 ;
  assign n7856 = ~n7854 & ~n7855 ;
  assign n7859 = n5377 & n7710 ;
  assign n7857 = ~n5377 & n7706 ;
  assign n7858 = n5095 & ~n7853 ;
  assign n7860 = n5446 & ~n7858 ;
  assign n7861 = ~n7857 & n7860 ;
  assign n7862 = ~n7859 & n7861 ;
  assign n7863 = ~n7856 & ~n7862 ;
  assign n7864 = \P1_InstQueue_reg[15][3]/NET0131  & ~n5291 ;
  assign n7865 = ~n2061 & n5326 ;
  assign n7866 = ~n7851 & ~n7865 ;
  assign n7867 = n3042 & ~n7866 ;
  assign n7868 = ~n7864 & ~n7867 ;
  assign n7869 = ~n7863 & n7868 ;
  assign n7870 = ~n5167 & ~n5462 ;
  assign n7871 = \P1_InstQueue_reg[1][3]/NET0131  & ~n5461 ;
  assign n7872 = ~n5324 & n7871 ;
  assign n7873 = ~n7870 & ~n7872 ;
  assign n7874 = ~n7697 & ~n7873 ;
  assign n7875 = n2436 & n5468 ;
  assign n7876 = ~n7874 & ~n7875 ;
  assign n7879 = n5336 & n7710 ;
  assign n7877 = ~n5336 & n7706 ;
  assign n7878 = n5095 & ~n7873 ;
  assign n7880 = n5468 & ~n7878 ;
  assign n7881 = ~n7877 & n7880 ;
  assign n7882 = ~n7879 & n7881 ;
  assign n7883 = ~n7876 & ~n7882 ;
  assign n7884 = \P1_InstQueue_reg[1][3]/NET0131  & ~n5291 ;
  assign n7885 = ~n2061 & n5461 ;
  assign n7886 = ~n7871 & ~n7885 ;
  assign n7887 = n3042 & ~n7886 ;
  assign n7888 = ~n7884 & ~n7887 ;
  assign n7889 = ~n7883 & n7888 ;
  assign n7890 = ~n5167 & ~n5506 ;
  assign n7891 = \P1_InstQueue_reg[2][3]/NET0131  & ~n5484 ;
  assign n7892 = ~n5461 & n7891 ;
  assign n7893 = ~n7890 & ~n7892 ;
  assign n7894 = ~n7697 & ~n7893 ;
  assign n7895 = n2436 & n5512 ;
  assign n7896 = ~n7894 & ~n7895 ;
  assign n7899 = n5326 & n7710 ;
  assign n7897 = ~n5326 & n7706 ;
  assign n7898 = n5095 & ~n7893 ;
  assign n7900 = n5512 & ~n7898 ;
  assign n7901 = ~n7897 & n7900 ;
  assign n7902 = ~n7899 & n7901 ;
  assign n7903 = ~n7896 & ~n7902 ;
  assign n7904 = \P1_InstQueue_reg[2][3]/NET0131  & ~n5291 ;
  assign n7905 = ~n2061 & n5484 ;
  assign n7906 = ~n7891 & ~n7905 ;
  assign n7907 = n3042 & ~n7906 ;
  assign n7908 = ~n7904 & ~n7907 ;
  assign n7909 = ~n7903 & n7908 ;
  assign n7910 = ~n5167 & ~n5485 ;
  assign n7911 = \P1_InstQueue_reg[3][3]/NET0131  & ~n5483 ;
  assign n7912 = ~n5484 & n7911 ;
  assign n7913 = ~n7910 & ~n7912 ;
  assign n7914 = ~n7697 & ~n7913 ;
  assign n7915 = n2436 & n5491 ;
  assign n7916 = ~n7914 & ~n7915 ;
  assign n7919 = n5324 & n7710 ;
  assign n7917 = ~n5324 & n7706 ;
  assign n7918 = n5095 & ~n7913 ;
  assign n7920 = n5491 & ~n7918 ;
  assign n7921 = ~n7917 & n7920 ;
  assign n7922 = ~n7919 & n7921 ;
  assign n7923 = ~n7916 & ~n7922 ;
  assign n7924 = \P1_InstQueue_reg[3][3]/NET0131  & ~n5291 ;
  assign n7925 = ~n2061 & n5483 ;
  assign n7926 = ~n7911 & ~n7925 ;
  assign n7927 = n3042 & ~n7926 ;
  assign n7928 = ~n7924 & ~n7927 ;
  assign n7929 = ~n7923 & n7928 ;
  assign n7930 = ~n5167 & ~n5528 ;
  assign n7931 = \P1_InstQueue_reg[4][3]/NET0131  & ~n5527 ;
  assign n7932 = ~n5483 & n7931 ;
  assign n7933 = ~n7930 & ~n7932 ;
  assign n7934 = ~n7697 & ~n7933 ;
  assign n7935 = n2436 & n5534 ;
  assign n7936 = ~n7934 & ~n7935 ;
  assign n7939 = n5461 & n7710 ;
  assign n7937 = ~n5461 & n7706 ;
  assign n7938 = n5095 & ~n7933 ;
  assign n7940 = n5534 & ~n7938 ;
  assign n7941 = ~n7937 & n7940 ;
  assign n7942 = ~n7939 & n7941 ;
  assign n7943 = ~n7936 & ~n7942 ;
  assign n7944 = \P1_InstQueue_reg[4][3]/NET0131  & ~n5291 ;
  assign n7945 = ~n2061 & n5527 ;
  assign n7946 = ~n7931 & ~n7945 ;
  assign n7947 = n3042 & ~n7946 ;
  assign n7948 = ~n7944 & ~n7947 ;
  assign n7949 = ~n7943 & n7948 ;
  assign n7950 = ~n5167 & ~n5550 ;
  assign n7951 = \P1_InstQueue_reg[5][3]/NET0131  & ~n5549 ;
  assign n7952 = ~n5527 & n7951 ;
  assign n7953 = ~n7950 & ~n7952 ;
  assign n7954 = ~n7697 & ~n7953 ;
  assign n7955 = n2436 & n5556 ;
  assign n7956 = ~n7954 & ~n7955 ;
  assign n7959 = n5484 & n7710 ;
  assign n7957 = ~n5484 & n7706 ;
  assign n7958 = n5095 & ~n7953 ;
  assign n7960 = n5556 & ~n7958 ;
  assign n7961 = ~n7957 & n7960 ;
  assign n7962 = ~n7959 & n7961 ;
  assign n7963 = ~n7956 & ~n7962 ;
  assign n7964 = \P1_InstQueue_reg[5][3]/NET0131  & ~n5291 ;
  assign n7965 = ~n2061 & n5549 ;
  assign n7966 = ~n7951 & ~n7965 ;
  assign n7967 = n3042 & ~n7966 ;
  assign n7968 = ~n7964 & ~n7967 ;
  assign n7969 = ~n7963 & n7968 ;
  assign n7970 = ~n5167 & ~n5572 ;
  assign n7971 = \P1_InstQueue_reg[6][3]/NET0131  & ~n5571 ;
  assign n7972 = ~n5549 & n7971 ;
  assign n7973 = ~n7970 & ~n7972 ;
  assign n7974 = ~n7697 & ~n7973 ;
  assign n7975 = n2436 & n5578 ;
  assign n7976 = ~n7974 & ~n7975 ;
  assign n7979 = n5483 & n7710 ;
  assign n7977 = ~n5483 & n7706 ;
  assign n7978 = n5095 & ~n7973 ;
  assign n7980 = n5578 & ~n7978 ;
  assign n7981 = ~n7977 & n7980 ;
  assign n7982 = ~n7979 & n7981 ;
  assign n7983 = ~n7976 & ~n7982 ;
  assign n7984 = \P1_InstQueue_reg[6][3]/NET0131  & ~n5291 ;
  assign n7985 = ~n2061 & n5571 ;
  assign n7986 = ~n7971 & ~n7985 ;
  assign n7987 = n3042 & ~n7986 ;
  assign n7988 = ~n7984 & ~n7987 ;
  assign n7989 = ~n7983 & n7988 ;
  assign n7990 = ~n5167 & ~n5593 ;
  assign n7991 = \P1_InstQueue_reg[7][3]/NET0131  & ~n5359 ;
  assign n7992 = ~n5571 & n7991 ;
  assign n7993 = ~n7990 & ~n7992 ;
  assign n7994 = ~n7697 & ~n7993 ;
  assign n7995 = n2436 & n5599 ;
  assign n7996 = ~n7994 & ~n7995 ;
  assign n7999 = n5527 & n7710 ;
  assign n7997 = ~n5527 & n7706 ;
  assign n7998 = n5095 & ~n7993 ;
  assign n8000 = n5599 & ~n7998 ;
  assign n8001 = ~n7997 & n8000 ;
  assign n8002 = ~n7999 & n8001 ;
  assign n8003 = ~n7996 & ~n8002 ;
  assign n8004 = \P1_InstQueue_reg[7][3]/NET0131  & ~n5291 ;
  assign n8005 = ~n2061 & n5359 ;
  assign n8006 = ~n7991 & ~n8005 ;
  assign n8007 = n3042 & ~n8006 ;
  assign n8008 = ~n8004 & ~n8007 ;
  assign n8009 = ~n8003 & n8008 ;
  assign n8010 = ~n5167 & ~n5360 ;
  assign n8011 = \P1_InstQueue_reg[8][3]/NET0131  & ~n5148 ;
  assign n8012 = ~n5359 & n8011 ;
  assign n8013 = ~n8010 & ~n8012 ;
  assign n8014 = ~n7697 & ~n8013 ;
  assign n8015 = n2436 & n5619 ;
  assign n8016 = ~n8014 & ~n8015 ;
  assign n8019 = n5549 & n7710 ;
  assign n8017 = ~n5549 & n7706 ;
  assign n8018 = n5095 & ~n8013 ;
  assign n8020 = n5619 & ~n8018 ;
  assign n8021 = ~n8017 & n8020 ;
  assign n8022 = ~n8019 & n8021 ;
  assign n8023 = ~n8016 & ~n8022 ;
  assign n8024 = \P1_InstQueue_reg[8][3]/NET0131  & ~n5291 ;
  assign n8025 = ~n2061 & n5148 ;
  assign n8026 = ~n8011 & ~n8025 ;
  assign n8027 = n3042 & ~n8026 ;
  assign n8028 = ~n8024 & ~n8027 ;
  assign n8029 = ~n8023 & n8028 ;
  assign n8030 = ~n5152 & ~n5167 ;
  assign n8031 = \P1_InstQueue_reg[9][3]/NET0131  & ~n5151 ;
  assign n8032 = ~n5148 & n8031 ;
  assign n8033 = ~n8030 & ~n8032 ;
  assign n8034 = ~n7697 & ~n8033 ;
  assign n8035 = n2436 & n5639 ;
  assign n8036 = ~n8034 & ~n8035 ;
  assign n8039 = n5571 & n7710 ;
  assign n8037 = ~n5571 & n7706 ;
  assign n8038 = n5095 & ~n8033 ;
  assign n8040 = n5639 & ~n8038 ;
  assign n8041 = ~n8037 & n8040 ;
  assign n8042 = ~n8039 & n8041 ;
  assign n8043 = ~n8036 & ~n8042 ;
  assign n8044 = \P1_InstQueue_reg[9][3]/NET0131  & ~n5291 ;
  assign n8045 = ~n2061 & n5151 ;
  assign n8046 = ~n8031 & ~n8045 ;
  assign n8047 = n3042 & ~n8046 ;
  assign n8048 = ~n8044 & ~n8047 ;
  assign n8049 = ~n8043 & n8048 ;
  assign n8055 = n3162 & ~n7732 ;
  assign n8056 = n3165 & ~n7736 ;
  assign n8057 = ~n8055 & ~n8056 ;
  assign n8058 = \P2_DataWidth_reg[1]/NET0131  & ~n8057 ;
  assign n8050 = ~n3155 & ~n7724 ;
  assign n8051 = \P2_InstQueue_reg[0][6]/NET0131  & ~n3152 ;
  assign n8052 = ~n3154 & n8051 ;
  assign n8053 = ~n8050 & ~n8052 ;
  assign n8059 = ~n3170 & ~n8053 ;
  assign n8060 = ~n8058 & ~n8059 ;
  assign n8061 = n1931 & ~n8060 ;
  assign n8054 = n3087 & ~n8053 ;
  assign n8062 = ~n1625 & n3152 ;
  assign n8063 = ~n8051 & ~n8062 ;
  assign n8064 = n3040 & ~n8063 ;
  assign n8065 = \P2_InstQueue_reg[0][6]/NET0131  & ~n3118 ;
  assign n8066 = ~n8064 & ~n8065 ;
  assign n8067 = ~n8054 & n8066 ;
  assign n8068 = ~n8061 & n8067 ;
  assign n8074 = n3091 & ~n7736 ;
  assign n8075 = n3198 & ~n7732 ;
  assign n8076 = ~n8074 & ~n8075 ;
  assign n8077 = \P2_DataWidth_reg[1]/NET0131  & ~n8076 ;
  assign n8069 = ~n3202 & ~n7724 ;
  assign n8070 = \P2_InstQueue_reg[10][6]/NET0131  & ~n3046 ;
  assign n8071 = ~n3098 & n8070 ;
  assign n8072 = ~n8069 & ~n8071 ;
  assign n8078 = ~n3200 & ~n8072 ;
  assign n8079 = ~n8077 & ~n8078 ;
  assign n8080 = n1931 & ~n8079 ;
  assign n8073 = n3087 & ~n8072 ;
  assign n8081 = ~n1625 & n3046 ;
  assign n8082 = ~n8070 & ~n8081 ;
  assign n8083 = n3040 & ~n8082 ;
  assign n8084 = \P2_InstQueue_reg[10][6]/NET0131  & ~n3118 ;
  assign n8085 = ~n8083 & ~n8084 ;
  assign n8086 = ~n8073 & n8085 ;
  assign n8087 = ~n8080 & n8086 ;
  assign n8093 = n3098 & ~n7732 ;
  assign n8094 = n3046 & ~n7736 ;
  assign n8095 = ~n8093 & ~n8094 ;
  assign n8096 = \P2_DataWidth_reg[1]/NET0131  & ~n8095 ;
  assign n8088 = ~n3238 & ~n7724 ;
  assign n8089 = \P2_InstQueue_reg[12][6]/NET0131  & ~n3237 ;
  assign n8090 = ~n3049 & n8089 ;
  assign n8091 = ~n8088 & ~n8090 ;
  assign n8097 = ~n3248 & ~n8091 ;
  assign n8098 = ~n8096 & ~n8097 ;
  assign n8099 = n1931 & ~n8098 ;
  assign n8092 = n3087 & ~n8091 ;
  assign n8100 = ~n1625 & n3237 ;
  assign n8101 = ~n8089 & ~n8100 ;
  assign n8102 = n3040 & ~n8101 ;
  assign n8103 = \P2_InstQueue_reg[12][6]/NET0131  & ~n3118 ;
  assign n8104 = ~n8102 & ~n8103 ;
  assign n8105 = ~n8092 & n8104 ;
  assign n8106 = ~n8099 & n8105 ;
  assign n8112 = n3046 & ~n7732 ;
  assign n8113 = n3049 & ~n7736 ;
  assign n8114 = ~n8112 & ~n8113 ;
  assign n8115 = \P2_DataWidth_reg[1]/NET0131  & ~n8114 ;
  assign n8107 = ~n3275 & ~n7724 ;
  assign n8108 = \P2_InstQueue_reg[13][6]/NET0131  & ~n3162 ;
  assign n8109 = ~n3237 & n8108 ;
  assign n8110 = ~n8107 & ~n8109 ;
  assign n8116 = ~n3285 & ~n8110 ;
  assign n8117 = ~n8115 & ~n8116 ;
  assign n8118 = n1931 & ~n8117 ;
  assign n8111 = n3087 & ~n8110 ;
  assign n8119 = ~n1625 & n3162 ;
  assign n8120 = ~n8108 & ~n8119 ;
  assign n8121 = n3040 & ~n8120 ;
  assign n8122 = \P2_InstQueue_reg[13][6]/NET0131  & ~n3118 ;
  assign n8123 = ~n8121 & ~n8122 ;
  assign n8124 = ~n8111 & n8123 ;
  assign n8125 = ~n8118 & n8124 ;
  assign n8131 = n3049 & ~n7732 ;
  assign n8132 = n3237 & ~n7736 ;
  assign n8133 = ~n8131 & ~n8132 ;
  assign n8134 = \P2_DataWidth_reg[1]/NET0131  & ~n8133 ;
  assign n8126 = ~n3169 & ~n7724 ;
  assign n8127 = \P2_InstQueue_reg[14][6]/NET0131  & ~n3165 ;
  assign n8128 = ~n3162 & n8127 ;
  assign n8129 = ~n8126 & ~n8128 ;
  assign n8135 = ~n3321 & ~n8129 ;
  assign n8136 = ~n8134 & ~n8135 ;
  assign n8137 = n1931 & ~n8136 ;
  assign n8130 = n3087 & ~n8129 ;
  assign n8138 = ~n1625 & n3165 ;
  assign n8139 = ~n8127 & ~n8138 ;
  assign n8140 = n3040 & ~n8139 ;
  assign n8141 = \P2_InstQueue_reg[14][6]/NET0131  & ~n3118 ;
  assign n8142 = ~n8140 & ~n8141 ;
  assign n8143 = ~n8130 & n8142 ;
  assign n8144 = ~n8137 & n8143 ;
  assign n8150 = n3237 & ~n7732 ;
  assign n8151 = n3162 & ~n7736 ;
  assign n8152 = ~n8150 & ~n8151 ;
  assign n8153 = \P2_DataWidth_reg[1]/NET0131  & ~n8152 ;
  assign n8145 = ~n3348 & ~n7724 ;
  assign n8146 = \P2_InstQueue_reg[15][6]/NET0131  & ~n3154 ;
  assign n8147 = ~n3165 & n8146 ;
  assign n8148 = ~n8145 & ~n8147 ;
  assign n8154 = ~n3358 & ~n8148 ;
  assign n8155 = ~n8153 & ~n8154 ;
  assign n8156 = n1931 & ~n8155 ;
  assign n8149 = n3087 & ~n8148 ;
  assign n8157 = ~n1625 & n3154 ;
  assign n8158 = ~n8146 & ~n8157 ;
  assign n8159 = n3040 & ~n8158 ;
  assign n8160 = \P2_InstQueue_reg[15][6]/NET0131  & ~n3118 ;
  assign n8161 = ~n8159 & ~n8160 ;
  assign n8162 = ~n8149 & n8161 ;
  assign n8163 = ~n8156 & n8162 ;
  assign n8169 = n3165 & ~n7732 ;
  assign n8170 = n3154 & ~n7736 ;
  assign n8171 = ~n8169 & ~n8170 ;
  assign n8172 = \P2_DataWidth_reg[1]/NET0131  & ~n8171 ;
  assign n8164 = ~n3389 & ~n7724 ;
  assign n8165 = \P2_InstQueue_reg[1][6]/NET0131  & ~n3388 ;
  assign n8166 = ~n3152 & n8165 ;
  assign n8167 = ~n8164 & ~n8166 ;
  assign n8173 = ~n3386 & ~n8167 ;
  assign n8174 = ~n8172 & ~n8173 ;
  assign n8175 = n1931 & ~n8174 ;
  assign n8168 = n3087 & ~n8167 ;
  assign n8176 = ~n1625 & n3388 ;
  assign n8177 = ~n8165 & ~n8176 ;
  assign n8178 = n3040 & ~n8177 ;
  assign n8179 = \P2_InstQueue_reg[1][6]/NET0131  & ~n3118 ;
  assign n8180 = ~n8178 & ~n8179 ;
  assign n8181 = ~n8168 & n8180 ;
  assign n8182 = ~n8175 & n8181 ;
  assign n8188 = n3152 & ~n7736 ;
  assign n8189 = n3154 & ~n7732 ;
  assign n8190 = ~n8188 & ~n8189 ;
  assign n8191 = \P2_DataWidth_reg[1]/NET0131  & ~n8190 ;
  assign n8183 = ~n3424 & ~n7724 ;
  assign n8184 = \P2_InstQueue_reg[2][6]/NET0131  & ~n3423 ;
  assign n8185 = ~n3388 & n8184 ;
  assign n8186 = ~n8183 & ~n8185 ;
  assign n8192 = ~n3434 & ~n8186 ;
  assign n8193 = ~n8191 & ~n8192 ;
  assign n8194 = n1931 & ~n8193 ;
  assign n8187 = n3087 & ~n8186 ;
  assign n8195 = ~n1625 & n3423 ;
  assign n8196 = ~n8184 & ~n8195 ;
  assign n8197 = n3040 & ~n8196 ;
  assign n8198 = \P2_InstQueue_reg[2][6]/NET0131  & ~n3118 ;
  assign n8199 = ~n8197 & ~n8198 ;
  assign n8200 = ~n8187 & n8199 ;
  assign n8201 = ~n8194 & n8200 ;
  assign n8207 = n3152 & ~n7732 ;
  assign n8208 = n3388 & ~n7736 ;
  assign n8209 = ~n8207 & ~n8208 ;
  assign n8210 = \P2_DataWidth_reg[1]/NET0131  & ~n8209 ;
  assign n8202 = ~n3462 & ~n7724 ;
  assign n8203 = \P2_InstQueue_reg[3][6]/NET0131  & ~n3461 ;
  assign n8204 = ~n3423 & n8203 ;
  assign n8205 = ~n8202 & ~n8204 ;
  assign n8211 = ~n3472 & ~n8205 ;
  assign n8212 = ~n8210 & ~n8211 ;
  assign n8213 = n1931 & ~n8212 ;
  assign n8206 = n3087 & ~n8205 ;
  assign n8214 = ~n1625 & n3461 ;
  assign n8215 = ~n8203 & ~n8214 ;
  assign n8216 = n3040 & ~n8215 ;
  assign n8217 = \P2_InstQueue_reg[3][6]/NET0131  & ~n3118 ;
  assign n8218 = ~n8216 & ~n8217 ;
  assign n8219 = ~n8206 & n8218 ;
  assign n8220 = ~n8213 & n8219 ;
  assign n8226 = n3388 & ~n7732 ;
  assign n8227 = n3423 & ~n7736 ;
  assign n8228 = ~n8226 & ~n8227 ;
  assign n8229 = \P2_DataWidth_reg[1]/NET0131  & ~n8228 ;
  assign n8221 = ~n3500 & ~n7724 ;
  assign n8222 = \P2_InstQueue_reg[4][6]/NET0131  & ~n3499 ;
  assign n8223 = ~n3461 & n8222 ;
  assign n8224 = ~n8221 & ~n8223 ;
  assign n8230 = ~n3510 & ~n8224 ;
  assign n8231 = ~n8229 & ~n8230 ;
  assign n8232 = n1931 & ~n8231 ;
  assign n8225 = n3087 & ~n8224 ;
  assign n8233 = ~n1625 & n3499 ;
  assign n8234 = ~n8222 & ~n8233 ;
  assign n8235 = n3040 & ~n8234 ;
  assign n8236 = \P2_InstQueue_reg[4][6]/NET0131  & ~n3118 ;
  assign n8237 = ~n8235 & ~n8236 ;
  assign n8238 = ~n8225 & n8237 ;
  assign n8239 = ~n8232 & n8238 ;
  assign n8245 = n3423 & ~n7732 ;
  assign n8246 = n3461 & ~n7736 ;
  assign n8247 = ~n8245 & ~n8246 ;
  assign n8248 = \P2_DataWidth_reg[1]/NET0131  & ~n8247 ;
  assign n8240 = ~n3538 & ~n7724 ;
  assign n8241 = \P2_InstQueue_reg[5][6]/NET0131  & ~n3537 ;
  assign n8242 = ~n3499 & n8241 ;
  assign n8243 = ~n8240 & ~n8242 ;
  assign n8249 = ~n3548 & ~n8243 ;
  assign n8250 = ~n8248 & ~n8249 ;
  assign n8251 = n1931 & ~n8250 ;
  assign n8244 = n3087 & ~n8243 ;
  assign n8252 = ~n1625 & n3537 ;
  assign n8253 = ~n8241 & ~n8252 ;
  assign n8254 = n3040 & ~n8253 ;
  assign n8255 = \P2_InstQueue_reg[5][6]/NET0131  & ~n3118 ;
  assign n8256 = ~n8254 & ~n8255 ;
  assign n8257 = ~n8244 & n8256 ;
  assign n8258 = ~n8251 & n8257 ;
  assign n8264 = n3461 & ~n7732 ;
  assign n8265 = n3499 & ~n7736 ;
  assign n8266 = ~n8264 & ~n8265 ;
  assign n8267 = \P2_DataWidth_reg[1]/NET0131  & ~n8266 ;
  assign n8259 = ~n3576 & ~n7724 ;
  assign n8260 = \P2_InstQueue_reg[6][6]/NET0131  & ~n3575 ;
  assign n8261 = ~n3537 & n8260 ;
  assign n8262 = ~n8259 & ~n8261 ;
  assign n8268 = ~n3586 & ~n8262 ;
  assign n8269 = ~n8267 & ~n8268 ;
  assign n8270 = n1931 & ~n8269 ;
  assign n8263 = n3087 & ~n8262 ;
  assign n8271 = ~n1625 & n3575 ;
  assign n8272 = ~n8260 & ~n8271 ;
  assign n8273 = n3040 & ~n8272 ;
  assign n8274 = \P2_InstQueue_reg[6][6]/NET0131  & ~n3118 ;
  assign n8275 = ~n8273 & ~n8274 ;
  assign n8276 = ~n8263 & n8275 ;
  assign n8277 = ~n8270 & n8276 ;
  assign n8283 = n3499 & ~n7732 ;
  assign n8284 = n3537 & ~n7736 ;
  assign n8285 = ~n8283 & ~n8284 ;
  assign n8286 = \P2_DataWidth_reg[1]/NET0131  & ~n8285 ;
  assign n8278 = ~n3613 & ~n7724 ;
  assign n8279 = \P2_InstQueue_reg[7][6]/NET0131  & ~n3198 ;
  assign n8280 = ~n3575 & n8279 ;
  assign n8281 = ~n8278 & ~n8280 ;
  assign n8287 = ~n3623 & ~n8281 ;
  assign n8288 = ~n8286 & ~n8287 ;
  assign n8289 = n1931 & ~n8288 ;
  assign n8282 = n3087 & ~n8281 ;
  assign n8290 = ~n1625 & n3198 ;
  assign n8291 = ~n8279 & ~n8290 ;
  assign n8292 = n3040 & ~n8291 ;
  assign n8293 = \P2_InstQueue_reg[7][6]/NET0131  & ~n3118 ;
  assign n8294 = ~n8292 & ~n8293 ;
  assign n8295 = ~n8282 & n8294 ;
  assign n8296 = ~n8289 & n8295 ;
  assign n8302 = n3537 & ~n7732 ;
  assign n8303 = n3575 & ~n7736 ;
  assign n8304 = ~n8302 & ~n8303 ;
  assign n8305 = \P2_DataWidth_reg[1]/NET0131  & ~n8304 ;
  assign n8297 = ~n3199 & ~n7724 ;
  assign n8298 = \P2_InstQueue_reg[8][6]/NET0131  & ~n3091 ;
  assign n8299 = ~n3198 & n8298 ;
  assign n8300 = ~n8297 & ~n8299 ;
  assign n8306 = ~n3659 & ~n8300 ;
  assign n8307 = ~n8305 & ~n8306 ;
  assign n8308 = n1931 & ~n8307 ;
  assign n8301 = n3087 & ~n8300 ;
  assign n8309 = ~n1625 & n3091 ;
  assign n8310 = ~n8298 & ~n8309 ;
  assign n8311 = n3040 & ~n8310 ;
  assign n8312 = \P2_InstQueue_reg[8][6]/NET0131  & ~n3118 ;
  assign n8313 = ~n8311 & ~n8312 ;
  assign n8314 = ~n8301 & n8313 ;
  assign n8315 = ~n8308 & n8314 ;
  assign n8321 = n3575 & ~n7732 ;
  assign n8322 = n3198 & ~n7736 ;
  assign n8323 = ~n8321 & ~n8322 ;
  assign n8324 = \P2_DataWidth_reg[1]/NET0131  & ~n8323 ;
  assign n8316 = ~n3105 & ~n7724 ;
  assign n8317 = \P2_InstQueue_reg[9][6]/NET0131  & ~n3098 ;
  assign n8318 = ~n3091 & n8317 ;
  assign n8319 = ~n8316 & ~n8318 ;
  assign n8325 = ~n3695 & ~n8319 ;
  assign n8326 = ~n8324 & ~n8325 ;
  assign n8327 = n1931 & ~n8326 ;
  assign n8320 = n3087 & ~n8319 ;
  assign n8328 = ~n1625 & n3098 ;
  assign n8329 = ~n8317 & ~n8328 ;
  assign n8330 = n3040 & ~n8329 ;
  assign n8331 = \P2_InstQueue_reg[9][6]/NET0131  & ~n3118 ;
  assign n8332 = ~n8330 & ~n8331 ;
  assign n8333 = ~n8320 & n8332 ;
  assign n8334 = ~n8327 & n8333 ;
  assign n8338 = \P3_InstAddrPointer_reg[21]/NET0131  & n2896 ;
  assign n8339 = n4167 & n4230 ;
  assign n8340 = n6042 & n6062 ;
  assign n8341 = ~n4254 & n8340 ;
  assign n8342 = n8339 & n8341 ;
  assign n8343 = n4257 & ~n8342 ;
  assign n8344 = ~n4257 & n8342 ;
  assign n8345 = ~n8343 & ~n8344 ;
  assign n8346 = ~n3753 & ~n8345 ;
  assign n8351 = n4061 & ~n4070 ;
  assign n8352 = ~n4055 & n8351 ;
  assign n8353 = ~\P3_InstAddrPointer_reg[9]/NET0131  & ~n3767 ;
  assign n8354 = ~n3778 & ~n8353 ;
  assign n8355 = \P3_InstAddrPointer_reg[12]/NET0131  & n8354 ;
  assign n8356 = n6072 & n8355 ;
  assign n8357 = n8352 & n8356 ;
  assign n8358 = ~n4095 & ~n4173 ;
  assign n8359 = n4079 & n8358 ;
  assign n8360 = n6089 & n8359 ;
  assign n8361 = n8357 & n8360 ;
  assign n8349 = ~\P3_InstAddrPointer_reg[17]/NET0131  & ~n4076 ;
  assign n8350 = ~n3784 & ~n8349 ;
  assign n8362 = n7381 & n8350 ;
  assign n8363 = n8361 & n8362 ;
  assign n8364 = ~n3789 & ~n8363 ;
  assign n8347 = n3792 & n6093 ;
  assign n8348 = n3789 & n8347 ;
  assign n8365 = n3753 & ~n8348 ;
  assign n8366 = ~n8364 & n8365 ;
  assign n8367 = ~n8346 & ~n8366 ;
  assign n8368 = ~n2896 & ~n8367 ;
  assign n8369 = ~n8338 & ~n8368 ;
  assign n8370 = n2894 & ~n8369 ;
  assign n8378 = n4362 & n4368 ;
  assign n8377 = ~n4362 & ~n4368 ;
  assign n8379 = n2905 & ~n8377 ;
  assign n8380 = ~n8378 & n8379 ;
  assign n8382 = ~\P3_InstAddrPointer_reg[21]/NET0131  & ~n2847 ;
  assign n8383 = ~n2841 & ~n8382 ;
  assign n8384 = n4368 & n8383 ;
  assign n8371 = ~n2823 & n2901 ;
  assign n8372 = ~n2819 & n3789 ;
  assign n8373 = ~n2890 & ~n7401 ;
  assign n8374 = ~n8372 & n8373 ;
  assign n8375 = n8371 & n8374 ;
  assign n8376 = \P3_InstAddrPointer_reg[21]/NET0131  & ~n8375 ;
  assign n8337 = ~n2777 & n4257 ;
  assign n8381 = ~n2923 & n3789 ;
  assign n8385 = ~n8337 & ~n8381 ;
  assign n8386 = ~n8376 & n8385 ;
  assign n8387 = ~n8384 & n8386 ;
  assign n8388 = ~n8380 & n8387 ;
  assign n8389 = ~n8370 & n8388 ;
  assign n8390 = n2453 & ~n8389 ;
  assign n8335 = \P3_InstAddrPointer_reg[21]/NET0131  & ~n4418 ;
  assign n8336 = \P3_rEIP_reg[21]/NET0131  & n4412 ;
  assign n8391 = ~n8335 & ~n8336 ;
  assign n8392 = ~n8390 & n8391 ;
  assign n8393 = n6059 & n8340 ;
  assign n8394 = n4258 & n4270 ;
  assign n8395 = n8393 & n8394 ;
  assign n8396 = ~n4263 & n8395 ;
  assign n8397 = n4274 & ~n8396 ;
  assign n8398 = n4271 & ~n4274 ;
  assign n8399 = n8344 & n8398 ;
  assign n8400 = ~n3753 & ~n8399 ;
  assign n8401 = ~n8397 & n8400 ;
  assign n8402 = n3790 & n4105 ;
  assign n8403 = n8363 & n8402 ;
  assign n8405 = n4100 & n8403 ;
  assign n8404 = ~n4100 & ~n8403 ;
  assign n8406 = n3753 & ~n8404 ;
  assign n8407 = ~n8405 & n8406 ;
  assign n8408 = ~n8401 & ~n8407 ;
  assign n8409 = ~n2896 & ~n8408 ;
  assign n8410 = \P3_InstAddrPointer_reg[25]/NET0131  & n2896 ;
  assign n8411 = ~n8409 & ~n8410 ;
  assign n8412 = n2894 & ~n8411 ;
  assign n8415 = n4374 & n4379 ;
  assign n8414 = ~n4374 & ~n4379 ;
  assign n8416 = n2905 & ~n8414 ;
  assign n8417 = ~n8415 & n8416 ;
  assign n8418 = ~n2835 & ~n4100 ;
  assign n8419 = n2820 & ~n8418 ;
  assign n8420 = n7404 & ~n8419 ;
  assign n8421 = \P3_InstAddrPointer_reg[25]/NET0131  & ~n8420 ;
  assign n8423 = ~n2923 & n4100 ;
  assign n8413 = n2918 & n4379 ;
  assign n8422 = ~n2777 & ~n4274 ;
  assign n8424 = ~n8413 & ~n8422 ;
  assign n8425 = ~n8423 & n8424 ;
  assign n8426 = ~n8421 & n8425 ;
  assign n8427 = ~n8417 & n8426 ;
  assign n8428 = ~n8412 & n8427 ;
  assign n8429 = n2453 & ~n8428 ;
  assign n8430 = \P3_rEIP_reg[25]/NET0131  & n4412 ;
  assign n8431 = \P3_InstAddrPointer_reg[25]/NET0131  & ~n4418 ;
  assign n8432 = ~n8430 & ~n8431 ;
  assign n8433 = ~n8429 & n8432 ;
  assign n8437 = \P2_InstAddrPointer_reg[11]/NET0131  & n1897 ;
  assign n8442 = ~n7439 & ~n7462 ;
  assign n8443 = n6603 & ~n7455 ;
  assign n8444 = n6646 & n8443 ;
  assign n8445 = ~n8442 & ~n8444 ;
  assign n8446 = n6188 & ~n8445 ;
  assign n8438 = ~n6485 & ~n7472 ;
  assign n8439 = n6485 & n7472 ;
  assign n8440 = ~n8438 & ~n8439 ;
  assign n8441 = ~n6188 & ~n8440 ;
  assign n8447 = ~n1897 & ~n8441 ;
  assign n8448 = ~n8446 & n8447 ;
  assign n8449 = ~n8437 & ~n8448 ;
  assign n8450 = n1734 & ~n8449 ;
  assign n8452 = n7485 & n7491 ;
  assign n8451 = ~n7485 & ~n7491 ;
  assign n8453 = n1890 & ~n8451 ;
  assign n8454 = ~n8452 & n8453 ;
  assign n8436 = \P2_InstAddrPointer_reg[11]/NET0131  & ~n7501 ;
  assign n8457 = ~n1798 & n6742 ;
  assign n8458 = n7491 & ~n8457 ;
  assign n8459 = ~n1727 & n8458 ;
  assign n8460 = ~n8436 & ~n8459 ;
  assign n8455 = ~n1771 & n6485 ;
  assign n8456 = ~n1831 & n7439 ;
  assign n8461 = ~n8455 & ~n8456 ;
  assign n8462 = n8460 & n8461 ;
  assign n8463 = ~n8454 & n8462 ;
  assign n8464 = ~n8450 & n8463 ;
  assign n8465 = n1927 & ~n8464 ;
  assign n8434 = \P2_rEIP_reg[11]/NET0131  & n3113 ;
  assign n8435 = \P2_InstAddrPointer_reg[11]/NET0131  & ~n6810 ;
  assign n8466 = ~n8434 & ~n8435 ;
  assign n8467 = ~n8465 & n8466 ;
  assign n8469 = \P2_InstAddrPointer_reg[18]/NET0131  & n1897 ;
  assign n8474 = ~n6524 & n7516 ;
  assign n8476 = ~n6527 & n8474 ;
  assign n8475 = n6527 & ~n8474 ;
  assign n8477 = ~n6188 & ~n8475 ;
  assign n8478 = ~n8476 & n8477 ;
  assign n8470 = n7457 & n7523 ;
  assign n8471 = ~n6663 & ~n8470 ;
  assign n8472 = ~n7592 & ~n8471 ;
  assign n8473 = n6188 & ~n8472 ;
  assign n8479 = ~n1897 & ~n8473 ;
  assign n8480 = ~n8478 & n8479 ;
  assign n8481 = ~n8469 & ~n8480 ;
  assign n8482 = n1734 & ~n8481 ;
  assign n8483 = ~n7538 & ~n7549 ;
  assign n8484 = n1890 & ~n7550 ;
  assign n8485 = ~n8483 & n8484 ;
  assign n8486 = \P2_InstAddrPointer_reg[18]/NET0131  & n1891 ;
  assign n8487 = n1831 & ~n8486 ;
  assign n8488 = n6663 & ~n8487 ;
  assign n8492 = ~n1798 & n6754 ;
  assign n8493 = \P2_InstAddrPointer_reg[17]/NET0131  & n8492 ;
  assign n8494 = ~n1727 & n7538 ;
  assign n8495 = ~n8493 & n8494 ;
  assign n8468 = ~n1771 & n6527 ;
  assign n8489 = ~n1821 & ~n1892 ;
  assign n8490 = n7500 & n8489 ;
  assign n8491 = \P2_InstAddrPointer_reg[18]/NET0131  & ~n8490 ;
  assign n8496 = ~n8468 & ~n8491 ;
  assign n8497 = ~n8495 & n8496 ;
  assign n8498 = ~n8488 & n8497 ;
  assign n8499 = ~n8485 & n8498 ;
  assign n8500 = ~n8482 & n8499 ;
  assign n8501 = n1927 & ~n8500 ;
  assign n8502 = \P2_rEIP_reg[18]/NET0131  & n3113 ;
  assign n8503 = \P2_InstAddrPointer_reg[18]/NET0131  & ~n6810 ;
  assign n8504 = ~n8502 & ~n8503 ;
  assign n8505 = ~n8501 & n8504 ;
  assign n8508 = \P2_InstAddrPointer_reg[25]/NET0131  & n1897 ;
  assign n8513 = ~n6671 & ~n6673 ;
  assign n8514 = ~n7588 & ~n8513 ;
  assign n8515 = n6188 & ~n8514 ;
  assign n8510 = n6563 & ~n6571 ;
  assign n8509 = ~n6563 & n6571 ;
  assign n8511 = ~n6188 & ~n8509 ;
  assign n8512 = ~n8510 & n8511 ;
  assign n8516 = ~n1897 & ~n8512 ;
  assign n8517 = ~n8515 & n8516 ;
  assign n8518 = ~n8508 & ~n8517 ;
  assign n8519 = n1734 & ~n8518 ;
  assign n8522 = n6772 & n6781 ;
  assign n8521 = ~n6772 & ~n6781 ;
  assign n8523 = n1890 & ~n8521 ;
  assign n8524 = ~n8522 & n8523 ;
  assign n8533 = n1870 & n6781 ;
  assign n8525 = ~n1727 & ~n6773 ;
  assign n8526 = ~n1747 & n1805 ;
  assign n8527 = ~n1852 & ~n8526 ;
  assign n8528 = ~n1810 & ~n8527 ;
  assign n8529 = n7500 & ~n8528 ;
  assign n8530 = ~n8525 & n8529 ;
  assign n8531 = \P2_InstAddrPointer_reg[25]/NET0131  & ~n8530 ;
  assign n8520 = ~n1831 & n6673 ;
  assign n8532 = ~n1771 & n6571 ;
  assign n8534 = ~n8520 & ~n8532 ;
  assign n8535 = ~n8531 & n8534 ;
  assign n8536 = ~n8533 & n8535 ;
  assign n8537 = ~n8524 & n8536 ;
  assign n8538 = ~n8519 & n8537 ;
  assign n8539 = n1927 & ~n8538 ;
  assign n8506 = \P2_rEIP_reg[25]/NET0131  & n3113 ;
  assign n8507 = \P2_InstAddrPointer_reg[25]/NET0131  & ~n6810 ;
  assign n8540 = ~n8506 & ~n8507 ;
  assign n8541 = ~n8539 & n8540 ;
  assign n8543 = \P1_InstAddrPointer_reg[18]/NET0131  & n2375 ;
  assign n8550 = ~n4918 & n7274 ;
  assign n8551 = ~n4916 & n8550 ;
  assign n8552 = n4887 & n8551 ;
  assign n8553 = n4921 & ~n8552 ;
  assign n8548 = n4887 & n7274 ;
  assign n8549 = n4923 & n8548 ;
  assign n8554 = ~n4453 & ~n8549 ;
  assign n8555 = ~n8553 & n8554 ;
  assign n8544 = ~n4776 & ~n5974 ;
  assign n8545 = \P1_InstAddrPointer_reg[18]/NET0131  & n5974 ;
  assign n8546 = ~n8544 & ~n8545 ;
  assign n8547 = n4453 & ~n8546 ;
  assign n8556 = ~n2375 & ~n8547 ;
  assign n8557 = ~n8555 & n8556 ;
  assign n8558 = ~n8543 & ~n8557 ;
  assign n8559 = n2244 & ~n8558 ;
  assign n8561 = n4970 & n5038 ;
  assign n8560 = ~n4970 & ~n5038 ;
  assign n8562 = n2385 & ~n8560 ;
  assign n8563 = ~n8561 & n8562 ;
  assign n8564 = n2387 & ~n4776 ;
  assign n8565 = n7308 & ~n8564 ;
  assign n8566 = n6026 & ~n8565 ;
  assign n8567 = \P1_InstAddrPointer_reg[18]/NET0131  & ~n8566 ;
  assign n8573 = ~\P1_InstAddrPointer_reg[18]/NET0131  & ~n2337 ;
  assign n8574 = ~n2332 & ~n8573 ;
  assign n8575 = n4970 & n8574 ;
  assign n8542 = ~n2271 & n4921 ;
  assign n8568 = n2237 & n4776 ;
  assign n8569 = ~\P1_InstAddrPointer_reg[18]/NET0131  & n2317 ;
  assign n8570 = ~n2317 & ~n4776 ;
  assign n8571 = ~n8569 & ~n8570 ;
  assign n8572 = ~n2314 & n8571 ;
  assign n8576 = ~n8568 & ~n8572 ;
  assign n8577 = ~n8542 & n8576 ;
  assign n8578 = ~n8575 & n8577 ;
  assign n8579 = ~n8567 & n8578 ;
  assign n8580 = ~n8563 & n8579 ;
  assign n8581 = ~n8559 & n8580 ;
  assign n8582 = n2432 & ~n8581 ;
  assign n8583 = \P1_InstAddrPointer_reg[18]/NET0131  & ~n5098 ;
  assign n8584 = \P1_rEIP_reg[18]/NET0131  & n5092 ;
  assign n8585 = ~n8583 & ~n8584 ;
  assign n8586 = ~n8582 & n8585 ;
  assign n8595 = \buf2_reg[26]/NET0131  & ~n3079 ;
  assign n8596 = \buf1_reg[26]/NET0131  & n3079 ;
  assign n8597 = ~n8595 & ~n8596 ;
  assign n8598 = n3091 & ~n8597 ;
  assign n8599 = \buf2_reg[18]/NET0131  & ~n3079 ;
  assign n8600 = \buf1_reg[18]/NET0131  & n3079 ;
  assign n8601 = ~n8599 & ~n8600 ;
  assign n8602 = n3098 & ~n8601 ;
  assign n8603 = ~n8598 & ~n8602 ;
  assign n8604 = \P2_DataWidth_reg[1]/NET0131  & ~n8603 ;
  assign n8587 = \buf2_reg[2]/NET0131  & ~n3079 ;
  assign n8588 = \buf1_reg[2]/NET0131  & n3079 ;
  assign n8589 = ~n8587 & ~n8588 ;
  assign n8590 = ~n3050 & ~n8589 ;
  assign n8591 = \P2_InstQueue_reg[11][2]/NET0131  & ~n3049 ;
  assign n8592 = ~n3046 & n8591 ;
  assign n8593 = ~n8590 & ~n8592 ;
  assign n8605 = ~n3106 & ~n8593 ;
  assign n8606 = ~n8604 & ~n8605 ;
  assign n8607 = n1931 & ~n8606 ;
  assign n8594 = n3087 & ~n8593 ;
  assign n8608 = ~n1561 & n3049 ;
  assign n8609 = ~n8591 & ~n8608 ;
  assign n8610 = n3040 & ~n8609 ;
  assign n8611 = \P2_InstQueue_reg[11][2]/NET0131  & ~n3118 ;
  assign n8612 = ~n8610 & ~n8611 ;
  assign n8613 = ~n8594 & n8612 ;
  assign n8614 = ~n8607 & n8613 ;
  assign n8620 = n3162 & ~n8597 ;
  assign n8621 = n3165 & ~n8601 ;
  assign n8622 = ~n8620 & ~n8621 ;
  assign n8623 = \P2_DataWidth_reg[1]/NET0131  & ~n8622 ;
  assign n8615 = ~n3155 & ~n8589 ;
  assign n8616 = \P2_InstQueue_reg[0][2]/NET0131  & ~n3152 ;
  assign n8617 = ~n3154 & n8616 ;
  assign n8618 = ~n8615 & ~n8617 ;
  assign n8624 = ~n3170 & ~n8618 ;
  assign n8625 = ~n8623 & ~n8624 ;
  assign n8626 = n1931 & ~n8625 ;
  assign n8619 = n3087 & ~n8618 ;
  assign n8627 = ~n1561 & n3152 ;
  assign n8628 = ~n8616 & ~n8627 ;
  assign n8629 = n3040 & ~n8628 ;
  assign n8630 = \P2_InstQueue_reg[0][2]/NET0131  & ~n3118 ;
  assign n8631 = ~n8629 & ~n8630 ;
  assign n8632 = ~n8619 & n8631 ;
  assign n8633 = ~n8626 & n8632 ;
  assign n8639 = n3091 & ~n8601 ;
  assign n8640 = n3198 & ~n8597 ;
  assign n8641 = ~n8639 & ~n8640 ;
  assign n8642 = \P2_DataWidth_reg[1]/NET0131  & ~n8641 ;
  assign n8634 = ~n3202 & ~n8589 ;
  assign n8635 = \P2_InstQueue_reg[10][2]/NET0131  & ~n3046 ;
  assign n8636 = ~n3098 & n8635 ;
  assign n8637 = ~n8634 & ~n8636 ;
  assign n8643 = ~n3200 & ~n8637 ;
  assign n8644 = ~n8642 & ~n8643 ;
  assign n8645 = n1931 & ~n8644 ;
  assign n8638 = n3087 & ~n8637 ;
  assign n8646 = ~n1561 & n3046 ;
  assign n8647 = ~n8635 & ~n8646 ;
  assign n8648 = n3040 & ~n8647 ;
  assign n8649 = \P2_InstQueue_reg[10][2]/NET0131  & ~n3118 ;
  assign n8650 = ~n8648 & ~n8649 ;
  assign n8651 = ~n8638 & n8650 ;
  assign n8652 = ~n8645 & n8651 ;
  assign n8658 = n3098 & ~n8597 ;
  assign n8659 = n3046 & ~n8601 ;
  assign n8660 = ~n8658 & ~n8659 ;
  assign n8661 = \P2_DataWidth_reg[1]/NET0131  & ~n8660 ;
  assign n8653 = ~n3238 & ~n8589 ;
  assign n8654 = \P2_InstQueue_reg[12][2]/NET0131  & ~n3237 ;
  assign n8655 = ~n3049 & n8654 ;
  assign n8656 = ~n8653 & ~n8655 ;
  assign n8662 = ~n3248 & ~n8656 ;
  assign n8663 = ~n8661 & ~n8662 ;
  assign n8664 = n1931 & ~n8663 ;
  assign n8657 = n3087 & ~n8656 ;
  assign n8665 = ~n1561 & n3237 ;
  assign n8666 = ~n8654 & ~n8665 ;
  assign n8667 = n3040 & ~n8666 ;
  assign n8668 = \P2_InstQueue_reg[12][2]/NET0131  & ~n3118 ;
  assign n8669 = ~n8667 & ~n8668 ;
  assign n8670 = ~n8657 & n8669 ;
  assign n8671 = ~n8664 & n8670 ;
  assign n8677 = n3046 & ~n8597 ;
  assign n8678 = n3049 & ~n8601 ;
  assign n8679 = ~n8677 & ~n8678 ;
  assign n8680 = \P2_DataWidth_reg[1]/NET0131  & ~n8679 ;
  assign n8672 = ~n3275 & ~n8589 ;
  assign n8673 = \P2_InstQueue_reg[13][2]/NET0131  & ~n3162 ;
  assign n8674 = ~n3237 & n8673 ;
  assign n8675 = ~n8672 & ~n8674 ;
  assign n8681 = ~n3285 & ~n8675 ;
  assign n8682 = ~n8680 & ~n8681 ;
  assign n8683 = n1931 & ~n8682 ;
  assign n8676 = n3087 & ~n8675 ;
  assign n8684 = ~n1561 & n3162 ;
  assign n8685 = ~n8673 & ~n8684 ;
  assign n8686 = n3040 & ~n8685 ;
  assign n8687 = \P2_InstQueue_reg[13][2]/NET0131  & ~n3118 ;
  assign n8688 = ~n8686 & ~n8687 ;
  assign n8689 = ~n8676 & n8688 ;
  assign n8690 = ~n8683 & n8689 ;
  assign n8696 = n3049 & ~n8597 ;
  assign n8697 = n3237 & ~n8601 ;
  assign n8698 = ~n8696 & ~n8697 ;
  assign n8699 = \P2_DataWidth_reg[1]/NET0131  & ~n8698 ;
  assign n8691 = ~n3169 & ~n8589 ;
  assign n8692 = \P2_InstQueue_reg[14][2]/NET0131  & ~n3165 ;
  assign n8693 = ~n3162 & n8692 ;
  assign n8694 = ~n8691 & ~n8693 ;
  assign n8700 = ~n3321 & ~n8694 ;
  assign n8701 = ~n8699 & ~n8700 ;
  assign n8702 = n1931 & ~n8701 ;
  assign n8695 = n3087 & ~n8694 ;
  assign n8703 = ~n1561 & n3165 ;
  assign n8704 = ~n8692 & ~n8703 ;
  assign n8705 = n3040 & ~n8704 ;
  assign n8706 = \P2_InstQueue_reg[14][2]/NET0131  & ~n3118 ;
  assign n8707 = ~n8705 & ~n8706 ;
  assign n8708 = ~n8695 & n8707 ;
  assign n8709 = ~n8702 & n8708 ;
  assign n8715 = n3237 & ~n8597 ;
  assign n8716 = n3162 & ~n8601 ;
  assign n8717 = ~n8715 & ~n8716 ;
  assign n8718 = \P2_DataWidth_reg[1]/NET0131  & ~n8717 ;
  assign n8710 = ~n3348 & ~n8589 ;
  assign n8711 = \P2_InstQueue_reg[15][2]/NET0131  & ~n3154 ;
  assign n8712 = ~n3165 & n8711 ;
  assign n8713 = ~n8710 & ~n8712 ;
  assign n8719 = ~n3358 & ~n8713 ;
  assign n8720 = ~n8718 & ~n8719 ;
  assign n8721 = n1931 & ~n8720 ;
  assign n8714 = n3087 & ~n8713 ;
  assign n8722 = ~n1561 & n3154 ;
  assign n8723 = ~n8711 & ~n8722 ;
  assign n8724 = n3040 & ~n8723 ;
  assign n8725 = \P2_InstQueue_reg[15][2]/NET0131  & ~n3118 ;
  assign n8726 = ~n8724 & ~n8725 ;
  assign n8727 = ~n8714 & n8726 ;
  assign n8728 = ~n8721 & n8727 ;
  assign n8734 = n3165 & ~n8597 ;
  assign n8735 = n3154 & ~n8601 ;
  assign n8736 = ~n8734 & ~n8735 ;
  assign n8737 = \P2_DataWidth_reg[1]/NET0131  & ~n8736 ;
  assign n8729 = ~n3389 & ~n8589 ;
  assign n8730 = \P2_InstQueue_reg[1][2]/NET0131  & ~n3388 ;
  assign n8731 = ~n3152 & n8730 ;
  assign n8732 = ~n8729 & ~n8731 ;
  assign n8738 = ~n3386 & ~n8732 ;
  assign n8739 = ~n8737 & ~n8738 ;
  assign n8740 = n1931 & ~n8739 ;
  assign n8733 = n3087 & ~n8732 ;
  assign n8741 = ~n1561 & n3388 ;
  assign n8742 = ~n8730 & ~n8741 ;
  assign n8743 = n3040 & ~n8742 ;
  assign n8744 = \P2_InstQueue_reg[1][2]/NET0131  & ~n3118 ;
  assign n8745 = ~n8743 & ~n8744 ;
  assign n8746 = ~n8733 & n8745 ;
  assign n8747 = ~n8740 & n8746 ;
  assign n8753 = n3152 & ~n8601 ;
  assign n8754 = n3154 & ~n8597 ;
  assign n8755 = ~n8753 & ~n8754 ;
  assign n8756 = \P2_DataWidth_reg[1]/NET0131  & ~n8755 ;
  assign n8748 = ~n3424 & ~n8589 ;
  assign n8749 = \P2_InstQueue_reg[2][2]/NET0131  & ~n3423 ;
  assign n8750 = ~n3388 & n8749 ;
  assign n8751 = ~n8748 & ~n8750 ;
  assign n8757 = ~n3434 & ~n8751 ;
  assign n8758 = ~n8756 & ~n8757 ;
  assign n8759 = n1931 & ~n8758 ;
  assign n8752 = n3087 & ~n8751 ;
  assign n8760 = ~n1561 & n3423 ;
  assign n8761 = ~n8749 & ~n8760 ;
  assign n8762 = n3040 & ~n8761 ;
  assign n8763 = \P2_InstQueue_reg[2][2]/NET0131  & ~n3118 ;
  assign n8764 = ~n8762 & ~n8763 ;
  assign n8765 = ~n8752 & n8764 ;
  assign n8766 = ~n8759 & n8765 ;
  assign n8772 = n3152 & ~n8597 ;
  assign n8773 = n3388 & ~n8601 ;
  assign n8774 = ~n8772 & ~n8773 ;
  assign n8775 = \P2_DataWidth_reg[1]/NET0131  & ~n8774 ;
  assign n8767 = ~n3462 & ~n8589 ;
  assign n8768 = \P2_InstQueue_reg[3][2]/NET0131  & ~n3461 ;
  assign n8769 = ~n3423 & n8768 ;
  assign n8770 = ~n8767 & ~n8769 ;
  assign n8776 = ~n3472 & ~n8770 ;
  assign n8777 = ~n8775 & ~n8776 ;
  assign n8778 = n1931 & ~n8777 ;
  assign n8771 = n3087 & ~n8770 ;
  assign n8779 = ~n1561 & n3461 ;
  assign n8780 = ~n8768 & ~n8779 ;
  assign n8781 = n3040 & ~n8780 ;
  assign n8782 = \P2_InstQueue_reg[3][2]/NET0131  & ~n3118 ;
  assign n8783 = ~n8781 & ~n8782 ;
  assign n8784 = ~n8771 & n8783 ;
  assign n8785 = ~n8778 & n8784 ;
  assign n8791 = n3388 & ~n8597 ;
  assign n8792 = n3423 & ~n8601 ;
  assign n8793 = ~n8791 & ~n8792 ;
  assign n8794 = \P2_DataWidth_reg[1]/NET0131  & ~n8793 ;
  assign n8786 = ~n3500 & ~n8589 ;
  assign n8787 = \P2_InstQueue_reg[4][2]/NET0131  & ~n3499 ;
  assign n8788 = ~n3461 & n8787 ;
  assign n8789 = ~n8786 & ~n8788 ;
  assign n8795 = ~n3510 & ~n8789 ;
  assign n8796 = ~n8794 & ~n8795 ;
  assign n8797 = n1931 & ~n8796 ;
  assign n8790 = n3087 & ~n8789 ;
  assign n8798 = ~n1561 & n3499 ;
  assign n8799 = ~n8787 & ~n8798 ;
  assign n8800 = n3040 & ~n8799 ;
  assign n8801 = \P2_InstQueue_reg[4][2]/NET0131  & ~n3118 ;
  assign n8802 = ~n8800 & ~n8801 ;
  assign n8803 = ~n8790 & n8802 ;
  assign n8804 = ~n8797 & n8803 ;
  assign n8810 = n3423 & ~n8597 ;
  assign n8811 = n3461 & ~n8601 ;
  assign n8812 = ~n8810 & ~n8811 ;
  assign n8813 = \P2_DataWidth_reg[1]/NET0131  & ~n8812 ;
  assign n8805 = ~n3538 & ~n8589 ;
  assign n8806 = \P2_InstQueue_reg[5][2]/NET0131  & ~n3537 ;
  assign n8807 = ~n3499 & n8806 ;
  assign n8808 = ~n8805 & ~n8807 ;
  assign n8814 = ~n3548 & ~n8808 ;
  assign n8815 = ~n8813 & ~n8814 ;
  assign n8816 = n1931 & ~n8815 ;
  assign n8809 = n3087 & ~n8808 ;
  assign n8817 = ~n1561 & n3537 ;
  assign n8818 = ~n8806 & ~n8817 ;
  assign n8819 = n3040 & ~n8818 ;
  assign n8820 = \P2_InstQueue_reg[5][2]/NET0131  & ~n3118 ;
  assign n8821 = ~n8819 & ~n8820 ;
  assign n8822 = ~n8809 & n8821 ;
  assign n8823 = ~n8816 & n8822 ;
  assign n8829 = n3461 & ~n8597 ;
  assign n8830 = n3499 & ~n8601 ;
  assign n8831 = ~n8829 & ~n8830 ;
  assign n8832 = \P2_DataWidth_reg[1]/NET0131  & ~n8831 ;
  assign n8824 = ~n3576 & ~n8589 ;
  assign n8825 = \P2_InstQueue_reg[6][2]/NET0131  & ~n3575 ;
  assign n8826 = ~n3537 & n8825 ;
  assign n8827 = ~n8824 & ~n8826 ;
  assign n8833 = ~n3586 & ~n8827 ;
  assign n8834 = ~n8832 & ~n8833 ;
  assign n8835 = n1931 & ~n8834 ;
  assign n8828 = n3087 & ~n8827 ;
  assign n8836 = ~n1561 & n3575 ;
  assign n8837 = ~n8825 & ~n8836 ;
  assign n8838 = n3040 & ~n8837 ;
  assign n8839 = \P2_InstQueue_reg[6][2]/NET0131  & ~n3118 ;
  assign n8840 = ~n8838 & ~n8839 ;
  assign n8841 = ~n8828 & n8840 ;
  assign n8842 = ~n8835 & n8841 ;
  assign n8848 = n3499 & ~n8597 ;
  assign n8849 = n3537 & ~n8601 ;
  assign n8850 = ~n8848 & ~n8849 ;
  assign n8851 = \P2_DataWidth_reg[1]/NET0131  & ~n8850 ;
  assign n8843 = ~n3613 & ~n8589 ;
  assign n8844 = \P2_InstQueue_reg[7][2]/NET0131  & ~n3198 ;
  assign n8845 = ~n3575 & n8844 ;
  assign n8846 = ~n8843 & ~n8845 ;
  assign n8852 = ~n3623 & ~n8846 ;
  assign n8853 = ~n8851 & ~n8852 ;
  assign n8854 = n1931 & ~n8853 ;
  assign n8847 = n3087 & ~n8846 ;
  assign n8855 = ~n1561 & n3198 ;
  assign n8856 = ~n8844 & ~n8855 ;
  assign n8857 = n3040 & ~n8856 ;
  assign n8858 = \P2_InstQueue_reg[7][2]/NET0131  & ~n3118 ;
  assign n8859 = ~n8857 & ~n8858 ;
  assign n8860 = ~n8847 & n8859 ;
  assign n8861 = ~n8854 & n8860 ;
  assign n8867 = n3537 & ~n8597 ;
  assign n8868 = n3575 & ~n8601 ;
  assign n8869 = ~n8867 & ~n8868 ;
  assign n8870 = \P2_DataWidth_reg[1]/NET0131  & ~n8869 ;
  assign n8862 = ~n3199 & ~n8589 ;
  assign n8863 = \P2_InstQueue_reg[8][2]/NET0131  & ~n3091 ;
  assign n8864 = ~n3198 & n8863 ;
  assign n8865 = ~n8862 & ~n8864 ;
  assign n8871 = ~n3659 & ~n8865 ;
  assign n8872 = ~n8870 & ~n8871 ;
  assign n8873 = n1931 & ~n8872 ;
  assign n8866 = n3087 & ~n8865 ;
  assign n8874 = ~n1561 & n3091 ;
  assign n8875 = ~n8863 & ~n8874 ;
  assign n8876 = n3040 & ~n8875 ;
  assign n8877 = \P2_InstQueue_reg[8][2]/NET0131  & ~n3118 ;
  assign n8878 = ~n8876 & ~n8877 ;
  assign n8879 = ~n8866 & n8878 ;
  assign n8880 = ~n8873 & n8879 ;
  assign n8886 = n3575 & ~n8597 ;
  assign n8887 = n3198 & ~n8601 ;
  assign n8888 = ~n8886 & ~n8887 ;
  assign n8889 = \P2_DataWidth_reg[1]/NET0131  & ~n8888 ;
  assign n8881 = ~n3105 & ~n8589 ;
  assign n8882 = \P2_InstQueue_reg[9][2]/NET0131  & ~n3098 ;
  assign n8883 = ~n3091 & n8882 ;
  assign n8884 = ~n8881 & ~n8883 ;
  assign n8890 = ~n3695 & ~n8884 ;
  assign n8891 = ~n8889 & ~n8890 ;
  assign n8892 = n1931 & ~n8891 ;
  assign n8885 = n3087 & ~n8884 ;
  assign n8893 = ~n1561 & n3098 ;
  assign n8894 = ~n8882 & ~n8893 ;
  assign n8895 = n3040 & ~n8894 ;
  assign n8896 = \P2_InstQueue_reg[9][2]/NET0131  & ~n3118 ;
  assign n8897 = ~n8895 & ~n8896 ;
  assign n8898 = ~n8885 & n8897 ;
  assign n8899 = ~n8892 & n8898 ;
  assign n8900 = \P2_PhyAddrPointer_reg[31]/NET0131  & n1897 ;
  assign n8912 = ~n6515 & n6528 ;
  assign n8913 = ~n6506 & n8912 ;
  assign n8914 = n7473 & n8913 ;
  assign n8915 = n6540 & n6551 ;
  assign n8916 = n8914 & n8915 ;
  assign n8920 = n6580 & ~n6588 ;
  assign n8917 = ~\P2_InstAddrPointer_reg[30]/NET0131  & ~n6587 ;
  assign n8918 = \P2_InstAddrPointer_reg[30]/NET0131  & n6587 ;
  assign n8919 = ~n8917 & ~n8918 ;
  assign n8921 = n6561 & n6572 ;
  assign n8922 = ~n8919 & n8921 ;
  assign n8923 = n8920 & n8922 ;
  assign n8924 = n8916 & n8923 ;
  assign n8925 = \P2_InstAddrPointer_reg[31]/NET0131  & ~n8918 ;
  assign n8926 = ~\P2_InstAddrPointer_reg[31]/NET0131  & n8918 ;
  assign n8927 = ~n8925 & ~n8926 ;
  assign n8929 = n8924 & n8927 ;
  assign n8928 = ~n8924 & ~n8927 ;
  assign n8930 = ~n6188 & ~n8928 ;
  assign n8931 = ~n8929 & n8930 ;
  assign n8901 = \P2_InstAddrPointer_reg[29]/NET0131  & \P2_InstAddrPointer_reg[30]/NET0131  ;
  assign n8902 = n6677 & n8901 ;
  assign n8903 = n7598 & n8902 ;
  assign n8904 = n6585 & n8901 ;
  assign n8905 = ~\P2_InstAddrPointer_reg[31]/NET0131  & ~n8904 ;
  assign n8906 = \P2_InstAddrPointer_reg[31]/NET0131  & n8904 ;
  assign n8907 = ~n8905 & ~n8906 ;
  assign n8909 = n8903 & ~n8907 ;
  assign n8908 = ~n8903 & n8907 ;
  assign n8910 = n6188 & ~n8908 ;
  assign n8911 = ~n8909 & n8910 ;
  assign n8932 = ~n1897 & ~n8911 ;
  assign n8933 = ~n8931 & n8932 ;
  assign n8934 = ~n8900 & ~n8933 ;
  assign n8935 = n1734 & ~n8934 ;
  assign n8936 = ~n1735 & ~n1902 ;
  assign n8937 = \P2_PhyAddrPointer_reg[31]/NET0131  & ~n8936 ;
  assign n8938 = \P2_InstAddrPointer_reg[16]/NET0131  & \P2_InstAddrPointer_reg[18]/NET0131  ;
  assign n8939 = n7483 & n8938 ;
  assign n8940 = n6757 & n8939 ;
  assign n8941 = n7494 & n8940 ;
  assign n8942 = n7553 & n8941 ;
  assign n8943 = n7627 & n8942 ;
  assign n8944 = n6779 & n8901 ;
  assign n8945 = n8943 & n8944 ;
  assign n8946 = n6785 & n8901 ;
  assign n8947 = \P2_InstAddrPointer_reg[31]/NET0131  & ~n8946 ;
  assign n8948 = ~\P2_InstAddrPointer_reg[31]/NET0131  & n8946 ;
  assign n8949 = ~n8947 & ~n8948 ;
  assign n8951 = n8945 & ~n8949 ;
  assign n8950 = ~n8945 & n8949 ;
  assign n8952 = n1890 & ~n8950 ;
  assign n8953 = ~n8951 & n8952 ;
  assign n8954 = ~n8937 & ~n8953 ;
  assign n8955 = ~n8935 & n8954 ;
  assign n8956 = n1927 & ~n8955 ;
  assign n8960 = \P2_PhyAddrPointer_reg[2]/NET0131  & \P2_PhyAddrPointer_reg[3]/NET0131  ;
  assign n8961 = \P2_PhyAddrPointer_reg[4]/NET0131  & n8960 ;
  assign n8962 = \P2_PhyAddrPointer_reg[5]/NET0131  & n8961 ;
  assign n8963 = \P2_PhyAddrPointer_reg[6]/NET0131  & n8962 ;
  assign n8964 = \P2_PhyAddrPointer_reg[7]/NET0131  & n8963 ;
  assign n8965 = \P2_PhyAddrPointer_reg[8]/NET0131  & n8964 ;
  assign n8966 = \P2_PhyAddrPointer_reg[9]/NET0131  & n8965 ;
  assign n8967 = \P2_PhyAddrPointer_reg[10]/NET0131  & \P2_PhyAddrPointer_reg[11]/NET0131  ;
  assign n8968 = n8966 & n8967 ;
  assign n8969 = \P2_PhyAddrPointer_reg[12]/NET0131  & \P2_PhyAddrPointer_reg[13]/NET0131  ;
  assign n8970 = \P2_PhyAddrPointer_reg[14]/NET0131  & n8969 ;
  assign n8971 = n8968 & n8970 ;
  assign n8972 = \P2_PhyAddrPointer_reg[15]/NET0131  & n8971 ;
  assign n8973 = \P2_PhyAddrPointer_reg[16]/NET0131  & \P2_PhyAddrPointer_reg[17]/NET0131  ;
  assign n8974 = \P2_PhyAddrPointer_reg[18]/NET0131  & n8973 ;
  assign n8975 = n8972 & n8974 ;
  assign n8976 = \P2_PhyAddrPointer_reg[19]/NET0131  & n8975 ;
  assign n8977 = \P2_PhyAddrPointer_reg[20]/NET0131  & n8976 ;
  assign n8978 = \P2_PhyAddrPointer_reg[21]/NET0131  & \P2_PhyAddrPointer_reg[22]/NET0131  ;
  assign n8979 = n8977 & n8978 ;
  assign n8980 = \P2_PhyAddrPointer_reg[23]/NET0131  & n8979 ;
  assign n8981 = \P2_PhyAddrPointer_reg[24]/NET0131  & n8980 ;
  assign n8982 = \P2_PhyAddrPointer_reg[25]/NET0131  & n8981 ;
  assign n8983 = \P2_PhyAddrPointer_reg[26]/NET0131  & n8982 ;
  assign n8984 = \P2_PhyAddrPointer_reg[27]/NET0131  & n8983 ;
  assign n8985 = \P2_PhyAddrPointer_reg[28]/NET0131  & n8984 ;
  assign n8986 = \P2_PhyAddrPointer_reg[29]/NET0131  & n8985 ;
  assign n8987 = \P2_PhyAddrPointer_reg[30]/NET0131  & n8986 ;
  assign n8989 = \P2_PhyAddrPointer_reg[31]/NET0131  & n8987 ;
  assign n8988 = ~\P2_PhyAddrPointer_reg[31]/NET0131  & ~n8987 ;
  assign n8990 = n3034 & ~n8988 ;
  assign n8991 = ~n8989 & n8990 ;
  assign n8993 = \P2_PhyAddrPointer_reg[26]/NET0131  & \P2_PhyAddrPointer_reg[27]/NET0131  ;
  assign n8994 = \P2_PhyAddrPointer_reg[1]/NET0131  & \P2_PhyAddrPointer_reg[24]/NET0131  ;
  assign n8995 = n8980 & n8994 ;
  assign n8996 = \P2_PhyAddrPointer_reg[25]/NET0131  & n8995 ;
  assign n8997 = n8993 & n8996 ;
  assign n8998 = \P2_PhyAddrPointer_reg[28]/NET0131  & n8997 ;
  assign n8999 = \P2_PhyAddrPointer_reg[29]/NET0131  & n8998 ;
  assign n9000 = \P2_PhyAddrPointer_reg[30]/NET0131  & n8999 ;
  assign n9001 = \P2_PhyAddrPointer_reg[31]/NET0131  & ~n9000 ;
  assign n9002 = ~\P2_PhyAddrPointer_reg[31]/NET0131  & n9000 ;
  assign n9003 = ~n9001 & ~n9002 ;
  assign n9004 = \P2_DataWidth_reg[1]/NET0131  & ~n3087 ;
  assign n9005 = ~n3125 & ~n9004 ;
  assign n9006 = ~n9003 & n9005 ;
  assign n8957 = ~n1933 & ~n2979 ;
  assign n8958 = ~n2986 & n8957 ;
  assign n8959 = \P2_PhyAddrPointer_reg[31]/NET0131  & ~n8958 ;
  assign n8992 = \P2_rEIP_reg[31]/NET0131  & n3113 ;
  assign n9007 = ~n8959 & ~n8992 ;
  assign n9008 = ~n9006 & n9007 ;
  assign n9009 = ~n8991 & n9008 ;
  assign n9010 = ~n8956 & n9009 ;
  assign n9011 = \P3_PhyAddrPointer_reg[31]/NET0131  & n2896 ;
  assign n9012 = ~n4290 & ~n9011 ;
  assign n9013 = n2894 & ~n9012 ;
  assign n9014 = n2762 & ~n2900 ;
  assign n9015 = \P3_PhyAddrPointer_reg[31]/NET0131  & ~n9014 ;
  assign n9016 = ~n4400 & ~n9015 ;
  assign n9017 = ~n9013 & n9016 ;
  assign n9018 = n2453 & ~n9017 ;
  assign n9019 = \P3_PhyAddrPointer_reg[28]/NET0131  & \P3_PhyAddrPointer_reg[29]/NET0131  ;
  assign n9020 = \P3_PhyAddrPointer_reg[2]/NET0131  & \P3_PhyAddrPointer_reg[3]/NET0131  ;
  assign n9021 = \P3_PhyAddrPointer_reg[4]/NET0131  & n9020 ;
  assign n9022 = \P3_PhyAddrPointer_reg[5]/NET0131  & n9021 ;
  assign n9023 = \P3_PhyAddrPointer_reg[6]/NET0131  & n9022 ;
  assign n9024 = \P3_PhyAddrPointer_reg[7]/NET0131  & n9023 ;
  assign n9025 = \P3_PhyAddrPointer_reg[8]/NET0131  & n9024 ;
  assign n9026 = \P3_PhyAddrPointer_reg[9]/NET0131  & n9025 ;
  assign n9027 = \P3_PhyAddrPointer_reg[10]/NET0131  & n9026 ;
  assign n9028 = \P3_PhyAddrPointer_reg[11]/NET0131  & n9027 ;
  assign n9029 = \P3_PhyAddrPointer_reg[12]/NET0131  & n9028 ;
  assign n9030 = \P3_PhyAddrPointer_reg[13]/NET0131  & n9029 ;
  assign n9031 = \P3_PhyAddrPointer_reg[14]/NET0131  & \P3_PhyAddrPointer_reg[15]/NET0131  ;
  assign n9032 = \P3_PhyAddrPointer_reg[16]/NET0131  & n9031 ;
  assign n9033 = n9030 & n9032 ;
  assign n9034 = \P3_PhyAddrPointer_reg[17]/NET0131  & n9033 ;
  assign n9035 = \P3_PhyAddrPointer_reg[18]/NET0131  & \P3_PhyAddrPointer_reg[19]/NET0131  ;
  assign n9036 = \P3_PhyAddrPointer_reg[20]/NET0131  & n9035 ;
  assign n9037 = n9034 & n9036 ;
  assign n9038 = \P3_PhyAddrPointer_reg[21]/NET0131  & n9037 ;
  assign n9039 = \P3_PhyAddrPointer_reg[22]/NET0131  & n9038 ;
  assign n9040 = \P3_PhyAddrPointer_reg[23]/NET0131  & \P3_PhyAddrPointer_reg[24]/NET0131  ;
  assign n9041 = \P3_PhyAddrPointer_reg[25]/NET0131  & n9040 ;
  assign n9042 = \P3_PhyAddrPointer_reg[26]/NET0131  & n9041 ;
  assign n9043 = n9039 & n9042 ;
  assign n9044 = \P3_PhyAddrPointer_reg[1]/NET0131  & n9043 ;
  assign n9045 = \P3_PhyAddrPointer_reg[27]/NET0131  & n9044 ;
  assign n9046 = n9019 & n9045 ;
  assign n9047 = \P3_PhyAddrPointer_reg[30]/NET0131  & n9046 ;
  assign n9048 = \P3_PhyAddrPointer_reg[31]/NET0131  & ~n9047 ;
  assign n9049 = \P3_PhyAddrPointer_reg[27]/NET0131  & n9043 ;
  assign n9050 = n9019 & n9049 ;
  assign n9051 = \P3_PhyAddrPointer_reg[30]/NET0131  & n9050 ;
  assign n9052 = ~\P3_PhyAddrPointer_reg[31]/NET0131  & n9051 ;
  assign n9053 = \P3_PhyAddrPointer_reg[1]/NET0131  & n9052 ;
  assign n9054 = ~n9048 & ~n9053 ;
  assign n9056 = ~\P3_DataWidth_reg[1]/NET0131  & ~n9054 ;
  assign n9057 = \P3_PhyAddrPointer_reg[31]/NET0131  & ~n9051 ;
  assign n9058 = ~n9052 & ~n9057 ;
  assign n9059 = \P3_DataWidth_reg[1]/NET0131  & ~n9058 ;
  assign n9060 = ~n9056 & ~n9059 ;
  assign n9061 = n2959 & ~n9060 ;
  assign n9055 = n4415 & ~n9054 ;
  assign n9062 = ~n2953 & ~n2996 ;
  assign n9063 = ~n2993 & n9062 ;
  assign n9064 = \P3_PhyAddrPointer_reg[31]/NET0131  & ~n9063 ;
  assign n9065 = ~n4413 & ~n9064 ;
  assign n9066 = ~n9055 & n9065 ;
  assign n9067 = ~n9061 & n9066 ;
  assign n9068 = ~n9018 & n9067 ;
  assign n9104 = n4304 & ~n6124 ;
  assign n9105 = \P3_InstAddrPointer_reg[9]/NET0131  & n9104 ;
  assign n9106 = n4301 & n9105 ;
  assign n9107 = \P3_InstAddrPointer_reg[11]/NET0131  & n9106 ;
  assign n9109 = \P3_InstAddrPointer_reg[12]/NET0131  & n9107 ;
  assign n9097 = \P3_InstAddrPointer_reg[11]/NET0131  & n4299 ;
  assign n9098 = ~\P3_InstAddrPointer_reg[12]/NET0131  & ~n9097 ;
  assign n9099 = ~n4350 & ~n9098 ;
  assign n9108 = ~n9099 & ~n9107 ;
  assign n9110 = n2905 & ~n9108 ;
  assign n9111 = ~n9109 & n9110 ;
  assign n9071 = \P3_InstAddrPointer_reg[12]/NET0131  & n2896 ;
  assign n9077 = ~n4058 & ~n6088 ;
  assign n9078 = n4058 & n6088 ;
  assign n9079 = ~n9077 & ~n9078 ;
  assign n9080 = n3753 & ~n9079 ;
  assign n9072 = ~n4158 & n6044 ;
  assign n9073 = n6058 & n9072 ;
  assign n9074 = n4166 & ~n9073 ;
  assign n9075 = ~n3753 & ~n6059 ;
  assign n9076 = ~n9074 & n9075 ;
  assign n9081 = ~n2896 & ~n9076 ;
  assign n9082 = ~n9080 & n9081 ;
  assign n9083 = ~n9071 & ~n9082 ;
  assign n9084 = n2894 & ~n9083 ;
  assign n9085 = \P3_InstAddrPointer_reg[12]/NET0131  & n2820 ;
  assign n9086 = n2834 & ~n9085 ;
  assign n9087 = n2819 & n9086 ;
  assign n9088 = ~n2816 & ~n2819 ;
  assign n9089 = ~n2835 & ~n4058 ;
  assign n9090 = ~n9088 & n9089 ;
  assign n9091 = ~n9087 & ~n9090 ;
  assign n9092 = n8371 & ~n9091 ;
  assign n9093 = \P3_InstAddrPointer_reg[12]/NET0131  & ~n9092 ;
  assign n9094 = ~n2835 & ~n9086 ;
  assign n9095 = ~n2767 & ~n9094 ;
  assign n9096 = n4058 & ~n9095 ;
  assign n9100 = ~\P3_InstAddrPointer_reg[12]/NET0131  & ~n2847 ;
  assign n9101 = n9099 & ~n9100 ;
  assign n9102 = ~n2841 & n9101 ;
  assign n9103 = ~n2777 & n4166 ;
  assign n9112 = ~n9102 & ~n9103 ;
  assign n9113 = ~n9096 & n9112 ;
  assign n9114 = ~n9093 & n9113 ;
  assign n9115 = ~n9084 & n9114 ;
  assign n9116 = ~n9111 & n9115 ;
  assign n9117 = n2453 & ~n9116 ;
  assign n9069 = \P3_InstAddrPointer_reg[12]/NET0131  & ~n4418 ;
  assign n9070 = \P3_rEIP_reg[12]/NET0131  & n4412 ;
  assign n9118 = ~n9069 & ~n9070 ;
  assign n9119 = ~n9117 & n9118 ;
  assign n9121 = \P3_InstAddrPointer_reg[8]/NET0131  & n2896 ;
  assign n9130 = ~n4061 & n6086 ;
  assign n9129 = n4061 & ~n6086 ;
  assign n9131 = n3753 & ~n9129 ;
  assign n9132 = ~n9130 & n9131 ;
  assign n9122 = ~n4182 & ~n4224 ;
  assign n9123 = ~n4211 & ~n9122 ;
  assign n9124 = ~n3753 & ~n4178 ;
  assign n9125 = n9123 & n9124 ;
  assign n9126 = ~n4220 & n9125 ;
  assign n9127 = ~n3753 & n4220 ;
  assign n9128 = ~n6058 & n9127 ;
  assign n9133 = ~n9126 & ~n9128 ;
  assign n9134 = ~n9132 & n9133 ;
  assign n9135 = ~n2896 & ~n9134 ;
  assign n9136 = ~n9121 & ~n9135 ;
  assign n9137 = n2894 & ~n9136 ;
  assign n9147 = ~n4304 & n6124 ;
  assign n9148 = n2905 & ~n9104 ;
  assign n9149 = ~n9147 & n9148 ;
  assign n9138 = ~n2835 & ~n4061 ;
  assign n9139 = ~n2824 & ~n9138 ;
  assign n9140 = n7404 & ~n9139 ;
  assign n9141 = \P3_InstAddrPointer_reg[8]/NET0131  & ~n9140 ;
  assign n9146 = ~n2923 & n4061 ;
  assign n9142 = ~\P3_InstAddrPointer_reg[8]/NET0131  & ~n2847 ;
  assign n9143 = n4304 & ~n9142 ;
  assign n9144 = ~n2841 & n9143 ;
  assign n9145 = ~n2777 & n4220 ;
  assign n9150 = ~n9144 & ~n9145 ;
  assign n9151 = ~n9146 & n9150 ;
  assign n9152 = ~n9141 & n9151 ;
  assign n9153 = ~n9149 & n9152 ;
  assign n9154 = ~n9137 & n9153 ;
  assign n9155 = n2453 & ~n9154 ;
  assign n9120 = \P3_rEIP_reg[8]/NET0131  & n4412 ;
  assign n9156 = \P3_InstAddrPointer_reg[8]/NET0131  & ~n4418 ;
  assign n9157 = ~n9120 & ~n9156 ;
  assign n9158 = ~n9155 & n9157 ;
  assign n9162 = \P2_InstAddrPointer_reg[10]/NET0131  & n1897 ;
  assign n9167 = ~n6634 & n6639 ;
  assign n9168 = n6600 & ~n9167 ;
  assign n9169 = n7441 & n9168 ;
  assign n9170 = ~\P2_InstAddrPointer_reg[10]/NET0131  & ~n6496 ;
  assign n9171 = ~n6471 & ~n9170 ;
  assign n9172 = \P2_InstAddrPointer_reg[9]/NET0131  & n8443 ;
  assign n9173 = ~n9171 & ~n9172 ;
  assign n9174 = ~n9169 & ~n9173 ;
  assign n9175 = n6188 & ~n9174 ;
  assign n9163 = ~n6480 & n7430 ;
  assign n9164 = n6482 & ~n9163 ;
  assign n9165 = ~n6188 & ~n7431 ;
  assign n9166 = ~n9164 & n9165 ;
  assign n9176 = ~n1897 & ~n9166 ;
  assign n9177 = ~n9175 & n9176 ;
  assign n9178 = ~n9162 & ~n9177 ;
  assign n9179 = n1734 & ~n9178 ;
  assign n9181 = n6743 & n7546 ;
  assign n9180 = ~n6743 & ~n7546 ;
  assign n9182 = n1890 & ~n9180 ;
  assign n9183 = ~n9181 & n9182 ;
  assign n9161 = n1870 & n6743 ;
  assign n9184 = ~n1771 & n6482 ;
  assign n9187 = ~n9161 & ~n9184 ;
  assign n9185 = ~n1831 & n9171 ;
  assign n9186 = \P2_InstAddrPointer_reg[10]/NET0131  & ~n7501 ;
  assign n9188 = ~n9185 & ~n9186 ;
  assign n9189 = n9187 & n9188 ;
  assign n9190 = ~n9183 & n9189 ;
  assign n9191 = ~n9179 & n9190 ;
  assign n9192 = n1927 & ~n9191 ;
  assign n9159 = \P2_rEIP_reg[10]/NET0131  & n3113 ;
  assign n9160 = \P2_InstAddrPointer_reg[10]/NET0131  & ~n6810 ;
  assign n9193 = ~n9159 & ~n9160 ;
  assign n9194 = ~n9192 & n9193 ;
  assign n9204 = \P1_InstAddrPointer_reg[10]/NET0131  & n2375 ;
  assign n9205 = ~n4766 & ~n4772 ;
  assign n9206 = ~n6843 & ~n9205 ;
  assign n9207 = n4453 & ~n9206 ;
  assign n9208 = n4824 & ~n4874 ;
  assign n9209 = ~n4453 & ~n4875 ;
  assign n9210 = ~n9208 & n9209 ;
  assign n9211 = ~n2375 & ~n9210 ;
  assign n9212 = ~n9207 & n9211 ;
  assign n9213 = ~n9204 & ~n9212 ;
  assign n9214 = n2244 & ~n9213 ;
  assign n9199 = ~n5020 & ~n5023 ;
  assign n9200 = n2385 & ~n5024 ;
  assign n9201 = ~n9199 & n9200 ;
  assign n9203 = \P1_InstAddrPointer_reg[10]/NET0131  & ~n6027 ;
  assign n9202 = ~n2402 & n4772 ;
  assign n9197 = n2397 & n5023 ;
  assign n9198 = ~n2271 & n4824 ;
  assign n9215 = ~n9197 & ~n9198 ;
  assign n9216 = ~n9202 & n9215 ;
  assign n9217 = ~n9203 & n9216 ;
  assign n9218 = ~n9201 & n9217 ;
  assign n9219 = ~n9214 & n9218 ;
  assign n9220 = n2432 & ~n9219 ;
  assign n9195 = \P1_rEIP_reg[10]/NET0131  & n5092 ;
  assign n9196 = \P1_InstAddrPointer_reg[10]/NET0131  & ~n5098 ;
  assign n9221 = ~n9195 & ~n9196 ;
  assign n9222 = ~n9220 & n9221 ;
  assign n9228 = \P2_InstAddrPointer_reg[12]/NET0131  & n1897 ;
  assign n9225 = ~\P2_InstAddrPointer_reg[12]/NET0131  & ~n6497 ;
  assign n9226 = ~n6489 & ~n9225 ;
  assign n9233 = ~n8444 & n9226 ;
  assign n9232 = n8444 & ~n9226 ;
  assign n9234 = n6188 & ~n9232 ;
  assign n9235 = ~n9233 & n9234 ;
  assign n9229 = n6477 & ~n7602 ;
  assign n9230 = ~n6188 & ~n7515 ;
  assign n9231 = ~n9229 & n9230 ;
  assign n9236 = ~n1897 & ~n9231 ;
  assign n9237 = ~n9235 & n9236 ;
  assign n9238 = ~n9228 & ~n9237 ;
  assign n9239 = n1734 & ~n9238 ;
  assign n9240 = ~\P2_InstAddrPointer_reg[12]/NET0131  & ~n7490 ;
  assign n9241 = ~n6747 & ~n9240 ;
  assign n9242 = n7484 & n7491 ;
  assign n9243 = ~n7545 & n9242 ;
  assign n9245 = n9241 & n9243 ;
  assign n9244 = ~n9241 & ~n9243 ;
  assign n9246 = n1890 & ~n9244 ;
  assign n9247 = ~n9245 & n9246 ;
  assign n9248 = ~n1727 & ~n7490 ;
  assign n9249 = n7501 & ~n9248 ;
  assign n9250 = \P2_InstAddrPointer_reg[12]/NET0131  & ~n9249 ;
  assign n9252 = ~n1771 & n6477 ;
  assign n9227 = ~n1831 & n9226 ;
  assign n9251 = n1870 & n9241 ;
  assign n9253 = ~n9227 & ~n9251 ;
  assign n9254 = ~n9252 & n9253 ;
  assign n9255 = ~n9250 & n9254 ;
  assign n9256 = ~n9247 & n9255 ;
  assign n9257 = ~n9239 & n9256 ;
  assign n9258 = n1927 & ~n9257 ;
  assign n9223 = \P2_rEIP_reg[12]/NET0131  & n3113 ;
  assign n9224 = \P2_InstAddrPointer_reg[12]/NET0131  & ~n6810 ;
  assign n9259 = ~n9223 & ~n9224 ;
  assign n9260 = ~n9258 & n9259 ;
  assign n9264 = \P2_InstAddrPointer_reg[13]/NET0131  & n1897 ;
  assign n9268 = ~n6648 & ~n6653 ;
  assign n9269 = ~n7457 & ~n9268 ;
  assign n9270 = n6188 & ~n9269 ;
  assign n9265 = ~n6488 & n6518 ;
  assign n9266 = ~n6188 & ~n7603 ;
  assign n9267 = ~n9265 & n9266 ;
  assign n9271 = ~n1897 & ~n9267 ;
  assign n9272 = ~n9270 & n9271 ;
  assign n9273 = ~n9264 & ~n9272 ;
  assign n9274 = n1734 & ~n9273 ;
  assign n9275 = n6739 & n6744 ;
  assign n9276 = ~n7487 & ~n9275 ;
  assign n9277 = n1890 & ~n6746 ;
  assign n9278 = ~n9276 & n9277 ;
  assign n9263 = ~n1831 & n6653 ;
  assign n9281 = ~n1798 & n6747 ;
  assign n9282 = ~n1727 & ~n9281 ;
  assign n9283 = n7487 & n9282 ;
  assign n9284 = ~n9263 & ~n9283 ;
  assign n9279 = ~n1771 & n6518 ;
  assign n9280 = \P2_InstAddrPointer_reg[13]/NET0131  & ~n7501 ;
  assign n9285 = ~n9279 & ~n9280 ;
  assign n9286 = n9284 & n9285 ;
  assign n9287 = ~n9278 & n9286 ;
  assign n9288 = ~n9274 & n9287 ;
  assign n9289 = n1927 & ~n9288 ;
  assign n9261 = \P2_rEIP_reg[13]/NET0131  & n3113 ;
  assign n9262 = \P2_InstAddrPointer_reg[13]/NET0131  & ~n6810 ;
  assign n9290 = ~n9261 & ~n9262 ;
  assign n9291 = ~n9289 & n9290 ;
  assign n9294 = \P1_InstAddrPointer_reg[12]/NET0131  & n2375 ;
  assign n9299 = ~n6828 & ~n6830 ;
  assign n9300 = n6828 & n6830 ;
  assign n9301 = ~n9299 & ~n9300 ;
  assign n9302 = n4453 & ~n9301 ;
  assign n9295 = ~n4884 & ~n7273 ;
  assign n9296 = n4884 & n7273 ;
  assign n9297 = ~n9295 & ~n9296 ;
  assign n9298 = ~n4453 & ~n9297 ;
  assign n9303 = ~n2375 & ~n9298 ;
  assign n9304 = ~n9302 & n9303 ;
  assign n9305 = ~n9294 & ~n9304 ;
  assign n9306 = n2244 & ~n9305 ;
  assign n9307 = n5026 & n7299 ;
  assign n9311 = \P1_InstAddrPointer_reg[12]/NET0131  & n9307 ;
  assign n9308 = ~\P1_InstAddrPointer_reg[12]/NET0131  & ~n4963 ;
  assign n9309 = ~n4964 & ~n9308 ;
  assign n9310 = ~n9307 & ~n9309 ;
  assign n9312 = n2385 & ~n9310 ;
  assign n9313 = ~n9311 & n9312 ;
  assign n9317 = ~n2402 & n6830 ;
  assign n9314 = ~n2325 & ~n2369 ;
  assign n9315 = n2390 & n9314 ;
  assign n9316 = \P1_InstAddrPointer_reg[12]/NET0131  & ~n9315 ;
  assign n9293 = ~n2271 & n4884 ;
  assign n9318 = ~\P1_InstAddrPointer_reg[12]/NET0131  & ~n2337 ;
  assign n9319 = n2337 & ~n9309 ;
  assign n9320 = ~n9318 & ~n9319 ;
  assign n9321 = ~n2332 & n9320 ;
  assign n9322 = ~n9293 & ~n9321 ;
  assign n9323 = ~n9316 & n9322 ;
  assign n9324 = ~n9317 & n9323 ;
  assign n9325 = ~n9313 & n9324 ;
  assign n9326 = ~n9306 & n9325 ;
  assign n9327 = n2432 & ~n9326 ;
  assign n9292 = \P1_rEIP_reg[12]/NET0131  & n5092 ;
  assign n9328 = \P1_InstAddrPointer_reg[12]/NET0131  & ~n5098 ;
  assign n9329 = ~n9292 & ~n9328 ;
  assign n9330 = ~n9327 & n9329 ;
  assign n9336 = n5957 & n8550 ;
  assign n9338 = n4916 & n9336 ;
  assign n9337 = ~n4916 & ~n9336 ;
  assign n9339 = ~n4453 & ~n9337 ;
  assign n9340 = ~n9338 & n9339 ;
  assign n9341 = ~n5968 & ~n5973 ;
  assign n9342 = n4453 & ~n5974 ;
  assign n9343 = ~n9341 & n9342 ;
  assign n9344 = ~n9340 & ~n9343 ;
  assign n9345 = ~n2375 & ~n9344 ;
  assign n9346 = \P1_InstAddrPointer_reg[17]/NET0131  & n2375 ;
  assign n9347 = ~n9345 & ~n9346 ;
  assign n9348 = n2244 & ~n9347 ;
  assign n9333 = ~\P1_InstAddrPointer_reg[17]/NET0131  & ~n4966 ;
  assign n9334 = ~n4967 & ~n9333 ;
  assign n9352 = n5032 & n6010 ;
  assign n9354 = ~n9334 & ~n9352 ;
  assign n9353 = \P1_InstAddrPointer_reg[17]/NET0131  & n9352 ;
  assign n9355 = n2385 & ~n9353 ;
  assign n9356 = ~n9354 & n9355 ;
  assign n9349 = ~n2332 & ~n4966 ;
  assign n9350 = n6026 & ~n9349 ;
  assign n9351 = \P1_InstAddrPointer_reg[17]/NET0131  & ~n9350 ;
  assign n9359 = \P1_InstAddrPointer_reg[17]/NET0131  & n2317 ;
  assign n9360 = ~n2317 & n5968 ;
  assign n9361 = ~n9359 & ~n9360 ;
  assign n9362 = ~n2303 & ~n9361 ;
  assign n9363 = \P1_InstAddrPointer_reg[17]/NET0131  & ~n2387 ;
  assign n9364 = ~n2311 & n9360 ;
  assign n9365 = ~n9363 & ~n9364 ;
  assign n9366 = ~n2306 & ~n9365 ;
  assign n9367 = ~n9362 & ~n9366 ;
  assign n9368 = ~n2301 & ~n9367 ;
  assign n9358 = ~n2271 & n4916 ;
  assign n9335 = n2397 & n9334 ;
  assign n9357 = n2237 & n5968 ;
  assign n9369 = ~n9335 & ~n9357 ;
  assign n9370 = ~n9358 & n9369 ;
  assign n9371 = ~n9368 & n9370 ;
  assign n9372 = ~n9351 & n9371 ;
  assign n9373 = ~n9356 & n9372 ;
  assign n9374 = ~n9348 & n9373 ;
  assign n9375 = n2432 & ~n9374 ;
  assign n9331 = \P1_InstAddrPointer_reg[17]/NET0131  & ~n5098 ;
  assign n9332 = \P1_rEIP_reg[17]/NET0131  & n5092 ;
  assign n9376 = ~n9331 & ~n9332 ;
  assign n9377 = ~n9375 & n9376 ;
  assign n9383 = ~n5269 & n6908 ;
  assign n9384 = ~n6909 & ~n9383 ;
  assign n9385 = n5148 & n9384 ;
  assign n9386 = n5227 & ~n5277 ;
  assign n9387 = ~n6918 & ~n9386 ;
  assign n9388 = n5151 & n9387 ;
  assign n9389 = ~n9385 & ~n9388 ;
  assign n9390 = \P1_DataWidth_reg[1]/NET0131  & ~n9389 ;
  assign n9378 = ~n5108 & ~n5164 ;
  assign n9379 = \P1_InstQueue_reg[11][5]/NET0131  & ~n5104 ;
  assign n9380 = ~n5107 & n9379 ;
  assign n9381 = ~n9378 & ~n9380 ;
  assign n9391 = ~n5153 & ~n9381 ;
  assign n9392 = ~n9390 & ~n9391 ;
  assign n9393 = n2436 & ~n9392 ;
  assign n9382 = n5095 & ~n9381 ;
  assign n9394 = ~n2219 & n5104 ;
  assign n9395 = ~n9379 & ~n9394 ;
  assign n9396 = n3042 & ~n9395 ;
  assign n9397 = \P1_InstQueue_reg[11][5]/NET0131  & ~n5291 ;
  assign n9398 = ~n9396 & ~n9397 ;
  assign n9399 = ~n9382 & n9398 ;
  assign n9400 = ~n9393 & n9399 ;
  assign n9406 = ~n6909 & n6912 ;
  assign n9407 = ~n6913 & ~n9406 ;
  assign n9408 = n5148 & n9407 ;
  assign n9409 = n5221 & ~n6918 ;
  assign n9410 = ~n6919 & ~n9409 ;
  assign n9411 = n5151 & n9410 ;
  assign n9412 = ~n9408 & ~n9411 ;
  assign n9413 = \P1_DataWidth_reg[1]/NET0131  & ~n9412 ;
  assign n9401 = ~n5108 & ~n5182 ;
  assign n9402 = \P1_InstQueue_reg[11][6]/NET0131  & ~n5104 ;
  assign n9403 = ~n5107 & n9402 ;
  assign n9404 = ~n9401 & ~n9403 ;
  assign n9414 = ~n5153 & ~n9404 ;
  assign n9415 = ~n9413 & ~n9414 ;
  assign n9416 = n2436 & ~n9415 ;
  assign n9405 = n5095 & ~n9404 ;
  assign n9417 = ~n2125 & n5104 ;
  assign n9418 = ~n9402 & ~n9417 ;
  assign n9419 = n3042 & ~n9418 ;
  assign n9420 = \P1_InstQueue_reg[11][6]/NET0131  & ~n5291 ;
  assign n9421 = ~n9419 & ~n9420 ;
  assign n9422 = ~n9405 & n9421 ;
  assign n9423 = ~n9416 & n9422 ;
  assign n9429 = n5334 & n9384 ;
  assign n9430 = n5336 & n9387 ;
  assign n9431 = ~n9429 & ~n9430 ;
  assign n9432 = \P1_DataWidth_reg[1]/NET0131  & ~n9431 ;
  assign n9424 = ~n5164 & ~n5327 ;
  assign n9425 = \P1_InstQueue_reg[0][5]/NET0131  & ~n5324 ;
  assign n9426 = ~n5326 & n9425 ;
  assign n9427 = ~n9424 & ~n9426 ;
  assign n9433 = ~n5338 & ~n9427 ;
  assign n9434 = ~n9432 & ~n9433 ;
  assign n9435 = n2436 & ~n9434 ;
  assign n9428 = n5095 & ~n9427 ;
  assign n9436 = ~n2219 & n5324 ;
  assign n9437 = ~n9425 & ~n9436 ;
  assign n9438 = n3042 & ~n9437 ;
  assign n9439 = \P1_InstQueue_reg[0][5]/NET0131  & ~n5291 ;
  assign n9440 = ~n9438 & ~n9439 ;
  assign n9441 = ~n9428 & n9440 ;
  assign n9442 = ~n9435 & n9441 ;
  assign n9448 = n5334 & n9407 ;
  assign n9449 = n5336 & n9410 ;
  assign n9450 = ~n9448 & ~n9449 ;
  assign n9451 = \P1_DataWidth_reg[1]/NET0131  & ~n9450 ;
  assign n9443 = ~n5182 & ~n5327 ;
  assign n9444 = \P1_InstQueue_reg[0][6]/NET0131  & ~n5324 ;
  assign n9445 = ~n5326 & n9444 ;
  assign n9446 = ~n9443 & ~n9445 ;
  assign n9452 = ~n5338 & ~n9446 ;
  assign n9453 = ~n9451 & ~n9452 ;
  assign n9454 = n2436 & ~n9453 ;
  assign n9447 = n5095 & ~n9446 ;
  assign n9455 = ~n2125 & n5324 ;
  assign n9456 = ~n9444 & ~n9455 ;
  assign n9457 = n3042 & ~n9456 ;
  assign n9458 = \P1_InstQueue_reg[0][6]/NET0131  & ~n5291 ;
  assign n9459 = ~n9457 & ~n9458 ;
  assign n9460 = ~n9447 & n9459 ;
  assign n9461 = ~n9454 & n9460 ;
  assign n9467 = n5148 & n9387 ;
  assign n9468 = n5359 & n9384 ;
  assign n9469 = ~n9467 & ~n9468 ;
  assign n9470 = \P1_DataWidth_reg[1]/NET0131  & ~n9469 ;
  assign n9462 = ~n5164 & ~n5353 ;
  assign n9463 = \P1_InstQueue_reg[10][5]/NET0131  & ~n5107 ;
  assign n9464 = ~n5151 & n9463 ;
  assign n9465 = ~n9462 & ~n9464 ;
  assign n9471 = ~n5361 & ~n9465 ;
  assign n9472 = ~n9470 & ~n9471 ;
  assign n9473 = n2436 & ~n9472 ;
  assign n9466 = n5095 & ~n9465 ;
  assign n9474 = ~n2219 & n5107 ;
  assign n9475 = ~n9463 & ~n9474 ;
  assign n9476 = n3042 & ~n9475 ;
  assign n9477 = \P1_InstQueue_reg[10][5]/NET0131  & ~n5291 ;
  assign n9478 = ~n9476 & ~n9477 ;
  assign n9479 = ~n9466 & n9478 ;
  assign n9480 = ~n9473 & n9479 ;
  assign n9486 = n5148 & n9410 ;
  assign n9487 = n5359 & n9407 ;
  assign n9488 = ~n9486 & ~n9487 ;
  assign n9489 = \P1_DataWidth_reg[1]/NET0131  & ~n9488 ;
  assign n9481 = ~n5182 & ~n5353 ;
  assign n9482 = \P1_InstQueue_reg[10][6]/NET0131  & ~n5107 ;
  assign n9483 = ~n5151 & n9482 ;
  assign n9484 = ~n9481 & ~n9483 ;
  assign n9490 = ~n5361 & ~n9484 ;
  assign n9491 = ~n9489 & ~n9490 ;
  assign n9492 = n2436 & ~n9491 ;
  assign n9485 = n5095 & ~n9484 ;
  assign n9493 = ~n2125 & n5107 ;
  assign n9494 = ~n9482 & ~n9493 ;
  assign n9495 = n3042 & ~n9494 ;
  assign n9496 = \P1_InstQueue_reg[10][6]/NET0131  & ~n5291 ;
  assign n9497 = ~n9495 & ~n9496 ;
  assign n9498 = ~n9485 & n9497 ;
  assign n9499 = ~n9492 & n9498 ;
  assign n9505 = n5151 & n9384 ;
  assign n9506 = n5107 & n9387 ;
  assign n9507 = ~n9505 & ~n9506 ;
  assign n9508 = \P1_DataWidth_reg[1]/NET0131  & ~n9507 ;
  assign n9500 = ~n5164 & ~n5378 ;
  assign n9501 = \P1_InstQueue_reg[12][5]/NET0131  & ~n5377 ;
  assign n9502 = ~n5104 & n9501 ;
  assign n9503 = ~n9500 & ~n9502 ;
  assign n9509 = ~n5384 & ~n9503 ;
  assign n9510 = ~n9508 & ~n9509 ;
  assign n9511 = n2436 & ~n9510 ;
  assign n9504 = n5095 & ~n9503 ;
  assign n9512 = ~n2219 & n5377 ;
  assign n9513 = ~n9501 & ~n9512 ;
  assign n9514 = n3042 & ~n9513 ;
  assign n9515 = \P1_InstQueue_reg[12][5]/NET0131  & ~n5291 ;
  assign n9516 = ~n9514 & ~n9515 ;
  assign n9517 = ~n9504 & n9516 ;
  assign n9518 = ~n9511 & n9517 ;
  assign n9524 = n5151 & n9407 ;
  assign n9525 = n5107 & n9410 ;
  assign n9526 = ~n9524 & ~n9525 ;
  assign n9527 = \P1_DataWidth_reg[1]/NET0131  & ~n9526 ;
  assign n9519 = ~n5182 & ~n5378 ;
  assign n9520 = \P1_InstQueue_reg[12][6]/NET0131  & ~n5377 ;
  assign n9521 = ~n5104 & n9520 ;
  assign n9522 = ~n9519 & ~n9521 ;
  assign n9528 = ~n5384 & ~n9522 ;
  assign n9529 = ~n9527 & ~n9528 ;
  assign n9530 = n2436 & ~n9529 ;
  assign n9523 = n5095 & ~n9522 ;
  assign n9531 = ~n2125 & n5377 ;
  assign n9532 = ~n9520 & ~n9531 ;
  assign n9533 = n3042 & ~n9532 ;
  assign n9534 = \P1_InstQueue_reg[12][6]/NET0131  & ~n5291 ;
  assign n9535 = ~n9533 & ~n9534 ;
  assign n9536 = ~n9523 & n9535 ;
  assign n9537 = ~n9530 & n9536 ;
  assign n9543 = n5107 & n9384 ;
  assign n9544 = n5104 & n9387 ;
  assign n9545 = ~n9543 & ~n9544 ;
  assign n9546 = \P1_DataWidth_reg[1]/NET0131  & ~n9545 ;
  assign n9538 = ~n5164 & ~n5399 ;
  assign n9539 = \P1_InstQueue_reg[13][5]/NET0131  & ~n5334 ;
  assign n9540 = ~n5377 & n9539 ;
  assign n9541 = ~n9538 & ~n9540 ;
  assign n9547 = ~n5405 & ~n9541 ;
  assign n9548 = ~n9546 & ~n9547 ;
  assign n9549 = n2436 & ~n9548 ;
  assign n9542 = n5095 & ~n9541 ;
  assign n9550 = ~n2219 & n5334 ;
  assign n9551 = ~n9539 & ~n9550 ;
  assign n9552 = n3042 & ~n9551 ;
  assign n9553 = \P1_InstQueue_reg[13][5]/NET0131  & ~n5291 ;
  assign n9554 = ~n9552 & ~n9553 ;
  assign n9555 = ~n9542 & n9554 ;
  assign n9556 = ~n9549 & n9555 ;
  assign n9562 = n5107 & n9407 ;
  assign n9563 = n5104 & n9410 ;
  assign n9564 = ~n9562 & ~n9563 ;
  assign n9565 = \P1_DataWidth_reg[1]/NET0131  & ~n9564 ;
  assign n9557 = ~n5182 & ~n5399 ;
  assign n9558 = \P1_InstQueue_reg[13][6]/NET0131  & ~n5334 ;
  assign n9559 = ~n5377 & n9558 ;
  assign n9560 = ~n9557 & ~n9559 ;
  assign n9566 = ~n5405 & ~n9560 ;
  assign n9567 = ~n9565 & ~n9566 ;
  assign n9568 = n2436 & ~n9567 ;
  assign n9561 = n5095 & ~n9560 ;
  assign n9569 = ~n2125 & n5334 ;
  assign n9570 = ~n9558 & ~n9569 ;
  assign n9571 = n3042 & ~n9570 ;
  assign n9572 = \P1_InstQueue_reg[13][6]/NET0131  & ~n5291 ;
  assign n9573 = ~n9571 & ~n9572 ;
  assign n9574 = ~n9561 & n9573 ;
  assign n9575 = ~n9568 & n9574 ;
  assign n9581 = n5104 & n9384 ;
  assign n9582 = n5377 & n9387 ;
  assign n9583 = ~n9581 & ~n9582 ;
  assign n9584 = \P1_DataWidth_reg[1]/NET0131  & ~n9583 ;
  assign n9576 = ~n5164 & ~n5337 ;
  assign n9577 = \P1_InstQueue_reg[14][5]/NET0131  & ~n5336 ;
  assign n9578 = ~n5334 & n9577 ;
  assign n9579 = ~n9576 & ~n9578 ;
  assign n9585 = ~n5425 & ~n9579 ;
  assign n9586 = ~n9584 & ~n9585 ;
  assign n9587 = n2436 & ~n9586 ;
  assign n9580 = n5095 & ~n9579 ;
  assign n9588 = ~n2219 & n5336 ;
  assign n9589 = ~n9577 & ~n9588 ;
  assign n9590 = n3042 & ~n9589 ;
  assign n9591 = \P1_InstQueue_reg[14][5]/NET0131  & ~n5291 ;
  assign n9592 = ~n9590 & ~n9591 ;
  assign n9593 = ~n9580 & n9592 ;
  assign n9594 = ~n9587 & n9593 ;
  assign n9600 = n5104 & n9407 ;
  assign n9601 = n5377 & n9410 ;
  assign n9602 = ~n9600 & ~n9601 ;
  assign n9603 = \P1_DataWidth_reg[1]/NET0131  & ~n9602 ;
  assign n9595 = ~n5182 & ~n5337 ;
  assign n9596 = \P1_InstQueue_reg[14][6]/NET0131  & ~n5336 ;
  assign n9597 = ~n5334 & n9596 ;
  assign n9598 = ~n9595 & ~n9597 ;
  assign n9604 = ~n5425 & ~n9598 ;
  assign n9605 = ~n9603 & ~n9604 ;
  assign n9606 = n2436 & ~n9605 ;
  assign n9599 = n5095 & ~n9598 ;
  assign n9607 = ~n2125 & n5336 ;
  assign n9608 = ~n9596 & ~n9607 ;
  assign n9609 = n3042 & ~n9608 ;
  assign n9610 = \P1_InstQueue_reg[14][6]/NET0131  & ~n5291 ;
  assign n9611 = ~n9609 & ~n9610 ;
  assign n9612 = ~n9599 & n9611 ;
  assign n9613 = ~n9606 & n9612 ;
  assign n9619 = n5377 & n9384 ;
  assign n9620 = n5334 & n9387 ;
  assign n9621 = ~n9619 & ~n9620 ;
  assign n9622 = \P1_DataWidth_reg[1]/NET0131  & ~n9621 ;
  assign n9614 = ~n5164 & ~n5440 ;
  assign n9615 = \P1_InstQueue_reg[15][5]/NET0131  & ~n5326 ;
  assign n9616 = ~n5336 & n9615 ;
  assign n9617 = ~n9614 & ~n9616 ;
  assign n9623 = ~n5446 & ~n9617 ;
  assign n9624 = ~n9622 & ~n9623 ;
  assign n9625 = n2436 & ~n9624 ;
  assign n9618 = n5095 & ~n9617 ;
  assign n9626 = ~n2219 & n5326 ;
  assign n9627 = ~n9615 & ~n9626 ;
  assign n9628 = n3042 & ~n9627 ;
  assign n9629 = \P1_InstQueue_reg[15][5]/NET0131  & ~n5291 ;
  assign n9630 = ~n9628 & ~n9629 ;
  assign n9631 = ~n9618 & n9630 ;
  assign n9632 = ~n9625 & n9631 ;
  assign n9638 = n5377 & n9407 ;
  assign n9639 = n5334 & n9410 ;
  assign n9640 = ~n9638 & ~n9639 ;
  assign n9641 = \P1_DataWidth_reg[1]/NET0131  & ~n9640 ;
  assign n9633 = ~n5182 & ~n5440 ;
  assign n9634 = \P1_InstQueue_reg[15][6]/NET0131  & ~n5326 ;
  assign n9635 = ~n5336 & n9634 ;
  assign n9636 = ~n9633 & ~n9635 ;
  assign n9642 = ~n5446 & ~n9636 ;
  assign n9643 = ~n9641 & ~n9642 ;
  assign n9644 = n2436 & ~n9643 ;
  assign n9637 = n5095 & ~n9636 ;
  assign n9645 = ~n2125 & n5326 ;
  assign n9646 = ~n9634 & ~n9645 ;
  assign n9647 = n3042 & ~n9646 ;
  assign n9648 = \P1_InstQueue_reg[15][6]/NET0131  & ~n5291 ;
  assign n9649 = ~n9647 & ~n9648 ;
  assign n9650 = ~n9637 & n9649 ;
  assign n9651 = ~n9644 & n9650 ;
  assign n9657 = n5336 & n9384 ;
  assign n9658 = n5326 & n9387 ;
  assign n9659 = ~n9657 & ~n9658 ;
  assign n9660 = \P1_DataWidth_reg[1]/NET0131  & ~n9659 ;
  assign n9652 = ~n5164 & ~n5462 ;
  assign n9653 = \P1_InstQueue_reg[1][5]/NET0131  & ~n5461 ;
  assign n9654 = ~n5324 & n9653 ;
  assign n9655 = ~n9652 & ~n9654 ;
  assign n9661 = ~n5468 & ~n9655 ;
  assign n9662 = ~n9660 & ~n9661 ;
  assign n9663 = n2436 & ~n9662 ;
  assign n9656 = n5095 & ~n9655 ;
  assign n9664 = ~n2219 & n5461 ;
  assign n9665 = ~n9653 & ~n9664 ;
  assign n9666 = n3042 & ~n9665 ;
  assign n9667 = \P1_InstQueue_reg[1][5]/NET0131  & ~n5291 ;
  assign n9668 = ~n9666 & ~n9667 ;
  assign n9669 = ~n9656 & n9668 ;
  assign n9670 = ~n9663 & n9669 ;
  assign n9676 = n5336 & n9407 ;
  assign n9677 = n5326 & n9410 ;
  assign n9678 = ~n9676 & ~n9677 ;
  assign n9679 = \P1_DataWidth_reg[1]/NET0131  & ~n9678 ;
  assign n9671 = ~n5182 & ~n5462 ;
  assign n9672 = \P1_InstQueue_reg[1][6]/NET0131  & ~n5461 ;
  assign n9673 = ~n5324 & n9672 ;
  assign n9674 = ~n9671 & ~n9673 ;
  assign n9680 = ~n5468 & ~n9674 ;
  assign n9681 = ~n9679 & ~n9680 ;
  assign n9682 = n2436 & ~n9681 ;
  assign n9675 = n5095 & ~n9674 ;
  assign n9683 = ~n2125 & n5461 ;
  assign n9684 = ~n9672 & ~n9683 ;
  assign n9685 = n3042 & ~n9684 ;
  assign n9686 = \P1_InstQueue_reg[1][6]/NET0131  & ~n5291 ;
  assign n9687 = ~n9685 & ~n9686 ;
  assign n9688 = ~n9675 & n9687 ;
  assign n9689 = ~n9682 & n9688 ;
  assign n9695 = n5324 & n9387 ;
  assign n9696 = n5326 & n9384 ;
  assign n9697 = ~n9695 & ~n9696 ;
  assign n9698 = \P1_DataWidth_reg[1]/NET0131  & ~n9697 ;
  assign n9690 = ~n5164 & ~n5506 ;
  assign n9691 = \P1_InstQueue_reg[2][5]/NET0131  & ~n5484 ;
  assign n9692 = ~n5461 & n9691 ;
  assign n9693 = ~n9690 & ~n9692 ;
  assign n9699 = ~n5512 & ~n9693 ;
  assign n9700 = ~n9698 & ~n9699 ;
  assign n9701 = n2436 & ~n9700 ;
  assign n9694 = n5095 & ~n9693 ;
  assign n9702 = ~n2219 & n5484 ;
  assign n9703 = ~n9691 & ~n9702 ;
  assign n9704 = n3042 & ~n9703 ;
  assign n9705 = \P1_InstQueue_reg[2][5]/NET0131  & ~n5291 ;
  assign n9706 = ~n9704 & ~n9705 ;
  assign n9707 = ~n9694 & n9706 ;
  assign n9708 = ~n9701 & n9707 ;
  assign n9714 = n5324 & n9410 ;
  assign n9715 = n5326 & n9407 ;
  assign n9716 = ~n9714 & ~n9715 ;
  assign n9717 = \P1_DataWidth_reg[1]/NET0131  & ~n9716 ;
  assign n9709 = ~n5182 & ~n5506 ;
  assign n9710 = \P1_InstQueue_reg[2][6]/NET0131  & ~n5484 ;
  assign n9711 = ~n5461 & n9710 ;
  assign n9712 = ~n9709 & ~n9711 ;
  assign n9718 = ~n5512 & ~n9712 ;
  assign n9719 = ~n9717 & ~n9718 ;
  assign n9720 = n2436 & ~n9719 ;
  assign n9713 = n5095 & ~n9712 ;
  assign n9721 = ~n2125 & n5484 ;
  assign n9722 = ~n9710 & ~n9721 ;
  assign n9723 = n3042 & ~n9722 ;
  assign n9724 = \P1_InstQueue_reg[2][6]/NET0131  & ~n5291 ;
  assign n9725 = ~n9723 & ~n9724 ;
  assign n9726 = ~n9713 & n9725 ;
  assign n9727 = ~n9720 & n9726 ;
  assign n9733 = n5324 & n9384 ;
  assign n9734 = n5461 & n9387 ;
  assign n9735 = ~n9733 & ~n9734 ;
  assign n9736 = \P1_DataWidth_reg[1]/NET0131  & ~n9735 ;
  assign n9728 = ~n5164 & ~n5485 ;
  assign n9729 = \P1_InstQueue_reg[3][5]/NET0131  & ~n5483 ;
  assign n9730 = ~n5484 & n9729 ;
  assign n9731 = ~n9728 & ~n9730 ;
  assign n9737 = ~n5491 & ~n9731 ;
  assign n9738 = ~n9736 & ~n9737 ;
  assign n9739 = n2436 & ~n9738 ;
  assign n9732 = n5095 & ~n9731 ;
  assign n9740 = ~n2219 & n5483 ;
  assign n9741 = ~n9729 & ~n9740 ;
  assign n9742 = n3042 & ~n9741 ;
  assign n9743 = \P1_InstQueue_reg[3][5]/NET0131  & ~n5291 ;
  assign n9744 = ~n9742 & ~n9743 ;
  assign n9745 = ~n9732 & n9744 ;
  assign n9746 = ~n9739 & n9745 ;
  assign n9752 = n5324 & n9407 ;
  assign n9753 = n5461 & n9410 ;
  assign n9754 = ~n9752 & ~n9753 ;
  assign n9755 = \P1_DataWidth_reg[1]/NET0131  & ~n9754 ;
  assign n9747 = ~n5182 & ~n5485 ;
  assign n9748 = \P1_InstQueue_reg[3][6]/NET0131  & ~n5483 ;
  assign n9749 = ~n5484 & n9748 ;
  assign n9750 = ~n9747 & ~n9749 ;
  assign n9756 = ~n5491 & ~n9750 ;
  assign n9757 = ~n9755 & ~n9756 ;
  assign n9758 = n2436 & ~n9757 ;
  assign n9751 = n5095 & ~n9750 ;
  assign n9759 = ~n2125 & n5483 ;
  assign n9760 = ~n9748 & ~n9759 ;
  assign n9761 = n3042 & ~n9760 ;
  assign n9762 = \P1_InstQueue_reg[3][6]/NET0131  & ~n5291 ;
  assign n9763 = ~n9761 & ~n9762 ;
  assign n9764 = ~n9751 & n9763 ;
  assign n9765 = ~n9758 & n9764 ;
  assign n9771 = n5461 & n9384 ;
  assign n9772 = n5484 & n9387 ;
  assign n9773 = ~n9771 & ~n9772 ;
  assign n9774 = \P1_DataWidth_reg[1]/NET0131  & ~n9773 ;
  assign n9766 = ~n5164 & ~n5528 ;
  assign n9767 = \P1_InstQueue_reg[4][5]/NET0131  & ~n5527 ;
  assign n9768 = ~n5483 & n9767 ;
  assign n9769 = ~n9766 & ~n9768 ;
  assign n9775 = ~n5534 & ~n9769 ;
  assign n9776 = ~n9774 & ~n9775 ;
  assign n9777 = n2436 & ~n9776 ;
  assign n9770 = n5095 & ~n9769 ;
  assign n9778 = ~n2219 & n5527 ;
  assign n9779 = ~n9767 & ~n9778 ;
  assign n9780 = n3042 & ~n9779 ;
  assign n9781 = \P1_InstQueue_reg[4][5]/NET0131  & ~n5291 ;
  assign n9782 = ~n9780 & ~n9781 ;
  assign n9783 = ~n9770 & n9782 ;
  assign n9784 = ~n9777 & n9783 ;
  assign n9790 = n5461 & n9407 ;
  assign n9791 = n5484 & n9410 ;
  assign n9792 = ~n9790 & ~n9791 ;
  assign n9793 = \P1_DataWidth_reg[1]/NET0131  & ~n9792 ;
  assign n9785 = ~n5182 & ~n5528 ;
  assign n9786 = \P1_InstQueue_reg[4][6]/NET0131  & ~n5527 ;
  assign n9787 = ~n5483 & n9786 ;
  assign n9788 = ~n9785 & ~n9787 ;
  assign n9794 = ~n5534 & ~n9788 ;
  assign n9795 = ~n9793 & ~n9794 ;
  assign n9796 = n2436 & ~n9795 ;
  assign n9789 = n5095 & ~n9788 ;
  assign n9797 = ~n2125 & n5527 ;
  assign n9798 = ~n9786 & ~n9797 ;
  assign n9799 = n3042 & ~n9798 ;
  assign n9800 = \P1_InstQueue_reg[4][6]/NET0131  & ~n5291 ;
  assign n9801 = ~n9799 & ~n9800 ;
  assign n9802 = ~n9789 & n9801 ;
  assign n9803 = ~n9796 & n9802 ;
  assign n9809 = n5484 & n9384 ;
  assign n9810 = n5483 & n9387 ;
  assign n9811 = ~n9809 & ~n9810 ;
  assign n9812 = \P1_DataWidth_reg[1]/NET0131  & ~n9811 ;
  assign n9804 = ~n5164 & ~n5550 ;
  assign n9805 = \P1_InstQueue_reg[5][5]/NET0131  & ~n5549 ;
  assign n9806 = ~n5527 & n9805 ;
  assign n9807 = ~n9804 & ~n9806 ;
  assign n9813 = ~n5556 & ~n9807 ;
  assign n9814 = ~n9812 & ~n9813 ;
  assign n9815 = n2436 & ~n9814 ;
  assign n9808 = n5095 & ~n9807 ;
  assign n9816 = ~n2219 & n5549 ;
  assign n9817 = ~n9805 & ~n9816 ;
  assign n9818 = n3042 & ~n9817 ;
  assign n9819 = \P1_InstQueue_reg[5][5]/NET0131  & ~n5291 ;
  assign n9820 = ~n9818 & ~n9819 ;
  assign n9821 = ~n9808 & n9820 ;
  assign n9822 = ~n9815 & n9821 ;
  assign n9828 = n5484 & n9407 ;
  assign n9829 = n5483 & n9410 ;
  assign n9830 = ~n9828 & ~n9829 ;
  assign n9831 = \P1_DataWidth_reg[1]/NET0131  & ~n9830 ;
  assign n9823 = ~n5182 & ~n5550 ;
  assign n9824 = \P1_InstQueue_reg[5][6]/NET0131  & ~n5549 ;
  assign n9825 = ~n5527 & n9824 ;
  assign n9826 = ~n9823 & ~n9825 ;
  assign n9832 = ~n5556 & ~n9826 ;
  assign n9833 = ~n9831 & ~n9832 ;
  assign n9834 = n2436 & ~n9833 ;
  assign n9827 = n5095 & ~n9826 ;
  assign n9835 = ~n2125 & n5549 ;
  assign n9836 = ~n9824 & ~n9835 ;
  assign n9837 = n3042 & ~n9836 ;
  assign n9838 = \P1_InstQueue_reg[5][6]/NET0131  & ~n5291 ;
  assign n9839 = ~n9837 & ~n9838 ;
  assign n9840 = ~n9827 & n9839 ;
  assign n9841 = ~n9834 & n9840 ;
  assign n9847 = n5483 & n9384 ;
  assign n9848 = n5527 & n9387 ;
  assign n9849 = ~n9847 & ~n9848 ;
  assign n9850 = \P1_DataWidth_reg[1]/NET0131  & ~n9849 ;
  assign n9842 = ~n5164 & ~n5572 ;
  assign n9843 = \P1_InstQueue_reg[6][5]/NET0131  & ~n5571 ;
  assign n9844 = ~n5549 & n9843 ;
  assign n9845 = ~n9842 & ~n9844 ;
  assign n9851 = ~n5578 & ~n9845 ;
  assign n9852 = ~n9850 & ~n9851 ;
  assign n9853 = n2436 & ~n9852 ;
  assign n9846 = n5095 & ~n9845 ;
  assign n9854 = ~n2219 & n5571 ;
  assign n9855 = ~n9843 & ~n9854 ;
  assign n9856 = n3042 & ~n9855 ;
  assign n9857 = \P1_InstQueue_reg[6][5]/NET0131  & ~n5291 ;
  assign n9858 = ~n9856 & ~n9857 ;
  assign n9859 = ~n9846 & n9858 ;
  assign n9860 = ~n9853 & n9859 ;
  assign n9866 = n5483 & n9407 ;
  assign n9867 = n5527 & n9410 ;
  assign n9868 = ~n9866 & ~n9867 ;
  assign n9869 = \P1_DataWidth_reg[1]/NET0131  & ~n9868 ;
  assign n9861 = ~n5182 & ~n5572 ;
  assign n9862 = \P1_InstQueue_reg[6][6]/NET0131  & ~n5571 ;
  assign n9863 = ~n5549 & n9862 ;
  assign n9864 = ~n9861 & ~n9863 ;
  assign n9870 = ~n5578 & ~n9864 ;
  assign n9871 = ~n9869 & ~n9870 ;
  assign n9872 = n2436 & ~n9871 ;
  assign n9865 = n5095 & ~n9864 ;
  assign n9873 = ~n2125 & n5571 ;
  assign n9874 = ~n9862 & ~n9873 ;
  assign n9875 = n3042 & ~n9874 ;
  assign n9876 = \P1_InstQueue_reg[6][6]/NET0131  & ~n5291 ;
  assign n9877 = ~n9875 & ~n9876 ;
  assign n9878 = ~n9865 & n9877 ;
  assign n9879 = ~n9872 & n9878 ;
  assign n9885 = n5527 & n9384 ;
  assign n9886 = n5549 & n9387 ;
  assign n9887 = ~n9885 & ~n9886 ;
  assign n9888 = \P1_DataWidth_reg[1]/NET0131  & ~n9887 ;
  assign n9880 = ~n5164 & ~n5593 ;
  assign n9881 = \P1_InstQueue_reg[7][5]/NET0131  & ~n5359 ;
  assign n9882 = ~n5571 & n9881 ;
  assign n9883 = ~n9880 & ~n9882 ;
  assign n9889 = ~n5599 & ~n9883 ;
  assign n9890 = ~n9888 & ~n9889 ;
  assign n9891 = n2436 & ~n9890 ;
  assign n9884 = n5095 & ~n9883 ;
  assign n9892 = ~n2219 & n5359 ;
  assign n9893 = ~n9881 & ~n9892 ;
  assign n9894 = n3042 & ~n9893 ;
  assign n9895 = \P1_InstQueue_reg[7][5]/NET0131  & ~n5291 ;
  assign n9896 = ~n9894 & ~n9895 ;
  assign n9897 = ~n9884 & n9896 ;
  assign n9898 = ~n9891 & n9897 ;
  assign n9904 = n5527 & n9407 ;
  assign n9905 = n5549 & n9410 ;
  assign n9906 = ~n9904 & ~n9905 ;
  assign n9907 = \P1_DataWidth_reg[1]/NET0131  & ~n9906 ;
  assign n9899 = ~n5182 & ~n5593 ;
  assign n9900 = \P1_InstQueue_reg[7][6]/NET0131  & ~n5359 ;
  assign n9901 = ~n5571 & n9900 ;
  assign n9902 = ~n9899 & ~n9901 ;
  assign n9908 = ~n5599 & ~n9902 ;
  assign n9909 = ~n9907 & ~n9908 ;
  assign n9910 = n2436 & ~n9909 ;
  assign n9903 = n5095 & ~n9902 ;
  assign n9911 = ~n2125 & n5359 ;
  assign n9912 = ~n9900 & ~n9911 ;
  assign n9913 = n3042 & ~n9912 ;
  assign n9914 = \P1_InstQueue_reg[7][6]/NET0131  & ~n5291 ;
  assign n9915 = ~n9913 & ~n9914 ;
  assign n9916 = ~n9903 & n9915 ;
  assign n9917 = ~n9910 & n9916 ;
  assign n9923 = n5549 & n9384 ;
  assign n9924 = n5571 & n9387 ;
  assign n9925 = ~n9923 & ~n9924 ;
  assign n9926 = \P1_DataWidth_reg[1]/NET0131  & ~n9925 ;
  assign n9918 = ~n5164 & ~n5360 ;
  assign n9919 = \P1_InstQueue_reg[8][5]/NET0131  & ~n5148 ;
  assign n9920 = ~n5359 & n9919 ;
  assign n9921 = ~n9918 & ~n9920 ;
  assign n9927 = ~n5619 & ~n9921 ;
  assign n9928 = ~n9926 & ~n9927 ;
  assign n9929 = n2436 & ~n9928 ;
  assign n9922 = n5095 & ~n9921 ;
  assign n9930 = ~n2219 & n5148 ;
  assign n9931 = ~n9919 & ~n9930 ;
  assign n9932 = n3042 & ~n9931 ;
  assign n9933 = \P1_InstQueue_reg[8][5]/NET0131  & ~n5291 ;
  assign n9934 = ~n9932 & ~n9933 ;
  assign n9935 = ~n9922 & n9934 ;
  assign n9936 = ~n9929 & n9935 ;
  assign n9942 = n5549 & n9407 ;
  assign n9943 = n5571 & n9410 ;
  assign n9944 = ~n9942 & ~n9943 ;
  assign n9945 = \P1_DataWidth_reg[1]/NET0131  & ~n9944 ;
  assign n9937 = ~n5182 & ~n5360 ;
  assign n9938 = \P1_InstQueue_reg[8][6]/NET0131  & ~n5148 ;
  assign n9939 = ~n5359 & n9938 ;
  assign n9940 = ~n9937 & ~n9939 ;
  assign n9946 = ~n5619 & ~n9940 ;
  assign n9947 = ~n9945 & ~n9946 ;
  assign n9948 = n2436 & ~n9947 ;
  assign n9941 = n5095 & ~n9940 ;
  assign n9949 = ~n2125 & n5148 ;
  assign n9950 = ~n9938 & ~n9949 ;
  assign n9951 = n3042 & ~n9950 ;
  assign n9952 = \P1_InstQueue_reg[8][6]/NET0131  & ~n5291 ;
  assign n9953 = ~n9951 & ~n9952 ;
  assign n9954 = ~n9941 & n9953 ;
  assign n9955 = ~n9948 & n9954 ;
  assign n9961 = n5571 & n9384 ;
  assign n9962 = n5359 & n9387 ;
  assign n9963 = ~n9961 & ~n9962 ;
  assign n9964 = \P1_DataWidth_reg[1]/NET0131  & ~n9963 ;
  assign n9956 = ~n5152 & ~n5164 ;
  assign n9957 = \P1_InstQueue_reg[9][5]/NET0131  & ~n5151 ;
  assign n9958 = ~n5148 & n9957 ;
  assign n9959 = ~n9956 & ~n9958 ;
  assign n9965 = ~n5639 & ~n9959 ;
  assign n9966 = ~n9964 & ~n9965 ;
  assign n9967 = n2436 & ~n9966 ;
  assign n9960 = n5095 & ~n9959 ;
  assign n9968 = ~n2219 & n5151 ;
  assign n9969 = ~n9957 & ~n9968 ;
  assign n9970 = n3042 & ~n9969 ;
  assign n9971 = \P1_InstQueue_reg[9][5]/NET0131  & ~n5291 ;
  assign n9972 = ~n9970 & ~n9971 ;
  assign n9973 = ~n9960 & n9972 ;
  assign n9974 = ~n9967 & n9973 ;
  assign n9980 = n5571 & n9407 ;
  assign n9981 = n5359 & n9410 ;
  assign n9982 = ~n9980 & ~n9981 ;
  assign n9983 = \P1_DataWidth_reg[1]/NET0131  & ~n9982 ;
  assign n9975 = ~n5152 & ~n5182 ;
  assign n9976 = \P1_InstQueue_reg[9][6]/NET0131  & ~n5151 ;
  assign n9977 = ~n5148 & n9976 ;
  assign n9978 = ~n9975 & ~n9977 ;
  assign n9984 = ~n5639 & ~n9978 ;
  assign n9985 = ~n9983 & ~n9984 ;
  assign n9986 = n2436 & ~n9985 ;
  assign n9979 = n5095 & ~n9978 ;
  assign n9987 = ~n2125 & n5151 ;
  assign n9988 = ~n9976 & ~n9987 ;
  assign n9989 = n3042 & ~n9988 ;
  assign n9990 = \P1_InstQueue_reg[9][6]/NET0131  & ~n5291 ;
  assign n9991 = ~n9989 & ~n9990 ;
  assign n9992 = ~n9979 & n9991 ;
  assign n9993 = ~n9986 & n9992 ;
  assign n9994 = \P2_PhyAddrPointer_reg[30]/NET0131  & n1897 ;
  assign n10004 = n7608 & n8920 ;
  assign n10006 = ~n8919 & n10004 ;
  assign n10005 = n8919 & ~n10004 ;
  assign n10007 = ~n6188 & ~n10005 ;
  assign n10008 = ~n10006 & n10007 ;
  assign n9995 = ~\P2_InstAddrPointer_reg[30]/NET0131  & ~n6586 ;
  assign n9996 = ~n8904 & ~n9995 ;
  assign n9997 = \P2_InstAddrPointer_reg[29]/NET0131  & n6598 ;
  assign n9998 = n6678 & n9997 ;
  assign n9999 = n7527 & n9998 ;
  assign n10001 = n9996 & ~n9999 ;
  assign n10000 = ~n9996 & n9999 ;
  assign n10002 = n6188 & ~n10000 ;
  assign n10003 = ~n10001 & n10002 ;
  assign n10009 = ~n1897 & ~n10003 ;
  assign n10010 = ~n10008 & n10009 ;
  assign n10011 = ~n9994 & ~n10010 ;
  assign n10012 = n1734 & ~n10011 ;
  assign n10013 = \P2_PhyAddrPointer_reg[30]/NET0131  & ~n8936 ;
  assign n10014 = ~\P2_InstAddrPointer_reg[30]/NET0131  & ~n6786 ;
  assign n10015 = ~n8946 & ~n10014 ;
  assign n10016 = \P2_InstAddrPointer_reg[29]/NET0131  & n6779 ;
  assign n10017 = n7628 & n10016 ;
  assign n10018 = ~n10015 & ~n10017 ;
  assign n10019 = n7628 & n8944 ;
  assign n10020 = n1890 & ~n10019 ;
  assign n10021 = ~n10018 & n10020 ;
  assign n10022 = ~n10013 & ~n10021 ;
  assign n10023 = ~n10012 & n10022 ;
  assign n10024 = n1927 & ~n10023 ;
  assign n10025 = ~\P2_PhyAddrPointer_reg[30]/NET0131  & ~n8986 ;
  assign n10026 = n3034 & ~n8987 ;
  assign n10027 = ~n10025 & n10026 ;
  assign n10028 = ~\P2_PhyAddrPointer_reg[30]/NET0131  & ~n8999 ;
  assign n10029 = ~n9000 & ~n10028 ;
  assign n10030 = n9005 & n10029 ;
  assign n10031 = \P2_rEIP_reg[30]/NET0131  & n3113 ;
  assign n10032 = \P2_PhyAddrPointer_reg[30]/NET0131  & ~n8958 ;
  assign n10033 = ~n10031 & ~n10032 ;
  assign n10034 = ~n10030 & n10033 ;
  assign n10035 = ~n10027 & n10034 ;
  assign n10036 = ~n10024 & n10035 ;
  assign n10037 = \P3_PhyAddrPointer_reg[30]/NET0131  & n2896 ;
  assign n10047 = n4100 & n7381 ;
  assign n10048 = n8402 & n10047 ;
  assign n10049 = n7382 & n10048 ;
  assign n10050 = n4093 & n4114 ;
  assign n10051 = n10049 & n10050 ;
  assign n10053 = n4120 & n10051 ;
  assign n10052 = ~n4120 & ~n10051 ;
  assign n10054 = n3753 & ~n10052 ;
  assign n10055 = ~n10053 & n10054 ;
  assign n10038 = n4275 & n7369 ;
  assign n10039 = n7373 & n10038 ;
  assign n10040 = n7371 & n10039 ;
  assign n10041 = ~n4277 & n10040 ;
  assign n10042 = n4147 & n10041 ;
  assign n10043 = n4153 & ~n10042 ;
  assign n10044 = n4154 & n10041 ;
  assign n10045 = ~n3753 & ~n10044 ;
  assign n10046 = ~n10043 & n10045 ;
  assign n10056 = ~n2896 & ~n10046 ;
  assign n10057 = ~n10055 & n10056 ;
  assign n10058 = ~n10037 & ~n10057 ;
  assign n10059 = n2894 & ~n10058 ;
  assign n10060 = \P3_PhyAddrPointer_reg[30]/NET0131  & ~n9014 ;
  assign n10061 = n4390 & n6130 ;
  assign n10062 = ~n4385 & ~n10061 ;
  assign n10063 = n4391 & n6130 ;
  assign n10064 = n2905 & ~n10063 ;
  assign n10065 = ~n10062 & n10064 ;
  assign n10066 = ~n10060 & ~n10065 ;
  assign n10067 = ~n10059 & n10066 ;
  assign n10068 = n2453 & ~n10067 ;
  assign n10072 = ~\P3_PhyAddrPointer_reg[30]/NET0131  & ~n9046 ;
  assign n10073 = ~n9047 & ~n10072 ;
  assign n10074 = ~n2959 & ~n4415 ;
  assign n10075 = \P3_DataWidth_reg[1]/NET0131  & ~n4415 ;
  assign n10076 = ~n10074 & ~n10075 ;
  assign n10077 = n10073 & n10076 ;
  assign n10069 = ~\P3_PhyAddrPointer_reg[30]/NET0131  & ~n9050 ;
  assign n10070 = n2970 & ~n9051 ;
  assign n10071 = ~n10069 & n10070 ;
  assign n10078 = \P3_rEIP_reg[30]/NET0131  & n4412 ;
  assign n10079 = \P3_PhyAddrPointer_reg[30]/NET0131  & ~n9063 ;
  assign n10080 = ~n10078 & ~n10079 ;
  assign n10081 = ~n10071 & n10080 ;
  assign n10082 = ~n10077 & n10081 ;
  assign n10083 = ~n10068 & n10082 ;
  assign n10084 = \P1_PhyAddrPointer_reg[30]/NET0131  & n2375 ;
  assign n10085 = ~n4954 & ~n10084 ;
  assign n10086 = n2244 & ~n10085 ;
  assign n10087 = ~n2245 & ~n2369 ;
  assign n10088 = \P1_PhyAddrPointer_reg[30]/NET0131  & ~n10087 ;
  assign n10089 = ~n5071 & ~n10088 ;
  assign n10090 = ~n10086 & n10089 ;
  assign n10091 = n2432 & ~n10090 ;
  assign n10116 = \P1_PhyAddrPointer_reg[27]/NET0131  & \P1_PhyAddrPointer_reg[28]/NET0131  ;
  assign n10117 = \P1_PhyAddrPointer_reg[29]/NET0131  & n10116 ;
  assign n10111 = \P1_PhyAddrPointer_reg[22]/NET0131  & \P1_PhyAddrPointer_reg[23]/NET0131  ;
  assign n10112 = \P1_PhyAddrPointer_reg[24]/NET0131  & \P1_PhyAddrPointer_reg[25]/NET0131  ;
  assign n10113 = n10111 & n10112 ;
  assign n10107 = \P1_PhyAddrPointer_reg[18]/NET0131  & \P1_PhyAddrPointer_reg[19]/NET0131  ;
  assign n10108 = \P1_PhyAddrPointer_reg[20]/NET0131  & \P1_PhyAddrPointer_reg[21]/NET0131  ;
  assign n10109 = n10107 & n10108 ;
  assign n10092 = \P1_PhyAddrPointer_reg[2]/NET0131  & \P1_PhyAddrPointer_reg[3]/NET0131  ;
  assign n10093 = \P1_PhyAddrPointer_reg[4]/NET0131  & n10092 ;
  assign n10094 = \P1_PhyAddrPointer_reg[5]/NET0131  & n10093 ;
  assign n10095 = \P1_PhyAddrPointer_reg[6]/NET0131  & n10094 ;
  assign n10096 = \P1_PhyAddrPointer_reg[7]/NET0131  & n10095 ;
  assign n10097 = \P1_PhyAddrPointer_reg[8]/NET0131  & n10096 ;
  assign n10098 = \P1_PhyAddrPointer_reg[9]/NET0131  & n10097 ;
  assign n10099 = \P1_PhyAddrPointer_reg[10]/NET0131  & n10098 ;
  assign n10100 = \P1_PhyAddrPointer_reg[11]/NET0131  & n10099 ;
  assign n10101 = \P1_PhyAddrPointer_reg[12]/NET0131  & n10100 ;
  assign n10102 = \P1_PhyAddrPointer_reg[13]/NET0131  & n10101 ;
  assign n10103 = \P1_PhyAddrPointer_reg[14]/NET0131  & n10102 ;
  assign n10104 = \P1_PhyAddrPointer_reg[15]/NET0131  & n10103 ;
  assign n10105 = \P1_PhyAddrPointer_reg[16]/NET0131  & n10104 ;
  assign n10123 = \P1_PhyAddrPointer_reg[1]/NET0131  & n10105 ;
  assign n10124 = \P1_PhyAddrPointer_reg[17]/NET0131  & n10123 ;
  assign n10125 = n10109 & n10124 ;
  assign n10126 = n10113 & n10125 ;
  assign n10127 = \P1_PhyAddrPointer_reg[26]/NET0131  & n10126 ;
  assign n10128 = n10117 & n10127 ;
  assign n10129 = ~\P1_PhyAddrPointer_reg[30]/NET0131  & ~n10128 ;
  assign n10130 = \P1_PhyAddrPointer_reg[30]/NET0131  & n10128 ;
  assign n10131 = ~n10129 & ~n10130 ;
  assign n10132 = \P1_DataWidth_reg[1]/NET0131  & ~n5095 ;
  assign n10133 = ~n7697 & ~n10132 ;
  assign n10134 = n10131 & n10133 ;
  assign n10106 = \P1_PhyAddrPointer_reg[17]/NET0131  & n10105 ;
  assign n10110 = n10106 & n10109 ;
  assign n10114 = n10110 & n10113 ;
  assign n10115 = \P1_PhyAddrPointer_reg[26]/NET0131  & n10114 ;
  assign n10118 = n10115 & n10117 ;
  assign n10120 = ~\P1_PhyAddrPointer_reg[30]/NET0131  & ~n10118 ;
  assign n10119 = \P1_PhyAddrPointer_reg[30]/NET0131  & n10118 ;
  assign n10121 = n3148 & ~n10119 ;
  assign n10122 = ~n10120 & n10121 ;
  assign n10135 = ~n2439 & ~n2445 ;
  assign n10136 = ~n3027 & n10135 ;
  assign n10137 = \P1_PhyAddrPointer_reg[30]/NET0131  & ~n10136 ;
  assign n10138 = ~n5093 & ~n10137 ;
  assign n10139 = ~n10122 & n10138 ;
  assign n10140 = ~n10134 & n10139 ;
  assign n10141 = ~n10091 & n10140 ;
  assign n10144 = \P3_InstAddrPointer_reg[7]/NET0131  & n2896 ;
  assign n10146 = ~n4046 & n4053 ;
  assign n10148 = n4048 & ~n10146 ;
  assign n10147 = ~n4048 & n10146 ;
  assign n10149 = n3753 & ~n10147 ;
  assign n10150 = ~n10148 & n10149 ;
  assign n10145 = n4218 & ~n9123 ;
  assign n10151 = ~n9125 & ~n10145 ;
  assign n10152 = ~n10150 & n10151 ;
  assign n10153 = ~n2896 & ~n10152 ;
  assign n10154 = ~n10144 & ~n10153 ;
  assign n10155 = n2894 & ~n10154 ;
  assign n10159 = ~n4310 & ~n4346 ;
  assign n10161 = n4345 & n10159 ;
  assign n10160 = ~n4345 & ~n10159 ;
  assign n10162 = n2905 & ~n10160 ;
  assign n10163 = ~n10161 & n10162 ;
  assign n10143 = n2918 & n4309 ;
  assign n10156 = ~n2777 & n4178 ;
  assign n10164 = ~n10143 & ~n10156 ;
  assign n10157 = \P3_InstAddrPointer_reg[7]/NET0131  & ~n4402 ;
  assign n10158 = ~n2923 & n4048 ;
  assign n10165 = ~n10157 & ~n10158 ;
  assign n10166 = n10164 & n10165 ;
  assign n10167 = ~n10163 & n10166 ;
  assign n10168 = ~n10155 & n10167 ;
  assign n10169 = n2453 & ~n10168 ;
  assign n10142 = \P3_InstAddrPointer_reg[7]/NET0131  & ~n4418 ;
  assign n10170 = \P3_rEIP_reg[7]/NET0131  & n4412 ;
  assign n10171 = ~n10142 & ~n10170 ;
  assign n10172 = ~n10169 & n10171 ;
  assign n10186 = \P3_InstAddrPointer_reg[9]/NET0131  & n2896 ;
  assign n10193 = n6043 & n6058 ;
  assign n10191 = ~n4212 & n4227 ;
  assign n10192 = n4217 & ~n10191 ;
  assign n10194 = ~n3753 & ~n10192 ;
  assign n10195 = ~n10193 & n10194 ;
  assign n10187 = ~n8352 & ~n8354 ;
  assign n10188 = \P3_InstAddrPointer_reg[9]/NET0131  & n9129 ;
  assign n10189 = ~n10187 & ~n10188 ;
  assign n10190 = n3753 & ~n10189 ;
  assign n10196 = ~n2896 & ~n10190 ;
  assign n10197 = ~n10195 & n10196 ;
  assign n10198 = ~n10186 & ~n10197 ;
  assign n10199 = n2894 & ~n10198 ;
  assign n10201 = n4304 & ~n4348 ;
  assign n10203 = \P3_InstAddrPointer_reg[9]/NET0131  & n10201 ;
  assign n10181 = ~\P3_InstAddrPointer_reg[9]/NET0131  & ~n4302 ;
  assign n10182 = ~n4298 & ~n10181 ;
  assign n10202 = ~n10182 & ~n10201 ;
  assign n10204 = n2905 & ~n10202 ;
  assign n10205 = ~n10203 & n10204 ;
  assign n10176 = ~n2835 & ~n8354 ;
  assign n10177 = ~n2819 & ~n10176 ;
  assign n10178 = n7402 & ~n10177 ;
  assign n10179 = \P3_InstAddrPointer_reg[9]/NET0131  & ~n10178 ;
  assign n10200 = ~n2777 & n4217 ;
  assign n10206 = ~\P3_InstAddrPointer_reg[9]/NET0131  & n2835 ;
  assign n10207 = ~n10176 & ~n10206 ;
  assign n10208 = ~n2834 & n10207 ;
  assign n10175 = n2767 & n8354 ;
  assign n10180 = ~\P3_InstAddrPointer_reg[9]/NET0131  & ~n2847 ;
  assign n10183 = n2847 & ~n10182 ;
  assign n10184 = ~n10180 & ~n10183 ;
  assign n10185 = ~n2841 & n10184 ;
  assign n10209 = ~n10175 & ~n10185 ;
  assign n10210 = ~n10208 & n10209 ;
  assign n10211 = ~n10200 & n10210 ;
  assign n10212 = ~n10179 & n10211 ;
  assign n10213 = ~n10205 & n10212 ;
  assign n10214 = ~n10199 & n10213 ;
  assign n10215 = n2453 & ~n10214 ;
  assign n10173 = \P3_rEIP_reg[9]/NET0131  & n4412 ;
  assign n10174 = \P3_InstAddrPointer_reg[9]/NET0131  & ~n4418 ;
  assign n10216 = ~n10173 & ~n10174 ;
  assign n10217 = ~n10215 & n10216 ;
  assign n10222 = \P2_InstAddrPointer_reg[7]/NET0131  & n1897 ;
  assign n10223 = ~n6197 & n7469 ;
  assign n10224 = n6197 & ~n7469 ;
  assign n10225 = ~n10223 & ~n10224 ;
  assign n10226 = ~n6188 & ~n10225 ;
  assign n10227 = ~n6600 & n9167 ;
  assign n10228 = n6188 & ~n9168 ;
  assign n10229 = ~n10227 & n10228 ;
  assign n10230 = ~n10226 & ~n10229 ;
  assign n10231 = ~n1897 & ~n10230 ;
  assign n10232 = ~n10222 & ~n10231 ;
  assign n10233 = n1734 & ~n10232 ;
  assign n10244 = ~n6697 & ~n6733 ;
  assign n10246 = ~n6731 & n10244 ;
  assign n10245 = n6731 & ~n10244 ;
  assign n10247 = n1890 & ~n10245 ;
  assign n10248 = ~n10246 & n10247 ;
  assign n10236 = n1742 & ~n1810 ;
  assign n10237 = ~n1803 & ~n10236 ;
  assign n10250 = ~n6468 & ~n10237 ;
  assign n10251 = n1831 & ~n10250 ;
  assign n10252 = n6600 & ~n10251 ;
  assign n10219 = n1798 & ~n6696 ;
  assign n10220 = ~n1727 & ~n10219 ;
  assign n10234 = ~n1742 & n1814 ;
  assign n10235 = n1810 & ~n10234 ;
  assign n10238 = ~n1811 & ~n10237 ;
  assign n10239 = ~n1902 & ~n10238 ;
  assign n10240 = ~n1893 & n10239 ;
  assign n10241 = ~n10235 & n10240 ;
  assign n10242 = ~n10220 & n10241 ;
  assign n10243 = \P2_InstAddrPointer_reg[7]/NET0131  & ~n10242 ;
  assign n10221 = n1798 & n10220 ;
  assign n10249 = ~n1771 & n6197 ;
  assign n10253 = ~n10221 & ~n10249 ;
  assign n10254 = ~n10243 & n10253 ;
  assign n10255 = ~n10252 & n10254 ;
  assign n10256 = ~n10248 & n10255 ;
  assign n10257 = ~n10233 & n10256 ;
  assign n10258 = n1927 & ~n10257 ;
  assign n10218 = \P2_rEIP_reg[7]/NET0131  & n3113 ;
  assign n10259 = \P2_InstAddrPointer_reg[7]/NET0131  & ~n6810 ;
  assign n10260 = ~n10218 & ~n10259 ;
  assign n10261 = ~n10258 & n10260 ;
  assign n10265 = \P2_InstAddrPointer_reg[9]/NET0131  & n1897 ;
  assign n10270 = ~n6643 & n6645 ;
  assign n10269 = n6643 & ~n6645 ;
  assign n10271 = n6188 & ~n10269 ;
  assign n10272 = ~n10270 & n10271 ;
  assign n10266 = ~n6462 & n6480 ;
  assign n10267 = ~n6188 & ~n10266 ;
  assign n10268 = ~n9163 & n10267 ;
  assign n10273 = ~n1897 & ~n10268 ;
  assign n10274 = ~n10272 & n10273 ;
  assign n10275 = ~n10265 & ~n10274 ;
  assign n10276 = n1734 & ~n10275 ;
  assign n10277 = ~\P2_InstAddrPointer_reg[9]/NET0131  & ~n6735 ;
  assign n10278 = ~n6740 & ~n10277 ;
  assign n10279 = ~n6732 & n6737 ;
  assign n10280 = ~n10278 & ~n10279 ;
  assign n10281 = n1890 & ~n6739 ;
  assign n10282 = ~n10280 & n10281 ;
  assign n10284 = ~n1771 & n6480 ;
  assign n10285 = \P2_InstAddrPointer_reg[9]/NET0131  & n1805 ;
  assign n10286 = ~n1805 & n6645 ;
  assign n10287 = ~n10285 & ~n10286 ;
  assign n10288 = ~n1804 & ~n10287 ;
  assign n10289 = \P2_InstAddrPointer_reg[9]/NET0131  & ~n1820 ;
  assign n10290 = ~n1819 & n10286 ;
  assign n10291 = ~n10289 & ~n10290 ;
  assign n10292 = ~n1814 & ~n10291 ;
  assign n10293 = ~n10288 & ~n10292 ;
  assign n10294 = ~n1810 & ~n10293 ;
  assign n10264 = \P2_InstAddrPointer_reg[9]/NET0131  & ~n7636 ;
  assign n10283 = n1739 & n6645 ;
  assign n10295 = ~\P2_InstAddrPointer_reg[9]/NET0131  & ~n1798 ;
  assign n10296 = n1798 & ~n10278 ;
  assign n10297 = ~n10295 & ~n10296 ;
  assign n10298 = ~n1727 & n10297 ;
  assign n10299 = ~n10283 & ~n10298 ;
  assign n10300 = ~n10264 & n10299 ;
  assign n10301 = ~n10294 & n10300 ;
  assign n10302 = ~n10284 & n10301 ;
  assign n10303 = ~n10282 & n10302 ;
  assign n10304 = ~n10276 & n10303 ;
  assign n10305 = n1927 & ~n10304 ;
  assign n10262 = \P2_rEIP_reg[9]/NET0131  & n3113 ;
  assign n10263 = \P2_InstAddrPointer_reg[9]/NET0131  & ~n6810 ;
  assign n10306 = ~n10262 & ~n10263 ;
  assign n10307 = ~n10305 & n10306 ;
  assign n10308 = ~n5108 & ~n5188 ;
  assign n10309 = \P1_InstQueue_reg[11][2]/NET0131  & ~n5104 ;
  assign n10310 = ~n5107 & n10309 ;
  assign n10311 = ~n10308 & ~n10310 ;
  assign n10312 = ~n7697 & ~n10311 ;
  assign n10313 = ~n7703 & ~n10312 ;
  assign n10318 = ~n5256 & n5259 ;
  assign n10319 = ~n5260 & ~n10318 ;
  assign n10320 = n5148 & n10319 ;
  assign n10314 = n5233 & ~n5274 ;
  assign n10315 = ~n5275 & ~n10314 ;
  assign n10316 = ~n5148 & n10315 ;
  assign n10317 = n5095 & ~n10311 ;
  assign n10321 = n5153 & ~n10317 ;
  assign n10322 = ~n10316 & n10321 ;
  assign n10323 = ~n10320 & n10322 ;
  assign n10324 = ~n10313 & ~n10323 ;
  assign n10325 = \P1_InstQueue_reg[11][2]/NET0131  & ~n5291 ;
  assign n10326 = ~n1998 & n5104 ;
  assign n10327 = ~n10309 & ~n10326 ;
  assign n10328 = n3042 & ~n10327 ;
  assign n10329 = ~n10325 & ~n10328 ;
  assign n10330 = ~n10324 & n10329 ;
  assign n10339 = \buf2_reg[29]/NET0131  & ~n3079 ;
  assign n10340 = \buf1_reg[29]/NET0131  & n3079 ;
  assign n10341 = ~n10339 & ~n10340 ;
  assign n10342 = n3091 & ~n10341 ;
  assign n10343 = \buf2_reg[21]/NET0131  & ~n3079 ;
  assign n10344 = \buf1_reg[21]/NET0131  & n3079 ;
  assign n10345 = ~n10343 & ~n10344 ;
  assign n10346 = n3098 & ~n10345 ;
  assign n10347 = ~n10342 & ~n10346 ;
  assign n10348 = \P2_DataWidth_reg[1]/NET0131  & ~n10347 ;
  assign n10331 = \buf2_reg[5]/NET0131  & ~n3079 ;
  assign n10332 = \buf1_reg[5]/NET0131  & n3079 ;
  assign n10333 = ~n10331 & ~n10332 ;
  assign n10334 = ~n3050 & ~n10333 ;
  assign n10335 = \P2_InstQueue_reg[11][5]/NET0131  & ~n3049 ;
  assign n10336 = ~n3046 & n10335 ;
  assign n10337 = ~n10334 & ~n10336 ;
  assign n10349 = ~n3106 & ~n10337 ;
  assign n10350 = ~n10348 & ~n10349 ;
  assign n10351 = n1931 & ~n10350 ;
  assign n10338 = n3087 & ~n10337 ;
  assign n10352 = ~n1720 & n3049 ;
  assign n10353 = ~n10335 & ~n10352 ;
  assign n10354 = n3040 & ~n10353 ;
  assign n10355 = \P2_InstQueue_reg[11][5]/NET0131  & ~n3118 ;
  assign n10356 = ~n10354 & ~n10355 ;
  assign n10357 = ~n10338 & n10356 ;
  assign n10358 = ~n10351 & n10357 ;
  assign n10359 = ~n5188 & ~n5327 ;
  assign n10360 = \P1_InstQueue_reg[0][2]/NET0131  & ~n5324 ;
  assign n10361 = ~n5326 & n10360 ;
  assign n10362 = ~n10359 & ~n10361 ;
  assign n10363 = ~n7697 & ~n10362 ;
  assign n10364 = ~n7755 & ~n10363 ;
  assign n10367 = n5334 & n10319 ;
  assign n10365 = ~n5334 & n10315 ;
  assign n10366 = n5095 & ~n10362 ;
  assign n10368 = n5338 & ~n10366 ;
  assign n10369 = ~n10365 & n10368 ;
  assign n10370 = ~n10367 & n10369 ;
  assign n10371 = ~n10364 & ~n10370 ;
  assign n10372 = \P1_InstQueue_reg[0][2]/NET0131  & ~n5291 ;
  assign n10373 = ~n1998 & n5324 ;
  assign n10374 = ~n10360 & ~n10373 ;
  assign n10375 = n3042 & ~n10374 ;
  assign n10376 = ~n10372 & ~n10375 ;
  assign n10377 = ~n10371 & n10376 ;
  assign n10378 = ~n5188 & ~n5353 ;
  assign n10379 = \P1_InstQueue_reg[10][2]/NET0131  & ~n5107 ;
  assign n10380 = ~n5151 & n10379 ;
  assign n10381 = ~n10378 & ~n10380 ;
  assign n10382 = ~n7697 & ~n10381 ;
  assign n10383 = ~n7775 & ~n10382 ;
  assign n10386 = n5359 & n10319 ;
  assign n10384 = ~n5359 & n10315 ;
  assign n10385 = n5095 & ~n10381 ;
  assign n10387 = n5361 & ~n10385 ;
  assign n10388 = ~n10384 & n10387 ;
  assign n10389 = ~n10386 & n10388 ;
  assign n10390 = ~n10383 & ~n10389 ;
  assign n10391 = \P1_InstQueue_reg[10][2]/NET0131  & ~n5291 ;
  assign n10392 = ~n1998 & n5107 ;
  assign n10393 = ~n10379 & ~n10392 ;
  assign n10394 = n3042 & ~n10393 ;
  assign n10395 = ~n10391 & ~n10394 ;
  assign n10396 = ~n10390 & n10395 ;
  assign n10397 = ~n5188 & ~n5378 ;
  assign n10398 = \P1_InstQueue_reg[12][2]/NET0131  & ~n5377 ;
  assign n10399 = ~n5104 & n10398 ;
  assign n10400 = ~n10397 & ~n10399 ;
  assign n10401 = ~n7697 & ~n10400 ;
  assign n10402 = ~n7795 & ~n10401 ;
  assign n10405 = n5151 & n10319 ;
  assign n10403 = ~n5151 & n10315 ;
  assign n10404 = n5095 & ~n10400 ;
  assign n10406 = n5384 & ~n10404 ;
  assign n10407 = ~n10403 & n10406 ;
  assign n10408 = ~n10405 & n10407 ;
  assign n10409 = ~n10402 & ~n10408 ;
  assign n10410 = \P1_InstQueue_reg[12][2]/NET0131  & ~n5291 ;
  assign n10411 = ~n1998 & n5377 ;
  assign n10412 = ~n10398 & ~n10411 ;
  assign n10413 = n3042 & ~n10412 ;
  assign n10414 = ~n10410 & ~n10413 ;
  assign n10415 = ~n10409 & n10414 ;
  assign n10416 = ~n5188 & ~n5399 ;
  assign n10417 = \P1_InstQueue_reg[13][2]/NET0131  & ~n5334 ;
  assign n10418 = ~n5377 & n10417 ;
  assign n10419 = ~n10416 & ~n10418 ;
  assign n10420 = ~n7697 & ~n10419 ;
  assign n10421 = ~n7815 & ~n10420 ;
  assign n10424 = n5107 & n10319 ;
  assign n10422 = ~n5107 & n10315 ;
  assign n10423 = n5095 & ~n10419 ;
  assign n10425 = n5405 & ~n10423 ;
  assign n10426 = ~n10422 & n10425 ;
  assign n10427 = ~n10424 & n10426 ;
  assign n10428 = ~n10421 & ~n10427 ;
  assign n10429 = \P1_InstQueue_reg[13][2]/NET0131  & ~n5291 ;
  assign n10430 = ~n1998 & n5334 ;
  assign n10431 = ~n10417 & ~n10430 ;
  assign n10432 = n3042 & ~n10431 ;
  assign n10433 = ~n10429 & ~n10432 ;
  assign n10434 = ~n10428 & n10433 ;
  assign n10435 = ~n5188 & ~n5337 ;
  assign n10436 = \P1_InstQueue_reg[14][2]/NET0131  & ~n5336 ;
  assign n10437 = ~n5334 & n10436 ;
  assign n10438 = ~n10435 & ~n10437 ;
  assign n10439 = ~n7697 & ~n10438 ;
  assign n10440 = ~n7835 & ~n10439 ;
  assign n10443 = n5104 & n10319 ;
  assign n10441 = ~n5104 & n10315 ;
  assign n10442 = n5095 & ~n10438 ;
  assign n10444 = n5425 & ~n10442 ;
  assign n10445 = ~n10441 & n10444 ;
  assign n10446 = ~n10443 & n10445 ;
  assign n10447 = ~n10440 & ~n10446 ;
  assign n10448 = \P1_InstQueue_reg[14][2]/NET0131  & ~n5291 ;
  assign n10449 = ~n1998 & n5336 ;
  assign n10450 = ~n10436 & ~n10449 ;
  assign n10451 = n3042 & ~n10450 ;
  assign n10452 = ~n10448 & ~n10451 ;
  assign n10453 = ~n10447 & n10452 ;
  assign n10454 = ~n5188 & ~n5440 ;
  assign n10455 = \P1_InstQueue_reg[15][2]/NET0131  & ~n5326 ;
  assign n10456 = ~n5336 & n10455 ;
  assign n10457 = ~n10454 & ~n10456 ;
  assign n10458 = ~n7697 & ~n10457 ;
  assign n10459 = ~n7855 & ~n10458 ;
  assign n10462 = n5377 & n10319 ;
  assign n10460 = ~n5377 & n10315 ;
  assign n10461 = n5095 & ~n10457 ;
  assign n10463 = n5446 & ~n10461 ;
  assign n10464 = ~n10460 & n10463 ;
  assign n10465 = ~n10462 & n10464 ;
  assign n10466 = ~n10459 & ~n10465 ;
  assign n10467 = \P1_InstQueue_reg[15][2]/NET0131  & ~n5291 ;
  assign n10468 = ~n1998 & n5326 ;
  assign n10469 = ~n10455 & ~n10468 ;
  assign n10470 = n3042 & ~n10469 ;
  assign n10471 = ~n10467 & ~n10470 ;
  assign n10472 = ~n10466 & n10471 ;
  assign n10473 = ~n5188 & ~n5462 ;
  assign n10474 = \P1_InstQueue_reg[1][2]/NET0131  & ~n5461 ;
  assign n10475 = ~n5324 & n10474 ;
  assign n10476 = ~n10473 & ~n10475 ;
  assign n10477 = ~n7697 & ~n10476 ;
  assign n10478 = ~n7875 & ~n10477 ;
  assign n10481 = n5336 & n10319 ;
  assign n10479 = ~n5336 & n10315 ;
  assign n10480 = n5095 & ~n10476 ;
  assign n10482 = n5468 & ~n10480 ;
  assign n10483 = ~n10479 & n10482 ;
  assign n10484 = ~n10481 & n10483 ;
  assign n10485 = ~n10478 & ~n10484 ;
  assign n10486 = \P1_InstQueue_reg[1][2]/NET0131  & ~n5291 ;
  assign n10487 = ~n1998 & n5461 ;
  assign n10488 = ~n10474 & ~n10487 ;
  assign n10489 = n3042 & ~n10488 ;
  assign n10490 = ~n10486 & ~n10489 ;
  assign n10491 = ~n10485 & n10490 ;
  assign n10492 = ~n5188 & ~n5506 ;
  assign n10493 = \P1_InstQueue_reg[2][2]/NET0131  & ~n5484 ;
  assign n10494 = ~n5461 & n10493 ;
  assign n10495 = ~n10492 & ~n10494 ;
  assign n10496 = ~n7697 & ~n10495 ;
  assign n10497 = ~n7895 & ~n10496 ;
  assign n10500 = n5326 & n10319 ;
  assign n10498 = ~n5326 & n10315 ;
  assign n10499 = n5095 & ~n10495 ;
  assign n10501 = n5512 & ~n10499 ;
  assign n10502 = ~n10498 & n10501 ;
  assign n10503 = ~n10500 & n10502 ;
  assign n10504 = ~n10497 & ~n10503 ;
  assign n10505 = \P1_InstQueue_reg[2][2]/NET0131  & ~n5291 ;
  assign n10506 = ~n1998 & n5484 ;
  assign n10507 = ~n10493 & ~n10506 ;
  assign n10508 = n3042 & ~n10507 ;
  assign n10509 = ~n10505 & ~n10508 ;
  assign n10510 = ~n10504 & n10509 ;
  assign n10511 = ~n5188 & ~n5485 ;
  assign n10512 = \P1_InstQueue_reg[3][2]/NET0131  & ~n5483 ;
  assign n10513 = ~n5484 & n10512 ;
  assign n10514 = ~n10511 & ~n10513 ;
  assign n10515 = ~n7697 & ~n10514 ;
  assign n10516 = ~n7915 & ~n10515 ;
  assign n10519 = n5324 & n10319 ;
  assign n10517 = ~n5324 & n10315 ;
  assign n10518 = n5095 & ~n10514 ;
  assign n10520 = n5491 & ~n10518 ;
  assign n10521 = ~n10517 & n10520 ;
  assign n10522 = ~n10519 & n10521 ;
  assign n10523 = ~n10516 & ~n10522 ;
  assign n10524 = \P1_InstQueue_reg[3][2]/NET0131  & ~n5291 ;
  assign n10525 = ~n1998 & n5483 ;
  assign n10526 = ~n10512 & ~n10525 ;
  assign n10527 = n3042 & ~n10526 ;
  assign n10528 = ~n10524 & ~n10527 ;
  assign n10529 = ~n10523 & n10528 ;
  assign n10530 = ~n5188 & ~n5528 ;
  assign n10531 = \P1_InstQueue_reg[4][2]/NET0131  & ~n5527 ;
  assign n10532 = ~n5483 & n10531 ;
  assign n10533 = ~n10530 & ~n10532 ;
  assign n10534 = ~n7697 & ~n10533 ;
  assign n10535 = ~n7935 & ~n10534 ;
  assign n10538 = n5461 & n10319 ;
  assign n10536 = ~n5461 & n10315 ;
  assign n10537 = n5095 & ~n10533 ;
  assign n10539 = n5534 & ~n10537 ;
  assign n10540 = ~n10536 & n10539 ;
  assign n10541 = ~n10538 & n10540 ;
  assign n10542 = ~n10535 & ~n10541 ;
  assign n10543 = \P1_InstQueue_reg[4][2]/NET0131  & ~n5291 ;
  assign n10544 = ~n1998 & n5527 ;
  assign n10545 = ~n10531 & ~n10544 ;
  assign n10546 = n3042 & ~n10545 ;
  assign n10547 = ~n10543 & ~n10546 ;
  assign n10548 = ~n10542 & n10547 ;
  assign n10549 = ~n5188 & ~n5550 ;
  assign n10550 = \P1_InstQueue_reg[5][2]/NET0131  & ~n5549 ;
  assign n10551 = ~n5527 & n10550 ;
  assign n10552 = ~n10549 & ~n10551 ;
  assign n10553 = ~n7697 & ~n10552 ;
  assign n10554 = ~n7955 & ~n10553 ;
  assign n10557 = n5484 & n10319 ;
  assign n10555 = ~n5484 & n10315 ;
  assign n10556 = n5095 & ~n10552 ;
  assign n10558 = n5556 & ~n10556 ;
  assign n10559 = ~n10555 & n10558 ;
  assign n10560 = ~n10557 & n10559 ;
  assign n10561 = ~n10554 & ~n10560 ;
  assign n10562 = \P1_InstQueue_reg[5][2]/NET0131  & ~n5291 ;
  assign n10563 = ~n1998 & n5549 ;
  assign n10564 = ~n10550 & ~n10563 ;
  assign n10565 = n3042 & ~n10564 ;
  assign n10566 = ~n10562 & ~n10565 ;
  assign n10567 = ~n10561 & n10566 ;
  assign n10568 = ~n5188 & ~n5572 ;
  assign n10569 = \P1_InstQueue_reg[6][2]/NET0131  & ~n5571 ;
  assign n10570 = ~n5549 & n10569 ;
  assign n10571 = ~n10568 & ~n10570 ;
  assign n10572 = ~n7697 & ~n10571 ;
  assign n10573 = ~n7975 & ~n10572 ;
  assign n10576 = n5483 & n10319 ;
  assign n10574 = ~n5483 & n10315 ;
  assign n10575 = n5095 & ~n10571 ;
  assign n10577 = n5578 & ~n10575 ;
  assign n10578 = ~n10574 & n10577 ;
  assign n10579 = ~n10576 & n10578 ;
  assign n10580 = ~n10573 & ~n10579 ;
  assign n10581 = \P1_InstQueue_reg[6][2]/NET0131  & ~n5291 ;
  assign n10582 = ~n1998 & n5571 ;
  assign n10583 = ~n10569 & ~n10582 ;
  assign n10584 = n3042 & ~n10583 ;
  assign n10585 = ~n10581 & ~n10584 ;
  assign n10586 = ~n10580 & n10585 ;
  assign n10587 = ~n5188 & ~n5593 ;
  assign n10588 = \P1_InstQueue_reg[7][2]/NET0131  & ~n5359 ;
  assign n10589 = ~n5571 & n10588 ;
  assign n10590 = ~n10587 & ~n10589 ;
  assign n10591 = ~n7697 & ~n10590 ;
  assign n10592 = ~n7995 & ~n10591 ;
  assign n10595 = n5527 & n10319 ;
  assign n10593 = ~n5527 & n10315 ;
  assign n10594 = n5095 & ~n10590 ;
  assign n10596 = n5599 & ~n10594 ;
  assign n10597 = ~n10593 & n10596 ;
  assign n10598 = ~n10595 & n10597 ;
  assign n10599 = ~n10592 & ~n10598 ;
  assign n10600 = \P1_InstQueue_reg[7][2]/NET0131  & ~n5291 ;
  assign n10601 = ~n1998 & n5359 ;
  assign n10602 = ~n10588 & ~n10601 ;
  assign n10603 = n3042 & ~n10602 ;
  assign n10604 = ~n10600 & ~n10603 ;
  assign n10605 = ~n10599 & n10604 ;
  assign n10606 = ~n5188 & ~n5360 ;
  assign n10607 = \P1_InstQueue_reg[8][2]/NET0131  & ~n5148 ;
  assign n10608 = ~n5359 & n10607 ;
  assign n10609 = ~n10606 & ~n10608 ;
  assign n10610 = ~n7697 & ~n10609 ;
  assign n10611 = ~n8015 & ~n10610 ;
  assign n10614 = n5549 & n10319 ;
  assign n10612 = ~n5549 & n10315 ;
  assign n10613 = n5095 & ~n10609 ;
  assign n10615 = n5619 & ~n10613 ;
  assign n10616 = ~n10612 & n10615 ;
  assign n10617 = ~n10614 & n10616 ;
  assign n10618 = ~n10611 & ~n10617 ;
  assign n10619 = \P1_InstQueue_reg[8][2]/NET0131  & ~n5291 ;
  assign n10620 = ~n1998 & n5148 ;
  assign n10621 = ~n10607 & ~n10620 ;
  assign n10622 = n3042 & ~n10621 ;
  assign n10623 = ~n10619 & ~n10622 ;
  assign n10624 = ~n10618 & n10623 ;
  assign n10625 = ~n5152 & ~n5188 ;
  assign n10626 = \P1_InstQueue_reg[9][2]/NET0131  & ~n5151 ;
  assign n10627 = ~n5148 & n10626 ;
  assign n10628 = ~n10625 & ~n10627 ;
  assign n10629 = ~n7697 & ~n10628 ;
  assign n10630 = ~n8035 & ~n10629 ;
  assign n10633 = n5571 & n10319 ;
  assign n10631 = ~n5571 & n10315 ;
  assign n10632 = n5095 & ~n10628 ;
  assign n10634 = n5639 & ~n10632 ;
  assign n10635 = ~n10631 & n10634 ;
  assign n10636 = ~n10633 & n10635 ;
  assign n10637 = ~n10630 & ~n10636 ;
  assign n10638 = \P1_InstQueue_reg[9][2]/NET0131  & ~n5291 ;
  assign n10639 = ~n1998 & n5151 ;
  assign n10640 = ~n10626 & ~n10639 ;
  assign n10641 = n3042 & ~n10640 ;
  assign n10642 = ~n10638 & ~n10641 ;
  assign n10643 = ~n10637 & n10642 ;
  assign n10649 = n3162 & ~n10341 ;
  assign n10650 = n3165 & ~n10345 ;
  assign n10651 = ~n10649 & ~n10650 ;
  assign n10652 = \P2_DataWidth_reg[1]/NET0131  & ~n10651 ;
  assign n10644 = ~n3155 & ~n10333 ;
  assign n10645 = \P2_InstQueue_reg[0][5]/NET0131  & ~n3152 ;
  assign n10646 = ~n3154 & n10645 ;
  assign n10647 = ~n10644 & ~n10646 ;
  assign n10653 = ~n3170 & ~n10647 ;
  assign n10654 = ~n10652 & ~n10653 ;
  assign n10655 = n1931 & ~n10654 ;
  assign n10648 = n3087 & ~n10647 ;
  assign n10656 = ~n1720 & n3152 ;
  assign n10657 = ~n10645 & ~n10656 ;
  assign n10658 = n3040 & ~n10657 ;
  assign n10659 = \P2_InstQueue_reg[0][5]/NET0131  & ~n3118 ;
  assign n10660 = ~n10658 & ~n10659 ;
  assign n10661 = ~n10648 & n10660 ;
  assign n10662 = ~n10655 & n10661 ;
  assign n10668 = n3091 & ~n10345 ;
  assign n10669 = n3198 & ~n10341 ;
  assign n10670 = ~n10668 & ~n10669 ;
  assign n10671 = \P2_DataWidth_reg[1]/NET0131  & ~n10670 ;
  assign n10663 = ~n3202 & ~n10333 ;
  assign n10664 = \P2_InstQueue_reg[10][5]/NET0131  & ~n3046 ;
  assign n10665 = ~n3098 & n10664 ;
  assign n10666 = ~n10663 & ~n10665 ;
  assign n10672 = ~n3200 & ~n10666 ;
  assign n10673 = ~n10671 & ~n10672 ;
  assign n10674 = n1931 & ~n10673 ;
  assign n10667 = n3087 & ~n10666 ;
  assign n10675 = ~n1720 & n3046 ;
  assign n10676 = ~n10664 & ~n10675 ;
  assign n10677 = n3040 & ~n10676 ;
  assign n10678 = \P2_InstQueue_reg[10][5]/NET0131  & ~n3118 ;
  assign n10679 = ~n10677 & ~n10678 ;
  assign n10680 = ~n10667 & n10679 ;
  assign n10681 = ~n10674 & n10680 ;
  assign n10687 = n3098 & ~n10341 ;
  assign n10688 = n3046 & ~n10345 ;
  assign n10689 = ~n10687 & ~n10688 ;
  assign n10690 = \P2_DataWidth_reg[1]/NET0131  & ~n10689 ;
  assign n10682 = ~n3238 & ~n10333 ;
  assign n10683 = \P2_InstQueue_reg[12][5]/NET0131  & ~n3237 ;
  assign n10684 = ~n3049 & n10683 ;
  assign n10685 = ~n10682 & ~n10684 ;
  assign n10691 = ~n3248 & ~n10685 ;
  assign n10692 = ~n10690 & ~n10691 ;
  assign n10693 = n1931 & ~n10692 ;
  assign n10686 = n3087 & ~n10685 ;
  assign n10694 = ~n1720 & n3237 ;
  assign n10695 = ~n10683 & ~n10694 ;
  assign n10696 = n3040 & ~n10695 ;
  assign n10697 = \P2_InstQueue_reg[12][5]/NET0131  & ~n3118 ;
  assign n10698 = ~n10696 & ~n10697 ;
  assign n10699 = ~n10686 & n10698 ;
  assign n10700 = ~n10693 & n10699 ;
  assign n10706 = n3046 & ~n10341 ;
  assign n10707 = n3049 & ~n10345 ;
  assign n10708 = ~n10706 & ~n10707 ;
  assign n10709 = \P2_DataWidth_reg[1]/NET0131  & ~n10708 ;
  assign n10701 = ~n3275 & ~n10333 ;
  assign n10702 = \P2_InstQueue_reg[13][5]/NET0131  & ~n3162 ;
  assign n10703 = ~n3237 & n10702 ;
  assign n10704 = ~n10701 & ~n10703 ;
  assign n10710 = ~n3285 & ~n10704 ;
  assign n10711 = ~n10709 & ~n10710 ;
  assign n10712 = n1931 & ~n10711 ;
  assign n10705 = n3087 & ~n10704 ;
  assign n10713 = ~n1720 & n3162 ;
  assign n10714 = ~n10702 & ~n10713 ;
  assign n10715 = n3040 & ~n10714 ;
  assign n10716 = \P2_InstQueue_reg[13][5]/NET0131  & ~n3118 ;
  assign n10717 = ~n10715 & ~n10716 ;
  assign n10718 = ~n10705 & n10717 ;
  assign n10719 = ~n10712 & n10718 ;
  assign n10725 = n3049 & ~n10341 ;
  assign n10726 = n3237 & ~n10345 ;
  assign n10727 = ~n10725 & ~n10726 ;
  assign n10728 = \P2_DataWidth_reg[1]/NET0131  & ~n10727 ;
  assign n10720 = ~n3169 & ~n10333 ;
  assign n10721 = \P2_InstQueue_reg[14][5]/NET0131  & ~n3165 ;
  assign n10722 = ~n3162 & n10721 ;
  assign n10723 = ~n10720 & ~n10722 ;
  assign n10729 = ~n3321 & ~n10723 ;
  assign n10730 = ~n10728 & ~n10729 ;
  assign n10731 = n1931 & ~n10730 ;
  assign n10724 = n3087 & ~n10723 ;
  assign n10732 = ~n1720 & n3165 ;
  assign n10733 = ~n10721 & ~n10732 ;
  assign n10734 = n3040 & ~n10733 ;
  assign n10735 = \P2_InstQueue_reg[14][5]/NET0131  & ~n3118 ;
  assign n10736 = ~n10734 & ~n10735 ;
  assign n10737 = ~n10724 & n10736 ;
  assign n10738 = ~n10731 & n10737 ;
  assign n10744 = n3237 & ~n10341 ;
  assign n10745 = n3162 & ~n10345 ;
  assign n10746 = ~n10744 & ~n10745 ;
  assign n10747 = \P2_DataWidth_reg[1]/NET0131  & ~n10746 ;
  assign n10739 = ~n3348 & ~n10333 ;
  assign n10740 = \P2_InstQueue_reg[15][5]/NET0131  & ~n3154 ;
  assign n10741 = ~n3165 & n10740 ;
  assign n10742 = ~n10739 & ~n10741 ;
  assign n10748 = ~n3358 & ~n10742 ;
  assign n10749 = ~n10747 & ~n10748 ;
  assign n10750 = n1931 & ~n10749 ;
  assign n10743 = n3087 & ~n10742 ;
  assign n10751 = ~n1720 & n3154 ;
  assign n10752 = ~n10740 & ~n10751 ;
  assign n10753 = n3040 & ~n10752 ;
  assign n10754 = \P2_InstQueue_reg[15][5]/NET0131  & ~n3118 ;
  assign n10755 = ~n10753 & ~n10754 ;
  assign n10756 = ~n10743 & n10755 ;
  assign n10757 = ~n10750 & n10756 ;
  assign n10763 = n3165 & ~n10341 ;
  assign n10764 = n3154 & ~n10345 ;
  assign n10765 = ~n10763 & ~n10764 ;
  assign n10766 = \P2_DataWidth_reg[1]/NET0131  & ~n10765 ;
  assign n10758 = ~n3389 & ~n10333 ;
  assign n10759 = \P2_InstQueue_reg[1][5]/NET0131  & ~n3388 ;
  assign n10760 = ~n3152 & n10759 ;
  assign n10761 = ~n10758 & ~n10760 ;
  assign n10767 = ~n3386 & ~n10761 ;
  assign n10768 = ~n10766 & ~n10767 ;
  assign n10769 = n1931 & ~n10768 ;
  assign n10762 = n3087 & ~n10761 ;
  assign n10770 = ~n1720 & n3388 ;
  assign n10771 = ~n10759 & ~n10770 ;
  assign n10772 = n3040 & ~n10771 ;
  assign n10773 = \P2_InstQueue_reg[1][5]/NET0131  & ~n3118 ;
  assign n10774 = ~n10772 & ~n10773 ;
  assign n10775 = ~n10762 & n10774 ;
  assign n10776 = ~n10769 & n10775 ;
  assign n10782 = n3152 & ~n10345 ;
  assign n10783 = n3154 & ~n10341 ;
  assign n10784 = ~n10782 & ~n10783 ;
  assign n10785 = \P2_DataWidth_reg[1]/NET0131  & ~n10784 ;
  assign n10777 = ~n3424 & ~n10333 ;
  assign n10778 = \P2_InstQueue_reg[2][5]/NET0131  & ~n3423 ;
  assign n10779 = ~n3388 & n10778 ;
  assign n10780 = ~n10777 & ~n10779 ;
  assign n10786 = ~n3434 & ~n10780 ;
  assign n10787 = ~n10785 & ~n10786 ;
  assign n10788 = n1931 & ~n10787 ;
  assign n10781 = n3087 & ~n10780 ;
  assign n10789 = ~n1720 & n3423 ;
  assign n10790 = ~n10778 & ~n10789 ;
  assign n10791 = n3040 & ~n10790 ;
  assign n10792 = \P2_InstQueue_reg[2][5]/NET0131  & ~n3118 ;
  assign n10793 = ~n10791 & ~n10792 ;
  assign n10794 = ~n10781 & n10793 ;
  assign n10795 = ~n10788 & n10794 ;
  assign n10801 = n3152 & ~n10341 ;
  assign n10802 = n3388 & ~n10345 ;
  assign n10803 = ~n10801 & ~n10802 ;
  assign n10804 = \P2_DataWidth_reg[1]/NET0131  & ~n10803 ;
  assign n10796 = ~n3462 & ~n10333 ;
  assign n10797 = \P2_InstQueue_reg[3][5]/NET0131  & ~n3461 ;
  assign n10798 = ~n3423 & n10797 ;
  assign n10799 = ~n10796 & ~n10798 ;
  assign n10805 = ~n3472 & ~n10799 ;
  assign n10806 = ~n10804 & ~n10805 ;
  assign n10807 = n1931 & ~n10806 ;
  assign n10800 = n3087 & ~n10799 ;
  assign n10808 = ~n1720 & n3461 ;
  assign n10809 = ~n10797 & ~n10808 ;
  assign n10810 = n3040 & ~n10809 ;
  assign n10811 = \P2_InstQueue_reg[3][5]/NET0131  & ~n3118 ;
  assign n10812 = ~n10810 & ~n10811 ;
  assign n10813 = ~n10800 & n10812 ;
  assign n10814 = ~n10807 & n10813 ;
  assign n10820 = n3388 & ~n10341 ;
  assign n10821 = n3423 & ~n10345 ;
  assign n10822 = ~n10820 & ~n10821 ;
  assign n10823 = \P2_DataWidth_reg[1]/NET0131  & ~n10822 ;
  assign n10815 = ~n3500 & ~n10333 ;
  assign n10816 = \P2_InstQueue_reg[4][5]/NET0131  & ~n3499 ;
  assign n10817 = ~n3461 & n10816 ;
  assign n10818 = ~n10815 & ~n10817 ;
  assign n10824 = ~n3510 & ~n10818 ;
  assign n10825 = ~n10823 & ~n10824 ;
  assign n10826 = n1931 & ~n10825 ;
  assign n10819 = n3087 & ~n10818 ;
  assign n10827 = ~n1720 & n3499 ;
  assign n10828 = ~n10816 & ~n10827 ;
  assign n10829 = n3040 & ~n10828 ;
  assign n10830 = \P2_InstQueue_reg[4][5]/NET0131  & ~n3118 ;
  assign n10831 = ~n10829 & ~n10830 ;
  assign n10832 = ~n10819 & n10831 ;
  assign n10833 = ~n10826 & n10832 ;
  assign n10839 = n3423 & ~n10341 ;
  assign n10840 = n3461 & ~n10345 ;
  assign n10841 = ~n10839 & ~n10840 ;
  assign n10842 = \P2_DataWidth_reg[1]/NET0131  & ~n10841 ;
  assign n10834 = ~n3538 & ~n10333 ;
  assign n10835 = \P2_InstQueue_reg[5][5]/NET0131  & ~n3537 ;
  assign n10836 = ~n3499 & n10835 ;
  assign n10837 = ~n10834 & ~n10836 ;
  assign n10843 = ~n3548 & ~n10837 ;
  assign n10844 = ~n10842 & ~n10843 ;
  assign n10845 = n1931 & ~n10844 ;
  assign n10838 = n3087 & ~n10837 ;
  assign n10846 = ~n1720 & n3537 ;
  assign n10847 = ~n10835 & ~n10846 ;
  assign n10848 = n3040 & ~n10847 ;
  assign n10849 = \P2_InstQueue_reg[5][5]/NET0131  & ~n3118 ;
  assign n10850 = ~n10848 & ~n10849 ;
  assign n10851 = ~n10838 & n10850 ;
  assign n10852 = ~n10845 & n10851 ;
  assign n10858 = n3461 & ~n10341 ;
  assign n10859 = n3499 & ~n10345 ;
  assign n10860 = ~n10858 & ~n10859 ;
  assign n10861 = \P2_DataWidth_reg[1]/NET0131  & ~n10860 ;
  assign n10853 = ~n3576 & ~n10333 ;
  assign n10854 = \P2_InstQueue_reg[6][5]/NET0131  & ~n3575 ;
  assign n10855 = ~n3537 & n10854 ;
  assign n10856 = ~n10853 & ~n10855 ;
  assign n10862 = ~n3586 & ~n10856 ;
  assign n10863 = ~n10861 & ~n10862 ;
  assign n10864 = n1931 & ~n10863 ;
  assign n10857 = n3087 & ~n10856 ;
  assign n10865 = ~n1720 & n3575 ;
  assign n10866 = ~n10854 & ~n10865 ;
  assign n10867 = n3040 & ~n10866 ;
  assign n10868 = \P2_InstQueue_reg[6][5]/NET0131  & ~n3118 ;
  assign n10869 = ~n10867 & ~n10868 ;
  assign n10870 = ~n10857 & n10869 ;
  assign n10871 = ~n10864 & n10870 ;
  assign n10877 = n3499 & ~n10341 ;
  assign n10878 = n3537 & ~n10345 ;
  assign n10879 = ~n10877 & ~n10878 ;
  assign n10880 = \P2_DataWidth_reg[1]/NET0131  & ~n10879 ;
  assign n10872 = ~n3613 & ~n10333 ;
  assign n10873 = \P2_InstQueue_reg[7][5]/NET0131  & ~n3198 ;
  assign n10874 = ~n3575 & n10873 ;
  assign n10875 = ~n10872 & ~n10874 ;
  assign n10881 = ~n3623 & ~n10875 ;
  assign n10882 = ~n10880 & ~n10881 ;
  assign n10883 = n1931 & ~n10882 ;
  assign n10876 = n3087 & ~n10875 ;
  assign n10884 = ~n1720 & n3198 ;
  assign n10885 = ~n10873 & ~n10884 ;
  assign n10886 = n3040 & ~n10885 ;
  assign n10887 = \P2_InstQueue_reg[7][5]/NET0131  & ~n3118 ;
  assign n10888 = ~n10886 & ~n10887 ;
  assign n10889 = ~n10876 & n10888 ;
  assign n10890 = ~n10883 & n10889 ;
  assign n10896 = n3537 & ~n10341 ;
  assign n10897 = n3575 & ~n10345 ;
  assign n10898 = ~n10896 & ~n10897 ;
  assign n10899 = \P2_DataWidth_reg[1]/NET0131  & ~n10898 ;
  assign n10891 = ~n3199 & ~n10333 ;
  assign n10892 = \P2_InstQueue_reg[8][5]/NET0131  & ~n3091 ;
  assign n10893 = ~n3198 & n10892 ;
  assign n10894 = ~n10891 & ~n10893 ;
  assign n10900 = ~n3659 & ~n10894 ;
  assign n10901 = ~n10899 & ~n10900 ;
  assign n10902 = n1931 & ~n10901 ;
  assign n10895 = n3087 & ~n10894 ;
  assign n10903 = ~n1720 & n3091 ;
  assign n10904 = ~n10892 & ~n10903 ;
  assign n10905 = n3040 & ~n10904 ;
  assign n10906 = \P2_InstQueue_reg[8][5]/NET0131  & ~n3118 ;
  assign n10907 = ~n10905 & ~n10906 ;
  assign n10908 = ~n10895 & n10907 ;
  assign n10909 = ~n10902 & n10908 ;
  assign n10915 = n3575 & ~n10341 ;
  assign n10916 = n3198 & ~n10345 ;
  assign n10917 = ~n10915 & ~n10916 ;
  assign n10918 = \P2_DataWidth_reg[1]/NET0131  & ~n10917 ;
  assign n10910 = ~n3105 & ~n10333 ;
  assign n10911 = \P2_InstQueue_reg[9][5]/NET0131  & ~n3098 ;
  assign n10912 = ~n3091 & n10911 ;
  assign n10913 = ~n10910 & ~n10912 ;
  assign n10919 = ~n3695 & ~n10913 ;
  assign n10920 = ~n10918 & ~n10919 ;
  assign n10921 = n1931 & ~n10920 ;
  assign n10914 = n3087 & ~n10913 ;
  assign n10922 = ~n1720 & n3098 ;
  assign n10923 = ~n10911 & ~n10922 ;
  assign n10924 = n3040 & ~n10923 ;
  assign n10925 = \P2_InstQueue_reg[9][5]/NET0131  & ~n3118 ;
  assign n10926 = ~n10924 & ~n10925 ;
  assign n10927 = ~n10914 & n10926 ;
  assign n10928 = ~n10921 & n10927 ;
  assign n10929 = \P2_PhyAddrPointer_reg[23]/NET0131  & n1897 ;
  assign n10943 = n6554 & ~n8916 ;
  assign n10939 = ~n6539 & n8914 ;
  assign n10940 = ~n6537 & ~n6554 ;
  assign n10941 = n6551 & n10940 ;
  assign n10942 = n10939 & n10941 ;
  assign n10944 = ~n6188 & ~n10942 ;
  assign n10945 = ~n10943 & n10944 ;
  assign n10930 = \P2_InstAddrPointer_reg[23]/NET0131  & n6556 ;
  assign n10931 = ~\P2_InstAddrPointer_reg[23]/NET0131  & ~n6556 ;
  assign n10932 = ~n10930 & ~n10931 ;
  assign n10933 = n6548 & n7594 ;
  assign n10934 = n7592 & n10933 ;
  assign n10936 = n10932 & ~n10934 ;
  assign n10935 = ~n10932 & n10934 ;
  assign n10937 = n6188 & ~n10935 ;
  assign n10938 = ~n10936 & n10937 ;
  assign n10946 = ~n1897 & ~n10938 ;
  assign n10947 = ~n10945 & n10946 ;
  assign n10948 = ~n10929 & ~n10947 ;
  assign n10949 = n1734 & ~n10948 ;
  assign n10950 = \P2_PhyAddrPointer_reg[23]/NET0131  & ~n8936 ;
  assign n10952 = n7623 & n8942 ;
  assign n10951 = ~n7623 & ~n8942 ;
  assign n10953 = n1890 & ~n10951 ;
  assign n10954 = ~n10952 & n10953 ;
  assign n10955 = ~n10950 & ~n10954 ;
  assign n10956 = ~n10949 & n10955 ;
  assign n10957 = n1927 & ~n10956 ;
  assign n10965 = ~\P2_DataWidth_reg[1]/NET0131  & ~\P2_PhyAddrPointer_reg[1]/NET0131  ;
  assign n10966 = n8979 & ~n10965 ;
  assign n10968 = \P2_PhyAddrPointer_reg[23]/NET0131  & n10966 ;
  assign n10967 = ~\P2_PhyAddrPointer_reg[23]/NET0131  & ~n10966 ;
  assign n10969 = n1931 & ~n10967 ;
  assign n10970 = ~n10968 & n10969 ;
  assign n10959 = \P2_PhyAddrPointer_reg[1]/NET0131  & n8979 ;
  assign n10960 = ~\P2_PhyAddrPointer_reg[23]/NET0131  & ~n10959 ;
  assign n10961 = \P2_PhyAddrPointer_reg[1]/NET0131  & n8980 ;
  assign n10962 = ~n10960 & ~n10961 ;
  assign n10963 = n3087 & n10962 ;
  assign n10958 = \P2_rEIP_reg[23]/NET0131  & n3113 ;
  assign n10964 = \P2_PhyAddrPointer_reg[23]/NET0131  & ~n8958 ;
  assign n10971 = ~n10958 & ~n10964 ;
  assign n10972 = ~n10963 & n10971 ;
  assign n10973 = ~n10970 & n10972 ;
  assign n10974 = ~n10957 & n10973 ;
  assign n10975 = \P2_PhyAddrPointer_reg[27]/NET0131  & n1897 ;
  assign n10976 = ~n6560 & n6572 ;
  assign n10977 = n6576 & n10976 ;
  assign n10978 = n10942 & n10977 ;
  assign n10979 = ~n6576 & ~n7608 ;
  assign n10980 = ~n6188 & ~n10979 ;
  assign n10981 = ~n10978 & n10980 ;
  assign n10983 = n6676 & n7598 ;
  assign n10982 = ~n6676 & ~n7598 ;
  assign n10984 = n6188 & ~n10982 ;
  assign n10985 = ~n10983 & n10984 ;
  assign n10986 = ~n10981 & ~n10985 ;
  assign n10987 = ~n1897 & ~n10986 ;
  assign n10988 = ~n10975 & ~n10987 ;
  assign n10989 = n1734 & ~n10988 ;
  assign n10990 = \P2_PhyAddrPointer_reg[27]/NET0131  & ~n8936 ;
  assign n10992 = n6778 & n8943 ;
  assign n10991 = ~n6778 & ~n8943 ;
  assign n10993 = n1890 & ~n10991 ;
  assign n10994 = ~n10992 & n10993 ;
  assign n10995 = ~n10990 & ~n10994 ;
  assign n10996 = ~n10989 & n10995 ;
  assign n10997 = n1927 & ~n10996 ;
  assign n11003 = \P2_PhyAddrPointer_reg[1]/NET0131  & n8983 ;
  assign n11004 = ~\P2_PhyAddrPointer_reg[27]/NET0131  & ~n11003 ;
  assign n11005 = ~n8997 & ~n11004 ;
  assign n11006 = n3087 & n11005 ;
  assign n10998 = n8983 & ~n10965 ;
  assign n11000 = ~\P2_PhyAddrPointer_reg[27]/NET0131  & ~n10998 ;
  assign n10999 = \P2_PhyAddrPointer_reg[27]/NET0131  & n10998 ;
  assign n11001 = n1931 & ~n10999 ;
  assign n11002 = ~n11000 & n11001 ;
  assign n11007 = \P2_PhyAddrPointer_reg[27]/NET0131  & ~n8958 ;
  assign n11008 = \P2_rEIP_reg[27]/NET0131  & n3113 ;
  assign n11009 = ~n11007 & ~n11008 ;
  assign n11010 = ~n11002 & n11009 ;
  assign n11011 = ~n11006 & n11010 ;
  assign n11012 = ~n10997 & n11011 ;
  assign n11013 = \P2_PhyAddrPointer_reg[28]/NET0131  & n1897 ;
  assign n11020 = n6507 & n7432 ;
  assign n11021 = n7602 & n11020 ;
  assign n11022 = ~n6539 & n8912 ;
  assign n11023 = n11021 & n11022 ;
  assign n11024 = n10941 & n11023 ;
  assign n11025 = ~n6576 & n10976 ;
  assign n11026 = n11024 & n11025 ;
  assign n11028 = ~n6579 & n11026 ;
  assign n11027 = n6579 & ~n11026 ;
  assign n11029 = ~n6188 & ~n11027 ;
  assign n11030 = ~n11028 & n11029 ;
  assign n11017 = ~\P2_InstAddrPointer_reg[28]/NET0131  & n10983 ;
  assign n11014 = ~\P2_InstAddrPointer_reg[28]/NET0131  & ~n6584 ;
  assign n11015 = ~n6585 & ~n11014 ;
  assign n11016 = ~n10983 & n11015 ;
  assign n11018 = n6188 & ~n11016 ;
  assign n11019 = ~n11017 & n11018 ;
  assign n11031 = ~n1897 & ~n11019 ;
  assign n11032 = ~n11030 & n11031 ;
  assign n11033 = ~n11013 & ~n11032 ;
  assign n11034 = n1734 & ~n11033 ;
  assign n11035 = \P2_PhyAddrPointer_reg[28]/NET0131  & ~n8936 ;
  assign n11036 = ~\P2_InstAddrPointer_reg[28]/NET0131  & ~n6777 ;
  assign n11037 = ~n6785 & ~n11036 ;
  assign n11038 = \P2_InstAddrPointer_reg[15]/NET0131  & n7488 ;
  assign n11039 = n9245 & n11038 ;
  assign n11040 = ~\P2_InstAddrPointer_reg[16]/NET0131  & ~n6753 ;
  assign n11041 = ~n6754 & ~n11040 ;
  assign n11042 = n11039 & n11041 ;
  assign n11043 = n6758 & n11042 ;
  assign n11044 = ~\P2_InstAddrPointer_reg[20]/NET0131  & ~n6762 ;
  assign n11045 = ~n6763 & ~n11044 ;
  assign n11046 = \P2_InstAddrPointer_reg[21]/NET0131  & \P2_InstAddrPointer_reg[23]/NET0131  ;
  assign n11047 = n11045 & n11046 ;
  assign n11048 = n6770 & n11047 ;
  assign n11049 = n6778 & n11048 ;
  assign n11050 = n7626 & n11049 ;
  assign n11051 = n11043 & n11050 ;
  assign n11053 = n11037 & n11051 ;
  assign n11052 = ~n11037 & ~n11051 ;
  assign n11054 = n1890 & ~n11052 ;
  assign n11055 = ~n11053 & n11054 ;
  assign n11056 = ~n11035 & ~n11055 ;
  assign n11057 = ~n11034 & n11056 ;
  assign n11058 = n1927 & ~n11057 ;
  assign n11059 = ~\P2_PhyAddrPointer_reg[28]/NET0131  & ~n8984 ;
  assign n11060 = n3034 & ~n8985 ;
  assign n11061 = ~n11059 & n11060 ;
  assign n11062 = ~\P2_PhyAddrPointer_reg[28]/NET0131  & ~n8997 ;
  assign n11063 = ~n8998 & ~n11062 ;
  assign n11064 = n9005 & n11063 ;
  assign n11065 = \P2_rEIP_reg[28]/NET0131  & n3113 ;
  assign n11066 = \P2_PhyAddrPointer_reg[28]/NET0131  & ~n8958 ;
  assign n11067 = ~n11065 & ~n11066 ;
  assign n11068 = ~n11064 & n11067 ;
  assign n11069 = ~n11061 & n11068 ;
  assign n11070 = ~n11058 & n11069 ;
  assign n11071 = \P2_PhyAddrPointer_reg[29]/NET0131  & n1897 ;
  assign n11072 = ~n6687 & ~n11071 ;
  assign n11073 = n1734 & ~n11072 ;
  assign n11074 = \P2_PhyAddrPointer_reg[29]/NET0131  & ~n8936 ;
  assign n11075 = ~n6792 & ~n11074 ;
  assign n11076 = ~n11073 & n11075 ;
  assign n11077 = n1927 & ~n11076 ;
  assign n11081 = n8985 & ~n10965 ;
  assign n11083 = \P2_PhyAddrPointer_reg[29]/NET0131  & n11081 ;
  assign n11082 = ~\P2_PhyAddrPointer_reg[29]/NET0131  & ~n11081 ;
  assign n11084 = n1931 & ~n11082 ;
  assign n11085 = ~n11083 & n11084 ;
  assign n11078 = ~\P2_PhyAddrPointer_reg[29]/NET0131  & ~n8998 ;
  assign n11079 = ~n8999 & ~n11078 ;
  assign n11080 = n3087 & n11079 ;
  assign n11086 = \P2_PhyAddrPointer_reg[29]/NET0131  & ~n8958 ;
  assign n11087 = ~n6806 & ~n11086 ;
  assign n11088 = ~n11080 & n11087 ;
  assign n11089 = ~n11085 & n11088 ;
  assign n11090 = ~n11077 & n11089 ;
  assign n11108 = \P3_InstAddrPointer_reg[22]/NET0131  & n8378 ;
  assign n11112 = \P3_InstAddrPointer_reg[23]/NET0131  & n11108 ;
  assign n11109 = ~\P3_InstAddrPointer_reg[23]/NET0131  & ~n4370 ;
  assign n11110 = ~n4375 & ~n11109 ;
  assign n11111 = ~n11108 & ~n11110 ;
  assign n11113 = n2905 & ~n11111 ;
  assign n11114 = ~n11112 & n11113 ;
  assign n11091 = \P3_PhyAddrPointer_reg[23]/NET0131  & n2896 ;
  assign n11092 = n4250 & ~n4281 ;
  assign n11093 = n4258 & ~n4269 ;
  assign n11094 = n11092 & n11093 ;
  assign n11095 = n4265 & ~n11094 ;
  assign n11096 = n8394 & n11092 ;
  assign n11097 = ~n3753 & ~n11096 ;
  assign n11098 = ~n11095 & n11097 ;
  assign n11100 = ~n4087 & n4104 ;
  assign n11099 = n4087 & ~n4104 ;
  assign n11101 = n3753 & ~n11099 ;
  assign n11102 = ~n11100 & n11101 ;
  assign n11103 = ~n2896 & ~n11102 ;
  assign n11104 = ~n11098 & n11103 ;
  assign n11105 = ~n11091 & ~n11104 ;
  assign n11106 = n2894 & ~n11105 ;
  assign n11107 = \P3_PhyAddrPointer_reg[23]/NET0131  & ~n9014 ;
  assign n11115 = ~n11106 & ~n11107 ;
  assign n11116 = ~n11114 & n11115 ;
  assign n11117 = n2453 & ~n11116 ;
  assign n11124 = ~\P3_DataWidth_reg[1]/NET0131  & ~\P3_PhyAddrPointer_reg[1]/NET0131  ;
  assign n11125 = n9039 & ~n11124 ;
  assign n11127 = \P3_PhyAddrPointer_reg[23]/NET0131  & n11125 ;
  assign n11126 = ~\P3_PhyAddrPointer_reg[23]/NET0131  & ~n11125 ;
  assign n11128 = n2959 & ~n11126 ;
  assign n11129 = ~n11127 & n11128 ;
  assign n11118 = \P3_PhyAddrPointer_reg[1]/NET0131  & n9039 ;
  assign n11119 = ~\P3_PhyAddrPointer_reg[23]/NET0131  & ~n11118 ;
  assign n11120 = \P3_PhyAddrPointer_reg[23]/NET0131  & n9039 ;
  assign n11121 = \P3_PhyAddrPointer_reg[1]/NET0131  & n11120 ;
  assign n11122 = ~n11119 & ~n11121 ;
  assign n11123 = n4415 & n11122 ;
  assign n11130 = \P3_rEIP_reg[23]/NET0131  & n4412 ;
  assign n11131 = \P3_PhyAddrPointer_reg[23]/NET0131  & ~n9063 ;
  assign n11132 = ~n11130 & ~n11131 ;
  assign n11133 = ~n11123 & n11132 ;
  assign n11134 = ~n11129 & n11133 ;
  assign n11135 = ~n11117 & n11134 ;
  assign n11150 = n4374 & n4380 ;
  assign n11152 = n4388 & n11150 ;
  assign n11151 = ~n4388 & ~n11150 ;
  assign n11153 = n2905 & ~n11151 ;
  assign n11154 = ~n11152 & n11153 ;
  assign n11136 = \P3_PhyAddrPointer_reg[27]/NET0131  & n2896 ;
  assign n11142 = ~n4139 & n4283 ;
  assign n11141 = n4139 & ~n4283 ;
  assign n11143 = ~n3753 & ~n11141 ;
  assign n11144 = ~n11142 & n11143 ;
  assign n11138 = ~n4107 & n4112 ;
  assign n11137 = n4107 & ~n4112 ;
  assign n11139 = n3753 & ~n11137 ;
  assign n11140 = ~n11138 & n11139 ;
  assign n11145 = ~n2896 & ~n11140 ;
  assign n11146 = ~n11144 & n11145 ;
  assign n11147 = ~n11136 & ~n11146 ;
  assign n11148 = n2894 & ~n11147 ;
  assign n11149 = \P3_PhyAddrPointer_reg[27]/NET0131  & ~n9014 ;
  assign n11155 = ~n11148 & ~n11149 ;
  assign n11156 = ~n11154 & n11155 ;
  assign n11157 = n2453 & ~n11156 ;
  assign n11165 = ~\P3_PhyAddrPointer_reg[27]/NET0131  & ~n9044 ;
  assign n11166 = ~n9045 & ~n11165 ;
  assign n11167 = n4415 & n11166 ;
  assign n11159 = n9042 & n11125 ;
  assign n11161 = \P3_PhyAddrPointer_reg[27]/NET0131  & n11159 ;
  assign n11160 = ~\P3_PhyAddrPointer_reg[27]/NET0131  & ~n11159 ;
  assign n11162 = n2959 & ~n11160 ;
  assign n11163 = ~n11161 & n11162 ;
  assign n11158 = \P3_PhyAddrPointer_reg[27]/NET0131  & ~n9063 ;
  assign n11164 = \P3_rEIP_reg[27]/NET0131  & n4412 ;
  assign n11168 = ~n11158 & ~n11164 ;
  assign n11169 = ~n11163 & n11168 ;
  assign n11170 = ~n11167 & n11169 ;
  assign n11171 = ~n11157 & n11170 ;
  assign n11172 = \P3_PhyAddrPointer_reg[28]/NET0131  & n2896 ;
  assign n11173 = ~n6109 & ~n11172 ;
  assign n11174 = n2894 & ~n11173 ;
  assign n11175 = \P3_PhyAddrPointer_reg[28]/NET0131  & ~n9014 ;
  assign n11176 = ~n6135 & ~n11175 ;
  assign n11177 = ~n11174 & n11176 ;
  assign n11178 = n2453 & ~n11177 ;
  assign n11183 = ~\P3_PhyAddrPointer_reg[28]/NET0131  & ~n9045 ;
  assign n11184 = \P3_PhyAddrPointer_reg[28]/NET0131  & n9045 ;
  assign n11185 = ~n11183 & ~n11184 ;
  assign n11186 = n10076 & n11185 ;
  assign n11180 = ~\P3_PhyAddrPointer_reg[28]/NET0131  & ~n9049 ;
  assign n11179 = \P3_PhyAddrPointer_reg[28]/NET0131  & n9049 ;
  assign n11181 = n2970 & ~n11179 ;
  assign n11182 = ~n11180 & n11181 ;
  assign n11187 = \P3_PhyAddrPointer_reg[28]/NET0131  & ~n9063 ;
  assign n11188 = ~n6151 & ~n11187 ;
  assign n11189 = ~n11182 & n11188 ;
  assign n11190 = ~n11186 & n11189 ;
  assign n11191 = ~n11178 & n11190 ;
  assign n11192 = \P3_PhyAddrPointer_reg[29]/NET0131  & n2896 ;
  assign n11203 = n4143 & n4278 ;
  assign n11204 = n8344 & n11203 ;
  assign n11206 = ~n4146 & n11204 ;
  assign n11205 = n4146 & ~n11204 ;
  assign n11207 = ~n3753 & ~n11205 ;
  assign n11208 = ~n11206 & n11207 ;
  assign n11193 = ~\P3_InstAddrPointer_reg[29]/NET0131  & ~n6102 ;
  assign n11194 = n4109 & n4116 ;
  assign n11195 = ~n11193 & ~n11194 ;
  assign n11196 = n3790 & n4113 ;
  assign n11197 = n4106 & n11196 ;
  assign n11198 = n8347 & n11197 ;
  assign n11200 = ~n11195 & n11198 ;
  assign n11199 = n11195 & ~n11198 ;
  assign n11201 = n3753 & ~n11199 ;
  assign n11202 = ~n11200 & n11201 ;
  assign n11209 = ~n2896 & ~n11202 ;
  assign n11210 = ~n11208 & n11209 ;
  assign n11211 = ~n11192 & ~n11210 ;
  assign n11212 = n2894 & ~n11211 ;
  assign n11213 = \P3_PhyAddrPointer_reg[29]/NET0131  & ~n9014 ;
  assign n11214 = n4389 & n11150 ;
  assign n11215 = ~\P3_InstAddrPointer_reg[29]/NET0131  & ~n6113 ;
  assign n11216 = ~n4382 & ~n11215 ;
  assign n11217 = ~n11214 & ~n11216 ;
  assign n11218 = n4390 & n11150 ;
  assign n11219 = n2905 & ~n11218 ;
  assign n11220 = ~n11217 & n11219 ;
  assign n11221 = ~n11213 & ~n11220 ;
  assign n11222 = ~n11212 & n11221 ;
  assign n11223 = n2453 & ~n11222 ;
  assign n11224 = ~\P3_PhyAddrPointer_reg[29]/NET0131  & ~n11184 ;
  assign n11225 = ~n9046 & ~n11224 ;
  assign n11227 = ~\P3_DataWidth_reg[1]/NET0131  & ~n11225 ;
  assign n11228 = ~\P3_PhyAddrPointer_reg[29]/NET0131  & ~n11179 ;
  assign n11229 = ~n9050 & ~n11228 ;
  assign n11230 = \P3_DataWidth_reg[1]/NET0131  & ~n11229 ;
  assign n11231 = n2959 & ~n11230 ;
  assign n11232 = ~n11227 & n11231 ;
  assign n11226 = n4415 & n11225 ;
  assign n11233 = \P3_rEIP_reg[29]/NET0131  & n4412 ;
  assign n11234 = \P3_PhyAddrPointer_reg[29]/NET0131  & ~n9063 ;
  assign n11235 = ~n11233 & ~n11234 ;
  assign n11236 = ~n11226 & n11235 ;
  assign n11237 = ~n11232 & n11236 ;
  assign n11238 = ~n11223 & n11237 ;
  assign n11239 = \P1_PhyAddrPointer_reg[23]/NET0131  & n2375 ;
  assign n11240 = ~n6870 & ~n11239 ;
  assign n11241 = n2244 & ~n11240 ;
  assign n11242 = \P1_PhyAddrPointer_reg[23]/NET0131  & ~n10087 ;
  assign n11243 = ~n6885 & ~n11242 ;
  assign n11244 = ~n11241 & n11243 ;
  assign n11245 = n2432 & ~n11244 ;
  assign n11252 = \P1_PhyAddrPointer_reg[22]/NET0131  & n10125 ;
  assign n11253 = ~\P1_PhyAddrPointer_reg[23]/NET0131  & ~n11252 ;
  assign n11254 = n10111 & n10125 ;
  assign n11255 = ~n11253 & ~n11254 ;
  assign n11256 = n10133 & n11255 ;
  assign n11246 = \P1_PhyAddrPointer_reg[22]/NET0131  & n10110 ;
  assign n11247 = n3148 & ~n11246 ;
  assign n11248 = n10136 & ~n11247 ;
  assign n11249 = \P1_PhyAddrPointer_reg[23]/NET0131  & ~n11248 ;
  assign n11250 = ~\P1_PhyAddrPointer_reg[23]/NET0131  & n3148 ;
  assign n11251 = n11246 & n11250 ;
  assign n11257 = ~n6902 & ~n11251 ;
  assign n11258 = ~n11249 & n11257 ;
  assign n11259 = ~n11256 & n11258 ;
  assign n11260 = ~n11245 & n11259 ;
  assign n11261 = \P1_PhyAddrPointer_reg[27]/NET0131  & n2375 ;
  assign n11262 = n4488 & n6847 ;
  assign n11263 = n8545 & n11262 ;
  assign n11264 = ~n4492 & ~n11263 ;
  assign n11265 = n4487 & n7288 ;
  assign n11266 = n4492 & n11265 ;
  assign n11267 = n6839 & n11266 ;
  assign n11268 = n4453 & ~n11267 ;
  assign n11269 = ~n11264 & n11268 ;
  assign n11270 = ~n4928 & ~n4940 ;
  assign n11271 = n4909 & n11270 ;
  assign n11272 = ~n4926 & n11271 ;
  assign n11273 = n6861 & n11272 ;
  assign n11275 = n4942 & n11273 ;
  assign n11274 = ~n4942 & ~n11273 ;
  assign n11276 = ~n4453 & ~n11274 ;
  assign n11277 = ~n11275 & n11276 ;
  assign n11278 = ~n11269 & ~n11277 ;
  assign n11279 = ~n2375 & ~n11278 ;
  assign n11280 = ~n11261 & ~n11279 ;
  assign n11281 = n2244 & ~n11280 ;
  assign n11282 = \P1_PhyAddrPointer_reg[27]/NET0131  & ~n10087 ;
  assign n11283 = n6015 & n7298 ;
  assign n11284 = n6883 & n11283 ;
  assign n11286 = n5060 & n11284 ;
  assign n11285 = ~n5060 & ~n11284 ;
  assign n11287 = n2385 & ~n11285 ;
  assign n11288 = ~n11286 & n11287 ;
  assign n11289 = ~n11282 & ~n11288 ;
  assign n11290 = ~n11281 & n11289 ;
  assign n11291 = n2432 & ~n11290 ;
  assign n11296 = ~\P1_PhyAddrPointer_reg[27]/NET0131  & ~n10127 ;
  assign n11292 = \P1_PhyAddrPointer_reg[27]/NET0131  & n10115 ;
  assign n11297 = \P1_PhyAddrPointer_reg[1]/NET0131  & n11292 ;
  assign n11298 = ~n11296 & ~n11297 ;
  assign n11299 = n10133 & n11298 ;
  assign n11293 = ~\P1_PhyAddrPointer_reg[27]/NET0131  & ~n10115 ;
  assign n11294 = n3148 & ~n11292 ;
  assign n11295 = ~n11293 & n11294 ;
  assign n11300 = \P1_PhyAddrPointer_reg[27]/NET0131  & ~n10136 ;
  assign n11301 = \P1_rEIP_reg[27]/NET0131  & n5092 ;
  assign n11302 = ~n11300 & ~n11301 ;
  assign n11303 = ~n11295 & n11302 ;
  assign n11304 = ~n11299 & n11303 ;
  assign n11305 = ~n11291 & n11304 ;
  assign n11306 = \P1_PhyAddrPointer_reg[28]/NET0131  & n2375 ;
  assign n11313 = ~\P1_InstAddrPointer_reg[28]/NET0131  & ~n4490 ;
  assign n11314 = ~n5964 & ~n11313 ;
  assign n11316 = n11267 & ~n11314 ;
  assign n11315 = ~n11267 & n11314 ;
  assign n11317 = n4453 & ~n11315 ;
  assign n11318 = ~n11316 & n11317 ;
  assign n11307 = ~n4942 & n11271 ;
  assign n11308 = n7278 & n11307 ;
  assign n11310 = n4937 & ~n11308 ;
  assign n11309 = ~n4937 & n11308 ;
  assign n11311 = ~n4453 & ~n11309 ;
  assign n11312 = ~n11310 & n11311 ;
  assign n11319 = ~n2375 & ~n11312 ;
  assign n11320 = ~n11318 & n11319 ;
  assign n11321 = ~n11306 & ~n11320 ;
  assign n11322 = n2244 & ~n11321 ;
  assign n11323 = \P1_PhyAddrPointer_reg[28]/NET0131  & ~n10087 ;
  assign n11324 = n6016 & n7305 ;
  assign n11326 = n6018 & n11324 ;
  assign n11325 = ~n6018 & ~n11324 ;
  assign n11327 = n2385 & ~n11325 ;
  assign n11328 = ~n11326 & n11327 ;
  assign n11329 = ~n11323 & ~n11328 ;
  assign n11330 = ~n11322 & n11329 ;
  assign n11331 = n2432 & ~n11330 ;
  assign n11338 = ~\P1_PhyAddrPointer_reg[28]/NET0131  & ~n11297 ;
  assign n11339 = \P1_PhyAddrPointer_reg[28]/NET0131  & n11297 ;
  assign n11340 = ~n11338 & ~n11339 ;
  assign n11341 = n5095 & n11340 ;
  assign n11332 = ~\P1_DataWidth_reg[1]/NET0131  & ~\P1_PhyAddrPointer_reg[1]/NET0131  ;
  assign n11333 = n11292 & ~n11332 ;
  assign n11335 = \P1_PhyAddrPointer_reg[28]/NET0131  & n11333 ;
  assign n11334 = ~\P1_PhyAddrPointer_reg[28]/NET0131  & ~n11333 ;
  assign n11336 = n2436 & ~n11334 ;
  assign n11337 = ~n11335 & n11336 ;
  assign n11342 = \P1_rEIP_reg[28]/NET0131  & n5092 ;
  assign n11343 = \P1_PhyAddrPointer_reg[28]/NET0131  & ~n10136 ;
  assign n11344 = ~n11342 & ~n11343 ;
  assign n11345 = ~n11337 & n11344 ;
  assign n11346 = ~n11341 & n11345 ;
  assign n11347 = ~n11331 & n11346 ;
  assign n11348 = \P1_PhyAddrPointer_reg[29]/NET0131  & n2375 ;
  assign n11349 = ~n5984 & ~n11348 ;
  assign n11350 = n2244 & ~n11349 ;
  assign n11351 = \P1_PhyAddrPointer_reg[29]/NET0131  & ~n10087 ;
  assign n11352 = ~n6024 & ~n11351 ;
  assign n11353 = ~n11350 & n11352 ;
  assign n11354 = n2432 & ~n11353 ;
  assign n11360 = ~\P1_PhyAddrPointer_reg[29]/NET0131  & ~n11339 ;
  assign n11361 = ~n10128 & ~n11360 ;
  assign n11362 = n10133 & n11361 ;
  assign n11356 = \P1_PhyAddrPointer_reg[28]/NET0131  & n11292 ;
  assign n11357 = ~\P1_PhyAddrPointer_reg[29]/NET0131  & ~n11356 ;
  assign n11358 = n3148 & ~n10118 ;
  assign n11359 = ~n11357 & n11358 ;
  assign n11355 = \P1_PhyAddrPointer_reg[29]/NET0131  & ~n10136 ;
  assign n11363 = ~n6037 & ~n11355 ;
  assign n11364 = ~n11359 & n11363 ;
  assign n11365 = ~n11362 & n11364 ;
  assign n11366 = ~n11354 & n11365 ;
  assign n11378 = \P1_InstAddrPointer_reg[4]/NET0131  & n2375 ;
  assign n11384 = ~n4608 & ~n4751 ;
  assign n11385 = ~n6817 & ~n11384 ;
  assign n11386 = n6817 & n11384 ;
  assign n11387 = ~n11385 & ~n11386 ;
  assign n11388 = n4453 & ~n11387 ;
  assign n11379 = ~n4838 & ~n4859 ;
  assign n11381 = n4857 & n11379 ;
  assign n11380 = ~n4857 & ~n11379 ;
  assign n11382 = ~n4453 & ~n11380 ;
  assign n11383 = ~n11381 & n11382 ;
  assign n11389 = ~n2375 & ~n11383 ;
  assign n11390 = ~n11388 & n11389 ;
  assign n11391 = ~n11378 & ~n11390 ;
  assign n11392 = n2244 & ~n11391 ;
  assign n11377 = ~n2402 & n4576 ;
  assign n11373 = ~n2303 & ~n4456 ;
  assign n11374 = ~n2369 & ~n11373 ;
  assign n11375 = ~n2379 & n11374 ;
  assign n11376 = \P1_InstAddrPointer_reg[4]/NET0131  & ~n11375 ;
  assign n11393 = ~n2271 & n4837 ;
  assign n11369 = ~\P1_InstAddrPointer_reg[4]/NET0131  & ~n2337 ;
  assign n11370 = n2337 & ~n4988 ;
  assign n11371 = ~n11369 & ~n11370 ;
  assign n11372 = ~n2332 & n11371 ;
  assign n11394 = ~n4989 & ~n5008 ;
  assign n11396 = ~n5005 & n11394 ;
  assign n11395 = n5005 & ~n11394 ;
  assign n11397 = n2385 & ~n11395 ;
  assign n11398 = ~n11396 & n11397 ;
  assign n11399 = ~n11372 & ~n11398 ;
  assign n11400 = ~n11393 & n11399 ;
  assign n11401 = ~n11376 & n11400 ;
  assign n11402 = ~n11377 & n11401 ;
  assign n11403 = ~n11392 & n11402 ;
  assign n11404 = n2432 & ~n11403 ;
  assign n11367 = \P1_rEIP_reg[4]/NET0131  & n5092 ;
  assign n11368 = \P1_InstAddrPointer_reg[4]/NET0131  & ~n5098 ;
  assign n11405 = ~n11367 & ~n11368 ;
  assign n11406 = ~n11404 & n11405 ;
  assign n11412 = ~n4833 & ~n4865 ;
  assign n11413 = ~n4830 & ~n4862 ;
  assign n11414 = ~n11412 & ~n11413 ;
  assign n11415 = n11412 & n11413 ;
  assign n11416 = ~n11414 & ~n11415 ;
  assign n11417 = ~n4453 & ~n11416 ;
  assign n11418 = ~n4540 & ~n4759 ;
  assign n11419 = n6814 & n6817 ;
  assign n11420 = n6821 & ~n11419 ;
  assign n11422 = n11418 & n11420 ;
  assign n11421 = ~n11418 & ~n11420 ;
  assign n11423 = n4453 & ~n11421 ;
  assign n11424 = ~n11422 & n11423 ;
  assign n11425 = ~n11417 & ~n11424 ;
  assign n11426 = n2384 & n11425 ;
  assign n11427 = n2373 & ~n2379 ;
  assign n11428 = ~n2376 & n11427 ;
  assign n11429 = \P1_InstAddrPointer_reg[6]/NET0131  & ~n11428 ;
  assign n11430 = ~n4983 & ~n5015 ;
  assign n11432 = ~n5011 & n11430 ;
  assign n11431 = n5011 & ~n11430 ;
  assign n11433 = n2385 & ~n11431 ;
  assign n11434 = ~n11432 & n11433 ;
  assign n11409 = ~n2402 & n4508 ;
  assign n11410 = n2397 & n4982 ;
  assign n11411 = ~n2271 & n4832 ;
  assign n11435 = ~n11410 & ~n11411 ;
  assign n11436 = ~n11409 & n11435 ;
  assign n11437 = ~n11434 & n11436 ;
  assign n11438 = ~n11429 & n11437 ;
  assign n11439 = ~n11426 & n11438 ;
  assign n11440 = n2432 & ~n11439 ;
  assign n11407 = \P1_rEIP_reg[6]/NET0131  & n5092 ;
  assign n11408 = \P1_InstAddrPointer_reg[6]/NET0131  & ~n5098 ;
  assign n11441 = ~n11407 & ~n11408 ;
  assign n11442 = ~n11440 & n11441 ;
  assign n11445 = ~n3865 & ~n4050 ;
  assign n11446 = ~n6081 & n11445 ;
  assign n11447 = n6081 & ~n11445 ;
  assign n11448 = ~n11446 & ~n11447 ;
  assign n11449 = n2904 & n11448 ;
  assign n11454 = n2918 & n4312 ;
  assign n11460 = ~n11449 & ~n11454 ;
  assign n11450 = ~n2923 & n3833 ;
  assign n11453 = ~n2777 & n4181 ;
  assign n11461 = ~n11450 & ~n11453 ;
  assign n11462 = n11460 & n11461 ;
  assign n11451 = ~n2897 & n4402 ;
  assign n11452 = \P3_InstAddrPointer_reg[6]/NET0131  & ~n11451 ;
  assign n11455 = ~n4313 & ~n4341 ;
  assign n11457 = ~n6119 & n11455 ;
  assign n11456 = n6119 & ~n11455 ;
  assign n11458 = n2905 & ~n11456 ;
  assign n11459 = ~n11457 & n11458 ;
  assign n11463 = ~n11452 & ~n11459 ;
  assign n11464 = n11462 & n11463 ;
  assign n11465 = n2453 & ~n11464 ;
  assign n11443 = \P3_rEIP_reg[6]/NET0131  & n4412 ;
  assign n11444 = \P3_InstAddrPointer_reg[6]/NET0131  & ~n4418 ;
  assign n11466 = ~n11443 & ~n11444 ;
  assign n11467 = ~n11465 & n11466 ;
  assign n11480 = \P2_InstAddrPointer_reg[4]/NET0131  & n1897 ;
  assign n11486 = ~n6620 & ~n6628 ;
  assign n11487 = ~n7445 & n11486 ;
  assign n11488 = n7445 & ~n11486 ;
  assign n11489 = ~n11487 & ~n11488 ;
  assign n11490 = n6188 & ~n11489 ;
  assign n11481 = ~n6406 & ~n6445 ;
  assign n11483 = n7422 & n11481 ;
  assign n11482 = ~n7422 & ~n11481 ;
  assign n11484 = ~n6188 & ~n11482 ;
  assign n11485 = ~n11483 & n11484 ;
  assign n11491 = ~n1897 & ~n11485 ;
  assign n11492 = ~n11490 & n11491 ;
  assign n11493 = ~n11480 & ~n11492 ;
  assign n11494 = n1734 & ~n11493 ;
  assign n11470 = \P2_InstAddrPointer_reg[4]/NET0131  & ~n7501 ;
  assign n11478 = n1870 & n6706 ;
  assign n11495 = ~n11470 & ~n11478 ;
  assign n11479 = ~n1831 & n6619 ;
  assign n11471 = ~n1771 & n6374 ;
  assign n11472 = ~n6707 & ~n6721 ;
  assign n11473 = ~n6710 & ~n7539 ;
  assign n11475 = n11472 & n11473 ;
  assign n11474 = ~n11472 & ~n11473 ;
  assign n11476 = n1890 & ~n11474 ;
  assign n11477 = ~n11475 & n11476 ;
  assign n11496 = ~n11471 & ~n11477 ;
  assign n11497 = ~n11479 & n11496 ;
  assign n11498 = n11495 & n11497 ;
  assign n11499 = ~n11494 & n11498 ;
  assign n11500 = n1927 & ~n11499 ;
  assign n11468 = \P2_rEIP_reg[4]/NET0131  & n3113 ;
  assign n11469 = \P2_InstAddrPointer_reg[4]/NET0131  & ~n6810 ;
  assign n11501 = ~n11468 & ~n11469 ;
  assign n11502 = ~n11500 & n11501 ;
  assign n11504 = \P2_InstAddrPointer_reg[6]/NET0131  & n1897 ;
  assign n11510 = ~n6232 & ~n6451 ;
  assign n11511 = ~n6266 & ~n7425 ;
  assign n11512 = ~n11510 & ~n11511 ;
  assign n11513 = n11510 & n11511 ;
  assign n11514 = ~n11512 & ~n11513 ;
  assign n11515 = ~n6188 & ~n11514 ;
  assign n11505 = ~n6606 & ~n6636 ;
  assign n11507 = n7450 & n11505 ;
  assign n11506 = ~n7450 & ~n11505 ;
  assign n11508 = n6188 & ~n11506 ;
  assign n11509 = ~n11507 & n11508 ;
  assign n11516 = ~n1897 & ~n11509 ;
  assign n11517 = ~n11515 & n11516 ;
  assign n11518 = ~n11504 & ~n11517 ;
  assign n11519 = n1734 & ~n11518 ;
  assign n11524 = ~n6700 & ~n6727 ;
  assign n11525 = ~n6703 & ~n7542 ;
  assign n11527 = n11524 & n11525 ;
  assign n11526 = ~n11524 & ~n11525 ;
  assign n11528 = n1890 & ~n11526 ;
  assign n11529 = ~n11527 & n11528 ;
  assign n11520 = ~n1771 & n6200 ;
  assign n11523 = n1870 & n6699 ;
  assign n11530 = ~n11520 & ~n11523 ;
  assign n11521 = ~n1831 & n6605 ;
  assign n11522 = \P2_InstAddrPointer_reg[6]/NET0131  & ~n7501 ;
  assign n11531 = ~n11521 & ~n11522 ;
  assign n11532 = n11530 & n11531 ;
  assign n11533 = ~n11529 & n11532 ;
  assign n11534 = ~n11519 & n11533 ;
  assign n11535 = n1927 & ~n11534 ;
  assign n11503 = \P2_rEIP_reg[6]/NET0131  & n3113 ;
  assign n11536 = \P2_InstAddrPointer_reg[6]/NET0131  & ~n6810 ;
  assign n11537 = ~n11503 & ~n11536 ;
  assign n11538 = ~n11535 & n11537 ;
  assign n11547 = \buf2_reg[25]/NET0131  & ~n3079 ;
  assign n11548 = \buf1_reg[25]/NET0131  & n3079 ;
  assign n11549 = ~n11547 & ~n11548 ;
  assign n11550 = n3091 & ~n11549 ;
  assign n11551 = \buf2_reg[17]/NET0131  & ~n3079 ;
  assign n11552 = \buf1_reg[17]/NET0131  & n3079 ;
  assign n11553 = ~n11551 & ~n11552 ;
  assign n11554 = n3098 & ~n11553 ;
  assign n11555 = ~n11550 & ~n11554 ;
  assign n11556 = \P2_DataWidth_reg[1]/NET0131  & ~n11555 ;
  assign n11539 = \buf2_reg[1]/NET0131  & ~n3079 ;
  assign n11540 = \buf1_reg[1]/NET0131  & n3079 ;
  assign n11541 = ~n11539 & ~n11540 ;
  assign n11542 = ~n3050 & ~n11541 ;
  assign n11543 = \P2_InstQueue_reg[11][1]/NET0131  & ~n3049 ;
  assign n11544 = ~n3046 & n11543 ;
  assign n11545 = ~n11542 & ~n11544 ;
  assign n11557 = ~n3106 & ~n11545 ;
  assign n11558 = ~n11556 & ~n11557 ;
  assign n11559 = n1931 & ~n11558 ;
  assign n11546 = n3087 & ~n11545 ;
  assign n11560 = ~n1592 & n3049 ;
  assign n11561 = ~n11543 & ~n11560 ;
  assign n11562 = n3040 & ~n11561 ;
  assign n11563 = \P2_InstQueue_reg[11][1]/NET0131  & ~n3118 ;
  assign n11564 = ~n11562 & ~n11563 ;
  assign n11565 = ~n11546 & n11564 ;
  assign n11566 = ~n11559 & n11565 ;
  assign n11572 = n3162 & ~n11549 ;
  assign n11573 = n3165 & ~n11553 ;
  assign n11574 = ~n11572 & ~n11573 ;
  assign n11575 = \P2_DataWidth_reg[1]/NET0131  & ~n11574 ;
  assign n11567 = ~n3155 & ~n11541 ;
  assign n11568 = \P2_InstQueue_reg[0][1]/NET0131  & ~n3152 ;
  assign n11569 = ~n3154 & n11568 ;
  assign n11570 = ~n11567 & ~n11569 ;
  assign n11576 = ~n3170 & ~n11570 ;
  assign n11577 = ~n11575 & ~n11576 ;
  assign n11578 = n1931 & ~n11577 ;
  assign n11571 = n3087 & ~n11570 ;
  assign n11579 = ~n1592 & n3152 ;
  assign n11580 = ~n11568 & ~n11579 ;
  assign n11581 = n3040 & ~n11580 ;
  assign n11582 = \P2_InstQueue_reg[0][1]/NET0131  & ~n3118 ;
  assign n11583 = ~n11581 & ~n11582 ;
  assign n11584 = ~n11571 & n11583 ;
  assign n11585 = ~n11578 & n11584 ;
  assign n11591 = n3091 & ~n11553 ;
  assign n11592 = n3198 & ~n11549 ;
  assign n11593 = ~n11591 & ~n11592 ;
  assign n11594 = \P2_DataWidth_reg[1]/NET0131  & ~n11593 ;
  assign n11586 = ~n3202 & ~n11541 ;
  assign n11587 = \P2_InstQueue_reg[10][1]/NET0131  & ~n3046 ;
  assign n11588 = ~n3098 & n11587 ;
  assign n11589 = ~n11586 & ~n11588 ;
  assign n11595 = ~n3200 & ~n11589 ;
  assign n11596 = ~n11594 & ~n11595 ;
  assign n11597 = n1931 & ~n11596 ;
  assign n11590 = n3087 & ~n11589 ;
  assign n11598 = ~n1592 & n3046 ;
  assign n11599 = ~n11587 & ~n11598 ;
  assign n11600 = n3040 & ~n11599 ;
  assign n11601 = \P2_InstQueue_reg[10][1]/NET0131  & ~n3118 ;
  assign n11602 = ~n11600 & ~n11601 ;
  assign n11603 = ~n11590 & n11602 ;
  assign n11604 = ~n11597 & n11603 ;
  assign n11610 = n3098 & ~n11549 ;
  assign n11611 = n3046 & ~n11553 ;
  assign n11612 = ~n11610 & ~n11611 ;
  assign n11613 = \P2_DataWidth_reg[1]/NET0131  & ~n11612 ;
  assign n11605 = ~n3238 & ~n11541 ;
  assign n11606 = \P2_InstQueue_reg[12][1]/NET0131  & ~n3237 ;
  assign n11607 = ~n3049 & n11606 ;
  assign n11608 = ~n11605 & ~n11607 ;
  assign n11614 = ~n3248 & ~n11608 ;
  assign n11615 = ~n11613 & ~n11614 ;
  assign n11616 = n1931 & ~n11615 ;
  assign n11609 = n3087 & ~n11608 ;
  assign n11617 = ~n1592 & n3237 ;
  assign n11618 = ~n11606 & ~n11617 ;
  assign n11619 = n3040 & ~n11618 ;
  assign n11620 = \P2_InstQueue_reg[12][1]/NET0131  & ~n3118 ;
  assign n11621 = ~n11619 & ~n11620 ;
  assign n11622 = ~n11609 & n11621 ;
  assign n11623 = ~n11616 & n11622 ;
  assign n11629 = n3046 & ~n11549 ;
  assign n11630 = n3049 & ~n11553 ;
  assign n11631 = ~n11629 & ~n11630 ;
  assign n11632 = \P2_DataWidth_reg[1]/NET0131  & ~n11631 ;
  assign n11624 = ~n3275 & ~n11541 ;
  assign n11625 = \P2_InstQueue_reg[13][1]/NET0131  & ~n3162 ;
  assign n11626 = ~n3237 & n11625 ;
  assign n11627 = ~n11624 & ~n11626 ;
  assign n11633 = ~n3285 & ~n11627 ;
  assign n11634 = ~n11632 & ~n11633 ;
  assign n11635 = n1931 & ~n11634 ;
  assign n11628 = n3087 & ~n11627 ;
  assign n11636 = ~n1592 & n3162 ;
  assign n11637 = ~n11625 & ~n11636 ;
  assign n11638 = n3040 & ~n11637 ;
  assign n11639 = \P2_InstQueue_reg[13][1]/NET0131  & ~n3118 ;
  assign n11640 = ~n11638 & ~n11639 ;
  assign n11641 = ~n11628 & n11640 ;
  assign n11642 = ~n11635 & n11641 ;
  assign n11648 = n3049 & ~n11549 ;
  assign n11649 = n3237 & ~n11553 ;
  assign n11650 = ~n11648 & ~n11649 ;
  assign n11651 = \P2_DataWidth_reg[1]/NET0131  & ~n11650 ;
  assign n11643 = ~n3169 & ~n11541 ;
  assign n11644 = \P2_InstQueue_reg[14][1]/NET0131  & ~n3165 ;
  assign n11645 = ~n3162 & n11644 ;
  assign n11646 = ~n11643 & ~n11645 ;
  assign n11652 = ~n3321 & ~n11646 ;
  assign n11653 = ~n11651 & ~n11652 ;
  assign n11654 = n1931 & ~n11653 ;
  assign n11647 = n3087 & ~n11646 ;
  assign n11655 = ~n1592 & n3165 ;
  assign n11656 = ~n11644 & ~n11655 ;
  assign n11657 = n3040 & ~n11656 ;
  assign n11658 = \P2_InstQueue_reg[14][1]/NET0131  & ~n3118 ;
  assign n11659 = ~n11657 & ~n11658 ;
  assign n11660 = ~n11647 & n11659 ;
  assign n11661 = ~n11654 & n11660 ;
  assign n11667 = n3237 & ~n11549 ;
  assign n11668 = n3162 & ~n11553 ;
  assign n11669 = ~n11667 & ~n11668 ;
  assign n11670 = \P2_DataWidth_reg[1]/NET0131  & ~n11669 ;
  assign n11662 = ~n3348 & ~n11541 ;
  assign n11663 = \P2_InstQueue_reg[15][1]/NET0131  & ~n3154 ;
  assign n11664 = ~n3165 & n11663 ;
  assign n11665 = ~n11662 & ~n11664 ;
  assign n11671 = ~n3358 & ~n11665 ;
  assign n11672 = ~n11670 & ~n11671 ;
  assign n11673 = n1931 & ~n11672 ;
  assign n11666 = n3087 & ~n11665 ;
  assign n11674 = ~n1592 & n3154 ;
  assign n11675 = ~n11663 & ~n11674 ;
  assign n11676 = n3040 & ~n11675 ;
  assign n11677 = \P2_InstQueue_reg[15][1]/NET0131  & ~n3118 ;
  assign n11678 = ~n11676 & ~n11677 ;
  assign n11679 = ~n11666 & n11678 ;
  assign n11680 = ~n11673 & n11679 ;
  assign n11686 = n3165 & ~n11549 ;
  assign n11687 = n3154 & ~n11553 ;
  assign n11688 = ~n11686 & ~n11687 ;
  assign n11689 = \P2_DataWidth_reg[1]/NET0131  & ~n11688 ;
  assign n11681 = ~n3389 & ~n11541 ;
  assign n11682 = \P2_InstQueue_reg[1][1]/NET0131  & ~n3388 ;
  assign n11683 = ~n3152 & n11682 ;
  assign n11684 = ~n11681 & ~n11683 ;
  assign n11690 = ~n3386 & ~n11684 ;
  assign n11691 = ~n11689 & ~n11690 ;
  assign n11692 = n1931 & ~n11691 ;
  assign n11685 = n3087 & ~n11684 ;
  assign n11693 = ~n1592 & n3388 ;
  assign n11694 = ~n11682 & ~n11693 ;
  assign n11695 = n3040 & ~n11694 ;
  assign n11696 = \P2_InstQueue_reg[1][1]/NET0131  & ~n3118 ;
  assign n11697 = ~n11695 & ~n11696 ;
  assign n11698 = ~n11685 & n11697 ;
  assign n11699 = ~n11692 & n11698 ;
  assign n11705 = n3152 & ~n11553 ;
  assign n11706 = n3154 & ~n11549 ;
  assign n11707 = ~n11705 & ~n11706 ;
  assign n11708 = \P2_DataWidth_reg[1]/NET0131  & ~n11707 ;
  assign n11700 = ~n3424 & ~n11541 ;
  assign n11701 = \P2_InstQueue_reg[2][1]/NET0131  & ~n3423 ;
  assign n11702 = ~n3388 & n11701 ;
  assign n11703 = ~n11700 & ~n11702 ;
  assign n11709 = ~n3434 & ~n11703 ;
  assign n11710 = ~n11708 & ~n11709 ;
  assign n11711 = n1931 & ~n11710 ;
  assign n11704 = n3087 & ~n11703 ;
  assign n11712 = ~n1592 & n3423 ;
  assign n11713 = ~n11701 & ~n11712 ;
  assign n11714 = n3040 & ~n11713 ;
  assign n11715 = \P2_InstQueue_reg[2][1]/NET0131  & ~n3118 ;
  assign n11716 = ~n11714 & ~n11715 ;
  assign n11717 = ~n11704 & n11716 ;
  assign n11718 = ~n11711 & n11717 ;
  assign n11724 = n3152 & ~n11549 ;
  assign n11725 = n3388 & ~n11553 ;
  assign n11726 = ~n11724 & ~n11725 ;
  assign n11727 = \P2_DataWidth_reg[1]/NET0131  & ~n11726 ;
  assign n11719 = ~n3462 & ~n11541 ;
  assign n11720 = \P2_InstQueue_reg[3][1]/NET0131  & ~n3461 ;
  assign n11721 = ~n3423 & n11720 ;
  assign n11722 = ~n11719 & ~n11721 ;
  assign n11728 = ~n3472 & ~n11722 ;
  assign n11729 = ~n11727 & ~n11728 ;
  assign n11730 = n1931 & ~n11729 ;
  assign n11723 = n3087 & ~n11722 ;
  assign n11731 = ~n1592 & n3461 ;
  assign n11732 = ~n11720 & ~n11731 ;
  assign n11733 = n3040 & ~n11732 ;
  assign n11734 = \P2_InstQueue_reg[3][1]/NET0131  & ~n3118 ;
  assign n11735 = ~n11733 & ~n11734 ;
  assign n11736 = ~n11723 & n11735 ;
  assign n11737 = ~n11730 & n11736 ;
  assign n11743 = n3388 & ~n11549 ;
  assign n11744 = n3423 & ~n11553 ;
  assign n11745 = ~n11743 & ~n11744 ;
  assign n11746 = \P2_DataWidth_reg[1]/NET0131  & ~n11745 ;
  assign n11738 = ~n3500 & ~n11541 ;
  assign n11739 = \P2_InstQueue_reg[4][1]/NET0131  & ~n3499 ;
  assign n11740 = ~n3461 & n11739 ;
  assign n11741 = ~n11738 & ~n11740 ;
  assign n11747 = ~n3510 & ~n11741 ;
  assign n11748 = ~n11746 & ~n11747 ;
  assign n11749 = n1931 & ~n11748 ;
  assign n11742 = n3087 & ~n11741 ;
  assign n11750 = ~n1592 & n3499 ;
  assign n11751 = ~n11739 & ~n11750 ;
  assign n11752 = n3040 & ~n11751 ;
  assign n11753 = \P2_InstQueue_reg[4][1]/NET0131  & ~n3118 ;
  assign n11754 = ~n11752 & ~n11753 ;
  assign n11755 = ~n11742 & n11754 ;
  assign n11756 = ~n11749 & n11755 ;
  assign n11762 = n3423 & ~n11549 ;
  assign n11763 = n3461 & ~n11553 ;
  assign n11764 = ~n11762 & ~n11763 ;
  assign n11765 = \P2_DataWidth_reg[1]/NET0131  & ~n11764 ;
  assign n11757 = ~n3538 & ~n11541 ;
  assign n11758 = \P2_InstQueue_reg[5][1]/NET0131  & ~n3537 ;
  assign n11759 = ~n3499 & n11758 ;
  assign n11760 = ~n11757 & ~n11759 ;
  assign n11766 = ~n3548 & ~n11760 ;
  assign n11767 = ~n11765 & ~n11766 ;
  assign n11768 = n1931 & ~n11767 ;
  assign n11761 = n3087 & ~n11760 ;
  assign n11769 = ~n1592 & n3537 ;
  assign n11770 = ~n11758 & ~n11769 ;
  assign n11771 = n3040 & ~n11770 ;
  assign n11772 = \P2_InstQueue_reg[5][1]/NET0131  & ~n3118 ;
  assign n11773 = ~n11771 & ~n11772 ;
  assign n11774 = ~n11761 & n11773 ;
  assign n11775 = ~n11768 & n11774 ;
  assign n11781 = n3461 & ~n11549 ;
  assign n11782 = n3499 & ~n11553 ;
  assign n11783 = ~n11781 & ~n11782 ;
  assign n11784 = \P2_DataWidth_reg[1]/NET0131  & ~n11783 ;
  assign n11776 = ~n3576 & ~n11541 ;
  assign n11777 = \P2_InstQueue_reg[6][1]/NET0131  & ~n3575 ;
  assign n11778 = ~n3537 & n11777 ;
  assign n11779 = ~n11776 & ~n11778 ;
  assign n11785 = ~n3586 & ~n11779 ;
  assign n11786 = ~n11784 & ~n11785 ;
  assign n11787 = n1931 & ~n11786 ;
  assign n11780 = n3087 & ~n11779 ;
  assign n11788 = ~n1592 & n3575 ;
  assign n11789 = ~n11777 & ~n11788 ;
  assign n11790 = n3040 & ~n11789 ;
  assign n11791 = \P2_InstQueue_reg[6][1]/NET0131  & ~n3118 ;
  assign n11792 = ~n11790 & ~n11791 ;
  assign n11793 = ~n11780 & n11792 ;
  assign n11794 = ~n11787 & n11793 ;
  assign n11800 = n3499 & ~n11549 ;
  assign n11801 = n3537 & ~n11553 ;
  assign n11802 = ~n11800 & ~n11801 ;
  assign n11803 = \P2_DataWidth_reg[1]/NET0131  & ~n11802 ;
  assign n11795 = ~n3613 & ~n11541 ;
  assign n11796 = \P2_InstQueue_reg[7][1]/NET0131  & ~n3198 ;
  assign n11797 = ~n3575 & n11796 ;
  assign n11798 = ~n11795 & ~n11797 ;
  assign n11804 = ~n3623 & ~n11798 ;
  assign n11805 = ~n11803 & ~n11804 ;
  assign n11806 = n1931 & ~n11805 ;
  assign n11799 = n3087 & ~n11798 ;
  assign n11807 = ~n1592 & n3198 ;
  assign n11808 = ~n11796 & ~n11807 ;
  assign n11809 = n3040 & ~n11808 ;
  assign n11810 = \P2_InstQueue_reg[7][1]/NET0131  & ~n3118 ;
  assign n11811 = ~n11809 & ~n11810 ;
  assign n11812 = ~n11799 & n11811 ;
  assign n11813 = ~n11806 & n11812 ;
  assign n11819 = n3537 & ~n11549 ;
  assign n11820 = n3575 & ~n11553 ;
  assign n11821 = ~n11819 & ~n11820 ;
  assign n11822 = \P2_DataWidth_reg[1]/NET0131  & ~n11821 ;
  assign n11814 = ~n3199 & ~n11541 ;
  assign n11815 = \P2_InstQueue_reg[8][1]/NET0131  & ~n3091 ;
  assign n11816 = ~n3198 & n11815 ;
  assign n11817 = ~n11814 & ~n11816 ;
  assign n11823 = ~n3659 & ~n11817 ;
  assign n11824 = ~n11822 & ~n11823 ;
  assign n11825 = n1931 & ~n11824 ;
  assign n11818 = n3087 & ~n11817 ;
  assign n11826 = ~n1592 & n3091 ;
  assign n11827 = ~n11815 & ~n11826 ;
  assign n11828 = n3040 & ~n11827 ;
  assign n11829 = \P2_InstQueue_reg[8][1]/NET0131  & ~n3118 ;
  assign n11830 = ~n11828 & ~n11829 ;
  assign n11831 = ~n11818 & n11830 ;
  assign n11832 = ~n11825 & n11831 ;
  assign n11838 = n3575 & ~n11549 ;
  assign n11839 = n3198 & ~n11553 ;
  assign n11840 = ~n11838 & ~n11839 ;
  assign n11841 = \P2_DataWidth_reg[1]/NET0131  & ~n11840 ;
  assign n11833 = ~n3105 & ~n11541 ;
  assign n11834 = \P2_InstQueue_reg[9][1]/NET0131  & ~n3098 ;
  assign n11835 = ~n3091 & n11834 ;
  assign n11836 = ~n11833 & ~n11835 ;
  assign n11842 = ~n3695 & ~n11836 ;
  assign n11843 = ~n11841 & ~n11842 ;
  assign n11844 = n1931 & ~n11843 ;
  assign n11837 = n3087 & ~n11836 ;
  assign n11845 = ~n1592 & n3098 ;
  assign n11846 = ~n11834 & ~n11845 ;
  assign n11847 = n3040 & ~n11846 ;
  assign n11848 = \P2_InstQueue_reg[9][1]/NET0131  & ~n3118 ;
  assign n11849 = ~n11847 & ~n11848 ;
  assign n11850 = ~n11837 & n11849 ;
  assign n11851 = ~n11844 & n11850 ;
  assign n11852 = \P2_PhyAddrPointer_reg[20]/NET0131  & n1897 ;
  assign n11853 = n6537 & ~n11023 ;
  assign n11854 = ~n6188 & ~n7517 ;
  assign n11855 = ~n11853 & n11854 ;
  assign n11856 = ~n6666 & ~n7525 ;
  assign n11857 = ~n6669 & ~n11856 ;
  assign n11858 = n6188 & ~n11857 ;
  assign n11859 = ~n1897 & ~n11858 ;
  assign n11860 = ~n11855 & n11859 ;
  assign n11861 = ~n11852 & ~n11860 ;
  assign n11862 = n1734 & ~n11861 ;
  assign n11863 = \P2_PhyAddrPointer_reg[20]/NET0131  & ~n8936 ;
  assign n11865 = ~n11043 & ~n11045 ;
  assign n11864 = n6759 & n11042 ;
  assign n11866 = n1890 & ~n11864 ;
  assign n11867 = ~n11865 & n11866 ;
  assign n11868 = ~n11863 & ~n11867 ;
  assign n11869 = ~n11862 & n11868 ;
  assign n11870 = n1927 & ~n11869 ;
  assign n11874 = \P2_PhyAddrPointer_reg[1]/NET0131  & n8976 ;
  assign n11875 = ~\P2_PhyAddrPointer_reg[20]/NET0131  & ~n11874 ;
  assign n11876 = \P2_PhyAddrPointer_reg[1]/NET0131  & n8977 ;
  assign n11877 = ~n11875 & ~n11876 ;
  assign n11878 = n9005 & n11877 ;
  assign n11871 = ~\P2_PhyAddrPointer_reg[20]/NET0131  & ~n8976 ;
  assign n11872 = n3034 & ~n8977 ;
  assign n11873 = ~n11871 & n11872 ;
  assign n11879 = \P2_PhyAddrPointer_reg[20]/NET0131  & ~n8958 ;
  assign n11880 = \P2_rEIP_reg[20]/NET0131  & n3113 ;
  assign n11881 = ~n11879 & ~n11880 ;
  assign n11882 = ~n11873 & n11881 ;
  assign n11883 = ~n11878 & n11882 ;
  assign n11884 = ~n11870 & n11883 ;
  assign n11885 = \P2_PhyAddrPointer_reg[22]/NET0131  & n1897 ;
  assign n11886 = ~n7533 & ~n11885 ;
  assign n11887 = n1734 & ~n11886 ;
  assign n11888 = \P2_PhyAddrPointer_reg[22]/NET0131  & ~n8936 ;
  assign n11889 = ~n7559 & ~n11888 ;
  assign n11890 = ~n11887 & n11889 ;
  assign n11891 = n1927 & ~n11890 ;
  assign n11892 = \P2_PhyAddrPointer_reg[21]/NET0131  & n8977 ;
  assign n11896 = \P2_PhyAddrPointer_reg[1]/NET0131  & n11892 ;
  assign n11897 = ~\P2_PhyAddrPointer_reg[22]/NET0131  & ~n11896 ;
  assign n11898 = ~n10959 & ~n11897 ;
  assign n11899 = n9005 & n11898 ;
  assign n11893 = ~\P2_PhyAddrPointer_reg[22]/NET0131  & ~n11892 ;
  assign n11894 = n3034 & ~n8979 ;
  assign n11895 = ~n11893 & n11894 ;
  assign n11900 = \P2_PhyAddrPointer_reg[22]/NET0131  & ~n8958 ;
  assign n11901 = ~n7581 & ~n11900 ;
  assign n11902 = ~n11895 & n11901 ;
  assign n11903 = ~n11899 & n11902 ;
  assign n11904 = ~n11891 & n11903 ;
  assign n11905 = \P2_PhyAddrPointer_reg[24]/NET0131  & n1897 ;
  assign n11910 = ~\P2_InstAddrPointer_reg[24]/NET0131  & ~n10930 ;
  assign n11911 = ~n6558 & ~n11910 ;
  assign n11912 = \P2_InstAddrPointer_reg[23]/NET0131  & n6597 ;
  assign n11913 = n7527 & n11912 ;
  assign n11914 = ~n11911 & ~n11913 ;
  assign n11915 = ~n6671 & ~n11914 ;
  assign n11916 = n6188 & ~n11915 ;
  assign n11906 = ~n6560 & ~n11024 ;
  assign n11907 = n6560 & n11024 ;
  assign n11908 = ~n11906 & ~n11907 ;
  assign n11909 = ~n6188 & ~n11908 ;
  assign n11917 = ~n1897 & ~n11909 ;
  assign n11918 = ~n11916 & n11917 ;
  assign n11919 = ~n11905 & ~n11918 ;
  assign n11920 = n1734 & ~n11919 ;
  assign n11921 = \P2_PhyAddrPointer_reg[24]/NET0131  & ~n8936 ;
  assign n11922 = n11043 & n11048 ;
  assign n11924 = n7625 & n11922 ;
  assign n11923 = ~n7625 & ~n11922 ;
  assign n11925 = n1890 & ~n11923 ;
  assign n11926 = ~n11924 & n11925 ;
  assign n11927 = ~n11921 & ~n11926 ;
  assign n11928 = ~n11920 & n11927 ;
  assign n11929 = n1927 & ~n11928 ;
  assign n11933 = ~\P2_PhyAddrPointer_reg[24]/NET0131  & ~n10961 ;
  assign n11934 = ~n8995 & ~n11933 ;
  assign n11935 = n9005 & n11934 ;
  assign n11930 = ~\P2_PhyAddrPointer_reg[24]/NET0131  & ~n8980 ;
  assign n11931 = n3034 & ~n8981 ;
  assign n11932 = ~n11930 & n11931 ;
  assign n11936 = \P2_PhyAddrPointer_reg[24]/NET0131  & ~n8958 ;
  assign n11937 = \P2_rEIP_reg[24]/NET0131  & n3113 ;
  assign n11938 = ~n11936 & ~n11937 ;
  assign n11939 = ~n11932 & n11938 ;
  assign n11940 = ~n11935 & n11939 ;
  assign n11941 = ~n11929 & n11940 ;
  assign n11942 = \P2_PhyAddrPointer_reg[26]/NET0131  & n1897 ;
  assign n11943 = ~n7613 & ~n11942 ;
  assign n11944 = n1734 & ~n11943 ;
  assign n11945 = \P2_PhyAddrPointer_reg[26]/NET0131  & ~n8936 ;
  assign n11946 = ~n7630 & ~n11945 ;
  assign n11947 = ~n11944 & n11946 ;
  assign n11948 = n1927 & ~n11947 ;
  assign n11952 = ~\P2_PhyAddrPointer_reg[26]/NET0131  & ~n8996 ;
  assign n11953 = ~n11003 & ~n11952 ;
  assign n11954 = n9005 & n11953 ;
  assign n11949 = ~\P2_PhyAddrPointer_reg[26]/NET0131  & ~n8982 ;
  assign n11950 = n3034 & ~n8983 ;
  assign n11951 = ~n11949 & n11950 ;
  assign n11955 = \P2_PhyAddrPointer_reg[26]/NET0131  & ~n8958 ;
  assign n11956 = ~n7654 & ~n11955 ;
  assign n11957 = ~n11951 & n11956 ;
  assign n11958 = ~n11954 & n11957 ;
  assign n11959 = ~n11948 & n11958 ;
  assign n11978 = n4301 & n10203 ;
  assign n11982 = \P3_InstAddrPointer_reg[11]/NET0131  & n11978 ;
  assign n11979 = ~\P3_InstAddrPointer_reg[11]/NET0131  & ~n4299 ;
  assign n11980 = ~n9097 & ~n11979 ;
  assign n11981 = ~n11978 & ~n11980 ;
  assign n11983 = n2905 & ~n11981 ;
  assign n11984 = ~n11982 & n11983 ;
  assign n11965 = ~n2897 & n9014 ;
  assign n11966 = \P3_PhyAddrPointer_reg[11]/NET0131  & ~n11965 ;
  assign n11971 = n4063 & n10148 ;
  assign n11972 = ~n4069 & ~n11971 ;
  assign n11973 = ~n6088 & ~n11972 ;
  assign n11974 = n3753 & ~n11973 ;
  assign n11967 = ~n4158 & ~n4230 ;
  assign n11968 = n4158 & n4230 ;
  assign n11969 = ~n11967 & ~n11968 ;
  assign n11970 = ~n3753 & ~n11969 ;
  assign n11975 = ~n2896 & ~n11970 ;
  assign n11976 = ~n11974 & n11975 ;
  assign n11977 = n2894 & n11976 ;
  assign n11985 = ~n11966 & ~n11977 ;
  assign n11986 = ~n11984 & n11985 ;
  assign n11987 = n2453 & ~n11986 ;
  assign n11960 = \P3_PhyAddrPointer_reg[1]/NET0131  & n9027 ;
  assign n11961 = ~\P3_PhyAddrPointer_reg[11]/NET0131  & ~n11960 ;
  assign n11962 = \P3_PhyAddrPointer_reg[1]/NET0131  & n9028 ;
  assign n11963 = ~n11961 & ~n11962 ;
  assign n11988 = ~\P3_DataWidth_reg[1]/NET0131  & ~n11963 ;
  assign n11989 = ~\P3_PhyAddrPointer_reg[11]/NET0131  & ~n9027 ;
  assign n11990 = ~n9028 & ~n11989 ;
  assign n11991 = \P3_DataWidth_reg[1]/NET0131  & ~n11990 ;
  assign n11992 = n2959 & ~n11991 ;
  assign n11993 = ~n11988 & n11992 ;
  assign n11964 = n4415 & n11963 ;
  assign n11994 = \P3_rEIP_reg[11]/NET0131  & n4412 ;
  assign n11995 = \P3_PhyAddrPointer_reg[11]/NET0131  & ~n9063 ;
  assign n11996 = ~n11994 & ~n11995 ;
  assign n11997 = ~n11964 & n11996 ;
  assign n11998 = ~n11993 & n11997 ;
  assign n11999 = ~n11987 & n11998 ;
  assign n12015 = \P3_PhyAddrPointer_reg[15]/NET0131  & n2896 ;
  assign n12016 = ~n7341 & ~n12015 ;
  assign n12017 = n2894 & ~n12016 ;
  assign n12018 = \P3_PhyAddrPointer_reg[15]/NET0131  & ~n9014 ;
  assign n12019 = ~n7355 & ~n12018 ;
  assign n12020 = ~n12017 & n12019 ;
  assign n12021 = n2453 & ~n12020 ;
  assign n12007 = \P3_PhyAddrPointer_reg[12]/NET0131  & n11962 ;
  assign n12008 = \P3_PhyAddrPointer_reg[13]/NET0131  & n12007 ;
  assign n12009 = \P3_PhyAddrPointer_reg[14]/NET0131  & n12008 ;
  assign n12010 = ~\P3_PhyAddrPointer_reg[15]/NET0131  & ~n12009 ;
  assign n12011 = n9030 & n9031 ;
  assign n12012 = \P3_PhyAddrPointer_reg[1]/NET0131  & n12011 ;
  assign n12013 = ~n12010 & ~n12012 ;
  assign n12014 = n4415 & n12013 ;
  assign n12000 = n9030 & ~n11124 ;
  assign n12001 = \P3_PhyAddrPointer_reg[14]/NET0131  & n12000 ;
  assign n12002 = n2959 & ~n12001 ;
  assign n12003 = n9063 & ~n12002 ;
  assign n12004 = \P3_PhyAddrPointer_reg[15]/NET0131  & ~n12003 ;
  assign n12005 = ~\P3_PhyAddrPointer_reg[15]/NET0131  & n2959 ;
  assign n12006 = n12001 & n12005 ;
  assign n12022 = ~n7328 & ~n12006 ;
  assign n12023 = ~n12004 & n12022 ;
  assign n12024 = ~n12014 & n12023 ;
  assign n12025 = ~n12021 & n12024 ;
  assign n12026 = \P3_PhyAddrPointer_reg[20]/NET0131  & n2896 ;
  assign n12030 = n4254 & ~n8393 ;
  assign n12031 = ~n3753 & ~n8342 ;
  assign n12032 = ~n12030 & n12031 ;
  assign n12027 = ~n3792 & ~n6093 ;
  assign n12028 = ~n8347 & ~n12027 ;
  assign n12029 = n3753 & ~n12028 ;
  assign n12033 = ~n2896 & ~n12029 ;
  assign n12034 = ~n12032 & n12033 ;
  assign n12035 = ~n12026 & ~n12034 ;
  assign n12036 = n2894 & ~n12035 ;
  assign n12037 = \P3_PhyAddrPointer_reg[20]/NET0131  & ~n9014 ;
  assign n12038 = ~\P3_InstAddrPointer_reg[20]/NET0131  & ~n4364 ;
  assign n12039 = ~n4365 & ~n12038 ;
  assign n12040 = n4360 & n6126 ;
  assign n12041 = n3754 & n12040 ;
  assign n12042 = ~n12039 & ~n12041 ;
  assign n12043 = n2905 & ~n6127 ;
  assign n12044 = ~n12042 & n12043 ;
  assign n12045 = ~n12037 & ~n12044 ;
  assign n12046 = ~n12036 & n12045 ;
  assign n12047 = n2453 & ~n12046 ;
  assign n12048 = n9034 & n9035 ;
  assign n12052 = \P3_PhyAddrPointer_reg[1]/NET0131  & n12048 ;
  assign n12053 = ~\P3_PhyAddrPointer_reg[20]/NET0131  & ~n12052 ;
  assign n12054 = \P3_PhyAddrPointer_reg[1]/NET0131  & n9037 ;
  assign n12055 = ~n12053 & ~n12054 ;
  assign n12056 = n10076 & n12055 ;
  assign n12049 = ~\P3_PhyAddrPointer_reg[20]/NET0131  & ~n12048 ;
  assign n12050 = n2970 & ~n9037 ;
  assign n12051 = ~n12049 & n12050 ;
  assign n12057 = \P3_PhyAddrPointer_reg[20]/NET0131  & ~n9063 ;
  assign n12058 = \P3_rEIP_reg[20]/NET0131  & n4412 ;
  assign n12059 = ~n12057 & ~n12058 ;
  assign n12060 = ~n12051 & n12059 ;
  assign n12061 = ~n12056 & n12060 ;
  assign n12062 = ~n12047 & n12061 ;
  assign n12063 = \P3_PhyAddrPointer_reg[22]/NET0131  & n2896 ;
  assign n12064 = ~n7390 & ~n12063 ;
  assign n12065 = n2894 & ~n12064 ;
  assign n12066 = \P3_PhyAddrPointer_reg[22]/NET0131  & ~n9014 ;
  assign n12067 = ~n7398 & ~n12066 ;
  assign n12068 = ~n12065 & n12067 ;
  assign n12069 = n2453 & ~n12068 ;
  assign n12073 = \P3_PhyAddrPointer_reg[1]/NET0131  & n9038 ;
  assign n12074 = ~\P3_PhyAddrPointer_reg[22]/NET0131  & ~n12073 ;
  assign n12075 = ~n11118 & ~n12074 ;
  assign n12076 = n10076 & n12075 ;
  assign n12070 = ~\P3_PhyAddrPointer_reg[22]/NET0131  & ~n9038 ;
  assign n12071 = n2970 & ~n9039 ;
  assign n12072 = ~n12070 & n12071 ;
  assign n12077 = \P3_PhyAddrPointer_reg[22]/NET0131  & ~n9063 ;
  assign n12078 = ~n7412 & ~n12077 ;
  assign n12079 = ~n12072 & n12078 ;
  assign n12080 = ~n12076 & n12079 ;
  assign n12081 = ~n12069 & n12080 ;
  assign n12089 = n4263 & ~n8395 ;
  assign n12090 = ~n8396 & ~n12089 ;
  assign n12091 = ~n3753 & ~n12090 ;
  assign n12092 = ~n6095 & ~n6097 ;
  assign n12093 = n3753 & ~n6098 ;
  assign n12094 = ~n12092 & n12093 ;
  assign n12095 = ~n12091 & ~n12094 ;
  assign n12096 = ~n2896 & ~n12095 ;
  assign n12097 = n2894 & n12096 ;
  assign n12082 = ~\P3_InstAddrPointer_reg[24]/NET0131  & ~n4375 ;
  assign n12083 = ~n4376 & ~n12082 ;
  assign n12084 = \P3_InstAddrPointer_reg[23]/NET0131  & n7395 ;
  assign n12085 = ~n12083 & ~n12084 ;
  assign n12086 = n2905 & ~n6128 ;
  assign n12087 = ~n12085 & n12086 ;
  assign n12088 = \P3_PhyAddrPointer_reg[24]/NET0131  & ~n11965 ;
  assign n12098 = ~n12087 & ~n12088 ;
  assign n12099 = ~n12097 & n12098 ;
  assign n12100 = n2453 & ~n12099 ;
  assign n12105 = ~\P3_PhyAddrPointer_reg[24]/NET0131  & ~n11121 ;
  assign n12106 = n9040 & n11118 ;
  assign n12107 = ~n12105 & ~n12106 ;
  assign n12108 = n10076 & n12107 ;
  assign n12102 = ~\P3_PhyAddrPointer_reg[24]/NET0131  & ~n11120 ;
  assign n12101 = n9039 & n9040 ;
  assign n12103 = n2970 & ~n12101 ;
  assign n12104 = ~n12102 & n12103 ;
  assign n12109 = \P3_PhyAddrPointer_reg[24]/NET0131  & ~n9063 ;
  assign n12110 = \P3_rEIP_reg[24]/NET0131  & n4412 ;
  assign n12111 = ~n12109 & ~n12110 ;
  assign n12112 = ~n12104 & n12111 ;
  assign n12113 = ~n12108 & n12112 ;
  assign n12114 = ~n12100 & n12113 ;
  assign n12116 = \P3_PhyAddrPointer_reg[26]/NET0131  & n2896 ;
  assign n12121 = ~n4093 & n10049 ;
  assign n12120 = n4093 & ~n10049 ;
  assign n12122 = n3753 & ~n12120 ;
  assign n12123 = ~n12121 & n12122 ;
  assign n12117 = n4277 & ~n10040 ;
  assign n12118 = ~n3753 & ~n10041 ;
  assign n12119 = ~n12117 & n12118 ;
  assign n12124 = ~n2896 & ~n12119 ;
  assign n12125 = ~n12123 & n12124 ;
  assign n12126 = ~n12116 & ~n12125 ;
  assign n12127 = n2894 & ~n12126 ;
  assign n12128 = \P3_PhyAddrPointer_reg[26]/NET0131  & ~n9014 ;
  assign n12129 = ~\P3_InstAddrPointer_reg[26]/NET0131  & ~n4378 ;
  assign n12130 = ~n4381 & ~n12129 ;
  assign n12131 = ~n6129 & ~n12130 ;
  assign n12132 = n2905 & ~n6130 ;
  assign n12133 = ~n12131 & n12132 ;
  assign n12134 = ~n12128 & ~n12133 ;
  assign n12135 = ~n12127 & n12134 ;
  assign n12136 = n2453 & ~n12135 ;
  assign n12142 = n9041 & n11118 ;
  assign n12143 = ~\P3_PhyAddrPointer_reg[26]/NET0131  & ~n12142 ;
  assign n12144 = ~n9044 & ~n12143 ;
  assign n12145 = n10076 & n12144 ;
  assign n12137 = n9039 & n9041 ;
  assign n12138 = ~\P3_PhyAddrPointer_reg[26]/NET0131  & ~n12137 ;
  assign n12139 = n2970 & ~n9043 ;
  assign n12140 = ~n12138 & n12139 ;
  assign n12115 = \P3_PhyAddrPointer_reg[26]/NET0131  & ~n9063 ;
  assign n12141 = \P3_rEIP_reg[26]/NET0131  & n4412 ;
  assign n12146 = ~n12115 & ~n12141 ;
  assign n12147 = ~n12140 & n12146 ;
  assign n12148 = ~n12145 & n12147 ;
  assign n12149 = ~n12136 & n12148 ;
  assign n12162 = \P1_PhyAddrPointer_reg[11]/NET0131  & n2375 ;
  assign n12163 = ~n4780 & n6844 ;
  assign n12164 = ~n6828 & ~n12163 ;
  assign n12165 = n4453 & ~n12164 ;
  assign n12167 = ~n4878 & n6858 ;
  assign n12166 = n4878 & ~n6858 ;
  assign n12168 = ~n4453 & ~n12166 ;
  assign n12169 = ~n12167 & n12168 ;
  assign n12170 = ~n2375 & ~n12169 ;
  assign n12171 = ~n12165 & n12170 ;
  assign n12172 = ~n12162 & ~n12171 ;
  assign n12173 = n2244 & ~n12172 ;
  assign n12159 = n5026 & n6005 ;
  assign n12158 = ~n5026 & ~n6005 ;
  assign n12160 = n2385 & ~n12158 ;
  assign n12161 = ~n12159 & n12160 ;
  assign n12174 = \P1_PhyAddrPointer_reg[11]/NET0131  & ~n10087 ;
  assign n12175 = ~n12161 & ~n12174 ;
  assign n12176 = ~n12173 & n12175 ;
  assign n12177 = n2432 & ~n12176 ;
  assign n12150 = \P1_PhyAddrPointer_reg[1]/NET0131  & n10096 ;
  assign n12151 = \P1_PhyAddrPointer_reg[8]/NET0131  & n12150 ;
  assign n12152 = \P1_PhyAddrPointer_reg[9]/NET0131  & n12151 ;
  assign n12153 = \P1_PhyAddrPointer_reg[10]/NET0131  & n12152 ;
  assign n12154 = ~\P1_PhyAddrPointer_reg[11]/NET0131  & ~n12153 ;
  assign n12155 = \P1_PhyAddrPointer_reg[11]/NET0131  & n12153 ;
  assign n12156 = ~n12154 & ~n12155 ;
  assign n12178 = ~\P1_DataWidth_reg[1]/NET0131  & ~n12156 ;
  assign n12179 = ~\P1_PhyAddrPointer_reg[11]/NET0131  & ~n10099 ;
  assign n12180 = ~n10100 & ~n12179 ;
  assign n12181 = \P1_DataWidth_reg[1]/NET0131  & ~n12180 ;
  assign n12182 = n2436 & ~n12181 ;
  assign n12183 = ~n12178 & n12182 ;
  assign n12157 = n5095 & n12156 ;
  assign n12184 = \P1_rEIP_reg[11]/NET0131  & n5092 ;
  assign n12185 = \P1_PhyAddrPointer_reg[11]/NET0131  & ~n10136 ;
  assign n12186 = ~n12184 & ~n12185 ;
  assign n12187 = ~n12157 & n12186 ;
  assign n12188 = ~n12183 & n12187 ;
  assign n12189 = ~n12177 & n12188 ;
  assign n12197 = \P1_InstAddrPointer_reg[14]/NET0131  & n4465 ;
  assign n12198 = ~\P1_InstAddrPointer_reg[15]/NET0131  & ~n12197 ;
  assign n12199 = ~n4782 & ~n12198 ;
  assign n12200 = n4765 & n5970 ;
  assign n12201 = n4788 & n12200 ;
  assign n12202 = \P1_InstAddrPointer_reg[14]/NET0131  & n12201 ;
  assign n12203 = ~n12199 & ~n12202 ;
  assign n12204 = ~n6832 & ~n12203 ;
  assign n12205 = n4453 & ~n12204 ;
  assign n12194 = n4913 & ~n6860 ;
  assign n12195 = ~n4453 & ~n8548 ;
  assign n12196 = ~n12194 & n12195 ;
  assign n12206 = ~n2375 & ~n12196 ;
  assign n12207 = ~n12205 & n12206 ;
  assign n12208 = n2244 & n12207 ;
  assign n12190 = n6005 & n6008 ;
  assign n12191 = ~n6007 & ~n12190 ;
  assign n12192 = n2385 & ~n6010 ;
  assign n12193 = ~n12191 & n12192 ;
  assign n12209 = ~n2376 & n10087 ;
  assign n12210 = \P1_PhyAddrPointer_reg[15]/NET0131  & ~n12209 ;
  assign n12211 = ~n12193 & ~n12210 ;
  assign n12212 = ~n12208 & n12211 ;
  assign n12213 = n2432 & ~n12212 ;
  assign n12217 = \P1_PhyAddrPointer_reg[12]/NET0131  & n12155 ;
  assign n12218 = \P1_PhyAddrPointer_reg[13]/NET0131  & n12217 ;
  assign n12219 = \P1_PhyAddrPointer_reg[14]/NET0131  & n12218 ;
  assign n12220 = ~\P1_PhyAddrPointer_reg[15]/NET0131  & ~n12219 ;
  assign n12221 = \P1_PhyAddrPointer_reg[15]/NET0131  & n12219 ;
  assign n12222 = ~n12220 & ~n12221 ;
  assign n12223 = n10133 & n12222 ;
  assign n12214 = ~\P1_PhyAddrPointer_reg[15]/NET0131  & ~n10103 ;
  assign n12215 = n3148 & ~n10104 ;
  assign n12216 = ~n12214 & n12215 ;
  assign n12224 = \P1_rEIP_reg[15]/NET0131  & n5092 ;
  assign n12225 = \P1_PhyAddrPointer_reg[15]/NET0131  & ~n10136 ;
  assign n12226 = ~n12224 & ~n12225 ;
  assign n12227 = ~n12216 & n12226 ;
  assign n12228 = ~n12223 & n12227 ;
  assign n12229 = ~n12213 & n12228 ;
  assign n12247 = \P1_PhyAddrPointer_reg[19]/NET0131  & n2375 ;
  assign n12252 = ~n6846 & ~n8545 ;
  assign n12253 = ~n6834 & ~n12252 ;
  assign n12254 = n4453 & ~n12253 ;
  assign n12248 = ~n4926 & ~n6861 ;
  assign n12249 = n4926 & n6861 ;
  assign n12250 = ~n12248 & ~n12249 ;
  assign n12251 = ~n4453 & ~n12250 ;
  assign n12255 = ~n2375 & ~n12251 ;
  assign n12256 = ~n12254 & n12255 ;
  assign n12257 = ~n12247 & ~n12256 ;
  assign n12258 = n2244 & ~n12257 ;
  assign n12243 = n4469 & n9352 ;
  assign n12244 = ~n4973 & ~n12243 ;
  assign n12245 = n2385 & ~n6012 ;
  assign n12246 = ~n12244 & n12245 ;
  assign n12259 = \P1_PhyAddrPointer_reg[19]/NET0131  & ~n10087 ;
  assign n12260 = ~n12246 & ~n12259 ;
  assign n12261 = ~n12258 & n12260 ;
  assign n12262 = n2432 & ~n12261 ;
  assign n12237 = \P1_PhyAddrPointer_reg[18]/NET0131  & n10124 ;
  assign n12238 = ~\P1_PhyAddrPointer_reg[19]/NET0131  & ~n12237 ;
  assign n12230 = \P1_PhyAddrPointer_reg[18]/NET0131  & n10106 ;
  assign n12239 = \P1_PhyAddrPointer_reg[19]/NET0131  & n12230 ;
  assign n12240 = \P1_PhyAddrPointer_reg[1]/NET0131  & n12239 ;
  assign n12241 = ~n12238 & ~n12240 ;
  assign n12242 = n10133 & n12241 ;
  assign n12231 = n3148 & ~n12230 ;
  assign n12232 = n10136 & ~n12231 ;
  assign n12233 = \P1_PhyAddrPointer_reg[19]/NET0131  & ~n12232 ;
  assign n12234 = ~\P1_PhyAddrPointer_reg[19]/NET0131  & n3148 ;
  assign n12235 = n12230 & n12234 ;
  assign n12236 = \P1_rEIP_reg[19]/NET0131  & n5092 ;
  assign n12263 = ~n12235 & ~n12236 ;
  assign n12264 = ~n12233 & n12263 ;
  assign n12265 = ~n12242 & n12264 ;
  assign n12266 = ~n12262 & n12265 ;
  assign n12267 = \P1_PhyAddrPointer_reg[20]/NET0131  & n2375 ;
  assign n12268 = ~n7669 & ~n12267 ;
  assign n12269 = n2244 & ~n12268 ;
  assign n12270 = \P1_PhyAddrPointer_reg[20]/NET0131  & ~n10087 ;
  assign n12271 = ~n7675 & ~n12270 ;
  assign n12272 = ~n12269 & n12271 ;
  assign n12273 = n2432 & ~n12272 ;
  assign n12275 = ~\P1_PhyAddrPointer_reg[20]/NET0131  & ~n12240 ;
  assign n12276 = \P1_PhyAddrPointer_reg[20]/NET0131  & n12239 ;
  assign n12277 = \P1_PhyAddrPointer_reg[1]/NET0131  & n12276 ;
  assign n12278 = ~n12275 & ~n12277 ;
  assign n12279 = n10133 & n12278 ;
  assign n12280 = n3148 & ~n12276 ;
  assign n12281 = ~\P1_PhyAddrPointer_reg[20]/NET0131  & ~n12239 ;
  assign n12282 = n12280 & ~n12281 ;
  assign n12274 = \P1_PhyAddrPointer_reg[20]/NET0131  & ~n10136 ;
  assign n12283 = ~n7658 & ~n12274 ;
  assign n12284 = ~n12282 & n12283 ;
  assign n12285 = ~n12279 & n12284 ;
  assign n12286 = ~n12273 & n12285 ;
  assign n12287 = \P1_PhyAddrPointer_reg[22]/NET0131  & n2375 ;
  assign n12289 = n6862 & n8549 ;
  assign n12290 = n4902 & ~n12289 ;
  assign n12288 = n6863 & n8549 ;
  assign n12291 = ~n4453 & ~n12288 ;
  assign n12292 = ~n12290 & n12291 ;
  assign n12294 = n4476 & ~n4795 ;
  assign n12293 = ~n4476 & n4795 ;
  assign n12295 = n4453 & ~n12293 ;
  assign n12296 = ~n12294 & n12295 ;
  assign n12297 = ~n2375 & ~n12296 ;
  assign n12298 = ~n12292 & n12297 ;
  assign n12299 = ~n12287 & ~n12298 ;
  assign n12300 = n2244 & ~n12299 ;
  assign n12301 = \P1_PhyAddrPointer_reg[22]/NET0131  & ~n10087 ;
  assign n12303 = n5040 & n5049 ;
  assign n12302 = ~n5040 & ~n5049 ;
  assign n12304 = n2385 & ~n12302 ;
  assign n12305 = ~n12303 & n12304 ;
  assign n12306 = ~n12301 & ~n12305 ;
  assign n12307 = ~n12300 & n12306 ;
  assign n12308 = n2432 & ~n12307 ;
  assign n12310 = ~\P1_PhyAddrPointer_reg[22]/NET0131  & ~n10125 ;
  assign n12311 = ~n11252 & ~n12310 ;
  assign n12312 = n10133 & n12311 ;
  assign n12313 = ~\P1_PhyAddrPointer_reg[22]/NET0131  & ~n10110 ;
  assign n12314 = n11247 & ~n12313 ;
  assign n12309 = \P1_PhyAddrPointer_reg[22]/NET0131  & ~n10136 ;
  assign n12315 = \P1_rEIP_reg[22]/NET0131  & n5092 ;
  assign n12316 = ~n12309 & ~n12315 ;
  assign n12317 = ~n12314 & n12316 ;
  assign n12318 = ~n12312 & n12317 ;
  assign n12319 = ~n12308 & n12318 ;
  assign n12320 = \P1_PhyAddrPointer_reg[24]/NET0131  & n2375 ;
  assign n12321 = ~n7293 & ~n12320 ;
  assign n12322 = n2244 & ~n12321 ;
  assign n12323 = \P1_PhyAddrPointer_reg[24]/NET0131  & ~n10087 ;
  assign n12324 = ~n7307 & ~n12323 ;
  assign n12325 = ~n12322 & n12324 ;
  assign n12326 = n2432 & ~n12325 ;
  assign n12332 = ~\P1_PhyAddrPointer_reg[24]/NET0131  & ~n11254 ;
  assign n12327 = \P1_PhyAddrPointer_reg[23]/NET0131  & n11246 ;
  assign n12328 = \P1_PhyAddrPointer_reg[24]/NET0131  & n12327 ;
  assign n12333 = \P1_PhyAddrPointer_reg[1]/NET0131  & n12328 ;
  assign n12334 = ~n12332 & ~n12333 ;
  assign n12335 = n10133 & n12334 ;
  assign n12329 = ~\P1_PhyAddrPointer_reg[24]/NET0131  & ~n12327 ;
  assign n12330 = n3148 & ~n12328 ;
  assign n12331 = ~n12329 & n12330 ;
  assign n12336 = \P1_PhyAddrPointer_reg[24]/NET0131  & ~n10136 ;
  assign n12337 = ~n7268 & ~n12336 ;
  assign n12338 = ~n12331 & n12337 ;
  assign n12339 = ~n12335 & n12338 ;
  assign n12340 = ~n12326 & n12339 ;
  assign n12341 = \P1_PhyAddrPointer_reg[26]/NET0131  & n2375 ;
  assign n12342 = ~n7243 & ~n12341 ;
  assign n12343 = n2244 & ~n12342 ;
  assign n12344 = \P1_PhyAddrPointer_reg[26]/NET0131  & ~n10087 ;
  assign n12345 = ~n7254 & ~n12344 ;
  assign n12346 = ~n12343 & n12345 ;
  assign n12347 = n2432 & ~n12346 ;
  assign n12353 = ~\P1_PhyAddrPointer_reg[26]/NET0131  & ~n10126 ;
  assign n12354 = ~n10127 & ~n12353 ;
  assign n12355 = n10133 & n12354 ;
  assign n12350 = n3148 & ~n10114 ;
  assign n12351 = n10136 & ~n12350 ;
  assign n12352 = \P1_PhyAddrPointer_reg[26]/NET0131  & ~n12351 ;
  assign n12348 = ~\P1_PhyAddrPointer_reg[26]/NET0131  & n3148 ;
  assign n12349 = n10114 & n12348 ;
  assign n12356 = ~n7226 & ~n12349 ;
  assign n12357 = ~n12352 & n12356 ;
  assign n12358 = ~n12355 & n12357 ;
  assign n12359 = ~n12347 & n12358 ;
  assign n12360 = \P2_PhyAddrPointer_reg[11]/NET0131  & n1897 ;
  assign n12361 = ~n8448 & ~n12360 ;
  assign n12362 = n1734 & ~n12361 ;
  assign n12363 = \P2_PhyAddrPointer_reg[11]/NET0131  & ~n8936 ;
  assign n12364 = ~n8454 & ~n12363 ;
  assign n12365 = ~n12362 & n12364 ;
  assign n12366 = n1927 & ~n12365 ;
  assign n12373 = \P2_PhyAddrPointer_reg[1]/NET0131  & n8966 ;
  assign n12374 = \P2_PhyAddrPointer_reg[10]/NET0131  & n12373 ;
  assign n12375 = ~\P2_PhyAddrPointer_reg[11]/NET0131  & ~n12374 ;
  assign n12376 = n8967 & n12373 ;
  assign n12377 = ~n12375 & ~n12376 ;
  assign n12378 = n3087 & n12377 ;
  assign n12367 = \P2_PhyAddrPointer_reg[10]/NET0131  & n8966 ;
  assign n12368 = ~n10965 & n12367 ;
  assign n12369 = ~\P2_PhyAddrPointer_reg[11]/NET0131  & ~n12368 ;
  assign n12370 = n8968 & ~n10965 ;
  assign n12371 = n1931 & ~n12370 ;
  assign n12372 = ~n12369 & n12371 ;
  assign n12379 = \P2_PhyAddrPointer_reg[11]/NET0131  & ~n8958 ;
  assign n12380 = ~n8434 & ~n12379 ;
  assign n12381 = ~n12372 & n12380 ;
  assign n12382 = ~n12378 & n12381 ;
  assign n12383 = ~n12366 & n12382 ;
  assign n12397 = n1734 & n7478 ;
  assign n12395 = ~n1901 & n8936 ;
  assign n12396 = \P2_PhyAddrPointer_reg[15]/NET0131  & ~n12395 ;
  assign n12398 = ~n7498 & ~n12396 ;
  assign n12399 = ~n12397 & n12398 ;
  assign n12400 = n1927 & ~n12399 ;
  assign n12390 = n8971 & ~n10965 ;
  assign n12391 = ~\P2_PhyAddrPointer_reg[15]/NET0131  & ~n12390 ;
  assign n12389 = n8972 & ~n10965 ;
  assign n12392 = n1931 & ~n12389 ;
  assign n12393 = ~n12391 & n12392 ;
  assign n12384 = \P2_PhyAddrPointer_reg[1]/NET0131  & n8971 ;
  assign n12385 = ~\P2_PhyAddrPointer_reg[15]/NET0131  & ~n12384 ;
  assign n12386 = \P2_PhyAddrPointer_reg[1]/NET0131  & n8972 ;
  assign n12387 = ~n12385 & ~n12386 ;
  assign n12388 = n3087 & n12387 ;
  assign n12394 = \P2_PhyAddrPointer_reg[15]/NET0131  & ~n8958 ;
  assign n12401 = ~n7416 & ~n12394 ;
  assign n12402 = ~n12388 & n12401 ;
  assign n12403 = ~n12393 & n12402 ;
  assign n12404 = ~n12400 & n12403 ;
  assign n12405 = \P2_PhyAddrPointer_reg[19]/NET0131  & n1897 ;
  assign n12409 = n6539 & ~n8914 ;
  assign n12410 = ~n6188 & ~n10939 ;
  assign n12411 = ~n12409 & n12410 ;
  assign n12406 = ~n7592 & ~n7594 ;
  assign n12407 = ~n7525 & ~n12406 ;
  assign n12408 = n6188 & ~n12407 ;
  assign n12412 = ~n1897 & ~n12408 ;
  assign n12413 = ~n12411 & n12412 ;
  assign n12414 = ~n12405 & ~n12413 ;
  assign n12415 = n1734 & ~n12414 ;
  assign n12416 = \P2_PhyAddrPointer_reg[19]/NET0131  & ~n8936 ;
  assign n12418 = n7552 & n8941 ;
  assign n12417 = ~n7552 & ~n8941 ;
  assign n12419 = n1890 & ~n12417 ;
  assign n12420 = ~n12418 & n12419 ;
  assign n12421 = ~n12416 & ~n12420 ;
  assign n12422 = ~n12415 & n12421 ;
  assign n12423 = n1927 & ~n12422 ;
  assign n12427 = \P2_PhyAddrPointer_reg[1]/NET0131  & n8975 ;
  assign n12428 = ~\P2_PhyAddrPointer_reg[19]/NET0131  & ~n12427 ;
  assign n12429 = ~n11874 & ~n12428 ;
  assign n12430 = n9005 & n12429 ;
  assign n12424 = ~\P2_PhyAddrPointer_reg[19]/NET0131  & ~n8975 ;
  assign n12425 = n3034 & ~n8976 ;
  assign n12426 = ~n12424 & n12425 ;
  assign n12431 = \P2_rEIP_reg[19]/NET0131  & n3113 ;
  assign n12432 = \P2_PhyAddrPointer_reg[19]/NET0131  & ~n8958 ;
  assign n12433 = ~n12431 & ~n12432 ;
  assign n12434 = ~n12426 & n12433 ;
  assign n12435 = ~n12430 & n12434 ;
  assign n12436 = ~n12423 & n12435 ;
  assign n12445 = ~n5001 & n5995 ;
  assign n12442 = ~n4993 & ~n5001 ;
  assign n12443 = ~n4994 & ~n5994 ;
  assign n12444 = ~n12442 & ~n12443 ;
  assign n12446 = n2385 & ~n12444 ;
  assign n12447 = ~n12445 & n12446 ;
  assign n12454 = ~n4642 & ~n4752 ;
  assign n12455 = n4748 & ~n12454 ;
  assign n12456 = ~n4748 & n12454 ;
  assign n12457 = ~n12455 & ~n12456 ;
  assign n12458 = n4453 & ~n12457 ;
  assign n12448 = ~n4850 & ~n5946 ;
  assign n12449 = ~n4847 & ~n4853 ;
  assign n12451 = n12448 & ~n12449 ;
  assign n12450 = ~n12448 & n12449 ;
  assign n12452 = ~n4453 & ~n12450 ;
  assign n12453 = ~n12451 & n12452 ;
  assign n12459 = n2384 & ~n12453 ;
  assign n12460 = ~n12458 & n12459 ;
  assign n12461 = ~n12447 & ~n12460 ;
  assign n12439 = \P1_InstAddrPointer_reg[3]/NET0131  & ~n11428 ;
  assign n12462 = ~n2402 & n4641 ;
  assign n12440 = ~n2271 & n4846 ;
  assign n12441 = n2397 & n4992 ;
  assign n12463 = ~n12440 & ~n12441 ;
  assign n12464 = ~n12462 & n12463 ;
  assign n12465 = ~n12439 & n12464 ;
  assign n12466 = n12461 & n12465 ;
  assign n12467 = n2432 & ~n12466 ;
  assign n12437 = \P1_rEIP_reg[3]/NET0131  & n5092 ;
  assign n12438 = \P1_InstAddrPointer_reg[3]/NET0131  & ~n5098 ;
  assign n12468 = ~n12437 & ~n12438 ;
  assign n12469 = ~n12467 & n12468 ;
  assign n12473 = \P1_InstAddrPointer_reg[5]/NET0131  & n2375 ;
  assign n12474 = ~n4574 & ~n4760 ;
  assign n12475 = ~n4755 & ~n12474 ;
  assign n12476 = n4755 & n12474 ;
  assign n12477 = ~n12475 & ~n12476 ;
  assign n12478 = ~n2375 & ~n12477 ;
  assign n12479 = ~n12473 & ~n12478 ;
  assign n12480 = n2244 & ~n12479 ;
  assign n12472 = \P1_InstAddrPointer_reg[5]/NET0131  & ~n11427 ;
  assign n12481 = ~n2271 & n4829 ;
  assign n12482 = n2397 & n4985 ;
  assign n12490 = ~n12481 & ~n12482 ;
  assign n12491 = ~n12472 & n12490 ;
  assign n12483 = ~n2402 & n4542 ;
  assign n12487 = ~n5007 & n5998 ;
  assign n12484 = ~n4986 & ~n5007 ;
  assign n12485 = ~n4989 & ~n5997 ;
  assign n12486 = ~n12484 & ~n12485 ;
  assign n12488 = n2385 & ~n12486 ;
  assign n12489 = ~n12487 & n12488 ;
  assign n12492 = ~n12483 & ~n12489 ;
  assign n12493 = n12491 & n12492 ;
  assign n12494 = ~n12480 & n12493 ;
  assign n12495 = n2432 & ~n12494 ;
  assign n12470 = \P1_rEIP_reg[5]/NET0131  & n5092 ;
  assign n12471 = \P1_InstAddrPointer_reg[5]/NET0131  & ~n5098 ;
  assign n12496 = ~n12470 & ~n12471 ;
  assign n12497 = ~n12495 & n12496 ;
  assign n12515 = ~n4198 & ~n4206 ;
  assign n12516 = ~n4193 & ~n4194 ;
  assign n12517 = ~n12515 & ~n12516 ;
  assign n12518 = n12515 & n12516 ;
  assign n12519 = ~n12517 & ~n12518 ;
  assign n12520 = ~n3753 & ~n12519 ;
  assign n12521 = ~n3967 & ~n4036 ;
  assign n12522 = ~n4035 & ~n4041 ;
  assign n12524 = ~n12521 & n12522 ;
  assign n12523 = n12521 & ~n12522 ;
  assign n12525 = n3753 & ~n12523 ;
  assign n12526 = ~n12524 & n12525 ;
  assign n12527 = ~n12520 & ~n12526 ;
  assign n12528 = ~n2896 & ~n12527 ;
  assign n12514 = ~\P3_InstAddrPointer_reg[3]/NET0131  & n2896 ;
  assign n12529 = n2894 & ~n12514 ;
  assign n12530 = ~n12528 & n12529 ;
  assign n12513 = ~n2923 & n4034 ;
  assign n12500 = ~n2777 & n4197 ;
  assign n12505 = n2891 & ~n2900 ;
  assign n12506 = \P3_InstAddrPointer_reg[3]/NET0131  & ~n12505 ;
  assign n12501 = n2847 & ~n4332 ;
  assign n12502 = ~\P3_InstAddrPointer_reg[3]/NET0131  & ~n2847 ;
  assign n12503 = ~n12501 & ~n12502 ;
  assign n12504 = ~n2841 & n12503 ;
  assign n12510 = n4335 & ~n4336 ;
  assign n12507 = ~n4333 & ~n4336 ;
  assign n12508 = ~n4329 & ~n4330 ;
  assign n12509 = ~n12507 & ~n12508 ;
  assign n12511 = n2905 & ~n12509 ;
  assign n12512 = ~n12510 & n12511 ;
  assign n12531 = ~n12504 & ~n12512 ;
  assign n12532 = ~n12506 & n12531 ;
  assign n12533 = ~n12500 & n12532 ;
  assign n12534 = ~n12513 & n12533 ;
  assign n12535 = ~n12530 & n12534 ;
  assign n12536 = n2453 & ~n12535 ;
  assign n12498 = \P3_rEIP_reg[3]/NET0131  & n4412 ;
  assign n12499 = \P3_InstAddrPointer_reg[3]/NET0131  & ~n4418 ;
  assign n12537 = ~n12498 & ~n12499 ;
  assign n12538 = ~n12536 & n12537 ;
  assign n12547 = \P3_InstAddrPointer_reg[5]/NET0131  & ~n11451 ;
  assign n12548 = ~n2923 & n3799 ;
  assign n12541 = ~n3831 & ~n4051 ;
  assign n12542 = n4044 & n12541 ;
  assign n12543 = ~n4044 & ~n12541 ;
  assign n12544 = ~n12542 & ~n12543 ;
  assign n12545 = n2904 & ~n12544 ;
  assign n12546 = n2918 & n4318 ;
  assign n12556 = ~n12545 & ~n12546 ;
  assign n12557 = ~n12548 & n12556 ;
  assign n12549 = ~n2777 & n4184 ;
  assign n12553 = n4340 & ~n4342 ;
  assign n12550 = ~n4319 & ~n4342 ;
  assign n12551 = ~n4316 & ~n4339 ;
  assign n12552 = ~n12550 & ~n12551 ;
  assign n12554 = n2905 & ~n12552 ;
  assign n12555 = ~n12553 & n12554 ;
  assign n12558 = ~n12549 & ~n12555 ;
  assign n12559 = n12557 & n12558 ;
  assign n12560 = ~n12547 & n12559 ;
  assign n12561 = n2453 & ~n12560 ;
  assign n12539 = \P3_rEIP_reg[5]/NET0131  & n4412 ;
  assign n12540 = \P3_InstAddrPointer_reg[5]/NET0131  & ~n4418 ;
  assign n12562 = ~n12539 & ~n12540 ;
  assign n12563 = ~n12561 & n12562 ;
  assign n12585 = ~n1771 & n6439 ;
  assign n12584 = ~n1831 & n6622 ;
  assign n12565 = n1870 & n6709 ;
  assign n12586 = ~n6710 & ~n6722 ;
  assign n12588 = ~n6719 & ~n12586 ;
  assign n12587 = n6719 & n12586 ;
  assign n12589 = n1890 & ~n12587 ;
  assign n12590 = ~n12588 & n12589 ;
  assign n12591 = ~n12565 & ~n12590 ;
  assign n12592 = ~n12584 & n12591 ;
  assign n12593 = ~n12585 & n12592 ;
  assign n12566 = n1824 & n1903 ;
  assign n12567 = ~n1901 & n12566 ;
  assign n12568 = \P2_InstAddrPointer_reg[3]/NET0131  & ~n12567 ;
  assign n12575 = ~n6623 & ~n6629 ;
  assign n12576 = ~n6617 & ~n6624 ;
  assign n12577 = ~n12575 & ~n12576 ;
  assign n12578 = n12575 & n12576 ;
  assign n12579 = ~n12577 & ~n12578 ;
  assign n12580 = n6188 & ~n12579 ;
  assign n12569 = ~n6372 & ~n6441 ;
  assign n12570 = ~n6440 & ~n6446 ;
  assign n12572 = n12569 & ~n12570 ;
  assign n12571 = ~n12569 & n12570 ;
  assign n12573 = ~n6188 & ~n12571 ;
  assign n12574 = ~n12572 & n12573 ;
  assign n12581 = ~n1897 & ~n12574 ;
  assign n12582 = ~n12580 & n12581 ;
  assign n12583 = n1734 & n12582 ;
  assign n12594 = ~n12568 & ~n12583 ;
  assign n12595 = n12593 & n12594 ;
  assign n12596 = n1927 & ~n12595 ;
  assign n12564 = \P2_rEIP_reg[3]/NET0131  & n3113 ;
  assign n12597 = \P2_InstAddrPointer_reg[3]/NET0131  & ~n6810 ;
  assign n12598 = ~n12564 & ~n12597 ;
  assign n12599 = ~n12596 & n12598 ;
  assign n12605 = ~n6703 & ~n6728 ;
  assign n12607 = ~n6725 & n12605 ;
  assign n12606 = n6725 & ~n12605 ;
  assign n12608 = n1890 & ~n12606 ;
  assign n12609 = ~n12607 & n12608 ;
  assign n12603 = ~n1831 & n6608 ;
  assign n12604 = \P2_InstAddrPointer_reg[5]/NET0131  & ~n10241 ;
  assign n12623 = ~n12603 & ~n12604 ;
  assign n12624 = ~n12609 & n12623 ;
  assign n12610 = \P2_InstAddrPointer_reg[5]/NET0131  & n1897 ;
  assign n12611 = ~n6609 & ~n6637 ;
  assign n12612 = ~n6632 & ~n12611 ;
  assign n12613 = n6632 & n12611 ;
  assign n12614 = ~n12612 & ~n12613 ;
  assign n12615 = ~n1897 & ~n12614 ;
  assign n12616 = ~n12610 & ~n12615 ;
  assign n12617 = n1734 & ~n12616 ;
  assign n12602 = ~n1771 & n6234 ;
  assign n12618 = ~\P2_InstAddrPointer_reg[5]/NET0131  & ~n1798 ;
  assign n12619 = n1798 & ~n6702 ;
  assign n12620 = ~n12618 & ~n12619 ;
  assign n12621 = ~n1727 & n12620 ;
  assign n12622 = ~n12602 & ~n12621 ;
  assign n12625 = ~n12617 & n12622 ;
  assign n12626 = n12624 & n12625 ;
  assign n12627 = n1927 & ~n12626 ;
  assign n12600 = \P2_rEIP_reg[5]/NET0131  & n3113 ;
  assign n12601 = \P2_InstAddrPointer_reg[5]/NET0131  & ~n6810 ;
  assign n12628 = ~n12600 & ~n12601 ;
  assign n12629 = ~n12627 & n12628 ;
  assign n12630 = ~n2980 & ~n2986 ;
  assign n12631 = ~n1933 & n12630 ;
  assign n12632 = ~n1935 & n12631 ;
  assign n12633 = \P2_EAX_reg[31]/NET0131  & ~n12632 ;
  assign n12634 = \P2_EAX_reg[0]/NET0131  & \P2_EAX_reg[1]/NET0131  ;
  assign n12635 = \P2_EAX_reg[2]/NET0131  & n12634 ;
  assign n12636 = \P2_EAX_reg[3]/NET0131  & n12635 ;
  assign n12637 = \P2_EAX_reg[4]/NET0131  & n12636 ;
  assign n12638 = \P2_EAX_reg[5]/NET0131  & n12637 ;
  assign n12639 = \P2_EAX_reg[6]/NET0131  & n12638 ;
  assign n12640 = \P2_EAX_reg[7]/NET0131  & n12639 ;
  assign n12641 = \P2_EAX_reg[8]/NET0131  & n12640 ;
  assign n12642 = \P2_EAX_reg[9]/NET0131  & n12641 ;
  assign n12643 = \P2_EAX_reg[10]/NET0131  & n12642 ;
  assign n12644 = \P2_EAX_reg[11]/NET0131  & n12643 ;
  assign n12645 = \P2_EAX_reg[12]/NET0131  & n12644 ;
  assign n12646 = \P2_EAX_reg[13]/NET0131  & n12645 ;
  assign n12647 = \P2_EAX_reg[14]/NET0131  & n12646 ;
  assign n12648 = \P2_EAX_reg[15]/NET0131  & n12647 ;
  assign n12649 = \P2_EAX_reg[16]/NET0131  & n12648 ;
  assign n12650 = \P2_EAX_reg[17]/NET0131  & \P2_EAX_reg[18]/NET0131  ;
  assign n12651 = n12649 & n12650 ;
  assign n12652 = \P2_EAX_reg[19]/NET0131  & n12651 ;
  assign n12653 = \P2_EAX_reg[20]/NET0131  & n12652 ;
  assign n12654 = \P2_EAX_reg[21]/NET0131  & \P2_EAX_reg[22]/NET0131  ;
  assign n12655 = n12653 & n12654 ;
  assign n12656 = \P2_EAX_reg[23]/NET0131  & \P2_EAX_reg[24]/NET0131  ;
  assign n12657 = \P2_EAX_reg[25]/NET0131  & n12656 ;
  assign n12658 = n12655 & n12657 ;
  assign n12659 = \P2_EAX_reg[26]/NET0131  & \P2_EAX_reg[27]/NET0131  ;
  assign n12660 = \P2_EAX_reg[28]/NET0131  & n12659 ;
  assign n12661 = n12658 & n12660 ;
  assign n12662 = \P2_EAX_reg[29]/NET0131  & n12661 ;
  assign n12663 = \P2_EAX_reg[30]/NET0131  & n12662 ;
  assign n12664 = n1737 & n1755 ;
  assign n12665 = ~n12663 & n12664 ;
  assign n12666 = ~n1726 & ~n12664 ;
  assign n12667 = n1804 & n12666 ;
  assign n12668 = ~n1876 & ~n12667 ;
  assign n12669 = ~n1812 & n12668 ;
  assign n12670 = ~n12665 & n12669 ;
  assign n12671 = \P2_EAX_reg[31]/NET0131  & ~n12670 ;
  assign n12672 = ~\P2_EAX_reg[31]/NET0131  & n12664 ;
  assign n12673 = n12663 & n12672 ;
  assign n12678 = \P2_InstQueue_reg[3][7]/NET0131  & n1464 ;
  assign n12679 = \P2_InstQueue_reg[0][7]/NET0131  & n1482 ;
  assign n12692 = ~n12678 & ~n12679 ;
  assign n12680 = \P2_InstQueue_reg[7][7]/NET0131  & n1474 ;
  assign n12681 = \P2_InstQueue_reg[4][7]/NET0131  & n1468 ;
  assign n12693 = ~n12680 & ~n12681 ;
  assign n12700 = n12692 & n12693 ;
  assign n12674 = \P2_InstQueue_reg[13][7]/NET0131  & n1459 ;
  assign n12675 = \P2_InstQueue_reg[9][7]/NET0131  & n1476 ;
  assign n12690 = ~n12674 & ~n12675 ;
  assign n12676 = \P2_InstQueue_reg[2][7]/NET0131  & n1456 ;
  assign n12677 = \P2_InstQueue_reg[15][7]/NET0131  & n1466 ;
  assign n12691 = ~n12676 & ~n12677 ;
  assign n12701 = n12690 & n12691 ;
  assign n12702 = n12700 & n12701 ;
  assign n12686 = \P2_InstQueue_reg[8][7]/NET0131  & n1447 ;
  assign n12687 = \P2_InstQueue_reg[6][7]/NET0131  & n1450 ;
  assign n12696 = ~n12686 & ~n12687 ;
  assign n12688 = \P2_InstQueue_reg[12][7]/NET0131  & n1453 ;
  assign n12689 = \P2_InstQueue_reg[14][7]/NET0131  & n1480 ;
  assign n12697 = ~n12688 & ~n12689 ;
  assign n12698 = n12696 & n12697 ;
  assign n12682 = \P2_InstQueue_reg[1][7]/NET0131  & n1478 ;
  assign n12683 = \P2_InstQueue_reg[11][7]/NET0131  & n1472 ;
  assign n12694 = ~n12682 & ~n12683 ;
  assign n12684 = \P2_InstQueue_reg[5][7]/NET0131  & n1470 ;
  assign n12685 = \P2_InstQueue_reg[10][7]/NET0131  & n1461 ;
  assign n12695 = ~n12684 & ~n12685 ;
  assign n12699 = n12694 & n12695 ;
  assign n12703 = n12698 & n12699 ;
  assign n12704 = n12702 & n12703 ;
  assign n12709 = \P2_InstQueue_reg[2][0]/NET0131  & n1478 ;
  assign n12710 = \P2_InstQueue_reg[0][0]/NET0131  & n1466 ;
  assign n12723 = ~n12709 & ~n12710 ;
  assign n12711 = \P2_InstQueue_reg[15][0]/NET0131  & n1480 ;
  assign n12712 = \P2_InstQueue_reg[14][0]/NET0131  & n1459 ;
  assign n12724 = ~n12711 & ~n12712 ;
  assign n12731 = n12723 & n12724 ;
  assign n12705 = \P2_InstQueue_reg[4][0]/NET0131  & n1464 ;
  assign n12706 = \P2_InstQueue_reg[10][0]/NET0131  & n1476 ;
  assign n12721 = ~n12705 & ~n12706 ;
  assign n12707 = \P2_InstQueue_reg[3][0]/NET0131  & n1456 ;
  assign n12708 = \P2_InstQueue_reg[6][0]/NET0131  & n1470 ;
  assign n12722 = ~n12707 & ~n12708 ;
  assign n12732 = n12721 & n12722 ;
  assign n12733 = n12731 & n12732 ;
  assign n12717 = \P2_InstQueue_reg[1][0]/NET0131  & n1482 ;
  assign n12718 = \P2_InstQueue_reg[7][0]/NET0131  & n1450 ;
  assign n12727 = ~n12717 & ~n12718 ;
  assign n12719 = \P2_InstQueue_reg[12][0]/NET0131  & n1472 ;
  assign n12720 = \P2_InstQueue_reg[8][0]/NET0131  & n1474 ;
  assign n12728 = ~n12719 & ~n12720 ;
  assign n12729 = n12727 & n12728 ;
  assign n12713 = \P2_InstQueue_reg[9][0]/NET0131  & n1447 ;
  assign n12714 = \P2_InstQueue_reg[13][0]/NET0131  & n1453 ;
  assign n12725 = ~n12713 & ~n12714 ;
  assign n12715 = \P2_InstQueue_reg[5][0]/NET0131  & n1468 ;
  assign n12716 = \P2_InstQueue_reg[11][0]/NET0131  & n1461 ;
  assign n12726 = ~n12715 & ~n12716 ;
  assign n12730 = n12725 & n12726 ;
  assign n12734 = n12729 & n12730 ;
  assign n12735 = n12733 & n12734 ;
  assign n12736 = ~n12704 & ~n12735 ;
  assign n12741 = \P2_InstQueue_reg[2][1]/NET0131  & n1478 ;
  assign n12742 = \P2_InstQueue_reg[0][1]/NET0131  & n1466 ;
  assign n12755 = ~n12741 & ~n12742 ;
  assign n12743 = \P2_InstQueue_reg[15][1]/NET0131  & n1480 ;
  assign n12744 = \P2_InstQueue_reg[14][1]/NET0131  & n1459 ;
  assign n12756 = ~n12743 & ~n12744 ;
  assign n12763 = n12755 & n12756 ;
  assign n12737 = \P2_InstQueue_reg[4][1]/NET0131  & n1464 ;
  assign n12738 = \P2_InstQueue_reg[10][1]/NET0131  & n1476 ;
  assign n12753 = ~n12737 & ~n12738 ;
  assign n12739 = \P2_InstQueue_reg[3][1]/NET0131  & n1456 ;
  assign n12740 = \P2_InstQueue_reg[6][1]/NET0131  & n1470 ;
  assign n12754 = ~n12739 & ~n12740 ;
  assign n12764 = n12753 & n12754 ;
  assign n12765 = n12763 & n12764 ;
  assign n12749 = \P2_InstQueue_reg[1][1]/NET0131  & n1482 ;
  assign n12750 = \P2_InstQueue_reg[7][1]/NET0131  & n1450 ;
  assign n12759 = ~n12749 & ~n12750 ;
  assign n12751 = \P2_InstQueue_reg[12][1]/NET0131  & n1472 ;
  assign n12752 = \P2_InstQueue_reg[8][1]/NET0131  & n1474 ;
  assign n12760 = ~n12751 & ~n12752 ;
  assign n12761 = n12759 & n12760 ;
  assign n12745 = \P2_InstQueue_reg[9][1]/NET0131  & n1447 ;
  assign n12746 = \P2_InstQueue_reg[13][1]/NET0131  & n1453 ;
  assign n12757 = ~n12745 & ~n12746 ;
  assign n12747 = \P2_InstQueue_reg[5][1]/NET0131  & n1468 ;
  assign n12748 = \P2_InstQueue_reg[11][1]/NET0131  & n1461 ;
  assign n12758 = ~n12747 & ~n12748 ;
  assign n12762 = n12757 & n12758 ;
  assign n12766 = n12761 & n12762 ;
  assign n12767 = n12765 & n12766 ;
  assign n12768 = n12736 & ~n12767 ;
  assign n12773 = \P2_InstQueue_reg[2][2]/NET0131  & n1478 ;
  assign n12774 = \P2_InstQueue_reg[0][2]/NET0131  & n1466 ;
  assign n12787 = ~n12773 & ~n12774 ;
  assign n12775 = \P2_InstQueue_reg[15][2]/NET0131  & n1480 ;
  assign n12776 = \P2_InstQueue_reg[14][2]/NET0131  & n1459 ;
  assign n12788 = ~n12775 & ~n12776 ;
  assign n12795 = n12787 & n12788 ;
  assign n12769 = \P2_InstQueue_reg[4][2]/NET0131  & n1464 ;
  assign n12770 = \P2_InstQueue_reg[10][2]/NET0131  & n1476 ;
  assign n12785 = ~n12769 & ~n12770 ;
  assign n12771 = \P2_InstQueue_reg[3][2]/NET0131  & n1456 ;
  assign n12772 = \P2_InstQueue_reg[6][2]/NET0131  & n1470 ;
  assign n12786 = ~n12771 & ~n12772 ;
  assign n12796 = n12785 & n12786 ;
  assign n12797 = n12795 & n12796 ;
  assign n12781 = \P2_InstQueue_reg[1][2]/NET0131  & n1482 ;
  assign n12782 = \P2_InstQueue_reg[7][2]/NET0131  & n1450 ;
  assign n12791 = ~n12781 & ~n12782 ;
  assign n12783 = \P2_InstQueue_reg[12][2]/NET0131  & n1472 ;
  assign n12784 = \P2_InstQueue_reg[8][2]/NET0131  & n1474 ;
  assign n12792 = ~n12783 & ~n12784 ;
  assign n12793 = n12791 & n12792 ;
  assign n12777 = \P2_InstQueue_reg[9][2]/NET0131  & n1447 ;
  assign n12778 = \P2_InstQueue_reg[13][2]/NET0131  & n1453 ;
  assign n12789 = ~n12777 & ~n12778 ;
  assign n12779 = \P2_InstQueue_reg[5][2]/NET0131  & n1468 ;
  assign n12780 = \P2_InstQueue_reg[11][2]/NET0131  & n1461 ;
  assign n12790 = ~n12779 & ~n12780 ;
  assign n12794 = n12789 & n12790 ;
  assign n12798 = n12793 & n12794 ;
  assign n12799 = n12797 & n12798 ;
  assign n12800 = n12768 & ~n12799 ;
  assign n12805 = \P2_InstQueue_reg[2][3]/NET0131  & n1478 ;
  assign n12806 = \P2_InstQueue_reg[0][3]/NET0131  & n1466 ;
  assign n12819 = ~n12805 & ~n12806 ;
  assign n12807 = \P2_InstQueue_reg[15][3]/NET0131  & n1480 ;
  assign n12808 = \P2_InstQueue_reg[14][3]/NET0131  & n1459 ;
  assign n12820 = ~n12807 & ~n12808 ;
  assign n12827 = n12819 & n12820 ;
  assign n12801 = \P2_InstQueue_reg[4][3]/NET0131  & n1464 ;
  assign n12802 = \P2_InstQueue_reg[10][3]/NET0131  & n1476 ;
  assign n12817 = ~n12801 & ~n12802 ;
  assign n12803 = \P2_InstQueue_reg[3][3]/NET0131  & n1456 ;
  assign n12804 = \P2_InstQueue_reg[6][3]/NET0131  & n1470 ;
  assign n12818 = ~n12803 & ~n12804 ;
  assign n12828 = n12817 & n12818 ;
  assign n12829 = n12827 & n12828 ;
  assign n12813 = \P2_InstQueue_reg[1][3]/NET0131  & n1482 ;
  assign n12814 = \P2_InstQueue_reg[7][3]/NET0131  & n1450 ;
  assign n12823 = ~n12813 & ~n12814 ;
  assign n12815 = \P2_InstQueue_reg[12][3]/NET0131  & n1472 ;
  assign n12816 = \P2_InstQueue_reg[8][3]/NET0131  & n1474 ;
  assign n12824 = ~n12815 & ~n12816 ;
  assign n12825 = n12823 & n12824 ;
  assign n12809 = \P2_InstQueue_reg[9][3]/NET0131  & n1447 ;
  assign n12810 = \P2_InstQueue_reg[13][3]/NET0131  & n1453 ;
  assign n12821 = ~n12809 & ~n12810 ;
  assign n12811 = \P2_InstQueue_reg[5][3]/NET0131  & n1468 ;
  assign n12812 = \P2_InstQueue_reg[11][3]/NET0131  & n1461 ;
  assign n12822 = ~n12811 & ~n12812 ;
  assign n12826 = n12821 & n12822 ;
  assign n12830 = n12825 & n12826 ;
  assign n12831 = n12829 & n12830 ;
  assign n12832 = n12800 & ~n12831 ;
  assign n12837 = \P2_InstQueue_reg[2][4]/NET0131  & n1478 ;
  assign n12838 = \P2_InstQueue_reg[0][4]/NET0131  & n1466 ;
  assign n12851 = ~n12837 & ~n12838 ;
  assign n12839 = \P2_InstQueue_reg[15][4]/NET0131  & n1480 ;
  assign n12840 = \P2_InstQueue_reg[14][4]/NET0131  & n1459 ;
  assign n12852 = ~n12839 & ~n12840 ;
  assign n12859 = n12851 & n12852 ;
  assign n12833 = \P2_InstQueue_reg[4][4]/NET0131  & n1464 ;
  assign n12834 = \P2_InstQueue_reg[10][4]/NET0131  & n1476 ;
  assign n12849 = ~n12833 & ~n12834 ;
  assign n12835 = \P2_InstQueue_reg[3][4]/NET0131  & n1456 ;
  assign n12836 = \P2_InstQueue_reg[6][4]/NET0131  & n1470 ;
  assign n12850 = ~n12835 & ~n12836 ;
  assign n12860 = n12849 & n12850 ;
  assign n12861 = n12859 & n12860 ;
  assign n12845 = \P2_InstQueue_reg[1][4]/NET0131  & n1482 ;
  assign n12846 = \P2_InstQueue_reg[7][4]/NET0131  & n1450 ;
  assign n12855 = ~n12845 & ~n12846 ;
  assign n12847 = \P2_InstQueue_reg[12][4]/NET0131  & n1472 ;
  assign n12848 = \P2_InstQueue_reg[8][4]/NET0131  & n1474 ;
  assign n12856 = ~n12847 & ~n12848 ;
  assign n12857 = n12855 & n12856 ;
  assign n12841 = \P2_InstQueue_reg[9][4]/NET0131  & n1447 ;
  assign n12842 = \P2_InstQueue_reg[13][4]/NET0131  & n1453 ;
  assign n12853 = ~n12841 & ~n12842 ;
  assign n12843 = \P2_InstQueue_reg[5][4]/NET0131  & n1468 ;
  assign n12844 = \P2_InstQueue_reg[11][4]/NET0131  & n1461 ;
  assign n12854 = ~n12843 & ~n12844 ;
  assign n12858 = n12853 & n12854 ;
  assign n12862 = n12857 & n12858 ;
  assign n12863 = n12861 & n12862 ;
  assign n12864 = n12832 & ~n12863 ;
  assign n12869 = \P2_InstQueue_reg[2][5]/NET0131  & n1478 ;
  assign n12870 = \P2_InstQueue_reg[0][5]/NET0131  & n1466 ;
  assign n12883 = ~n12869 & ~n12870 ;
  assign n12871 = \P2_InstQueue_reg[15][5]/NET0131  & n1480 ;
  assign n12872 = \P2_InstQueue_reg[14][5]/NET0131  & n1459 ;
  assign n12884 = ~n12871 & ~n12872 ;
  assign n12891 = n12883 & n12884 ;
  assign n12865 = \P2_InstQueue_reg[4][5]/NET0131  & n1464 ;
  assign n12866 = \P2_InstQueue_reg[10][5]/NET0131  & n1476 ;
  assign n12881 = ~n12865 & ~n12866 ;
  assign n12867 = \P2_InstQueue_reg[3][5]/NET0131  & n1456 ;
  assign n12868 = \P2_InstQueue_reg[6][5]/NET0131  & n1470 ;
  assign n12882 = ~n12867 & ~n12868 ;
  assign n12892 = n12881 & n12882 ;
  assign n12893 = n12891 & n12892 ;
  assign n12877 = \P2_InstQueue_reg[1][5]/NET0131  & n1482 ;
  assign n12878 = \P2_InstQueue_reg[7][5]/NET0131  & n1450 ;
  assign n12887 = ~n12877 & ~n12878 ;
  assign n12879 = \P2_InstQueue_reg[12][5]/NET0131  & n1472 ;
  assign n12880 = \P2_InstQueue_reg[8][5]/NET0131  & n1474 ;
  assign n12888 = ~n12879 & ~n12880 ;
  assign n12889 = n12887 & n12888 ;
  assign n12873 = \P2_InstQueue_reg[9][5]/NET0131  & n1447 ;
  assign n12874 = \P2_InstQueue_reg[13][5]/NET0131  & n1453 ;
  assign n12885 = ~n12873 & ~n12874 ;
  assign n12875 = \P2_InstQueue_reg[5][5]/NET0131  & n1468 ;
  assign n12876 = \P2_InstQueue_reg[11][5]/NET0131  & n1461 ;
  assign n12886 = ~n12875 & ~n12876 ;
  assign n12890 = n12885 & n12886 ;
  assign n12894 = n12889 & n12890 ;
  assign n12895 = n12893 & n12894 ;
  assign n12896 = n12864 & ~n12895 ;
  assign n12901 = \P2_InstQueue_reg[2][6]/NET0131  & n1478 ;
  assign n12902 = \P2_InstQueue_reg[0][6]/NET0131  & n1466 ;
  assign n12915 = ~n12901 & ~n12902 ;
  assign n12903 = \P2_InstQueue_reg[15][6]/NET0131  & n1480 ;
  assign n12904 = \P2_InstQueue_reg[14][6]/NET0131  & n1459 ;
  assign n12916 = ~n12903 & ~n12904 ;
  assign n12923 = n12915 & n12916 ;
  assign n12897 = \P2_InstQueue_reg[4][6]/NET0131  & n1464 ;
  assign n12898 = \P2_InstQueue_reg[10][6]/NET0131  & n1476 ;
  assign n12913 = ~n12897 & ~n12898 ;
  assign n12899 = \P2_InstQueue_reg[3][6]/NET0131  & n1456 ;
  assign n12900 = \P2_InstQueue_reg[6][6]/NET0131  & n1470 ;
  assign n12914 = ~n12899 & ~n12900 ;
  assign n12924 = n12913 & n12914 ;
  assign n12925 = n12923 & n12924 ;
  assign n12909 = \P2_InstQueue_reg[1][6]/NET0131  & n1482 ;
  assign n12910 = \P2_InstQueue_reg[7][6]/NET0131  & n1450 ;
  assign n12919 = ~n12909 & ~n12910 ;
  assign n12911 = \P2_InstQueue_reg[12][6]/NET0131  & n1472 ;
  assign n12912 = \P2_InstQueue_reg[8][6]/NET0131  & n1474 ;
  assign n12920 = ~n12911 & ~n12912 ;
  assign n12921 = n12919 & n12920 ;
  assign n12905 = \P2_InstQueue_reg[9][6]/NET0131  & n1447 ;
  assign n12906 = \P2_InstQueue_reg[13][6]/NET0131  & n1453 ;
  assign n12917 = ~n12905 & ~n12906 ;
  assign n12907 = \P2_InstQueue_reg[5][6]/NET0131  & n1468 ;
  assign n12908 = \P2_InstQueue_reg[11][6]/NET0131  & n1461 ;
  assign n12918 = ~n12907 & ~n12908 ;
  assign n12922 = n12917 & n12918 ;
  assign n12926 = n12921 & n12922 ;
  assign n12927 = n12925 & n12926 ;
  assign n12928 = n12896 & ~n12927 ;
  assign n12933 = \P2_InstQueue_reg[2][7]/NET0131  & n1478 ;
  assign n12934 = \P2_InstQueue_reg[4][7]/NET0131  & n1464 ;
  assign n12947 = ~n12933 & ~n12934 ;
  assign n12935 = \P2_InstQueue_reg[0][7]/NET0131  & n1466 ;
  assign n12936 = \P2_InstQueue_reg[14][7]/NET0131  & n1459 ;
  assign n12948 = ~n12935 & ~n12936 ;
  assign n12955 = n12947 & n12948 ;
  assign n12929 = \P2_InstQueue_reg[15][7]/NET0131  & n1480 ;
  assign n12930 = \P2_InstQueue_reg[10][7]/NET0131  & n1476 ;
  assign n12945 = ~n12929 & ~n12930 ;
  assign n12931 = \P2_InstQueue_reg[3][7]/NET0131  & n1456 ;
  assign n12932 = \P2_InstQueue_reg[6][7]/NET0131  & n1470 ;
  assign n12946 = ~n12931 & ~n12932 ;
  assign n12956 = n12945 & n12946 ;
  assign n12957 = n12955 & n12956 ;
  assign n12941 = \P2_InstQueue_reg[1][7]/NET0131  & n1482 ;
  assign n12942 = \P2_InstQueue_reg[7][7]/NET0131  & n1450 ;
  assign n12951 = ~n12941 & ~n12942 ;
  assign n12943 = \P2_InstQueue_reg[12][7]/NET0131  & n1472 ;
  assign n12944 = \P2_InstQueue_reg[8][7]/NET0131  & n1474 ;
  assign n12952 = ~n12943 & ~n12944 ;
  assign n12953 = n12951 & n12952 ;
  assign n12937 = \P2_InstQueue_reg[9][7]/NET0131  & n1447 ;
  assign n12938 = \P2_InstQueue_reg[13][7]/NET0131  & n1453 ;
  assign n12949 = ~n12937 & ~n12938 ;
  assign n12939 = \P2_InstQueue_reg[5][7]/NET0131  & n1468 ;
  assign n12940 = \P2_InstQueue_reg[11][7]/NET0131  & n1461 ;
  assign n12950 = ~n12939 & ~n12940 ;
  assign n12954 = n12949 & n12950 ;
  assign n12958 = n12953 & n12954 ;
  assign n12959 = n12957 & n12958 ;
  assign n12960 = n1798 & ~n12959 ;
  assign n12961 = n1726 & n12960 ;
  assign n12962 = n12928 & n12961 ;
  assign n12963 = ~n12673 & ~n12962 ;
  assign n12964 = ~n12671 & n12963 ;
  assign n12965 = n1927 & ~n12964 ;
  assign n12966 = ~n12633 & ~n12965 ;
  assign n12970 = \P2_PhyAddrPointer_reg[21]/NET0131  & n1897 ;
  assign n12975 = ~n6595 & ~n6669 ;
  assign n12976 = ~n7527 & ~n12975 ;
  assign n12977 = n6188 & ~n12976 ;
  assign n12971 = ~n6542 & ~n6546 ;
  assign n12972 = n6542 & n6546 ;
  assign n12973 = ~n12971 & ~n12972 ;
  assign n12974 = ~n6188 & ~n12973 ;
  assign n12978 = ~n1897 & ~n12974 ;
  assign n12979 = ~n12977 & n12978 ;
  assign n12980 = ~n12970 & ~n12979 ;
  assign n12981 = n1734 & ~n12980 ;
  assign n12982 = \P2_PhyAddrPointer_reg[21]/NET0131  & ~n8936 ;
  assign n12983 = ~n6761 & ~n6766 ;
  assign n12984 = n1890 & ~n6767 ;
  assign n12985 = ~n12983 & n12984 ;
  assign n12986 = ~n12982 & ~n12985 ;
  assign n12987 = ~n12981 & n12986 ;
  assign n12988 = n1927 & ~n12987 ;
  assign n12989 = n8977 & ~n10965 ;
  assign n12991 = \P2_PhyAddrPointer_reg[21]/NET0131  & n12989 ;
  assign n12990 = ~\P2_PhyAddrPointer_reg[21]/NET0131  & ~n12989 ;
  assign n12992 = n1931 & ~n12990 ;
  assign n12993 = ~n12991 & n12992 ;
  assign n12967 = ~\P2_PhyAddrPointer_reg[21]/NET0131  & ~n11876 ;
  assign n12968 = ~n11896 & ~n12967 ;
  assign n12969 = n3087 & n12968 ;
  assign n12994 = \P2_rEIP_reg[21]/NET0131  & n3113 ;
  assign n12995 = \P2_PhyAddrPointer_reg[21]/NET0131  & ~n8958 ;
  assign n12996 = ~n12994 & ~n12995 ;
  assign n12997 = ~n12969 & n12996 ;
  assign n12998 = ~n12993 & n12997 ;
  assign n12999 = ~n12988 & n12998 ;
  assign n13000 = \P2_PhyAddrPointer_reg[25]/NET0131  & n1897 ;
  assign n13001 = ~n8517 & ~n13000 ;
  assign n13002 = n1734 & ~n13001 ;
  assign n13003 = \P2_PhyAddrPointer_reg[25]/NET0131  & ~n8936 ;
  assign n13004 = ~n8524 & ~n13003 ;
  assign n13005 = ~n13002 & n13004 ;
  assign n13006 = n1927 & ~n13005 ;
  assign n13010 = ~\P2_PhyAddrPointer_reg[25]/NET0131  & ~n8995 ;
  assign n13011 = ~n8996 & ~n13010 ;
  assign n13012 = n9005 & n13011 ;
  assign n13007 = ~\P2_PhyAddrPointer_reg[25]/NET0131  & ~n8981 ;
  assign n13008 = n3034 & ~n8982 ;
  assign n13009 = ~n13007 & n13008 ;
  assign n13013 = \P2_PhyAddrPointer_reg[25]/NET0131  & ~n8958 ;
  assign n13014 = ~n8506 & ~n13013 ;
  assign n13015 = ~n13009 & n13014 ;
  assign n13016 = ~n13012 & n13015 ;
  assign n13017 = ~n13006 & n13016 ;
  assign n13018 = \P2_PhyAddrPointer_reg[8]/NET0131  & n1897 ;
  assign n13020 = ~n6459 & ~n10223 ;
  assign n13019 = n6459 & n7429 ;
  assign n13021 = ~n6188 & ~n13019 ;
  assign n13022 = ~n13020 & n13021 ;
  assign n13023 = ~n6603 & n7455 ;
  assign n13024 = n6188 & ~n8443 ;
  assign n13025 = ~n13023 & n13024 ;
  assign n13026 = ~n13022 & ~n13025 ;
  assign n13027 = ~n1897 & ~n13026 ;
  assign n13028 = ~n13018 & ~n13027 ;
  assign n13029 = n1734 & ~n13028 ;
  assign n13030 = \P2_PhyAddrPointer_reg[8]/NET0131  & ~n8936 ;
  assign n13031 = ~n6733 & ~n7545 ;
  assign n13033 = n6736 & n13031 ;
  assign n13032 = ~n6736 & ~n13031 ;
  assign n13034 = n1890 & ~n13032 ;
  assign n13035 = ~n13033 & n13034 ;
  assign n13036 = ~n13030 & ~n13035 ;
  assign n13037 = ~n13029 & n13036 ;
  assign n13038 = n1927 & ~n13037 ;
  assign n13042 = \P2_PhyAddrPointer_reg[1]/NET0131  & n8962 ;
  assign n13043 = \P2_PhyAddrPointer_reg[6]/NET0131  & n13042 ;
  assign n13044 = \P2_PhyAddrPointer_reg[7]/NET0131  & n13043 ;
  assign n13045 = ~\P2_PhyAddrPointer_reg[8]/NET0131  & ~n13044 ;
  assign n13046 = \P2_PhyAddrPointer_reg[8]/NET0131  & n13044 ;
  assign n13047 = ~n13045 & ~n13046 ;
  assign n13048 = n9005 & n13047 ;
  assign n13039 = ~\P2_PhyAddrPointer_reg[8]/NET0131  & ~n8964 ;
  assign n13040 = n3034 & ~n8965 ;
  assign n13041 = ~n13039 & n13040 ;
  assign n13049 = \P2_rEIP_reg[8]/NET0131  & n3113 ;
  assign n13050 = \P2_PhyAddrPointer_reg[8]/NET0131  & ~n8958 ;
  assign n13051 = ~n13049 & ~n13050 ;
  assign n13052 = ~n13041 & n13051 ;
  assign n13053 = ~n13048 & n13052 ;
  assign n13054 = ~n13038 & n13053 ;
  assign n13058 = \P3_PhyAddrPointer_reg[12]/NET0131  & n2896 ;
  assign n13059 = ~n9082 & ~n13058 ;
  assign n13060 = n2894 & ~n13059 ;
  assign n13061 = \P3_PhyAddrPointer_reg[12]/NET0131  & ~n9014 ;
  assign n13062 = ~n9111 & ~n13061 ;
  assign n13063 = ~n13060 & n13062 ;
  assign n13064 = n2453 & ~n13063 ;
  assign n13055 = ~\P3_PhyAddrPointer_reg[12]/NET0131  & ~n11962 ;
  assign n13056 = ~n12007 & ~n13055 ;
  assign n13065 = ~\P3_DataWidth_reg[1]/NET0131  & ~n13056 ;
  assign n13066 = ~\P3_PhyAddrPointer_reg[12]/NET0131  & ~n9028 ;
  assign n13067 = ~n9029 & ~n13066 ;
  assign n13068 = \P3_DataWidth_reg[1]/NET0131  & ~n13067 ;
  assign n13069 = n2959 & ~n13068 ;
  assign n13070 = ~n13065 & n13069 ;
  assign n13057 = n4415 & n13056 ;
  assign n13071 = \P3_PhyAddrPointer_reg[12]/NET0131  & ~n9063 ;
  assign n13072 = ~n9070 & ~n13071 ;
  assign n13073 = ~n13057 & n13072 ;
  assign n13074 = ~n13070 & n13073 ;
  assign n13075 = ~n13064 & n13074 ;
  assign n13076 = \P3_PhyAddrPointer_reg[13]/NET0131  & n2896 ;
  assign n13082 = n4175 & ~n8339 ;
  assign n13081 = ~n4175 & n8339 ;
  assign n13083 = ~n3753 & ~n13081 ;
  assign n13084 = ~n13082 & n13083 ;
  assign n13077 = ~n8357 & ~n8358 ;
  assign n13078 = n4059 & n6088 ;
  assign n13079 = ~n13077 & ~n13078 ;
  assign n13080 = n3753 & ~n13079 ;
  assign n13085 = ~n2896 & ~n13080 ;
  assign n13086 = ~n13084 & n13085 ;
  assign n13087 = ~n13076 & ~n13086 ;
  assign n13088 = n2894 & ~n13087 ;
  assign n13089 = \P3_PhyAddrPointer_reg[13]/NET0131  & ~n9014 ;
  assign n13090 = ~\P3_InstAddrPointer_reg[13]/NET0131  & ~n4350 ;
  assign n13091 = ~n4351 & ~n13090 ;
  assign n13092 = n4306 & ~n4348 ;
  assign n13093 = ~n13091 & ~n13092 ;
  assign n13094 = n2905 & ~n4349 ;
  assign n13095 = ~n13093 & n13094 ;
  assign n13096 = ~n13089 & ~n13095 ;
  assign n13097 = ~n13088 & n13096 ;
  assign n13098 = n2453 & ~n13097 ;
  assign n13103 = ~\P3_PhyAddrPointer_reg[13]/NET0131  & ~n12007 ;
  assign n13104 = ~n12008 & ~n13103 ;
  assign n13105 = n4415 & n13104 ;
  assign n13099 = n9029 & ~n11124 ;
  assign n13100 = ~\P3_PhyAddrPointer_reg[13]/NET0131  & ~n13099 ;
  assign n13101 = n2959 & ~n12000 ;
  assign n13102 = ~n13100 & n13101 ;
  assign n13106 = \P3_rEIP_reg[13]/NET0131  & n4412 ;
  assign n13107 = \P3_PhyAddrPointer_reg[13]/NET0131  & ~n9063 ;
  assign n13108 = ~n13106 & ~n13107 ;
  assign n13109 = ~n13102 & n13108 ;
  assign n13110 = ~n13105 & n13109 ;
  assign n13111 = ~n13098 & n13110 ;
  assign n13113 = ~n4066 & ~n13078 ;
  assign n13114 = ~n4075 & ~n13113 ;
  assign n13115 = n3753 & ~n13114 ;
  assign n13116 = n4171 & ~n7371 ;
  assign n13117 = ~n3753 & ~n4232 ;
  assign n13118 = ~n13116 & n13117 ;
  assign n13119 = ~n2896 & ~n13118 ;
  assign n13120 = ~n13115 & n13119 ;
  assign n13121 = n2894 & n13120 ;
  assign n13122 = \P3_PhyAddrPointer_reg[14]/NET0131  & ~n11965 ;
  assign n13124 = ~n4354 & ~n6125 ;
  assign n13123 = n4354 & n6125 ;
  assign n13125 = n2905 & ~n13123 ;
  assign n13126 = ~n13124 & n13125 ;
  assign n13127 = ~n13122 & ~n13126 ;
  assign n13128 = ~n13121 & n13127 ;
  assign n13129 = n2453 & ~n13128 ;
  assign n13133 = ~\P3_PhyAddrPointer_reg[14]/NET0131  & ~n12000 ;
  assign n13134 = n12002 & ~n13133 ;
  assign n13130 = ~\P3_PhyAddrPointer_reg[14]/NET0131  & ~n12008 ;
  assign n13131 = ~n12009 & ~n13130 ;
  assign n13132 = n4415 & n13131 ;
  assign n13112 = \P3_PhyAddrPointer_reg[14]/NET0131  & ~n9063 ;
  assign n13135 = \P3_rEIP_reg[14]/NET0131  & n4412 ;
  assign n13136 = ~n13112 & ~n13135 ;
  assign n13137 = ~n13132 & n13136 ;
  assign n13138 = ~n13134 & n13137 ;
  assign n13139 = ~n13129 & n13138 ;
  assign n13149 = ~n4237 & ~n6060 ;
  assign n13150 = n4237 & n6060 ;
  assign n13151 = ~n13149 & ~n13150 ;
  assign n13152 = ~n3753 & ~n13151 ;
  assign n13153 = ~n4079 & ~n7333 ;
  assign n13154 = n4079 & n7333 ;
  assign n13155 = ~n13153 & ~n13154 ;
  assign n13156 = n3753 & ~n13155 ;
  assign n13157 = ~n2896 & ~n13156 ;
  assign n13158 = ~n13152 & n13157 ;
  assign n13159 = n2894 & n13158 ;
  assign n13160 = \P3_PhyAddrPointer_reg[16]/NET0131  & ~n11965 ;
  assign n13161 = ~\P3_InstAddrPointer_reg[16]/NET0131  & ~n7345 ;
  assign n13162 = ~n4357 & ~n13161 ;
  assign n13163 = \P3_InstAddrPointer_reg[15]/NET0131  & n13123 ;
  assign n13164 = ~n13162 & ~n13163 ;
  assign n13165 = n2905 & ~n6126 ;
  assign n13166 = ~n13164 & n13165 ;
  assign n13167 = ~n13160 & ~n13166 ;
  assign n13168 = ~n13159 & n13167 ;
  assign n13169 = n2453 & ~n13168 ;
  assign n13143 = ~\P3_PhyAddrPointer_reg[16]/NET0131  & ~n12012 ;
  assign n13144 = n9032 & n12008 ;
  assign n13145 = ~n13143 & ~n13144 ;
  assign n13146 = n10076 & n13145 ;
  assign n13140 = ~\P3_PhyAddrPointer_reg[16]/NET0131  & ~n12011 ;
  assign n13141 = n2970 & ~n9033 ;
  assign n13142 = ~n13140 & n13141 ;
  assign n13147 = \P3_PhyAddrPointer_reg[16]/NET0131  & ~n9063 ;
  assign n13148 = \P3_rEIP_reg[16]/NET0131  & n4412 ;
  assign n13170 = ~n13147 & ~n13148 ;
  assign n13171 = ~n13142 & n13170 ;
  assign n13172 = ~n13146 & n13171 ;
  assign n13173 = ~n13169 & n13172 ;
  assign n13174 = ~n3794 & ~n7379 ;
  assign n13175 = ~n7382 & ~n13174 ;
  assign n13176 = ~n4085 & ~n13175 ;
  assign n13177 = n3753 & ~n13176 ;
  assign n13179 = ~n4248 & n7372 ;
  assign n13178 = n4248 & ~n7372 ;
  assign n13180 = ~n3753 & ~n13178 ;
  assign n13181 = ~n13179 & n13180 ;
  assign n13182 = ~n13177 & ~n13181 ;
  assign n13183 = n2904 & n13182 ;
  assign n13184 = \P3_PhyAddrPointer_reg[18]/NET0131  & ~n11965 ;
  assign n13186 = ~\P3_InstAddrPointer_reg[18]/NET0131  & ~n4359 ;
  assign n13187 = ~n4363 & ~n13186 ;
  assign n13188 = ~n12040 & ~n13187 ;
  assign n13185 = \P3_InstAddrPointer_reg[18]/NET0131  & n12040 ;
  assign n13189 = n2905 & ~n13185 ;
  assign n13190 = ~n13188 & n13189 ;
  assign n13191 = ~n13184 & ~n13190 ;
  assign n13192 = ~n13183 & n13191 ;
  assign n13193 = n2453 & ~n13192 ;
  assign n13198 = \P3_PhyAddrPointer_reg[1]/NET0131  & n9034 ;
  assign n13199 = ~\P3_PhyAddrPointer_reg[18]/NET0131  & ~n13198 ;
  assign n13200 = \P3_PhyAddrPointer_reg[18]/NET0131  & n13198 ;
  assign n13201 = ~n13199 & ~n13200 ;
  assign n13202 = n10076 & n13201 ;
  assign n13195 = ~\P3_PhyAddrPointer_reg[18]/NET0131  & ~n9034 ;
  assign n13194 = \P3_PhyAddrPointer_reg[18]/NET0131  & n9034 ;
  assign n13196 = n2970 & ~n13194 ;
  assign n13197 = ~n13195 & n13196 ;
  assign n13203 = \P3_PhyAddrPointer_reg[18]/NET0131  & ~n9063 ;
  assign n13204 = \P3_rEIP_reg[18]/NET0131  & n4412 ;
  assign n13205 = ~n13203 & ~n13204 ;
  assign n13206 = ~n13197 & n13205 ;
  assign n13207 = ~n13202 & n13206 ;
  assign n13208 = ~n13193 & n13207 ;
  assign n13210 = \P3_PhyAddrPointer_reg[21]/NET0131  & n2896 ;
  assign n13211 = ~n8368 & ~n13210 ;
  assign n13212 = n2894 & ~n13211 ;
  assign n13213 = \P3_PhyAddrPointer_reg[21]/NET0131  & ~n9014 ;
  assign n13214 = ~n8380 & ~n13213 ;
  assign n13215 = ~n13212 & n13214 ;
  assign n13216 = n2453 & ~n13215 ;
  assign n13221 = n9034 & ~n11124 ;
  assign n13222 = n9036 & n13221 ;
  assign n13223 = ~\P3_PhyAddrPointer_reg[21]/NET0131  & ~n13222 ;
  assign n13220 = n9038 & ~n11124 ;
  assign n13224 = n2959 & ~n13220 ;
  assign n13225 = ~n13223 & n13224 ;
  assign n13217 = ~\P3_PhyAddrPointer_reg[21]/NET0131  & ~n12054 ;
  assign n13218 = ~n12073 & ~n13217 ;
  assign n13219 = n4415 & n13218 ;
  assign n13209 = \P3_PhyAddrPointer_reg[21]/NET0131  & ~n9063 ;
  assign n13226 = ~n8336 & ~n13209 ;
  assign n13227 = ~n13219 & n13226 ;
  assign n13228 = ~n13225 & n13227 ;
  assign n13229 = ~n13216 & n13228 ;
  assign n13230 = \P3_PhyAddrPointer_reg[25]/NET0131  & n2896 ;
  assign n13231 = ~n8409 & ~n13230 ;
  assign n13232 = n2894 & ~n13231 ;
  assign n13233 = \P3_PhyAddrPointer_reg[25]/NET0131  & ~n9014 ;
  assign n13234 = ~n8417 & ~n13233 ;
  assign n13235 = ~n13232 & n13234 ;
  assign n13236 = n2453 & ~n13235 ;
  assign n13241 = ~\P3_PhyAddrPointer_reg[25]/NET0131  & ~n12106 ;
  assign n13242 = ~n12142 & ~n13241 ;
  assign n13243 = n10076 & n13242 ;
  assign n13238 = ~\P3_PhyAddrPointer_reg[25]/NET0131  & ~n12101 ;
  assign n13239 = n2970 & ~n12137 ;
  assign n13240 = ~n13238 & n13239 ;
  assign n13237 = \P3_PhyAddrPointer_reg[25]/NET0131  & ~n9063 ;
  assign n13244 = ~n8430 & ~n13237 ;
  assign n13245 = ~n13240 & n13244 ;
  assign n13246 = ~n13243 & n13245 ;
  assign n13247 = ~n13236 & n13246 ;
  assign n13256 = n2894 & n9135 ;
  assign n13255 = \P3_PhyAddrPointer_reg[8]/NET0131  & ~n11965 ;
  assign n13257 = ~n9149 & ~n13255 ;
  assign n13258 = ~n13256 & n13257 ;
  assign n13259 = n2453 & ~n13258 ;
  assign n13248 = \P3_PhyAddrPointer_reg[1]/NET0131  & n9022 ;
  assign n13249 = \P3_PhyAddrPointer_reg[6]/NET0131  & n13248 ;
  assign n13250 = \P3_PhyAddrPointer_reg[7]/NET0131  & n13249 ;
  assign n13251 = ~\P3_PhyAddrPointer_reg[8]/NET0131  & ~n13250 ;
  assign n13252 = \P3_PhyAddrPointer_reg[1]/NET0131  & n9025 ;
  assign n13253 = ~n13251 & ~n13252 ;
  assign n13260 = ~\P3_DataWidth_reg[1]/NET0131  & ~n13253 ;
  assign n13261 = ~\P3_PhyAddrPointer_reg[8]/NET0131  & ~n9024 ;
  assign n13262 = ~n9025 & ~n13261 ;
  assign n13263 = \P3_DataWidth_reg[1]/NET0131  & ~n13262 ;
  assign n13264 = n2959 & ~n13263 ;
  assign n13265 = ~n13260 & n13264 ;
  assign n13254 = n4415 & n13253 ;
  assign n13266 = \P3_PhyAddrPointer_reg[8]/NET0131  & ~n9063 ;
  assign n13267 = ~n9120 & ~n13266 ;
  assign n13268 = ~n13254 & n13267 ;
  assign n13269 = ~n13265 & n13268 ;
  assign n13270 = ~n13259 & n13269 ;
  assign n13271 = \P1_PhyAddrPointer_reg[12]/NET0131  & n2375 ;
  assign n13272 = ~n9304 & ~n13271 ;
  assign n13273 = n2244 & ~n13272 ;
  assign n13274 = \P1_PhyAddrPointer_reg[12]/NET0131  & ~n10087 ;
  assign n13275 = ~n9313 & ~n13274 ;
  assign n13276 = ~n13273 & n13275 ;
  assign n13277 = n2432 & ~n13276 ;
  assign n13283 = ~\P1_PhyAddrPointer_reg[12]/NET0131  & ~n12155 ;
  assign n13284 = ~n12217 & ~n13283 ;
  assign n13285 = n5095 & n13284 ;
  assign n13278 = n10100 & ~n11332 ;
  assign n13280 = \P1_PhyAddrPointer_reg[12]/NET0131  & n13278 ;
  assign n13279 = ~\P1_PhyAddrPointer_reg[12]/NET0131  & ~n13278 ;
  assign n13281 = n2436 & ~n13279 ;
  assign n13282 = ~n13280 & n13281 ;
  assign n13286 = \P1_PhyAddrPointer_reg[12]/NET0131  & ~n10136 ;
  assign n13287 = ~n9292 & ~n13286 ;
  assign n13288 = ~n13282 & n13287 ;
  assign n13289 = ~n13285 & n13288 ;
  assign n13290 = ~n13277 & n13289 ;
  assign n13298 = \P1_PhyAddrPointer_reg[13]/NET0131  & n2375 ;
  assign n13302 = ~n4788 & ~n12200 ;
  assign n13303 = ~n12201 & ~n13302 ;
  assign n13304 = n4453 & ~n13303 ;
  assign n13299 = n4882 & ~n5956 ;
  assign n13300 = ~n4453 & ~n5957 ;
  assign n13301 = ~n13299 & n13300 ;
  assign n13305 = ~n2375 & ~n13301 ;
  assign n13306 = ~n13304 & n13305 ;
  assign n13307 = ~n13298 & ~n13306 ;
  assign n13308 = n2244 & ~n13307 ;
  assign n13291 = ~\P1_InstAddrPointer_reg[13]/NET0131  & ~n4964 ;
  assign n13292 = ~n4965 & ~n13291 ;
  assign n13293 = \P1_InstAddrPointer_reg[12]/NET0131  & n12159 ;
  assign n13295 = n13292 & n13293 ;
  assign n13294 = ~n13292 & ~n13293 ;
  assign n13296 = n2385 & ~n13294 ;
  assign n13297 = ~n13295 & n13296 ;
  assign n13309 = \P1_PhyAddrPointer_reg[13]/NET0131  & ~n10087 ;
  assign n13310 = ~n13297 & ~n13309 ;
  assign n13311 = ~n13308 & n13310 ;
  assign n13312 = n2432 & ~n13311 ;
  assign n13316 = ~\P1_PhyAddrPointer_reg[13]/NET0131  & ~n12217 ;
  assign n13317 = ~n12218 & ~n13316 ;
  assign n13318 = n10133 & n13317 ;
  assign n13313 = ~\P1_PhyAddrPointer_reg[13]/NET0131  & ~n10101 ;
  assign n13314 = n3148 & ~n10102 ;
  assign n13315 = ~n13313 & n13314 ;
  assign n13319 = \P1_PhyAddrPointer_reg[13]/NET0131  & ~n10136 ;
  assign n13320 = \P1_rEIP_reg[13]/NET0131  & n5092 ;
  assign n13321 = ~n13319 & ~n13320 ;
  assign n13322 = ~n13315 & n13321 ;
  assign n13323 = ~n13318 & n13322 ;
  assign n13324 = ~n13312 & n13323 ;
  assign n13329 = \P1_PhyAddrPointer_reg[14]/NET0131  & n2375 ;
  assign n13334 = ~\P1_InstAddrPointer_reg[14]/NET0131  & ~n4465 ;
  assign n13335 = ~n12197 & ~n13334 ;
  assign n13336 = ~n12201 & ~n13335 ;
  assign n13337 = ~n12202 & ~n13336 ;
  assign n13338 = n4453 & ~n13337 ;
  assign n13331 = n4887 & ~n4931 ;
  assign n13330 = ~n4887 & n4931 ;
  assign n13332 = ~n4453 & ~n13330 ;
  assign n13333 = ~n13331 & n13332 ;
  assign n13339 = ~n2375 & ~n13333 ;
  assign n13340 = ~n13338 & n13339 ;
  assign n13341 = ~n13329 & ~n13340 ;
  assign n13342 = n2244 & ~n13341 ;
  assign n13326 = n5028 & n5034 ;
  assign n13325 = ~n5028 & ~n5034 ;
  assign n13327 = n2385 & ~n13325 ;
  assign n13328 = ~n13326 & n13327 ;
  assign n13343 = \P1_PhyAddrPointer_reg[14]/NET0131  & ~n10087 ;
  assign n13344 = ~n13328 & ~n13343 ;
  assign n13345 = ~n13342 & n13344 ;
  assign n13346 = n2432 & ~n13345 ;
  assign n13350 = ~\P1_PhyAddrPointer_reg[14]/NET0131  & ~n12218 ;
  assign n13351 = ~n12219 & ~n13350 ;
  assign n13352 = n10133 & n13351 ;
  assign n13347 = ~\P1_PhyAddrPointer_reg[14]/NET0131  & ~n10102 ;
  assign n13348 = n3148 & ~n10103 ;
  assign n13349 = ~n13347 & n13348 ;
  assign n13353 = \P1_rEIP_reg[14]/NET0131  & n5092 ;
  assign n13354 = \P1_PhyAddrPointer_reg[14]/NET0131  & ~n10136 ;
  assign n13355 = ~n13353 & ~n13354 ;
  assign n13356 = ~n13349 & n13355 ;
  assign n13357 = ~n13352 & n13356 ;
  assign n13358 = ~n13346 & n13357 ;
  assign n13366 = \P1_PhyAddrPointer_reg[16]/NET0131  & n2375 ;
  assign n13371 = ~n4784 & ~n6832 ;
  assign n13372 = n4784 & n6832 ;
  assign n13373 = ~n13371 & ~n13372 ;
  assign n13374 = n4453 & ~n13373 ;
  assign n13367 = ~n4918 & ~n7276 ;
  assign n13368 = n4918 & n7276 ;
  assign n13369 = ~n13367 & ~n13368 ;
  assign n13370 = ~n4453 & ~n13369 ;
  assign n13375 = ~n2375 & ~n13370 ;
  assign n13376 = ~n13374 & n13375 ;
  assign n13377 = ~n13366 & ~n13376 ;
  assign n13378 = n2244 & ~n13377 ;
  assign n13363 = n5032 & n7300 ;
  assign n13362 = ~n5032 & ~n7300 ;
  assign n13364 = n2385 & ~n13362 ;
  assign n13365 = ~n13363 & n13364 ;
  assign n13379 = \P1_PhyAddrPointer_reg[16]/NET0131  & ~n10087 ;
  assign n13380 = ~n13365 & ~n13379 ;
  assign n13381 = ~n13378 & n13380 ;
  assign n13382 = n2432 & ~n13381 ;
  assign n13385 = n10105 & ~n11332 ;
  assign n13383 = n10104 & ~n11332 ;
  assign n13384 = ~\P1_PhyAddrPointer_reg[16]/NET0131  & ~n13383 ;
  assign n13386 = n2436 & ~n13384 ;
  assign n13387 = ~n13385 & n13386 ;
  assign n13359 = ~\P1_PhyAddrPointer_reg[16]/NET0131  & ~n12221 ;
  assign n13360 = ~n10123 & ~n13359 ;
  assign n13361 = n5095 & n13360 ;
  assign n13388 = \P1_rEIP_reg[16]/NET0131  & n5092 ;
  assign n13389 = \P1_PhyAddrPointer_reg[16]/NET0131  & ~n10136 ;
  assign n13390 = ~n13388 & ~n13389 ;
  assign n13391 = ~n13361 & n13390 ;
  assign n13392 = ~n13387 & n13391 ;
  assign n13393 = ~n13382 & n13392 ;
  assign n13394 = \P1_PhyAddrPointer_reg[17]/NET0131  & n2375 ;
  assign n13395 = ~n9345 & ~n13394 ;
  assign n13396 = n2244 & ~n13395 ;
  assign n13397 = \P1_PhyAddrPointer_reg[17]/NET0131  & ~n10087 ;
  assign n13398 = ~n9356 & ~n13397 ;
  assign n13399 = ~n13396 & n13398 ;
  assign n13400 = n2432 & ~n13399 ;
  assign n13404 = ~\P1_PhyAddrPointer_reg[17]/NET0131  & ~n10123 ;
  assign n13405 = ~n10124 & ~n13404 ;
  assign n13406 = n10133 & n13405 ;
  assign n13401 = ~\P1_PhyAddrPointer_reg[17]/NET0131  & ~n10105 ;
  assign n13402 = n3148 & ~n10106 ;
  assign n13403 = ~n13401 & n13402 ;
  assign n13407 = \P1_PhyAddrPointer_reg[17]/NET0131  & ~n10136 ;
  assign n13408 = ~n9332 & ~n13407 ;
  assign n13409 = ~n13403 & n13408 ;
  assign n13410 = ~n13406 & n13409 ;
  assign n13411 = ~n13400 & n13410 ;
  assign n13412 = \P1_PhyAddrPointer_reg[18]/NET0131  & n2375 ;
  assign n13413 = ~n8557 & ~n13412 ;
  assign n13414 = n2244 & ~n13413 ;
  assign n13415 = \P1_PhyAddrPointer_reg[18]/NET0131  & ~n10087 ;
  assign n13416 = ~n8563 & ~n13415 ;
  assign n13417 = ~n13414 & n13416 ;
  assign n13418 = n2432 & ~n13417 ;
  assign n13420 = ~\P1_PhyAddrPointer_reg[18]/NET0131  & ~n10124 ;
  assign n13421 = ~n12237 & ~n13420 ;
  assign n13422 = n10133 & n13421 ;
  assign n13423 = ~\P1_PhyAddrPointer_reg[18]/NET0131  & ~n10106 ;
  assign n13424 = n12231 & ~n13423 ;
  assign n13419 = \P1_PhyAddrPointer_reg[18]/NET0131  & ~n10136 ;
  assign n13425 = ~n8584 & ~n13419 ;
  assign n13426 = ~n13424 & n13425 ;
  assign n13427 = ~n13422 & n13426 ;
  assign n13428 = ~n13418 & n13427 ;
  assign n13443 = \P1_PhyAddrPointer_reg[21]/NET0131  & n2375 ;
  assign n13448 = ~n4769 & ~n5975 ;
  assign n13449 = ~n4795 & ~n13448 ;
  assign n13450 = n4453 & ~n13449 ;
  assign n13444 = ~n4900 & ~n7282 ;
  assign n13445 = n4900 & n7282 ;
  assign n13446 = ~n13444 & ~n13445 ;
  assign n13447 = ~n4453 & ~n13446 ;
  assign n13451 = ~n2375 & ~n13447 ;
  assign n13452 = ~n13450 & n13451 ;
  assign n13453 = ~n13443 & ~n13452 ;
  assign n13454 = n2244 & ~n13453 ;
  assign n13437 = n5992 & n6012 ;
  assign n13438 = ~\P1_InstAddrPointer_reg[21]/NET0131  & ~n5990 ;
  assign n13439 = ~n5046 & ~n13438 ;
  assign n13440 = ~n13437 & ~n13439 ;
  assign n13441 = n2385 & ~n6013 ;
  assign n13442 = ~n13440 & n13441 ;
  assign n13455 = \P1_PhyAddrPointer_reg[21]/NET0131  & ~n10087 ;
  assign n13456 = ~n13442 & ~n13455 ;
  assign n13457 = ~n13454 & n13456 ;
  assign n13458 = n2432 & ~n13457 ;
  assign n13434 = ~\P1_PhyAddrPointer_reg[21]/NET0131  & ~n12277 ;
  assign n13435 = ~n10125 & ~n13434 ;
  assign n13436 = n10133 & n13435 ;
  assign n13429 = n10136 & ~n12280 ;
  assign n13430 = \P1_PhyAddrPointer_reg[21]/NET0131  & ~n13429 ;
  assign n13431 = ~\P1_PhyAddrPointer_reg[21]/NET0131  & n3148 ;
  assign n13432 = n12276 & n13431 ;
  assign n13433 = \P1_rEIP_reg[21]/NET0131  & n5092 ;
  assign n13459 = ~n13432 & ~n13433 ;
  assign n13460 = ~n13430 & n13459 ;
  assign n13461 = ~n13436 & n13460 ;
  assign n13462 = ~n13458 & n13461 ;
  assign n13463 = \P1_PhyAddrPointer_reg[25]/NET0131  & n2375 ;
  assign n13464 = ~n4486 & ~n7286 ;
  assign n13465 = ~n7237 & ~n13464 ;
  assign n13466 = n4453 & ~n13465 ;
  assign n13467 = n4908 & ~n7283 ;
  assign n13468 = ~n4453 & ~n5958 ;
  assign n13469 = ~n13467 & n13468 ;
  assign n13470 = ~n2375 & ~n13469 ;
  assign n13471 = ~n13466 & n13470 ;
  assign n13472 = ~n13463 & ~n13471 ;
  assign n13473 = n2244 & ~n13472 ;
  assign n13474 = \P1_PhyAddrPointer_reg[25]/NET0131  & ~n10087 ;
  assign n13476 = ~n5045 & ~n6014 ;
  assign n13475 = n5052 & n6013 ;
  assign n13477 = n2385 & ~n13475 ;
  assign n13478 = ~n13476 & n13477 ;
  assign n13479 = ~n13474 & ~n13478 ;
  assign n13480 = ~n13473 & n13479 ;
  assign n13481 = n2432 & ~n13480 ;
  assign n13485 = ~\P1_PhyAddrPointer_reg[25]/NET0131  & ~n12333 ;
  assign n13486 = ~n10126 & ~n13485 ;
  assign n13487 = n10133 & n13486 ;
  assign n13483 = \P1_PhyAddrPointer_reg[25]/NET0131  & ~n12351 ;
  assign n13482 = n12328 & n12350 ;
  assign n13484 = \P1_rEIP_reg[25]/NET0131  & n5092 ;
  assign n13488 = ~n13482 & ~n13484 ;
  assign n13489 = ~n13483 & n13488 ;
  assign n13490 = ~n13487 & n13489 ;
  assign n13491 = ~n13481 & n13490 ;
  assign n13499 = \P1_PhyAddrPointer_reg[8]/NET0131  & n2375 ;
  assign n13501 = ~n4502 & n6825 ;
  assign n13500 = n4502 & ~n6825 ;
  assign n13502 = n4453 & ~n13500 ;
  assign n13503 = ~n13501 & n13502 ;
  assign n13505 = ~n4826 & n6855 ;
  assign n13506 = ~n4869 & ~n13505 ;
  assign n13504 = n4869 & n7271 ;
  assign n13507 = ~n4453 & ~n13504 ;
  assign n13508 = ~n13506 & n13507 ;
  assign n13509 = ~n13503 & ~n13508 ;
  assign n13510 = ~n2375 & ~n13509 ;
  assign n13511 = ~n13499 & ~n13510 ;
  assign n13512 = n2244 & ~n13511 ;
  assign n13496 = ~n4977 & n5018 ;
  assign n13495 = n4977 & ~n5018 ;
  assign n13497 = n2385 & ~n13495 ;
  assign n13498 = ~n13496 & n13497 ;
  assign n13513 = \P1_PhyAddrPointer_reg[8]/NET0131  & ~n10087 ;
  assign n13514 = ~n13498 & ~n13513 ;
  assign n13515 = ~n13512 & n13514 ;
  assign n13516 = n2432 & ~n13515 ;
  assign n13492 = ~\P1_PhyAddrPointer_reg[8]/NET0131  & ~n12150 ;
  assign n13493 = ~n12151 & ~n13492 ;
  assign n13517 = ~\P1_DataWidth_reg[1]/NET0131  & ~n13493 ;
  assign n13518 = ~\P1_PhyAddrPointer_reg[8]/NET0131  & ~n10096 ;
  assign n13519 = ~n10097 & ~n13518 ;
  assign n13520 = \P1_DataWidth_reg[1]/NET0131  & ~n13519 ;
  assign n13521 = n2436 & ~n13520 ;
  assign n13522 = ~n13517 & n13521 ;
  assign n13494 = n5095 & n13493 ;
  assign n13523 = \P1_rEIP_reg[8]/NET0131  & n5092 ;
  assign n13524 = \P1_PhyAddrPointer_reg[8]/NET0131  & ~n10136 ;
  assign n13525 = ~n13523 & ~n13524 ;
  assign n13526 = ~n13494 & n13525 ;
  assign n13527 = ~n13522 & n13526 ;
  assign n13528 = ~n13516 & n13527 ;
  assign n13529 = \P2_PhyAddrPointer_reg[12]/NET0131  & n1897 ;
  assign n13530 = ~n9237 & ~n13529 ;
  assign n13531 = n1734 & ~n13530 ;
  assign n13532 = \P2_PhyAddrPointer_reg[12]/NET0131  & ~n8936 ;
  assign n13533 = ~n9247 & ~n13532 ;
  assign n13534 = ~n13531 & n13533 ;
  assign n13535 = n1927 & ~n13534 ;
  assign n13540 = ~\P2_PhyAddrPointer_reg[12]/NET0131  & ~n12376 ;
  assign n13541 = \P2_PhyAddrPointer_reg[12]/NET0131  & n12376 ;
  assign n13542 = ~n13540 & ~n13541 ;
  assign n13543 = n9005 & n13542 ;
  assign n13537 = ~\P2_PhyAddrPointer_reg[12]/NET0131  & ~n8968 ;
  assign n13536 = \P2_PhyAddrPointer_reg[12]/NET0131  & n8968 ;
  assign n13538 = n3034 & ~n13536 ;
  assign n13539 = ~n13537 & n13538 ;
  assign n13544 = \P2_PhyAddrPointer_reg[12]/NET0131  & ~n8958 ;
  assign n13545 = ~n9223 & ~n13544 ;
  assign n13546 = ~n13539 & n13545 ;
  assign n13547 = ~n13543 & n13546 ;
  assign n13548 = ~n13535 & n13547 ;
  assign n13550 = \P2_PhyAddrPointer_reg[13]/NET0131  & n1897 ;
  assign n13551 = ~n9272 & ~n13550 ;
  assign n13552 = n1734 & ~n13551 ;
  assign n13553 = \P2_PhyAddrPointer_reg[13]/NET0131  & ~n8936 ;
  assign n13554 = ~n9278 & ~n13553 ;
  assign n13555 = ~n13552 & n13554 ;
  assign n13556 = n1927 & ~n13555 ;
  assign n13557 = ~\P2_PhyAddrPointer_reg[13]/NET0131  & ~n13541 ;
  assign n13558 = n8968 & n8969 ;
  assign n13559 = \P2_PhyAddrPointer_reg[1]/NET0131  & n13558 ;
  assign n13560 = ~n13557 & ~n13559 ;
  assign n13561 = n3087 & n13560 ;
  assign n13563 = \P2_PhyAddrPointer_reg[12]/NET0131  & n12370 ;
  assign n13564 = ~\P2_PhyAddrPointer_reg[13]/NET0131  & ~n13563 ;
  assign n13562 = ~n10965 & n13558 ;
  assign n13565 = n1931 & ~n13562 ;
  assign n13566 = ~n13564 & n13565 ;
  assign n13549 = \P2_PhyAddrPointer_reg[13]/NET0131  & ~n8958 ;
  assign n13567 = ~n9261 & ~n13549 ;
  assign n13568 = ~n13566 & n13567 ;
  assign n13569 = ~n13561 & n13568 ;
  assign n13570 = ~n13556 & n13569 ;
  assign n13572 = \P2_PhyAddrPointer_reg[14]/NET0131  & n1897 ;
  assign n13574 = ~n6650 & ~n7457 ;
  assign n13575 = n6188 & ~n7464 ;
  assign n13576 = ~n13574 & n13575 ;
  assign n13573 = n6502 & n9266 ;
  assign n13577 = ~n7436 & ~n13573 ;
  assign n13578 = ~n13576 & n13577 ;
  assign n13579 = ~n1897 & ~n13578 ;
  assign n13580 = ~n13572 & ~n13579 ;
  assign n13581 = n1734 & ~n13580 ;
  assign n13582 = \P2_PhyAddrPointer_reg[14]/NET0131  & ~n8936 ;
  assign n13584 = n6751 & n7547 ;
  assign n13583 = ~n6751 & ~n7547 ;
  assign n13585 = n1890 & ~n13583 ;
  assign n13586 = ~n13584 & n13585 ;
  assign n13587 = ~n13582 & ~n13586 ;
  assign n13588 = ~n13581 & n13587 ;
  assign n13589 = n1927 & ~n13588 ;
  assign n13594 = ~\P2_PhyAddrPointer_reg[14]/NET0131  & ~n13559 ;
  assign n13595 = ~n12384 & ~n13594 ;
  assign n13596 = n9005 & n13595 ;
  assign n13590 = ~\P2_PhyAddrPointer_reg[14]/NET0131  & ~n13558 ;
  assign n13591 = n3034 & ~n8971 ;
  assign n13592 = ~n13590 & n13591 ;
  assign n13571 = \P2_PhyAddrPointer_reg[14]/NET0131  & ~n8958 ;
  assign n13593 = \P2_rEIP_reg[14]/NET0131  & n3113 ;
  assign n13597 = ~n13571 & ~n13593 ;
  assign n13598 = ~n13592 & n13597 ;
  assign n13599 = ~n13596 & n13598 ;
  assign n13600 = ~n13589 & n13599 ;
  assign n13602 = \P2_PhyAddrPointer_reg[16]/NET0131  & n1897 ;
  assign n13606 = ~\P2_InstAddrPointer_reg[16]/NET0131  & ~n7460 ;
  assign n13607 = ~n6657 & ~n13606 ;
  assign n13609 = ~n7458 & n13607 ;
  assign n13608 = n7458 & ~n13607 ;
  assign n13610 = n6188 & ~n13608 ;
  assign n13611 = ~n13609 & n13610 ;
  assign n13603 = n6515 & ~n11021 ;
  assign n13604 = ~n6188 & ~n7516 ;
  assign n13605 = ~n13603 & n13604 ;
  assign n13612 = ~n1897 & ~n13605 ;
  assign n13613 = ~n13611 & n13612 ;
  assign n13614 = ~n13602 & ~n13613 ;
  assign n13615 = n1734 & ~n13614 ;
  assign n13616 = \P2_PhyAddrPointer_reg[16]/NET0131  & ~n8936 ;
  assign n13617 = ~n11039 & ~n11041 ;
  assign n13618 = n1890 & ~n11042 ;
  assign n13619 = ~n13617 & n13618 ;
  assign n13620 = ~n13616 & ~n13619 ;
  assign n13621 = ~n13615 & n13620 ;
  assign n13622 = n1927 & ~n13621 ;
  assign n13623 = \P2_PhyAddrPointer_reg[16]/NET0131  & n8972 ;
  assign n13624 = ~\P2_PhyAddrPointer_reg[16]/NET0131  & ~n8972 ;
  assign n13625 = ~n13623 & ~n13624 ;
  assign n13626 = \P2_PhyAddrPointer_reg[1]/NET0131  & ~n13625 ;
  assign n13627 = ~\P2_PhyAddrPointer_reg[16]/NET0131  & ~\P2_PhyAddrPointer_reg[1]/NET0131  ;
  assign n13628 = ~n13626 & ~n13627 ;
  assign n13629 = n9005 & n13628 ;
  assign n13630 = n3034 & n13625 ;
  assign n13601 = \P2_rEIP_reg[16]/NET0131  & n3113 ;
  assign n13631 = \P2_PhyAddrPointer_reg[16]/NET0131  & ~n8958 ;
  assign n13632 = ~n13601 & ~n13631 ;
  assign n13633 = ~n13630 & n13632 ;
  assign n13634 = ~n13629 & n13633 ;
  assign n13635 = ~n13622 & n13634 ;
  assign n13636 = \P2_PhyAddrPointer_reg[17]/NET0131  & n1897 ;
  assign n13641 = ~n6656 & ~n6660 ;
  assign n13642 = n6656 & n6660 ;
  assign n13643 = ~n13641 & ~n13642 ;
  assign n13644 = n6188 & ~n13643 ;
  assign n13637 = ~n6520 & ~n6524 ;
  assign n13638 = n6520 & n6524 ;
  assign n13639 = ~n13637 & ~n13638 ;
  assign n13640 = ~n6188 & ~n13639 ;
  assign n13645 = ~n1897 & ~n13640 ;
  assign n13646 = ~n13644 & n13645 ;
  assign n13647 = ~n13636 & ~n13646 ;
  assign n13648 = n1734 & ~n13647 ;
  assign n13649 = \P2_PhyAddrPointer_reg[17]/NET0131  & ~n8936 ;
  assign n13650 = n6746 & n6752 ;
  assign n13652 = n6757 & n13650 ;
  assign n13651 = ~n6757 & ~n13650 ;
  assign n13653 = n1890 & ~n13651 ;
  assign n13654 = ~n13652 & n13653 ;
  assign n13655 = ~n13649 & ~n13654 ;
  assign n13656 = ~n13648 & n13655 ;
  assign n13657 = n1927 & ~n13656 ;
  assign n13662 = \P2_PhyAddrPointer_reg[16]/NET0131  & n12386 ;
  assign n13663 = ~\P2_PhyAddrPointer_reg[17]/NET0131  & ~n13662 ;
  assign n13664 = \P2_PhyAddrPointer_reg[17]/NET0131  & n13662 ;
  assign n13665 = ~n13663 & ~n13664 ;
  assign n13666 = n9005 & n13665 ;
  assign n13659 = ~\P2_PhyAddrPointer_reg[17]/NET0131  & ~n13623 ;
  assign n13658 = \P2_PhyAddrPointer_reg[17]/NET0131  & n13623 ;
  assign n13660 = n3034 & ~n13658 ;
  assign n13661 = ~n13659 & n13660 ;
  assign n13667 = \P2_PhyAddrPointer_reg[17]/NET0131  & ~n8958 ;
  assign n13668 = \P2_rEIP_reg[17]/NET0131  & n3113 ;
  assign n13669 = ~n13667 & ~n13668 ;
  assign n13670 = ~n13661 & n13669 ;
  assign n13671 = ~n13666 & n13670 ;
  assign n13672 = ~n13657 & n13671 ;
  assign n13676 = \P2_PhyAddrPointer_reg[18]/NET0131  & n1897 ;
  assign n13677 = ~n8480 & ~n13676 ;
  assign n13678 = n1734 & ~n13677 ;
  assign n13679 = \P2_PhyAddrPointer_reg[18]/NET0131  & ~n8936 ;
  assign n13680 = ~n8485 & ~n13679 ;
  assign n13681 = ~n13678 & n13680 ;
  assign n13682 = n1927 & ~n13681 ;
  assign n13673 = ~\P2_PhyAddrPointer_reg[18]/NET0131  & ~n13664 ;
  assign n13674 = ~n12427 & ~n13673 ;
  assign n13683 = ~\P2_DataWidth_reg[1]/NET0131  & ~n13674 ;
  assign n13684 = ~\P2_PhyAddrPointer_reg[18]/NET0131  & ~n13658 ;
  assign n13685 = ~n8975 & ~n13684 ;
  assign n13686 = \P2_DataWidth_reg[1]/NET0131  & ~n13685 ;
  assign n13687 = n1931 & ~n13686 ;
  assign n13688 = ~n13683 & n13687 ;
  assign n13675 = n3087 & n13674 ;
  assign n13689 = \P2_PhyAddrPointer_reg[18]/NET0131  & ~n8958 ;
  assign n13690 = ~n8502 & ~n13689 ;
  assign n13691 = ~n13675 & n13690 ;
  assign n13692 = ~n13688 & n13691 ;
  assign n13693 = ~n13682 & n13692 ;
  assign n13716 = ~\P1_InstAddrPointer_reg[1]/NET0131  & ~n2314 ;
  assign n13717 = n9315 & ~n13716 ;
  assign n13718 = \P1_InstAddrPointer_reg[2]/NET0131  & ~n13717 ;
  assign n13719 = ~n2402 & n4677 ;
  assign n13715 = ~n2271 & n4849 ;
  assign n13702 = ~n4850 & n5946 ;
  assign n13700 = ~n4850 & ~n4854 ;
  assign n13701 = n4844 & ~n13700 ;
  assign n13703 = ~n4453 & ~n13701 ;
  assign n13704 = ~n13702 & n13703 ;
  assign n13705 = ~n4678 & ~n4679 ;
  assign n13707 = n4746 & n13705 ;
  assign n13706 = ~n4746 & ~n13705 ;
  assign n13708 = n4453 & ~n13706 ;
  assign n13709 = ~n13707 & n13708 ;
  assign n13710 = ~n13704 & ~n13709 ;
  assign n13711 = ~n2375 & ~n13710 ;
  assign n13712 = ~\P1_InstAddrPointer_reg[2]/NET0131  & n2375 ;
  assign n13713 = n2244 & ~n13712 ;
  assign n13714 = ~n13711 & n13713 ;
  assign n13696 = ~\P1_InstAddrPointer_reg[2]/NET0131  & ~n2337 ;
  assign n13697 = n2337 & n4849 ;
  assign n13698 = ~n13696 & ~n13697 ;
  assign n13699 = ~n2332 & n13698 ;
  assign n13721 = ~n4999 & n13700 ;
  assign n13720 = n4999 & ~n13700 ;
  assign n13722 = n2385 & ~n13720 ;
  assign n13723 = ~n13721 & n13722 ;
  assign n13724 = ~n13699 & ~n13723 ;
  assign n13725 = ~n13714 & n13724 ;
  assign n13726 = ~n13715 & n13725 ;
  assign n13727 = ~n13719 & n13726 ;
  assign n13728 = ~n13718 & n13727 ;
  assign n13729 = n2432 & ~n13728 ;
  assign n13694 = \P1_rEIP_reg[2]/NET0131  & n5092 ;
  assign n13695 = \P1_InstAddrPointer_reg[2]/NET0131  & ~n5098 ;
  assign n13730 = ~n13694 & ~n13695 ;
  assign n13731 = ~n13729 & n13730 ;
  assign n13735 = \P3_InstAddrPointer_reg[2]/NET0131  & ~n11451 ;
  assign n13744 = ~n2777 & n4189 ;
  assign n13734 = ~n2923 & n3898 ;
  assign n13736 = ~n4190 & ~n4194 ;
  assign n13737 = n4328 & n13736 ;
  assign n13738 = ~n4328 & ~n13736 ;
  assign n13739 = ~n13737 & ~n13738 ;
  assign n13740 = n2899 & n13739 ;
  assign n13741 = ~n2841 & ~n4189 ;
  assign n13742 = ~n13740 & ~n13741 ;
  assign n13743 = n2847 & ~n13742 ;
  assign n13751 = n4192 & n13736 ;
  assign n13750 = ~n4192 & ~n13736 ;
  assign n13752 = ~n3753 & ~n13750 ;
  assign n13753 = ~n13751 & n13752 ;
  assign n13745 = ~n3899 & ~n4036 ;
  assign n13747 = n3966 & n13745 ;
  assign n13746 = ~n3966 & ~n13745 ;
  assign n13748 = n3753 & ~n13746 ;
  assign n13749 = ~n13747 & n13748 ;
  assign n13754 = n2904 & ~n13749 ;
  assign n13755 = ~n13753 & n13754 ;
  assign n13756 = ~n13743 & ~n13755 ;
  assign n13757 = ~n13734 & n13756 ;
  assign n13758 = ~n13744 & n13757 ;
  assign n13759 = ~n13735 & n13758 ;
  assign n13760 = n2453 & ~n13759 ;
  assign n13732 = \P3_rEIP_reg[2]/NET0131  & n4412 ;
  assign n13733 = \P3_InstAddrPointer_reg[2]/NET0131  & ~n4418 ;
  assign n13761 = ~n13732 & ~n13733 ;
  assign n13762 = ~n13760 & n13761 ;
  assign n13781 = \P2_InstAddrPointer_reg[2]/NET0131  & ~n7500 ;
  assign n13767 = ~n6302 & ~n6441 ;
  assign n13793 = ~n6717 & n13767 ;
  assign n13794 = n6717 & ~n13767 ;
  assign n13795 = ~n13793 & ~n13794 ;
  assign n13796 = n1732 & n13795 ;
  assign n13797 = ~n1727 & ~n6301 ;
  assign n13798 = ~n13796 & ~n13797 ;
  assign n13799 = n1798 & ~n13798 ;
  assign n13765 = n1739 & n6611 ;
  assign n13783 = ~\P2_InstAddrPointer_reg[2]/NET0131  & n1805 ;
  assign n13784 = ~n1805 & ~n6611 ;
  assign n13785 = ~n13783 & ~n13784 ;
  assign n13786 = ~n1804 & n13785 ;
  assign n13787 = ~\P2_InstAddrPointer_reg[2]/NET0131  & ~n1820 ;
  assign n13788 = n1820 & ~n6611 ;
  assign n13789 = ~n13787 & ~n13788 ;
  assign n13790 = ~n1814 & n13789 ;
  assign n13791 = ~n13786 & ~n13790 ;
  assign n13792 = ~n1810 & ~n13791 ;
  assign n13800 = ~n13765 & ~n13792 ;
  assign n13801 = ~n13799 & n13800 ;
  assign n13802 = ~n13781 & n13801 ;
  assign n13766 = \P2_InstAddrPointer_reg[2]/NET0131  & n1897 ;
  assign n13772 = ~n6612 & ~n6624 ;
  assign n13773 = n6616 & ~n13772 ;
  assign n13774 = ~n6616 & n13772 ;
  assign n13775 = ~n13773 & ~n13774 ;
  assign n13776 = n6188 & ~n13775 ;
  assign n13769 = n6371 & ~n13767 ;
  assign n13768 = ~n6371 & n13767 ;
  assign n13770 = ~n6188 & ~n13768 ;
  assign n13771 = ~n13769 & n13770 ;
  assign n13777 = ~n1897 & ~n13771 ;
  assign n13778 = ~n13776 & n13777 ;
  assign n13779 = ~n13766 & ~n13778 ;
  assign n13780 = n1734 & ~n13779 ;
  assign n13782 = ~n1771 & n6301 ;
  assign n13803 = ~n13780 & ~n13782 ;
  assign n13804 = n13802 & n13803 ;
  assign n13805 = n1927 & ~n13804 ;
  assign n13763 = \P2_rEIP_reg[2]/NET0131  & n3113 ;
  assign n13764 = \P2_InstAddrPointer_reg[2]/NET0131  & ~n6810 ;
  assign n13806 = ~n13763 & ~n13764 ;
  assign n13807 = ~n13805 & n13806 ;
  assign n13808 = ~n2993 & ~n2997 ;
  assign n13809 = ~n2951 & ~n2953 ;
  assign n13810 = n13808 & n13809 ;
  assign n13811 = \P3_EAX_reg[27]/NET0131  & ~n13810 ;
  assign n14017 = \P3_EAX_reg[0]/NET0131  & \P3_EAX_reg[1]/NET0131  ;
  assign n14018 = \P3_EAX_reg[2]/NET0131  & n14017 ;
  assign n14019 = \P3_EAX_reg[3]/NET0131  & n14018 ;
  assign n14020 = \P3_EAX_reg[4]/NET0131  & n14019 ;
  assign n14021 = \P3_EAX_reg[5]/NET0131  & n14020 ;
  assign n14022 = \P3_EAX_reg[6]/NET0131  & n14021 ;
  assign n14023 = \P3_EAX_reg[7]/NET0131  & n14022 ;
  assign n14024 = \P3_EAX_reg[8]/NET0131  & n14023 ;
  assign n14025 = \P3_EAX_reg[9]/NET0131  & n14024 ;
  assign n14026 = \P3_EAX_reg[10]/NET0131  & n14025 ;
  assign n14027 = \P3_EAX_reg[11]/NET0131  & n14026 ;
  assign n14028 = \P3_EAX_reg[12]/NET0131  & n14027 ;
  assign n14029 = \P3_EAX_reg[13]/NET0131  & n14028 ;
  assign n14030 = \P3_EAX_reg[14]/NET0131  & n14029 ;
  assign n14031 = \P3_EAX_reg[15]/NET0131  & n14030 ;
  assign n14032 = \P3_EAX_reg[16]/NET0131  & \P3_EAX_reg[17]/NET0131  ;
  assign n14033 = \P3_EAX_reg[18]/NET0131  & n14032 ;
  assign n14034 = n14031 & n14033 ;
  assign n14035 = \P3_EAX_reg[19]/NET0131  & n14034 ;
  assign n14036 = \P3_EAX_reg[20]/NET0131  & n14035 ;
  assign n14037 = \P3_EAX_reg[21]/NET0131  & n14036 ;
  assign n14038 = \P3_EAX_reg[22]/NET0131  & \P3_EAX_reg[23]/NET0131  ;
  assign n14039 = \P3_EAX_reg[24]/NET0131  & n14038 ;
  assign n14040 = \P3_EAX_reg[25]/NET0131  & n14039 ;
  assign n14041 = n14037 & n14040 ;
  assign n14042 = \P3_EAX_reg[26]/NET0131  & n14041 ;
  assign n14043 = ~\P3_EAX_reg[27]/NET0131  & ~n14042 ;
  assign n13813 = n2740 & n2742 ;
  assign n14044 = \P3_EAX_reg[26]/NET0131  & \P3_EAX_reg[27]/NET0131  ;
  assign n14045 = n14041 & n14044 ;
  assign n14046 = n13813 & ~n14045 ;
  assign n14047 = ~n14043 & n14046 ;
  assign n13812 = n2840 & n2847 ;
  assign n13814 = n2822 & ~n13813 ;
  assign n13815 = ~n2840 & ~n13814 ;
  assign n13816 = ~n13812 & ~n13815 ;
  assign n13817 = ~n2863 & ~n13816 ;
  assign n13818 = \P3_EAX_reg[27]/NET0131  & ~n13817 ;
  assign n14014 = ~\buf2_reg[27]/NET0131  & n2862 ;
  assign n14013 = ~\P3_EAX_reg[27]/NET0131  & ~n2862 ;
  assign n14015 = n2820 & ~n14013 ;
  assign n14016 = ~n14014 & n14015 ;
  assign n13823 = \P3_InstQueue_reg[14][0]/NET0131  & n2464 ;
  assign n13824 = \P3_InstQueue_reg[0][0]/NET0131  & n2472 ;
  assign n13837 = ~n13823 & ~n13824 ;
  assign n13825 = \P3_InstQueue_reg[13][0]/NET0131  & n2490 ;
  assign n13826 = \P3_InstQueue_reg[10][0]/NET0131  & n2474 ;
  assign n13838 = ~n13825 & ~n13826 ;
  assign n13845 = n13837 & n13838 ;
  assign n13819 = \P3_InstQueue_reg[4][0]/NET0131  & n2482 ;
  assign n13820 = \P3_InstQueue_reg[9][0]/NET0131  & n2492 ;
  assign n13835 = ~n13819 & ~n13820 ;
  assign n13821 = \P3_InstQueue_reg[3][0]/NET0131  & n2484 ;
  assign n13822 = \P3_InstQueue_reg[6][0]/NET0131  & n2466 ;
  assign n13836 = ~n13821 & ~n13822 ;
  assign n13846 = n13835 & n13836 ;
  assign n13847 = n13845 & n13846 ;
  assign n13831 = \P3_InstQueue_reg[1][0]/NET0131  & n2478 ;
  assign n13832 = \P3_InstQueue_reg[7][0]/NET0131  & n2480 ;
  assign n13841 = ~n13831 & ~n13832 ;
  assign n13833 = \P3_InstQueue_reg[11][0]/NET0131  & n2460 ;
  assign n13834 = \P3_InstQueue_reg[12][0]/NET0131  & n2476 ;
  assign n13842 = ~n13833 & ~n13834 ;
  assign n13843 = n13841 & n13842 ;
  assign n13827 = \P3_InstQueue_reg[15][0]/NET0131  & n2486 ;
  assign n13828 = \P3_InstQueue_reg[8][0]/NET0131  & n2469 ;
  assign n13839 = ~n13827 & ~n13828 ;
  assign n13829 = \P3_InstQueue_reg[5][0]/NET0131  & n2456 ;
  assign n13830 = \P3_InstQueue_reg[2][0]/NET0131  & n2488 ;
  assign n13840 = ~n13829 & ~n13830 ;
  assign n13844 = n13839 & n13840 ;
  assign n13848 = n13843 & n13844 ;
  assign n13849 = n13847 & n13848 ;
  assign n13854 = \P3_InstQueue_reg[5][7]/NET0131  & n2466 ;
  assign n13855 = \P3_InstQueue_reg[0][7]/NET0131  & n2478 ;
  assign n13868 = ~n13854 & ~n13855 ;
  assign n13856 = \P3_InstQueue_reg[7][7]/NET0131  & n2469 ;
  assign n13857 = \P3_InstQueue_reg[10][7]/NET0131  & n2460 ;
  assign n13869 = ~n13856 & ~n13857 ;
  assign n13876 = n13868 & n13869 ;
  assign n13850 = \P3_InstQueue_reg[15][7]/NET0131  & n2472 ;
  assign n13851 = \P3_InstQueue_reg[9][7]/NET0131  & n2474 ;
  assign n13866 = ~n13850 & ~n13851 ;
  assign n13852 = \P3_InstQueue_reg[11][7]/NET0131  & n2476 ;
  assign n13853 = \P3_InstQueue_reg[13][7]/NET0131  & n2464 ;
  assign n13867 = ~n13852 & ~n13853 ;
  assign n13877 = n13866 & n13867 ;
  assign n13878 = n13876 & n13877 ;
  assign n13862 = \P3_InstQueue_reg[4][7]/NET0131  & n2456 ;
  assign n13863 = \P3_InstQueue_reg[6][7]/NET0131  & n2480 ;
  assign n13872 = ~n13862 & ~n13863 ;
  assign n13864 = \P3_InstQueue_reg[3][7]/NET0131  & n2482 ;
  assign n13865 = \P3_InstQueue_reg[2][7]/NET0131  & n2484 ;
  assign n13873 = ~n13864 & ~n13865 ;
  assign n13874 = n13872 & n13873 ;
  assign n13858 = \P3_InstQueue_reg[12][7]/NET0131  & n2490 ;
  assign n13859 = \P3_InstQueue_reg[8][7]/NET0131  & n2492 ;
  assign n13870 = ~n13858 & ~n13859 ;
  assign n13860 = \P3_InstQueue_reg[14][7]/NET0131  & n2486 ;
  assign n13861 = \P3_InstQueue_reg[1][7]/NET0131  & n2488 ;
  assign n13871 = ~n13860 & ~n13861 ;
  assign n13875 = n13870 & n13871 ;
  assign n13879 = n13874 & n13875 ;
  assign n13880 = n13878 & n13879 ;
  assign n13881 = ~n13849 & ~n13880 ;
  assign n13886 = \P3_InstQueue_reg[14][1]/NET0131  & n2464 ;
  assign n13887 = \P3_InstQueue_reg[0][1]/NET0131  & n2472 ;
  assign n13900 = ~n13886 & ~n13887 ;
  assign n13888 = \P3_InstQueue_reg[13][1]/NET0131  & n2490 ;
  assign n13889 = \P3_InstQueue_reg[10][1]/NET0131  & n2474 ;
  assign n13901 = ~n13888 & ~n13889 ;
  assign n13908 = n13900 & n13901 ;
  assign n13882 = \P3_InstQueue_reg[4][1]/NET0131  & n2482 ;
  assign n13883 = \P3_InstQueue_reg[9][1]/NET0131  & n2492 ;
  assign n13898 = ~n13882 & ~n13883 ;
  assign n13884 = \P3_InstQueue_reg[3][1]/NET0131  & n2484 ;
  assign n13885 = \P3_InstQueue_reg[6][1]/NET0131  & n2466 ;
  assign n13899 = ~n13884 & ~n13885 ;
  assign n13909 = n13898 & n13899 ;
  assign n13910 = n13908 & n13909 ;
  assign n13894 = \P3_InstQueue_reg[1][1]/NET0131  & n2478 ;
  assign n13895 = \P3_InstQueue_reg[7][1]/NET0131  & n2480 ;
  assign n13904 = ~n13894 & ~n13895 ;
  assign n13896 = \P3_InstQueue_reg[11][1]/NET0131  & n2460 ;
  assign n13897 = \P3_InstQueue_reg[12][1]/NET0131  & n2476 ;
  assign n13905 = ~n13896 & ~n13897 ;
  assign n13906 = n13904 & n13905 ;
  assign n13890 = \P3_InstQueue_reg[15][1]/NET0131  & n2486 ;
  assign n13891 = \P3_InstQueue_reg[8][1]/NET0131  & n2469 ;
  assign n13902 = ~n13890 & ~n13891 ;
  assign n13892 = \P3_InstQueue_reg[5][1]/NET0131  & n2456 ;
  assign n13893 = \P3_InstQueue_reg[2][1]/NET0131  & n2488 ;
  assign n13903 = ~n13892 & ~n13893 ;
  assign n13907 = n13902 & n13903 ;
  assign n13911 = n13906 & n13907 ;
  assign n13912 = n13910 & n13911 ;
  assign n13913 = n13881 & ~n13912 ;
  assign n13918 = \P3_InstQueue_reg[14][2]/NET0131  & n2464 ;
  assign n13919 = \P3_InstQueue_reg[0][2]/NET0131  & n2472 ;
  assign n13932 = ~n13918 & ~n13919 ;
  assign n13920 = \P3_InstQueue_reg[13][2]/NET0131  & n2490 ;
  assign n13921 = \P3_InstQueue_reg[10][2]/NET0131  & n2474 ;
  assign n13933 = ~n13920 & ~n13921 ;
  assign n13940 = n13932 & n13933 ;
  assign n13914 = \P3_InstQueue_reg[4][2]/NET0131  & n2482 ;
  assign n13915 = \P3_InstQueue_reg[9][2]/NET0131  & n2492 ;
  assign n13930 = ~n13914 & ~n13915 ;
  assign n13916 = \P3_InstQueue_reg[3][2]/NET0131  & n2484 ;
  assign n13917 = \P3_InstQueue_reg[6][2]/NET0131  & n2466 ;
  assign n13931 = ~n13916 & ~n13917 ;
  assign n13941 = n13930 & n13931 ;
  assign n13942 = n13940 & n13941 ;
  assign n13926 = \P3_InstQueue_reg[1][2]/NET0131  & n2478 ;
  assign n13927 = \P3_InstQueue_reg[7][2]/NET0131  & n2480 ;
  assign n13936 = ~n13926 & ~n13927 ;
  assign n13928 = \P3_InstQueue_reg[11][2]/NET0131  & n2460 ;
  assign n13929 = \P3_InstQueue_reg[12][2]/NET0131  & n2476 ;
  assign n13937 = ~n13928 & ~n13929 ;
  assign n13938 = n13936 & n13937 ;
  assign n13922 = \P3_InstQueue_reg[15][2]/NET0131  & n2486 ;
  assign n13923 = \P3_InstQueue_reg[8][2]/NET0131  & n2469 ;
  assign n13934 = ~n13922 & ~n13923 ;
  assign n13924 = \P3_InstQueue_reg[5][2]/NET0131  & n2456 ;
  assign n13925 = \P3_InstQueue_reg[2][2]/NET0131  & n2488 ;
  assign n13935 = ~n13924 & ~n13925 ;
  assign n13939 = n13934 & n13935 ;
  assign n13943 = n13938 & n13939 ;
  assign n13944 = n13942 & n13943 ;
  assign n13945 = n13913 & ~n13944 ;
  assign n13950 = \P3_InstQueue_reg[14][3]/NET0131  & n2464 ;
  assign n13951 = \P3_InstQueue_reg[0][3]/NET0131  & n2472 ;
  assign n13964 = ~n13950 & ~n13951 ;
  assign n13952 = \P3_InstQueue_reg[13][3]/NET0131  & n2490 ;
  assign n13953 = \P3_InstQueue_reg[10][3]/NET0131  & n2474 ;
  assign n13965 = ~n13952 & ~n13953 ;
  assign n13972 = n13964 & n13965 ;
  assign n13946 = \P3_InstQueue_reg[4][3]/NET0131  & n2482 ;
  assign n13947 = \P3_InstQueue_reg[9][3]/NET0131  & n2492 ;
  assign n13962 = ~n13946 & ~n13947 ;
  assign n13948 = \P3_InstQueue_reg[3][3]/NET0131  & n2484 ;
  assign n13949 = \P3_InstQueue_reg[6][3]/NET0131  & n2466 ;
  assign n13963 = ~n13948 & ~n13949 ;
  assign n13973 = n13962 & n13963 ;
  assign n13974 = n13972 & n13973 ;
  assign n13958 = \P3_InstQueue_reg[1][3]/NET0131  & n2478 ;
  assign n13959 = \P3_InstQueue_reg[7][3]/NET0131  & n2480 ;
  assign n13968 = ~n13958 & ~n13959 ;
  assign n13960 = \P3_InstQueue_reg[11][3]/NET0131  & n2460 ;
  assign n13961 = \P3_InstQueue_reg[12][3]/NET0131  & n2476 ;
  assign n13969 = ~n13960 & ~n13961 ;
  assign n13970 = n13968 & n13969 ;
  assign n13954 = \P3_InstQueue_reg[15][3]/NET0131  & n2486 ;
  assign n13955 = \P3_InstQueue_reg[8][3]/NET0131  & n2469 ;
  assign n13966 = ~n13954 & ~n13955 ;
  assign n13956 = \P3_InstQueue_reg[5][3]/NET0131  & n2456 ;
  assign n13957 = \P3_InstQueue_reg[2][3]/NET0131  & n2488 ;
  assign n13967 = ~n13956 & ~n13957 ;
  assign n13971 = n13966 & n13967 ;
  assign n13975 = n13970 & n13971 ;
  assign n13976 = n13974 & n13975 ;
  assign n13977 = n13945 & ~n13976 ;
  assign n13982 = \P3_InstQueue_reg[14][4]/NET0131  & n2464 ;
  assign n13983 = \P3_InstQueue_reg[0][4]/NET0131  & n2472 ;
  assign n13996 = ~n13982 & ~n13983 ;
  assign n13984 = \P3_InstQueue_reg[13][4]/NET0131  & n2490 ;
  assign n13985 = \P3_InstQueue_reg[10][4]/NET0131  & n2474 ;
  assign n13997 = ~n13984 & ~n13985 ;
  assign n14004 = n13996 & n13997 ;
  assign n13978 = \P3_InstQueue_reg[4][4]/NET0131  & n2482 ;
  assign n13979 = \P3_InstQueue_reg[9][4]/NET0131  & n2492 ;
  assign n13994 = ~n13978 & ~n13979 ;
  assign n13980 = \P3_InstQueue_reg[3][4]/NET0131  & n2484 ;
  assign n13981 = \P3_InstQueue_reg[6][4]/NET0131  & n2466 ;
  assign n13995 = ~n13980 & ~n13981 ;
  assign n14005 = n13994 & n13995 ;
  assign n14006 = n14004 & n14005 ;
  assign n13990 = \P3_InstQueue_reg[1][4]/NET0131  & n2478 ;
  assign n13991 = \P3_InstQueue_reg[7][4]/NET0131  & n2480 ;
  assign n14000 = ~n13990 & ~n13991 ;
  assign n13992 = \P3_InstQueue_reg[11][4]/NET0131  & n2460 ;
  assign n13993 = \P3_InstQueue_reg[12][4]/NET0131  & n2476 ;
  assign n14001 = ~n13992 & ~n13993 ;
  assign n14002 = n14000 & n14001 ;
  assign n13986 = \P3_InstQueue_reg[15][4]/NET0131  & n2486 ;
  assign n13987 = \P3_InstQueue_reg[8][4]/NET0131  & n2469 ;
  assign n13998 = ~n13986 & ~n13987 ;
  assign n13988 = \P3_InstQueue_reg[5][4]/NET0131  & n2456 ;
  assign n13989 = \P3_InstQueue_reg[2][4]/NET0131  & n2488 ;
  assign n13999 = ~n13988 & ~n13989 ;
  assign n14003 = n13998 & n13999 ;
  assign n14007 = n14002 & n14003 ;
  assign n14008 = n14006 & n14007 ;
  assign n14009 = ~n13977 & n14008 ;
  assign n14010 = n13977 & ~n14008 ;
  assign n14011 = ~n14009 & ~n14010 ;
  assign n14012 = n13812 & n14011 ;
  assign n14048 = \buf2_reg[11]/NET0131  & n2862 ;
  assign n14049 = n2821 & n14048 ;
  assign n14050 = ~n14012 & ~n14049 ;
  assign n14051 = ~n14016 & n14050 ;
  assign n14052 = ~n13818 & n14051 ;
  assign n14053 = ~n14047 & n14052 ;
  assign n14054 = n2453 & ~n14053 ;
  assign n14055 = ~n13811 & ~n14054 ;
  assign n14056 = \P2_EAX_reg[27]/NET0131  & ~n12632 ;
  assign n14057 = \P2_EAX_reg[26]/NET0131  & n12658 ;
  assign n14058 = n12664 & ~n14057 ;
  assign n14059 = n12669 & ~n14058 ;
  assign n14060 = \P2_EAX_reg[27]/NET0131  & ~n14059 ;
  assign n14061 = ~\P2_EAX_reg[27]/NET0131  & n12664 ;
  assign n14062 = n14057 & n14061 ;
  assign n14063 = ~n12832 & n12863 ;
  assign n14064 = n1798 & ~n12864 ;
  assign n14065 = ~n14063 & n14064 ;
  assign n14066 = n1726 & n14065 ;
  assign n14067 = \buf2_reg[11]/NET0131  & ~n3079 ;
  assign n14068 = \buf1_reg[11]/NET0131  & n3079 ;
  assign n14069 = ~n14067 & ~n14068 ;
  assign n14070 = n1742 & ~n14069 ;
  assign n14071 = n1803 & ~n5306 ;
  assign n14072 = ~n14070 & ~n14071 ;
  assign n14073 = n1811 & ~n14072 ;
  assign n14074 = ~n14066 & ~n14073 ;
  assign n14075 = ~n14062 & n14074 ;
  assign n14076 = ~n14060 & n14075 ;
  assign n14077 = n1927 & ~n14076 ;
  assign n14078 = ~n14056 & ~n14077 ;
  assign n14080 = n2414 & n2432 ;
  assign n14081 = ~n2445 & ~n3017 ;
  assign n14082 = ~n3026 & ~n14081 ;
  assign n14083 = ~n2446 & ~n5092 ;
  assign n14084 = ~n3028 & n14083 ;
  assign n14085 = ~n14082 & n14084 ;
  assign n14086 = \P1_InstQueueRd_Addr_reg[0]/NET0131  & ~n14085 ;
  assign n14079 = ~\P1_InstQueueRd_Addr_reg[0]/NET0131  & n3042 ;
  assign n14087 = \P1_Flush_reg/NET0131  & \P1_InstAddrPointer_reg[0]/NET0131  ;
  assign n14088 = ~\P1_Flush_reg/NET0131  & ~\P1_InstQueueRd_Addr_reg[0]/NET0131  ;
  assign n14089 = ~n14087 & ~n14088 ;
  assign n14090 = n3020 & n14089 ;
  assign n14091 = ~n14079 & ~n14090 ;
  assign n14092 = ~n14086 & n14091 ;
  assign n14093 = ~n14080 & n14092 ;
  assign n14094 = ~n5108 & ~n5185 ;
  assign n14095 = \P1_InstQueue_reg[11][1]/NET0131  & ~n5104 ;
  assign n14096 = ~n5107 & n14095 ;
  assign n14097 = ~n14094 & ~n14096 ;
  assign n14098 = ~n7697 & ~n14097 ;
  assign n14099 = ~n7703 & ~n14098 ;
  assign n14104 = ~n5252 & n5255 ;
  assign n14105 = ~n5256 & ~n14104 ;
  assign n14106 = n5148 & n14105 ;
  assign n14100 = n5236 & ~n5273 ;
  assign n14101 = ~n5274 & ~n14100 ;
  assign n14102 = ~n5148 & n14101 ;
  assign n14103 = n5095 & ~n14097 ;
  assign n14107 = n5153 & ~n14103 ;
  assign n14108 = ~n14102 & n14107 ;
  assign n14109 = ~n14106 & n14108 ;
  assign n14110 = ~n14099 & ~n14109 ;
  assign n14111 = \P1_InstQueue_reg[11][1]/NET0131  & ~n5291 ;
  assign n14112 = ~n2029 & n5104 ;
  assign n14113 = ~n14095 & ~n14112 ;
  assign n14114 = n3042 & ~n14113 ;
  assign n14115 = ~n14111 & ~n14114 ;
  assign n14116 = ~n14110 & n14115 ;
  assign n14118 = n2453 & n2935 ;
  assign n14119 = ~n2962 & ~n4412 ;
  assign n14120 = ~n2952 & ~n2958 ;
  assign n14121 = n14119 & n14120 ;
  assign n14122 = \P3_InstQueueRd_Addr_reg[0]/NET0131  & ~n14121 ;
  assign n14117 = ~\P3_InstQueueRd_Addr_reg[0]/NET0131  & n2994 ;
  assign n14123 = \P3_Flush_reg/NET0131  & \P3_InstAddrPointer_reg[0]/NET0131  ;
  assign n14124 = ~\P3_Flush_reg/NET0131  & ~\P3_InstQueueRd_Addr_reg[0]/NET0131  ;
  assign n14125 = ~n14123 & ~n14124 ;
  assign n14126 = n2997 & n14125 ;
  assign n14127 = ~n14117 & ~n14126 ;
  assign n14128 = ~n14122 & n14127 ;
  assign n14129 = ~n14118 & n14128 ;
  assign n14131 = n1911 & n1927 ;
  assign n14132 = ~n1930 & ~n1936 ;
  assign n14133 = n3115 & n14132 ;
  assign n14134 = \P2_InstQueueRd_Addr_reg[0]/NET0131  & ~n14133 ;
  assign n14130 = ~\P2_InstQueueRd_Addr_reg[0]/NET0131  & n3040 ;
  assign n14135 = \P2_Flush_reg/NET0131  & \P2_InstAddrPointer_reg[0]/NET0131  ;
  assign n14136 = ~\P2_Flush_reg/NET0131  & ~\P2_InstQueueRd_Addr_reg[0]/NET0131  ;
  assign n14137 = ~n14135 & ~n14136 ;
  assign n14138 = n2980 & n14137 ;
  assign n14139 = ~n14130 & ~n14138 ;
  assign n14140 = ~n14134 & n14139 ;
  assign n14141 = ~n14131 & n14140 ;
  assign n14142 = ~n5185 & ~n5327 ;
  assign n14143 = \P1_InstQueue_reg[0][1]/NET0131  & ~n5324 ;
  assign n14144 = ~n5326 & n14143 ;
  assign n14145 = ~n14142 & ~n14144 ;
  assign n14146 = ~n7697 & ~n14145 ;
  assign n14147 = ~n7755 & ~n14146 ;
  assign n14150 = n5334 & n14105 ;
  assign n14148 = ~n5334 & n14101 ;
  assign n14149 = n5095 & ~n14145 ;
  assign n14151 = n5338 & ~n14149 ;
  assign n14152 = ~n14148 & n14151 ;
  assign n14153 = ~n14150 & n14152 ;
  assign n14154 = ~n14147 & ~n14153 ;
  assign n14155 = \P1_InstQueue_reg[0][1]/NET0131  & ~n5291 ;
  assign n14156 = ~n2029 & n5324 ;
  assign n14157 = ~n14143 & ~n14156 ;
  assign n14158 = n3042 & ~n14157 ;
  assign n14159 = ~n14155 & ~n14158 ;
  assign n14160 = ~n14154 & n14159 ;
  assign n14161 = ~n5185 & ~n5353 ;
  assign n14162 = \P1_InstQueue_reg[10][1]/NET0131  & ~n5107 ;
  assign n14163 = ~n5151 & n14162 ;
  assign n14164 = ~n14161 & ~n14163 ;
  assign n14165 = ~n7697 & ~n14164 ;
  assign n14166 = ~n7775 & ~n14165 ;
  assign n14169 = n5359 & n14105 ;
  assign n14167 = ~n5359 & n14101 ;
  assign n14168 = n5095 & ~n14164 ;
  assign n14170 = n5361 & ~n14168 ;
  assign n14171 = ~n14167 & n14170 ;
  assign n14172 = ~n14169 & n14171 ;
  assign n14173 = ~n14166 & ~n14172 ;
  assign n14174 = \P1_InstQueue_reg[10][1]/NET0131  & ~n5291 ;
  assign n14175 = ~n2029 & n5107 ;
  assign n14176 = ~n14162 & ~n14175 ;
  assign n14177 = n3042 & ~n14176 ;
  assign n14178 = ~n14174 & ~n14177 ;
  assign n14179 = ~n14173 & n14178 ;
  assign n14180 = ~n5185 & ~n5378 ;
  assign n14181 = \P1_InstQueue_reg[12][1]/NET0131  & ~n5377 ;
  assign n14182 = ~n5104 & n14181 ;
  assign n14183 = ~n14180 & ~n14182 ;
  assign n14184 = ~n7697 & ~n14183 ;
  assign n14185 = ~n7795 & ~n14184 ;
  assign n14188 = n5151 & n14105 ;
  assign n14186 = ~n5151 & n14101 ;
  assign n14187 = n5095 & ~n14183 ;
  assign n14189 = n5384 & ~n14187 ;
  assign n14190 = ~n14186 & n14189 ;
  assign n14191 = ~n14188 & n14190 ;
  assign n14192 = ~n14185 & ~n14191 ;
  assign n14193 = \P1_InstQueue_reg[12][1]/NET0131  & ~n5291 ;
  assign n14194 = ~n2029 & n5377 ;
  assign n14195 = ~n14181 & ~n14194 ;
  assign n14196 = n3042 & ~n14195 ;
  assign n14197 = ~n14193 & ~n14196 ;
  assign n14198 = ~n14192 & n14197 ;
  assign n14199 = ~n5185 & ~n5399 ;
  assign n14200 = \P1_InstQueue_reg[13][1]/NET0131  & ~n5334 ;
  assign n14201 = ~n5377 & n14200 ;
  assign n14202 = ~n14199 & ~n14201 ;
  assign n14203 = ~n7697 & ~n14202 ;
  assign n14204 = ~n7815 & ~n14203 ;
  assign n14207 = n5107 & n14105 ;
  assign n14205 = ~n5107 & n14101 ;
  assign n14206 = n5095 & ~n14202 ;
  assign n14208 = n5405 & ~n14206 ;
  assign n14209 = ~n14205 & n14208 ;
  assign n14210 = ~n14207 & n14209 ;
  assign n14211 = ~n14204 & ~n14210 ;
  assign n14212 = \P1_InstQueue_reg[13][1]/NET0131  & ~n5291 ;
  assign n14213 = ~n2029 & n5334 ;
  assign n14214 = ~n14200 & ~n14213 ;
  assign n14215 = n3042 & ~n14214 ;
  assign n14216 = ~n14212 & ~n14215 ;
  assign n14217 = ~n14211 & n14216 ;
  assign n14218 = ~n5185 & ~n5337 ;
  assign n14219 = \P1_InstQueue_reg[14][1]/NET0131  & ~n5336 ;
  assign n14220 = ~n5334 & n14219 ;
  assign n14221 = ~n14218 & ~n14220 ;
  assign n14222 = ~n7697 & ~n14221 ;
  assign n14223 = ~n7835 & ~n14222 ;
  assign n14226 = n5104 & n14105 ;
  assign n14224 = ~n5104 & n14101 ;
  assign n14225 = n5095 & ~n14221 ;
  assign n14227 = n5425 & ~n14225 ;
  assign n14228 = ~n14224 & n14227 ;
  assign n14229 = ~n14226 & n14228 ;
  assign n14230 = ~n14223 & ~n14229 ;
  assign n14231 = \P1_InstQueue_reg[14][1]/NET0131  & ~n5291 ;
  assign n14232 = ~n2029 & n5336 ;
  assign n14233 = ~n14219 & ~n14232 ;
  assign n14234 = n3042 & ~n14233 ;
  assign n14235 = ~n14231 & ~n14234 ;
  assign n14236 = ~n14230 & n14235 ;
  assign n14237 = ~n5185 & ~n5440 ;
  assign n14238 = \P1_InstQueue_reg[15][1]/NET0131  & ~n5326 ;
  assign n14239 = ~n5336 & n14238 ;
  assign n14240 = ~n14237 & ~n14239 ;
  assign n14241 = ~n7697 & ~n14240 ;
  assign n14242 = ~n7855 & ~n14241 ;
  assign n14245 = n5377 & n14105 ;
  assign n14243 = ~n5377 & n14101 ;
  assign n14244 = n5095 & ~n14240 ;
  assign n14246 = n5446 & ~n14244 ;
  assign n14247 = ~n14243 & n14246 ;
  assign n14248 = ~n14245 & n14247 ;
  assign n14249 = ~n14242 & ~n14248 ;
  assign n14250 = \P1_InstQueue_reg[15][1]/NET0131  & ~n5291 ;
  assign n14251 = ~n2029 & n5326 ;
  assign n14252 = ~n14238 & ~n14251 ;
  assign n14253 = n3042 & ~n14252 ;
  assign n14254 = ~n14250 & ~n14253 ;
  assign n14255 = ~n14249 & n14254 ;
  assign n14256 = ~n5185 & ~n5462 ;
  assign n14257 = \P1_InstQueue_reg[1][1]/NET0131  & ~n5461 ;
  assign n14258 = ~n5324 & n14257 ;
  assign n14259 = ~n14256 & ~n14258 ;
  assign n14260 = ~n7697 & ~n14259 ;
  assign n14261 = ~n7875 & ~n14260 ;
  assign n14264 = n5336 & n14105 ;
  assign n14262 = ~n5336 & n14101 ;
  assign n14263 = n5095 & ~n14259 ;
  assign n14265 = n5468 & ~n14263 ;
  assign n14266 = ~n14262 & n14265 ;
  assign n14267 = ~n14264 & n14266 ;
  assign n14268 = ~n14261 & ~n14267 ;
  assign n14269 = \P1_InstQueue_reg[1][1]/NET0131  & ~n5291 ;
  assign n14270 = ~n2029 & n5461 ;
  assign n14271 = ~n14257 & ~n14270 ;
  assign n14272 = n3042 & ~n14271 ;
  assign n14273 = ~n14269 & ~n14272 ;
  assign n14274 = ~n14268 & n14273 ;
  assign n14275 = ~n5185 & ~n5506 ;
  assign n14276 = \P1_InstQueue_reg[2][1]/NET0131  & ~n5484 ;
  assign n14277 = ~n5461 & n14276 ;
  assign n14278 = ~n14275 & ~n14277 ;
  assign n14279 = ~n7697 & ~n14278 ;
  assign n14280 = ~n7895 & ~n14279 ;
  assign n14283 = n5326 & n14105 ;
  assign n14281 = ~n5326 & n14101 ;
  assign n14282 = n5095 & ~n14278 ;
  assign n14284 = n5512 & ~n14282 ;
  assign n14285 = ~n14281 & n14284 ;
  assign n14286 = ~n14283 & n14285 ;
  assign n14287 = ~n14280 & ~n14286 ;
  assign n14288 = \P1_InstQueue_reg[2][1]/NET0131  & ~n5291 ;
  assign n14289 = ~n2029 & n5484 ;
  assign n14290 = ~n14276 & ~n14289 ;
  assign n14291 = n3042 & ~n14290 ;
  assign n14292 = ~n14288 & ~n14291 ;
  assign n14293 = ~n14287 & n14292 ;
  assign n14294 = ~n5185 & ~n5485 ;
  assign n14295 = \P1_InstQueue_reg[3][1]/NET0131  & ~n5483 ;
  assign n14296 = ~n5484 & n14295 ;
  assign n14297 = ~n14294 & ~n14296 ;
  assign n14298 = ~n7697 & ~n14297 ;
  assign n14299 = ~n7915 & ~n14298 ;
  assign n14302 = n5324 & n14105 ;
  assign n14300 = ~n5324 & n14101 ;
  assign n14301 = n5095 & ~n14297 ;
  assign n14303 = n5491 & ~n14301 ;
  assign n14304 = ~n14300 & n14303 ;
  assign n14305 = ~n14302 & n14304 ;
  assign n14306 = ~n14299 & ~n14305 ;
  assign n14307 = \P1_InstQueue_reg[3][1]/NET0131  & ~n5291 ;
  assign n14308 = ~n2029 & n5483 ;
  assign n14309 = ~n14295 & ~n14308 ;
  assign n14310 = n3042 & ~n14309 ;
  assign n14311 = ~n14307 & ~n14310 ;
  assign n14312 = ~n14306 & n14311 ;
  assign n14313 = ~n5185 & ~n5528 ;
  assign n14314 = \P1_InstQueue_reg[4][1]/NET0131  & ~n5527 ;
  assign n14315 = ~n5483 & n14314 ;
  assign n14316 = ~n14313 & ~n14315 ;
  assign n14317 = ~n7697 & ~n14316 ;
  assign n14318 = ~n7935 & ~n14317 ;
  assign n14321 = n5461 & n14105 ;
  assign n14319 = ~n5461 & n14101 ;
  assign n14320 = n5095 & ~n14316 ;
  assign n14322 = n5534 & ~n14320 ;
  assign n14323 = ~n14319 & n14322 ;
  assign n14324 = ~n14321 & n14323 ;
  assign n14325 = ~n14318 & ~n14324 ;
  assign n14326 = \P1_InstQueue_reg[4][1]/NET0131  & ~n5291 ;
  assign n14327 = ~n2029 & n5527 ;
  assign n14328 = ~n14314 & ~n14327 ;
  assign n14329 = n3042 & ~n14328 ;
  assign n14330 = ~n14326 & ~n14329 ;
  assign n14331 = ~n14325 & n14330 ;
  assign n14332 = ~n5185 & ~n5550 ;
  assign n14333 = \P1_InstQueue_reg[5][1]/NET0131  & ~n5549 ;
  assign n14334 = ~n5527 & n14333 ;
  assign n14335 = ~n14332 & ~n14334 ;
  assign n14336 = ~n7697 & ~n14335 ;
  assign n14337 = ~n7955 & ~n14336 ;
  assign n14340 = n5484 & n14105 ;
  assign n14338 = ~n5484 & n14101 ;
  assign n14339 = n5095 & ~n14335 ;
  assign n14341 = n5556 & ~n14339 ;
  assign n14342 = ~n14338 & n14341 ;
  assign n14343 = ~n14340 & n14342 ;
  assign n14344 = ~n14337 & ~n14343 ;
  assign n14345 = \P1_InstQueue_reg[5][1]/NET0131  & ~n5291 ;
  assign n14346 = ~n2029 & n5549 ;
  assign n14347 = ~n14333 & ~n14346 ;
  assign n14348 = n3042 & ~n14347 ;
  assign n14349 = ~n14345 & ~n14348 ;
  assign n14350 = ~n14344 & n14349 ;
  assign n14351 = ~n5185 & ~n5572 ;
  assign n14352 = \P1_InstQueue_reg[6][1]/NET0131  & ~n5571 ;
  assign n14353 = ~n5549 & n14352 ;
  assign n14354 = ~n14351 & ~n14353 ;
  assign n14355 = ~n7697 & ~n14354 ;
  assign n14356 = ~n7975 & ~n14355 ;
  assign n14359 = n5483 & n14105 ;
  assign n14357 = ~n5483 & n14101 ;
  assign n14358 = n5095 & ~n14354 ;
  assign n14360 = n5578 & ~n14358 ;
  assign n14361 = ~n14357 & n14360 ;
  assign n14362 = ~n14359 & n14361 ;
  assign n14363 = ~n14356 & ~n14362 ;
  assign n14364 = \P1_InstQueue_reg[6][1]/NET0131  & ~n5291 ;
  assign n14365 = ~n2029 & n5571 ;
  assign n14366 = ~n14352 & ~n14365 ;
  assign n14367 = n3042 & ~n14366 ;
  assign n14368 = ~n14364 & ~n14367 ;
  assign n14369 = ~n14363 & n14368 ;
  assign n14370 = ~n5185 & ~n5593 ;
  assign n14371 = \P1_InstQueue_reg[7][1]/NET0131  & ~n5359 ;
  assign n14372 = ~n5571 & n14371 ;
  assign n14373 = ~n14370 & ~n14372 ;
  assign n14374 = ~n7697 & ~n14373 ;
  assign n14375 = ~n7995 & ~n14374 ;
  assign n14378 = n5527 & n14105 ;
  assign n14376 = ~n5527 & n14101 ;
  assign n14377 = n5095 & ~n14373 ;
  assign n14379 = n5599 & ~n14377 ;
  assign n14380 = ~n14376 & n14379 ;
  assign n14381 = ~n14378 & n14380 ;
  assign n14382 = ~n14375 & ~n14381 ;
  assign n14383 = \P1_InstQueue_reg[7][1]/NET0131  & ~n5291 ;
  assign n14384 = ~n2029 & n5359 ;
  assign n14385 = ~n14371 & ~n14384 ;
  assign n14386 = n3042 & ~n14385 ;
  assign n14387 = ~n14383 & ~n14386 ;
  assign n14388 = ~n14382 & n14387 ;
  assign n14389 = ~n5185 & ~n5360 ;
  assign n14390 = \P1_InstQueue_reg[8][1]/NET0131  & ~n5148 ;
  assign n14391 = ~n5359 & n14390 ;
  assign n14392 = ~n14389 & ~n14391 ;
  assign n14393 = ~n7697 & ~n14392 ;
  assign n14394 = ~n8015 & ~n14393 ;
  assign n14397 = n5549 & n14105 ;
  assign n14395 = ~n5549 & n14101 ;
  assign n14396 = n5095 & ~n14392 ;
  assign n14398 = n5619 & ~n14396 ;
  assign n14399 = ~n14395 & n14398 ;
  assign n14400 = ~n14397 & n14399 ;
  assign n14401 = ~n14394 & ~n14400 ;
  assign n14402 = \P1_InstQueue_reg[8][1]/NET0131  & ~n5291 ;
  assign n14403 = ~n2029 & n5148 ;
  assign n14404 = ~n14390 & ~n14403 ;
  assign n14405 = n3042 & ~n14404 ;
  assign n14406 = ~n14402 & ~n14405 ;
  assign n14407 = ~n14401 & n14406 ;
  assign n14408 = ~n5152 & ~n5185 ;
  assign n14409 = \P1_InstQueue_reg[9][1]/NET0131  & ~n5151 ;
  assign n14410 = ~n5148 & n14409 ;
  assign n14411 = ~n14408 & ~n14410 ;
  assign n14412 = ~n7697 & ~n14411 ;
  assign n14413 = ~n8035 & ~n14412 ;
  assign n14416 = n5571 & n14105 ;
  assign n14414 = ~n5571 & n14101 ;
  assign n14415 = n5095 & ~n14411 ;
  assign n14417 = n5639 & ~n14415 ;
  assign n14418 = ~n14414 & n14417 ;
  assign n14419 = ~n14416 & n14418 ;
  assign n14420 = ~n14413 & ~n14419 ;
  assign n14421 = \P1_InstQueue_reg[9][1]/NET0131  & ~n5291 ;
  assign n14422 = ~n2029 & n5151 ;
  assign n14423 = ~n14409 & ~n14422 ;
  assign n14424 = n3042 & ~n14423 ;
  assign n14425 = ~n14421 & ~n14424 ;
  assign n14426 = ~n14420 & n14425 ;
  assign n14430 = \P2_PhyAddrPointer_reg[7]/NET0131  & n1897 ;
  assign n14431 = ~n10231 & ~n14430 ;
  assign n14432 = n1734 & ~n14431 ;
  assign n14433 = \P2_PhyAddrPointer_reg[7]/NET0131  & ~n8936 ;
  assign n14434 = ~n10248 & ~n14433 ;
  assign n14435 = ~n14432 & n14434 ;
  assign n14436 = n1927 & ~n14435 ;
  assign n14439 = n8964 & ~n10965 ;
  assign n14437 = n8963 & ~n10965 ;
  assign n14438 = ~\P2_PhyAddrPointer_reg[7]/NET0131  & ~n14437 ;
  assign n14440 = n1931 & ~n14438 ;
  assign n14441 = ~n14439 & n14440 ;
  assign n14427 = ~\P2_PhyAddrPointer_reg[7]/NET0131  & ~n13043 ;
  assign n14428 = ~n13044 & ~n14427 ;
  assign n14429 = n3087 & n14428 ;
  assign n14442 = \P2_PhyAddrPointer_reg[7]/NET0131  & ~n8958 ;
  assign n14443 = ~n10218 & ~n14442 ;
  assign n14444 = ~n14429 & n14443 ;
  assign n14445 = ~n14441 & n14444 ;
  assign n14446 = ~n14436 & n14445 ;
  assign n14450 = \P2_PhyAddrPointer_reg[9]/NET0131  & n1897 ;
  assign n14451 = ~n10274 & ~n14450 ;
  assign n14452 = n1734 & ~n14451 ;
  assign n14453 = \P2_PhyAddrPointer_reg[9]/NET0131  & ~n8936 ;
  assign n14454 = ~n10282 & ~n14453 ;
  assign n14455 = ~n14452 & n14454 ;
  assign n14456 = n1927 & ~n14455 ;
  assign n14447 = ~\P2_PhyAddrPointer_reg[9]/NET0131  & ~n13046 ;
  assign n14448 = ~n12373 & ~n14447 ;
  assign n14457 = ~\P2_DataWidth_reg[1]/NET0131  & ~n14448 ;
  assign n14458 = ~\P2_PhyAddrPointer_reg[9]/NET0131  & ~n8965 ;
  assign n14459 = ~n8966 & ~n14458 ;
  assign n14460 = \P2_DataWidth_reg[1]/NET0131  & ~n14459 ;
  assign n14461 = n1931 & ~n14460 ;
  assign n14462 = ~n14457 & n14461 ;
  assign n14449 = n3087 & n14448 ;
  assign n14463 = \P2_PhyAddrPointer_reg[9]/NET0131  & ~n8958 ;
  assign n14464 = ~n10262 & ~n14463 ;
  assign n14465 = ~n14449 & n14464 ;
  assign n14466 = ~n14462 & n14465 ;
  assign n14467 = ~n14456 & n14466 ;
  assign n14472 = ~n6071 & ~n10188 ;
  assign n14473 = ~n11971 & ~n14472 ;
  assign n14474 = n3753 & ~n14473 ;
  assign n14475 = n4215 & ~n10193 ;
  assign n14476 = ~n3753 & ~n4230 ;
  assign n14477 = ~n14475 & n14476 ;
  assign n14478 = ~n2896 & ~n14477 ;
  assign n14479 = ~n14474 & n14478 ;
  assign n14480 = n2894 & n14479 ;
  assign n14481 = \P3_PhyAddrPointer_reg[10]/NET0131  & ~n11965 ;
  assign n14482 = ~n4301 & ~n9105 ;
  assign n14483 = n2905 & ~n9106 ;
  assign n14484 = ~n14482 & n14483 ;
  assign n14485 = ~n14481 & ~n14484 ;
  assign n14486 = ~n14480 & n14485 ;
  assign n14487 = n2453 & ~n14486 ;
  assign n14468 = \P3_PhyAddrPointer_reg[1]/NET0131  & n9026 ;
  assign n14469 = ~\P3_PhyAddrPointer_reg[10]/NET0131  & ~n14468 ;
  assign n14470 = ~n11960 & ~n14469 ;
  assign n14488 = ~\P3_DataWidth_reg[1]/NET0131  & ~n14470 ;
  assign n14489 = ~\P3_PhyAddrPointer_reg[10]/NET0131  & ~n9026 ;
  assign n14490 = ~n9027 & ~n14489 ;
  assign n14491 = \P3_DataWidth_reg[1]/NET0131  & ~n14490 ;
  assign n14492 = n2959 & ~n14491 ;
  assign n14493 = ~n14488 & n14492 ;
  assign n14471 = n4415 & n14470 ;
  assign n14494 = \P3_rEIP_reg[10]/NET0131  & n4412 ;
  assign n14495 = \P3_PhyAddrPointer_reg[10]/NET0131  & ~n9063 ;
  assign n14496 = ~n14494 & ~n14495 ;
  assign n14497 = ~n14471 & n14496 ;
  assign n14498 = ~n14493 & n14497 ;
  assign n14499 = ~n14487 & n14498 ;
  assign n14503 = \P3_PhyAddrPointer_reg[7]/NET0131  & n2896 ;
  assign n14504 = ~n10153 & ~n14503 ;
  assign n14505 = n2894 & ~n14504 ;
  assign n14506 = \P3_PhyAddrPointer_reg[7]/NET0131  & ~n9014 ;
  assign n14507 = ~n10163 & ~n14506 ;
  assign n14508 = ~n14505 & n14507 ;
  assign n14509 = n2453 & ~n14508 ;
  assign n14500 = ~\P3_PhyAddrPointer_reg[7]/NET0131  & ~n13249 ;
  assign n14501 = ~n13250 & ~n14500 ;
  assign n14510 = ~\P3_DataWidth_reg[1]/NET0131  & ~n14501 ;
  assign n14511 = ~\P3_PhyAddrPointer_reg[7]/NET0131  & ~n9023 ;
  assign n14512 = ~n9024 & ~n14511 ;
  assign n14513 = \P3_DataWidth_reg[1]/NET0131  & ~n14512 ;
  assign n14514 = n2959 & ~n14513 ;
  assign n14515 = ~n14510 & n14514 ;
  assign n14502 = n4415 & n14501 ;
  assign n14516 = \P3_PhyAddrPointer_reg[7]/NET0131  & ~n9063 ;
  assign n14517 = ~n10170 & ~n14516 ;
  assign n14518 = ~n14502 & n14517 ;
  assign n14519 = ~n14515 & n14518 ;
  assign n14520 = ~n14509 & n14519 ;
  assign n14524 = \P3_PhyAddrPointer_reg[9]/NET0131  & n2896 ;
  assign n14525 = ~n10197 & ~n14524 ;
  assign n14526 = n2894 & ~n14525 ;
  assign n14527 = \P3_PhyAddrPointer_reg[9]/NET0131  & ~n9014 ;
  assign n14528 = ~n10205 & ~n14527 ;
  assign n14529 = ~n14526 & n14528 ;
  assign n14530 = n2453 & ~n14529 ;
  assign n14521 = ~\P3_PhyAddrPointer_reg[9]/NET0131  & ~n13252 ;
  assign n14522 = ~n14468 & ~n14521 ;
  assign n14531 = ~\P3_DataWidth_reg[1]/NET0131  & ~n14522 ;
  assign n14532 = ~\P3_PhyAddrPointer_reg[9]/NET0131  & ~n9025 ;
  assign n14533 = ~n9026 & ~n14532 ;
  assign n14534 = \P3_DataWidth_reg[1]/NET0131  & ~n14533 ;
  assign n14535 = n2959 & ~n14534 ;
  assign n14536 = ~n14531 & n14535 ;
  assign n14523 = n4415 & n14522 ;
  assign n14537 = \P3_PhyAddrPointer_reg[9]/NET0131  & ~n9063 ;
  assign n14538 = ~n10173 & ~n14537 ;
  assign n14539 = ~n14523 & n14538 ;
  assign n14540 = ~n14536 & n14539 ;
  assign n14541 = ~n14530 & n14540 ;
  assign n14545 = \P1_PhyAddrPointer_reg[10]/NET0131  & n2375 ;
  assign n14546 = ~n9212 & ~n14545 ;
  assign n14547 = n2244 & ~n14546 ;
  assign n14548 = \P1_PhyAddrPointer_reg[10]/NET0131  & ~n10087 ;
  assign n14549 = ~n9201 & ~n14548 ;
  assign n14550 = ~n14547 & n14549 ;
  assign n14551 = n2432 & ~n14550 ;
  assign n14542 = ~\P1_PhyAddrPointer_reg[10]/NET0131  & ~n12152 ;
  assign n14543 = ~n12153 & ~n14542 ;
  assign n14552 = ~\P1_DataWidth_reg[1]/NET0131  & ~n14543 ;
  assign n14553 = ~\P1_PhyAddrPointer_reg[10]/NET0131  & ~n10098 ;
  assign n14554 = ~n10099 & ~n14553 ;
  assign n14555 = \P1_DataWidth_reg[1]/NET0131  & ~n14554 ;
  assign n14556 = n2436 & ~n14555 ;
  assign n14557 = ~n14552 & n14556 ;
  assign n14544 = n5095 & n14543 ;
  assign n14558 = \P1_PhyAddrPointer_reg[10]/NET0131  & ~n10136 ;
  assign n14559 = ~n9195 & ~n14558 ;
  assign n14560 = ~n14544 & n14559 ;
  assign n14561 = ~n14557 & n14560 ;
  assign n14562 = ~n14551 & n14561 ;
  assign n14568 = \P1_PhyAddrPointer_reg[7]/NET0131  & n2375 ;
  assign n14569 = n4504 & ~n6841 ;
  assign n14570 = ~n4504 & n6841 ;
  assign n14571 = ~n14569 & ~n14570 ;
  assign n14572 = n4453 & ~n14571 ;
  assign n14573 = n4826 & ~n6855 ;
  assign n14574 = ~n4453 & ~n13505 ;
  assign n14575 = ~n14573 & n14574 ;
  assign n14576 = ~n2375 & ~n14575 ;
  assign n14577 = ~n14572 & n14576 ;
  assign n14578 = ~n14568 & ~n14577 ;
  assign n14579 = n2244 & ~n14578 ;
  assign n14563 = ~n4980 & ~n5014 ;
  assign n14565 = n6001 & n14563 ;
  assign n14564 = ~n6001 & ~n14563 ;
  assign n14566 = n2385 & ~n14564 ;
  assign n14567 = ~n14565 & n14566 ;
  assign n14580 = \P1_PhyAddrPointer_reg[7]/NET0131  & ~n10087 ;
  assign n14581 = ~n14567 & ~n14580 ;
  assign n14582 = ~n14579 & n14581 ;
  assign n14583 = n2432 & ~n14582 ;
  assign n14587 = \P1_PhyAddrPointer_reg[1]/NET0131  & n10094 ;
  assign n14588 = \P1_PhyAddrPointer_reg[6]/NET0131  & n14587 ;
  assign n14589 = ~\P1_PhyAddrPointer_reg[7]/NET0131  & ~n14588 ;
  assign n14590 = ~n12150 & ~n14589 ;
  assign n14591 = n10133 & n14590 ;
  assign n14584 = ~\P1_PhyAddrPointer_reg[7]/NET0131  & ~n10095 ;
  assign n14585 = n3148 & ~n10096 ;
  assign n14586 = ~n14584 & n14585 ;
  assign n14592 = \P1_rEIP_reg[7]/NET0131  & n5092 ;
  assign n14593 = \P1_PhyAddrPointer_reg[7]/NET0131  & ~n10136 ;
  assign n14594 = ~n14592 & ~n14593 ;
  assign n14595 = ~n14586 & n14594 ;
  assign n14596 = ~n14591 & n14595 ;
  assign n14597 = ~n14583 & n14596 ;
  assign n14608 = \P1_PhyAddrPointer_reg[9]/NET0131  & n2375 ;
  assign n14612 = ~n4499 & ~n4765 ;
  assign n14613 = ~n4766 & ~n14612 ;
  assign n14614 = n4453 & ~n14613 ;
  assign n14609 = n4871 & ~n5954 ;
  assign n14610 = ~n4453 & ~n4874 ;
  assign n14611 = ~n14609 & n14610 ;
  assign n14615 = ~n2375 & ~n14611 ;
  assign n14616 = ~n14614 & n14615 ;
  assign n14617 = ~n14608 & ~n14616 ;
  assign n14618 = n2244 & ~n14617 ;
  assign n14601 = ~\P1_InstAddrPointer_reg[9]/NET0131  & ~n4961 ;
  assign n14602 = ~n5021 & ~n14601 ;
  assign n14603 = ~n6002 & n6003 ;
  assign n14605 = n14602 & n14603 ;
  assign n14604 = ~n14602 & ~n14603 ;
  assign n14606 = n2385 & ~n14604 ;
  assign n14607 = ~n14605 & n14606 ;
  assign n14619 = \P1_PhyAddrPointer_reg[9]/NET0131  & ~n10087 ;
  assign n14620 = ~n14607 & ~n14619 ;
  assign n14621 = ~n14618 & n14620 ;
  assign n14622 = n2432 & ~n14621 ;
  assign n14598 = ~\P1_PhyAddrPointer_reg[9]/NET0131  & ~n12151 ;
  assign n14599 = ~n12152 & ~n14598 ;
  assign n14623 = ~\P1_DataWidth_reg[1]/NET0131  & ~n14599 ;
  assign n14624 = ~\P1_PhyAddrPointer_reg[9]/NET0131  & ~n10097 ;
  assign n14625 = ~n10098 & ~n14624 ;
  assign n14626 = \P1_DataWidth_reg[1]/NET0131  & ~n14625 ;
  assign n14627 = n2436 & ~n14626 ;
  assign n14628 = ~n14623 & n14627 ;
  assign n14600 = n5095 & n14599 ;
  assign n14629 = \P1_rEIP_reg[9]/NET0131  & n5092 ;
  assign n14630 = \P1_PhyAddrPointer_reg[9]/NET0131  & ~n10136 ;
  assign n14631 = ~n14629 & ~n14630 ;
  assign n14632 = ~n14600 & n14631 ;
  assign n14633 = ~n14628 & n14632 ;
  assign n14634 = ~n14622 & n14633 ;
  assign n14638 = \P2_PhyAddrPointer_reg[10]/NET0131  & n1897 ;
  assign n14639 = ~n9177 & ~n14638 ;
  assign n14640 = n1734 & ~n14639 ;
  assign n14641 = \P2_PhyAddrPointer_reg[10]/NET0131  & ~n8936 ;
  assign n14642 = ~n9183 & ~n14641 ;
  assign n14643 = ~n14640 & n14642 ;
  assign n14644 = n1927 & ~n14643 ;
  assign n14635 = ~\P2_PhyAddrPointer_reg[10]/NET0131  & ~n12373 ;
  assign n14636 = ~n12374 & ~n14635 ;
  assign n14645 = ~\P2_DataWidth_reg[1]/NET0131  & ~n14636 ;
  assign n14646 = ~\P2_PhyAddrPointer_reg[10]/NET0131  & ~n8966 ;
  assign n14647 = ~n12367 & ~n14646 ;
  assign n14648 = \P2_DataWidth_reg[1]/NET0131  & ~n14647 ;
  assign n14649 = n1931 & ~n14648 ;
  assign n14650 = ~n14645 & n14649 ;
  assign n14637 = n3087 & n14636 ;
  assign n14651 = \P2_PhyAddrPointer_reg[10]/NET0131  & ~n8958 ;
  assign n14652 = ~n9159 & ~n14651 ;
  assign n14653 = ~n14637 & n14652 ;
  assign n14654 = ~n14650 & n14653 ;
  assign n14655 = ~n14644 & n14654 ;
  assign n14657 = \P3_InstAddrPointer_reg[0]/NET0131  & n3963 ;
  assign n14658 = ~n4326 & ~n14657 ;
  assign n14659 = n2904 & ~n14658 ;
  assign n14660 = n2905 & n14658 ;
  assign n14661 = ~n14659 & ~n14660 ;
  assign n14662 = ~\P3_InstAddrPointer_reg[0]/NET0131  & n2919 ;
  assign n14663 = \P3_InstAddrPointer_reg[0]/NET0131  & n2768 ;
  assign n14664 = n2902 & n14663 ;
  assign n14665 = ~n14662 & ~n14664 ;
  assign n14666 = n14661 & ~n14665 ;
  assign n14667 = n2453 & ~n14666 ;
  assign n14656 = \P3_rEIP_reg[0]/NET0131  & n4412 ;
  assign n14668 = \P3_InstAddrPointer_reg[0]/NET0131  & ~n4418 ;
  assign n14669 = ~n14656 & ~n14668 ;
  assign n14670 = ~n14667 & n14669 ;
  assign n14672 = \P3_InstAddrPointer_reg[1]/NET0131  & ~n7403 ;
  assign n14697 = ~\P3_InstAddrPointer_reg[1]/NET0131  & ~n2923 ;
  assign n14696 = ~n2777 & ~n4323 ;
  assign n14673 = \P3_InstAddrPointer_reg[1]/NET0131  & n2896 ;
  assign n14676 = ~n3931 & ~n3932 ;
  assign n14677 = n14657 & ~n14676 ;
  assign n14674 = ~n4324 & ~n4325 ;
  assign n14675 = ~n14657 & n14674 ;
  assign n14678 = ~n3753 & ~n14675 ;
  assign n14679 = ~n14677 & n14678 ;
  assign n14681 = n3964 & n14676 ;
  assign n14680 = ~n3964 & ~n14676 ;
  assign n14682 = n3753 & ~n14680 ;
  assign n14683 = ~n14681 & n14682 ;
  assign n14684 = ~n14679 & ~n14683 ;
  assign n14685 = ~n2896 & ~n14684 ;
  assign n14686 = ~n14673 & ~n14685 ;
  assign n14687 = n2894 & ~n14686 ;
  assign n14688 = ~\P3_InstAddrPointer_reg[1]/NET0131  & ~n2847 ;
  assign n14689 = n2847 & n4323 ;
  assign n14690 = ~n14688 & ~n14689 ;
  assign n14691 = ~n2841 & n14690 ;
  assign n14692 = ~n4326 & ~n14674 ;
  assign n14693 = n4326 & ~n14676 ;
  assign n14694 = ~n14692 & ~n14693 ;
  assign n14695 = n2905 & n14694 ;
  assign n14698 = ~n14691 & ~n14695 ;
  assign n14699 = ~n14687 & n14698 ;
  assign n14700 = ~n14696 & n14699 ;
  assign n14701 = ~n14697 & n14700 ;
  assign n14702 = ~n14672 & n14701 ;
  assign n14703 = n2453 & ~n14702 ;
  assign n14671 = \P3_InstAddrPointer_reg[1]/NET0131  & ~n4418 ;
  assign n14704 = \P3_rEIP_reg[1]/NET0131  & n4412 ;
  assign n14705 = ~n14671 & ~n14704 ;
  assign n14706 = ~n14703 & n14705 ;
  assign n14715 = ~\P2_InstAddrPointer_reg[0]/NET0131  & n1871 ;
  assign n14716 = \P2_InstAddrPointer_reg[0]/NET0131  & n1748 ;
  assign n14717 = n1903 & n14716 ;
  assign n14718 = ~n14715 & ~n14717 ;
  assign n14709 = \P2_InstAddrPointer_reg[0]/NET0131  & n1897 ;
  assign n14710 = ~n6369 & ~n6715 ;
  assign n14711 = ~n1897 & ~n14710 ;
  assign n14712 = ~n14709 & ~n14711 ;
  assign n14713 = n1734 & ~n14712 ;
  assign n14714 = n1890 & n14710 ;
  assign n14719 = ~n14713 & ~n14714 ;
  assign n14720 = ~n14718 & n14719 ;
  assign n14721 = n1927 & ~n14720 ;
  assign n14707 = \P2_rEIP_reg[0]/NET0131  & n3113 ;
  assign n14708 = \P2_InstAddrPointer_reg[0]/NET0131  & ~n6810 ;
  assign n14722 = ~n14707 & ~n14708 ;
  assign n14723 = ~n14721 & n14722 ;
  assign n14732 = n2238 & n2373 ;
  assign n14733 = \P1_InstAddrPointer_reg[0]/NET0131  & ~n14732 ;
  assign n14731 = ~\P1_InstAddrPointer_reg[0]/NET0131  & ~n2398 ;
  assign n14726 = \P1_InstAddrPointer_reg[0]/NET0131  & n2375 ;
  assign n14727 = ~n4842 & ~n4997 ;
  assign n14728 = ~n2375 & ~n14727 ;
  assign n14729 = ~n14726 & ~n14728 ;
  assign n14730 = n2244 & ~n14729 ;
  assign n14734 = n2385 & n14727 ;
  assign n14735 = ~n14730 & ~n14734 ;
  assign n14736 = ~n14731 & n14735 ;
  assign n14737 = ~n14733 & n14736 ;
  assign n14738 = n2432 & ~n14737 ;
  assign n14724 = \P1_rEIP_reg[0]/NET0131  & n5092 ;
  assign n14725 = \P1_InstAddrPointer_reg[0]/NET0131  & ~n5098 ;
  assign n14739 = ~n14724 & ~n14725 ;
  assign n14740 = ~n14738 & n14739 ;
  assign n14743 = ~n1771 & n6335 ;
  assign n14771 = ~n1804 & n1811 ;
  assign n14772 = ~\P2_InstAddrPointer_reg[1]/NET0131  & ~n1739 ;
  assign n14773 = ~n14771 & n14772 ;
  assign n14774 = ~n1804 & n1805 ;
  assign n14775 = \P2_InstAddrPointer_reg[1]/NET0131  & ~n14774 ;
  assign n14776 = n7636 & n14775 ;
  assign n14777 = ~n14773 & ~n14776 ;
  assign n14748 = \P2_InstAddrPointer_reg[1]/NET0131  & n1897 ;
  assign n14751 = ~n6336 & ~n6714 ;
  assign n14752 = ~n6369 & n14751 ;
  assign n14749 = ~n6337 & ~n6613 ;
  assign n14750 = n6369 & ~n14749 ;
  assign n14753 = ~n6188 & ~n14750 ;
  assign n14754 = ~n14752 & n14753 ;
  assign n14756 = n6614 & n14749 ;
  assign n14755 = ~n6614 & ~n14749 ;
  assign n14757 = n6188 & ~n14755 ;
  assign n14758 = ~n14756 & n14757 ;
  assign n14759 = ~n14754 & ~n14758 ;
  assign n14760 = ~n1897 & ~n14759 ;
  assign n14761 = ~n14748 & ~n14760 ;
  assign n14762 = n1734 & ~n14761 ;
  assign n14744 = ~\P2_InstAddrPointer_reg[1]/NET0131  & ~n1820 ;
  assign n14745 = \P2_InstAddrPointer_reg[1]/NET0131  & n1820 ;
  assign n14746 = ~n14744 & ~n14745 ;
  assign n14747 = n7639 & n14746 ;
  assign n14763 = ~n6715 & ~n14751 ;
  assign n14764 = n6715 & ~n14749 ;
  assign n14765 = ~n14763 & ~n14764 ;
  assign n14766 = n1890 & n14765 ;
  assign n14767 = n1798 & ~n6335 ;
  assign n14768 = ~\P2_InstAddrPointer_reg[1]/NET0131  & ~n1798 ;
  assign n14769 = ~n14767 & ~n14768 ;
  assign n14770 = ~n1727 & n14769 ;
  assign n14778 = ~n14766 & ~n14770 ;
  assign n14779 = ~n14747 & n14778 ;
  assign n14780 = ~n14762 & n14779 ;
  assign n14781 = ~n14777 & n14780 ;
  assign n14782 = ~n14743 & n14781 ;
  assign n14783 = n1927 & ~n14782 ;
  assign n14741 = \P2_rEIP_reg[1]/NET0131  & n3113 ;
  assign n14742 = \P2_InstAddrPointer_reg[1]/NET0131  & ~n6810 ;
  assign n14784 = ~n14741 & ~n14742 ;
  assign n14785 = ~n14783 & n14784 ;
  assign n14809 = ~n2388 & ~n5080 ;
  assign n14810 = n2373 & n14809 ;
  assign n14811 = \P1_InstAddrPointer_reg[1]/NET0131  & ~n2376 ;
  assign n14812 = n14810 & n14811 ;
  assign n14813 = n2387 & n7308 ;
  assign n14814 = ~\P1_InstAddrPointer_reg[1]/NET0131  & ~n2237 ;
  assign n14815 = ~n14813 & n14814 ;
  assign n14816 = ~n14812 & ~n14815 ;
  assign n14787 = ~n2398 & n4840 ;
  assign n14790 = ~n4841 & ~n4996 ;
  assign n14791 = ~n4842 & n14790 ;
  assign n14788 = ~n4711 & ~n4712 ;
  assign n14789 = n4842 & ~n14788 ;
  assign n14792 = ~n4453 & ~n14789 ;
  assign n14793 = ~n14791 & n14792 ;
  assign n14795 = n4744 & n14788 ;
  assign n14794 = ~n4744 & ~n14788 ;
  assign n14796 = n4453 & ~n14794 ;
  assign n14797 = ~n14795 & n14796 ;
  assign n14798 = ~n14793 & ~n14797 ;
  assign n14799 = n2384 & ~n14798 ;
  assign n14800 = ~n4997 & ~n14790 ;
  assign n14801 = n4997 & ~n14788 ;
  assign n14802 = ~n14800 & ~n14801 ;
  assign n14803 = n2385 & n14802 ;
  assign n14804 = ~n14799 & ~n14803 ;
  assign n14806 = \P1_InstAddrPointer_reg[1]/NET0131  & n2377 ;
  assign n14805 = ~\P1_InstAddrPointer_reg[1]/NET0131  & ~n2377 ;
  assign n14807 = ~n7247 & ~n14805 ;
  assign n14808 = ~n14806 & n14807 ;
  assign n14817 = n14804 & ~n14808 ;
  assign n14818 = ~n14787 & n14817 ;
  assign n14819 = ~n14816 & n14818 ;
  assign n14820 = n2432 & ~n14819 ;
  assign n14786 = \P1_InstAddrPointer_reg[1]/NET0131  & ~n5098 ;
  assign n14821 = \P1_rEIP_reg[1]/NET0131  & n5092 ;
  assign n14822 = ~n14786 & ~n14821 ;
  assign n14823 = ~n14820 & n14822 ;
  assign n14824 = \P3_EAX_reg[31]/NET0131  & ~n13810 ;
  assign n14924 = \P3_EAX_reg[28]/NET0131  & n14045 ;
  assign n14925 = \P3_EAX_reg[29]/NET0131  & n14924 ;
  assign n14926 = \P3_EAX_reg[30]/NET0131  & n14925 ;
  assign n14928 = \P3_EAX_reg[31]/NET0131  & n14926 ;
  assign n14927 = ~\P3_EAX_reg[31]/NET0131  & ~n14926 ;
  assign n14929 = n13813 & ~n14927 ;
  assign n14930 = ~n14928 & n14929 ;
  assign n14829 = \P3_InstQueue_reg[14][5]/NET0131  & n2464 ;
  assign n14830 = \P3_InstQueue_reg[0][5]/NET0131  & n2472 ;
  assign n14843 = ~n14829 & ~n14830 ;
  assign n14831 = \P3_InstQueue_reg[13][5]/NET0131  & n2490 ;
  assign n14832 = \P3_InstQueue_reg[10][5]/NET0131  & n2474 ;
  assign n14844 = ~n14831 & ~n14832 ;
  assign n14851 = n14843 & n14844 ;
  assign n14825 = \P3_InstQueue_reg[4][5]/NET0131  & n2482 ;
  assign n14826 = \P3_InstQueue_reg[9][5]/NET0131  & n2492 ;
  assign n14841 = ~n14825 & ~n14826 ;
  assign n14827 = \P3_InstQueue_reg[3][5]/NET0131  & n2484 ;
  assign n14828 = \P3_InstQueue_reg[6][5]/NET0131  & n2466 ;
  assign n14842 = ~n14827 & ~n14828 ;
  assign n14852 = n14841 & n14842 ;
  assign n14853 = n14851 & n14852 ;
  assign n14837 = \P3_InstQueue_reg[1][5]/NET0131  & n2478 ;
  assign n14838 = \P3_InstQueue_reg[7][5]/NET0131  & n2480 ;
  assign n14847 = ~n14837 & ~n14838 ;
  assign n14839 = \P3_InstQueue_reg[11][5]/NET0131  & n2460 ;
  assign n14840 = \P3_InstQueue_reg[12][5]/NET0131  & n2476 ;
  assign n14848 = ~n14839 & ~n14840 ;
  assign n14849 = n14847 & n14848 ;
  assign n14833 = \P3_InstQueue_reg[15][5]/NET0131  & n2486 ;
  assign n14834 = \P3_InstQueue_reg[8][5]/NET0131  & n2469 ;
  assign n14845 = ~n14833 & ~n14834 ;
  assign n14835 = \P3_InstQueue_reg[5][5]/NET0131  & n2456 ;
  assign n14836 = \P3_InstQueue_reg[2][5]/NET0131  & n2488 ;
  assign n14846 = ~n14835 & ~n14836 ;
  assign n14850 = n14845 & n14846 ;
  assign n14854 = n14849 & n14850 ;
  assign n14855 = n14853 & n14854 ;
  assign n14856 = n14010 & ~n14855 ;
  assign n14861 = \P3_InstQueue_reg[14][6]/NET0131  & n2464 ;
  assign n14862 = \P3_InstQueue_reg[0][6]/NET0131  & n2472 ;
  assign n14875 = ~n14861 & ~n14862 ;
  assign n14863 = \P3_InstQueue_reg[13][6]/NET0131  & n2490 ;
  assign n14864 = \P3_InstQueue_reg[10][6]/NET0131  & n2474 ;
  assign n14876 = ~n14863 & ~n14864 ;
  assign n14883 = n14875 & n14876 ;
  assign n14857 = \P3_InstQueue_reg[4][6]/NET0131  & n2482 ;
  assign n14858 = \P3_InstQueue_reg[9][6]/NET0131  & n2492 ;
  assign n14873 = ~n14857 & ~n14858 ;
  assign n14859 = \P3_InstQueue_reg[3][6]/NET0131  & n2484 ;
  assign n14860 = \P3_InstQueue_reg[6][6]/NET0131  & n2466 ;
  assign n14874 = ~n14859 & ~n14860 ;
  assign n14884 = n14873 & n14874 ;
  assign n14885 = n14883 & n14884 ;
  assign n14869 = \P3_InstQueue_reg[1][6]/NET0131  & n2478 ;
  assign n14870 = \P3_InstQueue_reg[7][6]/NET0131  & n2480 ;
  assign n14879 = ~n14869 & ~n14870 ;
  assign n14871 = \P3_InstQueue_reg[11][6]/NET0131  & n2460 ;
  assign n14872 = \P3_InstQueue_reg[12][6]/NET0131  & n2476 ;
  assign n14880 = ~n14871 & ~n14872 ;
  assign n14881 = n14879 & n14880 ;
  assign n14865 = \P3_InstQueue_reg[15][6]/NET0131  & n2486 ;
  assign n14866 = \P3_InstQueue_reg[8][6]/NET0131  & n2469 ;
  assign n14877 = ~n14865 & ~n14866 ;
  assign n14867 = \P3_InstQueue_reg[5][6]/NET0131  & n2456 ;
  assign n14868 = \P3_InstQueue_reg[2][6]/NET0131  & n2488 ;
  assign n14878 = ~n14867 & ~n14868 ;
  assign n14882 = n14877 & n14878 ;
  assign n14886 = n14881 & n14882 ;
  assign n14887 = n14885 & n14886 ;
  assign n14888 = n14856 & ~n14887 ;
  assign n14893 = \P3_InstQueue_reg[14][7]/NET0131  & n2464 ;
  assign n14894 = \P3_InstQueue_reg[0][7]/NET0131  & n2472 ;
  assign n14907 = ~n14893 & ~n14894 ;
  assign n14895 = \P3_InstQueue_reg[13][7]/NET0131  & n2490 ;
  assign n14896 = \P3_InstQueue_reg[10][7]/NET0131  & n2474 ;
  assign n14908 = ~n14895 & ~n14896 ;
  assign n14915 = n14907 & n14908 ;
  assign n14889 = \P3_InstQueue_reg[4][7]/NET0131  & n2482 ;
  assign n14890 = \P3_InstQueue_reg[9][7]/NET0131  & n2492 ;
  assign n14905 = ~n14889 & ~n14890 ;
  assign n14891 = \P3_InstQueue_reg[3][7]/NET0131  & n2484 ;
  assign n14892 = \P3_InstQueue_reg[6][7]/NET0131  & n2466 ;
  assign n14906 = ~n14891 & ~n14892 ;
  assign n14916 = n14905 & n14906 ;
  assign n14917 = n14915 & n14916 ;
  assign n14901 = \P3_InstQueue_reg[1][7]/NET0131  & n2478 ;
  assign n14902 = \P3_InstQueue_reg[7][7]/NET0131  & n2480 ;
  assign n14911 = ~n14901 & ~n14902 ;
  assign n14903 = \P3_InstQueue_reg[11][7]/NET0131  & n2460 ;
  assign n14904 = \P3_InstQueue_reg[12][7]/NET0131  & n2476 ;
  assign n14912 = ~n14903 & ~n14904 ;
  assign n14913 = n14911 & n14912 ;
  assign n14897 = \P3_InstQueue_reg[15][7]/NET0131  & n2486 ;
  assign n14898 = \P3_InstQueue_reg[8][7]/NET0131  & n2469 ;
  assign n14909 = ~n14897 & ~n14898 ;
  assign n14899 = \P3_InstQueue_reg[5][7]/NET0131  & n2456 ;
  assign n14900 = \P3_InstQueue_reg[2][7]/NET0131  & n2488 ;
  assign n14910 = ~n14899 & ~n14900 ;
  assign n14914 = n14909 & n14910 ;
  assign n14918 = n14913 & n14914 ;
  assign n14919 = n14917 & n14918 ;
  assign n14920 = n14888 & ~n14919 ;
  assign n14921 = n13812 & n14920 ;
  assign n14922 = ~n2864 & n13817 ;
  assign n14923 = \P3_EAX_reg[31]/NET0131  & ~n14922 ;
  assign n14931 = ~n14921 & ~n14923 ;
  assign n14932 = ~n14930 & n14931 ;
  assign n14933 = n2453 & ~n14932 ;
  assign n14934 = ~n14824 & ~n14933 ;
  assign n14935 = \P3_EAX_reg[30]/NET0131  & ~n13810 ;
  assign n14939 = ~\P3_EAX_reg[30]/NET0131  & ~n14925 ;
  assign n14940 = n13813 & ~n14926 ;
  assign n14941 = ~n14939 & n14940 ;
  assign n14942 = \P3_EAX_reg[30]/NET0131  & ~n14922 ;
  assign n14936 = ~n14888 & n14919 ;
  assign n14937 = ~n14920 & ~n14936 ;
  assign n14938 = n13812 & n14937 ;
  assign n14943 = \buf2_reg[30]/NET0131  & n2820 ;
  assign n14944 = \buf2_reg[14]/NET0131  & n2821 ;
  assign n14945 = ~n14943 & ~n14944 ;
  assign n14946 = n2862 & ~n14945 ;
  assign n14947 = ~n14938 & ~n14946 ;
  assign n14948 = ~n14942 & n14947 ;
  assign n14949 = ~n14941 & n14948 ;
  assign n14950 = n2453 & ~n14949 ;
  assign n14951 = ~n14935 & ~n14950 ;
  assign n14957 = \P3_EBX_reg[0]/NET0131  & \P3_EBX_reg[1]/NET0131  ;
  assign n14958 = \P3_EBX_reg[2]/NET0131  & n14957 ;
  assign n14959 = \P3_EBX_reg[3]/NET0131  & n14958 ;
  assign n14960 = \P3_EBX_reg[4]/NET0131  & n14959 ;
  assign n14961 = \P3_EBX_reg[5]/NET0131  & n14960 ;
  assign n14962 = \P3_EBX_reg[6]/NET0131  & n14961 ;
  assign n14963 = \P3_EBX_reg[7]/NET0131  & n14962 ;
  assign n14964 = \P3_EBX_reg[8]/NET0131  & n14963 ;
  assign n14965 = \P3_EBX_reg[9]/NET0131  & n14964 ;
  assign n14966 = \P3_EBX_reg[10]/NET0131  & n14965 ;
  assign n14967 = \P3_EBX_reg[11]/NET0131  & n14966 ;
  assign n14968 = \P3_EBX_reg[12]/NET0131  & n14967 ;
  assign n14969 = \P3_EBX_reg[13]/NET0131  & n14968 ;
  assign n14970 = \P3_EBX_reg[14]/NET0131  & n14969 ;
  assign n14971 = \P3_EBX_reg[15]/NET0131  & n14970 ;
  assign n14972 = \P3_EBX_reg[16]/NET0131  & n14971 ;
  assign n14973 = \P3_EBX_reg[17]/NET0131  & n14972 ;
  assign n14974 = \P3_EBX_reg[18]/NET0131  & n14973 ;
  assign n14975 = \P3_EBX_reg[19]/NET0131  & n14974 ;
  assign n14976 = \P3_EBX_reg[20]/NET0131  & \P3_EBX_reg[21]/NET0131  ;
  assign n14977 = \P3_EBX_reg[22]/NET0131  & \P3_EBX_reg[23]/NET0131  ;
  assign n14978 = n14976 & n14977 ;
  assign n14979 = n14975 & n14978 ;
  assign n14980 = \P3_EBX_reg[24]/NET0131  & n14979 ;
  assign n14981 = \P3_EBX_reg[25]/NET0131  & n14980 ;
  assign n14982 = \P3_EBX_reg[26]/NET0131  & \P3_EBX_reg[27]/NET0131  ;
  assign n14983 = \P3_EBX_reg[28]/NET0131  & \P3_EBX_reg[29]/NET0131  ;
  assign n14984 = n14982 & n14983 ;
  assign n14985 = n14981 & n14984 ;
  assign n14986 = \P3_EBX_reg[30]/NET0131  & n14985 ;
  assign n14988 = \P3_EBX_reg[31]/NET0131  & n14986 ;
  assign n14987 = ~\P3_EBX_reg[31]/NET0131  & ~n14986 ;
  assign n14989 = n2748 & ~n14987 ;
  assign n14990 = ~n14988 & n14989 ;
  assign n14952 = n2771 & n2847 ;
  assign n14953 = n2748 & ~n2770 ;
  assign n14954 = ~n14952 & ~n14953 ;
  assign n14955 = \P3_EBX_reg[31]/NET0131  & n14954 ;
  assign n14956 = n14920 & n14952 ;
  assign n14991 = ~n14955 & ~n14956 ;
  assign n14992 = ~n14990 & n14991 ;
  assign n14993 = n2453 & ~n14992 ;
  assign n14994 = \P3_EBX_reg[31]/NET0131  & ~n13810 ;
  assign n14995 = ~n14993 & ~n14994 ;
  assign n14996 = \P2_EAX_reg[30]/NET0131  & ~n12632 ;
  assign n14997 = ~\P2_EAX_reg[30]/NET0131  & ~n12662 ;
  assign n14998 = n12665 & ~n14997 ;
  assign n15001 = ~n12928 & ~n12959 ;
  assign n15002 = n12928 & n12959 ;
  assign n15003 = ~n15001 & ~n15002 ;
  assign n15004 = n1798 & ~n15003 ;
  assign n15005 = n1726 & n15004 ;
  assign n15006 = \P2_EAX_reg[30]/NET0131  & ~n12669 ;
  assign n14999 = n1803 & ~n7732 ;
  assign n15000 = n1811 & n14999 ;
  assign n15007 = ~\buf2_reg[14]/NET0131  & ~n3079 ;
  assign n15008 = ~\buf1_reg[14]/NET0131  & n3079 ;
  assign n15009 = ~n15007 & ~n15008 ;
  assign n15010 = n1811 & n15009 ;
  assign n15011 = n1742 & n15010 ;
  assign n15012 = ~n15000 & ~n15011 ;
  assign n15013 = ~n15006 & n15012 ;
  assign n15014 = ~n15005 & n15013 ;
  assign n15015 = ~n14998 & n15014 ;
  assign n15016 = n1927 & ~n15015 ;
  assign n15017 = ~n14996 & ~n15016 ;
  assign n15022 = \P2_EBX_reg[0]/NET0131  & \P2_EBX_reg[1]/NET0131  ;
  assign n15023 = \P2_EBX_reg[2]/NET0131  & n15022 ;
  assign n15024 = \P2_EBX_reg[3]/NET0131  & n15023 ;
  assign n15025 = \P2_EBX_reg[4]/NET0131  & n15024 ;
  assign n15026 = \P2_EBX_reg[5]/NET0131  & n15025 ;
  assign n15027 = \P2_EBX_reg[6]/NET0131  & n15026 ;
  assign n15028 = \P2_EBX_reg[7]/NET0131  & n15027 ;
  assign n15029 = \P2_EBX_reg[8]/NET0131  & n15028 ;
  assign n15030 = \P2_EBX_reg[9]/NET0131  & n15029 ;
  assign n15031 = \P2_EBX_reg[10]/NET0131  & n15030 ;
  assign n15032 = \P2_EBX_reg[11]/NET0131  & n15031 ;
  assign n15033 = \P2_EBX_reg[12]/NET0131  & n15032 ;
  assign n15034 = \P2_EBX_reg[13]/NET0131  & \P2_EBX_reg[14]/NET0131  ;
  assign n15035 = n15033 & n15034 ;
  assign n15036 = \P2_EBX_reg[15]/NET0131  & n15035 ;
  assign n15037 = \P2_EBX_reg[16]/NET0131  & n15036 ;
  assign n15038 = \P2_EBX_reg[17]/NET0131  & \P2_EBX_reg[18]/NET0131  ;
  assign n15039 = n15037 & n15038 ;
  assign n15040 = \P2_EBX_reg[19]/NET0131  & n15039 ;
  assign n15041 = \P2_EBX_reg[20]/NET0131  & \P2_EBX_reg[21]/NET0131  ;
  assign n15042 = \P2_EBX_reg[22]/NET0131  & \P2_EBX_reg[23]/NET0131  ;
  assign n15043 = n15041 & n15042 ;
  assign n15044 = n15040 & n15043 ;
  assign n15045 = \P2_EBX_reg[24]/NET0131  & \P2_EBX_reg[25]/NET0131  ;
  assign n15046 = n15044 & n15045 ;
  assign n15047 = \P2_EBX_reg[26]/NET0131  & n15046 ;
  assign n15049 = ~\P2_EBX_reg[27]/NET0131  & ~n15047 ;
  assign n15048 = \P2_EBX_reg[27]/NET0131  & n15047 ;
  assign n15050 = n1766 & ~n15048 ;
  assign n15051 = ~n15049 & n15050 ;
  assign n15018 = ~n1722 & ~n1766 ;
  assign n15019 = ~n1877 & ~n15018 ;
  assign n15020 = \P2_EBX_reg[27]/NET0131  & ~n15019 ;
  assign n15021 = n1722 & n14065 ;
  assign n15052 = ~n15020 & ~n15021 ;
  assign n15053 = ~n15051 & n15052 ;
  assign n15054 = n1927 & ~n15053 ;
  assign n15055 = \P2_EBX_reg[27]/NET0131  & ~n12632 ;
  assign n15056 = ~n15054 & ~n15055 ;
  assign n15060 = \P2_EBX_reg[28]/NET0131  & n15048 ;
  assign n15061 = \P2_EBX_reg[29]/NET0131  & n15060 ;
  assign n15062 = \P2_EBX_reg[30]/NET0131  & n15061 ;
  assign n15064 = \P2_EBX_reg[31]/NET0131  & n15062 ;
  assign n15063 = ~\P2_EBX_reg[31]/NET0131  & ~n15062 ;
  assign n15065 = n1766 & ~n15063 ;
  assign n15066 = ~n15064 & n15065 ;
  assign n15057 = \P2_EBX_reg[31]/NET0131  & ~n15019 ;
  assign n15058 = n1722 & n12960 ;
  assign n15059 = n12928 & n15058 ;
  assign n15067 = ~n15057 & ~n15059 ;
  assign n15068 = ~n15066 & n15067 ;
  assign n15069 = n1927 & ~n15068 ;
  assign n15070 = \P2_EBX_reg[31]/NET0131  & ~n12632 ;
  assign n15071 = ~n15069 & ~n15070 ;
  assign n15364 = \P1_EBX_reg[0]/NET0131  & \P1_EBX_reg[1]/NET0131  ;
  assign n15365 = \P1_EBX_reg[2]/NET0131  & n15364 ;
  assign n15366 = \P1_EBX_reg[3]/NET0131  & n15365 ;
  assign n15367 = \P1_EBX_reg[4]/NET0131  & n15366 ;
  assign n15368 = \P1_EBX_reg[5]/NET0131  & n15367 ;
  assign n15369 = \P1_EBX_reg[6]/NET0131  & n15368 ;
  assign n15370 = \P1_EBX_reg[7]/NET0131  & n15369 ;
  assign n15371 = \P1_EBX_reg[8]/NET0131  & n15370 ;
  assign n15372 = \P1_EBX_reg[9]/NET0131  & n15371 ;
  assign n15373 = \P1_EBX_reg[10]/NET0131  & n15372 ;
  assign n15374 = \P1_EBX_reg[11]/NET0131  & n15373 ;
  assign n15375 = \P1_EBX_reg[12]/NET0131  & n15374 ;
  assign n15376 = \P1_EBX_reg[13]/NET0131  & n15375 ;
  assign n15377 = \P1_EBX_reg[14]/NET0131  & n15376 ;
  assign n15378 = \P1_EBX_reg[15]/NET0131  & n15377 ;
  assign n15379 = \P1_EBX_reg[16]/NET0131  & n15378 ;
  assign n15380 = \P1_EBX_reg[17]/NET0131  & n15379 ;
  assign n15381 = \P1_EBX_reg[18]/NET0131  & n15380 ;
  assign n15382 = \P1_EBX_reg[19]/NET0131  & n15381 ;
  assign n15383 = \P1_EBX_reg[20]/NET0131  & \P1_EBX_reg[21]/NET0131  ;
  assign n15384 = \P1_EBX_reg[22]/NET0131  & \P1_EBX_reg[23]/NET0131  ;
  assign n15385 = n15383 & n15384 ;
  assign n15386 = n15382 & n15385 ;
  assign n15387 = \P1_EBX_reg[24]/NET0131  & n15386 ;
  assign n15388 = \P1_EBX_reg[25]/NET0131  & n15387 ;
  assign n15389 = \P1_EBX_reg[26]/NET0131  & n15388 ;
  assign n15390 = \P1_EBX_reg[27]/NET0131  & \P1_EBX_reg[28]/NET0131  ;
  assign n15391 = \P1_EBX_reg[29]/NET0131  & \P1_EBX_reg[30]/NET0131  ;
  assign n15392 = n15390 & n15391 ;
  assign n15393 = n15389 & n15392 ;
  assign n15395 = \P1_EBX_reg[31]/NET0131  & n15393 ;
  assign n15394 = ~\P1_EBX_reg[31]/NET0131  & ~n15393 ;
  assign n15396 = n2262 & ~n15394 ;
  assign n15397 = ~n15395 & n15396 ;
  assign n15072 = ~n2242 & ~n2262 ;
  assign n15073 = ~n2370 & ~n15072 ;
  assign n15074 = \P1_EBX_reg[31]/NET0131  & ~n15073 ;
  assign n15110 = \P1_InstQueue_reg[7][7]/NET0131  & n1961 ;
  assign n15111 = \P1_InstQueue_reg[6][7]/NET0131  & n1976 ;
  assign n15124 = ~n15110 & ~n15111 ;
  assign n15112 = \P1_InstQueue_reg[5][7]/NET0131  & n1970 ;
  assign n15113 = \P1_InstQueue_reg[4][7]/NET0131  & n1966 ;
  assign n15125 = ~n15112 & ~n15113 ;
  assign n15132 = n15124 & n15125 ;
  assign n15106 = \P1_InstQueue_reg[8][7]/NET0131  & n1964 ;
  assign n15107 = \P1_InstQueue_reg[0][7]/NET0131  & n1980 ;
  assign n15122 = ~n15106 & ~n15107 ;
  assign n15108 = \P1_InstQueue_reg[13][7]/NET0131  & n1946 ;
  assign n15109 = \P1_InstQueue_reg[12][7]/NET0131  & n1978 ;
  assign n15123 = ~n15108 & ~n15109 ;
  assign n15133 = n15122 & n15123 ;
  assign n15134 = n15132 & n15133 ;
  assign n15118 = \P1_InstQueue_reg[9][7]/NET0131  & n1972 ;
  assign n15119 = \P1_InstQueue_reg[1][7]/NET0131  & n1955 ;
  assign n15128 = ~n15118 & ~n15119 ;
  assign n15120 = \P1_InstQueue_reg[15][7]/NET0131  & n1953 ;
  assign n15121 = \P1_InstQueue_reg[11][7]/NET0131  & n1974 ;
  assign n15129 = ~n15120 & ~n15121 ;
  assign n15130 = n15128 & n15129 ;
  assign n15114 = \P1_InstQueue_reg[3][7]/NET0131  & n1958 ;
  assign n15115 = \P1_InstQueue_reg[14][7]/NET0131  & n1949 ;
  assign n15126 = ~n15114 & ~n15115 ;
  assign n15116 = \P1_InstQueue_reg[10][7]/NET0131  & n1968 ;
  assign n15117 = \P1_InstQueue_reg[2][7]/NET0131  & n1982 ;
  assign n15127 = ~n15116 & ~n15117 ;
  assign n15131 = n15126 & n15127 ;
  assign n15135 = n15130 & n15131 ;
  assign n15136 = n15134 & n15135 ;
  assign n15141 = \P1_InstQueue_reg[6][0]/NET0131  & n1970 ;
  assign n15142 = \P1_InstQueue_reg[10][0]/NET0131  & n1972 ;
  assign n15155 = ~n15141 & ~n15142 ;
  assign n15143 = \P1_InstQueue_reg[14][0]/NET0131  & n1946 ;
  assign n15144 = \P1_InstQueue_reg[5][0]/NET0131  & n1966 ;
  assign n15156 = ~n15143 & ~n15144 ;
  assign n15163 = n15155 & n15156 ;
  assign n15137 = \P1_InstQueue_reg[13][0]/NET0131  & n1978 ;
  assign n15138 = \P1_InstQueue_reg[12][0]/NET0131  & n1974 ;
  assign n15153 = ~n15137 & ~n15138 ;
  assign n15139 = \P1_InstQueue_reg[9][0]/NET0131  & n1964 ;
  assign n15140 = \P1_InstQueue_reg[15][0]/NET0131  & n1949 ;
  assign n15154 = ~n15139 & ~n15140 ;
  assign n15164 = n15153 & n15154 ;
  assign n15165 = n15163 & n15164 ;
  assign n15149 = \P1_InstQueue_reg[4][0]/NET0131  & n1958 ;
  assign n15150 = \P1_InstQueue_reg[2][0]/NET0131  & n1955 ;
  assign n15159 = ~n15149 & ~n15150 ;
  assign n15151 = \P1_InstQueue_reg[7][0]/NET0131  & n1976 ;
  assign n15152 = \P1_InstQueue_reg[1][0]/NET0131  & n1980 ;
  assign n15160 = ~n15151 & ~n15152 ;
  assign n15161 = n15159 & n15160 ;
  assign n15145 = \P1_InstQueue_reg[11][0]/NET0131  & n1968 ;
  assign n15146 = \P1_InstQueue_reg[0][0]/NET0131  & n1953 ;
  assign n15157 = ~n15145 & ~n15146 ;
  assign n15147 = \P1_InstQueue_reg[8][0]/NET0131  & n1961 ;
  assign n15148 = \P1_InstQueue_reg[3][0]/NET0131  & n1982 ;
  assign n15158 = ~n15147 & ~n15148 ;
  assign n15162 = n15157 & n15158 ;
  assign n15166 = n15161 & n15162 ;
  assign n15167 = n15165 & n15166 ;
  assign n15168 = ~n15136 & ~n15167 ;
  assign n15173 = \P1_InstQueue_reg[9][1]/NET0131  & n1964 ;
  assign n15174 = \P1_InstQueue_reg[7][1]/NET0131  & n1976 ;
  assign n15187 = ~n15173 & ~n15174 ;
  assign n15175 = \P1_InstQueue_reg[4][1]/NET0131  & n1958 ;
  assign n15176 = \P1_InstQueue_reg[5][1]/NET0131  & n1966 ;
  assign n15188 = ~n15175 & ~n15176 ;
  assign n15195 = n15187 & n15188 ;
  assign n15169 = \P1_InstQueue_reg[6][1]/NET0131  & n1970 ;
  assign n15170 = \P1_InstQueue_reg[13][1]/NET0131  & n1978 ;
  assign n15185 = ~n15169 & ~n15170 ;
  assign n15171 = \P1_InstQueue_reg[12][1]/NET0131  & n1974 ;
  assign n15172 = \P1_InstQueue_reg[8][1]/NET0131  & n1961 ;
  assign n15186 = ~n15171 & ~n15172 ;
  assign n15196 = n15185 & n15186 ;
  assign n15197 = n15195 & n15196 ;
  assign n15181 = \P1_InstQueue_reg[11][1]/NET0131  & n1968 ;
  assign n15182 = \P1_InstQueue_reg[3][1]/NET0131  & n1982 ;
  assign n15191 = ~n15181 & ~n15182 ;
  assign n15183 = \P1_InstQueue_reg[1][1]/NET0131  & n1980 ;
  assign n15184 = \P1_InstQueue_reg[10][1]/NET0131  & n1972 ;
  assign n15192 = ~n15183 & ~n15184 ;
  assign n15193 = n15191 & n15192 ;
  assign n15177 = \P1_InstQueue_reg[0][1]/NET0131  & n1953 ;
  assign n15178 = \P1_InstQueue_reg[14][1]/NET0131  & n1946 ;
  assign n15189 = ~n15177 & ~n15178 ;
  assign n15179 = \P1_InstQueue_reg[15][1]/NET0131  & n1949 ;
  assign n15180 = \P1_InstQueue_reg[2][1]/NET0131  & n1955 ;
  assign n15190 = ~n15179 & ~n15180 ;
  assign n15194 = n15189 & n15190 ;
  assign n15198 = n15193 & n15194 ;
  assign n15199 = n15197 & n15198 ;
  assign n15200 = n15168 & ~n15199 ;
  assign n15205 = \P1_InstQueue_reg[6][2]/NET0131  & n1970 ;
  assign n15206 = \P1_InstQueue_reg[15][2]/NET0131  & n1949 ;
  assign n15219 = ~n15205 & ~n15206 ;
  assign n15207 = \P1_InstQueue_reg[14][2]/NET0131  & n1946 ;
  assign n15208 = \P1_InstQueue_reg[5][2]/NET0131  & n1966 ;
  assign n15220 = ~n15207 & ~n15208 ;
  assign n15227 = n15219 & n15220 ;
  assign n15201 = \P1_InstQueue_reg[9][2]/NET0131  & n1964 ;
  assign n15202 = \P1_InstQueue_reg[12][2]/NET0131  & n1974 ;
  assign n15217 = ~n15201 & ~n15202 ;
  assign n15203 = \P1_InstQueue_reg[13][2]/NET0131  & n1978 ;
  assign n15204 = \P1_InstQueue_reg[10][2]/NET0131  & n1972 ;
  assign n15218 = ~n15203 & ~n15204 ;
  assign n15228 = n15217 & n15218 ;
  assign n15229 = n15227 & n15228 ;
  assign n15213 = \P1_InstQueue_reg[4][2]/NET0131  & n1958 ;
  assign n15214 = \P1_InstQueue_reg[3][2]/NET0131  & n1982 ;
  assign n15223 = ~n15213 & ~n15214 ;
  assign n15215 = \P1_InstQueue_reg[7][2]/NET0131  & n1976 ;
  assign n15216 = \P1_InstQueue_reg[1][2]/NET0131  & n1980 ;
  assign n15224 = ~n15215 & ~n15216 ;
  assign n15225 = n15223 & n15224 ;
  assign n15209 = \P1_InstQueue_reg[11][2]/NET0131  & n1968 ;
  assign n15210 = \P1_InstQueue_reg[0][2]/NET0131  & n1953 ;
  assign n15221 = ~n15209 & ~n15210 ;
  assign n15211 = \P1_InstQueue_reg[8][2]/NET0131  & n1961 ;
  assign n15212 = \P1_InstQueue_reg[2][2]/NET0131  & n1955 ;
  assign n15222 = ~n15211 & ~n15212 ;
  assign n15226 = n15221 & n15222 ;
  assign n15230 = n15225 & n15226 ;
  assign n15231 = n15229 & n15230 ;
  assign n15232 = n15200 & ~n15231 ;
  assign n15237 = \P1_InstQueue_reg[9][3]/NET0131  & n1964 ;
  assign n15238 = \P1_InstQueue_reg[7][3]/NET0131  & n1976 ;
  assign n15251 = ~n15237 & ~n15238 ;
  assign n15239 = \P1_InstQueue_reg[4][3]/NET0131  & n1958 ;
  assign n15240 = \P1_InstQueue_reg[5][3]/NET0131  & n1966 ;
  assign n15252 = ~n15239 & ~n15240 ;
  assign n15259 = n15251 & n15252 ;
  assign n15233 = \P1_InstQueue_reg[6][3]/NET0131  & n1970 ;
  assign n15234 = \P1_InstQueue_reg[13][3]/NET0131  & n1978 ;
  assign n15249 = ~n15233 & ~n15234 ;
  assign n15235 = \P1_InstQueue_reg[12][3]/NET0131  & n1974 ;
  assign n15236 = \P1_InstQueue_reg[8][3]/NET0131  & n1961 ;
  assign n15250 = ~n15235 & ~n15236 ;
  assign n15260 = n15249 & n15250 ;
  assign n15261 = n15259 & n15260 ;
  assign n15245 = \P1_InstQueue_reg[11][3]/NET0131  & n1968 ;
  assign n15246 = \P1_InstQueue_reg[2][3]/NET0131  & n1955 ;
  assign n15255 = ~n15245 & ~n15246 ;
  assign n15247 = \P1_InstQueue_reg[1][3]/NET0131  & n1980 ;
  assign n15248 = \P1_InstQueue_reg[10][3]/NET0131  & n1972 ;
  assign n15256 = ~n15247 & ~n15248 ;
  assign n15257 = n15255 & n15256 ;
  assign n15241 = \P1_InstQueue_reg[0][3]/NET0131  & n1953 ;
  assign n15242 = \P1_InstQueue_reg[14][3]/NET0131  & n1946 ;
  assign n15253 = ~n15241 & ~n15242 ;
  assign n15243 = \P1_InstQueue_reg[15][3]/NET0131  & n1949 ;
  assign n15244 = \P1_InstQueue_reg[3][3]/NET0131  & n1982 ;
  assign n15254 = ~n15243 & ~n15244 ;
  assign n15258 = n15253 & n15254 ;
  assign n15262 = n15257 & n15258 ;
  assign n15263 = n15261 & n15262 ;
  assign n15264 = n15232 & ~n15263 ;
  assign n15269 = \P1_InstQueue_reg[13][4]/NET0131  & n1978 ;
  assign n15270 = \P1_InstQueue_reg[7][4]/NET0131  & n1976 ;
  assign n15283 = ~n15269 & ~n15270 ;
  assign n15271 = \P1_InstQueue_reg[4][4]/NET0131  & n1958 ;
  assign n15272 = \P1_InstQueue_reg[5][4]/NET0131  & n1966 ;
  assign n15284 = ~n15271 & ~n15272 ;
  assign n15291 = n15283 & n15284 ;
  assign n15265 = \P1_InstQueue_reg[6][4]/NET0131  & n1970 ;
  assign n15266 = \P1_InstQueue_reg[9][4]/NET0131  & n1964 ;
  assign n15281 = ~n15265 & ~n15266 ;
  assign n15267 = \P1_InstQueue_reg[12][4]/NET0131  & n1974 ;
  assign n15268 = \P1_InstQueue_reg[8][4]/NET0131  & n1961 ;
  assign n15282 = ~n15267 & ~n15268 ;
  assign n15292 = n15281 & n15282 ;
  assign n15293 = n15291 & n15292 ;
  assign n15277 = \P1_InstQueue_reg[11][4]/NET0131  & n1968 ;
  assign n15278 = \P1_InstQueue_reg[2][4]/NET0131  & n1955 ;
  assign n15287 = ~n15277 & ~n15278 ;
  assign n15279 = \P1_InstQueue_reg[1][4]/NET0131  & n1980 ;
  assign n15280 = \P1_InstQueue_reg[15][4]/NET0131  & n1949 ;
  assign n15288 = ~n15279 & ~n15280 ;
  assign n15289 = n15287 & n15288 ;
  assign n15273 = \P1_InstQueue_reg[0][4]/NET0131  & n1953 ;
  assign n15274 = \P1_InstQueue_reg[14][4]/NET0131  & n1946 ;
  assign n15285 = ~n15273 & ~n15274 ;
  assign n15275 = \P1_InstQueue_reg[10][4]/NET0131  & n1972 ;
  assign n15276 = \P1_InstQueue_reg[3][4]/NET0131  & n1982 ;
  assign n15286 = ~n15275 & ~n15276 ;
  assign n15290 = n15285 & n15286 ;
  assign n15294 = n15289 & n15290 ;
  assign n15295 = n15293 & n15294 ;
  assign n15296 = n15264 & ~n15295 ;
  assign n15301 = \P1_InstQueue_reg[13][5]/NET0131  & n1978 ;
  assign n15302 = \P1_InstQueue_reg[7][5]/NET0131  & n1976 ;
  assign n15315 = ~n15301 & ~n15302 ;
  assign n15303 = \P1_InstQueue_reg[4][5]/NET0131  & n1958 ;
  assign n15304 = \P1_InstQueue_reg[5][5]/NET0131  & n1966 ;
  assign n15316 = ~n15303 & ~n15304 ;
  assign n15323 = n15315 & n15316 ;
  assign n15297 = \P1_InstQueue_reg[6][5]/NET0131  & n1970 ;
  assign n15298 = \P1_InstQueue_reg[9][5]/NET0131  & n1964 ;
  assign n15313 = ~n15297 & ~n15298 ;
  assign n15299 = \P1_InstQueue_reg[12][5]/NET0131  & n1974 ;
  assign n15300 = \P1_InstQueue_reg[8][5]/NET0131  & n1961 ;
  assign n15314 = ~n15299 & ~n15300 ;
  assign n15324 = n15313 & n15314 ;
  assign n15325 = n15323 & n15324 ;
  assign n15309 = \P1_InstQueue_reg[11][5]/NET0131  & n1968 ;
  assign n15310 = \P1_InstQueue_reg[2][5]/NET0131  & n1955 ;
  assign n15319 = ~n15309 & ~n15310 ;
  assign n15311 = \P1_InstQueue_reg[1][5]/NET0131  & n1980 ;
  assign n15312 = \P1_InstQueue_reg[15][5]/NET0131  & n1949 ;
  assign n15320 = ~n15311 & ~n15312 ;
  assign n15321 = n15319 & n15320 ;
  assign n15305 = \P1_InstQueue_reg[0][5]/NET0131  & n1953 ;
  assign n15306 = \P1_InstQueue_reg[14][5]/NET0131  & n1946 ;
  assign n15317 = ~n15305 & ~n15306 ;
  assign n15307 = \P1_InstQueue_reg[10][5]/NET0131  & n1972 ;
  assign n15308 = \P1_InstQueue_reg[3][5]/NET0131  & n1982 ;
  assign n15318 = ~n15307 & ~n15308 ;
  assign n15322 = n15317 & n15318 ;
  assign n15326 = n15321 & n15322 ;
  assign n15327 = n15325 & n15326 ;
  assign n15328 = n15296 & ~n15327 ;
  assign n15333 = \P1_InstQueue_reg[13][6]/NET0131  & n1978 ;
  assign n15334 = \P1_InstQueue_reg[7][6]/NET0131  & n1976 ;
  assign n15347 = ~n15333 & ~n15334 ;
  assign n15335 = \P1_InstQueue_reg[4][6]/NET0131  & n1958 ;
  assign n15336 = \P1_InstQueue_reg[5][6]/NET0131  & n1966 ;
  assign n15348 = ~n15335 & ~n15336 ;
  assign n15355 = n15347 & n15348 ;
  assign n15329 = \P1_InstQueue_reg[6][6]/NET0131  & n1970 ;
  assign n15330 = \P1_InstQueue_reg[9][6]/NET0131  & n1964 ;
  assign n15345 = ~n15329 & ~n15330 ;
  assign n15331 = \P1_InstQueue_reg[12][6]/NET0131  & n1974 ;
  assign n15332 = \P1_InstQueue_reg[8][6]/NET0131  & n1961 ;
  assign n15346 = ~n15331 & ~n15332 ;
  assign n15356 = n15345 & n15346 ;
  assign n15357 = n15355 & n15356 ;
  assign n15341 = \P1_InstQueue_reg[11][6]/NET0131  & n1968 ;
  assign n15342 = \P1_InstQueue_reg[2][6]/NET0131  & n1955 ;
  assign n15351 = ~n15341 & ~n15342 ;
  assign n15343 = \P1_InstQueue_reg[1][6]/NET0131  & n1980 ;
  assign n15344 = \P1_InstQueue_reg[15][6]/NET0131  & n1949 ;
  assign n15352 = ~n15343 & ~n15344 ;
  assign n15353 = n15351 & n15352 ;
  assign n15337 = \P1_InstQueue_reg[0][6]/NET0131  & n1953 ;
  assign n15338 = \P1_InstQueue_reg[14][6]/NET0131  & n1946 ;
  assign n15349 = ~n15337 & ~n15338 ;
  assign n15339 = \P1_InstQueue_reg[10][6]/NET0131  & n1972 ;
  assign n15340 = \P1_InstQueue_reg[3][6]/NET0131  & n1982 ;
  assign n15350 = ~n15339 & ~n15340 ;
  assign n15354 = n15349 & n15350 ;
  assign n15358 = n15353 & n15354 ;
  assign n15359 = n15357 & n15358 ;
  assign n15360 = n15328 & ~n15359 ;
  assign n15079 = \P1_InstQueue_reg[13][7]/NET0131  & n1978 ;
  assign n15080 = \P1_InstQueue_reg[7][7]/NET0131  & n1976 ;
  assign n15093 = ~n15079 & ~n15080 ;
  assign n15081 = \P1_InstQueue_reg[4][7]/NET0131  & n1958 ;
  assign n15082 = \P1_InstQueue_reg[5][7]/NET0131  & n1966 ;
  assign n15094 = ~n15081 & ~n15082 ;
  assign n15101 = n15093 & n15094 ;
  assign n15075 = \P1_InstQueue_reg[6][7]/NET0131  & n1970 ;
  assign n15076 = \P1_InstQueue_reg[9][7]/NET0131  & n1964 ;
  assign n15091 = ~n15075 & ~n15076 ;
  assign n15077 = \P1_InstQueue_reg[12][7]/NET0131  & n1974 ;
  assign n15078 = \P1_InstQueue_reg[8][7]/NET0131  & n1961 ;
  assign n15092 = ~n15077 & ~n15078 ;
  assign n15102 = n15091 & n15092 ;
  assign n15103 = n15101 & n15102 ;
  assign n15087 = \P1_InstQueue_reg[11][7]/NET0131  & n1968 ;
  assign n15088 = \P1_InstQueue_reg[2][7]/NET0131  & n1955 ;
  assign n15097 = ~n15087 & ~n15088 ;
  assign n15089 = \P1_InstQueue_reg[1][7]/NET0131  & n1980 ;
  assign n15090 = \P1_InstQueue_reg[15][7]/NET0131  & n1949 ;
  assign n15098 = ~n15089 & ~n15090 ;
  assign n15099 = n15097 & n15098 ;
  assign n15083 = \P1_InstQueue_reg[0][7]/NET0131  & n1953 ;
  assign n15084 = \P1_InstQueue_reg[14][7]/NET0131  & n1946 ;
  assign n15095 = ~n15083 & ~n15084 ;
  assign n15085 = \P1_InstQueue_reg[10][7]/NET0131  & n1972 ;
  assign n15086 = \P1_InstQueue_reg[3][7]/NET0131  & n1982 ;
  assign n15096 = ~n15085 & ~n15086 ;
  assign n15100 = n15095 & n15096 ;
  assign n15104 = n15099 & n15100 ;
  assign n15105 = n15103 & n15104 ;
  assign n15361 = n2337 & ~n15105 ;
  assign n15362 = n15360 & n15361 ;
  assign n15363 = n2242 & n15362 ;
  assign n15398 = ~n15074 & ~n15363 ;
  assign n15399 = ~n15397 & n15398 ;
  assign n15400 = n2432 & ~n15399 ;
  assign n15401 = ~n3020 & ~n3027 ;
  assign n15402 = n14081 & n15401 ;
  assign n15403 = \P1_EBX_reg[31]/NET0131  & ~n15402 ;
  assign n15404 = ~n15400 & ~n15403 ;
  assign n15413 = \buf2_reg[24]/NET0131  & ~n3079 ;
  assign n15414 = \buf1_reg[24]/NET0131  & n3079 ;
  assign n15415 = ~n15413 & ~n15414 ;
  assign n15416 = n3091 & ~n15415 ;
  assign n15417 = \buf2_reg[16]/NET0131  & ~n3079 ;
  assign n15418 = \buf1_reg[16]/NET0131  & n3079 ;
  assign n15419 = ~n15417 & ~n15418 ;
  assign n15420 = n3098 & ~n15419 ;
  assign n15421 = ~n15416 & ~n15420 ;
  assign n15422 = \P2_DataWidth_reg[1]/NET0131  & ~n15421 ;
  assign n15405 = \buf2_reg[0]/NET0131  & ~n3079 ;
  assign n15406 = \buf1_reg[0]/NET0131  & n3079 ;
  assign n15407 = ~n15405 & ~n15406 ;
  assign n15408 = ~n3050 & ~n15407 ;
  assign n15409 = \P2_InstQueue_reg[11][0]/NET0131  & ~n3049 ;
  assign n15410 = ~n3046 & n15409 ;
  assign n15411 = ~n15408 & ~n15410 ;
  assign n15423 = ~n3106 & ~n15411 ;
  assign n15424 = ~n15422 & ~n15423 ;
  assign n15425 = n1931 & ~n15424 ;
  assign n15412 = n3087 & ~n15411 ;
  assign n15426 = ~n1498 & n3049 ;
  assign n15427 = ~n15409 & ~n15426 ;
  assign n15428 = n3040 & ~n15427 ;
  assign n15429 = \P2_InstQueue_reg[11][0]/NET0131  & ~n3118 ;
  assign n15430 = ~n15428 & ~n15429 ;
  assign n15431 = ~n15412 & n15430 ;
  assign n15432 = ~n15425 & n15431 ;
  assign n15437 = n2453 & ~n2855 ;
  assign n15438 = \P3_InstAddrPointer_reg[1]/NET0131  & ~\P3_InstAddrPointer_reg[31]/NET0131  ;
  assign n15439 = \P3_InstAddrPointer_reg[31]/NET0131  & ~n4323 ;
  assign n15440 = ~n15438 & ~n15439 ;
  assign n15441 = n14123 & ~n15440 ;
  assign n15442 = ~n3007 & ~n15441 ;
  assign n15443 = n2997 & ~n15442 ;
  assign n15433 = ~n2963 & ~n4412 ;
  assign n15434 = ~n3004 & n14120 ;
  assign n15435 = n15433 & n15434 ;
  assign n15436 = \P3_InstQueueRd_Addr_reg[2]/NET0131  & ~n15435 ;
  assign n15444 = n2780 & n2994 ;
  assign n15445 = ~n15436 & ~n15444 ;
  assign n15446 = ~n15443 & n15445 ;
  assign n15447 = ~n15437 & n15446 ;
  assign n15449 = ~n1837 & n1927 ;
  assign n15450 = \P2_InstAddrPointer_reg[31]/NET0131  & ~n6335 ;
  assign n15451 = ~\P2_InstAddrPointer_reg[1]/NET0131  & ~\P2_InstAddrPointer_reg[31]/NET0131  ;
  assign n15452 = ~n15450 & ~n15451 ;
  assign n15453 = n14135 & n15452 ;
  assign n15454 = ~n2981 & ~n15453 ;
  assign n15455 = n2980 & ~n15454 ;
  assign n15448 = \P2_InstQueueRd_Addr_reg[2]/NET0131  & ~n14133 ;
  assign n15456 = n1444 & n3040 ;
  assign n15457 = ~n15448 & ~n15456 ;
  assign n15458 = ~n15455 & n15457 ;
  assign n15459 = ~n15449 & n15458 ;
  assign n15465 = n3162 & ~n15415 ;
  assign n15466 = n3165 & ~n15419 ;
  assign n15467 = ~n15465 & ~n15466 ;
  assign n15468 = \P2_DataWidth_reg[1]/NET0131  & ~n15467 ;
  assign n15460 = ~n3155 & ~n15407 ;
  assign n15461 = \P2_InstQueue_reg[0][0]/NET0131  & ~n3152 ;
  assign n15462 = ~n3154 & n15461 ;
  assign n15463 = ~n15460 & ~n15462 ;
  assign n15469 = ~n3170 & ~n15463 ;
  assign n15470 = ~n15468 & ~n15469 ;
  assign n15471 = n1931 & ~n15470 ;
  assign n15464 = n3087 & ~n15463 ;
  assign n15472 = ~n1498 & n3152 ;
  assign n15473 = ~n15461 & ~n15472 ;
  assign n15474 = n3040 & ~n15473 ;
  assign n15475 = \P2_InstQueue_reg[0][0]/NET0131  & ~n3118 ;
  assign n15476 = ~n15474 & ~n15475 ;
  assign n15477 = ~n15464 & n15476 ;
  assign n15478 = ~n15471 & n15477 ;
  assign n15484 = n3091 & ~n15419 ;
  assign n15485 = n3198 & ~n15415 ;
  assign n15486 = ~n15484 & ~n15485 ;
  assign n15487 = \P2_DataWidth_reg[1]/NET0131  & ~n15486 ;
  assign n15479 = ~n3202 & ~n15407 ;
  assign n15480 = \P2_InstQueue_reg[10][0]/NET0131  & ~n3046 ;
  assign n15481 = ~n3098 & n15480 ;
  assign n15482 = ~n15479 & ~n15481 ;
  assign n15488 = ~n3200 & ~n15482 ;
  assign n15489 = ~n15487 & ~n15488 ;
  assign n15490 = n1931 & ~n15489 ;
  assign n15483 = n3087 & ~n15482 ;
  assign n15491 = ~n1498 & n3046 ;
  assign n15492 = ~n15480 & ~n15491 ;
  assign n15493 = n3040 & ~n15492 ;
  assign n15494 = \P2_InstQueue_reg[10][0]/NET0131  & ~n3118 ;
  assign n15495 = ~n15493 & ~n15494 ;
  assign n15496 = ~n15483 & n15495 ;
  assign n15497 = ~n15490 & n15496 ;
  assign n15503 = n3098 & ~n15415 ;
  assign n15504 = n3046 & ~n15419 ;
  assign n15505 = ~n15503 & ~n15504 ;
  assign n15506 = \P2_DataWidth_reg[1]/NET0131  & ~n15505 ;
  assign n15498 = ~n3238 & ~n15407 ;
  assign n15499 = \P2_InstQueue_reg[12][0]/NET0131  & ~n3237 ;
  assign n15500 = ~n3049 & n15499 ;
  assign n15501 = ~n15498 & ~n15500 ;
  assign n15507 = ~n3248 & ~n15501 ;
  assign n15508 = ~n15506 & ~n15507 ;
  assign n15509 = n1931 & ~n15508 ;
  assign n15502 = n3087 & ~n15501 ;
  assign n15510 = ~n1498 & n3237 ;
  assign n15511 = ~n15499 & ~n15510 ;
  assign n15512 = n3040 & ~n15511 ;
  assign n15513 = \P2_InstQueue_reg[12][0]/NET0131  & ~n3118 ;
  assign n15514 = ~n15512 & ~n15513 ;
  assign n15515 = ~n15502 & n15514 ;
  assign n15516 = ~n15509 & n15515 ;
  assign n15522 = n3046 & ~n15415 ;
  assign n15523 = n3049 & ~n15419 ;
  assign n15524 = ~n15522 & ~n15523 ;
  assign n15525 = \P2_DataWidth_reg[1]/NET0131  & ~n15524 ;
  assign n15517 = ~n3275 & ~n15407 ;
  assign n15518 = \P2_InstQueue_reg[13][0]/NET0131  & ~n3162 ;
  assign n15519 = ~n3237 & n15518 ;
  assign n15520 = ~n15517 & ~n15519 ;
  assign n15526 = ~n3285 & ~n15520 ;
  assign n15527 = ~n15525 & ~n15526 ;
  assign n15528 = n1931 & ~n15527 ;
  assign n15521 = n3087 & ~n15520 ;
  assign n15529 = ~n1498 & n3162 ;
  assign n15530 = ~n15518 & ~n15529 ;
  assign n15531 = n3040 & ~n15530 ;
  assign n15532 = \P2_InstQueue_reg[13][0]/NET0131  & ~n3118 ;
  assign n15533 = ~n15531 & ~n15532 ;
  assign n15534 = ~n15521 & n15533 ;
  assign n15535 = ~n15528 & n15534 ;
  assign n15541 = n3049 & ~n15415 ;
  assign n15542 = n3237 & ~n15419 ;
  assign n15543 = ~n15541 & ~n15542 ;
  assign n15544 = \P2_DataWidth_reg[1]/NET0131  & ~n15543 ;
  assign n15536 = ~n3169 & ~n15407 ;
  assign n15537 = \P2_InstQueue_reg[14][0]/NET0131  & ~n3165 ;
  assign n15538 = ~n3162 & n15537 ;
  assign n15539 = ~n15536 & ~n15538 ;
  assign n15545 = ~n3321 & ~n15539 ;
  assign n15546 = ~n15544 & ~n15545 ;
  assign n15547 = n1931 & ~n15546 ;
  assign n15540 = n3087 & ~n15539 ;
  assign n15548 = ~n1498 & n3165 ;
  assign n15549 = ~n15537 & ~n15548 ;
  assign n15550 = n3040 & ~n15549 ;
  assign n15551 = \P2_InstQueue_reg[14][0]/NET0131  & ~n3118 ;
  assign n15552 = ~n15550 & ~n15551 ;
  assign n15553 = ~n15540 & n15552 ;
  assign n15554 = ~n15547 & n15553 ;
  assign n15560 = n3237 & ~n15415 ;
  assign n15561 = n3162 & ~n15419 ;
  assign n15562 = ~n15560 & ~n15561 ;
  assign n15563 = \P2_DataWidth_reg[1]/NET0131  & ~n15562 ;
  assign n15555 = ~n3348 & ~n15407 ;
  assign n15556 = \P2_InstQueue_reg[15][0]/NET0131  & ~n3154 ;
  assign n15557 = ~n3165 & n15556 ;
  assign n15558 = ~n15555 & ~n15557 ;
  assign n15564 = ~n3358 & ~n15558 ;
  assign n15565 = ~n15563 & ~n15564 ;
  assign n15566 = n1931 & ~n15565 ;
  assign n15559 = n3087 & ~n15558 ;
  assign n15567 = ~n1498 & n3154 ;
  assign n15568 = ~n15556 & ~n15567 ;
  assign n15569 = n3040 & ~n15568 ;
  assign n15570 = \P2_InstQueue_reg[15][0]/NET0131  & ~n3118 ;
  assign n15571 = ~n15569 & ~n15570 ;
  assign n15572 = ~n15559 & n15571 ;
  assign n15573 = ~n15566 & n15572 ;
  assign n15579 = n3165 & ~n15415 ;
  assign n15580 = n3154 & ~n15419 ;
  assign n15581 = ~n15579 & ~n15580 ;
  assign n15582 = \P2_DataWidth_reg[1]/NET0131  & ~n15581 ;
  assign n15574 = ~n3389 & ~n15407 ;
  assign n15575 = \P2_InstQueue_reg[1][0]/NET0131  & ~n3388 ;
  assign n15576 = ~n3152 & n15575 ;
  assign n15577 = ~n15574 & ~n15576 ;
  assign n15583 = ~n3386 & ~n15577 ;
  assign n15584 = ~n15582 & ~n15583 ;
  assign n15585 = n1931 & ~n15584 ;
  assign n15578 = n3087 & ~n15577 ;
  assign n15586 = ~n1498 & n3388 ;
  assign n15587 = ~n15575 & ~n15586 ;
  assign n15588 = n3040 & ~n15587 ;
  assign n15589 = \P2_InstQueue_reg[1][0]/NET0131  & ~n3118 ;
  assign n15590 = ~n15588 & ~n15589 ;
  assign n15591 = ~n15578 & n15590 ;
  assign n15592 = ~n15585 & n15591 ;
  assign n15598 = n3152 & ~n15419 ;
  assign n15599 = n3154 & ~n15415 ;
  assign n15600 = ~n15598 & ~n15599 ;
  assign n15601 = \P2_DataWidth_reg[1]/NET0131  & ~n15600 ;
  assign n15593 = ~n3424 & ~n15407 ;
  assign n15594 = \P2_InstQueue_reg[2][0]/NET0131  & ~n3423 ;
  assign n15595 = ~n3388 & n15594 ;
  assign n15596 = ~n15593 & ~n15595 ;
  assign n15602 = ~n3434 & ~n15596 ;
  assign n15603 = ~n15601 & ~n15602 ;
  assign n15604 = n1931 & ~n15603 ;
  assign n15597 = n3087 & ~n15596 ;
  assign n15605 = ~n1498 & n3423 ;
  assign n15606 = ~n15594 & ~n15605 ;
  assign n15607 = n3040 & ~n15606 ;
  assign n15608 = \P2_InstQueue_reg[2][0]/NET0131  & ~n3118 ;
  assign n15609 = ~n15607 & ~n15608 ;
  assign n15610 = ~n15597 & n15609 ;
  assign n15611 = ~n15604 & n15610 ;
  assign n15617 = n3152 & ~n15415 ;
  assign n15618 = n3388 & ~n15419 ;
  assign n15619 = ~n15617 & ~n15618 ;
  assign n15620 = \P2_DataWidth_reg[1]/NET0131  & ~n15619 ;
  assign n15612 = ~n3462 & ~n15407 ;
  assign n15613 = \P2_InstQueue_reg[3][0]/NET0131  & ~n3461 ;
  assign n15614 = ~n3423 & n15613 ;
  assign n15615 = ~n15612 & ~n15614 ;
  assign n15621 = ~n3472 & ~n15615 ;
  assign n15622 = ~n15620 & ~n15621 ;
  assign n15623 = n1931 & ~n15622 ;
  assign n15616 = n3087 & ~n15615 ;
  assign n15624 = ~n1498 & n3461 ;
  assign n15625 = ~n15613 & ~n15624 ;
  assign n15626 = n3040 & ~n15625 ;
  assign n15627 = \P2_InstQueue_reg[3][0]/NET0131  & ~n3118 ;
  assign n15628 = ~n15626 & ~n15627 ;
  assign n15629 = ~n15616 & n15628 ;
  assign n15630 = ~n15623 & n15629 ;
  assign n15636 = n3388 & ~n15415 ;
  assign n15637 = n3423 & ~n15419 ;
  assign n15638 = ~n15636 & ~n15637 ;
  assign n15639 = \P2_DataWidth_reg[1]/NET0131  & ~n15638 ;
  assign n15631 = ~n3500 & ~n15407 ;
  assign n15632 = \P2_InstQueue_reg[4][0]/NET0131  & ~n3499 ;
  assign n15633 = ~n3461 & n15632 ;
  assign n15634 = ~n15631 & ~n15633 ;
  assign n15640 = ~n3510 & ~n15634 ;
  assign n15641 = ~n15639 & ~n15640 ;
  assign n15642 = n1931 & ~n15641 ;
  assign n15635 = n3087 & ~n15634 ;
  assign n15643 = ~n1498 & n3499 ;
  assign n15644 = ~n15632 & ~n15643 ;
  assign n15645 = n3040 & ~n15644 ;
  assign n15646 = \P2_InstQueue_reg[4][0]/NET0131  & ~n3118 ;
  assign n15647 = ~n15645 & ~n15646 ;
  assign n15648 = ~n15635 & n15647 ;
  assign n15649 = ~n15642 & n15648 ;
  assign n15655 = n3423 & ~n15415 ;
  assign n15656 = n3461 & ~n15419 ;
  assign n15657 = ~n15655 & ~n15656 ;
  assign n15658 = \P2_DataWidth_reg[1]/NET0131  & ~n15657 ;
  assign n15650 = ~n3538 & ~n15407 ;
  assign n15651 = \P2_InstQueue_reg[5][0]/NET0131  & ~n3537 ;
  assign n15652 = ~n3499 & n15651 ;
  assign n15653 = ~n15650 & ~n15652 ;
  assign n15659 = ~n3548 & ~n15653 ;
  assign n15660 = ~n15658 & ~n15659 ;
  assign n15661 = n1931 & ~n15660 ;
  assign n15654 = n3087 & ~n15653 ;
  assign n15662 = ~n1498 & n3537 ;
  assign n15663 = ~n15651 & ~n15662 ;
  assign n15664 = n3040 & ~n15663 ;
  assign n15665 = \P2_InstQueue_reg[5][0]/NET0131  & ~n3118 ;
  assign n15666 = ~n15664 & ~n15665 ;
  assign n15667 = ~n15654 & n15666 ;
  assign n15668 = ~n15661 & n15667 ;
  assign n15674 = n3461 & ~n15415 ;
  assign n15675 = n3499 & ~n15419 ;
  assign n15676 = ~n15674 & ~n15675 ;
  assign n15677 = \P2_DataWidth_reg[1]/NET0131  & ~n15676 ;
  assign n15669 = ~n3576 & ~n15407 ;
  assign n15670 = \P2_InstQueue_reg[6][0]/NET0131  & ~n3575 ;
  assign n15671 = ~n3537 & n15670 ;
  assign n15672 = ~n15669 & ~n15671 ;
  assign n15678 = ~n3586 & ~n15672 ;
  assign n15679 = ~n15677 & ~n15678 ;
  assign n15680 = n1931 & ~n15679 ;
  assign n15673 = n3087 & ~n15672 ;
  assign n15681 = ~n1498 & n3575 ;
  assign n15682 = ~n15670 & ~n15681 ;
  assign n15683 = n3040 & ~n15682 ;
  assign n15684 = \P2_InstQueue_reg[6][0]/NET0131  & ~n3118 ;
  assign n15685 = ~n15683 & ~n15684 ;
  assign n15686 = ~n15673 & n15685 ;
  assign n15687 = ~n15680 & n15686 ;
  assign n15693 = n3499 & ~n15415 ;
  assign n15694 = n3537 & ~n15419 ;
  assign n15695 = ~n15693 & ~n15694 ;
  assign n15696 = \P2_DataWidth_reg[1]/NET0131  & ~n15695 ;
  assign n15688 = ~n3613 & ~n15407 ;
  assign n15689 = \P2_InstQueue_reg[7][0]/NET0131  & ~n3198 ;
  assign n15690 = ~n3575 & n15689 ;
  assign n15691 = ~n15688 & ~n15690 ;
  assign n15697 = ~n3623 & ~n15691 ;
  assign n15698 = ~n15696 & ~n15697 ;
  assign n15699 = n1931 & ~n15698 ;
  assign n15692 = n3087 & ~n15691 ;
  assign n15700 = ~n1498 & n3198 ;
  assign n15701 = ~n15689 & ~n15700 ;
  assign n15702 = n3040 & ~n15701 ;
  assign n15703 = \P2_InstQueue_reg[7][0]/NET0131  & ~n3118 ;
  assign n15704 = ~n15702 & ~n15703 ;
  assign n15705 = ~n15692 & n15704 ;
  assign n15706 = ~n15699 & n15705 ;
  assign n15712 = n3537 & ~n15415 ;
  assign n15713 = n3575 & ~n15419 ;
  assign n15714 = ~n15712 & ~n15713 ;
  assign n15715 = \P2_DataWidth_reg[1]/NET0131  & ~n15714 ;
  assign n15707 = ~n3199 & ~n15407 ;
  assign n15708 = \P2_InstQueue_reg[8][0]/NET0131  & ~n3091 ;
  assign n15709 = ~n3198 & n15708 ;
  assign n15710 = ~n15707 & ~n15709 ;
  assign n15716 = ~n3659 & ~n15710 ;
  assign n15717 = ~n15715 & ~n15716 ;
  assign n15718 = n1931 & ~n15717 ;
  assign n15711 = n3087 & ~n15710 ;
  assign n15719 = ~n1498 & n3091 ;
  assign n15720 = ~n15708 & ~n15719 ;
  assign n15721 = n3040 & ~n15720 ;
  assign n15722 = \P2_InstQueue_reg[8][0]/NET0131  & ~n3118 ;
  assign n15723 = ~n15721 & ~n15722 ;
  assign n15724 = ~n15711 & n15723 ;
  assign n15725 = ~n15718 & n15724 ;
  assign n15731 = n3575 & ~n15415 ;
  assign n15732 = n3198 & ~n15419 ;
  assign n15733 = ~n15731 & ~n15732 ;
  assign n15734 = \P2_DataWidth_reg[1]/NET0131  & ~n15733 ;
  assign n15726 = ~n3105 & ~n15407 ;
  assign n15727 = \P2_InstQueue_reg[9][0]/NET0131  & ~n3098 ;
  assign n15728 = ~n3091 & n15727 ;
  assign n15729 = ~n15726 & ~n15728 ;
  assign n15735 = ~n3695 & ~n15729 ;
  assign n15736 = ~n15734 & ~n15735 ;
  assign n15737 = n1931 & ~n15736 ;
  assign n15730 = n3087 & ~n15729 ;
  assign n15738 = ~n1498 & n3098 ;
  assign n15739 = ~n15727 & ~n15738 ;
  assign n15740 = n3040 & ~n15739 ;
  assign n15741 = \P2_InstQueue_reg[9][0]/NET0131  & ~n3118 ;
  assign n15742 = ~n15740 & ~n15741 ;
  assign n15743 = ~n15730 & n15742 ;
  assign n15744 = ~n15737 & n15743 ;
  assign n15751 = \P2_PhyAddrPointer_reg[4]/NET0131  & n1897 ;
  assign n15752 = ~n11492 & ~n15751 ;
  assign n15753 = n1734 & ~n15752 ;
  assign n15754 = \P2_PhyAddrPointer_reg[4]/NET0131  & ~n8936 ;
  assign n15755 = ~n11477 & ~n15754 ;
  assign n15756 = ~n15753 & n15755 ;
  assign n15757 = n1927 & ~n15756 ;
  assign n15745 = \P2_PhyAddrPointer_reg[1]/NET0131  & \P2_PhyAddrPointer_reg[2]/NET0131  ;
  assign n15746 = \P2_PhyAddrPointer_reg[3]/NET0131  & n15745 ;
  assign n15747 = ~\P2_PhyAddrPointer_reg[4]/NET0131  & ~n15746 ;
  assign n15748 = \P2_PhyAddrPointer_reg[4]/NET0131  & n15746 ;
  assign n15749 = ~n15747 & ~n15748 ;
  assign n15758 = ~\P2_DataWidth_reg[1]/NET0131  & ~n15749 ;
  assign n15759 = ~\P2_PhyAddrPointer_reg[4]/NET0131  & ~n8960 ;
  assign n15760 = ~n8961 & ~n15759 ;
  assign n15761 = \P2_DataWidth_reg[1]/NET0131  & ~n15760 ;
  assign n15762 = n1931 & ~n15761 ;
  assign n15763 = ~n15758 & n15762 ;
  assign n15764 = \P2_PhyAddrPointer_reg[4]/NET0131  & ~n8958 ;
  assign n15750 = n3087 & n15749 ;
  assign n15765 = ~n11468 & ~n15750 ;
  assign n15766 = ~n15764 & n15765 ;
  assign n15767 = ~n15763 & n15766 ;
  assign n15768 = ~n15757 & n15767 ;
  assign n15774 = ~n2345 & n2432 ;
  assign n15775 = \P1_InstAddrPointer_reg[31]/NET0131  & ~n4840 ;
  assign n15776 = ~\P1_InstAddrPointer_reg[1]/NET0131  & ~\P1_InstAddrPointer_reg[31]/NET0131  ;
  assign n15777 = ~n15775 & ~n15776 ;
  assign n15778 = n14087 & n15777 ;
  assign n15779 = ~n3021 & ~n15778 ;
  assign n15780 = n3020 & ~n15779 ;
  assign n15769 = \P1_State2_reg[2]/NET0131  & n3017 ;
  assign n15770 = ~n3028 & ~n15769 ;
  assign n15771 = ~n2435 & n14083 ;
  assign n15772 = n15770 & n15771 ;
  assign n15773 = \P1_InstQueueRd_Addr_reg[2]/NET0131  & ~n15772 ;
  assign n15781 = n2274 & n3042 ;
  assign n15782 = ~n15773 & ~n15781 ;
  assign n15783 = ~n15780 & n15782 ;
  assign n15784 = ~n15774 & n15783 ;
  assign n15785 = \P3_PhyAddrPointer_reg[4]/NET0131  & ~n11965 ;
  assign n15786 = ~n4316 & ~n4337 ;
  assign n15788 = ~n6115 & n15786 ;
  assign n15787 = n6115 & ~n15786 ;
  assign n15789 = n2905 & ~n15787 ;
  assign n15790 = ~n15788 & n15789 ;
  assign n15791 = ~n4001 & ~n4040 ;
  assign n15793 = n6076 & ~n15791 ;
  assign n15792 = ~n6076 & n15791 ;
  assign n15794 = n2904 & ~n15792 ;
  assign n15795 = ~n15793 & n15794 ;
  assign n15796 = ~n15790 & ~n15795 ;
  assign n15797 = ~n15785 & n15796 ;
  assign n15798 = n2453 & ~n15797 ;
  assign n15803 = \P3_PhyAddrPointer_reg[1]/NET0131  & \P3_PhyAddrPointer_reg[2]/NET0131  ;
  assign n15804 = \P3_PhyAddrPointer_reg[3]/NET0131  & n15803 ;
  assign n15805 = ~\P3_PhyAddrPointer_reg[4]/NET0131  & ~n15804 ;
  assign n15806 = \P3_PhyAddrPointer_reg[4]/NET0131  & n15804 ;
  assign n15807 = ~n15805 & ~n15806 ;
  assign n15808 = n10076 & n15807 ;
  assign n15802 = \P3_PhyAddrPointer_reg[4]/NET0131  & ~n9063 ;
  assign n15799 = ~\P3_PhyAddrPointer_reg[4]/NET0131  & ~n9020 ;
  assign n15800 = ~n9021 & ~n15799 ;
  assign n15801 = n2970 & n15800 ;
  assign n15809 = \P3_rEIP_reg[4]/NET0131  & n4412 ;
  assign n15810 = ~n15801 & ~n15809 ;
  assign n15811 = ~n15802 & n15810 ;
  assign n15812 = ~n15808 & n15811 ;
  assign n15813 = ~n15798 & n15812 ;
  assign n15814 = \P1_PhyAddrPointer_reg[4]/NET0131  & n2375 ;
  assign n15815 = ~n11390 & ~n15814 ;
  assign n15816 = n2244 & ~n15815 ;
  assign n15817 = \P1_PhyAddrPointer_reg[4]/NET0131  & ~n10087 ;
  assign n15818 = ~n11398 & ~n15817 ;
  assign n15819 = ~n15816 & n15818 ;
  assign n15820 = n2432 & ~n15819 ;
  assign n15825 = \P1_PhyAddrPointer_reg[1]/NET0131  & \P1_PhyAddrPointer_reg[2]/NET0131  ;
  assign n15826 = \P1_PhyAddrPointer_reg[3]/NET0131  & n15825 ;
  assign n15827 = ~\P1_PhyAddrPointer_reg[4]/NET0131  & ~n15826 ;
  assign n15828 = \P1_PhyAddrPointer_reg[4]/NET0131  & n15826 ;
  assign n15829 = ~n15827 & ~n15828 ;
  assign n15830 = n10133 & n15829 ;
  assign n15824 = \P1_PhyAddrPointer_reg[4]/NET0131  & ~n10136 ;
  assign n15821 = ~\P1_PhyAddrPointer_reg[4]/NET0131  & ~n10092 ;
  assign n15822 = ~n10093 & ~n15821 ;
  assign n15823 = n3148 & n15822 ;
  assign n15831 = ~n11367 & ~n15823 ;
  assign n15832 = ~n15824 & n15831 ;
  assign n15833 = ~n15830 & n15832 ;
  assign n15834 = ~n15820 & n15833 ;
  assign n15836 = ~n2408 & n2432 ;
  assign n15837 = ~\P1_Flush_reg/NET0131  & \P1_InstQueueRd_Addr_reg[1]/NET0131  ;
  assign n15838 = n14087 & ~n15777 ;
  assign n15839 = ~n15837 & ~n15838 ;
  assign n15840 = n3020 & ~n15839 ;
  assign n15835 = \P1_InstQueueRd_Addr_reg[1]/NET0131  & ~n15772 ;
  assign n15841 = ~n2399 & n3042 ;
  assign n15842 = ~n15835 & ~n15841 ;
  assign n15843 = ~n15840 & n15842 ;
  assign n15844 = ~n15836 & n15843 ;
  assign n15846 = ~n2367 & n2432 ;
  assign n15847 = ~\P1_Flush_reg/NET0131  & \P1_InstQueueRd_Addr_reg[3]/NET0131  ;
  assign n15848 = ~n15778 & ~n15847 ;
  assign n15849 = n3020 & ~n15848 ;
  assign n15845 = \P1_InstQueueRd_Addr_reg[3]/NET0131  & ~n15772 ;
  assign n15850 = ~n2348 & n3042 ;
  assign n15851 = ~n15845 & ~n15850 ;
  assign n15852 = ~n15849 & n15851 ;
  assign n15853 = ~n15846 & n15852 ;
  assign n15855 = n2453 & ~n2888 ;
  assign n15856 = ~\P3_Flush_reg/NET0131  & \P3_InstQueueRd_Addr_reg[3]/NET0131  ;
  assign n15857 = ~n15441 & ~n15856 ;
  assign n15858 = n2997 & ~n15857 ;
  assign n15854 = \P3_InstQueueRd_Addr_reg[3]/NET0131  & ~n15435 ;
  assign n15859 = ~n2872 & n2994 ;
  assign n15860 = ~n15854 & ~n15859 ;
  assign n15861 = ~n15858 & n15860 ;
  assign n15862 = ~n15855 & n15861 ;
  assign n15864 = ~n1866 & n1927 ;
  assign n15865 = ~\P2_Flush_reg/NET0131  & \P2_InstQueueRd_Addr_reg[3]/NET0131  ;
  assign n15866 = ~n15453 & ~n15865 ;
  assign n15867 = n2980 & ~n15866 ;
  assign n15863 = \P2_InstQueueRd_Addr_reg[3]/NET0131  & ~n14133 ;
  assign n15868 = n1861 & n3040 ;
  assign n15869 = ~n15863 & ~n15868 ;
  assign n15870 = ~n15867 & n15869 ;
  assign n15871 = ~n15864 & n15870 ;
  assign n15873 = n2453 & ~n2929 ;
  assign n15874 = ~\P3_Flush_reg/NET0131  & \P3_InstQueueRd_Addr_reg[1]/NET0131  ;
  assign n15875 = n14123 & n15440 ;
  assign n15876 = ~n15874 & ~n15875 ;
  assign n15877 = n2997 & ~n15876 ;
  assign n15872 = \P3_InstQueueRd_Addr_reg[1]/NET0131  & ~n15435 ;
  assign n15878 = n2920 & n2994 ;
  assign n15879 = ~n15872 & ~n15878 ;
  assign n15880 = ~n15877 & n15879 ;
  assign n15881 = ~n15873 & n15880 ;
  assign n15883 = ~n1883 & n1927 ;
  assign n15884 = ~\P2_Flush_reg/NET0131  & \P2_InstQueueRd_Addr_reg[1]/NET0131  ;
  assign n15885 = n14135 & ~n15452 ;
  assign n15886 = ~n15884 & ~n15885 ;
  assign n15887 = n2980 & ~n15886 ;
  assign n15882 = \P2_InstQueueRd_Addr_reg[1]/NET0131  & ~n14133 ;
  assign n15888 = ~n1872 & n3040 ;
  assign n15889 = ~n15882 & ~n15888 ;
  assign n15890 = ~n15887 & n15889 ;
  assign n15891 = ~n15883 & n15890 ;
  assign n15892 = \P1_EAX_reg[26]/NET0131  & ~n15402 ;
  assign n15895 = \P1_EAX_reg[0]/NET0131  & \P1_EAX_reg[1]/NET0131  ;
  assign n15896 = \P1_EAX_reg[2]/NET0131  & n15895 ;
  assign n15897 = \P1_EAX_reg[3]/NET0131  & n15896 ;
  assign n15898 = \P1_EAX_reg[4]/NET0131  & n15897 ;
  assign n15899 = \P1_EAX_reg[5]/NET0131  & n15898 ;
  assign n15900 = \P1_EAX_reg[6]/NET0131  & n15899 ;
  assign n15901 = \P1_EAX_reg[7]/NET0131  & n15900 ;
  assign n15902 = \P1_EAX_reg[8]/NET0131  & n15901 ;
  assign n15903 = \P1_EAX_reg[9]/NET0131  & n15902 ;
  assign n15904 = \P1_EAX_reg[10]/NET0131  & n15903 ;
  assign n15905 = \P1_EAX_reg[11]/NET0131  & n15904 ;
  assign n15906 = \P1_EAX_reg[12]/NET0131  & n15905 ;
  assign n15907 = \P1_EAX_reg[13]/NET0131  & n15906 ;
  assign n15908 = \P1_EAX_reg[14]/NET0131  & n15907 ;
  assign n15909 = \P1_EAX_reg[15]/NET0131  & n15908 ;
  assign n15910 = \P1_EAX_reg[16]/NET0131  & n15909 ;
  assign n15911 = \P1_EAX_reg[17]/NET0131  & \P1_EAX_reg[18]/NET0131  ;
  assign n15912 = n15910 & n15911 ;
  assign n15913 = \P1_EAX_reg[19]/NET0131  & n15912 ;
  assign n15914 = \P1_EAX_reg[20]/NET0131  & \P1_EAX_reg[21]/NET0131  ;
  assign n15915 = \P1_EAX_reg[22]/NET0131  & n15914 ;
  assign n15916 = n15913 & n15915 ;
  assign n15917 = \P1_EAX_reg[23]/NET0131  & \P1_EAX_reg[24]/NET0131  ;
  assign n15918 = n15916 & n15917 ;
  assign n15919 = \P1_EAX_reg[25]/NET0131  & n15918 ;
  assign n15920 = n2260 & ~n15919 ;
  assign n15921 = ~n2303 & ~n2377 ;
  assign n15922 = ~n2260 & n2303 ;
  assign n15923 = ~n2331 & n15922 ;
  assign n15924 = ~n2371 & ~n15923 ;
  assign n15925 = ~n15921 & n15924 ;
  assign n15926 = ~n15920 & n15925 ;
  assign n15927 = \P1_EAX_reg[26]/NET0131  & ~n15926 ;
  assign n15934 = ~\P1_EAX_reg[26]/NET0131  & n2260 ;
  assign n15935 = n15919 & n15934 ;
  assign n15928 = ~n15232 & n15263 ;
  assign n15929 = n2337 & ~n15264 ;
  assign n15930 = ~n15928 & n15929 ;
  assign n15931 = n2331 & n15930 ;
  assign n15893 = n2302 & n2377 ;
  assign n15894 = ~n5259 & n15893 ;
  assign n15932 = n2222 & n2377 ;
  assign n15933 = ~n5161 & n15932 ;
  assign n15936 = ~n15894 & ~n15933 ;
  assign n15937 = ~n15931 & n15936 ;
  assign n15938 = ~n15935 & n15937 ;
  assign n15939 = ~n15927 & n15938 ;
  assign n15940 = n2432 & ~n15939 ;
  assign n15941 = ~n15892 & ~n15940 ;
  assign n15942 = ~n2985 & n6809 ;
  assign n15943 = \P2_uWord_reg[12]/NET0131  & ~n15942 ;
  assign n15945 = ~\buf1_reg[12]/NET0131  & n3079 ;
  assign n15944 = ~\buf2_reg[12]/NET0131  & ~n3079 ;
  assign n15946 = ~n1805 & ~n15944 ;
  assign n15947 = ~n15945 & n15946 ;
  assign n15948 = n1742 & n15947 ;
  assign n15951 = ~\P2_EAX_reg[13]/NET0131  & ~\P2_EAX_reg[14]/NET0131  ;
  assign n15952 = ~\P2_EAX_reg[15]/NET0131  & ~\P2_EAX_reg[1]/NET0131  ;
  assign n15959 = n15951 & n15952 ;
  assign n15949 = ~\P2_EAX_reg[0]/NET0131  & ~\P2_EAX_reg[10]/NET0131  ;
  assign n15950 = ~\P2_EAX_reg[11]/NET0131  & ~\P2_EAX_reg[12]/NET0131  ;
  assign n15960 = n15949 & n15950 ;
  assign n15961 = n15959 & n15960 ;
  assign n15955 = ~\P2_EAX_reg[6]/NET0131  & ~\P2_EAX_reg[7]/NET0131  ;
  assign n15956 = ~\P2_EAX_reg[8]/NET0131  & ~\P2_EAX_reg[9]/NET0131  ;
  assign n15957 = n15955 & n15956 ;
  assign n15953 = ~\P2_EAX_reg[2]/NET0131  & ~\P2_EAX_reg[3]/NET0131  ;
  assign n15954 = ~\P2_EAX_reg[4]/NET0131  & ~\P2_EAX_reg[5]/NET0131  ;
  assign n15958 = n15953 & n15954 ;
  assign n15962 = n15957 & n15958 ;
  assign n15963 = n15961 & n15962 ;
  assign n15964 = \P2_EAX_reg[31]/NET0131  & ~n15963 ;
  assign n15965 = \P2_EAX_reg[16]/NET0131  & n15964 ;
  assign n15966 = \P2_EAX_reg[17]/NET0131  & n15965 ;
  assign n15967 = \P2_EAX_reg[18]/NET0131  & n15966 ;
  assign n15968 = \P2_EAX_reg[19]/NET0131  & n15967 ;
  assign n15969 = \P2_EAX_reg[20]/NET0131  & n15968 ;
  assign n15970 = n12654 & n15969 ;
  assign n15971 = n12657 & n15970 ;
  assign n15972 = n12659 & n15971 ;
  assign n15974 = ~\P2_EAX_reg[28]/NET0131  & ~n15972 ;
  assign n15973 = \P2_EAX_reg[28]/NET0131  & n15972 ;
  assign n15975 = n1743 & ~n15973 ;
  assign n15976 = ~n15974 & n15975 ;
  assign n15977 = ~n15948 & ~n15976 ;
  assign n15978 = ~n1810 & ~n15977 ;
  assign n15979 = n1742 & n1805 ;
  assign n15980 = n1743 & ~n1810 ;
  assign n15981 = ~n10236 & ~n15980 ;
  assign n15982 = ~n15979 & ~n15981 ;
  assign n15983 = \P2_uWord_reg[12]/NET0131  & ~n15982 ;
  assign n15984 = ~n15978 & ~n15983 ;
  assign n15985 = n1927 & ~n15984 ;
  assign n15986 = ~n15943 & ~n15985 ;
  assign n15987 = ~n14082 & n15401 ;
  assign n15988 = n14083 & n15987 ;
  assign n15989 = n2222 & n2317 ;
  assign n15990 = n2225 & ~n2301 ;
  assign n15991 = ~n7246 & ~n15990 ;
  assign n15992 = ~n15989 & ~n15991 ;
  assign n15993 = n2432 & ~n15992 ;
  assign n15994 = n15988 & ~n15993 ;
  assign n15995 = \P1_uWord_reg[12]/NET0131  & ~n15994 ;
  assign n15996 = n2222 & ~n2317 ;
  assign n15997 = ~n5197 & n15996 ;
  assign n15998 = \P1_EAX_reg[25]/NET0131  & \P1_EAX_reg[26]/NET0131  ;
  assign n15999 = \P1_EAX_reg[27]/NET0131  & n15998 ;
  assign n16002 = ~\P1_EAX_reg[13]/NET0131  & ~\P1_EAX_reg[14]/NET0131  ;
  assign n16003 = ~\P1_EAX_reg[15]/NET0131  & ~\P1_EAX_reg[1]/NET0131  ;
  assign n16010 = n16002 & n16003 ;
  assign n16000 = ~\P1_EAX_reg[0]/NET0131  & ~\P1_EAX_reg[10]/NET0131  ;
  assign n16001 = ~\P1_EAX_reg[11]/NET0131  & ~\P1_EAX_reg[12]/NET0131  ;
  assign n16011 = n16000 & n16001 ;
  assign n16012 = n16010 & n16011 ;
  assign n16006 = ~\P1_EAX_reg[6]/NET0131  & ~\P1_EAX_reg[7]/NET0131  ;
  assign n16007 = ~\P1_EAX_reg[8]/NET0131  & ~\P1_EAX_reg[9]/NET0131  ;
  assign n16008 = n16006 & n16007 ;
  assign n16004 = ~\P1_EAX_reg[2]/NET0131  & ~\P1_EAX_reg[3]/NET0131  ;
  assign n16005 = ~\P1_EAX_reg[4]/NET0131  & ~\P1_EAX_reg[5]/NET0131  ;
  assign n16009 = n16004 & n16005 ;
  assign n16013 = n16008 & n16009 ;
  assign n16014 = n16012 & n16013 ;
  assign n16015 = \P1_EAX_reg[31]/NET0131  & ~n16014 ;
  assign n16016 = \P1_EAX_reg[16]/NET0131  & n16015 ;
  assign n16017 = \P1_EAX_reg[17]/NET0131  & n16016 ;
  assign n16018 = \P1_EAX_reg[18]/NET0131  & n16017 ;
  assign n16019 = \P1_EAX_reg[19]/NET0131  & n16018 ;
  assign n16020 = n15914 & n16019 ;
  assign n16021 = \P1_EAX_reg[22]/NET0131  & n16020 ;
  assign n16022 = n15917 & n16021 ;
  assign n16023 = n15999 & n16022 ;
  assign n16024 = ~\P1_EAX_reg[28]/NET0131  & ~n16023 ;
  assign n16025 = \P1_EAX_reg[28]/NET0131  & n16023 ;
  assign n16026 = ~n16024 & ~n16025 ;
  assign n16027 = n2225 & n16026 ;
  assign n16028 = ~n15997 & ~n16027 ;
  assign n16029 = ~n2301 & n2432 ;
  assign n16030 = ~n16028 & n16029 ;
  assign n16031 = ~n15995 & ~n16030 ;
  assign n16032 = \P3_EAX_reg[26]/NET0131  & ~n13810 ;
  assign n16037 = ~\P3_EAX_reg[26]/NET0131  & ~n14041 ;
  assign n16038 = n13813 & ~n14042 ;
  assign n16039 = ~n16037 & n16038 ;
  assign n16040 = \P3_EAX_reg[26]/NET0131  & ~n14922 ;
  assign n16033 = ~n13945 & n13976 ;
  assign n16034 = n2847 & ~n13977 ;
  assign n16035 = ~n16033 & n16034 ;
  assign n16036 = n2840 & n16035 ;
  assign n16041 = \buf2_reg[26]/NET0131  & n2820 ;
  assign n16042 = \buf2_reg[10]/NET0131  & n2821 ;
  assign n16043 = ~n16041 & ~n16042 ;
  assign n16044 = n2862 & ~n16043 ;
  assign n16045 = ~n16036 & ~n16044 ;
  assign n16046 = ~n16040 & n16045 ;
  assign n16047 = ~n16039 & n16046 ;
  assign n16048 = n2453 & ~n16047 ;
  assign n16049 = ~n16032 & ~n16048 ;
  assign n16051 = n2748 & ~n14985 ;
  assign n16052 = ~n14954 & ~n16051 ;
  assign n16053 = \P3_EBX_reg[30]/NET0131  & ~n16052 ;
  assign n16050 = n14937 & n14952 ;
  assign n16054 = ~\P3_EBX_reg[30]/NET0131  & n2748 ;
  assign n16055 = n14985 & n16054 ;
  assign n16056 = ~n16050 & ~n16055 ;
  assign n16057 = ~n16053 & n16056 ;
  assign n16058 = n2453 & ~n16057 ;
  assign n16059 = \P3_EBX_reg[30]/NET0131  & ~n13810 ;
  assign n16060 = ~n16058 & ~n16059 ;
  assign n16061 = \P2_EAX_reg[26]/NET0131  & ~n12632 ;
  assign n16066 = ~\P2_EAX_reg[26]/NET0131  & ~n12658 ;
  assign n16067 = n14058 & ~n16066 ;
  assign n16068 = \P2_EAX_reg[26]/NET0131  & ~n12668 ;
  assign n16069 = \P2_EAX_reg[26]/NET0131  & ~n1811 ;
  assign n16077 = n1811 & ~n8597 ;
  assign n16078 = ~n16069 & ~n16077 ;
  assign n16079 = n1803 & ~n16078 ;
  assign n16062 = ~n12800 & n12831 ;
  assign n16063 = n1798 & ~n12832 ;
  assign n16064 = ~n16062 & n16063 ;
  assign n16065 = n1726 & n16064 ;
  assign n16071 = ~\buf1_reg[10]/NET0131  & n3079 ;
  assign n16070 = ~\buf2_reg[10]/NET0131  & ~n3079 ;
  assign n16072 = ~n1805 & ~n16070 ;
  assign n16073 = ~n16071 & n16072 ;
  assign n16074 = ~n1810 & n16073 ;
  assign n16075 = ~n16069 & ~n16074 ;
  assign n16076 = n1742 & ~n16075 ;
  assign n16080 = ~n16065 & ~n16076 ;
  assign n16081 = ~n16079 & n16080 ;
  assign n16082 = ~n16068 & n16081 ;
  assign n16083 = ~n16067 & n16082 ;
  assign n16084 = n1927 & ~n16083 ;
  assign n16085 = ~n16061 & ~n16084 ;
  assign n16086 = ~n2961 & n4417 ;
  assign n16087 = ~n2698 & n2835 ;
  assign n16088 = n2908 & ~n16087 ;
  assign n16089 = n2453 & ~n16088 ;
  assign n16090 = n16086 & ~n16089 ;
  assign n16091 = \P3_uWord_reg[12]/NET0131  & ~n16090 ;
  assign n16092 = \buf2_reg[12]/NET0131  & n2862 ;
  assign n16093 = n2821 & n16092 ;
  assign n16097 = ~\P3_EAX_reg[13]/NET0131  & ~\P3_EAX_reg[14]/NET0131  ;
  assign n16098 = ~\P3_EAX_reg[15]/NET0131  & ~\P3_EAX_reg[1]/NET0131  ;
  assign n16105 = n16097 & n16098 ;
  assign n16095 = ~\P3_EAX_reg[0]/NET0131  & ~\P3_EAX_reg[10]/NET0131  ;
  assign n16096 = ~\P3_EAX_reg[11]/NET0131  & ~\P3_EAX_reg[12]/NET0131  ;
  assign n16106 = n16095 & n16096 ;
  assign n16107 = n16105 & n16106 ;
  assign n16101 = ~\P3_EAX_reg[6]/NET0131  & ~\P3_EAX_reg[7]/NET0131  ;
  assign n16102 = ~\P3_EAX_reg[8]/NET0131  & ~\P3_EAX_reg[9]/NET0131  ;
  assign n16103 = n16101 & n16102 ;
  assign n16099 = ~\P3_EAX_reg[2]/NET0131  & ~\P3_EAX_reg[3]/NET0131  ;
  assign n16100 = ~\P3_EAX_reg[4]/NET0131  & ~\P3_EAX_reg[5]/NET0131  ;
  assign n16104 = n16099 & n16100 ;
  assign n16108 = n16103 & n16104 ;
  assign n16109 = n16107 & n16108 ;
  assign n16110 = \P3_EAX_reg[31]/NET0131  & ~n16109 ;
  assign n16111 = n14032 & n16110 ;
  assign n16112 = \P3_EAX_reg[18]/NET0131  & n16111 ;
  assign n16113 = \P3_EAX_reg[19]/NET0131  & n16112 ;
  assign n16114 = \P3_EAX_reg[20]/NET0131  & n16113 ;
  assign n16115 = \P3_EAX_reg[21]/NET0131  & n16114 ;
  assign n16116 = n14038 & n16115 ;
  assign n16117 = \P3_EAX_reg[24]/NET0131  & n16116 ;
  assign n16118 = \P3_EAX_reg[25]/NET0131  & n16117 ;
  assign n16119 = n14044 & n16118 ;
  assign n16121 = ~\P3_EAX_reg[28]/NET0131  & ~n16119 ;
  assign n16094 = ~n2815 & n2818 ;
  assign n16120 = \P3_EAX_reg[28]/NET0131  & n16119 ;
  assign n16122 = n16094 & ~n16120 ;
  assign n16123 = ~n16121 & n16122 ;
  assign n16124 = ~n16093 & ~n16123 ;
  assign n16125 = n2453 & ~n16124 ;
  assign n16126 = ~n16091 & ~n16125 ;
  assign n16127 = \P2_PhyAddrPointer_reg[3]/NET0131  & n1897 ;
  assign n16128 = ~n12582 & ~n16127 ;
  assign n16129 = n1734 & ~n16128 ;
  assign n16130 = \P2_PhyAddrPointer_reg[3]/NET0131  & ~n8936 ;
  assign n16131 = ~n12590 & ~n16130 ;
  assign n16132 = ~n16129 & n16131 ;
  assign n16133 = n1927 & ~n16132 ;
  assign n16144 = \P2_PhyAddrPointer_reg[3]/NET0131  & n2987 ;
  assign n16141 = ~\P2_PhyAddrPointer_reg[3]/NET0131  & ~n15745 ;
  assign n16142 = ~n15746 & ~n16141 ;
  assign n16143 = n3087 & n16142 ;
  assign n16145 = ~n12564 & ~n16143 ;
  assign n16146 = ~n16144 & n16145 ;
  assign n16134 = \P2_PhyAddrPointer_reg[2]/NET0131  & ~n10965 ;
  assign n16135 = ~\P2_PhyAddrPointer_reg[3]/NET0131  & ~n16134 ;
  assign n16136 = n8960 & ~n10965 ;
  assign n16137 = n1931 & ~n16136 ;
  assign n16138 = ~n16135 & n16137 ;
  assign n16139 = ~n3040 & n8957 ;
  assign n16140 = \P2_PhyAddrPointer_reg[3]/NET0131  & ~n16139 ;
  assign n16147 = ~n16138 & ~n16140 ;
  assign n16148 = n16146 & n16147 ;
  assign n16149 = ~n16133 & n16148 ;
  assign n16150 = \P2_PhyAddrPointer_reg[5]/NET0131  & n1897 ;
  assign n16151 = ~n12615 & ~n16150 ;
  assign n16152 = n1734 & ~n16151 ;
  assign n16153 = \P2_PhyAddrPointer_reg[5]/NET0131  & ~n8936 ;
  assign n16154 = ~n12609 & ~n16153 ;
  assign n16155 = ~n16152 & n16154 ;
  assign n16156 = n1927 & ~n16155 ;
  assign n16160 = ~\P2_PhyAddrPointer_reg[5]/NET0131  & ~n15748 ;
  assign n16161 = ~n13042 & ~n16160 ;
  assign n16162 = n9005 & n16161 ;
  assign n16163 = \P2_PhyAddrPointer_reg[5]/NET0131  & ~n8958 ;
  assign n16157 = ~\P2_PhyAddrPointer_reg[5]/NET0131  & ~n8961 ;
  assign n16158 = ~n8962 & ~n16157 ;
  assign n16159 = n3034 & n16158 ;
  assign n16164 = ~n12600 & ~n16159 ;
  assign n16165 = ~n16163 & n16164 ;
  assign n16166 = ~n16162 & n16165 ;
  assign n16167 = ~n16156 & n16166 ;
  assign n16168 = \P2_PhyAddrPointer_reg[6]/NET0131  & n1897 ;
  assign n16169 = ~n11517 & ~n16168 ;
  assign n16170 = n1734 & ~n16169 ;
  assign n16171 = \P2_PhyAddrPointer_reg[6]/NET0131  & ~n8936 ;
  assign n16172 = ~n11529 & ~n16171 ;
  assign n16173 = ~n16170 & n16172 ;
  assign n16174 = n1927 & ~n16173 ;
  assign n16179 = ~\P2_PhyAddrPointer_reg[6]/NET0131  & ~n13042 ;
  assign n16180 = ~n13043 & ~n16179 ;
  assign n16181 = n3087 & n16180 ;
  assign n16175 = n8962 & ~n10965 ;
  assign n16176 = ~\P2_PhyAddrPointer_reg[6]/NET0131  & ~n16175 ;
  assign n16177 = n1931 & ~n14437 ;
  assign n16178 = ~n16176 & n16177 ;
  assign n16182 = \P2_PhyAddrPointer_reg[6]/NET0131  & ~n8958 ;
  assign n16183 = ~n11503 & ~n16182 ;
  assign n16184 = ~n16178 & n16183 ;
  assign n16185 = ~n16181 & n16184 ;
  assign n16186 = ~n16174 & n16185 ;
  assign n16187 = n2904 & n12527 ;
  assign n16188 = \P3_PhyAddrPointer_reg[3]/NET0131  & ~n11965 ;
  assign n16189 = ~n12512 & ~n16188 ;
  assign n16190 = ~n16187 & n16189 ;
  assign n16191 = n2453 & ~n16190 ;
  assign n16202 = \P3_PhyAddrPointer_reg[3]/NET0131  & n3004 ;
  assign n16199 = ~\P3_PhyAddrPointer_reg[3]/NET0131  & ~n15803 ;
  assign n16200 = ~n15804 & ~n16199 ;
  assign n16201 = n4415 & n16200 ;
  assign n16203 = ~n12498 & ~n16201 ;
  assign n16204 = ~n16202 & n16203 ;
  assign n16192 = \P3_PhyAddrPointer_reg[2]/NET0131  & ~n11124 ;
  assign n16193 = ~\P3_PhyAddrPointer_reg[3]/NET0131  & ~n16192 ;
  assign n16194 = n9020 & ~n11124 ;
  assign n16195 = n2959 & ~n16194 ;
  assign n16196 = ~n16193 & n16195 ;
  assign n16197 = ~n2994 & n9062 ;
  assign n16198 = \P3_PhyAddrPointer_reg[3]/NET0131  & ~n16197 ;
  assign n16205 = ~n16196 & ~n16198 ;
  assign n16206 = n16204 & n16205 ;
  assign n16207 = ~n16191 & n16206 ;
  assign n16213 = ~n2896 & n12544 ;
  assign n16212 = ~\P3_PhyAddrPointer_reg[5]/NET0131  & n2896 ;
  assign n16214 = n2894 & ~n16212 ;
  assign n16215 = ~n16213 & n16214 ;
  assign n16211 = \P3_PhyAddrPointer_reg[5]/NET0131  & ~n9014 ;
  assign n16216 = ~n12555 & ~n16211 ;
  assign n16217 = ~n16215 & n16216 ;
  assign n16218 = n2453 & ~n16217 ;
  assign n16208 = ~\P3_PhyAddrPointer_reg[5]/NET0131  & ~n15806 ;
  assign n16209 = ~n13248 & ~n16208 ;
  assign n16219 = ~\P3_DataWidth_reg[1]/NET0131  & ~n16209 ;
  assign n16220 = ~\P3_PhyAddrPointer_reg[5]/NET0131  & ~n9021 ;
  assign n16221 = ~n9022 & ~n16220 ;
  assign n16222 = \P3_DataWidth_reg[1]/NET0131  & ~n16221 ;
  assign n16223 = n2959 & ~n16222 ;
  assign n16224 = ~n16219 & n16223 ;
  assign n16210 = n4415 & n16209 ;
  assign n16225 = \P3_PhyAddrPointer_reg[5]/NET0131  & ~n9063 ;
  assign n16226 = ~n12539 & ~n16225 ;
  assign n16227 = ~n16210 & n16226 ;
  assign n16228 = ~n16224 & n16227 ;
  assign n16229 = ~n16218 & n16228 ;
  assign n16235 = ~n2896 & ~n11448 ;
  assign n16234 = ~\P3_PhyAddrPointer_reg[6]/NET0131  & n2896 ;
  assign n16236 = n2894 & ~n16234 ;
  assign n16237 = ~n16235 & n16236 ;
  assign n16233 = \P3_PhyAddrPointer_reg[6]/NET0131  & ~n9014 ;
  assign n16238 = ~n11459 & ~n16233 ;
  assign n16239 = ~n16237 & n16238 ;
  assign n16240 = n2453 & ~n16239 ;
  assign n16230 = ~\P3_PhyAddrPointer_reg[6]/NET0131  & ~n13248 ;
  assign n16231 = ~n13249 & ~n16230 ;
  assign n16241 = ~\P3_DataWidth_reg[1]/NET0131  & ~n16231 ;
  assign n16242 = ~\P3_PhyAddrPointer_reg[6]/NET0131  & ~n9022 ;
  assign n16243 = ~n9023 & ~n16242 ;
  assign n16244 = \P3_DataWidth_reg[1]/NET0131  & ~n16243 ;
  assign n16245 = n2959 & ~n16244 ;
  assign n16246 = ~n16241 & n16245 ;
  assign n16232 = n4415 & n16231 ;
  assign n16247 = \P3_PhyAddrPointer_reg[6]/NET0131  & ~n9063 ;
  assign n16248 = ~n11443 & ~n16247 ;
  assign n16249 = ~n16232 & n16248 ;
  assign n16250 = ~n16246 & n16249 ;
  assign n16251 = ~n16240 & n16250 ;
  assign n16252 = \P1_PhyAddrPointer_reg[3]/NET0131  & ~n12209 ;
  assign n16253 = n12461 & ~n16252 ;
  assign n16254 = n2432 & ~n16253 ;
  assign n16265 = \P1_PhyAddrPointer_reg[3]/NET0131  & n3028 ;
  assign n16262 = ~\P1_PhyAddrPointer_reg[3]/NET0131  & ~n15825 ;
  assign n16263 = ~n15826 & ~n16262 ;
  assign n16264 = n5095 & n16263 ;
  assign n16266 = ~n12437 & ~n16264 ;
  assign n16267 = ~n16265 & n16266 ;
  assign n16255 = \P1_PhyAddrPointer_reg[2]/NET0131  & ~n11332 ;
  assign n16256 = ~\P1_PhyAddrPointer_reg[3]/NET0131  & ~n16255 ;
  assign n16257 = n10092 & ~n11332 ;
  assign n16258 = n2436 & ~n16257 ;
  assign n16259 = ~n16256 & n16258 ;
  assign n16260 = ~n3042 & n10135 ;
  assign n16261 = \P1_PhyAddrPointer_reg[3]/NET0131  & ~n16260 ;
  assign n16268 = ~n16259 & ~n16261 ;
  assign n16269 = n16267 & n16268 ;
  assign n16270 = ~n16254 & n16269 ;
  assign n16271 = \P1_PhyAddrPointer_reg[5]/NET0131  & n2375 ;
  assign n16272 = ~n12478 & ~n16271 ;
  assign n16273 = n2244 & ~n16272 ;
  assign n16274 = \P1_PhyAddrPointer_reg[5]/NET0131  & ~n10087 ;
  assign n16275 = ~n12489 & ~n16274 ;
  assign n16276 = ~n16273 & n16275 ;
  assign n16277 = n2432 & ~n16276 ;
  assign n16281 = ~\P1_PhyAddrPointer_reg[5]/NET0131  & ~n15828 ;
  assign n16282 = ~n14587 & ~n16281 ;
  assign n16283 = n10133 & n16282 ;
  assign n16284 = \P1_PhyAddrPointer_reg[5]/NET0131  & ~n10136 ;
  assign n16278 = ~\P1_PhyAddrPointer_reg[5]/NET0131  & ~n10093 ;
  assign n16279 = ~n10094 & ~n16278 ;
  assign n16280 = n3148 & n16279 ;
  assign n16285 = ~n12470 & ~n16280 ;
  assign n16286 = ~n16284 & n16285 ;
  assign n16287 = ~n16283 & n16286 ;
  assign n16288 = ~n16277 & n16287 ;
  assign n16299 = ~n2375 & ~n11425 ;
  assign n16300 = n2244 & ~n16299 ;
  assign n16301 = n10087 & ~n16300 ;
  assign n16302 = \P1_PhyAddrPointer_reg[6]/NET0131  & ~n16301 ;
  assign n16303 = ~n2375 & n16300 ;
  assign n16304 = ~n11434 & ~n16303 ;
  assign n16305 = ~n16302 & n16304 ;
  assign n16306 = n2432 & ~n16305 ;
  assign n16289 = ~\P1_PhyAddrPointer_reg[6]/NET0131  & ~n14587 ;
  assign n16290 = ~n14588 & ~n16289 ;
  assign n16292 = ~\P1_DataWidth_reg[1]/NET0131  & ~n16290 ;
  assign n16293 = ~\P1_PhyAddrPointer_reg[6]/NET0131  & ~n10094 ;
  assign n16294 = ~n10095 & ~n16293 ;
  assign n16295 = \P1_DataWidth_reg[1]/NET0131  & ~n16294 ;
  assign n16296 = n2436 & ~n16295 ;
  assign n16297 = ~n16292 & n16296 ;
  assign n16291 = n5095 & n16290 ;
  assign n16298 = \P1_PhyAddrPointer_reg[6]/NET0131  & ~n10136 ;
  assign n16307 = ~n11407 & ~n16298 ;
  assign n16308 = ~n16291 & n16307 ;
  assign n16309 = ~n16297 & n16308 ;
  assign n16310 = ~n16306 & n16309 ;
  assign n16311 = \P1_EAX_reg[29]/NET0131  & ~n15402 ;
  assign n16319 = n15918 & n15999 ;
  assign n16320 = \P1_EAX_reg[28]/NET0131  & n16319 ;
  assign n16322 = ~\P1_EAX_reg[29]/NET0131  & ~n16320 ;
  assign n16321 = \P1_EAX_reg[29]/NET0131  & n16320 ;
  assign n16323 = n2260 & ~n16321 ;
  assign n16324 = ~n16322 & n16323 ;
  assign n16313 = ~n15328 & n15359 ;
  assign n16314 = n2337 & ~n15360 ;
  assign n16315 = ~n16313 & n16314 ;
  assign n16316 = n2331 & n16315 ;
  assign n16312 = \P1_EAX_reg[29]/NET0131  & ~n15925 ;
  assign n16317 = ~n6908 & n15893 ;
  assign n16318 = ~n5200 & n15932 ;
  assign n16325 = ~n16317 & ~n16318 ;
  assign n16326 = ~n16312 & n16325 ;
  assign n16327 = ~n16316 & n16326 ;
  assign n16328 = ~n16324 & n16327 ;
  assign n16329 = n2432 & ~n16328 ;
  assign n16330 = ~n16311 & ~n16329 ;
  assign n16331 = \P3_EAX_reg[29]/NET0131  & ~n13810 ;
  assign n16335 = ~\P3_EAX_reg[29]/NET0131  & ~n14924 ;
  assign n16336 = n13813 & ~n14925 ;
  assign n16337 = ~n16335 & n16336 ;
  assign n16338 = \P3_EAX_reg[29]/NET0131  & ~n14922 ;
  assign n16332 = ~n14856 & n14887 ;
  assign n16333 = ~n14888 & ~n16332 ;
  assign n16334 = n13812 & n16333 ;
  assign n16339 = \buf2_reg[29]/NET0131  & n2820 ;
  assign n16340 = \buf2_reg[13]/NET0131  & n2821 ;
  assign n16341 = ~n16339 & ~n16340 ;
  assign n16342 = n2862 & ~n16341 ;
  assign n16343 = ~n16334 & ~n16342 ;
  assign n16344 = ~n16338 & n16343 ;
  assign n16345 = ~n16337 & n16344 ;
  assign n16346 = n2453 & ~n16345 ;
  assign n16347 = ~n16331 & ~n16346 ;
  assign n16381 = ~\P2_EAX_reg[15]/NET0131  & ~n12647 ;
  assign n16382 = ~n12648 & n12664 ;
  assign n16383 = ~n16381 & n16382 ;
  assign n16389 = \P2_EAX_reg[15]/NET0131  & ~n12669 ;
  assign n16352 = \P2_InstQueue_reg[3][7]/NET0131  & n1468 ;
  assign n16353 = \P2_InstQueue_reg[10][7]/NET0131  & n1472 ;
  assign n16366 = ~n16352 & ~n16353 ;
  assign n16354 = \P2_InstQueue_reg[1][7]/NET0131  & n1456 ;
  assign n16355 = \P2_InstQueue_reg[14][7]/NET0131  & n1466 ;
  assign n16367 = ~n16354 & ~n16355 ;
  assign n16374 = n16366 & n16367 ;
  assign n16348 = \P2_InstQueue_reg[5][7]/NET0131  & n1450 ;
  assign n16349 = \P2_InstQueue_reg[2][7]/NET0131  & n1464 ;
  assign n16364 = ~n16348 & ~n16349 ;
  assign n16350 = \P2_InstQueue_reg[12][7]/NET0131  & n1459 ;
  assign n16351 = \P2_InstQueue_reg[6][7]/NET0131  & n1474 ;
  assign n16365 = ~n16350 & ~n16351 ;
  assign n16375 = n16364 & n16365 ;
  assign n16376 = n16374 & n16375 ;
  assign n16360 = \P2_InstQueue_reg[15][7]/NET0131  & n1482 ;
  assign n16361 = \P2_InstQueue_reg[4][7]/NET0131  & n1470 ;
  assign n16370 = ~n16360 & ~n16361 ;
  assign n16362 = \P2_InstQueue_reg[8][7]/NET0131  & n1476 ;
  assign n16363 = \P2_InstQueue_reg[11][7]/NET0131  & n1453 ;
  assign n16371 = ~n16362 & ~n16363 ;
  assign n16372 = n16370 & n16371 ;
  assign n16356 = \P2_InstQueue_reg[7][7]/NET0131  & n1447 ;
  assign n16357 = \P2_InstQueue_reg[0][7]/NET0131  & n1478 ;
  assign n16368 = ~n16356 & ~n16357 ;
  assign n16358 = \P2_InstQueue_reg[9][7]/NET0131  & n1461 ;
  assign n16359 = \P2_InstQueue_reg[13][7]/NET0131  & n1480 ;
  assign n16369 = ~n16358 & ~n16359 ;
  assign n16373 = n16368 & n16369 ;
  assign n16377 = n16372 & n16373 ;
  assign n16378 = n16376 & n16377 ;
  assign n16379 = n1798 & ~n16378 ;
  assign n16380 = n1726 & n16379 ;
  assign n16385 = ~\buf1_reg[15]/NET0131  & n3079 ;
  assign n16384 = ~\buf2_reg[15]/NET0131  & ~n3079 ;
  assign n16386 = ~n1805 & ~n16384 ;
  assign n16387 = ~n16385 & n16386 ;
  assign n16388 = n1891 & n16387 ;
  assign n16390 = ~n16380 & ~n16388 ;
  assign n16391 = ~n16389 & n16390 ;
  assign n16392 = ~n16383 & n16391 ;
  assign n16393 = n1927 & ~n16392 ;
  assign n16394 = \P2_EAX_reg[15]/NET0131  & ~n12632 ;
  assign n16395 = ~n16393 & ~n16394 ;
  assign n16396 = \P2_EAX_reg[29]/NET0131  & ~n12632 ;
  assign n16398 = ~\P2_EAX_reg[29]/NET0131  & ~n12661 ;
  assign n16399 = ~n12662 & n12664 ;
  assign n16400 = ~n16398 & n16399 ;
  assign n16401 = ~n12896 & n12927 ;
  assign n16402 = n1798 & ~n12928 ;
  assign n16403 = ~n16401 & n16402 ;
  assign n16404 = n1726 & n16403 ;
  assign n16397 = \P2_EAX_reg[29]/NET0131  & ~n12669 ;
  assign n16405 = \buf2_reg[13]/NET0131  & ~n3079 ;
  assign n16406 = \buf1_reg[13]/NET0131  & n3079 ;
  assign n16407 = ~n16405 & ~n16406 ;
  assign n16408 = n1742 & ~n16407 ;
  assign n16409 = n1803 & ~n10341 ;
  assign n16410 = ~n16408 & ~n16409 ;
  assign n16411 = n1811 & ~n16410 ;
  assign n16412 = ~n16397 & ~n16411 ;
  assign n16413 = ~n16404 & n16412 ;
  assign n16414 = ~n16400 & n16413 ;
  assign n16415 = n1927 & ~n16414 ;
  assign n16416 = ~n16396 & ~n16415 ;
  assign n16421 = ~\P1_EBX_reg[26]/NET0131  & ~n15388 ;
  assign n16422 = n2262 & ~n15389 ;
  assign n16423 = ~n16421 & n16422 ;
  assign n16417 = \P1_EBX_reg[26]/NET0131  & ~n2337 ;
  assign n16418 = ~n15930 & ~n16417 ;
  assign n16419 = n2242 & ~n16418 ;
  assign n16420 = \P1_EBX_reg[26]/NET0131  & n15072 ;
  assign n16424 = ~n16419 & ~n16420 ;
  assign n16425 = ~n16423 & n16424 ;
  assign n16426 = n2432 & ~n16425 ;
  assign n16427 = \P1_EBX_reg[26]/NET0131  & ~n15402 ;
  assign n16428 = ~n16426 & ~n16427 ;
  assign n16433 = ~\P2_EBX_reg[26]/NET0131  & ~n15046 ;
  assign n16434 = n1766 & ~n15047 ;
  assign n16435 = ~n16433 & n16434 ;
  assign n16429 = \P2_EBX_reg[26]/NET0131  & ~n1798 ;
  assign n16430 = ~n16064 & ~n16429 ;
  assign n16431 = n1722 & ~n16430 ;
  assign n16432 = \P2_EBX_reg[26]/NET0131  & n15018 ;
  assign n16436 = ~n16431 & ~n16432 ;
  assign n16437 = ~n16435 & n16436 ;
  assign n16438 = n1927 & ~n16437 ;
  assign n16439 = \P2_EBX_reg[26]/NET0131  & ~n12632 ;
  assign n16440 = ~n16438 & ~n16439 ;
  assign n16441 = \P1_EAX_reg[15]/NET0131  & ~n15402 ;
  assign n16444 = n2260 & ~n15908 ;
  assign n16445 = n15925 & ~n16444 ;
  assign n16446 = \P1_EAX_reg[15]/NET0131  & ~n16445 ;
  assign n16480 = n2260 & n15907 ;
  assign n16481 = \P1_EAX_reg[14]/NET0131  & ~\P1_EAX_reg[15]/NET0131  ;
  assign n16482 = n16480 & n16481 ;
  assign n16442 = n2304 & ~n2317 ;
  assign n16443 = ~n5194 & n16442 ;
  assign n16451 = \P1_InstQueue_reg[6][7]/NET0131  & n1961 ;
  assign n16452 = \P1_InstQueue_reg[2][7]/NET0131  & n1958 ;
  assign n16465 = ~n16451 & ~n16452 ;
  assign n16453 = \P1_InstQueue_reg[15][7]/NET0131  & n1980 ;
  assign n16454 = \P1_InstQueue_reg[9][7]/NET0131  & n1968 ;
  assign n16466 = ~n16453 & ~n16454 ;
  assign n16473 = n16465 & n16466 ;
  assign n16447 = \P1_InstQueue_reg[1][7]/NET0131  & n1982 ;
  assign n16448 = \P1_InstQueue_reg[3][7]/NET0131  & n1966 ;
  assign n16463 = ~n16447 & ~n16448 ;
  assign n16449 = \P1_InstQueue_reg[4][7]/NET0131  & n1970 ;
  assign n16450 = \P1_InstQueue_reg[13][7]/NET0131  & n1949 ;
  assign n16464 = ~n16449 & ~n16450 ;
  assign n16474 = n16463 & n16464 ;
  assign n16475 = n16473 & n16474 ;
  assign n16459 = \P1_InstQueue_reg[11][7]/NET0131  & n1978 ;
  assign n16460 = \P1_InstQueue_reg[7][7]/NET0131  & n1964 ;
  assign n16469 = ~n16459 & ~n16460 ;
  assign n16461 = \P1_InstQueue_reg[5][7]/NET0131  & n1976 ;
  assign n16462 = \P1_InstQueue_reg[10][7]/NET0131  & n1974 ;
  assign n16470 = ~n16461 & ~n16462 ;
  assign n16471 = n16469 & n16470 ;
  assign n16455 = \P1_InstQueue_reg[14][7]/NET0131  & n1953 ;
  assign n16456 = \P1_InstQueue_reg[8][7]/NET0131  & n1972 ;
  assign n16467 = ~n16455 & ~n16456 ;
  assign n16457 = \P1_InstQueue_reg[0][7]/NET0131  & n1955 ;
  assign n16458 = \P1_InstQueue_reg[12][7]/NET0131  & n1946 ;
  assign n16468 = ~n16457 & ~n16458 ;
  assign n16472 = n16467 & n16468 ;
  assign n16476 = n16471 & n16472 ;
  assign n16477 = n16475 & n16476 ;
  assign n16478 = n2337 & ~n16477 ;
  assign n16479 = n2331 & n16478 ;
  assign n16483 = ~n16443 & ~n16479 ;
  assign n16484 = ~n16482 & n16483 ;
  assign n16485 = ~n16446 & n16484 ;
  assign n16486 = n2432 & ~n16485 ;
  assign n16487 = ~n16441 & ~n16486 ;
  assign n16492 = ~n5248 & n5251 ;
  assign n16493 = ~n5252 & ~n16492 ;
  assign n16494 = n5148 & ~n16493 ;
  assign n16489 = n5218 & ~n5272 ;
  assign n16490 = ~n5273 & ~n16489 ;
  assign n16491 = ~n5148 & ~n16490 ;
  assign n16495 = n7703 & ~n16491 ;
  assign n16496 = ~n16494 & n16495 ;
  assign n16502 = ~n5108 & ~n5179 ;
  assign n16497 = \P1_InstQueue_reg[11][0]/NET0131  & ~n5104 ;
  assign n16503 = ~n5107 & n16497 ;
  assign n16504 = ~n16502 & ~n16503 ;
  assign n16501 = ~n5095 & n5153 ;
  assign n16505 = ~n7697 & ~n16501 ;
  assign n16506 = ~n16504 & n16505 ;
  assign n16488 = \P1_InstQueue_reg[11][0]/NET0131  & ~n5291 ;
  assign n16498 = ~n2092 & n5104 ;
  assign n16499 = ~n16497 & ~n16498 ;
  assign n16500 = n3042 & ~n16499 ;
  assign n16507 = ~n16488 & ~n16500 ;
  assign n16508 = ~n16506 & n16507 ;
  assign n16509 = ~n16496 & n16508 ;
  assign n16558 = ~\P2_DataWidth_reg[1]/NET0131  & n1820 ;
  assign n16559 = n15980 & ~n16558 ;
  assign n16560 = ~\P2_EBX_reg[0]/NET0131  & ~\P2_EBX_reg[1]/NET0131  ;
  assign n16561 = ~\P2_EBX_reg[2]/NET0131  & n16560 ;
  assign n16562 = ~\P2_EBX_reg[3]/NET0131  & n16561 ;
  assign n16563 = ~\P2_EBX_reg[4]/NET0131  & n16562 ;
  assign n16564 = ~\P2_EBX_reg[5]/NET0131  & n16563 ;
  assign n16565 = ~\P2_EBX_reg[6]/NET0131  & n16564 ;
  assign n16566 = ~\P2_EBX_reg[7]/NET0131  & n16565 ;
  assign n16567 = ~\P2_EBX_reg[8]/NET0131  & n16566 ;
  assign n16568 = ~\P2_EBX_reg[9]/NET0131  & n16567 ;
  assign n16569 = ~\P2_EBX_reg[10]/NET0131  & n16568 ;
  assign n16570 = ~\P2_EBX_reg[11]/NET0131  & n16569 ;
  assign n16571 = ~\P2_EBX_reg[12]/NET0131  & n16570 ;
  assign n16572 = ~\P2_EBX_reg[13]/NET0131  & n16571 ;
  assign n16573 = ~\P2_EBX_reg[14]/NET0131  & ~\P2_EBX_reg[15]/NET0131  ;
  assign n16574 = ~\P2_EBX_reg[16]/NET0131  & ~\P2_EBX_reg[17]/NET0131  ;
  assign n16575 = n16573 & n16574 ;
  assign n16576 = n16572 & n16575 ;
  assign n16577 = ~\P2_EBX_reg[18]/NET0131  & ~\P2_EBX_reg[19]/NET0131  ;
  assign n16578 = n16576 & n16577 ;
  assign n16579 = ~\P2_EBX_reg[20]/NET0131  & n16578 ;
  assign n16580 = ~\P2_EBX_reg[21]/NET0131  & n16579 ;
  assign n16581 = ~\P2_EBX_reg[22]/NET0131  & ~\P2_EBX_reg[23]/NET0131  ;
  assign n16582 = n16580 & n16581 ;
  assign n16583 = ~\P2_EBX_reg[24]/NET0131  & ~\P2_EBX_reg[25]/NET0131  ;
  assign n16584 = n16582 & n16583 ;
  assign n16585 = ~\P2_EBX_reg[26]/NET0131  & n16584 ;
  assign n16586 = ~\P2_EBX_reg[27]/NET0131  & ~\P2_EBX_reg[28]/NET0131  ;
  assign n16587 = n16585 & n16586 ;
  assign n16588 = ~\P2_EBX_reg[29]/NET0131  & n16587 ;
  assign n16589 = ~n1920 & n10236 ;
  assign n16590 = ~\P2_EBX_reg[30]/NET0131  & n16589 ;
  assign n16591 = n16588 & n16590 ;
  assign n16592 = ~n16559 & ~n16591 ;
  assign n16593 = \P2_EBX_reg[31]/NET0131  & ~n16592 ;
  assign n16524 = \P2_rEIP_reg[1]/NET0131  & \P2_rEIP_reg[2]/NET0131  ;
  assign n16525 = \P2_rEIP_reg[3]/NET0131  & n16524 ;
  assign n16526 = \P2_rEIP_reg[4]/NET0131  & n16525 ;
  assign n16527 = \P2_rEIP_reg[5]/NET0131  & \P2_rEIP_reg[6]/NET0131  ;
  assign n16528 = \P2_rEIP_reg[7]/NET0131  & n16527 ;
  assign n16529 = n16526 & n16528 ;
  assign n16530 = \P2_rEIP_reg[8]/NET0131  & n16529 ;
  assign n16531 = \P2_rEIP_reg[9]/NET0131  & n16530 ;
  assign n16523 = \P2_rEIP_reg[10]/NET0131  & \P2_rEIP_reg[11]/NET0131  ;
  assign n16532 = \P2_rEIP_reg[12]/NET0131  & n16523 ;
  assign n16533 = n16531 & n16532 ;
  assign n16534 = \P2_rEIP_reg[13]/NET0131  & \P2_rEIP_reg[14]/NET0131  ;
  assign n16535 = \P2_rEIP_reg[15]/NET0131  & n16534 ;
  assign n16536 = \P2_rEIP_reg[16]/NET0131  & n16535 ;
  assign n16537 = \P2_rEIP_reg[17]/NET0131  & n16536 ;
  assign n16538 = \P2_rEIP_reg[18]/NET0131  & n16537 ;
  assign n16539 = n16533 & n16538 ;
  assign n16540 = \P2_rEIP_reg[19]/NET0131  & n16539 ;
  assign n16541 = \P2_rEIP_reg[20]/NET0131  & n16540 ;
  assign n16542 = \P2_rEIP_reg[21]/NET0131  & n16541 ;
  assign n16543 = \P2_rEIP_reg[22]/NET0131  & n16542 ;
  assign n16544 = \P2_rEIP_reg[23]/NET0131  & n16543 ;
  assign n16545 = \P2_rEIP_reg[24]/NET0131  & n16544 ;
  assign n16546 = \P2_rEIP_reg[25]/NET0131  & n16545 ;
  assign n16547 = \P2_rEIP_reg[26]/NET0131  & n16546 ;
  assign n16548 = \P2_rEIP_reg[27]/NET0131  & n16547 ;
  assign n16549 = \P2_rEIP_reg[28]/NET0131  & n16548 ;
  assign n16550 = \P2_rEIP_reg[29]/NET0131  & n16549 ;
  assign n16551 = \P2_rEIP_reg[30]/NET0131  & n16550 ;
  assign n16552 = ~n1922 & ~n10236 ;
  assign n16553 = n1920 & ~n16552 ;
  assign n16554 = ~n16551 & n16553 ;
  assign n16555 = ~n1747 & ~n1810 ;
  assign n16556 = ~n16554 & n16555 ;
  assign n16557 = \P2_rEIP_reg[31]/NET0131  & ~n16556 ;
  assign n16594 = ~\P2_rEIP_reg[31]/NET0131  & n16553 ;
  assign n16595 = n16551 & n16594 ;
  assign n16596 = ~n16557 & ~n16595 ;
  assign n16597 = ~n16593 & n16596 ;
  assign n16598 = n1927 & ~n16597 ;
  assign n16513 = \P2_DataWidth_reg[1]/NET0131  & \P2_rEIP_reg[31]/NET0131  ;
  assign n16514 = ~\P2_PhyAddrPointer_reg[0]/NET0131  & \P2_PhyAddrPointer_reg[1]/NET0131  ;
  assign n16515 = n13658 & n16514 ;
  assign n16516 = n8981 & n16515 ;
  assign n16517 = \P2_PhyAddrPointer_reg[25]/NET0131  & n16516 ;
  assign n16518 = n8993 & n16517 ;
  assign n16519 = ~\P2_DataWidth_reg[1]/NET0131  & n16518 ;
  assign n16520 = n9002 & n16519 ;
  assign n16521 = ~n16513 & ~n16520 ;
  assign n16522 = n1931 & ~n16521 ;
  assign n16510 = \P2_PhyAddrPointer_reg[31]/NET0131  & n2987 ;
  assign n16511 = ~n3087 & n16139 ;
  assign n16512 = \P2_rEIP_reg[31]/NET0131  & ~n16511 ;
  assign n16599 = ~n16510 & ~n16512 ;
  assign n16600 = ~n16522 & n16599 ;
  assign n16601 = ~n16598 & n16600 ;
  assign n16604 = n5334 & ~n16493 ;
  assign n16603 = ~n5334 & ~n16490 ;
  assign n16605 = n7755 & ~n16603 ;
  assign n16606 = ~n16604 & n16605 ;
  assign n16612 = ~n5179 & ~n5327 ;
  assign n16607 = \P1_InstQueue_reg[0][0]/NET0131  & ~n5324 ;
  assign n16613 = ~n5326 & n16607 ;
  assign n16614 = ~n16612 & ~n16613 ;
  assign n16611 = ~n5095 & n5338 ;
  assign n16615 = ~n7697 & ~n16611 ;
  assign n16616 = ~n16614 & n16615 ;
  assign n16602 = \P1_InstQueue_reg[0][0]/NET0131  & ~n5291 ;
  assign n16608 = ~n2092 & n5324 ;
  assign n16609 = ~n16607 & ~n16608 ;
  assign n16610 = n3042 & ~n16609 ;
  assign n16617 = ~n16602 & ~n16610 ;
  assign n16618 = ~n16616 & n16617 ;
  assign n16619 = ~n16606 & n16618 ;
  assign n16622 = n5359 & ~n16493 ;
  assign n16621 = ~n5359 & ~n16490 ;
  assign n16623 = n7775 & ~n16621 ;
  assign n16624 = ~n16622 & n16623 ;
  assign n16630 = ~n5179 & ~n5353 ;
  assign n16625 = \P1_InstQueue_reg[10][0]/NET0131  & ~n5107 ;
  assign n16631 = ~n5151 & n16625 ;
  assign n16632 = ~n16630 & ~n16631 ;
  assign n16629 = ~n5095 & n5361 ;
  assign n16633 = ~n7697 & ~n16629 ;
  assign n16634 = ~n16632 & n16633 ;
  assign n16620 = \P1_InstQueue_reg[10][0]/NET0131  & ~n5291 ;
  assign n16626 = ~n2092 & n5107 ;
  assign n16627 = ~n16625 & ~n16626 ;
  assign n16628 = n3042 & ~n16627 ;
  assign n16635 = ~n16620 & ~n16628 ;
  assign n16636 = ~n16634 & n16635 ;
  assign n16637 = ~n16624 & n16636 ;
  assign n16640 = n5151 & ~n16493 ;
  assign n16639 = ~n5151 & ~n16490 ;
  assign n16641 = n7795 & ~n16639 ;
  assign n16642 = ~n16640 & n16641 ;
  assign n16648 = ~n5179 & ~n5378 ;
  assign n16643 = \P1_InstQueue_reg[12][0]/NET0131  & ~n5377 ;
  assign n16649 = ~n5104 & n16643 ;
  assign n16650 = ~n16648 & ~n16649 ;
  assign n16647 = ~n5095 & n5384 ;
  assign n16651 = ~n7697 & ~n16647 ;
  assign n16652 = ~n16650 & n16651 ;
  assign n16638 = \P1_InstQueue_reg[12][0]/NET0131  & ~n5291 ;
  assign n16644 = ~n2092 & n5377 ;
  assign n16645 = ~n16643 & ~n16644 ;
  assign n16646 = n3042 & ~n16645 ;
  assign n16653 = ~n16638 & ~n16646 ;
  assign n16654 = ~n16652 & n16653 ;
  assign n16655 = ~n16642 & n16654 ;
  assign n16658 = n5107 & ~n16493 ;
  assign n16657 = ~n5107 & ~n16490 ;
  assign n16659 = n7815 & ~n16657 ;
  assign n16660 = ~n16658 & n16659 ;
  assign n16666 = ~n5179 & ~n5399 ;
  assign n16661 = \P1_InstQueue_reg[13][0]/NET0131  & ~n5334 ;
  assign n16667 = ~n5377 & n16661 ;
  assign n16668 = ~n16666 & ~n16667 ;
  assign n16665 = ~n5095 & n5405 ;
  assign n16669 = ~n7697 & ~n16665 ;
  assign n16670 = ~n16668 & n16669 ;
  assign n16656 = \P1_InstQueue_reg[13][0]/NET0131  & ~n5291 ;
  assign n16662 = ~n2092 & n5334 ;
  assign n16663 = ~n16661 & ~n16662 ;
  assign n16664 = n3042 & ~n16663 ;
  assign n16671 = ~n16656 & ~n16664 ;
  assign n16672 = ~n16670 & n16671 ;
  assign n16673 = ~n16660 & n16672 ;
  assign n16676 = n5104 & ~n16493 ;
  assign n16675 = ~n5104 & ~n16490 ;
  assign n16677 = n7835 & ~n16675 ;
  assign n16678 = ~n16676 & n16677 ;
  assign n16684 = ~n5179 & ~n5337 ;
  assign n16679 = \P1_InstQueue_reg[14][0]/NET0131  & ~n5336 ;
  assign n16685 = ~n5334 & n16679 ;
  assign n16686 = ~n16684 & ~n16685 ;
  assign n16683 = ~n5095 & n5425 ;
  assign n16687 = ~n7697 & ~n16683 ;
  assign n16688 = ~n16686 & n16687 ;
  assign n16674 = \P1_InstQueue_reg[14][0]/NET0131  & ~n5291 ;
  assign n16680 = ~n2092 & n5336 ;
  assign n16681 = ~n16679 & ~n16680 ;
  assign n16682 = n3042 & ~n16681 ;
  assign n16689 = ~n16674 & ~n16682 ;
  assign n16690 = ~n16688 & n16689 ;
  assign n16691 = ~n16678 & n16690 ;
  assign n16694 = n5377 & ~n16493 ;
  assign n16693 = ~n5377 & ~n16490 ;
  assign n16695 = n7855 & ~n16693 ;
  assign n16696 = ~n16694 & n16695 ;
  assign n16702 = ~n5179 & ~n5440 ;
  assign n16697 = \P1_InstQueue_reg[15][0]/NET0131  & ~n5326 ;
  assign n16703 = ~n5336 & n16697 ;
  assign n16704 = ~n16702 & ~n16703 ;
  assign n16701 = ~n5095 & n5446 ;
  assign n16705 = ~n7697 & ~n16701 ;
  assign n16706 = ~n16704 & n16705 ;
  assign n16692 = \P1_InstQueue_reg[15][0]/NET0131  & ~n5291 ;
  assign n16698 = ~n2092 & n5326 ;
  assign n16699 = ~n16697 & ~n16698 ;
  assign n16700 = n3042 & ~n16699 ;
  assign n16707 = ~n16692 & ~n16700 ;
  assign n16708 = ~n16706 & n16707 ;
  assign n16709 = ~n16696 & n16708 ;
  assign n16712 = n5336 & ~n16493 ;
  assign n16711 = ~n5336 & ~n16490 ;
  assign n16713 = n7875 & ~n16711 ;
  assign n16714 = ~n16712 & n16713 ;
  assign n16720 = ~n5179 & ~n5462 ;
  assign n16715 = \P1_InstQueue_reg[1][0]/NET0131  & ~n5461 ;
  assign n16721 = ~n5324 & n16715 ;
  assign n16722 = ~n16720 & ~n16721 ;
  assign n16719 = ~n5095 & n5468 ;
  assign n16723 = ~n7697 & ~n16719 ;
  assign n16724 = ~n16722 & n16723 ;
  assign n16710 = \P1_InstQueue_reg[1][0]/NET0131  & ~n5291 ;
  assign n16716 = ~n2092 & n5461 ;
  assign n16717 = ~n16715 & ~n16716 ;
  assign n16718 = n3042 & ~n16717 ;
  assign n16725 = ~n16710 & ~n16718 ;
  assign n16726 = ~n16724 & n16725 ;
  assign n16727 = ~n16714 & n16726 ;
  assign n16730 = n5326 & ~n16493 ;
  assign n16729 = ~n5326 & ~n16490 ;
  assign n16731 = n7895 & ~n16729 ;
  assign n16732 = ~n16730 & n16731 ;
  assign n16738 = ~n5179 & ~n5506 ;
  assign n16733 = \P1_InstQueue_reg[2][0]/NET0131  & ~n5484 ;
  assign n16739 = ~n5461 & n16733 ;
  assign n16740 = ~n16738 & ~n16739 ;
  assign n16737 = ~n5095 & n5512 ;
  assign n16741 = ~n7697 & ~n16737 ;
  assign n16742 = ~n16740 & n16741 ;
  assign n16728 = \P1_InstQueue_reg[2][0]/NET0131  & ~n5291 ;
  assign n16734 = ~n2092 & n5484 ;
  assign n16735 = ~n16733 & ~n16734 ;
  assign n16736 = n3042 & ~n16735 ;
  assign n16743 = ~n16728 & ~n16736 ;
  assign n16744 = ~n16742 & n16743 ;
  assign n16745 = ~n16732 & n16744 ;
  assign n16748 = n5324 & ~n16493 ;
  assign n16747 = ~n5324 & ~n16490 ;
  assign n16749 = n7915 & ~n16747 ;
  assign n16750 = ~n16748 & n16749 ;
  assign n16756 = ~n5179 & ~n5485 ;
  assign n16751 = \P1_InstQueue_reg[3][0]/NET0131  & ~n5483 ;
  assign n16757 = ~n5484 & n16751 ;
  assign n16758 = ~n16756 & ~n16757 ;
  assign n16755 = ~n5095 & n5491 ;
  assign n16759 = ~n7697 & ~n16755 ;
  assign n16760 = ~n16758 & n16759 ;
  assign n16746 = \P1_InstQueue_reg[3][0]/NET0131  & ~n5291 ;
  assign n16752 = ~n2092 & n5483 ;
  assign n16753 = ~n16751 & ~n16752 ;
  assign n16754 = n3042 & ~n16753 ;
  assign n16761 = ~n16746 & ~n16754 ;
  assign n16762 = ~n16760 & n16761 ;
  assign n16763 = ~n16750 & n16762 ;
  assign n16766 = n5461 & ~n16493 ;
  assign n16765 = ~n5461 & ~n16490 ;
  assign n16767 = n7935 & ~n16765 ;
  assign n16768 = ~n16766 & n16767 ;
  assign n16774 = ~n5179 & ~n5528 ;
  assign n16769 = \P1_InstQueue_reg[4][0]/NET0131  & ~n5527 ;
  assign n16775 = ~n5483 & n16769 ;
  assign n16776 = ~n16774 & ~n16775 ;
  assign n16773 = ~n5095 & n5534 ;
  assign n16777 = ~n7697 & ~n16773 ;
  assign n16778 = ~n16776 & n16777 ;
  assign n16764 = \P1_InstQueue_reg[4][0]/NET0131  & ~n5291 ;
  assign n16770 = ~n2092 & n5527 ;
  assign n16771 = ~n16769 & ~n16770 ;
  assign n16772 = n3042 & ~n16771 ;
  assign n16779 = ~n16764 & ~n16772 ;
  assign n16780 = ~n16778 & n16779 ;
  assign n16781 = ~n16768 & n16780 ;
  assign n16784 = n5484 & ~n16493 ;
  assign n16783 = ~n5484 & ~n16490 ;
  assign n16785 = n7955 & ~n16783 ;
  assign n16786 = ~n16784 & n16785 ;
  assign n16792 = ~n5179 & ~n5550 ;
  assign n16787 = \P1_InstQueue_reg[5][0]/NET0131  & ~n5549 ;
  assign n16793 = ~n5527 & n16787 ;
  assign n16794 = ~n16792 & ~n16793 ;
  assign n16791 = ~n5095 & n5556 ;
  assign n16795 = ~n7697 & ~n16791 ;
  assign n16796 = ~n16794 & n16795 ;
  assign n16782 = \P1_InstQueue_reg[5][0]/NET0131  & ~n5291 ;
  assign n16788 = ~n2092 & n5549 ;
  assign n16789 = ~n16787 & ~n16788 ;
  assign n16790 = n3042 & ~n16789 ;
  assign n16797 = ~n16782 & ~n16790 ;
  assign n16798 = ~n16796 & n16797 ;
  assign n16799 = ~n16786 & n16798 ;
  assign n16802 = n5483 & ~n16493 ;
  assign n16801 = ~n5483 & ~n16490 ;
  assign n16803 = n7975 & ~n16801 ;
  assign n16804 = ~n16802 & n16803 ;
  assign n16810 = ~n5179 & ~n5572 ;
  assign n16805 = \P1_InstQueue_reg[6][0]/NET0131  & ~n5571 ;
  assign n16811 = ~n5549 & n16805 ;
  assign n16812 = ~n16810 & ~n16811 ;
  assign n16809 = ~n5095 & n5578 ;
  assign n16813 = ~n7697 & ~n16809 ;
  assign n16814 = ~n16812 & n16813 ;
  assign n16800 = \P1_InstQueue_reg[6][0]/NET0131  & ~n5291 ;
  assign n16806 = ~n2092 & n5571 ;
  assign n16807 = ~n16805 & ~n16806 ;
  assign n16808 = n3042 & ~n16807 ;
  assign n16815 = ~n16800 & ~n16808 ;
  assign n16816 = ~n16814 & n16815 ;
  assign n16817 = ~n16804 & n16816 ;
  assign n16820 = n5527 & ~n16493 ;
  assign n16819 = ~n5527 & ~n16490 ;
  assign n16821 = n7995 & ~n16819 ;
  assign n16822 = ~n16820 & n16821 ;
  assign n16828 = ~n5179 & ~n5593 ;
  assign n16823 = \P1_InstQueue_reg[7][0]/NET0131  & ~n5359 ;
  assign n16829 = ~n5571 & n16823 ;
  assign n16830 = ~n16828 & ~n16829 ;
  assign n16827 = ~n5095 & n5599 ;
  assign n16831 = ~n7697 & ~n16827 ;
  assign n16832 = ~n16830 & n16831 ;
  assign n16818 = \P1_InstQueue_reg[7][0]/NET0131  & ~n5291 ;
  assign n16824 = ~n2092 & n5359 ;
  assign n16825 = ~n16823 & ~n16824 ;
  assign n16826 = n3042 & ~n16825 ;
  assign n16833 = ~n16818 & ~n16826 ;
  assign n16834 = ~n16832 & n16833 ;
  assign n16835 = ~n16822 & n16834 ;
  assign n16838 = n5549 & ~n16493 ;
  assign n16837 = ~n5549 & ~n16490 ;
  assign n16839 = n8015 & ~n16837 ;
  assign n16840 = ~n16838 & n16839 ;
  assign n16846 = ~n5179 & ~n5360 ;
  assign n16841 = \P1_InstQueue_reg[8][0]/NET0131  & ~n5148 ;
  assign n16847 = ~n5359 & n16841 ;
  assign n16848 = ~n16846 & ~n16847 ;
  assign n16845 = ~n5095 & n5619 ;
  assign n16849 = ~n7697 & ~n16845 ;
  assign n16850 = ~n16848 & n16849 ;
  assign n16836 = \P1_InstQueue_reg[8][0]/NET0131  & ~n5291 ;
  assign n16842 = ~n2092 & n5148 ;
  assign n16843 = ~n16841 & ~n16842 ;
  assign n16844 = n3042 & ~n16843 ;
  assign n16851 = ~n16836 & ~n16844 ;
  assign n16852 = ~n16850 & n16851 ;
  assign n16853 = ~n16840 & n16852 ;
  assign n16856 = n5571 & ~n16493 ;
  assign n16855 = ~n5571 & ~n16490 ;
  assign n16857 = n8035 & ~n16855 ;
  assign n16858 = ~n16856 & n16857 ;
  assign n16864 = ~n5152 & ~n5179 ;
  assign n16859 = \P1_InstQueue_reg[9][0]/NET0131  & ~n5151 ;
  assign n16865 = ~n5148 & n16859 ;
  assign n16866 = ~n16864 & ~n16865 ;
  assign n16863 = ~n5095 & n5639 ;
  assign n16867 = ~n7697 & ~n16863 ;
  assign n16868 = ~n16866 & n16867 ;
  assign n16854 = \P1_InstQueue_reg[9][0]/NET0131  & ~n5291 ;
  assign n16860 = ~n2092 & n5151 ;
  assign n16861 = ~n16859 & ~n16860 ;
  assign n16862 = n3042 & ~n16861 ;
  assign n16869 = ~n16854 & ~n16862 ;
  assign n16870 = ~n16868 & n16869 ;
  assign n16871 = ~n16858 & n16870 ;
  assign n16873 = \P1_Datao_reg[24]/NET0131  & ~n2313 ;
  assign n16874 = \P1_EAX_reg[23]/NET0131  & n16021 ;
  assign n16875 = ~\P1_EAX_reg[24]/NET0131  & ~n16874 ;
  assign n16876 = n2225 & ~n16022 ;
  assign n16877 = ~n16875 & n16876 ;
  assign n16878 = n2312 & n16877 ;
  assign n16879 = ~n16873 & ~n16878 ;
  assign n16880 = n2432 & ~n16879 ;
  assign n16872 = \P1_uWord_reg[8]/NET0131  & n2440 ;
  assign n16882 = \P1_State2_reg[1]/NET0131  & n2444 ;
  assign n16881 = ~n2438 & n3017 ;
  assign n16883 = ~n3026 & ~n16881 ;
  assign n16884 = ~n16882 & n16883 ;
  assign n16885 = \P1_Datao_reg[24]/NET0131  & ~n16884 ;
  assign n16886 = ~n16872 & ~n16885 ;
  assign n16887 = ~n16880 & n16886 ;
  assign n16890 = \datao[24]_pad  & ~n2833 ;
  assign n16891 = ~\P3_EAX_reg[24]/NET0131  & ~n16116 ;
  assign n16892 = n2818 & ~n16117 ;
  assign n16893 = ~n16891 & n16892 ;
  assign n16894 = n2816 & n16893 ;
  assign n16895 = ~n16890 & ~n16894 ;
  assign n16896 = n2453 & ~n16895 ;
  assign n16888 = ~\P3_State2_reg[0]/NET0131  & n2996 ;
  assign n16889 = \P3_uWord_reg[8]/NET0131  & n16888 ;
  assign n16897 = \P3_State2_reg[1]/NET0131  & n2451 ;
  assign n16898 = ~n2961 & ~n16897 ;
  assign n16899 = n10074 & n16898 ;
  assign n16900 = \datao[24]_pad  & ~n16899 ;
  assign n16901 = ~n16889 & ~n16900 ;
  assign n16902 = ~n16896 & n16901 ;
  assign n16904 = \datao[28]_pad  & ~n2833 ;
  assign n16905 = ~n2786 & n16123 ;
  assign n16906 = ~n16904 & ~n16905 ;
  assign n16907 = n2453 & ~n16906 ;
  assign n16903 = \P3_uWord_reg[12]/NET0131  & n16888 ;
  assign n16908 = \datao[28]_pad  & ~n16899 ;
  assign n16909 = ~n16903 & ~n16908 ;
  assign n16910 = ~n16907 & n16909 ;
  assign n16912 = \P1_Datao_reg[28]/NET0131  & ~n2313 ;
  assign n16913 = n2426 & n16026 ;
  assign n16914 = ~n16912 & ~n16913 ;
  assign n16915 = n2432 & ~n16914 ;
  assign n16911 = \P1_uWord_reg[12]/NET0131  & n2440 ;
  assign n16916 = \P1_Datao_reg[28]/NET0131  & ~n16884 ;
  assign n16917 = ~n16911 & ~n16916 ;
  assign n16918 = ~n16915 & n16917 ;
  assign n16921 = n1813 & n1819 ;
  assign n16922 = n7639 & ~n16921 ;
  assign n16923 = \P2_EAX_reg[23]/NET0131  & n15970 ;
  assign n16924 = ~\P2_EAX_reg[24]/NET0131  & ~n16923 ;
  assign n16925 = \P2_EAX_reg[24]/NET0131  & n16923 ;
  assign n16926 = ~n16924 & ~n16925 ;
  assign n16927 = ~n1819 & ~n16926 ;
  assign n16928 = n15980 & ~n16927 ;
  assign n16929 = n16922 & ~n16928 ;
  assign n16930 = \P2_Datao_reg[24]/NET0131  & ~n16929 ;
  assign n16931 = n1922 & ~n16927 ;
  assign n16932 = ~n16930 & ~n16931 ;
  assign n16933 = n1927 & ~n16932 ;
  assign n16919 = ~\P2_State2_reg[0]/NET0131  & n2979 ;
  assign n16920 = \P2_uWord_reg[8]/NET0131  & n16919 ;
  assign n16934 = \P2_State2_reg[1]/NET0131  & n1925 ;
  assign n16935 = ~n2985 & ~n16934 ;
  assign n16936 = n3125 & n16935 ;
  assign n16937 = \P2_Datao_reg[24]/NET0131  & ~n16936 ;
  assign n16938 = ~n16920 & ~n16937 ;
  assign n16939 = ~n16933 & n16938 ;
  assign n16941 = ~n1810 & n1828 ;
  assign n16942 = \P2_Datao_reg[28]/NET0131  & ~n16941 ;
  assign n16943 = n1921 & n15976 ;
  assign n16944 = ~n16942 & ~n16943 ;
  assign n16945 = n1927 & ~n16944 ;
  assign n16940 = \P2_uWord_reg[12]/NET0131  & n16919 ;
  assign n16946 = \P2_Datao_reg[28]/NET0131  & ~n16936 ;
  assign n16947 = ~n16940 & ~n16946 ;
  assign n16948 = ~n16945 & n16947 ;
  assign n16949 = n1927 & ~n15982 ;
  assign n16950 = n15942 & ~n16949 ;
  assign n16951 = \P2_uWord_reg[8]/NET0131  & ~n16950 ;
  assign n16952 = n1743 & n16926 ;
  assign n16954 = ~\buf1_reg[8]/NET0131  & n3079 ;
  assign n16953 = ~\buf2_reg[8]/NET0131  & ~n3079 ;
  assign n16955 = ~n1805 & ~n16953 ;
  assign n16956 = ~n16954 & n16955 ;
  assign n16957 = n1742 & n16956 ;
  assign n16958 = ~n16952 & ~n16957 ;
  assign n16959 = ~n1810 & n1927 ;
  assign n16960 = ~n16958 & n16959 ;
  assign n16961 = ~n16951 & ~n16960 ;
  assign n16962 = \P1_uWord_reg[8]/NET0131  & ~n15994 ;
  assign n16963 = ~n5173 & n15996 ;
  assign n16964 = ~n16877 & ~n16963 ;
  assign n16965 = n16029 & ~n16964 ;
  assign n16966 = ~n16962 & ~n16965 ;
  assign n16967 = n2432 & ~n15925 ;
  assign n16968 = n15402 & ~n16967 ;
  assign n16969 = \P1_EAX_reg[2]/NET0131  & ~n16968 ;
  assign n16972 = n2337 & ~n4675 ;
  assign n16973 = n2331 & n16972 ;
  assign n16970 = n2377 & ~n5188 ;
  assign n16971 = ~n2303 & n16970 ;
  assign n16974 = ~\P1_EAX_reg[2]/NET0131  & ~n15895 ;
  assign n16975 = ~n15896 & ~n16974 ;
  assign n16976 = n2260 & n16975 ;
  assign n16977 = ~n16971 & ~n16976 ;
  assign n16978 = ~n16973 & n16977 ;
  assign n16979 = n2432 & ~n16978 ;
  assign n16980 = ~n16969 & ~n16979 ;
  assign n16981 = \P3_EAX_reg[10]/NET0131  & ~n13810 ;
  assign n16983 = n13813 & ~n14026 ;
  assign n16984 = n14922 & ~n16983 ;
  assign n16985 = \P3_EAX_reg[10]/NET0131  & ~n16984 ;
  assign n16982 = \buf2_reg[10]/NET0131  & n2857 ;
  assign n16990 = \P3_InstQueue_reg[0][2]/NET0131  & n2488 ;
  assign n16991 = \P3_InstQueue_reg[9][2]/NET0131  & n2460 ;
  assign n17004 = ~n16990 & ~n16991 ;
  assign n16992 = \P3_InstQueue_reg[14][2]/NET0131  & n2472 ;
  assign n16993 = \P3_InstQueue_reg[10][2]/NET0131  & n2476 ;
  assign n17005 = ~n16992 & ~n16993 ;
  assign n17012 = n17004 & n17005 ;
  assign n16986 = \P3_InstQueue_reg[5][2]/NET0131  & n2480 ;
  assign n16987 = \P3_InstQueue_reg[6][2]/NET0131  & n2469 ;
  assign n17002 = ~n16986 & ~n16987 ;
  assign n16988 = \P3_InstQueue_reg[2][2]/NET0131  & n2482 ;
  assign n16989 = \P3_InstQueue_reg[15][2]/NET0131  & n2478 ;
  assign n17003 = ~n16988 & ~n16989 ;
  assign n17013 = n17002 & n17003 ;
  assign n17014 = n17012 & n17013 ;
  assign n16998 = \P3_InstQueue_reg[4][2]/NET0131  & n2466 ;
  assign n16999 = \P3_InstQueue_reg[12][2]/NET0131  & n2464 ;
  assign n17008 = ~n16998 & ~n16999 ;
  assign n17000 = \P3_InstQueue_reg[3][2]/NET0131  & n2456 ;
  assign n17001 = \P3_InstQueue_reg[1][2]/NET0131  & n2484 ;
  assign n17009 = ~n17000 & ~n17001 ;
  assign n17010 = n17008 & n17009 ;
  assign n16994 = \P3_InstQueue_reg[7][2]/NET0131  & n2492 ;
  assign n16995 = \P3_InstQueue_reg[13][2]/NET0131  & n2486 ;
  assign n17006 = ~n16994 & ~n16995 ;
  assign n16996 = \P3_InstQueue_reg[11][2]/NET0131  & n2490 ;
  assign n16997 = \P3_InstQueue_reg[8][2]/NET0131  & n2474 ;
  assign n17007 = ~n16996 & ~n16997 ;
  assign n17011 = n17006 & n17007 ;
  assign n17015 = n17010 & n17011 ;
  assign n17016 = n17014 & n17015 ;
  assign n17017 = n13812 & ~n17016 ;
  assign n17018 = n14025 & n16983 ;
  assign n17019 = ~n17017 & ~n17018 ;
  assign n17020 = ~n16982 & n17019 ;
  assign n17021 = ~n16985 & n17020 ;
  assign n17022 = n2453 & ~n17021 ;
  assign n17023 = ~n16981 & ~n17022 ;
  assign n17024 = \P1_EAX_reg[3]/NET0131  & ~n16968 ;
  assign n17027 = n2337 & ~n4639 ;
  assign n17028 = n2331 & n17027 ;
  assign n17025 = n2377 & ~n5167 ;
  assign n17026 = ~n2303 & n17025 ;
  assign n17029 = ~\P1_EAX_reg[3]/NET0131  & ~n15896 ;
  assign n17030 = ~n15897 & ~n17029 ;
  assign n17031 = n2260 & n17030 ;
  assign n17032 = ~n17026 & ~n17031 ;
  assign n17033 = ~n17028 & n17032 ;
  assign n17034 = n2432 & ~n17033 ;
  assign n17035 = ~n17024 & ~n17034 ;
  assign n17036 = \P3_EAX_reg[11]/NET0131  & ~n13810 ;
  assign n17039 = \P3_EAX_reg[11]/NET0131  & ~n16984 ;
  assign n17044 = \P3_InstQueue_reg[0][3]/NET0131  & n2488 ;
  assign n17045 = \P3_InstQueue_reg[11][3]/NET0131  & n2490 ;
  assign n17058 = ~n17044 & ~n17045 ;
  assign n17046 = \P3_InstQueue_reg[12][3]/NET0131  & n2464 ;
  assign n17047 = \P3_InstQueue_reg[2][3]/NET0131  & n2482 ;
  assign n17059 = ~n17046 & ~n17047 ;
  assign n17066 = n17058 & n17059 ;
  assign n17040 = \P3_InstQueue_reg[5][3]/NET0131  & n2480 ;
  assign n17041 = \P3_InstQueue_reg[15][3]/NET0131  & n2478 ;
  assign n17056 = ~n17040 & ~n17041 ;
  assign n17042 = \P3_InstQueue_reg[10][3]/NET0131  & n2476 ;
  assign n17043 = \P3_InstQueue_reg[14][3]/NET0131  & n2472 ;
  assign n17057 = ~n17042 & ~n17043 ;
  assign n17067 = n17056 & n17057 ;
  assign n17068 = n17066 & n17067 ;
  assign n17052 = \P3_InstQueue_reg[4][3]/NET0131  & n2466 ;
  assign n17053 = \P3_InstQueue_reg[6][3]/NET0131  & n2469 ;
  assign n17062 = ~n17052 & ~n17053 ;
  assign n17054 = \P3_InstQueue_reg[1][3]/NET0131  & n2484 ;
  assign n17055 = \P3_InstQueue_reg[3][3]/NET0131  & n2456 ;
  assign n17063 = ~n17054 & ~n17055 ;
  assign n17064 = n17062 & n17063 ;
  assign n17048 = \P3_InstQueue_reg[8][3]/NET0131  & n2474 ;
  assign n17049 = \P3_InstQueue_reg[13][3]/NET0131  & n2486 ;
  assign n17060 = ~n17048 & ~n17049 ;
  assign n17050 = \P3_InstQueue_reg[9][3]/NET0131  & n2460 ;
  assign n17051 = \P3_InstQueue_reg[7][3]/NET0131  & n2492 ;
  assign n17061 = ~n17050 & ~n17051 ;
  assign n17065 = n17060 & n17061 ;
  assign n17069 = n17064 & n17065 ;
  assign n17070 = n17068 & n17069 ;
  assign n17071 = n13812 & ~n17070 ;
  assign n17037 = n13813 & ~n14027 ;
  assign n17038 = n14026 & n17037 ;
  assign n17072 = ~n2822 & n14048 ;
  assign n17073 = ~n17038 & ~n17072 ;
  assign n17074 = ~n17071 & n17073 ;
  assign n17075 = ~n17039 & n17074 ;
  assign n17076 = n2453 & ~n17075 ;
  assign n17077 = ~n17036 & ~n17076 ;
  assign n17078 = \P3_EAX_reg[12]/NET0131  & ~n13810 ;
  assign n17111 = ~n13816 & ~n17037 ;
  assign n17112 = \P3_EAX_reg[12]/NET0131  & ~n17111 ;
  assign n17113 = \P3_EAX_reg[12]/NET0131  & ~n2862 ;
  assign n17114 = ~n16092 & ~n17113 ;
  assign n17115 = ~n2822 & ~n17114 ;
  assign n17083 = \P3_InstQueue_reg[0][4]/NET0131  & n2488 ;
  assign n17084 = \P3_InstQueue_reg[11][4]/NET0131  & n2490 ;
  assign n17097 = ~n17083 & ~n17084 ;
  assign n17085 = \P3_InstQueue_reg[12][4]/NET0131  & n2464 ;
  assign n17086 = \P3_InstQueue_reg[2][4]/NET0131  & n2482 ;
  assign n17098 = ~n17085 & ~n17086 ;
  assign n17105 = n17097 & n17098 ;
  assign n17079 = \P3_InstQueue_reg[5][4]/NET0131  & n2480 ;
  assign n17080 = \P3_InstQueue_reg[15][4]/NET0131  & n2478 ;
  assign n17095 = ~n17079 & ~n17080 ;
  assign n17081 = \P3_InstQueue_reg[10][4]/NET0131  & n2476 ;
  assign n17082 = \P3_InstQueue_reg[14][4]/NET0131  & n2472 ;
  assign n17096 = ~n17081 & ~n17082 ;
  assign n17106 = n17095 & n17096 ;
  assign n17107 = n17105 & n17106 ;
  assign n17091 = \P3_InstQueue_reg[4][4]/NET0131  & n2466 ;
  assign n17092 = \P3_InstQueue_reg[6][4]/NET0131  & n2469 ;
  assign n17101 = ~n17091 & ~n17092 ;
  assign n17093 = \P3_InstQueue_reg[1][4]/NET0131  & n2484 ;
  assign n17094 = \P3_InstQueue_reg[3][4]/NET0131  & n2456 ;
  assign n17102 = ~n17093 & ~n17094 ;
  assign n17103 = n17101 & n17102 ;
  assign n17087 = \P3_InstQueue_reg[8][4]/NET0131  & n2474 ;
  assign n17088 = \P3_InstQueue_reg[13][4]/NET0131  & n2486 ;
  assign n17099 = ~n17087 & ~n17088 ;
  assign n17089 = \P3_InstQueue_reg[9][4]/NET0131  & n2460 ;
  assign n17090 = \P3_InstQueue_reg[7][4]/NET0131  & n2492 ;
  assign n17100 = ~n17089 & ~n17090 ;
  assign n17104 = n17099 & n17100 ;
  assign n17108 = n17103 & n17104 ;
  assign n17109 = n17107 & n17108 ;
  assign n17110 = n13812 & ~n17109 ;
  assign n17116 = ~\P3_EAX_reg[12]/NET0131  & n13813 ;
  assign n17117 = n14027 & n17116 ;
  assign n17118 = ~n17110 & ~n17117 ;
  assign n17119 = ~n17115 & n17118 ;
  assign n17120 = ~n17112 & n17119 ;
  assign n17121 = n2453 & ~n17120 ;
  assign n17122 = ~n17078 & ~n17121 ;
  assign n17123 = n2453 & ~n14922 ;
  assign n17124 = n13810 & ~n17123 ;
  assign n17125 = \P3_EAX_reg[13]/NET0131  & ~n17124 ;
  assign n17159 = ~\P3_EAX_reg[13]/NET0131  & ~n14028 ;
  assign n17160 = n13813 & ~n14029 ;
  assign n17161 = ~n17159 & n17160 ;
  assign n17130 = \P3_InstQueue_reg[0][5]/NET0131  & n2488 ;
  assign n17131 = \P3_InstQueue_reg[11][5]/NET0131  & n2490 ;
  assign n17144 = ~n17130 & ~n17131 ;
  assign n17132 = \P3_InstQueue_reg[12][5]/NET0131  & n2464 ;
  assign n17133 = \P3_InstQueue_reg[2][5]/NET0131  & n2482 ;
  assign n17145 = ~n17132 & ~n17133 ;
  assign n17152 = n17144 & n17145 ;
  assign n17126 = \P3_InstQueue_reg[5][5]/NET0131  & n2480 ;
  assign n17127 = \P3_InstQueue_reg[15][5]/NET0131  & n2478 ;
  assign n17142 = ~n17126 & ~n17127 ;
  assign n17128 = \P3_InstQueue_reg[10][5]/NET0131  & n2476 ;
  assign n17129 = \P3_InstQueue_reg[14][5]/NET0131  & n2472 ;
  assign n17143 = ~n17128 & ~n17129 ;
  assign n17153 = n17142 & n17143 ;
  assign n17154 = n17152 & n17153 ;
  assign n17138 = \P3_InstQueue_reg[4][5]/NET0131  & n2466 ;
  assign n17139 = \P3_InstQueue_reg[6][5]/NET0131  & n2469 ;
  assign n17148 = ~n17138 & ~n17139 ;
  assign n17140 = \P3_InstQueue_reg[1][5]/NET0131  & n2484 ;
  assign n17141 = \P3_InstQueue_reg[3][5]/NET0131  & n2456 ;
  assign n17149 = ~n17140 & ~n17141 ;
  assign n17150 = n17148 & n17149 ;
  assign n17134 = \P3_InstQueue_reg[8][5]/NET0131  & n2474 ;
  assign n17135 = \P3_InstQueue_reg[13][5]/NET0131  & n2486 ;
  assign n17146 = ~n17134 & ~n17135 ;
  assign n17136 = \P3_InstQueue_reg[9][5]/NET0131  & n2460 ;
  assign n17137 = \P3_InstQueue_reg[7][5]/NET0131  & n2492 ;
  assign n17147 = ~n17136 & ~n17137 ;
  assign n17151 = n17146 & n17147 ;
  assign n17155 = n17150 & n17151 ;
  assign n17156 = n17154 & n17155 ;
  assign n17157 = n13812 & ~n17156 ;
  assign n17158 = \buf2_reg[13]/NET0131  & n2857 ;
  assign n17162 = ~n17157 & ~n17158 ;
  assign n17163 = ~n17161 & n17162 ;
  assign n17164 = n2453 & ~n17163 ;
  assign n17165 = ~n17125 & ~n17164 ;
  assign n17166 = \P3_EAX_reg[14]/NET0131  & ~n17124 ;
  assign n17200 = ~\P3_EAX_reg[14]/NET0131  & ~n14029 ;
  assign n17201 = n13813 & ~n14030 ;
  assign n17202 = ~n17200 & n17201 ;
  assign n17167 = \buf2_reg[14]/NET0131  & n2857 ;
  assign n17172 = \P3_InstQueue_reg[0][6]/NET0131  & n2488 ;
  assign n17173 = \P3_InstQueue_reg[11][6]/NET0131  & n2490 ;
  assign n17186 = ~n17172 & ~n17173 ;
  assign n17174 = \P3_InstQueue_reg[12][6]/NET0131  & n2464 ;
  assign n17175 = \P3_InstQueue_reg[2][6]/NET0131  & n2482 ;
  assign n17187 = ~n17174 & ~n17175 ;
  assign n17194 = n17186 & n17187 ;
  assign n17168 = \P3_InstQueue_reg[5][6]/NET0131  & n2480 ;
  assign n17169 = \P3_InstQueue_reg[15][6]/NET0131  & n2478 ;
  assign n17184 = ~n17168 & ~n17169 ;
  assign n17170 = \P3_InstQueue_reg[10][6]/NET0131  & n2476 ;
  assign n17171 = \P3_InstQueue_reg[14][6]/NET0131  & n2472 ;
  assign n17185 = ~n17170 & ~n17171 ;
  assign n17195 = n17184 & n17185 ;
  assign n17196 = n17194 & n17195 ;
  assign n17180 = \P3_InstQueue_reg[4][6]/NET0131  & n2466 ;
  assign n17181 = \P3_InstQueue_reg[6][6]/NET0131  & n2469 ;
  assign n17190 = ~n17180 & ~n17181 ;
  assign n17182 = \P3_InstQueue_reg[1][6]/NET0131  & n2484 ;
  assign n17183 = \P3_InstQueue_reg[3][6]/NET0131  & n2456 ;
  assign n17191 = ~n17182 & ~n17183 ;
  assign n17192 = n17190 & n17191 ;
  assign n17176 = \P3_InstQueue_reg[8][6]/NET0131  & n2474 ;
  assign n17177 = \P3_InstQueue_reg[13][6]/NET0131  & n2486 ;
  assign n17188 = ~n17176 & ~n17177 ;
  assign n17178 = \P3_InstQueue_reg[9][6]/NET0131  & n2460 ;
  assign n17179 = \P3_InstQueue_reg[7][6]/NET0131  & n2492 ;
  assign n17189 = ~n17178 & ~n17179 ;
  assign n17193 = n17188 & n17189 ;
  assign n17197 = n17192 & n17193 ;
  assign n17198 = n17196 & n17197 ;
  assign n17199 = n13812 & ~n17198 ;
  assign n17203 = ~n17167 & ~n17199 ;
  assign n17204 = ~n17202 & n17203 ;
  assign n17205 = n2453 & ~n17204 ;
  assign n17206 = ~n17166 & ~n17205 ;
  assign n17207 = \P3_EAX_reg[15]/NET0131  & ~n17124 ;
  assign n17210 = ~\P3_EAX_reg[15]/NET0131  & ~n14030 ;
  assign n17211 = n13813 & ~n14031 ;
  assign n17212 = ~n17210 & n17211 ;
  assign n17208 = \buf2_reg[15]/NET0131  & n2862 ;
  assign n17209 = ~n2822 & n17208 ;
  assign n17217 = \P3_InstQueue_reg[0][7]/NET0131  & n2488 ;
  assign n17218 = \P3_InstQueue_reg[11][7]/NET0131  & n2490 ;
  assign n17231 = ~n17217 & ~n17218 ;
  assign n17219 = \P3_InstQueue_reg[12][7]/NET0131  & n2464 ;
  assign n17220 = \P3_InstQueue_reg[2][7]/NET0131  & n2482 ;
  assign n17232 = ~n17219 & ~n17220 ;
  assign n17239 = n17231 & n17232 ;
  assign n17213 = \P3_InstQueue_reg[5][7]/NET0131  & n2480 ;
  assign n17214 = \P3_InstQueue_reg[15][7]/NET0131  & n2478 ;
  assign n17229 = ~n17213 & ~n17214 ;
  assign n17215 = \P3_InstQueue_reg[10][7]/NET0131  & n2476 ;
  assign n17216 = \P3_InstQueue_reg[14][7]/NET0131  & n2472 ;
  assign n17230 = ~n17215 & ~n17216 ;
  assign n17240 = n17229 & n17230 ;
  assign n17241 = n17239 & n17240 ;
  assign n17225 = \P3_InstQueue_reg[4][7]/NET0131  & n2466 ;
  assign n17226 = \P3_InstQueue_reg[6][7]/NET0131  & n2469 ;
  assign n17235 = ~n17225 & ~n17226 ;
  assign n17227 = \P3_InstQueue_reg[1][7]/NET0131  & n2484 ;
  assign n17228 = \P3_InstQueue_reg[3][7]/NET0131  & n2456 ;
  assign n17236 = ~n17227 & ~n17228 ;
  assign n17237 = n17235 & n17236 ;
  assign n17221 = \P3_InstQueue_reg[8][7]/NET0131  & n2474 ;
  assign n17222 = \P3_InstQueue_reg[13][7]/NET0131  & n2486 ;
  assign n17233 = ~n17221 & ~n17222 ;
  assign n17223 = \P3_InstQueue_reg[9][7]/NET0131  & n2460 ;
  assign n17224 = \P3_InstQueue_reg[7][7]/NET0131  & n2492 ;
  assign n17234 = ~n17223 & ~n17224 ;
  assign n17238 = n17233 & n17234 ;
  assign n17242 = n17237 & n17238 ;
  assign n17243 = n17241 & n17242 ;
  assign n17244 = n13812 & ~n17243 ;
  assign n17245 = ~n17209 & ~n17244 ;
  assign n17246 = ~n17212 & n17245 ;
  assign n17247 = n2453 & ~n17246 ;
  assign n17248 = ~n17207 & ~n17247 ;
  assign n17249 = \P1_EAX_reg[4]/NET0131  & ~n16968 ;
  assign n17250 = ~n5140 & n16442 ;
  assign n17251 = n2337 & ~n4607 ;
  assign n17252 = n2331 & n17251 ;
  assign n17253 = ~\P1_EAX_reg[4]/NET0131  & ~n15897 ;
  assign n17254 = ~n15898 & ~n17253 ;
  assign n17255 = n2260 & n17254 ;
  assign n17256 = ~n17252 & ~n17255 ;
  assign n17257 = ~n17250 & n17256 ;
  assign n17258 = n2432 & ~n17257 ;
  assign n17259 = ~n17249 & ~n17258 ;
  assign n17260 = \P3_EAX_reg[1]/NET0131  & ~n13810 ;
  assign n17263 = ~\P3_EAX_reg[0]/NET0131  & n13813 ;
  assign n17264 = n14922 & ~n17263 ;
  assign n17265 = \P3_EAX_reg[1]/NET0131  & ~n17264 ;
  assign n17266 = ~n3930 & n13812 ;
  assign n17261 = \buf2_reg[1]/NET0131  & n2862 ;
  assign n17262 = ~n2822 & n17261 ;
  assign n17267 = \P3_EAX_reg[0]/NET0131  & ~\P3_EAX_reg[1]/NET0131  ;
  assign n17268 = n13813 & n17267 ;
  assign n17269 = ~n17262 & ~n17268 ;
  assign n17270 = ~n17266 & n17269 ;
  assign n17271 = ~n17265 & n17270 ;
  assign n17272 = n2453 & ~n17271 ;
  assign n17273 = ~n17260 & ~n17272 ;
  assign n17274 = \P1_EAX_reg[5]/NET0131  & ~n16968 ;
  assign n17275 = ~n5164 & n16442 ;
  assign n17276 = n2337 & ~n4573 ;
  assign n17277 = n2331 & n17276 ;
  assign n17278 = ~\P1_EAX_reg[5]/NET0131  & ~n15898 ;
  assign n17279 = ~n15899 & ~n17278 ;
  assign n17280 = n2260 & n17279 ;
  assign n17281 = ~n17277 & ~n17280 ;
  assign n17282 = ~n17275 & n17281 ;
  assign n17283 = n2432 & ~n17282 ;
  assign n17284 = ~n17274 & ~n17283 ;
  assign n17285 = \P3_EAX_reg[2]/NET0131  & ~n17124 ;
  assign n17286 = \buf2_reg[2]/NET0131  & n2857 ;
  assign n17287 = ~n3896 & n13812 ;
  assign n17288 = ~\P3_EAX_reg[2]/NET0131  & ~n14017 ;
  assign n17289 = ~n14018 & ~n17288 ;
  assign n17290 = n13813 & n17289 ;
  assign n17291 = ~n17287 & ~n17290 ;
  assign n17292 = ~n17286 & n17291 ;
  assign n17293 = n2453 & ~n17292 ;
  assign n17294 = ~n17285 & ~n17293 ;
  assign n17295 = \P3_EAX_reg[3]/NET0131  & ~n17124 ;
  assign n17296 = \buf2_reg[3]/NET0131  & n2857 ;
  assign n17297 = ~n4032 & n13812 ;
  assign n17298 = ~\P3_EAX_reg[3]/NET0131  & ~n14018 ;
  assign n17299 = ~n14019 & ~n17298 ;
  assign n17300 = n13813 & n17299 ;
  assign n17301 = ~n17297 & ~n17300 ;
  assign n17302 = ~n17296 & n17301 ;
  assign n17303 = n2453 & ~n17302 ;
  assign n17304 = ~n17295 & ~n17303 ;
  assign n17305 = \P1_EAX_reg[7]/NET0131  & ~n16968 ;
  assign n17306 = ~n5176 & n16442 ;
  assign n17307 = n2337 & ~n4453 ;
  assign n17308 = n2331 & n17307 ;
  assign n17309 = ~\P1_EAX_reg[7]/NET0131  & ~n15900 ;
  assign n17310 = ~n15901 & ~n17309 ;
  assign n17311 = n2260 & n17310 ;
  assign n17312 = ~n17308 & ~n17311 ;
  assign n17313 = ~n17306 & n17312 ;
  assign n17314 = n2432 & ~n17313 ;
  assign n17315 = ~n17305 & ~n17314 ;
  assign n17316 = \P3_EAX_reg[4]/NET0131  & ~n17124 ;
  assign n17317 = \buf2_reg[4]/NET0131  & n2857 ;
  assign n17318 = ~n4000 & n13812 ;
  assign n17319 = ~\P3_EAX_reg[4]/NET0131  & ~n14019 ;
  assign n17320 = ~n14020 & ~n17319 ;
  assign n17321 = n13813 & n17320 ;
  assign n17322 = ~n17318 & ~n17321 ;
  assign n17323 = ~n17317 & n17322 ;
  assign n17324 = n2453 & ~n17323 ;
  assign n17325 = ~n17316 & ~n17324 ;
  assign n17326 = \P3_EAX_reg[5]/NET0131  & ~n17124 ;
  assign n17327 = \buf2_reg[5]/NET0131  & n2857 ;
  assign n17328 = ~n3830 & n13812 ;
  assign n17329 = ~\P3_EAX_reg[5]/NET0131  & ~n14020 ;
  assign n17330 = ~n14021 & ~n17329 ;
  assign n17331 = n13813 & n17330 ;
  assign n17332 = ~n17328 & ~n17331 ;
  assign n17333 = ~n17327 & n17332 ;
  assign n17334 = n2453 & ~n17333 ;
  assign n17335 = ~n17326 & ~n17334 ;
  assign n17336 = \P3_EAX_reg[6]/NET0131  & ~n17124 ;
  assign n17337 = \buf2_reg[6]/NET0131  & n2857 ;
  assign n17338 = ~n3864 & n13812 ;
  assign n17339 = ~\P3_EAX_reg[6]/NET0131  & ~n14021 ;
  assign n17340 = ~n14022 & ~n17339 ;
  assign n17341 = n13813 & n17340 ;
  assign n17342 = ~n17338 & ~n17341 ;
  assign n17343 = ~n17337 & n17342 ;
  assign n17344 = n2453 & ~n17343 ;
  assign n17345 = ~n17336 & ~n17344 ;
  assign n17346 = \P3_EAX_reg[7]/NET0131  & ~n17124 ;
  assign n17347 = \buf2_reg[7]/NET0131  & n2857 ;
  assign n17348 = ~n3753 & n13812 ;
  assign n17349 = ~\P3_EAX_reg[7]/NET0131  & ~n14022 ;
  assign n17350 = ~n14023 & ~n17349 ;
  assign n17351 = n13813 & n17350 ;
  assign n17352 = ~n17348 & ~n17351 ;
  assign n17353 = ~n17347 & n17352 ;
  assign n17354 = n2453 & ~n17353 ;
  assign n17355 = ~n17346 & ~n17354 ;
  assign n17356 = \P3_EAX_reg[8]/NET0131  & ~n17124 ;
  assign n17357 = \buf2_reg[8]/NET0131  & n2857 ;
  assign n17362 = \P3_InstQueue_reg[0][0]/NET0131  & n2488 ;
  assign n17363 = \P3_InstQueue_reg[11][0]/NET0131  & n2490 ;
  assign n17376 = ~n17362 & ~n17363 ;
  assign n17364 = \P3_InstQueue_reg[12][0]/NET0131  & n2464 ;
  assign n17365 = \P3_InstQueue_reg[2][0]/NET0131  & n2482 ;
  assign n17377 = ~n17364 & ~n17365 ;
  assign n17384 = n17376 & n17377 ;
  assign n17358 = \P3_InstQueue_reg[5][0]/NET0131  & n2480 ;
  assign n17359 = \P3_InstQueue_reg[15][0]/NET0131  & n2478 ;
  assign n17374 = ~n17358 & ~n17359 ;
  assign n17360 = \P3_InstQueue_reg[10][0]/NET0131  & n2476 ;
  assign n17361 = \P3_InstQueue_reg[14][0]/NET0131  & n2472 ;
  assign n17375 = ~n17360 & ~n17361 ;
  assign n17385 = n17374 & n17375 ;
  assign n17386 = n17384 & n17385 ;
  assign n17370 = \P3_InstQueue_reg[4][0]/NET0131  & n2466 ;
  assign n17371 = \P3_InstQueue_reg[6][0]/NET0131  & n2469 ;
  assign n17380 = ~n17370 & ~n17371 ;
  assign n17372 = \P3_InstQueue_reg[1][0]/NET0131  & n2484 ;
  assign n17373 = \P3_InstQueue_reg[3][0]/NET0131  & n2456 ;
  assign n17381 = ~n17372 & ~n17373 ;
  assign n17382 = n17380 & n17381 ;
  assign n17366 = \P3_InstQueue_reg[8][0]/NET0131  & n2474 ;
  assign n17367 = \P3_InstQueue_reg[13][0]/NET0131  & n2486 ;
  assign n17378 = ~n17366 & ~n17367 ;
  assign n17368 = \P3_InstQueue_reg[9][0]/NET0131  & n2460 ;
  assign n17369 = \P3_InstQueue_reg[7][0]/NET0131  & n2492 ;
  assign n17379 = ~n17368 & ~n17369 ;
  assign n17383 = n17378 & n17379 ;
  assign n17387 = n17382 & n17383 ;
  assign n17388 = n17386 & n17387 ;
  assign n17389 = n13812 & ~n17388 ;
  assign n17390 = ~\P3_EAX_reg[8]/NET0131  & ~n14023 ;
  assign n17391 = ~n14024 & ~n17390 ;
  assign n17392 = n13813 & n17391 ;
  assign n17393 = ~n17389 & ~n17392 ;
  assign n17394 = ~n17357 & n17393 ;
  assign n17395 = n2453 & ~n17394 ;
  assign n17396 = ~n17356 & ~n17395 ;
  assign n17397 = \P3_EAX_reg[9]/NET0131  & ~n17124 ;
  assign n17398 = \buf2_reg[9]/NET0131  & n2857 ;
  assign n17403 = \P3_InstQueue_reg[0][1]/NET0131  & n2488 ;
  assign n17404 = \P3_InstQueue_reg[9][1]/NET0131  & n2460 ;
  assign n17417 = ~n17403 & ~n17404 ;
  assign n17405 = \P3_InstQueue_reg[2][1]/NET0131  & n2482 ;
  assign n17406 = \P3_InstQueue_reg[10][1]/NET0131  & n2476 ;
  assign n17418 = ~n17405 & ~n17406 ;
  assign n17425 = n17417 & n17418 ;
  assign n17399 = \P3_InstQueue_reg[5][1]/NET0131  & n2480 ;
  assign n17400 = \P3_InstQueue_reg[6][1]/NET0131  & n2469 ;
  assign n17415 = ~n17399 & ~n17400 ;
  assign n17401 = \P3_InstQueue_reg[11][1]/NET0131  & n2490 ;
  assign n17402 = \P3_InstQueue_reg[15][1]/NET0131  & n2478 ;
  assign n17416 = ~n17401 & ~n17402 ;
  assign n17426 = n17415 & n17416 ;
  assign n17427 = n17425 & n17426 ;
  assign n17411 = \P3_InstQueue_reg[4][1]/NET0131  & n2466 ;
  assign n17412 = \P3_InstQueue_reg[14][1]/NET0131  & n2472 ;
  assign n17421 = ~n17411 & ~n17412 ;
  assign n17413 = \P3_InstQueue_reg[1][1]/NET0131  & n2484 ;
  assign n17414 = \P3_InstQueue_reg[3][1]/NET0131  & n2456 ;
  assign n17422 = ~n17413 & ~n17414 ;
  assign n17423 = n17421 & n17422 ;
  assign n17407 = \P3_InstQueue_reg[7][1]/NET0131  & n2492 ;
  assign n17408 = \P3_InstQueue_reg[13][1]/NET0131  & n2486 ;
  assign n17419 = ~n17407 & ~n17408 ;
  assign n17409 = \P3_InstQueue_reg[8][1]/NET0131  & n2474 ;
  assign n17410 = \P3_InstQueue_reg[12][1]/NET0131  & n2464 ;
  assign n17420 = ~n17409 & ~n17410 ;
  assign n17424 = n17419 & n17420 ;
  assign n17428 = n17423 & n17424 ;
  assign n17429 = n17427 & n17428 ;
  assign n17430 = n13812 & ~n17429 ;
  assign n17431 = ~\P3_EAX_reg[9]/NET0131  & ~n14024 ;
  assign n17432 = ~n14025 & ~n17431 ;
  assign n17433 = n13813 & n17432 ;
  assign n17434 = ~n17430 & ~n17433 ;
  assign n17435 = ~n17398 & n17434 ;
  assign n17436 = n2453 & ~n17435 ;
  assign n17437 = ~n17397 & ~n17436 ;
  assign n17438 = n1927 & ~n12669 ;
  assign n17439 = n12632 & ~n17438 ;
  assign n17440 = \P2_EAX_reg[0]/NET0131  & ~n17439 ;
  assign n17444 = n1811 & ~n15407 ;
  assign n17445 = ~n1804 & n17444 ;
  assign n17441 = ~\P2_EAX_reg[0]/NET0131  & n12664 ;
  assign n17442 = n1798 & ~n6368 ;
  assign n17443 = n1726 & n17442 ;
  assign n17446 = ~n17441 & ~n17443 ;
  assign n17447 = ~n17445 & n17446 ;
  assign n17448 = n1927 & ~n17447 ;
  assign n17449 = ~n17440 & ~n17448 ;
  assign n17450 = \P3_EBX_reg[29]/NET0131  & ~n13810 ;
  assign n17453 = \P3_EBX_reg[26]/NET0131  & n14981 ;
  assign n17454 = \P3_EBX_reg[27]/NET0131  & n17453 ;
  assign n17455 = \P3_EBX_reg[28]/NET0131  & n16051 ;
  assign n17456 = n17454 & n17455 ;
  assign n17451 = \P3_EBX_reg[29]/NET0131  & ~n16052 ;
  assign n17452 = n14952 & n16333 ;
  assign n17457 = ~n17451 & ~n17452 ;
  assign n17458 = ~n17456 & n17457 ;
  assign n17459 = n2453 & ~n17458 ;
  assign n17460 = ~n17450 & ~n17459 ;
  assign n17461 = \P1_EAX_reg[8]/NET0131  & ~n16968 ;
  assign n17468 = \P1_InstQueue_reg[5][0]/NET0131  & n1976 ;
  assign n17469 = \P1_InstQueue_reg[10][0]/NET0131  & n1974 ;
  assign n17482 = ~n17468 & ~n17469 ;
  assign n17470 = \P1_InstQueue_reg[15][0]/NET0131  & n1980 ;
  assign n17471 = \P1_InstQueue_reg[8][0]/NET0131  & n1972 ;
  assign n17483 = ~n17470 & ~n17471 ;
  assign n17490 = n17482 & n17483 ;
  assign n17464 = \P1_InstQueue_reg[1][0]/NET0131  & n1982 ;
  assign n17465 = \P1_InstQueue_reg[13][0]/NET0131  & n1949 ;
  assign n17480 = ~n17464 & ~n17465 ;
  assign n17466 = \P1_InstQueue_reg[12][0]/NET0131  & n1946 ;
  assign n17467 = \P1_InstQueue_reg[3][0]/NET0131  & n1966 ;
  assign n17481 = ~n17466 & ~n17467 ;
  assign n17491 = n17480 & n17481 ;
  assign n17492 = n17490 & n17491 ;
  assign n17476 = \P1_InstQueue_reg[4][0]/NET0131  & n1970 ;
  assign n17477 = \P1_InstQueue_reg[14][0]/NET0131  & n1953 ;
  assign n17486 = ~n17476 & ~n17477 ;
  assign n17478 = \P1_InstQueue_reg[9][0]/NET0131  & n1968 ;
  assign n17479 = \P1_InstQueue_reg[11][0]/NET0131  & n1978 ;
  assign n17487 = ~n17478 & ~n17479 ;
  assign n17488 = n17486 & n17487 ;
  assign n17472 = \P1_InstQueue_reg[6][0]/NET0131  & n1961 ;
  assign n17473 = \P1_InstQueue_reg[2][0]/NET0131  & n1958 ;
  assign n17484 = ~n17472 & ~n17473 ;
  assign n17474 = \P1_InstQueue_reg[0][0]/NET0131  & n1955 ;
  assign n17475 = \P1_InstQueue_reg[7][0]/NET0131  & n1964 ;
  assign n17485 = ~n17474 & ~n17475 ;
  assign n17489 = n17484 & n17485 ;
  assign n17493 = n17488 & n17489 ;
  assign n17494 = n17492 & n17493 ;
  assign n17495 = n2337 & ~n17494 ;
  assign n17496 = n2331 & n17495 ;
  assign n17462 = n2377 & ~n5173 ;
  assign n17463 = ~n2303 & n17462 ;
  assign n17497 = ~\P1_EAX_reg[8]/NET0131  & ~n15901 ;
  assign n17498 = ~n15902 & ~n17497 ;
  assign n17499 = n2260 & n17498 ;
  assign n17500 = ~n17463 & ~n17499 ;
  assign n17501 = ~n17496 & n17500 ;
  assign n17502 = n2432 & ~n17501 ;
  assign n17503 = ~n17461 & ~n17502 ;
  assign n17504 = \P2_EAX_reg[10]/NET0131  & ~n12632 ;
  assign n17506 = ~n12643 & n12664 ;
  assign n17507 = n12669 & ~n17506 ;
  assign n17508 = \P2_EAX_reg[10]/NET0131  & ~n17507 ;
  assign n17505 = n1891 & n16073 ;
  assign n17513 = \P2_InstQueue_reg[3][2]/NET0131  & n1468 ;
  assign n17514 = \P2_InstQueue_reg[10][2]/NET0131  & n1472 ;
  assign n17527 = ~n17513 & ~n17514 ;
  assign n17515 = \P2_InstQueue_reg[1][2]/NET0131  & n1456 ;
  assign n17516 = \P2_InstQueue_reg[14][2]/NET0131  & n1466 ;
  assign n17528 = ~n17515 & ~n17516 ;
  assign n17535 = n17527 & n17528 ;
  assign n17509 = \P2_InstQueue_reg[5][2]/NET0131  & n1450 ;
  assign n17510 = \P2_InstQueue_reg[2][2]/NET0131  & n1464 ;
  assign n17525 = ~n17509 & ~n17510 ;
  assign n17511 = \P2_InstQueue_reg[12][2]/NET0131  & n1459 ;
  assign n17512 = \P2_InstQueue_reg[6][2]/NET0131  & n1474 ;
  assign n17526 = ~n17511 & ~n17512 ;
  assign n17536 = n17525 & n17526 ;
  assign n17537 = n17535 & n17536 ;
  assign n17521 = \P2_InstQueue_reg[15][2]/NET0131  & n1482 ;
  assign n17522 = \P2_InstQueue_reg[4][2]/NET0131  & n1470 ;
  assign n17531 = ~n17521 & ~n17522 ;
  assign n17523 = \P2_InstQueue_reg[8][2]/NET0131  & n1476 ;
  assign n17524 = \P2_InstQueue_reg[11][2]/NET0131  & n1453 ;
  assign n17532 = ~n17523 & ~n17524 ;
  assign n17533 = n17531 & n17532 ;
  assign n17517 = \P2_InstQueue_reg[7][2]/NET0131  & n1447 ;
  assign n17518 = \P2_InstQueue_reg[0][2]/NET0131  & n1478 ;
  assign n17529 = ~n17517 & ~n17518 ;
  assign n17519 = \P2_InstQueue_reg[9][2]/NET0131  & n1461 ;
  assign n17520 = \P2_InstQueue_reg[13][2]/NET0131  & n1480 ;
  assign n17530 = ~n17519 & ~n17520 ;
  assign n17534 = n17529 & n17530 ;
  assign n17538 = n17533 & n17534 ;
  assign n17539 = n17537 & n17538 ;
  assign n17540 = n1798 & ~n17539 ;
  assign n17541 = n1726 & n17540 ;
  assign n17542 = n12642 & n17506 ;
  assign n17543 = ~n17541 & ~n17542 ;
  assign n17544 = ~n17505 & n17543 ;
  assign n17545 = ~n17508 & n17544 ;
  assign n17546 = n1927 & ~n17545 ;
  assign n17547 = ~n17504 & ~n17546 ;
  assign n17548 = \P2_EAX_reg[11]/NET0131  & ~n12632 ;
  assign n17550 = \P2_EAX_reg[11]/NET0131  & ~n17507 ;
  assign n17549 = ~n14069 & n14771 ;
  assign n17555 = \P2_InstQueue_reg[3][3]/NET0131  & n1468 ;
  assign n17556 = \P2_InstQueue_reg[0][3]/NET0131  & n1478 ;
  assign n17569 = ~n17555 & ~n17556 ;
  assign n17557 = \P2_InstQueue_reg[1][3]/NET0131  & n1456 ;
  assign n17558 = \P2_InstQueue_reg[13][3]/NET0131  & n1480 ;
  assign n17570 = ~n17557 & ~n17558 ;
  assign n17577 = n17569 & n17570 ;
  assign n17551 = \P2_InstQueue_reg[5][3]/NET0131  & n1450 ;
  assign n17552 = \P2_InstQueue_reg[10][3]/NET0131  & n1472 ;
  assign n17567 = ~n17551 & ~n17552 ;
  assign n17553 = \P2_InstQueue_reg[15][3]/NET0131  & n1482 ;
  assign n17554 = \P2_InstQueue_reg[4][3]/NET0131  & n1470 ;
  assign n17568 = ~n17553 & ~n17554 ;
  assign n17578 = n17567 & n17568 ;
  assign n17579 = n17577 & n17578 ;
  assign n17563 = \P2_InstQueue_reg[12][3]/NET0131  & n1459 ;
  assign n17564 = \P2_InstQueue_reg[2][3]/NET0131  & n1464 ;
  assign n17573 = ~n17563 & ~n17564 ;
  assign n17565 = \P2_InstQueue_reg[7][3]/NET0131  & n1447 ;
  assign n17566 = \P2_InstQueue_reg[11][3]/NET0131  & n1453 ;
  assign n17574 = ~n17565 & ~n17566 ;
  assign n17575 = n17573 & n17574 ;
  assign n17559 = \P2_InstQueue_reg[6][3]/NET0131  & n1474 ;
  assign n17560 = \P2_InstQueue_reg[8][3]/NET0131  & n1476 ;
  assign n17571 = ~n17559 & ~n17560 ;
  assign n17561 = \P2_InstQueue_reg[9][3]/NET0131  & n1461 ;
  assign n17562 = \P2_InstQueue_reg[14][3]/NET0131  & n1466 ;
  assign n17572 = ~n17561 & ~n17562 ;
  assign n17576 = n17571 & n17572 ;
  assign n17580 = n17575 & n17576 ;
  assign n17581 = n17579 & n17580 ;
  assign n17582 = n1798 & ~n17581 ;
  assign n17583 = n1726 & n17582 ;
  assign n17584 = ~\P2_EAX_reg[11]/NET0131  & n12643 ;
  assign n17585 = n12664 & n17584 ;
  assign n17586 = ~n17583 & ~n17585 ;
  assign n17587 = ~n17549 & n17586 ;
  assign n17588 = ~n17550 & n17587 ;
  assign n17589 = n1927 & ~n17588 ;
  assign n17590 = ~n17548 & ~n17589 ;
  assign n17591 = \P2_EAX_reg[12]/NET0131  & ~n12632 ;
  assign n17593 = ~n12645 & n12664 ;
  assign n17594 = n12669 & ~n17593 ;
  assign n17595 = \P2_EAX_reg[12]/NET0131  & ~n17594 ;
  assign n17596 = n12644 & n17593 ;
  assign n17592 = n1891 & n15947 ;
  assign n17601 = \P2_InstQueue_reg[3][4]/NET0131  & n1468 ;
  assign n17602 = \P2_InstQueue_reg[10][4]/NET0131  & n1472 ;
  assign n17615 = ~n17601 & ~n17602 ;
  assign n17603 = \P2_InstQueue_reg[1][4]/NET0131  & n1456 ;
  assign n17604 = \P2_InstQueue_reg[14][4]/NET0131  & n1466 ;
  assign n17616 = ~n17603 & ~n17604 ;
  assign n17623 = n17615 & n17616 ;
  assign n17597 = \P2_InstQueue_reg[5][4]/NET0131  & n1450 ;
  assign n17598 = \P2_InstQueue_reg[2][4]/NET0131  & n1464 ;
  assign n17613 = ~n17597 & ~n17598 ;
  assign n17599 = \P2_InstQueue_reg[12][4]/NET0131  & n1459 ;
  assign n17600 = \P2_InstQueue_reg[6][4]/NET0131  & n1474 ;
  assign n17614 = ~n17599 & ~n17600 ;
  assign n17624 = n17613 & n17614 ;
  assign n17625 = n17623 & n17624 ;
  assign n17609 = \P2_InstQueue_reg[15][4]/NET0131  & n1482 ;
  assign n17610 = \P2_InstQueue_reg[4][4]/NET0131  & n1470 ;
  assign n17619 = ~n17609 & ~n17610 ;
  assign n17611 = \P2_InstQueue_reg[8][4]/NET0131  & n1476 ;
  assign n17612 = \P2_InstQueue_reg[11][4]/NET0131  & n1453 ;
  assign n17620 = ~n17611 & ~n17612 ;
  assign n17621 = n17619 & n17620 ;
  assign n17605 = \P2_InstQueue_reg[7][4]/NET0131  & n1447 ;
  assign n17606 = \P2_InstQueue_reg[0][4]/NET0131  & n1478 ;
  assign n17617 = ~n17605 & ~n17606 ;
  assign n17607 = \P2_InstQueue_reg[9][4]/NET0131  & n1461 ;
  assign n17608 = \P2_InstQueue_reg[13][4]/NET0131  & n1480 ;
  assign n17618 = ~n17607 & ~n17608 ;
  assign n17622 = n17617 & n17618 ;
  assign n17626 = n17621 & n17622 ;
  assign n17627 = n17625 & n17626 ;
  assign n17628 = n1798 & ~n17627 ;
  assign n17629 = n1726 & n17628 ;
  assign n17630 = ~n17592 & ~n17629 ;
  assign n17631 = ~n17596 & n17630 ;
  assign n17632 = ~n17595 & n17631 ;
  assign n17633 = n1927 & ~n17632 ;
  assign n17634 = ~n17591 & ~n17633 ;
  assign n17635 = \P1_EAX_reg[6]/NET0131  & ~n16968 ;
  assign n17636 = ~n5182 & n16442 ;
  assign n17637 = n2337 & ~n4539 ;
  assign n17638 = n2331 & n17637 ;
  assign n17639 = ~\P1_EAX_reg[6]/NET0131  & ~n15899 ;
  assign n17640 = ~n15900 & ~n17639 ;
  assign n17641 = n2260 & n17640 ;
  assign n17642 = ~n17638 & ~n17641 ;
  assign n17643 = ~n17636 & n17642 ;
  assign n17644 = n2432 & ~n17643 ;
  assign n17645 = ~n17635 & ~n17644 ;
  assign n17646 = \P1_EAX_reg[9]/NET0131  & ~n16968 ;
  assign n17647 = ~n5158 & n16442 ;
  assign n17652 = \P1_InstQueue_reg[11][1]/NET0131  & n1978 ;
  assign n17653 = \P1_InstQueue_reg[7][1]/NET0131  & n1964 ;
  assign n17666 = ~n17652 & ~n17653 ;
  assign n17654 = \P1_InstQueue_reg[15][1]/NET0131  & n1980 ;
  assign n17655 = \P1_InstQueue_reg[5][1]/NET0131  & n1976 ;
  assign n17667 = ~n17654 & ~n17655 ;
  assign n17674 = n17666 & n17667 ;
  assign n17648 = \P1_InstQueue_reg[1][1]/NET0131  & n1982 ;
  assign n17649 = \P1_InstQueue_reg[13][1]/NET0131  & n1949 ;
  assign n17664 = ~n17648 & ~n17649 ;
  assign n17650 = \P1_InstQueue_reg[12][1]/NET0131  & n1946 ;
  assign n17651 = \P1_InstQueue_reg[3][1]/NET0131  & n1966 ;
  assign n17665 = ~n17650 & ~n17651 ;
  assign n17675 = n17664 & n17665 ;
  assign n17676 = n17674 & n17675 ;
  assign n17660 = \P1_InstQueue_reg[6][1]/NET0131  & n1961 ;
  assign n17661 = \P1_InstQueue_reg[14][1]/NET0131  & n1953 ;
  assign n17670 = ~n17660 & ~n17661 ;
  assign n17662 = \P1_InstQueue_reg[10][1]/NET0131  & n1974 ;
  assign n17663 = \P1_InstQueue_reg[8][1]/NET0131  & n1972 ;
  assign n17671 = ~n17662 & ~n17663 ;
  assign n17672 = n17670 & n17671 ;
  assign n17656 = \P1_InstQueue_reg[9][1]/NET0131  & n1968 ;
  assign n17657 = \P1_InstQueue_reg[2][1]/NET0131  & n1958 ;
  assign n17668 = ~n17656 & ~n17657 ;
  assign n17658 = \P1_InstQueue_reg[0][1]/NET0131  & n1955 ;
  assign n17659 = \P1_InstQueue_reg[4][1]/NET0131  & n1970 ;
  assign n17669 = ~n17658 & ~n17659 ;
  assign n17673 = n17668 & n17669 ;
  assign n17677 = n17672 & n17673 ;
  assign n17678 = n17676 & n17677 ;
  assign n17679 = n2337 & ~n17678 ;
  assign n17680 = n2331 & n17679 ;
  assign n17681 = ~\P1_EAX_reg[9]/NET0131  & ~n15902 ;
  assign n17682 = ~n15903 & ~n17681 ;
  assign n17683 = n2260 & n17682 ;
  assign n17684 = ~n17680 & ~n17683 ;
  assign n17685 = ~n17647 & n17684 ;
  assign n17686 = n2432 & ~n17685 ;
  assign n17687 = ~n17646 & ~n17686 ;
  assign n17688 = \P2_EAX_reg[13]/NET0131  & ~n12632 ;
  assign n17691 = \P2_EAX_reg[13]/NET0131  & ~n17594 ;
  assign n17725 = ~\P2_EAX_reg[13]/NET0131  & n12664 ;
  assign n17726 = n12645 & n17725 ;
  assign n17689 = n1811 & ~n16407 ;
  assign n17690 = ~n1804 & n17689 ;
  assign n17696 = \P2_InstQueue_reg[3][5]/NET0131  & n1468 ;
  assign n17697 = \P2_InstQueue_reg[0][5]/NET0131  & n1478 ;
  assign n17710 = ~n17696 & ~n17697 ;
  assign n17698 = \P2_InstQueue_reg[1][5]/NET0131  & n1456 ;
  assign n17699 = \P2_InstQueue_reg[13][5]/NET0131  & n1480 ;
  assign n17711 = ~n17698 & ~n17699 ;
  assign n17718 = n17710 & n17711 ;
  assign n17692 = \P2_InstQueue_reg[5][5]/NET0131  & n1450 ;
  assign n17693 = \P2_InstQueue_reg[10][5]/NET0131  & n1472 ;
  assign n17708 = ~n17692 & ~n17693 ;
  assign n17694 = \P2_InstQueue_reg[15][5]/NET0131  & n1482 ;
  assign n17695 = \P2_InstQueue_reg[4][5]/NET0131  & n1470 ;
  assign n17709 = ~n17694 & ~n17695 ;
  assign n17719 = n17708 & n17709 ;
  assign n17720 = n17718 & n17719 ;
  assign n17704 = \P2_InstQueue_reg[12][5]/NET0131  & n1459 ;
  assign n17705 = \P2_InstQueue_reg[2][5]/NET0131  & n1464 ;
  assign n17714 = ~n17704 & ~n17705 ;
  assign n17706 = \P2_InstQueue_reg[7][5]/NET0131  & n1447 ;
  assign n17707 = \P2_InstQueue_reg[11][5]/NET0131  & n1453 ;
  assign n17715 = ~n17706 & ~n17707 ;
  assign n17716 = n17714 & n17715 ;
  assign n17700 = \P2_InstQueue_reg[6][5]/NET0131  & n1474 ;
  assign n17701 = \P2_InstQueue_reg[8][5]/NET0131  & n1476 ;
  assign n17712 = ~n17700 & ~n17701 ;
  assign n17702 = \P2_InstQueue_reg[9][5]/NET0131  & n1461 ;
  assign n17703 = \P2_InstQueue_reg[14][5]/NET0131  & n1466 ;
  assign n17713 = ~n17702 & ~n17703 ;
  assign n17717 = n17712 & n17713 ;
  assign n17721 = n17716 & n17717 ;
  assign n17722 = n17720 & n17721 ;
  assign n17723 = n1798 & ~n17722 ;
  assign n17724 = n1726 & n17723 ;
  assign n17727 = ~n17690 & ~n17724 ;
  assign n17728 = ~n17726 & n17727 ;
  assign n17729 = ~n17691 & n17728 ;
  assign n17730 = n1927 & ~n17729 ;
  assign n17731 = ~n17688 & ~n17730 ;
  assign n17732 = \P2_EAX_reg[14]/NET0131  & ~n12632 ;
  assign n17734 = ~n12646 & n12664 ;
  assign n17735 = n12669 & ~n17734 ;
  assign n17736 = \P2_EAX_reg[14]/NET0131  & ~n17735 ;
  assign n17770 = ~\P2_EAX_reg[14]/NET0131  & n12664 ;
  assign n17771 = n12646 & n17770 ;
  assign n17733 = ~n1804 & n15010 ;
  assign n17741 = \P2_InstQueue_reg[3][6]/NET0131  & n1468 ;
  assign n17742 = \P2_InstQueue_reg[0][6]/NET0131  & n1478 ;
  assign n17755 = ~n17741 & ~n17742 ;
  assign n17743 = \P2_InstQueue_reg[1][6]/NET0131  & n1456 ;
  assign n17744 = \P2_InstQueue_reg[13][6]/NET0131  & n1480 ;
  assign n17756 = ~n17743 & ~n17744 ;
  assign n17763 = n17755 & n17756 ;
  assign n17737 = \P2_InstQueue_reg[5][6]/NET0131  & n1450 ;
  assign n17738 = \P2_InstQueue_reg[10][6]/NET0131  & n1472 ;
  assign n17753 = ~n17737 & ~n17738 ;
  assign n17739 = \P2_InstQueue_reg[15][6]/NET0131  & n1482 ;
  assign n17740 = \P2_InstQueue_reg[4][6]/NET0131  & n1470 ;
  assign n17754 = ~n17739 & ~n17740 ;
  assign n17764 = n17753 & n17754 ;
  assign n17765 = n17763 & n17764 ;
  assign n17749 = \P2_InstQueue_reg[12][6]/NET0131  & n1459 ;
  assign n17750 = \P2_InstQueue_reg[2][6]/NET0131  & n1464 ;
  assign n17759 = ~n17749 & ~n17750 ;
  assign n17751 = \P2_InstQueue_reg[7][6]/NET0131  & n1447 ;
  assign n17752 = \P2_InstQueue_reg[11][6]/NET0131  & n1453 ;
  assign n17760 = ~n17751 & ~n17752 ;
  assign n17761 = n17759 & n17760 ;
  assign n17745 = \P2_InstQueue_reg[6][6]/NET0131  & n1474 ;
  assign n17746 = \P2_InstQueue_reg[8][6]/NET0131  & n1476 ;
  assign n17757 = ~n17745 & ~n17746 ;
  assign n17747 = \P2_InstQueue_reg[9][6]/NET0131  & n1461 ;
  assign n17748 = \P2_InstQueue_reg[14][6]/NET0131  & n1466 ;
  assign n17758 = ~n17747 & ~n17748 ;
  assign n17762 = n17757 & n17758 ;
  assign n17766 = n17761 & n17762 ;
  assign n17767 = n17765 & n17766 ;
  assign n17768 = n1798 & ~n17767 ;
  assign n17769 = n1726 & n17768 ;
  assign n17772 = ~n17733 & ~n17769 ;
  assign n17773 = ~n17771 & n17772 ;
  assign n17774 = ~n17736 & n17773 ;
  assign n17775 = n1927 & ~n17774 ;
  assign n17776 = ~n17732 & ~n17775 ;
  assign n17777 = \P2_EAX_reg[1]/NET0131  & ~n12632 ;
  assign n17780 = n12669 & ~n17441 ;
  assign n17781 = \P2_EAX_reg[1]/NET0131  & ~n17780 ;
  assign n17778 = n1811 & ~n11541 ;
  assign n17779 = ~n1804 & n17778 ;
  assign n17782 = n1798 & ~n6333 ;
  assign n17783 = n1726 & n17782 ;
  assign n17784 = \P2_EAX_reg[0]/NET0131  & ~\P2_EAX_reg[1]/NET0131  ;
  assign n17785 = n12664 & n17784 ;
  assign n17786 = ~n17783 & ~n17785 ;
  assign n17787 = ~n17779 & n17786 ;
  assign n17788 = ~n17781 & n17787 ;
  assign n17789 = n1927 & ~n17788 ;
  assign n17790 = ~n17777 & ~n17789 ;
  assign n17791 = \P2_EAX_reg[2]/NET0131  & ~n17439 ;
  assign n17792 = ~n8589 & n14771 ;
  assign n17793 = n1798 & ~n6299 ;
  assign n17794 = n1726 & n17793 ;
  assign n17795 = ~\P2_EAX_reg[2]/NET0131  & ~n12634 ;
  assign n17796 = ~n12635 & ~n17795 ;
  assign n17797 = n12664 & n17796 ;
  assign n17798 = ~n17794 & ~n17797 ;
  assign n17799 = ~n17792 & n17798 ;
  assign n17800 = n1927 & ~n17799 ;
  assign n17801 = ~n17791 & ~n17800 ;
  assign n17802 = \P2_EAX_reg[3]/NET0131  & ~n17439 ;
  assign n17803 = ~n5298 & n14771 ;
  assign n17804 = n1798 & ~n6437 ;
  assign n17805 = n1726 & n17804 ;
  assign n17806 = ~\P2_EAX_reg[3]/NET0131  & ~n12635 ;
  assign n17807 = ~n12636 & ~n17806 ;
  assign n17808 = n12664 & n17807 ;
  assign n17809 = ~n17805 & ~n17808 ;
  assign n17810 = ~n17803 & n17809 ;
  assign n17811 = n1927 & ~n17810 ;
  assign n17812 = ~n17802 & ~n17811 ;
  assign n17813 = \P2_EAX_reg[4]/NET0131  & ~n17439 ;
  assign n17814 = ~n3082 & n14771 ;
  assign n17815 = n1798 & ~n6405 ;
  assign n17816 = n1726 & n17815 ;
  assign n17817 = ~\P2_EAX_reg[4]/NET0131  & ~n12636 ;
  assign n17818 = ~n12637 & ~n17817 ;
  assign n17819 = n12664 & n17818 ;
  assign n17820 = ~n17816 & ~n17819 ;
  assign n17821 = ~n17814 & n17820 ;
  assign n17822 = n1927 & ~n17821 ;
  assign n17823 = ~n17813 & ~n17822 ;
  assign n17824 = \P1_EAX_reg[10]/NET0131  & ~n16968 ;
  assign n17831 = \P1_InstQueue_reg[7][2]/NET0131  & n1964 ;
  assign n17832 = \P1_InstQueue_reg[2][2]/NET0131  & n1958 ;
  assign n17845 = ~n17831 & ~n17832 ;
  assign n17833 = \P1_InstQueue_reg[15][2]/NET0131  & n1980 ;
  assign n17834 = \P1_InstQueue_reg[10][2]/NET0131  & n1974 ;
  assign n17846 = ~n17833 & ~n17834 ;
  assign n17853 = n17845 & n17846 ;
  assign n17827 = \P1_InstQueue_reg[1][2]/NET0131  & n1982 ;
  assign n17828 = \P1_InstQueue_reg[13][2]/NET0131  & n1949 ;
  assign n17843 = ~n17827 & ~n17828 ;
  assign n17829 = \P1_InstQueue_reg[14][2]/NET0131  & n1953 ;
  assign n17830 = \P1_InstQueue_reg[3][2]/NET0131  & n1966 ;
  assign n17844 = ~n17829 & ~n17830 ;
  assign n17854 = n17843 & n17844 ;
  assign n17855 = n17853 & n17854 ;
  assign n17839 = \P1_InstQueue_reg[8][2]/NET0131  & n1972 ;
  assign n17840 = \P1_InstQueue_reg[4][2]/NET0131  & n1970 ;
  assign n17849 = ~n17839 & ~n17840 ;
  assign n17841 = \P1_InstQueue_reg[11][2]/NET0131  & n1978 ;
  assign n17842 = \P1_InstQueue_reg[6][2]/NET0131  & n1961 ;
  assign n17850 = ~n17841 & ~n17842 ;
  assign n17851 = n17849 & n17850 ;
  assign n17835 = \P1_InstQueue_reg[5][2]/NET0131  & n1976 ;
  assign n17836 = \P1_InstQueue_reg[12][2]/NET0131  & n1946 ;
  assign n17847 = ~n17835 & ~n17836 ;
  assign n17837 = \P1_InstQueue_reg[0][2]/NET0131  & n1955 ;
  assign n17838 = \P1_InstQueue_reg[9][2]/NET0131  & n1968 ;
  assign n17848 = ~n17837 & ~n17838 ;
  assign n17852 = n17847 & n17848 ;
  assign n17856 = n17851 & n17852 ;
  assign n17857 = n17855 & n17856 ;
  assign n17858 = n2337 & ~n17857 ;
  assign n17859 = n2331 & n17858 ;
  assign n17825 = n2377 & ~n5161 ;
  assign n17826 = ~n2303 & n17825 ;
  assign n17860 = ~\P1_EAX_reg[10]/NET0131  & ~n15903 ;
  assign n17861 = ~n15904 & ~n17860 ;
  assign n17862 = n2260 & n17861 ;
  assign n17863 = ~n17826 & ~n17862 ;
  assign n17864 = ~n17859 & n17863 ;
  assign n17865 = n2432 & ~n17864 ;
  assign n17866 = ~n17824 & ~n17865 ;
  assign n17867 = \P2_EAX_reg[5]/NET0131  & ~n17439 ;
  assign n17868 = ~n10333 & n14771 ;
  assign n17869 = n1798 & ~n6265 ;
  assign n17870 = n1726 & n17869 ;
  assign n17871 = ~\P2_EAX_reg[5]/NET0131  & ~n12637 ;
  assign n17872 = ~n12638 & ~n17871 ;
  assign n17873 = n12664 & n17872 ;
  assign n17874 = ~n17870 & ~n17873 ;
  assign n17875 = ~n17868 & n17874 ;
  assign n17876 = n1927 & ~n17875 ;
  assign n17877 = ~n17867 & ~n17876 ;
  assign n17878 = \P2_EAX_reg[6]/NET0131  & ~n17439 ;
  assign n17879 = ~n7724 & n14771 ;
  assign n17880 = n1798 & ~n6231 ;
  assign n17881 = n1726 & n17880 ;
  assign n17882 = ~\P2_EAX_reg[6]/NET0131  & ~n12638 ;
  assign n17883 = ~n12639 & ~n17882 ;
  assign n17884 = n12664 & n17883 ;
  assign n17885 = ~n17881 & ~n17884 ;
  assign n17886 = ~n17879 & n17885 ;
  assign n17887 = n1927 & ~n17886 ;
  assign n17888 = ~n17878 & ~n17887 ;
  assign n17889 = \P2_EAX_reg[8]/NET0131  & ~n17439 ;
  assign n17890 = n1891 & n16956 ;
  assign n17895 = \P2_InstQueue_reg[3][0]/NET0131  & n1468 ;
  assign n17896 = \P2_InstQueue_reg[0][0]/NET0131  & n1478 ;
  assign n17909 = ~n17895 & ~n17896 ;
  assign n17897 = \P2_InstQueue_reg[1][0]/NET0131  & n1456 ;
  assign n17898 = \P2_InstQueue_reg[13][0]/NET0131  & n1480 ;
  assign n17910 = ~n17897 & ~n17898 ;
  assign n17917 = n17909 & n17910 ;
  assign n17891 = \P2_InstQueue_reg[5][0]/NET0131  & n1450 ;
  assign n17892 = \P2_InstQueue_reg[10][0]/NET0131  & n1472 ;
  assign n17907 = ~n17891 & ~n17892 ;
  assign n17893 = \P2_InstQueue_reg[15][0]/NET0131  & n1482 ;
  assign n17894 = \P2_InstQueue_reg[4][0]/NET0131  & n1470 ;
  assign n17908 = ~n17893 & ~n17894 ;
  assign n17918 = n17907 & n17908 ;
  assign n17919 = n17917 & n17918 ;
  assign n17903 = \P2_InstQueue_reg[12][0]/NET0131  & n1459 ;
  assign n17904 = \P2_InstQueue_reg[2][0]/NET0131  & n1464 ;
  assign n17913 = ~n17903 & ~n17904 ;
  assign n17905 = \P2_InstQueue_reg[7][0]/NET0131  & n1447 ;
  assign n17906 = \P2_InstQueue_reg[11][0]/NET0131  & n1453 ;
  assign n17914 = ~n17905 & ~n17906 ;
  assign n17915 = n17913 & n17914 ;
  assign n17899 = \P2_InstQueue_reg[6][0]/NET0131  & n1474 ;
  assign n17900 = \P2_InstQueue_reg[8][0]/NET0131  & n1476 ;
  assign n17911 = ~n17899 & ~n17900 ;
  assign n17901 = \P2_InstQueue_reg[9][0]/NET0131  & n1461 ;
  assign n17902 = \P2_InstQueue_reg[14][0]/NET0131  & n1466 ;
  assign n17912 = ~n17901 & ~n17902 ;
  assign n17916 = n17911 & n17912 ;
  assign n17920 = n17915 & n17916 ;
  assign n17921 = n17919 & n17920 ;
  assign n17922 = n1798 & ~n17921 ;
  assign n17923 = n1726 & n17922 ;
  assign n17924 = ~\P2_EAX_reg[8]/NET0131  & ~n12640 ;
  assign n17925 = ~n12641 & ~n17924 ;
  assign n17926 = n12664 & n17925 ;
  assign n17927 = ~n17923 & ~n17926 ;
  assign n17928 = ~n17890 & n17927 ;
  assign n17929 = n1927 & ~n17928 ;
  assign n17930 = ~n17889 & ~n17929 ;
  assign n17931 = \P2_EAX_reg[9]/NET0131  & ~n17439 ;
  assign n17932 = ~\buf2_reg[9]/NET0131  & ~n3079 ;
  assign n17933 = ~\buf1_reg[9]/NET0131  & n3079 ;
  assign n17934 = ~n17932 & ~n17933 ;
  assign n17935 = n1811 & n17934 ;
  assign n17936 = ~n1804 & n17935 ;
  assign n17941 = \P2_InstQueue_reg[3][1]/NET0131  & n1468 ;
  assign n17942 = \P2_InstQueue_reg[10][1]/NET0131  & n1472 ;
  assign n17955 = ~n17941 & ~n17942 ;
  assign n17943 = \P2_InstQueue_reg[1][1]/NET0131  & n1456 ;
  assign n17944 = \P2_InstQueue_reg[14][1]/NET0131  & n1466 ;
  assign n17956 = ~n17943 & ~n17944 ;
  assign n17963 = n17955 & n17956 ;
  assign n17937 = \P2_InstQueue_reg[5][1]/NET0131  & n1450 ;
  assign n17938 = \P2_InstQueue_reg[2][1]/NET0131  & n1464 ;
  assign n17953 = ~n17937 & ~n17938 ;
  assign n17939 = \P2_InstQueue_reg[12][1]/NET0131  & n1459 ;
  assign n17940 = \P2_InstQueue_reg[6][1]/NET0131  & n1474 ;
  assign n17954 = ~n17939 & ~n17940 ;
  assign n17964 = n17953 & n17954 ;
  assign n17965 = n17963 & n17964 ;
  assign n17949 = \P2_InstQueue_reg[15][1]/NET0131  & n1482 ;
  assign n17950 = \P2_InstQueue_reg[4][1]/NET0131  & n1470 ;
  assign n17959 = ~n17949 & ~n17950 ;
  assign n17951 = \P2_InstQueue_reg[8][1]/NET0131  & n1476 ;
  assign n17952 = \P2_InstQueue_reg[11][1]/NET0131  & n1453 ;
  assign n17960 = ~n17951 & ~n17952 ;
  assign n17961 = n17959 & n17960 ;
  assign n17945 = \P2_InstQueue_reg[7][1]/NET0131  & n1447 ;
  assign n17946 = \P2_InstQueue_reg[0][1]/NET0131  & n1478 ;
  assign n17957 = ~n17945 & ~n17946 ;
  assign n17947 = \P2_InstQueue_reg[9][1]/NET0131  & n1461 ;
  assign n17948 = \P2_InstQueue_reg[13][1]/NET0131  & n1480 ;
  assign n17958 = ~n17947 & ~n17948 ;
  assign n17962 = n17957 & n17958 ;
  assign n17966 = n17961 & n17962 ;
  assign n17967 = n17965 & n17966 ;
  assign n17968 = n1798 & ~n17967 ;
  assign n17969 = n1726 & n17968 ;
  assign n17970 = ~\P2_EAX_reg[9]/NET0131  & ~n12641 ;
  assign n17971 = ~n12642 & ~n17970 ;
  assign n17972 = n12664 & n17971 ;
  assign n17973 = ~n17969 & ~n17972 ;
  assign n17974 = ~n17936 & n17973 ;
  assign n17975 = n1927 & ~n17974 ;
  assign n17976 = ~n17931 & ~n17975 ;
  assign n17977 = \P1_EAX_reg[11]/NET0131  & ~n15402 ;
  assign n17980 = n2260 & ~n15905 ;
  assign n17981 = n15925 & ~n17980 ;
  assign n17982 = \P1_EAX_reg[11]/NET0131  & ~n17981 ;
  assign n18016 = n15904 & n17980 ;
  assign n17978 = n2377 & ~n5170 ;
  assign n17979 = ~n2303 & n17978 ;
  assign n17987 = \P1_InstQueue_reg[6][3]/NET0131  & n1961 ;
  assign n17988 = \P1_InstQueue_reg[2][3]/NET0131  & n1958 ;
  assign n18001 = ~n17987 & ~n17988 ;
  assign n17989 = \P1_InstQueue_reg[15][3]/NET0131  & n1980 ;
  assign n17990 = \P1_InstQueue_reg[9][3]/NET0131  & n1968 ;
  assign n18002 = ~n17989 & ~n17990 ;
  assign n18009 = n18001 & n18002 ;
  assign n17983 = \P1_InstQueue_reg[1][3]/NET0131  & n1982 ;
  assign n17984 = \P1_InstQueue_reg[3][3]/NET0131  & n1966 ;
  assign n17999 = ~n17983 & ~n17984 ;
  assign n17985 = \P1_InstQueue_reg[4][3]/NET0131  & n1970 ;
  assign n17986 = \P1_InstQueue_reg[13][3]/NET0131  & n1949 ;
  assign n18000 = ~n17985 & ~n17986 ;
  assign n18010 = n17999 & n18000 ;
  assign n18011 = n18009 & n18010 ;
  assign n17995 = \P1_InstQueue_reg[8][3]/NET0131  & n1972 ;
  assign n17996 = \P1_InstQueue_reg[7][3]/NET0131  & n1964 ;
  assign n18005 = ~n17995 & ~n17996 ;
  assign n17997 = \P1_InstQueue_reg[11][3]/NET0131  & n1978 ;
  assign n17998 = \P1_InstQueue_reg[10][3]/NET0131  & n1974 ;
  assign n18006 = ~n17997 & ~n17998 ;
  assign n18007 = n18005 & n18006 ;
  assign n17991 = \P1_InstQueue_reg[14][3]/NET0131  & n1953 ;
  assign n17992 = \P1_InstQueue_reg[5][3]/NET0131  & n1976 ;
  assign n18003 = ~n17991 & ~n17992 ;
  assign n17993 = \P1_InstQueue_reg[0][3]/NET0131  & n1955 ;
  assign n17994 = \P1_InstQueue_reg[12][3]/NET0131  & n1946 ;
  assign n18004 = ~n17993 & ~n17994 ;
  assign n18008 = n18003 & n18004 ;
  assign n18012 = n18007 & n18008 ;
  assign n18013 = n18011 & n18012 ;
  assign n18014 = n2337 & ~n18013 ;
  assign n18015 = n2331 & n18014 ;
  assign n18017 = ~n17979 & ~n18015 ;
  assign n18018 = ~n18016 & n18017 ;
  assign n18019 = ~n17982 & n18018 ;
  assign n18020 = n2432 & ~n18019 ;
  assign n18021 = ~n17977 & ~n18020 ;
  assign n18024 = n15389 & n15390 ;
  assign n18026 = \P1_EBX_reg[29]/NET0131  & n18024 ;
  assign n18025 = ~\P1_EBX_reg[29]/NET0131  & ~n18024 ;
  assign n18027 = n2262 & ~n18025 ;
  assign n18028 = ~n18026 & n18027 ;
  assign n18022 = \P1_EBX_reg[29]/NET0131  & ~n15073 ;
  assign n18023 = n2242 & n16315 ;
  assign n18029 = ~n18022 & ~n18023 ;
  assign n18030 = ~n18028 & n18029 ;
  assign n18031 = n2432 & ~n18030 ;
  assign n18032 = \P1_EBX_reg[29]/NET0131  & ~n15402 ;
  assign n18033 = ~n18031 & ~n18032 ;
  assign n18036 = ~\P2_EBX_reg[29]/NET0131  & ~n15060 ;
  assign n18037 = n1766 & ~n15061 ;
  assign n18038 = ~n18036 & n18037 ;
  assign n18034 = n1722 & n16403 ;
  assign n18035 = \P2_EBX_reg[29]/NET0131  & ~n15019 ;
  assign n18039 = ~n18034 & ~n18035 ;
  assign n18040 = ~n18038 & n18039 ;
  assign n18041 = n1927 & ~n18040 ;
  assign n18042 = \P2_EBX_reg[29]/NET0131  & ~n12632 ;
  assign n18043 = ~n18041 & ~n18042 ;
  assign n18044 = \P1_EAX_reg[14]/NET0131  & ~n15402 ;
  assign n18046 = n2260 & ~n15907 ;
  assign n18047 = n15925 & ~n18046 ;
  assign n18048 = \P1_EAX_reg[14]/NET0131  & ~n18047 ;
  assign n18082 = ~n5191 & n16442 ;
  assign n18045 = ~\P1_EAX_reg[14]/NET0131  & n16480 ;
  assign n18053 = \P1_InstQueue_reg[2][6]/NET0131  & n1958 ;
  assign n18054 = \P1_InstQueue_reg[7][6]/NET0131  & n1964 ;
  assign n18067 = ~n18053 & ~n18054 ;
  assign n18055 = \P1_InstQueue_reg[15][6]/NET0131  & n1980 ;
  assign n18056 = \P1_InstQueue_reg[8][6]/NET0131  & n1972 ;
  assign n18068 = ~n18055 & ~n18056 ;
  assign n18075 = n18067 & n18068 ;
  assign n18049 = \P1_InstQueue_reg[1][6]/NET0131  & n1982 ;
  assign n18050 = \P1_InstQueue_reg[3][6]/NET0131  & n1966 ;
  assign n18065 = ~n18049 & ~n18050 ;
  assign n18051 = \P1_InstQueue_reg[12][6]/NET0131  & n1946 ;
  assign n18052 = \P1_InstQueue_reg[13][6]/NET0131  & n1949 ;
  assign n18066 = ~n18051 & ~n18052 ;
  assign n18076 = n18065 & n18066 ;
  assign n18077 = n18075 & n18076 ;
  assign n18061 = \P1_InstQueue_reg[6][6]/NET0131  & n1961 ;
  assign n18062 = \P1_InstQueue_reg[14][6]/NET0131  & n1953 ;
  assign n18071 = ~n18061 & ~n18062 ;
  assign n18063 = \P1_InstQueue_reg[10][6]/NET0131  & n1974 ;
  assign n18064 = \P1_InstQueue_reg[11][6]/NET0131  & n1978 ;
  assign n18072 = ~n18063 & ~n18064 ;
  assign n18073 = n18071 & n18072 ;
  assign n18057 = \P1_InstQueue_reg[9][6]/NET0131  & n1968 ;
  assign n18058 = \P1_InstQueue_reg[5][6]/NET0131  & n1976 ;
  assign n18069 = ~n18057 & ~n18058 ;
  assign n18059 = \P1_InstQueue_reg[0][6]/NET0131  & n1955 ;
  assign n18060 = \P1_InstQueue_reg[4][6]/NET0131  & n1970 ;
  assign n18070 = ~n18059 & ~n18060 ;
  assign n18074 = n18069 & n18070 ;
  assign n18078 = n18073 & n18074 ;
  assign n18079 = n18077 & n18078 ;
  assign n18080 = n2337 & ~n18079 ;
  assign n18081 = n2331 & n18080 ;
  assign n18083 = ~n18045 & ~n18081 ;
  assign n18084 = ~n18082 & n18083 ;
  assign n18085 = ~n18048 & n18084 ;
  assign n18086 = n2432 & ~n18085 ;
  assign n18087 = ~n18044 & ~n18086 ;
  assign n18088 = \P1_EAX_reg[13]/NET0131  & ~n15402 ;
  assign n18090 = \P1_EAX_reg[13]/NET0131  & ~n18047 ;
  assign n18124 = n15906 & n18046 ;
  assign n18089 = ~n5200 & n16442 ;
  assign n18095 = \P1_InstQueue_reg[10][5]/NET0131  & n1974 ;
  assign n18096 = \P1_InstQueue_reg[2][5]/NET0131  & n1958 ;
  assign n18109 = ~n18095 & ~n18096 ;
  assign n18097 = \P1_InstQueue_reg[15][5]/NET0131  & n1980 ;
  assign n18098 = \P1_InstQueue_reg[7][5]/NET0131  & n1964 ;
  assign n18110 = ~n18097 & ~n18098 ;
  assign n18117 = n18109 & n18110 ;
  assign n18091 = \P1_InstQueue_reg[1][5]/NET0131  & n1982 ;
  assign n18092 = \P1_InstQueue_reg[13][5]/NET0131  & n1949 ;
  assign n18107 = ~n18091 & ~n18092 ;
  assign n18093 = \P1_InstQueue_reg[8][5]/NET0131  & n1972 ;
  assign n18094 = \P1_InstQueue_reg[3][5]/NET0131  & n1966 ;
  assign n18108 = ~n18093 & ~n18094 ;
  assign n18118 = n18107 & n18108 ;
  assign n18119 = n18117 & n18118 ;
  assign n18103 = \P1_InstQueue_reg[14][5]/NET0131  & n1953 ;
  assign n18104 = \P1_InstQueue_reg[4][5]/NET0131  & n1970 ;
  assign n18113 = ~n18103 & ~n18104 ;
  assign n18105 = \P1_InstQueue_reg[12][5]/NET0131  & n1946 ;
  assign n18106 = \P1_InstQueue_reg[9][5]/NET0131  & n1968 ;
  assign n18114 = ~n18105 & ~n18106 ;
  assign n18115 = n18113 & n18114 ;
  assign n18099 = \P1_InstQueue_reg[5][5]/NET0131  & n1976 ;
  assign n18100 = \P1_InstQueue_reg[11][5]/NET0131  & n1978 ;
  assign n18111 = ~n18099 & ~n18100 ;
  assign n18101 = \P1_InstQueue_reg[0][5]/NET0131  & n1955 ;
  assign n18102 = \P1_InstQueue_reg[6][5]/NET0131  & n1961 ;
  assign n18112 = ~n18101 & ~n18102 ;
  assign n18116 = n18111 & n18112 ;
  assign n18120 = n18115 & n18116 ;
  assign n18121 = n18119 & n18120 ;
  assign n18122 = n2337 & ~n18121 ;
  assign n18123 = n2331 & n18122 ;
  assign n18125 = ~n18089 & ~n18123 ;
  assign n18126 = ~n18124 & n18125 ;
  assign n18127 = ~n18090 & n18126 ;
  assign n18128 = n2432 & ~n18127 ;
  assign n18129 = ~n18088 & ~n18128 ;
  assign n18130 = \P1_EAX_reg[12]/NET0131  & ~n15402 ;
  assign n18131 = n15924 & ~n17980 ;
  assign n18132 = \P1_EAX_reg[12]/NET0131  & ~n18131 ;
  assign n18168 = \P1_EAX_reg[12]/NET0131  & ~n2377 ;
  assign n18169 = n2377 & ~n5197 ;
  assign n18170 = ~n18168 & ~n18169 ;
  assign n18171 = ~n2303 & ~n18170 ;
  assign n18133 = ~\P1_EAX_reg[12]/NET0131  & n2260 ;
  assign n18134 = n15905 & n18133 ;
  assign n18139 = \P1_InstQueue_reg[0][4]/NET0131  & n1955 ;
  assign n18140 = \P1_InstQueue_reg[12][4]/NET0131  & n1946 ;
  assign n18153 = ~n18139 & ~n18140 ;
  assign n18141 = \P1_InstQueue_reg[3][4]/NET0131  & n1966 ;
  assign n18142 = \P1_InstQueue_reg[9][4]/NET0131  & n1968 ;
  assign n18154 = ~n18141 & ~n18142 ;
  assign n18161 = n18153 & n18154 ;
  assign n18135 = \P1_InstQueue_reg[15][4]/NET0131  & n1980 ;
  assign n18136 = \P1_InstQueue_reg[13][4]/NET0131  & n1949 ;
  assign n18151 = ~n18135 & ~n18136 ;
  assign n18137 = \P1_InstQueue_reg[7][4]/NET0131  & n1964 ;
  assign n18138 = \P1_InstQueue_reg[8][4]/NET0131  & n1972 ;
  assign n18152 = ~n18137 & ~n18138 ;
  assign n18162 = n18151 & n18152 ;
  assign n18163 = n18161 & n18162 ;
  assign n18147 = \P1_InstQueue_reg[14][4]/NET0131  & n1953 ;
  assign n18148 = \P1_InstQueue_reg[6][4]/NET0131  & n1961 ;
  assign n18157 = ~n18147 & ~n18148 ;
  assign n18149 = \P1_InstQueue_reg[2][4]/NET0131  & n1958 ;
  assign n18150 = \P1_InstQueue_reg[10][4]/NET0131  & n1974 ;
  assign n18158 = ~n18149 & ~n18150 ;
  assign n18159 = n18157 & n18158 ;
  assign n18143 = \P1_InstQueue_reg[5][4]/NET0131  & n1976 ;
  assign n18144 = \P1_InstQueue_reg[4][4]/NET0131  & n1970 ;
  assign n18155 = ~n18143 & ~n18144 ;
  assign n18145 = \P1_InstQueue_reg[1][4]/NET0131  & n1982 ;
  assign n18146 = \P1_InstQueue_reg[11][4]/NET0131  & n1978 ;
  assign n18156 = ~n18145 & ~n18146 ;
  assign n18160 = n18155 & n18156 ;
  assign n18164 = n18159 & n18160 ;
  assign n18165 = n18163 & n18164 ;
  assign n18166 = n2337 & ~n18165 ;
  assign n18167 = n2331 & n18166 ;
  assign n18172 = ~n18134 & ~n18167 ;
  assign n18173 = ~n18171 & n18172 ;
  assign n18174 = ~n18132 & n18173 ;
  assign n18175 = n2432 & ~n18174 ;
  assign n18176 = ~n18130 & ~n18175 ;
  assign n18177 = \P3_uWord_reg[8]/NET0131  & ~n16090 ;
  assign n18178 = n2453 & ~n2815 ;
  assign n18179 = \buf2_reg[8]/NET0131  & ~n2835 ;
  assign n18180 = n2821 & n18179 ;
  assign n18181 = ~n16893 & ~n18180 ;
  assign n18182 = n18178 & ~n18181 ;
  assign n18183 = ~n18177 & ~n18182 ;
  assign n18184 = \P1_EAX_reg[1]/NET0131  & ~n15402 ;
  assign n18186 = ~\P1_EAX_reg[0]/NET0131  & n2260 ;
  assign n18187 = n15925 & ~n18186 ;
  assign n18188 = \P1_EAX_reg[1]/NET0131  & ~n18187 ;
  assign n18185 = ~n5185 & n16442 ;
  assign n18189 = n2337 & ~n4710 ;
  assign n18190 = n2331 & n18189 ;
  assign n18191 = \P1_EAX_reg[0]/NET0131  & ~\P1_EAX_reg[1]/NET0131  ;
  assign n18192 = n2260 & n18191 ;
  assign n18193 = ~n18190 & ~n18192 ;
  assign n18194 = ~n18185 & n18193 ;
  assign n18195 = ~n18188 & n18194 ;
  assign n18196 = n2432 & ~n18195 ;
  assign n18197 = ~n18184 & ~n18196 ;
  assign n18207 = ~\P3_InstQueueWr_Addr_reg[0]/NET0131  & ~\P3_InstQueueWr_Addr_reg[1]/NET0131  ;
  assign n18208 = ~\P3_InstQueueWr_Addr_reg[2]/NET0131  & ~\P3_InstQueueWr_Addr_reg[3]/NET0131  ;
  assign n18209 = n18207 & n18208 ;
  assign n18221 = n2571 & n18209 ;
  assign n18220 = ~\P3_InstQueue_reg[0][4]/NET0131  & ~n18209 ;
  assign n18222 = n2994 & ~n18220 ;
  assign n18223 = ~n18221 & n18222 ;
  assign n18198 = \P3_InstQueueWr_Addr_reg[0]/NET0131  & ~\P3_InstQueueWr_Addr_reg[1]/NET0131  ;
  assign n18199 = \P3_InstQueueWr_Addr_reg[2]/NET0131  & n18198 ;
  assign n18200 = \P3_InstQueueWr_Addr_reg[3]/NET0131  & n18199 ;
  assign n18201 = ~\P3_InstQueueWr_Addr_reg[0]/NET0131  & \P3_InstQueueWr_Addr_reg[1]/NET0131  ;
  assign n18202 = \P3_InstQueueWr_Addr_reg[2]/NET0131  & n18201 ;
  assign n18203 = \P3_InstQueueWr_Addr_reg[3]/NET0131  & n18202 ;
  assign n18204 = ~n18200 & ~n18203 ;
  assign n18205 = n2959 & n18204 ;
  assign n18206 = ~n10076 & ~n18205 ;
  assign n18210 = \P3_InstQueueWr_Addr_reg[0]/NET0131  & \P3_InstQueueWr_Addr_reg[1]/NET0131  ;
  assign n18211 = \P3_InstQueueWr_Addr_reg[2]/NET0131  & n18210 ;
  assign n18212 = \P3_InstQueueWr_Addr_reg[3]/NET0131  & n18211 ;
  assign n18213 = ~n18209 & ~n18212 ;
  assign n18214 = ~n18206 & n18213 ;
  assign n18215 = ~n2453 & ~n2996 ;
  assign n18216 = ~n2968 & n18215 ;
  assign n18217 = n14119 & n18216 ;
  assign n18218 = ~n18214 & n18217 ;
  assign n18219 = \P3_InstQueue_reg[0][4]/NET0131  & ~n18218 ;
  assign n18224 = \buf2_reg[28]/NET0131  & n18200 ;
  assign n18225 = \buf2_reg[20]/NET0131  & n18203 ;
  assign n18226 = ~n18224 & ~n18225 ;
  assign n18227 = n2970 & ~n18226 ;
  assign n18228 = ~n18206 & ~n18213 ;
  assign n18229 = \buf2_reg[4]/NET0131  & n18228 ;
  assign n18230 = ~n18227 & ~n18229 ;
  assign n18231 = ~n18219 & n18230 ;
  assign n18232 = ~n18223 & n18231 ;
  assign n18234 = ~\P3_InstQueueWr_Addr_reg[2]/NET0131  & \P3_InstQueueWr_Addr_reg[3]/NET0131  ;
  assign n18245 = \P3_InstQueueWr_Addr_reg[1]/NET0131  & n18234 ;
  assign n18246 = ~\P3_InstQueueWr_Addr_reg[0]/NET0131  & n18245 ;
  assign n18248 = n2571 & n18246 ;
  assign n18247 = ~\P3_InstQueue_reg[10][4]/NET0131  & ~n18246 ;
  assign n18249 = n2994 & ~n18247 ;
  assign n18250 = ~n18248 & n18249 ;
  assign n18233 = ~\P3_InstQueueWr_Addr_reg[3]/NET0131  & n18211 ;
  assign n18235 = ~\P3_InstQueueWr_Addr_reg[1]/NET0131  & n18234 ;
  assign n18236 = ~\P3_InstQueueWr_Addr_reg[0]/NET0131  & n18235 ;
  assign n18237 = ~n18233 & ~n18236 ;
  assign n18238 = n2959 & n18237 ;
  assign n18239 = ~n10076 & ~n18238 ;
  assign n18240 = ~n18198 & ~n18201 ;
  assign n18241 = n18234 & ~n18240 ;
  assign n18242 = ~n18239 & ~n18241 ;
  assign n18243 = n18217 & ~n18242 ;
  assign n18244 = \P3_InstQueue_reg[10][4]/NET0131  & ~n18243 ;
  assign n18251 = \buf2_reg[28]/NET0131  & n18233 ;
  assign n18252 = \buf2_reg[20]/NET0131  & n18236 ;
  assign n18253 = ~n18251 & ~n18252 ;
  assign n18254 = n2970 & ~n18253 ;
  assign n18255 = ~n18239 & n18241 ;
  assign n18256 = \buf2_reg[4]/NET0131  & n18255 ;
  assign n18257 = ~n18254 & ~n18256 ;
  assign n18258 = ~n18244 & n18257 ;
  assign n18259 = ~n18250 & n18258 ;
  assign n18266 = \P3_InstQueueWr_Addr_reg[0]/NET0131  & n18245 ;
  assign n18268 = n2571 & n18266 ;
  assign n18267 = ~\P3_InstQueue_reg[11][4]/NET0131  & ~n18266 ;
  assign n18269 = n2994 & ~n18267 ;
  assign n18270 = ~n18268 & n18269 ;
  assign n18260 = \P3_DataWidth_reg[1]/NET0131  & n18235 ;
  assign n18261 = ~n4415 & n18260 ;
  assign n18262 = ~n10074 & ~n18261 ;
  assign n18263 = ~n18245 & n18262 ;
  assign n18264 = n18217 & ~n18263 ;
  assign n18265 = \P3_InstQueue_reg[11][4]/NET0131  & ~n18264 ;
  assign n18271 = \P3_InstQueueWr_Addr_reg[0]/NET0131  & n18235 ;
  assign n18272 = \buf2_reg[20]/NET0131  & n18271 ;
  assign n18273 = \buf2_reg[28]/NET0131  & n18236 ;
  assign n18274 = ~n18272 & ~n18273 ;
  assign n18275 = n2970 & ~n18274 ;
  assign n18276 = \buf2_reg[4]/NET0131  & n18245 ;
  assign n18277 = n18262 & n18276 ;
  assign n18278 = ~n18275 & ~n18277 ;
  assign n18279 = ~n18265 & n18278 ;
  assign n18280 = ~n18270 & n18279 ;
  assign n18283 = \P3_InstQueueWr_Addr_reg[2]/NET0131  & n18207 ;
  assign n18284 = \P3_InstQueueWr_Addr_reg[3]/NET0131  & n18283 ;
  assign n18290 = n2571 & n18284 ;
  assign n18289 = ~\P3_InstQueue_reg[12][4]/NET0131  & ~n18284 ;
  assign n18291 = n2994 & ~n18289 ;
  assign n18292 = ~n18290 & n18291 ;
  assign n18281 = n2959 & ~n18241 ;
  assign n18282 = ~n10076 & ~n18281 ;
  assign n18285 = ~n18266 & ~n18284 ;
  assign n18286 = ~n18282 & n18285 ;
  assign n18287 = n18217 & ~n18286 ;
  assign n18288 = \P3_InstQueue_reg[12][4]/NET0131  & ~n18287 ;
  assign n18293 = \buf2_reg[20]/NET0131  & n18246 ;
  assign n18294 = \buf2_reg[28]/NET0131  & n18271 ;
  assign n18295 = ~n18293 & ~n18294 ;
  assign n18296 = n2970 & ~n18295 ;
  assign n18297 = ~n18282 & ~n18285 ;
  assign n18298 = \buf2_reg[4]/NET0131  & n18297 ;
  assign n18299 = ~n18296 & ~n18298 ;
  assign n18300 = ~n18288 & n18299 ;
  assign n18301 = ~n18292 & n18300 ;
  assign n18316 = n2571 & n18200 ;
  assign n18315 = ~\P3_InstQueue_reg[13][4]/NET0131  & ~n18200 ;
  assign n18317 = n2994 & ~n18315 ;
  assign n18318 = ~n18316 & n18317 ;
  assign n18302 = ~n18200 & ~n18284 ;
  assign n18303 = \P3_DataWidth_reg[1]/NET0131  & n18245 ;
  assign n18304 = ~n4415 & n18303 ;
  assign n18305 = ~n10074 & ~n18304 ;
  assign n18306 = n18302 & n18305 ;
  assign n18307 = n18217 & ~n18306 ;
  assign n18308 = \P3_InstQueue_reg[13][4]/NET0131  & ~n18307 ;
  assign n18309 = \buf2_reg[20]/NET0131  & n18266 ;
  assign n18310 = \buf2_reg[28]/NET0131  & n18246 ;
  assign n18311 = ~n18309 & ~n18310 ;
  assign n18312 = n2970 & ~n18311 ;
  assign n18313 = \buf2_reg[4]/NET0131  & ~n18302 ;
  assign n18314 = n18305 & n18313 ;
  assign n18319 = ~n18312 & ~n18314 ;
  assign n18320 = ~n18308 & n18319 ;
  assign n18321 = ~n18318 & n18320 ;
  assign n18328 = n2571 & n18203 ;
  assign n18327 = ~\P3_InstQueue_reg[14][4]/NET0131  & ~n18203 ;
  assign n18329 = n2994 & ~n18327 ;
  assign n18330 = ~n18328 & n18329 ;
  assign n18322 = n2959 & n18285 ;
  assign n18323 = ~n10076 & ~n18322 ;
  assign n18324 = n18204 & ~n18323 ;
  assign n18325 = n18217 & ~n18324 ;
  assign n18326 = \P3_InstQueue_reg[14][4]/NET0131  & ~n18325 ;
  assign n18331 = \buf2_reg[28]/NET0131  & n18266 ;
  assign n18332 = \buf2_reg[20]/NET0131  & n18284 ;
  assign n18333 = ~n18331 & ~n18332 ;
  assign n18334 = n2970 & ~n18333 ;
  assign n18335 = ~n18204 & ~n18323 ;
  assign n18336 = \buf2_reg[4]/NET0131  & n18335 ;
  assign n18337 = ~n18334 & ~n18336 ;
  assign n18338 = ~n18326 & n18337 ;
  assign n18339 = ~n18330 & n18338 ;
  assign n18347 = n2571 & n18212 ;
  assign n18346 = ~\P3_InstQueue_reg[15][4]/NET0131  & ~n18212 ;
  assign n18348 = n2994 & ~n18346 ;
  assign n18349 = ~n18347 & n18348 ;
  assign n18340 = n2959 & n18302 ;
  assign n18341 = ~n10076 & ~n18340 ;
  assign n18342 = ~n18203 & ~n18212 ;
  assign n18343 = ~n18341 & n18342 ;
  assign n18344 = n18217 & ~n18343 ;
  assign n18345 = \P3_InstQueue_reg[15][4]/NET0131  & ~n18344 ;
  assign n18350 = \buf2_reg[28]/NET0131  & n18284 ;
  assign n18351 = \buf2_reg[20]/NET0131  & n18200 ;
  assign n18352 = ~n18350 & ~n18351 ;
  assign n18353 = n2970 & ~n18352 ;
  assign n18354 = ~n18341 & ~n18342 ;
  assign n18355 = \buf2_reg[4]/NET0131  & n18354 ;
  assign n18356 = ~n18353 & ~n18355 ;
  assign n18357 = ~n18345 & n18356 ;
  assign n18358 = ~n18349 & n18357 ;
  assign n18361 = n18198 & n18208 ;
  assign n18367 = n2571 & n18361 ;
  assign n18366 = ~\P3_InstQueue_reg[1][4]/NET0131  & ~n18361 ;
  assign n18368 = n2994 & ~n18366 ;
  assign n18369 = ~n18367 & n18368 ;
  assign n18359 = n2959 & n18342 ;
  assign n18360 = ~n10076 & ~n18359 ;
  assign n18362 = ~n18209 & ~n18361 ;
  assign n18363 = ~n18360 & n18362 ;
  assign n18364 = n18217 & ~n18363 ;
  assign n18365 = \P3_InstQueue_reg[1][4]/NET0131  & ~n18364 ;
  assign n18370 = \buf2_reg[28]/NET0131  & n18203 ;
  assign n18371 = \buf2_reg[20]/NET0131  & n18212 ;
  assign n18372 = ~n18370 & ~n18371 ;
  assign n18373 = n2970 & ~n18372 ;
  assign n18374 = ~n18360 & ~n18362 ;
  assign n18375 = \buf2_reg[4]/NET0131  & n18374 ;
  assign n18376 = ~n18373 & ~n18375 ;
  assign n18377 = ~n18365 & n18376 ;
  assign n18378 = ~n18369 & n18377 ;
  assign n18385 = \P3_InstQueueWr_Addr_reg[1]/NET0131  & n18208 ;
  assign n18386 = ~\P3_InstQueueWr_Addr_reg[0]/NET0131  & n18385 ;
  assign n18388 = n2571 & n18386 ;
  assign n18387 = ~\P3_InstQueue_reg[2][4]/NET0131  & ~n18386 ;
  assign n18389 = n2994 & ~n18387 ;
  assign n18390 = ~n18388 & n18389 ;
  assign n18379 = n2959 & n18213 ;
  assign n18380 = ~n10076 & ~n18379 ;
  assign n18381 = n18208 & ~n18240 ;
  assign n18382 = ~n18380 & ~n18381 ;
  assign n18383 = n18217 & ~n18382 ;
  assign n18384 = \P3_InstQueue_reg[2][4]/NET0131  & ~n18383 ;
  assign n18391 = \buf2_reg[28]/NET0131  & n18212 ;
  assign n18392 = \buf2_reg[20]/NET0131  & n18209 ;
  assign n18393 = ~n18391 & ~n18392 ;
  assign n18394 = n2970 & ~n18393 ;
  assign n18395 = ~n18380 & n18381 ;
  assign n18396 = \buf2_reg[4]/NET0131  & n18395 ;
  assign n18397 = ~n18394 & ~n18396 ;
  assign n18398 = ~n18384 & n18397 ;
  assign n18399 = ~n18390 & n18398 ;
  assign n18405 = \P3_InstQueueWr_Addr_reg[0]/NET0131  & n18385 ;
  assign n18407 = n2571 & n18405 ;
  assign n18406 = ~\P3_InstQueue_reg[3][4]/NET0131  & ~n18405 ;
  assign n18408 = n2994 & ~n18406 ;
  assign n18409 = ~n18407 & n18408 ;
  assign n18400 = n2959 & n18362 ;
  assign n18401 = ~n10076 & ~n18400 ;
  assign n18402 = ~n18385 & ~n18401 ;
  assign n18403 = n18217 & ~n18402 ;
  assign n18404 = \P3_InstQueue_reg[3][4]/NET0131  & ~n18403 ;
  assign n18410 = \buf2_reg[20]/NET0131  & n18361 ;
  assign n18411 = \buf2_reg[28]/NET0131  & n18209 ;
  assign n18412 = ~n18410 & ~n18411 ;
  assign n18413 = n2970 & ~n18412 ;
  assign n18414 = n18385 & ~n18401 ;
  assign n18415 = \buf2_reg[4]/NET0131  & n18414 ;
  assign n18416 = ~n18413 & ~n18415 ;
  assign n18417 = ~n18404 & n18416 ;
  assign n18418 = ~n18409 & n18417 ;
  assign n18421 = ~\P3_InstQueueWr_Addr_reg[3]/NET0131  & n18283 ;
  assign n18427 = n2571 & n18421 ;
  assign n18426 = ~\P3_InstQueue_reg[4][4]/NET0131  & ~n18421 ;
  assign n18428 = n2994 & ~n18426 ;
  assign n18429 = ~n18427 & n18428 ;
  assign n18419 = n2959 & ~n18381 ;
  assign n18420 = ~n10076 & ~n18419 ;
  assign n18422 = ~n18405 & ~n18421 ;
  assign n18423 = ~n18420 & n18422 ;
  assign n18424 = n18217 & ~n18423 ;
  assign n18425 = \P3_InstQueue_reg[4][4]/NET0131  & ~n18424 ;
  assign n18430 = \buf2_reg[20]/NET0131  & n18386 ;
  assign n18431 = \buf2_reg[28]/NET0131  & n18361 ;
  assign n18432 = ~n18430 & ~n18431 ;
  assign n18433 = n2970 & ~n18432 ;
  assign n18434 = ~n18420 & ~n18422 ;
  assign n18435 = \buf2_reg[4]/NET0131  & n18434 ;
  assign n18436 = ~n18433 & ~n18435 ;
  assign n18437 = ~n18425 & n18436 ;
  assign n18438 = ~n18429 & n18437 ;
  assign n18439 = ~\P3_InstQueueWr_Addr_reg[3]/NET0131  & n18199 ;
  assign n18454 = n2571 & n18439 ;
  assign n18453 = ~\P3_InstQueue_reg[5][4]/NET0131  & ~n18439 ;
  assign n18455 = n2994 & ~n18453 ;
  assign n18456 = ~n18454 & n18455 ;
  assign n18440 = ~n18421 & ~n18439 ;
  assign n18441 = \P3_DataWidth_reg[1]/NET0131  & n18385 ;
  assign n18442 = ~n4415 & n18441 ;
  assign n18443 = ~n10074 & ~n18442 ;
  assign n18444 = n18440 & n18443 ;
  assign n18445 = n18217 & ~n18444 ;
  assign n18446 = \P3_InstQueue_reg[5][4]/NET0131  & ~n18445 ;
  assign n18447 = \buf2_reg[20]/NET0131  & n18405 ;
  assign n18448 = \buf2_reg[28]/NET0131  & n18386 ;
  assign n18449 = ~n18447 & ~n18448 ;
  assign n18450 = n2970 & ~n18449 ;
  assign n18451 = \buf2_reg[4]/NET0131  & ~n18440 ;
  assign n18452 = n18443 & n18451 ;
  assign n18457 = ~n18450 & ~n18452 ;
  assign n18458 = ~n18446 & n18457 ;
  assign n18459 = ~n18456 & n18458 ;
  assign n18462 = ~\P3_InstQueueWr_Addr_reg[3]/NET0131  & n18202 ;
  assign n18468 = n2571 & n18462 ;
  assign n18467 = ~\P3_InstQueue_reg[6][4]/NET0131  & ~n18462 ;
  assign n18469 = n2994 & ~n18467 ;
  assign n18470 = ~n18468 & n18469 ;
  assign n18460 = n2959 & n18422 ;
  assign n18461 = ~n10076 & ~n18460 ;
  assign n18463 = ~n18439 & ~n18462 ;
  assign n18464 = ~n18461 & n18463 ;
  assign n18465 = n18217 & ~n18464 ;
  assign n18466 = \P3_InstQueue_reg[6][4]/NET0131  & ~n18465 ;
  assign n18471 = \buf2_reg[28]/NET0131  & n18405 ;
  assign n18472 = \buf2_reg[20]/NET0131  & n18421 ;
  assign n18473 = ~n18471 & ~n18472 ;
  assign n18474 = n2970 & ~n18473 ;
  assign n18475 = ~n18461 & ~n18463 ;
  assign n18476 = \buf2_reg[4]/NET0131  & n18475 ;
  assign n18477 = ~n18474 & ~n18476 ;
  assign n18478 = ~n18466 & n18477 ;
  assign n18479 = ~n18470 & n18478 ;
  assign n18487 = n2571 & n18233 ;
  assign n18486 = ~\P3_InstQueue_reg[7][4]/NET0131  & ~n18233 ;
  assign n18488 = n2994 & ~n18486 ;
  assign n18489 = ~n18487 & n18488 ;
  assign n18480 = n2959 & n18440 ;
  assign n18481 = ~n10076 & ~n18480 ;
  assign n18482 = ~n18233 & ~n18462 ;
  assign n18483 = ~n18481 & n18482 ;
  assign n18484 = n18217 & ~n18483 ;
  assign n18485 = \P3_InstQueue_reg[7][4]/NET0131  & ~n18484 ;
  assign n18490 = \buf2_reg[28]/NET0131  & n18421 ;
  assign n18491 = \buf2_reg[20]/NET0131  & n18439 ;
  assign n18492 = ~n18490 & ~n18491 ;
  assign n18493 = n2970 & ~n18492 ;
  assign n18494 = ~n18481 & ~n18482 ;
  assign n18495 = \buf2_reg[4]/NET0131  & n18494 ;
  assign n18496 = ~n18493 & ~n18495 ;
  assign n18497 = ~n18485 & n18496 ;
  assign n18498 = ~n18489 & n18497 ;
  assign n18505 = n2571 & n18236 ;
  assign n18504 = ~\P3_InstQueue_reg[8][4]/NET0131  & ~n18236 ;
  assign n18506 = n2994 & ~n18504 ;
  assign n18507 = ~n18505 & n18506 ;
  assign n18499 = n2959 & n18463 ;
  assign n18500 = ~n10076 & ~n18499 ;
  assign n18501 = n18237 & ~n18500 ;
  assign n18502 = n18217 & ~n18501 ;
  assign n18503 = \P3_InstQueue_reg[8][4]/NET0131  & ~n18502 ;
  assign n18508 = \buf2_reg[28]/NET0131  & n18439 ;
  assign n18509 = \buf2_reg[20]/NET0131  & n18462 ;
  assign n18510 = ~n18508 & ~n18509 ;
  assign n18511 = n2970 & ~n18510 ;
  assign n18512 = ~n18237 & ~n18500 ;
  assign n18513 = \buf2_reg[4]/NET0131  & n18512 ;
  assign n18514 = ~n18511 & ~n18513 ;
  assign n18515 = ~n18503 & n18514 ;
  assign n18516 = ~n18507 & n18515 ;
  assign n18531 = n2571 & n18271 ;
  assign n18530 = ~\P3_InstQueue_reg[9][4]/NET0131  & ~n18271 ;
  assign n18532 = n2994 & ~n18530 ;
  assign n18533 = ~n18531 & n18532 ;
  assign n18521 = \buf2_reg[28]/NET0131  & n18462 ;
  assign n18522 = \buf2_reg[20]/NET0131  & n18233 ;
  assign n18523 = ~n18521 & ~n18522 ;
  assign n18524 = \P3_DataWidth_reg[1]/NET0131  & ~n18523 ;
  assign n18517 = \P3_InstQueue_reg[9][4]/NET0131  & ~n18235 ;
  assign n18518 = \buf2_reg[4]/NET0131  & n18235 ;
  assign n18519 = ~n18517 & ~n18518 ;
  assign n18525 = \P3_DataWidth_reg[1]/NET0131  & ~n18482 ;
  assign n18526 = ~n18519 & ~n18525 ;
  assign n18527 = ~n18524 & ~n18526 ;
  assign n18528 = n2959 & ~n18527 ;
  assign n18520 = n4415 & ~n18519 ;
  assign n18529 = \P3_InstQueue_reg[9][4]/NET0131  & ~n18217 ;
  assign n18534 = ~n18520 & ~n18529 ;
  assign n18535 = ~n18528 & n18534 ;
  assign n18536 = ~n18533 & n18535 ;
  assign n18538 = ~\P1_PhyAddrPointer_reg[31]/NET0131  & ~n10130 ;
  assign n18539 = \P1_PhyAddrPointer_reg[31]/NET0131  & n10130 ;
  assign n18540 = ~n18538 & ~n18539 ;
  assign n18541 = ~\P1_PhyAddrPointer_reg[0]/NET0131  & \P1_PhyAddrPointer_reg[1]/NET0131  ;
  assign n18542 = n10097 & n18541 ;
  assign n18543 = n10102 & n18542 ;
  assign n18544 = n18540 & ~n18543 ;
  assign n18546 = n13351 & ~n18544 ;
  assign n18545 = ~n13351 & n18544 ;
  assign n18547 = ~\P1_DataWidth_reg[1]/NET0131  & ~n18545 ;
  assign n18548 = ~n18546 & n18547 ;
  assign n18537 = \P1_DataWidth_reg[1]/NET0131  & ~\P1_rEIP_reg[14]/NET0131  ;
  assign n18549 = n2436 & ~n18537 ;
  assign n18550 = ~n18548 & n18549 ;
  assign n18554 = ~n2233 & ~n2301 ;
  assign n18555 = \P1_rEIP_reg[14]/NET0131  & ~n18554 ;
  assign n18558 = \P1_rEIP_reg[1]/NET0131  & \P1_rEIP_reg[2]/NET0131  ;
  assign n18559 = \P1_rEIP_reg[3]/NET0131  & n18558 ;
  assign n18560 = \P1_rEIP_reg[4]/NET0131  & n18559 ;
  assign n18561 = \P1_rEIP_reg[5]/NET0131  & n18560 ;
  assign n18562 = \P1_rEIP_reg[6]/NET0131  & n18561 ;
  assign n18563 = \P1_rEIP_reg[7]/NET0131  & n18562 ;
  assign n18564 = \P1_rEIP_reg[8]/NET0131  & n18563 ;
  assign n18565 = \P1_rEIP_reg[9]/NET0131  & n18564 ;
  assign n18566 = \P1_rEIP_reg[10]/NET0131  & n18565 ;
  assign n18567 = \P1_rEIP_reg[11]/NET0131  & n18566 ;
  assign n18568 = \P1_rEIP_reg[12]/NET0131  & n18567 ;
  assign n18569 = \P1_rEIP_reg[13]/NET0131  & n18568 ;
  assign n18570 = ~\P1_rEIP_reg[14]/NET0131  & ~n18569 ;
  assign n18571 = \P1_rEIP_reg[14]/NET0131  & n18569 ;
  assign n18572 = ~n18570 & ~n18571 ;
  assign n18573 = n2425 & ~n18572 ;
  assign n18574 = ~n2311 & n18573 ;
  assign n18556 = ~\P1_DataWidth_reg[1]/NET0131  & n2387 ;
  assign n18557 = ~\P1_EBX_reg[14]/NET0131  & ~n18556 ;
  assign n18575 = n2225 & ~n18557 ;
  assign n18576 = ~n18574 & n18575 ;
  assign n18577 = ~\P1_EBX_reg[0]/NET0131  & ~\P1_EBX_reg[1]/NET0131  ;
  assign n18578 = ~\P1_EBX_reg[2]/NET0131  & n18577 ;
  assign n18579 = ~\P1_EBX_reg[3]/NET0131  & n18578 ;
  assign n18580 = ~\P1_EBX_reg[4]/NET0131  & n18579 ;
  assign n18581 = ~\P1_EBX_reg[5]/NET0131  & n18580 ;
  assign n18582 = ~\P1_EBX_reg[6]/NET0131  & n18581 ;
  assign n18583 = ~\P1_EBX_reg[7]/NET0131  & n18582 ;
  assign n18584 = ~\P1_EBX_reg[8]/NET0131  & n18583 ;
  assign n18585 = ~\P1_EBX_reg[9]/NET0131  & n18584 ;
  assign n18586 = ~\P1_EBX_reg[10]/NET0131  & n18585 ;
  assign n18587 = ~\P1_EBX_reg[11]/NET0131  & n18586 ;
  assign n18588 = ~\P1_EBX_reg[12]/NET0131  & n18587 ;
  assign n18589 = ~\P1_EBX_reg[13]/NET0131  & n18588 ;
  assign n18590 = \P1_EBX_reg[31]/NET0131  & ~n18589 ;
  assign n18592 = \P1_EBX_reg[14]/NET0131  & ~n18590 ;
  assign n18591 = ~\P1_EBX_reg[14]/NET0131  & n18590 ;
  assign n18593 = ~n2425 & ~n18591 ;
  assign n18594 = ~n18592 & n18593 ;
  assign n18595 = n2222 & ~n18573 ;
  assign n18596 = ~n18594 & n18595 ;
  assign n18597 = ~n18576 & ~n18596 ;
  assign n18598 = ~n2301 & ~n18597 ;
  assign n18599 = ~n18555 & ~n18598 ;
  assign n18600 = n2432 & ~n18599 ;
  assign n18551 = ~n2445 & n3043 ;
  assign n18552 = ~n15769 & n18551 ;
  assign n18553 = \P1_rEIP_reg[14]/NET0131  & ~n18552 ;
  assign n18601 = \P1_PhyAddrPointer_reg[14]/NET0131  & n3028 ;
  assign n18602 = ~n5092 & ~n18601 ;
  assign n18603 = ~n18553 & n18602 ;
  assign n18604 = ~n18600 & n18603 ;
  assign n18605 = ~n18550 & n18604 ;
  assign n18607 = n10103 & n18542 ;
  assign n18608 = n18540 & ~n18607 ;
  assign n18610 = n12222 & ~n18608 ;
  assign n18609 = ~n12222 & n18608 ;
  assign n18611 = ~\P1_DataWidth_reg[1]/NET0131  & ~n18609 ;
  assign n18612 = ~n18610 & n18611 ;
  assign n18606 = \P1_DataWidth_reg[1]/NET0131  & ~\P1_rEIP_reg[15]/NET0131  ;
  assign n18613 = n2436 & ~n18606 ;
  assign n18614 = ~n18612 & n18613 ;
  assign n18616 = \P1_rEIP_reg[15]/NET0131  & ~n18554 ;
  assign n18618 = ~\P1_rEIP_reg[15]/NET0131  & ~n18571 ;
  assign n18619 = \P1_rEIP_reg[15]/NET0131  & n18571 ;
  assign n18620 = ~n18618 & ~n18619 ;
  assign n18621 = n2425 & ~n18620 ;
  assign n18622 = ~n2311 & n18621 ;
  assign n18617 = ~\P1_EBX_reg[15]/NET0131  & ~n18556 ;
  assign n18623 = n2225 & ~n18617 ;
  assign n18624 = ~n18622 & n18623 ;
  assign n18625 = ~\P1_EBX_reg[14]/NET0131  & n18589 ;
  assign n18626 = \P1_EBX_reg[31]/NET0131  & ~n18625 ;
  assign n18628 = \P1_EBX_reg[15]/NET0131  & ~n18626 ;
  assign n18627 = ~\P1_EBX_reg[15]/NET0131  & n18626 ;
  assign n18629 = ~n2425 & ~n18627 ;
  assign n18630 = ~n18628 & n18629 ;
  assign n18631 = n2222 & ~n18621 ;
  assign n18632 = ~n18630 & n18631 ;
  assign n18633 = ~n18624 & ~n18632 ;
  assign n18634 = ~n2301 & ~n18633 ;
  assign n18635 = ~n18616 & ~n18634 ;
  assign n18636 = n2432 & ~n18635 ;
  assign n18615 = \P1_rEIP_reg[15]/NET0131  & ~n18552 ;
  assign n18637 = \P1_PhyAddrPointer_reg[15]/NET0131  & n3028 ;
  assign n18638 = ~n5092 & ~n18637 ;
  assign n18639 = ~n18615 & n18638 ;
  assign n18640 = ~n18636 & n18639 ;
  assign n18641 = ~n18614 & n18640 ;
  assign n18643 = \P1_PhyAddrPointer_reg[15]/NET0131  & n18607 ;
  assign n18644 = n18540 & ~n18643 ;
  assign n18645 = ~n13360 & ~n18644 ;
  assign n18646 = n13360 & n18644 ;
  assign n18647 = ~n18645 & ~n18646 ;
  assign n18648 = ~\P1_DataWidth_reg[1]/NET0131  & ~n18647 ;
  assign n18642 = \P1_DataWidth_reg[1]/NET0131  & ~\P1_rEIP_reg[16]/NET0131  ;
  assign n18649 = n2436 & ~n18642 ;
  assign n18650 = ~n18648 & n18649 ;
  assign n18652 = \P1_rEIP_reg[16]/NET0131  & ~n18554 ;
  assign n18654 = ~\P1_rEIP_reg[16]/NET0131  & ~n18619 ;
  assign n18655 = \P1_rEIP_reg[16]/NET0131  & n18619 ;
  assign n18656 = ~n18654 & ~n18655 ;
  assign n18657 = n2425 & ~n18656 ;
  assign n18658 = ~n2311 & n18657 ;
  assign n18653 = ~\P1_EBX_reg[16]/NET0131  & ~n18556 ;
  assign n18659 = n2225 & ~n18653 ;
  assign n18660 = ~n18658 & n18659 ;
  assign n18661 = ~\P1_EBX_reg[14]/NET0131  & ~\P1_EBX_reg[15]/NET0131  ;
  assign n18662 = n18589 & n18661 ;
  assign n18663 = \P1_EBX_reg[31]/NET0131  & ~n18662 ;
  assign n18665 = ~\P1_EBX_reg[16]/NET0131  & n18663 ;
  assign n18664 = \P1_EBX_reg[16]/NET0131  & ~n18663 ;
  assign n18666 = ~n2425 & ~n18664 ;
  assign n18667 = ~n18665 & n18666 ;
  assign n18668 = n2222 & ~n18657 ;
  assign n18669 = ~n18667 & n18668 ;
  assign n18670 = ~n18660 & ~n18669 ;
  assign n18671 = ~n2301 & ~n18670 ;
  assign n18672 = ~n18652 & ~n18671 ;
  assign n18673 = n2432 & ~n18672 ;
  assign n18651 = \P1_rEIP_reg[16]/NET0131  & ~n18552 ;
  assign n18674 = \P1_PhyAddrPointer_reg[16]/NET0131  & n3028 ;
  assign n18675 = ~n5092 & ~n18674 ;
  assign n18676 = ~n18651 & n18675 ;
  assign n18677 = ~n18673 & n18676 ;
  assign n18678 = ~n18650 & n18677 ;
  assign n18680 = \P1_PhyAddrPointer_reg[16]/NET0131  & n18643 ;
  assign n18681 = n18540 & ~n18680 ;
  assign n18683 = ~n13405 & n18681 ;
  assign n18682 = n13405 & ~n18681 ;
  assign n18684 = ~\P1_DataWidth_reg[1]/NET0131  & ~n18682 ;
  assign n18685 = ~n18683 & n18684 ;
  assign n18679 = \P1_DataWidth_reg[1]/NET0131  & ~\P1_rEIP_reg[17]/NET0131  ;
  assign n18686 = n2436 & ~n18679 ;
  assign n18687 = ~n18685 & n18686 ;
  assign n18695 = ~\P1_rEIP_reg[17]/NET0131  & ~n18655 ;
  assign n18696 = \P1_rEIP_reg[17]/NET0131  & n18655 ;
  assign n18697 = ~n18695 & ~n18696 ;
  assign n18698 = n2425 & ~n18697 ;
  assign n18699 = ~\P1_EBX_reg[17]/NET0131  & ~n2425 ;
  assign n18700 = n2312 & ~n18699 ;
  assign n18701 = ~n18698 & n18700 ;
  assign n18692 = ~n2301 & n2311 ;
  assign n18693 = \P1_EBX_reg[17]/NET0131  & n18692 ;
  assign n18694 = \P1_rEIP_reg[17]/NET0131  & n2301 ;
  assign n18702 = ~n18693 & ~n18694 ;
  assign n18703 = ~n18701 & n18702 ;
  assign n18704 = n2225 & ~n18703 ;
  assign n18689 = n2225 & ~n2231 ;
  assign n18690 = ~n18554 & ~n18689 ;
  assign n18691 = \P1_rEIP_reg[17]/NET0131  & n18690 ;
  assign n18705 = ~\P1_EBX_reg[16]/NET0131  & n18662 ;
  assign n18706 = \P1_EBX_reg[31]/NET0131  & ~n18705 ;
  assign n18708 = ~\P1_EBX_reg[17]/NET0131  & n18706 ;
  assign n18707 = \P1_EBX_reg[17]/NET0131  & ~n18706 ;
  assign n18709 = ~n2425 & ~n18707 ;
  assign n18710 = ~n18708 & n18709 ;
  assign n18711 = n7246 & ~n18698 ;
  assign n18712 = ~n18710 & n18711 ;
  assign n18713 = ~n18691 & ~n18712 ;
  assign n18714 = ~n18704 & n18713 ;
  assign n18715 = n2432 & ~n18714 ;
  assign n18688 = \P1_rEIP_reg[17]/NET0131  & ~n18552 ;
  assign n18716 = \P1_PhyAddrPointer_reg[17]/NET0131  & n3028 ;
  assign n18717 = ~n5092 & ~n18716 ;
  assign n18718 = ~n18688 & n18717 ;
  assign n18719 = ~n18715 & n18718 ;
  assign n18720 = ~n18687 & n18719 ;
  assign n18744 = n10124 & n18643 ;
  assign n18745 = n18540 & ~n18744 ;
  assign n18746 = ~n13421 & ~n18745 ;
  assign n18747 = n13421 & n18745 ;
  assign n18748 = ~n18746 & ~n18747 ;
  assign n18749 = ~\P1_DataWidth_reg[1]/NET0131  & ~n18748 ;
  assign n18743 = \P1_DataWidth_reg[1]/NET0131  & ~\P1_rEIP_reg[18]/NET0131  ;
  assign n18750 = n2436 & ~n18743 ;
  assign n18751 = ~n18749 & n18750 ;
  assign n18722 = \P1_rEIP_reg[18]/NET0131  & ~n18554 ;
  assign n18723 = ~\P1_EBX_reg[18]/NET0131  & ~n18556 ;
  assign n18724 = n15990 & ~n18723 ;
  assign n18725 = ~\P1_EBX_reg[17]/NET0131  & n18705 ;
  assign n18726 = \P1_EBX_reg[31]/NET0131  & ~n18725 ;
  assign n18728 = ~\P1_EBX_reg[18]/NET0131  & n18726 ;
  assign n18727 = \P1_EBX_reg[18]/NET0131  & ~n18726 ;
  assign n18729 = ~n2425 & ~n18727 ;
  assign n18730 = ~n18728 & n18729 ;
  assign n18731 = n7246 & ~n18730 ;
  assign n18732 = ~n18724 & ~n18731 ;
  assign n18733 = ~\P1_rEIP_reg[18]/NET0131  & ~n18696 ;
  assign n18734 = \P1_rEIP_reg[18]/NET0131  & n18696 ;
  assign n18735 = ~n18733 & ~n18734 ;
  assign n18736 = n2311 & n18724 ;
  assign n18737 = n2425 & ~n18736 ;
  assign n18738 = ~n18735 & n18737 ;
  assign n18739 = ~n18732 & ~n18738 ;
  assign n18740 = ~n18722 & ~n18739 ;
  assign n18741 = n2432 & ~n18740 ;
  assign n18721 = \P1_rEIP_reg[18]/NET0131  & ~n18552 ;
  assign n18742 = \P1_PhyAddrPointer_reg[18]/NET0131  & n3028 ;
  assign n18752 = ~n5092 & ~n18742 ;
  assign n18753 = ~n18721 & n18752 ;
  assign n18754 = ~n18741 & n18753 ;
  assign n18755 = ~n18751 & n18754 ;
  assign n18757 = \P1_PhyAddrPointer_reg[18]/NET0131  & n18744 ;
  assign n18758 = n18540 & ~n18757 ;
  assign n18760 = n12241 & ~n18758 ;
  assign n18759 = ~n12241 & n18758 ;
  assign n18761 = ~\P1_DataWidth_reg[1]/NET0131  & ~n18759 ;
  assign n18762 = ~n18760 & n18761 ;
  assign n18756 = \P1_DataWidth_reg[1]/NET0131  & ~\P1_rEIP_reg[19]/NET0131  ;
  assign n18763 = n2436 & ~n18756 ;
  assign n18764 = ~n18762 & n18763 ;
  assign n18769 = \P1_rEIP_reg[19]/NET0131  & n18734 ;
  assign n18770 = ~\P1_rEIP_reg[19]/NET0131  & ~n18734 ;
  assign n18771 = ~n18769 & ~n18770 ;
  assign n18772 = n2425 & ~n18771 ;
  assign n18773 = ~\P1_EBX_reg[19]/NET0131  & ~n2425 ;
  assign n18774 = n2312 & ~n18773 ;
  assign n18775 = ~n18772 & n18774 ;
  assign n18767 = \P1_rEIP_reg[19]/NET0131  & n2301 ;
  assign n18768 = \P1_EBX_reg[19]/NET0131  & n18692 ;
  assign n18776 = ~n18767 & ~n18768 ;
  assign n18777 = ~n18775 & n18776 ;
  assign n18778 = n2225 & ~n18777 ;
  assign n18766 = \P1_rEIP_reg[19]/NET0131  & n18690 ;
  assign n18779 = ~\P1_EBX_reg[17]/NET0131  & ~\P1_EBX_reg[18]/NET0131  ;
  assign n18780 = n18705 & n18779 ;
  assign n18781 = \P1_EBX_reg[31]/NET0131  & ~n18780 ;
  assign n18783 = ~\P1_EBX_reg[19]/NET0131  & n18781 ;
  assign n18782 = \P1_EBX_reg[19]/NET0131  & ~n18781 ;
  assign n18784 = ~n2425 & ~n18782 ;
  assign n18785 = ~n18783 & n18784 ;
  assign n18786 = n7246 & ~n18772 ;
  assign n18787 = ~n18785 & n18786 ;
  assign n18788 = ~n18766 & ~n18787 ;
  assign n18789 = ~n18778 & n18788 ;
  assign n18790 = n2432 & ~n18789 ;
  assign n18765 = \P1_rEIP_reg[19]/NET0131  & ~n18552 ;
  assign n18791 = \P1_PhyAddrPointer_reg[19]/NET0131  & n3028 ;
  assign n18792 = ~n5092 & ~n18791 ;
  assign n18793 = ~n18765 & n18792 ;
  assign n18794 = ~n18790 & n18793 ;
  assign n18795 = ~n18764 & n18794 ;
  assign n18797 = \P1_PhyAddrPointer_reg[0]/NET0131  & n18540 ;
  assign n18798 = \P1_PhyAddrPointer_reg[1]/NET0131  & ~n18797 ;
  assign n18799 = ~\P1_PhyAddrPointer_reg[1]/NET0131  & n18797 ;
  assign n18800 = ~n18798 & ~n18799 ;
  assign n18801 = ~\P1_DataWidth_reg[1]/NET0131  & ~n18800 ;
  assign n18796 = \P1_DataWidth_reg[1]/NET0131  & ~\P1_rEIP_reg[1]/NET0131  ;
  assign n18802 = n2436 & ~n18796 ;
  assign n18803 = ~n18801 & n18802 ;
  assign n18809 = \P1_rEIP_reg[1]/NET0131  & ~n18554 ;
  assign n18816 = ~n15364 & ~n18577 ;
  assign n18817 = \P1_EBX_reg[31]/NET0131  & ~n18816 ;
  assign n18815 = ~\P1_EBX_reg[1]/NET0131  & ~\P1_EBX_reg[31]/NET0131  ;
  assign n18818 = ~n2425 & ~n18815 ;
  assign n18819 = ~n18817 & n18818 ;
  assign n18811 = ~\P1_DataWidth_reg[1]/NET0131  & ~\P1_rEIP_reg[1]/NET0131  ;
  assign n18820 = ~n2317 & n18811 ;
  assign n18821 = ~n18819 & ~n18820 ;
  assign n18822 = n7246 & ~n18821 ;
  assign n18807 = n2231 & ~n2301 ;
  assign n18808 = ~n2399 & n18807 ;
  assign n18810 = \P1_EBX_reg[1]/NET0131  & ~n18556 ;
  assign n18812 = n2387 & n18811 ;
  assign n18813 = ~n18810 & ~n18812 ;
  assign n18814 = n15990 & ~n18813 ;
  assign n18823 = ~n18808 & ~n18814 ;
  assign n18824 = ~n18822 & n18823 ;
  assign n18825 = ~n18809 & n18824 ;
  assign n18826 = n2432 & ~n18825 ;
  assign n18804 = \P1_PhyAddrPointer_reg[1]/NET0131  & n3028 ;
  assign n18805 = ~n5095 & n16260 ;
  assign n18806 = \P1_rEIP_reg[1]/NET0131  & ~n18805 ;
  assign n18827 = ~n18804 & ~n18806 ;
  assign n18828 = ~n18826 & n18827 ;
  assign n18829 = ~n18803 & n18828 ;
  assign n18831 = n12240 & n18643 ;
  assign n18832 = n18540 & ~n18831 ;
  assign n18834 = ~n12278 & n18832 ;
  assign n18833 = n12278 & ~n18832 ;
  assign n18835 = ~\P1_DataWidth_reg[1]/NET0131  & ~n18833 ;
  assign n18836 = ~n18834 & n18835 ;
  assign n18830 = \P1_DataWidth_reg[1]/NET0131  & ~\P1_rEIP_reg[20]/NET0131  ;
  assign n18837 = n2436 & ~n18830 ;
  assign n18838 = ~n18836 & n18837 ;
  assign n18840 = \P1_rEIP_reg[20]/NET0131  & ~n18554 ;
  assign n18841 = ~\P1_EBX_reg[20]/NET0131  & ~n18556 ;
  assign n18842 = n2225 & ~n18841 ;
  assign n18843 = ~\P1_EBX_reg[19]/NET0131  & n18780 ;
  assign n18844 = \P1_EBX_reg[31]/NET0131  & ~n18843 ;
  assign n18846 = ~\P1_EBX_reg[20]/NET0131  & n18844 ;
  assign n18845 = \P1_EBX_reg[20]/NET0131  & ~n18844 ;
  assign n18847 = ~n2425 & ~n18845 ;
  assign n18848 = ~n18846 & n18847 ;
  assign n18849 = n2222 & ~n18848 ;
  assign n18850 = ~n18842 & ~n18849 ;
  assign n18852 = ~\P1_rEIP_reg[20]/NET0131  & ~n18769 ;
  assign n18853 = \P1_rEIP_reg[19]/NET0131  & \P1_rEIP_reg[20]/NET0131  ;
  assign n18854 = n18734 & n18853 ;
  assign n18855 = ~n18852 & ~n18854 ;
  assign n18851 = n2311 & n18842 ;
  assign n18856 = n2425 & ~n18851 ;
  assign n18857 = ~n18855 & n18856 ;
  assign n18858 = ~n2301 & ~n18857 ;
  assign n18859 = ~n18850 & n18858 ;
  assign n18860 = ~n18840 & ~n18859 ;
  assign n18861 = n2432 & ~n18860 ;
  assign n18839 = \P1_PhyAddrPointer_reg[20]/NET0131  & n3028 ;
  assign n18862 = \P1_rEIP_reg[20]/NET0131  & ~n18805 ;
  assign n18863 = ~n18839 & ~n18862 ;
  assign n18864 = ~n18861 & n18863 ;
  assign n18865 = ~n18838 & n18864 ;
  assign n18893 = n12277 & n18643 ;
  assign n18894 = n18540 & ~n18893 ;
  assign n18896 = ~n13435 & n18894 ;
  assign n18895 = n13435 & ~n18894 ;
  assign n18897 = ~\P1_DataWidth_reg[1]/NET0131  & ~n18895 ;
  assign n18898 = ~n18896 & n18897 ;
  assign n18892 = \P1_DataWidth_reg[1]/NET0131  & ~\P1_rEIP_reg[21]/NET0131  ;
  assign n18899 = n2436 & ~n18892 ;
  assign n18900 = ~n18898 & n18899 ;
  assign n18871 = ~\P1_rEIP_reg[21]/NET0131  & ~n18854 ;
  assign n18872 = \P1_rEIP_reg[21]/NET0131  & n18854 ;
  assign n18873 = ~n18871 & ~n18872 ;
  assign n18874 = n2425 & ~n18873 ;
  assign n18875 = ~\P1_EBX_reg[21]/NET0131  & ~n2425 ;
  assign n18876 = n2312 & ~n18875 ;
  assign n18877 = ~n18874 & n18876 ;
  assign n18869 = \P1_EBX_reg[21]/NET0131  & n18692 ;
  assign n18870 = \P1_rEIP_reg[21]/NET0131  & n2301 ;
  assign n18878 = ~n18869 & ~n18870 ;
  assign n18879 = ~n18877 & n18878 ;
  assign n18880 = n2225 & ~n18879 ;
  assign n18868 = \P1_rEIP_reg[21]/NET0131  & n18690 ;
  assign n18881 = ~\P1_EBX_reg[20]/NET0131  & n18843 ;
  assign n18882 = \P1_EBX_reg[31]/NET0131  & ~n18881 ;
  assign n18884 = ~\P1_EBX_reg[21]/NET0131  & n18882 ;
  assign n18883 = \P1_EBX_reg[21]/NET0131  & ~n18882 ;
  assign n18885 = ~n2425 & ~n18883 ;
  assign n18886 = ~n18884 & n18885 ;
  assign n18887 = n7246 & ~n18874 ;
  assign n18888 = ~n18886 & n18887 ;
  assign n18889 = ~n18868 & ~n18888 ;
  assign n18890 = ~n18880 & n18889 ;
  assign n18891 = n2432 & ~n18890 ;
  assign n18866 = \P1_PhyAddrPointer_reg[21]/NET0131  & n3028 ;
  assign n18867 = \P1_rEIP_reg[21]/NET0131  & ~n18805 ;
  assign n18901 = ~n18866 & ~n18867 ;
  assign n18902 = ~n18891 & n18901 ;
  assign n18903 = ~n18900 & n18902 ;
  assign n18929 = n10125 & n18643 ;
  assign n18930 = n18540 & ~n18929 ;
  assign n18932 = n12311 & ~n18930 ;
  assign n18931 = ~n12311 & n18930 ;
  assign n18933 = ~\P1_DataWidth_reg[1]/NET0131  & ~n18931 ;
  assign n18934 = ~n18932 & n18933 ;
  assign n18928 = \P1_DataWidth_reg[1]/NET0131  & ~\P1_rEIP_reg[22]/NET0131  ;
  assign n18935 = n2436 & ~n18928 ;
  assign n18936 = ~n18934 & n18935 ;
  assign n18904 = \P1_rEIP_reg[22]/NET0131  & ~n18554 ;
  assign n18908 = ~\P1_EBX_reg[22]/NET0131  & ~n18556 ;
  assign n18909 = n2225 & ~n18908 ;
  assign n18913 = ~\P1_EBX_reg[20]/NET0131  & ~\P1_EBX_reg[21]/NET0131  ;
  assign n18914 = n18843 & n18913 ;
  assign n18915 = \P1_EBX_reg[31]/NET0131  & ~n18914 ;
  assign n18917 = ~\P1_EBX_reg[22]/NET0131  & n18915 ;
  assign n18916 = \P1_EBX_reg[22]/NET0131  & ~n18915 ;
  assign n18918 = ~n2425 & ~n18916 ;
  assign n18919 = ~n18917 & n18918 ;
  assign n18920 = n2222 & ~n18919 ;
  assign n18921 = ~n18909 & ~n18920 ;
  assign n18905 = ~\P1_rEIP_reg[22]/NET0131  & ~n18872 ;
  assign n18906 = \P1_rEIP_reg[22]/NET0131  & n18872 ;
  assign n18907 = ~n18905 & ~n18906 ;
  assign n18910 = n2311 & n18909 ;
  assign n18911 = n2425 & ~n18910 ;
  assign n18912 = ~n18907 & n18911 ;
  assign n18922 = ~n2301 & ~n18912 ;
  assign n18923 = ~n18921 & n18922 ;
  assign n18924 = ~n18904 & ~n18923 ;
  assign n18925 = n2432 & ~n18924 ;
  assign n18926 = \P1_PhyAddrPointer_reg[22]/NET0131  & n3028 ;
  assign n18927 = \P1_rEIP_reg[22]/NET0131  & ~n18805 ;
  assign n18937 = ~n18926 & ~n18927 ;
  assign n18938 = ~n18925 & n18937 ;
  assign n18939 = ~n18936 & n18938 ;
  assign n18969 = n11252 & n18643 ;
  assign n18970 = n18540 & ~n18969 ;
  assign n18972 = ~n11255 & n18970 ;
  assign n18971 = n11255 & ~n18970 ;
  assign n18973 = ~\P1_DataWidth_reg[1]/NET0131  & ~n18971 ;
  assign n18974 = ~n18972 & n18973 ;
  assign n18968 = \P1_DataWidth_reg[1]/NET0131  & ~\P1_rEIP_reg[23]/NET0131  ;
  assign n18975 = n2436 & ~n18968 ;
  assign n18976 = ~n18974 & n18975 ;
  assign n18947 = ~\P1_rEIP_reg[23]/NET0131  & ~n18906 ;
  assign n18948 = \P1_rEIP_reg[21]/NET0131  & \P1_rEIP_reg[22]/NET0131  ;
  assign n18949 = \P1_rEIP_reg[23]/NET0131  & n18948 ;
  assign n18950 = n18854 & n18949 ;
  assign n18951 = ~n18947 & ~n18950 ;
  assign n18952 = n2425 & ~n18951 ;
  assign n18953 = ~\P1_EBX_reg[23]/NET0131  & ~n2425 ;
  assign n18954 = n2426 & ~n18953 ;
  assign n18955 = ~\P1_EBX_reg[22]/NET0131  & n18913 ;
  assign n18956 = n18843 & n18955 ;
  assign n18957 = \P1_EBX_reg[31]/NET0131  & ~n18956 ;
  assign n18959 = ~\P1_EBX_reg[23]/NET0131  & n18957 ;
  assign n18958 = \P1_EBX_reg[23]/NET0131  & ~n18957 ;
  assign n18960 = ~n2425 & ~n18958 ;
  assign n18961 = ~n18959 & n18960 ;
  assign n18962 = n7246 & ~n18961 ;
  assign n18963 = ~n18954 & ~n18962 ;
  assign n18964 = ~n18952 & ~n18963 ;
  assign n18942 = \P1_rEIP_reg[23]/NET0131  & n18690 ;
  assign n18943 = \P1_EBX_reg[23]/NET0131  & n18692 ;
  assign n18944 = \P1_rEIP_reg[23]/NET0131  & n2301 ;
  assign n18945 = ~n18943 & ~n18944 ;
  assign n18946 = n2225 & ~n18945 ;
  assign n18965 = ~n18942 & ~n18946 ;
  assign n18966 = ~n18964 & n18965 ;
  assign n18967 = n2432 & ~n18966 ;
  assign n18940 = \P1_rEIP_reg[23]/NET0131  & ~n18805 ;
  assign n18941 = \P1_PhyAddrPointer_reg[23]/NET0131  & n3028 ;
  assign n18977 = ~n18940 & ~n18941 ;
  assign n18978 = ~n18967 & n18977 ;
  assign n18979 = ~n18976 & n18978 ;
  assign n18981 = ~\P2_PhyAddrPointer_reg[0]/NET0131  & n12373 ;
  assign n18982 = ~n9003 & ~n18981 ;
  assign n18984 = ~n14636 & n18982 ;
  assign n18983 = n14636 & ~n18982 ;
  assign n18985 = ~\P2_DataWidth_reg[1]/NET0131  & ~n18983 ;
  assign n18986 = ~n18984 & n18985 ;
  assign n18980 = \P2_DataWidth_reg[1]/NET0131  & ~\P2_rEIP_reg[10]/NET0131  ;
  assign n18987 = n1931 & ~n18980 ;
  assign n18988 = ~n18986 & n18987 ;
  assign n18991 = \P2_rEIP_reg[10]/NET0131  & ~n16555 ;
  assign n18992 = \P2_EBX_reg[31]/NET0131  & ~n16568 ;
  assign n18994 = \P2_EBX_reg[10]/NET0131  & n18992 ;
  assign n18993 = ~\P2_EBX_reg[10]/NET0131  & ~n18992 ;
  assign n18995 = ~n1920 & ~n18993 ;
  assign n18996 = ~n18994 & n18995 ;
  assign n18997 = \P2_rEIP_reg[10]/NET0131  & n16531 ;
  assign n18998 = ~\P2_rEIP_reg[10]/NET0131  & ~n16531 ;
  assign n18999 = ~n18997 & ~n18998 ;
  assign n19000 = ~\P2_DataWidth_reg[1]/NET0131  & n18999 ;
  assign n19001 = ~n1805 & n19000 ;
  assign n19002 = ~n18996 & ~n19001 ;
  assign n19003 = n1742 & ~n19002 ;
  assign n19004 = \P2_EBX_reg[10]/NET0131  & ~n16558 ;
  assign n19005 = n1820 & n19000 ;
  assign n19006 = ~n19004 & ~n19005 ;
  assign n19007 = n1743 & ~n19006 ;
  assign n19008 = ~n19003 & ~n19007 ;
  assign n19009 = ~n1810 & ~n19008 ;
  assign n19010 = ~n18991 & ~n19009 ;
  assign n19011 = n1927 & ~n19010 ;
  assign n18989 = n1937 & n3041 ;
  assign n18990 = \P2_rEIP_reg[10]/NET0131  & ~n18989 ;
  assign n19012 = \P2_PhyAddrPointer_reg[10]/NET0131  & n2987 ;
  assign n19013 = ~n3113 & ~n19012 ;
  assign n19014 = ~n18990 & n19013 ;
  assign n19015 = ~n19011 & n19014 ;
  assign n19016 = ~n18988 & n19015 ;
  assign n19044 = n10111 & n18929 ;
  assign n19045 = n18540 & ~n19044 ;
  assign n19046 = ~n12334 & ~n19045 ;
  assign n19047 = n12334 & n19045 ;
  assign n19048 = ~n19046 & ~n19047 ;
  assign n19049 = ~\P1_DataWidth_reg[1]/NET0131  & ~n19048 ;
  assign n19043 = \P1_DataWidth_reg[1]/NET0131  & ~\P1_rEIP_reg[24]/NET0131  ;
  assign n19050 = n2436 & ~n19043 ;
  assign n19051 = ~n19049 & n19050 ;
  assign n19019 = ~\P1_rEIP_reg[24]/NET0131  & ~n18950 ;
  assign n19020 = \P1_rEIP_reg[24]/NET0131  & n18950 ;
  assign n19021 = ~n19019 & ~n19020 ;
  assign n19022 = n2425 & ~n19021 ;
  assign n19032 = ~\P1_EBX_reg[24]/NET0131  & ~n2425 ;
  assign n19033 = n2312 & ~n19032 ;
  assign n19034 = ~n19022 & n19033 ;
  assign n19035 = \P1_EBX_reg[24]/NET0131  & n18692 ;
  assign n19036 = \P1_rEIP_reg[24]/NET0131  & n2301 ;
  assign n19037 = ~n19035 & ~n19036 ;
  assign n19038 = ~n19034 & n19037 ;
  assign n19039 = n2225 & ~n19038 ;
  assign n19023 = ~\P1_EBX_reg[23]/NET0131  & n18956 ;
  assign n19024 = \P1_EBX_reg[31]/NET0131  & ~n19023 ;
  assign n19026 = ~\P1_EBX_reg[24]/NET0131  & n19024 ;
  assign n19025 = \P1_EBX_reg[24]/NET0131  & ~n19024 ;
  assign n19027 = ~n2425 & ~n19025 ;
  assign n19028 = ~n19026 & n19027 ;
  assign n19029 = n7246 & ~n19022 ;
  assign n19030 = ~n19028 & n19029 ;
  assign n19031 = \P1_rEIP_reg[24]/NET0131  & n18690 ;
  assign n19040 = ~n19030 & ~n19031 ;
  assign n19041 = ~n19039 & n19040 ;
  assign n19042 = n2432 & ~n19041 ;
  assign n19017 = \P1_rEIP_reg[24]/NET0131  & ~n18805 ;
  assign n19018 = \P1_PhyAddrPointer_reg[24]/NET0131  & n3028 ;
  assign n19052 = ~n19017 & ~n19018 ;
  assign n19053 = ~n19042 & n19052 ;
  assign n19054 = ~n19051 & n19053 ;
  assign n19056 = ~n9003 & ~n16514 ;
  assign n19057 = ~n9003 & ~n12367 ;
  assign n19058 = ~n19056 & ~n19057 ;
  assign n19060 = ~n12377 & ~n19058 ;
  assign n19059 = n12377 & n19058 ;
  assign n19061 = ~\P2_DataWidth_reg[1]/NET0131  & ~n19059 ;
  assign n19062 = ~n19060 & n19061 ;
  assign n19055 = \P2_DataWidth_reg[1]/NET0131  & ~\P2_rEIP_reg[11]/NET0131  ;
  assign n19063 = n1931 & ~n19055 ;
  assign n19064 = ~n19062 & n19063 ;
  assign n19072 = \P2_EBX_reg[31]/NET0131  & ~n16569 ;
  assign n19073 = ~n16559 & n19072 ;
  assign n19071 = ~n16559 & ~n16589 ;
  assign n19074 = \P2_EBX_reg[11]/NET0131  & ~n19071 ;
  assign n19075 = ~n19073 & n19074 ;
  assign n19066 = ~\P2_rEIP_reg[11]/NET0131  & ~n18997 ;
  assign n19067 = n16523 & n16531 ;
  assign n19068 = ~n19066 & ~n19067 ;
  assign n19069 = n16553 & n19068 ;
  assign n19070 = \P2_rEIP_reg[11]/NET0131  & ~n16555 ;
  assign n19076 = ~\P2_EBX_reg[11]/NET0131  & n19072 ;
  assign n19077 = n16589 & n19076 ;
  assign n19078 = ~n19070 & ~n19077 ;
  assign n19079 = ~n19069 & n19078 ;
  assign n19080 = ~n19075 & n19079 ;
  assign n19081 = n1927 & ~n19080 ;
  assign n19065 = \P2_rEIP_reg[11]/NET0131  & ~n18989 ;
  assign n19082 = \P2_PhyAddrPointer_reg[11]/NET0131  & n2987 ;
  assign n19083 = ~n3113 & ~n19082 ;
  assign n19084 = ~n19065 & n19083 ;
  assign n19085 = ~n19081 & n19084 ;
  assign n19086 = ~n19064 & n19085 ;
  assign n19114 = \P1_PhyAddrPointer_reg[24]/NET0131  & n19044 ;
  assign n19115 = n18540 & ~n19114 ;
  assign n19117 = ~n13486 & n19115 ;
  assign n19116 = n13486 & ~n19115 ;
  assign n19118 = ~\P1_DataWidth_reg[1]/NET0131  & ~n19116 ;
  assign n19119 = ~n19117 & n19118 ;
  assign n19113 = \P1_DataWidth_reg[1]/NET0131  & ~\P1_rEIP_reg[25]/NET0131  ;
  assign n19120 = n2436 & ~n19113 ;
  assign n19121 = ~n19119 & n19120 ;
  assign n19101 = \P1_EBX_reg[24]/NET0131  & \P1_EBX_reg[31]/NET0131  ;
  assign n19102 = ~n19024 & ~n19101 ;
  assign n19103 = \P1_EBX_reg[25]/NET0131  & ~n19102 ;
  assign n19104 = ~\P1_EBX_reg[25]/NET0131  & n19102 ;
  assign n19105 = ~n19103 & ~n19104 ;
  assign n19106 = ~n2425 & ~n19105 ;
  assign n19091 = ~\P1_rEIP_reg[25]/NET0131  & ~n19020 ;
  assign n19092 = \P1_rEIP_reg[24]/NET0131  & n18949 ;
  assign n19093 = \P1_rEIP_reg[18]/NET0131  & \P1_rEIP_reg[25]/NET0131  ;
  assign n19094 = n18853 & n19093 ;
  assign n19095 = n19092 & n19094 ;
  assign n19096 = n18696 & n19095 ;
  assign n19097 = ~n19091 & ~n19096 ;
  assign n19107 = n2425 & ~n19097 ;
  assign n19108 = n7246 & ~n19107 ;
  assign n19109 = ~n19106 & n19108 ;
  assign n19089 = \P1_rEIP_reg[25]/NET0131  & ~n18554 ;
  assign n19098 = n18556 & ~n19097 ;
  assign n19090 = ~\P1_EBX_reg[25]/NET0131  & ~n18556 ;
  assign n19099 = n15990 & ~n19090 ;
  assign n19100 = ~n19098 & n19099 ;
  assign n19110 = ~n19089 & ~n19100 ;
  assign n19111 = ~n19109 & n19110 ;
  assign n19112 = n2432 & ~n19111 ;
  assign n19087 = \P1_rEIP_reg[25]/NET0131  & ~n18805 ;
  assign n19088 = \P1_PhyAddrPointer_reg[25]/NET0131  & n3028 ;
  assign n19122 = ~n19087 & ~n19088 ;
  assign n19123 = ~n19112 & n19122 ;
  assign n19124 = ~n19121 & n19123 ;
  assign n19126 = n8968 & n16514 ;
  assign n19127 = ~n9003 & ~n19126 ;
  assign n19129 = n13542 & ~n19127 ;
  assign n19128 = ~n13542 & n19127 ;
  assign n19130 = ~\P2_DataWidth_reg[1]/NET0131  & ~n19128 ;
  assign n19131 = ~n19129 & n19130 ;
  assign n19125 = \P2_DataWidth_reg[1]/NET0131  & ~\P2_rEIP_reg[12]/NET0131  ;
  assign n19132 = n1931 & ~n19125 ;
  assign n19133 = ~n19131 & n19132 ;
  assign n19135 = \P2_rEIP_reg[12]/NET0131  & ~n16555 ;
  assign n19136 = \P2_EBX_reg[12]/NET0131  & ~n16558 ;
  assign n19137 = ~\P2_rEIP_reg[12]/NET0131  & ~n19067 ;
  assign n19138 = ~n16533 & ~n19137 ;
  assign n19139 = n1920 & n19138 ;
  assign n19140 = ~n1819 & n19139 ;
  assign n19141 = ~n19136 & ~n19140 ;
  assign n19142 = n1743 & ~n19141 ;
  assign n19143 = \P2_EBX_reg[31]/NET0131  & ~n16570 ;
  assign n19145 = \P2_EBX_reg[12]/NET0131  & n19143 ;
  assign n19144 = ~\P2_EBX_reg[12]/NET0131  & ~n19143 ;
  assign n19146 = ~n1920 & ~n19144 ;
  assign n19147 = ~n19145 & n19146 ;
  assign n19148 = ~n19139 & ~n19147 ;
  assign n19149 = n1742 & ~n19148 ;
  assign n19150 = ~n19142 & ~n19149 ;
  assign n19151 = ~n1810 & ~n19150 ;
  assign n19152 = ~n19135 & ~n19151 ;
  assign n19153 = n1927 & ~n19152 ;
  assign n19134 = \P2_rEIP_reg[12]/NET0131  & ~n18989 ;
  assign n19154 = \P2_PhyAddrPointer_reg[12]/NET0131  & n2987 ;
  assign n19155 = ~n3113 & ~n19154 ;
  assign n19156 = ~n19134 & n19155 ;
  assign n19157 = ~n19153 & n19156 ;
  assign n19158 = ~n19133 & n19157 ;
  assign n19160 = n13536 & n16514 ;
  assign n19161 = ~n9003 & ~n19160 ;
  assign n19163 = n13560 & ~n19161 ;
  assign n19162 = ~n13560 & n19161 ;
  assign n19164 = ~\P2_DataWidth_reg[1]/NET0131  & ~n19162 ;
  assign n19165 = ~n19163 & n19164 ;
  assign n19159 = \P2_DataWidth_reg[1]/NET0131  & ~\P2_rEIP_reg[13]/NET0131  ;
  assign n19166 = n1931 & ~n19159 ;
  assign n19167 = ~n19165 & n19166 ;
  assign n19169 = \P2_rEIP_reg[13]/NET0131  & ~n16555 ;
  assign n19171 = ~\P2_rEIP_reg[13]/NET0131  & ~n16533 ;
  assign n19172 = \P2_rEIP_reg[13]/NET0131  & n16533 ;
  assign n19173 = ~n19171 & ~n19172 ;
  assign n19174 = n16558 & ~n19173 ;
  assign n19170 = ~\P2_EBX_reg[13]/NET0131  & ~n16558 ;
  assign n19175 = n1743 & ~n19170 ;
  assign n19176 = ~n19174 & n19175 ;
  assign n19178 = \P2_EBX_reg[31]/NET0131  & ~n16571 ;
  assign n19180 = ~\P2_EBX_reg[13]/NET0131  & n19178 ;
  assign n19179 = \P2_EBX_reg[13]/NET0131  & ~n19178 ;
  assign n19181 = ~n1920 & ~n19179 ;
  assign n19182 = ~n19180 & n19181 ;
  assign n19177 = n1920 & ~n19173 ;
  assign n19183 = n1742 & ~n19177 ;
  assign n19184 = ~n19182 & n19183 ;
  assign n19185 = ~n19176 & ~n19184 ;
  assign n19186 = ~n1810 & ~n19185 ;
  assign n19187 = ~n19169 & ~n19186 ;
  assign n19188 = n1927 & ~n19187 ;
  assign n19168 = \P2_rEIP_reg[13]/NET0131  & ~n18989 ;
  assign n19189 = \P2_PhyAddrPointer_reg[13]/NET0131  & n2987 ;
  assign n19190 = ~n3113 & ~n19189 ;
  assign n19191 = ~n19168 & n19190 ;
  assign n19192 = ~n19188 & n19191 ;
  assign n19193 = ~n19167 & n19192 ;
  assign n19195 = n10113 & n18929 ;
  assign n19196 = n18540 & ~n19195 ;
  assign n19197 = ~n12354 & ~n19196 ;
  assign n19198 = n12354 & n19196 ;
  assign n19199 = ~n19197 & ~n19198 ;
  assign n19200 = ~\P1_DataWidth_reg[1]/NET0131  & ~n19199 ;
  assign n19194 = \P1_DataWidth_reg[1]/NET0131  & ~\P1_rEIP_reg[26]/NET0131  ;
  assign n19201 = n2436 & ~n19194 ;
  assign n19202 = ~n19200 & n19201 ;
  assign n19209 = ~\P1_EBX_reg[24]/NET0131  & ~\P1_EBX_reg[25]/NET0131  ;
  assign n19210 = n19023 & n19209 ;
  assign n19211 = \P1_EBX_reg[31]/NET0131  & ~n19210 ;
  assign n19213 = ~\P1_EBX_reg[26]/NET0131  & n19211 ;
  assign n19212 = \P1_EBX_reg[26]/NET0131  & ~n19211 ;
  assign n19214 = ~n2425 & ~n19212 ;
  assign n19215 = ~n19213 & n19214 ;
  assign n19205 = ~\P1_rEIP_reg[26]/NET0131  & ~n19096 ;
  assign n19206 = \P1_rEIP_reg[26]/NET0131  & n19096 ;
  assign n19207 = ~n19205 & ~n19206 ;
  assign n19208 = n2425 & ~n19207 ;
  assign n19216 = n7246 & ~n19208 ;
  assign n19217 = ~n19215 & n19216 ;
  assign n19218 = \P1_rEIP_reg[26]/NET0131  & n18690 ;
  assign n19221 = ~\P1_EBX_reg[26]/NET0131  & ~n2425 ;
  assign n19222 = n2312 & ~n19221 ;
  assign n19223 = ~n19208 & n19222 ;
  assign n19219 = \P1_EBX_reg[26]/NET0131  & n18692 ;
  assign n19220 = \P1_rEIP_reg[26]/NET0131  & n2301 ;
  assign n19224 = ~n19219 & ~n19220 ;
  assign n19225 = ~n19223 & n19224 ;
  assign n19226 = n2225 & ~n19225 ;
  assign n19227 = ~n19218 & ~n19226 ;
  assign n19228 = ~n19217 & n19227 ;
  assign n19229 = n2432 & ~n19228 ;
  assign n19203 = \P1_rEIP_reg[26]/NET0131  & ~n18805 ;
  assign n19204 = \P1_PhyAddrPointer_reg[26]/NET0131  & n3028 ;
  assign n19230 = ~n19203 & ~n19204 ;
  assign n19231 = ~n19229 & n19230 ;
  assign n19232 = ~n19202 & n19231 ;
  assign n19234 = n8969 & n19126 ;
  assign n19235 = ~n9003 & ~n19234 ;
  assign n19237 = n13595 & ~n19235 ;
  assign n19236 = ~n13595 & n19235 ;
  assign n19238 = ~\P2_DataWidth_reg[1]/NET0131  & ~n19236 ;
  assign n19239 = ~n19237 & n19238 ;
  assign n19233 = \P2_DataWidth_reg[1]/NET0131  & ~\P2_rEIP_reg[14]/NET0131  ;
  assign n19240 = n1931 & ~n19233 ;
  assign n19241 = ~n19239 & n19240 ;
  assign n19243 = \P2_rEIP_reg[14]/NET0131  & ~n16555 ;
  assign n19245 = ~\P2_rEIP_reg[14]/NET0131  & ~n19172 ;
  assign n19246 = n16533 & n16534 ;
  assign n19247 = ~n19245 & ~n19246 ;
  assign n19248 = n16558 & ~n19247 ;
  assign n19244 = ~\P2_EBX_reg[14]/NET0131  & ~n16558 ;
  assign n19249 = n1743 & ~n19244 ;
  assign n19250 = ~n19248 & n19249 ;
  assign n19252 = \P2_EBX_reg[31]/NET0131  & ~n16572 ;
  assign n19254 = ~\P2_EBX_reg[14]/NET0131  & n19252 ;
  assign n19253 = \P2_EBX_reg[14]/NET0131  & ~n19252 ;
  assign n19255 = ~n1920 & ~n19253 ;
  assign n19256 = ~n19254 & n19255 ;
  assign n19251 = n1920 & ~n19247 ;
  assign n19257 = n1742 & ~n19251 ;
  assign n19258 = ~n19256 & n19257 ;
  assign n19259 = ~n19250 & ~n19258 ;
  assign n19260 = ~n1810 & ~n19259 ;
  assign n19261 = ~n19243 & ~n19260 ;
  assign n19262 = n1927 & ~n19261 ;
  assign n19242 = \P2_rEIP_reg[14]/NET0131  & ~n18989 ;
  assign n19263 = \P2_PhyAddrPointer_reg[14]/NET0131  & n2987 ;
  assign n19264 = ~n3113 & ~n19263 ;
  assign n19265 = ~n19242 & n19264 ;
  assign n19266 = ~n19262 & n19265 ;
  assign n19267 = ~n19241 & n19266 ;
  assign n19269 = n8971 & n16514 ;
  assign n19270 = ~n9003 & ~n19269 ;
  assign n19272 = ~n12387 & n19270 ;
  assign n19271 = n12387 & ~n19270 ;
  assign n19273 = ~\P2_DataWidth_reg[1]/NET0131  & ~n19271 ;
  assign n19274 = ~n19272 & n19273 ;
  assign n19268 = \P2_DataWidth_reg[1]/NET0131  & ~\P2_rEIP_reg[15]/NET0131  ;
  assign n19275 = n1931 & ~n19268 ;
  assign n19276 = ~n19274 & n19275 ;
  assign n19278 = \P2_rEIP_reg[15]/NET0131  & ~n16555 ;
  assign n19279 = ~\P2_EBX_reg[15]/NET0131  & ~n16558 ;
  assign n19280 = n1743 & ~n19279 ;
  assign n19287 = ~\P2_EBX_reg[14]/NET0131  & n16572 ;
  assign n19288 = \P2_EBX_reg[31]/NET0131  & ~n19287 ;
  assign n19290 = ~\P2_EBX_reg[15]/NET0131  & n19288 ;
  assign n19289 = \P2_EBX_reg[15]/NET0131  & ~n19288 ;
  assign n19291 = ~n1920 & ~n19289 ;
  assign n19292 = ~n19290 & n19291 ;
  assign n19293 = n1742 & ~n19292 ;
  assign n19294 = ~n19280 & ~n19293 ;
  assign n19281 = n1819 & n19280 ;
  assign n19282 = ~\P2_rEIP_reg[15]/NET0131  & ~n19246 ;
  assign n19283 = \P2_rEIP_reg[15]/NET0131  & n19246 ;
  assign n19284 = ~n19282 & ~n19283 ;
  assign n19285 = n1920 & ~n19284 ;
  assign n19286 = ~n19281 & n19285 ;
  assign n19295 = ~n1810 & ~n19286 ;
  assign n19296 = ~n19294 & n19295 ;
  assign n19297 = ~n19278 & ~n19296 ;
  assign n19298 = n1927 & ~n19297 ;
  assign n19277 = \P2_rEIP_reg[15]/NET0131  & ~n18989 ;
  assign n19299 = \P2_PhyAddrPointer_reg[15]/NET0131  & n2987 ;
  assign n19300 = ~n3113 & ~n19299 ;
  assign n19301 = ~n19277 & n19300 ;
  assign n19302 = ~n19298 & n19301 ;
  assign n19303 = ~n19276 & n19302 ;
  assign n19332 = \P1_PhyAddrPointer_reg[26]/NET0131  & n19195 ;
  assign n19333 = n18540 & ~n19332 ;
  assign n19335 = ~n11298 & n19333 ;
  assign n19334 = n11298 & ~n19333 ;
  assign n19336 = ~\P1_DataWidth_reg[1]/NET0131  & ~n19334 ;
  assign n19337 = ~n19335 & n19336 ;
  assign n19331 = \P1_DataWidth_reg[1]/NET0131  & ~\P1_rEIP_reg[27]/NET0131  ;
  assign n19338 = n2436 & ~n19331 ;
  assign n19339 = ~n19337 & n19338 ;
  assign n19319 = ~\P1_EBX_reg[26]/NET0131  & n19209 ;
  assign n19320 = n19023 & n19319 ;
  assign n19321 = \P1_EBX_reg[31]/NET0131  & ~n19320 ;
  assign n19323 = ~\P1_EBX_reg[27]/NET0131  & n19321 ;
  assign n19322 = \P1_EBX_reg[27]/NET0131  & ~n19321 ;
  assign n19324 = ~n2425 & ~n19322 ;
  assign n19325 = ~n19323 & n19324 ;
  assign n19309 = ~\P1_rEIP_reg[27]/NET0131  & ~n19206 ;
  assign n19310 = \P1_rEIP_reg[27]/NET0131  & n19206 ;
  assign n19311 = ~n19309 & ~n19310 ;
  assign n19312 = n2425 & ~n19311 ;
  assign n19326 = n7246 & ~n19312 ;
  assign n19327 = ~n19325 & n19326 ;
  assign n19306 = \P1_rEIP_reg[27]/NET0131  & n18690 ;
  assign n19313 = ~\P1_EBX_reg[27]/NET0131  & ~n2425 ;
  assign n19314 = n2312 & ~n19313 ;
  assign n19315 = ~n19312 & n19314 ;
  assign n19307 = \P1_EBX_reg[27]/NET0131  & n18692 ;
  assign n19308 = \P1_rEIP_reg[27]/NET0131  & n2301 ;
  assign n19316 = ~n19307 & ~n19308 ;
  assign n19317 = ~n19315 & n19316 ;
  assign n19318 = n2225 & ~n19317 ;
  assign n19328 = ~n19306 & ~n19318 ;
  assign n19329 = ~n19327 & n19328 ;
  assign n19330 = n2432 & ~n19329 ;
  assign n19304 = \P1_rEIP_reg[27]/NET0131  & ~n18805 ;
  assign n19305 = \P1_PhyAddrPointer_reg[27]/NET0131  & n3028 ;
  assign n19340 = ~n19304 & ~n19305 ;
  assign n19341 = ~n19330 & n19340 ;
  assign n19342 = ~n19339 & n19341 ;
  assign n19344 = n8972 & n16514 ;
  assign n19345 = ~n9003 & ~n19344 ;
  assign n19347 = ~n13628 & n19345 ;
  assign n19346 = n13628 & ~n19345 ;
  assign n19348 = ~\P2_DataWidth_reg[1]/NET0131  & ~n19346 ;
  assign n19349 = ~n19347 & n19348 ;
  assign n19343 = \P2_DataWidth_reg[1]/NET0131  & ~\P2_rEIP_reg[16]/NET0131  ;
  assign n19350 = n1931 & ~n19343 ;
  assign n19351 = ~n19349 & n19350 ;
  assign n19353 = \P2_rEIP_reg[16]/NET0131  & ~n16555 ;
  assign n19354 = ~\P2_EBX_reg[16]/NET0131  & ~n16558 ;
  assign n19355 = n1743 & ~n19354 ;
  assign n19362 = ~\P2_EBX_reg[15]/NET0131  & n19287 ;
  assign n19363 = \P2_EBX_reg[31]/NET0131  & ~n19362 ;
  assign n19365 = ~\P2_EBX_reg[16]/NET0131  & n19363 ;
  assign n19364 = \P2_EBX_reg[16]/NET0131  & ~n19363 ;
  assign n19366 = ~n1920 & ~n19364 ;
  assign n19367 = ~n19365 & n19366 ;
  assign n19368 = n1742 & ~n19367 ;
  assign n19369 = ~n19355 & ~n19368 ;
  assign n19356 = n1819 & n19355 ;
  assign n19357 = ~\P2_rEIP_reg[16]/NET0131  & ~n19283 ;
  assign n19358 = n16533 & n16536 ;
  assign n19359 = ~n19357 & ~n19358 ;
  assign n19360 = n1920 & ~n19359 ;
  assign n19361 = ~n19356 & n19360 ;
  assign n19370 = ~n1810 & ~n19361 ;
  assign n19371 = ~n19369 & n19370 ;
  assign n19372 = ~n19353 & ~n19371 ;
  assign n19373 = n1927 & ~n19372 ;
  assign n19352 = \P2_rEIP_reg[16]/NET0131  & ~n18989 ;
  assign n19374 = \P2_PhyAddrPointer_reg[16]/NET0131  & n2987 ;
  assign n19375 = ~n3113 & ~n19374 ;
  assign n19376 = ~n19352 & n19375 ;
  assign n19377 = ~n19373 & n19376 ;
  assign n19378 = ~n19351 & n19377 ;
  assign n19380 = \P2_PhyAddrPointer_reg[16]/NET0131  & n19344 ;
  assign n19381 = ~n9003 & ~n19380 ;
  assign n19383 = ~n13665 & n19381 ;
  assign n19382 = n13665 & ~n19381 ;
  assign n19384 = ~\P2_DataWidth_reg[1]/NET0131  & ~n19382 ;
  assign n19385 = ~n19383 & n19384 ;
  assign n19379 = \P2_DataWidth_reg[1]/NET0131  & ~\P2_rEIP_reg[17]/NET0131  ;
  assign n19386 = n1931 & ~n19379 ;
  assign n19387 = ~n19385 & n19386 ;
  assign n19389 = ~n1742 & ~n1745 ;
  assign n19390 = ~n1747 & n19389 ;
  assign n19391 = ~n16555 & ~n19390 ;
  assign n19393 = ~\P2_rEIP_reg[17]/NET0131  & ~n19358 ;
  assign n19394 = n16533 & n16537 ;
  assign n19395 = ~n19393 & ~n19394 ;
  assign n19396 = ~\P2_DataWidth_reg[1]/NET0131  & n19395 ;
  assign n19397 = n1820 & n19396 ;
  assign n19392 = \P2_EBX_reg[17]/NET0131  & ~n16558 ;
  assign n19398 = ~n1810 & ~n19392 ;
  assign n19399 = ~n19397 & n19398 ;
  assign n19400 = n1743 & ~n19399 ;
  assign n19401 = ~n19391 & ~n19400 ;
  assign n19402 = \P2_rEIP_reg[17]/NET0131  & ~n19401 ;
  assign n19403 = ~\P2_EBX_reg[16]/NET0131  & n19362 ;
  assign n19404 = \P2_EBX_reg[31]/NET0131  & ~n19403 ;
  assign n19406 = \P2_EBX_reg[17]/NET0131  & n19404 ;
  assign n19405 = ~\P2_EBX_reg[17]/NET0131  & ~n19404 ;
  assign n19407 = ~n1920 & ~n19405 ;
  assign n19408 = ~n19406 & n19407 ;
  assign n19409 = ~n1805 & n19396 ;
  assign n19410 = ~n19408 & ~n19409 ;
  assign n19411 = n1742 & ~n19410 ;
  assign n19412 = ~n19400 & ~n19411 ;
  assign n19413 = ~n1810 & ~n19412 ;
  assign n19414 = ~n19402 & ~n19413 ;
  assign n19415 = n1927 & ~n19414 ;
  assign n19388 = \P2_rEIP_reg[17]/NET0131  & ~n18989 ;
  assign n19416 = \P2_PhyAddrPointer_reg[17]/NET0131  & n2987 ;
  assign n19417 = ~n3113 & ~n19416 ;
  assign n19418 = ~n19388 & n19417 ;
  assign n19419 = ~n19415 & n19418 ;
  assign n19420 = ~n19387 & n19419 ;
  assign n19442 = n11292 & n19195 ;
  assign n19443 = n18540 & ~n19442 ;
  assign n19445 = ~n11340 & n19443 ;
  assign n19444 = n11340 & ~n19443 ;
  assign n19446 = ~\P1_DataWidth_reg[1]/NET0131  & ~n19444 ;
  assign n19447 = ~n19445 & n19446 ;
  assign n19441 = \P1_DataWidth_reg[1]/NET0131  & ~\P1_rEIP_reg[28]/NET0131  ;
  assign n19448 = n2436 & ~n19441 ;
  assign n19449 = ~n19447 & n19448 ;
  assign n19430 = ~\P1_EBX_reg[27]/NET0131  & n19320 ;
  assign n19431 = \P1_EBX_reg[31]/NET0131  & ~n19430 ;
  assign n19433 = ~\P1_EBX_reg[28]/NET0131  & n19431 ;
  assign n19432 = \P1_EBX_reg[28]/NET0131  & ~n19431 ;
  assign n19434 = ~n2425 & ~n19432 ;
  assign n19435 = ~n19433 & n19434 ;
  assign n19423 = ~\P1_rEIP_reg[28]/NET0131  & ~n19310 ;
  assign n19424 = \P1_rEIP_reg[28]/NET0131  & n19310 ;
  assign n19425 = ~n19423 & ~n19424 ;
  assign n19426 = n2425 & ~n19425 ;
  assign n19436 = n7246 & ~n19426 ;
  assign n19437 = ~n19435 & n19436 ;
  assign n19421 = \P1_rEIP_reg[28]/NET0131  & ~n18554 ;
  assign n19427 = ~n2311 & n19426 ;
  assign n19422 = ~\P1_EBX_reg[28]/NET0131  & ~n18556 ;
  assign n19428 = n15990 & ~n19422 ;
  assign n19429 = ~n19427 & n19428 ;
  assign n19438 = ~n19421 & ~n19429 ;
  assign n19439 = ~n19437 & n19438 ;
  assign n19440 = n2432 & ~n19439 ;
  assign n19450 = \P1_PhyAddrPointer_reg[28]/NET0131  & n3028 ;
  assign n19451 = \P1_rEIP_reg[28]/NET0131  & ~n18805 ;
  assign n19452 = ~n19450 & ~n19451 ;
  assign n19453 = ~n19440 & n19452 ;
  assign n19454 = ~n19449 & n19453 ;
  assign n19456 = ~n9003 & ~n16515 ;
  assign n19458 = ~n13674 & n19456 ;
  assign n19457 = n13674 & ~n19456 ;
  assign n19459 = ~\P2_DataWidth_reg[1]/NET0131  & ~n19457 ;
  assign n19460 = ~n19458 & n19459 ;
  assign n19455 = \P2_DataWidth_reg[1]/NET0131  & ~\P2_rEIP_reg[18]/NET0131  ;
  assign n19461 = n1931 & ~n19455 ;
  assign n19462 = ~n19460 & n19461 ;
  assign n19464 = \P2_rEIP_reg[18]/NET0131  & ~n16555 ;
  assign n19467 = ~\P2_EBX_reg[18]/NET0131  & ~n16558 ;
  assign n19468 = n1743 & ~n19467 ;
  assign n19472 = \P2_EBX_reg[31]/NET0131  & ~n16576 ;
  assign n19474 = ~\P2_EBX_reg[18]/NET0131  & n19472 ;
  assign n19473 = \P2_EBX_reg[18]/NET0131  & ~n19472 ;
  assign n19475 = ~n1920 & ~n19473 ;
  assign n19476 = ~n19474 & n19475 ;
  assign n19477 = n1742 & ~n19476 ;
  assign n19478 = ~n19468 & ~n19477 ;
  assign n19469 = n1819 & n19468 ;
  assign n19465 = ~\P2_rEIP_reg[18]/NET0131  & ~n19394 ;
  assign n19466 = ~n16539 & ~n19465 ;
  assign n19470 = n1920 & ~n19466 ;
  assign n19471 = ~n19469 & n19470 ;
  assign n19479 = ~n1810 & ~n19471 ;
  assign n19480 = ~n19478 & n19479 ;
  assign n19481 = ~n19464 & ~n19480 ;
  assign n19482 = n1927 & ~n19481 ;
  assign n19463 = \P2_rEIP_reg[18]/NET0131  & ~n18989 ;
  assign n19483 = \P2_PhyAddrPointer_reg[18]/NET0131  & n2987 ;
  assign n19484 = ~n3113 & ~n19483 ;
  assign n19485 = ~n19463 & n19484 ;
  assign n19486 = ~n19482 & n19485 ;
  assign n19487 = ~n19462 & n19486 ;
  assign n19489 = ~n8975 & ~n9003 ;
  assign n19490 = ~n19456 & ~n19489 ;
  assign n19492 = ~n12429 & ~n19490 ;
  assign n19491 = n12429 & n19490 ;
  assign n19493 = ~\P2_DataWidth_reg[1]/NET0131  & ~n19491 ;
  assign n19494 = ~n19492 & n19493 ;
  assign n19488 = \P2_DataWidth_reg[1]/NET0131  & ~\P2_rEIP_reg[19]/NET0131  ;
  assign n19495 = n1931 & ~n19488 ;
  assign n19496 = ~n19494 & n19495 ;
  assign n19498 = \P2_rEIP_reg[19]/NET0131  & ~n16555 ;
  assign n19500 = ~\P2_rEIP_reg[19]/NET0131  & ~n16539 ;
  assign n19501 = ~n16540 & ~n19500 ;
  assign n19502 = n16558 & ~n19501 ;
  assign n19499 = ~\P2_EBX_reg[19]/NET0131  & ~n16558 ;
  assign n19503 = n1743 & ~n19499 ;
  assign n19504 = ~n19502 & n19503 ;
  assign n19506 = ~\P2_EBX_reg[18]/NET0131  & n16576 ;
  assign n19507 = \P2_EBX_reg[31]/NET0131  & ~n19506 ;
  assign n19509 = ~\P2_EBX_reg[19]/NET0131  & n19507 ;
  assign n19508 = \P2_EBX_reg[19]/NET0131  & ~n19507 ;
  assign n19510 = ~n1920 & ~n19508 ;
  assign n19511 = ~n19509 & n19510 ;
  assign n19505 = n1920 & ~n19501 ;
  assign n19512 = n1742 & ~n19505 ;
  assign n19513 = ~n19511 & n19512 ;
  assign n19514 = ~n19504 & ~n19513 ;
  assign n19515 = ~n1810 & ~n19514 ;
  assign n19516 = ~n19498 & ~n19515 ;
  assign n19517 = n1927 & ~n19516 ;
  assign n19497 = \P2_rEIP_reg[19]/NET0131  & ~n18989 ;
  assign n19518 = \P2_PhyAddrPointer_reg[19]/NET0131  & n2987 ;
  assign n19519 = ~n3113 & ~n19518 ;
  assign n19520 = ~n19497 & n19519 ;
  assign n19521 = ~n19517 & n19520 ;
  assign n19522 = ~n19496 & n19521 ;
  assign n19536 = ~\P1_EBX_reg[27]/NET0131  & ~\P1_EBX_reg[28]/NET0131  ;
  assign n19537 = n19320 & n19536 ;
  assign n19538 = \P1_EBX_reg[31]/NET0131  & ~n19537 ;
  assign n19540 = ~\P1_EBX_reg[29]/NET0131  & n19538 ;
  assign n19539 = \P1_EBX_reg[29]/NET0131  & ~n19538 ;
  assign n19541 = ~n2425 & ~n19539 ;
  assign n19542 = ~n19540 & n19541 ;
  assign n19523 = ~\P1_rEIP_reg[29]/NET0131  & ~n19424 ;
  assign n19524 = \P1_rEIP_reg[29]/NET0131  & n19424 ;
  assign n19525 = ~n19523 & ~n19524 ;
  assign n19526 = n2425 & ~n19525 ;
  assign n19543 = n7246 & ~n19526 ;
  assign n19544 = ~n19542 & n19543 ;
  assign n19527 = ~\P1_EBX_reg[29]/NET0131  & ~n2425 ;
  assign n19528 = n2312 & ~n19527 ;
  assign n19529 = ~n19526 & n19528 ;
  assign n19530 = \P1_EBX_reg[29]/NET0131  & n18692 ;
  assign n19531 = \P1_rEIP_reg[29]/NET0131  & n2301 ;
  assign n19532 = ~n19530 & ~n19531 ;
  assign n19533 = ~n19529 & n19532 ;
  assign n19534 = n2225 & ~n19533 ;
  assign n19535 = \P1_rEIP_reg[29]/NET0131  & n18690 ;
  assign n19545 = ~n19534 & ~n19535 ;
  assign n19546 = ~n19544 & n19545 ;
  assign n19547 = n2432 & ~n19546 ;
  assign n19549 = \P1_PhyAddrPointer_reg[28]/NET0131  & n19442 ;
  assign n19550 = n18540 & ~n19549 ;
  assign n19552 = ~n11361 & n19550 ;
  assign n19551 = n11361 & ~n19550 ;
  assign n19553 = ~\P1_DataWidth_reg[1]/NET0131  & ~n19551 ;
  assign n19554 = ~n19552 & n19553 ;
  assign n19548 = \P1_DataWidth_reg[1]/NET0131  & ~\P1_rEIP_reg[29]/NET0131  ;
  assign n19555 = n2436 & ~n19548 ;
  assign n19556 = ~n19554 & n19555 ;
  assign n19557 = \P1_PhyAddrPointer_reg[29]/NET0131  & n3028 ;
  assign n19558 = \P1_rEIP_reg[29]/NET0131  & ~n18805 ;
  assign n19559 = ~n19557 & ~n19558 ;
  assign n19560 = ~n19556 & n19559 ;
  assign n19561 = ~n19547 & n19560 ;
  assign n19563 = \P2_PhyAddrPointer_reg[0]/NET0131  & ~n9003 ;
  assign n19565 = \P2_PhyAddrPointer_reg[1]/NET0131  & n19563 ;
  assign n19564 = ~\P2_PhyAddrPointer_reg[1]/NET0131  & ~n19563 ;
  assign n19566 = ~\P2_DataWidth_reg[1]/NET0131  & ~n19564 ;
  assign n19567 = ~n19565 & n19566 ;
  assign n19562 = \P2_DataWidth_reg[1]/NET0131  & ~\P2_rEIP_reg[1]/NET0131  ;
  assign n19568 = n1931 & ~n19562 ;
  assign n19569 = ~n19567 & n19568 ;
  assign n19572 = \P2_rEIP_reg[1]/NET0131  & ~n16555 ;
  assign n19580 = ~n15022 & ~n16560 ;
  assign n19581 = \P2_EBX_reg[31]/NET0131  & ~n19580 ;
  assign n19579 = ~\P2_EBX_reg[1]/NET0131  & ~\P2_EBX_reg[31]/NET0131  ;
  assign n19582 = ~n1920 & ~n19579 ;
  assign n19583 = ~n19581 & n19582 ;
  assign n19574 = ~\P2_DataWidth_reg[1]/NET0131  & ~\P2_rEIP_reg[1]/NET0131  ;
  assign n19584 = ~n1805 & n19574 ;
  assign n19585 = ~n19583 & ~n19584 ;
  assign n19586 = n1742 & ~n19585 ;
  assign n19573 = \P2_EBX_reg[1]/NET0131  & ~n16558 ;
  assign n19575 = n1820 & n19574 ;
  assign n19576 = ~n19573 & ~n19575 ;
  assign n19577 = n1743 & ~n19576 ;
  assign n19578 = n1745 & ~n1872 ;
  assign n19587 = ~n19577 & ~n19578 ;
  assign n19588 = ~n19586 & n19587 ;
  assign n19589 = ~n1810 & ~n19588 ;
  assign n19590 = ~n19572 & ~n19589 ;
  assign n19591 = n1927 & ~n19590 ;
  assign n19570 = \P2_PhyAddrPointer_reg[1]/NET0131  & n2987 ;
  assign n19571 = \P2_rEIP_reg[1]/NET0131  & ~n16511 ;
  assign n19592 = ~n19570 & ~n19571 ;
  assign n19593 = ~n19591 & n19592 ;
  assign n19594 = ~n19569 & n19593 ;
  assign n19596 = n8976 & n16515 ;
  assign n19597 = ~n9003 & ~n19596 ;
  assign n19599 = ~n11877 & n19597 ;
  assign n19598 = n11877 & ~n19597 ;
  assign n19600 = ~\P2_DataWidth_reg[1]/NET0131  & ~n19598 ;
  assign n19601 = ~n19599 & n19600 ;
  assign n19595 = \P2_DataWidth_reg[1]/NET0131  & ~\P2_rEIP_reg[20]/NET0131  ;
  assign n19602 = n1931 & ~n19595 ;
  assign n19603 = ~n19601 & n19602 ;
  assign n19606 = ~\P2_rEIP_reg[20]/NET0131  & ~n16540 ;
  assign n19607 = ~\P2_DataWidth_reg[1]/NET0131  & ~n16541 ;
  assign n19608 = ~n19606 & n19607 ;
  assign n19609 = n1820 & n19608 ;
  assign n19605 = \P2_EBX_reg[20]/NET0131  & ~n16558 ;
  assign n19610 = ~n1810 & ~n19605 ;
  assign n19611 = ~n19609 & n19610 ;
  assign n19612 = n1743 & ~n19611 ;
  assign n19613 = ~n19391 & ~n19612 ;
  assign n19614 = \P2_rEIP_reg[20]/NET0131  & ~n19613 ;
  assign n19615 = \P2_EBX_reg[31]/NET0131  & ~n16578 ;
  assign n19617 = \P2_EBX_reg[20]/NET0131  & n19615 ;
  assign n19616 = ~\P2_EBX_reg[20]/NET0131  & ~n19615 ;
  assign n19618 = ~n1920 & ~n19616 ;
  assign n19619 = ~n19617 & n19618 ;
  assign n19620 = ~n1805 & n19608 ;
  assign n19621 = ~n19619 & ~n19620 ;
  assign n19622 = n1742 & ~n19621 ;
  assign n19623 = ~n19612 & ~n19622 ;
  assign n19624 = ~n1810 & ~n19623 ;
  assign n19625 = ~n19614 & ~n19624 ;
  assign n19626 = n1927 & ~n19625 ;
  assign n19604 = \P2_rEIP_reg[20]/NET0131  & ~n16511 ;
  assign n19627 = \P2_PhyAddrPointer_reg[20]/NET0131  & n2987 ;
  assign n19628 = ~n19604 & ~n19627 ;
  assign n19629 = ~n19626 & n19628 ;
  assign n19630 = ~n19603 & n19629 ;
  assign n19632 = n8977 & n16515 ;
  assign n19633 = ~n9003 & ~n19632 ;
  assign n19635 = ~n12968 & n19633 ;
  assign n19634 = n12968 & ~n19633 ;
  assign n19636 = ~\P2_DataWidth_reg[1]/NET0131  & ~n19634 ;
  assign n19637 = ~n19635 & n19636 ;
  assign n19631 = \P2_DataWidth_reg[1]/NET0131  & ~\P2_rEIP_reg[21]/NET0131  ;
  assign n19638 = n1931 & ~n19631 ;
  assign n19639 = ~n19637 & n19638 ;
  assign n19641 = \P2_rEIP_reg[21]/NET0131  & ~n16555 ;
  assign n19642 = ~\P2_EBX_reg[21]/NET0131  & ~n16558 ;
  assign n19643 = n15980 & ~n19642 ;
  assign n19644 = \P2_EBX_reg[31]/NET0131  & ~n16579 ;
  assign n19646 = ~\P2_EBX_reg[21]/NET0131  & n19644 ;
  assign n19645 = \P2_EBX_reg[21]/NET0131  & ~n19644 ;
  assign n19647 = ~n1920 & ~n19645 ;
  assign n19648 = ~n19646 & n19647 ;
  assign n19649 = n10236 & ~n19648 ;
  assign n19650 = ~n19643 & ~n19649 ;
  assign n19653 = n1819 & n15980 ;
  assign n19654 = ~n19642 & n19653 ;
  assign n19651 = ~\P2_rEIP_reg[21]/NET0131  & ~n16541 ;
  assign n19652 = ~n16542 & ~n19651 ;
  assign n19655 = n1920 & ~n19652 ;
  assign n19656 = ~n19654 & n19655 ;
  assign n19657 = ~n19650 & ~n19656 ;
  assign n19658 = ~n19641 & ~n19657 ;
  assign n19659 = n1927 & ~n19658 ;
  assign n19640 = \P2_PhyAddrPointer_reg[21]/NET0131  & n2987 ;
  assign n19660 = \P2_rEIP_reg[21]/NET0131  & ~n16511 ;
  assign n19661 = ~n19640 & ~n19660 ;
  assign n19662 = ~n19659 & n19661 ;
  assign n19663 = ~n19639 & n19662 ;
  assign n19665 = n18540 & ~n18541 ;
  assign n19666 = ~\P1_PhyAddrPointer_reg[1]/NET0131  & ~\P1_PhyAddrPointer_reg[2]/NET0131  ;
  assign n19667 = ~n15825 & ~n19666 ;
  assign n19668 = ~n19665 & ~n19667 ;
  assign n19669 = n19665 & n19667 ;
  assign n19670 = ~n19668 & ~n19669 ;
  assign n19671 = ~\P1_DataWidth_reg[1]/NET0131  & ~n19670 ;
  assign n19664 = \P1_DataWidth_reg[1]/NET0131  & ~\P1_rEIP_reg[2]/NET0131  ;
  assign n19672 = n2436 & ~n19664 ;
  assign n19673 = ~n19671 & n19672 ;
  assign n19677 = \P1_rEIP_reg[2]/NET0131  & ~n18554 ;
  assign n19679 = ~\P1_rEIP_reg[1]/NET0131  & ~\P1_rEIP_reg[2]/NET0131  ;
  assign n19680 = ~\P1_DataWidth_reg[1]/NET0131  & ~n18558 ;
  assign n19681 = ~n19679 & n19680 ;
  assign n19685 = ~n2317 & n19681 ;
  assign n19686 = \P1_EBX_reg[31]/NET0131  & ~n18577 ;
  assign n19688 = \P1_EBX_reg[2]/NET0131  & n19686 ;
  assign n19687 = ~\P1_EBX_reg[2]/NET0131  & ~n19686 ;
  assign n19689 = ~n2425 & ~n19687 ;
  assign n19690 = ~n19688 & n19689 ;
  assign n19691 = ~n19685 & ~n19690 ;
  assign n19692 = n7246 & ~n19691 ;
  assign n19676 = n2274 & n18807 ;
  assign n19678 = \P1_EBX_reg[2]/NET0131  & ~n18556 ;
  assign n19682 = n2387 & n19681 ;
  assign n19683 = ~n19678 & ~n19682 ;
  assign n19684 = n15990 & ~n19683 ;
  assign n19693 = ~n19676 & ~n19684 ;
  assign n19694 = ~n19692 & n19693 ;
  assign n19695 = ~n19677 & n19694 ;
  assign n19696 = n2432 & ~n19695 ;
  assign n19674 = \P1_PhyAddrPointer_reg[2]/NET0131  & n3028 ;
  assign n19675 = \P1_rEIP_reg[2]/NET0131  & ~n18805 ;
  assign n19697 = ~n19674 & ~n19675 ;
  assign n19698 = ~n19696 & n19697 ;
  assign n19699 = ~n19673 & n19698 ;
  assign n19701 = \P2_PhyAddrPointer_reg[21]/NET0131  & n19632 ;
  assign n19702 = ~n9003 & ~n19701 ;
  assign n19704 = n11898 & ~n19702 ;
  assign n19703 = ~n11898 & n19702 ;
  assign n19705 = ~\P2_DataWidth_reg[1]/NET0131  & ~n19703 ;
  assign n19706 = ~n19704 & n19705 ;
  assign n19700 = \P2_DataWidth_reg[1]/NET0131  & ~\P2_rEIP_reg[22]/NET0131  ;
  assign n19707 = n1931 & ~n19700 ;
  assign n19708 = ~n19706 & n19707 ;
  assign n19710 = \P2_rEIP_reg[22]/NET0131  & ~n16555 ;
  assign n19713 = ~\P2_EBX_reg[22]/NET0131  & ~n16558 ;
  assign n19714 = n1743 & ~n19713 ;
  assign n19718 = \P2_EBX_reg[31]/NET0131  & ~n16580 ;
  assign n19720 = ~\P2_EBX_reg[22]/NET0131  & n19718 ;
  assign n19719 = \P2_EBX_reg[22]/NET0131  & ~n19718 ;
  assign n19721 = ~n1920 & ~n19719 ;
  assign n19722 = ~n19720 & n19721 ;
  assign n19723 = n1742 & ~n19722 ;
  assign n19724 = ~n19714 & ~n19723 ;
  assign n19711 = ~\P2_rEIP_reg[22]/NET0131  & ~n16542 ;
  assign n19712 = ~n16543 & ~n19711 ;
  assign n19715 = n1819 & n19714 ;
  assign n19716 = n1920 & ~n19715 ;
  assign n19717 = ~n19712 & n19716 ;
  assign n19725 = ~n1810 & ~n19717 ;
  assign n19726 = ~n19724 & n19725 ;
  assign n19727 = ~n19710 & ~n19726 ;
  assign n19728 = n1927 & ~n19727 ;
  assign n19709 = \P2_PhyAddrPointer_reg[22]/NET0131  & n2987 ;
  assign n19729 = \P2_rEIP_reg[22]/NET0131  & ~n16511 ;
  assign n19730 = ~n19709 & ~n19729 ;
  assign n19731 = ~n19728 & n19730 ;
  assign n19732 = ~n19708 & n19731 ;
  assign n19734 = n8978 & n19632 ;
  assign n19735 = ~n9003 & ~n19734 ;
  assign n19737 = ~n10962 & n19735 ;
  assign n19736 = n10962 & ~n19735 ;
  assign n19738 = ~\P2_DataWidth_reg[1]/NET0131  & ~n19736 ;
  assign n19739 = ~n19737 & n19738 ;
  assign n19733 = \P2_DataWidth_reg[1]/NET0131  & ~\P2_rEIP_reg[23]/NET0131  ;
  assign n19740 = n1931 & ~n19733 ;
  assign n19741 = ~n19739 & n19740 ;
  assign n19743 = \P2_rEIP_reg[23]/NET0131  & ~n16555 ;
  assign n19744 = ~\P2_EBX_reg[23]/NET0131  & ~n16558 ;
  assign n19745 = n15980 & ~n19744 ;
  assign n19746 = ~\P2_EBX_reg[22]/NET0131  & n16580 ;
  assign n19747 = \P2_EBX_reg[31]/NET0131  & ~n19746 ;
  assign n19749 = \P2_EBX_reg[23]/NET0131  & ~n19747 ;
  assign n19748 = ~\P2_EBX_reg[23]/NET0131  & n19747 ;
  assign n19750 = ~n1920 & ~n19748 ;
  assign n19751 = ~n19749 & n19750 ;
  assign n19752 = n10236 & ~n19751 ;
  assign n19753 = ~n19745 & ~n19752 ;
  assign n19755 = ~\P2_rEIP_reg[23]/NET0131  & ~n16543 ;
  assign n19756 = ~n16544 & ~n19755 ;
  assign n19754 = \P2_EBX_reg[23]/NET0131  & n19653 ;
  assign n19757 = n1920 & ~n19754 ;
  assign n19758 = ~n19756 & n19757 ;
  assign n19759 = ~n19753 & ~n19758 ;
  assign n19760 = ~n19743 & ~n19759 ;
  assign n19761 = n1927 & ~n19760 ;
  assign n19742 = \P2_rEIP_reg[23]/NET0131  & ~n16511 ;
  assign n19762 = \P2_PhyAddrPointer_reg[23]/NET0131  & n2987 ;
  assign n19763 = ~n19742 & ~n19762 ;
  assign n19764 = ~n19761 & n19763 ;
  assign n19765 = ~n19741 & n19764 ;
  assign n19767 = ~\P2_PhyAddrPointer_reg[23]/NET0131  & ~n9003 ;
  assign n19768 = ~n19735 & ~n19767 ;
  assign n19770 = n11934 & n19768 ;
  assign n19769 = ~n11934 & ~n19768 ;
  assign n19771 = ~\P2_DataWidth_reg[1]/NET0131  & ~n19769 ;
  assign n19772 = ~n19770 & n19771 ;
  assign n19766 = \P2_DataWidth_reg[1]/NET0131  & ~\P2_rEIP_reg[24]/NET0131  ;
  assign n19773 = n1931 & ~n19766 ;
  assign n19774 = ~n19772 & n19773 ;
  assign n19776 = \P2_rEIP_reg[24]/NET0131  & ~n16555 ;
  assign n19777 = \P2_EBX_reg[31]/NET0131  & ~n16582 ;
  assign n19780 = ~n15980 & n19777 ;
  assign n19781 = \P2_EBX_reg[24]/NET0131  & ~n15981 ;
  assign n19782 = ~n19780 & n19781 ;
  assign n19778 = ~\P2_EBX_reg[24]/NET0131  & n10236 ;
  assign n19779 = n19777 & n19778 ;
  assign n19783 = ~n16553 & ~n19779 ;
  assign n19784 = ~n19782 & n19783 ;
  assign n19786 = ~\P2_rEIP_reg[24]/NET0131  & ~n16544 ;
  assign n19787 = ~n16545 & ~n19786 ;
  assign n19785 = \P2_EBX_reg[24]/NET0131  & n19653 ;
  assign n19788 = n1920 & ~n19785 ;
  assign n19789 = ~n19787 & n19788 ;
  assign n19790 = ~n19784 & ~n19789 ;
  assign n19791 = ~n19776 & ~n19790 ;
  assign n19792 = n1927 & ~n19791 ;
  assign n19775 = \P2_PhyAddrPointer_reg[24]/NET0131  & n2987 ;
  assign n19793 = \P2_rEIP_reg[24]/NET0131  & ~n16511 ;
  assign n19794 = ~n19775 & ~n19793 ;
  assign n19795 = ~n19792 & n19794 ;
  assign n19796 = ~n19774 & n19795 ;
  assign n19817 = ~n9003 & ~n16516 ;
  assign n19819 = ~n13011 & n19817 ;
  assign n19818 = n13011 & ~n19817 ;
  assign n19820 = ~\P2_DataWidth_reg[1]/NET0131  & ~n19818 ;
  assign n19821 = ~n19819 & n19820 ;
  assign n19816 = \P2_DataWidth_reg[1]/NET0131  & ~\P2_rEIP_reg[25]/NET0131  ;
  assign n19822 = n1931 & ~n19816 ;
  assign n19823 = ~n19821 & n19822 ;
  assign n19797 = \P2_rEIP_reg[25]/NET0131  & ~n16555 ;
  assign n19798 = ~\P2_EBX_reg[25]/NET0131  & ~n16558 ;
  assign n19799 = n15980 & ~n19798 ;
  assign n19800 = ~\P2_EBX_reg[24]/NET0131  & n16582 ;
  assign n19801 = \P2_EBX_reg[31]/NET0131  & ~n19800 ;
  assign n19803 = \P2_EBX_reg[25]/NET0131  & ~n19801 ;
  assign n19802 = ~\P2_EBX_reg[25]/NET0131  & n19801 ;
  assign n19804 = ~n1920 & ~n19802 ;
  assign n19805 = ~n19803 & n19804 ;
  assign n19806 = n10236 & ~n19805 ;
  assign n19807 = ~n19799 & ~n19806 ;
  assign n19809 = ~\P2_rEIP_reg[25]/NET0131  & ~n16545 ;
  assign n19810 = ~n16546 & ~n19809 ;
  assign n19808 = \P2_EBX_reg[25]/NET0131  & n19653 ;
  assign n19811 = n1920 & ~n19808 ;
  assign n19812 = ~n19810 & n19811 ;
  assign n19813 = ~n19807 & ~n19812 ;
  assign n19814 = ~n19797 & ~n19813 ;
  assign n19815 = n1927 & ~n19814 ;
  assign n19824 = \P2_rEIP_reg[25]/NET0131  & ~n16511 ;
  assign n19825 = \P2_PhyAddrPointer_reg[25]/NET0131  & n2987 ;
  assign n19826 = ~n19824 & ~n19825 ;
  assign n19827 = ~n19815 & n19826 ;
  assign n19828 = ~n19823 & n19827 ;
  assign n19830 = ~\P1_PhyAddrPointer_reg[0]/NET0131  & n15825 ;
  assign n19831 = n18540 & ~n19830 ;
  assign n19833 = n16263 & ~n19831 ;
  assign n19832 = ~n16263 & n19831 ;
  assign n19834 = ~\P1_DataWidth_reg[1]/NET0131  & ~n19832 ;
  assign n19835 = ~n19833 & n19834 ;
  assign n19829 = \P1_DataWidth_reg[1]/NET0131  & ~\P1_rEIP_reg[3]/NET0131  ;
  assign n19836 = n2436 & ~n19829 ;
  assign n19837 = ~n19835 & n19836 ;
  assign n19839 = \P1_rEIP_reg[3]/NET0131  & ~n18554 ;
  assign n19852 = \P1_EBX_reg[3]/NET0131  & ~n18556 ;
  assign n19845 = ~\P1_rEIP_reg[3]/NET0131  & ~n18558 ;
  assign n19846 = ~\P1_DataWidth_reg[1]/NET0131  & ~n18559 ;
  assign n19847 = ~n19845 & n19846 ;
  assign n19853 = n2387 & n19847 ;
  assign n19854 = ~n19852 & ~n19853 ;
  assign n19855 = n2225 & ~n19854 ;
  assign n19840 = \P1_EBX_reg[31]/NET0131  & ~n18578 ;
  assign n19842 = \P1_EBX_reg[3]/NET0131  & n19840 ;
  assign n19841 = ~\P1_EBX_reg[3]/NET0131  & ~n19840 ;
  assign n19843 = ~n2425 & ~n19841 ;
  assign n19844 = ~n19842 & n19843 ;
  assign n19848 = ~n2317 & n19847 ;
  assign n19849 = ~n19844 & ~n19848 ;
  assign n19850 = n2222 & ~n19849 ;
  assign n19851 = n2231 & ~n2348 ;
  assign n19856 = ~n19850 & ~n19851 ;
  assign n19857 = ~n19855 & n19856 ;
  assign n19858 = ~n2301 & ~n19857 ;
  assign n19859 = ~n19839 & ~n19858 ;
  assign n19860 = n2432 & ~n19859 ;
  assign n19838 = \P1_rEIP_reg[3]/NET0131  & ~n18805 ;
  assign n19861 = ~n16265 & ~n19838 ;
  assign n19862 = ~n19860 & n19861 ;
  assign n19863 = ~n19837 & n19862 ;
  assign n19885 = ~n9003 & ~n16517 ;
  assign n19886 = ~n11953 & ~n19885 ;
  assign n19887 = n11953 & n19885 ;
  assign n19888 = ~n19886 & ~n19887 ;
  assign n19889 = ~\P2_DataWidth_reg[1]/NET0131  & ~n19888 ;
  assign n19884 = \P2_DataWidth_reg[1]/NET0131  & ~\P2_rEIP_reg[26]/NET0131  ;
  assign n19890 = n1931 & ~n19884 ;
  assign n19891 = ~n19889 & n19890 ;
  assign n19864 = \P2_rEIP_reg[26]/NET0131  & ~n16555 ;
  assign n19865 = ~\P2_EBX_reg[26]/NET0131  & ~n16558 ;
  assign n19866 = n15980 & ~n19865 ;
  assign n19867 = \P2_EBX_reg[31]/NET0131  & ~n16584 ;
  assign n19869 = ~\P2_EBX_reg[26]/NET0131  & n19867 ;
  assign n19868 = \P2_EBX_reg[26]/NET0131  & ~n19867 ;
  assign n19870 = ~n1920 & ~n19868 ;
  assign n19871 = ~n19869 & n19870 ;
  assign n19872 = n10236 & ~n19871 ;
  assign n19873 = ~n19866 & ~n19872 ;
  assign n19875 = ~\P2_rEIP_reg[26]/NET0131  & ~n16546 ;
  assign n19876 = ~n16547 & ~n19875 ;
  assign n19874 = \P2_EBX_reg[26]/NET0131  & n19653 ;
  assign n19877 = n1920 & ~n19874 ;
  assign n19878 = ~n19876 & n19877 ;
  assign n19879 = ~n19873 & ~n19878 ;
  assign n19880 = ~n19864 & ~n19879 ;
  assign n19881 = n1927 & ~n19880 ;
  assign n19882 = \P2_rEIP_reg[26]/NET0131  & ~n16511 ;
  assign n19883 = \P2_PhyAddrPointer_reg[26]/NET0131  & n2987 ;
  assign n19892 = ~n19882 & ~n19883 ;
  assign n19893 = ~n19881 & n19892 ;
  assign n19894 = ~n19891 & n19893 ;
  assign n19896 = ~n8983 & ~n9003 ;
  assign n19897 = ~n19456 & ~n19896 ;
  assign n19899 = ~n11005 & ~n19897 ;
  assign n19898 = n11005 & n19897 ;
  assign n19900 = ~\P2_DataWidth_reg[1]/NET0131  & ~n19898 ;
  assign n19901 = ~n19899 & n19900 ;
  assign n19895 = \P2_DataWidth_reg[1]/NET0131  & ~\P2_rEIP_reg[27]/NET0131  ;
  assign n19902 = n1931 & ~n19895 ;
  assign n19903 = ~n19901 & n19902 ;
  assign n19912 = \P2_EBX_reg[31]/NET0131  & ~n16585 ;
  assign n19914 = ~\P2_EBX_reg[27]/NET0131  & n19912 ;
  assign n19913 = \P2_EBX_reg[27]/NET0131  & ~n19912 ;
  assign n19915 = ~n1920 & ~n19913 ;
  assign n19916 = ~n19914 & n19915 ;
  assign n19906 = ~\P2_rEIP_reg[27]/NET0131  & ~n16547 ;
  assign n19907 = ~n16548 & ~n19906 ;
  assign n19908 = n1920 & ~n19907 ;
  assign n19917 = n10236 & ~n19908 ;
  assign n19918 = ~n19916 & n19917 ;
  assign n19904 = \P2_rEIP_reg[27]/NET0131  & ~n16555 ;
  assign n19909 = ~n1819 & n19908 ;
  assign n19905 = ~\P2_EBX_reg[27]/NET0131  & ~n16558 ;
  assign n19910 = n15980 & ~n19905 ;
  assign n19911 = ~n19909 & n19910 ;
  assign n19919 = ~n19904 & ~n19911 ;
  assign n19920 = ~n19918 & n19919 ;
  assign n19921 = n1927 & ~n19920 ;
  assign n19922 = \P2_rEIP_reg[27]/NET0131  & ~n16511 ;
  assign n19923 = \P2_PhyAddrPointer_reg[27]/NET0131  & n2987 ;
  assign n19924 = ~n19922 & ~n19923 ;
  assign n19925 = ~n19921 & n19924 ;
  assign n19926 = ~n19903 & n19925 ;
  assign n19927 = ~\P2_rEIP_reg[28]/NET0131  & ~n16548 ;
  assign n19928 = n1920 & ~n16549 ;
  assign n19929 = ~n19927 & n19928 ;
  assign n19930 = ~\P2_EBX_reg[27]/NET0131  & n16585 ;
  assign n19931 = \P2_EBX_reg[31]/NET0131  & ~n19930 ;
  assign n19933 = \P2_EBX_reg[28]/NET0131  & n19931 ;
  assign n19932 = ~\P2_EBX_reg[28]/NET0131  & ~n19931 ;
  assign n19934 = ~n1920 & ~n19932 ;
  assign n19935 = ~n19933 & n19934 ;
  assign n19936 = ~n19929 & ~n19935 ;
  assign n19937 = n10236 & ~n19936 ;
  assign n19938 = \P2_rEIP_reg[28]/NET0131  & n19391 ;
  assign n19940 = \P2_EBX_reg[28]/NET0131  & ~n1920 ;
  assign n19941 = ~n19929 & ~n19940 ;
  assign n19942 = n1921 & ~n19941 ;
  assign n19939 = \P2_rEIP_reg[28]/NET0131  & n1810 ;
  assign n19943 = \P2_EBX_reg[28]/NET0131  & n1819 ;
  assign n19944 = ~n1810 & n19943 ;
  assign n19945 = ~n19939 & ~n19944 ;
  assign n19946 = ~n19942 & n19945 ;
  assign n19947 = n1743 & ~n19946 ;
  assign n19948 = ~n19938 & ~n19947 ;
  assign n19949 = ~n19937 & n19948 ;
  assign n19950 = n1927 & ~n19949 ;
  assign n19952 = ~n9003 & ~n16518 ;
  assign n19954 = ~n11063 & n19952 ;
  assign n19953 = n11063 & ~n19952 ;
  assign n19955 = ~\P2_DataWidth_reg[1]/NET0131  & ~n19953 ;
  assign n19956 = ~n19954 & n19955 ;
  assign n19951 = \P2_DataWidth_reg[1]/NET0131  & ~\P2_rEIP_reg[28]/NET0131  ;
  assign n19957 = n1931 & ~n19951 ;
  assign n19958 = ~n19956 & n19957 ;
  assign n19959 = \P2_PhyAddrPointer_reg[28]/NET0131  & n2987 ;
  assign n19960 = \P2_rEIP_reg[28]/NET0131  & ~n16511 ;
  assign n19961 = ~n19959 & ~n19960 ;
  assign n19962 = ~n19958 & n19961 ;
  assign n19963 = ~n19950 & n19962 ;
  assign n19965 = \P1_PhyAddrPointer_reg[3]/NET0131  & n19830 ;
  assign n19966 = n18540 & ~n19965 ;
  assign n19968 = n15829 & ~n19966 ;
  assign n19967 = ~n15829 & n19966 ;
  assign n19969 = ~\P1_DataWidth_reg[1]/NET0131  & ~n19967 ;
  assign n19970 = ~n19968 & n19969 ;
  assign n19964 = \P1_DataWidth_reg[1]/NET0131  & ~\P1_rEIP_reg[4]/NET0131  ;
  assign n19971 = n2436 & ~n19964 ;
  assign n19972 = ~n19970 & n19971 ;
  assign n19974 = \P1_rEIP_reg[4]/NET0131  & ~n18554 ;
  assign n19975 = \P1_EBX_reg[31]/NET0131  & ~n18579 ;
  assign n19977 = ~\P1_EBX_reg[4]/NET0131  & n19975 ;
  assign n19976 = \P1_EBX_reg[4]/NET0131  & ~n19975 ;
  assign n19978 = ~n2425 & ~n19976 ;
  assign n19979 = ~n19977 & n19978 ;
  assign n19980 = ~\P1_rEIP_reg[4]/NET0131  & ~n18559 ;
  assign n19981 = ~n18560 & ~n19980 ;
  assign n19982 = n2425 & ~n19981 ;
  assign n19983 = ~n19979 & ~n19982 ;
  assign n19984 = n7246 & n19983 ;
  assign n19985 = ~\P1_EBX_reg[4]/NET0131  & ~n18556 ;
  assign n19986 = n18556 & ~n19981 ;
  assign n19987 = ~n19985 & ~n19986 ;
  assign n19988 = n15990 & n19987 ;
  assign n19989 = ~n19984 & ~n19988 ;
  assign n19990 = ~n19974 & n19989 ;
  assign n19991 = n2432 & ~n19990 ;
  assign n19973 = \P1_rEIP_reg[4]/NET0131  & ~n18552 ;
  assign n19992 = \P1_PhyAddrPointer_reg[4]/NET0131  & n3028 ;
  assign n19993 = ~n5092 & ~n19992 ;
  assign n19994 = ~n19973 & n19993 ;
  assign n19995 = ~n19991 & n19994 ;
  assign n19996 = ~n19972 & n19995 ;
  assign n19998 = \P2_PhyAddrPointer_reg[31]/NET0131  & ~n8998 ;
  assign n19999 = ~n19885 & ~n19998 ;
  assign n20001 = ~n11079 & ~n19999 ;
  assign n20000 = n11079 & n19999 ;
  assign n20002 = ~\P2_DataWidth_reg[1]/NET0131  & ~n20000 ;
  assign n20003 = ~n20001 & n20002 ;
  assign n19997 = \P2_DataWidth_reg[1]/NET0131  & ~\P2_rEIP_reg[29]/NET0131  ;
  assign n20004 = n1931 & ~n19997 ;
  assign n20005 = ~n20003 & n20004 ;
  assign n20009 = \P2_EBX_reg[31]/NET0131  & ~n16587 ;
  assign n20011 = ~\P2_EBX_reg[29]/NET0131  & n20009 ;
  assign n20010 = \P2_EBX_reg[29]/NET0131  & ~n20009 ;
  assign n20012 = ~n1920 & ~n20010 ;
  assign n20013 = ~n20011 & n20012 ;
  assign n20006 = ~\P2_rEIP_reg[29]/NET0131  & ~n16549 ;
  assign n20007 = ~n16550 & ~n20006 ;
  assign n20008 = n1920 & ~n20007 ;
  assign n20014 = n10236 & ~n20008 ;
  assign n20015 = ~n20013 & n20014 ;
  assign n20016 = n16558 & n20007 ;
  assign n20017 = \P2_EBX_reg[29]/NET0131  & ~n16558 ;
  assign n20018 = ~n1810 & ~n20017 ;
  assign n20019 = ~n20016 & n20018 ;
  assign n20020 = n1743 & ~n20019 ;
  assign n20021 = ~n19391 & ~n20020 ;
  assign n20022 = \P2_rEIP_reg[29]/NET0131  & ~n20021 ;
  assign n20023 = ~n1810 & n20020 ;
  assign n20024 = ~n20022 & ~n20023 ;
  assign n20025 = ~n20015 & n20024 ;
  assign n20026 = n1927 & ~n20025 ;
  assign n20027 = \P2_PhyAddrPointer_reg[29]/NET0131  & n2987 ;
  assign n20028 = \P2_rEIP_reg[29]/NET0131  & ~n16511 ;
  assign n20029 = ~n20027 & ~n20028 ;
  assign n20030 = ~n20026 & n20029 ;
  assign n20031 = ~n20005 & n20030 ;
  assign n20033 = ~\P2_PhyAddrPointer_reg[1]/NET0131  & ~\P2_PhyAddrPointer_reg[2]/NET0131  ;
  assign n20034 = ~n15745 & ~n20033 ;
  assign n20036 = n19056 & ~n20034 ;
  assign n20035 = ~n19056 & n20034 ;
  assign n20037 = ~\P2_DataWidth_reg[1]/NET0131  & ~n20035 ;
  assign n20038 = ~n20036 & n20037 ;
  assign n20032 = \P2_DataWidth_reg[1]/NET0131  & ~\P2_rEIP_reg[2]/NET0131  ;
  assign n20039 = n1931 & ~n20032 ;
  assign n20040 = ~n20038 & n20039 ;
  assign n20043 = \P2_rEIP_reg[2]/NET0131  & ~n16555 ;
  assign n20056 = \P2_EBX_reg[2]/NET0131  & ~n16558 ;
  assign n20045 = ~\P2_rEIP_reg[1]/NET0131  & ~\P2_rEIP_reg[2]/NET0131  ;
  assign n20046 = ~\P2_DataWidth_reg[1]/NET0131  & ~n16524 ;
  assign n20047 = ~n20045 & n20046 ;
  assign n20057 = n1820 & n20047 ;
  assign n20058 = ~n20056 & ~n20057 ;
  assign n20059 = n1743 & ~n20058 ;
  assign n20044 = n1444 & n1745 ;
  assign n20048 = ~n1805 & n20047 ;
  assign n20049 = \P2_EBX_reg[31]/NET0131  & ~n16560 ;
  assign n20051 = \P2_EBX_reg[2]/NET0131  & n20049 ;
  assign n20050 = ~\P2_EBX_reg[2]/NET0131  & ~n20049 ;
  assign n20052 = ~n1920 & ~n20050 ;
  assign n20053 = ~n20051 & n20052 ;
  assign n20054 = ~n20048 & ~n20053 ;
  assign n20055 = n1742 & ~n20054 ;
  assign n20060 = ~n20044 & ~n20055 ;
  assign n20061 = ~n20059 & n20060 ;
  assign n20062 = ~n1810 & ~n20061 ;
  assign n20063 = ~n20043 & ~n20062 ;
  assign n20064 = n1927 & ~n20063 ;
  assign n20041 = \P2_PhyAddrPointer_reg[2]/NET0131  & n2987 ;
  assign n20042 = \P2_rEIP_reg[2]/NET0131  & ~n16511 ;
  assign n20065 = ~n20041 & ~n20042 ;
  assign n20066 = ~n20064 & n20065 ;
  assign n20067 = ~n20040 & n20066 ;
  assign n20069 = n10094 & n18541 ;
  assign n20070 = n18540 & ~n20069 ;
  assign n20072 = n16290 & ~n20070 ;
  assign n20071 = ~n16290 & n20070 ;
  assign n20073 = ~\P1_DataWidth_reg[1]/NET0131  & ~n20071 ;
  assign n20074 = ~n20072 & n20073 ;
  assign n20068 = \P1_DataWidth_reg[1]/NET0131  & ~\P1_rEIP_reg[6]/NET0131  ;
  assign n20075 = n2436 & ~n20068 ;
  assign n20076 = ~n20074 & n20075 ;
  assign n20078 = \P1_rEIP_reg[6]/NET0131  & ~n18554 ;
  assign n20079 = ~\P1_rEIP_reg[6]/NET0131  & ~n18561 ;
  assign n20080 = ~n18562 & ~n20079 ;
  assign n20081 = n2425 & ~n20080 ;
  assign n20082 = ~n2311 & n20081 ;
  assign n20083 = ~\P1_EBX_reg[6]/NET0131  & ~n18556 ;
  assign n20084 = ~n20082 & ~n20083 ;
  assign n20085 = n15990 & n20084 ;
  assign n20086 = \P1_EBX_reg[31]/NET0131  & ~n18581 ;
  assign n20088 = \P1_EBX_reg[6]/NET0131  & ~n20086 ;
  assign n20087 = ~\P1_EBX_reg[6]/NET0131  & n20086 ;
  assign n20089 = ~n2425 & ~n20087 ;
  assign n20090 = ~n20088 & n20089 ;
  assign n20091 = ~n20081 & ~n20090 ;
  assign n20092 = n7246 & n20091 ;
  assign n20093 = ~n20085 & ~n20092 ;
  assign n20094 = ~n20078 & n20093 ;
  assign n20095 = n2432 & ~n20094 ;
  assign n20077 = \P1_rEIP_reg[6]/NET0131  & ~n18552 ;
  assign n20096 = \P1_PhyAddrPointer_reg[6]/NET0131  & n3028 ;
  assign n20097 = ~n5092 & ~n20096 ;
  assign n20098 = ~n20077 & n20097 ;
  assign n20099 = ~n20095 & n20098 ;
  assign n20100 = ~n20076 & n20099 ;
  assign n20102 = ~\P2_PhyAddrPointer_reg[0]/NET0131  & n15745 ;
  assign n20103 = ~n9003 & ~n20102 ;
  assign n20105 = ~n16142 & n20103 ;
  assign n20104 = n16142 & ~n20103 ;
  assign n20106 = ~\P2_DataWidth_reg[1]/NET0131  & ~n20104 ;
  assign n20107 = ~n20105 & n20106 ;
  assign n20101 = \P2_DataWidth_reg[1]/NET0131  & ~\P2_rEIP_reg[3]/NET0131  ;
  assign n20108 = n1931 & ~n20101 ;
  assign n20109 = ~n20107 & n20108 ;
  assign n20111 = \P2_rEIP_reg[3]/NET0131  & ~n16555 ;
  assign n20124 = \P2_EBX_reg[3]/NET0131  & ~n16558 ;
  assign n20118 = ~\P2_rEIP_reg[3]/NET0131  & ~n16524 ;
  assign n20119 = ~\P2_DataWidth_reg[1]/NET0131  & ~n16525 ;
  assign n20120 = ~n20118 & n20119 ;
  assign n20125 = n1820 & n20120 ;
  assign n20126 = ~n20124 & ~n20125 ;
  assign n20127 = n1743 & ~n20126 ;
  assign n20112 = n1745 & n1861 ;
  assign n20113 = \P2_EBX_reg[31]/NET0131  & ~n16561 ;
  assign n20115 = \P2_EBX_reg[3]/NET0131  & n20113 ;
  assign n20114 = ~\P2_EBX_reg[3]/NET0131  & ~n20113 ;
  assign n20116 = ~n1920 & ~n20114 ;
  assign n20117 = ~n20115 & n20116 ;
  assign n20121 = ~n1805 & n20120 ;
  assign n20122 = ~n20117 & ~n20121 ;
  assign n20123 = n1742 & ~n20122 ;
  assign n20128 = ~n20112 & ~n20123 ;
  assign n20129 = ~n20127 & n20128 ;
  assign n20130 = ~n1810 & ~n20129 ;
  assign n20131 = ~n20111 & ~n20130 ;
  assign n20132 = n1927 & ~n20131 ;
  assign n20110 = \P2_rEIP_reg[3]/NET0131  & ~n16511 ;
  assign n20133 = ~n16144 & ~n20110 ;
  assign n20134 = ~n20132 & n20133 ;
  assign n20135 = ~n20109 & n20134 ;
  assign n20137 = ~n8960 & ~n9003 ;
  assign n20138 = ~n19056 & ~n20137 ;
  assign n20140 = ~n15749 & ~n20138 ;
  assign n20139 = n15749 & n20138 ;
  assign n20141 = ~\P2_DataWidth_reg[1]/NET0131  & ~n20139 ;
  assign n20142 = ~n20140 & n20141 ;
  assign n20136 = \P2_DataWidth_reg[1]/NET0131  & ~\P2_rEIP_reg[4]/NET0131  ;
  assign n20143 = n1931 & ~n20136 ;
  assign n20144 = ~n20142 & n20143 ;
  assign n20149 = \P2_EBX_reg[31]/NET0131  & ~n16562 ;
  assign n20155 = ~n16559 & n20149 ;
  assign n20156 = \P2_EBX_reg[4]/NET0131  & ~n19071 ;
  assign n20157 = ~n20155 & n20156 ;
  assign n20150 = ~\P2_EBX_reg[4]/NET0131  & n20149 ;
  assign n20151 = n16589 & n20150 ;
  assign n20152 = ~\P2_rEIP_reg[4]/NET0131  & ~n16525 ;
  assign n20153 = ~n16526 & ~n20152 ;
  assign n20154 = n16553 & n20153 ;
  assign n20158 = ~n20151 & ~n20154 ;
  assign n20159 = ~n20157 & n20158 ;
  assign n20160 = n1927 & ~n20159 ;
  assign n20146 = n1927 & ~n16555 ;
  assign n20147 = n18989 & ~n20146 ;
  assign n20148 = \P2_rEIP_reg[4]/NET0131  & ~n20147 ;
  assign n20145 = \P2_PhyAddrPointer_reg[4]/NET0131  & n2987 ;
  assign n20161 = ~n3113 & ~n20145 ;
  assign n20162 = ~n20148 & n20161 ;
  assign n20163 = ~n20160 & n20162 ;
  assign n20164 = ~n20144 & n20163 ;
  assign n20166 = ~\P1_PhyAddrPointer_reg[0]/NET0131  & n14588 ;
  assign n20167 = n18540 & ~n20166 ;
  assign n20169 = n14590 & ~n20167 ;
  assign n20168 = ~n14590 & n20167 ;
  assign n20170 = ~\P1_DataWidth_reg[1]/NET0131  & ~n20168 ;
  assign n20171 = ~n20169 & n20170 ;
  assign n20165 = \P1_DataWidth_reg[1]/NET0131  & ~\P1_rEIP_reg[7]/NET0131  ;
  assign n20172 = n2436 & ~n20165 ;
  assign n20173 = ~n20171 & n20172 ;
  assign n20175 = \P1_rEIP_reg[7]/NET0131  & ~n18554 ;
  assign n20176 = ~\P1_EBX_reg[7]/NET0131  & ~n18556 ;
  assign n20177 = ~\P1_rEIP_reg[7]/NET0131  & ~n18562 ;
  assign n20178 = ~n18563 & ~n20177 ;
  assign n20179 = n18556 & ~n20178 ;
  assign n20180 = ~n20176 & ~n20179 ;
  assign n20181 = n2225 & n20180 ;
  assign n20183 = \P1_EBX_reg[31]/NET0131  & ~n18582 ;
  assign n20185 = ~\P1_EBX_reg[7]/NET0131  & n20183 ;
  assign n20184 = \P1_EBX_reg[7]/NET0131  & ~n20183 ;
  assign n20186 = ~n2425 & ~n20184 ;
  assign n20187 = ~n20185 & n20186 ;
  assign n20182 = n2425 & ~n20178 ;
  assign n20188 = n2222 & ~n20182 ;
  assign n20189 = ~n20187 & n20188 ;
  assign n20190 = ~n20181 & ~n20189 ;
  assign n20191 = ~n2301 & ~n20190 ;
  assign n20192 = ~n20175 & ~n20191 ;
  assign n20193 = n2432 & ~n20192 ;
  assign n20174 = \P1_rEIP_reg[7]/NET0131  & ~n18552 ;
  assign n20194 = \P1_PhyAddrPointer_reg[7]/NET0131  & n3028 ;
  assign n20195 = ~n5092 & ~n20194 ;
  assign n20196 = ~n20174 & n20195 ;
  assign n20197 = ~n20193 & n20196 ;
  assign n20198 = ~n20173 & n20197 ;
  assign n20200 = \P1_PhyAddrPointer_reg[7]/NET0131  & n20166 ;
  assign n20201 = n18540 & ~n20200 ;
  assign n20203 = ~n13493 & n20201 ;
  assign n20202 = n13493 & ~n20201 ;
  assign n20204 = ~\P1_DataWidth_reg[1]/NET0131  & ~n20202 ;
  assign n20205 = ~n20203 & n20204 ;
  assign n20199 = \P1_DataWidth_reg[1]/NET0131  & ~\P1_rEIP_reg[8]/NET0131  ;
  assign n20206 = n2436 & ~n20199 ;
  assign n20207 = ~n20205 & n20206 ;
  assign n20209 = \P1_rEIP_reg[8]/NET0131  & ~n18554 ;
  assign n20210 = ~\P1_EBX_reg[8]/NET0131  & ~n18556 ;
  assign n20211 = ~\P1_rEIP_reg[8]/NET0131  & ~n18563 ;
  assign n20212 = ~n18564 & ~n20211 ;
  assign n20213 = n18556 & ~n20212 ;
  assign n20214 = ~n20210 & ~n20213 ;
  assign n20215 = n2225 & n20214 ;
  assign n20217 = \P1_EBX_reg[31]/NET0131  & ~n18583 ;
  assign n20219 = ~\P1_EBX_reg[8]/NET0131  & n20217 ;
  assign n20218 = \P1_EBX_reg[8]/NET0131  & ~n20217 ;
  assign n20220 = ~n2425 & ~n20218 ;
  assign n20221 = ~n20219 & n20220 ;
  assign n20216 = n2425 & ~n20212 ;
  assign n20222 = n2222 & ~n20216 ;
  assign n20223 = ~n20221 & n20222 ;
  assign n20224 = ~n20215 & ~n20223 ;
  assign n20225 = ~n2301 & ~n20224 ;
  assign n20226 = ~n20209 & ~n20225 ;
  assign n20227 = n2432 & ~n20226 ;
  assign n20208 = \P1_rEIP_reg[8]/NET0131  & ~n18552 ;
  assign n20228 = \P1_PhyAddrPointer_reg[8]/NET0131  & n3028 ;
  assign n20229 = ~n5092 & ~n20228 ;
  assign n20230 = ~n20208 & n20229 ;
  assign n20231 = ~n20227 & n20230 ;
  assign n20232 = ~n20207 & n20231 ;
  assign n20234 = n8962 & n16514 ;
  assign n20235 = ~n9003 & ~n20234 ;
  assign n20237 = ~n16180 & n20235 ;
  assign n20236 = n16180 & ~n20235 ;
  assign n20238 = ~\P2_DataWidth_reg[1]/NET0131  & ~n20236 ;
  assign n20239 = ~n20237 & n20238 ;
  assign n20233 = \P2_DataWidth_reg[1]/NET0131  & ~\P2_rEIP_reg[6]/NET0131  ;
  assign n20240 = n1931 & ~n20233 ;
  assign n20241 = ~n20239 & n20240 ;
  assign n20250 = \P2_rEIP_reg[5]/NET0131  & n16526 ;
  assign n20251 = \P2_rEIP_reg[6]/NET0131  & n20250 ;
  assign n20252 = ~\P2_rEIP_reg[6]/NET0131  & ~n20250 ;
  assign n20253 = ~n20251 & ~n20252 ;
  assign n20254 = n16553 & n20253 ;
  assign n20244 = \P2_EBX_reg[31]/NET0131  & ~n16564 ;
  assign n20245 = ~n15980 & n20244 ;
  assign n20246 = \P2_EBX_reg[6]/NET0131  & ~n20245 ;
  assign n20247 = ~n19071 & n20246 ;
  assign n20243 = \P2_rEIP_reg[6]/NET0131  & ~n16555 ;
  assign n20248 = ~\P2_EBX_reg[6]/NET0131  & n20244 ;
  assign n20249 = n16589 & n20248 ;
  assign n20255 = ~n20243 & ~n20249 ;
  assign n20256 = ~n20247 & n20255 ;
  assign n20257 = ~n20254 & n20256 ;
  assign n20258 = n1927 & ~n20257 ;
  assign n20242 = \P2_rEIP_reg[6]/NET0131  & ~n18989 ;
  assign n20259 = \P2_PhyAddrPointer_reg[6]/NET0131  & n2987 ;
  assign n20260 = ~n3113 & ~n20259 ;
  assign n20261 = ~n20242 & n20260 ;
  assign n20262 = ~n20258 & n20261 ;
  assign n20263 = ~n20241 & n20262 ;
  assign n20265 = ~n9003 & ~n13043 ;
  assign n20266 = ~n19563 & ~n20265 ;
  assign n20268 = n14428 & n20266 ;
  assign n20267 = ~n14428 & ~n20266 ;
  assign n20269 = ~\P2_DataWidth_reg[1]/NET0131  & ~n20267 ;
  assign n20270 = ~n20268 & n20269 ;
  assign n20264 = \P2_DataWidth_reg[1]/NET0131  & ~\P2_rEIP_reg[7]/NET0131  ;
  assign n20271 = n1931 & ~n20264 ;
  assign n20272 = ~n20270 & n20271 ;
  assign n20274 = \P2_rEIP_reg[7]/NET0131  & ~n16555 ;
  assign n20275 = ~\P2_EBX_reg[7]/NET0131  & ~n16558 ;
  assign n20276 = ~\P2_rEIP_reg[7]/NET0131  & ~n20251 ;
  assign n20277 = ~n16529 & ~n20276 ;
  assign n20278 = n16558 & ~n20277 ;
  assign n20279 = ~n20275 & ~n20278 ;
  assign n20280 = n15980 & n20279 ;
  assign n20281 = n1920 & ~n20277 ;
  assign n20282 = \P2_EBX_reg[31]/NET0131  & ~n16565 ;
  assign n20284 = ~\P2_EBX_reg[7]/NET0131  & n20282 ;
  assign n20283 = \P2_EBX_reg[7]/NET0131  & ~n20282 ;
  assign n20285 = ~n1920 & ~n20283 ;
  assign n20286 = ~n20284 & n20285 ;
  assign n20287 = ~n20281 & ~n20286 ;
  assign n20288 = n10236 & n20287 ;
  assign n20289 = ~n20280 & ~n20288 ;
  assign n20290 = ~n20274 & n20289 ;
  assign n20291 = n1927 & ~n20290 ;
  assign n20273 = \P2_rEIP_reg[7]/NET0131  & ~n18989 ;
  assign n20292 = \P2_PhyAddrPointer_reg[7]/NET0131  & n2987 ;
  assign n20293 = ~n3113 & ~n20292 ;
  assign n20294 = ~n20273 & n20293 ;
  assign n20295 = ~n20291 & n20294 ;
  assign n20296 = ~n20272 & n20295 ;
  assign n20298 = n18540 & ~n18542 ;
  assign n20300 = ~n14599 & n20298 ;
  assign n20299 = n14599 & ~n20298 ;
  assign n20301 = ~\P1_DataWidth_reg[1]/NET0131  & ~n20299 ;
  assign n20302 = ~n20300 & n20301 ;
  assign n20297 = \P1_DataWidth_reg[1]/NET0131  & ~\P1_rEIP_reg[9]/NET0131  ;
  assign n20303 = n2436 & ~n20297 ;
  assign n20304 = ~n20302 & n20303 ;
  assign n20306 = \P1_rEIP_reg[9]/NET0131  & ~n18554 ;
  assign n20308 = ~\P1_rEIP_reg[9]/NET0131  & ~n18564 ;
  assign n20309 = ~n18565 & ~n20308 ;
  assign n20310 = n18556 & ~n20309 ;
  assign n20307 = ~\P1_EBX_reg[9]/NET0131  & ~n18556 ;
  assign n20311 = n2225 & ~n20307 ;
  assign n20312 = ~n20310 & n20311 ;
  assign n20314 = \P1_EBX_reg[31]/NET0131  & ~n18584 ;
  assign n20316 = ~\P1_EBX_reg[9]/NET0131  & n20314 ;
  assign n20315 = \P1_EBX_reg[9]/NET0131  & ~n20314 ;
  assign n20317 = ~n2425 & ~n20315 ;
  assign n20318 = ~n20316 & n20317 ;
  assign n20313 = n2425 & ~n20309 ;
  assign n20319 = n2222 & ~n20313 ;
  assign n20320 = ~n20318 & n20319 ;
  assign n20321 = ~n20312 & ~n20320 ;
  assign n20322 = ~n2301 & ~n20321 ;
  assign n20323 = ~n20306 & ~n20322 ;
  assign n20324 = n2432 & ~n20323 ;
  assign n20305 = \P1_rEIP_reg[9]/NET0131  & ~n18552 ;
  assign n20325 = \P1_PhyAddrPointer_reg[9]/NET0131  & n3028 ;
  assign n20326 = ~n5092 & ~n20325 ;
  assign n20327 = ~n20305 & n20326 ;
  assign n20328 = ~n20324 & n20327 ;
  assign n20329 = ~n20304 & n20328 ;
  assign n20331 = ~n8964 & ~n9003 ;
  assign n20332 = ~n19056 & ~n20331 ;
  assign n20334 = ~n13047 & ~n20332 ;
  assign n20333 = n13047 & n20332 ;
  assign n20335 = ~\P2_DataWidth_reg[1]/NET0131  & ~n20333 ;
  assign n20336 = ~n20334 & n20335 ;
  assign n20330 = \P2_DataWidth_reg[1]/NET0131  & ~\P2_rEIP_reg[8]/NET0131  ;
  assign n20337 = n1931 & ~n20330 ;
  assign n20338 = ~n20336 & n20337 ;
  assign n20340 = \P2_rEIP_reg[8]/NET0131  & ~n16555 ;
  assign n20341 = \P2_EBX_reg[31]/NET0131  & ~n16566 ;
  assign n20343 = \P2_EBX_reg[8]/NET0131  & n20341 ;
  assign n20342 = ~\P2_EBX_reg[8]/NET0131  & ~n20341 ;
  assign n20344 = ~n1920 & ~n20342 ;
  assign n20345 = ~n20343 & n20344 ;
  assign n20346 = ~\P2_rEIP_reg[8]/NET0131  & ~n16529 ;
  assign n20347 = ~n16530 & ~n20346 ;
  assign n20348 = ~\P2_DataWidth_reg[1]/NET0131  & n20347 ;
  assign n20349 = ~n1805 & n20348 ;
  assign n20350 = ~n20345 & ~n20349 ;
  assign n20351 = n1742 & ~n20350 ;
  assign n20352 = \P2_EBX_reg[8]/NET0131  & ~n16558 ;
  assign n20353 = n1820 & n20348 ;
  assign n20354 = ~n20352 & ~n20353 ;
  assign n20355 = n1743 & ~n20354 ;
  assign n20356 = ~n20351 & ~n20355 ;
  assign n20357 = ~n1810 & ~n20356 ;
  assign n20358 = ~n20340 & ~n20357 ;
  assign n20359 = n1927 & ~n20358 ;
  assign n20339 = \P2_rEIP_reg[8]/NET0131  & ~n18989 ;
  assign n20360 = \P2_PhyAddrPointer_reg[8]/NET0131  & n2987 ;
  assign n20361 = ~n3113 & ~n20360 ;
  assign n20362 = ~n20339 & n20361 ;
  assign n20363 = ~n20359 & n20362 ;
  assign n20364 = ~n20338 & n20363 ;
  assign n20366 = ~n8965 & ~n9003 ;
  assign n20367 = ~n19056 & ~n20366 ;
  assign n20369 = ~n14448 & ~n20367 ;
  assign n20368 = n14448 & n20367 ;
  assign n20370 = ~\P2_DataWidth_reg[1]/NET0131  & ~n20368 ;
  assign n20371 = ~n20369 & n20370 ;
  assign n20365 = \P2_DataWidth_reg[1]/NET0131  & ~\P2_rEIP_reg[9]/NET0131  ;
  assign n20372 = n1931 & ~n20365 ;
  assign n20373 = ~n20371 & n20372 ;
  assign n20375 = \P2_rEIP_reg[9]/NET0131  & ~n16555 ;
  assign n20376 = ~\P2_EBX_reg[9]/NET0131  & ~n16558 ;
  assign n20377 = ~\P2_rEIP_reg[9]/NET0131  & ~n16530 ;
  assign n20378 = ~n16531 & ~n20377 ;
  assign n20379 = n16558 & ~n20378 ;
  assign n20380 = ~n20376 & ~n20379 ;
  assign n20381 = n1743 & n20380 ;
  assign n20383 = \P2_EBX_reg[31]/NET0131  & ~n16567 ;
  assign n20385 = ~\P2_EBX_reg[9]/NET0131  & n20383 ;
  assign n20384 = \P2_EBX_reg[9]/NET0131  & ~n20383 ;
  assign n20386 = ~n1920 & ~n20384 ;
  assign n20387 = ~n20385 & n20386 ;
  assign n20382 = n1920 & ~n20378 ;
  assign n20388 = n1742 & ~n20382 ;
  assign n20389 = ~n20387 & n20388 ;
  assign n20390 = ~n20381 & ~n20389 ;
  assign n20391 = ~n1810 & ~n20390 ;
  assign n20392 = ~n20375 & ~n20391 ;
  assign n20393 = n1927 & ~n20392 ;
  assign n20374 = \P2_rEIP_reg[9]/NET0131  & ~n18989 ;
  assign n20394 = \P2_PhyAddrPointer_reg[9]/NET0131  & n2987 ;
  assign n20395 = ~n3113 & ~n20394 ;
  assign n20396 = ~n20374 & n20395 ;
  assign n20397 = ~n20393 & n20396 ;
  assign n20398 = ~n20373 & n20397 ;
  assign n20400 = ~\P3_PhyAddrPointer_reg[0]/NET0131  & n13249 ;
  assign n20401 = n9026 & n20400 ;
  assign n20402 = ~n9054 & ~n20401 ;
  assign n20404 = n14470 & ~n20402 ;
  assign n20403 = ~n14470 & n20402 ;
  assign n20405 = ~\P3_DataWidth_reg[1]/NET0131  & ~n20403 ;
  assign n20406 = ~n20404 & n20405 ;
  assign n20399 = \P3_DataWidth_reg[1]/NET0131  & ~\P3_rEIP_reg[10]/NET0131  ;
  assign n20407 = n2959 & ~n20399 ;
  assign n20408 = ~n20406 & n20407 ;
  assign n20411 = \P3_rEIP_reg[10]/NET0131  & n2910 ;
  assign n20412 = ~n2786 & n2946 ;
  assign n20414 = \P3_rEIP_reg[1]/NET0131  & \P3_rEIP_reg[2]/NET0131  ;
  assign n20415 = \P3_rEIP_reg[3]/NET0131  & n20414 ;
  assign n20416 = \P3_rEIP_reg[4]/NET0131  & n20415 ;
  assign n20417 = \P3_rEIP_reg[5]/NET0131  & n20416 ;
  assign n20418 = \P3_rEIP_reg[6]/NET0131  & n20417 ;
  assign n20419 = \P3_rEIP_reg[7]/NET0131  & n20418 ;
  assign n20420 = \P3_rEIP_reg[8]/NET0131  & n20419 ;
  assign n20421 = \P3_rEIP_reg[9]/NET0131  & n20420 ;
  assign n20422 = ~\P3_rEIP_reg[10]/NET0131  & ~n20421 ;
  assign n20423 = \P3_rEIP_reg[10]/NET0131  & n20421 ;
  assign n20424 = ~n20422 & ~n20423 ;
  assign n20425 = n20412 & ~n20424 ;
  assign n20413 = ~\P3_EBX_reg[10]/NET0131  & ~n20412 ;
  assign n20426 = n2818 & ~n20413 ;
  assign n20427 = ~n20425 & n20426 ;
  assign n20429 = ~\P3_EBX_reg[0]/NET0131  & ~\P3_EBX_reg[1]/NET0131  ;
  assign n20430 = ~\P3_EBX_reg[2]/NET0131  & n20429 ;
  assign n20431 = ~\P3_EBX_reg[3]/NET0131  & n20430 ;
  assign n20432 = ~\P3_EBX_reg[4]/NET0131  & n20431 ;
  assign n20433 = ~\P3_EBX_reg[5]/NET0131  & n20432 ;
  assign n20434 = ~\P3_EBX_reg[6]/NET0131  & n20433 ;
  assign n20435 = ~\P3_EBX_reg[7]/NET0131  & n20434 ;
  assign n20436 = ~\P3_EBX_reg[8]/NET0131  & n20435 ;
  assign n20437 = ~\P3_EBX_reg[9]/NET0131  & n20436 ;
  assign n20438 = \P3_EBX_reg[31]/NET0131  & ~n20437 ;
  assign n20440 = ~\P3_EBX_reg[10]/NET0131  & n20438 ;
  assign n20439 = \P3_EBX_reg[10]/NET0131  & ~n20438 ;
  assign n20441 = ~n2946 & ~n20439 ;
  assign n20442 = ~n20440 & n20441 ;
  assign n20428 = n2946 & ~n20424 ;
  assign n20443 = n2821 & ~n20428 ;
  assign n20444 = ~n20442 & n20443 ;
  assign n20445 = ~n20427 & ~n20444 ;
  assign n20446 = ~n2815 & ~n20445 ;
  assign n20447 = ~n20411 & ~n20446 ;
  assign n20448 = n2453 & ~n20447 ;
  assign n20409 = n2954 & n2998 ;
  assign n20410 = \P3_rEIP_reg[10]/NET0131  & ~n20409 ;
  assign n20449 = \P3_PhyAddrPointer_reg[10]/NET0131  & n3004 ;
  assign n20450 = ~n4412 & ~n20449 ;
  assign n20451 = ~n20410 & n20450 ;
  assign n20452 = ~n20448 & n20451 ;
  assign n20453 = ~n20408 & n20452 ;
  assign n20455 = ~n14470 & n20401 ;
  assign n20456 = ~n9054 & ~n20455 ;
  assign n20458 = n11963 & ~n20456 ;
  assign n20457 = ~n11963 & n20456 ;
  assign n20459 = ~\P3_DataWidth_reg[1]/NET0131  & ~n20457 ;
  assign n20460 = ~n20458 & n20459 ;
  assign n20454 = \P3_DataWidth_reg[1]/NET0131  & ~\P3_rEIP_reg[11]/NET0131  ;
  assign n20461 = n2959 & ~n20454 ;
  assign n20462 = ~n20460 & n20461 ;
  assign n20474 = ~\P3_EBX_reg[10]/NET0131  & n20437 ;
  assign n20475 = \P3_EBX_reg[31]/NET0131  & ~n20474 ;
  assign n20477 = \P3_EBX_reg[11]/NET0131  & ~n20475 ;
  assign n20476 = ~\P3_EBX_reg[11]/NET0131  & n20475 ;
  assign n20478 = ~n2946 & ~n20476 ;
  assign n20479 = ~n20477 & n20478 ;
  assign n20466 = ~\P3_rEIP_reg[11]/NET0131  & ~n20423 ;
  assign n20467 = \P3_rEIP_reg[11]/NET0131  & n20423 ;
  assign n20468 = ~n20466 & ~n20467 ;
  assign n20469 = n2946 & ~n20468 ;
  assign n20473 = ~n2815 & n2821 ;
  assign n20480 = ~n20469 & n20473 ;
  assign n20481 = ~n20479 & n20480 ;
  assign n20464 = \P3_rEIP_reg[11]/NET0131  & n2910 ;
  assign n20470 = ~n2786 & n20469 ;
  assign n20465 = ~\P3_EBX_reg[11]/NET0131  & ~n20412 ;
  assign n20471 = n16094 & ~n20465 ;
  assign n20472 = ~n20470 & n20471 ;
  assign n20482 = ~n20464 & ~n20472 ;
  assign n20483 = ~n20481 & n20482 ;
  assign n20484 = n2453 & ~n20483 ;
  assign n20463 = \P3_rEIP_reg[11]/NET0131  & ~n20409 ;
  assign n20485 = \P3_PhyAddrPointer_reg[11]/NET0131  & n3004 ;
  assign n20486 = ~n4412 & ~n20485 ;
  assign n20487 = ~n20463 & n20486 ;
  assign n20488 = ~n20484 & n20487 ;
  assign n20489 = ~n20462 & n20488 ;
  assign n20491 = ~n11963 & n20455 ;
  assign n20492 = ~n9054 & ~n20491 ;
  assign n20494 = n13056 & ~n20492 ;
  assign n20493 = ~n13056 & n20492 ;
  assign n20495 = ~\P3_DataWidth_reg[1]/NET0131  & ~n20493 ;
  assign n20496 = ~n20494 & n20495 ;
  assign n20490 = \P3_DataWidth_reg[1]/NET0131  & ~\P3_rEIP_reg[12]/NET0131  ;
  assign n20497 = n2959 & ~n20490 ;
  assign n20498 = ~n20496 & n20497 ;
  assign n20500 = \P3_rEIP_reg[12]/NET0131  & n2910 ;
  assign n20501 = ~\P3_rEIP_reg[12]/NET0131  & ~n20467 ;
  assign n20502 = \P3_rEIP_reg[12]/NET0131  & n20467 ;
  assign n20503 = ~n20501 & ~n20502 ;
  assign n20504 = n2946 & ~n20503 ;
  assign n20505 = ~\P3_EBX_reg[12]/NET0131  & ~n20412 ;
  assign n20506 = n2818 & ~n20505 ;
  assign n20507 = ~\P3_EBX_reg[11]/NET0131  & n20474 ;
  assign n20508 = \P3_EBX_reg[31]/NET0131  & ~n20507 ;
  assign n20510 = ~\P3_EBX_reg[12]/NET0131  & n20508 ;
  assign n20509 = \P3_EBX_reg[12]/NET0131  & ~n20508 ;
  assign n20511 = ~n2946 & ~n20509 ;
  assign n20512 = ~n20510 & n20511 ;
  assign n20513 = n2821 & ~n20512 ;
  assign n20514 = ~n20506 & ~n20513 ;
  assign n20515 = ~n20504 & ~n20514 ;
  assign n20516 = n2786 & n20506 ;
  assign n20517 = ~n20515 & ~n20516 ;
  assign n20518 = ~n2815 & ~n20517 ;
  assign n20519 = ~n20500 & ~n20518 ;
  assign n20520 = n2453 & ~n20519 ;
  assign n20499 = \P3_rEIP_reg[12]/NET0131  & ~n20409 ;
  assign n20521 = \P3_PhyAddrPointer_reg[12]/NET0131  & n3004 ;
  assign n20522 = ~n4412 & ~n20521 ;
  assign n20523 = ~n20499 & n20522 ;
  assign n20524 = ~n20520 & n20523 ;
  assign n20525 = ~n20498 & n20524 ;
  assign n20527 = ~n13056 & n20491 ;
  assign n20528 = ~n9054 & ~n20527 ;
  assign n20530 = n13104 & ~n20528 ;
  assign n20529 = ~n13104 & n20528 ;
  assign n20531 = ~\P3_DataWidth_reg[1]/NET0131  & ~n20529 ;
  assign n20532 = ~n20530 & n20531 ;
  assign n20526 = \P3_DataWidth_reg[1]/NET0131  & ~\P3_rEIP_reg[13]/NET0131  ;
  assign n20533 = n2959 & ~n20526 ;
  assign n20534 = ~n20532 & n20533 ;
  assign n20536 = \P3_rEIP_reg[13]/NET0131  & n2910 ;
  assign n20540 = ~\P3_EBX_reg[13]/NET0131  & ~n20412 ;
  assign n20541 = n2818 & ~n20540 ;
  assign n20545 = ~\P3_EBX_reg[12]/NET0131  & n20507 ;
  assign n20546 = \P3_EBX_reg[31]/NET0131  & ~n20545 ;
  assign n20548 = \P3_EBX_reg[13]/NET0131  & ~n20546 ;
  assign n20547 = ~\P3_EBX_reg[13]/NET0131  & n20546 ;
  assign n20549 = ~n2946 & ~n20547 ;
  assign n20550 = ~n20548 & n20549 ;
  assign n20551 = n2821 & ~n20550 ;
  assign n20552 = ~n20541 & ~n20551 ;
  assign n20542 = n2786 & n20541 ;
  assign n20537 = ~\P3_rEIP_reg[13]/NET0131  & ~n20502 ;
  assign n20538 = \P3_rEIP_reg[13]/NET0131  & n20502 ;
  assign n20539 = ~n20537 & ~n20538 ;
  assign n20543 = n2946 & ~n20539 ;
  assign n20544 = ~n20542 & n20543 ;
  assign n20553 = ~n2815 & ~n20544 ;
  assign n20554 = ~n20552 & n20553 ;
  assign n20555 = ~n20536 & ~n20554 ;
  assign n20556 = n2453 & ~n20555 ;
  assign n20535 = \P3_rEIP_reg[13]/NET0131  & ~n20409 ;
  assign n20557 = \P3_PhyAddrPointer_reg[13]/NET0131  & n3004 ;
  assign n20558 = ~n4412 & ~n20557 ;
  assign n20559 = ~n20535 & n20558 ;
  assign n20560 = ~n20556 & n20559 ;
  assign n20561 = ~n20534 & n20560 ;
  assign n20563 = ~n13104 & n20527 ;
  assign n20564 = ~n9054 & ~n20563 ;
  assign n20566 = n13131 & ~n20564 ;
  assign n20565 = ~n13131 & n20564 ;
  assign n20567 = ~\P3_DataWidth_reg[1]/NET0131  & ~n20565 ;
  assign n20568 = ~n20566 & n20567 ;
  assign n20562 = \P3_DataWidth_reg[1]/NET0131  & ~\P3_rEIP_reg[14]/NET0131  ;
  assign n20569 = n2959 & ~n20562 ;
  assign n20570 = ~n20568 & n20569 ;
  assign n20572 = \P3_rEIP_reg[14]/NET0131  & n2910 ;
  assign n20574 = ~\P3_rEIP_reg[14]/NET0131  & ~n20538 ;
  assign n20575 = \P3_rEIP_reg[14]/NET0131  & n20538 ;
  assign n20576 = ~n20574 & ~n20575 ;
  assign n20577 = n20412 & ~n20576 ;
  assign n20573 = ~\P3_EBX_reg[14]/NET0131  & ~n20412 ;
  assign n20578 = n2818 & ~n20573 ;
  assign n20579 = ~n20577 & n20578 ;
  assign n20581 = ~\P3_EBX_reg[13]/NET0131  & n20545 ;
  assign n20582 = \P3_EBX_reg[31]/NET0131  & ~n20581 ;
  assign n20583 = ~\P3_EBX_reg[14]/NET0131  & ~n20582 ;
  assign n20584 = \P3_EBX_reg[14]/NET0131  & n20582 ;
  assign n20585 = ~n20583 & ~n20584 ;
  assign n20586 = ~n2946 & ~n20585 ;
  assign n20580 = n2946 & ~n20576 ;
  assign n20587 = n2821 & ~n20580 ;
  assign n20588 = ~n20586 & n20587 ;
  assign n20589 = ~n20579 & ~n20588 ;
  assign n20590 = ~n2815 & ~n20589 ;
  assign n20591 = ~n20572 & ~n20590 ;
  assign n20592 = n2453 & ~n20591 ;
  assign n20571 = \P3_rEIP_reg[14]/NET0131  & ~n20409 ;
  assign n20593 = \P3_PhyAddrPointer_reg[14]/NET0131  & n3004 ;
  assign n20594 = ~n4412 & ~n20593 ;
  assign n20595 = ~n20571 & n20594 ;
  assign n20596 = ~n20592 & n20595 ;
  assign n20597 = ~n20570 & n20596 ;
  assign n20599 = ~n13131 & n20563 ;
  assign n20600 = ~n9054 & ~n20599 ;
  assign n20602 = n12013 & ~n20600 ;
  assign n20601 = ~n12013 & n20600 ;
  assign n20603 = ~\P3_DataWidth_reg[1]/NET0131  & ~n20601 ;
  assign n20604 = ~n20602 & n20603 ;
  assign n20598 = \P3_DataWidth_reg[1]/NET0131  & ~\P3_rEIP_reg[15]/NET0131  ;
  assign n20605 = n2959 & ~n20598 ;
  assign n20606 = ~n20604 & n20605 ;
  assign n20608 = \P3_rEIP_reg[15]/NET0131  & n2910 ;
  assign n20612 = ~\P3_EBX_reg[15]/NET0131  & ~n20412 ;
  assign n20617 = n2818 & ~n20612 ;
  assign n20618 = ~\P3_EBX_reg[14]/NET0131  & n20581 ;
  assign n20619 = \P3_EBX_reg[31]/NET0131  & ~n20618 ;
  assign n20621 = ~\P3_EBX_reg[15]/NET0131  & n20619 ;
  assign n20620 = \P3_EBX_reg[15]/NET0131  & ~n20619 ;
  assign n20622 = ~n2946 & ~n20620 ;
  assign n20623 = ~n20621 & n20622 ;
  assign n20624 = n2821 & ~n20623 ;
  assign n20625 = ~n20617 & ~n20624 ;
  assign n20609 = ~\P3_rEIP_reg[15]/NET0131  & ~n20575 ;
  assign n20610 = \P3_rEIP_reg[15]/NET0131  & n20575 ;
  assign n20611 = ~n20609 & ~n20610 ;
  assign n20613 = n2786 & n2818 ;
  assign n20614 = ~n20612 & n20613 ;
  assign n20615 = n2946 & ~n20614 ;
  assign n20616 = ~n20611 & n20615 ;
  assign n20626 = ~n2815 & ~n20616 ;
  assign n20627 = ~n20625 & n20626 ;
  assign n20628 = ~n20608 & ~n20627 ;
  assign n20629 = n2453 & ~n20628 ;
  assign n20607 = \P3_rEIP_reg[15]/NET0131  & ~n20409 ;
  assign n20630 = \P3_PhyAddrPointer_reg[15]/NET0131  & n3004 ;
  assign n20631 = ~n4412 & ~n20630 ;
  assign n20632 = ~n20607 & n20631 ;
  assign n20633 = ~n20629 & n20632 ;
  assign n20634 = ~n20606 & n20633 ;
  assign n20636 = ~n12013 & n20599 ;
  assign n20637 = ~n9054 & ~n20636 ;
  assign n20639 = ~n13145 & n20637 ;
  assign n20638 = n13145 & ~n20637 ;
  assign n20640 = ~\P3_DataWidth_reg[1]/NET0131  & ~n20638 ;
  assign n20641 = ~n20639 & n20640 ;
  assign n20635 = \P3_DataWidth_reg[1]/NET0131  & ~\P3_rEIP_reg[16]/NET0131  ;
  assign n20642 = n2959 & ~n20635 ;
  assign n20643 = ~n20641 & n20642 ;
  assign n20653 = \P3_EBX_reg[15]/NET0131  & \P3_EBX_reg[31]/NET0131  ;
  assign n20654 = ~n20619 & ~n20653 ;
  assign n20655 = \P3_EBX_reg[16]/NET0131  & ~n20654 ;
  assign n20656 = ~\P3_EBX_reg[16]/NET0131  & n20654 ;
  assign n20657 = ~n20655 & ~n20656 ;
  assign n20658 = ~n2946 & ~n20657 ;
  assign n20646 = ~\P3_rEIP_reg[16]/NET0131  & ~n20610 ;
  assign n20647 = \P3_rEIP_reg[16]/NET0131  & n20610 ;
  assign n20648 = ~n20646 & ~n20647 ;
  assign n20659 = n2946 & ~n20648 ;
  assign n20660 = n20473 & ~n20659 ;
  assign n20661 = ~n20658 & n20660 ;
  assign n20645 = \P3_rEIP_reg[16]/NET0131  & n2910 ;
  assign n20649 = n20412 & ~n20648 ;
  assign n20650 = ~\P3_EBX_reg[16]/NET0131  & ~n20412 ;
  assign n20651 = n16094 & ~n20650 ;
  assign n20652 = ~n20649 & n20651 ;
  assign n20662 = ~n20645 & ~n20652 ;
  assign n20663 = ~n20661 & n20662 ;
  assign n20664 = n2453 & ~n20663 ;
  assign n20644 = \P3_rEIP_reg[16]/NET0131  & ~n20409 ;
  assign n20665 = \P3_PhyAddrPointer_reg[16]/NET0131  & n3004 ;
  assign n20666 = ~n4412 & ~n20665 ;
  assign n20667 = ~n20644 & n20666 ;
  assign n20668 = ~n20664 & n20667 ;
  assign n20669 = ~n20643 & n20668 ;
  assign n20671 = ~n13145 & n20636 ;
  assign n20672 = ~n9054 & ~n20671 ;
  assign n20673 = ~\P3_PhyAddrPointer_reg[17]/NET0131  & ~n13144 ;
  assign n20674 = ~n13198 & ~n20673 ;
  assign n20676 = n20672 & ~n20674 ;
  assign n20675 = ~n20672 & n20674 ;
  assign n20677 = ~\P3_DataWidth_reg[1]/NET0131  & ~n20675 ;
  assign n20678 = ~n20676 & n20677 ;
  assign n20670 = \P3_DataWidth_reg[1]/NET0131  & ~\P3_rEIP_reg[17]/NET0131  ;
  assign n20679 = n2959 & ~n20670 ;
  assign n20680 = ~n20678 & n20679 ;
  assign n20688 = ~\P3_rEIP_reg[17]/NET0131  & ~n20647 ;
  assign n20689 = \P3_rEIP_reg[17]/NET0131  & n20647 ;
  assign n20690 = ~n20688 & ~n20689 ;
  assign n20691 = n2946 & ~n20690 ;
  assign n20692 = ~\P3_EBX_reg[17]/NET0131  & ~n2946 ;
  assign n20693 = n2816 & ~n20692 ;
  assign n20694 = ~n20691 & n20693 ;
  assign n20685 = \P3_rEIP_reg[17]/NET0131  & n2815 ;
  assign n20686 = n2786 & ~n2815 ;
  assign n20687 = \P3_EBX_reg[17]/NET0131  & n20686 ;
  assign n20695 = ~n20685 & ~n20687 ;
  assign n20696 = ~n20694 & n20695 ;
  assign n20697 = n2818 & ~n20696 ;
  assign n20682 = ~n2763 & n2818 ;
  assign n20683 = n2910 & ~n20682 ;
  assign n20684 = \P3_rEIP_reg[17]/NET0131  & n20683 ;
  assign n20698 = ~\P3_EBX_reg[15]/NET0131  & ~\P3_EBX_reg[16]/NET0131  ;
  assign n20699 = n20618 & n20698 ;
  assign n20700 = \P3_EBX_reg[31]/NET0131  & ~n20699 ;
  assign n20702 = ~\P3_EBX_reg[17]/NET0131  & n20700 ;
  assign n20701 = \P3_EBX_reg[17]/NET0131  & ~n20700 ;
  assign n20703 = ~n2946 & ~n20701 ;
  assign n20704 = ~n20702 & n20703 ;
  assign n20705 = n20473 & ~n20691 ;
  assign n20706 = ~n20704 & n20705 ;
  assign n20707 = ~n20684 & ~n20706 ;
  assign n20708 = ~n20697 & n20707 ;
  assign n20709 = n2453 & ~n20708 ;
  assign n20681 = \P3_rEIP_reg[17]/NET0131  & ~n20409 ;
  assign n20710 = \P3_PhyAddrPointer_reg[17]/NET0131  & n3004 ;
  assign n20711 = ~n4412 & ~n20710 ;
  assign n20712 = ~n20681 & n20711 ;
  assign n20713 = ~n20709 & n20712 ;
  assign n20714 = ~n20680 & n20713 ;
  assign n20716 = n20671 & ~n20674 ;
  assign n20717 = ~n9054 & ~n20716 ;
  assign n20719 = n13201 & ~n20717 ;
  assign n20718 = ~n13201 & n20717 ;
  assign n20720 = ~\P3_DataWidth_reg[1]/NET0131  & ~n20718 ;
  assign n20721 = ~n20719 & n20720 ;
  assign n20715 = \P3_DataWidth_reg[1]/NET0131  & ~\P3_rEIP_reg[18]/NET0131  ;
  assign n20722 = n2959 & ~n20715 ;
  assign n20723 = ~n20721 & n20722 ;
  assign n20725 = \P3_rEIP_reg[18]/NET0131  & n2910 ;
  assign n20730 = ~\P3_EBX_reg[18]/NET0131  & ~n20412 ;
  assign n20734 = n2818 & ~n20730 ;
  assign n20735 = \P3_EBX_reg[17]/NET0131  & \P3_EBX_reg[31]/NET0131  ;
  assign n20736 = ~n20700 & ~n20735 ;
  assign n20738 = \P3_EBX_reg[18]/NET0131  & n20736 ;
  assign n20737 = ~\P3_EBX_reg[18]/NET0131  & ~n20736 ;
  assign n20739 = ~n2946 & ~n20737 ;
  assign n20740 = ~n20738 & n20739 ;
  assign n20741 = n2821 & ~n20740 ;
  assign n20742 = ~n20734 & ~n20741 ;
  assign n20726 = ~\P3_rEIP_reg[18]/NET0131  & ~n20689 ;
  assign n20727 = \P3_rEIP_reg[17]/NET0131  & \P3_rEIP_reg[18]/NET0131  ;
  assign n20728 = n20647 & n20727 ;
  assign n20729 = ~n20726 & ~n20728 ;
  assign n20731 = n20613 & ~n20730 ;
  assign n20732 = n2946 & ~n20731 ;
  assign n20733 = ~n20729 & n20732 ;
  assign n20743 = ~n2815 & ~n20733 ;
  assign n20744 = ~n20742 & n20743 ;
  assign n20745 = ~n20725 & ~n20744 ;
  assign n20746 = n2453 & ~n20745 ;
  assign n20724 = \P3_rEIP_reg[18]/NET0131  & ~n20409 ;
  assign n20747 = \P3_PhyAddrPointer_reg[18]/NET0131  & n3004 ;
  assign n20748 = ~n4412 & ~n20747 ;
  assign n20749 = ~n20724 & n20748 ;
  assign n20750 = ~n20746 & n20749 ;
  assign n20751 = ~n20723 & n20750 ;
  assign n20753 = ~\P3_PhyAddrPointer_reg[19]/NET0131  & ~n13200 ;
  assign n20754 = ~n12052 & ~n20753 ;
  assign n20755 = ~n9054 & n13201 ;
  assign n20756 = ~n20717 & ~n20755 ;
  assign n20758 = n20754 & n20756 ;
  assign n20757 = ~n20754 & ~n20756 ;
  assign n20759 = ~\P3_DataWidth_reg[1]/NET0131  & ~n20757 ;
  assign n20760 = ~n20758 & n20759 ;
  assign n20752 = \P3_DataWidth_reg[1]/NET0131  & ~\P3_rEIP_reg[19]/NET0131  ;
  assign n20761 = n2959 & ~n20752 ;
  assign n20762 = ~n20760 & n20761 ;
  assign n20764 = \P3_rEIP_reg[19]/NET0131  & n2910 ;
  assign n20768 = ~\P3_EBX_reg[19]/NET0131  & ~n20412 ;
  assign n20772 = n2818 & ~n20768 ;
  assign n20773 = ~\P3_EBX_reg[17]/NET0131  & ~\P3_EBX_reg[18]/NET0131  ;
  assign n20774 = n20699 & n20773 ;
  assign n20775 = \P3_EBX_reg[31]/NET0131  & ~n20774 ;
  assign n20777 = ~\P3_EBX_reg[19]/NET0131  & n20775 ;
  assign n20776 = \P3_EBX_reg[19]/NET0131  & ~n20775 ;
  assign n20778 = ~n2946 & ~n20776 ;
  assign n20779 = ~n20777 & n20778 ;
  assign n20780 = n2821 & ~n20779 ;
  assign n20781 = ~n20772 & ~n20780 ;
  assign n20765 = ~\P3_rEIP_reg[19]/NET0131  & ~n20728 ;
  assign n20766 = \P3_rEIP_reg[19]/NET0131  & n20728 ;
  assign n20767 = ~n20765 & ~n20766 ;
  assign n20769 = n20613 & ~n20768 ;
  assign n20770 = n2946 & ~n20769 ;
  assign n20771 = ~n20767 & n20770 ;
  assign n20782 = ~n2815 & ~n20771 ;
  assign n20783 = ~n20781 & n20782 ;
  assign n20784 = ~n20764 & ~n20783 ;
  assign n20785 = n2453 & ~n20784 ;
  assign n20763 = \P3_rEIP_reg[19]/NET0131  & ~n20409 ;
  assign n20786 = \P3_PhyAddrPointer_reg[19]/NET0131  & n3004 ;
  assign n20787 = ~n4412 & ~n20786 ;
  assign n20788 = ~n20763 & n20787 ;
  assign n20789 = ~n20785 & n20788 ;
  assign n20790 = ~n20762 & n20789 ;
  assign n20792 = \P3_PhyAddrPointer_reg[0]/NET0131  & ~n9054 ;
  assign n20794 = \P3_PhyAddrPointer_reg[1]/NET0131  & n20792 ;
  assign n20793 = ~\P3_PhyAddrPointer_reg[1]/NET0131  & ~n20792 ;
  assign n20795 = ~\P3_DataWidth_reg[1]/NET0131  & ~n20793 ;
  assign n20796 = ~n20794 & n20795 ;
  assign n20791 = \P3_DataWidth_reg[1]/NET0131  & ~\P3_rEIP_reg[1]/NET0131  ;
  assign n20797 = n2959 & ~n20791 ;
  assign n20798 = ~n20796 & n20797 ;
  assign n20802 = \P3_rEIP_reg[1]/NET0131  & n2910 ;
  assign n20810 = ~n14957 & ~n20429 ;
  assign n20811 = \P3_EBX_reg[31]/NET0131  & ~n20810 ;
  assign n20809 = ~\P3_EBX_reg[1]/NET0131  & ~\P3_EBX_reg[31]/NET0131  ;
  assign n20812 = ~n2946 & ~n20809 ;
  assign n20813 = ~n20811 & n20812 ;
  assign n20805 = ~\P3_DataWidth_reg[1]/NET0131  & ~\P3_rEIP_reg[1]/NET0131  ;
  assign n20814 = ~n2835 & n20805 ;
  assign n20815 = ~n20813 & ~n20814 ;
  assign n20816 = n2821 & ~n20815 ;
  assign n20803 = n2763 & n2920 ;
  assign n20804 = \P3_EBX_reg[1]/NET0131  & ~n20412 ;
  assign n20806 = n2874 & n20805 ;
  assign n20807 = ~n20804 & ~n20806 ;
  assign n20808 = n2818 & ~n20807 ;
  assign n20817 = ~n20803 & ~n20808 ;
  assign n20818 = ~n20816 & n20817 ;
  assign n20819 = ~n2815 & ~n20818 ;
  assign n20820 = ~n20802 & ~n20819 ;
  assign n20821 = n2453 & ~n20820 ;
  assign n20799 = \P3_PhyAddrPointer_reg[1]/NET0131  & n3004 ;
  assign n20800 = ~n4415 & n16197 ;
  assign n20801 = \P3_rEIP_reg[1]/NET0131  & ~n20800 ;
  assign n20822 = ~n20799 & ~n20801 ;
  assign n20823 = ~n20821 & n20822 ;
  assign n20824 = ~n20798 & n20823 ;
  assign n20826 = ~n13201 & ~n20754 ;
  assign n20827 = n20716 & n20826 ;
  assign n20828 = ~n9054 & ~n20827 ;
  assign n20830 = ~n12055 & n20828 ;
  assign n20829 = n12055 & ~n20828 ;
  assign n20831 = ~\P3_DataWidth_reg[1]/NET0131  & ~n20829 ;
  assign n20832 = ~n20830 & n20831 ;
  assign n20825 = \P3_DataWidth_reg[1]/NET0131  & ~\P3_rEIP_reg[20]/NET0131  ;
  assign n20833 = n2959 & ~n20825 ;
  assign n20834 = ~n20832 & n20833 ;
  assign n20840 = ~\P3_rEIP_reg[20]/NET0131  & ~n20766 ;
  assign n20841 = \P3_rEIP_reg[19]/NET0131  & n20727 ;
  assign n20842 = \P3_rEIP_reg[20]/NET0131  & n20841 ;
  assign n20843 = n20647 & n20842 ;
  assign n20844 = ~n20840 & ~n20843 ;
  assign n20845 = n2946 & ~n20844 ;
  assign n20846 = ~\P3_EBX_reg[20]/NET0131  & ~n2946 ;
  assign n20847 = n2816 & ~n20846 ;
  assign n20848 = ~n20845 & n20847 ;
  assign n20838 = \P3_rEIP_reg[20]/NET0131  & n2815 ;
  assign n20839 = \P3_EBX_reg[20]/NET0131  & n20686 ;
  assign n20849 = ~n20838 & ~n20839 ;
  assign n20850 = ~n20848 & n20849 ;
  assign n20851 = n2818 & ~n20850 ;
  assign n20837 = \P3_rEIP_reg[20]/NET0131  & n20683 ;
  assign n20852 = ~\P3_EBX_reg[19]/NET0131  & n20774 ;
  assign n20853 = \P3_EBX_reg[31]/NET0131  & ~n20852 ;
  assign n20855 = ~\P3_EBX_reg[20]/NET0131  & n20853 ;
  assign n20854 = \P3_EBX_reg[20]/NET0131  & ~n20853 ;
  assign n20856 = ~n2946 & ~n20854 ;
  assign n20857 = ~n20855 & n20856 ;
  assign n20858 = n20473 & ~n20845 ;
  assign n20859 = ~n20857 & n20858 ;
  assign n20860 = ~n20837 & ~n20859 ;
  assign n20861 = ~n20851 & n20860 ;
  assign n20862 = n2453 & ~n20861 ;
  assign n20835 = \P3_PhyAddrPointer_reg[20]/NET0131  & n3004 ;
  assign n20836 = \P3_rEIP_reg[20]/NET0131  & ~n20800 ;
  assign n20863 = ~n20835 & ~n20836 ;
  assign n20864 = ~n20862 & n20863 ;
  assign n20865 = ~n20834 & n20864 ;
  assign n20867 = ~n9054 & n12055 ;
  assign n20868 = ~n20828 & ~n20867 ;
  assign n20870 = n13218 & n20868 ;
  assign n20869 = ~n13218 & ~n20868 ;
  assign n20871 = ~\P3_DataWidth_reg[1]/NET0131  & ~n20869 ;
  assign n20872 = ~n20870 & n20871 ;
  assign n20866 = \P3_DataWidth_reg[1]/NET0131  & ~\P3_rEIP_reg[21]/NET0131  ;
  assign n20873 = n2959 & ~n20866 ;
  assign n20874 = ~n20872 & n20873 ;
  assign n20886 = ~\P3_EBX_reg[19]/NET0131  & ~\P3_EBX_reg[20]/NET0131  ;
  assign n20887 = n20774 & n20886 ;
  assign n20888 = \P3_EBX_reg[31]/NET0131  & ~n20887 ;
  assign n20889 = ~\P3_EBX_reg[21]/NET0131  & ~n20888 ;
  assign n20890 = \P3_EBX_reg[21]/NET0131  & n20888 ;
  assign n20891 = ~n20889 & ~n20890 ;
  assign n20892 = ~n2946 & ~n20891 ;
  assign n20878 = ~\P3_rEIP_reg[21]/NET0131  & ~n20843 ;
  assign n20879 = \P3_rEIP_reg[21]/NET0131  & n20843 ;
  assign n20880 = ~n20878 & ~n20879 ;
  assign n20885 = n2946 & ~n20880 ;
  assign n20893 = n20473 & ~n20885 ;
  assign n20894 = ~n20892 & n20893 ;
  assign n20877 = \P3_rEIP_reg[21]/NET0131  & n2910 ;
  assign n20881 = n20412 & ~n20880 ;
  assign n20882 = ~\P3_EBX_reg[21]/NET0131  & ~n20412 ;
  assign n20883 = n16094 & ~n20882 ;
  assign n20884 = ~n20881 & n20883 ;
  assign n20895 = ~n20877 & ~n20884 ;
  assign n20896 = ~n20894 & n20895 ;
  assign n20897 = n2453 & ~n20896 ;
  assign n20875 = \P3_PhyAddrPointer_reg[21]/NET0131  & n3004 ;
  assign n20876 = \P3_rEIP_reg[21]/NET0131  & ~n20800 ;
  assign n20898 = ~n20875 & ~n20876 ;
  assign n20899 = ~n20897 & n20898 ;
  assign n20900 = ~n20874 & n20899 ;
  assign n20926 = ~n12055 & ~n13218 ;
  assign n20927 = n20827 & n20926 ;
  assign n20928 = ~n9054 & ~n20927 ;
  assign n20930 = ~n12075 & n20928 ;
  assign n20929 = n12075 & ~n20928 ;
  assign n20931 = ~\P3_DataWidth_reg[1]/NET0131  & ~n20929 ;
  assign n20932 = ~n20930 & n20931 ;
  assign n20925 = \P3_DataWidth_reg[1]/NET0131  & ~\P3_rEIP_reg[22]/NET0131  ;
  assign n20933 = n2959 & ~n20925 ;
  assign n20934 = ~n20932 & n20933 ;
  assign n20903 = \P3_rEIP_reg[22]/NET0131  & n2910 ;
  assign n20908 = ~\P3_EBX_reg[22]/NET0131  & ~n20412 ;
  assign n20912 = n2818 & ~n20908 ;
  assign n20913 = ~\P3_EBX_reg[21]/NET0131  & n20887 ;
  assign n20914 = \P3_EBX_reg[31]/NET0131  & ~n20913 ;
  assign n20916 = ~\P3_EBX_reg[22]/NET0131  & n20914 ;
  assign n20915 = \P3_EBX_reg[22]/NET0131  & ~n20914 ;
  assign n20917 = ~n2946 & ~n20915 ;
  assign n20918 = ~n20916 & n20917 ;
  assign n20919 = n2821 & ~n20918 ;
  assign n20920 = ~n20912 & ~n20919 ;
  assign n20904 = ~\P3_rEIP_reg[22]/NET0131  & ~n20879 ;
  assign n20905 = \P3_rEIP_reg[21]/NET0131  & \P3_rEIP_reg[22]/NET0131  ;
  assign n20906 = n20843 & n20905 ;
  assign n20907 = ~n20904 & ~n20906 ;
  assign n20909 = n20613 & ~n20908 ;
  assign n20910 = n2946 & ~n20909 ;
  assign n20911 = ~n20907 & n20910 ;
  assign n20921 = ~n2815 & ~n20911 ;
  assign n20922 = ~n20920 & n20921 ;
  assign n20923 = ~n20903 & ~n20922 ;
  assign n20924 = n2453 & ~n20923 ;
  assign n20901 = \P3_rEIP_reg[22]/NET0131  & ~n20800 ;
  assign n20902 = \P3_PhyAddrPointer_reg[22]/NET0131  & n3004 ;
  assign n20935 = ~n20901 & ~n20902 ;
  assign n20936 = ~n20924 & n20935 ;
  assign n20937 = ~n20934 & n20936 ;
  assign n20960 = ~n12075 & n20927 ;
  assign n20961 = ~n9054 & ~n20960 ;
  assign n20963 = ~n11122 & n20961 ;
  assign n20962 = n11122 & ~n20961 ;
  assign n20964 = ~\P3_DataWidth_reg[1]/NET0131  & ~n20962 ;
  assign n20965 = ~n20963 & n20964 ;
  assign n20959 = \P3_DataWidth_reg[1]/NET0131  & ~\P3_rEIP_reg[23]/NET0131  ;
  assign n20966 = n2959 & ~n20959 ;
  assign n20967 = ~n20965 & n20966 ;
  assign n20938 = \P3_rEIP_reg[23]/NET0131  & n2910 ;
  assign n20940 = ~\P3_rEIP_reg[23]/NET0131  & ~n20906 ;
  assign n20941 = \P3_rEIP_reg[23]/NET0131  & n20906 ;
  assign n20942 = ~n20940 & ~n20941 ;
  assign n20943 = n20412 & ~n20942 ;
  assign n20939 = ~\P3_EBX_reg[23]/NET0131  & ~n20412 ;
  assign n20944 = n2818 & ~n20939 ;
  assign n20945 = ~n20943 & n20944 ;
  assign n20947 = ~\P3_EBX_reg[22]/NET0131  & n20913 ;
  assign n20948 = \P3_EBX_reg[31]/NET0131  & ~n20947 ;
  assign n20950 = ~\P3_EBX_reg[23]/NET0131  & n20948 ;
  assign n20949 = \P3_EBX_reg[23]/NET0131  & ~n20948 ;
  assign n20951 = ~n2946 & ~n20949 ;
  assign n20952 = ~n20950 & n20951 ;
  assign n20946 = n2946 & ~n20942 ;
  assign n20953 = n2821 & ~n20946 ;
  assign n20954 = ~n20952 & n20953 ;
  assign n20955 = ~n20945 & ~n20954 ;
  assign n20956 = ~n2815 & ~n20955 ;
  assign n20957 = ~n20938 & ~n20956 ;
  assign n20958 = n2453 & ~n20957 ;
  assign n20968 = \P3_rEIP_reg[23]/NET0131  & ~n20800 ;
  assign n20969 = \P3_PhyAddrPointer_reg[23]/NET0131  & n3004 ;
  assign n20970 = ~n20968 & ~n20969 ;
  assign n20971 = ~n20958 & n20970 ;
  assign n20972 = ~n20967 & n20971 ;
  assign n21001 = ~n11122 & ~n12075 ;
  assign n21002 = n20927 & n21001 ;
  assign n21003 = ~n9054 & ~n21002 ;
  assign n21005 = ~n12107 & n21003 ;
  assign n21004 = n12107 & ~n21003 ;
  assign n21006 = ~\P3_DataWidth_reg[1]/NET0131  & ~n21004 ;
  assign n21007 = ~n21005 & n21006 ;
  assign n21000 = \P3_DataWidth_reg[1]/NET0131  & ~\P3_rEIP_reg[24]/NET0131  ;
  assign n21008 = n2959 & ~n21000 ;
  assign n21009 = ~n21007 & n21008 ;
  assign n20988 = ~\P3_EBX_reg[22]/NET0131  & ~\P3_EBX_reg[23]/NET0131  ;
  assign n20989 = n20913 & n20988 ;
  assign n20990 = \P3_EBX_reg[31]/NET0131  & ~n20989 ;
  assign n20992 = ~\P3_EBX_reg[24]/NET0131  & n20990 ;
  assign n20991 = \P3_EBX_reg[24]/NET0131  & ~n20990 ;
  assign n20993 = ~n2946 & ~n20991 ;
  assign n20994 = ~n20992 & n20993 ;
  assign n20977 = ~\P3_rEIP_reg[24]/NET0131  & ~n20941 ;
  assign n20978 = \P3_rEIP_reg[24]/NET0131  & n20941 ;
  assign n20979 = ~n20977 & ~n20978 ;
  assign n20980 = n2946 & ~n20979 ;
  assign n20995 = n20473 & ~n20980 ;
  assign n20996 = ~n20994 & n20995 ;
  assign n20981 = ~\P3_EBX_reg[24]/NET0131  & ~n2946 ;
  assign n20982 = n2816 & ~n20981 ;
  assign n20983 = ~n20980 & n20982 ;
  assign n20975 = \P3_rEIP_reg[24]/NET0131  & n2815 ;
  assign n20976 = \P3_EBX_reg[24]/NET0131  & n20686 ;
  assign n20984 = ~n20975 & ~n20976 ;
  assign n20985 = ~n20983 & n20984 ;
  assign n20986 = n2818 & ~n20985 ;
  assign n20987 = \P3_rEIP_reg[24]/NET0131  & n20683 ;
  assign n20997 = ~n20986 & ~n20987 ;
  assign n20998 = ~n20996 & n20997 ;
  assign n20999 = n2453 & ~n20998 ;
  assign n20973 = \P3_rEIP_reg[24]/NET0131  & ~n20800 ;
  assign n20974 = \P3_PhyAddrPointer_reg[24]/NET0131  & n3004 ;
  assign n21010 = ~n20973 & ~n20974 ;
  assign n21011 = ~n20999 & n21010 ;
  assign n21012 = ~n21009 & n21011 ;
  assign n21014 = ~n9054 & n12107 ;
  assign n21015 = ~n21003 & ~n21014 ;
  assign n21017 = ~n13242 & ~n21015 ;
  assign n21016 = n13242 & n21015 ;
  assign n21018 = ~\P3_DataWidth_reg[1]/NET0131  & ~n21016 ;
  assign n21019 = ~n21017 & n21018 ;
  assign n21013 = \P3_DataWidth_reg[1]/NET0131  & ~\P3_rEIP_reg[25]/NET0131  ;
  assign n21020 = n2959 & ~n21013 ;
  assign n21021 = ~n21019 & n21020 ;
  assign n21025 = ~\P3_rEIP_reg[25]/NET0131  & ~n20978 ;
  assign n21026 = \P3_rEIP_reg[23]/NET0131  & \P3_rEIP_reg[24]/NET0131  ;
  assign n21027 = \P3_rEIP_reg[25]/NET0131  & n21026 ;
  assign n21028 = n20906 & n21027 ;
  assign n21029 = ~n21025 & ~n21028 ;
  assign n21030 = n2946 & ~n21029 ;
  assign n21031 = ~\P3_EBX_reg[25]/NET0131  & ~n2946 ;
  assign n21032 = n2816 & ~n21031 ;
  assign n21033 = ~n21030 & n21032 ;
  assign n21034 = \P3_rEIP_reg[25]/NET0131  & n2815 ;
  assign n21035 = \P3_EBX_reg[25]/NET0131  & n20686 ;
  assign n21036 = ~n21034 & ~n21035 ;
  assign n21037 = ~n21033 & n21036 ;
  assign n21038 = n2818 & ~n21037 ;
  assign n21024 = \P3_rEIP_reg[25]/NET0131  & n20683 ;
  assign n21039 = ~\P3_EBX_reg[24]/NET0131  & n20988 ;
  assign n21040 = n20913 & n21039 ;
  assign n21041 = \P3_EBX_reg[31]/NET0131  & ~n21040 ;
  assign n21043 = ~\P3_EBX_reg[25]/NET0131  & n21041 ;
  assign n21042 = \P3_EBX_reg[25]/NET0131  & ~n21041 ;
  assign n21044 = ~n2946 & ~n21042 ;
  assign n21045 = ~n21043 & n21044 ;
  assign n21046 = n20473 & ~n21030 ;
  assign n21047 = ~n21045 & n21046 ;
  assign n21048 = ~n21024 & ~n21047 ;
  assign n21049 = ~n21038 & n21048 ;
  assign n21050 = n2453 & ~n21049 ;
  assign n21022 = \P3_rEIP_reg[25]/NET0131  & ~n20800 ;
  assign n21023 = \P3_PhyAddrPointer_reg[25]/NET0131  & n3004 ;
  assign n21051 = ~n21022 & ~n21023 ;
  assign n21052 = ~n21050 & n21051 ;
  assign n21053 = ~n21021 & n21052 ;
  assign n21075 = ~n12107 & ~n13242 ;
  assign n21076 = n21002 & n21075 ;
  assign n21077 = ~n9054 & ~n21076 ;
  assign n21079 = ~n12144 & n21077 ;
  assign n21078 = n12144 & ~n21077 ;
  assign n21080 = ~\P3_DataWidth_reg[1]/NET0131  & ~n21078 ;
  assign n21081 = ~n21079 & n21080 ;
  assign n21074 = \P3_DataWidth_reg[1]/NET0131  & ~\P3_rEIP_reg[26]/NET0131  ;
  assign n21082 = n2959 & ~n21074 ;
  assign n21083 = ~n21081 & n21082 ;
  assign n21063 = ~\P3_EBX_reg[25]/NET0131  & n21040 ;
  assign n21064 = \P3_EBX_reg[31]/NET0131  & ~n21063 ;
  assign n21065 = ~\P3_EBX_reg[26]/NET0131  & ~n21064 ;
  assign n21066 = \P3_EBX_reg[26]/NET0131  & n21064 ;
  assign n21067 = ~n21065 & ~n21066 ;
  assign n21068 = ~n2946 & ~n21067 ;
  assign n21055 = \P3_rEIP_reg[26]/NET0131  & n21028 ;
  assign n21056 = ~\P3_rEIP_reg[26]/NET0131  & ~n21028 ;
  assign n21057 = ~n21055 & ~n21056 ;
  assign n21062 = n2946 & ~n21057 ;
  assign n21069 = n20473 & ~n21062 ;
  assign n21070 = ~n21068 & n21069 ;
  assign n21054 = \P3_rEIP_reg[26]/NET0131  & n2910 ;
  assign n21058 = n20412 & ~n21057 ;
  assign n21059 = ~\P3_EBX_reg[26]/NET0131  & ~n20412 ;
  assign n21060 = n16094 & ~n21059 ;
  assign n21061 = ~n21058 & n21060 ;
  assign n21071 = ~n21054 & ~n21061 ;
  assign n21072 = ~n21070 & n21071 ;
  assign n21073 = n2453 & ~n21072 ;
  assign n21084 = \P3_PhyAddrPointer_reg[26]/NET0131  & n3004 ;
  assign n21085 = \P3_rEIP_reg[26]/NET0131  & ~n20800 ;
  assign n21086 = ~n21084 & ~n21085 ;
  assign n21087 = ~n21073 & n21086 ;
  assign n21088 = ~n21083 & n21087 ;
  assign n21116 = ~n12144 & n21076 ;
  assign n21117 = ~n9054 & ~n21116 ;
  assign n21119 = ~n11166 & n21117 ;
  assign n21118 = n11166 & ~n21117 ;
  assign n21120 = ~\P3_DataWidth_reg[1]/NET0131  & ~n21118 ;
  assign n21121 = ~n21119 & n21120 ;
  assign n21115 = \P3_DataWidth_reg[1]/NET0131  & ~\P3_rEIP_reg[27]/NET0131  ;
  assign n21122 = n2959 & ~n21115 ;
  assign n21123 = ~n21121 & n21122 ;
  assign n21094 = ~\P3_EBX_reg[26]/NET0131  & n21063 ;
  assign n21095 = \P3_EBX_reg[31]/NET0131  & ~n21094 ;
  assign n21097 = ~\P3_EBX_reg[27]/NET0131  & n21095 ;
  assign n21096 = \P3_EBX_reg[27]/NET0131  & ~n21095 ;
  assign n21098 = ~n2946 & ~n21096 ;
  assign n21099 = ~n21097 & n21098 ;
  assign n21089 = ~\P3_rEIP_reg[27]/NET0131  & ~n21055 ;
  assign n21090 = \P3_rEIP_reg[26]/NET0131  & \P3_rEIP_reg[27]/NET0131  ;
  assign n21091 = n21028 & n21090 ;
  assign n21092 = ~n21089 & ~n21091 ;
  assign n21093 = n2946 & ~n21092 ;
  assign n21100 = n20473 & ~n21093 ;
  assign n21101 = ~n21099 & n21100 ;
  assign n21102 = \P3_rEIP_reg[27]/NET0131  & n20683 ;
  assign n21104 = n20412 & n21092 ;
  assign n21105 = \P3_EBX_reg[27]/NET0131  & ~n20412 ;
  assign n21106 = ~n2815 & ~n21105 ;
  assign n21107 = ~n21104 & n21106 ;
  assign n21103 = ~\P3_rEIP_reg[27]/NET0131  & n2815 ;
  assign n21108 = n2818 & ~n21103 ;
  assign n21109 = ~n21107 & n21108 ;
  assign n21110 = ~n21102 & ~n21109 ;
  assign n21111 = ~n21101 & n21110 ;
  assign n21112 = n2453 & ~n21111 ;
  assign n21113 = \P3_PhyAddrPointer_reg[27]/NET0131  & n3004 ;
  assign n21114 = \P3_rEIP_reg[27]/NET0131  & ~n20800 ;
  assign n21124 = ~n21113 & ~n21114 ;
  assign n21125 = ~n21112 & n21124 ;
  assign n21126 = ~n21123 & n21125 ;
  assign n21131 = ~\P3_EBX_reg[27]/NET0131  & n21094 ;
  assign n21132 = \P3_EBX_reg[31]/NET0131  & ~n21131 ;
  assign n21134 = \P3_EBX_reg[28]/NET0131  & ~n21132 ;
  assign n21133 = ~\P3_EBX_reg[28]/NET0131  & n21132 ;
  assign n21135 = ~n2946 & ~n21133 ;
  assign n21136 = ~n21134 & n21135 ;
  assign n21127 = ~\P3_rEIP_reg[28]/NET0131  & ~n21091 ;
  assign n21128 = \P3_rEIP_reg[28]/NET0131  & n21091 ;
  assign n21129 = ~n21127 & ~n21128 ;
  assign n21130 = n2946 & ~n21129 ;
  assign n21137 = n20473 & ~n21130 ;
  assign n21138 = ~n21136 & n21137 ;
  assign n21140 = n20412 & n21129 ;
  assign n21139 = \P3_EBX_reg[28]/NET0131  & ~n20412 ;
  assign n21141 = ~n2815 & ~n21139 ;
  assign n21142 = ~n21140 & n21141 ;
  assign n21143 = n2818 & ~n21142 ;
  assign n21144 = ~n20683 & ~n21143 ;
  assign n21145 = \P3_rEIP_reg[28]/NET0131  & ~n21144 ;
  assign n21146 = ~n2815 & n21143 ;
  assign n21147 = ~n21145 & ~n21146 ;
  assign n21148 = ~n21138 & n21147 ;
  assign n21149 = n2453 & ~n21148 ;
  assign n21151 = ~n11166 & ~n12144 ;
  assign n21152 = n21076 & n21151 ;
  assign n21153 = ~n9054 & ~n21152 ;
  assign n21155 = ~n11185 & n21153 ;
  assign n21154 = n11185 & ~n21153 ;
  assign n21156 = ~\P3_DataWidth_reg[1]/NET0131  & ~n21154 ;
  assign n21157 = ~n21155 & n21156 ;
  assign n21150 = \P3_DataWidth_reg[1]/NET0131  & ~\P3_rEIP_reg[28]/NET0131  ;
  assign n21158 = n2959 & ~n21150 ;
  assign n21159 = ~n21157 & n21158 ;
  assign n21160 = \P3_PhyAddrPointer_reg[28]/NET0131  & n3004 ;
  assign n21161 = \P3_rEIP_reg[28]/NET0131  & ~n20800 ;
  assign n21162 = ~n21160 & ~n21161 ;
  assign n21163 = ~n21159 & n21162 ;
  assign n21164 = ~n21149 & n21163 ;
  assign n21171 = ~\P3_EBX_reg[27]/NET0131  & ~\P3_EBX_reg[28]/NET0131  ;
  assign n21172 = n21094 & n21171 ;
  assign n21173 = \P3_EBX_reg[31]/NET0131  & ~n21172 ;
  assign n21175 = ~\P3_EBX_reg[29]/NET0131  & n21173 ;
  assign n21174 = \P3_EBX_reg[29]/NET0131  & ~n21173 ;
  assign n21176 = ~n2946 & ~n21174 ;
  assign n21177 = ~n21175 & n21176 ;
  assign n21165 = ~\P3_rEIP_reg[29]/NET0131  & ~n21128 ;
  assign n21166 = \P3_rEIP_reg[28]/NET0131  & n21090 ;
  assign n21167 = \P3_rEIP_reg[29]/NET0131  & n21166 ;
  assign n21168 = n21028 & n21167 ;
  assign n21169 = ~n21165 & ~n21168 ;
  assign n21170 = n2946 & ~n21169 ;
  assign n21178 = n20473 & ~n21170 ;
  assign n21179 = ~n21177 & n21178 ;
  assign n21180 = \P3_rEIP_reg[29]/NET0131  & n20683 ;
  assign n21182 = n20412 & n21169 ;
  assign n21183 = \P3_EBX_reg[29]/NET0131  & ~n20412 ;
  assign n21184 = ~n2815 & ~n21183 ;
  assign n21185 = ~n21182 & n21184 ;
  assign n21181 = ~\P3_rEIP_reg[29]/NET0131  & n2815 ;
  assign n21186 = n2818 & ~n21181 ;
  assign n21187 = ~n21185 & n21186 ;
  assign n21188 = ~n21180 & ~n21187 ;
  assign n21189 = ~n21179 & n21188 ;
  assign n21190 = n2453 & ~n21189 ;
  assign n21192 = ~n11185 & n21151 ;
  assign n21193 = n21076 & n21192 ;
  assign n21194 = ~n9054 & ~n21193 ;
  assign n21196 = ~n11225 & n21194 ;
  assign n21195 = n11225 & ~n21194 ;
  assign n21197 = ~\P3_DataWidth_reg[1]/NET0131  & ~n21195 ;
  assign n21198 = ~n21196 & n21197 ;
  assign n21191 = \P3_DataWidth_reg[1]/NET0131  & ~\P3_rEIP_reg[29]/NET0131  ;
  assign n21199 = n2959 & ~n21191 ;
  assign n21200 = ~n21198 & n21199 ;
  assign n21201 = \P3_rEIP_reg[29]/NET0131  & ~n20800 ;
  assign n21202 = \P3_PhyAddrPointer_reg[29]/NET0131  & n3004 ;
  assign n21203 = ~n21201 & ~n21202 ;
  assign n21204 = ~n21200 & n21203 ;
  assign n21205 = ~n21190 & n21204 ;
  assign n21207 = ~\P3_PhyAddrPointer_reg[0]/NET0131  & \P3_PhyAddrPointer_reg[1]/NET0131  ;
  assign n21208 = ~n9054 & ~n21207 ;
  assign n21209 = ~\P3_PhyAddrPointer_reg[1]/NET0131  & ~\P3_PhyAddrPointer_reg[2]/NET0131  ;
  assign n21210 = ~n15803 & ~n21209 ;
  assign n21212 = ~n21208 & n21210 ;
  assign n21211 = n21208 & ~n21210 ;
  assign n21213 = ~\P3_DataWidth_reg[1]/NET0131  & ~n21211 ;
  assign n21214 = ~n21212 & n21213 ;
  assign n21206 = \P3_DataWidth_reg[1]/NET0131  & ~\P3_rEIP_reg[2]/NET0131  ;
  assign n21215 = n2959 & ~n21206 ;
  assign n21216 = ~n21214 & n21215 ;
  assign n21219 = \P3_rEIP_reg[2]/NET0131  & n2910 ;
  assign n21222 = ~\P3_rEIP_reg[1]/NET0131  & ~\P3_rEIP_reg[2]/NET0131  ;
  assign n21223 = ~\P3_DataWidth_reg[1]/NET0131  & ~n20414 ;
  assign n21224 = ~n21222 & n21223 ;
  assign n21228 = ~n2835 & n21224 ;
  assign n21229 = \P3_EBX_reg[31]/NET0131  & ~n20429 ;
  assign n21231 = \P3_EBX_reg[2]/NET0131  & n21229 ;
  assign n21230 = ~\P3_EBX_reg[2]/NET0131  & ~n21229 ;
  assign n21232 = ~n2946 & ~n21230 ;
  assign n21233 = ~n21231 & n21232 ;
  assign n21234 = ~n21228 & ~n21233 ;
  assign n21235 = n2821 & ~n21234 ;
  assign n21220 = n2763 & n2780 ;
  assign n21221 = \P3_EBX_reg[2]/NET0131  & ~n20412 ;
  assign n21225 = n2874 & n21224 ;
  assign n21226 = ~n21221 & ~n21225 ;
  assign n21227 = n2818 & ~n21226 ;
  assign n21236 = ~n21220 & ~n21227 ;
  assign n21237 = ~n21235 & n21236 ;
  assign n21238 = ~n2815 & ~n21237 ;
  assign n21239 = ~n21219 & ~n21238 ;
  assign n21240 = n2453 & ~n21239 ;
  assign n21217 = \P3_PhyAddrPointer_reg[2]/NET0131  & n3004 ;
  assign n21218 = \P3_rEIP_reg[2]/NET0131  & ~n20800 ;
  assign n21241 = ~n21217 & ~n21218 ;
  assign n21242 = ~n21240 & n21241 ;
  assign n21243 = ~n21216 & n21242 ;
  assign n21244 = \P3_EBX_reg[31]/NET0131  & ~n2946 ;
  assign n21245 = ~\P3_EBX_reg[29]/NET0131  & ~\P3_EBX_reg[30]/NET0131  ;
  assign n21246 = n21244 & n21245 ;
  assign n21247 = n21172 & n21246 ;
  assign n21248 = \P3_rEIP_reg[30]/NET0131  & n21168 ;
  assign n21250 = \P3_rEIP_reg[31]/NET0131  & n21248 ;
  assign n21249 = ~\P3_rEIP_reg[31]/NET0131  & ~n21248 ;
  assign n21251 = n2946 & ~n21249 ;
  assign n21252 = ~n21250 & n21251 ;
  assign n21253 = ~n21247 & ~n21252 ;
  assign n21254 = n2821 & ~n21253 ;
  assign n21255 = ~n21244 & ~n21252 ;
  assign n21256 = ~n2786 & n2818 ;
  assign n21257 = ~n21255 & n21256 ;
  assign n21258 = ~n21254 & ~n21257 ;
  assign n21259 = ~n2815 & ~n21258 ;
  assign n21260 = \P3_rEIP_reg[31]/NET0131  & n2910 ;
  assign n21261 = ~n2815 & n20613 ;
  assign n21262 = \P3_EBX_reg[31]/NET0131  & n21261 ;
  assign n21263 = ~n21260 & ~n21262 ;
  assign n21264 = ~n21259 & n21263 ;
  assign n21265 = n2453 & ~n21264 ;
  assign n21268 = \P3_DataWidth_reg[1]/NET0131  & \P3_rEIP_reg[31]/NET0131  ;
  assign n21269 = ~n11166 & ~n11185 ;
  assign n21270 = ~n10073 & n21269 ;
  assign n21271 = ~n11225 & n21270 ;
  assign n21272 = n21116 & n21271 ;
  assign n21273 = n9056 & n21272 ;
  assign n21274 = ~n21268 & ~n21273 ;
  assign n21275 = n2959 & ~n21274 ;
  assign n21266 = \P3_PhyAddrPointer_reg[31]/NET0131  & n3004 ;
  assign n21267 = \P3_rEIP_reg[31]/NET0131  & ~n20800 ;
  assign n21276 = ~n21266 & ~n21267 ;
  assign n21277 = ~n21275 & n21276 ;
  assign n21278 = ~n21265 & n21277 ;
  assign n21280 = \P3_PhyAddrPointer_reg[2]/NET0131  & n21207 ;
  assign n21281 = ~n9054 & ~n21280 ;
  assign n21283 = n16200 & ~n21281 ;
  assign n21282 = ~n16200 & n21281 ;
  assign n21284 = ~\P3_DataWidth_reg[1]/NET0131  & ~n21282 ;
  assign n21285 = ~n21283 & n21284 ;
  assign n21279 = \P3_DataWidth_reg[1]/NET0131  & ~\P3_rEIP_reg[3]/NET0131  ;
  assign n21286 = n2959 & ~n21279 ;
  assign n21287 = ~n21285 & n21286 ;
  assign n21289 = \P3_rEIP_reg[3]/NET0131  & n2910 ;
  assign n21302 = \P3_EBX_reg[3]/NET0131  & ~n20412 ;
  assign n21296 = ~\P3_rEIP_reg[3]/NET0131  & ~n20414 ;
  assign n21297 = ~\P3_DataWidth_reg[1]/NET0131  & ~n20415 ;
  assign n21298 = ~n21296 & n21297 ;
  assign n21303 = n2874 & n21298 ;
  assign n21304 = ~n21302 & ~n21303 ;
  assign n21305 = n2818 & ~n21304 ;
  assign n21290 = n2763 & ~n2872 ;
  assign n21291 = \P3_EBX_reg[31]/NET0131  & ~n20430 ;
  assign n21293 = \P3_EBX_reg[3]/NET0131  & n21291 ;
  assign n21292 = ~\P3_EBX_reg[3]/NET0131  & ~n21291 ;
  assign n21294 = ~n2946 & ~n21292 ;
  assign n21295 = ~n21293 & n21294 ;
  assign n21299 = ~n2835 & n21298 ;
  assign n21300 = ~n21295 & ~n21299 ;
  assign n21301 = n2821 & ~n21300 ;
  assign n21306 = ~n21290 & ~n21301 ;
  assign n21307 = ~n21305 & n21306 ;
  assign n21308 = ~n2815 & ~n21307 ;
  assign n21309 = ~n21289 & ~n21308 ;
  assign n21310 = n2453 & ~n21309 ;
  assign n21288 = \P3_rEIP_reg[3]/NET0131  & ~n20800 ;
  assign n21311 = ~n16202 & ~n21288 ;
  assign n21312 = ~n21310 & n21311 ;
  assign n21313 = ~n21287 & n21312 ;
  assign n21315 = ~n9054 & ~n15804 ;
  assign n21316 = ~n20792 & ~n21315 ;
  assign n21318 = ~n15807 & ~n21316 ;
  assign n21317 = n15807 & n21316 ;
  assign n21319 = ~\P3_DataWidth_reg[1]/NET0131  & ~n21317 ;
  assign n21320 = ~n21318 & n21319 ;
  assign n21314 = \P3_DataWidth_reg[1]/NET0131  & ~\P3_rEIP_reg[4]/NET0131  ;
  assign n21321 = n2959 & ~n21314 ;
  assign n21322 = ~n21320 & n21321 ;
  assign n21330 = \P3_EBX_reg[31]/NET0131  & ~n20431 ;
  assign n21333 = ~n21256 & n21330 ;
  assign n21334 = \P3_EBX_reg[4]/NET0131  & ~n21333 ;
  assign n21331 = ~\P3_EBX_reg[4]/NET0131  & n21330 ;
  assign n21332 = n2821 & n21331 ;
  assign n21335 = ~n2946 & ~n21332 ;
  assign n21336 = ~n21334 & n21335 ;
  assign n21326 = ~n2821 & ~n21256 ;
  assign n21327 = ~\P3_rEIP_reg[4]/NET0131  & ~n20415 ;
  assign n21328 = ~n20416 & ~n21327 ;
  assign n21329 = n2946 & ~n21328 ;
  assign n21337 = ~n2815 & ~n21329 ;
  assign n21338 = ~n21326 & n21337 ;
  assign n21339 = ~n21336 & n21338 ;
  assign n21324 = \P3_EBX_reg[4]/NET0131  & n21261 ;
  assign n21325 = \P3_rEIP_reg[4]/NET0131  & n2910 ;
  assign n21340 = ~n21324 & ~n21325 ;
  assign n21341 = ~n21339 & n21340 ;
  assign n21342 = n2453 & ~n21341 ;
  assign n21323 = \P3_rEIP_reg[4]/NET0131  & ~n20409 ;
  assign n21343 = \P3_PhyAddrPointer_reg[4]/NET0131  & n3004 ;
  assign n21344 = ~n4412 & ~n21343 ;
  assign n21345 = ~n21323 & n21344 ;
  assign n21346 = ~n21342 & n21345 ;
  assign n21347 = ~n21322 & n21346 ;
  assign n21349 = ~\P3_PhyAddrPointer_reg[0]/NET0131  & n13248 ;
  assign n21350 = ~n9054 & ~n21349 ;
  assign n21352 = ~n16231 & n21350 ;
  assign n21351 = n16231 & ~n21350 ;
  assign n21353 = ~\P3_DataWidth_reg[1]/NET0131  & ~n21351 ;
  assign n21354 = ~n21352 & n21353 ;
  assign n21348 = \P3_DataWidth_reg[1]/NET0131  & ~\P3_rEIP_reg[6]/NET0131  ;
  assign n21355 = n2959 & ~n21348 ;
  assign n21356 = ~n21354 & n21355 ;
  assign n21359 = ~\P3_rEIP_reg[6]/NET0131  & ~n20417 ;
  assign n21360 = ~n20418 & ~n21359 ;
  assign n21369 = n20412 & ~n21360 ;
  assign n21370 = ~\P3_EBX_reg[6]/NET0131  & ~n20412 ;
  assign n21371 = ~n21369 & ~n21370 ;
  assign n21372 = n16094 & n21371 ;
  assign n21358 = \P3_rEIP_reg[6]/NET0131  & n2910 ;
  assign n21361 = n2946 & ~n21360 ;
  assign n21362 = \P3_EBX_reg[31]/NET0131  & ~n20433 ;
  assign n21364 = ~\P3_EBX_reg[6]/NET0131  & n21362 ;
  assign n21363 = \P3_EBX_reg[6]/NET0131  & ~n21362 ;
  assign n21365 = ~n2946 & ~n21363 ;
  assign n21366 = ~n21364 & n21365 ;
  assign n21367 = ~n21361 & ~n21366 ;
  assign n21368 = n20473 & n21367 ;
  assign n21373 = ~n21358 & ~n21368 ;
  assign n21374 = ~n21372 & n21373 ;
  assign n21375 = n2453 & ~n21374 ;
  assign n21357 = \P3_rEIP_reg[6]/NET0131  & ~n20409 ;
  assign n21376 = \P3_PhyAddrPointer_reg[6]/NET0131  & n3004 ;
  assign n21377 = ~n4412 & ~n21376 ;
  assign n21378 = ~n21357 & n21377 ;
  assign n21379 = ~n21375 & n21378 ;
  assign n21380 = ~n21356 & n21379 ;
  assign n21382 = ~n9054 & ~n20400 ;
  assign n21384 = ~n14501 & n21382 ;
  assign n21383 = n14501 & ~n21382 ;
  assign n21385 = ~\P3_DataWidth_reg[1]/NET0131  & ~n21383 ;
  assign n21386 = ~n21384 & n21385 ;
  assign n21381 = \P3_DataWidth_reg[1]/NET0131  & ~\P3_rEIP_reg[7]/NET0131  ;
  assign n21387 = n2959 & ~n21381 ;
  assign n21388 = ~n21386 & n21387 ;
  assign n21391 = ~\P3_rEIP_reg[7]/NET0131  & ~n20418 ;
  assign n21392 = ~n20419 & ~n21391 ;
  assign n21401 = n20412 & ~n21392 ;
  assign n21402 = ~\P3_EBX_reg[7]/NET0131  & ~n20412 ;
  assign n21403 = ~n21401 & ~n21402 ;
  assign n21404 = n16094 & n21403 ;
  assign n21390 = \P3_rEIP_reg[7]/NET0131  & n2910 ;
  assign n21393 = n2946 & ~n21392 ;
  assign n21394 = \P3_EBX_reg[31]/NET0131  & ~n20434 ;
  assign n21396 = ~\P3_EBX_reg[7]/NET0131  & n21394 ;
  assign n21395 = \P3_EBX_reg[7]/NET0131  & ~n21394 ;
  assign n21397 = ~n2946 & ~n21395 ;
  assign n21398 = ~n21396 & n21397 ;
  assign n21399 = ~n21393 & ~n21398 ;
  assign n21400 = n20473 & n21399 ;
  assign n21405 = ~n21390 & ~n21400 ;
  assign n21406 = ~n21404 & n21405 ;
  assign n21407 = n2453 & ~n21406 ;
  assign n21389 = \P3_rEIP_reg[7]/NET0131  & ~n20409 ;
  assign n21408 = \P3_PhyAddrPointer_reg[7]/NET0131  & n3004 ;
  assign n21409 = ~n4412 & ~n21408 ;
  assign n21410 = ~n21389 & n21409 ;
  assign n21411 = ~n21407 & n21410 ;
  assign n21412 = ~n21388 & n21411 ;
  assign n21414 = n9024 & n21207 ;
  assign n21415 = ~n9054 & ~n21414 ;
  assign n21417 = ~n13253 & n21415 ;
  assign n21416 = n13253 & ~n21415 ;
  assign n21418 = ~\P3_DataWidth_reg[1]/NET0131  & ~n21416 ;
  assign n21419 = ~n21417 & n21418 ;
  assign n21413 = \P3_DataWidth_reg[1]/NET0131  & ~\P3_rEIP_reg[8]/NET0131  ;
  assign n21420 = n2959 & ~n21413 ;
  assign n21421 = ~n21419 & n21420 ;
  assign n21423 = \P3_rEIP_reg[8]/NET0131  & n2910 ;
  assign n21424 = ~\P3_rEIP_reg[8]/NET0131  & ~n20419 ;
  assign n21425 = ~n20420 & ~n21424 ;
  assign n21426 = n2946 & ~n21425 ;
  assign n21427 = ~\P3_EBX_reg[8]/NET0131  & ~n20412 ;
  assign n21428 = n2818 & ~n21427 ;
  assign n21429 = \P3_EBX_reg[31]/NET0131  & ~n20435 ;
  assign n21431 = \P3_EBX_reg[8]/NET0131  & ~n21429 ;
  assign n21430 = ~\P3_EBX_reg[8]/NET0131  & n21429 ;
  assign n21432 = ~n2946 & ~n21430 ;
  assign n21433 = ~n21431 & n21432 ;
  assign n21434 = n2821 & ~n21433 ;
  assign n21435 = ~n21428 & ~n21434 ;
  assign n21436 = ~n21426 & ~n21435 ;
  assign n21437 = n2786 & n21428 ;
  assign n21438 = ~n21436 & ~n21437 ;
  assign n21439 = ~n2815 & ~n21438 ;
  assign n21440 = ~n21423 & ~n21439 ;
  assign n21441 = n2453 & ~n21440 ;
  assign n21422 = \P3_rEIP_reg[8]/NET0131  & ~n20409 ;
  assign n21442 = \P3_PhyAddrPointer_reg[8]/NET0131  & n3004 ;
  assign n21443 = ~n4412 & ~n21442 ;
  assign n21444 = ~n21422 & n21443 ;
  assign n21445 = ~n21441 & n21444 ;
  assign n21446 = ~n21421 & n21445 ;
  assign n21448 = ~\P3_PhyAddrPointer_reg[0]/NET0131  & n13252 ;
  assign n21449 = ~n9054 & ~n21448 ;
  assign n21451 = ~n14522 & n21449 ;
  assign n21450 = n14522 & ~n21449 ;
  assign n21452 = ~\P3_DataWidth_reg[1]/NET0131  & ~n21450 ;
  assign n21453 = ~n21451 & n21452 ;
  assign n21447 = \P3_DataWidth_reg[1]/NET0131  & ~\P3_rEIP_reg[9]/NET0131  ;
  assign n21454 = n2959 & ~n21447 ;
  assign n21455 = ~n21453 & n21454 ;
  assign n21457 = \P3_rEIP_reg[9]/NET0131  & n2910 ;
  assign n21458 = ~\P3_rEIP_reg[9]/NET0131  & ~n20420 ;
  assign n21459 = ~n20421 & ~n21458 ;
  assign n21460 = n2946 & ~n21459 ;
  assign n21461 = ~n2786 & n21460 ;
  assign n21462 = ~\P3_EBX_reg[9]/NET0131  & ~n20412 ;
  assign n21463 = n2818 & ~n21462 ;
  assign n21464 = ~n21461 & n21463 ;
  assign n21465 = \P3_EBX_reg[31]/NET0131  & ~n20436 ;
  assign n21467 = ~\P3_EBX_reg[9]/NET0131  & n21465 ;
  assign n21466 = \P3_EBX_reg[9]/NET0131  & ~n21465 ;
  assign n21468 = ~n2946 & ~n21466 ;
  assign n21469 = ~n21467 & n21468 ;
  assign n21470 = n2821 & ~n21460 ;
  assign n21471 = ~n21469 & n21470 ;
  assign n21472 = ~n21464 & ~n21471 ;
  assign n21473 = ~n2815 & ~n21472 ;
  assign n21474 = ~n21457 & ~n21473 ;
  assign n21475 = n2453 & ~n21474 ;
  assign n21456 = \P3_rEIP_reg[9]/NET0131  & ~n20409 ;
  assign n21476 = \P3_PhyAddrPointer_reg[9]/NET0131  & n3004 ;
  assign n21477 = ~n4412 & ~n21476 ;
  assign n21478 = ~n21456 & n21477 ;
  assign n21479 = ~n21475 & n21478 ;
  assign n21480 = ~n21455 & n21479 ;
  assign n21482 = \P1_PhyAddrPointer_reg[9]/NET0131  & n18542 ;
  assign n21483 = n18540 & ~n21482 ;
  assign n21485 = ~n14543 & n21483 ;
  assign n21484 = n14543 & ~n21483 ;
  assign n21486 = ~\P1_DataWidth_reg[1]/NET0131  & ~n21484 ;
  assign n21487 = ~n21485 & n21486 ;
  assign n21481 = \P1_DataWidth_reg[1]/NET0131  & ~\P1_rEIP_reg[10]/NET0131  ;
  assign n21488 = n2436 & ~n21481 ;
  assign n21489 = ~n21487 & n21488 ;
  assign n21491 = \P1_rEIP_reg[10]/NET0131  & ~n18554 ;
  assign n21493 = ~\P1_rEIP_reg[10]/NET0131  & ~n18565 ;
  assign n21494 = ~n18566 & ~n21493 ;
  assign n21495 = n18556 & ~n21494 ;
  assign n21492 = ~\P1_EBX_reg[10]/NET0131  & ~n18556 ;
  assign n21496 = n2225 & ~n21492 ;
  assign n21497 = ~n21495 & n21496 ;
  assign n21499 = \P1_EBX_reg[31]/NET0131  & ~n18585 ;
  assign n21501 = ~\P1_EBX_reg[10]/NET0131  & n21499 ;
  assign n21500 = \P1_EBX_reg[10]/NET0131  & ~n21499 ;
  assign n21502 = ~n2425 & ~n21500 ;
  assign n21503 = ~n21501 & n21502 ;
  assign n21498 = n2425 & ~n21494 ;
  assign n21504 = n2222 & ~n21498 ;
  assign n21505 = ~n21503 & n21504 ;
  assign n21506 = ~n21497 & ~n21505 ;
  assign n21507 = ~n2301 & ~n21506 ;
  assign n21508 = ~n21491 & ~n21507 ;
  assign n21509 = n2432 & ~n21508 ;
  assign n21490 = \P1_rEIP_reg[10]/NET0131  & ~n18552 ;
  assign n21510 = \P1_PhyAddrPointer_reg[10]/NET0131  & n3028 ;
  assign n21511 = ~n5092 & ~n21510 ;
  assign n21512 = ~n21490 & n21511 ;
  assign n21513 = ~n21509 & n21512 ;
  assign n21514 = ~n21489 & n21513 ;
  assign n21516 = \P1_PhyAddrPointer_reg[10]/NET0131  & n21482 ;
  assign n21517 = n18540 & ~n21516 ;
  assign n21519 = n12156 & ~n21517 ;
  assign n21518 = ~n12156 & n21517 ;
  assign n21520 = ~\P1_DataWidth_reg[1]/NET0131  & ~n21518 ;
  assign n21521 = ~n21519 & n21520 ;
  assign n21515 = \P1_DataWidth_reg[1]/NET0131  & ~\P1_rEIP_reg[11]/NET0131  ;
  assign n21522 = n2436 & ~n21515 ;
  assign n21523 = ~n21521 & n21522 ;
  assign n21525 = \P1_rEIP_reg[11]/NET0131  & ~n18554 ;
  assign n21527 = ~\P1_rEIP_reg[11]/NET0131  & ~n18566 ;
  assign n21528 = ~n18567 & ~n21527 ;
  assign n21529 = n18556 & ~n21528 ;
  assign n21526 = ~\P1_EBX_reg[11]/NET0131  & ~n18556 ;
  assign n21530 = n2225 & ~n21526 ;
  assign n21531 = ~n21529 & n21530 ;
  assign n21533 = \P1_EBX_reg[31]/NET0131  & ~n18586 ;
  assign n21535 = \P1_EBX_reg[11]/NET0131  & ~n21533 ;
  assign n21534 = ~\P1_EBX_reg[11]/NET0131  & n21533 ;
  assign n21536 = ~n2425 & ~n21534 ;
  assign n21537 = ~n21535 & n21536 ;
  assign n21532 = n2425 & ~n21528 ;
  assign n21538 = n2222 & ~n21532 ;
  assign n21539 = ~n21537 & n21538 ;
  assign n21540 = ~n21531 & ~n21539 ;
  assign n21541 = ~n2301 & ~n21540 ;
  assign n21542 = ~n21525 & ~n21541 ;
  assign n21543 = n2432 & ~n21542 ;
  assign n21524 = \P1_rEIP_reg[11]/NET0131  & ~n18552 ;
  assign n21544 = \P1_PhyAddrPointer_reg[11]/NET0131  & n3028 ;
  assign n21545 = ~n5092 & ~n21544 ;
  assign n21546 = ~n21524 & n21545 ;
  assign n21547 = ~n21543 & n21546 ;
  assign n21548 = ~n21523 & n21547 ;
  assign n21550 = ~\P1_PhyAddrPointer_reg[0]/NET0131  & n12155 ;
  assign n21551 = n18540 & ~n21550 ;
  assign n21553 = n13284 & ~n21551 ;
  assign n21552 = ~n13284 & n21551 ;
  assign n21554 = ~\P1_DataWidth_reg[1]/NET0131  & ~n21552 ;
  assign n21555 = ~n21553 & n21554 ;
  assign n21549 = \P1_DataWidth_reg[1]/NET0131  & ~\P1_rEIP_reg[12]/NET0131  ;
  assign n21556 = n2436 & ~n21549 ;
  assign n21557 = ~n21555 & n21556 ;
  assign n21559 = \P1_rEIP_reg[12]/NET0131  & ~n18554 ;
  assign n21561 = ~\P1_rEIP_reg[12]/NET0131  & ~n18567 ;
  assign n21562 = ~n18568 & ~n21561 ;
  assign n21563 = n2425 & ~n21562 ;
  assign n21564 = ~n2311 & n21563 ;
  assign n21560 = ~\P1_EBX_reg[12]/NET0131  & ~n18556 ;
  assign n21565 = n2225 & ~n21560 ;
  assign n21566 = ~n21564 & n21565 ;
  assign n21567 = \P1_EBX_reg[31]/NET0131  & ~n18587 ;
  assign n21569 = \P1_EBX_reg[12]/NET0131  & ~n21567 ;
  assign n21568 = ~\P1_EBX_reg[12]/NET0131  & n21567 ;
  assign n21570 = ~n2425 & ~n21568 ;
  assign n21571 = ~n21569 & n21570 ;
  assign n21572 = n2222 & ~n21563 ;
  assign n21573 = ~n21571 & n21572 ;
  assign n21574 = ~n21566 & ~n21573 ;
  assign n21575 = ~n2301 & ~n21574 ;
  assign n21576 = ~n21559 & ~n21575 ;
  assign n21577 = n2432 & ~n21576 ;
  assign n21558 = \P1_rEIP_reg[12]/NET0131  & ~n18552 ;
  assign n21578 = \P1_PhyAddrPointer_reg[12]/NET0131  & n3028 ;
  assign n21579 = ~n5092 & ~n21578 ;
  assign n21580 = ~n21558 & n21579 ;
  assign n21581 = ~n21577 & n21580 ;
  assign n21582 = ~n21557 & n21581 ;
  assign n21584 = n10101 & n18542 ;
  assign n21585 = n18540 & ~n21584 ;
  assign n21587 = n13317 & ~n21585 ;
  assign n21586 = ~n13317 & n21585 ;
  assign n21588 = ~\P1_DataWidth_reg[1]/NET0131  & ~n21586 ;
  assign n21589 = ~n21587 & n21588 ;
  assign n21583 = \P1_DataWidth_reg[1]/NET0131  & ~\P1_rEIP_reg[13]/NET0131  ;
  assign n21590 = n2436 & ~n21583 ;
  assign n21591 = ~n21589 & n21590 ;
  assign n21593 = \P1_rEIP_reg[13]/NET0131  & ~n18554 ;
  assign n21595 = ~\P1_rEIP_reg[13]/NET0131  & ~n18568 ;
  assign n21596 = ~n18569 & ~n21595 ;
  assign n21597 = n2425 & ~n21596 ;
  assign n21598 = ~n2311 & n21597 ;
  assign n21594 = ~\P1_EBX_reg[13]/NET0131  & ~n18556 ;
  assign n21599 = n2225 & ~n21594 ;
  assign n21600 = ~n21598 & n21599 ;
  assign n21601 = \P1_EBX_reg[31]/NET0131  & ~n18588 ;
  assign n21603 = ~\P1_EBX_reg[13]/NET0131  & n21601 ;
  assign n21602 = \P1_EBX_reg[13]/NET0131  & ~n21601 ;
  assign n21604 = ~n2425 & ~n21602 ;
  assign n21605 = ~n21603 & n21604 ;
  assign n21606 = n2222 & ~n21597 ;
  assign n21607 = ~n21605 & n21606 ;
  assign n21608 = ~n21600 & ~n21607 ;
  assign n21609 = ~n2301 & ~n21608 ;
  assign n21610 = ~n21593 & ~n21609 ;
  assign n21611 = n2432 & ~n21610 ;
  assign n21592 = \P1_rEIP_reg[13]/NET0131  & ~n18552 ;
  assign n21612 = \P1_PhyAddrPointer_reg[13]/NET0131  & n3028 ;
  assign n21613 = ~n5092 & ~n21612 ;
  assign n21614 = ~n21592 & n21613 ;
  assign n21615 = ~n21611 & n21614 ;
  assign n21616 = ~n21591 & n21615 ;
  assign n21619 = n1734 & n13778 ;
  assign n21618 = n1890 & n13795 ;
  assign n21620 = \P2_PhyAddrPointer_reg[2]/NET0131  & ~n12395 ;
  assign n21621 = ~n21618 & ~n21620 ;
  assign n21622 = ~n21619 & n21621 ;
  assign n21623 = n1927 & ~n21622 ;
  assign n21624 = n9005 & n20034 ;
  assign n21625 = \P2_PhyAddrPointer_reg[2]/NET0131  & ~n8958 ;
  assign n21617 = ~\P2_PhyAddrPointer_reg[2]/NET0131  & n3034 ;
  assign n21626 = ~n13763 & ~n21617 ;
  assign n21627 = ~n21625 & n21626 ;
  assign n21628 = ~n21624 & n21627 ;
  assign n21629 = ~n21623 & n21628 ;
  assign n21632 = ~\P2_RequestPending_reg/NET0131  & n1810 ;
  assign n21633 = ~n1824 & ~n21632 ;
  assign n21630 = \P2_RequestPending_reg/NET0131  & n1747 ;
  assign n21631 = ~\P2_DataWidth_reg[1]/NET0131  & n15980 ;
  assign n21634 = ~n21630 & ~n21631 ;
  assign n21635 = ~n21633 & n21634 ;
  assign n21636 = n1927 & ~n21635 ;
  assign n21639 = \P2_RequestPending_reg/NET0131  & ~n12630 ;
  assign n21637 = \P2_RequestPending_reg/NET0131  & n1935 ;
  assign n21638 = n2977 & n21637 ;
  assign n21640 = ~n1933 & ~n3113 ;
  assign n21641 = ~n21638 & n21640 ;
  assign n21642 = ~n21639 & n21641 ;
  assign n21643 = ~n21636 & n21642 ;
  assign n21645 = \P3_PhyAddrPointer_reg[2]/NET0131  & ~n11965 ;
  assign n21646 = n2905 & n13739 ;
  assign n21647 = ~n13755 & ~n21646 ;
  assign n21648 = ~n21645 & n21647 ;
  assign n21649 = n2453 & ~n21648 ;
  assign n21651 = ~n2997 & ~n4414 ;
  assign n21652 = ~n2955 & n21651 ;
  assign n21653 = \P3_PhyAddrPointer_reg[2]/NET0131  & ~n21652 ;
  assign n21644 = n10076 & n21210 ;
  assign n21650 = ~\P3_PhyAddrPointer_reg[2]/NET0131  & n2970 ;
  assign n21654 = ~n13732 & ~n21650 ;
  assign n21655 = ~n21644 & n21654 ;
  assign n21656 = ~n21653 & n21655 ;
  assign n21657 = ~n21649 & n21656 ;
  assign n21661 = ~\P3_DataWidth_reg[1]/NET0131  & n2818 ;
  assign n21662 = n2891 & ~n21661 ;
  assign n21663 = ~n2766 & n21662 ;
  assign n21664 = \P3_RequestPending_reg/NET0131  & ~n21663 ;
  assign n21665 = ~n2815 & ~n21662 ;
  assign n21666 = ~n21664 & ~n21665 ;
  assign n21667 = n2453 & ~n21666 ;
  assign n21658 = n2835 & n16888 ;
  assign n21659 = n13808 & ~n21658 ;
  assign n21660 = \P3_RequestPending_reg/NET0131  & ~n21659 ;
  assign n21668 = ~n2953 & ~n4412 ;
  assign n21669 = ~n21660 & n21668 ;
  assign n21670 = ~n21667 & n21669 ;
  assign n21672 = n2384 & n13710 ;
  assign n21673 = \P1_PhyAddrPointer_reg[2]/NET0131  & ~n12209 ;
  assign n21674 = ~n13723 & ~n21673 ;
  assign n21675 = ~n21672 & n21674 ;
  assign n21676 = n2432 & ~n21675 ;
  assign n21677 = n10133 & n19667 ;
  assign n21678 = \P1_PhyAddrPointer_reg[2]/NET0131  & ~n10136 ;
  assign n21671 = ~\P1_PhyAddrPointer_reg[2]/NET0131  & n3148 ;
  assign n21679 = ~n13694 & ~n21671 ;
  assign n21680 = ~n21678 & n21679 ;
  assign n21681 = ~n21677 & n21680 ;
  assign n21682 = ~n21676 & n21681 ;
  assign n21688 = ~\P1_RequestPending_reg/NET0131  & n2301 ;
  assign n21689 = n2379 & ~n21688 ;
  assign n21686 = \P1_RequestPending_reg/NET0131  & n2233 ;
  assign n21687 = ~\P1_DataWidth_reg[1]/NET0131  & n15990 ;
  assign n21690 = ~n21686 & ~n21687 ;
  assign n21691 = ~n21689 & n21690 ;
  assign n21692 = n2432 & ~n21691 ;
  assign n21683 = n2317 & n2440 ;
  assign n21684 = n15401 & ~n21683 ;
  assign n21685 = \P1_RequestPending_reg/NET0131  & ~n21684 ;
  assign n21693 = n5288 & ~n21685 ;
  assign n21694 = ~n21692 & n21693 ;
  assign n21696 = \P1_Datao_reg[20]/NET0131  & n2306 ;
  assign n21697 = ~n2225 & n2312 ;
  assign n21698 = ~n2306 & ~n21697 ;
  assign n21699 = ~\P1_Datao_reg[20]/NET0131  & ~n2312 ;
  assign n21700 = ~\P1_EAX_reg[20]/NET0131  & ~n16019 ;
  assign n21701 = \P1_EAX_reg[20]/NET0131  & n16019 ;
  assign n21702 = ~n21700 & ~n21701 ;
  assign n21703 = n2312 & ~n21702 ;
  assign n21704 = ~n21699 & ~n21703 ;
  assign n21705 = n21698 & n21704 ;
  assign n21706 = ~n21696 & ~n21705 ;
  assign n21707 = n2432 & ~n21706 ;
  assign n21695 = \P1_uWord_reg[4]/NET0131  & n2440 ;
  assign n21708 = \P1_Datao_reg[20]/NET0131  & ~n16884 ;
  assign n21709 = ~n21695 & ~n21708 ;
  assign n21710 = ~n21707 & n21709 ;
  assign n21712 = \datao[20]_pad  & ~n2833 ;
  assign n21713 = ~\P3_EAX_reg[20]/NET0131  & ~n16113 ;
  assign n21714 = ~n16114 & ~n21713 ;
  assign n21715 = n16094 & n21714 ;
  assign n21716 = ~n2786 & n21715 ;
  assign n21717 = ~n21712 & ~n21716 ;
  assign n21718 = n2453 & ~n21717 ;
  assign n21711 = \P3_uWord_reg[4]/NET0131  & n16888 ;
  assign n21719 = \datao[20]_pad  & ~n16899 ;
  assign n21720 = ~n21711 & ~n21719 ;
  assign n21721 = ~n21718 & n21720 ;
  assign n21723 = ~\P2_EAX_reg[20]/NET0131  & ~n15968 ;
  assign n21724 = ~n15969 & ~n21723 ;
  assign n21725 = ~n1819 & ~n21724 ;
  assign n21726 = n15980 & ~n21725 ;
  assign n21727 = n16922 & ~n21726 ;
  assign n21728 = \P2_Datao_reg[20]/NET0131  & ~n21727 ;
  assign n21729 = n1922 & n21724 ;
  assign n21730 = ~n21728 & ~n21729 ;
  assign n21731 = n1927 & ~n21730 ;
  assign n21722 = \P2_uWord_reg[4]/NET0131  & n16919 ;
  assign n21732 = \P2_Datao_reg[20]/NET0131  & ~n16936 ;
  assign n21733 = ~n21722 & ~n21732 ;
  assign n21734 = ~n21731 & n21733 ;
  assign n21735 = \P1_EAX_reg[25]/NET0131  & ~n15402 ;
  assign n21737 = ~\P1_EAX_reg[25]/NET0131  & ~n15918 ;
  assign n21738 = n15920 & ~n21737 ;
  assign n21736 = \P1_EAX_reg[25]/NET0131  & ~n15925 ;
  assign n21739 = n2302 & ~n5255 ;
  assign n21740 = n2222 & ~n5158 ;
  assign n21741 = ~n21739 & ~n21740 ;
  assign n21742 = n2377 & ~n21741 ;
  assign n21743 = ~n15200 & n15231 ;
  assign n21744 = n2337 & ~n15232 ;
  assign n21745 = ~n21743 & n21744 ;
  assign n21746 = n2331 & n21745 ;
  assign n21747 = ~n21742 & ~n21746 ;
  assign n21748 = ~n21736 & n21747 ;
  assign n21749 = ~n21738 & n21748 ;
  assign n21750 = n2432 & ~n21749 ;
  assign n21751 = ~n21735 & ~n21750 ;
  assign n21752 = \P2_uWord_reg[4]/NET0131  & ~n15942 ;
  assign n21755 = n1811 & ~n3082 ;
  assign n21756 = \P2_uWord_reg[4]/NET0131  & n1805 ;
  assign n21757 = ~n21755 & ~n21756 ;
  assign n21758 = n1742 & ~n21757 ;
  assign n21753 = \P2_uWord_reg[4]/NET0131  & n15981 ;
  assign n21754 = n15980 & n21724 ;
  assign n21759 = ~n21753 & ~n21754 ;
  assign n21760 = ~n21758 & n21759 ;
  assign n21761 = n1927 & ~n21760 ;
  assign n21762 = ~n21752 & ~n21761 ;
  assign n21763 = \P1_uWord_reg[4]/NET0131  & ~n15994 ;
  assign n21764 = n15990 & n21702 ;
  assign n21765 = ~n5140 & n15932 ;
  assign n21766 = ~n21764 & ~n21765 ;
  assign n21767 = n2432 & ~n21766 ;
  assign n21768 = ~n21763 & ~n21767 ;
  assign n21769 = \P3_EAX_reg[25]/NET0131  & ~n13810 ;
  assign n21773 = n14037 & n14039 ;
  assign n21774 = ~\P3_EAX_reg[25]/NET0131  & ~n21773 ;
  assign n21775 = n13813 & ~n14041 ;
  assign n21776 = ~n21774 & n21775 ;
  assign n21777 = \P3_EAX_reg[25]/NET0131  & ~n14922 ;
  assign n21770 = ~n13913 & n13944 ;
  assign n21771 = ~n13945 & ~n21770 ;
  assign n21772 = n13812 & n21771 ;
  assign n21778 = \buf2_reg[25]/NET0131  & n2820 ;
  assign n21779 = \buf2_reg[9]/NET0131  & n2821 ;
  assign n21780 = ~n21778 & ~n21779 ;
  assign n21781 = n2862 & ~n21780 ;
  assign n21782 = ~n21772 & ~n21781 ;
  assign n21783 = ~n21777 & n21782 ;
  assign n21784 = ~n21776 & n21783 ;
  assign n21785 = n2453 & ~n21784 ;
  assign n21786 = ~n21769 & ~n21785 ;
  assign n21787 = \P2_EAX_reg[25]/NET0131  & ~n12632 ;
  assign n21792 = \P2_EAX_reg[23]/NET0131  & n12655 ;
  assign n21793 = \P2_EAX_reg[24]/NET0131  & n21792 ;
  assign n21794 = n12664 & ~n21793 ;
  assign n21795 = n12668 & ~n21794 ;
  assign n21796 = \P2_EAX_reg[25]/NET0131  & ~n21795 ;
  assign n21803 = ~\P2_EAX_reg[25]/NET0131  & n12664 ;
  assign n21804 = n21793 & n21803 ;
  assign n21797 = \P2_EAX_reg[25]/NET0131  & ~n1811 ;
  assign n21800 = n1811 & ~n11549 ;
  assign n21801 = ~n21797 & ~n21800 ;
  assign n21802 = n1803 & ~n21801 ;
  assign n21788 = ~n12768 & n12799 ;
  assign n21789 = n1798 & ~n12800 ;
  assign n21790 = ~n21788 & n21789 ;
  assign n21791 = n1726 & n21790 ;
  assign n21798 = ~n17935 & ~n21797 ;
  assign n21799 = n1742 & ~n21798 ;
  assign n21805 = ~n21791 & ~n21799 ;
  assign n21806 = ~n21802 & n21805 ;
  assign n21807 = ~n21804 & n21806 ;
  assign n21808 = ~n21796 & n21807 ;
  assign n21809 = n1927 & ~n21808 ;
  assign n21810 = ~n21787 & ~n21809 ;
  assign n21811 = \P3_uWord_reg[4]/NET0131  & ~n16086 ;
  assign n21812 = \buf2_reg[4]/NET0131  & n2862 ;
  assign n21813 = \P3_uWord_reg[4]/NET0131  & n2835 ;
  assign n21814 = ~n21812 & ~n21813 ;
  assign n21815 = n2821 & ~n21814 ;
  assign n21816 = \P3_uWord_reg[4]/NET0131  & ~n2908 ;
  assign n21817 = ~n21715 & ~n21816 ;
  assign n21818 = ~n21815 & n21817 ;
  assign n21819 = n2453 & ~n21818 ;
  assign n21820 = ~n21811 & ~n21819 ;
  assign n21828 = \P3_InstQueue_reg[0][7]/NET0131  & ~n18218 ;
  assign n21823 = n2539 & n18209 ;
  assign n21822 = ~\P3_InstQueue_reg[0][7]/NET0131  & ~n18209 ;
  assign n21824 = n2994 & ~n21822 ;
  assign n21825 = ~n21823 & n21824 ;
  assign n21821 = \buf2_reg[7]/NET0131  & n18228 ;
  assign n21826 = \buf2_reg[23]/NET0131  & n2970 ;
  assign n21827 = n18203 & n21826 ;
  assign n21829 = ~n21821 & ~n21827 ;
  assign n21830 = ~n21825 & n21829 ;
  assign n21831 = ~n21828 & n21830 ;
  assign n21838 = \P3_InstQueue_reg[10][7]/NET0131  & ~n18243 ;
  assign n21834 = n2539 & n18246 ;
  assign n21833 = ~\P3_InstQueue_reg[10][7]/NET0131  & ~n18246 ;
  assign n21835 = n2994 & ~n21833 ;
  assign n21836 = ~n21834 & n21835 ;
  assign n21832 = \buf2_reg[7]/NET0131  & n18255 ;
  assign n21837 = n18236 & n21826 ;
  assign n21839 = ~n21832 & ~n21837 ;
  assign n21840 = ~n21836 & n21839 ;
  assign n21841 = ~n21838 & n21840 ;
  assign n21843 = n2539 & n18266 ;
  assign n21842 = ~\P3_InstQueue_reg[11][7]/NET0131  & ~n18266 ;
  assign n21844 = n2994 & ~n21842 ;
  assign n21845 = ~n21843 & n21844 ;
  assign n21847 = \P3_InstQueue_reg[11][7]/NET0131  & ~n18264 ;
  assign n21846 = n18271 & n21826 ;
  assign n21848 = \buf2_reg[7]/NET0131  & n18245 ;
  assign n21849 = n18262 & n21848 ;
  assign n21850 = ~n21846 & ~n21849 ;
  assign n21851 = ~n21847 & n21850 ;
  assign n21852 = ~n21845 & n21851 ;
  assign n21859 = \P3_InstQueue_reg[12][7]/NET0131  & ~n18287 ;
  assign n21855 = n2539 & n18284 ;
  assign n21854 = ~\P3_InstQueue_reg[12][7]/NET0131  & ~n18284 ;
  assign n21856 = n2994 & ~n21854 ;
  assign n21857 = ~n21855 & n21856 ;
  assign n21853 = \buf2_reg[7]/NET0131  & n18297 ;
  assign n21858 = n18246 & n21826 ;
  assign n21860 = ~n21853 & ~n21858 ;
  assign n21861 = ~n21857 & n21860 ;
  assign n21862 = ~n21859 & n21861 ;
  assign n21870 = n2539 & n18200 ;
  assign n21869 = ~\P3_InstQueue_reg[13][7]/NET0131  & ~n18200 ;
  assign n21871 = n2994 & ~n21869 ;
  assign n21872 = ~n21870 & n21871 ;
  assign n21866 = ~\P3_InstQueue_reg[13][7]/NET0131  & n18302 ;
  assign n21865 = ~\buf2_reg[7]/NET0131  & ~n18302 ;
  assign n21867 = n18305 & ~n21865 ;
  assign n21868 = ~n21866 & n21867 ;
  assign n21863 = n18266 & n21826 ;
  assign n21864 = \P3_InstQueue_reg[13][7]/NET0131  & ~n18217 ;
  assign n21873 = ~n21863 & ~n21864 ;
  assign n21874 = ~n21868 & n21873 ;
  assign n21875 = ~n21872 & n21874 ;
  assign n21882 = \P3_InstQueue_reg[14][7]/NET0131  & ~n18325 ;
  assign n21878 = n2539 & n18203 ;
  assign n21877 = ~\P3_InstQueue_reg[14][7]/NET0131  & ~n18203 ;
  assign n21879 = n2994 & ~n21877 ;
  assign n21880 = ~n21878 & n21879 ;
  assign n21876 = \buf2_reg[7]/NET0131  & n18335 ;
  assign n21881 = n18284 & n21826 ;
  assign n21883 = ~n21876 & ~n21881 ;
  assign n21884 = ~n21880 & n21883 ;
  assign n21885 = ~n21882 & n21884 ;
  assign n21893 = n2539 & n18212 ;
  assign n21892 = ~\P3_InstQueue_reg[15][7]/NET0131  & ~n18212 ;
  assign n21894 = n2994 & ~n21892 ;
  assign n21895 = ~n21893 & n21894 ;
  assign n21888 = ~\buf2_reg[7]/NET0131  & ~n18342 ;
  assign n21889 = ~\P3_InstQueue_reg[15][7]/NET0131  & n18342 ;
  assign n21890 = ~n21888 & ~n21889 ;
  assign n21891 = ~n18341 & n21890 ;
  assign n21886 = n18200 & n21826 ;
  assign n21887 = \P3_InstQueue_reg[15][7]/NET0131  & ~n18217 ;
  assign n21896 = ~n21886 & ~n21887 ;
  assign n21897 = ~n21891 & n21896 ;
  assign n21898 = ~n21895 & n21897 ;
  assign n21905 = \P3_InstQueue_reg[1][7]/NET0131  & ~n18364 ;
  assign n21901 = n2539 & n18361 ;
  assign n21900 = ~\P3_InstQueue_reg[1][7]/NET0131  & ~n18361 ;
  assign n21902 = n2994 & ~n21900 ;
  assign n21903 = ~n21901 & n21902 ;
  assign n21899 = \buf2_reg[7]/NET0131  & n18374 ;
  assign n21904 = n18212 & n21826 ;
  assign n21906 = ~n21899 & ~n21904 ;
  assign n21907 = ~n21903 & n21906 ;
  assign n21908 = ~n21905 & n21907 ;
  assign n21915 = \P3_InstQueue_reg[2][7]/NET0131  & ~n18383 ;
  assign n21911 = n2539 & n18386 ;
  assign n21910 = ~\P3_InstQueue_reg[2][7]/NET0131  & ~n18386 ;
  assign n21912 = n2994 & ~n21910 ;
  assign n21913 = ~n21911 & n21912 ;
  assign n21909 = \buf2_reg[7]/NET0131  & n18395 ;
  assign n21914 = n18209 & n21826 ;
  assign n21916 = ~n21909 & ~n21914 ;
  assign n21917 = ~n21913 & n21916 ;
  assign n21918 = ~n21915 & n21917 ;
  assign n21925 = \P3_InstQueue_reg[3][7]/NET0131  & ~n18403 ;
  assign n21921 = n2539 & n18405 ;
  assign n21920 = ~\P3_InstQueue_reg[3][7]/NET0131  & ~n18405 ;
  assign n21922 = n2994 & ~n21920 ;
  assign n21923 = ~n21921 & n21922 ;
  assign n21919 = \buf2_reg[7]/NET0131  & n18414 ;
  assign n21924 = n18361 & n21826 ;
  assign n21926 = ~n21919 & ~n21924 ;
  assign n21927 = ~n21923 & n21926 ;
  assign n21928 = ~n21925 & n21927 ;
  assign n21935 = \P3_InstQueue_reg[4][7]/NET0131  & ~n18424 ;
  assign n21931 = n2539 & n18421 ;
  assign n21930 = ~\P3_InstQueue_reg[4][7]/NET0131  & ~n18421 ;
  assign n21932 = n2994 & ~n21930 ;
  assign n21933 = ~n21931 & n21932 ;
  assign n21929 = \buf2_reg[7]/NET0131  & n18434 ;
  assign n21934 = n18386 & n21826 ;
  assign n21936 = ~n21929 & ~n21934 ;
  assign n21937 = ~n21933 & n21936 ;
  assign n21938 = ~n21935 & n21937 ;
  assign n21946 = n2539 & n18439 ;
  assign n21945 = ~\P3_InstQueue_reg[5][7]/NET0131  & ~n18439 ;
  assign n21947 = n2994 & ~n21945 ;
  assign n21948 = ~n21946 & n21947 ;
  assign n21942 = ~\P3_InstQueue_reg[5][7]/NET0131  & n18440 ;
  assign n21941 = ~\buf2_reg[7]/NET0131  & ~n18440 ;
  assign n21943 = n18443 & ~n21941 ;
  assign n21944 = ~n21942 & n21943 ;
  assign n21939 = n18405 & n21826 ;
  assign n21940 = \P3_InstQueue_reg[5][7]/NET0131  & ~n18217 ;
  assign n21949 = ~n21939 & ~n21940 ;
  assign n21950 = ~n21944 & n21949 ;
  assign n21951 = ~n21948 & n21950 ;
  assign n21958 = \P3_InstQueue_reg[6][7]/NET0131  & ~n18465 ;
  assign n21954 = n2539 & n18462 ;
  assign n21953 = ~\P3_InstQueue_reg[6][7]/NET0131  & ~n18462 ;
  assign n21955 = n2994 & ~n21953 ;
  assign n21956 = ~n21954 & n21955 ;
  assign n21952 = \buf2_reg[7]/NET0131  & n18475 ;
  assign n21957 = n18421 & n21826 ;
  assign n21959 = ~n21952 & ~n21957 ;
  assign n21960 = ~n21956 & n21959 ;
  assign n21961 = ~n21958 & n21960 ;
  assign n21969 = n2539 & n18233 ;
  assign n21968 = ~\P3_InstQueue_reg[7][7]/NET0131  & ~n18233 ;
  assign n21970 = n2994 & ~n21968 ;
  assign n21971 = ~n21969 & n21970 ;
  assign n21964 = ~\buf2_reg[7]/NET0131  & ~n18482 ;
  assign n21965 = ~\P3_InstQueue_reg[7][7]/NET0131  & n18482 ;
  assign n21966 = ~n21964 & ~n21965 ;
  assign n21967 = ~n18481 & n21966 ;
  assign n21962 = n18439 & n21826 ;
  assign n21963 = \P3_InstQueue_reg[7][7]/NET0131  & ~n18217 ;
  assign n21972 = ~n21962 & ~n21963 ;
  assign n21973 = ~n21967 & n21972 ;
  assign n21974 = ~n21971 & n21973 ;
  assign n21981 = \P3_InstQueue_reg[8][7]/NET0131  & ~n18502 ;
  assign n21977 = n2539 & n18236 ;
  assign n21976 = ~\P3_InstQueue_reg[8][7]/NET0131  & ~n18236 ;
  assign n21978 = n2994 & ~n21976 ;
  assign n21979 = ~n21977 & n21978 ;
  assign n21975 = \buf2_reg[7]/NET0131  & n18512 ;
  assign n21980 = n18462 & n21826 ;
  assign n21982 = ~n21975 & ~n21980 ;
  assign n21983 = ~n21979 & n21982 ;
  assign n21984 = ~n21981 & n21983 ;
  assign n21987 = n2539 & n18271 ;
  assign n21986 = ~\P3_InstQueue_reg[9][7]/NET0131  & ~n18271 ;
  assign n21988 = n2994 & ~n21986 ;
  assign n21989 = ~n21987 & n21988 ;
  assign n21991 = ~n4415 & n18525 ;
  assign n21992 = \buf2_reg[7]/NET0131  & n18235 ;
  assign n21993 = \P3_InstQueue_reg[9][7]/NET0131  & ~n18235 ;
  assign n21994 = ~n21992 & ~n21993 ;
  assign n21995 = ~n10074 & ~n21994 ;
  assign n21996 = ~n21991 & n21995 ;
  assign n21985 = n18233 & n21826 ;
  assign n21990 = \P3_InstQueue_reg[9][7]/NET0131  & ~n18217 ;
  assign n21997 = ~n21985 & ~n21990 ;
  assign n21998 = ~n21996 & n21997 ;
  assign n21999 = ~n21989 & n21998 ;
  assign n22002 = \P3_MemoryFetch_reg/NET0131  & ~n2909 ;
  assign n22003 = ~n2908 & ~n22002 ;
  assign n22004 = n2453 & ~n22003 ;
  assign n22000 = ~n2993 & n4417 ;
  assign n22001 = \P3_MemoryFetch_reg/NET0131  & ~n22000 ;
  assign n22005 = n15433 & ~n22001 ;
  assign n22006 = ~n22004 & n22005 ;
  assign n22008 = \P1_MemoryFetch_reg/NET0131  & ~n18807 ;
  assign n22009 = n15991 & ~n22008 ;
  assign n22010 = n2432 & ~n22009 ;
  assign n22007 = \P1_MemoryFetch_reg/NET0131  & ~n15987 ;
  assign n22011 = n14083 & ~n22007 ;
  assign n22012 = ~n22010 & n22011 ;
  assign n22015 = n1745 & ~n1810 ;
  assign n22016 = \P2_MemoryFetch_reg/NET0131  & ~n22015 ;
  assign n22017 = n15981 & ~n22016 ;
  assign n22018 = n1927 & ~n22017 ;
  assign n22013 = ~n2986 & n6809 ;
  assign n22014 = \P2_MemoryFetch_reg/NET0131  & ~n22013 ;
  assign n22019 = n3114 & ~n22014 ;
  assign n22020 = ~n22018 & n22019 ;
  assign n22022 = ~n16553 & n16555 ;
  assign n22023 = \P2_rEIP_reg[0]/NET0131  & ~n22022 ;
  assign n22021 = \P2_EBX_reg[0]/NET0131  & ~n19071 ;
  assign n22024 = ~\P2_InstQueueRd_Addr_reg[0]/NET0131  & n22015 ;
  assign n22025 = ~n22021 & ~n22024 ;
  assign n22026 = ~n22023 & n22025 ;
  assign n22027 = n1927 & ~n22026 ;
  assign n22028 = ~n1932 & ~n2987 ;
  assign n22029 = \P2_PhyAddrPointer_reg[0]/NET0131  & ~n22028 ;
  assign n22030 = ~n3034 & n16511 ;
  assign n22031 = \P2_rEIP_reg[0]/NET0131  & ~n22030 ;
  assign n22032 = ~n22029 & ~n22031 ;
  assign n22033 = ~n22027 & n22032 ;
  assign n22038 = ~\P1_EBX_reg[29]/NET0131  & n19537 ;
  assign n22039 = \P1_EBX_reg[31]/NET0131  & ~n22038 ;
  assign n22041 = ~\P1_EBX_reg[30]/NET0131  & n22039 ;
  assign n22040 = \P1_EBX_reg[30]/NET0131  & ~n22039 ;
  assign n22042 = ~n2425 & ~n22040 ;
  assign n22043 = ~n22041 & n22042 ;
  assign n22034 = ~\P1_rEIP_reg[30]/NET0131  & ~n19524 ;
  assign n22035 = \P1_rEIP_reg[30]/NET0131  & n19524 ;
  assign n22036 = ~n22034 & ~n22035 ;
  assign n22037 = n2425 & ~n22036 ;
  assign n22044 = n7246 & ~n22037 ;
  assign n22045 = ~n22043 & n22044 ;
  assign n22046 = \P1_rEIP_reg[30]/NET0131  & ~n18554 ;
  assign n22048 = n18556 & ~n22036 ;
  assign n22047 = ~\P1_EBX_reg[30]/NET0131  & ~n18556 ;
  assign n22049 = n15990 & ~n22047 ;
  assign n22050 = ~n22048 & n22049 ;
  assign n22051 = ~n22046 & ~n22050 ;
  assign n22052 = ~n22045 & n22051 ;
  assign n22053 = n2432 & ~n22052 ;
  assign n22055 = \P1_PhyAddrPointer_reg[29]/NET0131  & n19549 ;
  assign n22056 = n18540 & ~n22055 ;
  assign n22058 = ~n10131 & n22056 ;
  assign n22057 = n10131 & ~n22056 ;
  assign n22059 = ~\P1_DataWidth_reg[1]/NET0131  & ~n22057 ;
  assign n22060 = ~n22058 & n22059 ;
  assign n22054 = \P1_DataWidth_reg[1]/NET0131  & ~\P1_rEIP_reg[30]/NET0131  ;
  assign n22061 = n2436 & ~n22054 ;
  assign n22062 = ~n22060 & n22061 ;
  assign n22063 = \P1_PhyAddrPointer_reg[30]/NET0131  & n3028 ;
  assign n22064 = \P1_rEIP_reg[30]/NET0131  & ~n18805 ;
  assign n22065 = ~n22063 & ~n22064 ;
  assign n22066 = ~n22062 & n22065 ;
  assign n22067 = ~n22053 & n22066 ;
  assign n22068 = ~\P1_rEIP_reg[31]/NET0131  & ~n22035 ;
  assign n22069 = \P1_rEIP_reg[31]/NET0131  & n22035 ;
  assign n22070 = ~n22068 & ~n22069 ;
  assign n22071 = n2425 & n22070 ;
  assign n22072 = ~\P1_EBX_reg[30]/NET0131  & \P1_EBX_reg[31]/NET0131  ;
  assign n22073 = n19527 & n22072 ;
  assign n22074 = n19537 & n22073 ;
  assign n22075 = ~n22071 & ~n22074 ;
  assign n22076 = n7246 & ~n22075 ;
  assign n22077 = \P1_rEIP_reg[31]/NET0131  & ~n18554 ;
  assign n22078 = n18556 & ~n22070 ;
  assign n22079 = ~\P1_EBX_reg[31]/NET0131  & ~n18556 ;
  assign n22080 = n15990 & ~n22079 ;
  assign n22081 = ~n22078 & n22080 ;
  assign n22082 = ~n22077 & ~n22081 ;
  assign n22083 = ~n22076 & n22082 ;
  assign n22084 = n2432 & ~n22083 ;
  assign n22085 = \P1_DataWidth_reg[1]/NET0131  & \P1_rEIP_reg[31]/NET0131  ;
  assign n22086 = ~\P1_DataWidth_reg[1]/NET0131  & ~n10131 ;
  assign n22087 = n22055 & n22086 ;
  assign n22088 = n18540 & n22087 ;
  assign n22089 = ~n22085 & ~n22088 ;
  assign n22090 = n2436 & ~n22089 ;
  assign n22091 = \P1_PhyAddrPointer_reg[31]/NET0131  & n3028 ;
  assign n22092 = \P1_rEIP_reg[31]/NET0131  & ~n18805 ;
  assign n22093 = ~n22091 & ~n22092 ;
  assign n22094 = ~n22090 & n22093 ;
  assign n22095 = ~n22084 & n22094 ;
  assign n22097 = n10093 & n18541 ;
  assign n22098 = n18540 & ~n22097 ;
  assign n22100 = ~n16282 & n22098 ;
  assign n22099 = n16282 & ~n22098 ;
  assign n22101 = ~\P1_DataWidth_reg[1]/NET0131  & ~n22099 ;
  assign n22102 = ~n22100 & n22101 ;
  assign n22096 = \P1_DataWidth_reg[1]/NET0131  & ~\P1_rEIP_reg[5]/NET0131  ;
  assign n22103 = n2436 & ~n22096 ;
  assign n22104 = ~n22102 & n22103 ;
  assign n22106 = \P1_rEIP_reg[5]/NET0131  & ~n18554 ;
  assign n22107 = ~\P1_rEIP_reg[5]/NET0131  & ~n18560 ;
  assign n22108 = ~n18561 & ~n22107 ;
  assign n22109 = n2425 & ~n22108 ;
  assign n22110 = ~n2311 & n22109 ;
  assign n22111 = ~\P1_EBX_reg[5]/NET0131  & ~n18556 ;
  assign n22112 = ~n22110 & ~n22111 ;
  assign n22113 = n15990 & n22112 ;
  assign n22114 = \P1_EBX_reg[31]/NET0131  & ~n18580 ;
  assign n22116 = ~\P1_EBX_reg[5]/NET0131  & n22114 ;
  assign n22115 = \P1_EBX_reg[5]/NET0131  & ~n22114 ;
  assign n22117 = ~n2425 & ~n22115 ;
  assign n22118 = ~n22116 & n22117 ;
  assign n22119 = ~n22109 & ~n22118 ;
  assign n22120 = n7246 & n22119 ;
  assign n22121 = ~n22113 & ~n22120 ;
  assign n22122 = ~n22106 & n22121 ;
  assign n22123 = n2432 & ~n22122 ;
  assign n22105 = \P1_rEIP_reg[5]/NET0131  & ~n18552 ;
  assign n22124 = \P1_PhyAddrPointer_reg[5]/NET0131  & n3028 ;
  assign n22125 = ~n5092 & ~n22124 ;
  assign n22126 = ~n22105 & n22125 ;
  assign n22127 = ~n22123 & n22126 ;
  assign n22128 = ~n22104 & n22127 ;
  assign n22132 = \P2_EBX_reg[31]/NET0131  & ~n16588 ;
  assign n22134 = ~\P2_EBX_reg[30]/NET0131  & n22132 ;
  assign n22133 = \P2_EBX_reg[30]/NET0131  & ~n22132 ;
  assign n22135 = ~n1920 & ~n22133 ;
  assign n22136 = ~n22134 & n22135 ;
  assign n22129 = ~\P2_rEIP_reg[30]/NET0131  & ~n16550 ;
  assign n22130 = ~n16551 & ~n22129 ;
  assign n22131 = n1920 & ~n22130 ;
  assign n22137 = n10236 & ~n22131 ;
  assign n22138 = ~n22136 & n22137 ;
  assign n22139 = \P2_rEIP_reg[30]/NET0131  & ~n16555 ;
  assign n22141 = n16558 & ~n22130 ;
  assign n22140 = ~\P2_EBX_reg[30]/NET0131  & ~n16558 ;
  assign n22142 = n15980 & ~n22140 ;
  assign n22143 = ~n22141 & n22142 ;
  assign n22144 = ~n22139 & ~n22143 ;
  assign n22145 = ~n22138 & n22144 ;
  assign n22146 = n1927 & ~n22145 ;
  assign n22148 = n8999 & n16518 ;
  assign n22149 = ~n9003 & ~n22148 ;
  assign n22151 = n10029 & ~n22149 ;
  assign n22150 = ~n10029 & n22149 ;
  assign n22152 = ~\P2_DataWidth_reg[1]/NET0131  & ~n22150 ;
  assign n22153 = ~n22151 & n22152 ;
  assign n22147 = \P2_DataWidth_reg[1]/NET0131  & ~\P2_rEIP_reg[30]/NET0131  ;
  assign n22154 = n1931 & ~n22147 ;
  assign n22155 = ~n22153 & n22154 ;
  assign n22156 = \P2_PhyAddrPointer_reg[30]/NET0131  & n2987 ;
  assign n22157 = \P2_rEIP_reg[30]/NET0131  & ~n16511 ;
  assign n22158 = ~n22156 & ~n22157 ;
  assign n22159 = ~n22155 & n22158 ;
  assign n22160 = ~n22146 & n22159 ;
  assign n22162 = ~n8961 & ~n9003 ;
  assign n22163 = ~n19056 & ~n22162 ;
  assign n22165 = ~n16161 & ~n22163 ;
  assign n22164 = n16161 & n22163 ;
  assign n22166 = ~\P2_DataWidth_reg[1]/NET0131  & ~n22164 ;
  assign n22167 = ~n22165 & n22166 ;
  assign n22161 = \P2_DataWidth_reg[1]/NET0131  & ~\P2_rEIP_reg[5]/NET0131  ;
  assign n22168 = n1931 & ~n22161 ;
  assign n22169 = ~n22167 & n22168 ;
  assign n22171 = \P2_rEIP_reg[5]/NET0131  & ~n16555 ;
  assign n22172 = \P2_EBX_reg[31]/NET0131  & ~n16563 ;
  assign n22174 = ~\P2_EBX_reg[5]/NET0131  & n22172 ;
  assign n22173 = \P2_EBX_reg[5]/NET0131  & ~n22172 ;
  assign n22175 = ~n1920 & ~n22173 ;
  assign n22176 = ~n22174 & n22175 ;
  assign n22177 = ~\P2_rEIP_reg[5]/NET0131  & ~n16526 ;
  assign n22178 = ~n20250 & ~n22177 ;
  assign n22179 = n1920 & ~n22178 ;
  assign n22180 = ~n22176 & ~n22179 ;
  assign n22181 = n10236 & n22180 ;
  assign n22182 = ~\P2_EBX_reg[5]/NET0131  & ~n16558 ;
  assign n22183 = n16558 & ~n22178 ;
  assign n22184 = ~n22182 & ~n22183 ;
  assign n22185 = n15980 & n22184 ;
  assign n22186 = ~n22181 & ~n22185 ;
  assign n22187 = ~n22171 & n22186 ;
  assign n22188 = n1927 & ~n22187 ;
  assign n22170 = \P2_rEIP_reg[5]/NET0131  & ~n18989 ;
  assign n22189 = \P2_PhyAddrPointer_reg[5]/NET0131  & n2987 ;
  assign n22190 = ~n3113 & ~n22189 ;
  assign n22191 = ~n22170 & n22190 ;
  assign n22192 = ~n22188 & n22191 ;
  assign n22193 = ~n22169 & n22192 ;
  assign n22194 = n2946 & ~n21326 ;
  assign n22195 = ~n2910 & ~n22194 ;
  assign n22196 = \P3_rEIP_reg[0]/NET0131  & ~n22195 ;
  assign n22197 = ~\P3_InstQueueRd_Addr_reg[0]/NET0131  & n2763 ;
  assign n22198 = n2765 & ~n2946 ;
  assign n22199 = ~n20613 & ~n22198 ;
  assign n22200 = \P3_EBX_reg[0]/NET0131  & ~n22199 ;
  assign n22201 = ~n22197 & ~n22200 ;
  assign n22202 = ~n2815 & ~n22201 ;
  assign n22203 = ~n22196 & ~n22202 ;
  assign n22204 = n2453 & ~n22203 ;
  assign n22205 = ~n2960 & ~n3004 ;
  assign n22206 = \P3_PhyAddrPointer_reg[0]/NET0131  & ~n22205 ;
  assign n22207 = ~n2970 & n20800 ;
  assign n22208 = \P3_rEIP_reg[0]/NET0131  & ~n22207 ;
  assign n22209 = ~n22206 & ~n22208 ;
  assign n22210 = ~n22204 & n22209 ;
  assign n22212 = ~n9054 & n11225 ;
  assign n22213 = ~n21194 & ~n22212 ;
  assign n22215 = n10073 & n22213 ;
  assign n22214 = ~n10073 & ~n22213 ;
  assign n22216 = ~\P3_DataWidth_reg[1]/NET0131  & ~n22214 ;
  assign n22217 = ~n22215 & n22216 ;
  assign n22211 = \P3_DataWidth_reg[1]/NET0131  & ~\P3_rEIP_reg[30]/NET0131  ;
  assign n22218 = n2959 & ~n22211 ;
  assign n22219 = ~n22217 & n22218 ;
  assign n22223 = ~\P3_EBX_reg[26]/NET0131  & ~\P3_EBX_reg[29]/NET0131  ;
  assign n22224 = n21171 & n22223 ;
  assign n22225 = n21063 & n22224 ;
  assign n22226 = \P3_EBX_reg[31]/NET0131  & ~n22225 ;
  assign n22228 = \P3_EBX_reg[30]/NET0131  & ~n22226 ;
  assign n22227 = ~\P3_EBX_reg[30]/NET0131  & n22226 ;
  assign n22229 = ~n2946 & ~n22227 ;
  assign n22230 = ~n22228 & n22229 ;
  assign n22220 = ~\P3_rEIP_reg[30]/NET0131  & ~n21168 ;
  assign n22221 = ~n21248 & ~n22220 ;
  assign n22222 = n2946 & ~n22221 ;
  assign n22231 = n20473 & ~n22222 ;
  assign n22232 = ~n22230 & n22231 ;
  assign n22233 = \P3_rEIP_reg[30]/NET0131  & n2910 ;
  assign n22235 = ~n2786 & n22222 ;
  assign n22234 = ~\P3_EBX_reg[30]/NET0131  & ~n20412 ;
  assign n22236 = n16094 & ~n22234 ;
  assign n22237 = ~n22235 & n22236 ;
  assign n22238 = ~n22233 & ~n22237 ;
  assign n22239 = ~n22232 & n22238 ;
  assign n22240 = n2453 & ~n22239 ;
  assign n22241 = \P3_PhyAddrPointer_reg[30]/NET0131  & n3004 ;
  assign n22242 = \P3_rEIP_reg[30]/NET0131  & ~n20800 ;
  assign n22243 = ~n22241 & ~n22242 ;
  assign n22244 = ~n22240 & n22243 ;
  assign n22245 = ~n22219 & n22244 ;
  assign n22247 = ~n9021 & ~n9054 ;
  assign n22248 = ~n21208 & ~n22247 ;
  assign n22250 = n16209 & n22248 ;
  assign n22249 = ~n16209 & ~n22248 ;
  assign n22251 = ~\P3_DataWidth_reg[1]/NET0131  & ~n22249 ;
  assign n22252 = ~n22250 & n22251 ;
  assign n22246 = \P3_DataWidth_reg[1]/NET0131  & ~\P3_rEIP_reg[5]/NET0131  ;
  assign n22253 = n2959 & ~n22246 ;
  assign n22254 = ~n22252 & n22253 ;
  assign n22257 = ~\P3_rEIP_reg[5]/NET0131  & ~n20416 ;
  assign n22258 = ~n20417 & ~n22257 ;
  assign n22267 = n20412 & ~n22258 ;
  assign n22268 = ~\P3_EBX_reg[5]/NET0131  & ~n20412 ;
  assign n22269 = ~n22267 & ~n22268 ;
  assign n22270 = n16094 & n22269 ;
  assign n22256 = \P3_rEIP_reg[5]/NET0131  & n2910 ;
  assign n22259 = n2946 & ~n22258 ;
  assign n22260 = \P3_EBX_reg[31]/NET0131  & ~n20432 ;
  assign n22262 = ~\P3_EBX_reg[5]/NET0131  & n22260 ;
  assign n22261 = \P3_EBX_reg[5]/NET0131  & ~n22260 ;
  assign n22263 = ~n2946 & ~n22261 ;
  assign n22264 = ~n22262 & n22263 ;
  assign n22265 = ~n22259 & ~n22264 ;
  assign n22266 = n20473 & n22265 ;
  assign n22271 = ~n22256 & ~n22266 ;
  assign n22272 = ~n22270 & n22271 ;
  assign n22273 = n2453 & ~n22272 ;
  assign n22255 = \P3_rEIP_reg[5]/NET0131  & ~n20409 ;
  assign n22274 = \P3_PhyAddrPointer_reg[5]/NET0131  & n3004 ;
  assign n22275 = ~n4412 & ~n22274 ;
  assign n22276 = ~n22255 & n22275 ;
  assign n22277 = ~n22273 & n22276 ;
  assign n22278 = ~n22254 & n22277 ;
  assign n22284 = n2225 & n18556 ;
  assign n22285 = n18554 & ~n22284 ;
  assign n22286 = \P1_rEIP_reg[0]/NET0131  & ~n22285 ;
  assign n22279 = \P1_rEIP_reg[0]/NET0131  & n2425 ;
  assign n22280 = \P1_EBX_reg[0]/NET0131  & ~n2425 ;
  assign n22281 = ~n2301 & n22280 ;
  assign n22282 = ~n22279 & ~n22281 ;
  assign n22283 = n2222 & ~n22282 ;
  assign n22287 = ~\P1_InstQueueRd_Addr_reg[0]/NET0131  & n2231 ;
  assign n22288 = \P1_EBX_reg[0]/NET0131  & ~n18556 ;
  assign n22289 = n2225 & n22288 ;
  assign n22290 = ~n22287 & ~n22289 ;
  assign n22291 = ~n2301 & ~n22290 ;
  assign n22292 = ~n22283 & ~n22291 ;
  assign n22293 = ~n22286 & n22292 ;
  assign n22294 = n2432 & ~n22293 ;
  assign n22295 = ~n2437 & ~n3028 ;
  assign n22296 = \P1_PhyAddrPointer_reg[0]/NET0131  & ~n22295 ;
  assign n22297 = ~n3148 & n18805 ;
  assign n22298 = \P1_rEIP_reg[0]/NET0131  & ~n22297 ;
  assign n22299 = ~n22296 & ~n22298 ;
  assign n22300 = ~n22294 & n22299 ;
  assign n22302 = \datao[27]_pad  & ~n2833 ;
  assign n22303 = \P3_EAX_reg[26]/NET0131  & n16118 ;
  assign n22304 = ~\P3_EAX_reg[27]/NET0131  & ~n22303 ;
  assign n22305 = n16094 & ~n16119 ;
  assign n22306 = ~n22304 & n22305 ;
  assign n22307 = ~n2786 & n22306 ;
  assign n22308 = ~n22302 & ~n22307 ;
  assign n22309 = n2453 & ~n22308 ;
  assign n22301 = \P3_uWord_reg[11]/NET0131  & n16888 ;
  assign n22310 = \datao[27]_pad  & ~n16899 ;
  assign n22311 = ~n22301 & ~n22310 ;
  assign n22312 = ~n22309 & n22311 ;
  assign n22314 = \P1_Datao_reg[27]/NET0131  & ~n2313 ;
  assign n22315 = \P1_EAX_reg[25]/NET0131  & n16022 ;
  assign n22316 = \P1_EAX_reg[26]/NET0131  & n22315 ;
  assign n22317 = ~\P1_EAX_reg[27]/NET0131  & ~n22316 ;
  assign n22318 = n2225 & ~n16023 ;
  assign n22319 = ~n22317 & n22318 ;
  assign n22320 = n2312 & n22319 ;
  assign n22321 = ~n22314 & ~n22320 ;
  assign n22322 = n2432 & ~n22321 ;
  assign n22313 = \P1_uWord_reg[11]/NET0131  & n2440 ;
  assign n22323 = \P1_Datao_reg[27]/NET0131  & ~n16884 ;
  assign n22324 = ~n22313 & ~n22323 ;
  assign n22325 = ~n22322 & n22324 ;
  assign n22327 = \P2_EAX_reg[26]/NET0131  & n15971 ;
  assign n22328 = ~\P2_EAX_reg[27]/NET0131  & ~n22327 ;
  assign n22329 = ~n15972 & ~n22328 ;
  assign n22330 = ~n1819 & ~n22329 ;
  assign n22331 = ~\P2_Datao_reg[27]/NET0131  & n1819 ;
  assign n22332 = n15980 & ~n22331 ;
  assign n22333 = ~n22330 & n22332 ;
  assign n22334 = \P2_Datao_reg[27]/NET0131  & ~n16922 ;
  assign n22335 = ~n22333 & ~n22334 ;
  assign n22336 = n1927 & ~n22335 ;
  assign n22326 = \P2_uWord_reg[11]/NET0131  & n16919 ;
  assign n22337 = \P2_Datao_reg[27]/NET0131  & ~n16936 ;
  assign n22338 = ~n22326 & ~n22337 ;
  assign n22339 = ~n22336 & n22338 ;
  assign n22340 = \P1_EAX_reg[23]/NET0131  & ~n15402 ;
  assign n22345 = ~\P1_EAX_reg[23]/NET0131  & ~n15916 ;
  assign n22346 = \P1_EAX_reg[23]/NET0131  & n15916 ;
  assign n22347 = n2260 & ~n22346 ;
  assign n22348 = ~n22345 & n22347 ;
  assign n22349 = \P1_EAX_reg[23]/NET0131  & ~n15925 ;
  assign n22351 = ~n5224 & n15893 ;
  assign n22341 = n15136 & n15167 ;
  assign n22342 = ~n15168 & ~n22341 ;
  assign n22343 = n2337 & n22342 ;
  assign n22344 = n2331 & n22343 ;
  assign n22350 = ~n5176 & n15932 ;
  assign n22352 = ~n22344 & ~n22350 ;
  assign n22353 = ~n22351 & n22352 ;
  assign n22354 = ~n22349 & n22353 ;
  assign n22355 = ~n22348 & n22354 ;
  assign n22356 = n2432 & ~n22355 ;
  assign n22357 = ~n22340 & ~n22356 ;
  assign n22359 = \P2_lWord_reg[0]/NET0131  & n1805 ;
  assign n22360 = ~n17444 & ~n22359 ;
  assign n22361 = n1742 & ~n22360 ;
  assign n22358 = \P2_lWord_reg[0]/NET0131  & n15981 ;
  assign n22362 = \P2_EAX_reg[0]/NET0131  & n15980 ;
  assign n22363 = ~n22358 & ~n22362 ;
  assign n22364 = ~n22361 & n22363 ;
  assign n22365 = n1927 & ~n22364 ;
  assign n22366 = \P2_lWord_reg[0]/NET0131  & ~n15942 ;
  assign n22367 = ~n22365 & ~n22366 ;
  assign n22368 = \P2_lWord_reg[10]/NET0131  & ~n15942 ;
  assign n22371 = \P2_lWord_reg[10]/NET0131  & n1805 ;
  assign n22372 = ~n16074 & ~n22371 ;
  assign n22373 = n1742 & ~n22372 ;
  assign n22369 = \P2_EAX_reg[10]/NET0131  & n15980 ;
  assign n22370 = \P2_lWord_reg[10]/NET0131  & n15981 ;
  assign n22374 = ~n22369 & ~n22370 ;
  assign n22375 = ~n22373 & n22374 ;
  assign n22376 = n1927 & ~n22375 ;
  assign n22377 = ~n22368 & ~n22376 ;
  assign n22378 = \P2_lWord_reg[11]/NET0131  & ~n15942 ;
  assign n22381 = \P2_lWord_reg[11]/NET0131  & n1805 ;
  assign n22382 = ~n1805 & ~n14069 ;
  assign n22383 = ~n1810 & n22382 ;
  assign n22384 = ~n22381 & ~n22383 ;
  assign n22385 = n1742 & ~n22384 ;
  assign n22379 = \P2_EAX_reg[11]/NET0131  & n15980 ;
  assign n22380 = \P2_lWord_reg[11]/NET0131  & n15981 ;
  assign n22386 = ~n22379 & ~n22380 ;
  assign n22387 = ~n22385 & n22386 ;
  assign n22388 = n1927 & ~n22387 ;
  assign n22389 = ~n22378 & ~n22388 ;
  assign n22390 = \P1_EAX_reg[24]/NET0131  & ~n15402 ;
  assign n22395 = n15924 & ~n22347 ;
  assign n22396 = \P1_EAX_reg[24]/NET0131  & ~n22395 ;
  assign n22403 = ~\P1_EAX_reg[24]/NET0131  & n2260 ;
  assign n22404 = n22346 & n22403 ;
  assign n22397 = \P1_EAX_reg[24]/NET0131  & ~n2377 ;
  assign n22401 = ~n17462 & ~n22397 ;
  assign n22402 = n2222 & ~n22401 ;
  assign n22391 = ~n15168 & n15199 ;
  assign n22392 = ~n15200 & ~n22391 ;
  assign n22393 = n2337 & n22392 ;
  assign n22394 = n2331 & n22393 ;
  assign n22398 = n2377 & ~n5251 ;
  assign n22399 = ~n22397 & ~n22398 ;
  assign n22400 = n2302 & ~n22399 ;
  assign n22405 = ~n22394 & ~n22400 ;
  assign n22406 = ~n22402 & n22405 ;
  assign n22407 = ~n22404 & n22406 ;
  assign n22408 = ~n22396 & n22407 ;
  assign n22409 = n2432 & ~n22408 ;
  assign n22410 = ~n22390 & ~n22409 ;
  assign n22411 = \P2_lWord_reg[12]/NET0131  & ~n15942 ;
  assign n22414 = \P2_lWord_reg[12]/NET0131  & n1805 ;
  assign n22415 = ~n1810 & n15947 ;
  assign n22416 = ~n22414 & ~n22415 ;
  assign n22417 = n1742 & ~n22416 ;
  assign n22412 = \P2_EAX_reg[12]/NET0131  & n15980 ;
  assign n22413 = \P2_lWord_reg[12]/NET0131  & n15981 ;
  assign n22418 = ~n22412 & ~n22413 ;
  assign n22419 = ~n22417 & n22418 ;
  assign n22420 = n1927 & ~n22419 ;
  assign n22421 = ~n22411 & ~n22420 ;
  assign n22422 = \P2_lWord_reg[13]/NET0131  & ~n15942 ;
  assign n22424 = \P2_lWord_reg[13]/NET0131  & n1805 ;
  assign n22425 = ~n17689 & ~n22424 ;
  assign n22426 = n1742 & ~n22425 ;
  assign n22423 = \P2_lWord_reg[13]/NET0131  & n15981 ;
  assign n22427 = \P2_EAX_reg[13]/NET0131  & n15980 ;
  assign n22428 = ~n22423 & ~n22427 ;
  assign n22429 = ~n22426 & n22428 ;
  assign n22430 = n1927 & ~n22429 ;
  assign n22431 = ~n22422 & ~n22430 ;
  assign n22432 = \P2_lWord_reg[14]/NET0131  & ~n15942 ;
  assign n22434 = \P2_lWord_reg[14]/NET0131  & n1805 ;
  assign n22435 = ~n15010 & ~n22434 ;
  assign n22436 = n1742 & ~n22435 ;
  assign n22433 = \P2_lWord_reg[14]/NET0131  & n15981 ;
  assign n22437 = \P2_EAX_reg[14]/NET0131  & n15980 ;
  assign n22438 = ~n22433 & ~n22437 ;
  assign n22439 = ~n22436 & n22438 ;
  assign n22440 = n1927 & ~n22439 ;
  assign n22441 = ~n22432 & ~n22440 ;
  assign n22442 = \P2_lWord_reg[15]/NET0131  & ~n16950 ;
  assign n22443 = n1742 & n16387 ;
  assign n22444 = \P2_EAX_reg[15]/NET0131  & n1743 ;
  assign n22445 = ~n22443 & ~n22444 ;
  assign n22446 = n16959 & ~n22445 ;
  assign n22447 = ~n22442 & ~n22446 ;
  assign n22449 = \P2_lWord_reg[1]/NET0131  & n1805 ;
  assign n22450 = ~n17778 & ~n22449 ;
  assign n22451 = n1742 & ~n22450 ;
  assign n22448 = \P2_lWord_reg[1]/NET0131  & n15981 ;
  assign n22452 = \P2_EAX_reg[1]/NET0131  & n15980 ;
  assign n22453 = ~n22448 & ~n22452 ;
  assign n22454 = ~n22451 & n22453 ;
  assign n22455 = n1927 & ~n22454 ;
  assign n22456 = \P2_lWord_reg[1]/NET0131  & ~n15942 ;
  assign n22457 = ~n22455 & ~n22456 ;
  assign n22459 = n1811 & ~n8589 ;
  assign n22460 = \P2_lWord_reg[2]/NET0131  & n1805 ;
  assign n22461 = ~n22459 & ~n22460 ;
  assign n22462 = n1742 & ~n22461 ;
  assign n22458 = \P2_lWord_reg[2]/NET0131  & n15981 ;
  assign n22463 = \P2_EAX_reg[2]/NET0131  & n15980 ;
  assign n22464 = ~n22458 & ~n22463 ;
  assign n22465 = ~n22462 & n22464 ;
  assign n22466 = n1927 & ~n22465 ;
  assign n22467 = \P2_lWord_reg[2]/NET0131  & ~n15942 ;
  assign n22468 = ~n22466 & ~n22467 ;
  assign n22470 = n1811 & ~n5298 ;
  assign n22471 = \P2_lWord_reg[3]/NET0131  & n1805 ;
  assign n22472 = ~n22470 & ~n22471 ;
  assign n22473 = n1742 & ~n22472 ;
  assign n22469 = \P2_lWord_reg[3]/NET0131  & n15981 ;
  assign n22474 = \P2_EAX_reg[3]/NET0131  & n15980 ;
  assign n22475 = ~n22469 & ~n22474 ;
  assign n22476 = ~n22473 & n22475 ;
  assign n22477 = n1927 & ~n22476 ;
  assign n22478 = \P2_lWord_reg[3]/NET0131  & ~n15942 ;
  assign n22479 = ~n22477 & ~n22478 ;
  assign n22481 = \P2_lWord_reg[4]/NET0131  & n1805 ;
  assign n22482 = ~n21755 & ~n22481 ;
  assign n22483 = n1742 & ~n22482 ;
  assign n22480 = \P2_lWord_reg[4]/NET0131  & n15981 ;
  assign n22484 = \P2_EAX_reg[4]/NET0131  & n15980 ;
  assign n22485 = ~n22480 & ~n22484 ;
  assign n22486 = ~n22483 & n22485 ;
  assign n22487 = n1927 & ~n22486 ;
  assign n22488 = \P2_lWord_reg[4]/NET0131  & ~n15942 ;
  assign n22489 = ~n22487 & ~n22488 ;
  assign n22491 = n1811 & ~n10333 ;
  assign n22492 = \P2_lWord_reg[5]/NET0131  & n1805 ;
  assign n22493 = ~n22491 & ~n22492 ;
  assign n22494 = n1742 & ~n22493 ;
  assign n22490 = \P2_lWord_reg[5]/NET0131  & n15981 ;
  assign n22495 = \P2_EAX_reg[5]/NET0131  & n15980 ;
  assign n22496 = ~n22490 & ~n22495 ;
  assign n22497 = ~n22494 & n22496 ;
  assign n22498 = n1927 & ~n22497 ;
  assign n22499 = \P2_lWord_reg[5]/NET0131  & ~n15942 ;
  assign n22500 = ~n22498 & ~n22499 ;
  assign n22503 = \P2_lWord_reg[6]/NET0131  & n1805 ;
  assign n22504 = ~n1805 & ~n7724 ;
  assign n22505 = ~n1810 & n22504 ;
  assign n22506 = ~n22503 & ~n22505 ;
  assign n22507 = n1742 & ~n22506 ;
  assign n22501 = \P2_EAX_reg[6]/NET0131  & n15980 ;
  assign n22502 = \P2_lWord_reg[6]/NET0131  & n15981 ;
  assign n22508 = ~n22501 & ~n22502 ;
  assign n22509 = ~n22507 & n22508 ;
  assign n22510 = n1927 & ~n22509 ;
  assign n22511 = \P2_lWord_reg[6]/NET0131  & ~n15942 ;
  assign n22512 = ~n22510 & ~n22511 ;
  assign n22514 = \P2_lWord_reg[7]/NET0131  & n1805 ;
  assign n22515 = n1811 & ~n3128 ;
  assign n22516 = ~n22514 & ~n22515 ;
  assign n22517 = n1742 & ~n22516 ;
  assign n22513 = \P2_lWord_reg[7]/NET0131  & n15981 ;
  assign n22518 = \P2_EAX_reg[7]/NET0131  & n15980 ;
  assign n22519 = ~n22513 & ~n22518 ;
  assign n22520 = ~n22517 & n22519 ;
  assign n22521 = n1927 & ~n22520 ;
  assign n22522 = \P2_lWord_reg[7]/NET0131  & ~n15942 ;
  assign n22523 = ~n22521 & ~n22522 ;
  assign n22524 = \P2_lWord_reg[8]/NET0131  & ~n15942 ;
  assign n22527 = ~n1810 & n16956 ;
  assign n22528 = \P2_lWord_reg[8]/NET0131  & n1805 ;
  assign n22529 = ~n22527 & ~n22528 ;
  assign n22530 = n1742 & ~n22529 ;
  assign n22525 = \P2_EAX_reg[8]/NET0131  & n15980 ;
  assign n22526 = \P2_lWord_reg[8]/NET0131  & n15981 ;
  assign n22531 = ~n22525 & ~n22526 ;
  assign n22532 = ~n22530 & n22531 ;
  assign n22533 = n1927 & ~n22532 ;
  assign n22534 = ~n22524 & ~n22533 ;
  assign n22535 = \P2_lWord_reg[9]/NET0131  & ~n15942 ;
  assign n22537 = \P2_lWord_reg[9]/NET0131  & n1805 ;
  assign n22538 = ~n17935 & ~n22537 ;
  assign n22539 = n1742 & ~n22538 ;
  assign n22536 = \P2_lWord_reg[9]/NET0131  & n15981 ;
  assign n22540 = \P2_EAX_reg[9]/NET0131  & n15980 ;
  assign n22541 = ~n22536 & ~n22540 ;
  assign n22542 = ~n22539 & n22541 ;
  assign n22543 = n1927 & ~n22542 ;
  assign n22544 = ~n22535 & ~n22543 ;
  assign n22545 = \P2_uWord_reg[11]/NET0131  & ~n16950 ;
  assign n22546 = n1743 & n22329 ;
  assign n22547 = n1742 & n22382 ;
  assign n22548 = ~n22546 & ~n22547 ;
  assign n22549 = n16959 & ~n22548 ;
  assign n22550 = ~n22545 & ~n22549 ;
  assign n22551 = \P1_uWord_reg[11]/NET0131  & ~n15994 ;
  assign n22552 = ~n5170 & n15996 ;
  assign n22553 = ~n22319 & ~n22552 ;
  assign n22554 = n16029 & ~n22553 ;
  assign n22555 = ~n22551 & ~n22554 ;
  assign n22556 = \P1_EAX_reg[28]/NET0131  & ~n15402 ;
  assign n22558 = ~\P1_EAX_reg[28]/NET0131  & ~n16319 ;
  assign n22559 = n2260 & ~n16320 ;
  assign n22560 = ~n22558 & n22559 ;
  assign n22561 = n2222 & ~n2377 ;
  assign n22562 = n15924 & ~n22561 ;
  assign n22563 = \P1_EAX_reg[28]/NET0131  & ~n22562 ;
  assign n22564 = ~n15296 & n15327 ;
  assign n22565 = n2337 & ~n15328 ;
  assign n22566 = ~n22564 & n22565 ;
  assign n22567 = n2331 & n22566 ;
  assign n22557 = n2222 & n18169 ;
  assign n22569 = n2377 & n5267 ;
  assign n22568 = ~\P1_EAX_reg[28]/NET0131  & ~n2377 ;
  assign n22570 = n2302 & ~n22568 ;
  assign n22571 = ~n22569 & n22570 ;
  assign n22572 = ~n22557 & ~n22571 ;
  assign n22573 = ~n22567 & n22572 ;
  assign n22574 = ~n22563 & n22573 ;
  assign n22575 = ~n22560 & n22574 ;
  assign n22576 = n2432 & ~n22575 ;
  assign n22577 = ~n22556 & ~n22576 ;
  assign n22578 = \P3_EAX_reg[0]/NET0131  & ~n17124 ;
  assign n22580 = \buf2_reg[0]/NET0131  & n2857 ;
  assign n22579 = ~n3963 & n13812 ;
  assign n22581 = ~n17263 & ~n22579 ;
  assign n22582 = ~n22580 & n22581 ;
  assign n22583 = n2453 & ~n22582 ;
  assign n22584 = ~n22578 & ~n22583 ;
  assign n22585 = \P3_EAX_reg[16]/NET0131  & ~n13810 ;
  assign n22621 = ~n13816 & ~n17211 ;
  assign n22622 = \P3_EAX_reg[16]/NET0131  & ~n22621 ;
  assign n22618 = \P3_EAX_reg[16]/NET0131  & n14031 ;
  assign n22619 = n13813 & ~n22618 ;
  assign n22620 = n14031 & n22619 ;
  assign n22623 = \P3_EAX_reg[16]/NET0131  & ~n2862 ;
  assign n22627 = \buf2_reg[0]/NET0131  & n2862 ;
  assign n22628 = ~n22623 & ~n22627 ;
  assign n22629 = n2821 & ~n22628 ;
  assign n22590 = \P3_InstQueue_reg[13][0]/NET0131  & n2464 ;
  assign n22591 = \P3_InstQueue_reg[15][0]/NET0131  & n2472 ;
  assign n22604 = ~n22590 & ~n22591 ;
  assign n22592 = \P3_InstQueue_reg[7][0]/NET0131  & n2469 ;
  assign n22593 = \P3_InstQueue_reg[11][0]/NET0131  & n2476 ;
  assign n22605 = ~n22592 & ~n22593 ;
  assign n22612 = n22604 & n22605 ;
  assign n22586 = \P3_InstQueue_reg[12][0]/NET0131  & n2490 ;
  assign n22587 = \P3_InstQueue_reg[3][0]/NET0131  & n2482 ;
  assign n22602 = ~n22586 & ~n22587 ;
  assign n22588 = \P3_InstQueue_reg[6][0]/NET0131  & n2480 ;
  assign n22589 = \P3_InstQueue_reg[0][0]/NET0131  & n2478 ;
  assign n22603 = ~n22588 & ~n22589 ;
  assign n22613 = n22602 & n22603 ;
  assign n22614 = n22612 & n22613 ;
  assign n22598 = \P3_InstQueue_reg[10][0]/NET0131  & n2460 ;
  assign n22599 = \P3_InstQueue_reg[14][0]/NET0131  & n2486 ;
  assign n22608 = ~n22598 & ~n22599 ;
  assign n22600 = \P3_InstQueue_reg[9][0]/NET0131  & n2474 ;
  assign n22601 = \P3_InstQueue_reg[5][0]/NET0131  & n2466 ;
  assign n22609 = ~n22600 & ~n22601 ;
  assign n22610 = n22608 & n22609 ;
  assign n22594 = \P3_InstQueue_reg[8][0]/NET0131  & n2492 ;
  assign n22595 = \P3_InstQueue_reg[2][0]/NET0131  & n2484 ;
  assign n22606 = ~n22594 & ~n22595 ;
  assign n22596 = \P3_InstQueue_reg[1][0]/NET0131  & n2488 ;
  assign n22597 = \P3_InstQueue_reg[4][0]/NET0131  & n2456 ;
  assign n22607 = ~n22596 & ~n22597 ;
  assign n22611 = n22606 & n22607 ;
  assign n22615 = n22610 & n22611 ;
  assign n22616 = n22614 & n22615 ;
  assign n22617 = n13812 & ~n22616 ;
  assign n22624 = \buf2_reg[16]/NET0131  & n2862 ;
  assign n22625 = ~n22623 & ~n22624 ;
  assign n22626 = n2820 & ~n22625 ;
  assign n22630 = ~n22617 & ~n22626 ;
  assign n22631 = ~n22629 & n22630 ;
  assign n22632 = ~n22620 & n22631 ;
  assign n22633 = ~n22622 & n22632 ;
  assign n22634 = n2453 & ~n22633 ;
  assign n22635 = ~n22585 & ~n22634 ;
  assign n22636 = \P3_EAX_reg[17]/NET0131  & ~n13810 ;
  assign n22637 = n14922 & ~n22619 ;
  assign n22638 = \P3_EAX_reg[17]/NET0131  & ~n22637 ;
  assign n22639 = ~\P3_EAX_reg[17]/NET0131  & n13813 ;
  assign n22640 = n22618 & n22639 ;
  assign n22645 = \P3_InstQueue_reg[1][1]/NET0131  & n2488 ;
  assign n22646 = \P3_InstQueue_reg[4][1]/NET0131  & n2456 ;
  assign n22659 = ~n22645 & ~n22646 ;
  assign n22647 = \P3_InstQueue_reg[13][1]/NET0131  & n2464 ;
  assign n22648 = \P3_InstQueue_reg[12][1]/NET0131  & n2490 ;
  assign n22660 = ~n22647 & ~n22648 ;
  assign n22667 = n22659 & n22660 ;
  assign n22641 = \P3_InstQueue_reg[6][1]/NET0131  & n2480 ;
  assign n22642 = \P3_InstQueue_reg[11][1]/NET0131  & n2476 ;
  assign n22657 = ~n22641 & ~n22642 ;
  assign n22643 = \P3_InstQueue_reg[15][1]/NET0131  & n2472 ;
  assign n22644 = \P3_InstQueue_reg[14][1]/NET0131  & n2486 ;
  assign n22658 = ~n22643 & ~n22644 ;
  assign n22668 = n22657 & n22658 ;
  assign n22669 = n22667 & n22668 ;
  assign n22653 = \P3_InstQueue_reg[9][1]/NET0131  & n2474 ;
  assign n22654 = \P3_InstQueue_reg[5][1]/NET0131  & n2466 ;
  assign n22663 = ~n22653 & ~n22654 ;
  assign n22655 = \P3_InstQueue_reg[2][1]/NET0131  & n2484 ;
  assign n22656 = \P3_InstQueue_reg[3][1]/NET0131  & n2482 ;
  assign n22664 = ~n22655 & ~n22656 ;
  assign n22665 = n22663 & n22664 ;
  assign n22649 = \P3_InstQueue_reg[8][1]/NET0131  & n2492 ;
  assign n22650 = \P3_InstQueue_reg[10][1]/NET0131  & n2460 ;
  assign n22661 = ~n22649 & ~n22650 ;
  assign n22651 = \P3_InstQueue_reg[0][1]/NET0131  & n2478 ;
  assign n22652 = \P3_InstQueue_reg[7][1]/NET0131  & n2469 ;
  assign n22662 = ~n22651 & ~n22652 ;
  assign n22666 = n22661 & n22662 ;
  assign n22670 = n22665 & n22666 ;
  assign n22671 = n22669 & n22670 ;
  assign n22672 = n13812 & ~n22671 ;
  assign n22673 = \buf2_reg[1]/NET0131  & n2821 ;
  assign n22674 = \buf2_reg[17]/NET0131  & n2820 ;
  assign n22675 = ~n22673 & ~n22674 ;
  assign n22676 = n2862 & ~n22675 ;
  assign n22677 = ~n22672 & ~n22676 ;
  assign n22678 = ~n22640 & n22677 ;
  assign n22679 = ~n22638 & n22678 ;
  assign n22680 = n2453 & ~n22679 ;
  assign n22681 = ~n22636 & ~n22680 ;
  assign n22682 = n2453 & n13816 ;
  assign n22683 = n13810 & ~n22682 ;
  assign n22684 = \P3_EAX_reg[18]/NET0131  & ~n22683 ;
  assign n22724 = \P3_EAX_reg[17]/NET0131  & n22618 ;
  assign n22725 = ~\P3_EAX_reg[18]/NET0131  & ~n22724 ;
  assign n22726 = n13813 & ~n14034 ;
  assign n22727 = ~n22725 & n22726 ;
  assign n22686 = \P3_EAX_reg[18]/NET0131  & ~n2862 ;
  assign n22721 = \buf2_reg[18]/NET0131  & n2862 ;
  assign n22722 = ~n22686 & ~n22721 ;
  assign n22723 = n2820 & ~n22722 ;
  assign n22685 = \buf2_reg[2]/NET0131  & n2862 ;
  assign n22687 = ~n22685 & ~n22686 ;
  assign n22688 = n2821 & ~n22687 ;
  assign n22693 = \P3_InstQueue_reg[6][2]/NET0131  & n2480 ;
  assign n22694 = \P3_InstQueue_reg[5][2]/NET0131  & n2466 ;
  assign n22707 = ~n22693 & ~n22694 ;
  assign n22695 = \P3_InstQueue_reg[9][2]/NET0131  & n2474 ;
  assign n22696 = \P3_InstQueue_reg[4][2]/NET0131  & n2456 ;
  assign n22708 = ~n22695 & ~n22696 ;
  assign n22715 = n22707 & n22708 ;
  assign n22689 = \P3_InstQueue_reg[1][2]/NET0131  & n2488 ;
  assign n22690 = \P3_InstQueue_reg[8][2]/NET0131  & n2492 ;
  assign n22705 = ~n22689 & ~n22690 ;
  assign n22691 = \P3_InstQueue_reg[11][2]/NET0131  & n2476 ;
  assign n22692 = \P3_InstQueue_reg[10][2]/NET0131  & n2460 ;
  assign n22706 = ~n22691 & ~n22692 ;
  assign n22716 = n22705 & n22706 ;
  assign n22717 = n22715 & n22716 ;
  assign n22701 = \P3_InstQueue_reg[12][2]/NET0131  & n2490 ;
  assign n22702 = \P3_InstQueue_reg[13][2]/NET0131  & n2464 ;
  assign n22711 = ~n22701 & ~n22702 ;
  assign n22703 = \P3_InstQueue_reg[2][2]/NET0131  & n2484 ;
  assign n22704 = \P3_InstQueue_reg[0][2]/NET0131  & n2478 ;
  assign n22712 = ~n22703 & ~n22704 ;
  assign n22713 = n22711 & n22712 ;
  assign n22697 = \P3_InstQueue_reg[7][2]/NET0131  & n2469 ;
  assign n22698 = \P3_InstQueue_reg[14][2]/NET0131  & n2486 ;
  assign n22709 = ~n22697 & ~n22698 ;
  assign n22699 = \P3_InstQueue_reg[3][2]/NET0131  & n2482 ;
  assign n22700 = \P3_InstQueue_reg[15][2]/NET0131  & n2472 ;
  assign n22710 = ~n22699 & ~n22700 ;
  assign n22714 = n22709 & n22710 ;
  assign n22718 = n22713 & n22714 ;
  assign n22719 = n22717 & n22718 ;
  assign n22720 = n13812 & ~n22719 ;
  assign n22728 = ~n22688 & ~n22720 ;
  assign n22729 = ~n22723 & n22728 ;
  assign n22730 = ~n22727 & n22729 ;
  assign n22731 = n2453 & ~n22730 ;
  assign n22732 = ~n22684 & ~n22731 ;
  assign n22733 = \P3_EAX_reg[19]/NET0131  & ~n13810 ;
  assign n22735 = ~\P3_EAX_reg[19]/NET0131  & ~n14034 ;
  assign n22736 = n13813 & ~n14035 ;
  assign n22737 = ~n22735 & n22736 ;
  assign n22734 = \P3_EAX_reg[19]/NET0131  & ~n14922 ;
  assign n22742 = \P3_InstQueue_reg[13][3]/NET0131  & n2464 ;
  assign n22743 = \P3_InstQueue_reg[15][3]/NET0131  & n2472 ;
  assign n22756 = ~n22742 & ~n22743 ;
  assign n22744 = \P3_InstQueue_reg[7][3]/NET0131  & n2469 ;
  assign n22745 = \P3_InstQueue_reg[11][3]/NET0131  & n2476 ;
  assign n22757 = ~n22744 & ~n22745 ;
  assign n22764 = n22756 & n22757 ;
  assign n22738 = \P3_InstQueue_reg[12][3]/NET0131  & n2490 ;
  assign n22739 = \P3_InstQueue_reg[3][3]/NET0131  & n2482 ;
  assign n22754 = ~n22738 & ~n22739 ;
  assign n22740 = \P3_InstQueue_reg[6][3]/NET0131  & n2480 ;
  assign n22741 = \P3_InstQueue_reg[0][3]/NET0131  & n2478 ;
  assign n22755 = ~n22740 & ~n22741 ;
  assign n22765 = n22754 & n22755 ;
  assign n22766 = n22764 & n22765 ;
  assign n22750 = \P3_InstQueue_reg[10][3]/NET0131  & n2460 ;
  assign n22751 = \P3_InstQueue_reg[14][3]/NET0131  & n2486 ;
  assign n22760 = ~n22750 & ~n22751 ;
  assign n22752 = \P3_InstQueue_reg[9][3]/NET0131  & n2474 ;
  assign n22753 = \P3_InstQueue_reg[5][3]/NET0131  & n2466 ;
  assign n22761 = ~n22752 & ~n22753 ;
  assign n22762 = n22760 & n22761 ;
  assign n22746 = \P3_InstQueue_reg[8][3]/NET0131  & n2492 ;
  assign n22747 = \P3_InstQueue_reg[2][3]/NET0131  & n2484 ;
  assign n22758 = ~n22746 & ~n22747 ;
  assign n22748 = \P3_InstQueue_reg[1][3]/NET0131  & n2488 ;
  assign n22749 = \P3_InstQueue_reg[4][3]/NET0131  & n2456 ;
  assign n22759 = ~n22748 & ~n22749 ;
  assign n22763 = n22758 & n22759 ;
  assign n22767 = n22762 & n22763 ;
  assign n22768 = n22766 & n22767 ;
  assign n22769 = n13812 & ~n22768 ;
  assign n22770 = \buf2_reg[19]/NET0131  & n2820 ;
  assign n22771 = \buf2_reg[3]/NET0131  & n2821 ;
  assign n22772 = ~n22770 & ~n22771 ;
  assign n22773 = n2862 & ~n22772 ;
  assign n22774 = ~n22769 & ~n22773 ;
  assign n22775 = ~n22734 & n22774 ;
  assign n22776 = ~n22737 & n22775 ;
  assign n22777 = n2453 & ~n22776 ;
  assign n22778 = ~n22733 & ~n22777 ;
  assign n22779 = ~n2864 & ~n13816 ;
  assign n22780 = n2453 & ~n22779 ;
  assign n22781 = n13810 & ~n22780 ;
  assign n22782 = \P3_EAX_reg[20]/NET0131  & ~n22781 ;
  assign n22815 = ~\P3_EAX_reg[20]/NET0131  & ~n14035 ;
  assign n22816 = n13813 & ~n14036 ;
  assign n22817 = ~n22815 & n22816 ;
  assign n22818 = \P3_EAX_reg[20]/NET0131  & ~n2862 ;
  assign n22819 = ~n21812 & ~n22818 ;
  assign n22820 = n2821 & ~n22819 ;
  assign n22787 = \P3_InstQueue_reg[6][4]/NET0131  & n2480 ;
  assign n22788 = \P3_InstQueue_reg[5][4]/NET0131  & n2466 ;
  assign n22801 = ~n22787 & ~n22788 ;
  assign n22789 = \P3_InstQueue_reg[9][4]/NET0131  & n2474 ;
  assign n22790 = \P3_InstQueue_reg[4][4]/NET0131  & n2456 ;
  assign n22802 = ~n22789 & ~n22790 ;
  assign n22809 = n22801 & n22802 ;
  assign n22783 = \P3_InstQueue_reg[1][4]/NET0131  & n2488 ;
  assign n22784 = \P3_InstQueue_reg[8][4]/NET0131  & n2492 ;
  assign n22799 = ~n22783 & ~n22784 ;
  assign n22785 = \P3_InstQueue_reg[11][4]/NET0131  & n2476 ;
  assign n22786 = \P3_InstQueue_reg[10][4]/NET0131  & n2460 ;
  assign n22800 = ~n22785 & ~n22786 ;
  assign n22810 = n22799 & n22800 ;
  assign n22811 = n22809 & n22810 ;
  assign n22795 = \P3_InstQueue_reg[12][4]/NET0131  & n2490 ;
  assign n22796 = \P3_InstQueue_reg[13][4]/NET0131  & n2464 ;
  assign n22805 = ~n22795 & ~n22796 ;
  assign n22797 = \P3_InstQueue_reg[2][4]/NET0131  & n2484 ;
  assign n22798 = \P3_InstQueue_reg[0][4]/NET0131  & n2478 ;
  assign n22806 = ~n22797 & ~n22798 ;
  assign n22807 = n22805 & n22806 ;
  assign n22791 = \P3_InstQueue_reg[7][4]/NET0131  & n2469 ;
  assign n22792 = \P3_InstQueue_reg[14][4]/NET0131  & n2486 ;
  assign n22803 = ~n22791 & ~n22792 ;
  assign n22793 = \P3_InstQueue_reg[3][4]/NET0131  & n2482 ;
  assign n22794 = \P3_InstQueue_reg[15][4]/NET0131  & n2472 ;
  assign n22804 = ~n22793 & ~n22794 ;
  assign n22808 = n22803 & n22804 ;
  assign n22812 = n22807 & n22808 ;
  assign n22813 = n22811 & n22812 ;
  assign n22814 = n13812 & ~n22813 ;
  assign n22821 = \buf2_reg[20]/NET0131  & n2820 ;
  assign n22822 = n2862 & n22821 ;
  assign n22823 = ~n22814 & ~n22822 ;
  assign n22824 = ~n22820 & n22823 ;
  assign n22825 = ~n22817 & n22824 ;
  assign n22826 = n2453 & ~n22825 ;
  assign n22827 = ~n22782 & ~n22826 ;
  assign n22828 = \P3_EAX_reg[21]/NET0131  & ~n13810 ;
  assign n22830 = ~\P3_EAX_reg[21]/NET0131  & ~n14036 ;
  assign n22831 = n13813 & ~n14037 ;
  assign n22832 = ~n22830 & n22831 ;
  assign n22829 = \P3_EAX_reg[21]/NET0131  & ~n14922 ;
  assign n22837 = \P3_InstQueue_reg[13][5]/NET0131  & n2464 ;
  assign n22838 = \P3_InstQueue_reg[15][5]/NET0131  & n2472 ;
  assign n22851 = ~n22837 & ~n22838 ;
  assign n22839 = \P3_InstQueue_reg[7][5]/NET0131  & n2469 ;
  assign n22840 = \P3_InstQueue_reg[11][5]/NET0131  & n2476 ;
  assign n22852 = ~n22839 & ~n22840 ;
  assign n22859 = n22851 & n22852 ;
  assign n22833 = \P3_InstQueue_reg[12][5]/NET0131  & n2490 ;
  assign n22834 = \P3_InstQueue_reg[3][5]/NET0131  & n2482 ;
  assign n22849 = ~n22833 & ~n22834 ;
  assign n22835 = \P3_InstQueue_reg[6][5]/NET0131  & n2480 ;
  assign n22836 = \P3_InstQueue_reg[0][5]/NET0131  & n2478 ;
  assign n22850 = ~n22835 & ~n22836 ;
  assign n22860 = n22849 & n22850 ;
  assign n22861 = n22859 & n22860 ;
  assign n22845 = \P3_InstQueue_reg[10][5]/NET0131  & n2460 ;
  assign n22846 = \P3_InstQueue_reg[14][5]/NET0131  & n2486 ;
  assign n22855 = ~n22845 & ~n22846 ;
  assign n22847 = \P3_InstQueue_reg[9][5]/NET0131  & n2474 ;
  assign n22848 = \P3_InstQueue_reg[5][5]/NET0131  & n2466 ;
  assign n22856 = ~n22847 & ~n22848 ;
  assign n22857 = n22855 & n22856 ;
  assign n22841 = \P3_InstQueue_reg[8][5]/NET0131  & n2492 ;
  assign n22842 = \P3_InstQueue_reg[2][5]/NET0131  & n2484 ;
  assign n22853 = ~n22841 & ~n22842 ;
  assign n22843 = \P3_InstQueue_reg[1][5]/NET0131  & n2488 ;
  assign n22844 = \P3_InstQueue_reg[4][5]/NET0131  & n2456 ;
  assign n22854 = ~n22843 & ~n22844 ;
  assign n22858 = n22853 & n22854 ;
  assign n22862 = n22857 & n22858 ;
  assign n22863 = n22861 & n22862 ;
  assign n22864 = n13812 & ~n22863 ;
  assign n22865 = \buf2_reg[21]/NET0131  & n2820 ;
  assign n22866 = \buf2_reg[5]/NET0131  & n2821 ;
  assign n22867 = ~n22865 & ~n22866 ;
  assign n22868 = n2862 & ~n22867 ;
  assign n22869 = ~n22864 & ~n22868 ;
  assign n22870 = ~n22829 & n22869 ;
  assign n22871 = ~n22832 & n22870 ;
  assign n22872 = n2453 & ~n22871 ;
  assign n22873 = ~n22828 & ~n22872 ;
  assign n22874 = \P3_EAX_reg[22]/NET0131  & ~n22683 ;
  assign n22907 = ~\P3_EAX_reg[22]/NET0131  & ~n14037 ;
  assign n22908 = \P3_EAX_reg[22]/NET0131  & n14037 ;
  assign n22909 = n13813 & ~n22908 ;
  assign n22910 = ~n22907 & n22909 ;
  assign n22911 = \P3_EAX_reg[22]/NET0131  & ~n2862 ;
  assign n22915 = \buf2_reg[6]/NET0131  & n2862 ;
  assign n22916 = ~n22911 & ~n22915 ;
  assign n22917 = n2821 & ~n22916 ;
  assign n22879 = \P3_InstQueue_reg[5][6]/NET0131  & n2466 ;
  assign n22880 = \P3_InstQueue_reg[7][6]/NET0131  & n2469 ;
  assign n22893 = ~n22879 & ~n22880 ;
  assign n22881 = \P3_InstQueue_reg[8][6]/NET0131  & n2492 ;
  assign n22882 = \P3_InstQueue_reg[15][6]/NET0131  & n2472 ;
  assign n22894 = ~n22881 & ~n22882 ;
  assign n22901 = n22893 & n22894 ;
  assign n22875 = \P3_InstQueue_reg[9][6]/NET0131  & n2474 ;
  assign n22876 = \P3_InstQueue_reg[0][6]/NET0131  & n2478 ;
  assign n22891 = ~n22875 & ~n22876 ;
  assign n22877 = \P3_InstQueue_reg[1][6]/NET0131  & n2488 ;
  assign n22878 = \P3_InstQueue_reg[3][6]/NET0131  & n2482 ;
  assign n22892 = ~n22877 & ~n22878 ;
  assign n22902 = n22891 & n22892 ;
  assign n22903 = n22901 & n22902 ;
  assign n22887 = \P3_InstQueue_reg[14][6]/NET0131  & n2486 ;
  assign n22888 = \P3_InstQueue_reg[10][6]/NET0131  & n2460 ;
  assign n22897 = ~n22887 & ~n22888 ;
  assign n22889 = \P3_InstQueue_reg[13][6]/NET0131  & n2464 ;
  assign n22890 = \P3_InstQueue_reg[4][6]/NET0131  & n2456 ;
  assign n22898 = ~n22889 & ~n22890 ;
  assign n22899 = n22897 & n22898 ;
  assign n22883 = \P3_InstQueue_reg[11][6]/NET0131  & n2476 ;
  assign n22884 = \P3_InstQueue_reg[2][6]/NET0131  & n2484 ;
  assign n22895 = ~n22883 & ~n22884 ;
  assign n22885 = \P3_InstQueue_reg[6][6]/NET0131  & n2480 ;
  assign n22886 = \P3_InstQueue_reg[12][6]/NET0131  & n2490 ;
  assign n22896 = ~n22885 & ~n22886 ;
  assign n22900 = n22895 & n22896 ;
  assign n22904 = n22899 & n22900 ;
  assign n22905 = n22903 & n22904 ;
  assign n22906 = n13812 & ~n22905 ;
  assign n22912 = \buf2_reg[22]/NET0131  & n2862 ;
  assign n22913 = ~n22911 & ~n22912 ;
  assign n22914 = n2820 & ~n22913 ;
  assign n22918 = ~n22906 & ~n22914 ;
  assign n22919 = ~n22917 & n22918 ;
  assign n22920 = ~n22910 & n22919 ;
  assign n22921 = n2453 & ~n22920 ;
  assign n22922 = ~n22874 & ~n22921 ;
  assign n22923 = \P3_EAX_reg[23]/NET0131  & ~n13810 ;
  assign n22927 = ~n13816 & ~n22909 ;
  assign n22928 = \P3_EAX_reg[23]/NET0131  & ~n22927 ;
  assign n22936 = ~\P3_EAX_reg[23]/NET0131  & n13813 ;
  assign n22937 = n22908 & n22936 ;
  assign n22929 = \P3_EAX_reg[23]/NET0131  & ~n2862 ;
  assign n22933 = \buf2_reg[7]/NET0131  & n2862 ;
  assign n22934 = ~n22929 & ~n22933 ;
  assign n22935 = n2821 & ~n22934 ;
  assign n22924 = n13849 & n13880 ;
  assign n22925 = ~n13881 & ~n22924 ;
  assign n22926 = n13812 & n22925 ;
  assign n22930 = \buf2_reg[23]/NET0131  & n2862 ;
  assign n22931 = ~n22929 & ~n22930 ;
  assign n22932 = n2820 & ~n22931 ;
  assign n22938 = ~n22926 & ~n22932 ;
  assign n22939 = ~n22935 & n22938 ;
  assign n22940 = ~n22937 & n22939 ;
  assign n22941 = ~n22928 & n22940 ;
  assign n22942 = n2453 & ~n22941 ;
  assign n22943 = ~n22923 & ~n22942 ;
  assign n22944 = \P3_EAX_reg[24]/NET0131  & ~n13810 ;
  assign n22948 = \P3_EAX_reg[23]/NET0131  & n22908 ;
  assign n22949 = n13813 & ~n22948 ;
  assign n22950 = ~n13816 & ~n22949 ;
  assign n22951 = \P3_EAX_reg[24]/NET0131  & ~n22950 ;
  assign n22959 = ~\P3_EAX_reg[24]/NET0131  & n13813 ;
  assign n22960 = n22948 & n22959 ;
  assign n22952 = \P3_EAX_reg[24]/NET0131  & ~n2862 ;
  assign n22956 = \buf2_reg[8]/NET0131  & n2862 ;
  assign n22957 = ~n22952 & ~n22956 ;
  assign n22958 = n2821 & ~n22957 ;
  assign n22945 = ~n13881 & n13912 ;
  assign n22946 = ~n13913 & ~n22945 ;
  assign n22947 = n13812 & n22946 ;
  assign n22953 = \buf2_reg[24]/NET0131  & n2862 ;
  assign n22954 = ~n22952 & ~n22953 ;
  assign n22955 = n2820 & ~n22954 ;
  assign n22961 = ~n22947 & ~n22955 ;
  assign n22962 = ~n22958 & n22961 ;
  assign n22963 = ~n22960 & n22962 ;
  assign n22964 = ~n22951 & n22963 ;
  assign n22965 = n2453 & ~n22964 ;
  assign n22966 = ~n22944 & ~n22965 ;
  assign n22967 = \P3_EAX_reg[28]/NET0131  & ~n13810 ;
  assign n22968 = ~n14046 & n14922 ;
  assign n22969 = \P3_EAX_reg[28]/NET0131  & ~n22968 ;
  assign n22970 = ~\P3_EAX_reg[28]/NET0131  & n13813 ;
  assign n22971 = n14045 & n22970 ;
  assign n22972 = ~n14010 & n14855 ;
  assign n22973 = ~n14856 & ~n22972 ;
  assign n22974 = n13812 & n22973 ;
  assign n22975 = \buf2_reg[12]/NET0131  & n2821 ;
  assign n22976 = \buf2_reg[28]/NET0131  & n2820 ;
  assign n22977 = ~n22975 & ~n22976 ;
  assign n22978 = n2862 & ~n22977 ;
  assign n22979 = ~n22974 & ~n22978 ;
  assign n22980 = ~n22971 & n22979 ;
  assign n22981 = ~n22969 & n22980 ;
  assign n22982 = n2453 & ~n22981 ;
  assign n22983 = ~n22967 & ~n22982 ;
  assign n22984 = n2453 & ~n2914 ;
  assign n22985 = \P3_Flush_reg/NET0131  & ~n13810 ;
  assign n22986 = ~n22984 & ~n22985 ;
  assign n22987 = \P2_EAX_reg[16]/NET0131  & ~n12632 ;
  assign n23021 = n12669 & ~n16382 ;
  assign n23022 = \P2_EAX_reg[16]/NET0131  & ~n23021 ;
  assign n23027 = ~\P2_EAX_reg[16]/NET0131  & n12664 ;
  assign n23028 = n12648 & n23027 ;
  assign n22992 = \P2_InstQueue_reg[0][0]/NET0131  & n1482 ;
  assign n22993 = \P2_InstQueue_reg[11][0]/NET0131  & n1472 ;
  assign n23006 = ~n22992 & ~n22993 ;
  assign n22994 = \P2_InstQueue_reg[3][0]/NET0131  & n1464 ;
  assign n22995 = \P2_InstQueue_reg[1][0]/NET0131  & n1478 ;
  assign n23007 = ~n22994 & ~n22995 ;
  assign n23014 = n23006 & n23007 ;
  assign n22988 = \P2_InstQueue_reg[6][0]/NET0131  & n1450 ;
  assign n22989 = \P2_InstQueue_reg[12][0]/NET0131  & n1453 ;
  assign n23004 = ~n22988 & ~n22989 ;
  assign n22990 = \P2_InstQueue_reg[13][0]/NET0131  & n1459 ;
  assign n22991 = \P2_InstQueue_reg[4][0]/NET0131  & n1468 ;
  assign n23005 = ~n22990 & ~n22991 ;
  assign n23015 = n23004 & n23005 ;
  assign n23016 = n23014 & n23015 ;
  assign n23000 = \P2_InstQueue_reg[2][0]/NET0131  & n1456 ;
  assign n23001 = \P2_InstQueue_reg[9][0]/NET0131  & n1476 ;
  assign n23010 = ~n23000 & ~n23001 ;
  assign n23002 = \P2_InstQueue_reg[8][0]/NET0131  & n1447 ;
  assign n23003 = \P2_InstQueue_reg[7][0]/NET0131  & n1474 ;
  assign n23011 = ~n23002 & ~n23003 ;
  assign n23012 = n23010 & n23011 ;
  assign n22996 = \P2_InstQueue_reg[14][0]/NET0131  & n1480 ;
  assign n22997 = \P2_InstQueue_reg[15][0]/NET0131  & n1466 ;
  assign n23008 = ~n22996 & ~n22997 ;
  assign n22998 = \P2_InstQueue_reg[10][0]/NET0131  & n1461 ;
  assign n22999 = \P2_InstQueue_reg[5][0]/NET0131  & n1470 ;
  assign n23009 = ~n22998 & ~n22999 ;
  assign n23013 = n23008 & n23009 ;
  assign n23017 = n23012 & n23013 ;
  assign n23018 = n23016 & n23017 ;
  assign n23019 = n1798 & ~n23018 ;
  assign n23020 = n1726 & n23019 ;
  assign n23023 = n1803 & ~n15419 ;
  assign n23024 = n1742 & ~n15407 ;
  assign n23025 = ~n23023 & ~n23024 ;
  assign n23026 = n1811 & ~n23025 ;
  assign n23029 = ~n23020 & ~n23026 ;
  assign n23030 = ~n23028 & n23029 ;
  assign n23031 = ~n23022 & n23030 ;
  assign n23032 = n1927 & ~n23031 ;
  assign n23033 = ~n22987 & ~n23032 ;
  assign n23034 = \P2_EAX_reg[17]/NET0131  & ~n12632 ;
  assign n23069 = \P2_EAX_reg[17]/NET0131  & n12649 ;
  assign n23068 = ~\P2_EAX_reg[17]/NET0131  & ~n12649 ;
  assign n23070 = n12664 & ~n23068 ;
  assign n23071 = ~n23069 & n23070 ;
  assign n23076 = n1742 & ~n1811 ;
  assign n23077 = n12668 & ~n23076 ;
  assign n23078 = \P2_EAX_reg[17]/NET0131  & ~n23077 ;
  assign n23073 = n1811 & n11553 ;
  assign n23072 = ~\P2_EAX_reg[17]/NET0131  & ~n1811 ;
  assign n23074 = n1803 & ~n23072 ;
  assign n23075 = ~n23073 & n23074 ;
  assign n23039 = \P2_InstQueue_reg[3][1]/NET0131  & n1464 ;
  assign n23040 = \P2_InstQueue_reg[13][1]/NET0131  & n1459 ;
  assign n23053 = ~n23039 & ~n23040 ;
  assign n23041 = \P2_InstQueue_reg[9][1]/NET0131  & n1476 ;
  assign n23042 = \P2_InstQueue_reg[7][1]/NET0131  & n1474 ;
  assign n23054 = ~n23041 & ~n23042 ;
  assign n23061 = n23053 & n23054 ;
  assign n23035 = \P2_InstQueue_reg[6][1]/NET0131  & n1450 ;
  assign n23036 = \P2_InstQueue_reg[12][1]/NET0131  & n1453 ;
  assign n23051 = ~n23035 & ~n23036 ;
  assign n23037 = \P2_InstQueue_reg[11][1]/NET0131  & n1472 ;
  assign n23038 = \P2_InstQueue_reg[5][1]/NET0131  & n1470 ;
  assign n23052 = ~n23037 & ~n23038 ;
  assign n23062 = n23051 & n23052 ;
  assign n23063 = n23061 & n23062 ;
  assign n23047 = \P2_InstQueue_reg[15][1]/NET0131  & n1466 ;
  assign n23048 = \P2_InstQueue_reg[8][1]/NET0131  & n1447 ;
  assign n23057 = ~n23047 & ~n23048 ;
  assign n23049 = \P2_InstQueue_reg[1][1]/NET0131  & n1478 ;
  assign n23050 = \P2_InstQueue_reg[0][1]/NET0131  & n1482 ;
  assign n23058 = ~n23049 & ~n23050 ;
  assign n23059 = n23057 & n23058 ;
  assign n23043 = \P2_InstQueue_reg[4][1]/NET0131  & n1468 ;
  assign n23044 = \P2_InstQueue_reg[2][1]/NET0131  & n1456 ;
  assign n23055 = ~n23043 & ~n23044 ;
  assign n23045 = \P2_InstQueue_reg[10][1]/NET0131  & n1461 ;
  assign n23046 = \P2_InstQueue_reg[14][1]/NET0131  & n1480 ;
  assign n23056 = ~n23045 & ~n23046 ;
  assign n23060 = n23055 & n23056 ;
  assign n23064 = n23059 & n23060 ;
  assign n23065 = n23063 & n23064 ;
  assign n23066 = n1798 & ~n23065 ;
  assign n23067 = n1726 & n23066 ;
  assign n23079 = n1742 & n17778 ;
  assign n23080 = ~n23067 & ~n23079 ;
  assign n23081 = ~n23075 & n23080 ;
  assign n23082 = ~n23078 & n23081 ;
  assign n23083 = ~n23071 & n23082 ;
  assign n23084 = n1927 & ~n23083 ;
  assign n23085 = ~n23034 & ~n23084 ;
  assign n23086 = \P2_EAX_reg[18]/NET0131  & ~n12632 ;
  assign n23120 = ~n12651 & n12664 ;
  assign n23121 = n12668 & ~n23120 ;
  assign n23122 = \P2_EAX_reg[18]/NET0131  & ~n23121 ;
  assign n23123 = n23069 & n23120 ;
  assign n23124 = \P2_EAX_reg[18]/NET0131  & ~n1811 ;
  assign n23127 = n1811 & ~n8601 ;
  assign n23128 = ~n23124 & ~n23127 ;
  assign n23129 = n1803 & ~n23128 ;
  assign n23091 = \P2_InstQueue_reg[3][2]/NET0131  & n1464 ;
  assign n23092 = \P2_InstQueue_reg[9][2]/NET0131  & n1476 ;
  assign n23105 = ~n23091 & ~n23092 ;
  assign n23093 = \P2_InstQueue_reg[12][2]/NET0131  & n1453 ;
  assign n23094 = \P2_InstQueue_reg[7][2]/NET0131  & n1474 ;
  assign n23106 = ~n23093 & ~n23094 ;
  assign n23113 = n23105 & n23106 ;
  assign n23087 = \P2_InstQueue_reg[10][2]/NET0131  & n1461 ;
  assign n23088 = \P2_InstQueue_reg[5][2]/NET0131  & n1470 ;
  assign n23103 = ~n23087 & ~n23088 ;
  assign n23089 = \P2_InstQueue_reg[11][2]/NET0131  & n1472 ;
  assign n23090 = \P2_InstQueue_reg[4][2]/NET0131  & n1468 ;
  assign n23104 = ~n23089 & ~n23090 ;
  assign n23114 = n23103 & n23104 ;
  assign n23115 = n23113 & n23114 ;
  assign n23099 = \P2_InstQueue_reg[15][2]/NET0131  & n1466 ;
  assign n23100 = \P2_InstQueue_reg[8][2]/NET0131  & n1447 ;
  assign n23109 = ~n23099 & ~n23100 ;
  assign n23101 = \P2_InstQueue_reg[13][2]/NET0131  & n1459 ;
  assign n23102 = \P2_InstQueue_reg[0][2]/NET0131  & n1482 ;
  assign n23110 = ~n23101 & ~n23102 ;
  assign n23111 = n23109 & n23110 ;
  assign n23095 = \P2_InstQueue_reg[1][2]/NET0131  & n1478 ;
  assign n23096 = \P2_InstQueue_reg[2][2]/NET0131  & n1456 ;
  assign n23107 = ~n23095 & ~n23096 ;
  assign n23097 = \P2_InstQueue_reg[6][2]/NET0131  & n1450 ;
  assign n23098 = \P2_InstQueue_reg[14][2]/NET0131  & n1480 ;
  assign n23108 = ~n23097 & ~n23098 ;
  assign n23112 = n23107 & n23108 ;
  assign n23116 = n23111 & n23112 ;
  assign n23117 = n23115 & n23116 ;
  assign n23118 = n1798 & ~n23117 ;
  assign n23119 = n1726 & n23118 ;
  assign n23125 = ~n22459 & ~n23124 ;
  assign n23126 = n1742 & ~n23125 ;
  assign n23130 = ~n23119 & ~n23126 ;
  assign n23131 = ~n23129 & n23130 ;
  assign n23132 = ~n23123 & n23131 ;
  assign n23133 = ~n23122 & n23132 ;
  assign n23134 = n1927 & ~n23133 ;
  assign n23135 = ~n23086 & ~n23134 ;
  assign n23136 = \P2_EAX_reg[19]/NET0131  & ~n12632 ;
  assign n23170 = \P2_EAX_reg[19]/NET0131  & ~n23121 ;
  assign n23177 = ~\P2_EAX_reg[19]/NET0131  & n12664 ;
  assign n23178 = n12651 & n23177 ;
  assign n23171 = \P2_EAX_reg[19]/NET0131  & ~n1811 ;
  assign n23175 = ~n22470 & ~n23171 ;
  assign n23176 = n1742 & ~n23175 ;
  assign n23141 = \P2_InstQueue_reg[3][3]/NET0131  & n1464 ;
  assign n23142 = \P2_InstQueue_reg[9][3]/NET0131  & n1476 ;
  assign n23155 = ~n23141 & ~n23142 ;
  assign n23143 = \P2_InstQueue_reg[12][3]/NET0131  & n1453 ;
  assign n23144 = \P2_InstQueue_reg[7][3]/NET0131  & n1474 ;
  assign n23156 = ~n23143 & ~n23144 ;
  assign n23163 = n23155 & n23156 ;
  assign n23137 = \P2_InstQueue_reg[10][3]/NET0131  & n1461 ;
  assign n23138 = \P2_InstQueue_reg[5][3]/NET0131  & n1470 ;
  assign n23153 = ~n23137 & ~n23138 ;
  assign n23139 = \P2_InstQueue_reg[11][3]/NET0131  & n1472 ;
  assign n23140 = \P2_InstQueue_reg[4][3]/NET0131  & n1468 ;
  assign n23154 = ~n23139 & ~n23140 ;
  assign n23164 = n23153 & n23154 ;
  assign n23165 = n23163 & n23164 ;
  assign n23149 = \P2_InstQueue_reg[15][3]/NET0131  & n1466 ;
  assign n23150 = \P2_InstQueue_reg[8][3]/NET0131  & n1447 ;
  assign n23159 = ~n23149 & ~n23150 ;
  assign n23151 = \P2_InstQueue_reg[13][3]/NET0131  & n1459 ;
  assign n23152 = \P2_InstQueue_reg[0][3]/NET0131  & n1482 ;
  assign n23160 = ~n23151 & ~n23152 ;
  assign n23161 = n23159 & n23160 ;
  assign n23145 = \P2_InstQueue_reg[1][3]/NET0131  & n1478 ;
  assign n23146 = \P2_InstQueue_reg[2][3]/NET0131  & n1456 ;
  assign n23157 = ~n23145 & ~n23146 ;
  assign n23147 = \P2_InstQueue_reg[6][3]/NET0131  & n1450 ;
  assign n23148 = \P2_InstQueue_reg[14][3]/NET0131  & n1480 ;
  assign n23158 = ~n23147 & ~n23148 ;
  assign n23162 = n23157 & n23158 ;
  assign n23166 = n23161 & n23162 ;
  assign n23167 = n23165 & n23166 ;
  assign n23168 = n1798 & ~n23167 ;
  assign n23169 = n1726 & n23168 ;
  assign n23172 = n1811 & ~n5310 ;
  assign n23173 = ~n23171 & ~n23172 ;
  assign n23174 = n1803 & ~n23173 ;
  assign n23179 = ~n23169 & ~n23174 ;
  assign n23180 = ~n23176 & n23179 ;
  assign n23181 = ~n23178 & n23180 ;
  assign n23182 = ~n23170 & n23181 ;
  assign n23183 = n1927 & ~n23182 ;
  assign n23184 = ~n23136 & ~n23183 ;
  assign n23185 = n1927 & ~n12668 ;
  assign n23186 = n12632 & ~n23185 ;
  assign n23187 = \P2_EAX_reg[20]/NET0131  & ~n23186 ;
  assign n23221 = ~n12653 & n12664 ;
  assign n23222 = ~n1812 & ~n23221 ;
  assign n23223 = \P2_EAX_reg[20]/NET0131  & ~n23222 ;
  assign n23224 = n12652 & n23221 ;
  assign n23192 = \P2_InstQueue_reg[7][4]/NET0131  & n1474 ;
  assign n23193 = \P2_InstQueue_reg[1][4]/NET0131  & n1478 ;
  assign n23206 = ~n23192 & ~n23193 ;
  assign n23194 = \P2_InstQueue_reg[11][4]/NET0131  & n1472 ;
  assign n23195 = \P2_InstQueue_reg[14][4]/NET0131  & n1480 ;
  assign n23207 = ~n23194 & ~n23195 ;
  assign n23214 = n23206 & n23207 ;
  assign n23188 = \P2_InstQueue_reg[10][4]/NET0131  & n1461 ;
  assign n23189 = \P2_InstQueue_reg[4][4]/NET0131  & n1468 ;
  assign n23204 = ~n23188 & ~n23189 ;
  assign n23190 = \P2_InstQueue_reg[9][4]/NET0131  & n1476 ;
  assign n23191 = \P2_InstQueue_reg[13][4]/NET0131  & n1459 ;
  assign n23205 = ~n23190 & ~n23191 ;
  assign n23215 = n23204 & n23205 ;
  assign n23216 = n23214 & n23215 ;
  assign n23200 = \P2_InstQueue_reg[8][4]/NET0131  & n1447 ;
  assign n23201 = \P2_InstQueue_reg[2][4]/NET0131  & n1456 ;
  assign n23210 = ~n23200 & ~n23201 ;
  assign n23202 = \P2_InstQueue_reg[5][4]/NET0131  & n1470 ;
  assign n23203 = \P2_InstQueue_reg[3][4]/NET0131  & n1464 ;
  assign n23211 = ~n23202 & ~n23203 ;
  assign n23212 = n23210 & n23211 ;
  assign n23196 = \P2_InstQueue_reg[12][4]/NET0131  & n1453 ;
  assign n23197 = \P2_InstQueue_reg[15][4]/NET0131  & n1466 ;
  assign n23208 = ~n23196 & ~n23197 ;
  assign n23198 = \P2_InstQueue_reg[6][4]/NET0131  & n1450 ;
  assign n23199 = \P2_InstQueue_reg[0][4]/NET0131  & n1482 ;
  assign n23209 = ~n23198 & ~n23199 ;
  assign n23213 = n23208 & n23209 ;
  assign n23217 = n23212 & n23213 ;
  assign n23218 = n23216 & n23217 ;
  assign n23219 = n1798 & ~n23218 ;
  assign n23220 = n1726 & n23219 ;
  assign n23225 = n1803 & ~n3101 ;
  assign n23226 = n1742 & ~n3082 ;
  assign n23227 = ~n23225 & ~n23226 ;
  assign n23228 = n1811 & ~n23227 ;
  assign n23229 = ~n23220 & ~n23228 ;
  assign n23230 = ~n23224 & n23229 ;
  assign n23231 = ~n23223 & n23230 ;
  assign n23232 = n1927 & ~n23231 ;
  assign n23233 = ~n23187 & ~n23232 ;
  assign n23234 = \P2_EAX_reg[21]/NET0131  & ~n12632 ;
  assign n23236 = ~\P2_EAX_reg[21]/NET0131  & ~n12653 ;
  assign n23237 = \P2_EAX_reg[21]/NET0131  & n12653 ;
  assign n23238 = n12664 & ~n23237 ;
  assign n23239 = ~n23236 & n23238 ;
  assign n23235 = \P2_EAX_reg[21]/NET0131  & ~n12669 ;
  assign n23240 = n1742 & ~n10333 ;
  assign n23241 = n1803 & ~n10345 ;
  assign n23242 = ~n23240 & ~n23241 ;
  assign n23243 = n1811 & ~n23242 ;
  assign n23248 = \P2_InstQueue_reg[5][5]/NET0131  & n1470 ;
  assign n23249 = \P2_InstQueue_reg[9][5]/NET0131  & n1476 ;
  assign n23262 = ~n23248 & ~n23249 ;
  assign n23250 = \P2_InstQueue_reg[12][5]/NET0131  & n1453 ;
  assign n23251 = \P2_InstQueue_reg[7][5]/NET0131  & n1474 ;
  assign n23263 = ~n23250 & ~n23251 ;
  assign n23270 = n23262 & n23263 ;
  assign n23244 = \P2_InstQueue_reg[10][5]/NET0131  & n1461 ;
  assign n23245 = \P2_InstQueue_reg[8][5]/NET0131  & n1447 ;
  assign n23260 = ~n23244 & ~n23245 ;
  assign n23246 = \P2_InstQueue_reg[14][5]/NET0131  & n1480 ;
  assign n23247 = \P2_InstQueue_reg[4][5]/NET0131  & n1468 ;
  assign n23261 = ~n23246 & ~n23247 ;
  assign n23271 = n23260 & n23261 ;
  assign n23272 = n23270 & n23271 ;
  assign n23256 = \P2_InstQueue_reg[15][5]/NET0131  & n1466 ;
  assign n23257 = \P2_InstQueue_reg[3][5]/NET0131  & n1464 ;
  assign n23266 = ~n23256 & ~n23257 ;
  assign n23258 = \P2_InstQueue_reg[13][5]/NET0131  & n1459 ;
  assign n23259 = \P2_InstQueue_reg[0][5]/NET0131  & n1482 ;
  assign n23267 = ~n23258 & ~n23259 ;
  assign n23268 = n23266 & n23267 ;
  assign n23252 = \P2_InstQueue_reg[11][5]/NET0131  & n1472 ;
  assign n23253 = \P2_InstQueue_reg[2][5]/NET0131  & n1456 ;
  assign n23264 = ~n23252 & ~n23253 ;
  assign n23254 = \P2_InstQueue_reg[6][5]/NET0131  & n1450 ;
  assign n23255 = \P2_InstQueue_reg[1][5]/NET0131  & n1478 ;
  assign n23265 = ~n23254 & ~n23255 ;
  assign n23269 = n23264 & n23265 ;
  assign n23273 = n23268 & n23269 ;
  assign n23274 = n23272 & n23273 ;
  assign n23275 = n1798 & ~n23274 ;
  assign n23276 = n1726 & n23275 ;
  assign n23277 = ~n23243 & ~n23276 ;
  assign n23278 = ~n23235 & n23277 ;
  assign n23279 = ~n23239 & n23278 ;
  assign n23280 = n1927 & ~n23279 ;
  assign n23281 = ~n23234 & ~n23280 ;
  assign n23282 = \P2_EAX_reg[22]/NET0131  & ~n12632 ;
  assign n23316 = n12669 & ~n23238 ;
  assign n23317 = \P2_EAX_reg[22]/NET0131  & ~n23316 ;
  assign n23322 = ~\P2_EAX_reg[22]/NET0131  & n12664 ;
  assign n23323 = n23237 & n23322 ;
  assign n23287 = \P2_InstQueue_reg[5][6]/NET0131  & n1470 ;
  assign n23288 = \P2_InstQueue_reg[2][6]/NET0131  & n1456 ;
  assign n23301 = ~n23287 & ~n23288 ;
  assign n23289 = \P2_InstQueue_reg[13][6]/NET0131  & n1459 ;
  assign n23290 = \P2_InstQueue_reg[0][6]/NET0131  & n1482 ;
  assign n23302 = ~n23289 & ~n23290 ;
  assign n23309 = n23301 & n23302 ;
  assign n23283 = \P2_InstQueue_reg[6][6]/NET0131  & n1450 ;
  assign n23284 = \P2_InstQueue_reg[12][6]/NET0131  & n1453 ;
  assign n23299 = ~n23283 & ~n23284 ;
  assign n23285 = \P2_InstQueue_reg[1][6]/NET0131  & n1478 ;
  assign n23286 = \P2_InstQueue_reg[3][6]/NET0131  & n1464 ;
  assign n23300 = ~n23285 & ~n23286 ;
  assign n23310 = n23299 & n23300 ;
  assign n23311 = n23309 & n23310 ;
  assign n23295 = \P2_InstQueue_reg[15][6]/NET0131  & n1466 ;
  assign n23296 = \P2_InstQueue_reg[11][6]/NET0131  & n1472 ;
  assign n23305 = ~n23295 & ~n23296 ;
  assign n23297 = \P2_InstQueue_reg[9][6]/NET0131  & n1476 ;
  assign n23298 = \P2_InstQueue_reg[14][6]/NET0131  & n1480 ;
  assign n23306 = ~n23297 & ~n23298 ;
  assign n23307 = n23305 & n23306 ;
  assign n23291 = \P2_InstQueue_reg[4][6]/NET0131  & n1468 ;
  assign n23292 = \P2_InstQueue_reg[8][6]/NET0131  & n1447 ;
  assign n23303 = ~n23291 & ~n23292 ;
  assign n23293 = \P2_InstQueue_reg[10][6]/NET0131  & n1461 ;
  assign n23294 = \P2_InstQueue_reg[7][6]/NET0131  & n1474 ;
  assign n23304 = ~n23293 & ~n23294 ;
  assign n23308 = n23303 & n23304 ;
  assign n23312 = n23307 & n23308 ;
  assign n23313 = n23311 & n23312 ;
  assign n23314 = n1798 & ~n23313 ;
  assign n23315 = n1726 & n23314 ;
  assign n23318 = n1742 & ~n7724 ;
  assign n23319 = n1803 & ~n7736 ;
  assign n23320 = ~n23318 & ~n23319 ;
  assign n23321 = n1811 & ~n23320 ;
  assign n23324 = ~n23315 & ~n23321 ;
  assign n23325 = ~n23323 & n23324 ;
  assign n23326 = ~n23317 & n23325 ;
  assign n23327 = n1927 & ~n23326 ;
  assign n23328 = ~n23282 & ~n23327 ;
  assign n23329 = \P2_EAX_reg[23]/NET0131  & ~n12632 ;
  assign n23331 = ~\P2_EAX_reg[23]/NET0131  & ~n12655 ;
  assign n23332 = n12664 & ~n21792 ;
  assign n23333 = ~n23331 & n23332 ;
  assign n23330 = \P2_EAX_reg[23]/NET0131  & ~n12669 ;
  assign n23334 = n1803 & ~n3140 ;
  assign n23335 = n1742 & ~n3128 ;
  assign n23336 = ~n23334 & ~n23335 ;
  assign n23337 = n1811 & ~n23336 ;
  assign n23338 = n12704 & n12735 ;
  assign n23339 = ~n12736 & ~n23338 ;
  assign n23340 = n1798 & n23339 ;
  assign n23341 = n1726 & n23340 ;
  assign n23342 = ~n23337 & ~n23341 ;
  assign n23343 = ~n23330 & n23342 ;
  assign n23344 = ~n23333 & n23343 ;
  assign n23345 = n1927 & ~n23344 ;
  assign n23346 = ~n23329 & ~n23345 ;
  assign n23347 = \P2_EAX_reg[24]/NET0131  & ~n23186 ;
  assign n23352 = ~\P2_EAX_reg[24]/NET0131  & ~n21792 ;
  assign n23353 = n21794 & ~n23352 ;
  assign n23355 = ~n1805 & ~n15415 ;
  assign n23356 = n1803 & n23355 ;
  assign n23357 = ~n16957 & ~n23356 ;
  assign n23358 = ~n1810 & ~n23357 ;
  assign n23348 = ~n12736 & n12767 ;
  assign n23349 = ~n12768 & ~n23348 ;
  assign n23350 = n1798 & n23349 ;
  assign n23351 = n1726 & n23350 ;
  assign n23354 = \P2_EAX_reg[24]/NET0131  & n1812 ;
  assign n23359 = ~n23351 & ~n23354 ;
  assign n23360 = ~n23358 & n23359 ;
  assign n23361 = ~n23353 & n23360 ;
  assign n23362 = n1927 & ~n23361 ;
  assign n23363 = ~n23347 & ~n23362 ;
  assign n23364 = \P2_EAX_reg[28]/NET0131  & ~n23186 ;
  assign n23366 = n12658 & n12659 ;
  assign n23367 = ~\P2_EAX_reg[28]/NET0131  & ~n23366 ;
  assign n23368 = ~n12661 & n12664 ;
  assign n23369 = ~n23367 & n23368 ;
  assign n23370 = ~n12864 & n12895 ;
  assign n23371 = n1798 & ~n12896 ;
  assign n23372 = ~n23370 & n23371 ;
  assign n23373 = n1726 & n23372 ;
  assign n23365 = \P2_EAX_reg[28]/NET0131  & n1812 ;
  assign n23374 = ~n1805 & ~n3094 ;
  assign n23375 = n1803 & n23374 ;
  assign n23376 = ~n15948 & ~n23375 ;
  assign n23377 = ~n1810 & ~n23376 ;
  assign n23378 = ~n23365 & ~n23377 ;
  assign n23379 = ~n23373 & n23378 ;
  assign n23380 = ~n23369 & n23379 ;
  assign n23381 = n1927 & ~n23380 ;
  assign n23382 = ~n23364 & ~n23381 ;
  assign n23383 = \P1_EAX_reg[0]/NET0131  & ~n16968 ;
  assign n23386 = n2377 & ~n5179 ;
  assign n23387 = ~n2303 & n23386 ;
  assign n23384 = n2337 & ~n4743 ;
  assign n23385 = n2331 & n23384 ;
  assign n23388 = ~n18186 & ~n23385 ;
  assign n23389 = ~n23387 & n23388 ;
  assign n23390 = n2432 & ~n23389 ;
  assign n23391 = ~n23383 & ~n23390 ;
  assign n23394 = ~\P1_EBX_reg[25]/NET0131  & ~n15387 ;
  assign n23395 = n2262 & ~n15388 ;
  assign n23396 = ~n23394 & n23395 ;
  assign n23392 = n2242 & n21745 ;
  assign n23393 = \P1_EBX_reg[25]/NET0131  & ~n15073 ;
  assign n23397 = ~n23392 & ~n23393 ;
  assign n23398 = ~n23396 & n23397 ;
  assign n23399 = n2432 & ~n23398 ;
  assign n23400 = \P1_EBX_reg[25]/NET0131  & ~n15402 ;
  assign n23401 = ~n23399 & ~n23400 ;
  assign n23402 = \P2_EBX_reg[25]/NET0131  & ~n12632 ;
  assign n23404 = \P2_EBX_reg[24]/NET0131  & n15044 ;
  assign n23405 = n1766 & ~n23404 ;
  assign n23406 = n15019 & ~n23405 ;
  assign n23407 = \P2_EBX_reg[25]/NET0131  & ~n23406 ;
  assign n23403 = n1722 & n21790 ;
  assign n23408 = ~\P2_EBX_reg[25]/NET0131  & n1766 ;
  assign n23409 = n23404 & n23408 ;
  assign n23410 = ~n23403 & ~n23409 ;
  assign n23411 = ~n23407 & n23410 ;
  assign n23412 = n1927 & ~n23411 ;
  assign n23413 = ~n23402 & ~n23412 ;
  assign n23414 = ~n1900 & n1927 ;
  assign n23415 = \P2_Flush_reg/NET0131  & ~n12632 ;
  assign n23416 = ~n23414 & ~n23415 ;
  assign n23417 = ~n2393 & n2432 ;
  assign n23418 = \P1_Flush_reg/NET0131  & ~n15402 ;
  assign n23419 = ~n23417 & ~n23418 ;
  assign n23420 = n2453 & ~n2903 ;
  assign n23421 = \P3_More_reg/NET0131  & ~n13810 ;
  assign n23422 = ~n23420 & ~n23421 ;
  assign n23423 = \P3_uWord_reg[11]/NET0131  & ~n16090 ;
  assign n23424 = ~n14049 & ~n22306 ;
  assign n23425 = n2453 & ~n23424 ;
  assign n23426 = ~n23423 & ~n23425 ;
  assign n23428 = ~\P1_EAX_reg[16]/NET0131  & ~n15909 ;
  assign n23429 = n2260 & ~n15910 ;
  assign n23430 = ~n23428 & n23429 ;
  assign n23427 = \P1_EAX_reg[16]/NET0131  & ~n15925 ;
  assign n23431 = n2222 & ~n5179 ;
  assign n23432 = n2302 & ~n5218 ;
  assign n23433 = ~n23431 & ~n23432 ;
  assign n23434 = n2377 & ~n23433 ;
  assign n23439 = \P1_InstQueue_reg[3][0]/NET0131  & n1958 ;
  assign n23440 = \P1_InstQueue_reg[15][0]/NET0131  & n1953 ;
  assign n23453 = ~n23439 & ~n23440 ;
  assign n23441 = \P1_InstQueue_reg[7][0]/NET0131  & n1961 ;
  assign n23442 = \P1_InstQueue_reg[5][0]/NET0131  & n1970 ;
  assign n23454 = ~n23441 & ~n23442 ;
  assign n23461 = n23453 & n23454 ;
  assign n23435 = \P1_InstQueue_reg[2][0]/NET0131  & n1982 ;
  assign n23436 = \P1_InstQueue_reg[11][0]/NET0131  & n1974 ;
  assign n23451 = ~n23435 & ~n23436 ;
  assign n23437 = \P1_InstQueue_reg[6][0]/NET0131  & n1976 ;
  assign n23438 = \P1_InstQueue_reg[4][0]/NET0131  & n1966 ;
  assign n23452 = ~n23437 & ~n23438 ;
  assign n23462 = n23451 & n23452 ;
  assign n23463 = n23461 & n23462 ;
  assign n23447 = \P1_InstQueue_reg[14][0]/NET0131  & n1949 ;
  assign n23448 = \P1_InstQueue_reg[12][0]/NET0131  & n1978 ;
  assign n23457 = ~n23447 & ~n23448 ;
  assign n23449 = \P1_InstQueue_reg[10][0]/NET0131  & n1968 ;
  assign n23450 = \P1_InstQueue_reg[8][0]/NET0131  & n1964 ;
  assign n23458 = ~n23449 & ~n23450 ;
  assign n23459 = n23457 & n23458 ;
  assign n23443 = \P1_InstQueue_reg[9][0]/NET0131  & n1972 ;
  assign n23444 = \P1_InstQueue_reg[13][0]/NET0131  & n1946 ;
  assign n23455 = ~n23443 & ~n23444 ;
  assign n23445 = \P1_InstQueue_reg[1][0]/NET0131  & n1955 ;
  assign n23446 = \P1_InstQueue_reg[0][0]/NET0131  & n1980 ;
  assign n23456 = ~n23445 & ~n23446 ;
  assign n23460 = n23455 & n23456 ;
  assign n23464 = n23459 & n23460 ;
  assign n23465 = n23463 & n23464 ;
  assign n23466 = n2337 & ~n23465 ;
  assign n23467 = n2331 & n23466 ;
  assign n23468 = ~n23434 & ~n23467 ;
  assign n23469 = ~n23427 & n23468 ;
  assign n23470 = ~n23430 & n23469 ;
  assign n23471 = n2432 & ~n23470 ;
  assign n23472 = \P1_EAX_reg[16]/NET0131  & ~n15402 ;
  assign n23473 = ~n23471 & ~n23472 ;
  assign n23474 = \P1_EAX_reg[17]/NET0131  & ~n15402 ;
  assign n23475 = n15925 & ~n23429 ;
  assign n23476 = \P1_EAX_reg[17]/NET0131  & ~n23475 ;
  assign n23477 = ~\P1_EAX_reg[17]/NET0131  & n2260 ;
  assign n23478 = n15910 & n23477 ;
  assign n23483 = \P1_InstQueue_reg[3][1]/NET0131  & n1958 ;
  assign n23484 = \P1_InstQueue_reg[10][1]/NET0131  & n1968 ;
  assign n23497 = ~n23483 & ~n23484 ;
  assign n23485 = \P1_InstQueue_reg[15][1]/NET0131  & n1953 ;
  assign n23486 = \P1_InstQueue_reg[8][1]/NET0131  & n1964 ;
  assign n23498 = ~n23485 & ~n23486 ;
  assign n23505 = n23497 & n23498 ;
  assign n23479 = \P1_InstQueue_reg[2][1]/NET0131  & n1982 ;
  assign n23480 = \P1_InstQueue_reg[11][1]/NET0131  & n1974 ;
  assign n23495 = ~n23479 & ~n23480 ;
  assign n23481 = \P1_InstQueue_reg[6][1]/NET0131  & n1976 ;
  assign n23482 = \P1_InstQueue_reg[4][1]/NET0131  & n1966 ;
  assign n23496 = ~n23481 & ~n23482 ;
  assign n23506 = n23495 & n23496 ;
  assign n23507 = n23505 & n23506 ;
  assign n23491 = \P1_InstQueue_reg[14][1]/NET0131  & n1949 ;
  assign n23492 = \P1_InstQueue_reg[12][1]/NET0131  & n1978 ;
  assign n23501 = ~n23491 & ~n23492 ;
  assign n23493 = \P1_InstQueue_reg[9][1]/NET0131  & n1972 ;
  assign n23494 = \P1_InstQueue_reg[5][1]/NET0131  & n1970 ;
  assign n23502 = ~n23493 & ~n23494 ;
  assign n23503 = n23501 & n23502 ;
  assign n23487 = \P1_InstQueue_reg[7][1]/NET0131  & n1961 ;
  assign n23488 = \P1_InstQueue_reg[13][1]/NET0131  & n1946 ;
  assign n23499 = ~n23487 & ~n23488 ;
  assign n23489 = \P1_InstQueue_reg[1][1]/NET0131  & n1955 ;
  assign n23490 = \P1_InstQueue_reg[0][1]/NET0131  & n1980 ;
  assign n23500 = ~n23489 & ~n23490 ;
  assign n23504 = n23499 & n23500 ;
  assign n23508 = n23503 & n23504 ;
  assign n23509 = n23507 & n23508 ;
  assign n23510 = n2337 & ~n23509 ;
  assign n23511 = n2331 & n23510 ;
  assign n23512 = n2302 & ~n5236 ;
  assign n23513 = n2222 & ~n5185 ;
  assign n23514 = ~n23512 & ~n23513 ;
  assign n23515 = n2377 & ~n23514 ;
  assign n23516 = ~n23511 & ~n23515 ;
  assign n23517 = ~n23478 & n23516 ;
  assign n23518 = ~n23476 & n23517 ;
  assign n23519 = n2432 & ~n23518 ;
  assign n23520 = ~n23474 & ~n23519 ;
  assign n23521 = ~n2383 & n2432 ;
  assign n23522 = \P1_More_reg/NET0131  & ~n15402 ;
  assign n23523 = ~n23521 & ~n23522 ;
  assign n23524 = \P1_EAX_reg[19]/NET0131  & ~n15402 ;
  assign n23527 = n2260 & ~n15912 ;
  assign n23528 = n15925 & ~n23527 ;
  assign n23529 = \P1_EAX_reg[19]/NET0131  & ~n23528 ;
  assign n23525 = ~\P1_EAX_reg[19]/NET0131  & n2260 ;
  assign n23526 = n15912 & n23525 ;
  assign n23534 = \P1_InstQueue_reg[3][3]/NET0131  & n1958 ;
  assign n23535 = \P1_InstQueue_reg[10][3]/NET0131  & n1968 ;
  assign n23548 = ~n23534 & ~n23535 ;
  assign n23536 = \P1_InstQueue_reg[6][3]/NET0131  & n1976 ;
  assign n23537 = \P1_InstQueue_reg[5][3]/NET0131  & n1970 ;
  assign n23549 = ~n23536 & ~n23537 ;
  assign n23556 = n23548 & n23549 ;
  assign n23530 = \P1_InstQueue_reg[2][3]/NET0131  & n1982 ;
  assign n23531 = \P1_InstQueue_reg[4][3]/NET0131  & n1966 ;
  assign n23546 = ~n23530 & ~n23531 ;
  assign n23532 = \P1_InstQueue_reg[15][3]/NET0131  & n1953 ;
  assign n23533 = \P1_InstQueue_reg[11][3]/NET0131  & n1974 ;
  assign n23547 = ~n23532 & ~n23533 ;
  assign n23557 = n23546 & n23547 ;
  assign n23558 = n23556 & n23557 ;
  assign n23542 = \P1_InstQueue_reg[12][3]/NET0131  & n1978 ;
  assign n23543 = \P1_InstQueue_reg[13][3]/NET0131  & n1946 ;
  assign n23552 = ~n23542 & ~n23543 ;
  assign n23544 = \P1_InstQueue_reg[9][3]/NET0131  & n1972 ;
  assign n23545 = \P1_InstQueue_reg[8][3]/NET0131  & n1964 ;
  assign n23553 = ~n23544 & ~n23545 ;
  assign n23554 = n23552 & n23553 ;
  assign n23538 = \P1_InstQueue_reg[7][3]/NET0131  & n1961 ;
  assign n23539 = \P1_InstQueue_reg[14][3]/NET0131  & n1949 ;
  assign n23550 = ~n23538 & ~n23539 ;
  assign n23540 = \P1_InstQueue_reg[1][3]/NET0131  & n1955 ;
  assign n23541 = \P1_InstQueue_reg[0][3]/NET0131  & n1980 ;
  assign n23551 = ~n23540 & ~n23541 ;
  assign n23555 = n23550 & n23551 ;
  assign n23559 = n23554 & n23555 ;
  assign n23560 = n23558 & n23559 ;
  assign n23561 = n2337 & ~n23560 ;
  assign n23562 = n2331 & n23561 ;
  assign n23563 = n2302 & ~n5230 ;
  assign n23564 = n2222 & ~n5167 ;
  assign n23565 = ~n23563 & ~n23564 ;
  assign n23566 = n2377 & ~n23565 ;
  assign n23567 = ~n23562 & ~n23566 ;
  assign n23568 = ~n23526 & n23567 ;
  assign n23569 = ~n23529 & n23568 ;
  assign n23570 = n2432 & ~n23569 ;
  assign n23571 = ~n23524 & ~n23570 ;
  assign n23572 = \P1_EAX_reg[18]/NET0131  & ~n15402 ;
  assign n23606 = \P1_EAX_reg[18]/NET0131  & ~n23528 ;
  assign n23611 = \P1_EAX_reg[17]/NET0131  & n15910 ;
  assign n23612 = n23527 & n23611 ;
  assign n23577 = \P1_InstQueue_reg[1][2]/NET0131  & n1955 ;
  assign n23578 = \P1_InstQueue_reg[14][2]/NET0131  & n1949 ;
  assign n23591 = ~n23577 & ~n23578 ;
  assign n23579 = \P1_InstQueue_reg[4][2]/NET0131  & n1966 ;
  assign n23580 = \P1_InstQueue_reg[8][2]/NET0131  & n1964 ;
  assign n23592 = ~n23579 & ~n23580 ;
  assign n23599 = n23591 & n23592 ;
  assign n23573 = \P1_InstQueue_reg[6][2]/NET0131  & n1976 ;
  assign n23574 = \P1_InstQueue_reg[11][2]/NET0131  & n1974 ;
  assign n23589 = ~n23573 & ~n23574 ;
  assign n23575 = \P1_InstQueue_reg[0][2]/NET0131  & n1980 ;
  assign n23576 = \P1_InstQueue_reg[3][2]/NET0131  & n1958 ;
  assign n23590 = ~n23575 & ~n23576 ;
  assign n23600 = n23589 & n23590 ;
  assign n23601 = n23599 & n23600 ;
  assign n23585 = \P1_InstQueue_reg[13][2]/NET0131  & n1946 ;
  assign n23586 = \P1_InstQueue_reg[9][2]/NET0131  & n1972 ;
  assign n23595 = ~n23585 & ~n23586 ;
  assign n23587 = \P1_InstQueue_reg[7][2]/NET0131  & n1961 ;
  assign n23588 = \P1_InstQueue_reg[5][2]/NET0131  & n1970 ;
  assign n23596 = ~n23587 & ~n23588 ;
  assign n23597 = n23595 & n23596 ;
  assign n23581 = \P1_InstQueue_reg[15][2]/NET0131  & n1953 ;
  assign n23582 = \P1_InstQueue_reg[12][2]/NET0131  & n1978 ;
  assign n23593 = ~n23581 & ~n23582 ;
  assign n23583 = \P1_InstQueue_reg[2][2]/NET0131  & n1982 ;
  assign n23584 = \P1_InstQueue_reg[10][2]/NET0131  & n1968 ;
  assign n23594 = ~n23583 & ~n23584 ;
  assign n23598 = n23593 & n23594 ;
  assign n23602 = n23597 & n23598 ;
  assign n23603 = n23601 & n23602 ;
  assign n23604 = n2337 & ~n23603 ;
  assign n23605 = n2331 & n23604 ;
  assign n23607 = n2302 & ~n5233 ;
  assign n23608 = n2222 & ~n5188 ;
  assign n23609 = ~n23607 & ~n23608 ;
  assign n23610 = n2377 & ~n23609 ;
  assign n23613 = ~n23605 & ~n23610 ;
  assign n23614 = ~n23612 & n23613 ;
  assign n23615 = ~n23606 & n23614 ;
  assign n23616 = n2432 & ~n23615 ;
  assign n23617 = ~n23572 & ~n23616 ;
  assign n23618 = \P1_EAX_reg[20]/NET0131  & ~n15402 ;
  assign n23621 = \P1_EAX_reg[20]/NET0131  & n15913 ;
  assign n23620 = ~\P1_EAX_reg[20]/NET0131  & ~n15913 ;
  assign n23622 = n2260 & ~n23620 ;
  assign n23623 = ~n23621 & n23622 ;
  assign n23619 = \P1_EAX_reg[20]/NET0131  & ~n15925 ;
  assign n23624 = n2222 & ~n5140 ;
  assign n23625 = n2302 & ~n5239 ;
  assign n23626 = ~n23624 & ~n23625 ;
  assign n23627 = n2377 & ~n23626 ;
  assign n23632 = \P1_InstQueue_reg[6][4]/NET0131  & n1976 ;
  assign n23633 = \P1_InstQueue_reg[12][4]/NET0131  & n1978 ;
  assign n23646 = ~n23632 & ~n23633 ;
  assign n23634 = \P1_InstQueue_reg[4][4]/NET0131  & n1966 ;
  assign n23635 = \P1_InstQueue_reg[10][4]/NET0131  & n1968 ;
  assign n23647 = ~n23634 & ~n23635 ;
  assign n23654 = n23646 & n23647 ;
  assign n23628 = \P1_InstQueue_reg[1][4]/NET0131  & n1955 ;
  assign n23629 = \P1_InstQueue_reg[11][4]/NET0131  & n1974 ;
  assign n23644 = ~n23628 & ~n23629 ;
  assign n23630 = \P1_InstQueue_reg[0][4]/NET0131  & n1980 ;
  assign n23631 = \P1_InstQueue_reg[7][4]/NET0131  & n1961 ;
  assign n23645 = ~n23630 & ~n23631 ;
  assign n23655 = n23644 & n23645 ;
  assign n23656 = n23654 & n23655 ;
  assign n23640 = \P1_InstQueue_reg[14][4]/NET0131  & n1949 ;
  assign n23641 = \P1_InstQueue_reg[8][4]/NET0131  & n1964 ;
  assign n23650 = ~n23640 & ~n23641 ;
  assign n23642 = \P1_InstQueue_reg[5][4]/NET0131  & n1970 ;
  assign n23643 = \P1_InstQueue_reg[15][4]/NET0131  & n1953 ;
  assign n23651 = ~n23642 & ~n23643 ;
  assign n23652 = n23650 & n23651 ;
  assign n23636 = \P1_InstQueue_reg[3][4]/NET0131  & n1958 ;
  assign n23637 = \P1_InstQueue_reg[13][4]/NET0131  & n1946 ;
  assign n23648 = ~n23636 & ~n23637 ;
  assign n23638 = \P1_InstQueue_reg[2][4]/NET0131  & n1982 ;
  assign n23639 = \P1_InstQueue_reg[9][4]/NET0131  & n1972 ;
  assign n23649 = ~n23638 & ~n23639 ;
  assign n23653 = n23648 & n23649 ;
  assign n23657 = n23652 & n23653 ;
  assign n23658 = n23656 & n23657 ;
  assign n23659 = n2337 & ~n23658 ;
  assign n23660 = n2331 & n23659 ;
  assign n23661 = ~n23627 & ~n23660 ;
  assign n23662 = ~n23619 & n23661 ;
  assign n23663 = ~n23623 & n23662 ;
  assign n23664 = n2432 & ~n23663 ;
  assign n23665 = ~n23618 & ~n23664 ;
  assign n23666 = \P1_EAX_reg[21]/NET0131  & ~n15402 ;
  assign n23668 = ~\P1_EAX_reg[21]/NET0131  & ~n23621 ;
  assign n23669 = n15913 & n15914 ;
  assign n23670 = n2260 & ~n23669 ;
  assign n23671 = ~n23668 & n23670 ;
  assign n23667 = \P1_EAX_reg[21]/NET0131  & ~n15925 ;
  assign n23672 = n2302 & ~n5227 ;
  assign n23673 = n2222 & ~n5164 ;
  assign n23674 = ~n23672 & ~n23673 ;
  assign n23675 = n2377 & ~n23674 ;
  assign n23680 = \P1_InstQueue_reg[1][5]/NET0131  & n1955 ;
  assign n23681 = \P1_InstQueue_reg[14][5]/NET0131  & n1949 ;
  assign n23694 = ~n23680 & ~n23681 ;
  assign n23682 = \P1_InstQueue_reg[11][5]/NET0131  & n1974 ;
  assign n23683 = \P1_InstQueue_reg[3][5]/NET0131  & n1958 ;
  assign n23695 = ~n23682 & ~n23683 ;
  assign n23702 = n23694 & n23695 ;
  assign n23676 = \P1_InstQueue_reg[15][5]/NET0131  & n1953 ;
  assign n23677 = \P1_InstQueue_reg[4][5]/NET0131  & n1966 ;
  assign n23692 = ~n23676 & ~n23677 ;
  assign n23678 = \P1_InstQueue_reg[0][5]/NET0131  & n1980 ;
  assign n23679 = \P1_InstQueue_reg[9][5]/NET0131  & n1972 ;
  assign n23693 = ~n23678 & ~n23679 ;
  assign n23703 = n23692 & n23693 ;
  assign n23704 = n23702 & n23703 ;
  assign n23688 = \P1_InstQueue_reg[13][5]/NET0131  & n1946 ;
  assign n23689 = \P1_InstQueue_reg[6][5]/NET0131  & n1976 ;
  assign n23698 = ~n23688 & ~n23689 ;
  assign n23690 = \P1_InstQueue_reg[7][5]/NET0131  & n1961 ;
  assign n23691 = \P1_InstQueue_reg[5][5]/NET0131  & n1970 ;
  assign n23699 = ~n23690 & ~n23691 ;
  assign n23700 = n23698 & n23699 ;
  assign n23684 = \P1_InstQueue_reg[10][5]/NET0131  & n1968 ;
  assign n23685 = \P1_InstQueue_reg[12][5]/NET0131  & n1978 ;
  assign n23696 = ~n23684 & ~n23685 ;
  assign n23686 = \P1_InstQueue_reg[2][5]/NET0131  & n1982 ;
  assign n23687 = \P1_InstQueue_reg[8][5]/NET0131  & n1964 ;
  assign n23697 = ~n23686 & ~n23687 ;
  assign n23701 = n23696 & n23697 ;
  assign n23705 = n23700 & n23701 ;
  assign n23706 = n23704 & n23705 ;
  assign n23707 = n2337 & ~n23706 ;
  assign n23708 = n2331 & n23707 ;
  assign n23709 = ~n23675 & ~n23708 ;
  assign n23710 = ~n23667 & n23709 ;
  assign n23711 = ~n23671 & n23710 ;
  assign n23712 = n2432 & ~n23711 ;
  assign n23713 = ~n23666 & ~n23712 ;
  assign n23714 = \P1_EAX_reg[22]/NET0131  & ~n15402 ;
  assign n23748 = ~\P1_EAX_reg[22]/NET0131  & ~n23669 ;
  assign n23749 = n2260 & ~n15916 ;
  assign n23750 = ~n23748 & n23749 ;
  assign n23751 = \P1_EAX_reg[22]/NET0131  & ~n15925 ;
  assign n23719 = \P1_InstQueue_reg[1][6]/NET0131  & n1955 ;
  assign n23720 = \P1_InstQueue_reg[14][6]/NET0131  & n1949 ;
  assign n23733 = ~n23719 & ~n23720 ;
  assign n23721 = \P1_InstQueue_reg[4][6]/NET0131  & n1966 ;
  assign n23722 = \P1_InstQueue_reg[3][6]/NET0131  & n1958 ;
  assign n23734 = ~n23721 & ~n23722 ;
  assign n23741 = n23733 & n23734 ;
  assign n23715 = \P1_InstQueue_reg[6][6]/NET0131  & n1976 ;
  assign n23716 = \P1_InstQueue_reg[11][6]/NET0131  & n1974 ;
  assign n23731 = ~n23715 & ~n23716 ;
  assign n23717 = \P1_InstQueue_reg[0][6]/NET0131  & n1980 ;
  assign n23718 = \P1_InstQueue_reg[9][6]/NET0131  & n1972 ;
  assign n23732 = ~n23717 & ~n23718 ;
  assign n23742 = n23731 & n23732 ;
  assign n23743 = n23741 & n23742 ;
  assign n23727 = \P1_InstQueue_reg[13][6]/NET0131  & n1946 ;
  assign n23728 = \P1_InstQueue_reg[7][6]/NET0131  & n1961 ;
  assign n23737 = ~n23727 & ~n23728 ;
  assign n23729 = \P1_InstQueue_reg[15][6]/NET0131  & n1953 ;
  assign n23730 = \P1_InstQueue_reg[5][6]/NET0131  & n1970 ;
  assign n23738 = ~n23729 & ~n23730 ;
  assign n23739 = n23737 & n23738 ;
  assign n23723 = \P1_InstQueue_reg[10][6]/NET0131  & n1968 ;
  assign n23724 = \P1_InstQueue_reg[12][6]/NET0131  & n1978 ;
  assign n23735 = ~n23723 & ~n23724 ;
  assign n23725 = \P1_InstQueue_reg[2][6]/NET0131  & n1982 ;
  assign n23726 = \P1_InstQueue_reg[8][6]/NET0131  & n1964 ;
  assign n23736 = ~n23725 & ~n23726 ;
  assign n23740 = n23735 & n23736 ;
  assign n23744 = n23739 & n23740 ;
  assign n23745 = n23743 & n23744 ;
  assign n23746 = n2337 & ~n23745 ;
  assign n23747 = n2331 & n23746 ;
  assign n23752 = n2302 & ~n5221 ;
  assign n23753 = n2222 & ~n5182 ;
  assign n23754 = ~n23752 & ~n23753 ;
  assign n23755 = n2377 & ~n23754 ;
  assign n23756 = ~n23747 & ~n23755 ;
  assign n23757 = ~n23751 & n23756 ;
  assign n23758 = ~n23750 & n23757 ;
  assign n23759 = n2432 & ~n23758 ;
  assign n23760 = ~n23714 & ~n23759 ;
  assign n23761 = ~n1907 & n1927 ;
  assign n23762 = \P2_More_reg/NET0131  & ~n12632 ;
  assign n23763 = ~n23761 & ~n23762 ;
  assign n23767 = ~\P2_ReadRequest_reg/NET0131  & ~n1891 ;
  assign n23765 = ~n1746 & n1804 ;
  assign n23766 = ~n1822 & n23765 ;
  assign n23768 = n1927 & ~n23766 ;
  assign n23769 = ~n23767 & n23768 ;
  assign n23764 = \P2_ReadRequest_reg/NET0131  & ~n22013 ;
  assign n23770 = n3114 & ~n23764 ;
  assign n23771 = ~n23769 & n23770 ;
  assign n23774 = n2737 & n18209 ;
  assign n23773 = ~\P3_InstQueue_reg[0][3]/NET0131  & ~n18209 ;
  assign n23775 = n2994 & ~n23773 ;
  assign n23776 = ~n23774 & n23775 ;
  assign n23772 = \P3_InstQueue_reg[0][3]/NET0131  & ~n18218 ;
  assign n23777 = \buf2_reg[27]/NET0131  & n18200 ;
  assign n23778 = \buf2_reg[19]/NET0131  & n18203 ;
  assign n23779 = ~n23777 & ~n23778 ;
  assign n23780 = n2970 & ~n23779 ;
  assign n23781 = \buf2_reg[3]/NET0131  & n18228 ;
  assign n23782 = ~n23780 & ~n23781 ;
  assign n23783 = ~n23772 & n23782 ;
  assign n23784 = ~n23776 & n23783 ;
  assign n23787 = n2508 & n18209 ;
  assign n23786 = ~\P3_InstQueue_reg[0][6]/NET0131  & ~n18209 ;
  assign n23788 = n2994 & ~n23786 ;
  assign n23789 = ~n23787 & n23788 ;
  assign n23785 = \P3_InstQueue_reg[0][6]/NET0131  & ~n18218 ;
  assign n23790 = \buf2_reg[30]/NET0131  & n18200 ;
  assign n23791 = \buf2_reg[22]/NET0131  & n18203 ;
  assign n23792 = ~n23790 & ~n23791 ;
  assign n23793 = n2970 & ~n23792 ;
  assign n23794 = \buf2_reg[6]/NET0131  & n18228 ;
  assign n23795 = ~n23793 & ~n23794 ;
  assign n23796 = ~n23785 & n23795 ;
  assign n23797 = ~n23789 & n23796 ;
  assign n23800 = n2737 & n18246 ;
  assign n23799 = ~\P3_InstQueue_reg[10][3]/NET0131  & ~n18246 ;
  assign n23801 = n2994 & ~n23799 ;
  assign n23802 = ~n23800 & n23801 ;
  assign n23798 = \P3_InstQueue_reg[10][3]/NET0131  & ~n18243 ;
  assign n23803 = \buf2_reg[27]/NET0131  & n18233 ;
  assign n23804 = \buf2_reg[19]/NET0131  & n18236 ;
  assign n23805 = ~n23803 & ~n23804 ;
  assign n23806 = n2970 & ~n23805 ;
  assign n23807 = \buf2_reg[3]/NET0131  & n18255 ;
  assign n23808 = ~n23806 & ~n23807 ;
  assign n23809 = ~n23798 & n23808 ;
  assign n23810 = ~n23802 & n23809 ;
  assign n23813 = n2508 & n18246 ;
  assign n23812 = ~\P3_InstQueue_reg[10][6]/NET0131  & ~n18246 ;
  assign n23814 = n2994 & ~n23812 ;
  assign n23815 = ~n23813 & n23814 ;
  assign n23811 = \P3_InstQueue_reg[10][6]/NET0131  & ~n18243 ;
  assign n23816 = \buf2_reg[30]/NET0131  & n18233 ;
  assign n23817 = \buf2_reg[22]/NET0131  & n18236 ;
  assign n23818 = ~n23816 & ~n23817 ;
  assign n23819 = n2970 & ~n23818 ;
  assign n23820 = \buf2_reg[6]/NET0131  & n18255 ;
  assign n23821 = ~n23819 & ~n23820 ;
  assign n23822 = ~n23811 & n23821 ;
  assign n23823 = ~n23815 & n23822 ;
  assign n23825 = n2737 & n18266 ;
  assign n23824 = ~\P3_InstQueue_reg[11][3]/NET0131  & ~n18266 ;
  assign n23826 = n2994 & ~n23824 ;
  assign n23827 = ~n23825 & n23826 ;
  assign n23833 = \P3_InstQueue_reg[11][3]/NET0131  & ~n18264 ;
  assign n23828 = ~\P3_InstQueueWr_Addr_reg[0]/NET0131  & ~\buf2_reg[27]/NET0131  ;
  assign n23829 = \P3_InstQueueWr_Addr_reg[0]/NET0131  & ~\buf2_reg[19]/NET0131  ;
  assign n23830 = ~n23828 & ~n23829 ;
  assign n23831 = n2959 & n23830 ;
  assign n23832 = n18260 & n23831 ;
  assign n23834 = \buf2_reg[3]/NET0131  & n18245 ;
  assign n23835 = n18262 & n23834 ;
  assign n23836 = ~n23832 & ~n23835 ;
  assign n23837 = ~n23833 & n23836 ;
  assign n23838 = ~n23827 & n23837 ;
  assign n23840 = n2508 & n18266 ;
  assign n23839 = ~\P3_InstQueue_reg[11][6]/NET0131  & ~n18266 ;
  assign n23841 = n2994 & ~n23839 ;
  assign n23842 = ~n23840 & n23841 ;
  assign n23848 = \P3_InstQueue_reg[11][6]/NET0131  & ~n18264 ;
  assign n23843 = ~\P3_InstQueueWr_Addr_reg[0]/NET0131  & ~\buf2_reg[30]/NET0131  ;
  assign n23844 = \P3_InstQueueWr_Addr_reg[0]/NET0131  & ~\buf2_reg[22]/NET0131  ;
  assign n23845 = ~n23843 & ~n23844 ;
  assign n23846 = n2959 & n23845 ;
  assign n23847 = n18260 & n23846 ;
  assign n23849 = \buf2_reg[6]/NET0131  & n18245 ;
  assign n23850 = n18262 & n23849 ;
  assign n23851 = ~n23847 & ~n23850 ;
  assign n23852 = ~n23848 & n23851 ;
  assign n23853 = ~n23842 & n23852 ;
  assign n23856 = n2737 & n18284 ;
  assign n23855 = ~\P3_InstQueue_reg[12][3]/NET0131  & ~n18284 ;
  assign n23857 = n2994 & ~n23855 ;
  assign n23858 = ~n23856 & n23857 ;
  assign n23854 = \P3_InstQueue_reg[12][3]/NET0131  & ~n18287 ;
  assign n23859 = \buf2_reg[19]/NET0131  & n18246 ;
  assign n23860 = \buf2_reg[27]/NET0131  & n18271 ;
  assign n23861 = ~n23859 & ~n23860 ;
  assign n23862 = n2970 & ~n23861 ;
  assign n23863 = \buf2_reg[3]/NET0131  & n18297 ;
  assign n23864 = ~n23862 & ~n23863 ;
  assign n23865 = ~n23854 & n23864 ;
  assign n23866 = ~n23858 & n23865 ;
  assign n23869 = n2508 & n18284 ;
  assign n23868 = ~\P3_InstQueue_reg[12][6]/NET0131  & ~n18284 ;
  assign n23870 = n2994 & ~n23868 ;
  assign n23871 = ~n23869 & n23870 ;
  assign n23867 = \P3_InstQueue_reg[12][6]/NET0131  & ~n18287 ;
  assign n23872 = \buf2_reg[22]/NET0131  & n18246 ;
  assign n23873 = \buf2_reg[30]/NET0131  & n18271 ;
  assign n23874 = ~n23872 & ~n23873 ;
  assign n23875 = n2970 & ~n23874 ;
  assign n23876 = \buf2_reg[6]/NET0131  & n18297 ;
  assign n23877 = ~n23875 & ~n23876 ;
  assign n23878 = ~n23867 & n23877 ;
  assign n23879 = ~n23871 & n23878 ;
  assign n23887 = n2737 & n18200 ;
  assign n23886 = ~\P3_InstQueue_reg[13][3]/NET0131  & ~n18200 ;
  assign n23888 = n2994 & ~n23886 ;
  assign n23889 = ~n23887 & n23888 ;
  assign n23883 = ~\P3_InstQueue_reg[13][3]/NET0131  & n18302 ;
  assign n23882 = ~\buf2_reg[3]/NET0131  & ~n18302 ;
  assign n23884 = n18305 & ~n23882 ;
  assign n23885 = ~n23883 & n23884 ;
  assign n23880 = n18303 & n23831 ;
  assign n23881 = \P3_InstQueue_reg[13][3]/NET0131  & ~n18217 ;
  assign n23890 = ~n23880 & ~n23881 ;
  assign n23891 = ~n23885 & n23890 ;
  assign n23892 = ~n23889 & n23891 ;
  assign n23900 = n2508 & n18200 ;
  assign n23899 = ~\P3_InstQueue_reg[13][6]/NET0131  & ~n18200 ;
  assign n23901 = n2994 & ~n23899 ;
  assign n23902 = ~n23900 & n23901 ;
  assign n23896 = ~\P3_InstQueue_reg[13][6]/NET0131  & n18302 ;
  assign n23895 = ~\buf2_reg[6]/NET0131  & ~n18302 ;
  assign n23897 = n18305 & ~n23895 ;
  assign n23898 = ~n23896 & n23897 ;
  assign n23893 = \P3_InstQueue_reg[13][6]/NET0131  & ~n18217 ;
  assign n23894 = n18303 & n23846 ;
  assign n23903 = ~n23893 & ~n23894 ;
  assign n23904 = ~n23898 & n23903 ;
  assign n23905 = ~n23902 & n23904 ;
  assign n23908 = n2737 & n18203 ;
  assign n23907 = ~\P3_InstQueue_reg[14][3]/NET0131  & ~n18203 ;
  assign n23909 = n2994 & ~n23907 ;
  assign n23910 = ~n23908 & n23909 ;
  assign n23906 = \P3_InstQueue_reg[14][3]/NET0131  & ~n18325 ;
  assign n23911 = \buf2_reg[27]/NET0131  & n18266 ;
  assign n23912 = \buf2_reg[19]/NET0131  & n18284 ;
  assign n23913 = ~n23911 & ~n23912 ;
  assign n23914 = n2970 & ~n23913 ;
  assign n23915 = \buf2_reg[3]/NET0131  & n18335 ;
  assign n23916 = ~n23914 & ~n23915 ;
  assign n23917 = ~n23906 & n23916 ;
  assign n23918 = ~n23910 & n23917 ;
  assign n23921 = n2508 & n18203 ;
  assign n23920 = ~\P3_InstQueue_reg[14][6]/NET0131  & ~n18203 ;
  assign n23922 = n2994 & ~n23920 ;
  assign n23923 = ~n23921 & n23922 ;
  assign n23919 = \P3_InstQueue_reg[14][6]/NET0131  & ~n18325 ;
  assign n23924 = \buf2_reg[30]/NET0131  & n18266 ;
  assign n23925 = \buf2_reg[22]/NET0131  & n18284 ;
  assign n23926 = ~n23924 & ~n23925 ;
  assign n23927 = n2970 & ~n23926 ;
  assign n23928 = \buf2_reg[6]/NET0131  & n18335 ;
  assign n23929 = ~n23927 & ~n23928 ;
  assign n23930 = ~n23919 & n23929 ;
  assign n23931 = ~n23923 & n23930 ;
  assign n23934 = n2737 & n18212 ;
  assign n23933 = ~\P3_InstQueue_reg[15][3]/NET0131  & ~n18212 ;
  assign n23935 = n2994 & ~n23933 ;
  assign n23936 = ~n23934 & n23935 ;
  assign n23932 = \P3_InstQueue_reg[15][3]/NET0131  & ~n18344 ;
  assign n23937 = \buf2_reg[27]/NET0131  & n18284 ;
  assign n23938 = \buf2_reg[19]/NET0131  & n18200 ;
  assign n23939 = ~n23937 & ~n23938 ;
  assign n23940 = n2970 & ~n23939 ;
  assign n23941 = \buf2_reg[3]/NET0131  & n18354 ;
  assign n23942 = ~n23940 & ~n23941 ;
  assign n23943 = ~n23932 & n23942 ;
  assign n23944 = ~n23936 & n23943 ;
  assign n23947 = n2508 & n18212 ;
  assign n23946 = ~\P3_InstQueue_reg[15][6]/NET0131  & ~n18212 ;
  assign n23948 = n2994 & ~n23946 ;
  assign n23949 = ~n23947 & n23948 ;
  assign n23945 = \P3_InstQueue_reg[15][6]/NET0131  & ~n18344 ;
  assign n23950 = \buf2_reg[30]/NET0131  & n18284 ;
  assign n23951 = \buf2_reg[22]/NET0131  & n18200 ;
  assign n23952 = ~n23950 & ~n23951 ;
  assign n23953 = n2970 & ~n23952 ;
  assign n23954 = \buf2_reg[6]/NET0131  & n18354 ;
  assign n23955 = ~n23953 & ~n23954 ;
  assign n23956 = ~n23945 & n23955 ;
  assign n23957 = ~n23949 & n23956 ;
  assign n23960 = n2737 & n18361 ;
  assign n23959 = ~\P3_InstQueue_reg[1][3]/NET0131  & ~n18361 ;
  assign n23961 = n2994 & ~n23959 ;
  assign n23962 = ~n23960 & n23961 ;
  assign n23958 = \P3_InstQueue_reg[1][3]/NET0131  & ~n18364 ;
  assign n23963 = \buf2_reg[27]/NET0131  & n18203 ;
  assign n23964 = \buf2_reg[19]/NET0131  & n18212 ;
  assign n23965 = ~n23963 & ~n23964 ;
  assign n23966 = n2970 & ~n23965 ;
  assign n23967 = \buf2_reg[3]/NET0131  & n18374 ;
  assign n23968 = ~n23966 & ~n23967 ;
  assign n23969 = ~n23958 & n23968 ;
  assign n23970 = ~n23962 & n23969 ;
  assign n23973 = n2508 & n18361 ;
  assign n23972 = ~\P3_InstQueue_reg[1][6]/NET0131  & ~n18361 ;
  assign n23974 = n2994 & ~n23972 ;
  assign n23975 = ~n23973 & n23974 ;
  assign n23971 = \P3_InstQueue_reg[1][6]/NET0131  & ~n18364 ;
  assign n23976 = \buf2_reg[30]/NET0131  & n18203 ;
  assign n23977 = \buf2_reg[22]/NET0131  & n18212 ;
  assign n23978 = ~n23976 & ~n23977 ;
  assign n23979 = n2970 & ~n23978 ;
  assign n23980 = \buf2_reg[6]/NET0131  & n18374 ;
  assign n23981 = ~n23979 & ~n23980 ;
  assign n23982 = ~n23971 & n23981 ;
  assign n23983 = ~n23975 & n23982 ;
  assign n23986 = n2737 & n18386 ;
  assign n23985 = ~\P3_InstQueue_reg[2][3]/NET0131  & ~n18386 ;
  assign n23987 = n2994 & ~n23985 ;
  assign n23988 = ~n23986 & n23987 ;
  assign n23984 = \P3_InstQueue_reg[2][3]/NET0131  & ~n18383 ;
  assign n23989 = \buf2_reg[27]/NET0131  & n18212 ;
  assign n23990 = \buf2_reg[19]/NET0131  & n18209 ;
  assign n23991 = ~n23989 & ~n23990 ;
  assign n23992 = n2970 & ~n23991 ;
  assign n23993 = \buf2_reg[3]/NET0131  & n18395 ;
  assign n23994 = ~n23992 & ~n23993 ;
  assign n23995 = ~n23984 & n23994 ;
  assign n23996 = ~n23988 & n23995 ;
  assign n23999 = n2508 & n18386 ;
  assign n23998 = ~\P3_InstQueue_reg[2][6]/NET0131  & ~n18386 ;
  assign n24000 = n2994 & ~n23998 ;
  assign n24001 = ~n23999 & n24000 ;
  assign n23997 = \P3_InstQueue_reg[2][6]/NET0131  & ~n18383 ;
  assign n24002 = \buf2_reg[30]/NET0131  & n18212 ;
  assign n24003 = \buf2_reg[22]/NET0131  & n18209 ;
  assign n24004 = ~n24002 & ~n24003 ;
  assign n24005 = n2970 & ~n24004 ;
  assign n24006 = \buf2_reg[6]/NET0131  & n18395 ;
  assign n24007 = ~n24005 & ~n24006 ;
  assign n24008 = ~n23997 & n24007 ;
  assign n24009 = ~n24001 & n24008 ;
  assign n24012 = n2737 & n18405 ;
  assign n24011 = ~\P3_InstQueue_reg[3][3]/NET0131  & ~n18405 ;
  assign n24013 = n2994 & ~n24011 ;
  assign n24014 = ~n24012 & n24013 ;
  assign n24010 = \P3_InstQueue_reg[3][3]/NET0131  & ~n18403 ;
  assign n24015 = \buf2_reg[19]/NET0131  & n18361 ;
  assign n24016 = \buf2_reg[27]/NET0131  & n18209 ;
  assign n24017 = ~n24015 & ~n24016 ;
  assign n24018 = n2970 & ~n24017 ;
  assign n24019 = \buf2_reg[3]/NET0131  & n18414 ;
  assign n24020 = ~n24018 & ~n24019 ;
  assign n24021 = ~n24010 & n24020 ;
  assign n24022 = ~n24014 & n24021 ;
  assign n24025 = n2508 & n18405 ;
  assign n24024 = ~\P3_InstQueue_reg[3][6]/NET0131  & ~n18405 ;
  assign n24026 = n2994 & ~n24024 ;
  assign n24027 = ~n24025 & n24026 ;
  assign n24023 = \P3_InstQueue_reg[3][6]/NET0131  & ~n18403 ;
  assign n24028 = \buf2_reg[22]/NET0131  & n18361 ;
  assign n24029 = \buf2_reg[30]/NET0131  & n18209 ;
  assign n24030 = ~n24028 & ~n24029 ;
  assign n24031 = n2970 & ~n24030 ;
  assign n24032 = \buf2_reg[6]/NET0131  & n18414 ;
  assign n24033 = ~n24031 & ~n24032 ;
  assign n24034 = ~n24023 & n24033 ;
  assign n24035 = ~n24027 & n24034 ;
  assign n24038 = n2737 & n18421 ;
  assign n24037 = ~\P3_InstQueue_reg[4][3]/NET0131  & ~n18421 ;
  assign n24039 = n2994 & ~n24037 ;
  assign n24040 = ~n24038 & n24039 ;
  assign n24036 = \P3_InstQueue_reg[4][3]/NET0131  & ~n18424 ;
  assign n24041 = \buf2_reg[19]/NET0131  & n18386 ;
  assign n24042 = \buf2_reg[27]/NET0131  & n18361 ;
  assign n24043 = ~n24041 & ~n24042 ;
  assign n24044 = n2970 & ~n24043 ;
  assign n24045 = \buf2_reg[3]/NET0131  & n18434 ;
  assign n24046 = ~n24044 & ~n24045 ;
  assign n24047 = ~n24036 & n24046 ;
  assign n24048 = ~n24040 & n24047 ;
  assign n24051 = n2508 & n18421 ;
  assign n24050 = ~\P3_InstQueue_reg[4][6]/NET0131  & ~n18421 ;
  assign n24052 = n2994 & ~n24050 ;
  assign n24053 = ~n24051 & n24052 ;
  assign n24049 = \P3_InstQueue_reg[4][6]/NET0131  & ~n18424 ;
  assign n24054 = \buf2_reg[22]/NET0131  & n18386 ;
  assign n24055 = \buf2_reg[30]/NET0131  & n18361 ;
  assign n24056 = ~n24054 & ~n24055 ;
  assign n24057 = n2970 & ~n24056 ;
  assign n24058 = \buf2_reg[6]/NET0131  & n18434 ;
  assign n24059 = ~n24057 & ~n24058 ;
  assign n24060 = ~n24049 & n24059 ;
  assign n24061 = ~n24053 & n24060 ;
  assign n24069 = n2737 & n18439 ;
  assign n24068 = ~\P3_InstQueue_reg[5][3]/NET0131  & ~n18439 ;
  assign n24070 = n2994 & ~n24068 ;
  assign n24071 = ~n24069 & n24070 ;
  assign n24065 = ~\P3_InstQueue_reg[5][3]/NET0131  & n18440 ;
  assign n24064 = ~\buf2_reg[3]/NET0131  & ~n18440 ;
  assign n24066 = n18443 & ~n24064 ;
  assign n24067 = ~n24065 & n24066 ;
  assign n24062 = n18441 & n23831 ;
  assign n24063 = \P3_InstQueue_reg[5][3]/NET0131  & ~n18217 ;
  assign n24072 = ~n24062 & ~n24063 ;
  assign n24073 = ~n24067 & n24072 ;
  assign n24074 = ~n24071 & n24073 ;
  assign n24082 = n2508 & n18439 ;
  assign n24081 = ~\P3_InstQueue_reg[5][6]/NET0131  & ~n18439 ;
  assign n24083 = n2994 & ~n24081 ;
  assign n24084 = ~n24082 & n24083 ;
  assign n24078 = ~\P3_InstQueue_reg[5][6]/NET0131  & n18440 ;
  assign n24077 = ~\buf2_reg[6]/NET0131  & ~n18440 ;
  assign n24079 = n18443 & ~n24077 ;
  assign n24080 = ~n24078 & n24079 ;
  assign n24075 = \P3_InstQueue_reg[5][6]/NET0131  & ~n18217 ;
  assign n24076 = n18441 & n23846 ;
  assign n24085 = ~n24075 & ~n24076 ;
  assign n24086 = ~n24080 & n24085 ;
  assign n24087 = ~n24084 & n24086 ;
  assign n24090 = n2737 & n18462 ;
  assign n24089 = ~\P3_InstQueue_reg[6][3]/NET0131  & ~n18462 ;
  assign n24091 = n2994 & ~n24089 ;
  assign n24092 = ~n24090 & n24091 ;
  assign n24088 = \P3_InstQueue_reg[6][3]/NET0131  & ~n18465 ;
  assign n24093 = \buf2_reg[27]/NET0131  & n18405 ;
  assign n24094 = \buf2_reg[19]/NET0131  & n18421 ;
  assign n24095 = ~n24093 & ~n24094 ;
  assign n24096 = n2970 & ~n24095 ;
  assign n24097 = \buf2_reg[3]/NET0131  & n18475 ;
  assign n24098 = ~n24096 & ~n24097 ;
  assign n24099 = ~n24088 & n24098 ;
  assign n24100 = ~n24092 & n24099 ;
  assign n24103 = n2508 & n18462 ;
  assign n24102 = ~\P3_InstQueue_reg[6][6]/NET0131  & ~n18462 ;
  assign n24104 = n2994 & ~n24102 ;
  assign n24105 = ~n24103 & n24104 ;
  assign n24101 = \P3_InstQueue_reg[6][6]/NET0131  & ~n18465 ;
  assign n24106 = \buf2_reg[30]/NET0131  & n18405 ;
  assign n24107 = \buf2_reg[22]/NET0131  & n18421 ;
  assign n24108 = ~n24106 & ~n24107 ;
  assign n24109 = n2970 & ~n24108 ;
  assign n24110 = \buf2_reg[6]/NET0131  & n18475 ;
  assign n24111 = ~n24109 & ~n24110 ;
  assign n24112 = ~n24101 & n24111 ;
  assign n24113 = ~n24105 & n24112 ;
  assign n24116 = n2737 & n18233 ;
  assign n24115 = ~\P3_InstQueue_reg[7][3]/NET0131  & ~n18233 ;
  assign n24117 = n2994 & ~n24115 ;
  assign n24118 = ~n24116 & n24117 ;
  assign n24114 = \P3_InstQueue_reg[7][3]/NET0131  & ~n18484 ;
  assign n24119 = \buf2_reg[27]/NET0131  & n18421 ;
  assign n24120 = \buf2_reg[19]/NET0131  & n18439 ;
  assign n24121 = ~n24119 & ~n24120 ;
  assign n24122 = n2970 & ~n24121 ;
  assign n24123 = \buf2_reg[3]/NET0131  & n18494 ;
  assign n24124 = ~n24122 & ~n24123 ;
  assign n24125 = ~n24114 & n24124 ;
  assign n24126 = ~n24118 & n24125 ;
  assign n24129 = n2508 & n18233 ;
  assign n24128 = ~\P3_InstQueue_reg[7][6]/NET0131  & ~n18233 ;
  assign n24130 = n2994 & ~n24128 ;
  assign n24131 = ~n24129 & n24130 ;
  assign n24127 = \P3_InstQueue_reg[7][6]/NET0131  & ~n18484 ;
  assign n24132 = \buf2_reg[30]/NET0131  & n18421 ;
  assign n24133 = \buf2_reg[22]/NET0131  & n18439 ;
  assign n24134 = ~n24132 & ~n24133 ;
  assign n24135 = n2970 & ~n24134 ;
  assign n24136 = \buf2_reg[6]/NET0131  & n18494 ;
  assign n24137 = ~n24135 & ~n24136 ;
  assign n24138 = ~n24127 & n24137 ;
  assign n24139 = ~n24131 & n24138 ;
  assign n24142 = n2737 & n18236 ;
  assign n24141 = ~\P3_InstQueue_reg[8][3]/NET0131  & ~n18236 ;
  assign n24143 = n2994 & ~n24141 ;
  assign n24144 = ~n24142 & n24143 ;
  assign n24140 = \P3_InstQueue_reg[8][3]/NET0131  & ~n18502 ;
  assign n24145 = \buf2_reg[27]/NET0131  & n18439 ;
  assign n24146 = \buf2_reg[19]/NET0131  & n18462 ;
  assign n24147 = ~n24145 & ~n24146 ;
  assign n24148 = n2970 & ~n24147 ;
  assign n24149 = \buf2_reg[3]/NET0131  & n18512 ;
  assign n24150 = ~n24148 & ~n24149 ;
  assign n24151 = ~n24140 & n24150 ;
  assign n24152 = ~n24144 & n24151 ;
  assign n24155 = n2508 & n18236 ;
  assign n24154 = ~\P3_InstQueue_reg[8][6]/NET0131  & ~n18236 ;
  assign n24156 = n2994 & ~n24154 ;
  assign n24157 = ~n24155 & n24156 ;
  assign n24153 = \P3_InstQueue_reg[8][6]/NET0131  & ~n18502 ;
  assign n24158 = \buf2_reg[30]/NET0131  & n18439 ;
  assign n24159 = \buf2_reg[22]/NET0131  & n18462 ;
  assign n24160 = ~n24158 & ~n24159 ;
  assign n24161 = n2970 & ~n24160 ;
  assign n24162 = \buf2_reg[6]/NET0131  & n18512 ;
  assign n24163 = ~n24161 & ~n24162 ;
  assign n24164 = ~n24153 & n24163 ;
  assign n24165 = ~n24157 & n24164 ;
  assign n24179 = n2737 & n18271 ;
  assign n24178 = ~\P3_InstQueue_reg[9][3]/NET0131  & ~n18271 ;
  assign n24180 = n2994 & ~n24178 ;
  assign n24181 = ~n24179 & n24180 ;
  assign n24170 = \buf2_reg[27]/NET0131  & n18462 ;
  assign n24171 = \buf2_reg[19]/NET0131  & n18233 ;
  assign n24172 = ~n24170 & ~n24171 ;
  assign n24173 = \P3_DataWidth_reg[1]/NET0131  & ~n24172 ;
  assign n24166 = \P3_InstQueue_reg[9][3]/NET0131  & ~n18235 ;
  assign n24167 = \buf2_reg[3]/NET0131  & n18235 ;
  assign n24168 = ~n24166 & ~n24167 ;
  assign n24174 = ~n18525 & ~n24168 ;
  assign n24175 = ~n24173 & ~n24174 ;
  assign n24176 = n2959 & ~n24175 ;
  assign n24169 = n4415 & ~n24168 ;
  assign n24177 = \P3_InstQueue_reg[9][3]/NET0131  & ~n18217 ;
  assign n24182 = ~n24169 & ~n24177 ;
  assign n24183 = ~n24176 & n24182 ;
  assign n24184 = ~n24181 & n24183 ;
  assign n24198 = n2508 & n18271 ;
  assign n24197 = ~\P3_InstQueue_reg[9][6]/NET0131  & ~n18271 ;
  assign n24199 = n2994 & ~n24197 ;
  assign n24200 = ~n24198 & n24199 ;
  assign n24189 = \buf2_reg[30]/NET0131  & n18462 ;
  assign n24190 = \buf2_reg[22]/NET0131  & n18233 ;
  assign n24191 = ~n24189 & ~n24190 ;
  assign n24192 = \P3_DataWidth_reg[1]/NET0131  & ~n24191 ;
  assign n24185 = \P3_InstQueue_reg[9][6]/NET0131  & ~n18235 ;
  assign n24186 = \buf2_reg[6]/NET0131  & n18235 ;
  assign n24187 = ~n24185 & ~n24186 ;
  assign n24193 = ~n18525 & ~n24187 ;
  assign n24194 = ~n24192 & ~n24193 ;
  assign n24195 = n2959 & ~n24194 ;
  assign n24188 = n4415 & ~n24187 ;
  assign n24196 = \P3_InstQueue_reg[9][6]/NET0131  & ~n18217 ;
  assign n24201 = ~n24188 & ~n24196 ;
  assign n24202 = ~n24195 & n24201 ;
  assign n24203 = ~n24200 & n24202 ;
  assign n24207 = \P3_PhyAddrPointer_reg[0]/NET0131  & ~n11965 ;
  assign n24208 = n14661 & ~n24207 ;
  assign n24209 = n2453 & ~n24208 ;
  assign n24204 = ~n2959 & ~n3004 ;
  assign n24205 = n20409 & n24204 ;
  assign n24206 = \P3_PhyAddrPointer_reg[0]/NET0131  & ~n24205 ;
  assign n24210 = ~n14656 & ~n24206 ;
  assign n24211 = ~n24209 & n24210 ;
  assign n24213 = ~n2815 & ~n2819 ;
  assign n24214 = \P3_ReadRequest_reg/NET0131  & ~n24213 ;
  assign n24215 = ~n2832 & ~n24214 ;
  assign n24216 = n2453 & ~n24215 ;
  assign n24212 = \P3_ReadRequest_reg/NET0131  & ~n22000 ;
  assign n24217 = n15433 & ~n24212 ;
  assign n24218 = ~n24216 & n24217 ;
  assign n24222 = n2432 & ~n12209 ;
  assign n24223 = ~n2436 & n15770 ;
  assign n24224 = n18551 & n24223 ;
  assign n24225 = ~n24222 & n24224 ;
  assign n24226 = \P1_PhyAddrPointer_reg[0]/NET0131  & ~n24225 ;
  assign n24219 = n2244 & n14728 ;
  assign n24220 = ~n14734 & ~n24219 ;
  assign n24221 = n2432 & ~n24220 ;
  assign n24227 = ~n14724 & ~n24221 ;
  assign n24228 = ~n24226 & n24227 ;
  assign n24230 = \P1_ReadRequest_reg/NET0131  & ~n7308 ;
  assign n24231 = ~n2304 & ~n24230 ;
  assign n24232 = n2432 & ~n24231 ;
  assign n24229 = \P1_ReadRequest_reg/NET0131  & ~n15987 ;
  assign n24233 = n14083 & ~n24229 ;
  assign n24234 = ~n24232 & n24233 ;
  assign n24238 = n1927 & ~n12395 ;
  assign n24239 = n1935 & ~n2985 ;
  assign n24240 = n12631 & ~n24239 ;
  assign n24241 = ~n24238 & n24240 ;
  assign n24242 = \P2_PhyAddrPointer_reg[0]/NET0131  & ~n24241 ;
  assign n24235 = n1734 & n14711 ;
  assign n24236 = ~n14714 & ~n24235 ;
  assign n24237 = n1927 & ~n24236 ;
  assign n24243 = ~n14707 & ~n24237 ;
  assign n24244 = ~n24242 & n24243 ;
  assign n24247 = n1734 & n14760 ;
  assign n24246 = \P2_PhyAddrPointer_reg[1]/NET0131  & ~n12395 ;
  assign n24248 = ~n14766 & ~n24246 ;
  assign n24249 = ~n24247 & n24248 ;
  assign n24250 = n1927 & ~n24249 ;
  assign n24251 = ~n3034 & n8958 ;
  assign n24252 = \P2_PhyAddrPointer_reg[1]/NET0131  & ~n24251 ;
  assign n24245 = ~\P2_PhyAddrPointer_reg[1]/NET0131  & n9005 ;
  assign n24253 = ~n14741 & ~n24245 ;
  assign n24254 = ~n24252 & n24253 ;
  assign n24255 = ~n24250 & n24254 ;
  assign n24258 = n2894 & n14685 ;
  assign n24257 = \P3_PhyAddrPointer_reg[1]/NET0131  & ~n11965 ;
  assign n24259 = ~n14695 & ~n24257 ;
  assign n24260 = ~n24258 & n24259 ;
  assign n24261 = n2453 & ~n24260 ;
  assign n24262 = ~n2970 & n9063 ;
  assign n24263 = \P3_PhyAddrPointer_reg[1]/NET0131  & ~n24262 ;
  assign n24256 = ~\P3_PhyAddrPointer_reg[1]/NET0131  & n10076 ;
  assign n24264 = ~n14704 & ~n24256 ;
  assign n24265 = ~n24263 & n24264 ;
  assign n24266 = ~n24261 & n24265 ;
  assign n24268 = \P1_PhyAddrPointer_reg[1]/NET0131  & ~n12209 ;
  assign n24269 = n14804 & ~n24268 ;
  assign n24270 = n2432 & ~n24269 ;
  assign n24271 = ~n3148 & n10136 ;
  assign n24272 = \P1_PhyAddrPointer_reg[1]/NET0131  & ~n24271 ;
  assign n24267 = ~\P1_PhyAddrPointer_reg[1]/NET0131  & n10133 ;
  assign n24273 = ~n14821 & ~n24267 ;
  assign n24274 = ~n24272 & n24273 ;
  assign n24275 = ~n24270 & n24274 ;
  assign n24277 = \P1_Datao_reg[19]/NET0131  & n2306 ;
  assign n24278 = ~\P1_Datao_reg[19]/NET0131  & ~n2312 ;
  assign n24279 = ~\P1_EAX_reg[19]/NET0131  & ~n16018 ;
  assign n24280 = ~n16019 & ~n24279 ;
  assign n24281 = n2312 & ~n24280 ;
  assign n24282 = ~n24278 & ~n24281 ;
  assign n24283 = n21698 & n24282 ;
  assign n24284 = ~n24277 & ~n24283 ;
  assign n24285 = n2432 & ~n24284 ;
  assign n24276 = \P1_uWord_reg[3]/NET0131  & n2440 ;
  assign n24286 = \P1_Datao_reg[19]/NET0131  & ~n16884 ;
  assign n24287 = ~n24276 & ~n24286 ;
  assign n24288 = ~n24285 & n24287 ;
  assign n24290 = \P1_Datao_reg[23]/NET0131  & ~n2313 ;
  assign n24291 = ~\P1_EAX_reg[23]/NET0131  & ~n16021 ;
  assign n24292 = n15990 & ~n16874 ;
  assign n24293 = ~n24291 & n24292 ;
  assign n24294 = ~n2311 & n24293 ;
  assign n24295 = ~n24290 & ~n24294 ;
  assign n24296 = n2432 & ~n24295 ;
  assign n24289 = \P1_uWord_reg[7]/NET0131  & n2440 ;
  assign n24297 = \P1_Datao_reg[23]/NET0131  & ~n16884 ;
  assign n24298 = ~n24289 & ~n24297 ;
  assign n24299 = ~n24296 & n24298 ;
  assign n24301 = n2453 & ~n2833 ;
  assign n24302 = n16899 & ~n24301 ;
  assign n24303 = \datao[19]_pad  & ~n24302 ;
  assign n24300 = \P3_uWord_reg[3]/NET0131  & n16888 ;
  assign n24304 = n2453 & ~n2786 ;
  assign n24305 = ~\P3_EAX_reg[19]/NET0131  & ~n16112 ;
  assign n24306 = ~n16113 & ~n24305 ;
  assign n24307 = n16094 & n24306 ;
  assign n24308 = n24304 & n24307 ;
  assign n24309 = ~n24300 & ~n24308 ;
  assign n24310 = ~n24303 & n24309 ;
  assign n24312 = \datao[23]_pad  & ~n2833 ;
  assign n24313 = \P3_EAX_reg[22]/NET0131  & n16115 ;
  assign n24314 = ~\P3_EAX_reg[23]/NET0131  & ~n24313 ;
  assign n24315 = n16094 & ~n16116 ;
  assign n24316 = ~n24314 & n24315 ;
  assign n24317 = ~n2786 & n24316 ;
  assign n24318 = ~n24312 & ~n24317 ;
  assign n24319 = n2453 & ~n24318 ;
  assign n24311 = \P3_uWord_reg[7]/NET0131  & n16888 ;
  assign n24320 = \datao[23]_pad  & ~n16899 ;
  assign n24321 = ~n24311 & ~n24320 ;
  assign n24322 = ~n24319 & n24321 ;
  assign n24324 = \P2_Datao_reg[19]/NET0131  & ~n16941 ;
  assign n24325 = ~\P2_EAX_reg[19]/NET0131  & ~n15967 ;
  assign n24326 = ~n15968 & ~n24325 ;
  assign n24327 = n15980 & n24326 ;
  assign n24328 = ~n1819 & n24327 ;
  assign n24329 = ~n24324 & ~n24328 ;
  assign n24330 = n1927 & ~n24329 ;
  assign n24323 = \P2_uWord_reg[3]/NET0131  & n16919 ;
  assign n24331 = \P2_Datao_reg[19]/NET0131  & ~n16936 ;
  assign n24332 = ~n24323 & ~n24331 ;
  assign n24333 = ~n24330 & n24332 ;
  assign n24335 = \P2_Datao_reg[23]/NET0131  & ~n16941 ;
  assign n24336 = ~\P2_EAX_reg[23]/NET0131  & ~n15970 ;
  assign n24337 = ~n16923 & ~n24336 ;
  assign n24338 = n1922 & n24337 ;
  assign n24339 = ~n24335 & ~n24338 ;
  assign n24340 = n1927 & ~n24339 ;
  assign n24334 = \P2_uWord_reg[7]/NET0131  & n16919 ;
  assign n24341 = \P2_Datao_reg[23]/NET0131  & ~n16936 ;
  assign n24342 = ~n24334 & ~n24341 ;
  assign n24343 = ~n24340 & n24342 ;
  assign n24344 = \P2_uWord_reg[3]/NET0131  & ~n15942 ;
  assign n24345 = \P2_uWord_reg[3]/NET0131  & n1805 ;
  assign n24346 = ~n22470 & ~n24345 ;
  assign n24347 = n1742 & ~n24346 ;
  assign n24348 = \P2_uWord_reg[3]/NET0131  & n15981 ;
  assign n24349 = ~n24327 & ~n24348 ;
  assign n24350 = ~n24347 & n24349 ;
  assign n24351 = n1927 & ~n24350 ;
  assign n24352 = ~n24344 & ~n24351 ;
  assign n24353 = \P2_uWord_reg[7]/NET0131  & ~n15942 ;
  assign n24355 = \P2_uWord_reg[7]/NET0131  & n1805 ;
  assign n24356 = ~n22515 & ~n24355 ;
  assign n24357 = n1742 & ~n24356 ;
  assign n24354 = n15980 & n24337 ;
  assign n24358 = \P2_uWord_reg[7]/NET0131  & n15981 ;
  assign n24359 = ~n24354 & ~n24358 ;
  assign n24360 = ~n24357 & n24359 ;
  assign n24361 = n1927 & ~n24360 ;
  assign n24362 = ~n24353 & ~n24361 ;
  assign n24363 = \P1_uWord_reg[3]/NET0131  & ~n15988 ;
  assign n24365 = \P1_uWord_reg[3]/NET0131  & n2317 ;
  assign n24366 = ~n17025 & ~n24365 ;
  assign n24367 = n2222 & ~n24366 ;
  assign n24364 = \P1_uWord_reg[3]/NET0131  & n15991 ;
  assign n24368 = n15990 & n24280 ;
  assign n24369 = ~n24364 & ~n24368 ;
  assign n24370 = ~n24367 & n24369 ;
  assign n24371 = n2432 & ~n24370 ;
  assign n24372 = ~n24363 & ~n24371 ;
  assign n24373 = \P1_uWord_reg[7]/NET0131  & ~n15988 ;
  assign n24374 = \P1_uWord_reg[7]/NET0131  & ~n15992 ;
  assign n24375 = ~n22350 & ~n24293 ;
  assign n24376 = ~n24374 & n24375 ;
  assign n24377 = n2432 & ~n24376 ;
  assign n24378 = ~n24373 & ~n24377 ;
  assign n24379 = n2453 & n14954 ;
  assign n24380 = n13810 & ~n24379 ;
  assign n24381 = \P3_EBX_reg[0]/NET0131  & ~n24380 ;
  assign n24382 = ~\P3_EBX_reg[0]/NET0131  & n2748 ;
  assign n24383 = ~n3963 & n14952 ;
  assign n24384 = ~n24382 & ~n24383 ;
  assign n24385 = n2453 & ~n24384 ;
  assign n24386 = ~n24381 & ~n24385 ;
  assign n24388 = \P3_EBX_reg[10]/NET0131  & n14954 ;
  assign n24387 = n14952 & ~n17016 ;
  assign n24389 = ~\P3_EBX_reg[10]/NET0131  & ~n14965 ;
  assign n24390 = n2748 & ~n14966 ;
  assign n24391 = ~n24389 & n24390 ;
  assign n24392 = ~n24387 & ~n24391 ;
  assign n24393 = ~n24388 & n24392 ;
  assign n24394 = n2453 & ~n24393 ;
  assign n24395 = \P3_EBX_reg[10]/NET0131  & ~n13810 ;
  assign n24396 = ~n24394 & ~n24395 ;
  assign n24397 = \P3_EBX_reg[11]/NET0131  & ~n13810 ;
  assign n24399 = ~n14954 & ~n24390 ;
  assign n24400 = \P3_EBX_reg[11]/NET0131  & ~n24399 ;
  assign n24398 = n14952 & ~n17070 ;
  assign n24401 = ~\P3_EBX_reg[11]/NET0131  & n14966 ;
  assign n24402 = n2748 & n24401 ;
  assign n24403 = ~n24398 & ~n24402 ;
  assign n24404 = ~n24400 & n24403 ;
  assign n24405 = n2453 & ~n24404 ;
  assign n24406 = ~n24397 & ~n24405 ;
  assign n24408 = \P3_EBX_reg[12]/NET0131  & n14954 ;
  assign n24407 = n14952 & ~n17109 ;
  assign n24409 = ~\P3_EBX_reg[12]/NET0131  & ~n14967 ;
  assign n24410 = n2748 & ~n14968 ;
  assign n24411 = ~n24409 & n24410 ;
  assign n24412 = ~n24407 & ~n24411 ;
  assign n24413 = ~n24408 & n24412 ;
  assign n24414 = n2453 & ~n24413 ;
  assign n24415 = \P3_EBX_reg[12]/NET0131  & ~n13810 ;
  assign n24416 = ~n24414 & ~n24415 ;
  assign n24417 = \P3_EBX_reg[13]/NET0131  & ~n13810 ;
  assign n24419 = ~n14954 & ~n24410 ;
  assign n24420 = \P3_EBX_reg[13]/NET0131  & ~n24419 ;
  assign n24418 = n14952 & ~n17156 ;
  assign n24421 = ~\P3_EBX_reg[13]/NET0131  & n2748 ;
  assign n24422 = n14968 & n24421 ;
  assign n24423 = ~n24418 & ~n24422 ;
  assign n24424 = ~n24420 & n24423 ;
  assign n24425 = n2453 & ~n24424 ;
  assign n24426 = ~n24417 & ~n24425 ;
  assign n24429 = ~\P3_EBX_reg[14]/NET0131  & ~n14969 ;
  assign n24430 = n2748 & ~n14970 ;
  assign n24431 = ~n24429 & n24430 ;
  assign n24427 = \P3_EBX_reg[14]/NET0131  & n14954 ;
  assign n24428 = n14952 & ~n17198 ;
  assign n24432 = ~n24427 & ~n24428 ;
  assign n24433 = ~n24431 & n24432 ;
  assign n24434 = n2453 & ~n24433 ;
  assign n24435 = \P3_EBX_reg[14]/NET0131  & ~n13810 ;
  assign n24436 = ~n24434 & ~n24435 ;
  assign n24439 = ~\P3_EBX_reg[15]/NET0131  & ~n14970 ;
  assign n24440 = n2748 & ~n14971 ;
  assign n24441 = ~n24439 & n24440 ;
  assign n24437 = \P3_EBX_reg[15]/NET0131  & n14954 ;
  assign n24438 = n14952 & ~n17243 ;
  assign n24442 = ~n24437 & ~n24438 ;
  assign n24443 = ~n24441 & n24442 ;
  assign n24444 = n2453 & ~n24443 ;
  assign n24445 = \P3_EBX_reg[15]/NET0131  & ~n13810 ;
  assign n24446 = ~n24444 & ~n24445 ;
  assign n24449 = ~\P3_EBX_reg[16]/NET0131  & ~n14971 ;
  assign n24450 = n2748 & ~n14972 ;
  assign n24451 = ~n24449 & n24450 ;
  assign n24447 = \P3_EBX_reg[16]/NET0131  & n14954 ;
  assign n24448 = n14952 & ~n22616 ;
  assign n24452 = ~n24447 & ~n24448 ;
  assign n24453 = ~n24451 & n24452 ;
  assign n24454 = n2453 & ~n24453 ;
  assign n24455 = \P3_EBX_reg[16]/NET0131  & ~n13810 ;
  assign n24456 = ~n24454 & ~n24455 ;
  assign n24458 = ~\P3_EBX_reg[17]/NET0131  & ~n14972 ;
  assign n24459 = n2748 & ~n14973 ;
  assign n24460 = ~n24458 & n24459 ;
  assign n24457 = n14952 & ~n22671 ;
  assign n24461 = \P3_EBX_reg[17]/NET0131  & n14954 ;
  assign n24462 = ~n24457 & ~n24461 ;
  assign n24463 = ~n24460 & n24462 ;
  assign n24464 = n2453 & ~n24463 ;
  assign n24465 = \P3_EBX_reg[17]/NET0131  & ~n13810 ;
  assign n24466 = ~n24464 & ~n24465 ;
  assign n24467 = \P3_EBX_reg[18]/NET0131  & ~n13810 ;
  assign n24469 = ~n14954 & ~n24459 ;
  assign n24470 = \P3_EBX_reg[18]/NET0131  & ~n24469 ;
  assign n24468 = n14952 & ~n22719 ;
  assign n24471 = ~\P3_EBX_reg[18]/NET0131  & n2748 ;
  assign n24472 = n14973 & n24471 ;
  assign n24473 = ~n24468 & ~n24472 ;
  assign n24474 = ~n24470 & n24473 ;
  assign n24475 = n2453 & ~n24474 ;
  assign n24476 = ~n24467 & ~n24475 ;
  assign n24479 = ~\P3_EBX_reg[19]/NET0131  & ~n14974 ;
  assign n24480 = n2748 & ~n14975 ;
  assign n24481 = ~n24479 & n24480 ;
  assign n24477 = \P3_EBX_reg[19]/NET0131  & n14954 ;
  assign n24478 = n14952 & ~n22768 ;
  assign n24482 = ~n24477 & ~n24478 ;
  assign n24483 = ~n24481 & n24482 ;
  assign n24484 = n2453 & ~n24483 ;
  assign n24485 = \P3_EBX_reg[19]/NET0131  & ~n13810 ;
  assign n24486 = ~n24484 & ~n24485 ;
  assign n24488 = \P3_EBX_reg[1]/NET0131  & n14954 ;
  assign n24487 = n2748 & n20810 ;
  assign n24489 = ~n3930 & n14952 ;
  assign n24490 = ~n24487 & ~n24489 ;
  assign n24491 = ~n24488 & n24490 ;
  assign n24492 = n2453 & ~n24491 ;
  assign n24493 = \P3_EBX_reg[1]/NET0131  & ~n13810 ;
  assign n24494 = ~n24492 & ~n24493 ;
  assign n24498 = ~\P3_EBX_reg[20]/NET0131  & ~n14975 ;
  assign n24497 = \P3_EBX_reg[20]/NET0131  & n14975 ;
  assign n24499 = n2748 & ~n24497 ;
  assign n24500 = ~n24498 & n24499 ;
  assign n24495 = \P3_EBX_reg[20]/NET0131  & n14954 ;
  assign n24496 = n14952 & ~n22813 ;
  assign n24501 = ~n24495 & ~n24496 ;
  assign n24502 = ~n24500 & n24501 ;
  assign n24503 = n2453 & ~n24502 ;
  assign n24504 = \P3_EBX_reg[20]/NET0131  & ~n13810 ;
  assign n24505 = ~n24503 & ~n24504 ;
  assign n24509 = \P3_EBX_reg[21]/NET0131  & n24497 ;
  assign n24508 = ~\P3_EBX_reg[21]/NET0131  & ~n24497 ;
  assign n24510 = n2748 & ~n24508 ;
  assign n24511 = ~n24509 & n24510 ;
  assign n24506 = \P3_EBX_reg[21]/NET0131  & n14954 ;
  assign n24507 = n14952 & ~n22863 ;
  assign n24512 = ~n24506 & ~n24507 ;
  assign n24513 = ~n24511 & n24512 ;
  assign n24514 = n2453 & ~n24513 ;
  assign n24515 = \P3_EBX_reg[21]/NET0131  & ~n13810 ;
  assign n24516 = ~n24514 & ~n24515 ;
  assign n24520 = \P3_EBX_reg[22]/NET0131  & n24509 ;
  assign n24519 = ~\P3_EBX_reg[22]/NET0131  & ~n24509 ;
  assign n24521 = n2748 & ~n24519 ;
  assign n24522 = ~n24520 & n24521 ;
  assign n24517 = \P3_EBX_reg[22]/NET0131  & n14954 ;
  assign n24518 = n14952 & ~n22905 ;
  assign n24523 = ~n24517 & ~n24518 ;
  assign n24524 = ~n24522 & n24523 ;
  assign n24525 = n2453 & ~n24524 ;
  assign n24526 = \P3_EBX_reg[22]/NET0131  & ~n13810 ;
  assign n24527 = ~n24525 & ~n24526 ;
  assign n24528 = \P3_EBX_reg[23]/NET0131  & ~n13810 ;
  assign n24531 = ~\P3_EBX_reg[23]/NET0131  & ~n24520 ;
  assign n24532 = n2748 & ~n14979 ;
  assign n24533 = ~n24531 & n24532 ;
  assign n24529 = \P3_EBX_reg[23]/NET0131  & n14954 ;
  assign n24530 = n14952 & n22925 ;
  assign n24534 = ~n24529 & ~n24530 ;
  assign n24535 = ~n24533 & n24534 ;
  assign n24536 = n2453 & ~n24535 ;
  assign n24537 = ~n24528 & ~n24536 ;
  assign n24540 = ~\P3_EBX_reg[24]/NET0131  & ~n14979 ;
  assign n24541 = n2748 & ~n14980 ;
  assign n24542 = ~n24540 & n24541 ;
  assign n24538 = \P3_EBX_reg[24]/NET0131  & n14954 ;
  assign n24539 = n14952 & n22946 ;
  assign n24543 = ~n24538 & ~n24539 ;
  assign n24544 = ~n24542 & n24543 ;
  assign n24545 = n2453 & ~n24544 ;
  assign n24546 = \P3_EBX_reg[24]/NET0131  & ~n13810 ;
  assign n24547 = ~n24545 & ~n24546 ;
  assign n24548 = \P3_EBX_reg[28]/NET0131  & ~n13810 ;
  assign n24549 = n2748 & ~n17454 ;
  assign n24550 = ~n14954 & ~n24549 ;
  assign n24551 = \P3_EBX_reg[28]/NET0131  & ~n24550 ;
  assign n24552 = n14952 & n22973 ;
  assign n24553 = ~\P3_EBX_reg[28]/NET0131  & n2748 ;
  assign n24554 = n17454 & n24553 ;
  assign n24555 = ~n24552 & ~n24554 ;
  assign n24556 = ~n24551 & n24555 ;
  assign n24557 = n2453 & ~n24556 ;
  assign n24558 = ~n24548 & ~n24557 ;
  assign n24560 = \P3_EBX_reg[2]/NET0131  & n14954 ;
  assign n24559 = ~n3896 & n14952 ;
  assign n24561 = ~\P3_EBX_reg[2]/NET0131  & ~n14957 ;
  assign n24562 = ~n14958 & ~n24561 ;
  assign n24563 = n2748 & n24562 ;
  assign n24564 = ~n24559 & ~n24563 ;
  assign n24565 = ~n24560 & n24564 ;
  assign n24566 = n2453 & ~n24565 ;
  assign n24567 = \P3_EBX_reg[2]/NET0131  & ~n13810 ;
  assign n24568 = ~n24566 & ~n24567 ;
  assign n24570 = \P3_EBX_reg[3]/NET0131  & n14954 ;
  assign n24569 = ~n4032 & n14952 ;
  assign n24571 = ~\P3_EBX_reg[3]/NET0131  & ~n14958 ;
  assign n24572 = ~n14959 & ~n24571 ;
  assign n24573 = n2748 & n24572 ;
  assign n24574 = ~n24569 & ~n24573 ;
  assign n24575 = ~n24570 & n24574 ;
  assign n24576 = n2453 & ~n24575 ;
  assign n24577 = \P3_EBX_reg[3]/NET0131  & ~n13810 ;
  assign n24578 = ~n24576 & ~n24577 ;
  assign n24580 = \P3_EBX_reg[4]/NET0131  & n14954 ;
  assign n24579 = ~n4000 & n14952 ;
  assign n24581 = ~\P3_EBX_reg[4]/NET0131  & ~n14959 ;
  assign n24582 = ~n14960 & ~n24581 ;
  assign n24583 = n2748 & n24582 ;
  assign n24584 = ~n24579 & ~n24583 ;
  assign n24585 = ~n24580 & n24584 ;
  assign n24586 = n2453 & ~n24585 ;
  assign n24587 = \P3_EBX_reg[4]/NET0131  & ~n13810 ;
  assign n24588 = ~n24586 & ~n24587 ;
  assign n24590 = \P3_EBX_reg[5]/NET0131  & n14954 ;
  assign n24589 = ~n3830 & n14952 ;
  assign n24591 = ~\P3_EBX_reg[5]/NET0131  & ~n14960 ;
  assign n24592 = ~n14961 & ~n24591 ;
  assign n24593 = n2748 & n24592 ;
  assign n24594 = ~n24589 & ~n24593 ;
  assign n24595 = ~n24590 & n24594 ;
  assign n24596 = n2453 & ~n24595 ;
  assign n24597 = \P3_EBX_reg[5]/NET0131  & ~n13810 ;
  assign n24598 = ~n24596 & ~n24597 ;
  assign n24600 = \P3_EBX_reg[6]/NET0131  & n14954 ;
  assign n24599 = ~n3864 & n14952 ;
  assign n24601 = ~\P3_EBX_reg[6]/NET0131  & ~n14961 ;
  assign n24602 = ~n14962 & ~n24601 ;
  assign n24603 = n2748 & n24602 ;
  assign n24604 = ~n24599 & ~n24603 ;
  assign n24605 = ~n24600 & n24604 ;
  assign n24606 = n2453 & ~n24605 ;
  assign n24607 = \P3_EBX_reg[6]/NET0131  & ~n13810 ;
  assign n24608 = ~n24606 & ~n24607 ;
  assign n24610 = \P3_EBX_reg[7]/NET0131  & n14954 ;
  assign n24609 = ~n3753 & n14952 ;
  assign n24611 = ~\P3_EBX_reg[7]/NET0131  & ~n14962 ;
  assign n24612 = ~n14963 & ~n24611 ;
  assign n24613 = n2748 & n24612 ;
  assign n24614 = ~n24609 & ~n24613 ;
  assign n24615 = ~n24610 & n24614 ;
  assign n24616 = n2453 & ~n24615 ;
  assign n24617 = \P3_EBX_reg[7]/NET0131  & ~n13810 ;
  assign n24618 = ~n24616 & ~n24617 ;
  assign n24620 = \P3_EBX_reg[8]/NET0131  & n14954 ;
  assign n24619 = n14952 & ~n17388 ;
  assign n24621 = ~\P3_EBX_reg[8]/NET0131  & ~n14963 ;
  assign n24622 = ~n14964 & ~n24621 ;
  assign n24623 = n2748 & n24622 ;
  assign n24624 = ~n24619 & ~n24623 ;
  assign n24625 = ~n24620 & n24624 ;
  assign n24626 = n2453 & ~n24625 ;
  assign n24627 = \P3_EBX_reg[8]/NET0131  & ~n13810 ;
  assign n24628 = ~n24626 & ~n24627 ;
  assign n24630 = \P3_EBX_reg[9]/NET0131  & n14954 ;
  assign n24629 = n14952 & ~n17429 ;
  assign n24631 = ~\P3_EBX_reg[9]/NET0131  & ~n14964 ;
  assign n24632 = ~n14965 & ~n24631 ;
  assign n24633 = n2748 & n24632 ;
  assign n24634 = ~n24629 & ~n24633 ;
  assign n24635 = ~n24630 & n24634 ;
  assign n24636 = n2453 & ~n24635 ;
  assign n24637 = \P3_EBX_reg[9]/NET0131  & ~n13810 ;
  assign n24638 = ~n24636 & ~n24637 ;
  assign n24639 = n2432 & ~n15073 ;
  assign n24640 = n15402 & ~n24639 ;
  assign n24641 = \P1_EBX_reg[0]/NET0131  & ~n24640 ;
  assign n24642 = ~\P1_EBX_reg[0]/NET0131  & n2262 ;
  assign n24643 = n2242 & n23384 ;
  assign n24644 = ~n24642 & ~n24643 ;
  assign n24645 = n2432 & ~n24644 ;
  assign n24646 = ~n24641 & ~n24645 ;
  assign n24648 = \P1_EBX_reg[10]/NET0131  & ~n15073 ;
  assign n24647 = n2242 & n17858 ;
  assign n24649 = ~\P1_EBX_reg[10]/NET0131  & ~n15372 ;
  assign n24650 = ~n15373 & ~n24649 ;
  assign n24651 = n2262 & n24650 ;
  assign n24652 = ~n24647 & ~n24651 ;
  assign n24653 = ~n24648 & n24652 ;
  assign n24654 = n2432 & ~n24653 ;
  assign n24655 = \P1_EBX_reg[10]/NET0131  & ~n15402 ;
  assign n24656 = ~n24654 & ~n24655 ;
  assign n24658 = \P1_EBX_reg[11]/NET0131  & ~n15073 ;
  assign n24657 = n2242 & n18014 ;
  assign n24659 = ~\P1_EBX_reg[11]/NET0131  & ~n15373 ;
  assign n24660 = n2262 & ~n15374 ;
  assign n24661 = ~n24659 & n24660 ;
  assign n24662 = ~n24657 & ~n24661 ;
  assign n24663 = ~n24658 & n24662 ;
  assign n24664 = n2432 & ~n24663 ;
  assign n24665 = \P1_EBX_reg[11]/NET0131  & ~n15402 ;
  assign n24666 = ~n24664 & ~n24665 ;
  assign n24667 = \P1_EBX_reg[12]/NET0131  & ~n15402 ;
  assign n24669 = n15073 & ~n24660 ;
  assign n24670 = \P1_EBX_reg[12]/NET0131  & ~n24669 ;
  assign n24668 = n2242 & n18166 ;
  assign n24671 = ~\P1_EBX_reg[12]/NET0131  & n2262 ;
  assign n24672 = n15374 & n24671 ;
  assign n24673 = ~n24668 & ~n24672 ;
  assign n24674 = ~n24670 & n24673 ;
  assign n24675 = n2432 & ~n24674 ;
  assign n24676 = ~n24667 & ~n24675 ;
  assign n24678 = n2262 & ~n15376 ;
  assign n24679 = n15073 & ~n24678 ;
  assign n24680 = \P1_EBX_reg[14]/NET0131  & ~n24679 ;
  assign n24677 = n2242 & n18080 ;
  assign n24681 = ~\P1_EBX_reg[14]/NET0131  & n2262 ;
  assign n24682 = n15376 & n24681 ;
  assign n24683 = ~n24677 & ~n24682 ;
  assign n24684 = ~n24680 & n24683 ;
  assign n24685 = n2432 & ~n24684 ;
  assign n24686 = \P1_EBX_reg[14]/NET0131  & ~n15402 ;
  assign n24687 = ~n24685 & ~n24686 ;
  assign n24689 = ~\P1_EBX_reg[13]/NET0131  & ~n15375 ;
  assign n24690 = n24678 & ~n24689 ;
  assign n24688 = \P1_EBX_reg[13]/NET0131  & ~n15073 ;
  assign n24691 = n2242 & n18122 ;
  assign n24692 = ~n24688 & ~n24691 ;
  assign n24693 = ~n24690 & n24692 ;
  assign n24694 = n2432 & ~n24693 ;
  assign n24695 = \P1_EBX_reg[13]/NET0131  & ~n15402 ;
  assign n24696 = ~n24694 & ~n24695 ;
  assign n24699 = ~\P1_EBX_reg[15]/NET0131  & ~n15377 ;
  assign n24700 = n2262 & ~n15378 ;
  assign n24701 = ~n24699 & n24700 ;
  assign n24697 = \P1_EBX_reg[15]/NET0131  & ~n15073 ;
  assign n24698 = n2242 & n16478 ;
  assign n24702 = ~n24697 & ~n24698 ;
  assign n24703 = ~n24701 & n24702 ;
  assign n24704 = n2432 & ~n24703 ;
  assign n24705 = \P1_EBX_reg[15]/NET0131  & ~n15402 ;
  assign n24706 = ~n24704 & ~n24705 ;
  assign n24709 = ~\P1_EBX_reg[16]/NET0131  & ~n15378 ;
  assign n24710 = n2262 & ~n15379 ;
  assign n24711 = ~n24709 & n24710 ;
  assign n24707 = n2242 & n23466 ;
  assign n24708 = \P1_EBX_reg[16]/NET0131  & ~n15073 ;
  assign n24712 = ~n24707 & ~n24708 ;
  assign n24713 = ~n24711 & n24712 ;
  assign n24714 = n2432 & ~n24713 ;
  assign n24715 = \P1_EBX_reg[16]/NET0131  & ~n15402 ;
  assign n24716 = ~n24714 & ~n24715 ;
  assign n24719 = ~\P1_EBX_reg[17]/NET0131  & ~n15379 ;
  assign n24720 = n2262 & ~n15380 ;
  assign n24721 = ~n24719 & n24720 ;
  assign n24717 = \P1_EBX_reg[17]/NET0131  & ~n15073 ;
  assign n24718 = n2242 & n23510 ;
  assign n24722 = ~n24717 & ~n24718 ;
  assign n24723 = ~n24721 & n24722 ;
  assign n24724 = n2432 & ~n24723 ;
  assign n24725 = \P1_EBX_reg[17]/NET0131  & ~n15402 ;
  assign n24726 = ~n24724 & ~n24725 ;
  assign n24728 = ~\P1_EBX_reg[19]/NET0131  & ~n15381 ;
  assign n24729 = n2262 & ~n15382 ;
  assign n24730 = ~n24728 & n24729 ;
  assign n24727 = \P1_EBX_reg[19]/NET0131  & ~n15073 ;
  assign n24731 = n2242 & n23561 ;
  assign n24732 = ~n24727 & ~n24731 ;
  assign n24733 = ~n24730 & n24732 ;
  assign n24734 = n2432 & ~n24733 ;
  assign n24735 = \P1_EBX_reg[19]/NET0131  & ~n15402 ;
  assign n24736 = ~n24734 & ~n24735 ;
  assign n24739 = ~\P1_EBX_reg[18]/NET0131  & ~n15380 ;
  assign n24740 = n2262 & ~n15381 ;
  assign n24741 = ~n24739 & n24740 ;
  assign n24737 = \P1_EBX_reg[18]/NET0131  & ~n15073 ;
  assign n24738 = n2242 & n23604 ;
  assign n24742 = ~n24737 & ~n24738 ;
  assign n24743 = ~n24741 & n24742 ;
  assign n24744 = n2432 & ~n24743 ;
  assign n24745 = \P1_EBX_reg[18]/NET0131  & ~n15402 ;
  assign n24746 = ~n24744 & ~n24745 ;
  assign n24748 = \P1_EBX_reg[1]/NET0131  & ~n15073 ;
  assign n24747 = n2242 & n18189 ;
  assign n24749 = n2262 & n18816 ;
  assign n24750 = ~n24747 & ~n24749 ;
  assign n24751 = ~n24748 & n24750 ;
  assign n24752 = n2432 & ~n24751 ;
  assign n24753 = \P1_EBX_reg[1]/NET0131  & ~n15402 ;
  assign n24754 = ~n24752 & ~n24753 ;
  assign n24755 = \P1_EBX_reg[20]/NET0131  & ~n15402 ;
  assign n24757 = n15073 & ~n24729 ;
  assign n24758 = \P1_EBX_reg[20]/NET0131  & ~n24757 ;
  assign n24756 = n2242 & n23659 ;
  assign n24759 = ~\P1_EBX_reg[20]/NET0131  & n2262 ;
  assign n24760 = n15382 & n24759 ;
  assign n24761 = ~n24756 & ~n24760 ;
  assign n24762 = ~n24758 & n24761 ;
  assign n24763 = n2432 & ~n24762 ;
  assign n24764 = ~n24755 & ~n24763 ;
  assign n24767 = \P1_EBX_reg[20]/NET0131  & n15382 ;
  assign n24769 = \P1_EBX_reg[21]/NET0131  & n24767 ;
  assign n24768 = ~\P1_EBX_reg[21]/NET0131  & ~n24767 ;
  assign n24770 = n2262 & ~n24768 ;
  assign n24771 = ~n24769 & n24770 ;
  assign n24765 = \P1_EBX_reg[21]/NET0131  & ~n15073 ;
  assign n24766 = n2242 & n23707 ;
  assign n24772 = ~n24765 & ~n24766 ;
  assign n24773 = ~n24771 & n24772 ;
  assign n24774 = n2432 & ~n24773 ;
  assign n24775 = \P1_EBX_reg[21]/NET0131  & ~n15402 ;
  assign n24776 = ~n24774 & ~n24775 ;
  assign n24780 = \P1_EBX_reg[22]/NET0131  & n24769 ;
  assign n24779 = ~\P1_EBX_reg[22]/NET0131  & ~n24769 ;
  assign n24781 = n2262 & ~n24779 ;
  assign n24782 = ~n24780 & n24781 ;
  assign n24777 = \P1_EBX_reg[22]/NET0131  & ~n15073 ;
  assign n24778 = n2242 & n23746 ;
  assign n24783 = ~n24777 & ~n24778 ;
  assign n24784 = ~n24782 & n24783 ;
  assign n24785 = n2432 & ~n24784 ;
  assign n24786 = \P1_EBX_reg[22]/NET0131  & ~n15402 ;
  assign n24787 = ~n24785 & ~n24786 ;
  assign n24790 = ~\P1_EBX_reg[23]/NET0131  & ~n24780 ;
  assign n24791 = n2262 & ~n15386 ;
  assign n24792 = ~n24790 & n24791 ;
  assign n24788 = n2242 & n22343 ;
  assign n24789 = \P1_EBX_reg[23]/NET0131  & ~n15073 ;
  assign n24793 = ~n24788 & ~n24789 ;
  assign n24794 = ~n24792 & n24793 ;
  assign n24795 = n2432 & ~n24794 ;
  assign n24796 = \P1_EBX_reg[23]/NET0131  & ~n15402 ;
  assign n24797 = ~n24795 & ~n24796 ;
  assign n24800 = ~\P1_EBX_reg[24]/NET0131  & ~n15386 ;
  assign n24801 = n2262 & ~n15387 ;
  assign n24802 = ~n24800 & n24801 ;
  assign n24798 = \P1_EBX_reg[24]/NET0131  & ~n15073 ;
  assign n24799 = n2242 & n22393 ;
  assign n24803 = ~n24798 & ~n24799 ;
  assign n24804 = ~n24802 & n24803 ;
  assign n24805 = n2432 & ~n24804 ;
  assign n24806 = \P1_EBX_reg[24]/NET0131  & ~n15402 ;
  assign n24807 = ~n24805 & ~n24806 ;
  assign n24808 = n1927 & ~n15019 ;
  assign n24809 = n12632 & ~n24808 ;
  assign n24810 = \P2_EBX_reg[0]/NET0131  & ~n24809 ;
  assign n24811 = ~\P2_EBX_reg[0]/NET0131  & n1766 ;
  assign n24812 = n1722 & n17442 ;
  assign n24813 = ~n24811 & ~n24812 ;
  assign n24814 = n1927 & ~n24813 ;
  assign n24815 = ~n24810 & ~n24814 ;
  assign n24817 = \P2_EBX_reg[10]/NET0131  & ~n15019 ;
  assign n24816 = n1722 & n17540 ;
  assign n24818 = ~\P2_EBX_reg[10]/NET0131  & ~n15030 ;
  assign n24819 = n1766 & ~n15031 ;
  assign n24820 = ~n24818 & n24819 ;
  assign n24821 = ~n24816 & ~n24820 ;
  assign n24822 = ~n24817 & n24821 ;
  assign n24823 = n1927 & ~n24822 ;
  assign n24824 = \P2_EBX_reg[10]/NET0131  & ~n12632 ;
  assign n24825 = ~n24823 & ~n24824 ;
  assign n24827 = n15019 & ~n24819 ;
  assign n24828 = \P2_EBX_reg[11]/NET0131  & ~n24827 ;
  assign n24826 = n1722 & n17582 ;
  assign n24829 = ~\P2_EBX_reg[11]/NET0131  & n1766 ;
  assign n24830 = n15031 & n24829 ;
  assign n24831 = ~n24826 & ~n24830 ;
  assign n24832 = ~n24828 & n24831 ;
  assign n24833 = n1927 & ~n24832 ;
  assign n24834 = \P2_EBX_reg[11]/NET0131  & ~n12632 ;
  assign n24835 = ~n24833 & ~n24834 ;
  assign n24838 = ~\P2_EBX_reg[12]/NET0131  & ~n15032 ;
  assign n24839 = n1766 & ~n15033 ;
  assign n24840 = ~n24838 & n24839 ;
  assign n24836 = n1722 & n17628 ;
  assign n24837 = \P2_EBX_reg[12]/NET0131  & ~n15019 ;
  assign n24841 = ~n24836 & ~n24837 ;
  assign n24842 = ~n24840 & n24841 ;
  assign n24843 = n1927 & ~n24842 ;
  assign n24844 = \P2_EBX_reg[12]/NET0131  & ~n12632 ;
  assign n24845 = ~n24843 & ~n24844 ;
  assign n24847 = n15019 & ~n24839 ;
  assign n24848 = \P2_EBX_reg[13]/NET0131  & ~n24847 ;
  assign n24846 = n1722 & n17723 ;
  assign n24849 = ~\P2_EBX_reg[13]/NET0131  & n1766 ;
  assign n24850 = n15033 & n24849 ;
  assign n24851 = ~n24846 & ~n24850 ;
  assign n24852 = ~n24848 & n24851 ;
  assign n24853 = n1927 & ~n24852 ;
  assign n24854 = \P2_EBX_reg[13]/NET0131  & ~n12632 ;
  assign n24855 = ~n24853 & ~n24854 ;
  assign n24858 = \P2_EBX_reg[13]/NET0131  & n15033 ;
  assign n24859 = ~\P2_EBX_reg[14]/NET0131  & ~n24858 ;
  assign n24860 = n1766 & ~n15035 ;
  assign n24861 = ~n24859 & n24860 ;
  assign n24856 = n1722 & n17768 ;
  assign n24857 = \P2_EBX_reg[14]/NET0131  & ~n15019 ;
  assign n24862 = ~n24856 & ~n24857 ;
  assign n24863 = ~n24861 & n24862 ;
  assign n24864 = n1927 & ~n24863 ;
  assign n24865 = \P2_EBX_reg[14]/NET0131  & ~n12632 ;
  assign n24866 = ~n24864 & ~n24865 ;
  assign n24869 = ~\P2_EBX_reg[15]/NET0131  & ~n15035 ;
  assign n24870 = n1766 & ~n15036 ;
  assign n24871 = ~n24869 & n24870 ;
  assign n24867 = \P2_EBX_reg[15]/NET0131  & ~n15019 ;
  assign n24868 = n1722 & n16379 ;
  assign n24872 = ~n24867 & ~n24868 ;
  assign n24873 = ~n24871 & n24872 ;
  assign n24874 = n1927 & ~n24873 ;
  assign n24875 = \P2_EBX_reg[15]/NET0131  & ~n12632 ;
  assign n24876 = ~n24874 & ~n24875 ;
  assign n24879 = ~\P2_EBX_reg[16]/NET0131  & ~n15036 ;
  assign n24880 = n1766 & ~n15037 ;
  assign n24881 = ~n24879 & n24880 ;
  assign n24877 = n1722 & n23019 ;
  assign n24878 = \P2_EBX_reg[16]/NET0131  & ~n15019 ;
  assign n24882 = ~n24877 & ~n24878 ;
  assign n24883 = ~n24881 & n24882 ;
  assign n24884 = n1927 & ~n24883 ;
  assign n24885 = \P2_EBX_reg[16]/NET0131  & ~n12632 ;
  assign n24886 = ~n24884 & ~n24885 ;
  assign n24887 = \P1_EBX_reg[28]/NET0131  & ~n15402 ;
  assign n24888 = \P1_EBX_reg[27]/NET0131  & n15389 ;
  assign n24889 = n2262 & ~n24888 ;
  assign n24890 = n15073 & ~n24889 ;
  assign n24891 = \P1_EBX_reg[28]/NET0131  & ~n24890 ;
  assign n24892 = n2242 & n22566 ;
  assign n24893 = ~\P1_EBX_reg[28]/NET0131  & n2262 ;
  assign n24894 = n24888 & n24893 ;
  assign n24895 = ~n24892 & ~n24894 ;
  assign n24896 = ~n24891 & n24895 ;
  assign n24897 = n2432 & ~n24896 ;
  assign n24898 = ~n24887 & ~n24897 ;
  assign n24900 = ~\P2_EBX_reg[17]/NET0131  & ~n15037 ;
  assign n24901 = \P2_EBX_reg[17]/NET0131  & n15037 ;
  assign n24902 = n1766 & ~n24901 ;
  assign n24903 = ~n24900 & n24902 ;
  assign n24899 = n1722 & n23066 ;
  assign n24904 = \P2_EBX_reg[17]/NET0131  & ~n15019 ;
  assign n24905 = ~n24899 & ~n24904 ;
  assign n24906 = ~n24903 & n24905 ;
  assign n24907 = n1927 & ~n24906 ;
  assign n24908 = \P2_EBX_reg[17]/NET0131  & ~n12632 ;
  assign n24909 = ~n24907 & ~n24908 ;
  assign n24910 = \P2_EBX_reg[18]/NET0131  & ~n12632 ;
  assign n24912 = n15019 & ~n24902 ;
  assign n24913 = \P2_EBX_reg[18]/NET0131  & ~n24912 ;
  assign n24911 = n1722 & n23118 ;
  assign n24914 = ~\P2_EBX_reg[18]/NET0131  & n1766 ;
  assign n24915 = n24901 & n24914 ;
  assign n24916 = ~n24911 & ~n24915 ;
  assign n24917 = ~n24913 & n24916 ;
  assign n24918 = n1927 & ~n24917 ;
  assign n24919 = ~n24910 & ~n24918 ;
  assign n24922 = ~\P2_EBX_reg[19]/NET0131  & ~n15039 ;
  assign n24923 = n1766 & ~n15040 ;
  assign n24924 = ~n24922 & n24923 ;
  assign n24920 = n1722 & n23168 ;
  assign n24921 = \P2_EBX_reg[19]/NET0131  & ~n15019 ;
  assign n24925 = ~n24920 & ~n24921 ;
  assign n24926 = ~n24924 & n24925 ;
  assign n24927 = n1927 & ~n24926 ;
  assign n24928 = \P2_EBX_reg[19]/NET0131  & ~n12632 ;
  assign n24929 = ~n24927 & ~n24928 ;
  assign n24931 = \P2_EBX_reg[1]/NET0131  & ~n15019 ;
  assign n24930 = n1722 & n17782 ;
  assign n24932 = n1766 & n19580 ;
  assign n24933 = ~n24930 & ~n24932 ;
  assign n24934 = ~n24931 & n24933 ;
  assign n24935 = n1927 & ~n24934 ;
  assign n24936 = \P2_EBX_reg[1]/NET0131  & ~n12632 ;
  assign n24937 = ~n24935 & ~n24936 ;
  assign n24941 = \P2_EBX_reg[20]/NET0131  & n15040 ;
  assign n24940 = ~\P2_EBX_reg[20]/NET0131  & ~n15040 ;
  assign n24942 = n1766 & ~n24940 ;
  assign n24943 = ~n24941 & n24942 ;
  assign n24938 = \P2_EBX_reg[20]/NET0131  & ~n15019 ;
  assign n24939 = n1722 & n23219 ;
  assign n24944 = ~n24938 & ~n24939 ;
  assign n24945 = ~n24943 & n24944 ;
  assign n24946 = n1927 & ~n24945 ;
  assign n24947 = \P2_EBX_reg[20]/NET0131  & ~n12632 ;
  assign n24948 = ~n24946 & ~n24947 ;
  assign n24952 = \P2_EBX_reg[21]/NET0131  & n24941 ;
  assign n24951 = ~\P2_EBX_reg[21]/NET0131  & ~n24941 ;
  assign n24953 = n1766 & ~n24951 ;
  assign n24954 = ~n24952 & n24953 ;
  assign n24949 = \P2_EBX_reg[21]/NET0131  & ~n15019 ;
  assign n24950 = n1722 & n23275 ;
  assign n24955 = ~n24949 & ~n24950 ;
  assign n24956 = ~n24954 & n24955 ;
  assign n24957 = n1927 & ~n24956 ;
  assign n24958 = \P2_EBX_reg[21]/NET0131  & ~n12632 ;
  assign n24959 = ~n24957 & ~n24958 ;
  assign n24963 = \P2_EBX_reg[22]/NET0131  & n24952 ;
  assign n24962 = ~\P2_EBX_reg[22]/NET0131  & ~n24952 ;
  assign n24964 = n1766 & ~n24962 ;
  assign n24965 = ~n24963 & n24964 ;
  assign n24960 = n1722 & n23314 ;
  assign n24961 = \P2_EBX_reg[22]/NET0131  & ~n15019 ;
  assign n24966 = ~n24960 & ~n24961 ;
  assign n24967 = ~n24965 & n24966 ;
  assign n24968 = n1927 & ~n24967 ;
  assign n24969 = \P2_EBX_reg[22]/NET0131  & ~n12632 ;
  assign n24970 = ~n24968 & ~n24969 ;
  assign n24973 = ~\P2_EBX_reg[23]/NET0131  & ~n24963 ;
  assign n24974 = n1766 & ~n15044 ;
  assign n24975 = ~n24973 & n24974 ;
  assign n24971 = n1722 & n23340 ;
  assign n24972 = \P2_EBX_reg[23]/NET0131  & ~n15019 ;
  assign n24976 = ~n24971 & ~n24972 ;
  assign n24977 = ~n24975 & n24976 ;
  assign n24978 = n1927 & ~n24977 ;
  assign n24979 = \P2_EBX_reg[23]/NET0131  & ~n12632 ;
  assign n24980 = ~n24978 & ~n24979 ;
  assign n24982 = ~\P2_EBX_reg[24]/NET0131  & ~n15044 ;
  assign n24983 = n23405 & ~n24982 ;
  assign n24981 = \P2_EBX_reg[24]/NET0131  & n15018 ;
  assign n24984 = \P2_EBX_reg[24]/NET0131  & ~n1798 ;
  assign n24985 = ~n23350 & ~n24984 ;
  assign n24986 = n1722 & ~n24985 ;
  assign n24987 = ~n24981 & ~n24986 ;
  assign n24988 = ~n24983 & n24987 ;
  assign n24989 = n1927 & ~n24988 ;
  assign n24990 = \P2_EBX_reg[24]/NET0131  & ~n12632 ;
  assign n24991 = ~n24989 & ~n24990 ;
  assign n24993 = \P1_EBX_reg[2]/NET0131  & ~n15073 ;
  assign n24992 = n2242 & n16972 ;
  assign n24994 = ~\P1_EBX_reg[2]/NET0131  & ~n15364 ;
  assign n24995 = ~n15365 & ~n24994 ;
  assign n24996 = n2262 & n24995 ;
  assign n24997 = ~n24992 & ~n24996 ;
  assign n24998 = ~n24993 & n24997 ;
  assign n24999 = n2432 & ~n24998 ;
  assign n25000 = \P1_EBX_reg[2]/NET0131  & ~n15402 ;
  assign n25001 = ~n24999 & ~n25000 ;
  assign n25004 = ~\P2_EBX_reg[28]/NET0131  & ~n15048 ;
  assign n25005 = n1766 & ~n15060 ;
  assign n25006 = ~n25004 & n25005 ;
  assign n25002 = n1722 & n23372 ;
  assign n25003 = \P2_EBX_reg[28]/NET0131  & ~n15019 ;
  assign n25007 = ~n25002 & ~n25003 ;
  assign n25008 = ~n25006 & n25007 ;
  assign n25009 = n1927 & ~n25008 ;
  assign n25010 = \P2_EBX_reg[28]/NET0131  & ~n12632 ;
  assign n25011 = ~n25009 & ~n25010 ;
  assign n25013 = \P2_EBX_reg[2]/NET0131  & ~n15019 ;
  assign n25012 = n1722 & n17793 ;
  assign n25014 = ~\P2_EBX_reg[2]/NET0131  & ~n15022 ;
  assign n25015 = ~n15023 & ~n25014 ;
  assign n25016 = n1766 & n25015 ;
  assign n25017 = ~n25012 & ~n25016 ;
  assign n25018 = ~n25013 & n25017 ;
  assign n25019 = n1927 & ~n25018 ;
  assign n25020 = \P2_EBX_reg[2]/NET0131  & ~n12632 ;
  assign n25021 = ~n25019 & ~n25020 ;
  assign n25023 = \P2_EBX_reg[3]/NET0131  & ~n15019 ;
  assign n25022 = n1722 & n17804 ;
  assign n25024 = ~\P2_EBX_reg[3]/NET0131  & ~n15023 ;
  assign n25025 = ~n15024 & ~n25024 ;
  assign n25026 = n1766 & n25025 ;
  assign n25027 = ~n25022 & ~n25026 ;
  assign n25028 = ~n25023 & n25027 ;
  assign n25029 = n1927 & ~n25028 ;
  assign n25030 = \P2_EBX_reg[3]/NET0131  & ~n12632 ;
  assign n25031 = ~n25029 & ~n25030 ;
  assign n25033 = \P2_EBX_reg[4]/NET0131  & ~n15019 ;
  assign n25032 = n1722 & n17815 ;
  assign n25034 = ~\P2_EBX_reg[4]/NET0131  & ~n15024 ;
  assign n25035 = ~n15025 & ~n25034 ;
  assign n25036 = n1766 & n25035 ;
  assign n25037 = ~n25032 & ~n25036 ;
  assign n25038 = ~n25033 & n25037 ;
  assign n25039 = n1927 & ~n25038 ;
  assign n25040 = \P2_EBX_reg[4]/NET0131  & ~n12632 ;
  assign n25041 = ~n25039 & ~n25040 ;
  assign n25043 = \P2_EBX_reg[5]/NET0131  & ~n15019 ;
  assign n25042 = n1722 & n17869 ;
  assign n25044 = ~\P2_EBX_reg[5]/NET0131  & ~n15025 ;
  assign n25045 = ~n15026 & ~n25044 ;
  assign n25046 = n1766 & n25045 ;
  assign n25047 = ~n25042 & ~n25046 ;
  assign n25048 = ~n25043 & n25047 ;
  assign n25049 = n1927 & ~n25048 ;
  assign n25050 = \P2_EBX_reg[5]/NET0131  & ~n12632 ;
  assign n25051 = ~n25049 & ~n25050 ;
  assign n25053 = \P1_EBX_reg[3]/NET0131  & ~n15073 ;
  assign n25052 = n2242 & n17027 ;
  assign n25054 = ~\P1_EBX_reg[3]/NET0131  & ~n15365 ;
  assign n25055 = ~n15366 & ~n25054 ;
  assign n25056 = n2262 & n25055 ;
  assign n25057 = ~n25052 & ~n25056 ;
  assign n25058 = ~n25053 & n25057 ;
  assign n25059 = n2432 & ~n25058 ;
  assign n25060 = \P1_EBX_reg[3]/NET0131  & ~n15402 ;
  assign n25061 = ~n25059 & ~n25060 ;
  assign n25063 = \P2_EBX_reg[6]/NET0131  & ~n15019 ;
  assign n25062 = n1722 & n17880 ;
  assign n25064 = ~\P2_EBX_reg[6]/NET0131  & ~n15026 ;
  assign n25065 = ~n15027 & ~n25064 ;
  assign n25066 = n1766 & n25065 ;
  assign n25067 = ~n25062 & ~n25066 ;
  assign n25068 = ~n25063 & n25067 ;
  assign n25069 = n1927 & ~n25068 ;
  assign n25070 = \P2_EBX_reg[6]/NET0131  & ~n12632 ;
  assign n25071 = ~n25069 & ~n25070 ;
  assign n25074 = \P2_EBX_reg[7]/NET0131  & ~n15019 ;
  assign n25072 = n1798 & ~n6188 ;
  assign n25073 = n1722 & n25072 ;
  assign n25075 = ~\P2_EBX_reg[7]/NET0131  & ~n15027 ;
  assign n25076 = ~n15028 & ~n25075 ;
  assign n25077 = n1766 & n25076 ;
  assign n25078 = ~n25073 & ~n25077 ;
  assign n25079 = ~n25074 & n25078 ;
  assign n25080 = n1927 & ~n25079 ;
  assign n25081 = \P2_EBX_reg[7]/NET0131  & ~n12632 ;
  assign n25082 = ~n25080 & ~n25081 ;
  assign n25084 = \P2_EBX_reg[8]/NET0131  & ~n15019 ;
  assign n25083 = n1722 & n17922 ;
  assign n25085 = ~\P2_EBX_reg[8]/NET0131  & ~n15028 ;
  assign n25086 = ~n15029 & ~n25085 ;
  assign n25087 = n1766 & n25086 ;
  assign n25088 = ~n25083 & ~n25087 ;
  assign n25089 = ~n25084 & n25088 ;
  assign n25090 = n1927 & ~n25089 ;
  assign n25091 = \P2_EBX_reg[8]/NET0131  & ~n12632 ;
  assign n25092 = ~n25090 & ~n25091 ;
  assign n25094 = \P2_EBX_reg[9]/NET0131  & ~n15019 ;
  assign n25093 = n1722 & n17968 ;
  assign n25095 = ~\P2_EBX_reg[9]/NET0131  & ~n15029 ;
  assign n25096 = ~n15030 & ~n25095 ;
  assign n25097 = n1766 & n25096 ;
  assign n25098 = ~n25093 & ~n25097 ;
  assign n25099 = ~n25094 & n25098 ;
  assign n25100 = n1927 & ~n25099 ;
  assign n25101 = \P2_EBX_reg[9]/NET0131  & ~n12632 ;
  assign n25102 = ~n25100 & ~n25101 ;
  assign n25104 = \P1_EBX_reg[4]/NET0131  & ~n15073 ;
  assign n25103 = n2242 & n17251 ;
  assign n25105 = ~\P1_EBX_reg[4]/NET0131  & ~n15366 ;
  assign n25106 = ~n15367 & ~n25105 ;
  assign n25107 = n2262 & n25106 ;
  assign n25108 = ~n25103 & ~n25107 ;
  assign n25109 = ~n25104 & n25108 ;
  assign n25110 = n2432 & ~n25109 ;
  assign n25111 = \P1_EBX_reg[4]/NET0131  & ~n15402 ;
  assign n25112 = ~n25110 & ~n25111 ;
  assign n25114 = \P1_EBX_reg[5]/NET0131  & ~n15073 ;
  assign n25113 = n2242 & n17276 ;
  assign n25115 = ~\P1_EBX_reg[5]/NET0131  & ~n15367 ;
  assign n25116 = ~n15368 & ~n25115 ;
  assign n25117 = n2262 & n25116 ;
  assign n25118 = ~n25113 & ~n25117 ;
  assign n25119 = ~n25114 & n25118 ;
  assign n25120 = n2432 & ~n25119 ;
  assign n25121 = \P1_EBX_reg[5]/NET0131  & ~n15402 ;
  assign n25122 = ~n25120 & ~n25121 ;
  assign n25124 = \P1_EBX_reg[6]/NET0131  & ~n15073 ;
  assign n25123 = n2242 & n17637 ;
  assign n25125 = ~\P1_EBX_reg[6]/NET0131  & ~n15368 ;
  assign n25126 = ~n15369 & ~n25125 ;
  assign n25127 = n2262 & n25126 ;
  assign n25128 = ~n25123 & ~n25127 ;
  assign n25129 = ~n25124 & n25128 ;
  assign n25130 = n2432 & ~n25129 ;
  assign n25131 = \P1_EBX_reg[6]/NET0131  & ~n15402 ;
  assign n25132 = ~n25130 & ~n25131 ;
  assign n25134 = \P1_EBX_reg[7]/NET0131  & ~n15073 ;
  assign n25133 = n2242 & n17307 ;
  assign n25135 = ~\P1_EBX_reg[7]/NET0131  & ~n15369 ;
  assign n25136 = ~n15370 & ~n25135 ;
  assign n25137 = n2262 & n25136 ;
  assign n25138 = ~n25133 & ~n25137 ;
  assign n25139 = ~n25134 & n25138 ;
  assign n25140 = n2432 & ~n25139 ;
  assign n25141 = \P1_EBX_reg[7]/NET0131  & ~n15402 ;
  assign n25142 = ~n25140 & ~n25141 ;
  assign n25144 = \P1_EBX_reg[8]/NET0131  & ~n15073 ;
  assign n25143 = n2242 & n17495 ;
  assign n25145 = ~\P1_EBX_reg[8]/NET0131  & ~n15370 ;
  assign n25146 = ~n15371 & ~n25145 ;
  assign n25147 = n2262 & n25146 ;
  assign n25148 = ~n25143 & ~n25147 ;
  assign n25149 = ~n25144 & n25148 ;
  assign n25150 = n2432 & ~n25149 ;
  assign n25151 = \P1_EBX_reg[8]/NET0131  & ~n15402 ;
  assign n25152 = ~n25150 & ~n25151 ;
  assign n25154 = \P1_EBX_reg[9]/NET0131  & ~n15073 ;
  assign n25153 = n2242 & n17679 ;
  assign n25155 = ~\P1_EBX_reg[9]/NET0131  & ~n15371 ;
  assign n25156 = ~n15372 & ~n25155 ;
  assign n25157 = n2262 & n25156 ;
  assign n25158 = ~n25153 & ~n25157 ;
  assign n25159 = ~n25154 & n25158 ;
  assign n25160 = n2432 & ~n25159 ;
  assign n25161 = \P1_EBX_reg[9]/NET0131  & ~n15402 ;
  assign n25162 = ~n25160 & ~n25161 ;
  assign n25163 = \P3_uWord_reg[3]/NET0131  & ~n16086 ;
  assign n25164 = \buf2_reg[3]/NET0131  & n2862 ;
  assign n25165 = \P3_uWord_reg[3]/NET0131  & n2835 ;
  assign n25166 = ~n25164 & ~n25165 ;
  assign n25167 = n2821 & ~n25166 ;
  assign n25168 = \P3_uWord_reg[3]/NET0131  & ~n2908 ;
  assign n25169 = ~n24307 & ~n25168 ;
  assign n25170 = ~n25167 & n25169 ;
  assign n25171 = n2453 & ~n25170 ;
  assign n25172 = ~n25163 & ~n25171 ;
  assign n25173 = \P3_uWord_reg[7]/NET0131  & ~n16090 ;
  assign n25174 = n2821 & n22933 ;
  assign n25175 = ~n24316 & ~n25174 ;
  assign n25176 = n2453 & ~n25175 ;
  assign n25177 = ~n25173 & ~n25176 ;
  assign n25178 = n2453 & n2910 ;
  assign n25179 = n16086 & ~n25178 ;
  assign n25180 = \P3_CodeFetch_reg/NET0131  & ~n25179 ;
  assign n25181 = ~n2963 & ~n25180 ;
  assign n25182 = n15942 & ~n20146 ;
  assign n25183 = \P2_CodeFetch_reg/NET0131  & ~n25182 ;
  assign n25184 = ~n1934 & ~n25183 ;
  assign n25186 = \datao[30]_pad  & ~n2833 ;
  assign n25187 = \P3_EAX_reg[29]/NET0131  & n16120 ;
  assign n25189 = \P3_EAX_reg[30]/NET0131  & n25187 ;
  assign n25188 = ~\P3_EAX_reg[30]/NET0131  & ~n25187 ;
  assign n25190 = n16094 & ~n25188 ;
  assign n25191 = ~n25189 & n25190 ;
  assign n25192 = ~n2786 & n25191 ;
  assign n25193 = ~n25186 & ~n25192 ;
  assign n25194 = n2453 & ~n25193 ;
  assign n25185 = \P3_uWord_reg[14]/NET0131  & n16888 ;
  assign n25195 = \datao[30]_pad  & ~n16899 ;
  assign n25196 = ~n25185 & ~n25195 ;
  assign n25197 = ~n25194 & n25196 ;
  assign n25199 = \P2_Datao_reg[30]/NET0131  & ~n16941 ;
  assign n25200 = \P2_EAX_reg[29]/NET0131  & n15973 ;
  assign n25201 = ~\P2_EAX_reg[30]/NET0131  & ~n25200 ;
  assign n25202 = \P2_EAX_reg[30]/NET0131  & n25200 ;
  assign n25203 = ~n25201 & ~n25202 ;
  assign n25204 = n1922 & n25203 ;
  assign n25205 = ~n25199 & ~n25204 ;
  assign n25206 = n1927 & ~n25205 ;
  assign n25198 = \P2_uWord_reg[14]/NET0131  & n16919 ;
  assign n25207 = \P2_Datao_reg[30]/NET0131  & ~n16936 ;
  assign n25208 = ~n25198 & ~n25207 ;
  assign n25209 = ~n25206 & n25208 ;
  assign n25211 = ~n2311 & n2432 ;
  assign n25212 = \P1_EAX_reg[29]/NET0131  & n16025 ;
  assign n25214 = \P1_EAX_reg[30]/NET0131  & n25212 ;
  assign n25213 = ~\P1_EAX_reg[30]/NET0131  & ~n25212 ;
  assign n25215 = n15990 & ~n25213 ;
  assign n25216 = ~n25214 & n25215 ;
  assign n25217 = n25211 & n25216 ;
  assign n25210 = \P1_uWord_reg[14]/NET0131  & n2440 ;
  assign n25218 = ~n2313 & n2432 ;
  assign n25219 = n16884 & ~n25218 ;
  assign n25220 = \P1_Datao_reg[30]/NET0131  & ~n25219 ;
  assign n25221 = ~n25210 & ~n25220 ;
  assign n25222 = ~n25217 & n25221 ;
  assign n25225 = \P1_CodeFetch_reg/NET0131  & n2432 ;
  assign n25226 = ~n18554 & n25225 ;
  assign n25223 = ~n3026 & n5097 ;
  assign n25224 = \P1_CodeFetch_reg/NET0131  & ~n25223 ;
  assign n25227 = ~n2446 & ~n25224 ;
  assign n25228 = ~n25226 & n25227 ;
  assign n25229 = \P1_uWord_reg[0]/NET0131  & ~n15988 ;
  assign n25233 = \P1_uWord_reg[0]/NET0131  & n2317 ;
  assign n25234 = ~n23386 & ~n25233 ;
  assign n25235 = n2222 & ~n25234 ;
  assign n25230 = ~\P1_EAX_reg[16]/NET0131  & ~n16015 ;
  assign n25231 = ~n16016 & ~n25230 ;
  assign n25232 = n15990 & n25231 ;
  assign n25236 = \P1_uWord_reg[0]/NET0131  & n15991 ;
  assign n25237 = ~n25232 & ~n25236 ;
  assign n25238 = ~n25235 & n25237 ;
  assign n25239 = n2432 & ~n25238 ;
  assign n25240 = ~n25229 & ~n25239 ;
  assign n25241 = \P2_uWord_reg[0]/NET0131  & ~n15942 ;
  assign n25242 = \P2_uWord_reg[0]/NET0131  & n1805 ;
  assign n25243 = ~n17444 & ~n25242 ;
  assign n25244 = n1742 & ~n25243 ;
  assign n25245 = \P2_uWord_reg[0]/NET0131  & n15981 ;
  assign n25246 = ~\P2_EAX_reg[16]/NET0131  & ~n15964 ;
  assign n25247 = ~n15965 & ~n25246 ;
  assign n25248 = n15980 & n25247 ;
  assign n25249 = ~n25245 & ~n25248 ;
  assign n25250 = ~n25244 & n25249 ;
  assign n25251 = n1927 & ~n25250 ;
  assign n25252 = ~n25241 & ~n25251 ;
  assign n25253 = \P2_uWord_reg[10]/NET0131  & ~n16950 ;
  assign n25254 = n1742 & n16073 ;
  assign n25255 = ~\P2_EAX_reg[26]/NET0131  & ~n15971 ;
  assign n25256 = n1743 & ~n22327 ;
  assign n25257 = ~n25255 & n25256 ;
  assign n25258 = ~n25254 & ~n25257 ;
  assign n25259 = n16959 & ~n25258 ;
  assign n25260 = ~n25253 & ~n25259 ;
  assign n25261 = \P1_uWord_reg[10]/NET0131  & ~n15994 ;
  assign n25262 = ~n5161 & n15996 ;
  assign n25263 = ~\P1_EAX_reg[26]/NET0131  & ~n22315 ;
  assign n25264 = n2225 & ~n22316 ;
  assign n25265 = ~n25263 & n25264 ;
  assign n25266 = ~n25262 & ~n25265 ;
  assign n25267 = n16029 & ~n25266 ;
  assign n25268 = ~n25261 & ~n25267 ;
  assign n25269 = \P2_uWord_reg[14]/NET0131  & ~n15942 ;
  assign n25271 = n15980 & n25203 ;
  assign n25270 = \P2_uWord_reg[14]/NET0131  & ~n15982 ;
  assign n25272 = ~n15011 & ~n25270 ;
  assign n25273 = ~n25271 & n25272 ;
  assign n25274 = n1927 & ~n25273 ;
  assign n25275 = ~n25269 & ~n25274 ;
  assign n25276 = \P2_uWord_reg[1]/NET0131  & ~n15942 ;
  assign n25277 = \P2_uWord_reg[1]/NET0131  & n1805 ;
  assign n25278 = ~n17778 & ~n25277 ;
  assign n25279 = n1742 & ~n25278 ;
  assign n25280 = \P2_uWord_reg[1]/NET0131  & n15981 ;
  assign n25281 = ~\P2_EAX_reg[17]/NET0131  & ~n15965 ;
  assign n25282 = ~n15966 & ~n25281 ;
  assign n25283 = n15980 & n25282 ;
  assign n25284 = ~n25280 & ~n25283 ;
  assign n25285 = ~n25279 & n25284 ;
  assign n25286 = n1927 & ~n25285 ;
  assign n25287 = ~n25276 & ~n25286 ;
  assign n25288 = \P2_uWord_reg[2]/NET0131  & ~n15942 ;
  assign n25289 = \P2_uWord_reg[2]/NET0131  & n1805 ;
  assign n25290 = ~n22459 & ~n25289 ;
  assign n25291 = n1742 & ~n25290 ;
  assign n25292 = \P2_uWord_reg[2]/NET0131  & n15981 ;
  assign n25293 = ~\P2_EAX_reg[18]/NET0131  & ~n15966 ;
  assign n25294 = ~n15967 & ~n25293 ;
  assign n25295 = n15980 & n25294 ;
  assign n25296 = ~n25292 & ~n25295 ;
  assign n25297 = ~n25291 & n25296 ;
  assign n25298 = n1927 & ~n25297 ;
  assign n25299 = ~n25288 & ~n25298 ;
  assign n25300 = \P1_uWord_reg[13]/NET0131  & ~n15988 ;
  assign n25301 = ~\P1_EAX_reg[29]/NET0131  & ~n16025 ;
  assign n25302 = ~n25212 & ~n25301 ;
  assign n25303 = n15990 & n25302 ;
  assign n25304 = \P1_uWord_reg[13]/NET0131  & ~n15992 ;
  assign n25305 = ~n16318 & ~n25304 ;
  assign n25306 = ~n25303 & n25305 ;
  assign n25307 = n2432 & ~n25306 ;
  assign n25308 = ~n25300 & ~n25307 ;
  assign n25309 = \P2_uWord_reg[5]/NET0131  & ~n15942 ;
  assign n25310 = \P2_uWord_reg[5]/NET0131  & n1805 ;
  assign n25311 = ~n22491 & ~n25310 ;
  assign n25312 = n1742 & ~n25311 ;
  assign n25313 = \P2_uWord_reg[5]/NET0131  & n15981 ;
  assign n25315 = \P2_EAX_reg[21]/NET0131  & n15969 ;
  assign n25314 = ~\P2_EAX_reg[21]/NET0131  & ~n15969 ;
  assign n25316 = n15980 & ~n25314 ;
  assign n25317 = ~n25315 & n25316 ;
  assign n25318 = ~n25313 & ~n25317 ;
  assign n25319 = ~n25312 & n25318 ;
  assign n25320 = n1927 & ~n25319 ;
  assign n25321 = ~n25309 & ~n25320 ;
  assign n25322 = \P1_uWord_reg[14]/NET0131  & ~n15988 ;
  assign n25323 = \P1_uWord_reg[14]/NET0131  & ~n15992 ;
  assign n25324 = ~n5191 & n15932 ;
  assign n25325 = ~n25323 & ~n25324 ;
  assign n25326 = ~n25216 & n25325 ;
  assign n25327 = n2432 & ~n25326 ;
  assign n25328 = ~n25322 & ~n25327 ;
  assign n25329 = \P2_uWord_reg[6]/NET0131  & ~n16950 ;
  assign n25330 = ~\P2_EAX_reg[22]/NET0131  & ~n25315 ;
  assign n25331 = ~n15970 & ~n25330 ;
  assign n25332 = n1743 & n25331 ;
  assign n25333 = n1742 & n22504 ;
  assign n25334 = ~n25332 & ~n25333 ;
  assign n25335 = n16959 & ~n25334 ;
  assign n25336 = ~n25329 & ~n25335 ;
  assign n25337 = \P1_uWord_reg[1]/NET0131  & ~n15994 ;
  assign n25338 = ~\P1_EAX_reg[17]/NET0131  & ~n16016 ;
  assign n25339 = ~n16017 & ~n25338 ;
  assign n25340 = n15990 & n25339 ;
  assign n25341 = n2377 & n23513 ;
  assign n25342 = ~n25340 & ~n25341 ;
  assign n25343 = n2432 & ~n25342 ;
  assign n25344 = ~n25337 & ~n25343 ;
  assign n25345 = \P1_uWord_reg[2]/NET0131  & ~n15988 ;
  assign n25347 = \P1_uWord_reg[2]/NET0131  & n2317 ;
  assign n25348 = ~n16970 & ~n25347 ;
  assign n25349 = n2222 & ~n25348 ;
  assign n25346 = \P1_uWord_reg[2]/NET0131  & n15991 ;
  assign n25350 = ~\P1_EAX_reg[18]/NET0131  & ~n16017 ;
  assign n25351 = ~n16018 & ~n25350 ;
  assign n25352 = n15990 & n25351 ;
  assign n25353 = ~n25346 & ~n25352 ;
  assign n25354 = ~n25349 & n25353 ;
  assign n25355 = n2432 & ~n25354 ;
  assign n25356 = ~n25345 & ~n25355 ;
  assign n25357 = \P2_uWord_reg[9]/NET0131  & ~n15942 ;
  assign n25360 = ~\P2_EAX_reg[25]/NET0131  & ~n16925 ;
  assign n25361 = ~n15971 & n15980 ;
  assign n25362 = ~n25360 & n25361 ;
  assign n25358 = \P2_uWord_reg[9]/NET0131  & ~n15982 ;
  assign n25359 = n1742 & n17935 ;
  assign n25363 = ~n25358 & ~n25359 ;
  assign n25364 = ~n25362 & n25363 ;
  assign n25365 = n1927 & ~n25364 ;
  assign n25366 = ~n25357 & ~n25365 ;
  assign n25367 = \P1_uWord_reg[5]/NET0131  & ~n15994 ;
  assign n25368 = ~\P1_EAX_reg[21]/NET0131  & ~n21701 ;
  assign n25369 = n15990 & ~n16020 ;
  assign n25370 = ~n25368 & n25369 ;
  assign n25371 = n2377 & n23673 ;
  assign n25372 = ~n25370 & ~n25371 ;
  assign n25373 = n2432 & ~n25372 ;
  assign n25374 = ~n25367 & ~n25373 ;
  assign n25375 = \P1_uWord_reg[6]/NET0131  & ~n15994 ;
  assign n25376 = n2377 & n23753 ;
  assign n25377 = ~\P1_EAX_reg[22]/NET0131  & ~n16020 ;
  assign n25378 = n15990 & ~n16021 ;
  assign n25379 = ~n25377 & n25378 ;
  assign n25380 = ~n25376 & ~n25379 ;
  assign n25381 = n2432 & ~n25380 ;
  assign n25382 = ~n25375 & ~n25381 ;
  assign n25383 = \P1_uWord_reg[9]/NET0131  & ~n15994 ;
  assign n25384 = ~\P1_EAX_reg[25]/NET0131  & ~n16022 ;
  assign n25385 = n2225 & ~n22315 ;
  assign n25386 = ~n25384 & n25385 ;
  assign n25387 = ~n5158 & n15996 ;
  assign n25388 = ~n25386 & ~n25387 ;
  assign n25389 = n16029 & ~n25388 ;
  assign n25390 = ~n25383 & ~n25389 ;
  assign n25391 = \P3_uWord_reg[0]/NET0131  & ~n16086 ;
  assign n25392 = \P3_uWord_reg[0]/NET0131  & n2835 ;
  assign n25393 = ~n22627 & ~n25392 ;
  assign n25394 = n2821 & ~n25393 ;
  assign n25395 = \P3_uWord_reg[0]/NET0131  & ~n2908 ;
  assign n25396 = \P3_EAX_reg[16]/NET0131  & n16110 ;
  assign n25397 = ~\P3_EAX_reg[16]/NET0131  & ~n16110 ;
  assign n25398 = ~n25396 & ~n25397 ;
  assign n25399 = n16094 & n25398 ;
  assign n25400 = ~n25395 & ~n25399 ;
  assign n25401 = ~n25394 & n25400 ;
  assign n25402 = n2453 & ~n25401 ;
  assign n25403 = ~n25391 & ~n25402 ;
  assign n25404 = \P3_uWord_reg[10]/NET0131  & ~n16090 ;
  assign n25405 = ~n2835 & n16042 ;
  assign n25406 = ~\P3_EAX_reg[26]/NET0131  & ~n16118 ;
  assign n25407 = n2818 & ~n22303 ;
  assign n25408 = ~n25406 & n25407 ;
  assign n25409 = ~n25405 & ~n25408 ;
  assign n25410 = n18178 & ~n25409 ;
  assign n25411 = ~n25404 & ~n25410 ;
  assign n25412 = \P3_uWord_reg[13]/NET0131  & ~n16086 ;
  assign n25413 = ~\P3_EAX_reg[29]/NET0131  & ~n16120 ;
  assign n25414 = n16094 & ~n25187 ;
  assign n25415 = ~n25413 & n25414 ;
  assign n25416 = \P3_uWord_reg[13]/NET0131  & ~n16088 ;
  assign n25417 = \buf2_reg[13]/NET0131  & n2862 ;
  assign n25418 = n2821 & n25417 ;
  assign n25419 = ~n25416 & ~n25418 ;
  assign n25420 = ~n25415 & n25419 ;
  assign n25421 = n2453 & ~n25420 ;
  assign n25422 = ~n25412 & ~n25421 ;
  assign n25423 = \P3_uWord_reg[14]/NET0131  & ~n16086 ;
  assign n25424 = \P3_uWord_reg[14]/NET0131  & ~n16088 ;
  assign n25425 = n2862 & n14944 ;
  assign n25426 = ~n25424 & ~n25425 ;
  assign n25427 = ~n25191 & n25426 ;
  assign n25428 = n2453 & ~n25427 ;
  assign n25429 = ~n25423 & ~n25428 ;
  assign n25430 = \P3_uWord_reg[1]/NET0131  & ~n16086 ;
  assign n25431 = \P3_uWord_reg[1]/NET0131  & n2835 ;
  assign n25432 = ~n17261 & ~n25431 ;
  assign n25433 = n2821 & ~n25432 ;
  assign n25434 = \P3_uWord_reg[1]/NET0131  & ~n2908 ;
  assign n25435 = ~\P3_EAX_reg[17]/NET0131  & ~n25396 ;
  assign n25436 = ~n16111 & ~n25435 ;
  assign n25437 = n16094 & n25436 ;
  assign n25438 = ~n25434 & ~n25437 ;
  assign n25439 = ~n25433 & n25438 ;
  assign n25440 = n2453 & ~n25439 ;
  assign n25441 = ~n25430 & ~n25440 ;
  assign n25442 = \P3_uWord_reg[2]/NET0131  & ~n16086 ;
  assign n25443 = \P3_uWord_reg[2]/NET0131  & n2835 ;
  assign n25444 = ~n22685 & ~n25443 ;
  assign n25445 = n2821 & ~n25444 ;
  assign n25446 = \P3_uWord_reg[2]/NET0131  & ~n2908 ;
  assign n25447 = ~\P3_EAX_reg[18]/NET0131  & ~n16111 ;
  assign n25448 = ~n16112 & ~n25447 ;
  assign n25449 = n16094 & n25448 ;
  assign n25450 = ~n25446 & ~n25449 ;
  assign n25451 = ~n25445 & n25450 ;
  assign n25452 = n2453 & ~n25451 ;
  assign n25453 = ~n25442 & ~n25452 ;
  assign n25454 = \P3_uWord_reg[5]/NET0131  & ~n16086 ;
  assign n25455 = \buf2_reg[5]/NET0131  & n2862 ;
  assign n25456 = \P3_uWord_reg[5]/NET0131  & n2835 ;
  assign n25457 = ~n25455 & ~n25456 ;
  assign n25458 = n2821 & ~n25457 ;
  assign n25459 = \P3_uWord_reg[5]/NET0131  & ~n2908 ;
  assign n25460 = ~\P3_EAX_reg[21]/NET0131  & ~n16114 ;
  assign n25461 = ~n16115 & ~n25460 ;
  assign n25462 = n16094 & n25461 ;
  assign n25463 = ~n25459 & ~n25462 ;
  assign n25464 = ~n25458 & n25463 ;
  assign n25465 = n2453 & ~n25464 ;
  assign n25466 = ~n25454 & ~n25465 ;
  assign n25467 = \P3_uWord_reg[6]/NET0131  & ~n16086 ;
  assign n25468 = \P3_uWord_reg[6]/NET0131  & n2835 ;
  assign n25469 = ~n22915 & ~n25468 ;
  assign n25470 = n2821 & ~n25469 ;
  assign n25471 = \P3_uWord_reg[6]/NET0131  & ~n2908 ;
  assign n25472 = ~\P3_EAX_reg[22]/NET0131  & ~n16115 ;
  assign n25473 = ~n24313 & ~n25472 ;
  assign n25474 = n16094 & n25473 ;
  assign n25475 = ~n25471 & ~n25474 ;
  assign n25476 = ~n25470 & n25475 ;
  assign n25477 = n2453 & ~n25476 ;
  assign n25478 = ~n25467 & ~n25477 ;
  assign n25479 = \P3_uWord_reg[9]/NET0131  & ~n16090 ;
  assign n25480 = ~\P3_EAX_reg[25]/NET0131  & ~n16117 ;
  assign n25481 = n16094 & ~n16118 ;
  assign n25482 = ~n25480 & n25481 ;
  assign n25483 = \buf2_reg[9]/NET0131  & n2862 ;
  assign n25484 = n2821 & n25483 ;
  assign n25485 = ~n25482 & ~n25484 ;
  assign n25486 = n2453 & ~n25485 ;
  assign n25487 = ~n25479 & ~n25486 ;
  assign n25489 = \P1_lWord_reg[0]/NET0131  & n2317 ;
  assign n25490 = ~n23386 & ~n25489 ;
  assign n25491 = n2222 & ~n25490 ;
  assign n25488 = \P1_lWord_reg[0]/NET0131  & n15991 ;
  assign n25492 = \P1_EAX_reg[0]/NET0131  & n15990 ;
  assign n25493 = ~n25488 & ~n25492 ;
  assign n25494 = ~n25491 & n25493 ;
  assign n25495 = n2432 & ~n25494 ;
  assign n25496 = \P1_lWord_reg[0]/NET0131  & ~n15988 ;
  assign n25497 = ~n25495 & ~n25496 ;
  assign n25499 = \P1_lWord_reg[10]/NET0131  & n2317 ;
  assign n25500 = ~n17825 & ~n25499 ;
  assign n25501 = n2222 & ~n25500 ;
  assign n25498 = \P1_lWord_reg[10]/NET0131  & n15991 ;
  assign n25502 = \P1_EAX_reg[10]/NET0131  & n15990 ;
  assign n25503 = ~n25498 & ~n25502 ;
  assign n25504 = ~n25501 & n25503 ;
  assign n25505 = n2432 & ~n25504 ;
  assign n25506 = \P1_lWord_reg[10]/NET0131  & ~n15988 ;
  assign n25507 = ~n25505 & ~n25506 ;
  assign n25509 = \P1_lWord_reg[11]/NET0131  & n2317 ;
  assign n25510 = ~n17978 & ~n25509 ;
  assign n25511 = n2222 & ~n25510 ;
  assign n25508 = \P1_lWord_reg[11]/NET0131  & n15991 ;
  assign n25512 = \P1_EAX_reg[11]/NET0131  & n15990 ;
  assign n25513 = ~n25508 & ~n25512 ;
  assign n25514 = ~n25511 & n25513 ;
  assign n25515 = n2432 & ~n25514 ;
  assign n25516 = \P1_lWord_reg[11]/NET0131  & ~n15988 ;
  assign n25517 = ~n25515 & ~n25516 ;
  assign n25519 = \P1_lWord_reg[12]/NET0131  & n2317 ;
  assign n25520 = ~n18169 & ~n25519 ;
  assign n25521 = n2222 & ~n25520 ;
  assign n25518 = \P1_lWord_reg[12]/NET0131  & n15991 ;
  assign n25522 = \P1_EAX_reg[12]/NET0131  & n15990 ;
  assign n25523 = ~n25518 & ~n25522 ;
  assign n25524 = ~n25521 & n25523 ;
  assign n25525 = n2432 & ~n25524 ;
  assign n25526 = \P1_lWord_reg[12]/NET0131  & ~n15988 ;
  assign n25527 = ~n25525 & ~n25526 ;
  assign n25528 = \P1_lWord_reg[13]/NET0131  & ~n15994 ;
  assign n25529 = \P1_EAX_reg[13]/NET0131  & n15990 ;
  assign n25530 = ~n16318 & ~n25529 ;
  assign n25531 = n2432 & ~n25530 ;
  assign n25532 = ~n25528 & ~n25531 ;
  assign n25533 = \P1_lWord_reg[14]/NET0131  & ~n15994 ;
  assign n25534 = \P1_EAX_reg[14]/NET0131  & n15990 ;
  assign n25535 = ~n25324 & ~n25534 ;
  assign n25536 = n2432 & ~n25535 ;
  assign n25537 = ~n25533 & ~n25536 ;
  assign n25538 = \P1_lWord_reg[15]/NET0131  & ~n15994 ;
  assign n25539 = \P1_EAX_reg[15]/NET0131  & n2225 ;
  assign n25540 = ~n5194 & n15996 ;
  assign n25541 = ~n25539 & ~n25540 ;
  assign n25542 = n16029 & ~n25541 ;
  assign n25543 = ~n25538 & ~n25542 ;
  assign n25544 = \P1_lWord_reg[1]/NET0131  & ~n15994 ;
  assign n25545 = \P1_EAX_reg[1]/NET0131  & n15990 ;
  assign n25546 = ~n25341 & ~n25545 ;
  assign n25547 = n2432 & ~n25546 ;
  assign n25548 = ~n25544 & ~n25547 ;
  assign n25549 = \P1_lWord_reg[3]/NET0131  & ~n15994 ;
  assign n25550 = \P1_EAX_reg[3]/NET0131  & n15990 ;
  assign n25551 = n2377 & n23564 ;
  assign n25552 = ~n25550 & ~n25551 ;
  assign n25553 = n2432 & ~n25552 ;
  assign n25554 = ~n25549 & ~n25553 ;
  assign n25555 = \P1_lWord_reg[2]/NET0131  & ~n15994 ;
  assign n25556 = \P1_EAX_reg[2]/NET0131  & n15990 ;
  assign n25557 = n2377 & n23608 ;
  assign n25558 = ~n25556 & ~n25557 ;
  assign n25559 = n2432 & ~n25558 ;
  assign n25560 = ~n25555 & ~n25559 ;
  assign n25561 = \P1_lWord_reg[4]/NET0131  & ~n15994 ;
  assign n25562 = \P1_EAX_reg[4]/NET0131  & n15990 ;
  assign n25563 = ~n21765 & ~n25562 ;
  assign n25564 = n2432 & ~n25563 ;
  assign n25565 = ~n25561 & ~n25564 ;
  assign n25566 = \P1_lWord_reg[5]/NET0131  & ~n15994 ;
  assign n25567 = \P1_EAX_reg[5]/NET0131  & n15990 ;
  assign n25568 = ~n25371 & ~n25567 ;
  assign n25569 = n2432 & ~n25568 ;
  assign n25570 = ~n25566 & ~n25569 ;
  assign n25571 = \P1_lWord_reg[6]/NET0131  & ~n15994 ;
  assign n25572 = \P1_EAX_reg[6]/NET0131  & n15990 ;
  assign n25573 = ~n25376 & ~n25572 ;
  assign n25574 = n2432 & ~n25573 ;
  assign n25575 = ~n25571 & ~n25574 ;
  assign n25576 = \P1_lWord_reg[7]/NET0131  & ~n15994 ;
  assign n25577 = \P1_EAX_reg[7]/NET0131  & n15990 ;
  assign n25578 = ~n22350 & ~n25577 ;
  assign n25579 = n2432 & ~n25578 ;
  assign n25580 = ~n25576 & ~n25579 ;
  assign n25581 = \P1_EAX_reg[8]/NET0131  & n2225 ;
  assign n25582 = ~n16963 & ~n25581 ;
  assign n25583 = ~n2301 & ~n25582 ;
  assign n25584 = \P1_lWord_reg[8]/NET0131  & ~n15992 ;
  assign n25585 = ~n25583 & ~n25584 ;
  assign n25586 = n2432 & ~n25585 ;
  assign n25587 = \P1_lWord_reg[8]/NET0131  & ~n15988 ;
  assign n25588 = ~n25586 & ~n25587 ;
  assign n25589 = \P1_lWord_reg[9]/NET0131  & ~n15994 ;
  assign n25590 = \P1_EAX_reg[9]/NET0131  & n2225 ;
  assign n25591 = ~n25387 & ~n25590 ;
  assign n25592 = n16029 & ~n25591 ;
  assign n25593 = ~n25589 & ~n25592 ;
  assign n25597 = ~\P3_EAX_reg[12]/NET0131  & n2833 ;
  assign n25596 = ~\datao[12]_pad  & ~n2833 ;
  assign n25598 = n2453 & ~n25596 ;
  assign n25599 = ~n25597 & n25598 ;
  assign n25594 = \P3_lWord_reg[12]/NET0131  & n16888 ;
  assign n25595 = \datao[12]_pad  & ~n16899 ;
  assign n25600 = ~n25594 & ~n25595 ;
  assign n25601 = ~n25599 & n25600 ;
  assign n25605 = ~\P3_EAX_reg[13]/NET0131  & n2833 ;
  assign n25604 = ~\datao[13]_pad  & ~n2833 ;
  assign n25606 = n2453 & ~n25604 ;
  assign n25607 = ~n25605 & n25606 ;
  assign n25602 = \P3_lWord_reg[13]/NET0131  & n16888 ;
  assign n25603 = \datao[13]_pad  & ~n16899 ;
  assign n25608 = ~n25602 & ~n25603 ;
  assign n25609 = ~n25607 & n25608 ;
  assign n25613 = ~\P3_EAX_reg[14]/NET0131  & n2833 ;
  assign n25612 = ~\datao[14]_pad  & ~n2833 ;
  assign n25614 = n2453 & ~n25612 ;
  assign n25615 = ~n25613 & n25614 ;
  assign n25610 = \P3_lWord_reg[14]/NET0131  & n16888 ;
  assign n25611 = \datao[14]_pad  & ~n16899 ;
  assign n25616 = ~n25610 & ~n25611 ;
  assign n25617 = ~n25615 & n25616 ;
  assign n25621 = ~\P3_EAX_reg[2]/NET0131  & n2833 ;
  assign n25620 = ~\datao[2]_pad  & ~n2833 ;
  assign n25622 = n2453 & ~n25620 ;
  assign n25623 = ~n25621 & n25622 ;
  assign n25618 = \P3_lWord_reg[2]/NET0131  & n16888 ;
  assign n25619 = \datao[2]_pad  & ~n16899 ;
  assign n25624 = ~n25618 & ~n25619 ;
  assign n25625 = ~n25623 & n25624 ;
  assign n25629 = ~\P3_EAX_reg[3]/NET0131  & n2833 ;
  assign n25628 = ~\datao[3]_pad  & ~n2833 ;
  assign n25630 = n2453 & ~n25628 ;
  assign n25631 = ~n25629 & n25630 ;
  assign n25626 = \P3_lWord_reg[3]/NET0131  & n16888 ;
  assign n25627 = \datao[3]_pad  & ~n16899 ;
  assign n25632 = ~n25626 & ~n25627 ;
  assign n25633 = ~n25631 & n25632 ;
  assign n25637 = ~\P2_EAX_reg[0]/NET0131  & n16941 ;
  assign n25636 = ~\P2_Datao_reg[0]/NET0131  & ~n16941 ;
  assign n25638 = n1927 & ~n25636 ;
  assign n25639 = ~n25637 & n25638 ;
  assign n25634 = \P2_lWord_reg[0]/NET0131  & n16919 ;
  assign n25635 = \P2_Datao_reg[0]/NET0131  & ~n16936 ;
  assign n25640 = ~n25634 & ~n25635 ;
  assign n25641 = ~n25639 & n25640 ;
  assign n25645 = ~\P2_EAX_reg[10]/NET0131  & n16941 ;
  assign n25644 = ~\P2_Datao_reg[10]/NET0131  & ~n16941 ;
  assign n25646 = n1927 & ~n25644 ;
  assign n25647 = ~n25645 & n25646 ;
  assign n25642 = \P2_lWord_reg[10]/NET0131  & n16919 ;
  assign n25643 = \P2_Datao_reg[10]/NET0131  & ~n16936 ;
  assign n25648 = ~n25642 & ~n25643 ;
  assign n25649 = ~n25647 & n25648 ;
  assign n25653 = ~\P2_EAX_reg[11]/NET0131  & n16941 ;
  assign n25652 = ~\P2_Datao_reg[11]/NET0131  & ~n16941 ;
  assign n25654 = n1927 & ~n25652 ;
  assign n25655 = ~n25653 & n25654 ;
  assign n25650 = \P2_lWord_reg[11]/NET0131  & n16919 ;
  assign n25651 = \P2_Datao_reg[11]/NET0131  & ~n16936 ;
  assign n25656 = ~n25650 & ~n25651 ;
  assign n25657 = ~n25655 & n25656 ;
  assign n25661 = ~\P2_EAX_reg[12]/NET0131  & n16941 ;
  assign n25660 = ~\P2_Datao_reg[12]/NET0131  & ~n16941 ;
  assign n25662 = n1927 & ~n25660 ;
  assign n25663 = ~n25661 & n25662 ;
  assign n25658 = \P2_lWord_reg[12]/NET0131  & n16919 ;
  assign n25659 = \P2_Datao_reg[12]/NET0131  & ~n16936 ;
  assign n25664 = ~n25658 & ~n25659 ;
  assign n25665 = ~n25663 & n25664 ;
  assign n25669 = ~\P1_EAX_reg[2]/NET0131  & n2313 ;
  assign n25668 = ~\P1_Datao_reg[2]/NET0131  & ~n2313 ;
  assign n25670 = n2432 & ~n25668 ;
  assign n25671 = ~n25669 & n25670 ;
  assign n25666 = \P1_lWord_reg[2]/NET0131  & n2440 ;
  assign n25667 = \P1_Datao_reg[2]/NET0131  & ~n16884 ;
  assign n25672 = ~n25666 & ~n25667 ;
  assign n25673 = ~n25671 & n25672 ;
  assign n25677 = ~\P2_EAX_reg[5]/NET0131  & n16941 ;
  assign n25676 = ~\P2_Datao_reg[5]/NET0131  & ~n16941 ;
  assign n25678 = n1927 & ~n25676 ;
  assign n25679 = ~n25677 & n25678 ;
  assign n25674 = \P2_lWord_reg[5]/NET0131  & n16919 ;
  assign n25675 = \P2_Datao_reg[5]/NET0131  & ~n16936 ;
  assign n25680 = ~n25674 & ~n25675 ;
  assign n25681 = ~n25679 & n25680 ;
  assign n25685 = ~\P2_EAX_reg[7]/NET0131  & n16941 ;
  assign n25684 = ~\P2_Datao_reg[7]/NET0131  & ~n16941 ;
  assign n25686 = n1927 & ~n25684 ;
  assign n25687 = ~n25685 & n25686 ;
  assign n25682 = \P2_lWord_reg[7]/NET0131  & n16919 ;
  assign n25683 = \P2_Datao_reg[7]/NET0131  & ~n16936 ;
  assign n25688 = ~n25682 & ~n25683 ;
  assign n25689 = ~n25687 & n25688 ;
  assign n25693 = ~\P2_EAX_reg[8]/NET0131  & n16941 ;
  assign n25692 = ~\P2_Datao_reg[8]/NET0131  & ~n16941 ;
  assign n25694 = n1927 & ~n25692 ;
  assign n25695 = ~n25693 & n25694 ;
  assign n25690 = \P2_lWord_reg[8]/NET0131  & n16919 ;
  assign n25691 = \P2_Datao_reg[8]/NET0131  & ~n16936 ;
  assign n25696 = ~n25690 & ~n25691 ;
  assign n25697 = ~n25695 & n25696 ;
  assign n25701 = ~\P1_EAX_reg[4]/NET0131  & n2313 ;
  assign n25700 = ~\P1_Datao_reg[4]/NET0131  & ~n2313 ;
  assign n25702 = n2432 & ~n25700 ;
  assign n25703 = ~n25701 & n25702 ;
  assign n25698 = \P1_lWord_reg[4]/NET0131  & n2440 ;
  assign n25699 = \P1_Datao_reg[4]/NET0131  & ~n16884 ;
  assign n25704 = ~n25698 & ~n25699 ;
  assign n25705 = ~n25703 & n25704 ;
  assign n25709 = ~\P1_EAX_reg[6]/NET0131  & n2313 ;
  assign n25708 = ~\P1_Datao_reg[6]/NET0131  & ~n2313 ;
  assign n25710 = n2432 & ~n25708 ;
  assign n25711 = ~n25709 & n25710 ;
  assign n25706 = \P1_lWord_reg[6]/NET0131  & n2440 ;
  assign n25707 = \P1_Datao_reg[6]/NET0131  & ~n16884 ;
  assign n25712 = ~n25706 & ~n25707 ;
  assign n25713 = ~n25711 & n25712 ;
  assign n25717 = ~\P1_EAX_reg[8]/NET0131  & n2313 ;
  assign n25716 = ~\P1_Datao_reg[8]/NET0131  & ~n2313 ;
  assign n25718 = n2432 & ~n25716 ;
  assign n25719 = ~n25717 & n25718 ;
  assign n25714 = \P1_lWord_reg[8]/NET0131  & n2440 ;
  assign n25715 = \P1_Datao_reg[8]/NET0131  & ~n16884 ;
  assign n25720 = ~n25714 & ~n25715 ;
  assign n25721 = ~n25719 & n25720 ;
  assign n25725 = ~\P1_EAX_reg[14]/NET0131  & n2313 ;
  assign n25724 = ~\P1_Datao_reg[14]/NET0131  & ~n2313 ;
  assign n25726 = n2432 & ~n25724 ;
  assign n25727 = ~n25725 & n25726 ;
  assign n25722 = \P1_lWord_reg[14]/NET0131  & n2440 ;
  assign n25723 = \P1_Datao_reg[14]/NET0131  & ~n16884 ;
  assign n25728 = ~n25722 & ~n25723 ;
  assign n25729 = ~n25727 & n25728 ;
  assign n25733 = ~\P1_EAX_reg[15]/NET0131  & n2313 ;
  assign n25732 = ~\P1_Datao_reg[15]/NET0131  & ~n2313 ;
  assign n25734 = n2432 & ~n25732 ;
  assign n25735 = ~n25733 & n25734 ;
  assign n25730 = \P1_lWord_reg[15]/NET0131  & n2440 ;
  assign n25731 = \P1_Datao_reg[15]/NET0131  & ~n16884 ;
  assign n25736 = ~n25730 & ~n25731 ;
  assign n25737 = ~n25735 & n25736 ;
  assign n25739 = \P1_Datao_reg[18]/NET0131  & n2306 ;
  assign n25740 = ~\P1_Datao_reg[18]/NET0131  & ~n2312 ;
  assign n25741 = n2312 & ~n25351 ;
  assign n25742 = ~n25740 & ~n25741 ;
  assign n25743 = n21698 & n25742 ;
  assign n25744 = ~n25739 & ~n25743 ;
  assign n25745 = n2432 & ~n25744 ;
  assign n25738 = \P1_uWord_reg[2]/NET0131  & n2440 ;
  assign n25746 = \P1_Datao_reg[18]/NET0131  & ~n16884 ;
  assign n25747 = ~n25738 & ~n25746 ;
  assign n25748 = ~n25745 & n25747 ;
  assign n25750 = \P1_Datao_reg[17]/NET0131  & ~n2313 ;
  assign n25751 = ~n2311 & n25340 ;
  assign n25752 = ~n25750 & ~n25751 ;
  assign n25753 = n2432 & ~n25752 ;
  assign n25749 = \P1_uWord_reg[1]/NET0131  & n2440 ;
  assign n25754 = \P1_Datao_reg[17]/NET0131  & ~n16884 ;
  assign n25755 = ~n25749 & ~n25754 ;
  assign n25756 = ~n25753 & n25755 ;
  assign n25758 = \P1_Datao_reg[21]/NET0131  & ~n2313 ;
  assign n25759 = ~n2311 & n25370 ;
  assign n25760 = ~n25758 & ~n25759 ;
  assign n25761 = n2432 & ~n25760 ;
  assign n25757 = \P1_uWord_reg[5]/NET0131  & n2440 ;
  assign n25762 = \P1_Datao_reg[21]/NET0131  & ~n16884 ;
  assign n25763 = ~n25757 & ~n25762 ;
  assign n25764 = ~n25761 & n25763 ;
  assign n25766 = \P1_Datao_reg[22]/NET0131  & ~n25219 ;
  assign n25765 = \P1_uWord_reg[6]/NET0131  & n2440 ;
  assign n25767 = n25211 & n25379 ;
  assign n25768 = ~n25765 & ~n25767 ;
  assign n25769 = ~n25766 & n25768 ;
  assign n25771 = \datao[16]_pad  & ~n2833 ;
  assign n25772 = ~n2786 & n25399 ;
  assign n25773 = ~n25771 & ~n25772 ;
  assign n25774 = n2453 & ~n25773 ;
  assign n25770 = \P3_uWord_reg[0]/NET0131  & n16888 ;
  assign n25775 = \datao[16]_pad  & ~n16899 ;
  assign n25776 = ~n25770 & ~n25775 ;
  assign n25777 = ~n25774 & n25776 ;
  assign n25779 = \datao[17]_pad  & ~n24302 ;
  assign n25778 = \P3_uWord_reg[1]/NET0131  & n16888 ;
  assign n25780 = n24304 & n25437 ;
  assign n25781 = ~n25778 & ~n25780 ;
  assign n25782 = ~n25779 & n25781 ;
  assign n25784 = \datao[18]_pad  & ~n2833 ;
  assign n25785 = ~n2786 & n25449 ;
  assign n25786 = ~n25784 & ~n25785 ;
  assign n25787 = n2453 & ~n25786 ;
  assign n25783 = \P3_uWord_reg[2]/NET0131  & n16888 ;
  assign n25788 = \datao[18]_pad  & ~n16899 ;
  assign n25789 = ~n25783 & ~n25788 ;
  assign n25790 = ~n25787 & n25789 ;
  assign n25792 = \P1_Datao_reg[25]/NET0131  & ~n2313 ;
  assign n25793 = n2312 & n25386 ;
  assign n25794 = ~n25792 & ~n25793 ;
  assign n25795 = n2432 & ~n25794 ;
  assign n25791 = \P1_uWord_reg[9]/NET0131  & n2440 ;
  assign n25796 = \P1_Datao_reg[25]/NET0131  & ~n16884 ;
  assign n25797 = ~n25791 & ~n25796 ;
  assign n25798 = ~n25795 & n25797 ;
  assign n25800 = \datao[21]_pad  & ~n2833 ;
  assign n25801 = ~n2786 & n25462 ;
  assign n25802 = ~n25800 & ~n25801 ;
  assign n25803 = n2453 & ~n25802 ;
  assign n25799 = \P3_uWord_reg[5]/NET0131  & n16888 ;
  assign n25804 = \datao[21]_pad  & ~n16899 ;
  assign n25805 = ~n25799 & ~n25804 ;
  assign n25806 = ~n25803 & n25805 ;
  assign n25808 = \P1_Datao_reg[26]/NET0131  & ~n2313 ;
  assign n25809 = n2312 & n25265 ;
  assign n25810 = ~n25808 & ~n25809 ;
  assign n25811 = n2432 & ~n25810 ;
  assign n25807 = \P1_uWord_reg[10]/NET0131  & n2440 ;
  assign n25812 = \P1_Datao_reg[26]/NET0131  & ~n16884 ;
  assign n25813 = ~n25807 & ~n25812 ;
  assign n25814 = ~n25811 & n25813 ;
  assign n25816 = \datao[22]_pad  & ~n2833 ;
  assign n25817 = ~n2786 & n25474 ;
  assign n25818 = ~n25816 & ~n25817 ;
  assign n25819 = n2453 & ~n25818 ;
  assign n25815 = \P3_uWord_reg[6]/NET0131  & n16888 ;
  assign n25820 = \datao[22]_pad  & ~n16899 ;
  assign n25821 = ~n25815 & ~n25820 ;
  assign n25822 = ~n25819 & n25821 ;
  assign n25824 = \datao[25]_pad  & ~n2833 ;
  assign n25825 = ~n2786 & n25482 ;
  assign n25826 = ~n25824 & ~n25825 ;
  assign n25827 = n2453 & ~n25826 ;
  assign n25823 = \P3_uWord_reg[9]/NET0131  & n16888 ;
  assign n25828 = \datao[25]_pad  & ~n16899 ;
  assign n25829 = ~n25823 & ~n25828 ;
  assign n25830 = ~n25827 & n25829 ;
  assign n25833 = ~n2815 & n24304 ;
  assign n25834 = n25408 & n25833 ;
  assign n25831 = \P3_uWord_reg[10]/NET0131  & n16888 ;
  assign n25832 = \datao[26]_pad  & ~n24302 ;
  assign n25835 = ~n25831 & ~n25832 ;
  assign n25836 = ~n25834 & n25835 ;
  assign n25838 = \datao[29]_pad  & ~n2833 ;
  assign n25839 = ~n2786 & n25415 ;
  assign n25840 = ~n25838 & ~n25839 ;
  assign n25841 = n2453 & ~n25840 ;
  assign n25837 = \P3_uWord_reg[13]/NET0131  & n16888 ;
  assign n25842 = \datao[29]_pad  & ~n16899 ;
  assign n25843 = ~n25837 & ~n25842 ;
  assign n25844 = ~n25841 & n25843 ;
  assign n25846 = \P1_Datao_reg[29]/NET0131  & ~n2313 ;
  assign n25847 = n2426 & n25302 ;
  assign n25848 = ~n25846 & ~n25847 ;
  assign n25849 = n2432 & ~n25848 ;
  assign n25845 = \P1_uWord_reg[13]/NET0131  & n2440 ;
  assign n25850 = \P1_Datao_reg[29]/NET0131  & ~n16884 ;
  assign n25851 = ~n25845 & ~n25850 ;
  assign n25852 = ~n25849 & n25851 ;
  assign n25854 = \P2_Datao_reg[16]/NET0131  & ~n16941 ;
  assign n25855 = ~n1819 & n25248 ;
  assign n25856 = ~n25854 & ~n25855 ;
  assign n25857 = n1927 & ~n25856 ;
  assign n25853 = \P2_uWord_reg[0]/NET0131  & n16919 ;
  assign n25858 = \P2_Datao_reg[16]/NET0131  & ~n16936 ;
  assign n25859 = ~n25853 & ~n25858 ;
  assign n25860 = ~n25857 & n25859 ;
  assign n25862 = ~n1819 & n25283 ;
  assign n25863 = \P2_Datao_reg[17]/NET0131  & ~n16941 ;
  assign n25864 = ~n25862 & ~n25863 ;
  assign n25865 = n1927 & ~n25864 ;
  assign n25861 = \P2_uWord_reg[1]/NET0131  & n16919 ;
  assign n25866 = \P2_Datao_reg[17]/NET0131  & ~n16936 ;
  assign n25867 = ~n25861 & ~n25866 ;
  assign n25868 = ~n25865 & n25867 ;
  assign n25870 = \P2_Datao_reg[18]/NET0131  & ~n16941 ;
  assign n25871 = ~n1819 & n25295 ;
  assign n25872 = ~n25870 & ~n25871 ;
  assign n25873 = n1927 & ~n25872 ;
  assign n25869 = \P2_uWord_reg[2]/NET0131  & n16919 ;
  assign n25874 = \P2_Datao_reg[18]/NET0131  & ~n16936 ;
  assign n25875 = ~n25869 & ~n25874 ;
  assign n25876 = ~n25873 & n25875 ;
  assign n25878 = \P2_Datao_reg[21]/NET0131  & ~n16941 ;
  assign n25879 = ~n1819 & n25317 ;
  assign n25880 = ~n25878 & ~n25879 ;
  assign n25881 = n1927 & ~n25880 ;
  assign n25877 = \P2_uWord_reg[5]/NET0131  & n16919 ;
  assign n25882 = \P2_Datao_reg[21]/NET0131  & ~n16936 ;
  assign n25883 = ~n25877 & ~n25882 ;
  assign n25884 = ~n25881 & n25883 ;
  assign n25886 = ~n1819 & ~n25331 ;
  assign n25887 = ~\P2_Datao_reg[22]/NET0131  & n1819 ;
  assign n25888 = n15980 & ~n25887 ;
  assign n25889 = ~n25886 & n25888 ;
  assign n25890 = \P2_Datao_reg[22]/NET0131  & ~n16922 ;
  assign n25891 = ~n25889 & ~n25890 ;
  assign n25892 = n1927 & ~n25891 ;
  assign n25885 = \P2_uWord_reg[6]/NET0131  & n16919 ;
  assign n25893 = \P2_Datao_reg[22]/NET0131  & ~n16936 ;
  assign n25894 = ~n25885 & ~n25893 ;
  assign n25895 = ~n25892 & n25894 ;
  assign n25897 = \P2_Datao_reg[25]/NET0131  & ~n16941 ;
  assign n25898 = ~n1819 & n25362 ;
  assign n25899 = ~n25897 & ~n25898 ;
  assign n25900 = n1927 & ~n25899 ;
  assign n25896 = \P2_uWord_reg[9]/NET0131  & n16919 ;
  assign n25901 = \P2_Datao_reg[25]/NET0131  & ~n16936 ;
  assign n25902 = ~n25896 & ~n25901 ;
  assign n25903 = ~n25900 & n25902 ;
  assign n25905 = n1927 & ~n16941 ;
  assign n25906 = n16936 & ~n25905 ;
  assign n25907 = \P2_Datao_reg[26]/NET0131  & ~n25906 ;
  assign n25904 = \P2_uWord_reg[10]/NET0131  & n16919 ;
  assign n25908 = ~n1819 & n16959 ;
  assign n25909 = n25257 & n25908 ;
  assign n25910 = ~n25904 & ~n25909 ;
  assign n25911 = ~n25907 & n25910 ;
  assign n25913 = \P2_Datao_reg[29]/NET0131  & ~n16941 ;
  assign n25914 = ~\P2_EAX_reg[29]/NET0131  & ~n15973 ;
  assign n25915 = n15980 & ~n25200 ;
  assign n25916 = ~n25914 & n25915 ;
  assign n25917 = ~n1819 & n25916 ;
  assign n25918 = ~n25913 & ~n25917 ;
  assign n25919 = n1927 & ~n25918 ;
  assign n25912 = \P2_uWord_reg[13]/NET0131  & n16919 ;
  assign n25920 = \P2_Datao_reg[29]/NET0131  & ~n16936 ;
  assign n25921 = ~n25912 & ~n25920 ;
  assign n25922 = ~n25919 & n25921 ;
  assign n25924 = \P1_Datao_reg[16]/NET0131  & ~n2313 ;
  assign n25925 = ~n2311 & n25232 ;
  assign n25926 = ~n25924 & ~n25925 ;
  assign n25927 = n2432 & ~n25926 ;
  assign n25923 = \P1_uWord_reg[0]/NET0131  & n2440 ;
  assign n25928 = \P1_Datao_reg[16]/NET0131  & ~n16884 ;
  assign n25929 = ~n25923 & ~n25928 ;
  assign n25930 = ~n25927 & n25929 ;
  assign n25932 = \P3_lWord_reg[0]/NET0131  & n2835 ;
  assign n25933 = ~n22627 & ~n25932 ;
  assign n25934 = n2821 & ~n25933 ;
  assign n25931 = \P3_EAX_reg[0]/NET0131  & n16094 ;
  assign n25935 = \P3_lWord_reg[0]/NET0131  & ~n2908 ;
  assign n25936 = ~n25931 & ~n25935 ;
  assign n25937 = ~n25934 & n25936 ;
  assign n25938 = n2453 & ~n25937 ;
  assign n25939 = \P3_lWord_reg[0]/NET0131  & ~n16086 ;
  assign n25940 = ~n25938 & ~n25939 ;
  assign n25941 = \P3_lWord_reg[10]/NET0131  & ~n16090 ;
  assign n25942 = \P3_EAX_reg[10]/NET0131  & n16094 ;
  assign n25943 = n2862 & n16042 ;
  assign n25944 = ~n25942 & ~n25943 ;
  assign n25945 = n2453 & ~n25944 ;
  assign n25946 = ~n25941 & ~n25945 ;
  assign n25948 = \P3_lWord_reg[11]/NET0131  & n2835 ;
  assign n25949 = ~n14048 & ~n25948 ;
  assign n25950 = n2821 & ~n25949 ;
  assign n25947 = \P3_EAX_reg[11]/NET0131  & n16094 ;
  assign n25951 = \P3_lWord_reg[11]/NET0131  & ~n2908 ;
  assign n25952 = ~n25947 & ~n25951 ;
  assign n25953 = ~n25950 & n25952 ;
  assign n25954 = n2453 & ~n25953 ;
  assign n25955 = \P3_lWord_reg[11]/NET0131  & ~n16086 ;
  assign n25956 = ~n25954 & ~n25955 ;
  assign n25957 = \P3_lWord_reg[12]/NET0131  & ~n16090 ;
  assign n25958 = \P3_EAX_reg[12]/NET0131  & n16094 ;
  assign n25959 = ~n16093 & ~n25958 ;
  assign n25960 = n2453 & ~n25959 ;
  assign n25961 = ~n25957 & ~n25960 ;
  assign n25963 = \P3_lWord_reg[13]/NET0131  & n2835 ;
  assign n25964 = ~n25417 & ~n25963 ;
  assign n25965 = n2821 & ~n25964 ;
  assign n25962 = \P3_EAX_reg[13]/NET0131  & n16094 ;
  assign n25966 = \P3_lWord_reg[13]/NET0131  & ~n2908 ;
  assign n25967 = ~n25962 & ~n25966 ;
  assign n25968 = ~n25965 & n25967 ;
  assign n25969 = n2453 & ~n25968 ;
  assign n25970 = \P3_lWord_reg[13]/NET0131  & ~n16086 ;
  assign n25971 = ~n25969 & ~n25970 ;
  assign n25972 = \P3_lWord_reg[14]/NET0131  & ~n16090 ;
  assign n25973 = \P3_EAX_reg[14]/NET0131  & n16094 ;
  assign n25974 = ~n25425 & ~n25973 ;
  assign n25975 = n2453 & ~n25974 ;
  assign n25976 = ~n25972 & ~n25975 ;
  assign n25978 = \P3_lWord_reg[15]/NET0131  & n2835 ;
  assign n25979 = ~n17208 & ~n25978 ;
  assign n25980 = n2821 & ~n25979 ;
  assign n25977 = \P3_EAX_reg[15]/NET0131  & n16094 ;
  assign n25981 = \P3_lWord_reg[15]/NET0131  & ~n2908 ;
  assign n25982 = ~n25977 & ~n25981 ;
  assign n25983 = ~n25980 & n25982 ;
  assign n25984 = n2453 & ~n25983 ;
  assign n25985 = \P3_lWord_reg[15]/NET0131  & ~n16086 ;
  assign n25986 = ~n25984 & ~n25985 ;
  assign n25988 = \P3_lWord_reg[1]/NET0131  & n2835 ;
  assign n25989 = ~n17261 & ~n25988 ;
  assign n25990 = n2821 & ~n25989 ;
  assign n25987 = \P3_EAX_reg[1]/NET0131  & n16094 ;
  assign n25991 = \P3_lWord_reg[1]/NET0131  & ~n2908 ;
  assign n25992 = ~n25987 & ~n25991 ;
  assign n25993 = ~n25990 & n25992 ;
  assign n25994 = n2453 & ~n25993 ;
  assign n25995 = \P3_lWord_reg[1]/NET0131  & ~n16086 ;
  assign n25996 = ~n25994 & ~n25995 ;
  assign n25998 = \P3_lWord_reg[2]/NET0131  & n2835 ;
  assign n25999 = ~n22685 & ~n25998 ;
  assign n26000 = n2821 & ~n25999 ;
  assign n25997 = \P3_EAX_reg[2]/NET0131  & n16094 ;
  assign n26001 = \P3_lWord_reg[2]/NET0131  & ~n2908 ;
  assign n26002 = ~n25997 & ~n26001 ;
  assign n26003 = ~n26000 & n26002 ;
  assign n26004 = n2453 & ~n26003 ;
  assign n26005 = \P3_lWord_reg[2]/NET0131  & ~n16086 ;
  assign n26006 = ~n26004 & ~n26005 ;
  assign n26008 = \P3_lWord_reg[3]/NET0131  & n2835 ;
  assign n26009 = ~n25164 & ~n26008 ;
  assign n26010 = n2821 & ~n26009 ;
  assign n26007 = \P3_EAX_reg[3]/NET0131  & n16094 ;
  assign n26011 = \P3_lWord_reg[3]/NET0131  & ~n2908 ;
  assign n26012 = ~n26007 & ~n26011 ;
  assign n26013 = ~n26010 & n26012 ;
  assign n26014 = n2453 & ~n26013 ;
  assign n26015 = \P3_lWord_reg[3]/NET0131  & ~n16086 ;
  assign n26016 = ~n26014 & ~n26015 ;
  assign n26018 = \P3_lWord_reg[4]/NET0131  & n2835 ;
  assign n26019 = ~n21812 & ~n26018 ;
  assign n26020 = n2821 & ~n26019 ;
  assign n26017 = \P3_EAX_reg[4]/NET0131  & n16094 ;
  assign n26021 = \P3_lWord_reg[4]/NET0131  & ~n2908 ;
  assign n26022 = ~n26017 & ~n26021 ;
  assign n26023 = ~n26020 & n26022 ;
  assign n26024 = n2453 & ~n26023 ;
  assign n26025 = \P3_lWord_reg[4]/NET0131  & ~n16086 ;
  assign n26026 = ~n26024 & ~n26025 ;
  assign n26028 = \P3_lWord_reg[5]/NET0131  & n2835 ;
  assign n26029 = ~n25455 & ~n26028 ;
  assign n26030 = n2821 & ~n26029 ;
  assign n26027 = \P3_EAX_reg[5]/NET0131  & n16094 ;
  assign n26031 = \P3_lWord_reg[5]/NET0131  & ~n2908 ;
  assign n26032 = ~n26027 & ~n26031 ;
  assign n26033 = ~n26030 & n26032 ;
  assign n26034 = n2453 & ~n26033 ;
  assign n26035 = \P3_lWord_reg[5]/NET0131  & ~n16086 ;
  assign n26036 = ~n26034 & ~n26035 ;
  assign n26038 = \P3_lWord_reg[6]/NET0131  & n2835 ;
  assign n26039 = ~n22915 & ~n26038 ;
  assign n26040 = n2821 & ~n26039 ;
  assign n26037 = \P3_EAX_reg[6]/NET0131  & n16094 ;
  assign n26041 = \P3_lWord_reg[6]/NET0131  & ~n2908 ;
  assign n26042 = ~n26037 & ~n26041 ;
  assign n26043 = ~n26040 & n26042 ;
  assign n26044 = n2453 & ~n26043 ;
  assign n26045 = \P3_lWord_reg[6]/NET0131  & ~n16086 ;
  assign n26046 = ~n26044 & ~n26045 ;
  assign n26048 = \P3_lWord_reg[7]/NET0131  & n2835 ;
  assign n26049 = ~n22933 & ~n26048 ;
  assign n26050 = n2821 & ~n26049 ;
  assign n26047 = \P3_EAX_reg[7]/NET0131  & n16094 ;
  assign n26051 = \P3_lWord_reg[7]/NET0131  & ~n2908 ;
  assign n26052 = ~n26047 & ~n26051 ;
  assign n26053 = ~n26050 & n26052 ;
  assign n26054 = n2453 & ~n26053 ;
  assign n26055 = \P3_lWord_reg[7]/NET0131  & ~n16086 ;
  assign n26056 = ~n26054 & ~n26055 ;
  assign n26058 = \P3_lWord_reg[8]/NET0131  & n2835 ;
  assign n26059 = ~n22956 & ~n26058 ;
  assign n26060 = n2821 & ~n26059 ;
  assign n26057 = \P3_lWord_reg[8]/NET0131  & ~n2908 ;
  assign n26061 = \P3_EAX_reg[8]/NET0131  & n16094 ;
  assign n26062 = ~n26057 & ~n26061 ;
  assign n26063 = ~n26060 & n26062 ;
  assign n26064 = n2453 & ~n26063 ;
  assign n26065 = \P3_lWord_reg[8]/NET0131  & ~n16086 ;
  assign n26066 = ~n26064 & ~n26065 ;
  assign n26068 = \P3_lWord_reg[9]/NET0131  & n2835 ;
  assign n26069 = ~n25483 & ~n26068 ;
  assign n26070 = n2821 & ~n26069 ;
  assign n26067 = \P3_EAX_reg[9]/NET0131  & n16094 ;
  assign n26071 = \P3_lWord_reg[9]/NET0131  & ~n2908 ;
  assign n26072 = ~n26067 & ~n26071 ;
  assign n26073 = ~n26070 & n26072 ;
  assign n26074 = n2453 & ~n26073 ;
  assign n26075 = \P3_lWord_reg[9]/NET0131  & ~n16086 ;
  assign n26076 = ~n26074 & ~n26075 ;
  assign n26079 = n2635 & n18209 ;
  assign n26078 = ~\P3_InstQueue_reg[0][2]/NET0131  & ~n18209 ;
  assign n26080 = n2994 & ~n26078 ;
  assign n26081 = ~n26079 & n26080 ;
  assign n26077 = \P3_InstQueue_reg[0][2]/NET0131  & ~n18218 ;
  assign n26082 = \buf2_reg[26]/NET0131  & n18200 ;
  assign n26083 = \buf2_reg[18]/NET0131  & n18203 ;
  assign n26084 = ~n26082 & ~n26083 ;
  assign n26085 = n2970 & ~n26084 ;
  assign n26086 = \buf2_reg[2]/NET0131  & n18228 ;
  assign n26087 = ~n26085 & ~n26086 ;
  assign n26088 = ~n26077 & n26087 ;
  assign n26089 = ~n26081 & n26088 ;
  assign n26092 = n2635 & n18246 ;
  assign n26091 = ~\P3_InstQueue_reg[10][2]/NET0131  & ~n18246 ;
  assign n26093 = n2994 & ~n26091 ;
  assign n26094 = ~n26092 & n26093 ;
  assign n26090 = \P3_InstQueue_reg[10][2]/NET0131  & ~n18243 ;
  assign n26095 = \buf2_reg[26]/NET0131  & n18233 ;
  assign n26096 = \buf2_reg[18]/NET0131  & n18236 ;
  assign n26097 = ~n26095 & ~n26096 ;
  assign n26098 = n2970 & ~n26097 ;
  assign n26099 = \buf2_reg[2]/NET0131  & n18255 ;
  assign n26100 = ~n26098 & ~n26099 ;
  assign n26101 = ~n26090 & n26100 ;
  assign n26102 = ~n26094 & n26101 ;
  assign n26104 = n2635 & n18266 ;
  assign n26103 = ~\P3_InstQueue_reg[11][2]/NET0131  & ~n18266 ;
  assign n26105 = n2994 & ~n26103 ;
  assign n26106 = ~n26104 & n26105 ;
  assign n26112 = \P3_InstQueue_reg[11][2]/NET0131  & ~n18264 ;
  assign n26107 = ~\P3_InstQueueWr_Addr_reg[0]/NET0131  & ~\buf2_reg[26]/NET0131  ;
  assign n26108 = \P3_InstQueueWr_Addr_reg[0]/NET0131  & ~\buf2_reg[18]/NET0131  ;
  assign n26109 = ~n26107 & ~n26108 ;
  assign n26110 = n2959 & n26109 ;
  assign n26111 = n18260 & n26110 ;
  assign n26113 = \buf2_reg[2]/NET0131  & n18245 ;
  assign n26114 = n18262 & n26113 ;
  assign n26115 = ~n26111 & ~n26114 ;
  assign n26116 = ~n26112 & n26115 ;
  assign n26117 = ~n26106 & n26116 ;
  assign n26120 = n2635 & n18284 ;
  assign n26119 = ~\P3_InstQueue_reg[12][2]/NET0131  & ~n18284 ;
  assign n26121 = n2994 & ~n26119 ;
  assign n26122 = ~n26120 & n26121 ;
  assign n26118 = \P3_InstQueue_reg[12][2]/NET0131  & ~n18287 ;
  assign n26123 = \buf2_reg[18]/NET0131  & n18246 ;
  assign n26124 = \buf2_reg[26]/NET0131  & n18271 ;
  assign n26125 = ~n26123 & ~n26124 ;
  assign n26126 = n2970 & ~n26125 ;
  assign n26127 = \buf2_reg[2]/NET0131  & n18297 ;
  assign n26128 = ~n26126 & ~n26127 ;
  assign n26129 = ~n26118 & n26128 ;
  assign n26130 = ~n26122 & n26129 ;
  assign n26138 = n2635 & n18200 ;
  assign n26137 = ~\P3_InstQueue_reg[13][2]/NET0131  & ~n18200 ;
  assign n26139 = n2994 & ~n26137 ;
  assign n26140 = ~n26138 & n26139 ;
  assign n26134 = ~\P3_InstQueue_reg[13][2]/NET0131  & n18302 ;
  assign n26133 = ~\buf2_reg[2]/NET0131  & ~n18302 ;
  assign n26135 = n18305 & ~n26133 ;
  assign n26136 = ~n26134 & n26135 ;
  assign n26131 = \P3_InstQueue_reg[13][2]/NET0131  & ~n18217 ;
  assign n26132 = n18303 & n26110 ;
  assign n26141 = ~n26131 & ~n26132 ;
  assign n26142 = ~n26136 & n26141 ;
  assign n26143 = ~n26140 & n26142 ;
  assign n26146 = n2635 & n18203 ;
  assign n26145 = ~\P3_InstQueue_reg[14][2]/NET0131  & ~n18203 ;
  assign n26147 = n2994 & ~n26145 ;
  assign n26148 = ~n26146 & n26147 ;
  assign n26144 = \P3_InstQueue_reg[14][2]/NET0131  & ~n18325 ;
  assign n26149 = \buf2_reg[26]/NET0131  & n18266 ;
  assign n26150 = \buf2_reg[18]/NET0131  & n18284 ;
  assign n26151 = ~n26149 & ~n26150 ;
  assign n26152 = n2970 & ~n26151 ;
  assign n26153 = \buf2_reg[2]/NET0131  & n18335 ;
  assign n26154 = ~n26152 & ~n26153 ;
  assign n26155 = ~n26144 & n26154 ;
  assign n26156 = ~n26148 & n26155 ;
  assign n26159 = n2635 & n18212 ;
  assign n26158 = ~\P3_InstQueue_reg[15][2]/NET0131  & ~n18212 ;
  assign n26160 = n2994 & ~n26158 ;
  assign n26161 = ~n26159 & n26160 ;
  assign n26157 = \P3_InstQueue_reg[15][2]/NET0131  & ~n18344 ;
  assign n26162 = \buf2_reg[26]/NET0131  & n18284 ;
  assign n26163 = \buf2_reg[18]/NET0131  & n18200 ;
  assign n26164 = ~n26162 & ~n26163 ;
  assign n26165 = n2970 & ~n26164 ;
  assign n26166 = \buf2_reg[2]/NET0131  & n18354 ;
  assign n26167 = ~n26165 & ~n26166 ;
  assign n26168 = ~n26157 & n26167 ;
  assign n26169 = ~n26161 & n26168 ;
  assign n26172 = n2635 & n18361 ;
  assign n26171 = ~\P3_InstQueue_reg[1][2]/NET0131  & ~n18361 ;
  assign n26173 = n2994 & ~n26171 ;
  assign n26174 = ~n26172 & n26173 ;
  assign n26170 = \P3_InstQueue_reg[1][2]/NET0131  & ~n18364 ;
  assign n26175 = \buf2_reg[26]/NET0131  & n18203 ;
  assign n26176 = \buf2_reg[18]/NET0131  & n18212 ;
  assign n26177 = ~n26175 & ~n26176 ;
  assign n26178 = n2970 & ~n26177 ;
  assign n26179 = \buf2_reg[2]/NET0131  & n18374 ;
  assign n26180 = ~n26178 & ~n26179 ;
  assign n26181 = ~n26170 & n26180 ;
  assign n26182 = ~n26174 & n26181 ;
  assign n26185 = n2635 & n18386 ;
  assign n26184 = ~\P3_InstQueue_reg[2][2]/NET0131  & ~n18386 ;
  assign n26186 = n2994 & ~n26184 ;
  assign n26187 = ~n26185 & n26186 ;
  assign n26183 = \P3_InstQueue_reg[2][2]/NET0131  & ~n18383 ;
  assign n26188 = \buf2_reg[26]/NET0131  & n18212 ;
  assign n26189 = \buf2_reg[18]/NET0131  & n18209 ;
  assign n26190 = ~n26188 & ~n26189 ;
  assign n26191 = n2970 & ~n26190 ;
  assign n26192 = \buf2_reg[2]/NET0131  & n18395 ;
  assign n26193 = ~n26191 & ~n26192 ;
  assign n26194 = ~n26183 & n26193 ;
  assign n26195 = ~n26187 & n26194 ;
  assign n26198 = n2635 & n18405 ;
  assign n26197 = ~\P3_InstQueue_reg[3][2]/NET0131  & ~n18405 ;
  assign n26199 = n2994 & ~n26197 ;
  assign n26200 = ~n26198 & n26199 ;
  assign n26196 = \P3_InstQueue_reg[3][2]/NET0131  & ~n18403 ;
  assign n26201 = \buf2_reg[18]/NET0131  & n18361 ;
  assign n26202 = \buf2_reg[26]/NET0131  & n18209 ;
  assign n26203 = ~n26201 & ~n26202 ;
  assign n26204 = n2970 & ~n26203 ;
  assign n26205 = \buf2_reg[2]/NET0131  & n18414 ;
  assign n26206 = ~n26204 & ~n26205 ;
  assign n26207 = ~n26196 & n26206 ;
  assign n26208 = ~n26200 & n26207 ;
  assign n26211 = n2635 & n18421 ;
  assign n26210 = ~\P3_InstQueue_reg[4][2]/NET0131  & ~n18421 ;
  assign n26212 = n2994 & ~n26210 ;
  assign n26213 = ~n26211 & n26212 ;
  assign n26209 = \P3_InstQueue_reg[4][2]/NET0131  & ~n18424 ;
  assign n26214 = \buf2_reg[18]/NET0131  & n18386 ;
  assign n26215 = \buf2_reg[26]/NET0131  & n18361 ;
  assign n26216 = ~n26214 & ~n26215 ;
  assign n26217 = n2970 & ~n26216 ;
  assign n26218 = \buf2_reg[2]/NET0131  & n18434 ;
  assign n26219 = ~n26217 & ~n26218 ;
  assign n26220 = ~n26209 & n26219 ;
  assign n26221 = ~n26213 & n26220 ;
  assign n26229 = n2635 & n18439 ;
  assign n26228 = ~\P3_InstQueue_reg[5][2]/NET0131  & ~n18439 ;
  assign n26230 = n2994 & ~n26228 ;
  assign n26231 = ~n26229 & n26230 ;
  assign n26225 = ~\P3_InstQueue_reg[5][2]/NET0131  & n18440 ;
  assign n26224 = ~\buf2_reg[2]/NET0131  & ~n18440 ;
  assign n26226 = n18443 & ~n26224 ;
  assign n26227 = ~n26225 & n26226 ;
  assign n26222 = \P3_InstQueue_reg[5][2]/NET0131  & ~n18217 ;
  assign n26223 = n18441 & n26110 ;
  assign n26232 = ~n26222 & ~n26223 ;
  assign n26233 = ~n26227 & n26232 ;
  assign n26234 = ~n26231 & n26233 ;
  assign n26237 = n2635 & n18462 ;
  assign n26236 = ~\P3_InstQueue_reg[6][2]/NET0131  & ~n18462 ;
  assign n26238 = n2994 & ~n26236 ;
  assign n26239 = ~n26237 & n26238 ;
  assign n26235 = \P3_InstQueue_reg[6][2]/NET0131  & ~n18465 ;
  assign n26240 = \buf2_reg[26]/NET0131  & n18405 ;
  assign n26241 = \buf2_reg[18]/NET0131  & n18421 ;
  assign n26242 = ~n26240 & ~n26241 ;
  assign n26243 = n2970 & ~n26242 ;
  assign n26244 = \buf2_reg[2]/NET0131  & n18475 ;
  assign n26245 = ~n26243 & ~n26244 ;
  assign n26246 = ~n26235 & n26245 ;
  assign n26247 = ~n26239 & n26246 ;
  assign n26250 = n2635 & n18233 ;
  assign n26249 = ~\P3_InstQueue_reg[7][2]/NET0131  & ~n18233 ;
  assign n26251 = n2994 & ~n26249 ;
  assign n26252 = ~n26250 & n26251 ;
  assign n26248 = \P3_InstQueue_reg[7][2]/NET0131  & ~n18484 ;
  assign n26253 = \buf2_reg[26]/NET0131  & n18421 ;
  assign n26254 = \buf2_reg[18]/NET0131  & n18439 ;
  assign n26255 = ~n26253 & ~n26254 ;
  assign n26256 = n2970 & ~n26255 ;
  assign n26257 = \buf2_reg[2]/NET0131  & n18494 ;
  assign n26258 = ~n26256 & ~n26257 ;
  assign n26259 = ~n26248 & n26258 ;
  assign n26260 = ~n26252 & n26259 ;
  assign n26263 = n2635 & n18236 ;
  assign n26262 = ~\P3_InstQueue_reg[8][2]/NET0131  & ~n18236 ;
  assign n26264 = n2994 & ~n26262 ;
  assign n26265 = ~n26263 & n26264 ;
  assign n26261 = \P3_InstQueue_reg[8][2]/NET0131  & ~n18502 ;
  assign n26266 = \buf2_reg[26]/NET0131  & n18439 ;
  assign n26267 = \buf2_reg[18]/NET0131  & n18462 ;
  assign n26268 = ~n26266 & ~n26267 ;
  assign n26269 = n2970 & ~n26268 ;
  assign n26270 = \buf2_reg[2]/NET0131  & n18512 ;
  assign n26271 = ~n26269 & ~n26270 ;
  assign n26272 = ~n26261 & n26271 ;
  assign n26273 = ~n26265 & n26272 ;
  assign n26287 = n2635 & n18271 ;
  assign n26286 = ~\P3_InstQueue_reg[9][2]/NET0131  & ~n18271 ;
  assign n26288 = n2994 & ~n26286 ;
  assign n26289 = ~n26287 & n26288 ;
  assign n26278 = \buf2_reg[26]/NET0131  & n18462 ;
  assign n26279 = \buf2_reg[18]/NET0131  & n18233 ;
  assign n26280 = ~n26278 & ~n26279 ;
  assign n26281 = \P3_DataWidth_reg[1]/NET0131  & ~n26280 ;
  assign n26274 = \P3_InstQueue_reg[9][2]/NET0131  & ~n18235 ;
  assign n26275 = \buf2_reg[2]/NET0131  & n18235 ;
  assign n26276 = ~n26274 & ~n26275 ;
  assign n26282 = ~n18525 & ~n26276 ;
  assign n26283 = ~n26281 & ~n26282 ;
  assign n26284 = n2959 & ~n26283 ;
  assign n26277 = n4415 & ~n26276 ;
  assign n26285 = \P3_InstQueue_reg[9][2]/NET0131  & ~n18217 ;
  assign n26290 = ~n26277 & ~n26285 ;
  assign n26291 = ~n26284 & n26290 ;
  assign n26292 = ~n26289 & n26291 ;
  assign n26296 = ~\P1_EAX_reg[1]/NET0131  & n2313 ;
  assign n26295 = ~\P1_Datao_reg[1]/NET0131  & ~n2313 ;
  assign n26297 = n2432 & ~n26295 ;
  assign n26298 = ~n26296 & n26297 ;
  assign n26293 = \P1_lWord_reg[1]/NET0131  & n2440 ;
  assign n26294 = \P1_Datao_reg[1]/NET0131  & ~n16884 ;
  assign n26299 = ~n26293 & ~n26294 ;
  assign n26300 = ~n26298 & n26299 ;
  assign n26304 = ~\P3_EAX_reg[0]/NET0131  & n2833 ;
  assign n26303 = ~\datao[0]_pad  & ~n2833 ;
  assign n26305 = n2453 & ~n26303 ;
  assign n26306 = ~n26304 & n26305 ;
  assign n26301 = \P3_lWord_reg[0]/NET0131  & n16888 ;
  assign n26302 = \datao[0]_pad  & ~n16899 ;
  assign n26307 = ~n26301 & ~n26302 ;
  assign n26308 = ~n26306 & n26307 ;
  assign n26312 = ~\P3_EAX_reg[10]/NET0131  & n2833 ;
  assign n26311 = ~\datao[10]_pad  & ~n2833 ;
  assign n26313 = n2453 & ~n26311 ;
  assign n26314 = ~n26312 & n26313 ;
  assign n26309 = \P3_lWord_reg[10]/NET0131  & n16888 ;
  assign n26310 = \datao[10]_pad  & ~n16899 ;
  assign n26315 = ~n26309 & ~n26310 ;
  assign n26316 = ~n26314 & n26315 ;
  assign n26320 = ~\P3_EAX_reg[11]/NET0131  & n2833 ;
  assign n26319 = ~\datao[11]_pad  & ~n2833 ;
  assign n26321 = n2453 & ~n26319 ;
  assign n26322 = ~n26320 & n26321 ;
  assign n26317 = \P3_lWord_reg[11]/NET0131  & n16888 ;
  assign n26318 = \datao[11]_pad  & ~n16899 ;
  assign n26323 = ~n26317 & ~n26318 ;
  assign n26324 = ~n26322 & n26323 ;
  assign n26328 = ~\P3_EAX_reg[15]/NET0131  & n2833 ;
  assign n26327 = ~\datao[15]_pad  & ~n2833 ;
  assign n26329 = n2453 & ~n26327 ;
  assign n26330 = ~n26328 & n26329 ;
  assign n26325 = \P3_lWord_reg[15]/NET0131  & n16888 ;
  assign n26326 = \datao[15]_pad  & ~n16899 ;
  assign n26331 = ~n26325 & ~n26326 ;
  assign n26332 = ~n26330 & n26331 ;
  assign n26336 = ~\P3_EAX_reg[1]/NET0131  & n2833 ;
  assign n26335 = ~\datao[1]_pad  & ~n2833 ;
  assign n26337 = n2453 & ~n26335 ;
  assign n26338 = ~n26336 & n26337 ;
  assign n26333 = \P3_lWord_reg[1]/NET0131  & n16888 ;
  assign n26334 = \datao[1]_pad  & ~n16899 ;
  assign n26339 = ~n26333 & ~n26334 ;
  assign n26340 = ~n26338 & n26339 ;
  assign n26344 = ~\P3_EAX_reg[4]/NET0131  & n2833 ;
  assign n26343 = ~\datao[4]_pad  & ~n2833 ;
  assign n26345 = n2453 & ~n26343 ;
  assign n26346 = ~n26344 & n26345 ;
  assign n26341 = \P3_lWord_reg[4]/NET0131  & n16888 ;
  assign n26342 = \datao[4]_pad  & ~n16899 ;
  assign n26347 = ~n26341 & ~n26342 ;
  assign n26348 = ~n26346 & n26347 ;
  assign n26352 = ~\P3_EAX_reg[5]/NET0131  & n2833 ;
  assign n26351 = ~\datao[5]_pad  & ~n2833 ;
  assign n26353 = n2453 & ~n26351 ;
  assign n26354 = ~n26352 & n26353 ;
  assign n26349 = \P3_lWord_reg[5]/NET0131  & n16888 ;
  assign n26350 = \datao[5]_pad  & ~n16899 ;
  assign n26355 = ~n26349 & ~n26350 ;
  assign n26356 = ~n26354 & n26355 ;
  assign n26360 = ~\P3_EAX_reg[6]/NET0131  & n2833 ;
  assign n26359 = ~\datao[6]_pad  & ~n2833 ;
  assign n26361 = n2453 & ~n26359 ;
  assign n26362 = ~n26360 & n26361 ;
  assign n26357 = \P3_lWord_reg[6]/NET0131  & n16888 ;
  assign n26358 = \datao[6]_pad  & ~n16899 ;
  assign n26363 = ~n26357 & ~n26358 ;
  assign n26364 = ~n26362 & n26363 ;
  assign n26368 = ~\P3_EAX_reg[7]/NET0131  & n2833 ;
  assign n26367 = ~\datao[7]_pad  & ~n2833 ;
  assign n26369 = n2453 & ~n26367 ;
  assign n26370 = ~n26368 & n26369 ;
  assign n26365 = \P3_lWord_reg[7]/NET0131  & n16888 ;
  assign n26366 = \datao[7]_pad  & ~n16899 ;
  assign n26371 = ~n26365 & ~n26366 ;
  assign n26372 = ~n26370 & n26371 ;
  assign n26376 = ~\P3_EAX_reg[8]/NET0131  & n2833 ;
  assign n26375 = ~\datao[8]_pad  & ~n2833 ;
  assign n26377 = n2453 & ~n26375 ;
  assign n26378 = ~n26376 & n26377 ;
  assign n26373 = \P3_lWord_reg[8]/NET0131  & n16888 ;
  assign n26374 = \datao[8]_pad  & ~n16899 ;
  assign n26379 = ~n26373 & ~n26374 ;
  assign n26380 = ~n26378 & n26379 ;
  assign n26384 = ~\P3_EAX_reg[9]/NET0131  & n2833 ;
  assign n26383 = ~\datao[9]_pad  & ~n2833 ;
  assign n26385 = n2453 & ~n26383 ;
  assign n26386 = ~n26384 & n26385 ;
  assign n26381 = \P3_lWord_reg[9]/NET0131  & n16888 ;
  assign n26382 = \datao[9]_pad  & ~n16899 ;
  assign n26387 = ~n26381 & ~n26382 ;
  assign n26388 = ~n26386 & n26387 ;
  assign n26392 = ~\P2_EAX_reg[13]/NET0131  & n16941 ;
  assign n26391 = ~\P2_Datao_reg[13]/NET0131  & ~n16941 ;
  assign n26393 = n1927 & ~n26391 ;
  assign n26394 = ~n26392 & n26393 ;
  assign n26389 = \P2_lWord_reg[13]/NET0131  & n16919 ;
  assign n26390 = \P2_Datao_reg[13]/NET0131  & ~n16936 ;
  assign n26395 = ~n26389 & ~n26390 ;
  assign n26396 = ~n26394 & n26395 ;
  assign n26400 = ~\P2_EAX_reg[14]/NET0131  & n16941 ;
  assign n26399 = ~\P2_Datao_reg[14]/NET0131  & ~n16941 ;
  assign n26401 = n1927 & ~n26399 ;
  assign n26402 = ~n26400 & n26401 ;
  assign n26397 = \P2_lWord_reg[14]/NET0131  & n16919 ;
  assign n26398 = \P2_Datao_reg[14]/NET0131  & ~n16936 ;
  assign n26403 = ~n26397 & ~n26398 ;
  assign n26404 = ~n26402 & n26403 ;
  assign n26408 = ~\P2_EAX_reg[15]/NET0131  & n16941 ;
  assign n26407 = ~\P2_Datao_reg[15]/NET0131  & ~n16941 ;
  assign n26409 = n1927 & ~n26407 ;
  assign n26410 = ~n26408 & n26409 ;
  assign n26405 = \P2_lWord_reg[15]/NET0131  & n16919 ;
  assign n26406 = \P2_Datao_reg[15]/NET0131  & ~n16936 ;
  assign n26411 = ~n26405 & ~n26406 ;
  assign n26412 = ~n26410 & n26411 ;
  assign n26416 = ~\P2_EAX_reg[1]/NET0131  & n16941 ;
  assign n26415 = ~\P2_Datao_reg[1]/NET0131  & ~n16941 ;
  assign n26417 = n1927 & ~n26415 ;
  assign n26418 = ~n26416 & n26417 ;
  assign n26413 = \P2_lWord_reg[1]/NET0131  & n16919 ;
  assign n26414 = \P2_Datao_reg[1]/NET0131  & ~n16936 ;
  assign n26419 = ~n26413 & ~n26414 ;
  assign n26420 = ~n26418 & n26419 ;
  assign n26424 = ~\P2_EAX_reg[2]/NET0131  & n16941 ;
  assign n26423 = ~\P2_Datao_reg[2]/NET0131  & ~n16941 ;
  assign n26425 = n1927 & ~n26423 ;
  assign n26426 = ~n26424 & n26425 ;
  assign n26421 = \P2_lWord_reg[2]/NET0131  & n16919 ;
  assign n26422 = \P2_Datao_reg[2]/NET0131  & ~n16936 ;
  assign n26427 = ~n26421 & ~n26422 ;
  assign n26428 = ~n26426 & n26427 ;
  assign n26432 = ~\P2_EAX_reg[3]/NET0131  & n16941 ;
  assign n26431 = ~\P2_Datao_reg[3]/NET0131  & ~n16941 ;
  assign n26433 = n1927 & ~n26431 ;
  assign n26434 = ~n26432 & n26433 ;
  assign n26429 = \P2_lWord_reg[3]/NET0131  & n16919 ;
  assign n26430 = \P2_Datao_reg[3]/NET0131  & ~n16936 ;
  assign n26435 = ~n26429 & ~n26430 ;
  assign n26436 = ~n26434 & n26435 ;
  assign n26440 = ~\P2_EAX_reg[4]/NET0131  & n16941 ;
  assign n26439 = ~\P2_Datao_reg[4]/NET0131  & ~n16941 ;
  assign n26441 = n1927 & ~n26439 ;
  assign n26442 = ~n26440 & n26441 ;
  assign n26437 = \P2_lWord_reg[4]/NET0131  & n16919 ;
  assign n26438 = \P2_Datao_reg[4]/NET0131  & ~n16936 ;
  assign n26443 = ~n26437 & ~n26438 ;
  assign n26444 = ~n26442 & n26443 ;
  assign n26448 = ~\P2_EAX_reg[6]/NET0131  & n16941 ;
  assign n26447 = ~\P2_Datao_reg[6]/NET0131  & ~n16941 ;
  assign n26449 = n1927 & ~n26447 ;
  assign n26450 = ~n26448 & n26449 ;
  assign n26445 = \P2_lWord_reg[6]/NET0131  & n16919 ;
  assign n26446 = \P2_Datao_reg[6]/NET0131  & ~n16936 ;
  assign n26451 = ~n26445 & ~n26446 ;
  assign n26452 = ~n26450 & n26451 ;
  assign n26456 = ~\P2_EAX_reg[9]/NET0131  & n16941 ;
  assign n26455 = ~\P2_Datao_reg[9]/NET0131  & ~n16941 ;
  assign n26457 = n1927 & ~n26455 ;
  assign n26458 = ~n26456 & n26457 ;
  assign n26453 = \P2_lWord_reg[9]/NET0131  & n16919 ;
  assign n26454 = \P2_Datao_reg[9]/NET0131  & ~n16936 ;
  assign n26459 = ~n26453 & ~n26454 ;
  assign n26460 = ~n26458 & n26459 ;
  assign n26464 = ~\P1_EAX_reg[3]/NET0131  & n2313 ;
  assign n26463 = ~\P1_Datao_reg[3]/NET0131  & ~n2313 ;
  assign n26465 = n2432 & ~n26463 ;
  assign n26466 = ~n26464 & n26465 ;
  assign n26461 = \P1_lWord_reg[3]/NET0131  & n2440 ;
  assign n26462 = \P1_Datao_reg[3]/NET0131  & ~n16884 ;
  assign n26467 = ~n26461 & ~n26462 ;
  assign n26468 = ~n26466 & n26467 ;
  assign n26472 = ~\P1_EAX_reg[5]/NET0131  & n2313 ;
  assign n26471 = ~\P1_Datao_reg[5]/NET0131  & ~n2313 ;
  assign n26473 = n2432 & ~n26471 ;
  assign n26474 = ~n26472 & n26473 ;
  assign n26469 = \P1_lWord_reg[5]/NET0131  & n2440 ;
  assign n26470 = \P1_Datao_reg[5]/NET0131  & ~n16884 ;
  assign n26475 = ~n26469 & ~n26470 ;
  assign n26476 = ~n26474 & n26475 ;
  assign n26480 = ~\P1_EAX_reg[7]/NET0131  & n2313 ;
  assign n26479 = ~\P1_Datao_reg[7]/NET0131  & ~n2313 ;
  assign n26481 = n2432 & ~n26479 ;
  assign n26482 = ~n26480 & n26481 ;
  assign n26477 = \P1_lWord_reg[7]/NET0131  & n2440 ;
  assign n26478 = \P1_Datao_reg[7]/NET0131  & ~n16884 ;
  assign n26483 = ~n26477 & ~n26478 ;
  assign n26484 = ~n26482 & n26483 ;
  assign n26488 = ~\P1_EAX_reg[9]/NET0131  & n2313 ;
  assign n26487 = ~\P1_Datao_reg[9]/NET0131  & ~n2313 ;
  assign n26489 = n2432 & ~n26487 ;
  assign n26490 = ~n26488 & n26489 ;
  assign n26485 = \P1_lWord_reg[9]/NET0131  & n2440 ;
  assign n26486 = \P1_Datao_reg[9]/NET0131  & ~n16884 ;
  assign n26491 = ~n26485 & ~n26486 ;
  assign n26492 = ~n26490 & n26491 ;
  assign n26496 = ~\P1_EAX_reg[0]/NET0131  & n2313 ;
  assign n26495 = ~\P1_Datao_reg[0]/NET0131  & ~n2313 ;
  assign n26497 = n2432 & ~n26495 ;
  assign n26498 = ~n26496 & n26497 ;
  assign n26493 = \P1_lWord_reg[0]/NET0131  & n2440 ;
  assign n26494 = \P1_Datao_reg[0]/NET0131  & ~n16884 ;
  assign n26499 = ~n26493 & ~n26494 ;
  assign n26500 = ~n26498 & n26499 ;
  assign n26504 = ~\P1_EAX_reg[10]/NET0131  & n2313 ;
  assign n26503 = ~\P1_Datao_reg[10]/NET0131  & ~n2313 ;
  assign n26505 = n2432 & ~n26503 ;
  assign n26506 = ~n26504 & n26505 ;
  assign n26501 = \P1_lWord_reg[10]/NET0131  & n2440 ;
  assign n26502 = \P1_Datao_reg[10]/NET0131  & ~n16884 ;
  assign n26507 = ~n26501 & ~n26502 ;
  assign n26508 = ~n26506 & n26507 ;
  assign n26512 = ~\P1_EAX_reg[11]/NET0131  & n2313 ;
  assign n26511 = ~\P1_Datao_reg[11]/NET0131  & ~n2313 ;
  assign n26513 = n2432 & ~n26511 ;
  assign n26514 = ~n26512 & n26513 ;
  assign n26509 = \P1_lWord_reg[11]/NET0131  & n2440 ;
  assign n26510 = \P1_Datao_reg[11]/NET0131  & ~n16884 ;
  assign n26515 = ~n26509 & ~n26510 ;
  assign n26516 = ~n26514 & n26515 ;
  assign n26520 = ~\P1_EAX_reg[12]/NET0131  & n2313 ;
  assign n26519 = ~\P1_Datao_reg[12]/NET0131  & ~n2313 ;
  assign n26521 = n2432 & ~n26519 ;
  assign n26522 = ~n26520 & n26521 ;
  assign n26517 = \P1_lWord_reg[12]/NET0131  & n2440 ;
  assign n26518 = \P1_Datao_reg[12]/NET0131  & ~n16884 ;
  assign n26523 = ~n26517 & ~n26518 ;
  assign n26524 = ~n26522 & n26523 ;
  assign n26528 = ~\P1_EAX_reg[13]/NET0131  & n2313 ;
  assign n26527 = ~\P1_Datao_reg[13]/NET0131  & ~n2313 ;
  assign n26529 = n2432 & ~n26527 ;
  assign n26530 = ~n26528 & n26529 ;
  assign n26525 = \P1_lWord_reg[13]/NET0131  & n2440 ;
  assign n26526 = \P1_Datao_reg[13]/NET0131  & ~n16884 ;
  assign n26531 = ~n26525 & ~n26526 ;
  assign n26532 = ~n26530 & n26531 ;
  assign n26543 = ~\P3_rEIP_reg[0]/NET0131  & ~\P3_rEIP_reg[1]/NET0131  ;
  assign n26544 = \P3_rEIP_reg[31]/NET0131  & ~n26543 ;
  assign n26545 = \P3_rEIP_reg[2]/NET0131  & n26544 ;
  assign n26546 = \P3_rEIP_reg[3]/NET0131  & n26545 ;
  assign n26547 = \P3_rEIP_reg[4]/NET0131  & n26546 ;
  assign n26548 = \P3_rEIP_reg[5]/NET0131  & n26547 ;
  assign n26549 = \P3_rEIP_reg[6]/NET0131  & n26548 ;
  assign n26550 = \P3_rEIP_reg[7]/NET0131  & n26549 ;
  assign n26551 = \P3_rEIP_reg[8]/NET0131  & n26550 ;
  assign n26552 = \P3_rEIP_reg[9]/NET0131  & n26551 ;
  assign n26553 = \P3_rEIP_reg[10]/NET0131  & n26552 ;
  assign n26554 = \P3_rEIP_reg[11]/NET0131  & n26553 ;
  assign n26555 = \P3_rEIP_reg[12]/NET0131  & n26554 ;
  assign n26556 = \P3_rEIP_reg[13]/NET0131  & n26555 ;
  assign n26557 = \P3_rEIP_reg[14]/NET0131  & n26556 ;
  assign n26558 = \P3_rEIP_reg[15]/NET0131  & n26557 ;
  assign n26559 = \P3_rEIP_reg[16]/NET0131  & n26558 ;
  assign n26560 = n20842 & n26559 ;
  assign n26561 = \P3_rEIP_reg[21]/NET0131  & n26560 ;
  assign n26562 = \P3_rEIP_reg[22]/NET0131  & n26561 ;
  assign n26563 = \P3_rEIP_reg[23]/NET0131  & n26562 ;
  assign n26564 = \P3_rEIP_reg[24]/NET0131  & n26563 ;
  assign n26565 = \P3_rEIP_reg[25]/NET0131  & n26564 ;
  assign n26566 = n21166 & n26565 ;
  assign n26567 = \P3_rEIP_reg[29]/NET0131  & n26566 ;
  assign n26569 = \P3_rEIP_reg[30]/NET0131  & n26567 ;
  assign n26568 = ~\P3_rEIP_reg[30]/NET0131  & ~n26567 ;
  assign n26570 = n2783 & ~n26568 ;
  assign n26571 = ~n26569 & n26570 ;
  assign n26533 = \P3_Address_reg[28]/NET0131  & ~n2782 ;
  assign n26534 = \P3_rEIP_reg[0]/NET0131  & \P3_rEIP_reg[31]/NET0131  ;
  assign n26536 = n20906 & n26534 ;
  assign n26537 = n21027 & n26536 ;
  assign n26538 = n21166 & n26537 ;
  assign n26539 = ~\P3_rEIP_reg[29]/NET0131  & ~n26538 ;
  assign n26535 = n21168 & n26534 ;
  assign n26540 = \P3_State_reg[2]/NET0131  & n2782 ;
  assign n26541 = ~n26535 & n26540 ;
  assign n26542 = ~n26539 & n26541 ;
  assign n26572 = ~n26533 & ~n26542 ;
  assign n26573 = ~n26571 & n26572 ;
  assign n26585 = ~\P2_rEIP_reg[0]/NET0131  & ~\P2_rEIP_reg[1]/NET0131  ;
  assign n26586 = \P2_rEIP_reg[31]/NET0131  & ~n26585 ;
  assign n26587 = \P2_rEIP_reg[2]/NET0131  & n26586 ;
  assign n26588 = \P2_rEIP_reg[3]/NET0131  & n26587 ;
  assign n26589 = \P2_rEIP_reg[4]/NET0131  & n26588 ;
  assign n26590 = n16528 & n26589 ;
  assign n26591 = \P2_rEIP_reg[8]/NET0131  & n26590 ;
  assign n26592 = \P2_rEIP_reg[9]/NET0131  & n26591 ;
  assign n26593 = \P2_rEIP_reg[10]/NET0131  & n26592 ;
  assign n26594 = \P2_rEIP_reg[11]/NET0131  & n26593 ;
  assign n26595 = \P2_rEIP_reg[12]/NET0131  & n26594 ;
  assign n26596 = n16538 & n26595 ;
  assign n26597 = \P2_rEIP_reg[19]/NET0131  & n26596 ;
  assign n26598 = \P2_rEIP_reg[20]/NET0131  & n26597 ;
  assign n26599 = \P2_rEIP_reg[21]/NET0131  & n26598 ;
  assign n26600 = \P2_rEIP_reg[22]/NET0131  & n26599 ;
  assign n26601 = \P2_rEIP_reg[23]/NET0131  & n26600 ;
  assign n26602 = \P2_rEIP_reg[24]/NET0131  & n26601 ;
  assign n26603 = \P2_rEIP_reg[25]/NET0131  & n26602 ;
  assign n26604 = \P2_rEIP_reg[26]/NET0131  & n26603 ;
  assign n26605 = \P2_rEIP_reg[27]/NET0131  & n26604 ;
  assign n26606 = \P2_rEIP_reg[28]/NET0131  & n26605 ;
  assign n26607 = \P2_rEIP_reg[29]/NET0131  & n26606 ;
  assign n26609 = \P2_rEIP_reg[30]/NET0131  & n26607 ;
  assign n26608 = ~\P2_rEIP_reg[30]/NET0131  & ~n26607 ;
  assign n26610 = n1816 & ~n26608 ;
  assign n26611 = ~n26609 & n26610 ;
  assign n26574 = \P2_Address_reg[28]/NET0131  & ~n1815 ;
  assign n26576 = \P2_rEIP_reg[0]/NET0131  & \P2_rEIP_reg[31]/NET0131  ;
  assign n26577 = n16546 & n26576 ;
  assign n26578 = \P2_rEIP_reg[26]/NET0131  & n26577 ;
  assign n26579 = \P2_rEIP_reg[27]/NET0131  & n26578 ;
  assign n26580 = \P2_rEIP_reg[28]/NET0131  & n26579 ;
  assign n26582 = \P2_rEIP_reg[29]/NET0131  & n26580 ;
  assign n26575 = \P2_State_reg[2]/NET0131  & n1815 ;
  assign n26581 = ~\P2_rEIP_reg[29]/NET0131  & ~n26580 ;
  assign n26583 = n26575 & ~n26581 ;
  assign n26584 = ~n26582 & n26583 ;
  assign n26612 = ~n26574 & ~n26584 ;
  assign n26613 = ~n26611 & n26612 ;
  assign n26615 = ~\P1_rEIP_reg[0]/NET0131  & ~\P1_rEIP_reg[1]/NET0131  ;
  assign n26616 = \P1_rEIP_reg[31]/NET0131  & ~n26615 ;
  assign n26617 = \P1_rEIP_reg[2]/NET0131  & n26616 ;
  assign n26618 = \P1_rEIP_reg[3]/NET0131  & n26617 ;
  assign n26619 = \P1_rEIP_reg[4]/NET0131  & n26618 ;
  assign n26620 = \P1_rEIP_reg[5]/NET0131  & n26619 ;
  assign n26621 = \P1_rEIP_reg[6]/NET0131  & n26620 ;
  assign n26622 = \P1_rEIP_reg[7]/NET0131  & n26621 ;
  assign n26623 = \P1_rEIP_reg[8]/NET0131  & n26622 ;
  assign n26624 = \P1_rEIP_reg[9]/NET0131  & n26623 ;
  assign n26625 = \P1_rEIP_reg[10]/NET0131  & n26624 ;
  assign n26626 = \P1_rEIP_reg[11]/NET0131  & n26625 ;
  assign n26627 = \P1_rEIP_reg[12]/NET0131  & n26626 ;
  assign n26628 = \P1_rEIP_reg[13]/NET0131  & n26627 ;
  assign n26629 = \P1_rEIP_reg[14]/NET0131  & n26628 ;
  assign n26630 = \P1_rEIP_reg[15]/NET0131  & n26629 ;
  assign n26631 = \P1_rEIP_reg[16]/NET0131  & n26630 ;
  assign n26632 = \P1_rEIP_reg[17]/NET0131  & n26631 ;
  assign n26633 = n19095 & n26632 ;
  assign n26634 = \P1_rEIP_reg[26]/NET0131  & n26633 ;
  assign n26635 = \P1_rEIP_reg[27]/NET0131  & n26634 ;
  assign n26636 = \P1_rEIP_reg[28]/NET0131  & n26635 ;
  assign n26637 = \P1_rEIP_reg[29]/NET0131  & n26636 ;
  assign n26639 = \P1_rEIP_reg[30]/NET0131  & n26637 ;
  assign n26638 = ~\P1_rEIP_reg[30]/NET0131  & ~n26637 ;
  assign n26640 = n2308 & ~n26638 ;
  assign n26641 = ~n26639 & n26640 ;
  assign n26614 = \address1[28]_pad  & ~n2307 ;
  assign n26642 = \P1_rEIP_reg[0]/NET0131  & \P1_rEIP_reg[31]/NET0131  ;
  assign n26643 = n19206 & n26642 ;
  assign n26644 = \P1_rEIP_reg[27]/NET0131  & n26643 ;
  assign n26645 = \P1_rEIP_reg[28]/NET0131  & n26644 ;
  assign n26648 = \P1_rEIP_reg[29]/NET0131  & n26645 ;
  assign n26646 = ~\P1_rEIP_reg[29]/NET0131  & ~n26645 ;
  assign n26647 = \P1_State_reg[2]/NET0131  & n2307 ;
  assign n26649 = ~n26646 & n26647 ;
  assign n26650 = ~n26648 & n26649 ;
  assign n26651 = ~n26614 & ~n26650 ;
  assign n26652 = ~n26641 & n26651 ;
  assign n26653 = ~\P1_Flush_reg/NET0131  & n3024 ;
  assign n26654 = ~n2432 & ~n2440 ;
  assign n26655 = ~n3028 & n26654 ;
  assign n26656 = ~n26653 & n26655 ;
  assign n26657 = n5288 & n26656 ;
  assign n26658 = \P1_InstQueueWr_Addr_reg[2]/NET0131  & ~n26657 ;
  assign n26659 = ~n5105 & ~n10132 ;
  assign n26660 = \P1_InstQueueWr_Addr_reg[2]/NET0131  & ~n26659 ;
  assign n26661 = ~n7697 & ~n26660 ;
  assign n26662 = ~n3042 & ~n26661 ;
  assign n26663 = n5105 & ~n7697 ;
  assign n26664 = ~\P1_InstQueueWr_Addr_reg[2]/NET0131  & ~n5102 ;
  assign n26665 = ~n3148 & n26664 ;
  assign n26666 = ~n26663 & n26665 ;
  assign n26667 = ~n5325 & ~n26666 ;
  assign n26668 = ~n26662 & n26667 ;
  assign n26669 = ~n26658 & ~n26668 ;
  assign n26672 = ~\P3_Flush_reg/NET0131  & n3010 ;
  assign n26670 = ~n2453 & ~n3004 ;
  assign n26671 = ~n16888 & n26670 ;
  assign n26673 = n21668 & n26671 ;
  assign n26674 = ~n26672 & n26673 ;
  assign n26675 = \P3_InstQueueWr_Addr_reg[2]/NET0131  & ~n26674 ;
  assign n26680 = ~n10075 & ~n18201 ;
  assign n26681 = \P3_InstQueueWr_Addr_reg[2]/NET0131  & ~n26680 ;
  assign n26682 = ~n10074 & ~n26681 ;
  assign n26683 = ~n2994 & ~n26682 ;
  assign n26676 = ~\P3_InstQueueWr_Addr_reg[0]/NET0131  & n10074 ;
  assign n26677 = \P3_InstQueueWr_Addr_reg[1]/NET0131  & ~n26676 ;
  assign n26678 = ~\P3_InstQueueWr_Addr_reg[2]/NET0131  & ~n2970 ;
  assign n26679 = ~n26677 & n26678 ;
  assign n26684 = ~n18211 & ~n26679 ;
  assign n26685 = ~n26683 & n26684 ;
  assign n26686 = ~n26675 & ~n26685 ;
  assign n26689 = n2603 & n18209 ;
  assign n26688 = ~\P3_InstQueue_reg[0][5]/NET0131  & ~n18209 ;
  assign n26690 = n2994 & ~n26688 ;
  assign n26691 = ~n26689 & n26690 ;
  assign n26687 = \P3_InstQueue_reg[0][5]/NET0131  & ~n18218 ;
  assign n26692 = \buf2_reg[29]/NET0131  & n18200 ;
  assign n26693 = \buf2_reg[21]/NET0131  & n18203 ;
  assign n26694 = ~n26692 & ~n26693 ;
  assign n26695 = n2970 & ~n26694 ;
  assign n26696 = \buf2_reg[5]/NET0131  & n18228 ;
  assign n26697 = ~n26695 & ~n26696 ;
  assign n26698 = ~n26687 & n26697 ;
  assign n26699 = ~n26691 & n26698 ;
  assign n26702 = n2603 & n18246 ;
  assign n26701 = ~\P3_InstQueue_reg[10][5]/NET0131  & ~n18246 ;
  assign n26703 = n2994 & ~n26701 ;
  assign n26704 = ~n26702 & n26703 ;
  assign n26700 = \P3_InstQueue_reg[10][5]/NET0131  & ~n18243 ;
  assign n26705 = \buf2_reg[29]/NET0131  & n18233 ;
  assign n26706 = \buf2_reg[21]/NET0131  & n18236 ;
  assign n26707 = ~n26705 & ~n26706 ;
  assign n26708 = n2970 & ~n26707 ;
  assign n26709 = \buf2_reg[5]/NET0131  & n18255 ;
  assign n26710 = ~n26708 & ~n26709 ;
  assign n26711 = ~n26700 & n26710 ;
  assign n26712 = ~n26704 & n26711 ;
  assign n26714 = n2603 & n18266 ;
  assign n26713 = ~\P3_InstQueue_reg[11][5]/NET0131  & ~n18266 ;
  assign n26715 = n2994 & ~n26713 ;
  assign n26716 = ~n26714 & n26715 ;
  assign n26722 = \P3_InstQueue_reg[11][5]/NET0131  & ~n18264 ;
  assign n26717 = ~\P3_InstQueueWr_Addr_reg[0]/NET0131  & ~\buf2_reg[29]/NET0131  ;
  assign n26718 = \P3_InstQueueWr_Addr_reg[0]/NET0131  & ~\buf2_reg[21]/NET0131  ;
  assign n26719 = ~n26717 & ~n26718 ;
  assign n26720 = n2959 & n26719 ;
  assign n26721 = n18260 & n26720 ;
  assign n26723 = \buf2_reg[5]/NET0131  & n18245 ;
  assign n26724 = n18262 & n26723 ;
  assign n26725 = ~n26721 & ~n26724 ;
  assign n26726 = ~n26722 & n26725 ;
  assign n26727 = ~n26716 & n26726 ;
  assign n26730 = n2603 & n18284 ;
  assign n26729 = ~\P3_InstQueue_reg[12][5]/NET0131  & ~n18284 ;
  assign n26731 = n2994 & ~n26729 ;
  assign n26732 = ~n26730 & n26731 ;
  assign n26728 = \P3_InstQueue_reg[12][5]/NET0131  & ~n18287 ;
  assign n26733 = \buf2_reg[21]/NET0131  & n18246 ;
  assign n26734 = \buf2_reg[29]/NET0131  & n18271 ;
  assign n26735 = ~n26733 & ~n26734 ;
  assign n26736 = n2970 & ~n26735 ;
  assign n26737 = \buf2_reg[5]/NET0131  & n18297 ;
  assign n26738 = ~n26736 & ~n26737 ;
  assign n26739 = ~n26728 & n26738 ;
  assign n26740 = ~n26732 & n26739 ;
  assign n26748 = n2603 & n18200 ;
  assign n26747 = ~\P3_InstQueue_reg[13][5]/NET0131  & ~n18200 ;
  assign n26749 = n2994 & ~n26747 ;
  assign n26750 = ~n26748 & n26749 ;
  assign n26744 = ~\P3_InstQueue_reg[13][5]/NET0131  & n18302 ;
  assign n26743 = ~\buf2_reg[5]/NET0131  & ~n18302 ;
  assign n26745 = n18305 & ~n26743 ;
  assign n26746 = ~n26744 & n26745 ;
  assign n26741 = \P3_InstQueue_reg[13][5]/NET0131  & ~n18217 ;
  assign n26742 = n18303 & n26720 ;
  assign n26751 = ~n26741 & ~n26742 ;
  assign n26752 = ~n26746 & n26751 ;
  assign n26753 = ~n26750 & n26752 ;
  assign n26756 = n2603 & n18203 ;
  assign n26755 = ~\P3_InstQueue_reg[14][5]/NET0131  & ~n18203 ;
  assign n26757 = n2994 & ~n26755 ;
  assign n26758 = ~n26756 & n26757 ;
  assign n26754 = \P3_InstQueue_reg[14][5]/NET0131  & ~n18325 ;
  assign n26759 = \buf2_reg[29]/NET0131  & n18266 ;
  assign n26760 = \buf2_reg[21]/NET0131  & n18284 ;
  assign n26761 = ~n26759 & ~n26760 ;
  assign n26762 = n2970 & ~n26761 ;
  assign n26763 = \buf2_reg[5]/NET0131  & n18335 ;
  assign n26764 = ~n26762 & ~n26763 ;
  assign n26765 = ~n26754 & n26764 ;
  assign n26766 = ~n26758 & n26765 ;
  assign n26769 = n2603 & n18212 ;
  assign n26768 = ~\P3_InstQueue_reg[15][5]/NET0131  & ~n18212 ;
  assign n26770 = n2994 & ~n26768 ;
  assign n26771 = ~n26769 & n26770 ;
  assign n26767 = \P3_InstQueue_reg[15][5]/NET0131  & ~n18344 ;
  assign n26772 = \buf2_reg[29]/NET0131  & n18284 ;
  assign n26773 = \buf2_reg[21]/NET0131  & n18200 ;
  assign n26774 = ~n26772 & ~n26773 ;
  assign n26775 = n2970 & ~n26774 ;
  assign n26776 = \buf2_reg[5]/NET0131  & n18354 ;
  assign n26777 = ~n26775 & ~n26776 ;
  assign n26778 = ~n26767 & n26777 ;
  assign n26779 = ~n26771 & n26778 ;
  assign n26782 = n2603 & n18361 ;
  assign n26781 = ~\P3_InstQueue_reg[1][5]/NET0131  & ~n18361 ;
  assign n26783 = n2994 & ~n26781 ;
  assign n26784 = ~n26782 & n26783 ;
  assign n26780 = \P3_InstQueue_reg[1][5]/NET0131  & ~n18364 ;
  assign n26785 = \buf2_reg[29]/NET0131  & n18203 ;
  assign n26786 = \buf2_reg[21]/NET0131  & n18212 ;
  assign n26787 = ~n26785 & ~n26786 ;
  assign n26788 = n2970 & ~n26787 ;
  assign n26789 = \buf2_reg[5]/NET0131  & n18374 ;
  assign n26790 = ~n26788 & ~n26789 ;
  assign n26791 = ~n26780 & n26790 ;
  assign n26792 = ~n26784 & n26791 ;
  assign n26795 = n2603 & n18386 ;
  assign n26794 = ~\P3_InstQueue_reg[2][5]/NET0131  & ~n18386 ;
  assign n26796 = n2994 & ~n26794 ;
  assign n26797 = ~n26795 & n26796 ;
  assign n26793 = \P3_InstQueue_reg[2][5]/NET0131  & ~n18383 ;
  assign n26798 = \buf2_reg[29]/NET0131  & n18212 ;
  assign n26799 = \buf2_reg[21]/NET0131  & n18209 ;
  assign n26800 = ~n26798 & ~n26799 ;
  assign n26801 = n2970 & ~n26800 ;
  assign n26802 = \buf2_reg[5]/NET0131  & n18395 ;
  assign n26803 = ~n26801 & ~n26802 ;
  assign n26804 = ~n26793 & n26803 ;
  assign n26805 = ~n26797 & n26804 ;
  assign n26808 = n2603 & n18405 ;
  assign n26807 = ~\P3_InstQueue_reg[3][5]/NET0131  & ~n18405 ;
  assign n26809 = n2994 & ~n26807 ;
  assign n26810 = ~n26808 & n26809 ;
  assign n26806 = \P3_InstQueue_reg[3][5]/NET0131  & ~n18403 ;
  assign n26811 = \buf2_reg[21]/NET0131  & n18361 ;
  assign n26812 = \buf2_reg[29]/NET0131  & n18209 ;
  assign n26813 = ~n26811 & ~n26812 ;
  assign n26814 = n2970 & ~n26813 ;
  assign n26815 = \buf2_reg[5]/NET0131  & n18414 ;
  assign n26816 = ~n26814 & ~n26815 ;
  assign n26817 = ~n26806 & n26816 ;
  assign n26818 = ~n26810 & n26817 ;
  assign n26821 = n2603 & n18421 ;
  assign n26820 = ~\P3_InstQueue_reg[4][5]/NET0131  & ~n18421 ;
  assign n26822 = n2994 & ~n26820 ;
  assign n26823 = ~n26821 & n26822 ;
  assign n26819 = \P3_InstQueue_reg[4][5]/NET0131  & ~n18424 ;
  assign n26824 = \buf2_reg[21]/NET0131  & n18386 ;
  assign n26825 = \buf2_reg[29]/NET0131  & n18361 ;
  assign n26826 = ~n26824 & ~n26825 ;
  assign n26827 = n2970 & ~n26826 ;
  assign n26828 = \buf2_reg[5]/NET0131  & n18434 ;
  assign n26829 = ~n26827 & ~n26828 ;
  assign n26830 = ~n26819 & n26829 ;
  assign n26831 = ~n26823 & n26830 ;
  assign n26839 = n2603 & n18439 ;
  assign n26838 = ~\P3_InstQueue_reg[5][5]/NET0131  & ~n18439 ;
  assign n26840 = n2994 & ~n26838 ;
  assign n26841 = ~n26839 & n26840 ;
  assign n26835 = ~\P3_InstQueue_reg[5][5]/NET0131  & n18440 ;
  assign n26834 = ~\buf2_reg[5]/NET0131  & ~n18440 ;
  assign n26836 = n18443 & ~n26834 ;
  assign n26837 = ~n26835 & n26836 ;
  assign n26832 = \P3_InstQueue_reg[5][5]/NET0131  & ~n18217 ;
  assign n26833 = n18441 & n26720 ;
  assign n26842 = ~n26832 & ~n26833 ;
  assign n26843 = ~n26837 & n26842 ;
  assign n26844 = ~n26841 & n26843 ;
  assign n26847 = n2603 & n18462 ;
  assign n26846 = ~\P3_InstQueue_reg[6][5]/NET0131  & ~n18462 ;
  assign n26848 = n2994 & ~n26846 ;
  assign n26849 = ~n26847 & n26848 ;
  assign n26845 = \P3_InstQueue_reg[6][5]/NET0131  & ~n18465 ;
  assign n26850 = \buf2_reg[29]/NET0131  & n18405 ;
  assign n26851 = \buf2_reg[21]/NET0131  & n18421 ;
  assign n26852 = ~n26850 & ~n26851 ;
  assign n26853 = n2970 & ~n26852 ;
  assign n26854 = \buf2_reg[5]/NET0131  & n18475 ;
  assign n26855 = ~n26853 & ~n26854 ;
  assign n26856 = ~n26845 & n26855 ;
  assign n26857 = ~n26849 & n26856 ;
  assign n26860 = n2603 & n18233 ;
  assign n26859 = ~\P3_InstQueue_reg[7][5]/NET0131  & ~n18233 ;
  assign n26861 = n2994 & ~n26859 ;
  assign n26862 = ~n26860 & n26861 ;
  assign n26858 = \P3_InstQueue_reg[7][5]/NET0131  & ~n18484 ;
  assign n26863 = \buf2_reg[29]/NET0131  & n18421 ;
  assign n26864 = \buf2_reg[21]/NET0131  & n18439 ;
  assign n26865 = ~n26863 & ~n26864 ;
  assign n26866 = n2970 & ~n26865 ;
  assign n26867 = \buf2_reg[5]/NET0131  & n18494 ;
  assign n26868 = ~n26866 & ~n26867 ;
  assign n26869 = ~n26858 & n26868 ;
  assign n26870 = ~n26862 & n26869 ;
  assign n26873 = n2603 & n18236 ;
  assign n26872 = ~\P3_InstQueue_reg[8][5]/NET0131  & ~n18236 ;
  assign n26874 = n2994 & ~n26872 ;
  assign n26875 = ~n26873 & n26874 ;
  assign n26871 = \P3_InstQueue_reg[8][5]/NET0131  & ~n18502 ;
  assign n26876 = \buf2_reg[29]/NET0131  & n18439 ;
  assign n26877 = \buf2_reg[21]/NET0131  & n18462 ;
  assign n26878 = ~n26876 & ~n26877 ;
  assign n26879 = n2970 & ~n26878 ;
  assign n26880 = \buf2_reg[5]/NET0131  & n18512 ;
  assign n26881 = ~n26879 & ~n26880 ;
  assign n26882 = ~n26871 & n26881 ;
  assign n26883 = ~n26875 & n26882 ;
  assign n26897 = n2603 & n18271 ;
  assign n26896 = ~\P3_InstQueue_reg[9][5]/NET0131  & ~n18271 ;
  assign n26898 = n2994 & ~n26896 ;
  assign n26899 = ~n26897 & n26898 ;
  assign n26888 = \buf2_reg[29]/NET0131  & n18462 ;
  assign n26889 = \buf2_reg[21]/NET0131  & n18233 ;
  assign n26890 = ~n26888 & ~n26889 ;
  assign n26891 = \P3_DataWidth_reg[1]/NET0131  & ~n26890 ;
  assign n26884 = \P3_InstQueue_reg[9][5]/NET0131  & ~n18235 ;
  assign n26885 = \buf2_reg[5]/NET0131  & n18235 ;
  assign n26886 = ~n26884 & ~n26885 ;
  assign n26892 = ~n18525 & ~n26886 ;
  assign n26893 = ~n26891 & ~n26892 ;
  assign n26894 = n2959 & ~n26893 ;
  assign n26887 = n4415 & ~n26886 ;
  assign n26895 = \P3_InstQueue_reg[9][5]/NET0131  & ~n18217 ;
  assign n26900 = ~n26887 & ~n26895 ;
  assign n26901 = ~n26894 & n26900 ;
  assign n26902 = ~n26899 & n26901 ;
  assign n26903 = ~\P2_Flush_reg/NET0131  & n2984 ;
  assign n26904 = ~n1927 & ~n2987 ;
  assign n26905 = ~n16919 & n26904 ;
  assign n26906 = ~n26903 & n26905 ;
  assign n26907 = n21640 & n26906 ;
  assign n26908 = \P2_InstQueueWr_Addr_reg[2]/NET0131  & ~n26907 ;
  assign n26909 = ~n3044 & ~n9004 ;
  assign n26910 = \P2_InstQueueWr_Addr_reg[2]/NET0131  & ~n26909 ;
  assign n26911 = ~n3125 & ~n26910 ;
  assign n26912 = ~n3040 & ~n26911 ;
  assign n26913 = n3044 & ~n3125 ;
  assign n26914 = ~\P2_InstQueueWr_Addr_reg[2]/NET0131  & ~n3047 ;
  assign n26915 = ~n3034 & n26914 ;
  assign n26916 = ~n26913 & n26915 ;
  assign n26917 = ~n3153 & ~n26916 ;
  assign n26918 = ~n26912 & n26917 ;
  assign n26919 = ~n26908 & ~n26918 ;
  assign n26922 = \P3_rEIP_reg[17]/NET0131  & n26559 ;
  assign n26923 = ~\P3_rEIP_reg[18]/NET0131  & ~n26922 ;
  assign n26921 = n20727 & n26559 ;
  assign n26924 = n2783 & ~n26921 ;
  assign n26925 = ~n26923 & n26924 ;
  assign n26920 = \P3_Address_reg[16]/NET0131  & ~n2782 ;
  assign n26926 = n20575 & n26534 ;
  assign n26927 = \P3_rEIP_reg[15]/NET0131  & n26926 ;
  assign n26928 = \P3_rEIP_reg[16]/NET0131  & n26927 ;
  assign n26930 = ~\P3_rEIP_reg[17]/NET0131  & ~n26928 ;
  assign n26929 = \P3_rEIP_reg[17]/NET0131  & n26928 ;
  assign n26931 = n26540 & ~n26929 ;
  assign n26932 = ~n26930 & n26931 ;
  assign n26933 = ~n26920 & ~n26932 ;
  assign n26934 = ~n26925 & n26933 ;
  assign n26940 = n16537 & n26595 ;
  assign n26941 = ~\P2_rEIP_reg[18]/NET0131  & ~n26940 ;
  assign n26942 = n1816 & ~n26596 ;
  assign n26943 = ~n26941 & n26942 ;
  assign n26935 = \P2_Address_reg[16]/NET0131  & ~n1815 ;
  assign n26937 = ~n19395 & n26576 ;
  assign n26936 = ~\P2_rEIP_reg[17]/NET0131  & ~n26576 ;
  assign n26938 = n26575 & ~n26936 ;
  assign n26939 = ~n26937 & n26938 ;
  assign n26944 = ~n26935 & ~n26939 ;
  assign n26945 = ~n26943 & n26944 ;
  assign n26952 = ~\P1_rEIP_reg[18]/NET0131  & ~n26632 ;
  assign n26951 = \P1_rEIP_reg[18]/NET0131  & n26632 ;
  assign n26953 = n2308 & ~n26951 ;
  assign n26954 = ~n26952 & n26953 ;
  assign n26946 = \address1[16]_pad  & ~n2307 ;
  assign n26948 = ~n18697 & n26642 ;
  assign n26947 = ~\P1_rEIP_reg[17]/NET0131  & ~n26642 ;
  assign n26949 = n26647 & ~n26947 ;
  assign n26950 = ~n26948 & n26949 ;
  assign n26955 = ~n26946 & ~n26950 ;
  assign n26956 = ~n26954 & n26955 ;
  assign n26957 = ~\P1_InstQueueWr_Addr_reg[3]/NET0131  & ~n5325 ;
  assign n26958 = ~n5326 & ~n26957 ;
  assign n26960 = ~n5335 & n26958 ;
  assign n26961 = ~n5571 & ~n26960 ;
  assign n26962 = ~n5333 & ~n26961 ;
  assign n26963 = ~n5376 & ~n5549 ;
  assign n26964 = ~n26962 & n26963 ;
  assign n26965 = n3148 & ~n5377 ;
  assign n26966 = ~n26964 & n26965 ;
  assign n26967 = \P1_InstQueueWr_Addr_reg[3]/NET0131  & ~n26657 ;
  assign n26959 = n3042 & n26958 ;
  assign n26968 = n10133 & ~n26961 ;
  assign n26969 = ~n26959 & ~n26968 ;
  assign n26970 = ~n26967 & n26969 ;
  assign n26971 = ~n26966 & n26970 ;
  assign n26972 = ~\P3_InstQueueWr_Addr_reg[3]/NET0131  & ~n18211 ;
  assign n26973 = ~n18212 & ~n26972 ;
  assign n26975 = ~n18202 & n26973 ;
  assign n26976 = ~n18462 & ~n26975 ;
  assign n26977 = ~n18199 & ~n26976 ;
  assign n26978 = ~n18283 & ~n18439 ;
  assign n26979 = ~n26977 & n26978 ;
  assign n26980 = n2970 & ~n18284 ;
  assign n26981 = ~n26979 & n26980 ;
  assign n26982 = \P3_InstQueueWr_Addr_reg[3]/NET0131  & ~n26674 ;
  assign n26974 = n2994 & n26973 ;
  assign n26983 = n10076 & ~n26976 ;
  assign n26984 = ~n26974 & ~n26983 ;
  assign n26985 = ~n26982 & n26984 ;
  assign n26986 = ~n26981 & n26985 ;
  assign n26987 = \P2_InstQueueWr_Addr_reg[3]/NET0131  & ~n3153 ;
  assign n26988 = ~n3198 & ~n26987 ;
  assign n26990 = ~n3164 & ~n26988 ;
  assign n26991 = ~n3575 & ~n26990 ;
  assign n26992 = ~n3161 & ~n26991 ;
  assign n26993 = ~n3236 & ~n3537 ;
  assign n26994 = ~n26992 & n26993 ;
  assign n26995 = n3034 & ~n3237 ;
  assign n26996 = ~n26994 & n26995 ;
  assign n26997 = \P2_InstQueueWr_Addr_reg[3]/NET0131  & ~n26907 ;
  assign n26989 = n3040 & ~n26988 ;
  assign n26998 = n9005 & ~n26991 ;
  assign n26999 = ~n26989 & ~n26998 ;
  assign n27000 = ~n26997 & n26999 ;
  assign n27001 = ~n26996 & n27000 ;
  assign n27002 = \P1_InstQueueWr_Addr_reg[1]/NET0131  & ~n26656 ;
  assign n27003 = ~\P1_InstQueueWr_Addr_reg[0]/NET0131  & n3042 ;
  assign n27004 = \P1_InstQueueWr_Addr_reg[1]/NET0131  & n5288 ;
  assign n27005 = ~n3148 & n27004 ;
  assign n27006 = ~n27003 & n27005 ;
  assign n27007 = \P1_InstQueueWr_Addr_reg[0]/NET0131  & n3042 ;
  assign n27008 = ~\P1_InstQueueWr_Addr_reg[1]/NET0131  & ~n27007 ;
  assign n27009 = ~n10133 & n27008 ;
  assign n27010 = ~n27006 & ~n27009 ;
  assign n27011 = ~n27002 & ~n27010 ;
  assign n27013 = ~n2970 & n26674 ;
  assign n27014 = \P3_InstQueueWr_Addr_reg[1]/NET0131  & ~n27013 ;
  assign n27012 = ~\P3_InstQueueWr_Addr_reg[1]/NET0131  & n10076 ;
  assign n27015 = n2994 & ~n18240 ;
  assign n27016 = ~n27012 & ~n27015 ;
  assign n27017 = ~n27014 & n27016 ;
  assign n27018 = \P2_InstQueueWr_Addr_reg[1]/NET0131  & ~n26906 ;
  assign n27019 = ~\P2_InstQueueWr_Addr_reg[0]/NET0131  & n3040 ;
  assign n27020 = \P2_InstQueueWr_Addr_reg[1]/NET0131  & n21640 ;
  assign n27021 = ~n3034 & n27020 ;
  assign n27022 = ~n27019 & n27021 ;
  assign n27023 = \P2_InstQueueWr_Addr_reg[0]/NET0131  & n3040 ;
  assign n27024 = ~\P2_InstQueueWr_Addr_reg[1]/NET0131  & ~n27023 ;
  assign n27025 = ~n9005 & n27024 ;
  assign n27026 = ~n27022 & ~n27025 ;
  assign n27027 = ~n27018 & ~n27026 ;
  assign n27030 = ~n2435 & n3146 ;
  assign n27031 = n14084 & n27030 ;
  assign n27032 = \P1_InstQueueWr_Addr_reg[0]/NET0131  & ~n27031 ;
  assign n27028 = ~\P1_Flush_reg/NET0131  & ~\P1_InstQueueWr_Addr_reg[0]/NET0131  ;
  assign n27029 = n3024 & ~n27028 ;
  assign n27033 = ~n27003 & ~n27029 ;
  assign n27034 = ~n27032 & n27033 ;
  assign n27038 = n4416 & n15433 ;
  assign n27039 = n26671 & n27038 ;
  assign n27040 = \P3_InstQueueWr_Addr_reg[0]/NET0131  & ~n27039 ;
  assign n27035 = ~\P3_InstQueueWr_Addr_reg[0]/NET0131  & n2994 ;
  assign n27036 = ~\P3_Flush_reg/NET0131  & ~\P3_InstQueueWr_Addr_reg[0]/NET0131  ;
  assign n27037 = n3010 & ~n27036 ;
  assign n27041 = ~n27035 & ~n27037 ;
  assign n27042 = ~n27040 & n27041 ;
  assign n27045 = n2698 & n18209 ;
  assign n27044 = ~\P3_InstQueue_reg[0][1]/NET0131  & ~n18209 ;
  assign n27046 = n2994 & ~n27044 ;
  assign n27047 = ~n27045 & n27046 ;
  assign n27043 = \P3_InstQueue_reg[0][1]/NET0131  & ~n18218 ;
  assign n27048 = \buf2_reg[25]/NET0131  & n18200 ;
  assign n27049 = \buf2_reg[17]/NET0131  & n18203 ;
  assign n27050 = ~n27048 & ~n27049 ;
  assign n27051 = n2970 & ~n27050 ;
  assign n27052 = \buf2_reg[1]/NET0131  & n18228 ;
  assign n27053 = ~n27051 & ~n27052 ;
  assign n27054 = ~n27043 & n27053 ;
  assign n27055 = ~n27047 & n27054 ;
  assign n27058 = n2698 & n18246 ;
  assign n27057 = ~\P3_InstQueue_reg[10][1]/NET0131  & ~n18246 ;
  assign n27059 = n2994 & ~n27057 ;
  assign n27060 = ~n27058 & n27059 ;
  assign n27056 = \P3_InstQueue_reg[10][1]/NET0131  & ~n18243 ;
  assign n27061 = \buf2_reg[25]/NET0131  & n18233 ;
  assign n27062 = \buf2_reg[17]/NET0131  & n18236 ;
  assign n27063 = ~n27061 & ~n27062 ;
  assign n27064 = n2970 & ~n27063 ;
  assign n27065 = \buf2_reg[1]/NET0131  & n18255 ;
  assign n27066 = ~n27064 & ~n27065 ;
  assign n27067 = ~n27056 & n27066 ;
  assign n27068 = ~n27060 & n27067 ;
  assign n27070 = n2666 & n18266 ;
  assign n27069 = ~\P3_InstQueue_reg[11][0]/NET0131  & ~n18266 ;
  assign n27071 = n2994 & ~n27069 ;
  assign n27072 = ~n27070 & n27071 ;
  assign n27078 = \P3_InstQueue_reg[11][0]/NET0131  & ~n18264 ;
  assign n27073 = ~\P3_InstQueueWr_Addr_reg[0]/NET0131  & ~\buf2_reg[24]/NET0131  ;
  assign n27074 = \P3_InstQueueWr_Addr_reg[0]/NET0131  & ~\buf2_reg[16]/NET0131  ;
  assign n27075 = ~n27073 & ~n27074 ;
  assign n27076 = n2959 & n27075 ;
  assign n27077 = n18260 & n27076 ;
  assign n27079 = \buf2_reg[0]/NET0131  & n18245 ;
  assign n27080 = n18262 & n27079 ;
  assign n27081 = ~n27077 & ~n27080 ;
  assign n27082 = ~n27078 & n27081 ;
  assign n27083 = ~n27072 & n27082 ;
  assign n27085 = n2698 & n18266 ;
  assign n27084 = ~\P3_InstQueue_reg[11][1]/NET0131  & ~n18266 ;
  assign n27086 = n2994 & ~n27084 ;
  assign n27087 = ~n27085 & n27086 ;
  assign n27093 = \P3_InstQueue_reg[11][1]/NET0131  & ~n18264 ;
  assign n27088 = ~\P3_InstQueueWr_Addr_reg[0]/NET0131  & ~\buf2_reg[25]/NET0131  ;
  assign n27089 = \P3_InstQueueWr_Addr_reg[0]/NET0131  & ~\buf2_reg[17]/NET0131  ;
  assign n27090 = ~n27088 & ~n27089 ;
  assign n27091 = n2959 & n27090 ;
  assign n27092 = n18260 & n27091 ;
  assign n27094 = \buf2_reg[1]/NET0131  & n18245 ;
  assign n27095 = n18262 & n27094 ;
  assign n27096 = ~n27092 & ~n27095 ;
  assign n27097 = ~n27093 & n27096 ;
  assign n27098 = ~n27087 & n27097 ;
  assign n27101 = n2698 & n18284 ;
  assign n27100 = ~\P3_InstQueue_reg[12][1]/NET0131  & ~n18284 ;
  assign n27102 = n2994 & ~n27100 ;
  assign n27103 = ~n27101 & n27102 ;
  assign n27099 = \P3_InstQueue_reg[12][1]/NET0131  & ~n18287 ;
  assign n27104 = \buf2_reg[17]/NET0131  & n18246 ;
  assign n27105 = \buf2_reg[25]/NET0131  & n18271 ;
  assign n27106 = ~n27104 & ~n27105 ;
  assign n27107 = n2970 & ~n27106 ;
  assign n27108 = \buf2_reg[1]/NET0131  & n18297 ;
  assign n27109 = ~n27107 & ~n27108 ;
  assign n27110 = ~n27099 & n27109 ;
  assign n27111 = ~n27103 & n27110 ;
  assign n27119 = n2698 & n18200 ;
  assign n27118 = ~\P3_InstQueue_reg[13][1]/NET0131  & ~n18200 ;
  assign n27120 = n2994 & ~n27118 ;
  assign n27121 = ~n27119 & n27120 ;
  assign n27115 = ~\P3_InstQueue_reg[13][1]/NET0131  & n18302 ;
  assign n27114 = ~\buf2_reg[1]/NET0131  & ~n18302 ;
  assign n27116 = n18305 & ~n27114 ;
  assign n27117 = ~n27115 & n27116 ;
  assign n27112 = \P3_InstQueue_reg[13][1]/NET0131  & ~n18217 ;
  assign n27113 = n18303 & n27091 ;
  assign n27122 = ~n27112 & ~n27113 ;
  assign n27123 = ~n27117 & n27122 ;
  assign n27124 = ~n27121 & n27123 ;
  assign n27127 = n2698 & n18203 ;
  assign n27126 = ~\P3_InstQueue_reg[14][1]/NET0131  & ~n18203 ;
  assign n27128 = n2994 & ~n27126 ;
  assign n27129 = ~n27127 & n27128 ;
  assign n27125 = \P3_InstQueue_reg[14][1]/NET0131  & ~n18325 ;
  assign n27130 = \buf2_reg[25]/NET0131  & n18266 ;
  assign n27131 = \buf2_reg[17]/NET0131  & n18284 ;
  assign n27132 = ~n27130 & ~n27131 ;
  assign n27133 = n2970 & ~n27132 ;
  assign n27134 = \buf2_reg[1]/NET0131  & n18335 ;
  assign n27135 = ~n27133 & ~n27134 ;
  assign n27136 = ~n27125 & n27135 ;
  assign n27137 = ~n27129 & n27136 ;
  assign n27140 = n2698 & n18212 ;
  assign n27139 = ~\P3_InstQueue_reg[15][1]/NET0131  & ~n18212 ;
  assign n27141 = n2994 & ~n27139 ;
  assign n27142 = ~n27140 & n27141 ;
  assign n27138 = \P3_InstQueue_reg[15][1]/NET0131  & ~n18344 ;
  assign n27143 = \buf2_reg[25]/NET0131  & n18284 ;
  assign n27144 = \buf2_reg[17]/NET0131  & n18200 ;
  assign n27145 = ~n27143 & ~n27144 ;
  assign n27146 = n2970 & ~n27145 ;
  assign n27147 = \buf2_reg[1]/NET0131  & n18354 ;
  assign n27148 = ~n27146 & ~n27147 ;
  assign n27149 = ~n27138 & n27148 ;
  assign n27150 = ~n27142 & n27149 ;
  assign n27153 = n2698 & n18361 ;
  assign n27152 = ~\P3_InstQueue_reg[1][1]/NET0131  & ~n18361 ;
  assign n27154 = n2994 & ~n27152 ;
  assign n27155 = ~n27153 & n27154 ;
  assign n27151 = \P3_InstQueue_reg[1][1]/NET0131  & ~n18364 ;
  assign n27156 = \buf2_reg[25]/NET0131  & n18203 ;
  assign n27157 = \buf2_reg[17]/NET0131  & n18212 ;
  assign n27158 = ~n27156 & ~n27157 ;
  assign n27159 = n2970 & ~n27158 ;
  assign n27160 = \buf2_reg[1]/NET0131  & n18374 ;
  assign n27161 = ~n27159 & ~n27160 ;
  assign n27162 = ~n27151 & n27161 ;
  assign n27163 = ~n27155 & n27162 ;
  assign n27166 = n2698 & n18386 ;
  assign n27165 = ~\P3_InstQueue_reg[2][1]/NET0131  & ~n18386 ;
  assign n27167 = n2994 & ~n27165 ;
  assign n27168 = ~n27166 & n27167 ;
  assign n27164 = \P3_InstQueue_reg[2][1]/NET0131  & ~n18383 ;
  assign n27169 = \buf2_reg[25]/NET0131  & n18212 ;
  assign n27170 = \buf2_reg[17]/NET0131  & n18209 ;
  assign n27171 = ~n27169 & ~n27170 ;
  assign n27172 = n2970 & ~n27171 ;
  assign n27173 = \buf2_reg[1]/NET0131  & n18395 ;
  assign n27174 = ~n27172 & ~n27173 ;
  assign n27175 = ~n27164 & n27174 ;
  assign n27176 = ~n27168 & n27175 ;
  assign n27179 = n2666 & n18405 ;
  assign n27178 = ~\P3_InstQueue_reg[3][0]/NET0131  & ~n18405 ;
  assign n27180 = n2994 & ~n27178 ;
  assign n27181 = ~n27179 & n27180 ;
  assign n27177 = \P3_InstQueue_reg[3][0]/NET0131  & ~n18403 ;
  assign n27182 = \buf2_reg[16]/NET0131  & n18361 ;
  assign n27183 = \buf2_reg[24]/NET0131  & n18209 ;
  assign n27184 = ~n27182 & ~n27183 ;
  assign n27185 = n2970 & ~n27184 ;
  assign n27186 = \buf2_reg[0]/NET0131  & n18414 ;
  assign n27187 = ~n27185 & ~n27186 ;
  assign n27188 = ~n27177 & n27187 ;
  assign n27189 = ~n27181 & n27188 ;
  assign n27192 = n2698 & n18405 ;
  assign n27191 = ~\P3_InstQueue_reg[3][1]/NET0131  & ~n18405 ;
  assign n27193 = n2994 & ~n27191 ;
  assign n27194 = ~n27192 & n27193 ;
  assign n27190 = \P3_InstQueue_reg[3][1]/NET0131  & ~n18403 ;
  assign n27195 = \buf2_reg[17]/NET0131  & n18361 ;
  assign n27196 = \buf2_reg[25]/NET0131  & n18209 ;
  assign n27197 = ~n27195 & ~n27196 ;
  assign n27198 = n2970 & ~n27197 ;
  assign n27199 = \buf2_reg[1]/NET0131  & n18414 ;
  assign n27200 = ~n27198 & ~n27199 ;
  assign n27201 = ~n27190 & n27200 ;
  assign n27202 = ~n27194 & n27201 ;
  assign n27205 = n2698 & n18421 ;
  assign n27204 = ~\P3_InstQueue_reg[4][1]/NET0131  & ~n18421 ;
  assign n27206 = n2994 & ~n27204 ;
  assign n27207 = ~n27205 & n27206 ;
  assign n27203 = \P3_InstQueue_reg[4][1]/NET0131  & ~n18424 ;
  assign n27208 = \buf2_reg[17]/NET0131  & n18386 ;
  assign n27209 = \buf2_reg[25]/NET0131  & n18361 ;
  assign n27210 = ~n27208 & ~n27209 ;
  assign n27211 = n2970 & ~n27210 ;
  assign n27212 = \buf2_reg[1]/NET0131  & n18434 ;
  assign n27213 = ~n27211 & ~n27212 ;
  assign n27214 = ~n27203 & n27213 ;
  assign n27215 = ~n27207 & n27214 ;
  assign n27223 = n2698 & n18439 ;
  assign n27222 = ~\P3_InstQueue_reg[5][1]/NET0131  & ~n18439 ;
  assign n27224 = n2994 & ~n27222 ;
  assign n27225 = ~n27223 & n27224 ;
  assign n27219 = ~\P3_InstQueue_reg[5][1]/NET0131  & n18440 ;
  assign n27218 = ~\buf2_reg[1]/NET0131  & ~n18440 ;
  assign n27220 = n18443 & ~n27218 ;
  assign n27221 = ~n27219 & n27220 ;
  assign n27216 = \P3_InstQueue_reg[5][1]/NET0131  & ~n18217 ;
  assign n27217 = n18441 & n27091 ;
  assign n27226 = ~n27216 & ~n27217 ;
  assign n27227 = ~n27221 & n27226 ;
  assign n27228 = ~n27225 & n27227 ;
  assign n27231 = n2698 & n18462 ;
  assign n27230 = ~\P3_InstQueue_reg[6][1]/NET0131  & ~n18462 ;
  assign n27232 = n2994 & ~n27230 ;
  assign n27233 = ~n27231 & n27232 ;
  assign n27229 = \P3_InstQueue_reg[6][1]/NET0131  & ~n18465 ;
  assign n27234 = \buf2_reg[25]/NET0131  & n18405 ;
  assign n27235 = \buf2_reg[17]/NET0131  & n18421 ;
  assign n27236 = ~n27234 & ~n27235 ;
  assign n27237 = n2970 & ~n27236 ;
  assign n27238 = \buf2_reg[1]/NET0131  & n18475 ;
  assign n27239 = ~n27237 & ~n27238 ;
  assign n27240 = ~n27229 & n27239 ;
  assign n27241 = ~n27233 & n27240 ;
  assign n27244 = n2666 & n18233 ;
  assign n27243 = ~\P3_InstQueue_reg[7][0]/NET0131  & ~n18233 ;
  assign n27245 = n2994 & ~n27243 ;
  assign n27246 = ~n27244 & n27245 ;
  assign n27242 = \P3_InstQueue_reg[7][0]/NET0131  & ~n18484 ;
  assign n27247 = \buf2_reg[24]/NET0131  & n18421 ;
  assign n27248 = \buf2_reg[16]/NET0131  & n18439 ;
  assign n27249 = ~n27247 & ~n27248 ;
  assign n27250 = n2970 & ~n27249 ;
  assign n27251 = \buf2_reg[0]/NET0131  & n18494 ;
  assign n27252 = ~n27250 & ~n27251 ;
  assign n27253 = ~n27242 & n27252 ;
  assign n27254 = ~n27246 & n27253 ;
  assign n27257 = n2698 & n18233 ;
  assign n27256 = ~\P3_InstQueue_reg[7][1]/NET0131  & ~n18233 ;
  assign n27258 = n2994 & ~n27256 ;
  assign n27259 = ~n27257 & n27258 ;
  assign n27255 = \P3_InstQueue_reg[7][1]/NET0131  & ~n18484 ;
  assign n27260 = \buf2_reg[25]/NET0131  & n18421 ;
  assign n27261 = \buf2_reg[17]/NET0131  & n18439 ;
  assign n27262 = ~n27260 & ~n27261 ;
  assign n27263 = n2970 & ~n27262 ;
  assign n27264 = \buf2_reg[1]/NET0131  & n18494 ;
  assign n27265 = ~n27263 & ~n27264 ;
  assign n27266 = ~n27255 & n27265 ;
  assign n27267 = ~n27259 & n27266 ;
  assign n27270 = n2698 & n18236 ;
  assign n27269 = ~\P3_InstQueue_reg[8][1]/NET0131  & ~n18236 ;
  assign n27271 = n2994 & ~n27269 ;
  assign n27272 = ~n27270 & n27271 ;
  assign n27268 = \P3_InstQueue_reg[8][1]/NET0131  & ~n18502 ;
  assign n27273 = \buf2_reg[25]/NET0131  & n18439 ;
  assign n27274 = \buf2_reg[17]/NET0131  & n18462 ;
  assign n27275 = ~n27273 & ~n27274 ;
  assign n27276 = n2970 & ~n27275 ;
  assign n27277 = \buf2_reg[1]/NET0131  & n18512 ;
  assign n27278 = ~n27276 & ~n27277 ;
  assign n27279 = ~n27268 & n27278 ;
  assign n27280 = ~n27272 & n27279 ;
  assign n27294 = n2698 & n18271 ;
  assign n27293 = ~\P3_InstQueue_reg[9][1]/NET0131  & ~n18271 ;
  assign n27295 = n2994 & ~n27293 ;
  assign n27296 = ~n27294 & n27295 ;
  assign n27285 = \buf2_reg[25]/NET0131  & n18462 ;
  assign n27286 = \buf2_reg[17]/NET0131  & n18233 ;
  assign n27287 = ~n27285 & ~n27286 ;
  assign n27288 = \P3_DataWidth_reg[1]/NET0131  & ~n27287 ;
  assign n27281 = \P3_InstQueue_reg[9][1]/NET0131  & ~n18235 ;
  assign n27282 = \buf2_reg[1]/NET0131  & n18235 ;
  assign n27283 = ~n27281 & ~n27282 ;
  assign n27289 = ~n18525 & ~n27283 ;
  assign n27290 = ~n27288 & ~n27289 ;
  assign n27291 = n2959 & ~n27290 ;
  assign n27284 = n4415 & ~n27283 ;
  assign n27292 = \P3_InstQueue_reg[9][1]/NET0131  & ~n18217 ;
  assign n27297 = ~n27284 & ~n27292 ;
  assign n27298 = ~n27291 & n27297 ;
  assign n27299 = ~n27296 & n27298 ;
  assign n27302 = ~n1927 & n14133 ;
  assign n27303 = \P2_InstQueueWr_Addr_reg[0]/NET0131  & ~n27302 ;
  assign n27300 = ~\P2_Flush_reg/NET0131  & ~\P2_InstQueueWr_Addr_reg[0]/NET0131  ;
  assign n27301 = n2984 & ~n27300 ;
  assign n27304 = ~n27019 & ~n27301 ;
  assign n27305 = ~n27303 & n27304 ;
  assign n27308 = \P3_rEIP_reg[26]/NET0131  & n26565 ;
  assign n27307 = ~\P3_rEIP_reg[26]/NET0131  & ~n26565 ;
  assign n27309 = n2783 & ~n27307 ;
  assign n27310 = ~n27308 & n27309 ;
  assign n27306 = \P3_Address_reg[24]/NET0131  & ~n2782 ;
  assign n27311 = n21026 & n26536 ;
  assign n27312 = ~\P3_rEIP_reg[25]/NET0131  & ~n27311 ;
  assign n27313 = ~n26537 & n26540 ;
  assign n27314 = ~n27312 & n27313 ;
  assign n27315 = ~n27306 & ~n27314 ;
  assign n27316 = ~n27310 & n27315 ;
  assign n27318 = ~\P2_rEIP_reg[26]/NET0131  & ~n26603 ;
  assign n27319 = n1816 & ~n26604 ;
  assign n27320 = ~n27318 & n27319 ;
  assign n27317 = \P2_Address_reg[24]/NET0131  & ~n1815 ;
  assign n27321 = n16545 & n26576 ;
  assign n27322 = ~\P2_rEIP_reg[25]/NET0131  & ~n27321 ;
  assign n27323 = n26575 & ~n26577 ;
  assign n27324 = ~n27322 & n27323 ;
  assign n27325 = ~n27317 & ~n27324 ;
  assign n27326 = ~n27320 & n27325 ;
  assign n27332 = ~n19097 & n26642 ;
  assign n27331 = ~\P1_rEIP_reg[25]/NET0131  & ~n26642 ;
  assign n27333 = n26647 & ~n27331 ;
  assign n27334 = ~n27332 & n27333 ;
  assign n27327 = \address1[24]_pad  & ~n2307 ;
  assign n27328 = ~\P1_rEIP_reg[26]/NET0131  & ~n26633 ;
  assign n27329 = n2308 & ~n26634 ;
  assign n27330 = ~n27328 & n27329 ;
  assign n27335 = ~n27327 & ~n27330 ;
  assign n27336 = ~n27334 & n27335 ;
  assign n27338 = ~\P3_rEIP_reg[14]/NET0131  & ~n26556 ;
  assign n27339 = n2783 & ~n26557 ;
  assign n27340 = ~n27338 & n27339 ;
  assign n27337 = \P3_Address_reg[12]/NET0131  & ~n2782 ;
  assign n27341 = n20423 & n26534 ;
  assign n27342 = \P3_rEIP_reg[11]/NET0131  & n27341 ;
  assign n27343 = \P3_rEIP_reg[12]/NET0131  & n27342 ;
  assign n27345 = ~\P3_rEIP_reg[13]/NET0131  & ~n27343 ;
  assign n27344 = \P3_rEIP_reg[13]/NET0131  & n27343 ;
  assign n27346 = n26540 & ~n27344 ;
  assign n27347 = ~n27345 & n27346 ;
  assign n27348 = ~n27337 & ~n27347 ;
  assign n27349 = ~n27340 & n27348 ;
  assign n27351 = \P2_rEIP_reg[13]/NET0131  & n26595 ;
  assign n27353 = \P2_rEIP_reg[14]/NET0131  & n27351 ;
  assign n27352 = ~\P2_rEIP_reg[14]/NET0131  & ~n27351 ;
  assign n27354 = n1816 & ~n27352 ;
  assign n27355 = ~n27353 & n27354 ;
  assign n27350 = \P2_Address_reg[12]/NET0131  & ~n1815 ;
  assign n27356 = n16533 & n26576 ;
  assign n27358 = ~\P2_rEIP_reg[13]/NET0131  & ~n27356 ;
  assign n27357 = \P2_rEIP_reg[13]/NET0131  & n27356 ;
  assign n27359 = n26575 & ~n27357 ;
  assign n27360 = ~n27358 & n27359 ;
  assign n27361 = ~n27350 & ~n27360 ;
  assign n27362 = ~n27355 & n27361 ;
  assign n27364 = ~\P1_rEIP_reg[14]/NET0131  & ~n26628 ;
  assign n27365 = n2308 & ~n26629 ;
  assign n27366 = ~n27364 & n27365 ;
  assign n27363 = \address1[12]_pad  & ~n2307 ;
  assign n27369 = n18569 & n26642 ;
  assign n27367 = n18568 & n26642 ;
  assign n27368 = ~\P1_rEIP_reg[13]/NET0131  & ~n27367 ;
  assign n27370 = n26647 & ~n27368 ;
  assign n27371 = ~n27369 & n27370 ;
  assign n27372 = ~n27363 & ~n27371 ;
  assign n27373 = ~n27366 & n27372 ;
  assign n27376 = n2666 & n18209 ;
  assign n27375 = ~\P3_InstQueue_reg[0][0]/NET0131  & ~n18209 ;
  assign n27377 = n2994 & ~n27375 ;
  assign n27378 = ~n27376 & n27377 ;
  assign n27374 = \P3_InstQueue_reg[0][0]/NET0131  & ~n18218 ;
  assign n27379 = \buf2_reg[24]/NET0131  & n18200 ;
  assign n27380 = \buf2_reg[16]/NET0131  & n18203 ;
  assign n27381 = ~n27379 & ~n27380 ;
  assign n27382 = n2970 & ~n27381 ;
  assign n27383 = \buf2_reg[0]/NET0131  & n18228 ;
  assign n27384 = ~n27382 & ~n27383 ;
  assign n27385 = ~n27374 & n27384 ;
  assign n27386 = ~n27378 & n27385 ;
  assign n27389 = n2666 & n18246 ;
  assign n27388 = ~\P3_InstQueue_reg[10][0]/NET0131  & ~n18246 ;
  assign n27390 = n2994 & ~n27388 ;
  assign n27391 = ~n27389 & n27390 ;
  assign n27387 = \P3_InstQueue_reg[10][0]/NET0131  & ~n18243 ;
  assign n27392 = \buf2_reg[24]/NET0131  & n18233 ;
  assign n27393 = \buf2_reg[16]/NET0131  & n18236 ;
  assign n27394 = ~n27392 & ~n27393 ;
  assign n27395 = n2970 & ~n27394 ;
  assign n27396 = \buf2_reg[0]/NET0131  & n18255 ;
  assign n27397 = ~n27395 & ~n27396 ;
  assign n27398 = ~n27387 & n27397 ;
  assign n27399 = ~n27391 & n27398 ;
  assign n27402 = n2666 & n18284 ;
  assign n27401 = ~\P3_InstQueue_reg[12][0]/NET0131  & ~n18284 ;
  assign n27403 = n2994 & ~n27401 ;
  assign n27404 = ~n27402 & n27403 ;
  assign n27400 = \P3_InstQueue_reg[12][0]/NET0131  & ~n18287 ;
  assign n27405 = \buf2_reg[16]/NET0131  & n18246 ;
  assign n27406 = \buf2_reg[24]/NET0131  & n18271 ;
  assign n27407 = ~n27405 & ~n27406 ;
  assign n27408 = n2970 & ~n27407 ;
  assign n27409 = \buf2_reg[0]/NET0131  & n18297 ;
  assign n27410 = ~n27408 & ~n27409 ;
  assign n27411 = ~n27400 & n27410 ;
  assign n27412 = ~n27404 & n27411 ;
  assign n27420 = n2666 & n18200 ;
  assign n27419 = ~\P3_InstQueue_reg[13][0]/NET0131  & ~n18200 ;
  assign n27421 = n2994 & ~n27419 ;
  assign n27422 = ~n27420 & n27421 ;
  assign n27416 = ~\P3_InstQueue_reg[13][0]/NET0131  & n18302 ;
  assign n27415 = ~\buf2_reg[0]/NET0131  & ~n18302 ;
  assign n27417 = n18305 & ~n27415 ;
  assign n27418 = ~n27416 & n27417 ;
  assign n27413 = \P3_InstQueue_reg[13][0]/NET0131  & ~n18217 ;
  assign n27414 = n18303 & n27076 ;
  assign n27423 = ~n27413 & ~n27414 ;
  assign n27424 = ~n27418 & n27423 ;
  assign n27425 = ~n27422 & n27424 ;
  assign n27428 = n2666 & n18203 ;
  assign n27427 = ~\P3_InstQueue_reg[14][0]/NET0131  & ~n18203 ;
  assign n27429 = n2994 & ~n27427 ;
  assign n27430 = ~n27428 & n27429 ;
  assign n27426 = \P3_InstQueue_reg[14][0]/NET0131  & ~n18325 ;
  assign n27431 = \buf2_reg[24]/NET0131  & n18266 ;
  assign n27432 = \buf2_reg[16]/NET0131  & n18284 ;
  assign n27433 = ~n27431 & ~n27432 ;
  assign n27434 = n2970 & ~n27433 ;
  assign n27435 = \buf2_reg[0]/NET0131  & n18335 ;
  assign n27436 = ~n27434 & ~n27435 ;
  assign n27437 = ~n27426 & n27436 ;
  assign n27438 = ~n27430 & n27437 ;
  assign n27441 = n2666 & n18212 ;
  assign n27440 = ~\P3_InstQueue_reg[15][0]/NET0131  & ~n18212 ;
  assign n27442 = n2994 & ~n27440 ;
  assign n27443 = ~n27441 & n27442 ;
  assign n27439 = \P3_InstQueue_reg[15][0]/NET0131  & ~n18344 ;
  assign n27444 = \buf2_reg[24]/NET0131  & n18284 ;
  assign n27445 = \buf2_reg[16]/NET0131  & n18200 ;
  assign n27446 = ~n27444 & ~n27445 ;
  assign n27447 = n2970 & ~n27446 ;
  assign n27448 = \buf2_reg[0]/NET0131  & n18354 ;
  assign n27449 = ~n27447 & ~n27448 ;
  assign n27450 = ~n27439 & n27449 ;
  assign n27451 = ~n27443 & n27450 ;
  assign n27454 = n2666 & n18361 ;
  assign n27453 = ~\P3_InstQueue_reg[1][0]/NET0131  & ~n18361 ;
  assign n27455 = n2994 & ~n27453 ;
  assign n27456 = ~n27454 & n27455 ;
  assign n27452 = \P3_InstQueue_reg[1][0]/NET0131  & ~n18364 ;
  assign n27457 = \buf2_reg[24]/NET0131  & n18203 ;
  assign n27458 = \buf2_reg[16]/NET0131  & n18212 ;
  assign n27459 = ~n27457 & ~n27458 ;
  assign n27460 = n2970 & ~n27459 ;
  assign n27461 = \buf2_reg[0]/NET0131  & n18374 ;
  assign n27462 = ~n27460 & ~n27461 ;
  assign n27463 = ~n27452 & n27462 ;
  assign n27464 = ~n27456 & n27463 ;
  assign n27467 = n2666 & n18386 ;
  assign n27466 = ~\P3_InstQueue_reg[2][0]/NET0131  & ~n18386 ;
  assign n27468 = n2994 & ~n27466 ;
  assign n27469 = ~n27467 & n27468 ;
  assign n27465 = \P3_InstQueue_reg[2][0]/NET0131  & ~n18383 ;
  assign n27470 = \buf2_reg[24]/NET0131  & n18212 ;
  assign n27471 = \buf2_reg[16]/NET0131  & n18209 ;
  assign n27472 = ~n27470 & ~n27471 ;
  assign n27473 = n2970 & ~n27472 ;
  assign n27474 = \buf2_reg[0]/NET0131  & n18395 ;
  assign n27475 = ~n27473 & ~n27474 ;
  assign n27476 = ~n27465 & n27475 ;
  assign n27477 = ~n27469 & n27476 ;
  assign n27480 = n2666 & n18421 ;
  assign n27479 = ~\P3_InstQueue_reg[4][0]/NET0131  & ~n18421 ;
  assign n27481 = n2994 & ~n27479 ;
  assign n27482 = ~n27480 & n27481 ;
  assign n27478 = \P3_InstQueue_reg[4][0]/NET0131  & ~n18424 ;
  assign n27483 = \buf2_reg[16]/NET0131  & n18386 ;
  assign n27484 = \buf2_reg[24]/NET0131  & n18361 ;
  assign n27485 = ~n27483 & ~n27484 ;
  assign n27486 = n2970 & ~n27485 ;
  assign n27487 = \buf2_reg[0]/NET0131  & n18434 ;
  assign n27488 = ~n27486 & ~n27487 ;
  assign n27489 = ~n27478 & n27488 ;
  assign n27490 = ~n27482 & n27489 ;
  assign n27498 = n2666 & n18439 ;
  assign n27497 = ~\P3_InstQueue_reg[5][0]/NET0131  & ~n18439 ;
  assign n27499 = n2994 & ~n27497 ;
  assign n27500 = ~n27498 & n27499 ;
  assign n27494 = ~\P3_InstQueue_reg[5][0]/NET0131  & n18440 ;
  assign n27493 = ~\buf2_reg[0]/NET0131  & ~n18440 ;
  assign n27495 = n18443 & ~n27493 ;
  assign n27496 = ~n27494 & n27495 ;
  assign n27491 = \P3_InstQueue_reg[5][0]/NET0131  & ~n18217 ;
  assign n27492 = n18441 & n27076 ;
  assign n27501 = ~n27491 & ~n27492 ;
  assign n27502 = ~n27496 & n27501 ;
  assign n27503 = ~n27500 & n27502 ;
  assign n27506 = n2666 & n18462 ;
  assign n27505 = ~\P3_InstQueue_reg[6][0]/NET0131  & ~n18462 ;
  assign n27507 = n2994 & ~n27505 ;
  assign n27508 = ~n27506 & n27507 ;
  assign n27504 = \P3_InstQueue_reg[6][0]/NET0131  & ~n18465 ;
  assign n27509 = \buf2_reg[24]/NET0131  & n18405 ;
  assign n27510 = \buf2_reg[16]/NET0131  & n18421 ;
  assign n27511 = ~n27509 & ~n27510 ;
  assign n27512 = n2970 & ~n27511 ;
  assign n27513 = \buf2_reg[0]/NET0131  & n18475 ;
  assign n27514 = ~n27512 & ~n27513 ;
  assign n27515 = ~n27504 & n27514 ;
  assign n27516 = ~n27508 & n27515 ;
  assign n27519 = n2666 & n18236 ;
  assign n27518 = ~\P3_InstQueue_reg[8][0]/NET0131  & ~n18236 ;
  assign n27520 = n2994 & ~n27518 ;
  assign n27521 = ~n27519 & n27520 ;
  assign n27517 = \P3_InstQueue_reg[8][0]/NET0131  & ~n18502 ;
  assign n27522 = \buf2_reg[24]/NET0131  & n18439 ;
  assign n27523 = \buf2_reg[16]/NET0131  & n18462 ;
  assign n27524 = ~n27522 & ~n27523 ;
  assign n27525 = n2970 & ~n27524 ;
  assign n27526 = \buf2_reg[0]/NET0131  & n18512 ;
  assign n27527 = ~n27525 & ~n27526 ;
  assign n27528 = ~n27517 & n27527 ;
  assign n27529 = ~n27521 & n27528 ;
  assign n27543 = n2666 & n18271 ;
  assign n27542 = ~\P3_InstQueue_reg[9][0]/NET0131  & ~n18271 ;
  assign n27544 = n2994 & ~n27542 ;
  assign n27545 = ~n27543 & n27544 ;
  assign n27534 = \buf2_reg[24]/NET0131  & n18462 ;
  assign n27535 = \buf2_reg[16]/NET0131  & n18233 ;
  assign n27536 = ~n27534 & ~n27535 ;
  assign n27537 = \P3_DataWidth_reg[1]/NET0131  & ~n27536 ;
  assign n27530 = \P3_InstQueue_reg[9][0]/NET0131  & ~n18235 ;
  assign n27531 = \buf2_reg[0]/NET0131  & n18235 ;
  assign n27532 = ~n27530 & ~n27531 ;
  assign n27538 = ~n18525 & ~n27532 ;
  assign n27539 = ~n27537 & ~n27538 ;
  assign n27540 = n2959 & ~n27539 ;
  assign n27533 = n4415 & ~n27532 ;
  assign n27541 = \P3_InstQueue_reg[9][0]/NET0131  & ~n18217 ;
  assign n27546 = ~n27533 & ~n27541 ;
  assign n27547 = ~n27540 & n27546 ;
  assign n27548 = ~n27545 & n27547 ;
  assign n27550 = ~\P3_rEIP_reg[22]/NET0131  & ~n26561 ;
  assign n27551 = n2783 & ~n26562 ;
  assign n27552 = ~n27550 & n27551 ;
  assign n27549 = \P3_Address_reg[20]/NET0131  & ~n2782 ;
  assign n27553 = n20842 & n26928 ;
  assign n27555 = ~\P3_rEIP_reg[21]/NET0131  & ~n27553 ;
  assign n27554 = \P3_rEIP_reg[21]/NET0131  & n27553 ;
  assign n27556 = n26540 & ~n27554 ;
  assign n27557 = ~n27555 & n27556 ;
  assign n27558 = ~n27549 & ~n27557 ;
  assign n27559 = ~n27552 & n27558 ;
  assign n27561 = ~\P2_rEIP_reg[22]/NET0131  & ~n26599 ;
  assign n27562 = n1816 & ~n26600 ;
  assign n27563 = ~n27561 & n27562 ;
  assign n27560 = \P2_Address_reg[20]/NET0131  & ~n1815 ;
  assign n27567 = n16542 & n26576 ;
  assign n27564 = n16540 & n26576 ;
  assign n27565 = \P2_rEIP_reg[20]/NET0131  & n27564 ;
  assign n27566 = ~\P2_rEIP_reg[21]/NET0131  & ~n27565 ;
  assign n27568 = n26575 & ~n27566 ;
  assign n27569 = ~n27567 & n27568 ;
  assign n27570 = ~n27560 & ~n27569 ;
  assign n27571 = ~n27563 & n27570 ;
  assign n27573 = \P1_rEIP_reg[19]/NET0131  & n26951 ;
  assign n27574 = \P1_rEIP_reg[20]/NET0131  & n27573 ;
  assign n27575 = \P1_rEIP_reg[21]/NET0131  & n27574 ;
  assign n27577 = \P1_rEIP_reg[22]/NET0131  & n27575 ;
  assign n27576 = ~\P1_rEIP_reg[22]/NET0131  & ~n27575 ;
  assign n27578 = n2308 & ~n27576 ;
  assign n27579 = ~n27577 & n27578 ;
  assign n27572 = \address1[20]_pad  & ~n2307 ;
  assign n27580 = n18734 & n26642 ;
  assign n27581 = n18853 & n27580 ;
  assign n27583 = ~\P1_rEIP_reg[21]/NET0131  & ~n27581 ;
  assign n27582 = \P1_rEIP_reg[21]/NET0131  & n27581 ;
  assign n27584 = n26647 & ~n27582 ;
  assign n27585 = ~n27583 & n27584 ;
  assign n27586 = ~n27572 & ~n27585 ;
  assign n27587 = ~n27579 & n27586 ;
  assign n27593 = ~\P3_rEIP_reg[10]/NET0131  & ~n26552 ;
  assign n27594 = n2783 & ~n26553 ;
  assign n27595 = ~n27593 & n27594 ;
  assign n27588 = \P3_Address_reg[8]/NET0131  & ~n2782 ;
  assign n27590 = ~n21459 & n26534 ;
  assign n27589 = ~\P3_rEIP_reg[9]/NET0131  & ~n26534 ;
  assign n27591 = n26540 & ~n27589 ;
  assign n27592 = ~n27590 & n27591 ;
  assign n27596 = ~n27588 & ~n27592 ;
  assign n27597 = ~n27595 & n27596 ;
  assign n27603 = ~\P2_rEIP_reg[10]/NET0131  & ~n26592 ;
  assign n27604 = n1816 & ~n26593 ;
  assign n27605 = ~n27603 & n27604 ;
  assign n27598 = \P2_Address_reg[8]/NET0131  & ~n1815 ;
  assign n27600 = ~n20378 & n26576 ;
  assign n27599 = ~\P2_rEIP_reg[9]/NET0131  & ~n26576 ;
  assign n27601 = n26575 & ~n27599 ;
  assign n27602 = ~n27600 & n27601 ;
  assign n27606 = ~n27598 & ~n27602 ;
  assign n27607 = ~n27605 & n27606 ;
  assign n27616 = ~\P1_rEIP_reg[10]/NET0131  & ~n26624 ;
  assign n27617 = n2308 & ~n26625 ;
  assign n27618 = ~n27616 & n27617 ;
  assign n27608 = \address1[8]_pad  & ~n2307 ;
  assign n27609 = n18562 & n26642 ;
  assign n27610 = \P1_rEIP_reg[7]/NET0131  & n27609 ;
  assign n27611 = \P1_rEIP_reg[8]/NET0131  & n27610 ;
  assign n27613 = \P1_rEIP_reg[9]/NET0131  & n27611 ;
  assign n27612 = ~\P1_rEIP_reg[9]/NET0131  & ~n27611 ;
  assign n27614 = n26647 & ~n27612 ;
  assign n27615 = ~n27613 & n27614 ;
  assign n27619 = ~n27608 & ~n27615 ;
  assign n27620 = ~n27618 & n27619 ;
  assign n27622 = ~\P3_rEIP_reg[6]/NET0131  & ~n26548 ;
  assign n27623 = n2783 & ~n26549 ;
  assign n27624 = ~n27622 & n27623 ;
  assign n27621 = \P3_Address_reg[4]/NET0131  & ~n2782 ;
  assign n27625 = \P3_rEIP_reg[1]/NET0131  & n26534 ;
  assign n27626 = \P3_rEIP_reg[2]/NET0131  & n27625 ;
  assign n27627 = \P3_rEIP_reg[3]/NET0131  & n27626 ;
  assign n27628 = \P3_rEIP_reg[4]/NET0131  & n27627 ;
  assign n27629 = ~\P3_rEIP_reg[5]/NET0131  & ~n27628 ;
  assign n27630 = n20417 & n26534 ;
  assign n27631 = n26540 & ~n27630 ;
  assign n27632 = ~n27629 & n27631 ;
  assign n27633 = ~n27621 & ~n27632 ;
  assign n27634 = ~n27624 & n27633 ;
  assign n27636 = \P2_rEIP_reg[5]/NET0131  & n26589 ;
  assign n27638 = ~\P2_rEIP_reg[6]/NET0131  & ~n27636 ;
  assign n27637 = \P2_rEIP_reg[6]/NET0131  & n27636 ;
  assign n27639 = n1816 & ~n27637 ;
  assign n27640 = ~n27638 & n27639 ;
  assign n27635 = \P2_Address_reg[4]/NET0131  & ~n1815 ;
  assign n27641 = \P2_rEIP_reg[1]/NET0131  & n26576 ;
  assign n27642 = \P2_rEIP_reg[2]/NET0131  & n27641 ;
  assign n27643 = \P2_rEIP_reg[3]/NET0131  & n27642 ;
  assign n27644 = \P2_rEIP_reg[4]/NET0131  & n27643 ;
  assign n27646 = ~\P2_rEIP_reg[5]/NET0131  & ~n27644 ;
  assign n27645 = \P2_rEIP_reg[5]/NET0131  & n27644 ;
  assign n27647 = n26575 & ~n27645 ;
  assign n27648 = ~n27646 & n27647 ;
  assign n27649 = ~n27635 & ~n27648 ;
  assign n27650 = ~n27640 & n27649 ;
  assign n27652 = ~\P1_rEIP_reg[6]/NET0131  & ~n26620 ;
  assign n27653 = n2308 & ~n26621 ;
  assign n27654 = ~n27652 & n27653 ;
  assign n27651 = \address1[4]_pad  & ~n2307 ;
  assign n27655 = \P1_rEIP_reg[1]/NET0131  & n26642 ;
  assign n27656 = \P1_rEIP_reg[2]/NET0131  & n27655 ;
  assign n27657 = \P1_rEIP_reg[3]/NET0131  & n27656 ;
  assign n27658 = \P1_rEIP_reg[4]/NET0131  & n27657 ;
  assign n27660 = ~\P1_rEIP_reg[5]/NET0131  & ~n27658 ;
  assign n27659 = \P1_rEIP_reg[5]/NET0131  & n27658 ;
  assign n27661 = n26647 & ~n27659 ;
  assign n27662 = ~n27660 & n27661 ;
  assign n27663 = ~n27651 & ~n27662 ;
  assign n27664 = ~n27654 & n27663 ;
  assign n27672 = ~\P1_rEIP_reg[17]/NET0131  & ~n26631 ;
  assign n27673 = n2308 & ~n26632 ;
  assign n27674 = ~n27672 & n27673 ;
  assign n27665 = \address1[15]_pad  & ~n2307 ;
  assign n27666 = \P1_rEIP_reg[14]/NET0131  & n27369 ;
  assign n27667 = \P1_rEIP_reg[15]/NET0131  & n27666 ;
  assign n27669 = \P1_rEIP_reg[16]/NET0131  & n27667 ;
  assign n27668 = ~\P1_rEIP_reg[16]/NET0131  & ~n27667 ;
  assign n27670 = n26647 & ~n27668 ;
  assign n27671 = ~n27669 & n27670 ;
  assign n27675 = ~n27665 & ~n27671 ;
  assign n27676 = ~n27674 & n27675 ;
  assign n27678 = ~\P3_rEIP_reg[17]/NET0131  & ~n26559 ;
  assign n27679 = n2783 & ~n26922 ;
  assign n27680 = ~n27678 & n27679 ;
  assign n27677 = \P3_Address_reg[15]/NET0131  & ~n2782 ;
  assign n27681 = ~\P3_rEIP_reg[16]/NET0131  & ~n26927 ;
  assign n27682 = n26540 & ~n26928 ;
  assign n27683 = ~n27681 & n27682 ;
  assign n27684 = ~n27677 & ~n27683 ;
  assign n27685 = ~n27680 & n27684 ;
  assign n27687 = ~\P3_rEIP_reg[29]/NET0131  & ~n26566 ;
  assign n27688 = n2783 & ~n26567 ;
  assign n27689 = ~n27687 & n27688 ;
  assign n27686 = \P3_Address_reg[27]/NET0131  & ~n2782 ;
  assign n27690 = \P3_rEIP_reg[26]/NET0131  & n26537 ;
  assign n27691 = \P3_rEIP_reg[27]/NET0131  & n27690 ;
  assign n27692 = ~\P3_rEIP_reg[28]/NET0131  & ~n27691 ;
  assign n27693 = ~n26538 & n26540 ;
  assign n27694 = ~n27692 & n27693 ;
  assign n27695 = ~n27686 & ~n27694 ;
  assign n27696 = ~n27689 & n27695 ;
  assign n27703 = n16536 & n26595 ;
  assign n27704 = ~\P2_rEIP_reg[17]/NET0131  & ~n27703 ;
  assign n27705 = n1816 & ~n26940 ;
  assign n27706 = ~n27704 & n27705 ;
  assign n27697 = \P2_Address_reg[15]/NET0131  & ~n1815 ;
  assign n27699 = n16535 & n27356 ;
  assign n27700 = ~\P2_rEIP_reg[16]/NET0131  & ~n27699 ;
  assign n27698 = n16536 & n27356 ;
  assign n27701 = n26575 & ~n27698 ;
  assign n27702 = ~n27700 & n27701 ;
  assign n27707 = ~n27697 & ~n27702 ;
  assign n27708 = ~n27706 & n27707 ;
  assign n27710 = ~\P2_rEIP_reg[29]/NET0131  & ~n26606 ;
  assign n27711 = n1816 & ~n26607 ;
  assign n27712 = ~n27710 & n27711 ;
  assign n27709 = \P2_Address_reg[27]/NET0131  & ~n1815 ;
  assign n27713 = ~\P2_rEIP_reg[28]/NET0131  & ~n26579 ;
  assign n27714 = n26575 & ~n26580 ;
  assign n27715 = ~n27713 & n27714 ;
  assign n27716 = ~n27709 & ~n27715 ;
  assign n27717 = ~n27712 & n27716 ;
  assign n27719 = ~\P1_rEIP_reg[29]/NET0131  & ~n26636 ;
  assign n27720 = n2308 & ~n26637 ;
  assign n27721 = ~n27719 & n27720 ;
  assign n27718 = \address1[27]_pad  & ~n2307 ;
  assign n27722 = ~\P1_rEIP_reg[28]/NET0131  & ~n26644 ;
  assign n27723 = ~n26645 & n26647 ;
  assign n27724 = ~n27722 & n27723 ;
  assign n27725 = ~n27718 & ~n27724 ;
  assign n27726 = ~n27721 & n27725 ;
  assign n27728 = ~\P3_rEIP_reg[25]/NET0131  & ~n26564 ;
  assign n27729 = n2783 & ~n26565 ;
  assign n27730 = ~n27728 & n27729 ;
  assign n27727 = \P3_Address_reg[23]/NET0131  & ~n2782 ;
  assign n27731 = \P3_rEIP_reg[23]/NET0131  & n26536 ;
  assign n27732 = ~\P3_rEIP_reg[24]/NET0131  & ~n27731 ;
  assign n27733 = n26540 & ~n27311 ;
  assign n27734 = ~n27732 & n27733 ;
  assign n27735 = ~n27727 & ~n27734 ;
  assign n27736 = ~n27730 & n27735 ;
  assign n27738 = ~\P2_rEIP_reg[25]/NET0131  & ~n26602 ;
  assign n27739 = n1816 & ~n26603 ;
  assign n27740 = ~n27738 & n27739 ;
  assign n27737 = \P2_Address_reg[23]/NET0131  & ~n1815 ;
  assign n27741 = n16544 & n26576 ;
  assign n27742 = ~\P2_rEIP_reg[24]/NET0131  & ~n27741 ;
  assign n27743 = n26575 & ~n27321 ;
  assign n27744 = ~n27742 & n27743 ;
  assign n27745 = ~n27737 & ~n27744 ;
  assign n27746 = ~n27740 & n27745 ;
  assign n27753 = n19092 & n27574 ;
  assign n27754 = ~\P1_rEIP_reg[25]/NET0131  & ~n27753 ;
  assign n27755 = n2308 & ~n26633 ;
  assign n27756 = ~n27754 & n27755 ;
  assign n27747 = \address1[23]_pad  & ~n2307 ;
  assign n27748 = n18949 & n27581 ;
  assign n27750 = \P1_rEIP_reg[24]/NET0131  & n27748 ;
  assign n27749 = ~\P1_rEIP_reg[24]/NET0131  & ~n27748 ;
  assign n27751 = n26647 & ~n27749 ;
  assign n27752 = ~n27750 & n27751 ;
  assign n27757 = ~n27747 & ~n27752 ;
  assign n27758 = ~n27756 & n27757 ;
  assign n27760 = ~\P3_rEIP_reg[13]/NET0131  & ~n26555 ;
  assign n27761 = n2783 & ~n26556 ;
  assign n27762 = ~n27760 & n27761 ;
  assign n27759 = \P3_Address_reg[11]/NET0131  & ~n2782 ;
  assign n27763 = ~\P3_rEIP_reg[12]/NET0131  & ~n27342 ;
  assign n27764 = n26540 & ~n27343 ;
  assign n27765 = ~n27763 & n27764 ;
  assign n27766 = ~n27759 & ~n27765 ;
  assign n27767 = ~n27762 & n27766 ;
  assign n27773 = ~\P2_rEIP_reg[13]/NET0131  & ~n26595 ;
  assign n27774 = n1816 & ~n27351 ;
  assign n27775 = ~n27773 & n27774 ;
  assign n27768 = \P2_Address_reg[11]/NET0131  & ~n1815 ;
  assign n27770 = ~n19138 & n26576 ;
  assign n27769 = ~\P2_rEIP_reg[12]/NET0131  & ~n26576 ;
  assign n27771 = n26575 & ~n27769 ;
  assign n27772 = ~n27770 & n27771 ;
  assign n27776 = ~n27768 & ~n27772 ;
  assign n27777 = ~n27775 & n27776 ;
  assign n27783 = ~\P1_rEIP_reg[13]/NET0131  & ~n26627 ;
  assign n27784 = n2308 & ~n26628 ;
  assign n27785 = ~n27783 & n27784 ;
  assign n27778 = \address1[11]_pad  & ~n2307 ;
  assign n27780 = ~n21562 & n26642 ;
  assign n27779 = ~\P1_rEIP_reg[12]/NET0131  & ~n26642 ;
  assign n27781 = n26647 & ~n27779 ;
  assign n27782 = ~n27780 & n27781 ;
  assign n27786 = ~n27778 & ~n27782 ;
  assign n27787 = ~n27785 & n27786 ;
  assign n27789 = ~\P3_rEIP_reg[5]/NET0131  & ~n26547 ;
  assign n27790 = n2783 & ~n26548 ;
  assign n27791 = ~n27789 & n27790 ;
  assign n27788 = \P3_Address_reg[3]/NET0131  & ~n2782 ;
  assign n27792 = ~\P3_rEIP_reg[4]/NET0131  & ~n27627 ;
  assign n27793 = n26540 & ~n27628 ;
  assign n27794 = ~n27792 & n27793 ;
  assign n27795 = ~n27788 & ~n27794 ;
  assign n27796 = ~n27791 & n27795 ;
  assign n27798 = ~\P2_rEIP_reg[5]/NET0131  & ~n26589 ;
  assign n27799 = n1816 & ~n27636 ;
  assign n27800 = ~n27798 & n27799 ;
  assign n27797 = \P2_Address_reg[3]/NET0131  & ~n1815 ;
  assign n27801 = ~\P2_rEIP_reg[4]/NET0131  & ~n27643 ;
  assign n27802 = n26575 & ~n27644 ;
  assign n27803 = ~n27801 & n27802 ;
  assign n27804 = ~n27797 & ~n27803 ;
  assign n27805 = ~n27800 & n27804 ;
  assign n27807 = ~\P1_rEIP_reg[5]/NET0131  & ~n26619 ;
  assign n27808 = n2308 & ~n26620 ;
  assign n27809 = ~n27807 & n27808 ;
  assign n27806 = \address1[3]_pad  & ~n2307 ;
  assign n27810 = ~\P1_rEIP_reg[4]/NET0131  & ~n27657 ;
  assign n27811 = n26647 & ~n27658 ;
  assign n27812 = ~n27810 & n27811 ;
  assign n27813 = ~n27806 & ~n27812 ;
  assign n27814 = ~n27809 & n27813 ;
  assign n27816 = ~\P3_rEIP_reg[21]/NET0131  & ~n26560 ;
  assign n27817 = n2783 & ~n26561 ;
  assign n27818 = ~n27816 & n27817 ;
  assign n27815 = \P3_Address_reg[19]/NET0131  & ~n2782 ;
  assign n27819 = n20766 & n26534 ;
  assign n27820 = ~\P3_rEIP_reg[20]/NET0131  & ~n27819 ;
  assign n27821 = n26540 & ~n27553 ;
  assign n27822 = ~n27820 & n27821 ;
  assign n27823 = ~n27815 & ~n27822 ;
  assign n27824 = ~n27818 & n27823 ;
  assign n27826 = ~\P2_rEIP_reg[21]/NET0131  & ~n26598 ;
  assign n27827 = n1816 & ~n26599 ;
  assign n27828 = ~n27826 & n27827 ;
  assign n27825 = \P2_Address_reg[19]/NET0131  & ~n1815 ;
  assign n27829 = ~\P2_rEIP_reg[20]/NET0131  & ~n27564 ;
  assign n27830 = n26575 & ~n27565 ;
  assign n27831 = ~n27829 & n27830 ;
  assign n27832 = ~n27825 & ~n27831 ;
  assign n27833 = ~n27828 & n27832 ;
  assign n27835 = ~\P1_rEIP_reg[21]/NET0131  & ~n27574 ;
  assign n27836 = n2308 & ~n27575 ;
  assign n27837 = ~n27835 & n27836 ;
  assign n27834 = \address1[19]_pad  & ~n2307 ;
  assign n27838 = n18769 & n26642 ;
  assign n27839 = ~\P1_rEIP_reg[20]/NET0131  & ~n27838 ;
  assign n27840 = n26647 & ~n27581 ;
  assign n27841 = ~n27839 & n27840 ;
  assign n27842 = ~n27834 & ~n27841 ;
  assign n27843 = ~n27837 & n27842 ;
  assign n27849 = ~\P3_rEIP_reg[9]/NET0131  & ~n26551 ;
  assign n27850 = n2783 & ~n26552 ;
  assign n27851 = ~n27849 & n27850 ;
  assign n27844 = \P3_Address_reg[7]/NET0131  & ~n2782 ;
  assign n27846 = ~n21425 & n26534 ;
  assign n27845 = ~\P3_rEIP_reg[8]/NET0131  & ~n26534 ;
  assign n27847 = n26540 & ~n27845 ;
  assign n27848 = ~n27846 & n27847 ;
  assign n27852 = ~n27844 & ~n27848 ;
  assign n27853 = ~n27851 & n27852 ;
  assign n27859 = ~\P2_rEIP_reg[9]/NET0131  & ~n26591 ;
  assign n27860 = n1816 & ~n26592 ;
  assign n27861 = ~n27859 & n27860 ;
  assign n27854 = \P2_Address_reg[7]/NET0131  & ~n1815 ;
  assign n27856 = ~n20347 & n26576 ;
  assign n27855 = ~\P2_rEIP_reg[8]/NET0131  & ~n26576 ;
  assign n27857 = n26575 & ~n27855 ;
  assign n27858 = ~n27856 & n27857 ;
  assign n27862 = ~n27854 & ~n27858 ;
  assign n27863 = ~n27861 & n27862 ;
  assign n27865 = ~\P1_rEIP_reg[9]/NET0131  & ~n26623 ;
  assign n27866 = n2308 & ~n26624 ;
  assign n27867 = ~n27865 & n27866 ;
  assign n27864 = \address1[7]_pad  & ~n2307 ;
  assign n27868 = ~\P1_rEIP_reg[8]/NET0131  & ~n27610 ;
  assign n27869 = n26647 & ~n27611 ;
  assign n27870 = ~n27868 & n27869 ;
  assign n27871 = ~n27864 & ~n27870 ;
  assign n27872 = ~n27867 & n27871 ;
  assign n27875 = ~\P1_D_C_n_reg/NET0131  & \P1_M_IO_n_reg/NET0131  ;
  assign n27876 = \P1_W_R_n_reg/NET0131  & ~\ast1_pad  ;
  assign n27877 = n27875 & n27876 ;
  assign n27873 = ~\P1_BE_n_reg[0]/NET0131  & ~\P1_BE_n_reg[1]/NET0131  ;
  assign n27874 = ~\P1_BE_n_reg[2]/NET0131  & ~\P1_BE_n_reg[3]/NET0131  ;
  assign n27878 = n27873 & n27874 ;
  assign n27879 = n27877 & n27878 ;
  assign n27880 = n5137 & n27879 ;
  assign n27883 = ~\P2_BE_n_reg[3]/NET0131  & ~\P2_D_C_n_reg/NET0131  ;
  assign n27884 = \P2_M_IO_n_reg/NET0131  & \P2_W_R_n_reg/NET0131  ;
  assign n27885 = n27883 & n27884 ;
  assign n27881 = ~\P2_ADS_n_reg/NET0131  & ~\P2_BE_n_reg[0]/NET0131  ;
  assign n27882 = ~\P2_BE_n_reg[1]/NET0131  & ~\P2_BE_n_reg[2]/NET0131  ;
  assign n27886 = n27881 & n27882 ;
  assign n27887 = n27885 & n27886 ;
  assign n27888 = n3079 & n27887 ;
  assign n27889 = \buf1_reg[16]/NET0131  & ~n27888 ;
  assign n27890 = \P2_Datao_reg[16]/NET0131  & n27888 ;
  assign n27891 = ~n27889 & ~n27890 ;
  assign n27892 = ~n27880 & ~n27891 ;
  assign n27893 = \P1_Datao_reg[16]/NET0131  & n27880 ;
  assign n27894 = ~n27892 & ~n27893 ;
  assign n27895 = \buf1_reg[27]/NET0131  & ~n27888 ;
  assign n27896 = \P2_Datao_reg[27]/NET0131  & n27888 ;
  assign n27897 = ~n27895 & ~n27896 ;
  assign n27898 = ~n27880 & ~n27897 ;
  assign n27899 = \P1_Datao_reg[27]/NET0131  & n27880 ;
  assign n27900 = ~n27898 & ~n27899 ;
  assign n27901 = \buf1_reg[3]/NET0131  & ~n27888 ;
  assign n27902 = \P2_Datao_reg[3]/NET0131  & n27888 ;
  assign n27903 = ~n27901 & ~n27902 ;
  assign n27904 = ~n27880 & ~n27903 ;
  assign n27905 = \P1_Datao_reg[3]/NET0131  & n27880 ;
  assign n27906 = ~n27904 & ~n27905 ;
  assign n27907 = \buf1_reg[14]/NET0131  & ~n27888 ;
  assign n27908 = \P2_Datao_reg[14]/NET0131  & n27888 ;
  assign n27909 = ~n27907 & ~n27908 ;
  assign n27910 = ~n27880 & ~n27909 ;
  assign n27911 = \P1_Datao_reg[14]/NET0131  & n27880 ;
  assign n27912 = ~n27910 & ~n27911 ;
  assign n27913 = \buf1_reg[30]/NET0131  & ~n27888 ;
  assign n27914 = \P2_Datao_reg[30]/NET0131  & n27888 ;
  assign n27915 = ~n27913 & ~n27914 ;
  assign n27916 = ~n27880 & ~n27915 ;
  assign n27917 = \P1_Datao_reg[30]/NET0131  & n27880 ;
  assign n27918 = ~n27916 & ~n27917 ;
  assign n27919 = \buf1_reg[25]/NET0131  & ~n27888 ;
  assign n27920 = \P2_Datao_reg[25]/NET0131  & n27888 ;
  assign n27921 = ~n27919 & ~n27920 ;
  assign n27922 = ~n27880 & ~n27921 ;
  assign n27923 = \P1_Datao_reg[25]/NET0131  & n27880 ;
  assign n27924 = ~n27922 & ~n27923 ;
  assign n27925 = \buf1_reg[26]/NET0131  & ~n27888 ;
  assign n27926 = \P2_Datao_reg[26]/NET0131  & n27888 ;
  assign n27927 = ~n27925 & ~n27926 ;
  assign n27928 = ~n27880 & ~n27927 ;
  assign n27929 = \P1_Datao_reg[26]/NET0131  & n27880 ;
  assign n27930 = ~n27928 & ~n27929 ;
  assign n27931 = \buf1_reg[15]/NET0131  & ~n27888 ;
  assign n27932 = \P2_Datao_reg[15]/NET0131  & n27888 ;
  assign n27933 = ~n27931 & ~n27932 ;
  assign n27934 = ~n27880 & ~n27933 ;
  assign n27935 = \P1_Datao_reg[15]/NET0131  & n27880 ;
  assign n27936 = ~n27934 & ~n27935 ;
  assign n27937 = \buf1_reg[19]/NET0131  & ~n27888 ;
  assign n27938 = \P2_Datao_reg[19]/NET0131  & n27888 ;
  assign n27939 = ~n27937 & ~n27938 ;
  assign n27940 = ~n27880 & ~n27939 ;
  assign n27941 = \P1_Datao_reg[19]/NET0131  & n27880 ;
  assign n27942 = ~n27940 & ~n27941 ;
  assign n27943 = \buf1_reg[0]/NET0131  & ~n27888 ;
  assign n27944 = \P2_Datao_reg[0]/NET0131  & n27888 ;
  assign n27945 = ~n27943 & ~n27944 ;
  assign n27946 = ~n27880 & ~n27945 ;
  assign n27947 = \P1_Datao_reg[0]/NET0131  & n27880 ;
  assign n27948 = ~n27946 & ~n27947 ;
  assign n27949 = \buf1_reg[10]/NET0131  & ~n27888 ;
  assign n27950 = \P2_Datao_reg[10]/NET0131  & n27888 ;
  assign n27951 = ~n27949 & ~n27950 ;
  assign n27952 = ~n27880 & ~n27951 ;
  assign n27953 = \P1_Datao_reg[10]/NET0131  & n27880 ;
  assign n27954 = ~n27952 & ~n27953 ;
  assign n27955 = \buf1_reg[11]/NET0131  & ~n27888 ;
  assign n27956 = \P2_Datao_reg[11]/NET0131  & n27888 ;
  assign n27957 = ~n27955 & ~n27956 ;
  assign n27958 = ~n27880 & ~n27957 ;
  assign n27959 = \P1_Datao_reg[11]/NET0131  & n27880 ;
  assign n27960 = ~n27958 & ~n27959 ;
  assign n27961 = \buf1_reg[12]/NET0131  & ~n27888 ;
  assign n27962 = \P2_Datao_reg[12]/NET0131  & n27888 ;
  assign n27963 = ~n27961 & ~n27962 ;
  assign n27964 = ~n27880 & ~n27963 ;
  assign n27965 = \P1_Datao_reg[12]/NET0131  & n27880 ;
  assign n27966 = ~n27964 & ~n27965 ;
  assign n27967 = \buf1_reg[13]/NET0131  & ~n27888 ;
  assign n27968 = \P2_Datao_reg[13]/NET0131  & n27888 ;
  assign n27969 = ~n27967 & ~n27968 ;
  assign n27970 = ~n27880 & ~n27969 ;
  assign n27971 = \P1_Datao_reg[13]/NET0131  & n27880 ;
  assign n27972 = ~n27970 & ~n27971 ;
  assign n27973 = \buf1_reg[17]/NET0131  & ~n27888 ;
  assign n27974 = \P2_Datao_reg[17]/NET0131  & n27888 ;
  assign n27975 = ~n27973 & ~n27974 ;
  assign n27976 = ~n27880 & ~n27975 ;
  assign n27977 = \P1_Datao_reg[17]/NET0131  & n27880 ;
  assign n27978 = ~n27976 & ~n27977 ;
  assign n27979 = \buf1_reg[1]/NET0131  & ~n27888 ;
  assign n27980 = \P2_Datao_reg[1]/NET0131  & n27888 ;
  assign n27981 = ~n27979 & ~n27980 ;
  assign n27982 = ~n27880 & ~n27981 ;
  assign n27983 = \P1_Datao_reg[1]/NET0131  & n27880 ;
  assign n27984 = ~n27982 & ~n27983 ;
  assign n27985 = \buf1_reg[20]/NET0131  & ~n27888 ;
  assign n27986 = \P2_Datao_reg[20]/NET0131  & n27888 ;
  assign n27987 = ~n27985 & ~n27986 ;
  assign n27988 = ~n27880 & ~n27987 ;
  assign n27989 = \P1_Datao_reg[20]/NET0131  & n27880 ;
  assign n27990 = ~n27988 & ~n27989 ;
  assign n27991 = \buf1_reg[21]/NET0131  & ~n27888 ;
  assign n27992 = \P2_Datao_reg[21]/NET0131  & n27888 ;
  assign n27993 = ~n27991 & ~n27992 ;
  assign n27994 = ~n27880 & ~n27993 ;
  assign n27995 = \P1_Datao_reg[21]/NET0131  & n27880 ;
  assign n27996 = ~n27994 & ~n27995 ;
  assign n27997 = \buf1_reg[22]/NET0131  & ~n27888 ;
  assign n27998 = \P2_Datao_reg[22]/NET0131  & n27888 ;
  assign n27999 = ~n27997 & ~n27998 ;
  assign n28000 = ~n27880 & ~n27999 ;
  assign n28001 = \P1_Datao_reg[22]/NET0131  & n27880 ;
  assign n28002 = ~n28000 & ~n28001 ;
  assign n28003 = \buf1_reg[23]/NET0131  & ~n27888 ;
  assign n28004 = \P2_Datao_reg[23]/NET0131  & n27888 ;
  assign n28005 = ~n28003 & ~n28004 ;
  assign n28006 = ~n27880 & ~n28005 ;
  assign n28007 = \P1_Datao_reg[23]/NET0131  & n27880 ;
  assign n28008 = ~n28006 & ~n28007 ;
  assign n28009 = \buf1_reg[24]/NET0131  & ~n27888 ;
  assign n28010 = \P2_Datao_reg[24]/NET0131  & n27888 ;
  assign n28011 = ~n28009 & ~n28010 ;
  assign n28012 = ~n27880 & ~n28011 ;
  assign n28013 = \P1_Datao_reg[24]/NET0131  & n27880 ;
  assign n28014 = ~n28012 & ~n28013 ;
  assign n28015 = \buf1_reg[28]/NET0131  & ~n27888 ;
  assign n28016 = \P2_Datao_reg[28]/NET0131  & n27888 ;
  assign n28017 = ~n28015 & ~n28016 ;
  assign n28018 = ~n27880 & ~n28017 ;
  assign n28019 = \P1_Datao_reg[28]/NET0131  & n27880 ;
  assign n28020 = ~n28018 & ~n28019 ;
  assign n28021 = \buf1_reg[2]/NET0131  & ~n27888 ;
  assign n28022 = \P2_Datao_reg[2]/NET0131  & n27888 ;
  assign n28023 = ~n28021 & ~n28022 ;
  assign n28024 = ~n27880 & ~n28023 ;
  assign n28025 = \P1_Datao_reg[2]/NET0131  & n27880 ;
  assign n28026 = ~n28024 & ~n28025 ;
  assign n28027 = \buf1_reg[4]/NET0131  & ~n27888 ;
  assign n28028 = \P2_Datao_reg[4]/NET0131  & n27888 ;
  assign n28029 = ~n28027 & ~n28028 ;
  assign n28030 = ~n27880 & ~n28029 ;
  assign n28031 = \P1_Datao_reg[4]/NET0131  & n27880 ;
  assign n28032 = ~n28030 & ~n28031 ;
  assign n28033 = \buf1_reg[6]/NET0131  & ~n27888 ;
  assign n28034 = \P2_Datao_reg[6]/NET0131  & n27888 ;
  assign n28035 = ~n28033 & ~n28034 ;
  assign n28036 = ~n27880 & ~n28035 ;
  assign n28037 = \P1_Datao_reg[6]/NET0131  & n27880 ;
  assign n28038 = ~n28036 & ~n28037 ;
  assign n28039 = \buf1_reg[9]/NET0131  & ~n27888 ;
  assign n28040 = \P2_Datao_reg[9]/NET0131  & n27888 ;
  assign n28041 = ~n28039 & ~n28040 ;
  assign n28042 = ~n27880 & ~n28041 ;
  assign n28043 = \P1_Datao_reg[9]/NET0131  & n27880 ;
  assign n28044 = ~n28042 & ~n28043 ;
  assign n28045 = \buf1_reg[29]/NET0131  & ~n27888 ;
  assign n28046 = \P2_Datao_reg[29]/NET0131  & n27888 ;
  assign n28047 = ~n28045 & ~n28046 ;
  assign n28048 = ~n27880 & ~n28047 ;
  assign n28049 = \P1_Datao_reg[29]/NET0131  & n27880 ;
  assign n28050 = ~n28048 & ~n28049 ;
  assign n28051 = \buf1_reg[18]/NET0131  & ~n27888 ;
  assign n28052 = \P2_Datao_reg[18]/NET0131  & n27888 ;
  assign n28053 = ~n28051 & ~n28052 ;
  assign n28054 = ~n27880 & ~n28053 ;
  assign n28055 = \P1_Datao_reg[18]/NET0131  & n27880 ;
  assign n28056 = ~n28054 & ~n28055 ;
  assign n28057 = \buf1_reg[7]/NET0131  & ~n27888 ;
  assign n28058 = \P2_Datao_reg[7]/NET0131  & n27888 ;
  assign n28059 = ~n28057 & ~n28058 ;
  assign n28060 = ~n27880 & ~n28059 ;
  assign n28061 = \P1_Datao_reg[7]/NET0131  & n27880 ;
  assign n28062 = ~n28060 & ~n28061 ;
  assign n28063 = \buf1_reg[8]/NET0131  & ~n27888 ;
  assign n28064 = \P2_Datao_reg[8]/NET0131  & n27888 ;
  assign n28065 = ~n28063 & ~n28064 ;
  assign n28066 = ~n27880 & ~n28065 ;
  assign n28067 = \P1_Datao_reg[8]/NET0131  & n27880 ;
  assign n28068 = ~n28066 & ~n28067 ;
  assign n28069 = \buf1_reg[5]/NET0131  & ~n27888 ;
  assign n28070 = \P2_Datao_reg[5]/NET0131  & n27888 ;
  assign n28071 = ~n28069 & ~n28070 ;
  assign n28072 = ~n27880 & ~n28071 ;
  assign n28073 = \P1_Datao_reg[5]/NET0131  & n27880 ;
  assign n28074 = ~n28072 & ~n28073 ;
  assign n28076 = ~\P3_rEIP_reg[16]/NET0131  & ~n26558 ;
  assign n28077 = n2783 & ~n26559 ;
  assign n28078 = ~n28076 & n28077 ;
  assign n28075 = \P3_Address_reg[14]/NET0131  & ~n2782 ;
  assign n28079 = ~\P3_rEIP_reg[15]/NET0131  & ~n26926 ;
  assign n28080 = n26540 & ~n26927 ;
  assign n28081 = ~n28079 & n28080 ;
  assign n28082 = ~n28075 & ~n28081 ;
  assign n28083 = ~n28078 & n28082 ;
  assign n28085 = \P2_rEIP_reg[15]/NET0131  & n27353 ;
  assign n28086 = ~\P2_rEIP_reg[16]/NET0131  & ~n28085 ;
  assign n28087 = n1816 & ~n27703 ;
  assign n28088 = ~n28086 & n28087 ;
  assign n28084 = \P2_Address_reg[14]/NET0131  & ~n1815 ;
  assign n28089 = n16534 & n27356 ;
  assign n28090 = ~\P2_rEIP_reg[15]/NET0131  & ~n28089 ;
  assign n28091 = n26575 & ~n27699 ;
  assign n28092 = ~n28090 & n28091 ;
  assign n28093 = ~n28084 & ~n28092 ;
  assign n28094 = ~n28088 & n28093 ;
  assign n28096 = ~\P1_rEIP_reg[16]/NET0131  & ~n26630 ;
  assign n28097 = n2308 & ~n26631 ;
  assign n28098 = ~n28096 & n28097 ;
  assign n28095 = \address1[14]_pad  & ~n2307 ;
  assign n28099 = ~\P1_rEIP_reg[15]/NET0131  & ~n27666 ;
  assign n28100 = n26647 & ~n27667 ;
  assign n28101 = ~n28099 & n28100 ;
  assign n28102 = ~n28095 & ~n28101 ;
  assign n28103 = ~n28098 & n28102 ;
  assign n28105 = ~\P1_rEIP_reg[28]/NET0131  & ~n26635 ;
  assign n28106 = n2308 & ~n26636 ;
  assign n28107 = ~n28105 & n28106 ;
  assign n28104 = \address1[26]_pad  & ~n2307 ;
  assign n28108 = ~\P1_rEIP_reg[27]/NET0131  & ~n26643 ;
  assign n28109 = ~n26644 & n26647 ;
  assign n28110 = ~n28108 & n28109 ;
  assign n28111 = ~n28104 & ~n28110 ;
  assign n28112 = ~n28107 & n28111 ;
  assign n28114 = \P3_rEIP_reg[27]/NET0131  & n27308 ;
  assign n28115 = ~\P3_rEIP_reg[28]/NET0131  & ~n28114 ;
  assign n28116 = n2783 & ~n26566 ;
  assign n28117 = ~n28115 & n28116 ;
  assign n28113 = \P3_Address_reg[26]/NET0131  & ~n2782 ;
  assign n28118 = ~\P3_rEIP_reg[27]/NET0131  & ~n27690 ;
  assign n28119 = n26540 & ~n27691 ;
  assign n28120 = ~n28118 & n28119 ;
  assign n28121 = ~n28113 & ~n28120 ;
  assign n28122 = ~n28117 & n28121 ;
  assign n28124 = ~\P2_rEIP_reg[28]/NET0131  & ~n26605 ;
  assign n28125 = n1816 & ~n26606 ;
  assign n28126 = ~n28124 & n28125 ;
  assign n28123 = \P2_Address_reg[26]/NET0131  & ~n1815 ;
  assign n28127 = ~\P2_rEIP_reg[27]/NET0131  & ~n26578 ;
  assign n28128 = n26575 & ~n26579 ;
  assign n28129 = ~n28127 & n28128 ;
  assign n28130 = ~n28123 & ~n28129 ;
  assign n28131 = ~n28126 & n28130 ;
  assign n28133 = ~\P3_rEIP_reg[24]/NET0131  & ~n26563 ;
  assign n28134 = n2783 & ~n26564 ;
  assign n28135 = ~n28133 & n28134 ;
  assign n28132 = \P3_Address_reg[22]/NET0131  & ~n2782 ;
  assign n28136 = ~\P3_rEIP_reg[23]/NET0131  & ~n26536 ;
  assign n28137 = n26540 & ~n27731 ;
  assign n28138 = ~n28136 & n28137 ;
  assign n28139 = ~n28132 & ~n28138 ;
  assign n28140 = ~n28135 & n28139 ;
  assign n28142 = ~\P2_rEIP_reg[24]/NET0131  & ~n26601 ;
  assign n28143 = n1816 & ~n26602 ;
  assign n28144 = ~n28142 & n28143 ;
  assign n28141 = \P2_Address_reg[22]/NET0131  & ~n1815 ;
  assign n28145 = n16543 & n26576 ;
  assign n28146 = ~\P2_rEIP_reg[23]/NET0131  & ~n28145 ;
  assign n28147 = n26575 & ~n27741 ;
  assign n28148 = ~n28146 & n28147 ;
  assign n28149 = ~n28141 & ~n28148 ;
  assign n28150 = ~n28144 & n28149 ;
  assign n28152 = n18949 & n27574 ;
  assign n28153 = ~\P1_rEIP_reg[24]/NET0131  & ~n28152 ;
  assign n28154 = n2308 & ~n27753 ;
  assign n28155 = ~n28153 & n28154 ;
  assign n28151 = \address1[22]_pad  & ~n2307 ;
  assign n28156 = \P1_rEIP_reg[22]/NET0131  & n27582 ;
  assign n28157 = ~\P1_rEIP_reg[23]/NET0131  & ~n28156 ;
  assign n28158 = n26647 & ~n27748 ;
  assign n28159 = ~n28157 & n28158 ;
  assign n28160 = ~n28151 & ~n28159 ;
  assign n28161 = ~n28155 & n28160 ;
  assign n28163 = ~\P3_rEIP_reg[12]/NET0131  & ~n26554 ;
  assign n28164 = n2783 & ~n26555 ;
  assign n28165 = ~n28163 & n28164 ;
  assign n28162 = \P3_Address_reg[10]/NET0131  & ~n2782 ;
  assign n28166 = ~\P3_rEIP_reg[11]/NET0131  & ~n27341 ;
  assign n28167 = n26540 & ~n27342 ;
  assign n28168 = ~n28166 & n28167 ;
  assign n28169 = ~n28162 & ~n28168 ;
  assign n28170 = ~n28165 & n28169 ;
  assign n28176 = ~\P2_rEIP_reg[12]/NET0131  & ~n26594 ;
  assign n28177 = n1816 & ~n26595 ;
  assign n28178 = ~n28176 & n28177 ;
  assign n28171 = \P2_Address_reg[10]/NET0131  & ~n1815 ;
  assign n28173 = ~n19068 & n26576 ;
  assign n28172 = ~\P2_rEIP_reg[11]/NET0131  & ~n26576 ;
  assign n28174 = n26575 & ~n28172 ;
  assign n28175 = ~n28173 & n28174 ;
  assign n28179 = ~n28171 & ~n28175 ;
  assign n28180 = ~n28178 & n28179 ;
  assign n28186 = ~\P1_rEIP_reg[12]/NET0131  & ~n26626 ;
  assign n28187 = n2308 & ~n26627 ;
  assign n28188 = ~n28186 & n28187 ;
  assign n28181 = \address1[10]_pad  & ~n2307 ;
  assign n28183 = ~n21528 & n26642 ;
  assign n28182 = ~\P1_rEIP_reg[11]/NET0131  & ~n26642 ;
  assign n28184 = n26647 & ~n28182 ;
  assign n28185 = ~n28183 & n28184 ;
  assign n28189 = ~n28181 & ~n28185 ;
  assign n28190 = ~n28188 & n28189 ;
  assign n28191 = ~n27880 & n27888 ;
  assign n28193 = ~\P3_rEIP_reg[4]/NET0131  & ~n26546 ;
  assign n28194 = n2783 & ~n26547 ;
  assign n28195 = ~n28193 & n28194 ;
  assign n28192 = \P3_Address_reg[2]/NET0131  & ~n2782 ;
  assign n28196 = ~\P3_rEIP_reg[3]/NET0131  & ~n27626 ;
  assign n28197 = n26540 & ~n27627 ;
  assign n28198 = ~n28196 & n28197 ;
  assign n28199 = ~n28192 & ~n28198 ;
  assign n28200 = ~n28195 & n28199 ;
  assign n28202 = ~\P2_rEIP_reg[4]/NET0131  & ~n26588 ;
  assign n28203 = n1816 & ~n26589 ;
  assign n28204 = ~n28202 & n28203 ;
  assign n28201 = \P2_Address_reg[2]/NET0131  & ~n1815 ;
  assign n28205 = ~\P2_rEIP_reg[3]/NET0131  & ~n27642 ;
  assign n28206 = n26575 & ~n27643 ;
  assign n28207 = ~n28205 & n28206 ;
  assign n28208 = ~n28201 & ~n28207 ;
  assign n28209 = ~n28204 & n28208 ;
  assign n28211 = ~\P1_rEIP_reg[4]/NET0131  & ~n26618 ;
  assign n28212 = n2308 & ~n26619 ;
  assign n28213 = ~n28211 & n28212 ;
  assign n28210 = \address1[2]_pad  & ~n2307 ;
  assign n28214 = ~\P1_rEIP_reg[3]/NET0131  & ~n27656 ;
  assign n28215 = n26647 & ~n27657 ;
  assign n28216 = ~n28214 & n28215 ;
  assign n28217 = ~n28210 & ~n28216 ;
  assign n28218 = ~n28213 & n28217 ;
  assign n28224 = n20728 & n26534 ;
  assign n28225 = ~\P3_rEIP_reg[19]/NET0131  & ~n28224 ;
  assign n28226 = n26540 & ~n27819 ;
  assign n28227 = ~n28225 & n28226 ;
  assign n28219 = \P3_Address_reg[18]/NET0131  & ~n2782 ;
  assign n28220 = n20841 & n26559 ;
  assign n28221 = ~\P3_rEIP_reg[20]/NET0131  & ~n28220 ;
  assign n28222 = n2783 & ~n26560 ;
  assign n28223 = ~n28221 & n28222 ;
  assign n28228 = ~n28219 & ~n28223 ;
  assign n28229 = ~n28227 & n28228 ;
  assign n28235 = ~\P2_rEIP_reg[20]/NET0131  & ~n26597 ;
  assign n28236 = n1816 & ~n26598 ;
  assign n28237 = ~n28235 & n28236 ;
  assign n28230 = \P2_Address_reg[18]/NET0131  & ~n1815 ;
  assign n28232 = ~n19501 & n26576 ;
  assign n28231 = ~\P2_rEIP_reg[19]/NET0131  & ~n26576 ;
  assign n28233 = n26575 & ~n28231 ;
  assign n28234 = ~n28232 & n28233 ;
  assign n28238 = ~n28230 & ~n28234 ;
  assign n28239 = ~n28237 & n28238 ;
  assign n28241 = ~\P1_rEIP_reg[20]/NET0131  & ~n27573 ;
  assign n28242 = n2308 & ~n27574 ;
  assign n28243 = ~n28241 & n28242 ;
  assign n28240 = \address1[18]_pad  & ~n2307 ;
  assign n28244 = ~\P1_rEIP_reg[19]/NET0131  & ~n27580 ;
  assign n28245 = n26647 & ~n27838 ;
  assign n28246 = ~n28244 & n28245 ;
  assign n28247 = ~n28240 & ~n28246 ;
  assign n28248 = ~n28243 & n28247 ;
  assign n28255 = ~\P3_rEIP_reg[8]/NET0131  & ~n26550 ;
  assign n28256 = n2783 & ~n26551 ;
  assign n28257 = ~n28255 & n28256 ;
  assign n28249 = \P3_Address_reg[6]/NET0131  & ~n2782 ;
  assign n28250 = \P3_rEIP_reg[6]/NET0131  & n27630 ;
  assign n28252 = \P3_rEIP_reg[7]/NET0131  & n28250 ;
  assign n28251 = ~\P3_rEIP_reg[7]/NET0131  & ~n28250 ;
  assign n28253 = n26540 & ~n28251 ;
  assign n28254 = ~n28252 & n28253 ;
  assign n28258 = ~n28249 & ~n28254 ;
  assign n28259 = ~n28257 & n28258 ;
  assign n28265 = ~\P2_rEIP_reg[8]/NET0131  & ~n26590 ;
  assign n28266 = n1816 & ~n26591 ;
  assign n28267 = ~n28265 & n28266 ;
  assign n28260 = \P2_Address_reg[6]/NET0131  & ~n1815 ;
  assign n28262 = ~n20277 & n26576 ;
  assign n28261 = ~\P2_rEIP_reg[7]/NET0131  & ~n26576 ;
  assign n28263 = n26575 & ~n28261 ;
  assign n28264 = ~n28262 & n28263 ;
  assign n28268 = ~n28260 & ~n28264 ;
  assign n28269 = ~n28267 & n28268 ;
  assign n28271 = ~\P1_rEIP_reg[8]/NET0131  & ~n26622 ;
  assign n28272 = n2308 & ~n26623 ;
  assign n28273 = ~n28271 & n28272 ;
  assign n28270 = \address1[6]_pad  & ~n2307 ;
  assign n28274 = ~\P1_rEIP_reg[7]/NET0131  & ~n27609 ;
  assign n28275 = n26647 & ~n27610 ;
  assign n28276 = ~n28274 & n28275 ;
  assign n28277 = ~n28270 & ~n28276 ;
  assign n28278 = ~n28273 & n28277 ;
  assign n28280 = ~\P3_rEIP_reg[27]/NET0131  & ~n27308 ;
  assign n28281 = n2783 & ~n28114 ;
  assign n28282 = ~n28280 & n28281 ;
  assign n28279 = \P3_Address_reg[25]/NET0131  & ~n2782 ;
  assign n28283 = ~\P3_rEIP_reg[26]/NET0131  & ~n26537 ;
  assign n28284 = n26540 & ~n27690 ;
  assign n28285 = ~n28283 & n28284 ;
  assign n28286 = ~n28279 & ~n28285 ;
  assign n28287 = ~n28282 & n28286 ;
  assign n28289 = ~\P2_rEIP_reg[27]/NET0131  & ~n26604 ;
  assign n28290 = n1816 & ~n26605 ;
  assign n28291 = ~n28289 & n28290 ;
  assign n28288 = \P2_Address_reg[25]/NET0131  & ~n1815 ;
  assign n28292 = ~\P2_rEIP_reg[26]/NET0131  & ~n26577 ;
  assign n28293 = n26575 & ~n26578 ;
  assign n28294 = ~n28292 & n28293 ;
  assign n28295 = ~n28288 & ~n28294 ;
  assign n28296 = ~n28291 & n28295 ;
  assign n28298 = ~\P1_rEIP_reg[27]/NET0131  & ~n26634 ;
  assign n28299 = n2308 & ~n26635 ;
  assign n28300 = ~n28298 & n28299 ;
  assign n28297 = \address1[25]_pad  & ~n2307 ;
  assign n28301 = n19096 & n26642 ;
  assign n28302 = ~\P1_rEIP_reg[26]/NET0131  & ~n28301 ;
  assign n28303 = ~n26643 & n26647 ;
  assign n28304 = ~n28302 & n28303 ;
  assign n28305 = ~n28297 & ~n28304 ;
  assign n28306 = ~n28300 & n28305 ;
  assign n28313 = \P3_rEIP_reg[31]/NET0131  & n26569 ;
  assign n28312 = ~\P3_rEIP_reg[31]/NET0131  & ~n26569 ;
  assign n28314 = n2783 & ~n28312 ;
  assign n28315 = ~n28313 & n28314 ;
  assign n28307 = \P3_Address_reg[29]/NET0131  & ~n2782 ;
  assign n28309 = ~n22221 & n26534 ;
  assign n28308 = ~\P3_rEIP_reg[30]/NET0131  & ~n26534 ;
  assign n28310 = n26540 & ~n28308 ;
  assign n28311 = ~n28309 & n28310 ;
  assign n28316 = ~n28307 & ~n28311 ;
  assign n28317 = ~n28315 & n28316 ;
  assign n28324 = \P2_rEIP_reg[31]/NET0131  & n26609 ;
  assign n28323 = ~\P2_rEIP_reg[31]/NET0131  & ~n26609 ;
  assign n28325 = n1816 & ~n28323 ;
  assign n28326 = ~n28324 & n28325 ;
  assign n28318 = \P2_Address_reg[29]/NET0131  & ~n1815 ;
  assign n28320 = ~n22130 & n26576 ;
  assign n28319 = ~\P2_rEIP_reg[30]/NET0131  & ~n26576 ;
  assign n28321 = n26575 & ~n28319 ;
  assign n28322 = ~n28320 & n28321 ;
  assign n28327 = ~n28318 & ~n28322 ;
  assign n28328 = ~n28326 & n28327 ;
  assign n28335 = \P1_rEIP_reg[31]/NET0131  & n26639 ;
  assign n28334 = ~\P1_rEIP_reg[31]/NET0131  & ~n26639 ;
  assign n28336 = n2308 & ~n28334 ;
  assign n28337 = ~n28335 & n28336 ;
  assign n28329 = \address1[29]_pad  & ~n2307 ;
  assign n28331 = \P1_rEIP_reg[30]/NET0131  & n26648 ;
  assign n28330 = ~\P1_rEIP_reg[30]/NET0131  & ~n26648 ;
  assign n28332 = n26647 & ~n28330 ;
  assign n28333 = ~n28331 & n28332 ;
  assign n28338 = ~n28329 & ~n28333 ;
  assign n28339 = ~n28337 & n28338 ;
  assign n28342 = \P2_State_reg[1]/NET0131  & hold_pad ;
  assign n28343 = ~\P2_RequestPending_reg/NET0131  & ~n28342 ;
  assign n28344 = ~\P2_State_reg[2]/NET0131  & ~n28343 ;
  assign n28340 = \P2_State_reg[1]/NET0131  & n1805 ;
  assign n28345 = \P2_RequestPending_reg/NET0131  & ~hold_pad ;
  assign n28346 = ~n28340 & ~n28345 ;
  assign n28347 = ~n28344 & n28346 ;
  assign n28348 = \P2_State_reg[0]/NET0131  & ~n28347 ;
  assign n28341 = \P2_State_reg[2]/NET0131  & n28340 ;
  assign n28349 = n1819 & ~n28341 ;
  assign n28350 = ~n28348 & n28349 ;
  assign n28353 = \P3_State_reg[1]/NET0131  & hold_pad ;
  assign n28354 = ~\P3_RequestPending_reg/NET0131  & ~n28353 ;
  assign n28355 = ~\P3_State_reg[2]/NET0131  & ~n28354 ;
  assign n28351 = \P3_State_reg[1]/NET0131  & n2835 ;
  assign n28356 = \P3_RequestPending_reg/NET0131  & ~hold_pad ;
  assign n28357 = ~n28351 & ~n28356 ;
  assign n28358 = ~n28355 & n28357 ;
  assign n28359 = \P3_State_reg[0]/NET0131  & ~n28358 ;
  assign n28352 = \P3_State_reg[2]/NET0131  & n28351 ;
  assign n28360 = n2786 & ~n28352 ;
  assign n28361 = ~n28359 & n28360 ;
  assign n28366 = ~\P1_State_reg[2]/NET0131  & hold_pad ;
  assign n28367 = ~n2317 & ~n28366 ;
  assign n28365 = ~\P1_State_reg[0]/NET0131  & ~\P1_State_reg[2]/NET0131  ;
  assign n28368 = \P1_State_reg[1]/NET0131  & ~n28365 ;
  assign n28369 = ~n28367 & n28368 ;
  assign n28362 = \P1_State_reg[2]/NET0131  & hold_pad ;
  assign n28363 = \P1_RequestPending_reg/NET0131  & \P1_State_reg[0]/NET0131  ;
  assign n28364 = ~n28362 & n28363 ;
  assign n28370 = n2311 & ~n28364 ;
  assign n28371 = ~n28369 & n28370 ;
  assign n28372 = \P2_State_reg[0]/NET0131  & ~n1805 ;
  assign n28373 = ~\P2_State_reg[0]/NET0131  & na_pad ;
  assign n28374 = \P2_State_reg[2]/NET0131  & ~n28373 ;
  assign n28375 = ~n28372 & ~n28374 ;
  assign n28376 = ~hold_pad & ~n28375 ;
  assign n28377 = \P2_State_reg[0]/NET0131  & ~\P2_State_reg[1]/NET0131  ;
  assign n28378 = ~\P2_State_reg[2]/NET0131  & n28377 ;
  assign n28379 = ~n28376 & ~n28378 ;
  assign n28380 = \P2_RequestPending_reg/NET0131  & ~n28379 ;
  assign n28381 = ~n26575 & ~n28380 ;
  assign n28382 = ~\P3_RequestPending_reg/NET0131  & ~\P3_State_reg[1]/NET0131  ;
  assign n28383 = ~\P3_State_reg[2]/NET0131  & ~n28382 ;
  assign n28384 = \P3_State_reg[0]/NET0131  & ~n28383 ;
  assign n28385 = ~n28356 & n28384 ;
  assign n28386 = ~n2835 & n28356 ;
  assign n28387 = \P3_State_reg[1]/NET0131  & ~n28386 ;
  assign n28388 = \P3_State_reg[0]/NET0131  & ~n28387 ;
  assign n28389 = ~na_pad & n28356 ;
  assign n28390 = ~\P3_State_reg[1]/NET0131  & ~n28389 ;
  assign n28391 = \P3_State_reg[2]/NET0131  & ~n28390 ;
  assign n28392 = ~n28388 & ~n28391 ;
  assign n28393 = ~n28385 & ~n28392 ;
  assign n28394 = \P1_State_reg[0]/NET0131  & ~\P1_State_reg[1]/NET0131  ;
  assign n28395 = ~\P1_State_reg[2]/NET0131  & n28394 ;
  assign n28396 = \P1_State_reg[0]/NET0131  & ~n2317 ;
  assign n28397 = ~\P1_State_reg[0]/NET0131  & na_pad ;
  assign n28398 = \P1_State_reg[2]/NET0131  & ~n28397 ;
  assign n28399 = ~n28396 & ~n28398 ;
  assign n28400 = ~hold_pad & ~n28399 ;
  assign n28401 = ~n28395 & ~n28400 ;
  assign n28402 = \P1_RequestPending_reg/NET0131  & ~n28401 ;
  assign n28403 = ~n26647 & ~n28402 ;
  assign n28405 = ~\P3_rEIP_reg[15]/NET0131  & ~n26557 ;
  assign n28406 = n2783 & ~n26558 ;
  assign n28407 = ~n28405 & n28406 ;
  assign n28404 = \P3_Address_reg[13]/NET0131  & ~n2782 ;
  assign n28408 = ~\P3_rEIP_reg[14]/NET0131  & ~n27344 ;
  assign n28409 = n26540 & ~n26926 ;
  assign n28410 = ~n28408 & n28409 ;
  assign n28411 = ~n28404 & ~n28410 ;
  assign n28412 = ~n28407 & n28411 ;
  assign n28414 = ~\P2_rEIP_reg[15]/NET0131  & ~n27353 ;
  assign n28415 = n1816 & ~n28085 ;
  assign n28416 = ~n28414 & n28415 ;
  assign n28413 = \P2_Address_reg[13]/NET0131  & ~n1815 ;
  assign n28417 = ~\P2_rEIP_reg[14]/NET0131  & ~n27357 ;
  assign n28418 = n26575 & ~n28089 ;
  assign n28419 = ~n28417 & n28418 ;
  assign n28420 = ~n28413 & ~n28419 ;
  assign n28421 = ~n28416 & n28420 ;
  assign n28423 = ~\P1_rEIP_reg[15]/NET0131  & ~n26629 ;
  assign n28424 = n2308 & ~n26630 ;
  assign n28425 = ~n28423 & n28424 ;
  assign n28422 = \address1[13]_pad  & ~n2307 ;
  assign n28426 = ~\P1_rEIP_reg[14]/NET0131  & ~n27369 ;
  assign n28427 = n26647 & ~n27666 ;
  assign n28428 = ~n28426 & n28427 ;
  assign n28429 = ~n28422 & ~n28428 ;
  assign n28430 = ~n28425 & n28429 ;
  assign n28436 = ~\P2_rEIP_reg[11]/NET0131  & ~n26593 ;
  assign n28437 = n1816 & ~n26594 ;
  assign n28438 = ~n28436 & n28437 ;
  assign n28431 = \P2_Address_reg[9]/NET0131  & ~n1815 ;
  assign n28433 = ~n18999 & n26576 ;
  assign n28432 = ~\P2_rEIP_reg[10]/NET0131  & ~n26576 ;
  assign n28434 = n26575 & ~n28432 ;
  assign n28435 = ~n28433 & n28434 ;
  assign n28439 = ~n28431 & ~n28435 ;
  assign n28440 = ~n28438 & n28439 ;
  assign n28442 = ~\P3_rEIP_reg[11]/NET0131  & ~n26553 ;
  assign n28443 = n2783 & ~n26554 ;
  assign n28444 = ~n28442 & n28443 ;
  assign n28441 = \P3_Address_reg[9]/NET0131  & ~n2782 ;
  assign n28445 = n20421 & n26534 ;
  assign n28446 = ~\P3_rEIP_reg[10]/NET0131  & ~n28445 ;
  assign n28447 = n26540 & ~n27341 ;
  assign n28448 = ~n28446 & n28447 ;
  assign n28449 = ~n28441 & ~n28448 ;
  assign n28450 = ~n28444 & n28449 ;
  assign n28456 = ~\P1_rEIP_reg[11]/NET0131  & ~n26625 ;
  assign n28457 = n2308 & ~n26626 ;
  assign n28458 = ~n28456 & n28457 ;
  assign n28451 = \address1[9]_pad  & ~n2307 ;
  assign n28453 = ~n21494 & n26642 ;
  assign n28452 = ~\P1_rEIP_reg[10]/NET0131  & ~n26642 ;
  assign n28454 = n26647 & ~n28452 ;
  assign n28455 = ~n28453 & n28454 ;
  assign n28459 = ~n28451 & ~n28455 ;
  assign n28460 = ~n28458 & n28459 ;
  assign n28462 = ~\P3_rEIP_reg[23]/NET0131  & ~n26562 ;
  assign n28463 = n2783 & ~n26563 ;
  assign n28464 = ~n28462 & n28463 ;
  assign n28461 = \P3_Address_reg[21]/NET0131  & ~n2782 ;
  assign n28465 = ~\P3_rEIP_reg[22]/NET0131  & ~n27554 ;
  assign n28466 = ~n26536 & n26540 ;
  assign n28467 = ~n28465 & n28466 ;
  assign n28468 = ~n28461 & ~n28467 ;
  assign n28469 = ~n28464 & n28468 ;
  assign n28471 = ~\P2_rEIP_reg[23]/NET0131  & ~n26600 ;
  assign n28472 = n1816 & ~n26601 ;
  assign n28473 = ~n28471 & n28472 ;
  assign n28470 = \P2_Address_reg[21]/NET0131  & ~n1815 ;
  assign n28474 = ~\P2_rEIP_reg[22]/NET0131  & ~n27567 ;
  assign n28475 = n26575 & ~n28145 ;
  assign n28476 = ~n28474 & n28475 ;
  assign n28477 = ~n28470 & ~n28476 ;
  assign n28478 = ~n28473 & n28477 ;
  assign n28480 = ~\P1_rEIP_reg[23]/NET0131  & ~n27577 ;
  assign n28481 = n2308 & ~n28152 ;
  assign n28482 = ~n28480 & n28481 ;
  assign n28479 = \address1[21]_pad  & ~n2307 ;
  assign n28483 = ~\P1_rEIP_reg[22]/NET0131  & ~n27582 ;
  assign n28484 = n26647 & ~n28156 ;
  assign n28485 = ~n28483 & n28484 ;
  assign n28486 = ~n28479 & ~n28485 ;
  assign n28487 = ~n28482 & n28486 ;
  assign n28488 = \P2_State_reg[0]/NET0131  & \P2_State_reg[1]/NET0131  ;
  assign n28489 = ~\P2_State_reg[2]/NET0131  & n28488 ;
  assign n28490 = ~\P2_RequestPending_reg/NET0131  & ~hold_pad ;
  assign n28491 = n1805 & ~n28490 ;
  assign n28492 = n28489 & n28491 ;
  assign n28493 = ~n1818 & ~n28492 ;
  assign n28494 = ~na_pad & ~n28493 ;
  assign n28495 = ~\P2_RequestPending_reg/NET0131  & ~\P2_State_reg[1]/NET0131  ;
  assign n28496 = ~\P2_State_reg[2]/NET0131  & ~n28495 ;
  assign n28497 = \P2_State_reg[0]/NET0131  & hold_pad ;
  assign n28498 = ~n28496 & n28497 ;
  assign n28499 = \P2_State_reg[1]/NET0131  & \P2_State_reg[2]/NET0131  ;
  assign n28500 = ~n28372 & n28499 ;
  assign n28501 = ~n28498 & ~n28500 ;
  assign n28502 = ~n28494 & n28501 ;
  assign n28508 = \P3_State_reg[0]/NET0131  & \P3_State_reg[1]/NET0131  ;
  assign n28509 = ~\P3_State_reg[2]/NET0131  & n28508 ;
  assign n28510 = ~\P3_RequestPending_reg/NET0131  & ~hold_pad ;
  assign n28511 = ~na_pad & n2835 ;
  assign n28512 = ~n28510 & n28511 ;
  assign n28513 = n28509 & n28512 ;
  assign n28503 = hold_pad & n28384 ;
  assign n28504 = ~\P3_State_reg[1]/NET0131  & na_pad ;
  assign n28505 = ~\P3_State_reg[0]/NET0131  & ~n28504 ;
  assign n28506 = ~n28351 & ~n28505 ;
  assign n28507 = \P3_State_reg[2]/NET0131  & ~n28506 ;
  assign n28514 = ~n28503 & ~n28507 ;
  assign n28515 = ~n28513 & n28514 ;
  assign n28516 = \P1_State_reg[0]/NET0131  & \P1_State_reg[1]/NET0131  ;
  assign n28517 = ~\P1_State_reg[2]/NET0131  & n28516 ;
  assign n28518 = ~\P1_RequestPending_reg/NET0131  & ~hold_pad ;
  assign n28519 = n2317 & ~n28518 ;
  assign n28520 = n28517 & n28519 ;
  assign n28521 = ~n2310 & ~n28520 ;
  assign n28522 = ~na_pad & ~n28521 ;
  assign n28523 = \P1_RequestPending_reg/NET0131  & ~\P1_State_reg[2]/NET0131  ;
  assign n28524 = hold_pad & n28394 ;
  assign n28525 = ~n28523 & n28524 ;
  assign n28526 = ~hold_pad & n28396 ;
  assign n28527 = \P1_State_reg[1]/NET0131  & \P1_State_reg[2]/NET0131  ;
  assign n28528 = ~n28526 & n28527 ;
  assign n28529 = ~n28525 & ~n28528 ;
  assign n28530 = ~n28522 & n28529 ;
  assign n28532 = ~\P2_DataWidth_reg[0]/NET0131  & ~\P2_DataWidth_reg[1]/NET0131  ;
  assign n28533 = \P2_DataWidth_reg[0]/NET0131  & \P2_DataWidth_reg[1]/NET0131  ;
  assign n28534 = \P2_rEIP_reg[1]/NET0131  & ~n28533 ;
  assign n28535 = ~n28532 & ~n28534 ;
  assign n28536 = \P2_rEIP_reg[0]/NET0131  & ~n28535 ;
  assign n28531 = ~\P2_rEIP_reg[0]/NET0131  & n19574 ;
  assign n28537 = \P2_ByteEnable_reg[2]/NET0131  & n28533 ;
  assign n28538 = ~n28531 & ~n28537 ;
  assign n28539 = ~n28536 & n28538 ;
  assign n28540 = \P1_DataWidth_reg[0]/NET0131  & \P1_DataWidth_reg[1]/NET0131  ;
  assign n28542 = \P1_rEIP_reg[1]/NET0131  & ~n28540 ;
  assign n28543 = \P1_rEIP_reg[0]/NET0131  & n28542 ;
  assign n28541 = \P1_ByteEnable_reg[2]/NET0131  & n28540 ;
  assign n28544 = \P1_DataWidth_reg[0]/NET0131  & \P1_rEIP_reg[0]/NET0131  ;
  assign n28545 = n18811 & ~n28544 ;
  assign n28546 = ~n28541 & ~n28545 ;
  assign n28547 = ~n28543 & n28546 ;
  assign n28549 = ~\P3_DataWidth_reg[0]/NET0131  & ~\P3_DataWidth_reg[1]/NET0131  ;
  assign n28550 = \P3_DataWidth_reg[0]/NET0131  & \P3_DataWidth_reg[1]/NET0131  ;
  assign n28551 = \P3_rEIP_reg[1]/NET0131  & ~n28550 ;
  assign n28552 = ~n28549 & ~n28551 ;
  assign n28553 = \P3_rEIP_reg[0]/NET0131  & ~n28552 ;
  assign n28548 = ~\P3_rEIP_reg[0]/NET0131  & n20805 ;
  assign n28554 = \P3_ByteEnable_reg[2]/NET0131  & n28550 ;
  assign n28555 = ~n28548 & ~n28554 ;
  assign n28556 = ~n28553 & n28555 ;
  assign n28558 = ~\P3_DataWidth_reg[0]/NET0131  & ~\P3_rEIP_reg[0]/NET0131  ;
  assign n28559 = ~\P3_DataWidth_reg[1]/NET0131  & n28558 ;
  assign n28557 = \P3_ByteEnable_reg[1]/NET0131  & n28550 ;
  assign n28560 = ~n28551 & ~n28557 ;
  assign n28561 = ~n28559 & n28560 ;
  assign n28563 = ~\P1_DataWidth_reg[0]/NET0131  & ~\P1_rEIP_reg[0]/NET0131  ;
  assign n28564 = ~\P1_DataWidth_reg[1]/NET0131  & n28563 ;
  assign n28562 = \P1_ByteEnable_reg[1]/NET0131  & n28540 ;
  assign n28565 = ~n28542 & ~n28562 ;
  assign n28566 = ~n28564 & n28565 ;
  assign n28568 = ~\P2_DataWidth_reg[0]/NET0131  & ~\P2_rEIP_reg[0]/NET0131  ;
  assign n28569 = ~\P2_DataWidth_reg[1]/NET0131  & n28568 ;
  assign n28567 = \P2_ByteEnable_reg[1]/NET0131  & n28533 ;
  assign n28570 = ~n28534 & ~n28567 ;
  assign n28571 = ~n28569 & n28570 ;
  assign n28573 = ~\P3_rEIP_reg[3]/NET0131  & ~n26545 ;
  assign n28574 = n2783 & ~n26546 ;
  assign n28575 = ~n28573 & n28574 ;
  assign n28572 = \P3_Address_reg[1]/NET0131  & ~n2782 ;
  assign n28576 = ~\P3_rEIP_reg[2]/NET0131  & ~n27625 ;
  assign n28577 = n26540 & ~n27626 ;
  assign n28578 = ~n28576 & n28577 ;
  assign n28579 = ~n28572 & ~n28578 ;
  assign n28580 = ~n28575 & n28579 ;
  assign n28582 = ~\P2_rEIP_reg[3]/NET0131  & ~n26587 ;
  assign n28583 = n1816 & ~n26588 ;
  assign n28584 = ~n28582 & n28583 ;
  assign n28581 = \P2_Address_reg[1]/NET0131  & ~n1815 ;
  assign n28585 = ~\P2_rEIP_reg[2]/NET0131  & ~n27641 ;
  assign n28586 = n26575 & ~n27642 ;
  assign n28587 = ~n28585 & n28586 ;
  assign n28588 = ~n28581 & ~n28587 ;
  assign n28589 = ~n28584 & n28588 ;
  assign n28591 = ~\P1_rEIP_reg[3]/NET0131  & ~n26617 ;
  assign n28592 = n2308 & ~n26618 ;
  assign n28593 = ~n28591 & n28592 ;
  assign n28590 = \address1[1]_pad  & ~n2307 ;
  assign n28594 = ~\P1_rEIP_reg[2]/NET0131  & ~n27655 ;
  assign n28595 = n26647 & ~n27656 ;
  assign n28596 = ~n28594 & n28595 ;
  assign n28597 = ~n28590 & ~n28596 ;
  assign n28598 = ~n28593 & n28597 ;
  assign n28600 = ~\P3_rEIP_reg[19]/NET0131  & ~n26921 ;
  assign n28601 = n2783 & ~n28220 ;
  assign n28602 = ~n28600 & n28601 ;
  assign n28599 = \P3_Address_reg[17]/NET0131  & ~n2782 ;
  assign n28603 = ~\P3_rEIP_reg[18]/NET0131  & ~n26929 ;
  assign n28604 = n26540 & ~n28224 ;
  assign n28605 = ~n28603 & n28604 ;
  assign n28606 = ~n28599 & ~n28605 ;
  assign n28607 = ~n28602 & n28606 ;
  assign n28613 = ~\P1_rEIP_reg[19]/NET0131  & ~n26951 ;
  assign n28614 = n2308 & ~n27573 ;
  assign n28615 = ~n28613 & n28614 ;
  assign n28608 = \address1[17]_pad  & ~n2307 ;
  assign n28610 = ~n18735 & n26642 ;
  assign n28609 = ~\P1_rEIP_reg[18]/NET0131  & ~n26642 ;
  assign n28611 = n26647 & ~n28609 ;
  assign n28612 = ~n28610 & n28611 ;
  assign n28616 = ~n28608 & ~n28612 ;
  assign n28617 = ~n28615 & n28616 ;
  assign n28623 = ~\P2_rEIP_reg[19]/NET0131  & ~n26596 ;
  assign n28624 = n1816 & ~n26597 ;
  assign n28625 = ~n28623 & n28624 ;
  assign n28618 = \P2_Address_reg[17]/NET0131  & ~n1815 ;
  assign n28620 = ~n19466 & n26576 ;
  assign n28619 = ~\P2_rEIP_reg[18]/NET0131  & ~n26576 ;
  assign n28621 = n26575 & ~n28619 ;
  assign n28622 = ~n28620 & n28621 ;
  assign n28626 = ~n28618 & ~n28622 ;
  assign n28627 = ~n28625 & n28626 ;
  assign n28629 = ~\P3_rEIP_reg[7]/NET0131  & ~n26549 ;
  assign n28630 = n2783 & ~n26550 ;
  assign n28631 = ~n28629 & n28630 ;
  assign n28628 = \P3_Address_reg[5]/NET0131  & ~n2782 ;
  assign n28632 = ~\P3_rEIP_reg[6]/NET0131  & ~n27630 ;
  assign n28633 = n26540 & ~n28250 ;
  assign n28634 = ~n28632 & n28633 ;
  assign n28635 = ~n28628 & ~n28634 ;
  assign n28636 = ~n28631 & n28635 ;
  assign n28642 = ~\P2_rEIP_reg[7]/NET0131  & ~n27637 ;
  assign n28643 = n1816 & ~n26590 ;
  assign n28644 = ~n28642 & n28643 ;
  assign n28637 = \P2_Address_reg[5]/NET0131  & ~n1815 ;
  assign n28639 = \P2_rEIP_reg[6]/NET0131  & n27645 ;
  assign n28638 = ~\P2_rEIP_reg[6]/NET0131  & ~n27645 ;
  assign n28640 = n26575 & ~n28638 ;
  assign n28641 = ~n28639 & n28640 ;
  assign n28645 = ~n28637 & ~n28641 ;
  assign n28646 = ~n28644 & n28645 ;
  assign n28648 = ~\P1_rEIP_reg[7]/NET0131  & ~n26621 ;
  assign n28649 = n2308 & ~n26622 ;
  assign n28650 = ~n28648 & n28649 ;
  assign n28647 = \address1[5]_pad  & ~n2307 ;
  assign n28651 = ~\P1_rEIP_reg[6]/NET0131  & ~n27659 ;
  assign n28652 = n26647 & ~n27609 ;
  assign n28653 = ~n28651 & n28652 ;
  assign n28654 = ~n28647 & ~n28653 ;
  assign n28655 = ~n28650 & n28654 ;
  assign n28656 = \P1_ByteEnable_reg[3]/NET0131  & n28540 ;
  assign n28657 = \P1_rEIP_reg[1]/NET0131  & ~n28563 ;
  assign n28658 = ~\P1_DataWidth_reg[1]/NET0131  & ~n28657 ;
  assign n28659 = ~n28656 & ~n28658 ;
  assign n28660 = \P3_ByteEnable_reg[3]/NET0131  & n28550 ;
  assign n28661 = \P3_rEIP_reg[1]/NET0131  & ~n28558 ;
  assign n28662 = ~\P3_DataWidth_reg[1]/NET0131  & ~n28661 ;
  assign n28663 = ~n28660 & ~n28662 ;
  assign n28664 = \P2_ByteEnable_reg[3]/NET0131  & n28533 ;
  assign n28665 = \P2_rEIP_reg[1]/NET0131  & ~n28568 ;
  assign n28666 = ~\P2_DataWidth_reg[1]/NET0131  & ~n28665 ;
  assign n28667 = ~n28664 & ~n28666 ;
  assign n28669 = ~\P1_rEIP_reg[2]/NET0131  & ~n26616 ;
  assign n28670 = n2308 & ~n26617 ;
  assign n28671 = ~n28669 & n28670 ;
  assign n28668 = \address1[0]_pad  & ~n2307 ;
  assign n28672 = ~\P1_rEIP_reg[1]/NET0131  & ~n26642 ;
  assign n28673 = n26647 & ~n27655 ;
  assign n28674 = ~n28672 & n28673 ;
  assign n28675 = ~n28668 & ~n28674 ;
  assign n28676 = ~n28671 & n28675 ;
  assign n28677 = ~\P2_rEIP_reg[2]/NET0131  & ~n26586 ;
  assign n28678 = ~\P2_State_reg[2]/NET0131  & ~n26587 ;
  assign n28679 = ~n28677 & n28678 ;
  assign n28680 = ~\P2_rEIP_reg[1]/NET0131  & ~n26576 ;
  assign n28681 = \P2_State_reg[2]/NET0131  & ~n27641 ;
  assign n28682 = ~n28680 & n28681 ;
  assign n28683 = ~n28679 & ~n28682 ;
  assign n28684 = n1815 & ~n28683 ;
  assign n28685 = \P2_Address_reg[0]/NET0131  & ~n1815 ;
  assign n28686 = ~n28684 & ~n28685 ;
  assign n28687 = ~\P3_rEIP_reg[2]/NET0131  & ~n26544 ;
  assign n28688 = ~\P3_State_reg[2]/NET0131  & ~n26545 ;
  assign n28689 = ~n28687 & n28688 ;
  assign n28690 = ~\P3_rEIP_reg[1]/NET0131  & ~n26534 ;
  assign n28691 = \P3_State_reg[2]/NET0131  & ~n27625 ;
  assign n28692 = ~n28690 & n28691 ;
  assign n28693 = ~n28689 & ~n28692 ;
  assign n28694 = n2782 & ~n28693 ;
  assign n28695 = \P3_Address_reg[0]/NET0131  & ~n2782 ;
  assign n28696 = ~n28694 & ~n28695 ;
  assign n28697 = ~\P2_Address_reg[29]/NET0131  & n27887 ;
  assign n28700 = ~\ast2_pad  & ~dc_pad ;
  assign n28701 = mio_pad & ~wr_pad ;
  assign n28702 = n28700 & n28701 ;
  assign n28698 = ~\P3_BE_n_reg[0]/NET0131  & ~\P3_BE_n_reg[1]/NET0131  ;
  assign n28699 = ~\P3_BE_n_reg[2]/NET0131  & ~\P3_BE_n_reg[3]/NET0131  ;
  assign n28703 = n28698 & n28699 ;
  assign n28704 = n28702 & n28703 ;
  assign n28705 = ~n28697 & n28704 ;
  assign n28706 = ~n2784 & ~n28509 ;
  assign n28707 = ~\P3_DataWidth_reg[1]/NET0131  & n28706 ;
  assign n28708 = ~n2785 & ~n28509 ;
  assign n28709 = ~\bs16_pad  & ~n28708 ;
  assign n28710 = ~n28707 & ~n28709 ;
  assign n28711 = ~n1818 & ~n28489 ;
  assign n28712 = ~\bs16_pad  & ~n28711 ;
  assign n28713 = ~n1817 & ~n28489 ;
  assign n28714 = ~\P2_DataWidth_reg[1]/NET0131  & n28713 ;
  assign n28715 = ~n28712 & ~n28714 ;
  assign n28716 = ~n2310 & ~n28517 ;
  assign n28717 = ~\bs16_pad  & ~n28716 ;
  assign n28718 = ~n2309 & ~n28517 ;
  assign n28719 = ~\P1_DataWidth_reg[1]/NET0131  & n28718 ;
  assign n28720 = ~n28717 & ~n28719 ;
  assign n28721 = \P1_BE_n_reg[2]/NET0131  & ~n2307 ;
  assign n28722 = \P1_ByteEnable_reg[2]/NET0131  & n2307 ;
  assign n28723 = ~n28721 & ~n28722 ;
  assign n28724 = \P1_BE_n_reg[3]/NET0131  & ~n2307 ;
  assign n28725 = \P1_ByteEnable_reg[3]/NET0131  & n2307 ;
  assign n28726 = ~n28724 & ~n28725 ;
  assign n28727 = \P3_State_reg[0]/NET0131  & \ast2_pad  ;
  assign n28728 = n28706 & ~n28727 ;
  assign n28729 = \P3_DataWidth_reg[0]/NET0131  & n28706 ;
  assign n28730 = ~n28709 & ~n28729 ;
  assign n28731 = \P2_BE_n_reg[0]/NET0131  & ~n1815 ;
  assign n28732 = \P2_ByteEnable_reg[0]/NET0131  & n1815 ;
  assign n28733 = ~n28731 & ~n28732 ;
  assign n28734 = \P2_BE_n_reg[3]/NET0131  & ~n1815 ;
  assign n28735 = \P2_ByteEnable_reg[3]/NET0131  & n1815 ;
  assign n28736 = ~n28734 & ~n28735 ;
  assign n28737 = \P2_DataWidth_reg[0]/NET0131  & n28713 ;
  assign n28738 = ~n28712 & ~n28737 ;
  assign n28739 = \P3_BE_n_reg[3]/NET0131  & ~n2782 ;
  assign n28740 = \P3_ByteEnable_reg[3]/NET0131  & n2782 ;
  assign n28741 = ~n28739 & ~n28740 ;
  assign n28742 = \P3_BE_n_reg[1]/NET0131  & ~n2782 ;
  assign n28743 = \P3_ByteEnable_reg[1]/NET0131  & n2782 ;
  assign n28744 = ~n28742 & ~n28743 ;
  assign n28745 = \P3_BE_n_reg[2]/NET0131  & ~n2782 ;
  assign n28746 = \P3_ByteEnable_reg[2]/NET0131  & n2782 ;
  assign n28747 = ~n28745 & ~n28746 ;
  assign n28748 = \P3_BE_n_reg[0]/NET0131  & ~n2782 ;
  assign n28749 = \P3_ByteEnable_reg[0]/NET0131  & n2782 ;
  assign n28750 = ~n28748 & ~n28749 ;
  assign n28751 = \P1_State_reg[0]/NET0131  & \ast1_pad  ;
  assign n28752 = n28718 & ~n28751 ;
  assign n28753 = \P2_ADS_n_reg/NET0131  & \P2_State_reg[0]/NET0131  ;
  assign n28754 = n28713 & ~n28753 ;
  assign n28755 = mio_pad & ~n2782 ;
  assign n28756 = \P3_MemoryFetch_reg/NET0131  & n2782 ;
  assign n28757 = ~n28755 & ~n28756 ;
  assign n28758 = wr_pad & ~n2782 ;
  assign n28759 = ~\P3_ReadRequest_reg/NET0131  & n2782 ;
  assign n28760 = ~n28758 & ~n28759 ;
  assign n28761 = \P1_DataWidth_reg[0]/NET0131  & n28718 ;
  assign n28762 = ~n28717 & ~n28761 ;
  assign n28763 = \P1_M_IO_n_reg/NET0131  & ~n2307 ;
  assign n28764 = \P1_MemoryFetch_reg/NET0131  & n2307 ;
  assign n28765 = ~n28763 & ~n28764 ;
  assign n28766 = \P2_BE_n_reg[2]/NET0131  & ~n1815 ;
  assign n28767 = \P2_ByteEnable_reg[2]/NET0131  & n1815 ;
  assign n28768 = ~n28766 & ~n28767 ;
  assign n28769 = \P2_W_R_n_reg/NET0131  & ~n1815 ;
  assign n28770 = ~\P2_ReadRequest_reg/NET0131  & n1815 ;
  assign n28771 = ~n28769 & ~n28770 ;
  assign n28772 = \P2_BE_n_reg[1]/NET0131  & ~n1815 ;
  assign n28773 = \P2_ByteEnable_reg[1]/NET0131  & n1815 ;
  assign n28774 = ~n28772 & ~n28773 ;
  assign n28775 = \P1_W_R_n_reg/NET0131  & ~n2307 ;
  assign n28776 = ~\P1_ReadRequest_reg/NET0131  & n2307 ;
  assign n28777 = ~n28775 & ~n28776 ;
  assign n28778 = \P1_BE_n_reg[0]/NET0131  & ~n2307 ;
  assign n28779 = \P1_ByteEnable_reg[0]/NET0131  & n2307 ;
  assign n28780 = ~n28778 & ~n28779 ;
  assign n28781 = \P2_M_IO_n_reg/NET0131  & ~n1815 ;
  assign n28782 = \P2_MemoryFetch_reg/NET0131  & n1815 ;
  assign n28783 = ~n28781 & ~n28782 ;
  assign n28784 = \P1_BE_n_reg[1]/NET0131  & ~n2307 ;
  assign n28785 = \P1_ByteEnable_reg[1]/NET0131  & n2307 ;
  assign n28786 = ~n28784 & ~n28785 ;
  assign n28787 = ~\P3_State_reg[1]/NET0131  & \P3_State_reg[2]/NET0131  ;
  assign n28788 = ~\P3_State_reg[0]/NET0131  & ~n28787 ;
  assign n28789 = ~dc_pad & ~n28788 ;
  assign n28790 = \P3_CodeFetch_reg/NET0131  & n2782 ;
  assign n28791 = ~n28789 & ~n28790 ;
  assign n28792 = ~\P2_State_reg[1]/NET0131  & \P2_State_reg[2]/NET0131  ;
  assign n28793 = ~\P2_State_reg[0]/NET0131  & ~n28792 ;
  assign n28794 = ~\P2_D_C_n_reg/NET0131  & ~n28793 ;
  assign n28795 = \P2_CodeFetch_reg/NET0131  & n1815 ;
  assign n28796 = ~n28794 & ~n28795 ;
  assign n28797 = ~\P1_State_reg[1]/NET0131  & \P1_State_reg[2]/NET0131  ;
  assign n28798 = ~\P1_State_reg[0]/NET0131  & ~n28797 ;
  assign n28799 = ~\P1_D_C_n_reg/NET0131  & ~n28798 ;
  assign n28800 = \P1_CodeFetch_reg/NET0131  & n2307 ;
  assign n28801 = ~n28799 & ~n28800 ;
  assign n28804 = \P3_InstAddrPointer_reg[10]/NET0131  & n2896 ;
  assign n28805 = ~n14479 & ~n28804 ;
  assign n28806 = n2894 & ~n28805 ;
  assign n28803 = ~n2777 & n4215 ;
  assign n28807 = n2918 & n4301 ;
  assign n28810 = ~n28803 & ~n28807 ;
  assign n28808 = \P3_InstAddrPointer_reg[10]/NET0131  & ~n4402 ;
  assign n28809 = ~n2923 & n6071 ;
  assign n28811 = ~n28808 & ~n28809 ;
  assign n28812 = n28810 & n28811 ;
  assign n28813 = ~n14484 & n28812 ;
  assign n28814 = ~n28806 & n28813 ;
  assign n28815 = n2453 & ~n28814 ;
  assign n28802 = \P3_InstAddrPointer_reg[10]/NET0131  & ~n4418 ;
  assign n28816 = ~n14494 & ~n28802 ;
  assign n28817 = ~n28815 & n28816 ;
  assign n28818 = \P3_InstAddrPointer_reg[29]/NET0131  & n2896 ;
  assign n28819 = ~n11210 & ~n28818 ;
  assign n28820 = n2894 & ~n28819 ;
  assign n28825 = n2918 & n11216 ;
  assign n28822 = ~n2841 & ~n6113 ;
  assign n28823 = n4402 & ~n28822 ;
  assign n28824 = \P3_InstAddrPointer_reg[29]/NET0131  & ~n28823 ;
  assign n28821 = ~n2777 & n4146 ;
  assign n28826 = \P3_InstAddrPointer_reg[29]/NET0131  & n20473 ;
  assign n28827 = n2923 & ~n28826 ;
  assign n28828 = n11195 & ~n28827 ;
  assign n28829 = ~n28821 & ~n28828 ;
  assign n28830 = ~n28824 & n28829 ;
  assign n28831 = ~n28825 & n28830 ;
  assign n28832 = ~n11220 & n28831 ;
  assign n28833 = ~n28820 & n28832 ;
  assign n28834 = n2453 & ~n28833 ;
  assign n28835 = \P3_InstAddrPointer_reg[29]/NET0131  & ~n4418 ;
  assign n28836 = ~n11233 & ~n28835 ;
  assign n28837 = ~n28834 & n28836 ;
  assign n28839 = \P2_InstAddrPointer_reg[20]/NET0131  & n1897 ;
  assign n28840 = ~n11860 & ~n28839 ;
  assign n28841 = n1734 & ~n28840 ;
  assign n28838 = ~n1771 & n6537 ;
  assign n28842 = n1870 & n11045 ;
  assign n28845 = ~n28838 & ~n28842 ;
  assign n28843 = \P2_InstAddrPointer_reg[20]/NET0131  & ~n12566 ;
  assign n28844 = ~n1831 & n6666 ;
  assign n28846 = ~n28843 & ~n28844 ;
  assign n28847 = n28845 & n28846 ;
  assign n28848 = ~n11867 & n28847 ;
  assign n28849 = ~n28841 & n28848 ;
  assign n28850 = n1927 & ~n28849 ;
  assign n28851 = \P2_InstAddrPointer_reg[20]/NET0131  & ~n6810 ;
  assign n28852 = ~n11880 & ~n28851 ;
  assign n28853 = ~n28850 & n28852 ;
  assign n28854 = \P2_InstAddrPointer_reg[31]/NET0131  & n1897 ;
  assign n28855 = ~n8933 & ~n28854 ;
  assign n28856 = n1734 & ~n28855 ;
  assign n28860 = n1870 & ~n8949 ;
  assign n28857 = ~n1771 & ~n8927 ;
  assign n28858 = ~n1831 & n8907 ;
  assign n28859 = \P2_InstAddrPointer_reg[31]/NET0131  & ~n12566 ;
  assign n28861 = ~n28858 & ~n28859 ;
  assign n28862 = ~n28857 & n28861 ;
  assign n28863 = ~n28860 & n28862 ;
  assign n28864 = ~n8953 & n28863 ;
  assign n28865 = ~n28856 & n28864 ;
  assign n28866 = n1927 & ~n28865 ;
  assign n28867 = \P2_InstAddrPointer_reg[31]/NET0131  & ~n6810 ;
  assign n28868 = ~n8992 & ~n28867 ;
  assign n28869 = ~n28866 & n28868 ;
  assign n28872 = \P3_InstAddrPointer_reg[13]/NET0131  & n2896 ;
  assign n28873 = ~n13086 & ~n28872 ;
  assign n28874 = n2894 & ~n28873 ;
  assign n28871 = n2918 & n13091 ;
  assign n28875 = ~n2923 & n8358 ;
  assign n28878 = ~n28871 & ~n28875 ;
  assign n28876 = \P3_InstAddrPointer_reg[13]/NET0131  & ~n4402 ;
  assign n28877 = ~n2777 & n4175 ;
  assign n28879 = ~n28876 & ~n28877 ;
  assign n28880 = n28878 & n28879 ;
  assign n28881 = ~n13095 & n28880 ;
  assign n28882 = ~n28874 & n28881 ;
  assign n28883 = n2453 & ~n28882 ;
  assign n28870 = \P3_InstAddrPointer_reg[13]/NET0131  & ~n4418 ;
  assign n28884 = ~n13106 & ~n28870 ;
  assign n28885 = ~n28883 & n28884 ;
  assign n28888 = \P2_InstAddrPointer_reg[19]/NET0131  & n1897 ;
  assign n28889 = ~n12413 & ~n28888 ;
  assign n28890 = n1734 & ~n28889 ;
  assign n28887 = \P2_InstAddrPointer_reg[19]/NET0131  & ~n12566 ;
  assign n28891 = n1870 & n7552 ;
  assign n28894 = ~n28887 & ~n28891 ;
  assign n28892 = ~n1771 & n6539 ;
  assign n28893 = ~n1831 & n7594 ;
  assign n28895 = ~n28892 & ~n28893 ;
  assign n28896 = n28894 & n28895 ;
  assign n28897 = ~n12420 & n28896 ;
  assign n28898 = ~n28890 & n28897 ;
  assign n28899 = n1927 & ~n28898 ;
  assign n28886 = \P2_InstAddrPointer_reg[19]/NET0131  & ~n6810 ;
  assign n28900 = ~n12431 & ~n28886 ;
  assign n28901 = ~n28899 & n28900 ;
  assign n28902 = \P3_InstAddrPointer_reg[30]/NET0131  & n2896 ;
  assign n28903 = ~n10057 & ~n28902 ;
  assign n28904 = n2894 & ~n28903 ;
  assign n28908 = n2918 & n4385 ;
  assign n28907 = ~n2923 & ~n4120 ;
  assign n28905 = ~n2777 & n4153 ;
  assign n28906 = \P3_InstAddrPointer_reg[30]/NET0131  & ~n4402 ;
  assign n28909 = ~n28905 & ~n28906 ;
  assign n28910 = ~n28907 & n28909 ;
  assign n28911 = ~n28908 & n28910 ;
  assign n28912 = ~n10065 & n28911 ;
  assign n28913 = ~n28904 & n28912 ;
  assign n28914 = n2453 & ~n28913 ;
  assign n28915 = \P3_InstAddrPointer_reg[30]/NET0131  & ~n4418 ;
  assign n28916 = ~n10078 & ~n28915 ;
  assign n28917 = ~n28914 & n28916 ;
  assign n28918 = \P2_InstAddrPointer_reg[30]/NET0131  & n1897 ;
  assign n28919 = ~n10010 & ~n28918 ;
  assign n28920 = n1734 & ~n28919 ;
  assign n28921 = ~n1727 & n10015 ;
  assign n28922 = n12566 & ~n28921 ;
  assign n28923 = \P2_InstAddrPointer_reg[30]/NET0131  & ~n28922 ;
  assign n28926 = n1798 & n28921 ;
  assign n28924 = ~n1831 & n9996 ;
  assign n28925 = ~n1771 & n8919 ;
  assign n28927 = ~n28924 & ~n28925 ;
  assign n28928 = ~n28926 & n28927 ;
  assign n28929 = ~n28923 & n28928 ;
  assign n28930 = ~n10021 & n28929 ;
  assign n28931 = ~n28920 & n28930 ;
  assign n28932 = n1927 & ~n28931 ;
  assign n28933 = \P2_InstAddrPointer_reg[30]/NET0131  & ~n6810 ;
  assign n28934 = ~n10031 & ~n28933 ;
  assign n28935 = ~n28932 & n28934 ;
  assign n28950 = ~\P3_InstAddrPointer_reg[19]/NET0131  & ~n4363 ;
  assign n28951 = ~n4364 & ~n28950 ;
  assign n28953 = n4356 & n4360 ;
  assign n28955 = \P3_InstAddrPointer_reg[18]/NET0131  & n28953 ;
  assign n28956 = ~n28951 & ~n28955 ;
  assign n28954 = n3754 & n28953 ;
  assign n28957 = n2905 & ~n28954 ;
  assign n28958 = ~n28956 & n28957 ;
  assign n28941 = ~n4250 & n4281 ;
  assign n28942 = ~n3753 & ~n11092 ;
  assign n28943 = ~n28941 & n28942 ;
  assign n28938 = n3797 & ~n4085 ;
  assign n28939 = ~n6093 & ~n28938 ;
  assign n28940 = n3753 & ~n28939 ;
  assign n28944 = ~n2896 & ~n28940 ;
  assign n28945 = ~n28943 & n28944 ;
  assign n28946 = n2894 & n28945 ;
  assign n28952 = n2918 & n28951 ;
  assign n28948 = \P3_InstAddrPointer_reg[19]/NET0131  & ~n11451 ;
  assign n28947 = ~n2923 & ~n3797 ;
  assign n28949 = ~n2777 & n4281 ;
  assign n28959 = ~n28947 & ~n28949 ;
  assign n28960 = ~n28948 & n28959 ;
  assign n28961 = ~n28952 & n28960 ;
  assign n28962 = ~n28946 & n28961 ;
  assign n28963 = ~n28958 & n28962 ;
  assign n28964 = n2453 & ~n28963 ;
  assign n28936 = \P3_rEIP_reg[19]/NET0131  & n4412 ;
  assign n28937 = \P3_InstAddrPointer_reg[19]/NET0131  & ~n4418 ;
  assign n28965 = ~n28936 & ~n28937 ;
  assign n28966 = ~n28964 & n28965 ;
  assign n28970 = ~n2896 & ~n13182 ;
  assign n28969 = ~\P3_InstAddrPointer_reg[18]/NET0131  & n2896 ;
  assign n28971 = n2894 & ~n28969 ;
  assign n28972 = ~n28970 & n28971 ;
  assign n28968 = n2918 & n13187 ;
  assign n28973 = ~n2923 & n13174 ;
  assign n28976 = ~n28968 & ~n28973 ;
  assign n28974 = \P3_InstAddrPointer_reg[18]/NET0131  & ~n4402 ;
  assign n28975 = ~n2777 & n4248 ;
  assign n28977 = ~n28974 & ~n28975 ;
  assign n28978 = n28976 & n28977 ;
  assign n28979 = ~n13190 & n28978 ;
  assign n28980 = ~n28972 & n28979 ;
  assign n28981 = n2453 & ~n28980 ;
  assign n28967 = \P3_InstAddrPointer_reg[18]/NET0131  & ~n4418 ;
  assign n28982 = ~n13204 & ~n28967 ;
  assign n28983 = ~n28981 & n28982 ;
  assign n28986 = \P3_InstAddrPointer_reg[14]/NET0131  & n2896 ;
  assign n28987 = ~n13120 & ~n28986 ;
  assign n28988 = n2894 & ~n28987 ;
  assign n28985 = ~n2777 & n4171 ;
  assign n28989 = n2918 & n4354 ;
  assign n28992 = ~n28985 & ~n28989 ;
  assign n28990 = \P3_InstAddrPointer_reg[14]/NET0131  & ~n4402 ;
  assign n28991 = ~n2923 & n4066 ;
  assign n28993 = ~n28990 & ~n28991 ;
  assign n28994 = n28992 & n28993 ;
  assign n28995 = ~n13126 & n28994 ;
  assign n28996 = ~n28988 & n28995 ;
  assign n28997 = n2453 & ~n28996 ;
  assign n28984 = \P3_InstAddrPointer_reg[14]/NET0131  & ~n4418 ;
  assign n28998 = ~n13135 & ~n28984 ;
  assign n28999 = ~n28997 & n28998 ;
  assign n29001 = \P3_InstAddrPointer_reg[26]/NET0131  & n2896 ;
  assign n29002 = ~n12125 & ~n29001 ;
  assign n29003 = n2894 & ~n29002 ;
  assign n29000 = n2918 & n12130 ;
  assign n29006 = \P3_InstAddrPointer_reg[26]/NET0131  & ~n4402 ;
  assign n29004 = ~n2923 & n4093 ;
  assign n29005 = ~n2777 & n4277 ;
  assign n29007 = ~n29004 & ~n29005 ;
  assign n29008 = ~n29006 & n29007 ;
  assign n29009 = ~n29000 & n29008 ;
  assign n29010 = ~n12133 & n29009 ;
  assign n29011 = ~n29003 & n29010 ;
  assign n29012 = n2453 & ~n29011 ;
  assign n29013 = \P3_InstAddrPointer_reg[26]/NET0131  & ~n4418 ;
  assign n29014 = ~n12141 & ~n29013 ;
  assign n29015 = ~n29012 & n29014 ;
  assign n29016 = \P1_InstAddrPointer_reg[31]/NET0131  & n2375 ;
  assign n29026 = \P1_InstAddrPointer_reg[31]/NET0131  & ~n4811 ;
  assign n29027 = ~\P1_InstAddrPointer_reg[31]/NET0131  & n4811 ;
  assign n29028 = ~n29026 & ~n29027 ;
  assign n29030 = n4950 & n29028 ;
  assign n29029 = ~n4950 & ~n29028 ;
  assign n29031 = ~n4453 & ~n29029 ;
  assign n29032 = ~n29030 & n29031 ;
  assign n29017 = \P1_InstAddrPointer_reg[30]/NET0131  & n4495 ;
  assign n29018 = n6850 & n29017 ;
  assign n29019 = ~\P1_InstAddrPointer_reg[31]/NET0131  & ~n4800 ;
  assign n29020 = \P1_InstAddrPointer_reg[31]/NET0131  & n4800 ;
  assign n29021 = ~n29019 & ~n29020 ;
  assign n29023 = n29018 & ~n29021 ;
  assign n29022 = ~n29018 & n29021 ;
  assign n29024 = n4453 & ~n29022 ;
  assign n29025 = ~n29023 & n29024 ;
  assign n29033 = ~n2375 & ~n29025 ;
  assign n29034 = ~n29032 & n29033 ;
  assign n29035 = ~n29016 & ~n29034 ;
  assign n29036 = n2244 & ~n29035 ;
  assign n29037 = n5068 & n11284 ;
  assign n29038 = \P1_InstAddrPointer_reg[31]/NET0131  & ~n5065 ;
  assign n29039 = ~\P1_InstAddrPointer_reg[31]/NET0131  & n5065 ;
  assign n29040 = ~n29038 & ~n29039 ;
  assign n29042 = ~n29037 & n29040 ;
  assign n29041 = n29037 & ~n29040 ;
  assign n29043 = n2385 & ~n29041 ;
  assign n29044 = ~n29042 & n29043 ;
  assign n29047 = n2397 & ~n29040 ;
  assign n29046 = ~n2271 & ~n29028 ;
  assign n29045 = ~n2402 & n29021 ;
  assign n29048 = ~n2377 & ~n7247 ;
  assign n29049 = n14810 & ~n29048 ;
  assign n29050 = \P1_InstAddrPointer_reg[31]/NET0131  & ~n29049 ;
  assign n29051 = ~n29045 & ~n29050 ;
  assign n29052 = ~n29046 & n29051 ;
  assign n29053 = ~n29047 & n29052 ;
  assign n29054 = ~n29044 & n29053 ;
  assign n29055 = ~n29036 & n29054 ;
  assign n29056 = n2432 & ~n29055 ;
  assign n29057 = \P1_rEIP_reg[31]/NET0131  & n5092 ;
  assign n29058 = \P1_InstAddrPointer_reg[31]/NET0131  & ~n5098 ;
  assign n29059 = ~n29057 & ~n29058 ;
  assign n29060 = ~n29056 & n29059 ;
  assign n29061 = \P1_InstAddrPointer_reg[27]/NET0131  & n2375 ;
  assign n29062 = ~n11279 & ~n29061 ;
  assign n29063 = n2244 & ~n29062 ;
  assign n29067 = n2397 & n5060 ;
  assign n29064 = \P1_InstAddrPointer_reg[27]/NET0131  & ~n6027 ;
  assign n29065 = ~n2271 & n4942 ;
  assign n29066 = ~n2402 & n4492 ;
  assign n29068 = ~n29065 & ~n29066 ;
  assign n29069 = ~n29064 & n29068 ;
  assign n29070 = ~n29067 & n29069 ;
  assign n29071 = ~n11288 & n29070 ;
  assign n29072 = ~n29063 & n29071 ;
  assign n29073 = n2432 & ~n29072 ;
  assign n29074 = \P1_InstAddrPointer_reg[27]/NET0131  & ~n5098 ;
  assign n29075 = ~n11301 & ~n29074 ;
  assign n29076 = ~n29073 & n29075 ;
  assign n29079 = \P3_InstAddrPointer_reg[17]/NET0131  & n2896 ;
  assign n29085 = ~n4237 & n7337 ;
  assign n29086 = n4240 & ~n29085 ;
  assign n29084 = n4241 & n7337 ;
  assign n29087 = ~n3753 & ~n29084 ;
  assign n29088 = ~n29086 & n29087 ;
  assign n29081 = ~n8350 & n8361 ;
  assign n29080 = n8350 & ~n8361 ;
  assign n29082 = n3753 & ~n29080 ;
  assign n29083 = ~n29081 & n29082 ;
  assign n29089 = ~n2896 & ~n29083 ;
  assign n29090 = ~n29088 & n29089 ;
  assign n29091 = ~n29079 & ~n29090 ;
  assign n29092 = n2894 & ~n29091 ;
  assign n29097 = ~n4356 & ~n4360 ;
  assign n29098 = n2905 & ~n28953 ;
  assign n29099 = ~n29097 & n29098 ;
  assign n29093 = n2918 & n4360 ;
  assign n29094 = ~n2777 & n4240 ;
  assign n29100 = ~n29093 & ~n29094 ;
  assign n29095 = ~n2923 & n8350 ;
  assign n29096 = \P3_InstAddrPointer_reg[17]/NET0131  & ~n4402 ;
  assign n29101 = ~n29095 & ~n29096 ;
  assign n29102 = n29100 & n29101 ;
  assign n29103 = ~n29099 & n29102 ;
  assign n29104 = ~n29092 & n29103 ;
  assign n29105 = n2453 & ~n29104 ;
  assign n29077 = \P3_rEIP_reg[17]/NET0131  & n4412 ;
  assign n29078 = \P3_InstAddrPointer_reg[17]/NET0131  & ~n4418 ;
  assign n29106 = ~n29077 & ~n29078 ;
  assign n29107 = ~n29105 & n29106 ;
  assign n29123 = \P3_InstAddrPointer_reg[23]/NET0131  & n2896 ;
  assign n29124 = ~n11104 & ~n29123 ;
  assign n29125 = n2894 & ~n29124 ;
  assign n29110 = ~n2763 & ~n2818 ;
  assign n29111 = \P3_InstAddrPointer_reg[23]/NET0131  & ~n29110 ;
  assign n29112 = n2834 & ~n29111 ;
  assign n29117 = n2835 & ~n29112 ;
  assign n29118 = ~n2841 & ~n4370 ;
  assign n29119 = ~n2898 & ~n29118 ;
  assign n29120 = n7402 & n29119 ;
  assign n29121 = ~n29117 & n29120 ;
  assign n29122 = \P3_InstAddrPointer_reg[23]/NET0131  & ~n29121 ;
  assign n29113 = ~n2835 & ~n29112 ;
  assign n29114 = ~n2767 & ~n29113 ;
  assign n29115 = n4104 & ~n29114 ;
  assign n29109 = ~n2777 & n4265 ;
  assign n29116 = n2918 & n11110 ;
  assign n29126 = ~n29109 & ~n29116 ;
  assign n29127 = ~n29115 & n29126 ;
  assign n29128 = ~n29122 & n29127 ;
  assign n29129 = ~n11114 & n29128 ;
  assign n29130 = ~n29125 & n29129 ;
  assign n29131 = n2453 & ~n29130 ;
  assign n29108 = \P3_InstAddrPointer_reg[23]/NET0131  & ~n4418 ;
  assign n29132 = ~n11130 & ~n29108 ;
  assign n29133 = ~n29131 & n29132 ;
  assign n29135 = ~\P3_EBX_reg[27]/NET0131  & ~n17453 ;
  assign n29136 = n24549 & ~n29135 ;
  assign n29134 = \P3_EBX_reg[27]/NET0131  & n14954 ;
  assign n29137 = n14011 & n14952 ;
  assign n29138 = ~n29134 & ~n29137 ;
  assign n29139 = ~n29136 & n29138 ;
  assign n29140 = n2453 & ~n29139 ;
  assign n29141 = \P3_EBX_reg[27]/NET0131  & ~n13810 ;
  assign n29142 = ~n29140 & ~n29141 ;
  assign n29145 = \P2_InstAddrPointer_reg[14]/NET0131  & n1897 ;
  assign n29146 = ~n13579 & ~n29145 ;
  assign n29147 = n1734 & ~n29146 ;
  assign n29144 = n1870 & n6751 ;
  assign n29148 = ~n1831 & n6650 ;
  assign n29151 = ~n29144 & ~n29148 ;
  assign n29149 = ~n1771 & n6502 ;
  assign n29150 = \P2_InstAddrPointer_reg[14]/NET0131  & ~n7501 ;
  assign n29152 = ~n29149 & ~n29150 ;
  assign n29153 = n29151 & n29152 ;
  assign n29154 = ~n13586 & n29153 ;
  assign n29155 = ~n29147 & n29154 ;
  assign n29156 = n1927 & ~n29155 ;
  assign n29143 = \P2_InstAddrPointer_reg[14]/NET0131  & ~n6810 ;
  assign n29157 = ~n13593 & ~n29143 ;
  assign n29158 = ~n29156 & n29157 ;
  assign n29161 = \P3_InstAddrPointer_reg[20]/NET0131  & n2896 ;
  assign n29162 = ~n12034 & ~n29161 ;
  assign n29163 = n2894 & ~n29162 ;
  assign n29160 = n2918 & n12039 ;
  assign n29166 = ~n2777 & n4254 ;
  assign n29164 = ~n2923 & n3792 ;
  assign n29165 = \P3_InstAddrPointer_reg[20]/NET0131  & ~n4402 ;
  assign n29167 = ~n29164 & ~n29165 ;
  assign n29168 = ~n29166 & n29167 ;
  assign n29169 = ~n29160 & n29168 ;
  assign n29170 = ~n12044 & n29169 ;
  assign n29171 = ~n29163 & n29170 ;
  assign n29172 = n2453 & ~n29171 ;
  assign n29159 = \P3_InstAddrPointer_reg[20]/NET0131  & ~n4418 ;
  assign n29173 = ~n12058 & ~n29159 ;
  assign n29174 = ~n29172 & n29173 ;
  assign n29177 = \P1_InstAddrPointer_reg[9]/NET0131  & n2375 ;
  assign n29178 = ~n14616 & ~n29177 ;
  assign n29179 = n2244 & ~n29178 ;
  assign n29180 = ~n2332 & ~n4961 ;
  assign n29181 = n11427 & ~n29180 ;
  assign n29182 = \P1_InstAddrPointer_reg[9]/NET0131  & ~n29181 ;
  assign n29183 = ~n2402 & n4499 ;
  assign n29176 = ~n2271 & n4871 ;
  assign n29184 = n2397 & n14602 ;
  assign n29185 = ~n29176 & ~n29184 ;
  assign n29186 = ~n29183 & n29185 ;
  assign n29187 = ~n29182 & n29186 ;
  assign n29188 = ~n14607 & n29187 ;
  assign n29189 = ~n29179 & n29188 ;
  assign n29190 = n2432 & ~n29189 ;
  assign n29175 = \P1_InstAddrPointer_reg[9]/NET0131  & ~n5098 ;
  assign n29191 = ~n14629 & ~n29175 ;
  assign n29192 = ~n29190 & n29191 ;
  assign n29193 = \P2_InstAddrPointer_reg[27]/NET0131  & n1897 ;
  assign n29194 = ~n10987 & ~n29193 ;
  assign n29195 = n1734 & ~n29194 ;
  assign n29196 = n1870 & n6778 ;
  assign n29198 = n10237 & ~n16941 ;
  assign n29202 = ~n1811 & ~n29198 ;
  assign n29203 = ~n1852 & n1903 ;
  assign n29204 = ~n10235 & n29203 ;
  assign n29205 = ~n29202 & n29204 ;
  assign n29206 = \P2_InstAddrPointer_reg[27]/NET0131  & ~n29205 ;
  assign n29197 = ~n1771 & n6576 ;
  assign n29199 = n1811 & ~n29198 ;
  assign n29200 = ~n1739 & ~n29199 ;
  assign n29201 = n6676 & ~n29200 ;
  assign n29207 = ~n29197 & ~n29201 ;
  assign n29208 = ~n29206 & n29207 ;
  assign n29209 = ~n29196 & n29208 ;
  assign n29210 = ~n10994 & n29209 ;
  assign n29211 = ~n29195 & n29210 ;
  assign n29212 = n1927 & ~n29211 ;
  assign n29213 = \P2_InstAddrPointer_reg[27]/NET0131  & ~n6810 ;
  assign n29214 = ~n11008 & ~n29213 ;
  assign n29215 = ~n29212 & n29214 ;
  assign n29218 = \P3_InstAddrPointer_reg[16]/NET0131  & n2896 ;
  assign n29219 = ~n13158 & ~n29218 ;
  assign n29220 = n2894 & ~n29219 ;
  assign n29216 = ~n2841 & n13162 ;
  assign n29222 = n4402 & ~n29216 ;
  assign n29223 = \P3_InstAddrPointer_reg[16]/NET0131  & ~n29222 ;
  assign n29224 = ~n2777 & n4237 ;
  assign n29217 = n2847 & n29216 ;
  assign n29221 = ~n2923 & n4079 ;
  assign n29225 = ~n29217 & ~n29221 ;
  assign n29226 = ~n29224 & n29225 ;
  assign n29227 = ~n29223 & n29226 ;
  assign n29228 = ~n13166 & n29227 ;
  assign n29229 = ~n29220 & n29228 ;
  assign n29230 = n2453 & ~n29229 ;
  assign n29231 = \P3_InstAddrPointer_reg[16]/NET0131  & ~n4418 ;
  assign n29232 = ~n13148 & ~n29231 ;
  assign n29233 = ~n29230 & n29232 ;
  assign n29239 = \P3_InstAddrPointer_reg[27]/NET0131  & n2896 ;
  assign n29240 = ~n11146 & ~n29239 ;
  assign n29241 = n2894 & ~n29240 ;
  assign n29238 = n2918 & n4388 ;
  assign n29237 = \P3_InstAddrPointer_reg[27]/NET0131  & ~n4402 ;
  assign n29235 = ~n2777 & n4139 ;
  assign n29236 = ~n2923 & n4112 ;
  assign n29242 = ~n29235 & ~n29236 ;
  assign n29243 = ~n29237 & n29242 ;
  assign n29244 = ~n29238 & n29243 ;
  assign n29245 = ~n11154 & n29244 ;
  assign n29246 = ~n29241 & n29245 ;
  assign n29247 = n2453 & ~n29246 ;
  assign n29234 = \P3_InstAddrPointer_reg[27]/NET0131  & ~n4418 ;
  assign n29248 = ~n11164 & ~n29234 ;
  assign n29249 = ~n29247 & n29248 ;
  assign n29250 = \P2_InstAddrPointer_reg[28]/NET0131  & n1897 ;
  assign n29251 = ~n11032 & ~n29250 ;
  assign n29252 = n1734 & ~n29251 ;
  assign n29254 = ~\P2_InstAddrPointer_reg[28]/NET0131  & ~n1798 ;
  assign n29255 = ~n1727 & ~n29254 ;
  assign n29256 = n11037 & n29255 ;
  assign n29258 = \P2_InstAddrPointer_reg[28]/NET0131  & ~n8490 ;
  assign n29253 = ~n1831 & n11015 ;
  assign n29257 = ~n1771 & n6579 ;
  assign n29259 = ~n29253 & ~n29257 ;
  assign n29260 = ~n29258 & n29259 ;
  assign n29261 = ~n29256 & n29260 ;
  assign n29262 = ~n11055 & n29261 ;
  assign n29263 = ~n29252 & n29262 ;
  assign n29264 = n1927 & ~n29263 ;
  assign n29265 = \P2_InstAddrPointer_reg[28]/NET0131  & ~n6810 ;
  assign n29266 = ~n11065 & ~n29265 ;
  assign n29267 = ~n29264 & n29266 ;
  assign n29269 = \P1_InstAddrPointer_reg[25]/NET0131  & n2375 ;
  assign n29270 = ~n13471 & ~n29269 ;
  assign n29271 = n2244 & ~n29270 ;
  assign n29275 = \P1_InstAddrPointer_reg[25]/NET0131  & ~n6027 ;
  assign n29274 = n2397 & n5045 ;
  assign n29272 = ~n2402 & n4486 ;
  assign n29273 = ~n2271 & n4908 ;
  assign n29276 = ~n29272 & ~n29273 ;
  assign n29277 = ~n29274 & n29276 ;
  assign n29278 = ~n29275 & n29277 ;
  assign n29279 = ~n13478 & n29278 ;
  assign n29280 = ~n29271 & n29279 ;
  assign n29281 = n2432 & ~n29280 ;
  assign n29268 = \P1_InstAddrPointer_reg[25]/NET0131  & ~n5098 ;
  assign n29282 = ~n13484 & ~n29268 ;
  assign n29283 = ~n29281 & n29282 ;
  assign n29286 = \P2_InstAddrPointer_reg[16]/NET0131  & n1897 ;
  assign n29287 = ~n13613 & ~n29286 ;
  assign n29288 = n1734 & ~n29287 ;
  assign n29285 = ~n1831 & n13607 ;
  assign n29289 = n1870 & n11041 ;
  assign n29292 = ~n29285 & ~n29289 ;
  assign n29290 = \P2_InstAddrPointer_reg[16]/NET0131  & ~n12566 ;
  assign n29291 = ~n1771 & n6515 ;
  assign n29293 = ~n29290 & ~n29291 ;
  assign n29294 = n29292 & n29293 ;
  assign n29295 = ~n13619 & n29294 ;
  assign n29296 = ~n29288 & n29295 ;
  assign n29297 = n1927 & ~n29296 ;
  assign n29284 = \P2_InstAddrPointer_reg[16]/NET0131  & ~n6810 ;
  assign n29298 = ~n13601 & ~n29284 ;
  assign n29299 = ~n29297 & n29298 ;
  assign n29300 = \P3_InstAddrPointer_reg[24]/NET0131  & n2896 ;
  assign n29301 = ~n12096 & ~n29300 ;
  assign n29302 = n2894 & ~n29301 ;
  assign n29303 = n2918 & n12083 ;
  assign n29304 = ~n2923 & n6097 ;
  assign n29307 = ~n29303 & ~n29304 ;
  assign n29305 = \P3_InstAddrPointer_reg[24]/NET0131  & ~n4402 ;
  assign n29306 = ~n2777 & n4263 ;
  assign n29308 = ~n29305 & ~n29306 ;
  assign n29309 = n29307 & n29308 ;
  assign n29310 = ~n12087 & n29309 ;
  assign n29311 = ~n29302 & n29310 ;
  assign n29312 = n2453 & ~n29311 ;
  assign n29313 = \P3_InstAddrPointer_reg[24]/NET0131  & ~n4418 ;
  assign n29314 = ~n12110 & ~n29313 ;
  assign n29315 = ~n29312 & n29314 ;
  assign n29321 = \P1_InstAddrPointer_reg[11]/NET0131  & n2375 ;
  assign n29322 = ~n12171 & ~n29321 ;
  assign n29323 = n2244 & ~n29322 ;
  assign n29318 = ~n2402 & n4780 ;
  assign n29317 = \P1_InstAddrPointer_reg[11]/NET0131  & ~n11427 ;
  assign n29319 = n2397 & n5026 ;
  assign n29320 = ~n2271 & n4878 ;
  assign n29324 = ~n29319 & ~n29320 ;
  assign n29325 = ~n29317 & n29324 ;
  assign n29326 = ~n29318 & n29325 ;
  assign n29327 = ~n12161 & n29326 ;
  assign n29328 = ~n29323 & n29327 ;
  assign n29329 = n2432 & ~n29328 ;
  assign n29316 = \P1_InstAddrPointer_reg[11]/NET0131  & ~n5098 ;
  assign n29330 = ~n12184 & ~n29316 ;
  assign n29331 = ~n29329 & n29330 ;
  assign n29332 = \P1_InstAddrPointer_reg[28]/NET0131  & n2375 ;
  assign n29333 = ~n11320 & ~n29332 ;
  assign n29334 = n2244 & ~n29333 ;
  assign n29337 = n2397 & n6018 ;
  assign n29338 = \P1_InstAddrPointer_reg[28]/NET0131  & ~n6027 ;
  assign n29335 = ~n2402 & n11314 ;
  assign n29336 = ~n2271 & n4937 ;
  assign n29339 = ~n29335 & ~n29336 ;
  assign n29340 = ~n29338 & n29339 ;
  assign n29341 = ~n29337 & n29340 ;
  assign n29342 = ~n11328 & n29341 ;
  assign n29343 = ~n29334 & n29342 ;
  assign n29344 = n2432 & ~n29343 ;
  assign n29345 = \P1_InstAddrPointer_reg[28]/NET0131  & ~n5098 ;
  assign n29346 = ~n11342 & ~n29345 ;
  assign n29347 = ~n29344 & n29346 ;
  assign n29353 = ~\P3_EBX_reg[26]/NET0131  & ~n14981 ;
  assign n29354 = n2748 & ~n17453 ;
  assign n29355 = ~n29353 & n29354 ;
  assign n29348 = \P3_EBX_reg[26]/NET0131  & ~n2847 ;
  assign n29349 = ~n16035 & ~n29348 ;
  assign n29350 = n2771 & ~n29349 ;
  assign n29351 = \P3_EBX_reg[26]/NET0131  & ~n2748 ;
  assign n29352 = ~n2771 & n29351 ;
  assign n29356 = ~n29350 & ~n29352 ;
  assign n29357 = ~n29355 & n29356 ;
  assign n29358 = n2453 & ~n29357 ;
  assign n29359 = \P3_EBX_reg[26]/NET0131  & ~n13810 ;
  assign n29360 = ~n29358 & ~n29359 ;
  assign n29361 = \P2_InstAddrPointer_reg[24]/NET0131  & n1897 ;
  assign n29362 = ~n11918 & ~n29361 ;
  assign n29363 = n1734 & ~n29362 ;
  assign n29365 = n1870 & n7625 ;
  assign n29367 = ~n1831 & n11911 ;
  assign n29364 = ~n1771 & n6560 ;
  assign n29366 = \P2_InstAddrPointer_reg[24]/NET0131  & ~n7501 ;
  assign n29368 = ~n29364 & ~n29366 ;
  assign n29369 = ~n29367 & n29368 ;
  assign n29370 = ~n29365 & n29369 ;
  assign n29371 = ~n11926 & n29370 ;
  assign n29372 = ~n29363 & n29371 ;
  assign n29373 = n1927 & ~n29372 ;
  assign n29374 = \P2_InstAddrPointer_reg[24]/NET0131  & ~n6810 ;
  assign n29375 = ~n11937 & ~n29374 ;
  assign n29376 = ~n29373 & n29375 ;
  assign n29379 = \P1_InstAddrPointer_reg[13]/NET0131  & n2375 ;
  assign n29380 = ~n13306 & ~n29379 ;
  assign n29381 = n2244 & ~n29380 ;
  assign n29383 = \P1_InstAddrPointer_reg[13]/NET0131  & ~n11427 ;
  assign n29382 = ~n2402 & n4788 ;
  assign n29378 = ~n2271 & n4882 ;
  assign n29384 = n2397 & n13292 ;
  assign n29385 = ~n29378 & ~n29384 ;
  assign n29386 = ~n29382 & n29385 ;
  assign n29387 = ~n29383 & n29386 ;
  assign n29388 = ~n13297 & n29387 ;
  assign n29389 = ~n29381 & n29388 ;
  assign n29390 = n2432 & ~n29389 ;
  assign n29377 = \P1_InstAddrPointer_reg[13]/NET0131  & ~n5098 ;
  assign n29391 = ~n13320 & ~n29377 ;
  assign n29392 = ~n29390 & n29391 ;
  assign n29393 = \P1_InstAddrPointer_reg[15]/NET0131  & n2375 ;
  assign n29394 = ~n12207 & ~n29393 ;
  assign n29395 = n2244 & ~n29394 ;
  assign n29397 = ~n2332 & ~n5029 ;
  assign n29398 = n11427 & ~n29397 ;
  assign n29399 = \P1_InstAddrPointer_reg[15]/NET0131  & ~n29398 ;
  assign n29401 = ~n2402 & n12199 ;
  assign n29396 = ~n2271 & n4913 ;
  assign n29400 = n2397 & n6007 ;
  assign n29402 = ~n29396 & ~n29400 ;
  assign n29403 = ~n29401 & n29402 ;
  assign n29404 = ~n29399 & n29403 ;
  assign n29405 = ~n12193 & n29404 ;
  assign n29406 = ~n29395 & n29405 ;
  assign n29407 = n2432 & ~n29406 ;
  assign n29408 = \P1_InstAddrPointer_reg[15]/NET0131  & ~n5098 ;
  assign n29409 = ~n12224 & ~n29408 ;
  assign n29410 = ~n29407 & n29409 ;
  assign n29415 = ~\P1_EBX_reg[27]/NET0131  & ~n15389 ;
  assign n29416 = n24889 & ~n29415 ;
  assign n29411 = ~n15264 & n15295 ;
  assign n29412 = n2337 & ~n15296 ;
  assign n29413 = ~n29411 & n29412 ;
  assign n29414 = n2242 & n29413 ;
  assign n29417 = \P1_EBX_reg[27]/NET0131  & ~n15073 ;
  assign n29418 = ~n29414 & ~n29417 ;
  assign n29419 = ~n29416 & n29418 ;
  assign n29420 = n2432 & ~n29419 ;
  assign n29421 = \P1_EBX_reg[27]/NET0131  & ~n15402 ;
  assign n29422 = ~n29420 & ~n29421 ;
  assign n29425 = \P2_InstAddrPointer_reg[17]/NET0131  & n1897 ;
  assign n29426 = ~n13646 & ~n29425 ;
  assign n29427 = n1734 & ~n29426 ;
  assign n29428 = ~n1805 & n6660 ;
  assign n29429 = \P2_InstAddrPointer_reg[17]/NET0131  & n1805 ;
  assign n29430 = ~n29428 & ~n29429 ;
  assign n29431 = ~n1810 & n29430 ;
  assign n29432 = n1803 & ~n29431 ;
  assign n29433 = n29204 & ~n29432 ;
  assign n29434 = \P2_InstAddrPointer_reg[17]/NET0131  & ~n29433 ;
  assign n29437 = ~n1727 & ~n8492 ;
  assign n29438 = n6757 & n29437 ;
  assign n29435 = ~n1771 & n6524 ;
  assign n29424 = n1739 & n6660 ;
  assign n29436 = n1845 & ~n29430 ;
  assign n29439 = ~n29424 & ~n29436 ;
  assign n29440 = ~n29435 & n29439 ;
  assign n29441 = ~n29438 & n29440 ;
  assign n29442 = ~n29434 & n29441 ;
  assign n29443 = ~n13654 & n29442 ;
  assign n29444 = ~n29427 & n29443 ;
  assign n29445 = n1927 & ~n29444 ;
  assign n29423 = \P2_InstAddrPointer_reg[17]/NET0131  & ~n6810 ;
  assign n29446 = ~n13668 & ~n29423 ;
  assign n29447 = ~n29445 & n29446 ;
  assign n29448 = ~\P1_EBX_reg[30]/NET0131  & ~n18026 ;
  assign n29449 = n2262 & ~n15393 ;
  assign n29450 = ~n29448 & n29449 ;
  assign n29451 = ~n15105 & ~n15360 ;
  assign n29452 = n15105 & n15360 ;
  assign n29453 = ~n29451 & ~n29452 ;
  assign n29454 = n2337 & ~n29453 ;
  assign n29455 = n2242 & n29454 ;
  assign n29456 = \P1_EBX_reg[30]/NET0131  & ~n15073 ;
  assign n29457 = ~n29455 & ~n29456 ;
  assign n29458 = ~n29450 & n29457 ;
  assign n29459 = n2432 & ~n29458 ;
  assign n29460 = \P1_EBX_reg[30]/NET0131  & ~n15402 ;
  assign n29461 = ~n29459 & ~n29460 ;
  assign n29462 = \P1_EAX_reg[27]/NET0131  & ~n15402 ;
  assign n29471 = n15918 & n15998 ;
  assign n29472 = ~\P1_EAX_reg[27]/NET0131  & ~n29471 ;
  assign n29473 = n2260 & ~n16319 ;
  assign n29474 = ~n29472 & n29473 ;
  assign n29466 = \P1_EAX_reg[27]/NET0131  & ~n15924 ;
  assign n29467 = n2331 & n29413 ;
  assign n29463 = \P1_EAX_reg[27]/NET0131  & ~n2377 ;
  assign n29464 = ~n17978 & ~n29463 ;
  assign n29465 = n2222 & ~n29464 ;
  assign n29468 = n2377 & ~n5263 ;
  assign n29469 = ~n29463 & ~n29468 ;
  assign n29470 = n2302 & ~n29469 ;
  assign n29475 = ~n29465 & ~n29470 ;
  assign n29476 = ~n29467 & n29475 ;
  assign n29477 = ~n29466 & n29476 ;
  assign n29478 = ~n29474 & n29477 ;
  assign n29479 = n2432 & ~n29478 ;
  assign n29480 = ~n29462 & ~n29479 ;
  assign n29482 = \P2_InstAddrPointer_reg[23]/NET0131  & n1897 ;
  assign n29483 = ~n10947 & ~n29482 ;
  assign n29484 = n1734 & ~n29483 ;
  assign n29488 = ~n1798 & n6769 ;
  assign n29489 = ~n1727 & ~n29488 ;
  assign n29490 = n7623 & n29489 ;
  assign n29487 = ~n1831 & n10932 ;
  assign n29485 = \P2_InstAddrPointer_reg[23]/NET0131  & ~n7501 ;
  assign n29486 = ~n1771 & n6554 ;
  assign n29491 = ~n29485 & ~n29486 ;
  assign n29492 = ~n29487 & n29491 ;
  assign n29493 = ~n29490 & n29492 ;
  assign n29494 = ~n10954 & n29493 ;
  assign n29495 = ~n29484 & n29494 ;
  assign n29496 = n1927 & ~n29495 ;
  assign n29481 = \P2_InstAddrPointer_reg[23]/NET0131  & ~n6810 ;
  assign n29497 = ~n10958 & ~n29481 ;
  assign n29498 = ~n29496 & n29497 ;
  assign n29501 = \P1_InstAddrPointer_reg[14]/NET0131  & n2375 ;
  assign n29502 = ~n13340 & ~n29501 ;
  assign n29503 = n2244 & ~n29502 ;
  assign n29506 = ~n2402 & n13335 ;
  assign n29500 = \P1_InstAddrPointer_reg[14]/NET0131  & ~n11427 ;
  assign n29504 = ~n2271 & n4931 ;
  assign n29505 = n2397 & n5034 ;
  assign n29507 = ~n29504 & ~n29505 ;
  assign n29508 = ~n29500 & n29507 ;
  assign n29509 = ~n29506 & n29508 ;
  assign n29510 = ~n13328 & n29509 ;
  assign n29511 = ~n29503 & n29510 ;
  assign n29512 = n2432 & ~n29511 ;
  assign n29499 = \P1_InstAddrPointer_reg[14]/NET0131  & ~n5098 ;
  assign n29513 = ~n13353 & ~n29499 ;
  assign n29514 = ~n29512 & n29513 ;
  assign n29517 = \P1_InstAddrPointer_reg[21]/NET0131  & n2375 ;
  assign n29518 = ~n13452 & ~n29517 ;
  assign n29519 = n2244 & ~n29518 ;
  assign n29520 = \P1_InstAddrPointer_reg[21]/NET0131  & n7308 ;
  assign n29521 = n2402 & ~n29520 ;
  assign n29522 = n4769 & ~n29521 ;
  assign n29524 = n2397 & n13439 ;
  assign n29516 = ~n2271 & n4900 ;
  assign n29523 = \P1_InstAddrPointer_reg[21]/NET0131  & ~n11427 ;
  assign n29525 = ~n29516 & ~n29523 ;
  assign n29526 = ~n29524 & n29525 ;
  assign n29527 = ~n29522 & n29526 ;
  assign n29528 = ~n13442 & n29527 ;
  assign n29529 = ~n29519 & n29528 ;
  assign n29530 = n2432 & ~n29529 ;
  assign n29515 = \P1_InstAddrPointer_reg[21]/NET0131  & ~n5098 ;
  assign n29531 = ~n13433 & ~n29515 ;
  assign n29532 = ~n29530 & n29531 ;
  assign n29537 = \P2_InstAddrPointer_reg[8]/NET0131  & n1897 ;
  assign n29538 = ~n13027 & ~n29537 ;
  assign n29539 = n1734 & ~n29538 ;
  assign n29534 = n1798 & ~n6736 ;
  assign n29535 = ~n1727 & ~n29534 ;
  assign n29536 = n1798 & n29535 ;
  assign n29540 = ~n1771 & n6459 ;
  assign n29545 = ~n29536 & ~n29540 ;
  assign n29541 = ~n1831 & n6603 ;
  assign n29542 = ~n1892 & ~n29535 ;
  assign n29543 = n7637 & n29542 ;
  assign n29544 = \P2_InstAddrPointer_reg[8]/NET0131  & ~n29543 ;
  assign n29546 = ~n29541 & ~n29544 ;
  assign n29547 = n29545 & n29546 ;
  assign n29548 = ~n13035 & n29547 ;
  assign n29549 = ~n29539 & n29548 ;
  assign n29550 = n1927 & ~n29549 ;
  assign n29533 = \P2_InstAddrPointer_reg[8]/NET0131  & ~n6810 ;
  assign n29551 = ~n13049 & ~n29533 ;
  assign n29552 = ~n29550 & n29551 ;
  assign n29554 = \P1_InstAddrPointer_reg[22]/NET0131  & n2375 ;
  assign n29555 = ~n12298 & ~n29554 ;
  assign n29556 = n2244 & ~n29555 ;
  assign n29558 = \P1_InstAddrPointer_reg[22]/NET0131  & ~n7316 ;
  assign n29559 = n2397 & n5049 ;
  assign n29564 = ~n2271 & n4902 ;
  assign n29557 = n2237 & n4476 ;
  assign n29560 = ~\P1_InstAddrPointer_reg[22]/NET0131  & n2317 ;
  assign n29561 = ~n2317 & ~n4476 ;
  assign n29562 = ~n29560 & ~n29561 ;
  assign n29563 = ~n2314 & n29562 ;
  assign n29565 = ~n29557 & ~n29563 ;
  assign n29566 = ~n29564 & n29565 ;
  assign n29567 = ~n29559 & n29566 ;
  assign n29568 = ~n29558 & n29567 ;
  assign n29569 = ~n12305 & n29568 ;
  assign n29570 = ~n29556 & n29569 ;
  assign n29571 = n2432 & ~n29570 ;
  assign n29553 = \P1_InstAddrPointer_reg[22]/NET0131  & ~n5098 ;
  assign n29572 = ~n12315 & ~n29553 ;
  assign n29573 = ~n29571 & n29572 ;
  assign n29576 = \P3_InstAddrPointer_reg[11]/NET0131  & n2896 ;
  assign n29577 = ~n11976 & ~n29576 ;
  assign n29578 = n2894 & ~n29577 ;
  assign n29575 = n2918 & n11980 ;
  assign n29579 = ~n2923 & n4069 ;
  assign n29582 = ~n29575 & ~n29579 ;
  assign n29580 = \P3_InstAddrPointer_reg[11]/NET0131  & ~n4402 ;
  assign n29581 = ~n2777 & n4158 ;
  assign n29583 = ~n29580 & ~n29581 ;
  assign n29584 = n29582 & n29583 ;
  assign n29585 = ~n11984 & n29584 ;
  assign n29586 = ~n29578 & n29585 ;
  assign n29587 = n2453 & ~n29586 ;
  assign n29574 = \P3_InstAddrPointer_reg[11]/NET0131  & ~n4418 ;
  assign n29588 = ~n11994 & ~n29574 ;
  assign n29589 = ~n29587 & n29588 ;
  assign n29592 = ~\P3_EBX_reg[25]/NET0131  & ~n14980 ;
  assign n29593 = n2748 & ~n14981 ;
  assign n29594 = ~n29592 & n29593 ;
  assign n29590 = \P3_EBX_reg[25]/NET0131  & n14954 ;
  assign n29591 = n14952 & n21771 ;
  assign n29595 = ~n29590 & ~n29591 ;
  assign n29596 = ~n29594 & n29595 ;
  assign n29597 = n2453 & ~n29596 ;
  assign n29598 = \P3_EBX_reg[25]/NET0131  & ~n13810 ;
  assign n29599 = ~n29597 & ~n29598 ;
  assign n29601 = \P1_InstAddrPointer_reg[19]/NET0131  & n2375 ;
  assign n29602 = ~n12256 & ~n29601 ;
  assign n29603 = n2244 & ~n29602 ;
  assign n29604 = ~n2402 & n6846 ;
  assign n29600 = \P1_InstAddrPointer_reg[19]/NET0131  & ~n11427 ;
  assign n29605 = n2397 & n4973 ;
  assign n29606 = ~n2271 & n4926 ;
  assign n29607 = ~n29605 & ~n29606 ;
  assign n29608 = ~n29600 & n29607 ;
  assign n29609 = ~n29604 & n29608 ;
  assign n29610 = ~n12246 & n29609 ;
  assign n29611 = ~n29603 & n29610 ;
  assign n29612 = n2432 & ~n29611 ;
  assign n29613 = \P1_InstAddrPointer_reg[19]/NET0131  & ~n5098 ;
  assign n29614 = ~n12236 & ~n29613 ;
  assign n29615 = ~n29612 & n29614 ;
  assign n29618 = \P1_InstAddrPointer_reg[16]/NET0131  & n2375 ;
  assign n29619 = ~n13376 & ~n29618 ;
  assign n29620 = n2244 & ~n29619 ;
  assign n29623 = ~n2402 & n4784 ;
  assign n29622 = \P1_InstAddrPointer_reg[16]/NET0131  & ~n11427 ;
  assign n29617 = n2397 & n5032 ;
  assign n29621 = ~n2271 & n4918 ;
  assign n29624 = ~n29617 & ~n29621 ;
  assign n29625 = ~n29622 & n29624 ;
  assign n29626 = ~n29623 & n29625 ;
  assign n29627 = ~n13365 & n29626 ;
  assign n29628 = ~n29620 & n29627 ;
  assign n29629 = n2432 & ~n29628 ;
  assign n29616 = \P1_InstAddrPointer_reg[16]/NET0131  & ~n5098 ;
  assign n29630 = ~n13388 & ~n29616 ;
  assign n29631 = ~n29629 & n29630 ;
  assign n29632 = \P1_PhyAddrPointer_reg[31]/NET0131  & n2375 ;
  assign n29633 = ~n29034 & ~n29632 ;
  assign n29634 = n2244 & ~n29633 ;
  assign n29635 = \P1_PhyAddrPointer_reg[31]/NET0131  & ~n10087 ;
  assign n29636 = ~n29044 & ~n29635 ;
  assign n29637 = ~n29634 & n29636 ;
  assign n29638 = n2432 & ~n29637 ;
  assign n29639 = n10133 & n18540 ;
  assign n29641 = \P1_PhyAddrPointer_reg[31]/NET0131  & n10119 ;
  assign n29640 = ~\P1_PhyAddrPointer_reg[31]/NET0131  & ~n10119 ;
  assign n29642 = n3148 & ~n29640 ;
  assign n29643 = ~n29641 & n29642 ;
  assign n29644 = \P1_PhyAddrPointer_reg[31]/NET0131  & ~n10136 ;
  assign n29645 = ~n29057 & ~n29644 ;
  assign n29646 = ~n29643 & n29645 ;
  assign n29647 = ~n29639 & n29646 ;
  assign n29648 = ~n29638 & n29647 ;
  assign n29649 = \P3_PhyAddrPointer_reg[17]/NET0131  & n2896 ;
  assign n29650 = ~n29090 & ~n29649 ;
  assign n29651 = n2894 & ~n29650 ;
  assign n29652 = \P3_PhyAddrPointer_reg[17]/NET0131  & ~n9014 ;
  assign n29653 = ~n29099 & ~n29652 ;
  assign n29654 = ~n29651 & n29653 ;
  assign n29655 = n2453 & ~n29654 ;
  assign n29660 = n4415 & n20674 ;
  assign n29656 = n9032 & n12000 ;
  assign n29657 = ~\P3_PhyAddrPointer_reg[17]/NET0131  & ~n29656 ;
  assign n29658 = n2959 & ~n13221 ;
  assign n29659 = ~n29657 & n29658 ;
  assign n29661 = \P3_PhyAddrPointer_reg[17]/NET0131  & ~n9063 ;
  assign n29662 = ~n29077 & ~n29661 ;
  assign n29663 = ~n29659 & n29662 ;
  assign n29664 = ~n29660 & n29663 ;
  assign n29665 = ~n29655 & n29664 ;
  assign n29668 = \P1_InstAddrPointer_reg[7]/NET0131  & n2375 ;
  assign n29669 = ~n14577 & ~n29668 ;
  assign n29670 = n2244 & ~n29669 ;
  assign n29671 = ~n2332 & ~n4960 ;
  assign n29672 = n11427 & ~n29671 ;
  assign n29673 = \P1_InstAddrPointer_reg[7]/NET0131  & ~n29672 ;
  assign n29667 = ~n2402 & n4504 ;
  assign n29674 = ~n2271 & n4826 ;
  assign n29675 = n2397 & n4979 ;
  assign n29676 = ~n29674 & ~n29675 ;
  assign n29677 = ~n29667 & n29676 ;
  assign n29678 = ~n29673 & n29677 ;
  assign n29679 = ~n14567 & n29678 ;
  assign n29680 = ~n29670 & n29679 ;
  assign n29681 = n2432 & ~n29680 ;
  assign n29666 = \P1_InstAddrPointer_reg[7]/NET0131  & ~n5098 ;
  assign n29682 = ~n14592 & ~n29666 ;
  assign n29683 = ~n29681 & n29682 ;
  assign n29684 = \P2_EBX_reg[30]/NET0131  & ~n12632 ;
  assign n29687 = ~\P2_EBX_reg[30]/NET0131  & ~n15061 ;
  assign n29688 = n1766 & ~n15062 ;
  assign n29689 = ~n29687 & n29688 ;
  assign n29685 = \P2_EBX_reg[30]/NET0131  & ~n15019 ;
  assign n29686 = n1722 & n15004 ;
  assign n29690 = ~n29685 & ~n29686 ;
  assign n29691 = ~n29689 & n29690 ;
  assign n29692 = n1927 & ~n29691 ;
  assign n29693 = ~n29684 & ~n29692 ;
  assign n29696 = \P1_EAX_reg[30]/NET0131  & n16321 ;
  assign n29695 = ~\P1_EAX_reg[30]/NET0131  & ~n16321 ;
  assign n29697 = n2260 & ~n29695 ;
  assign n29698 = ~n29696 & n29697 ;
  assign n29699 = n2331 & n29454 ;
  assign n29694 = \P1_EAX_reg[30]/NET0131  & ~n15925 ;
  assign n29700 = n2222 & ~n5191 ;
  assign n29701 = n2302 & ~n6912 ;
  assign n29702 = ~n29700 & ~n29701 ;
  assign n29703 = n2377 & ~n29702 ;
  assign n29704 = ~n29694 & ~n29703 ;
  assign n29705 = ~n29699 & n29704 ;
  assign n29706 = ~n29698 & n29705 ;
  assign n29707 = n2432 & ~n29706 ;
  assign n29708 = \P1_EAX_reg[30]/NET0131  & ~n15402 ;
  assign n29709 = ~n29707 & ~n29708 ;
  assign n29712 = \P1_InstAddrPointer_reg[8]/NET0131  & n2375 ;
  assign n29713 = ~n13510 & ~n29712 ;
  assign n29714 = n2244 & ~n29713 ;
  assign n29717 = ~n2402 & n4502 ;
  assign n29711 = \P1_InstAddrPointer_reg[8]/NET0131  & ~n11427 ;
  assign n29715 = ~n2271 & n4869 ;
  assign n29716 = n2397 & n4977 ;
  assign n29718 = ~n29715 & ~n29716 ;
  assign n29719 = ~n29711 & n29718 ;
  assign n29720 = ~n29717 & n29719 ;
  assign n29721 = ~n13498 & n29720 ;
  assign n29722 = ~n29714 & n29721 ;
  assign n29723 = n2432 & ~n29722 ;
  assign n29710 = \P1_InstAddrPointer_reg[8]/NET0131  & ~n5098 ;
  assign n29724 = ~n13523 & ~n29710 ;
  assign n29725 = ~n29723 & n29724 ;
  assign n29726 = \P2_uWord_reg[13]/NET0131  & ~n15942 ;
  assign n29727 = \P2_uWord_reg[13]/NET0131  & ~n15982 ;
  assign n29728 = n1742 & n17689 ;
  assign n29729 = ~n29727 & ~n29728 ;
  assign n29730 = ~n25916 & n29729 ;
  assign n29731 = n1927 & ~n29730 ;
  assign n29732 = ~n29726 & ~n29731 ;
  assign n29733 = \P2_EAX_reg[7]/NET0131  & ~n17439 ;
  assign n29734 = ~n3128 & n14771 ;
  assign n29735 = n1726 & n25072 ;
  assign n29736 = ~\P2_EAX_reg[7]/NET0131  & ~n12639 ;
  assign n29737 = ~n12640 & ~n29736 ;
  assign n29738 = n12664 & n29737 ;
  assign n29739 = ~n29735 & ~n29738 ;
  assign n29740 = ~n29734 & n29739 ;
  assign n29741 = n1927 & ~n29740 ;
  assign n29742 = ~n29733 & ~n29741 ;
  assign n29747 = n2847 & ~n4315 ;
  assign n29748 = ~\P3_InstAddrPointer_reg[4]/NET0131  & ~n2847 ;
  assign n29749 = ~n29747 & ~n29748 ;
  assign n29750 = ~n2841 & n29749 ;
  assign n29752 = n15796 & ~n29750 ;
  assign n29751 = ~n2777 & n4201 ;
  assign n29744 = ~n2923 & n3969 ;
  assign n29745 = ~n2897 & n12505 ;
  assign n29746 = \P3_InstAddrPointer_reg[4]/NET0131  & ~n29745 ;
  assign n29753 = ~n29744 & ~n29746 ;
  assign n29754 = ~n29751 & n29753 ;
  assign n29755 = n29752 & n29754 ;
  assign n29756 = n2453 & ~n29755 ;
  assign n29743 = \P3_InstAddrPointer_reg[4]/NET0131  & ~n4418 ;
  assign n29757 = ~n15809 & ~n29743 ;
  assign n29758 = ~n29756 & n29757 ;
  assign n29760 = \P3_PhyAddrPointer_reg[19]/NET0131  & n2896 ;
  assign n29761 = ~n28945 & ~n29760 ;
  assign n29762 = n2894 & ~n29761 ;
  assign n29763 = \P3_PhyAddrPointer_reg[19]/NET0131  & ~n9014 ;
  assign n29764 = ~n28958 & ~n29763 ;
  assign n29765 = ~n29762 & n29764 ;
  assign n29766 = n2453 & ~n29765 ;
  assign n29767 = ~\P3_DataWidth_reg[1]/NET0131  & ~n20754 ;
  assign n29768 = ~\P3_PhyAddrPointer_reg[19]/NET0131  & ~n13194 ;
  assign n29769 = ~n12048 & ~n29768 ;
  assign n29770 = \P3_DataWidth_reg[1]/NET0131  & ~n29769 ;
  assign n29771 = n2959 & ~n29770 ;
  assign n29772 = ~n29767 & n29771 ;
  assign n29759 = n4415 & n20754 ;
  assign n29773 = \P3_PhyAddrPointer_reg[19]/NET0131  & ~n9063 ;
  assign n29774 = ~n28936 & ~n29773 ;
  assign n29775 = ~n29759 & n29774 ;
  assign n29776 = ~n29772 & n29775 ;
  assign n29777 = ~n29766 & n29776 ;
  assign n29778 = \P1_EAX_reg[31]/NET0131  & ~n15402 ;
  assign n29780 = \P1_EAX_reg[31]/NET0131  & n29696 ;
  assign n29779 = ~\P1_EAX_reg[31]/NET0131  & ~n29696 ;
  assign n29781 = n2260 & ~n29779 ;
  assign n29782 = ~n29780 & n29781 ;
  assign n29783 = \P1_EAX_reg[31]/NET0131  & ~n15925 ;
  assign n29784 = n2331 & n15362 ;
  assign n29785 = n5155 & n15893 ;
  assign n29786 = ~n29784 & ~n29785 ;
  assign n29787 = ~n29783 & n29786 ;
  assign n29788 = ~n29782 & n29787 ;
  assign n29789 = n2432 & ~n29788 ;
  assign n29790 = ~n29778 & ~n29789 ;
  assign n29793 = \P2_InstAddrPointer_reg[21]/NET0131  & n1897 ;
  assign n29794 = ~n12979 & ~n29793 ;
  assign n29795 = n1734 & ~n29794 ;
  assign n29792 = \P2_InstAddrPointer_reg[21]/NET0131  & ~n12566 ;
  assign n29796 = n1870 & n6766 ;
  assign n29799 = ~n29792 & ~n29796 ;
  assign n29797 = ~n1831 & n6595 ;
  assign n29798 = ~n1771 & n6546 ;
  assign n29800 = ~n29797 & ~n29798 ;
  assign n29801 = n29799 & n29800 ;
  assign n29802 = ~n12985 & n29801 ;
  assign n29803 = ~n29795 & n29802 ;
  assign n29804 = n1927 & ~n29803 ;
  assign n29791 = \P2_InstAddrPointer_reg[21]/NET0131  & ~n6810 ;
  assign n29805 = ~n12994 & ~n29791 ;
  assign n29806 = ~n29804 & n29805 ;
  assign \_al_n0  = 1'b0 ;
  assign \_al_n1  = ~1'b0 ;
  assign \address2[0]_pad  = ~n1353 ;
  assign \address2[10]_pad  = ~n1356 ;
  assign \address2[11]_pad  = ~n1359 ;
  assign \address2[12]_pad  = ~n1362 ;
  assign \address2[13]_pad  = ~n1365 ;
  assign \address2[14]_pad  = ~n1368 ;
  assign \address2[15]_pad  = ~n1371 ;
  assign \address2[16]_pad  = ~n1374 ;
  assign \address2[17]_pad  = ~n1377 ;
  assign \address2[18]_pad  = ~n1380 ;
  assign \address2[19]_pad  = ~n1383 ;
  assign \address2[1]_pad  = ~n1386 ;
  assign \address2[20]_pad  = ~n1389 ;
  assign \address2[21]_pad  = ~n1392 ;
  assign \address2[22]_pad  = ~n1395 ;
  assign \address2[23]_pad  = ~n1398 ;
  assign \address2[24]_pad  = ~n1401 ;
  assign \address2[25]_pad  = ~n1404 ;
  assign \address2[26]_pad  = ~n1407 ;
  assign \address2[27]_pad  = ~n1410 ;
  assign \address2[28]_pad  = ~n1413 ;
  assign \address2[29]_pad  = ~n1416 ;
  assign \address2[2]_pad  = ~n1419 ;
  assign \address2[3]_pad  = ~n1422 ;
  assign \address2[4]_pad  = ~n1425 ;
  assign \address2[5]_pad  = ~n1428 ;
  assign \address2[6]_pad  = ~n1431 ;
  assign \address2[7]_pad  = ~n1434 ;
  assign \address2[8]_pad  = ~n1437 ;
  assign \address2[9]_pad  = ~n1440 ;
  assign \g133468/_2_  = ~n1943 ;
  assign \g133469/_2_  = ~n2450 ;
  assign \g133470/_2_  = ~n2967 ;
  assign \g133475/_0_  = ~n2973 ;
  assign \g133476/_2_  = ~n2992 ;
  assign \g133515/_0_  = ~n2998 ;
  assign \g133516/_0_  = ~n3014 ;
  assign \g133517/_0_  = ~n3033 ;
  assign \g133518/_0_  = ~n3039 ;
  assign \g133523/_0_  = ~n3041 ;
  assign \g133524/_0_  = ~n3043 ;
  assign \g133528/_0_  = ~n3122 ;
  assign \g133529/_0_  = ~n3145 ;
  assign \g133531/_0_  = ~n3151 ;
  assign \g133532/_0_  = ~n3180 ;
  assign \g133533/_0_  = ~n3196 ;
  assign \g133534/_0_  = ~n3216 ;
  assign \g133535/_0_  = ~n3235 ;
  assign \g133536/_0_  = ~n3258 ;
  assign \g133537/_0_  = ~n3274 ;
  assign \g133538/_0_  = ~n3295 ;
  assign \g133539/_0_  = ~n3311 ;
  assign \g133540/_0_  = ~n3331 ;
  assign \g133541/_0_  = ~n3347 ;
  assign \g133542/_0_  = ~n3368 ;
  assign \g133543/_0_  = ~n3384 ;
  assign \g133544/_0_  = ~n3403 ;
  assign \g133545/_0_  = ~n3422 ;
  assign \g133546/_0_  = ~n3444 ;
  assign \g133547/_0_  = ~n3460 ;
  assign \g133548/_0_  = ~n3482 ;
  assign \g133549/_0_  = ~n3498 ;
  assign \g133550/_0_  = ~n3520 ;
  assign \g133551/_0_  = ~n3536 ;
  assign \g133552/_0_  = ~n3558 ;
  assign \g133553/_0_  = ~n3574 ;
  assign \g133554/_0_  = ~n3596 ;
  assign \g133555/_0_  = ~n3612 ;
  assign \g133556/_0_  = ~n3633 ;
  assign \g133557/_0_  = ~n3649 ;
  assign \g133558/_0_  = ~n3669 ;
  assign \g133559/_0_  = ~n3685 ;
  assign \g133560/_0_  = ~n3705 ;
  assign \g133561/_0_  = ~n3721 ;
  assign \g133566/_0_  = ~n4421 ;
  assign \g133619/_0_  = ~n5101 ;
  assign \g133659/_0_  = ~n5295 ;
  assign \g133660/_0_  = ~n5323 ;
  assign \g133662/_0_  = ~n5352 ;
  assign \g133663/_0_  = ~n5375 ;
  assign \g133664/_0_  = ~n5398 ;
  assign \g133665/_0_  = ~n5419 ;
  assign \g133666/_0_  = ~n5439 ;
  assign \g133667/_0_  = ~n5460 ;
  assign \g133668/_0_  = ~n5482 ;
  assign \g133669/_0_  = ~n5505 ;
  assign \g133670/_0_  = ~n5526 ;
  assign \g133671/_0_  = ~n5548 ;
  assign \g133672/_0_  = ~n5570 ;
  assign \g133673/_0_  = ~n5592 ;
  assign \g133674/_0_  = ~n5613 ;
  assign \g133675/_0_  = ~n5633 ;
  assign \g133676/_0_  = ~n5653 ;
  assign \g133677/_0_  = ~n5672 ;
  assign \g133678/_0_  = ~n5691 ;
  assign \g133679/_0_  = ~n5710 ;
  assign \g133680/_0_  = ~n5729 ;
  assign \g133681/_0_  = ~n5748 ;
  assign \g133682/_0_  = ~n5767 ;
  assign \g133683/_0_  = ~n5786 ;
  assign \g133684/_0_  = ~n5805 ;
  assign \g133685/_0_  = ~n5824 ;
  assign \g133686/_0_  = ~n5843 ;
  assign \g133687/_0_  = ~n5862 ;
  assign \g133688/_0_  = ~n5881 ;
  assign \g133689/_0_  = ~n5900 ;
  assign \g133690/_0_  = ~n5919 ;
  assign \g133691/_0_  = ~n5938 ;
  assign \g133694/_0_  = ~n6040 ;
  assign \g133697/_0_  = ~n6154 ;
  assign \g133702/_0_  = ~n6813 ;
  assign \g133703/_0_  = ~n6905 ;
  assign \g133756/_0_  = ~n6940 ;
  assign \g133792/_0_  = ~n6959 ;
  assign \g133793/_0_  = ~n6978 ;
  assign \g133794/_0_  = ~n6997 ;
  assign \g133796/_0_  = ~n7016 ;
  assign \g133797/_0_  = ~n7035 ;
  assign \g133798/_0_  = ~n7054 ;
  assign \g133799/_0_  = ~n7073 ;
  assign \g133800/_0_  = ~n7092 ;
  assign \g133801/_0_  = ~n7111 ;
  assign \g133802/_0_  = ~n7130 ;
  assign \g133803/_0_  = ~n7149 ;
  assign \g133804/_0_  = ~n7168 ;
  assign \g133806/_0_  = ~n7187 ;
  assign \g133807/_0_  = ~n7206 ;
  assign \g133808/_0_  = ~n7225 ;
  assign \g133812/_0_  = ~n7267 ;
  assign \g133813/_0_  = ~n7327 ;
  assign \g133814/_0_  = ~n7367 ;
  assign \g133817/_0_  = ~n7415 ;
  assign \g133821/_0_  = ~n7513 ;
  assign \g133824/_0_  = ~n7584 ;
  assign \g133826/_0_  = ~n7657 ;
  assign \g133828/_0_  = ~n7696 ;
  assign \g133864/_0_  = ~n7721 ;
  assign \g133865/_0_  = ~n7749 ;
  assign \g133867/_0_  = ~n7769 ;
  assign \g133868/_0_  = ~n7789 ;
  assign \g133869/_0_  = ~n7809 ;
  assign \g133871/_0_  = ~n7829 ;
  assign \g133872/_0_  = ~n7849 ;
  assign \g133873/_0_  = ~n7869 ;
  assign \g133874/_0_  = ~n7889 ;
  assign \g133875/_0_  = ~n7909 ;
  assign \g133876/_0_  = ~n7929 ;
  assign \g133877/_0_  = ~n7949 ;
  assign \g133878/_0_  = ~n7969 ;
  assign \g133879/_0_  = ~n7989 ;
  assign \g133881/_0_  = ~n8009 ;
  assign \g133882/_0_  = ~n8029 ;
  assign \g133883/_0_  = ~n8049 ;
  assign \g133884/_0_  = ~n8068 ;
  assign \g133885/_0_  = ~n8087 ;
  assign \g133886/_0_  = ~n8106 ;
  assign \g133887/_0_  = ~n8125 ;
  assign \g133888/_0_  = ~n8144 ;
  assign \g133889/_0_  = ~n8163 ;
  assign \g133890/_0_  = ~n8182 ;
  assign \g133891/_0_  = ~n8201 ;
  assign \g133892/_0_  = ~n8220 ;
  assign \g133893/_0_  = ~n8239 ;
  assign \g133894/_0_  = ~n8258 ;
  assign \g133895/_0_  = ~n8277 ;
  assign \g133896/_0_  = ~n8296 ;
  assign \g133897/_0_  = ~n8315 ;
  assign \g133898/_0_  = ~n8334 ;
  assign \g133910/_0_  = ~n8392 ;
  assign \g133911/_0_  = ~n8433 ;
  assign \g133912/_0_  = ~n8467 ;
  assign \g133915/_0_  = ~n8505 ;
  assign \g133917/_0_  = ~n8541 ;
  assign \g133929/_0_  = ~n8586 ;
  assign \g134014/_0_  = ~n8614 ;
  assign \g134040/_0_  = ~n8633 ;
  assign \g134041/_0_  = ~n8652 ;
  assign \g134042/_0_  = ~n8671 ;
  assign \g134043/_0_  = ~n8690 ;
  assign \g134044/_0_  = ~n8709 ;
  assign \g134045/_0_  = ~n8728 ;
  assign \g134046/_0_  = ~n8747 ;
  assign \g134047/_0_  = ~n8766 ;
  assign \g134048/_0_  = ~n8785 ;
  assign \g134049/_0_  = ~n8804 ;
  assign \g134050/_0_  = ~n8823 ;
  assign \g134051/_0_  = ~n8842 ;
  assign \g134052/_0_  = ~n8861 ;
  assign \g134053/_0_  = ~n8880 ;
  assign \g134054/_0_  = ~n8899 ;
  assign \g134056/_0_  = ~n9010 ;
  assign \g134059/_0_  = ~n9068 ;
  assign \g134064/_0_  = ~n9119 ;
  assign \g134067/_0_  = ~n9158 ;
  assign \g134068/_0_  = ~n9194 ;
  assign \g134069/_0_  = ~n9222 ;
  assign \g134070/_0_  = ~n9260 ;
  assign \g134071/_0_  = ~n9291 ;
  assign \g134073/_0_  = ~n9330 ;
  assign \g134076/_0_  = ~n9377 ;
  assign \g134131/_0_  = ~n9400 ;
  assign \g134132/_0_  = ~n9423 ;
  assign \g134156/_0_  = ~n9442 ;
  assign \g134157/_0_  = ~n9461 ;
  assign \g134158/_0_  = ~n9480 ;
  assign \g134159/_0_  = ~n9499 ;
  assign \g134163/_0_  = ~n9518 ;
  assign \g134164/_0_  = ~n9537 ;
  assign \g134165/_0_  = ~n9556 ;
  assign \g134166/_0_  = ~n9575 ;
  assign \g134167/_0_  = ~n9594 ;
  assign \g134168/_0_  = ~n9613 ;
  assign \g134169/_0_  = ~n9632 ;
  assign \g134170/_0_  = ~n9651 ;
  assign \g134171/_0_  = ~n9670 ;
  assign \g134172/_0_  = ~n9689 ;
  assign \g134173/_0_  = ~n9708 ;
  assign \g134174/_0_  = ~n9727 ;
  assign \g134176/_0_  = ~n9746 ;
  assign \g134177/_0_  = ~n9765 ;
  assign \g134178/_0_  = ~n9784 ;
  assign \g134179/_0_  = ~n9803 ;
  assign \g134181/_0_  = ~n9822 ;
  assign \g134183/_0_  = ~n9841 ;
  assign \g134184/_0_  = ~n9860 ;
  assign \g134185/_0_  = ~n9879 ;
  assign \g134186/_0_  = ~n9898 ;
  assign \g134187/_0_  = ~n9917 ;
  assign \g134188/_0_  = ~n9936 ;
  assign \g134189/_0_  = ~n9955 ;
  assign \g134190/_0_  = ~n9974 ;
  assign \g134191/_0_  = ~n9993 ;
  assign \g134194/_0_  = ~n10036 ;
  assign \g134202/_0_  = ~n10083 ;
  assign \g134207/_0_  = ~n10141 ;
  assign \g134214/_0_  = ~n10172 ;
  assign \g134216/_0_  = ~n10217 ;
  assign \g134226/_0_  = ~n10261 ;
  assign \g134228/_0_  = ~n10307 ;
  assign \g134360/_0_  = ~n10330 ;
  assign \g134383/_0_  = ~n10358 ;
  assign \g134412/_0_  = ~n10377 ;
  assign \g134413/_0_  = ~n10396 ;
  assign \g134419/_0_  = ~n10415 ;
  assign \g134420/_0_  = ~n10434 ;
  assign \g134421/_0_  = ~n10453 ;
  assign \g134422/_0_  = ~n10472 ;
  assign \g134423/_0_  = ~n10491 ;
  assign \g134424/_0_  = ~n10510 ;
  assign \g134426/_0_  = ~n10529 ;
  assign \g134429/_0_  = ~n10548 ;
  assign \g134431/_0_  = ~n10567 ;
  assign \g134433/_0_  = ~n10586 ;
  assign \g134434/_0_  = ~n10605 ;
  assign \g134435/_0_  = ~n10624 ;
  assign \g134436/_0_  = ~n10643 ;
  assign \g134438/_0_  = ~n10662 ;
  assign \g134439/_0_  = ~n10681 ;
  assign \g134441/_0_  = ~n10700 ;
  assign \g134442/_0_  = ~n10719 ;
  assign \g134443/_0_  = ~n10738 ;
  assign \g134445/_0_  = ~n10757 ;
  assign \g134446/_0_  = ~n10776 ;
  assign \g134447/_0_  = ~n10795 ;
  assign \g134448/_0_  = ~n10814 ;
  assign \g134449/_0_  = ~n10833 ;
  assign \g134450/_0_  = ~n10852 ;
  assign \g134451/_0_  = ~n10871 ;
  assign \g134453/_0_  = ~n10890 ;
  assign \g134454/_0_  = ~n10909 ;
  assign \g134455/_0_  = ~n10928 ;
  assign \g134457/_0_  = ~n10974 ;
  assign \g134458/_0_  = ~n11012 ;
  assign \g134459/_0_  = ~n11070 ;
  assign \g134460/_0_  = ~n11090 ;
  assign \g134469/_0_  = ~n11135 ;
  assign \g134470/_0_  = ~n11171 ;
  assign \g134471/_0_  = ~n11191 ;
  assign \g134472/_0_  = ~n11238 ;
  assign \g134479/_0_  = ~n11260 ;
  assign \g134480/_0_  = ~n11305 ;
  assign \g134481/_0_  = ~n11347 ;
  assign \g134482/_0_  = ~n11366 ;
  assign \g134490/_0_  = ~n11406 ;
  assign \g134491/_0_  = ~n11442 ;
  assign \g134496/_0_  = ~n11467 ;
  assign \g134506/_0_  = ~n11502 ;
  assign \g134508/_0_  = ~n11538 ;
  assign \g134579/_0_  = ~n11566 ;
  assign \g134603/_0_  = ~n11585 ;
  assign \g134604/_0_  = ~n11604 ;
  assign \g134605/_0_  = ~n11623 ;
  assign \g134606/_0_  = ~n11642 ;
  assign \g134607/_0_  = ~n11661 ;
  assign \g134608/_0_  = ~n11680 ;
  assign \g134609/_0_  = ~n11699 ;
  assign \g134610/_0_  = ~n11718 ;
  assign \g134611/_0_  = ~n11737 ;
  assign \g134612/_0_  = ~n11756 ;
  assign \g134613/_0_  = ~n11775 ;
  assign \g134614/_0_  = ~n11794 ;
  assign \g134615/_0_  = ~n11813 ;
  assign \g134616/_0_  = ~n11832 ;
  assign \g134617/_0_  = ~n11851 ;
  assign \g134618/_0_  = ~n11884 ;
  assign \g134619/_0_  = ~n11904 ;
  assign \g134620/_0_  = ~n11941 ;
  assign \g134621/_0_  = ~n11959 ;
  assign \g134632/_0_  = ~n11999 ;
  assign \g134633/_0_  = ~n12025 ;
  assign \g134636/_0_  = ~n12062 ;
  assign \g134637/_0_  = ~n12081 ;
  assign \g134638/_0_  = ~n12114 ;
  assign \g134639/_0_  = ~n12149 ;
  assign \g134645/_0_  = ~n12189 ;
  assign \g134646/_0_  = ~n12229 ;
  assign \g134648/_0_  = ~n12266 ;
  assign \g134649/_0_  = ~n12286 ;
  assign \g134650/_0_  = ~n12319 ;
  assign \g134651/_0_  = ~n12340 ;
  assign \g134652/_0_  = ~n12359 ;
  assign \g134656/_0_  = ~n12383 ;
  assign \g134657/_0_  = ~n12404 ;
  assign \g134658/_0_  = ~n12436 ;
  assign \g134664/_0_  = ~n12469 ;
  assign \g134665/_0_  = ~n12497 ;
  assign \g134671/_0_  = ~n12538 ;
  assign \g134672/_0_  = ~n12563 ;
  assign \g134686/_0_  = ~n12599 ;
  assign \g134687/_0_  = ~n12629 ;
  assign \g134735/_0_  = ~n12966 ;
  assign \g134908/_0_  = ~n12999 ;
  assign \g134909/_0_  = ~n13017 ;
  assign \g134910/_0_  = ~n13054 ;
  assign \g134920/_0_  = ~n13075 ;
  assign \g134921/_0_  = ~n13111 ;
  assign \g134922/_0_  = ~n13139 ;
  assign \g134923/_0_  = ~n13173 ;
  assign \g134925/_0_  = ~n13208 ;
  assign \g134926/_0_  = ~n13229 ;
  assign \g134928/_0_  = ~n13247 ;
  assign \g134929/_0_  = ~n13270 ;
  assign \g134933/_0_  = ~n13290 ;
  assign \g134934/_0_  = ~n13324 ;
  assign \g134935/_0_  = ~n13358 ;
  assign \g134936/_0_  = ~n13393 ;
  assign \g134937/_0_  = ~n13411 ;
  assign \g134938/_0_  = ~n13428 ;
  assign \g134940/_0_  = ~n13462 ;
  assign \g134941/_0_  = ~n13491 ;
  assign \g134943/_0_  = ~n13528 ;
  assign \g134945/_0_  = ~n13548 ;
  assign \g134946/_0_  = ~n13570 ;
  assign \g134947/_0_  = ~n13600 ;
  assign \g134948/_0_  = ~n13635 ;
  assign \g134949/_0_  = ~n13672 ;
  assign \g134950/_0_  = ~n13693 ;
  assign \g134959/_0_  = ~n13731 ;
  assign \g134960/_0_  = ~n13762 ;
  assign \g134961/_0_  = ~n13807 ;
  assign \g134979/_0_  = ~n14055 ;
  assign \g134980/_0_  = ~n14078 ;
  assign \g135054/_0_  = ~n14093 ;
  assign \g135061/_0_  = ~n14116 ;
  assign \g135072/_0_  = ~n14129 ;
  assign \g135100/_0_  = ~n14141 ;
  assign \g135127/_0_  = ~n14160 ;
  assign \g135128/_0_  = ~n14179 ;
  assign \g135129/_0_  = ~n14198 ;
  assign \g135130/_0_  = ~n14217 ;
  assign \g135132/_0_  = ~n14236 ;
  assign \g135133/_0_  = ~n14255 ;
  assign \g135134/_0_  = ~n14274 ;
  assign \g135135/_0_  = ~n14293 ;
  assign \g135136/_0_  = ~n14312 ;
  assign \g135137/_0_  = ~n14331 ;
  assign \g135138/_0_  = ~n14350 ;
  assign \g135139/_0_  = ~n14369 ;
  assign \g135140/_0_  = ~n14388 ;
  assign \g135141/_0_  = ~n14407 ;
  assign \g135142/_0_  = ~n14426 ;
  assign \g135145/_0_  = ~n14446 ;
  assign \g135146/_0_  = ~n14467 ;
  assign \g135151/_0_  = ~n14499 ;
  assign \g135154/_0_  = ~n14520 ;
  assign \g135155/_0_  = ~n14541 ;
  assign \g135158/_0_  = ~n14562 ;
  assign \g135163/_0_  = ~n14597 ;
  assign \g135164/_0_  = ~n14634 ;
  assign \g135165/_0_  = ~n14655 ;
  assign \g135192/_0_  = ~n14670 ;
  assign \g135197/_0_  = ~n14706 ;
  assign \g135217/_0_  = ~n14723 ;
  assign \g135225/_0_  = ~n14740 ;
  assign \g135231/_0_  = ~n14785 ;
  assign \g135272/_0_  = ~n14823 ;
  assign \g135290/_0_  = ~n14934 ;
  assign \g135291/_0_  = ~n14951 ;
  assign \g135293/_0_  = ~n14995 ;
  assign \g135294/_0_  = ~n15017 ;
  assign \g135295/_0_  = ~n15056 ;
  assign \g135296/_0_  = ~n15071 ;
  assign \g135297/_0_  = ~n15404 ;
  assign \g135412/_0_  = ~n15432 ;
  assign \g135437/_0_  = ~n15447 ;
  assign \g135438/_0_  = ~n15459 ;
  assign \g135443/_0_  = ~n15478 ;
  assign \g135444/_0_  = ~n15497 ;
  assign \g135445/_0_  = ~n15516 ;
  assign \g135446/_0_  = ~n15535 ;
  assign \g135447/_0_  = ~n15554 ;
  assign \g135448/_0_  = ~n15573 ;
  assign \g135449/_0_  = ~n15592 ;
  assign \g135450/_0_  = ~n15611 ;
  assign \g135451/_0_  = ~n15630 ;
  assign \g135452/_0_  = ~n15649 ;
  assign \g135454/_0_  = ~n15668 ;
  assign \g135455/_0_  = ~n15687 ;
  assign \g135456/_0_  = ~n15706 ;
  assign \g135457/_0_  = ~n15725 ;
  assign \g135458/_0_  = ~n15744 ;
  assign \g135463/_0_  = ~n15768 ;
  assign \g135466/_0_  = ~n15784 ;
  assign \g135473/_0_  = ~n15813 ;
  assign \g135481/_0_  = ~n15834 ;
  assign \g135497/_0_  = ~n15844 ;
  assign \g135503/_0_  = ~n15853 ;
  assign \g135505/_0_  = ~n15862 ;
  assign \g135506/_0_  = ~n15871 ;
  assign \g135557/_0_  = ~n15881 ;
  assign \g135558/_0_  = ~n15891 ;
  assign \g135569/_0_  = ~n15941 ;
  assign \g135570/_0_  = ~n15986 ;
  assign \g135571/_0_  = ~n16031 ;
  assign \g135572/_0_  = ~n16049 ;
  assign \g135573/_0_  = ~n16060 ;
  assign \g135575/_0_  = ~n16085 ;
  assign \g135578/_0_  = ~n16126 ;
  assign \g135754/_0_  = ~n16149 ;
  assign \g135755/_0_  = ~n16167 ;
  assign \g135756/_0_  = ~n16186 ;
  assign \g135767/_0_  = ~n16207 ;
  assign \g135768/_0_  = ~n16229 ;
  assign \g135769/_0_  = ~n16251 ;
  assign \g135777/_0_  = ~n16270 ;
  assign \g135778/_0_  = ~n16288 ;
  assign \g135779/_0_  = ~n16310 ;
  assign \g135872/_0_  = ~n16330 ;
  assign \g135873/_0_  = ~n16347 ;
  assign \g135875/_0_  = ~n16395 ;
  assign \g135877/_0_  = ~n16416 ;
  assign \g135878/_0_  = ~n16428 ;
  assign \g135879/_0_  = ~n16440 ;
  assign \g135880/_0_  = ~n16487 ;
  assign \g136087/_0_  = ~n16509 ;
  assign \g136118/_0_  = ~n16601 ;
  assign \g136119/_0_  = ~n16619 ;
  assign \g136120/_0_  = ~n16637 ;
  assign \g136121/_0_  = ~n16655 ;
  assign \g136122/_0_  = ~n16673 ;
  assign \g136123/_0_  = ~n16691 ;
  assign \g136124/_0_  = ~n16709 ;
  assign \g136125/_0_  = ~n16727 ;
  assign \g136126/_0_  = ~n16745 ;
  assign \g136127/_0_  = ~n16763 ;
  assign \g136128/_0_  = ~n16781 ;
  assign \g136129/_0_  = ~n16799 ;
  assign \g136130/_0_  = ~n16817 ;
  assign \g136131/_0_  = ~n16835 ;
  assign \g136132/_0_  = ~n16853 ;
  assign \g136133/_0_  = ~n16871 ;
  assign \g136172/_0_  = ~n16887 ;
  assign \g136173/_0_  = ~n16902 ;
  assign \g136174/_0_  = ~n16910 ;
  assign \g136175/_0_  = ~n16918 ;
  assign \g136177/_0_  = ~n16939 ;
  assign \g136178/_0_  = ~n16948 ;
  assign \g136242/_0_  = ~n16961 ;
  assign \g136243/_0_  = ~n16966 ;
  assign \g136244/_0_  = ~n16980 ;
  assign \g136246/_0_  = ~n17023 ;
  assign \g136248/_0_  = ~n17035 ;
  assign \g136249/_0_  = ~n17077 ;
  assign \g136250/_0_  = ~n17122 ;
  assign \g136251/_0_  = ~n17165 ;
  assign \g136252/_0_  = ~n17206 ;
  assign \g136253/_0_  = ~n17248 ;
  assign \g136254/_0_  = ~n17259 ;
  assign \g136255/_0_  = ~n17273 ;
  assign \g136256/_0_  = ~n17284 ;
  assign \g136257/_0_  = ~n17294 ;
  assign \g136258/_0_  = ~n17304 ;
  assign \g136259/_0_  = ~n17315 ;
  assign \g136260/_0_  = ~n17325 ;
  assign \g136261/_0_  = ~n17335 ;
  assign \g136262/_0_  = ~n17345 ;
  assign \g136263/_0_  = ~n17355 ;
  assign \g136264/_0_  = ~n17396 ;
  assign \g136265/_0_  = ~n17437 ;
  assign \g136266/_0_  = ~n17449 ;
  assign \g136267/_0_  = ~n17460 ;
  assign \g136268/_0_  = ~n17503 ;
  assign \g136269/_0_  = ~n17547 ;
  assign \g136270/_0_  = ~n17590 ;
  assign \g136271/_0_  = ~n17634 ;
  assign \g136272/_0_  = ~n17645 ;
  assign \g136273/_0_  = ~n17687 ;
  assign \g136274/_0_  = ~n17731 ;
  assign \g136275/_0_  = ~n17776 ;
  assign \g136276/_0_  = ~n17790 ;
  assign \g136277/_0_  = ~n17801 ;
  assign \g136279/_0_  = ~n17812 ;
  assign \g136280/_0_  = ~n17823 ;
  assign \g136281/_0_  = ~n17866 ;
  assign \g136282/_0_  = ~n17877 ;
  assign \g136283/_0_  = ~n17888 ;
  assign \g136285/_0_  = ~n17930 ;
  assign \g136286/_0_  = ~n17976 ;
  assign \g136287/_0_  = ~n18021 ;
  assign \g136288/_0_  = ~n18033 ;
  assign \g136289/_0_  = ~n18043 ;
  assign \g136290/_0_  = ~n18087 ;
  assign \g136291/_0_  = ~n18129 ;
  assign \g136292/_0_  = ~n18176 ;
  assign \g136293/_0_  = ~n18183 ;
  assign \g136295/_0_  = ~n18197 ;
  assign \g136467/_0_  = ~n18232 ;
  assign \g136468/_0_  = ~n18259 ;
  assign \g136469/_0_  = ~n18280 ;
  assign \g136470/_0_  = ~n18301 ;
  assign \g136472/_0_  = ~n18321 ;
  assign \g136473/_0_  = ~n18339 ;
  assign \g136474/_0_  = ~n18358 ;
  assign \g136476/_0_  = ~n18378 ;
  assign \g136479/_0_  = ~n18399 ;
  assign \g136480/_0_  = ~n18418 ;
  assign \g136481/_0_  = ~n18438 ;
  assign \g136482/_0_  = ~n18459 ;
  assign \g136483/_0_  = ~n18479 ;
  assign \g136484/_0_  = ~n18498 ;
  assign \g136485/_0_  = ~n18516 ;
  assign \g136486/_0_  = ~n18536 ;
  assign \g136528/_0_  = ~n18605 ;
  assign \g136529/_0_  = ~n18641 ;
  assign \g136530/_0_  = ~n18678 ;
  assign \g136531/_0_  = ~n18720 ;
  assign \g136532/_0_  = ~n18755 ;
  assign \g136533/_0_  = ~n18795 ;
  assign \g136534/_0_  = ~n18829 ;
  assign \g136535/_0_  = ~n18865 ;
  assign \g136536/_0_  = ~n18903 ;
  assign \g136537/_0_  = ~n18939 ;
  assign \g136538/_0_  = ~n18979 ;
  assign \g136539/_0_  = ~n19016 ;
  assign \g136540/_0_  = ~n19054 ;
  assign \g136541/_0_  = ~n19086 ;
  assign \g136542/_0_  = ~n19124 ;
  assign \g136543/_0_  = ~n19158 ;
  assign \g136544/_0_  = ~n19193 ;
  assign \g136545/_0_  = ~n19232 ;
  assign \g136546/_0_  = ~n19267 ;
  assign \g136547/_0_  = ~n19303 ;
  assign \g136548/_0_  = ~n19342 ;
  assign \g136549/_0_  = ~n19378 ;
  assign \g136550/_0_  = ~n19420 ;
  assign \g136551/_0_  = ~n19454 ;
  assign \g136552/_0_  = ~n19487 ;
  assign \g136553/_0_  = ~n19522 ;
  assign \g136554/_0_  = ~n19561 ;
  assign \g136555/_0_  = ~n19594 ;
  assign \g136556/_0_  = ~n19630 ;
  assign \g136557/_0_  = ~n19663 ;
  assign \g136558/_0_  = ~n19699 ;
  assign \g136559/_0_  = ~n19732 ;
  assign \g136560/_0_  = ~n19765 ;
  assign \g136561/_0_  = ~n19796 ;
  assign \g136562/_0_  = ~n19828 ;
  assign \g136563/_0_  = ~n19863 ;
  assign \g136564/_0_  = ~n19894 ;
  assign \g136565/_0_  = ~n19926 ;
  assign \g136566/_0_  = ~n19963 ;
  assign \g136567/_0_  = ~n19996 ;
  assign \g136568/_0_  = ~n20031 ;
  assign \g136570/_0_  = ~n20067 ;
  assign \g136571/_0_  = ~n20100 ;
  assign \g136572/_0_  = ~n20135 ;
  assign \g136573/_0_  = ~n20164 ;
  assign \g136574/_0_  = ~n20198 ;
  assign \g136575/_0_  = ~n20232 ;
  assign \g136576/_0_  = ~n20263 ;
  assign \g136577/_0_  = ~n20296 ;
  assign \g136578/_0_  = ~n20329 ;
  assign \g136579/_0_  = ~n20364 ;
  assign \g136580/_0_  = ~n20398 ;
  assign \g136582/_0_  = ~n20453 ;
  assign \g136583/_0_  = ~n20489 ;
  assign \g136584/_0_  = ~n20525 ;
  assign \g136585/_0_  = ~n20561 ;
  assign \g136586/_0_  = ~n20597 ;
  assign \g136587/_0_  = ~n20634 ;
  assign \g136588/_0_  = ~n20669 ;
  assign \g136589/_0_  = ~n20714 ;
  assign \g136590/_0_  = ~n20751 ;
  assign \g136591/_0_  = ~n20790 ;
  assign \g136592/_0_  = ~n20824 ;
  assign \g136593/_0_  = ~n20865 ;
  assign \g136594/_0_  = ~n20900 ;
  assign \g136595/_0_  = ~n20937 ;
  assign \g136596/_0_  = ~n20972 ;
  assign \g136597/_0_  = ~n21012 ;
  assign \g136598/_0_  = ~n21053 ;
  assign \g136599/_0_  = ~n21088 ;
  assign \g136600/_0_  = ~n21126 ;
  assign \g136601/_0_  = ~n21164 ;
  assign \g136602/_0_  = ~n21205 ;
  assign \g136603/_0_  = ~n21243 ;
  assign \g136604/_0_  = ~n21278 ;
  assign \g136605/_0_  = ~n21313 ;
  assign \g136606/_0_  = ~n21347 ;
  assign \g136607/_0_  = ~n21380 ;
  assign \g136609/_0_  = ~n21412 ;
  assign \g136610/_0_  = ~n21446 ;
  assign \g136611/_0_  = ~n21480 ;
  assign \g136616/_0_  = ~n21514 ;
  assign \g136617/_0_  = ~n21548 ;
  assign \g136618/_0_  = ~n21582 ;
  assign \g136619/_0_  = ~n21616 ;
  assign \g136626/_0_  = ~n21629 ;
  assign \g136628/_0_  = ~n21643 ;
  assign \g136646/_0_  = ~n21657 ;
  assign \g136649/_0_  = ~n21670 ;
  assign \g136662/_0_  = ~n21682 ;
  assign \g136666/_0_  = ~n21694 ;
  assign \g136695/_0_  = ~n21710 ;
  assign \g136696/_0_  = ~n21721 ;
  assign \g136699/_0_  = ~n21734 ;
  assign \g136762/_0_  = ~n21751 ;
  assign \g136763/_0_  = ~n21762 ;
  assign \g136764/_0_  = ~n21768 ;
  assign \g136765/_0_  = ~n21786 ;
  assign \g136768/_0_  = ~n21810 ;
  assign \g136769/_0_  = ~n21820 ;
  assign \g137051/_0_  = ~n21831 ;
  assign \g137052/_0_  = ~n21841 ;
  assign \g137053/_0_  = ~n21852 ;
  assign \g137054/_0_  = ~n21862 ;
  assign \g137055/_0_  = ~n21875 ;
  assign \g137056/_0_  = ~n21885 ;
  assign \g137057/_0_  = ~n21898 ;
  assign \g137060/_0_  = ~n21908 ;
  assign \g137061/_0_  = ~n21918 ;
  assign \g137063/_0_  = ~n21928 ;
  assign \g137064/_0_  = ~n21938 ;
  assign \g137065/_0_  = ~n21951 ;
  assign \g137067/_0_  = ~n21961 ;
  assign \g137069/_0_  = ~n21974 ;
  assign \g137072/_0_  = ~n21984 ;
  assign \g137073/_0_  = ~n21999 ;
  assign \g137075/_0_  = ~n22006 ;
  assign \g137111/_0_  = ~n22012 ;
  assign \g137122/_0_  = ~n22020 ;
  assign \g137133/_0_  = ~n22033 ;
  assign \g137134/_0_  = ~n22067 ;
  assign \g137135/_0_  = ~n22095 ;
  assign \g137136/_0_  = ~n22128 ;
  assign \g137137/_0_  = ~n22160 ;
  assign \g137138/_0_  = ~n22193 ;
  assign \g137144/_0_  = ~n22210 ;
  assign \g137145/_0_  = ~n22245 ;
  assign \g137146/_0_  = ~n22278 ;
  assign \g137149/_0_  = ~n22300 ;
  assign \g137234/_0_  = ~n22312 ;
  assign \g137237/_0_  = ~n22325 ;
  assign \g137238/_0_  = ~n22339 ;
  assign \g137294/_0_  = ~n22357 ;
  assign \g137295/_0_  = ~n22367 ;
  assign \g137296/_0_  = ~n22377 ;
  assign \g137297/_0_  = ~n22389 ;
  assign \g137298/_0_  = ~n22410 ;
  assign \g137299/_0_  = ~n22421 ;
  assign \g137300/_0_  = ~n22431 ;
  assign \g137301/_0_  = ~n22441 ;
  assign \g137302/_0_  = ~n22447 ;
  assign \g137303/_0_  = ~n22457 ;
  assign \g137304/_0_  = ~n22468 ;
  assign \g137305/_0_  = ~n22479 ;
  assign \g137306/_0_  = ~n22489 ;
  assign \g137307/_0_  = ~n22500 ;
  assign \g137308/_0_  = ~n22512 ;
  assign \g137309/_0_  = ~n22523 ;
  assign \g137310/_0_  = ~n22534 ;
  assign \g137311/_0_  = ~n22544 ;
  assign \g137312/_0_  = ~n22550 ;
  assign \g137313/_0_  = ~n22555 ;
  assign \g137314/_0_  = ~n22577 ;
  assign \g137315/_0_  = ~n22584 ;
  assign \g137316/_0_  = ~n22635 ;
  assign \g137317/_0_  = ~n22681 ;
  assign \g137318/_0_  = ~n22732 ;
  assign \g137319/_0_  = ~n22778 ;
  assign \g137320/_0_  = ~n22827 ;
  assign \g137321/_0_  = ~n22873 ;
  assign \g137322/_0_  = ~n22922 ;
  assign \g137323/_0_  = ~n22943 ;
  assign \g137324/_0_  = ~n22966 ;
  assign \g137325/_0_  = ~n22983 ;
  assign \g137327/_0_  = ~n22986 ;
  assign \g137328/_0_  = ~n23033 ;
  assign \g137329/_0_  = ~n23085 ;
  assign \g137330/_0_  = ~n23135 ;
  assign \g137331/_0_  = ~n23184 ;
  assign \g137332/_0_  = ~n23233 ;
  assign \g137333/_0_  = ~n23281 ;
  assign \g137334/_0_  = ~n23328 ;
  assign \g137335/_0_  = ~n23346 ;
  assign \g137336/_0_  = ~n23363 ;
  assign \g137337/_0_  = ~n23382 ;
  assign \g137338/_0_  = ~n23391 ;
  assign \g137339/_0_  = ~n23401 ;
  assign \g137340/_0_  = ~n23413 ;
  assign \g137341/_0_  = ~n23416 ;
  assign \g137342/_0_  = ~n23419 ;
  assign \g137343/_0_  = ~n23422 ;
  assign \g137344/_0_  = ~n23426 ;
  assign \g137345/_0_  = ~n23473 ;
  assign \g137346/_0_  = ~n23520 ;
  assign \g137347/_0_  = ~n23523 ;
  assign \g137349/_0_  = ~n23571 ;
  assign \g137350/_0_  = ~n23617 ;
  assign \g137351/_0_  = ~n23665 ;
  assign \g137352/_0_  = ~n23713 ;
  assign \g137353/_0_  = ~n23760 ;
  assign \g137354/_0_  = ~n23763 ;
  assign \g137448/_0_  = ~n23771 ;
  assign \g137483/_0_  = ~n23784 ;
  assign \g137484/_0_  = ~n23797 ;
  assign \g137485/_0_  = ~n23810 ;
  assign \g137486/_0_  = ~n23823 ;
  assign \g137487/_0_  = ~n23838 ;
  assign \g137488/_0_  = ~n23853 ;
  assign \g137491/_0_  = ~n23866 ;
  assign \g137492/_0_  = ~n23879 ;
  assign \g137493/_0_  = ~n23892 ;
  assign \g137494/_0_  = ~n23905 ;
  assign \g137495/_0_  = ~n23918 ;
  assign \g137496/_0_  = ~n23931 ;
  assign \g137497/_0_  = ~n23944 ;
  assign \g137499/_0_  = ~n23957 ;
  assign \g137501/_0_  = ~n23970 ;
  assign \g137502/_0_  = ~n23983 ;
  assign \g137503/_0_  = ~n23996 ;
  assign \g137504/_0_  = ~n24009 ;
  assign \g137505/_0_  = ~n24022 ;
  assign \g137506/_0_  = ~n24035 ;
  assign \g137507/_0_  = ~n24048 ;
  assign \g137508/_0_  = ~n24061 ;
  assign \g137509/_0_  = ~n24074 ;
  assign \g137511/_0_  = ~n24087 ;
  assign \g137512/_0_  = ~n24100 ;
  assign \g137513/_0_  = ~n24113 ;
  assign \g137514/_0_  = ~n24126 ;
  assign \g137515/_0_  = ~n24139 ;
  assign \g137516/_0_  = ~n24152 ;
  assign \g137517/_0_  = ~n24165 ;
  assign \g137519/_0_  = ~n24184 ;
  assign \g137520/_0_  = ~n24203 ;
  assign \g137521/_0_  = ~n24211 ;
  assign \g137524/_0_  = ~n24218 ;
  assign \g137541/_0_  = ~n24228 ;
  assign \g137547/_0_  = ~n24234 ;
  assign \g137554/_0_  = ~n24244 ;
  assign \g137559/_0_  = ~n24255 ;
  assign \g137566/_0_  = ~n24266 ;
  assign \g137571/_0_  = ~n24275 ;
  assign \g137778/_0_  = ~n24288 ;
  assign \g137782/_0_  = ~n24299 ;
  assign \g137783/_0_  = ~n24310 ;
  assign \g137784/_0_  = ~n24322 ;
  assign \g137785/_0_  = ~n24333 ;
  assign \g137786/_0_  = ~n24343 ;
  assign \g137820/_0_  = ~n24352 ;
  assign \g137821/_0_  = ~n24362 ;
  assign \g137822/_0_  = ~n24372 ;
  assign \g137823/_0_  = ~n24378 ;
  assign \g137824/_0_  = ~n24386 ;
  assign \g137825/_0_  = ~n24396 ;
  assign \g137826/_0_  = ~n24406 ;
  assign \g137827/_0_  = ~n24416 ;
  assign \g137828/_0_  = ~n24426 ;
  assign \g137829/_0_  = ~n24436 ;
  assign \g137830/_0_  = ~n24446 ;
  assign \g137831/_0_  = ~n24456 ;
  assign \g137832/_0_  = ~n24466 ;
  assign \g137833/_0_  = ~n24476 ;
  assign \g137834/_0_  = ~n24486 ;
  assign \g137835/_0_  = ~n24494 ;
  assign \g137836/_0_  = ~n24505 ;
  assign \g137837/_0_  = ~n24516 ;
  assign \g137838/_0_  = ~n24527 ;
  assign \g137839/_0_  = ~n24537 ;
  assign \g137840/_0_  = ~n24547 ;
  assign \g137841/_0_  = ~n24558 ;
  assign \g137842/_0_  = ~n24568 ;
  assign \g137843/_0_  = ~n24578 ;
  assign \g137844/_0_  = ~n24588 ;
  assign \g137845/_0_  = ~n24598 ;
  assign \g137846/_0_  = ~n24608 ;
  assign \g137847/_0_  = ~n24618 ;
  assign \g137848/_0_  = ~n24628 ;
  assign \g137849/_0_  = ~n24638 ;
  assign \g137850/_0_  = ~n24646 ;
  assign \g137851/_0_  = ~n24656 ;
  assign \g137852/_0_  = ~n24666 ;
  assign \g137853/_0_  = ~n24676 ;
  assign \g137854/_0_  = ~n24687 ;
  assign \g137855/_0_  = ~n24696 ;
  assign \g137856/_0_  = ~n24706 ;
  assign \g137857/_0_  = ~n24716 ;
  assign \g137858/_0_  = ~n24726 ;
  assign \g137859/_0_  = ~n24736 ;
  assign \g137860/_0_  = ~n24746 ;
  assign \g137861/_0_  = ~n24754 ;
  assign \g137862/_0_  = ~n24764 ;
  assign \g137863/_0_  = ~n24776 ;
  assign \g137864/_0_  = ~n24787 ;
  assign \g137865/_0_  = ~n24797 ;
  assign \g137866/_0_  = ~n24807 ;
  assign \g137867/_0_  = ~n24815 ;
  assign \g137868/_0_  = ~n24825 ;
  assign \g137869/_0_  = ~n24835 ;
  assign \g137870/_0_  = ~n24845 ;
  assign \g137871/_0_  = ~n24855 ;
  assign \g137872/_0_  = ~n24866 ;
  assign \g137873/_0_  = ~n24876 ;
  assign \g137874/_0_  = ~n24886 ;
  assign \g137875/_0_  = ~n24898 ;
  assign \g137876/_0_  = ~n24909 ;
  assign \g137877/_0_  = ~n24919 ;
  assign \g137878/_0_  = ~n24929 ;
  assign \g137879/_0_  = ~n24937 ;
  assign \g137880/_0_  = ~n24948 ;
  assign \g137881/_0_  = ~n24959 ;
  assign \g137882/_0_  = ~n24970 ;
  assign \g137883/_0_  = ~n24980 ;
  assign \g137884/_0_  = ~n24991 ;
  assign \g137885/_0_  = ~n25001 ;
  assign \g137886/_0_  = ~n25011 ;
  assign \g137887/_0_  = ~n25021 ;
  assign \g137888/_0_  = ~n25031 ;
  assign \g137889/_0_  = ~n25041 ;
  assign \g137890/_0_  = ~n25051 ;
  assign \g137891/_0_  = ~n25061 ;
  assign \g137892/_0_  = ~n25071 ;
  assign \g137893/_0_  = ~n25082 ;
  assign \g137894/_0_  = ~n25092 ;
  assign \g137895/_0_  = ~n25102 ;
  assign \g137896/_0_  = ~n25112 ;
  assign \g137897/_0_  = ~n25122 ;
  assign \g137898/_0_  = ~n25132 ;
  assign \g137899/_0_  = ~n25142 ;
  assign \g137900/_0_  = ~n25152 ;
  assign \g137901/_0_  = ~n25162 ;
  assign \g137902/_0_  = ~n25172 ;
  assign \g137903/_0_  = ~n25177 ;
  assign \g138338/_0_  = ~n25181 ;
  assign \g138340/_0_  = ~n25184 ;
  assign \g138341/_0_  = ~n25197 ;
  assign \g138346/_0_  = ~n25209 ;
  assign \g138347/_0_  = ~n25222 ;
  assign \g138375/_0_  = ~n25228 ;
  assign \g138395/_0_  = ~n25240 ;
  assign \g138396/_0_  = ~n25252 ;
  assign \g138397/_0_  = ~n25260 ;
  assign \g138398/_0_  = ~n25268 ;
  assign \g138400/_0_  = ~n25275 ;
  assign \g138401/_0_  = ~n25287 ;
  assign \g138402/_0_  = ~n25299 ;
  assign \g138403/_0_  = ~n25308 ;
  assign \g138404/_0_  = ~n25321 ;
  assign \g138405/_0_  = ~n25328 ;
  assign \g138406/_0_  = ~n25336 ;
  assign \g138407/_0_  = ~n25344 ;
  assign \g138408/_0_  = ~n25356 ;
  assign \g138409/_0_  = ~n25366 ;
  assign \g138410/_0_  = ~n25374 ;
  assign \g138411/_0_  = ~n25382 ;
  assign \g138412/_0_  = ~n25390 ;
  assign \g138419/_0_  = ~n25403 ;
  assign \g138420/_0_  = ~n25411 ;
  assign \g138421/_0_  = ~n25422 ;
  assign \g138422/_0_  = ~n25429 ;
  assign \g138423/_0_  = ~n25441 ;
  assign \g138424/_0_  = ~n25453 ;
  assign \g138425/_0_  = ~n25466 ;
  assign \g138426/_0_  = ~n25478 ;
  assign \g138427/_0_  = ~n25487 ;
  assign \g138428/_0_  = ~n25497 ;
  assign \g138429/_0_  = ~n25507 ;
  assign \g138430/_0_  = ~n25517 ;
  assign \g138431/_0_  = ~n25527 ;
  assign \g138432/_0_  = ~n25532 ;
  assign \g138433/_0_  = ~n25537 ;
  assign \g138434/_0_  = ~n25543 ;
  assign \g138435/_0_  = ~n25548 ;
  assign \g138436/_0_  = ~n25554 ;
  assign \g138437/_0_  = ~n25560 ;
  assign \g138438/_0_  = ~n25565 ;
  assign \g138439/_0_  = ~n25570 ;
  assign \g138440/_0_  = ~n25575 ;
  assign \g138441/_0_  = ~n25580 ;
  assign \g138442/_0_  = ~n25588 ;
  assign \g138443/_0_  = ~n25593 ;
  assign \g138908/_0_  = ~n25601 ;
  assign \g138909/_0_  = ~n25609 ;
  assign \g138910/_0_  = ~n25617 ;
  assign \g138914/_0_  = ~n25625 ;
  assign \g138915/_0_  = ~n25633 ;
  assign \g138917/_0_  = ~n25641 ;
  assign \g138918/_0_  = ~n25649 ;
  assign \g138919/_0_  = ~n25657 ;
  assign \g138920/_0_  = ~n25665 ;
  assign \g138921/_0_  = ~n25673 ;
  assign \g138925/_0_  = ~n25681 ;
  assign \g138926/_0_  = ~n25689 ;
  assign \g138927/_0_  = ~n25697 ;
  assign \g138930/_0_  = ~n25705 ;
  assign \g138931/_0_  = ~n25713 ;
  assign \g138932/_0_  = ~n25721 ;
  assign \g138960/_0_  = ~n25729 ;
  assign \g138962/_0_  = ~n25737 ;
  assign \g139037/_0_  = ~n25748 ;
  assign \g139038/_0_  = ~n25756 ;
  assign \g139040/_0_  = ~n25764 ;
  assign \g139043/_0_  = ~n25769 ;
  assign \g139044/_0_  = ~n25777 ;
  assign \g139045/_0_  = ~n25782 ;
  assign \g139046/_0_  = ~n25790 ;
  assign \g139047/_0_  = ~n25798 ;
  assign \g139048/_0_  = ~n25806 ;
  assign \g139049/_0_  = ~n25814 ;
  assign \g139050/_0_  = ~n25822 ;
  assign \g139051/_0_  = ~n25830 ;
  assign \g139053/_0_  = ~n25836 ;
  assign \g139054/_0_  = ~n25844 ;
  assign \g139055/_0_  = ~n25852 ;
  assign \g139056/_0_  = ~n25860 ;
  assign \g139057/_0_  = ~n25868 ;
  assign \g139058/_0_  = ~n25876 ;
  assign \g139059/_0_  = ~n25884 ;
  assign \g139060/_0_  = ~n25895 ;
  assign \g139062/_0_  = ~n25903 ;
  assign \g139063/_0_  = ~n25911 ;
  assign \g139064/_0_  = ~n25922 ;
  assign \g139099/_0_  = ~n25930 ;
  assign \g139126/_0_  = ~n25940 ;
  assign \g139127/_0_  = ~n25946 ;
  assign \g139128/_0_  = ~n25956 ;
  assign \g139129/_0_  = ~n25961 ;
  assign \g139130/_0_  = ~n25971 ;
  assign \g139131/_0_  = ~n25976 ;
  assign \g139132/_0_  = ~n25986 ;
  assign \g139133/_0_  = ~n25996 ;
  assign \g139134/_0_  = ~n26006 ;
  assign \g139135/_0_  = ~n26016 ;
  assign \g139136/_0_  = ~n26026 ;
  assign \g139137/_0_  = ~n26036 ;
  assign \g139138/_0_  = ~n26046 ;
  assign \g139139/_0_  = ~n26056 ;
  assign \g139140/_0_  = ~n26066 ;
  assign \g139141/_0_  = ~n26076 ;
  assign \g139260/_0_  = ~n26089 ;
  assign \g139263/_0_  = ~n26102 ;
  assign \g139267/_0_  = ~n26117 ;
  assign \g139270/_0_  = ~n26130 ;
  assign \g139273/_0_  = ~n26143 ;
  assign \g139276/_0_  = ~n26156 ;
  assign \g139279/_0_  = ~n26169 ;
  assign \g139283/_0_  = ~n26182 ;
  assign \g139286/_0_  = ~n26195 ;
  assign \g139289/_0_  = ~n26208 ;
  assign \g139292/_0_  = ~n26221 ;
  assign \g139295/_0_  = ~n26234 ;
  assign \g139298/_0_  = ~n26247 ;
  assign \g139302/_0_  = ~n26260 ;
  assign \g139305/_0_  = ~n26273 ;
  assign \g139309/_0_  = ~n26292 ;
  assign \g139871/_0_  = ~n26300 ;
  assign \g139872/_0_  = ~n26308 ;
  assign \g139873/_0_  = ~n26316 ;
  assign \g139874/_0_  = ~n26324 ;
  assign \g139875/_0_  = ~n26332 ;
  assign \g139876/_0_  = ~n26340 ;
  assign \g139877/_0_  = ~n26348 ;
  assign \g139878/_0_  = ~n26356 ;
  assign \g139879/_0_  = ~n26364 ;
  assign \g139880/_0_  = ~n26372 ;
  assign \g139881/_0_  = ~n26380 ;
  assign \g139882/_0_  = ~n26388 ;
  assign \g139883/_0_  = ~n26396 ;
  assign \g139884/_0_  = ~n26404 ;
  assign \g139885/_0_  = ~n26412 ;
  assign \g139886/_0_  = ~n26420 ;
  assign \g139887/_0_  = ~n26428 ;
  assign \g139888/_0_  = ~n26436 ;
  assign \g139889/_0_  = ~n26444 ;
  assign \g139890/_0_  = ~n26452 ;
  assign \g139891/_0_  = ~n26460 ;
  assign \g139892/_0_  = ~n26468 ;
  assign \g139893/_0_  = ~n26476 ;
  assign \g139895/_0_  = ~n26484 ;
  assign \g139896/_0_  = ~n26492 ;
  assign \g139899/_0_  = ~n26500 ;
  assign \g139901/_0_  = ~n26508 ;
  assign \g139902/_0_  = ~n26516 ;
  assign \g139903/_0_  = ~n26524 ;
  assign \g139904/_0_  = ~n26532 ;
  assign \g140285/_0_  = ~n26573 ;
  assign \g140288/_0_  = ~n26613 ;
  assign \g140329/_0_  = ~n26652 ;
  assign \g140774/_0_  = ~n26669 ;
  assign \g140832/_0_  = ~n26686 ;
  assign \g140834/_0_  = ~n26699 ;
  assign \g140836/_0_  = ~n26712 ;
  assign \g140838/_0_  = ~n26727 ;
  assign \g140840/_0_  = ~n26740 ;
  assign \g140842/_0_  = ~n26753 ;
  assign \g140844/_0_  = ~n26766 ;
  assign \g140846/_0_  = ~n26779 ;
  assign \g140847/_0_  = ~n26792 ;
  assign \g140848/_0_  = ~n26805 ;
  assign \g140850/_0_  = ~n26818 ;
  assign \g140851/_0_  = ~n26831 ;
  assign \g140852/_0_  = ~n26844 ;
  assign \g140853/_0_  = ~n26857 ;
  assign \g140855/_0_  = ~n26870 ;
  assign \g140857/_0_  = ~n26883 ;
  assign \g140861/_0_  = ~n26902 ;
  assign \g140923/_0_  = ~n26919 ;
  assign \g141178/_0_  = ~n26934 ;
  assign \g141179/_0_  = ~n26945 ;
  assign \g141180/_0_  = ~n26956 ;
  assign \g141480/_0_  = ~n26971 ;
  assign \g141495/_0_  = ~n26986 ;
  assign \g141497/_0_  = ~n27001 ;
  assign \g141562/_0_  = ~n27011 ;
  assign \g141563/_0_  = ~n27017 ;
  assign \g141564/_0_  = ~n27027 ;
  assign \g141589/_0_  = ~n27034 ;
  assign \g141617/_0_  = ~n27042 ;
  assign \g141618/_0_  = ~n27055 ;
  assign \g141621/_0_  = ~n27068 ;
  assign \g141625/_0_  = ~n27083 ;
  assign \g141626/_0_  = ~n27098 ;
  assign \g141630/_0_  = ~n27111 ;
  assign \g141634/_0_  = ~n27124 ;
  assign \g141638/_0_  = ~n27137 ;
  assign \g141642/_0_  = ~n27150 ;
  assign \g141646/_0_  = ~n27163 ;
  assign \g141649/_0_  = ~n27176 ;
  assign \g141651/_0_  = ~n27189 ;
  assign \g141652/_0_  = ~n27202 ;
  assign \g141655/_0_  = ~n27215 ;
  assign \g141658/_0_  = ~n27228 ;
  assign \g141661/_0_  = ~n27241 ;
  assign \g141663/_0_  = ~n27254 ;
  assign \g141664/_0_  = ~n27267 ;
  assign \g141667/_0_  = ~n27280 ;
  assign \g141671/_0_  = ~n27299 ;
  assign \g141706/_0_  = ~n27305 ;
  assign \g141976/_0_  = ~n27316 ;
  assign \g141977/_0_  = ~n27326 ;
  assign \g141994/_0_  = ~n27336 ;
  assign \g142246/_0_  = ~n27349 ;
  assign \g142247/_0_  = ~n27362 ;
  assign \g142253/_0_  = ~n27373 ;
  assign \g142689/_0_  = ~n27386 ;
  assign \g142693/_0_  = ~n27399 ;
  assign \g142701/_0_  = ~n27412 ;
  assign \g142704/_0_  = ~n27425 ;
  assign \g142707/_0_  = ~n27438 ;
  assign \g142710/_0_  = ~n27451 ;
  assign \g142713/_0_  = ~n27464 ;
  assign \g142714/_0_  = ~n27477 ;
  assign \g142717/_0_  = ~n27490 ;
  assign \g142720/_0_  = ~n27503 ;
  assign \g142723/_0_  = ~n27516 ;
  assign \g142727/_0_  = ~n27529 ;
  assign \g142734/_0_  = ~n27548 ;
  assign \g143080/_0_  = ~n27559 ;
  assign \g143081/_0_  = ~n27571 ;
  assign \g143083/_0_  = ~n27587 ;
  assign \g143149/_0_  = ~n27597 ;
  assign \g143150/_0_  = ~n27607 ;
  assign \g143153/_0_  = ~n27620 ;
  assign \g143752/_0_  = ~n27634 ;
  assign \g143753/_0_  = ~n27650 ;
  assign \g143759/_0_  = ~n27664 ;
  assign \g144242/_0_  = ~n27676 ;
  assign \g144243/_0_  = ~n27685 ;
  assign \g144244/_0_  = ~n27696 ;
  assign \g144245/_0_  = ~n27708 ;
  assign \g144246/_0_  = ~n27717 ;
  assign \g144249/_0_  = ~n27726 ;
  assign \g145699/_0_  = ~n27736 ;
  assign \g145700/_0_  = ~n27746 ;
  assign \g145702/_0_  = ~n27758 ;
  assign \g145756/_0_  = ~n27767 ;
  assign \g145757/_0_  = ~n27777 ;
  assign \g145758/_0_  = ~n27787 ;
  assign \g146850/_0_  = ~n27796 ;
  assign \g146851/_0_  = ~n27805 ;
  assign \g146864/_0_  = ~n27814 ;
  assign \g147277/_0_  = ~n27824 ;
  assign \g147278/_0_  = ~n27833 ;
  assign \g147279/_0_  = ~n27843 ;
  assign \g147304/_0_  = ~n27853 ;
  assign \g147305/_0_  = ~n27863 ;
  assign \g147306/_0_  = ~n27872 ;
  assign \g147338/_3_  = ~n27894 ;
  assign \g147339/_3_  = ~n27900 ;
  assign \g147340/_3_  = ~n27906 ;
  assign \g147341/_3_  = ~n27912 ;
  assign \g147342/_3_  = ~n27918 ;
  assign \g147343/_3_  = ~n27924 ;
  assign \g147344/_3_  = ~n27930 ;
  assign \g147345/_3_  = ~n27936 ;
  assign \g147346/_3_  = ~n27942 ;
  assign \g147347/_3_  = ~n27948 ;
  assign \g147348/_3_  = ~n27954 ;
  assign \g147349/_3_  = ~n27960 ;
  assign \g147350/_3_  = ~n27966 ;
  assign \g147351/_3_  = ~n27972 ;
  assign \g147352/_3_  = ~n27978 ;
  assign \g147353/_3_  = ~n27984 ;
  assign \g147354/_3_  = ~n27990 ;
  assign \g147355/_3_  = ~n27996 ;
  assign \g147356/_3_  = ~n28002 ;
  assign \g147357/_3_  = ~n28008 ;
  assign \g147358/_3_  = ~n28014 ;
  assign \g147359/_3_  = ~n28020 ;
  assign \g147360/_3_  = ~n28026 ;
  assign \g147362/_3_  = ~n28032 ;
  assign \g147363/_3_  = ~n28038 ;
  assign \g147364/_3_  = ~n28044 ;
  assign \g147365/_3_  = ~n28050 ;
  assign \g147366/_3_  = ~n28056 ;
  assign \g147367/_3_  = ~n28062 ;
  assign \g147368/_3_  = ~n28068 ;
  assign \g147369/_3_  = ~n28074 ;
  assign \g148630/_0_  = ~n28083 ;
  assign \g148631/_0_  = ~n28094 ;
  assign \g148676/_0_  = ~n28103 ;
  assign \g148785/_0_  = ~n28112 ;
  assign \g148788/_0_  = ~n28122 ;
  assign \g148789/_0_  = ~n28131 ;
  assign \g148834/_0_  = ~n28140 ;
  assign \g148836/_0_  = ~n28150 ;
  assign \g148838/_0_  = ~n28161 ;
  assign \g149836/_0_  = ~n28170 ;
  assign \g149837/_0_  = ~n28180 ;
  assign \g149838/_0_  = ~n28190 ;
  assign \g150142/_0_  = ~n28191 ;
  assign \g152366/_0_  = ~n28200 ;
  assign \g152367/_0_  = ~n28209 ;
  assign \g152368/_0_  = ~n28218 ;
  assign \g152426/_0_  = ~n28229 ;
  assign \g152427/_0_  = ~n28239 ;
  assign \g152428/_0_  = ~n28248 ;
  assign \g152586/_0_  = ~n28259 ;
  assign \g152587/_0_  = ~n28269 ;
  assign \g152588/_0_  = ~n28278 ;
  assign \g153217/_0_  = ~n27880 ;
  assign \g154117/_0_  = ~n28287 ;
  assign \g154118/_0_  = ~n28296 ;
  assign \g154130/_0_  = ~n28306 ;
  assign \g154269/_0_  = ~n28317 ;
  assign \g154270/_0_  = ~n28328 ;
  assign \g154284/_0_  = ~n28339 ;
  assign \g154682/_0_  = ~n28350 ;
  assign \g155004/_0_  = ~n28361 ;
  assign \g155020/_0_  = ~n28371 ;
  assign \g155121/_0_  = n28381 ;
  assign \g155124/_0_  = ~n28393 ;
  assign \g155126/_0_  = n28403 ;
  assign \g155228/_0_  = ~n28412 ;
  assign \g155229/_0_  = ~n28421 ;
  assign \g155230/_0_  = ~n28430 ;
  assign \g155326/_0_  = ~n28440 ;
  assign \g155327/_0_  = ~n28450 ;
  assign \g155330/_0_  = ~n28460 ;
  assign \g155353/_0_  = ~n28469 ;
  assign \g155354/_0_  = ~n28478 ;
  assign \g155356/_0_  = ~n28487 ;
  assign \g155602/_0_  = ~n28502 ;
  assign \g155633/_0_  = ~n28515 ;
  assign \g155634/_0_  = ~n28530 ;
  assign \g155699/_0_  = ~n28539 ;
  assign \g155708/_0_  = ~n28547 ;
  assign \g155715/_0_  = ~n28556 ;
  assign \g156008/_0_  = ~n28561 ;
  assign \g156013/_0_  = ~n28566 ;
  assign \g156019/_0_  = ~n28571 ;
  assign \g156352/_0_  = ~n28580 ;
  assign \g156353/_0_  = ~n28589 ;
  assign \g156356/_0_  = ~n28598 ;
  assign \g156359/_0_  = ~n28607 ;
  assign \g156360/_0_  = ~n28617 ;
  assign \g156361/_0_  = ~n28627 ;
  assign \g156464/_0_  = ~n28636 ;
  assign \g156465/_0_  = ~n28646 ;
  assign \g156469/_0_  = ~n28655 ;
  assign \g156777/_0_  = ~n28659 ;
  assign \g156778/_0_  = ~n28663 ;
  assign \g156789/_0_  = ~n28667 ;
  assign \g158956/_0_  = ~n28676 ;
  assign \g158957/_0_  = ~n28686 ;
  assign \g158966/_0_  = ~n28696 ;
  assign \g159429/_1_  = ~n28550 ;
  assign \g159477/_1_  = ~n28533 ;
  assign \g159500/_1_  = ~n28540 ;
  assign \g159681/_0_  = ~n28705 ;
  assign \g159890/_0_  = n28710 ;
  assign \g159950/_0_  = n28715 ;
  assign \g160246/_0_  = n28720 ;
  assign \g160846/_0_  = ~n28723 ;
  assign \g160860/_0_  = ~n28726 ;
  assign \g160961/_0_  = ~n28728 ;
  assign \g160987/_0_  = ~n28730 ;
  assign \g161000/_0_  = ~n28733 ;
  assign \g161005/_0_  = ~n28736 ;
  assign \g161042/_0_  = ~n28738 ;
  assign \g161119/_0_  = ~n28741 ;
  assign \g161143/_0_  = ~n28744 ;
  assign \g161150/_0_  = ~n28747 ;
  assign \g161172/_0_  = ~n28750 ;
  assign \g161207/_0_  = ~n28752 ;
  assign \g161315/_0_  = ~n28754 ;
  assign \g161332/_0_  = ~n28757 ;
  assign \g161421/_0_  = ~n28760 ;
  assign \g161492/_0_  = ~n28762 ;
  assign \g161541/_0_  = ~n28765 ;
  assign \g161623/_0_  = ~n28768 ;
  assign \g161655/_0_  = ~n28771 ;
  assign \g161678/_0_  = ~n28774 ;
  assign \g161709/_0_  = ~n28777 ;
  assign \g161737/_0_  = ~n28780 ;
  assign \g161751/_0_  = ~n28783 ;
  assign \g161756/_0_  = ~n28786 ;
  assign \g162016/_0_  = n28791 ;
  assign \g162020/_0_  = n28796 ;
  assign \g162024/_0_  = n28801 ;
  assign \g163326/_0_  = ~n28697 ;
  assign \g163326/_3_  = n28697 ;
  assign \g174072/_1_  = ~n26585 ;
  assign \g174360/_1_  = ~n26543 ;
  assign \g174391/_0_  = ~n26615 ;
  assign \g180307/_0_  = ~n28817 ;
  assign \g180335/_0_  = ~n28837 ;
  assign \g180369/_0_  = ~n28853 ;
  assign \g180385/_0_  = ~n28869 ;
  assign \g180395/_0_  = ~n28885 ;
  assign \g180442/_0_  = ~n28901 ;
  assign \g180453/_0_  = ~n28917 ;
  assign \g180524/_0_  = ~n28935 ;
  assign \g180586/_0_  = ~n28966 ;
  assign \g180596/_0_  = ~n28983 ;
  assign \g180606/_0_  = ~n28999 ;
  assign \g180654/_0_  = ~n29015 ;
  assign \g180715/_0_  = ~n29060 ;
  assign \g180805/_0_  = ~n29076 ;
  assign \g180836/_0_  = ~n29107 ;
  assign \g180929/_0_  = ~n29133 ;
  assign \g180944/_0_  = ~n29142 ;
  assign \g180975/_0_  = ~n29158 ;
  assign \g181036/_0_  = ~n29174 ;
  assign \g181072/_0_  = ~n29192 ;
  assign \g181083/_0_  = ~n29215 ;
  assign \g181093/_0_  = ~n29233 ;
  assign \g181127/_0_  = ~n29249 ;
  assign \g181137/_0_  = ~n29267 ;
  assign \g181150/_0_  = ~n29283 ;
  assign \g181160/_0_  = ~n29299 ;
  assign \g181180/_0_  = ~n29315 ;
  assign \g181191/_0_  = ~n29331 ;
  assign \g181238/_0_  = ~n29347 ;
  assign \g181262/_0_  = ~n29360 ;
  assign \g181270/_0_  = ~n29376 ;
  assign \g181280/_0_  = ~n29392 ;
  assign \g181315/_0_  = ~n29410 ;
  assign \g181366/_0_  = ~n29422 ;
  assign \g181385/_0_  = ~n29447 ;
  assign \g181458/_0_  = ~n29461 ;
  assign \g181464/_0_  = ~n29480 ;
  assign \g181478/_0_  = ~n29498 ;
  assign \g181522/_0_  = ~n29514 ;
  assign \g181537/_0_  = ~n29532 ;
  assign \g181584/_0_  = ~n29552 ;
  assign \g181669/_0_  = ~n29573 ;
  assign \g181681/_0_  = ~n29589 ;
  assign \g181719/_0_  = ~n29599 ;
  assign \g181778/_0_  = ~n29615 ;
  assign \g181840/_0_  = ~n29631 ;
  assign \g181936/_0_  = ~n29648 ;
  assign \g181986/_0_  = ~n29665 ;
  assign \g182000/_0_  = ~n29683 ;
  assign \g182083/_0_  = ~n29693 ;
  assign \g182179/_0_  = ~n29709 ;
  assign \g182201/_0_  = ~n29725 ;
  assign \g182227/_0_  = ~n29732 ;
  assign \g182316/_0_  = ~n29742 ;
  assign \g182358/_0_  = ~n29758 ;
  assign \g182473/_0_  = ~n29777 ;
  assign \g182678/_0_  = ~n29790 ;
  assign \g53/_0_  = ~n29806 ;
endmodule
