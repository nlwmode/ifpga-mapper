module top (\a0_pad , a_pad, \b0_pad , \c0_pad , c_pad, \d0_pad , d_pad, \e0_pad , e_pad, \f0_pad , f_pad, \g0_pad , g_pad, \h0_pad , h_pad, \i0_pad , i_pad, \j0_pad , j_pad, \k0_pad , k_pad, \l0_pad , l_pad, \m0_pad , m_pad, \n0_pad , n_pad, \o0_pad , o_pad, \p0_pad , p_pad, \q0_pad , q_pad, \r0_pad , r_pad, \s0_pad , s_pad, \t0_pad , t_pad, \u0_pad , u_pad, \v0_pad , v_pad, w_pad, x_pad, y_pad, z_pad, \a1_pad , \a2_pad , \b1_pad , \b2_pad , \c1_pad , \c2_pad , \d1_pad , \d2_pad , \e1_pad , \e2_pad , \f1_pad , \f2_pad , \g1_pad , \h1_pad , \i1_pad , \j1_pad , \k1_pad , \l1_pad , \m1_pad , \n1_pad , \o1_pad , \p1_pad , \q1_pad , \r1_pad , \s1_pad , \t1_pad , \u1_pad , \v1_pad , \w0_pad , \w1_pad , \x0_pad , \x1_pad , \y0_pad , \y1_pad , \z0_pad , \z1_pad );
	input \a0_pad  ;
	input a_pad ;
	input \b0_pad  ;
	input \c0_pad  ;
	input c_pad ;
	input \d0_pad  ;
	input d_pad ;
	input \e0_pad  ;
	input e_pad ;
	input \f0_pad  ;
	input f_pad ;
	input \g0_pad  ;
	input g_pad ;
	input \h0_pad  ;
	input h_pad ;
	input \i0_pad  ;
	input i_pad ;
	input \j0_pad  ;
	input j_pad ;
	input \k0_pad  ;
	input k_pad ;
	input \l0_pad  ;
	input l_pad ;
	input \m0_pad  ;
	input m_pad ;
	input \n0_pad  ;
	input n_pad ;
	input \o0_pad  ;
	input o_pad ;
	input \p0_pad  ;
	input p_pad ;
	input \q0_pad  ;
	input q_pad ;
	input \r0_pad  ;
	input r_pad ;
	input \s0_pad  ;
	input s_pad ;
	input \t0_pad  ;
	input t_pad ;
	input \u0_pad  ;
	input u_pad ;
	input \v0_pad  ;
	input v_pad ;
	input w_pad ;
	input x_pad ;
	input y_pad ;
	input z_pad ;
	output \a1_pad  ;
	output \a2_pad  ;
	output \b1_pad  ;
	output \b2_pad  ;
	output \c1_pad  ;
	output \c2_pad  ;
	output \d1_pad  ;
	output \d2_pad  ;
	output \e1_pad  ;
	output \e2_pad  ;
	output \f1_pad  ;
	output \f2_pad  ;
	output \g1_pad  ;
	output \h1_pad  ;
	output \i1_pad  ;
	output \j1_pad  ;
	output \k1_pad  ;
	output \l1_pad  ;
	output \m1_pad  ;
	output \n1_pad  ;
	output \o1_pad  ;
	output \p1_pad  ;
	output \q1_pad  ;
	output \r1_pad  ;
	output \s1_pad  ;
	output \t1_pad  ;
	output \u1_pad  ;
	output \v1_pad  ;
	output \w0_pad  ;
	output \w1_pad  ;
	output \x0_pad  ;
	output \x1_pad  ;
	output \y0_pad  ;
	output \y1_pad  ;
	output \z0_pad  ;
	output \z1_pad  ;
	wire _w102_ ;
	wire _w101_ ;
	wire _w100_ ;
	wire _w99_ ;
	wire _w98_ ;
	wire _w97_ ;
	wire _w96_ ;
	wire _w95_ ;
	wire _w94_ ;
	wire _w93_ ;
	wire _w92_ ;
	wire _w91_ ;
	wire _w90_ ;
	wire _w89_ ;
	wire _w88_ ;
	wire _w87_ ;
	wire _w86_ ;
	wire _w85_ ;
	wire _w84_ ;
	wire _w83_ ;
	wire _w82_ ;
	wire _w81_ ;
	wire _w80_ ;
	wire _w79_ ;
	wire _w78_ ;
	wire _w61_ ;
	wire _w60_ ;
	wire _w59_ ;
	wire _w58_ ;
	wire _w57_ ;
	wire _w56_ ;
	wire _w55_ ;
	wire _w54_ ;
	wire _w53_ ;
	wire _w52_ ;
	wire _w51_ ;
	wire _w50_ ;
	wire _w49_ ;
	wire _w62_ ;
	wire _w63_ ;
	wire _w64_ ;
	wire _w65_ ;
	wire _w66_ ;
	wire _w67_ ;
	wire _w68_ ;
	wire _w69_ ;
	wire _w70_ ;
	wire _w71_ ;
	wire _w72_ ;
	wire _w73_ ;
	wire _w74_ ;
	wire _w75_ ;
	wire _w76_ ;
	wire _w77_ ;
	LUT4 #(
		.INIT('h0b08)
	) name0 (
		d_pad,
		i_pad,
		l_pad,
		q_pad,
		_w49_
	);
	LUT3 #(
		.INIT('h02)
	) name1 (
		k_pad,
		p_pad,
		\r0_pad ,
		_w50_
	);
	LUT4 #(
		.INIT('h3302)
	) name2 (
		k_pad,
		l_pad,
		p_pad,
		\q0_pad ,
		_w51_
	);
	LUT2 #(
		.INIT('h4)
	) name3 (
		_w50_,
		_w51_,
		_w52_
	);
	LUT4 #(
		.INIT('h0b08)
	) name4 (
		e_pad,
		i_pad,
		l_pad,
		r_pad,
		_w53_
	);
	LUT3 #(
		.INIT('h02)
	) name5 (
		k_pad,
		p_pad,
		\s0_pad ,
		_w54_
	);
	LUT4 #(
		.INIT('h3302)
	) name6 (
		k_pad,
		l_pad,
		p_pad,
		\r0_pad ,
		_w55_
	);
	LUT2 #(
		.INIT('h4)
	) name7 (
		_w54_,
		_w55_,
		_w56_
	);
	LUT4 #(
		.INIT('h3210)
	) name8 (
		j_pad,
		l_pad,
		s_pad,
		t_pad,
		_w57_
	);
	LUT3 #(
		.INIT('h02)
	) name9 (
		k_pad,
		p_pad,
		\t0_pad ,
		_w58_
	);
	LUT4 #(
		.INIT('h3302)
	) name10 (
		k_pad,
		l_pad,
		p_pad,
		\s0_pad ,
		_w59_
	);
	LUT2 #(
		.INIT('h4)
	) name11 (
		_w58_,
		_w59_,
		_w60_
	);
	LUT4 #(
		.INIT('h3210)
	) name12 (
		j_pad,
		l_pad,
		t_pad,
		u_pad,
		_w61_
	);
	LUT3 #(
		.INIT('h02)
	) name13 (
		k_pad,
		p_pad,
		\u0_pad ,
		_w62_
	);
	LUT4 #(
		.INIT('h3302)
	) name14 (
		k_pad,
		l_pad,
		p_pad,
		\t0_pad ,
		_w63_
	);
	LUT2 #(
		.INIT('h4)
	) name15 (
		_w62_,
		_w63_,
		_w64_
	);
	LUT4 #(
		.INIT('h3210)
	) name16 (
		j_pad,
		l_pad,
		u_pad,
		v_pad,
		_w65_
	);
	LUT3 #(
		.INIT('h02)
	) name17 (
		k_pad,
		p_pad,
		\v0_pad ,
		_w66_
	);
	LUT4 #(
		.INIT('h3302)
	) name18 (
		k_pad,
		l_pad,
		p_pad,
		\u0_pad ,
		_w67_
	);
	LUT2 #(
		.INIT('h4)
	) name19 (
		_w66_,
		_w67_,
		_w68_
	);
	LUT4 #(
		.INIT('h3210)
	) name20 (
		j_pad,
		l_pad,
		v_pad,
		w_pad,
		_w69_
	);
	LUT3 #(
		.INIT('h04)
	) name21 (
		a_pad,
		k_pad,
		p_pad,
		_w70_
	);
	LUT4 #(
		.INIT('h3302)
	) name22 (
		k_pad,
		l_pad,
		p_pad,
		\v0_pad ,
		_w71_
	);
	LUT2 #(
		.INIT('h4)
	) name23 (
		_w70_,
		_w71_,
		_w72_
	);
	LUT4 #(
		.INIT('h3210)
	) name24 (
		j_pad,
		l_pad,
		w_pad,
		x_pad,
		_w73_
	);
	LUT4 #(
		.INIT('h3210)
	) name25 (
		j_pad,
		l_pad,
		x_pad,
		y_pad,
		_w74_
	);
	LUT4 #(
		.INIT('h3210)
	) name26 (
		j_pad,
		l_pad,
		y_pad,
		z_pad,
		_w75_
	);
	LUT4 #(
		.INIT('h0b08)
	) name27 (
		\a0_pad ,
		j_pad,
		l_pad,
		z_pad,
		_w76_
	);
	LUT4 #(
		.INIT('h00ca)
	) name28 (
		\a0_pad ,
		\b0_pad ,
		j_pad,
		l_pad,
		_w77_
	);
	LUT4 #(
		.INIT('h00ca)
	) name29 (
		\b0_pad ,
		\c0_pad ,
		j_pad,
		l_pad,
		_w78_
	);
	LUT4 #(
		.INIT('h00ca)
	) name30 (
		\c0_pad ,
		\d0_pad ,
		j_pad,
		l_pad,
		_w79_
	);
	LUT4 #(
		.INIT('h00ca)
	) name31 (
		\d0_pad ,
		\e0_pad ,
		j_pad,
		l_pad,
		_w80_
	);
	LUT4 #(
		.INIT('h00ca)
	) name32 (
		\e0_pad ,
		\f0_pad ,
		j_pad,
		l_pad,
		_w81_
	);
	LUT4 #(
		.INIT('h00ac)
	) name33 (
		a_pad,
		\f0_pad ,
		j_pad,
		l_pad,
		_w82_
	);
	LUT4 #(
		.INIT('h00ca)
	) name34 (
		\g0_pad ,
		\h0_pad ,
		k_pad,
		l_pad,
		_w83_
	);
	LUT4 #(
		.INIT('h00ca)
	) name35 (
		\h0_pad ,
		\i0_pad ,
		k_pad,
		l_pad,
		_w84_
	);
	LUT4 #(
		.INIT('h00ca)
	) name36 (
		\i0_pad ,
		\j0_pad ,
		k_pad,
		l_pad,
		_w85_
	);
	LUT4 #(
		.INIT('h00ca)
	) name37 (
		\j0_pad ,
		\k0_pad ,
		k_pad,
		l_pad,
		_w86_
	);
	LUT4 #(
		.INIT('h00e2)
	) name38 (
		\k0_pad ,
		k_pad,
		\l0_pad ,
		l_pad,
		_w87_
	);
	LUT4 #(
		.INIT('h0e04)
	) name39 (
		k_pad,
		\l0_pad ,
		l_pad,
		\m0_pad ,
		_w88_
	);
	LUT4 #(
		.INIT('h0b08)
	) name40 (
		f_pad,
		i_pad,
		l_pad,
		m_pad,
		_w89_
	);
	LUT4 #(
		.INIT('h3210)
	) name41 (
		k_pad,
		l_pad,
		\m0_pad ,
		\n0_pad ,
		_w90_
	);
	LUT4 #(
		.INIT('h0b08)
	) name42 (
		g_pad,
		i_pad,
		l_pad,
		n_pad,
		_w91_
	);
	LUT4 #(
		.INIT('h440c)
	) name43 (
		a_pad,
		k_pad,
		\o0_pad ,
		p_pad,
		_w92_
	);
	LUT3 #(
		.INIT('h32)
	) name44 (
		k_pad,
		l_pad,
		\n0_pad ,
		_w93_
	);
	LUT2 #(
		.INIT('h4)
	) name45 (
		_w92_,
		_w93_,
		_w94_
	);
	LUT4 #(
		.INIT('h0b08)
	) name46 (
		h_pad,
		i_pad,
		l_pad,
		o_pad,
		_w95_
	);
	LUT3 #(
		.INIT('h02)
	) name47 (
		k_pad,
		\p0_pad ,
		p_pad,
		_w96_
	);
	LUT4 #(
		.INIT('h3032)
	) name48 (
		k_pad,
		l_pad,
		\o0_pad ,
		p_pad,
		_w97_
	);
	LUT2 #(
		.INIT('h4)
	) name49 (
		_w96_,
		_w97_,
		_w98_
	);
	LUT4 #(
		.INIT('h0b08)
	) name50 (
		c_pad,
		i_pad,
		l_pad,
		p_pad,
		_w99_
	);
	LUT3 #(
		.INIT('h02)
	) name51 (
		k_pad,
		p_pad,
		\q0_pad ,
		_w100_
	);
	LUT4 #(
		.INIT('h3032)
	) name52 (
		k_pad,
		l_pad,
		\p0_pad ,
		p_pad,
		_w101_
	);
	LUT2 #(
		.INIT('h4)
	) name53 (
		_w100_,
		_w101_,
		_w102_
	);
	assign \a1_pad  = _w49_ ;
	assign \a2_pad  = _w52_ ;
	assign \b1_pad  = _w53_ ;
	assign \b2_pad  = _w56_ ;
	assign \c1_pad  = _w57_ ;
	assign \c2_pad  = _w60_ ;
	assign \d1_pad  = _w61_ ;
	assign \d2_pad  = _w64_ ;
	assign \e1_pad  = _w65_ ;
	assign \e2_pad  = _w68_ ;
	assign \f1_pad  = _w69_ ;
	assign \f2_pad  = _w72_ ;
	assign \g1_pad  = _w73_ ;
	assign \h1_pad  = _w74_ ;
	assign \i1_pad  = _w75_ ;
	assign \j1_pad  = _w76_ ;
	assign \k1_pad  = _w77_ ;
	assign \l1_pad  = _w78_ ;
	assign \m1_pad  = _w79_ ;
	assign \n1_pad  = _w80_ ;
	assign \o1_pad  = _w81_ ;
	assign \p1_pad  = _w82_ ;
	assign \q1_pad  = _w83_ ;
	assign \r1_pad  = _w84_ ;
	assign \s1_pad  = _w85_ ;
	assign \t1_pad  = _w86_ ;
	assign \u1_pad  = _w87_ ;
	assign \v1_pad  = _w88_ ;
	assign \w0_pad  = _w89_ ;
	assign \w1_pad  = _w90_ ;
	assign \x0_pad  = _w91_ ;
	assign \x1_pad  = _w94_ ;
	assign \y0_pad  = _w95_ ;
	assign \y1_pad  = _w98_ ;
	assign \z0_pad  = _w99_ ;
	assign \z1_pad  = _w102_ ;
endmodule;