module top (\a0_pad , a_pad, \b0_pad , b_pad, \c0_pad , c_pad, \d0_pad , d_pad, \e0_pad , e_pad, \f0_pad , f_pad, \g0_pad , g_pad, h_pad, i_pad, j_pad, k_pad, l_pad, m_pad, n_pad, o_pad, p_pad, q_pad, r_pad, s_pad, t_pad, u_pad, v_pad, w_pad, x_pad, y_pad, z_pad, \h0_pad , \i0_pad , \j0_pad , \k0_pad , \l0_pad , \m0_pad , \n0_pad , \o0_pad , \p0_pad , \q0_pad , \r0_pad , \s0_pad , \t0_pad , \u0_pad , \v0_pad , \w0_pad , \x0_pad );
	input \a0_pad  ;
	input a_pad ;
	input \b0_pad  ;
	input b_pad ;
	input \c0_pad  ;
	input c_pad ;
	input \d0_pad  ;
	input d_pad ;
	input \e0_pad  ;
	input e_pad ;
	input \f0_pad  ;
	input f_pad ;
	input \g0_pad  ;
	input g_pad ;
	input h_pad ;
	input i_pad ;
	input j_pad ;
	input k_pad ;
	input l_pad ;
	input m_pad ;
	input n_pad ;
	input o_pad ;
	input p_pad ;
	input q_pad ;
	input r_pad ;
	input s_pad ;
	input t_pad ;
	input u_pad ;
	input v_pad ;
	input w_pad ;
	input x_pad ;
	input y_pad ;
	input z_pad ;
	output \h0_pad  ;
	output \i0_pad  ;
	output \j0_pad  ;
	output \k0_pad  ;
	output \l0_pad  ;
	output \m0_pad  ;
	output \n0_pad  ;
	output \o0_pad  ;
	output \p0_pad  ;
	output \q0_pad  ;
	output \r0_pad  ;
	output \s0_pad  ;
	output \t0_pad  ;
	output \u0_pad  ;
	output \v0_pad  ;
	output \w0_pad  ;
	output \x0_pad  ;
	wire _w161_ ;
	wire _w92_ ;
	wire _w91_ ;
	wire _w90_ ;
	wire _w89_ ;
	wire _w88_ ;
	wire _w87_ ;
	wire _w86_ ;
	wire _w85_ ;
	wire _w84_ ;
	wire _w83_ ;
	wire _w82_ ;
	wire _w81_ ;
	wire _w80_ ;
	wire _w79_ ;
	wire _w78_ ;
	wire _w77_ ;
	wire _w76_ ;
	wire _w75_ ;
	wire _w74_ ;
	wire _w73_ ;
	wire _w72_ ;
	wire _w71_ ;
	wire _w70_ ;
	wire _w69_ ;
	wire _w68_ ;
	wire _w67_ ;
	wire _w66_ ;
	wire _w65_ ;
	wire _w64_ ;
	wire _w63_ ;
	wire _w46_ ;
	wire _w45_ ;
	wire _w44_ ;
	wire _w43_ ;
	wire _w42_ ;
	wire _w41_ ;
	wire _w40_ ;
	wire _w39_ ;
	wire _w38_ ;
	wire _w37_ ;
	wire _w36_ ;
	wire _w35_ ;
	wire _w34_ ;
	wire _w47_ ;
	wire _w48_ ;
	wire _w49_ ;
	wire _w50_ ;
	wire _w51_ ;
	wire _w52_ ;
	wire _w53_ ;
	wire _w54_ ;
	wire _w55_ ;
	wire _w56_ ;
	wire _w57_ ;
	wire _w58_ ;
	wire _w59_ ;
	wire _w60_ ;
	wire _w61_ ;
	wire _w62_ ;
	wire _w93_ ;
	wire _w94_ ;
	wire _w95_ ;
	wire _w96_ ;
	wire _w97_ ;
	wire _w98_ ;
	wire _w99_ ;
	wire _w100_ ;
	wire _w101_ ;
	wire _w102_ ;
	wire _w103_ ;
	wire _w104_ ;
	wire _w105_ ;
	wire _w106_ ;
	wire _w107_ ;
	wire _w108_ ;
	wire _w109_ ;
	wire _w110_ ;
	wire _w111_ ;
	wire _w112_ ;
	wire _w113_ ;
	wire _w114_ ;
	wire _w115_ ;
	wire _w116_ ;
	wire _w117_ ;
	wire _w118_ ;
	wire _w119_ ;
	wire _w120_ ;
	wire _w121_ ;
	wire _w122_ ;
	wire _w123_ ;
	wire _w124_ ;
	wire _w125_ ;
	wire _w126_ ;
	wire _w127_ ;
	wire _w128_ ;
	wire _w129_ ;
	wire _w130_ ;
	wire _w131_ ;
	wire _w132_ ;
	wire _w133_ ;
	wire _w134_ ;
	wire _w135_ ;
	wire _w136_ ;
	wire _w137_ ;
	wire _w138_ ;
	wire _w139_ ;
	wire _w140_ ;
	wire _w141_ ;
	wire _w142_ ;
	wire _w143_ ;
	wire _w144_ ;
	wire _w145_ ;
	wire _w146_ ;
	wire _w147_ ;
	wire _w148_ ;
	wire _w149_ ;
	wire _w150_ ;
	wire _w151_ ;
	wire _w152_ ;
	wire _w153_ ;
	wire _w154_ ;
	wire _w155_ ;
	wire _w156_ ;
	wire _w157_ ;
	wire _w158_ ;
	wire _w159_ ;
	wire _w160_ ;
	LUT2 #(
		.INIT('h1)
	) name0 (
		a_pad,
		q_pad,
		_w34_
	);
	LUT2 #(
		.INIT('h8)
	) name1 (
		a_pad,
		q_pad,
		_w35_
	);
	LUT2 #(
		.INIT('h1)
	) name2 (
		_w34_,
		_w35_,
		_w36_
	);
	LUT2 #(
		.INIT('h8)
	) name3 (
		b_pad,
		r_pad,
		_w37_
	);
	LUT2 #(
		.INIT('h1)
	) name4 (
		b_pad,
		r_pad,
		_w38_
	);
	LUT2 #(
		.INIT('h8)
	) name5 (
		c_pad,
		s_pad,
		_w39_
	);
	LUT2 #(
		.INIT('h1)
	) name6 (
		c_pad,
		s_pad,
		_w40_
	);
	LUT2 #(
		.INIT('h8)
	) name7 (
		d_pad,
		t_pad,
		_w41_
	);
	LUT2 #(
		.INIT('h1)
	) name8 (
		d_pad,
		t_pad,
		_w42_
	);
	LUT2 #(
		.INIT('h8)
	) name9 (
		e_pad,
		u_pad,
		_w43_
	);
	LUT2 #(
		.INIT('h1)
	) name10 (
		e_pad,
		u_pad,
		_w44_
	);
	LUT2 #(
		.INIT('h8)
	) name11 (
		f_pad,
		v_pad,
		_w45_
	);
	LUT2 #(
		.INIT('h1)
	) name12 (
		f_pad,
		v_pad,
		_w46_
	);
	LUT2 #(
		.INIT('h8)
	) name13 (
		g_pad,
		w_pad,
		_w47_
	);
	LUT2 #(
		.INIT('h1)
	) name14 (
		g_pad,
		w_pad,
		_w48_
	);
	LUT2 #(
		.INIT('h8)
	) name15 (
		h_pad,
		x_pad,
		_w49_
	);
	LUT2 #(
		.INIT('h1)
	) name16 (
		h_pad,
		x_pad,
		_w50_
	);
	LUT2 #(
		.INIT('h8)
	) name17 (
		i_pad,
		y_pad,
		_w51_
	);
	LUT2 #(
		.INIT('h1)
	) name18 (
		i_pad,
		y_pad,
		_w52_
	);
	LUT2 #(
		.INIT('h8)
	) name19 (
		j_pad,
		z_pad,
		_w53_
	);
	LUT2 #(
		.INIT('h1)
	) name20 (
		j_pad,
		z_pad,
		_w54_
	);
	LUT2 #(
		.INIT('h8)
	) name21 (
		\a0_pad ,
		k_pad,
		_w55_
	);
	LUT2 #(
		.INIT('h1)
	) name22 (
		\a0_pad ,
		k_pad,
		_w56_
	);
	LUT2 #(
		.INIT('h8)
	) name23 (
		\b0_pad ,
		l_pad,
		_w57_
	);
	LUT2 #(
		.INIT('h1)
	) name24 (
		\b0_pad ,
		l_pad,
		_w58_
	);
	LUT2 #(
		.INIT('h8)
	) name25 (
		\c0_pad ,
		m_pad,
		_w59_
	);
	LUT2 #(
		.INIT('h1)
	) name26 (
		\c0_pad ,
		m_pad,
		_w60_
	);
	LUT2 #(
		.INIT('h8)
	) name27 (
		\d0_pad ,
		n_pad,
		_w61_
	);
	LUT2 #(
		.INIT('h1)
	) name28 (
		\d0_pad ,
		n_pad,
		_w62_
	);
	LUT2 #(
		.INIT('h8)
	) name29 (
		\e0_pad ,
		o_pad,
		_w63_
	);
	LUT2 #(
		.INIT('h1)
	) name30 (
		\e0_pad ,
		o_pad,
		_w64_
	);
	LUT2 #(
		.INIT('h8)
	) name31 (
		\f0_pad ,
		p_pad,
		_w65_
	);
	LUT2 #(
		.INIT('h1)
	) name32 (
		\f0_pad ,
		p_pad,
		_w66_
	);
	LUT2 #(
		.INIT('h2)
	) name33 (
		\g0_pad ,
		_w66_,
		_w67_
	);
	LUT2 #(
		.INIT('h1)
	) name34 (
		_w65_,
		_w67_,
		_w68_
	);
	LUT2 #(
		.INIT('h1)
	) name35 (
		_w64_,
		_w68_,
		_w69_
	);
	LUT2 #(
		.INIT('h1)
	) name36 (
		_w63_,
		_w69_,
		_w70_
	);
	LUT2 #(
		.INIT('h1)
	) name37 (
		_w62_,
		_w70_,
		_w71_
	);
	LUT2 #(
		.INIT('h1)
	) name38 (
		_w61_,
		_w71_,
		_w72_
	);
	LUT2 #(
		.INIT('h1)
	) name39 (
		_w60_,
		_w72_,
		_w73_
	);
	LUT2 #(
		.INIT('h1)
	) name40 (
		_w59_,
		_w73_,
		_w74_
	);
	LUT2 #(
		.INIT('h1)
	) name41 (
		_w58_,
		_w74_,
		_w75_
	);
	LUT2 #(
		.INIT('h1)
	) name42 (
		_w57_,
		_w75_,
		_w76_
	);
	LUT2 #(
		.INIT('h1)
	) name43 (
		_w56_,
		_w76_,
		_w77_
	);
	LUT2 #(
		.INIT('h1)
	) name44 (
		_w55_,
		_w77_,
		_w78_
	);
	LUT2 #(
		.INIT('h1)
	) name45 (
		_w54_,
		_w78_,
		_w79_
	);
	LUT2 #(
		.INIT('h1)
	) name46 (
		_w53_,
		_w79_,
		_w80_
	);
	LUT2 #(
		.INIT('h1)
	) name47 (
		_w52_,
		_w80_,
		_w81_
	);
	LUT2 #(
		.INIT('h1)
	) name48 (
		_w51_,
		_w81_,
		_w82_
	);
	LUT2 #(
		.INIT('h1)
	) name49 (
		_w50_,
		_w82_,
		_w83_
	);
	LUT2 #(
		.INIT('h1)
	) name50 (
		_w49_,
		_w83_,
		_w84_
	);
	LUT2 #(
		.INIT('h1)
	) name51 (
		_w48_,
		_w84_,
		_w85_
	);
	LUT2 #(
		.INIT('h1)
	) name52 (
		_w47_,
		_w85_,
		_w86_
	);
	LUT2 #(
		.INIT('h1)
	) name53 (
		_w46_,
		_w86_,
		_w87_
	);
	LUT2 #(
		.INIT('h1)
	) name54 (
		_w45_,
		_w87_,
		_w88_
	);
	LUT2 #(
		.INIT('h1)
	) name55 (
		_w44_,
		_w88_,
		_w89_
	);
	LUT2 #(
		.INIT('h1)
	) name56 (
		_w43_,
		_w89_,
		_w90_
	);
	LUT2 #(
		.INIT('h1)
	) name57 (
		_w42_,
		_w90_,
		_w91_
	);
	LUT2 #(
		.INIT('h1)
	) name58 (
		_w41_,
		_w91_,
		_w92_
	);
	LUT2 #(
		.INIT('h1)
	) name59 (
		_w40_,
		_w92_,
		_w93_
	);
	LUT2 #(
		.INIT('h1)
	) name60 (
		_w39_,
		_w93_,
		_w94_
	);
	LUT2 #(
		.INIT('h1)
	) name61 (
		_w38_,
		_w94_,
		_w95_
	);
	LUT2 #(
		.INIT('h1)
	) name62 (
		_w37_,
		_w95_,
		_w96_
	);
	LUT2 #(
		.INIT('h2)
	) name63 (
		_w36_,
		_w96_,
		_w97_
	);
	LUT2 #(
		.INIT('h4)
	) name64 (
		_w36_,
		_w96_,
		_w98_
	);
	LUT2 #(
		.INIT('h1)
	) name65 (
		_w97_,
		_w98_,
		_w99_
	);
	LUT2 #(
		.INIT('h1)
	) name66 (
		_w37_,
		_w38_,
		_w100_
	);
	LUT2 #(
		.INIT('h4)
	) name67 (
		_w94_,
		_w100_,
		_w101_
	);
	LUT2 #(
		.INIT('h2)
	) name68 (
		_w94_,
		_w100_,
		_w102_
	);
	LUT2 #(
		.INIT('h1)
	) name69 (
		_w101_,
		_w102_,
		_w103_
	);
	LUT2 #(
		.INIT('h1)
	) name70 (
		_w39_,
		_w40_,
		_w104_
	);
	LUT2 #(
		.INIT('h4)
	) name71 (
		_w92_,
		_w104_,
		_w105_
	);
	LUT2 #(
		.INIT('h2)
	) name72 (
		_w92_,
		_w104_,
		_w106_
	);
	LUT2 #(
		.INIT('h1)
	) name73 (
		_w105_,
		_w106_,
		_w107_
	);
	LUT2 #(
		.INIT('h1)
	) name74 (
		_w41_,
		_w42_,
		_w108_
	);
	LUT2 #(
		.INIT('h4)
	) name75 (
		_w90_,
		_w108_,
		_w109_
	);
	LUT2 #(
		.INIT('h2)
	) name76 (
		_w90_,
		_w108_,
		_w110_
	);
	LUT2 #(
		.INIT('h1)
	) name77 (
		_w109_,
		_w110_,
		_w111_
	);
	LUT2 #(
		.INIT('h1)
	) name78 (
		_w43_,
		_w44_,
		_w112_
	);
	LUT2 #(
		.INIT('h4)
	) name79 (
		_w88_,
		_w112_,
		_w113_
	);
	LUT2 #(
		.INIT('h2)
	) name80 (
		_w88_,
		_w112_,
		_w114_
	);
	LUT2 #(
		.INIT('h1)
	) name81 (
		_w113_,
		_w114_,
		_w115_
	);
	LUT2 #(
		.INIT('h1)
	) name82 (
		_w45_,
		_w46_,
		_w116_
	);
	LUT2 #(
		.INIT('h4)
	) name83 (
		_w86_,
		_w116_,
		_w117_
	);
	LUT2 #(
		.INIT('h2)
	) name84 (
		_w86_,
		_w116_,
		_w118_
	);
	LUT2 #(
		.INIT('h1)
	) name85 (
		_w117_,
		_w118_,
		_w119_
	);
	LUT2 #(
		.INIT('h1)
	) name86 (
		_w47_,
		_w48_,
		_w120_
	);
	LUT2 #(
		.INIT('h4)
	) name87 (
		_w84_,
		_w120_,
		_w121_
	);
	LUT2 #(
		.INIT('h2)
	) name88 (
		_w84_,
		_w120_,
		_w122_
	);
	LUT2 #(
		.INIT('h1)
	) name89 (
		_w121_,
		_w122_,
		_w123_
	);
	LUT2 #(
		.INIT('h1)
	) name90 (
		_w49_,
		_w50_,
		_w124_
	);
	LUT2 #(
		.INIT('h4)
	) name91 (
		_w82_,
		_w124_,
		_w125_
	);
	LUT2 #(
		.INIT('h2)
	) name92 (
		_w82_,
		_w124_,
		_w126_
	);
	LUT2 #(
		.INIT('h1)
	) name93 (
		_w125_,
		_w126_,
		_w127_
	);
	LUT2 #(
		.INIT('h1)
	) name94 (
		_w51_,
		_w52_,
		_w128_
	);
	LUT2 #(
		.INIT('h4)
	) name95 (
		_w80_,
		_w128_,
		_w129_
	);
	LUT2 #(
		.INIT('h2)
	) name96 (
		_w80_,
		_w128_,
		_w130_
	);
	LUT2 #(
		.INIT('h1)
	) name97 (
		_w129_,
		_w130_,
		_w131_
	);
	LUT2 #(
		.INIT('h1)
	) name98 (
		_w53_,
		_w54_,
		_w132_
	);
	LUT2 #(
		.INIT('h4)
	) name99 (
		_w78_,
		_w132_,
		_w133_
	);
	LUT2 #(
		.INIT('h2)
	) name100 (
		_w78_,
		_w132_,
		_w134_
	);
	LUT2 #(
		.INIT('h1)
	) name101 (
		_w133_,
		_w134_,
		_w135_
	);
	LUT2 #(
		.INIT('h1)
	) name102 (
		_w55_,
		_w56_,
		_w136_
	);
	LUT2 #(
		.INIT('h4)
	) name103 (
		_w76_,
		_w136_,
		_w137_
	);
	LUT2 #(
		.INIT('h2)
	) name104 (
		_w76_,
		_w136_,
		_w138_
	);
	LUT2 #(
		.INIT('h1)
	) name105 (
		_w137_,
		_w138_,
		_w139_
	);
	LUT2 #(
		.INIT('h1)
	) name106 (
		_w57_,
		_w58_,
		_w140_
	);
	LUT2 #(
		.INIT('h4)
	) name107 (
		_w74_,
		_w140_,
		_w141_
	);
	LUT2 #(
		.INIT('h2)
	) name108 (
		_w74_,
		_w140_,
		_w142_
	);
	LUT2 #(
		.INIT('h1)
	) name109 (
		_w141_,
		_w142_,
		_w143_
	);
	LUT2 #(
		.INIT('h1)
	) name110 (
		_w59_,
		_w60_,
		_w144_
	);
	LUT2 #(
		.INIT('h4)
	) name111 (
		_w72_,
		_w144_,
		_w145_
	);
	LUT2 #(
		.INIT('h2)
	) name112 (
		_w72_,
		_w144_,
		_w146_
	);
	LUT2 #(
		.INIT('h1)
	) name113 (
		_w145_,
		_w146_,
		_w147_
	);
	LUT2 #(
		.INIT('h1)
	) name114 (
		_w61_,
		_w62_,
		_w148_
	);
	LUT2 #(
		.INIT('h4)
	) name115 (
		_w70_,
		_w148_,
		_w149_
	);
	LUT2 #(
		.INIT('h2)
	) name116 (
		_w70_,
		_w148_,
		_w150_
	);
	LUT2 #(
		.INIT('h1)
	) name117 (
		_w149_,
		_w150_,
		_w151_
	);
	LUT2 #(
		.INIT('h1)
	) name118 (
		_w63_,
		_w64_,
		_w152_
	);
	LUT2 #(
		.INIT('h4)
	) name119 (
		_w68_,
		_w152_,
		_w153_
	);
	LUT2 #(
		.INIT('h2)
	) name120 (
		_w68_,
		_w152_,
		_w154_
	);
	LUT2 #(
		.INIT('h1)
	) name121 (
		_w153_,
		_w154_,
		_w155_
	);
	LUT2 #(
		.INIT('h1)
	) name122 (
		_w65_,
		_w66_,
		_w156_
	);
	LUT2 #(
		.INIT('h1)
	) name123 (
		\g0_pad ,
		_w156_,
		_w157_
	);
	LUT2 #(
		.INIT('h8)
	) name124 (
		\g0_pad ,
		_w156_,
		_w158_
	);
	LUT2 #(
		.INIT('h1)
	) name125 (
		_w157_,
		_w158_,
		_w159_
	);
	LUT2 #(
		.INIT('h1)
	) name126 (
		_w34_,
		_w96_,
		_w160_
	);
	LUT2 #(
		.INIT('h1)
	) name127 (
		_w35_,
		_w160_,
		_w161_
	);
	assign \h0_pad  = _w99_ ;
	assign \i0_pad  = _w103_ ;
	assign \j0_pad  = _w107_ ;
	assign \k0_pad  = _w111_ ;
	assign \l0_pad  = _w115_ ;
	assign \m0_pad  = _w119_ ;
	assign \n0_pad  = _w123_ ;
	assign \o0_pad  = _w127_ ;
	assign \p0_pad  = _w131_ ;
	assign \q0_pad  = _w135_ ;
	assign \r0_pad  = _w139_ ;
	assign \s0_pad  = _w143_ ;
	assign \t0_pad  = _w147_ ;
	assign \u0_pad  = _w151_ ;
	assign \v0_pad  = _w155_ ;
	assign \w0_pad  = _w159_ ;
	assign \x0_pad  = _w161_ ;
endmodule;