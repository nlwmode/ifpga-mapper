module top (CLR_pad, \v0_pad , \v10_reg/NET0131 , \v11_reg/NET0131 , \v12_reg/NET0131 , \v1_pad , \v2_pad , \v3_pad , \v4_pad , \v5_pad , \v6_pad , \v7_reg/NET0131 , \v8_reg/NET0131 , \v9_reg/NET0131 , \_al_n0 , \_al_n1 , \g1759/_1_ , \g1762/_1_ , \g1764/_1_ , \g1765/_0_ , \g1786/_2_ , \g1791/_3_ , \g1808/_3_ , \g1822/_2_ , \g1929/_3_ , \g2713/_1_ , \g2744/_0_ , \v13_D_11_pad , \v13_D_12_pad , \v13_D_13_pad , \v13_D_14_pad , \v13_D_16_pad , \v13_D_18_pad , \v13_D_19_pad , \v13_D_21_pad , \v13_D_22_pad , \v13_D_23_pad , \v13_D_24_pad , \v13_D_7_pad , \v13_D_8_pad , \v13_D_9_pad );
	input CLR_pad ;
	input \v0_pad  ;
	input \v10_reg/NET0131  ;
	input \v11_reg/NET0131  ;
	input \v12_reg/NET0131  ;
	input \v1_pad  ;
	input \v2_pad  ;
	input \v3_pad  ;
	input \v4_pad  ;
	input \v5_pad  ;
	input \v6_pad  ;
	input \v7_reg/NET0131  ;
	input \v8_reg/NET0131  ;
	input \v9_reg/NET0131  ;
	output \_al_n0  ;
	output \_al_n1  ;
	output \g1759/_1_  ;
	output \g1762/_1_  ;
	output \g1764/_1_  ;
	output \g1765/_0_  ;
	output \g1786/_2_  ;
	output \g1791/_3_  ;
	output \g1808/_3_  ;
	output \g1822/_2_  ;
	output \g1929/_3_  ;
	output \g2713/_1_  ;
	output \g2744/_0_  ;
	output \v13_D_11_pad  ;
	output \v13_D_12_pad  ;
	output \v13_D_13_pad  ;
	output \v13_D_14_pad  ;
	output \v13_D_16_pad  ;
	output \v13_D_18_pad  ;
	output \v13_D_19_pad  ;
	output \v13_D_21_pad  ;
	output \v13_D_22_pad  ;
	output \v13_D_23_pad  ;
	output \v13_D_24_pad  ;
	output \v13_D_7_pad  ;
	output \v13_D_8_pad  ;
	output \v13_D_9_pad  ;
	wire _w580_ ;
	wire _w579_ ;
	wire _w578_ ;
	wire _w577_ ;
	wire _w576_ ;
	wire _w575_ ;
	wire _w574_ ;
	wire _w573_ ;
	wire _w572_ ;
	wire _w571_ ;
	wire _w570_ ;
	wire _w569_ ;
	wire _w568_ ;
	wire _w567_ ;
	wire _w566_ ;
	wire _w565_ ;
	wire _w564_ ;
	wire _w563_ ;
	wire _w562_ ;
	wire _w561_ ;
	wire _w560_ ;
	wire _w559_ ;
	wire _w558_ ;
	wire _w557_ ;
	wire _w556_ ;
	wire _w271_ ;
	wire _w270_ ;
	wire _w269_ ;
	wire _w268_ ;
	wire _w267_ ;
	wire _w266_ ;
	wire _w265_ ;
	wire _w264_ ;
	wire _w263_ ;
	wire _w262_ ;
	wire _w261_ ;
	wire _w260_ ;
	wire _w259_ ;
	wire _w258_ ;
	wire _w257_ ;
	wire _w256_ ;
	wire _w255_ ;
	wire _w254_ ;
	wire _w253_ ;
	wire _w252_ ;
	wire _w251_ ;
	wire _w250_ ;
	wire _w249_ ;
	wire _w248_ ;
	wire _w247_ ;
	wire _w246_ ;
	wire _w245_ ;
	wire _w244_ ;
	wire _w243_ ;
	wire _w242_ ;
	wire _w241_ ;
	wire _w240_ ;
	wire _w239_ ;
	wire _w238_ ;
	wire _w237_ ;
	wire _w236_ ;
	wire _w235_ ;
	wire _w234_ ;
	wire _w233_ ;
	wire _w232_ ;
	wire _w231_ ;
	wire _w230_ ;
	wire _w229_ ;
	wire _w228_ ;
	wire _w227_ ;
	wire _w226_ ;
	wire _w225_ ;
	wire _w224_ ;
	wire _w223_ ;
	wire _w222_ ;
	wire _w221_ ;
	wire _w220_ ;
	wire _w219_ ;
	wire _w218_ ;
	wire _w217_ ;
	wire _w216_ ;
	wire _w215_ ;
	wire _w214_ ;
	wire _w213_ ;
	wire _w212_ ;
	wire _w211_ ;
	wire _w210_ ;
	wire _w209_ ;
	wire _w208_ ;
	wire _w207_ ;
	wire _w206_ ;
	wire _w205_ ;
	wire _w204_ ;
	wire _w203_ ;
	wire _w202_ ;
	wire _w201_ ;
	wire _w200_ ;
	wire _w199_ ;
	wire _w198_ ;
	wire _w197_ ;
	wire _w196_ ;
	wire _w195_ ;
	wire _w194_ ;
	wire _w193_ ;
	wire _w192_ ;
	wire _w191_ ;
	wire _w190_ ;
	wire _w189_ ;
	wire _w188_ ;
	wire _w187_ ;
	wire _w186_ ;
	wire _w185_ ;
	wire _w184_ ;
	wire _w183_ ;
	wire _w182_ ;
	wire _w181_ ;
	wire _w180_ ;
	wire _w179_ ;
	wire _w178_ ;
	wire _w177_ ;
	wire _w176_ ;
	wire _w175_ ;
	wire _w174_ ;
	wire _w173_ ;
	wire _w172_ ;
	wire _w171_ ;
	wire _w170_ ;
	wire _w169_ ;
	wire _w168_ ;
	wire _w167_ ;
	wire _w166_ ;
	wire _w165_ ;
	wire _w164_ ;
	wire _w163_ ;
	wire _w162_ ;
	wire _w161_ ;
	wire _w160_ ;
	wire _w159_ ;
	wire _w158_ ;
	wire _w157_ ;
	wire _w156_ ;
	wire _w155_ ;
	wire _w154_ ;
	wire _w153_ ;
	wire _w152_ ;
	wire _w151_ ;
	wire _w150_ ;
	wire _w149_ ;
	wire _w148_ ;
	wire _w147_ ;
	wire _w146_ ;
	wire _w145_ ;
	wire _w144_ ;
	wire _w143_ ;
	wire _w142_ ;
	wire _w73_ ;
	wire _w72_ ;
	wire _w71_ ;
	wire _w70_ ;
	wire _w69_ ;
	wire _w68_ ;
	wire _w67_ ;
	wire _w66_ ;
	wire _w65_ ;
	wire _w64_ ;
	wire _w63_ ;
	wire _w62_ ;
	wire _w61_ ;
	wire _w60_ ;
	wire _w59_ ;
	wire _w58_ ;
	wire _w57_ ;
	wire _w56_ ;
	wire _w55_ ;
	wire _w54_ ;
	wire _w53_ ;
	wire _w52_ ;
	wire _w51_ ;
	wire _w50_ ;
	wire _w49_ ;
	wire _w48_ ;
	wire _w47_ ;
	wire _w46_ ;
	wire _w45_ ;
	wire _w44_ ;
	wire _w27_ ;
	wire _w26_ ;
	wire _w25_ ;
	wire _w24_ ;
	wire _w23_ ;
	wire _w22_ ;
	wire _w21_ ;
	wire _w20_ ;
	wire _w19_ ;
	wire _w18_ ;
	wire _w17_ ;
	wire _w16_ ;
	wire _w15_ ;
	wire _w28_ ;
	wire _w29_ ;
	wire _w30_ ;
	wire _w31_ ;
	wire _w32_ ;
	wire _w33_ ;
	wire _w34_ ;
	wire _w35_ ;
	wire _w36_ ;
	wire _w37_ ;
	wire _w38_ ;
	wire _w39_ ;
	wire _w40_ ;
	wire _w41_ ;
	wire _w42_ ;
	wire _w43_ ;
	wire _w74_ ;
	wire _w75_ ;
	wire _w76_ ;
	wire _w77_ ;
	wire _w78_ ;
	wire _w79_ ;
	wire _w80_ ;
	wire _w81_ ;
	wire _w82_ ;
	wire _w83_ ;
	wire _w84_ ;
	wire _w85_ ;
	wire _w86_ ;
	wire _w87_ ;
	wire _w88_ ;
	wire _w89_ ;
	wire _w90_ ;
	wire _w91_ ;
	wire _w92_ ;
	wire _w93_ ;
	wire _w94_ ;
	wire _w95_ ;
	wire _w96_ ;
	wire _w97_ ;
	wire _w98_ ;
	wire _w99_ ;
	wire _w100_ ;
	wire _w101_ ;
	wire _w102_ ;
	wire _w103_ ;
	wire _w104_ ;
	wire _w105_ ;
	wire _w106_ ;
	wire _w107_ ;
	wire _w108_ ;
	wire _w109_ ;
	wire _w110_ ;
	wire _w111_ ;
	wire _w112_ ;
	wire _w113_ ;
	wire _w114_ ;
	wire _w115_ ;
	wire _w116_ ;
	wire _w117_ ;
	wire _w118_ ;
	wire _w119_ ;
	wire _w120_ ;
	wire _w121_ ;
	wire _w122_ ;
	wire _w123_ ;
	wire _w124_ ;
	wire _w125_ ;
	wire _w126_ ;
	wire _w127_ ;
	wire _w128_ ;
	wire _w129_ ;
	wire _w130_ ;
	wire _w131_ ;
	wire _w132_ ;
	wire _w133_ ;
	wire _w134_ ;
	wire _w135_ ;
	wire _w136_ ;
	wire _w137_ ;
	wire _w138_ ;
	wire _w139_ ;
	wire _w140_ ;
	wire _w141_ ;
	wire _w272_ ;
	wire _w273_ ;
	wire _w274_ ;
	wire _w275_ ;
	wire _w276_ ;
	wire _w277_ ;
	wire _w278_ ;
	wire _w279_ ;
	wire _w280_ ;
	wire _w281_ ;
	wire _w282_ ;
	wire _w283_ ;
	wire _w284_ ;
	wire _w285_ ;
	wire _w286_ ;
	wire _w287_ ;
	wire _w288_ ;
	wire _w289_ ;
	wire _w290_ ;
	wire _w291_ ;
	wire _w292_ ;
	wire _w293_ ;
	wire _w294_ ;
	wire _w295_ ;
	wire _w296_ ;
	wire _w297_ ;
	wire _w298_ ;
	wire _w299_ ;
	wire _w300_ ;
	wire _w301_ ;
	wire _w302_ ;
	wire _w303_ ;
	wire _w304_ ;
	wire _w305_ ;
	wire _w306_ ;
	wire _w307_ ;
	wire _w308_ ;
	wire _w309_ ;
	wire _w310_ ;
	wire _w311_ ;
	wire _w312_ ;
	wire _w313_ ;
	wire _w314_ ;
	wire _w315_ ;
	wire _w316_ ;
	wire _w317_ ;
	wire _w318_ ;
	wire _w319_ ;
	wire _w320_ ;
	wire _w321_ ;
	wire _w322_ ;
	wire _w323_ ;
	wire _w324_ ;
	wire _w325_ ;
	wire _w326_ ;
	wire _w327_ ;
	wire _w328_ ;
	wire _w329_ ;
	wire _w330_ ;
	wire _w331_ ;
	wire _w332_ ;
	wire _w333_ ;
	wire _w334_ ;
	wire _w335_ ;
	wire _w336_ ;
	wire _w337_ ;
	wire _w338_ ;
	wire _w339_ ;
	wire _w340_ ;
	wire _w341_ ;
	wire _w342_ ;
	wire _w343_ ;
	wire _w344_ ;
	wire _w345_ ;
	wire _w346_ ;
	wire _w347_ ;
	wire _w348_ ;
	wire _w349_ ;
	wire _w350_ ;
	wire _w351_ ;
	wire _w352_ ;
	wire _w353_ ;
	wire _w354_ ;
	wire _w355_ ;
	wire _w356_ ;
	wire _w357_ ;
	wire _w358_ ;
	wire _w359_ ;
	wire _w360_ ;
	wire _w361_ ;
	wire _w362_ ;
	wire _w363_ ;
	wire _w364_ ;
	wire _w365_ ;
	wire _w366_ ;
	wire _w367_ ;
	wire _w368_ ;
	wire _w369_ ;
	wire _w370_ ;
	wire _w371_ ;
	wire _w372_ ;
	wire _w373_ ;
	wire _w374_ ;
	wire _w375_ ;
	wire _w376_ ;
	wire _w377_ ;
	wire _w378_ ;
	wire _w379_ ;
	wire _w380_ ;
	wire _w381_ ;
	wire _w382_ ;
	wire _w383_ ;
	wire _w384_ ;
	wire _w385_ ;
	wire _w386_ ;
	wire _w387_ ;
	wire _w388_ ;
	wire _w389_ ;
	wire _w390_ ;
	wire _w391_ ;
	wire _w392_ ;
	wire _w393_ ;
	wire _w394_ ;
	wire _w395_ ;
	wire _w396_ ;
	wire _w397_ ;
	wire _w398_ ;
	wire _w399_ ;
	wire _w400_ ;
	wire _w401_ ;
	wire _w402_ ;
	wire _w403_ ;
	wire _w404_ ;
	wire _w405_ ;
	wire _w406_ ;
	wire _w407_ ;
	wire _w408_ ;
	wire _w409_ ;
	wire _w410_ ;
	wire _w411_ ;
	wire _w412_ ;
	wire _w413_ ;
	wire _w414_ ;
	wire _w415_ ;
	wire _w416_ ;
	wire _w417_ ;
	wire _w418_ ;
	wire _w419_ ;
	wire _w420_ ;
	wire _w421_ ;
	wire _w422_ ;
	wire _w423_ ;
	wire _w424_ ;
	wire _w425_ ;
	wire _w426_ ;
	wire _w427_ ;
	wire _w428_ ;
	wire _w429_ ;
	wire _w430_ ;
	wire _w431_ ;
	wire _w432_ ;
	wire _w433_ ;
	wire _w434_ ;
	wire _w435_ ;
	wire _w436_ ;
	wire _w437_ ;
	wire _w438_ ;
	wire _w439_ ;
	wire _w440_ ;
	wire _w441_ ;
	wire _w442_ ;
	wire _w443_ ;
	wire _w444_ ;
	wire _w445_ ;
	wire _w446_ ;
	wire _w447_ ;
	wire _w448_ ;
	wire _w449_ ;
	wire _w450_ ;
	wire _w451_ ;
	wire _w452_ ;
	wire _w453_ ;
	wire _w454_ ;
	wire _w455_ ;
	wire _w456_ ;
	wire _w457_ ;
	wire _w458_ ;
	wire _w459_ ;
	wire _w460_ ;
	wire _w461_ ;
	wire _w462_ ;
	wire _w463_ ;
	wire _w464_ ;
	wire _w465_ ;
	wire _w466_ ;
	wire _w467_ ;
	wire _w468_ ;
	wire _w469_ ;
	wire _w470_ ;
	wire _w471_ ;
	wire _w472_ ;
	wire _w473_ ;
	wire _w474_ ;
	wire _w475_ ;
	wire _w476_ ;
	wire _w477_ ;
	wire _w478_ ;
	wire _w479_ ;
	wire _w480_ ;
	wire _w481_ ;
	wire _w482_ ;
	wire _w483_ ;
	wire _w484_ ;
	wire _w485_ ;
	wire _w486_ ;
	wire _w487_ ;
	wire _w488_ ;
	wire _w489_ ;
	wire _w490_ ;
	wire _w491_ ;
	wire _w492_ ;
	wire _w493_ ;
	wire _w494_ ;
	wire _w495_ ;
	wire _w496_ ;
	wire _w497_ ;
	wire _w498_ ;
	wire _w499_ ;
	wire _w500_ ;
	wire _w501_ ;
	wire _w502_ ;
	wire _w503_ ;
	wire _w504_ ;
	wire _w505_ ;
	wire _w506_ ;
	wire _w507_ ;
	wire _w508_ ;
	wire _w509_ ;
	wire _w510_ ;
	wire _w511_ ;
	wire _w512_ ;
	wire _w513_ ;
	wire _w514_ ;
	wire _w515_ ;
	wire _w516_ ;
	wire _w517_ ;
	wire _w518_ ;
	wire _w519_ ;
	wire _w520_ ;
	wire _w521_ ;
	wire _w522_ ;
	wire _w523_ ;
	wire _w524_ ;
	wire _w525_ ;
	wire _w526_ ;
	wire _w527_ ;
	wire _w528_ ;
	wire _w529_ ;
	wire _w530_ ;
	wire _w531_ ;
	wire _w532_ ;
	wire _w533_ ;
	wire _w534_ ;
	wire _w535_ ;
	wire _w536_ ;
	wire _w537_ ;
	wire _w538_ ;
	wire _w539_ ;
	wire _w540_ ;
	wire _w541_ ;
	wire _w542_ ;
	wire _w543_ ;
	wire _w544_ ;
	wire _w545_ ;
	wire _w546_ ;
	wire _w547_ ;
	wire _w548_ ;
	wire _w549_ ;
	wire _w550_ ;
	wire _w551_ ;
	wire _w552_ ;
	wire _w553_ ;
	wire _w554_ ;
	wire _w555_ ;
	LUT2 #(
		.INIT('h4)
	) name0 (
		\v0_pad ,
		\v10_reg/NET0131 ,
		_w15_
	);
	LUT2 #(
		.INIT('h1)
	) name1 (
		\v12_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w16_
	);
	LUT2 #(
		.INIT('h8)
	) name2 (
		\v4_pad ,
		\v5_pad ,
		_w17_
	);
	LUT2 #(
		.INIT('h8)
	) name3 (
		_w16_,
		_w17_,
		_w18_
	);
	LUT2 #(
		.INIT('h8)
	) name4 (
		\v11_reg/NET0131 ,
		\v12_reg/NET0131 ,
		_w19_
	);
	LUT2 #(
		.INIT('h8)
	) name5 (
		\v8_reg/NET0131 ,
		_w19_,
		_w20_
	);
	LUT2 #(
		.INIT('h4)
	) name6 (
		\v1_pad ,
		\v6_pad ,
		_w21_
	);
	LUT2 #(
		.INIT('h8)
	) name7 (
		\v3_pad ,
		_w21_,
		_w22_
	);
	LUT2 #(
		.INIT('h8)
	) name8 (
		_w20_,
		_w22_,
		_w23_
	);
	LUT2 #(
		.INIT('h1)
	) name9 (
		_w18_,
		_w23_,
		_w24_
	);
	LUT2 #(
		.INIT('h2)
	) name10 (
		_w15_,
		_w24_,
		_w25_
	);
	LUT2 #(
		.INIT('h8)
	) name11 (
		\v12_reg/NET0131 ,
		\v3_pad ,
		_w26_
	);
	LUT2 #(
		.INIT('h8)
	) name12 (
		\v0_pad ,
		\v11_reg/NET0131 ,
		_w27_
	);
	LUT2 #(
		.INIT('h8)
	) name13 (
		\v10_reg/NET0131 ,
		\v8_reg/NET0131 ,
		_w28_
	);
	LUT2 #(
		.INIT('h4)
	) name14 (
		_w21_,
		_w28_,
		_w29_
	);
	LUT2 #(
		.INIT('h8)
	) name15 (
		_w27_,
		_w29_,
		_w30_
	);
	LUT2 #(
		.INIT('h1)
	) name16 (
		\v11_reg/NET0131 ,
		\v8_reg/NET0131 ,
		_w31_
	);
	LUT2 #(
		.INIT('h4)
	) name17 (
		\v9_reg/NET0131 ,
		_w31_,
		_w32_
	);
	LUT2 #(
		.INIT('h4)
	) name18 (
		\v10_reg/NET0131 ,
		_w32_,
		_w33_
	);
	LUT2 #(
		.INIT('h1)
	) name19 (
		_w30_,
		_w33_,
		_w34_
	);
	LUT2 #(
		.INIT('h2)
	) name20 (
		_w26_,
		_w34_,
		_w35_
	);
	LUT2 #(
		.INIT('h8)
	) name21 (
		\v10_reg/NET0131 ,
		\v11_reg/NET0131 ,
		_w36_
	);
	LUT2 #(
		.INIT('h4)
	) name22 (
		\v8_reg/NET0131 ,
		_w36_,
		_w37_
	);
	LUT2 #(
		.INIT('h8)
	) name23 (
		\v9_reg/NET0131 ,
		_w37_,
		_w38_
	);
	LUT2 #(
		.INIT('h2)
	) name24 (
		\v6_pad ,
		\v8_reg/NET0131 ,
		_w39_
	);
	LUT2 #(
		.INIT('h2)
	) name25 (
		\v12_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w40_
	);
	LUT2 #(
		.INIT('h4)
	) name26 (
		\v10_reg/NET0131 ,
		_w40_,
		_w41_
	);
	LUT2 #(
		.INIT('h4)
	) name27 (
		\v11_reg/NET0131 ,
		_w41_,
		_w42_
	);
	LUT2 #(
		.INIT('h8)
	) name28 (
		_w39_,
		_w42_,
		_w43_
	);
	LUT2 #(
		.INIT('h2)
	) name29 (
		\v10_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w44_
	);
	LUT2 #(
		.INIT('h1)
	) name30 (
		\v11_reg/NET0131 ,
		\v12_reg/NET0131 ,
		_w45_
	);
	LUT2 #(
		.INIT('h8)
	) name31 (
		_w44_,
		_w45_,
		_w46_
	);
	LUT2 #(
		.INIT('h1)
	) name32 (
		\v10_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w47_
	);
	LUT2 #(
		.INIT('h2)
	) name33 (
		\v11_reg/NET0131 ,
		\v12_reg/NET0131 ,
		_w48_
	);
	LUT2 #(
		.INIT('h2)
	) name34 (
		\v10_reg/NET0131 ,
		\v2_pad ,
		_w49_
	);
	LUT2 #(
		.INIT('h4)
	) name35 (
		_w17_,
		_w49_,
		_w50_
	);
	LUT2 #(
		.INIT('h2)
	) name36 (
		_w48_,
		_w50_,
		_w51_
	);
	LUT2 #(
		.INIT('h2)
	) name37 (
		\v9_reg/NET0131 ,
		_w51_,
		_w52_
	);
	LUT2 #(
		.INIT('h2)
	) name38 (
		\v8_reg/NET0131 ,
		_w47_,
		_w53_
	);
	LUT2 #(
		.INIT('h4)
	) name39 (
		_w52_,
		_w53_,
		_w54_
	);
	LUT2 #(
		.INIT('h1)
	) name40 (
		_w38_,
		_w46_,
		_w55_
	);
	LUT2 #(
		.INIT('h4)
	) name41 (
		_w43_,
		_w55_,
		_w56_
	);
	LUT2 #(
		.INIT('h4)
	) name42 (
		_w25_,
		_w56_,
		_w57_
	);
	LUT2 #(
		.INIT('h1)
	) name43 (
		_w35_,
		_w54_,
		_w58_
	);
	LUT2 #(
		.INIT('h8)
	) name44 (
		_w57_,
		_w58_,
		_w59_
	);
	LUT2 #(
		.INIT('h1)
	) name45 (
		\v7_reg/NET0131 ,
		_w59_,
		_w60_
	);
	LUT2 #(
		.INIT('h4)
	) name46 (
		\v2_pad ,
		\v8_reg/NET0131 ,
		_w61_
	);
	LUT2 #(
		.INIT('h4)
	) name47 (
		\v9_reg/NET0131 ,
		_w36_,
		_w62_
	);
	LUT2 #(
		.INIT('h8)
	) name48 (
		_w61_,
		_w62_,
		_w63_
	);
	LUT2 #(
		.INIT('h8)
	) name49 (
		\v10_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w64_
	);
	LUT2 #(
		.INIT('h8)
	) name50 (
		_w48_,
		_w64_,
		_w65_
	);
	LUT2 #(
		.INIT('h8)
	) name51 (
		\v7_reg/NET0131 ,
		_w65_,
		_w66_
	);
	LUT2 #(
		.INIT('h8)
	) name52 (
		_w16_,
		_w28_,
		_w67_
	);
	LUT2 #(
		.INIT('h4)
	) name53 (
		\v10_reg/NET0131 ,
		\v7_reg/NET0131 ,
		_w68_
	);
	LUT2 #(
		.INIT('h4)
	) name54 (
		\v11_reg/NET0131 ,
		\v8_reg/NET0131 ,
		_w69_
	);
	LUT2 #(
		.INIT('h4)
	) name55 (
		_w16_,
		_w69_,
		_w70_
	);
	LUT2 #(
		.INIT('h2)
	) name56 (
		\v11_reg/NET0131 ,
		\v8_reg/NET0131 ,
		_w71_
	);
	LUT2 #(
		.INIT('h4)
	) name57 (
		\v12_reg/NET0131 ,
		_w71_,
		_w72_
	);
	LUT2 #(
		.INIT('h1)
	) name58 (
		_w70_,
		_w72_,
		_w73_
	);
	LUT2 #(
		.INIT('h2)
	) name59 (
		_w68_,
		_w73_,
		_w74_
	);
	LUT2 #(
		.INIT('h1)
	) name60 (
		\v10_reg/NET0131 ,
		\v11_reg/NET0131 ,
		_w75_
	);
	LUT2 #(
		.INIT('h4)
	) name61 (
		\v12_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w76_
	);
	LUT2 #(
		.INIT('h4)
	) name62 (
		\v7_reg/NET0131 ,
		_w76_,
		_w77_
	);
	LUT2 #(
		.INIT('h2)
	) name63 (
		\v1_pad ,
		\v2_pad ,
		_w78_
	);
	LUT2 #(
		.INIT('h8)
	) name64 (
		_w39_,
		_w78_,
		_w79_
	);
	LUT2 #(
		.INIT('h8)
	) name65 (
		_w75_,
		_w79_,
		_w80_
	);
	LUT2 #(
		.INIT('h8)
	) name66 (
		_w77_,
		_w80_,
		_w81_
	);
	LUT2 #(
		.INIT('h1)
	) name67 (
		_w63_,
		_w67_,
		_w82_
	);
	LUT2 #(
		.INIT('h4)
	) name68 (
		_w66_,
		_w82_,
		_w83_
	);
	LUT2 #(
		.INIT('h1)
	) name69 (
		_w74_,
		_w81_,
		_w84_
	);
	LUT2 #(
		.INIT('h8)
	) name70 (
		_w83_,
		_w84_,
		_w85_
	);
	LUT2 #(
		.INIT('h4)
	) name71 (
		_w60_,
		_w85_,
		_w86_
	);
	LUT2 #(
		.INIT('h2)
	) name72 (
		CLR_pad,
		_w86_,
		_w87_
	);
	LUT2 #(
		.INIT('h4)
	) name73 (
		\v12_reg/NET0131 ,
		_w17_,
		_w88_
	);
	LUT2 #(
		.INIT('h4)
	) name74 (
		\v0_pad ,
		_w36_,
		_w89_
	);
	LUT2 #(
		.INIT('h1)
	) name75 (
		_w75_,
		_w89_,
		_w90_
	);
	LUT2 #(
		.INIT('h2)
	) name76 (
		_w88_,
		_w90_,
		_w91_
	);
	LUT2 #(
		.INIT('h8)
	) name77 (
		\v10_reg/NET0131 ,
		\v12_reg/NET0131 ,
		_w92_
	);
	LUT2 #(
		.INIT('h4)
	) name78 (
		\v3_pad ,
		_w92_,
		_w93_
	);
	LUT2 #(
		.INIT('h1)
	) name79 (
		\v9_reg/NET0131 ,
		_w93_,
		_w94_
	);
	LUT2 #(
		.INIT('h2)
	) name80 (
		\v2_pad ,
		_w94_,
		_w95_
	);
	LUT2 #(
		.INIT('h1)
	) name81 (
		_w36_,
		_w75_,
		_w96_
	);
	LUT2 #(
		.INIT('h8)
	) name82 (
		\v12_reg/NET0131 ,
		_w96_,
		_w97_
	);
	LUT2 #(
		.INIT('h2)
	) name83 (
		\v12_reg/NET0131 ,
		\v6_pad ,
		_w98_
	);
	LUT2 #(
		.INIT('h4)
	) name84 (
		\v3_pad ,
		_w98_,
		_w99_
	);
	LUT2 #(
		.INIT('h4)
	) name85 (
		\v10_reg/NET0131 ,
		_w99_,
		_w100_
	);
	LUT2 #(
		.INIT('h2)
	) name86 (
		\v10_reg/NET0131 ,
		\v12_reg/NET0131 ,
		_w101_
	);
	LUT2 #(
		.INIT('h4)
	) name87 (
		\v11_reg/NET0131 ,
		_w101_,
		_w102_
	);
	LUT2 #(
		.INIT('h2)
	) name88 (
		\v9_reg/NET0131 ,
		_w102_,
		_w103_
	);
	LUT2 #(
		.INIT('h1)
	) name89 (
		_w97_,
		_w100_,
		_w104_
	);
	LUT2 #(
		.INIT('h4)
	) name90 (
		_w103_,
		_w104_,
		_w105_
	);
	LUT2 #(
		.INIT('h1)
	) name91 (
		_w91_,
		_w95_,
		_w106_
	);
	LUT2 #(
		.INIT('h8)
	) name92 (
		_w105_,
		_w106_,
		_w107_
	);
	LUT2 #(
		.INIT('h1)
	) name93 (
		\v8_reg/NET0131 ,
		_w107_,
		_w108_
	);
	LUT2 #(
		.INIT('h1)
	) name94 (
		\v10_reg/NET0131 ,
		\v1_pad ,
		_w109_
	);
	LUT2 #(
		.INIT('h8)
	) name95 (
		\v2_pad ,
		_w109_,
		_w110_
	);
	LUT2 #(
		.INIT('h1)
	) name96 (
		\v9_reg/NET0131 ,
		_w110_,
		_w111_
	);
	LUT2 #(
		.INIT('h2)
	) name97 (
		_w19_,
		_w111_,
		_w112_
	);
	LUT2 #(
		.INIT('h4)
	) name98 (
		\v12_reg/NET0131 ,
		\v8_reg/NET0131 ,
		_w113_
	);
	LUT2 #(
		.INIT('h8)
	) name99 (
		_w47_,
		_w113_,
		_w114_
	);
	LUT2 #(
		.INIT('h1)
	) name100 (
		_w112_,
		_w114_,
		_w115_
	);
	LUT2 #(
		.INIT('h4)
	) name101 (
		_w108_,
		_w115_,
		_w116_
	);
	LUT2 #(
		.INIT('h1)
	) name102 (
		\v7_reg/NET0131 ,
		_w116_,
		_w117_
	);
	LUT2 #(
		.INIT('h1)
	) name103 (
		\v10_reg/NET0131 ,
		\v12_reg/NET0131 ,
		_w118_
	);
	LUT2 #(
		.INIT('h8)
	) name104 (
		\v3_pad ,
		_w118_,
		_w119_
	);
	LUT2 #(
		.INIT('h1)
	) name105 (
		_w40_,
		_w119_,
		_w120_
	);
	LUT2 #(
		.INIT('h2)
	) name106 (
		_w69_,
		_w120_,
		_w121_
	);
	LUT2 #(
		.INIT('h8)
	) name107 (
		\v10_reg/NET0131 ,
		_w48_,
		_w122_
	);
	LUT2 #(
		.INIT('h8)
	) name108 (
		\v7_reg/NET0131 ,
		_w40_,
		_w123_
	);
	LUT2 #(
		.INIT('h1)
	) name109 (
		_w122_,
		_w123_,
		_w124_
	);
	LUT2 #(
		.INIT('h2)
	) name110 (
		_w61_,
		_w124_,
		_w125_
	);
	LUT2 #(
		.INIT('h1)
	) name111 (
		\v2_pad ,
		\v7_reg/NET0131 ,
		_w126_
	);
	LUT2 #(
		.INIT('h8)
	) name112 (
		\v12_reg/NET0131 ,
		\v1_pad ,
		_w127_
	);
	LUT2 #(
		.INIT('h4)
	) name113 (
		\v10_reg/NET0131 ,
		_w127_,
		_w128_
	);
	LUT2 #(
		.INIT('h8)
	) name114 (
		_w17_,
		_w113_,
		_w129_
	);
	LUT2 #(
		.INIT('h1)
	) name115 (
		_w128_,
		_w129_,
		_w130_
	);
	LUT2 #(
		.INIT('h8)
	) name116 (
		\v11_reg/NET0131 ,
		_w126_,
		_w131_
	);
	LUT2 #(
		.INIT('h4)
	) name117 (
		_w130_,
		_w131_,
		_w132_
	);
	LUT2 #(
		.INIT('h4)
	) name118 (
		\v10_reg/NET0131 ,
		\v8_reg/NET0131 ,
		_w133_
	);
	LUT2 #(
		.INIT('h2)
	) name119 (
		\v11_reg/NET0131 ,
		_w40_,
		_w134_
	);
	LUT2 #(
		.INIT('h2)
	) name120 (
		_w133_,
		_w134_,
		_w135_
	);
	LUT2 #(
		.INIT('h1)
	) name121 (
		\v8_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w136_
	);
	LUT2 #(
		.INIT('h2)
	) name122 (
		_w122_,
		_w136_,
		_w137_
	);
	LUT2 #(
		.INIT('h1)
	) name123 (
		\v10_reg/NET0131 ,
		\v8_reg/NET0131 ,
		_w138_
	);
	LUT2 #(
		.INIT('h8)
	) name124 (
		_w48_,
		_w138_,
		_w139_
	);
	LUT2 #(
		.INIT('h1)
	) name125 (
		_w135_,
		_w139_,
		_w140_
	);
	LUT2 #(
		.INIT('h4)
	) name126 (
		_w137_,
		_w140_,
		_w141_
	);
	LUT2 #(
		.INIT('h2)
	) name127 (
		\v7_reg/NET0131 ,
		_w141_,
		_w142_
	);
	LUT2 #(
		.INIT('h1)
	) name128 (
		_w121_,
		_w125_,
		_w143_
	);
	LUT2 #(
		.INIT('h4)
	) name129 (
		_w132_,
		_w143_,
		_w144_
	);
	LUT2 #(
		.INIT('h4)
	) name130 (
		_w142_,
		_w144_,
		_w145_
	);
	LUT2 #(
		.INIT('h4)
	) name131 (
		_w117_,
		_w145_,
		_w146_
	);
	LUT2 #(
		.INIT('h2)
	) name132 (
		CLR_pad,
		_w146_,
		_w147_
	);
	LUT2 #(
		.INIT('h4)
	) name133 (
		\v11_reg/NET0131 ,
		\v3_pad ,
		_w148_
	);
	LUT2 #(
		.INIT('h8)
	) name134 (
		_w113_,
		_w148_,
		_w149_
	);
	LUT2 #(
		.INIT('h8)
	) name135 (
		_w31_,
		_w76_,
		_w150_
	);
	LUT2 #(
		.INIT('h8)
	) name136 (
		_w19_,
		_w61_,
		_w151_
	);
	LUT2 #(
		.INIT('h1)
	) name137 (
		_w150_,
		_w151_,
		_w152_
	);
	LUT2 #(
		.INIT('h1)
	) name138 (
		\v1_pad ,
		_w152_,
		_w153_
	);
	LUT2 #(
		.INIT('h4)
	) name139 (
		\v6_pad ,
		\v9_reg/NET0131 ,
		_w154_
	);
	LUT2 #(
		.INIT('h8)
	) name140 (
		_w45_,
		_w154_,
		_w155_
	);
	LUT2 #(
		.INIT('h4)
	) name141 (
		\v8_reg/NET0131 ,
		_w155_,
		_w156_
	);
	LUT2 #(
		.INIT('h1)
	) name142 (
		_w149_,
		_w156_,
		_w157_
	);
	LUT2 #(
		.INIT('h4)
	) name143 (
		_w153_,
		_w157_,
		_w158_
	);
	LUT2 #(
		.INIT('h1)
	) name144 (
		\v10_reg/NET0131 ,
		_w158_,
		_w159_
	);
	LUT2 #(
		.INIT('h4)
	) name145 (
		\v10_reg/NET0131 ,
		_w150_,
		_w160_
	);
	LUT2 #(
		.INIT('h8)
	) name146 (
		\v11_reg/NET0131 ,
		_w133_,
		_w161_
	);
	LUT2 #(
		.INIT('h1)
	) name147 (
		\v9_reg/NET0131 ,
		_w127_,
		_w162_
	);
	LUT2 #(
		.INIT('h2)
	) name148 (
		_w161_,
		_w162_,
		_w163_
	);
	LUT2 #(
		.INIT('h1)
	) name149 (
		_w160_,
		_w163_,
		_w164_
	);
	LUT2 #(
		.INIT('h2)
	) name150 (
		\v2_pad ,
		_w164_,
		_w165_
	);
	LUT2 #(
		.INIT('h1)
	) name151 (
		\v12_reg/NET0131 ,
		\v8_reg/NET0131 ,
		_w166_
	);
	LUT2 #(
		.INIT('h8)
	) name152 (
		_w44_,
		_w166_,
		_w167_
	);
	LUT2 #(
		.INIT('h8)
	) name153 (
		\v9_reg/NET0131 ,
		_w161_,
		_w168_
	);
	LUT2 #(
		.INIT('h1)
	) name154 (
		_w167_,
		_w168_,
		_w169_
	);
	LUT2 #(
		.INIT('h1)
	) name155 (
		_w17_,
		_w169_,
		_w170_
	);
	LUT2 #(
		.INIT('h1)
	) name156 (
		\v9_reg/NET0131 ,
		_w92_,
		_w171_
	);
	LUT2 #(
		.INIT('h1)
	) name157 (
		\v8_reg/NET0131 ,
		_w118_,
		_w172_
	);
	LUT2 #(
		.INIT('h8)
	) name158 (
		_w171_,
		_w172_,
		_w173_
	);
	LUT2 #(
		.INIT('h8)
	) name159 (
		_w90_,
		_w173_,
		_w174_
	);
	LUT2 #(
		.INIT('h8)
	) name160 (
		_w18_,
		_w75_,
		_w175_
	);
	LUT2 #(
		.INIT('h8)
	) name161 (
		\v8_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w176_
	);
	LUT2 #(
		.INIT('h2)
	) name162 (
		\v12_reg/NET0131 ,
		_w36_,
		_w177_
	);
	LUT2 #(
		.INIT('h8)
	) name163 (
		_w176_,
		_w177_,
		_w178_
	);
	LUT2 #(
		.INIT('h4)
	) name164 (
		\v11_reg/NET0131 ,
		_w92_,
		_w179_
	);
	LUT2 #(
		.INIT('h8)
	) name165 (
		\v9_reg/NET0131 ,
		_w179_,
		_w180_
	);
	LUT2 #(
		.INIT('h2)
	) name166 (
		\v10_reg/NET0131 ,
		\v11_reg/NET0131 ,
		_w181_
	);
	LUT2 #(
		.INIT('h8)
	) name167 (
		\v2_pad ,
		_w181_,
		_w182_
	);
	LUT2 #(
		.INIT('h8)
	) name168 (
		_w16_,
		_w182_,
		_w183_
	);
	LUT2 #(
		.INIT('h1)
	) name169 (
		_w175_,
		_w178_,
		_w184_
	);
	LUT2 #(
		.INIT('h1)
	) name170 (
		_w180_,
		_w183_,
		_w185_
	);
	LUT2 #(
		.INIT('h8)
	) name171 (
		_w184_,
		_w185_,
		_w186_
	);
	LUT2 #(
		.INIT('h4)
	) name172 (
		_w174_,
		_w186_,
		_w187_
	);
	LUT2 #(
		.INIT('h1)
	) name173 (
		_w165_,
		_w170_,
		_w188_
	);
	LUT2 #(
		.INIT('h8)
	) name174 (
		_w187_,
		_w188_,
		_w189_
	);
	LUT2 #(
		.INIT('h4)
	) name175 (
		_w159_,
		_w189_,
		_w190_
	);
	LUT2 #(
		.INIT('h1)
	) name176 (
		\v7_reg/NET0131 ,
		_w190_,
		_w191_
	);
	LUT2 #(
		.INIT('h8)
	) name177 (
		\v7_reg/NET0131 ,
		\v8_reg/NET0131 ,
		_w192_
	);
	LUT2 #(
		.INIT('h4)
	) name178 (
		_w75_,
		_w192_,
		_w193_
	);
	LUT2 #(
		.INIT('h8)
	) name179 (
		\v2_pad ,
		_w36_,
		_w194_
	);
	LUT2 #(
		.INIT('h1)
	) name180 (
		\v9_reg/NET0131 ,
		_w194_,
		_w195_
	);
	LUT2 #(
		.INIT('h2)
	) name181 (
		\v12_reg/NET0131 ,
		_w195_,
		_w196_
	);
	LUT2 #(
		.INIT('h2)
	) name182 (
		_w193_,
		_w196_,
		_w197_
	);
	LUT2 #(
		.INIT('h8)
	) name183 (
		\v11_reg/NET0131 ,
		\v3_pad ,
		_w198_
	);
	LUT2 #(
		.INIT('h2)
	) name184 (
		_w114_,
		_w198_,
		_w199_
	);
	LUT2 #(
		.INIT('h4)
	) name185 (
		\v12_reg/NET0131 ,
		\v7_reg/NET0131 ,
		_w200_
	);
	LUT2 #(
		.INIT('h2)
	) name186 (
		\v11_reg/NET0131 ,
		_w44_,
		_w201_
	);
	LUT2 #(
		.INIT('h8)
	) name187 (
		_w200_,
		_w201_,
		_w202_
	);
	LUT2 #(
		.INIT('h1)
	) name188 (
		\v7_reg/NET0131 ,
		\v8_reg/NET0131 ,
		_w203_
	);
	LUT2 #(
		.INIT('h8)
	) name189 (
		_w47_,
		_w203_,
		_w204_
	);
	LUT2 #(
		.INIT('h8)
	) name190 (
		_w99_,
		_w204_,
		_w205_
	);
	LUT2 #(
		.INIT('h1)
	) name191 (
		_w199_,
		_w202_,
		_w206_
	);
	LUT2 #(
		.INIT('h4)
	) name192 (
		_w205_,
		_w206_,
		_w207_
	);
	LUT2 #(
		.INIT('h4)
	) name193 (
		_w197_,
		_w207_,
		_w208_
	);
	LUT2 #(
		.INIT('h4)
	) name194 (
		_w191_,
		_w208_,
		_w209_
	);
	LUT2 #(
		.INIT('h2)
	) name195 (
		CLR_pad,
		_w209_,
		_w210_
	);
	LUT2 #(
		.INIT('h8)
	) name196 (
		\v2_pad ,
		_w77_,
		_w211_
	);
	LUT2 #(
		.INIT('h1)
	) name197 (
		_w19_,
		_w31_,
		_w212_
	);
	LUT2 #(
		.INIT('h1)
	) name198 (
		_w113_,
		_w136_,
		_w213_
	);
	LUT2 #(
		.INIT('h8)
	) name199 (
		_w212_,
		_w213_,
		_w214_
	);
	LUT2 #(
		.INIT('h1)
	) name200 (
		_w211_,
		_w214_,
		_w215_
	);
	LUT2 #(
		.INIT('h1)
	) name201 (
		\v10_reg/NET0131 ,
		_w215_,
		_w216_
	);
	LUT2 #(
		.INIT('h8)
	) name202 (
		\v9_reg/NET0131 ,
		_w109_,
		_w217_
	);
	LUT2 #(
		.INIT('h1)
	) name203 (
		_w62_,
		_w217_,
		_w218_
	);
	LUT2 #(
		.INIT('h2)
	) name204 (
		_w166_,
		_w218_,
		_w219_
	);
	LUT2 #(
		.INIT('h4)
	) name205 (
		\v12_reg/NET0131 ,
		_w176_,
		_w220_
	);
	LUT2 #(
		.INIT('h8)
	) name206 (
		_w17_,
		_w220_,
		_w221_
	);
	LUT2 #(
		.INIT('h1)
	) name207 (
		_w67_,
		_w221_,
		_w222_
	);
	LUT2 #(
		.INIT('h1)
	) name208 (
		\v2_pad ,
		_w222_,
		_w223_
	);
	LUT2 #(
		.INIT('h1)
	) name209 (
		\v3_pad ,
		\v9_reg/NET0131 ,
		_w224_
	);
	LUT2 #(
		.INIT('h2)
	) name210 (
		_w48_,
		_w224_,
		_w225_
	);
	LUT2 #(
		.INIT('h2)
	) name211 (
		_w133_,
		_w225_,
		_w226_
	);
	LUT2 #(
		.INIT('h4)
	) name212 (
		\v9_reg/NET0131 ,
		_w98_,
		_w227_
	);
	LUT2 #(
		.INIT('h1)
	) name213 (
		_w92_,
		_w227_,
		_w228_
	);
	LUT2 #(
		.INIT('h1)
	) name214 (
		\v11_reg/NET0131 ,
		_w228_,
		_w229_
	);
	LUT2 #(
		.INIT('h8)
	) name215 (
		\v0_pad ,
		_w21_,
		_w230_
	);
	LUT2 #(
		.INIT('h8)
	) name216 (
		_w26_,
		_w176_,
		_w231_
	);
	LUT2 #(
		.INIT('h4)
	) name217 (
		_w230_,
		_w231_,
		_w232_
	);
	LUT2 #(
		.INIT('h2)
	) name218 (
		\v9_reg/NET0131 ,
		_w48_,
		_w233_
	);
	LUT2 #(
		.INIT('h8)
	) name219 (
		_w96_,
		_w233_,
		_w234_
	);
	LUT2 #(
		.INIT('h4)
	) name220 (
		\v8_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w235_
	);
	LUT2 #(
		.INIT('h4)
	) name221 (
		\v6_pad ,
		_w118_,
		_w236_
	);
	LUT2 #(
		.INIT('h8)
	) name222 (
		_w235_,
		_w236_,
		_w237_
	);
	LUT2 #(
		.INIT('h1)
	) name223 (
		\v7_reg/NET0131 ,
		_w226_,
		_w238_
	);
	LUT2 #(
		.INIT('h1)
	) name224 (
		_w232_,
		_w234_,
		_w239_
	);
	LUT2 #(
		.INIT('h4)
	) name225 (
		_w237_,
		_w239_,
		_w240_
	);
	LUT2 #(
		.INIT('h4)
	) name226 (
		_w219_,
		_w238_,
		_w241_
	);
	LUT2 #(
		.INIT('h4)
	) name227 (
		_w229_,
		_w241_,
		_w242_
	);
	LUT2 #(
		.INIT('h4)
	) name228 (
		_w223_,
		_w240_,
		_w243_
	);
	LUT2 #(
		.INIT('h8)
	) name229 (
		_w242_,
		_w243_,
		_w244_
	);
	LUT2 #(
		.INIT('h8)
	) name230 (
		\v2_pad ,
		_w44_,
		_w245_
	);
	LUT2 #(
		.INIT('h8)
	) name231 (
		_w20_,
		_w245_,
		_w246_
	);
	LUT2 #(
		.INIT('h2)
	) name232 (
		\v11_reg/NET0131 ,
		_w138_,
		_w247_
	);
	LUT2 #(
		.INIT('h1)
	) name233 (
		\v12_reg/NET0131 ,
		_w31_,
		_w248_
	);
	LUT2 #(
		.INIT('h1)
	) name234 (
		_w64_,
		_w133_,
		_w249_
	);
	LUT2 #(
		.INIT('h4)
	) name235 (
		_w247_,
		_w249_,
		_w250_
	);
	LUT2 #(
		.INIT('h8)
	) name236 (
		_w248_,
		_w250_,
		_w251_
	);
	LUT2 #(
		.INIT('h2)
	) name237 (
		\v7_reg/NET0131 ,
		_w246_,
		_w252_
	);
	LUT2 #(
		.INIT('h4)
	) name238 (
		_w251_,
		_w252_,
		_w253_
	);
	LUT2 #(
		.INIT('h1)
	) name239 (
		_w244_,
		_w253_,
		_w254_
	);
	LUT2 #(
		.INIT('h1)
	) name240 (
		_w216_,
		_w254_,
		_w255_
	);
	LUT2 #(
		.INIT('h2)
	) name241 (
		CLR_pad,
		_w255_,
		_w256_
	);
	LUT2 #(
		.INIT('h8)
	) name242 (
		\v12_reg/NET0131 ,
		_w44_,
		_w257_
	);
	LUT2 #(
		.INIT('h1)
	) name243 (
		\v12_reg/NET0131 ,
		_w47_,
		_w258_
	);
	LUT2 #(
		.INIT('h4)
	) name244 (
		_w126_,
		_w258_,
		_w259_
	);
	LUT2 #(
		.INIT('h1)
	) name245 (
		_w257_,
		_w259_,
		_w260_
	);
	LUT2 #(
		.INIT('h2)
	) name246 (
		\v11_reg/NET0131 ,
		_w260_,
		_w261_
	);
	LUT2 #(
		.INIT('h1)
	) name247 (
		_w118_,
		_w171_,
		_w262_
	);
	LUT2 #(
		.INIT('h4)
	) name248 (
		\v11_reg/NET0131 ,
		\v7_reg/NET0131 ,
		_w263_
	);
	LUT2 #(
		.INIT('h4)
	) name249 (
		_w262_,
		_w263_,
		_w264_
	);
	LUT2 #(
		.INIT('h1)
	) name250 (
		_w261_,
		_w264_,
		_w265_
	);
	LUT2 #(
		.INIT('h2)
	) name251 (
		\v8_reg/NET0131 ,
		_w265_,
		_w266_
	);
	LUT2 #(
		.INIT('h1)
	) name252 (
		_w47_,
		_w64_,
		_w267_
	);
	LUT2 #(
		.INIT('h2)
	) name253 (
		_w71_,
		_w267_,
		_w268_
	);
	LUT2 #(
		.INIT('h8)
	) name254 (
		\v11_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w269_
	);
	LUT2 #(
		.INIT('h1)
	) name255 (
		_w203_,
		_w269_,
		_w270_
	);
	LUT2 #(
		.INIT('h2)
	) name256 (
		_w17_,
		_w235_,
		_w271_
	);
	LUT2 #(
		.INIT('h4)
	) name257 (
		_w270_,
		_w271_,
		_w272_
	);
	LUT2 #(
		.INIT('h1)
	) name258 (
		\v7_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w273_
	);
	LUT2 #(
		.INIT('h2)
	) name259 (
		\v8_reg/NET0131 ,
		_w182_,
		_w274_
	);
	LUT2 #(
		.INIT('h1)
	) name260 (
		_w27_,
		_w181_,
		_w275_
	);
	LUT2 #(
		.INIT('h2)
	) name261 (
		_w273_,
		_w275_,
		_w276_
	);
	LUT2 #(
		.INIT('h4)
	) name262 (
		_w274_,
		_w276_,
		_w277_
	);
	LUT2 #(
		.INIT('h1)
	) name263 (
		_w268_,
		_w272_,
		_w278_
	);
	LUT2 #(
		.INIT('h4)
	) name264 (
		_w277_,
		_w278_,
		_w279_
	);
	LUT2 #(
		.INIT('h1)
	) name265 (
		\v12_reg/NET0131 ,
		_w279_,
		_w280_
	);
	LUT2 #(
		.INIT('h1)
	) name266 (
		_w266_,
		_w280_,
		_w281_
	);
	LUT2 #(
		.INIT('h8)
	) name267 (
		_w175_,
		_w203_,
		_w282_
	);
	LUT2 #(
		.INIT('h2)
	) name268 (
		\v12_reg/NET0131 ,
		_w62_,
		_w283_
	);
	LUT2 #(
		.INIT('h2)
	) name269 (
		\v8_reg/NET0131 ,
		_w283_,
		_w284_
	);
	LUT2 #(
		.INIT('h4)
	) name270 (
		\v10_reg/NET0131 ,
		_w48_,
		_w285_
	);
	LUT2 #(
		.INIT('h1)
	) name271 (
		_w284_,
		_w285_,
		_w286_
	);
	LUT2 #(
		.INIT('h2)
	) name272 (
		\v7_reg/NET0131 ,
		_w286_,
		_w287_
	);
	LUT2 #(
		.INIT('h4)
	) name273 (
		_w27_,
		_w273_,
		_w288_
	);
	LUT2 #(
		.INIT('h1)
	) name274 (
		_w269_,
		_w288_,
		_w289_
	);
	LUT2 #(
		.INIT('h2)
	) name275 (
		\v10_reg/NET0131 ,
		_w289_,
		_w290_
	);
	LUT2 #(
		.INIT('h8)
	) name276 (
		\v11_reg/NET0131 ,
		\v8_reg/NET0131 ,
		_w291_
	);
	LUT2 #(
		.INIT('h4)
	) name277 (
		_w47_,
		_w291_,
		_w292_
	);
	LUT2 #(
		.INIT('h1)
	) name278 (
		_w290_,
		_w292_,
		_w293_
	);
	LUT2 #(
		.INIT('h1)
	) name279 (
		\v12_reg/NET0131 ,
		_w293_,
		_w294_
	);
	LUT2 #(
		.INIT('h1)
	) name280 (
		_w287_,
		_w294_,
		_w295_
	);
	LUT2 #(
		.INIT('h2)
	) name281 (
		\v2_pad ,
		_w295_,
		_w296_
	);
	LUT2 #(
		.INIT('h1)
	) name282 (
		_w282_,
		_w296_,
		_w297_
	);
	LUT2 #(
		.INIT('h4)
	) name283 (
		\v4_pad ,
		\v5_pad ,
		_w298_
	);
	LUT2 #(
		.INIT('h1)
	) name284 (
		\v10_reg/NET0131 ,
		_w298_,
		_w299_
	);
	LUT2 #(
		.INIT('h1)
	) name285 (
		\v9_reg/NET0131 ,
		_w299_,
		_w300_
	);
	LUT2 #(
		.INIT('h1)
	) name286 (
		_w247_,
		_w300_,
		_w301_
	);
	LUT2 #(
		.INIT('h1)
	) name287 (
		\v12_reg/NET0131 ,
		_w301_,
		_w302_
	);
	LUT2 #(
		.INIT('h8)
	) name288 (
		\v11_reg/NET0131 ,
		_w47_,
		_w303_
	);
	LUT2 #(
		.INIT('h1)
	) name289 (
		_w302_,
		_w303_,
		_w304_
	);
	LUT2 #(
		.INIT('h2)
	) name290 (
		\v11_reg/NET0131 ,
		\v2_pad ,
		_w305_
	);
	LUT2 #(
		.INIT('h8)
	) name291 (
		\v9_reg/NET0131 ,
		_w305_,
		_w306_
	);
	LUT2 #(
		.INIT('h2)
	) name292 (
		_w274_,
		_w306_,
		_w307_
	);
	LUT2 #(
		.INIT('h1)
	) name293 (
		_w304_,
		_w307_,
		_w308_
	);
	LUT2 #(
		.INIT('h1)
	) name294 (
		\v7_reg/NET0131 ,
		_w308_,
		_w309_
	);
	LUT2 #(
		.INIT('h2)
	) name295 (
		\v9_reg/NET0131 ,
		_w75_,
		_w310_
	);
	LUT2 #(
		.INIT('h2)
	) name296 (
		\v8_reg/NET0131 ,
		_w310_,
		_w311_
	);
	LUT2 #(
		.INIT('h8)
	) name297 (
		\v7_reg/NET0131 ,
		_w47_,
		_w312_
	);
	LUT2 #(
		.INIT('h1)
	) name298 (
		\v12_reg/NET0131 ,
		_w312_,
		_w313_
	);
	LUT2 #(
		.INIT('h4)
	) name299 (
		_w42_,
		_w311_,
		_w314_
	);
	LUT2 #(
		.INIT('h4)
	) name300 (
		_w313_,
		_w314_,
		_w315_
	);
	LUT2 #(
		.INIT('h1)
	) name301 (
		_w309_,
		_w315_,
		_w316_
	);
	LUT2 #(
		.INIT('h4)
	) name302 (
		_w90_,
		_w136_,
		_w317_
	);
	LUT2 #(
		.INIT('h8)
	) name303 (
		_w176_,
		_w305_,
		_w318_
	);
	LUT2 #(
		.INIT('h1)
	) name304 (
		_w317_,
		_w318_,
		_w319_
	);
	LUT2 #(
		.INIT('h1)
	) name305 (
		\v12_reg/NET0131 ,
		\v7_reg/NET0131 ,
		_w320_
	);
	LUT2 #(
		.INIT('h2)
	) name306 (
		\v4_pad ,
		\v5_pad ,
		_w321_
	);
	LUT2 #(
		.INIT('h8)
	) name307 (
		_w320_,
		_w321_,
		_w322_
	);
	LUT2 #(
		.INIT('h4)
	) name308 (
		_w319_,
		_w322_,
		_w323_
	);
	LUT2 #(
		.INIT('h8)
	) name309 (
		_w26_,
		_w269_,
		_w324_
	);
	LUT2 #(
		.INIT('h4)
	) name310 (
		\v7_reg/NET0131 ,
		_w29_,
		_w325_
	);
	LUT2 #(
		.INIT('h8)
	) name311 (
		_w324_,
		_w325_,
		_w326_
	);
	LUT2 #(
		.INIT('h8)
	) name312 (
		_w17_,
		_w291_,
		_w327_
	);
	LUT2 #(
		.INIT('h1)
	) name313 (
		_w31_,
		_w327_,
		_w328_
	);
	LUT2 #(
		.INIT('h2)
	) name314 (
		_w77_,
		_w328_,
		_w329_
	);
	LUT2 #(
		.INIT('h8)
	) name315 (
		_w40_,
		_w192_,
		_w330_
	);
	LUT2 #(
		.INIT('h1)
	) name316 (
		_w329_,
		_w330_,
		_w331_
	);
	LUT2 #(
		.INIT('h1)
	) name317 (
		\v2_pad ,
		_w331_,
		_w332_
	);
	LUT2 #(
		.INIT('h8)
	) name318 (
		_w15_,
		_w136_,
		_w333_
	);
	LUT2 #(
		.INIT('h8)
	) name319 (
		_w88_,
		_w333_,
		_w334_
	);
	LUT2 #(
		.INIT('h1)
	) name320 (
		\v8_reg/NET0131 ,
		_w101_,
		_w335_
	);
	LUT2 #(
		.INIT('h8)
	) name321 (
		\v9_reg/NET0131 ,
		_w335_,
		_w336_
	);
	LUT2 #(
		.INIT('h1)
	) name322 (
		_w334_,
		_w336_,
		_w337_
	);
	LUT2 #(
		.INIT('h2)
	) name323 (
		\v11_reg/NET0131 ,
		_w337_,
		_w338_
	);
	LUT2 #(
		.INIT('h8)
	) name324 (
		_w76_,
		_w181_,
		_w339_
	);
	LUT2 #(
		.INIT('h1)
	) name325 (
		_w155_,
		_w339_,
		_w340_
	);
	LUT2 #(
		.INIT('h1)
	) name326 (
		\v8_reg/NET0131 ,
		_w340_,
		_w341_
	);
	LUT2 #(
		.INIT('h4)
	) name327 (
		\v12_reg/NET0131 ,
		\v1_pad ,
		_w342_
	);
	LUT2 #(
		.INIT('h4)
	) name328 (
		_w21_,
		_w36_,
		_w343_
	);
	LUT2 #(
		.INIT('h1)
	) name329 (
		_w342_,
		_w343_,
		_w344_
	);
	LUT2 #(
		.INIT('h2)
	) name330 (
		\v3_pad ,
		_w344_,
		_w345_
	);
	LUT2 #(
		.INIT('h8)
	) name331 (
		_w31_,
		_w92_,
		_w346_
	);
	LUT2 #(
		.INIT('h2)
	) name332 (
		\v9_reg/NET0131 ,
		_w248_,
		_w347_
	);
	LUT2 #(
		.INIT('h4)
	) name333 (
		_w346_,
		_w347_,
		_w348_
	);
	LUT2 #(
		.INIT('h4)
	) name334 (
		_w345_,
		_w348_,
		_w349_
	);
	LUT2 #(
		.INIT('h1)
	) name335 (
		_w338_,
		_w341_,
		_w350_
	);
	LUT2 #(
		.INIT('h4)
	) name336 (
		_w349_,
		_w350_,
		_w351_
	);
	LUT2 #(
		.INIT('h1)
	) name337 (
		\v7_reg/NET0131 ,
		_w351_,
		_w352_
	);
	LUT2 #(
		.INIT('h4)
	) name338 (
		_w16_,
		_w192_,
		_w353_
	);
	LUT2 #(
		.INIT('h4)
	) name339 (
		_w62_,
		_w353_,
		_w354_
	);
	LUT2 #(
		.INIT('h4)
	) name340 (
		_w310_,
		_w354_,
		_w355_
	);
	LUT2 #(
		.INIT('h1)
	) name341 (
		_w332_,
		_w355_,
		_w356_
	);
	LUT2 #(
		.INIT('h4)
	) name342 (
		_w352_,
		_w356_,
		_w357_
	);
	LUT2 #(
		.INIT('h2)
	) name343 (
		CLR_pad,
		_w357_,
		_w358_
	);
	LUT2 #(
		.INIT('h4)
	) name344 (
		\v12_reg/NET0131 ,
		\v2_pad ,
		_w359_
	);
	LUT2 #(
		.INIT('h1)
	) name345 (
		\v11_reg/NET0131 ,
		_w359_,
		_w360_
	);
	LUT2 #(
		.INIT('h2)
	) name346 (
		\v10_reg/NET0131 ,
		_w360_,
		_w361_
	);
	LUT2 #(
		.INIT('h1)
	) name347 (
		\v9_reg/NET0131 ,
		_w361_,
		_w362_
	);
	LUT2 #(
		.INIT('h2)
	) name348 (
		_w17_,
		_w19_,
		_w363_
	);
	LUT2 #(
		.INIT('h1)
	) name349 (
		\v10_reg/NET0131 ,
		_w363_,
		_w364_
	);
	LUT2 #(
		.INIT('h4)
	) name350 (
		_w230_,
		_w324_,
		_w365_
	);
	LUT2 #(
		.INIT('h1)
	) name351 (
		_w155_,
		_w364_,
		_w366_
	);
	LUT2 #(
		.INIT('h4)
	) name352 (
		_w365_,
		_w366_,
		_w367_
	);
	LUT2 #(
		.INIT('h4)
	) name353 (
		_w362_,
		_w367_,
		_w368_
	);
	LUT2 #(
		.INIT('h2)
	) name354 (
		\v8_reg/NET0131 ,
		_w368_,
		_w369_
	);
	LUT2 #(
		.INIT('h4)
	) name355 (
		\v10_reg/NET0131 ,
		\v12_reg/NET0131 ,
		_w370_
	);
	LUT2 #(
		.INIT('h1)
	) name356 (
		_w220_,
		_w370_,
		_w371_
	);
	LUT2 #(
		.INIT('h1)
	) name357 (
		\v3_pad ,
		_w371_,
		_w372_
	);
	LUT2 #(
		.INIT('h4)
	) name358 (
		\v10_reg/NET0131 ,
		_w18_,
		_w373_
	);
	LUT2 #(
		.INIT('h1)
	) name359 (
		_w372_,
		_w373_,
		_w374_
	);
	LUT2 #(
		.INIT('h1)
	) name360 (
		\v11_reg/NET0131 ,
		_w374_,
		_w375_
	);
	LUT2 #(
		.INIT('h8)
	) name361 (
		_w37_,
		_w40_,
		_w376_
	);
	LUT2 #(
		.INIT('h2)
	) name362 (
		\v10_reg/NET0131 ,
		_w235_,
		_w377_
	);
	LUT2 #(
		.INIT('h4)
	) name363 (
		_w138_,
		_w359_,
		_w378_
	);
	LUT2 #(
		.INIT('h4)
	) name364 (
		_w377_,
		_w378_,
		_w379_
	);
	LUT2 #(
		.INIT('h4)
	) name365 (
		\v11_reg/NET0131 ,
		\v6_pad ,
		_w380_
	);
	LUT2 #(
		.INIT('h1)
	) name366 (
		\v9_reg/NET0131 ,
		_w380_,
		_w381_
	);
	LUT2 #(
		.INIT('h8)
	) name367 (
		\v12_reg/NET0131 ,
		_w138_,
		_w382_
	);
	LUT2 #(
		.INIT('h4)
	) name368 (
		_w381_,
		_w382_,
		_w383_
	);
	LUT2 #(
		.INIT('h1)
	) name369 (
		_w376_,
		_w379_,
		_w384_
	);
	LUT2 #(
		.INIT('h4)
	) name370 (
		_w383_,
		_w384_,
		_w385_
	);
	LUT2 #(
		.INIT('h4)
	) name371 (
		_w375_,
		_w385_,
		_w386_
	);
	LUT2 #(
		.INIT('h4)
	) name372 (
		_w369_,
		_w386_,
		_w387_
	);
	LUT2 #(
		.INIT('h1)
	) name373 (
		\v7_reg/NET0131 ,
		_w387_,
		_w388_
	);
	LUT2 #(
		.INIT('h8)
	) name374 (
		_w200_,
		_w269_,
		_w389_
	);
	LUT2 #(
		.INIT('h2)
	) name375 (
		\v10_reg/NET0131 ,
		_w40_,
		_w390_
	);
	LUT2 #(
		.INIT('h4)
	) name376 (
		_w41_,
		_w69_,
		_w391_
	);
	LUT2 #(
		.INIT('h4)
	) name377 (
		_w390_,
		_w391_,
		_w392_
	);
	LUT2 #(
		.INIT('h1)
	) name378 (
		_w389_,
		_w392_,
		_w393_
	);
	LUT2 #(
		.INIT('h4)
	) name379 (
		_w388_,
		_w393_,
		_w394_
	);
	LUT2 #(
		.INIT('h2)
	) name380 (
		CLR_pad,
		_w394_,
		_w395_
	);
	LUT2 #(
		.INIT('h8)
	) name381 (
		\v3_pad ,
		_w380_,
		_w396_
	);
	LUT2 #(
		.INIT('h1)
	) name382 (
		_w305_,
		_w396_,
		_w397_
	);
	LUT2 #(
		.INIT('h2)
	) name383 (
		\v8_reg/NET0131 ,
		_w397_,
		_w398_
	);
	LUT2 #(
		.INIT('h8)
	) name384 (
		_w136_,
		_w275_,
		_w399_
	);
	LUT2 #(
		.INIT('h1)
	) name385 (
		_w398_,
		_w399_,
		_w400_
	);
	LUT2 #(
		.INIT('h2)
	) name386 (
		_w17_,
		_w69_,
		_w401_
	);
	LUT2 #(
		.INIT('h1)
	) name387 (
		\v12_reg/NET0131 ,
		_w401_,
		_w402_
	);
	LUT2 #(
		.INIT('h4)
	) name388 (
		_w400_,
		_w402_,
		_w403_
	);
	LUT2 #(
		.INIT('h1)
	) name389 (
		\v7_reg/NET0131 ,
		_w403_,
		_w404_
	);
	LUT2 #(
		.INIT('h1)
	) name390 (
		_w139_,
		_w311_,
		_w405_
	);
	LUT2 #(
		.INIT('h4)
	) name391 (
		_w404_,
		_w405_,
		_w406_
	);
	LUT2 #(
		.INIT('h4)
	) name392 (
		\v10_reg/NET0131 ,
		_w17_,
		_w407_
	);
	LUT2 #(
		.INIT('h1)
	) name393 (
		_w27_,
		_w407_,
		_w408_
	);
	LUT2 #(
		.INIT('h1)
	) name394 (
		\v12_reg/NET0131 ,
		_w408_,
		_w409_
	);
	LUT2 #(
		.INIT('h1)
	) name395 (
		_w179_,
		_w409_,
		_w410_
	);
	LUT2 #(
		.INIT('h1)
	) name396 (
		\v9_reg/NET0131 ,
		_w410_,
		_w411_
	);
	LUT2 #(
		.INIT('h1)
	) name397 (
		_w65_,
		_w411_,
		_w412_
	);
	LUT2 #(
		.INIT('h1)
	) name398 (
		\v7_reg/NET0131 ,
		_w412_,
		_w413_
	);
	LUT2 #(
		.INIT('h4)
	) name399 (
		\v9_reg/NET0131 ,
		_w285_,
		_w414_
	);
	LUT2 #(
		.INIT('h1)
	) name400 (
		_w413_,
		_w414_,
		_w415_
	);
	LUT2 #(
		.INIT('h1)
	) name401 (
		\v8_reg/NET0131 ,
		_w415_,
		_w416_
	);
	LUT2 #(
		.INIT('h4)
	) name402 (
		_w47_,
		_w359_,
		_w417_
	);
	LUT2 #(
		.INIT('h1)
	) name403 (
		_w257_,
		_w417_,
		_w418_
	);
	LUT2 #(
		.INIT('h2)
	) name404 (
		\v11_reg/NET0131 ,
		_w418_,
		_w419_
	);
	LUT2 #(
		.INIT('h1)
	) name405 (
		_w200_,
		_w419_,
		_w420_
	);
	LUT2 #(
		.INIT('h2)
	) name406 (
		\v8_reg/NET0131 ,
		_w420_,
		_w421_
	);
	LUT2 #(
		.INIT('h1)
	) name407 (
		_w416_,
		_w421_,
		_w422_
	);
	LUT2 #(
		.INIT('h1)
	) name408 (
		_w291_,
		_w320_,
		_w423_
	);
	LUT2 #(
		.INIT('h1)
	) name409 (
		\v1_pad ,
		_w423_,
		_w424_
	);
	LUT2 #(
		.INIT('h1)
	) name410 (
		_w20_,
		_w424_,
		_w425_
	);
	LUT2 #(
		.INIT('h1)
	) name411 (
		\v9_reg/NET0131 ,
		_w425_,
		_w426_
	);
	LUT2 #(
		.INIT('h8)
	) name412 (
		\v9_reg/NET0131 ,
		_w48_,
		_w427_
	);
	LUT2 #(
		.INIT('h8)
	) name413 (
		\v1_pad ,
		_w427_,
		_w428_
	);
	LUT2 #(
		.INIT('h1)
	) name414 (
		_w426_,
		_w428_,
		_w429_
	);
	LUT2 #(
		.INIT('h2)
	) name415 (
		\v10_reg/NET0131 ,
		_w429_,
		_w430_
	);
	LUT2 #(
		.INIT('h4)
	) name416 (
		_w19_,
		_w47_,
		_w431_
	);
	LUT2 #(
		.INIT('h1)
	) name417 (
		_w339_,
		_w431_,
		_w432_
	);
	LUT2 #(
		.INIT('h2)
	) name418 (
		\v8_reg/NET0131 ,
		_w432_,
		_w433_
	);
	LUT2 #(
		.INIT('h2)
	) name419 (
		\v7_reg/NET0131 ,
		_w139_,
		_w434_
	);
	LUT2 #(
		.INIT('h4)
	) name420 (
		_w433_,
		_w434_,
		_w435_
	);
	LUT2 #(
		.INIT('h2)
	) name421 (
		\v11_reg/NET0131 ,
		_w15_,
		_w436_
	);
	LUT2 #(
		.INIT('h2)
	) name422 (
		_w136_,
		_w436_,
		_w437_
	);
	LUT2 #(
		.INIT('h1)
	) name423 (
		_w318_,
		_w437_,
		_w438_
	);
	LUT2 #(
		.INIT('h2)
	) name424 (
		_w17_,
		_w438_,
		_w439_
	);
	LUT2 #(
		.INIT('h8)
	) name425 (
		\v2_pad ,
		_w292_,
		_w440_
	);
	LUT2 #(
		.INIT('h1)
	) name426 (
		_w439_,
		_w440_,
		_w441_
	);
	LUT2 #(
		.INIT('h1)
	) name427 (
		\v12_reg/NET0131 ,
		_w441_,
		_w442_
	);
	LUT2 #(
		.INIT('h1)
	) name428 (
		_w45_,
		_w172_,
		_w443_
	);
	LUT2 #(
		.INIT('h4)
	) name429 (
		\v9_reg/NET0131 ,
		_w96_,
		_w444_
	);
	LUT2 #(
		.INIT('h4)
	) name430 (
		_w443_,
		_w444_,
		_w445_
	);
	LUT2 #(
		.INIT('h1)
	) name431 (
		\v7_reg/NET0131 ,
		_w445_,
		_w446_
	);
	LUT2 #(
		.INIT('h4)
	) name432 (
		_w442_,
		_w446_,
		_w447_
	);
	LUT2 #(
		.INIT('h1)
	) name433 (
		_w435_,
		_w447_,
		_w448_
	);
	LUT2 #(
		.INIT('h1)
	) name434 (
		_w430_,
		_w448_,
		_w449_
	);
	LUT2 #(
		.INIT('h4)
	) name435 (
		_w200_,
		_w310_,
		_w450_
	);
	LUT2 #(
		.INIT('h2)
	) name436 (
		\v8_reg/NET0131 ,
		_w450_,
		_w451_
	);
	LUT2 #(
		.INIT('h1)
	) name437 (
		\v9_reg/NET0131 ,
		_w436_,
		_w452_
	);
	LUT2 #(
		.INIT('h1)
	) name438 (
		\v8_reg/NET0131 ,
		_w452_,
		_w453_
	);
	LUT2 #(
		.INIT('h1)
	) name439 (
		\v4_pad ,
		\v5_pad ,
		_w454_
	);
	LUT2 #(
		.INIT('h8)
	) name440 (
		\v2_pad ,
		\v8_reg/NET0131 ,
		_w455_
	);
	LUT2 #(
		.INIT('h1)
	) name441 (
		\v12_reg/NET0131 ,
		_w17_,
		_w456_
	);
	LUT2 #(
		.INIT('h1)
	) name442 (
		_w181_,
		_w454_,
		_w457_
	);
	LUT2 #(
		.INIT('h4)
	) name443 (
		_w455_,
		_w457_,
		_w458_
	);
	LUT2 #(
		.INIT('h8)
	) name444 (
		_w456_,
		_w458_,
		_w459_
	);
	LUT2 #(
		.INIT('h4)
	) name445 (
		_w453_,
		_w459_,
		_w460_
	);
	LUT2 #(
		.INIT('h1)
	) name446 (
		\v7_reg/NET0131 ,
		_w460_,
		_w461_
	);
	LUT2 #(
		.INIT('h1)
	) name447 (
		_w202_,
		_w451_,
		_w462_
	);
	LUT2 #(
		.INIT('h4)
	) name448 (
		_w461_,
		_w462_,
		_w463_
	);
	LUT2 #(
		.INIT('h8)
	) name449 (
		_w77_,
		_w396_,
		_w464_
	);
	LUT2 #(
		.INIT('h8)
	) name450 (
		\v11_reg/NET0131 ,
		\v2_pad ,
		_w465_
	);
	LUT2 #(
		.INIT('h8)
	) name451 (
		_w123_,
		_w465_,
		_w466_
	);
	LUT2 #(
		.INIT('h1)
	) name452 (
		_w464_,
		_w466_,
		_w467_
	);
	LUT2 #(
		.INIT('h2)
	) name453 (
		_w28_,
		_w467_,
		_w468_
	);
	LUT2 #(
		.INIT('h4)
	) name454 (
		\v2_pad ,
		\v9_reg/NET0131 ,
		_w469_
	);
	LUT2 #(
		.INIT('h8)
	) name455 (
		\v8_reg/NET0131 ,
		_w469_,
		_w470_
	);
	LUT2 #(
		.INIT('h1)
	) name456 (
		_w333_,
		_w470_,
		_w471_
	);
	LUT2 #(
		.INIT('h2)
	) name457 (
		\v11_reg/NET0131 ,
		_w454_,
		_w472_
	);
	LUT2 #(
		.INIT('h4)
	) name458 (
		_w471_,
		_w472_,
		_w473_
	);
	LUT2 #(
		.INIT('h8)
	) name459 (
		_w32_,
		_w407_,
		_w474_
	);
	LUT2 #(
		.INIT('h1)
	) name460 (
		_w473_,
		_w474_,
		_w475_
	);
	LUT2 #(
		.INIT('h2)
	) name461 (
		_w320_,
		_w475_,
		_w476_
	);
	LUT2 #(
		.INIT('h8)
	) name462 (
		_w28_,
		_w466_,
		_w477_
	);
	LUT2 #(
		.INIT('h8)
	) name463 (
		_w138_,
		_w227_,
		_w478_
	);
	LUT2 #(
		.INIT('h8)
	) name464 (
		\v6_pad ,
		_w101_,
		_w479_
	);
	LUT2 #(
		.INIT('h8)
	) name465 (
		_w176_,
		_w479_,
		_w480_
	);
	LUT2 #(
		.INIT('h1)
	) name466 (
		_w478_,
		_w480_,
		_w481_
	);
	LUT2 #(
		.INIT('h4)
	) name467 (
		\v7_reg/NET0131 ,
		_w148_,
		_w482_
	);
	LUT2 #(
		.INIT('h4)
	) name468 (
		_w481_,
		_w482_,
		_w483_
	);
	LUT2 #(
		.INIT('h1)
	) name469 (
		_w477_,
		_w483_,
		_w484_
	);
	LUT2 #(
		.INIT('h8)
	) name470 (
		_w17_,
		_w32_,
		_w485_
	);
	LUT2 #(
		.INIT('h8)
	) name471 (
		\v2_pad ,
		_w176_,
		_w486_
	);
	LUT2 #(
		.INIT('h1)
	) name472 (
		_w485_,
		_w486_,
		_w487_
	);
	LUT2 #(
		.INIT('h4)
	) name473 (
		\v7_reg/NET0131 ,
		_w118_,
		_w488_
	);
	LUT2 #(
		.INIT('h4)
	) name474 (
		_w487_,
		_w488_,
		_w489_
	);
	LUT2 #(
		.INIT('h8)
	) name475 (
		\v7_reg/NET0131 ,
		_w176_,
		_w490_
	);
	LUT2 #(
		.INIT('h8)
	) name476 (
		_w102_,
		_w490_,
		_w491_
	);
	LUT2 #(
		.INIT('h8)
	) name477 (
		_w45_,
		_w61_,
		_w492_
	);
	LUT2 #(
		.INIT('h8)
	) name478 (
		\v12_reg/NET0131 ,
		_w235_,
		_w493_
	);
	LUT2 #(
		.INIT('h1)
	) name479 (
		_w492_,
		_w493_,
		_w494_
	);
	LUT2 #(
		.INIT('h1)
	) name480 (
		\v10_reg/NET0131 ,
		\v7_reg/NET0131 ,
		_w495_
	);
	LUT2 #(
		.INIT('h4)
	) name481 (
		_w494_,
		_w495_,
		_w496_
	);
	LUT2 #(
		.INIT('h1)
	) name482 (
		_w491_,
		_w496_,
		_w497_
	);
	LUT2 #(
		.INIT('h8)
	) name483 (
		_w370_,
		_w380_,
		_w498_
	);
	LUT2 #(
		.INIT('h8)
	) name484 (
		\v0_pad ,
		_w122_,
		_w499_
	);
	LUT2 #(
		.INIT('h1)
	) name485 (
		_w498_,
		_w499_,
		_w500_
	);
	LUT2 #(
		.INIT('h1)
	) name486 (
		\v9_reg/NET0131 ,
		_w500_,
		_w501_
	);
	LUT2 #(
		.INIT('h8)
	) name487 (
		_w19_,
		_w64_,
		_w502_
	);
	LUT2 #(
		.INIT('h1)
	) name488 (
		_w501_,
		_w502_,
		_w503_
	);
	LUT2 #(
		.INIT('h2)
	) name489 (
		_w203_,
		_w503_,
		_w504_
	);
	LUT2 #(
		.INIT('h4)
	) name490 (
		\v5_pad ,
		_w45_,
		_w505_
	);
	LUT2 #(
		.INIT('h1)
	) name491 (
		_w19_,
		_w505_,
		_w506_
	);
	LUT2 #(
		.INIT('h1)
	) name492 (
		\v10_reg/NET0131 ,
		_w506_,
		_w507_
	);
	LUT2 #(
		.INIT('h1)
	) name493 (
		_w179_,
		_w507_,
		_w508_
	);
	LUT2 #(
		.INIT('h2)
	) name494 (
		_w136_,
		_w508_,
		_w509_
	);
	LUT2 #(
		.INIT('h8)
	) name495 (
		_w148_,
		_w480_,
		_w510_
	);
	LUT2 #(
		.INIT('h1)
	) name496 (
		_w509_,
		_w510_,
		_w511_
	);
	LUT2 #(
		.INIT('h1)
	) name497 (
		\v7_reg/NET0131 ,
		_w511_,
		_w512_
	);
	LUT2 #(
		.INIT('h2)
	) name498 (
		\v10_reg/NET0131 ,
		_w176_,
		_w513_
	);
	LUT2 #(
		.INIT('h4)
	) name499 (
		\v10_reg/NET0131 ,
		_w176_,
		_w514_
	);
	LUT2 #(
		.INIT('h2)
	) name500 (
		_w200_,
		_w513_,
		_w515_
	);
	LUT2 #(
		.INIT('h4)
	) name501 (
		_w514_,
		_w515_,
		_w516_
	);
	LUT2 #(
		.INIT('h4)
	) name502 (
		\v5_pad ,
		_w76_,
		_w517_
	);
	LUT2 #(
		.INIT('h1)
	) name503 (
		_w123_,
		_w517_,
		_w518_
	);
	LUT2 #(
		.INIT('h2)
	) name504 (
		_w61_,
		_w68_,
		_w519_
	);
	LUT2 #(
		.INIT('h4)
	) name505 (
		_w518_,
		_w519_,
		_w520_
	);
	LUT2 #(
		.INIT('h1)
	) name506 (
		_w516_,
		_w520_,
		_w521_
	);
	LUT2 #(
		.INIT('h2)
	) name507 (
		\v11_reg/NET0131 ,
		_w521_,
		_w522_
	);
	LUT2 #(
		.INIT('h8)
	) name508 (
		_w61_,
		_w68_,
		_w523_
	);
	LUT2 #(
		.INIT('h4)
	) name509 (
		\v5_pad ,
		_w36_,
		_w524_
	);
	LUT2 #(
		.INIT('h8)
	) name510 (
		_w203_,
		_w524_,
		_w525_
	);
	LUT2 #(
		.INIT('h1)
	) name511 (
		_w523_,
		_w525_,
		_w526_
	);
	LUT2 #(
		.INIT('h4)
	) name512 (
		\v0_pad ,
		_w16_,
		_w527_
	);
	LUT2 #(
		.INIT('h4)
	) name513 (
		_w526_,
		_w527_,
		_w528_
	);
	LUT2 #(
		.INIT('h1)
	) name514 (
		_w522_,
		_w528_,
		_w529_
	);
	LUT2 #(
		.INIT('h4)
	) name515 (
		_w512_,
		_w529_,
		_w530_
	);
	LUT2 #(
		.INIT('h1)
	) name516 (
		_w41_,
		_w258_,
		_w531_
	);
	LUT2 #(
		.INIT('h2)
	) name517 (
		_w69_,
		_w531_,
		_w532_
	);
	LUT2 #(
		.INIT('h4)
	) name518 (
		_w133_,
		_w427_,
		_w533_
	);
	LUT2 #(
		.INIT('h1)
	) name519 (
		_w532_,
		_w533_,
		_w534_
	);
	LUT2 #(
		.INIT('h2)
	) name520 (
		\v7_reg/NET0131 ,
		_w534_,
		_w535_
	);
	LUT2 #(
		.INIT('h8)
	) name521 (
		_w181_,
		_w359_,
		_w536_
	);
	LUT2 #(
		.INIT('h1)
	) name522 (
		_w19_,
		_w101_,
		_w537_
	);
	LUT2 #(
		.INIT('h1)
	) name523 (
		\v8_reg/NET0131 ,
		_w36_,
		_w538_
	);
	LUT2 #(
		.INIT('h4)
	) name524 (
		_w537_,
		_w538_,
		_w539_
	);
	LUT2 #(
		.INIT('h1)
	) name525 (
		_w536_,
		_w539_,
		_w540_
	);
	LUT2 #(
		.INIT('h1)
	) name526 (
		\v9_reg/NET0131 ,
		_w540_,
		_w541_
	);
	LUT2 #(
		.INIT('h1)
	) name527 (
		_w318_,
		_w333_,
		_w542_
	);
	LUT2 #(
		.INIT('h1)
	) name528 (
		\v12_reg/NET0131 ,
		_w298_,
		_w543_
	);
	LUT2 #(
		.INIT('h4)
	) name529 (
		_w542_,
		_w543_,
		_w544_
	);
	LUT2 #(
		.INIT('h1)
	) name530 (
		_w541_,
		_w544_,
		_w545_
	);
	LUT2 #(
		.INIT('h1)
	) name531 (
		\v7_reg/NET0131 ,
		_w545_,
		_w546_
	);
	LUT2 #(
		.INIT('h1)
	) name532 (
		_w535_,
		_w546_,
		_w547_
	);
	LUT2 #(
		.INIT('h1)
	) name533 (
		_w71_,
		_w469_,
		_w548_
	);
	LUT2 #(
		.INIT('h1)
	) name534 (
		_w298_,
		_w548_,
		_w549_
	);
	LUT2 #(
		.INIT('h1)
	) name535 (
		\v0_pad ,
		\v12_reg/NET0131 ,
		_w550_
	);
	LUT2 #(
		.INIT('h2)
	) name536 (
		\v11_reg/NET0131 ,
		_w550_,
		_w551_
	);
	LUT2 #(
		.INIT('h1)
	) name537 (
		\v9_reg/NET0131 ,
		_w102_,
		_w552_
	);
	LUT2 #(
		.INIT('h4)
	) name538 (
		_w551_,
		_w552_,
		_w553_
	);
	LUT2 #(
		.INIT('h1)
	) name539 (
		\v8_reg/NET0131 ,
		_w553_,
		_w554_
	);
	LUT2 #(
		.INIT('h4)
	) name540 (
		_w45_,
		_w47_,
		_w555_
	);
	LUT2 #(
		.INIT('h4)
	) name541 (
		\v2_pad ,
		_w101_,
		_w556_
	);
	LUT2 #(
		.INIT('h1)
	) name542 (
		\v11_reg/NET0131 ,
		_w335_,
		_w557_
	);
	LUT2 #(
		.INIT('h4)
	) name543 (
		_w556_,
		_w557_,
		_w558_
	);
	LUT2 #(
		.INIT('h1)
	) name544 (
		\v7_reg/NET0131 ,
		_w233_,
		_w559_
	);
	LUT2 #(
		.INIT('h4)
	) name545 (
		_w555_,
		_w559_,
		_w560_
	);
	LUT2 #(
		.INIT('h4)
	) name546 (
		_w549_,
		_w560_,
		_w561_
	);
	LUT2 #(
		.INIT('h4)
	) name547 (
		_w558_,
		_w561_,
		_w562_
	);
	LUT2 #(
		.INIT('h4)
	) name548 (
		_w554_,
		_w562_,
		_w563_
	);
	LUT2 #(
		.INIT('h2)
	) name549 (
		\v9_reg/NET0131 ,
		_w45_,
		_w564_
	);
	LUT2 #(
		.INIT('h4)
	) name550 (
		_w19_,
		_w28_,
		_w565_
	);
	LUT2 #(
		.INIT('h4)
	) name551 (
		_w564_,
		_w565_,
		_w566_
	);
	LUT2 #(
		.INIT('h2)
	) name552 (
		_w434_,
		_w566_,
		_w567_
	);
	LUT2 #(
		.INIT('h1)
	) name553 (
		_w563_,
		_w567_,
		_w568_
	);
	LUT2 #(
		.INIT('h4)
	) name554 (
		_w16_,
		_w133_,
		_w569_
	);
	LUT2 #(
		.INIT('h4)
	) name555 (
		_w269_,
		_w569_,
		_w570_
	);
	LUT2 #(
		.INIT('h1)
	) name556 (
		_w568_,
		_w570_,
		_w571_
	);
	LUT2 #(
		.INIT('h1)
	) name557 (
		_w37_,
		_w193_,
		_w572_
	);
	LUT2 #(
		.INIT('h2)
	) name558 (
		\v9_reg/NET0131 ,
		_w572_,
		_w573_
	);
	LUT2 #(
		.INIT('h4)
	) name559 (
		\v9_reg/NET0131 ,
		_w61_,
		_w574_
	);
	LUT2 #(
		.INIT('h8)
	) name560 (
		\v0_pad ,
		_w71_,
		_w575_
	);
	LUT2 #(
		.INIT('h1)
	) name561 (
		_w574_,
		_w575_,
		_w576_
	);
	LUT2 #(
		.INIT('h2)
	) name562 (
		\v10_reg/NET0131 ,
		\v7_reg/NET0131 ,
		_w577_
	);
	LUT2 #(
		.INIT('h4)
	) name563 (
		_w576_,
		_w577_,
		_w578_
	);
	LUT2 #(
		.INIT('h1)
	) name564 (
		_w573_,
		_w578_,
		_w579_
	);
	LUT2 #(
		.INIT('h1)
	) name565 (
		\v12_reg/NET0131 ,
		_w579_,
		_w580_
	);
	assign \_al_n0  = 1'b0;
	assign \_al_n1  = 1'b0;
	assign \g1759/_1_  = _w87_ ;
	assign \g1762/_1_  = _w147_ ;
	assign \g1764/_1_  = _w210_ ;
	assign \g1765/_0_  = _w256_ ;
	assign \g1786/_2_  = _w281_ ;
	assign \g1791/_3_  = _w297_ ;
	assign \g1808/_3_  = _w316_ ;
	assign \g1822/_2_  = _w323_ ;
	assign \g1929/_3_  = _w326_ ;
	assign \g2713/_1_  = _w358_ ;
	assign \g2744/_0_  = _w395_ ;
	assign \v13_D_11_pad  = _w406_ ;
	assign \v13_D_12_pad  = _w422_ ;
	assign \v13_D_13_pad  = _w449_ ;
	assign \v13_D_14_pad  = _w463_ ;
	assign \v13_D_16_pad  = _w468_ ;
	assign \v13_D_18_pad  = _w476_ ;
	assign \v13_D_19_pad  = _w484_ ;
	assign \v13_D_21_pad  = _w489_ ;
	assign \v13_D_22_pad  = _w497_ ;
	assign \v13_D_23_pad  = _w504_ ;
	assign \v13_D_24_pad  = _w530_ ;
	assign \v13_D_7_pad  = _w547_ ;
	assign \v13_D_8_pad  = _w571_ ;
	assign \v13_D_9_pad  = _w580_ ;
endmodule;