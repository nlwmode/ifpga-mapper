module top (\G0_pad , \G10_reg/NET0131 , \G117_pad , \G118_pad , \G11_reg/NET0131 , \G12_reg/NET0131 , \G132_pad , \G133_pad , \G13_reg/NET0131 , \G14_reg/NET0131 , \G15_reg/NET0131 , \G1_pad , \G22_reg/NET0131 , \G23_reg/NET0131 , \G2_pad , \G66_pad , \G67_pad , \_al_n0 , \_al_n1 , \g14/_0_ , \g22/_2_ , \g29/_0_ , \g37/_2_ , \g528/_2_ , \g535/_0_ , \g561/_0_ , \g572/_0_ , \g573/_0_ , \g612/_0_ , \g750/_2_ , \g757/_0_ , \g771/_0_ , \g818/_0_ );
	input \G0_pad  ;
	input \G10_reg/NET0131  ;
	input \G117_pad  ;
	input \G118_pad  ;
	input \G11_reg/NET0131  ;
	input \G12_reg/NET0131  ;
	input \G132_pad  ;
	input \G133_pad  ;
	input \G13_reg/NET0131  ;
	input \G14_reg/NET0131  ;
	input \G15_reg/NET0131  ;
	input \G1_pad  ;
	input \G22_reg/NET0131  ;
	input \G23_reg/NET0131  ;
	input \G2_pad  ;
	input \G66_pad  ;
	input \G67_pad  ;
	output \_al_n0  ;
	output \_al_n1  ;
	output \g14/_0_  ;
	output \g22/_2_  ;
	output \g29/_0_  ;
	output \g37/_2_  ;
	output \g528/_2_  ;
	output \g535/_0_  ;
	output \g561/_0_  ;
	output \g572/_0_  ;
	output \g573/_0_  ;
	output \g612/_0_  ;
	output \g750/_2_  ;
	output \g757/_0_  ;
	output \g771/_0_  ;
	output \g818/_0_  ;
	wire _w95_ ;
	wire _w94_ ;
	wire _w93_ ;
	wire _w92_ ;
	wire _w91_ ;
	wire _w90_ ;
	wire _w89_ ;
	wire _w88_ ;
	wire _w87_ ;
	wire _w86_ ;
	wire _w85_ ;
	wire _w84_ ;
	wire _w83_ ;
	wire _w82_ ;
	wire _w81_ ;
	wire _w80_ ;
	wire _w79_ ;
	wire _w78_ ;
	wire _w77_ ;
	wire _w46_ ;
	wire _w45_ ;
	wire _w44_ ;
	wire _w43_ ;
	wire _w42_ ;
	wire _w41_ ;
	wire _w40_ ;
	wire _w39_ ;
	wire _w38_ ;
	wire _w37_ ;
	wire _w36_ ;
	wire _w35_ ;
	wire _w34_ ;
	wire _w33_ ;
	wire _w32_ ;
	wire _w31_ ;
	wire _w18_ ;
	wire _w19_ ;
	wire _w20_ ;
	wire _w21_ ;
	wire _w22_ ;
	wire _w23_ ;
	wire _w24_ ;
	wire _w25_ ;
	wire _w26_ ;
	wire _w27_ ;
	wire _w28_ ;
	wire _w29_ ;
	wire _w30_ ;
	wire _w47_ ;
	wire _w48_ ;
	wire _w49_ ;
	wire _w50_ ;
	wire _w51_ ;
	wire _w52_ ;
	wire _w53_ ;
	wire _w54_ ;
	wire _w55_ ;
	wire _w56_ ;
	wire _w57_ ;
	wire _w58_ ;
	wire _w59_ ;
	wire _w60_ ;
	wire _w61_ ;
	wire _w62_ ;
	wire _w63_ ;
	wire _w64_ ;
	wire _w65_ ;
	wire _w66_ ;
	wire _w67_ ;
	wire _w68_ ;
	wire _w69_ ;
	wire _w70_ ;
	wire _w71_ ;
	wire _w72_ ;
	wire _w73_ ;
	wire _w74_ ;
	wire _w75_ ;
	wire _w76_ ;
	LUT2 #(
		.INIT('h2)
	) name0 (
		\G11_reg/NET0131 ,
		\G14_reg/NET0131 ,
		_w18_
	);
	LUT2 #(
		.INIT('h4)
	) name1 (
		\G12_reg/NET0131 ,
		\G13_reg/NET0131 ,
		_w19_
	);
	LUT2 #(
		.INIT('h4)
	) name2 (
		\G22_reg/NET0131 ,
		_w18_,
		_w20_
	);
	LUT2 #(
		.INIT('h8)
	) name3 (
		_w19_,
		_w20_,
		_w21_
	);
	LUT2 #(
		.INIT('h2)
	) name4 (
		\G15_reg/NET0131 ,
		_w21_,
		_w22_
	);
	LUT2 #(
		.INIT('h2)
	) name5 (
		\G13_reg/NET0131 ,
		\G14_reg/NET0131 ,
		_w23_
	);
	LUT2 #(
		.INIT('h1)
	) name6 (
		\G11_reg/NET0131 ,
		\G12_reg/NET0131 ,
		_w24_
	);
	LUT2 #(
		.INIT('h8)
	) name7 (
		\G22_reg/NET0131 ,
		_w23_,
		_w25_
	);
	LUT2 #(
		.INIT('h8)
	) name8 (
		_w24_,
		_w25_,
		_w26_
	);
	LUT2 #(
		.INIT('h1)
	) name9 (
		_w22_,
		_w26_,
		_w27_
	);
	LUT2 #(
		.INIT('h1)
	) name10 (
		\G0_pad ,
		_w27_,
		_w28_
	);
	LUT2 #(
		.INIT('h1)
	) name11 (
		\G10_reg/NET0131 ,
		_w27_,
		_w29_
	);
	LUT2 #(
		.INIT('h8)
	) name12 (
		\G12_reg/NET0131 ,
		\G14_reg/NET0131 ,
		_w30_
	);
	LUT2 #(
		.INIT('h8)
	) name13 (
		\G118_pad ,
		_w30_,
		_w31_
	);
	LUT2 #(
		.INIT('h8)
	) name14 (
		\G14_reg/NET0131 ,
		_w24_,
		_w32_
	);
	LUT2 #(
		.INIT('h1)
	) name15 (
		\G13_reg/NET0131 ,
		_w31_,
		_w33_
	);
	LUT2 #(
		.INIT('h4)
	) name16 (
		_w32_,
		_w33_,
		_w34_
	);
	LUT2 #(
		.INIT('h2)
	) name17 (
		_w27_,
		_w34_,
		_w35_
	);
	LUT2 #(
		.INIT('h1)
	) name18 (
		_w29_,
		_w35_,
		_w36_
	);
	LUT2 #(
		.INIT('h2)
	) name19 (
		\G14_reg/NET0131 ,
		\G15_reg/NET0131 ,
		_w37_
	);
	LUT2 #(
		.INIT('h4)
	) name20 (
		\G118_pad ,
		\G13_reg/NET0131 ,
		_w38_
	);
	LUT2 #(
		.INIT('h8)
	) name21 (
		_w37_,
		_w38_,
		_w39_
	);
	LUT2 #(
		.INIT('h1)
	) name22 (
		_w36_,
		_w39_,
		_w40_
	);
	LUT2 #(
		.INIT('h8)
	) name23 (
		\G10_reg/NET0131 ,
		_w24_,
		_w41_
	);
	LUT2 #(
		.INIT('h8)
	) name24 (
		\G13_reg/NET0131 ,
		_w41_,
		_w42_
	);
	LUT2 #(
		.INIT('h1)
	) name25 (
		\G23_reg/NET0131 ,
		_w42_,
		_w43_
	);
	LUT2 #(
		.INIT('h2)
	) name26 (
		\G14_reg/NET0131 ,
		_w43_,
		_w44_
	);
	LUT2 #(
		.INIT('h4)
	) name27 (
		\G14_reg/NET0131 ,
		_w43_,
		_w45_
	);
	LUT2 #(
		.INIT('h1)
	) name28 (
		\G0_pad ,
		_w44_,
		_w46_
	);
	LUT2 #(
		.INIT('h4)
	) name29 (
		_w45_,
		_w46_,
		_w47_
	);
	LUT2 #(
		.INIT('h1)
	) name30 (
		\G13_reg/NET0131 ,
		_w30_,
		_w48_
	);
	LUT2 #(
		.INIT('h1)
	) name31 (
		\G117_pad ,
		_w48_,
		_w49_
	);
	LUT2 #(
		.INIT('h4)
	) name32 (
		\G13_reg/NET0131 ,
		_w32_,
		_w50_
	);
	LUT2 #(
		.INIT('h1)
	) name33 (
		\G15_reg/NET0131 ,
		_w23_,
		_w51_
	);
	LUT2 #(
		.INIT('h4)
	) name34 (
		_w50_,
		_w51_,
		_w52_
	);
	LUT2 #(
		.INIT('h4)
	) name35 (
		_w49_,
		_w52_,
		_w53_
	);
	LUT2 #(
		.INIT('h2)
	) name36 (
		\G11_reg/NET0131 ,
		\G13_reg/NET0131 ,
		_w54_
	);
	LUT2 #(
		.INIT('h1)
	) name37 (
		\G14_reg/NET0131 ,
		_w54_,
		_w55_
	);
	LUT2 #(
		.INIT('h1)
	) name38 (
		\G12_reg/NET0131 ,
		\G13_reg/NET0131 ,
		_w56_
	);
	LUT2 #(
		.INIT('h4)
	) name39 (
		\G133_pad ,
		\G14_reg/NET0131 ,
		_w57_
	);
	LUT2 #(
		.INIT('h1)
	) name40 (
		_w56_,
		_w57_,
		_w58_
	);
	LUT2 #(
		.INIT('h4)
	) name41 (
		_w55_,
		_w58_,
		_w59_
	);
	LUT2 #(
		.INIT('h8)
	) name42 (
		_w27_,
		_w59_,
		_w60_
	);
	LUT2 #(
		.INIT('h2)
	) name43 (
		\G14_reg/NET0131 ,
		\G66_pad ,
		_w61_
	);
	LUT2 #(
		.INIT('h1)
	) name44 (
		_w48_,
		_w61_,
		_w62_
	);
	LUT2 #(
		.INIT('h8)
	) name45 (
		_w27_,
		_w62_,
		_w63_
	);
	LUT2 #(
		.INIT('h8)
	) name46 (
		\G10_reg/NET0131 ,
		\G11_reg/NET0131 ,
		_w64_
	);
	LUT2 #(
		.INIT('h8)
	) name47 (
		\G12_reg/NET0131 ,
		_w64_,
		_w65_
	);
	LUT2 #(
		.INIT('h1)
	) name48 (
		\G13_reg/NET0131 ,
		_w65_,
		_w66_
	);
	LUT2 #(
		.INIT('h8)
	) name49 (
		\G13_reg/NET0131 ,
		_w65_,
		_w67_
	);
	LUT2 #(
		.INIT('h1)
	) name50 (
		\G0_pad ,
		_w41_,
		_w68_
	);
	LUT2 #(
		.INIT('h4)
	) name51 (
		_w66_,
		_w68_,
		_w69_
	);
	LUT2 #(
		.INIT('h4)
	) name52 (
		_w67_,
		_w69_,
		_w70_
	);
	LUT2 #(
		.INIT('h2)
	) name53 (
		\G1_pad ,
		\G23_reg/NET0131 ,
		_w71_
	);
	LUT2 #(
		.INIT('h4)
	) name54 (
		\G1_pad ,
		\G23_reg/NET0131 ,
		_w72_
	);
	LUT2 #(
		.INIT('h1)
	) name55 (
		_w71_,
		_w72_,
		_w73_
	);
	LUT2 #(
		.INIT('h1)
	) name56 (
		\G0_pad ,
		_w73_,
		_w74_
	);
	LUT2 #(
		.INIT('h2)
	) name57 (
		\G22_reg/NET0131 ,
		\G2_pad ,
		_w75_
	);
	LUT2 #(
		.INIT('h4)
	) name58 (
		\G22_reg/NET0131 ,
		\G2_pad ,
		_w76_
	);
	LUT2 #(
		.INIT('h1)
	) name59 (
		_w75_,
		_w76_,
		_w77_
	);
	LUT2 #(
		.INIT('h1)
	) name60 (
		\G0_pad ,
		_w77_,
		_w78_
	);
	LUT2 #(
		.INIT('h1)
	) name61 (
		\G0_pad ,
		\G10_reg/NET0131 ,
		_w79_
	);
	LUT2 #(
		.INIT('h8)
	) name62 (
		\G12_reg/NET0131 ,
		_w18_,
		_w80_
	);
	LUT2 #(
		.INIT('h1)
	) name63 (
		\G67_pad ,
		_w48_,
		_w81_
	);
	LUT2 #(
		.INIT('h1)
	) name64 (
		_w80_,
		_w81_,
		_w82_
	);
	LUT2 #(
		.INIT('h8)
	) name65 (
		_w52_,
		_w82_,
		_w83_
	);
	LUT2 #(
		.INIT('h1)
	) name66 (
		\G12_reg/NET0131 ,
		_w64_,
		_w84_
	);
	LUT2 #(
		.INIT('h1)
	) name67 (
		\G0_pad ,
		_w65_,
		_w85_
	);
	LUT2 #(
		.INIT('h4)
	) name68 (
		_w84_,
		_w85_,
		_w86_
	);
	LUT2 #(
		.INIT('h2)
	) name69 (
		\G10_reg/NET0131 ,
		_w19_,
		_w87_
	);
	LUT2 #(
		.INIT('h1)
	) name70 (
		\G11_reg/NET0131 ,
		_w87_,
		_w88_
	);
	LUT2 #(
		.INIT('h1)
	) name71 (
		\G0_pad ,
		_w64_,
		_w89_
	);
	LUT2 #(
		.INIT('h4)
	) name72 (
		_w88_,
		_w89_,
		_w90_
	);
	LUT2 #(
		.INIT('h1)
	) name73 (
		\G132_pad ,
		_w56_,
		_w91_
	);
	LUT2 #(
		.INIT('h8)
	) name74 (
		\G11_reg/NET0131 ,
		_w56_,
		_w92_
	);
	LUT2 #(
		.INIT('h2)
	) name75 (
		_w37_,
		_w91_,
		_w93_
	);
	LUT2 #(
		.INIT('h4)
	) name76 (
		_w92_,
		_w93_,
		_w94_
	);
	LUT2 #(
		.INIT('h1)
	) name77 (
		_w29_,
		_w94_,
		_w95_
	);
	assign \_al_n0  = 1'b0;
	assign \_al_n1  = 1'b0;
	assign \g14/_0_  = _w28_ ;
	assign \g22/_2_  = _w40_ ;
	assign \g29/_0_  = _w47_ ;
	assign \g37/_2_  = _w53_ ;
	assign \g528/_2_  = _w60_ ;
	assign \g535/_0_  = _w63_ ;
	assign \g561/_0_  = _w70_ ;
	assign \g572/_0_  = _w74_ ;
	assign \g573/_0_  = _w78_ ;
	assign \g612/_0_  = _w79_ ;
	assign \g750/_2_  = _w83_ ;
	assign \g757/_0_  = _w86_ ;
	assign \g771/_0_  = _w90_ ;
	assign \g818/_0_  = _w95_ ;
endmodule;