module top (\G0_pad , \G10_reg/NET0131 , \G11_reg/NET0131 , \G12_reg/NET0131 , \G13_reg/NET0131 , \G147_pad , \G148_pad , \G14_reg/NET0131 , \G15_reg/NET0131 , \G16_reg/NET0131 , \G17_reg/NET0131 , \G18_reg/NET0131 , \G198_pad , \G199_pad , \G19_reg/NET0131 , \G1_pad , \G20_reg/NET0131 , \G213_pad , \G214_pad , \G21_reg/NET0131 , \G22_reg/NET0131 , \G29_reg/NET0131 , \G2_pad , \G30_reg/NET0131 , \_al_n0 , \_al_n1 , \g1001/_0_ , \g1006/_0_ , \g1008/_0_ , \g1012/_0_ , \g1020/_0_ , \g1036/_0_ , \g1056/_0_ , \g1068/_0_ , \g1070/_0_ , \g1152/_0_ , \g1298/_0_ , \g1331/_2_ , \g971/_2_ , \g973/_2_ , \g975/_2_ , \g983/_0_ , \g984/_0_ , \g985/_0_ , \g991/_2_ , \g993/_0_ , \g997/_0_ );
	input \G0_pad  ;
	input \G10_reg/NET0131  ;
	input \G11_reg/NET0131  ;
	input \G12_reg/NET0131  ;
	input \G13_reg/NET0131  ;
	input \G147_pad  ;
	input \G148_pad  ;
	input \G14_reg/NET0131  ;
	input \G15_reg/NET0131  ;
	input \G16_reg/NET0131  ;
	input \G17_reg/NET0131  ;
	input \G18_reg/NET0131  ;
	input \G198_pad  ;
	input \G199_pad  ;
	input \G19_reg/NET0131  ;
	input \G1_pad  ;
	input \G20_reg/NET0131  ;
	input \G213_pad  ;
	input \G214_pad  ;
	input \G21_reg/NET0131  ;
	input \G22_reg/NET0131  ;
	input \G29_reg/NET0131  ;
	input \G2_pad  ;
	input \G30_reg/NET0131  ;
	output \_al_n0  ;
	output \_al_n1  ;
	output \g1001/_0_  ;
	output \g1006/_0_  ;
	output \g1008/_0_  ;
	output \g1012/_0_  ;
	output \g1020/_0_  ;
	output \g1036/_0_  ;
	output \g1056/_0_  ;
	output \g1068/_0_  ;
	output \g1070/_0_  ;
	output \g1152/_0_  ;
	output \g1298/_0_  ;
	output \g1331/_2_  ;
	output \g971/_2_  ;
	output \g973/_2_  ;
	output \g975/_2_  ;
	output \g983/_0_  ;
	output \g984/_0_  ;
	output \g985/_0_  ;
	output \g991/_2_  ;
	output \g993/_0_  ;
	output \g997/_0_  ;
	wire _w150_ ;
	wire _w149_ ;
	wire _w148_ ;
	wire _w147_ ;
	wire _w146_ ;
	wire _w145_ ;
	wire _w144_ ;
	wire _w143_ ;
	wire _w142_ ;
	wire _w141_ ;
	wire _w140_ ;
	wire _w139_ ;
	wire _w138_ ;
	wire _w137_ ;
	wire _w136_ ;
	wire _w135_ ;
	wire _w134_ ;
	wire _w133_ ;
	wire _w132_ ;
	wire _w131_ ;
	wire _w130_ ;
	wire _w129_ ;
	wire _w128_ ;
	wire _w127_ ;
	wire _w126_ ;
	wire _w125_ ;
	wire _w124_ ;
	wire _w123_ ;
	wire _w122_ ;
	wire _w121_ ;
	wire _w120_ ;
	wire _w119_ ;
	wire _w118_ ;
	wire _w117_ ;
	wire _w116_ ;
	wire _w115_ ;
	wire _w114_ ;
	wire _w113_ ;
	wire _w112_ ;
	wire _w111_ ;
	wire _w110_ ;
	wire _w109_ ;
	wire _w108_ ;
	wire _w107_ ;
	wire _w106_ ;
	wire _w105_ ;
	wire _w104_ ;
	wire _w103_ ;
	wire _w102_ ;
	wire _w101_ ;
	wire _w100_ ;
	wire _w99_ ;
	wire _w98_ ;
	wire _w97_ ;
	wire _w96_ ;
	wire _w95_ ;
	wire _w94_ ;
	wire _w93_ ;
	wire _w92_ ;
	wire _w91_ ;
	wire _w90_ ;
	wire _w89_ ;
	wire _w88_ ;
	wire _w87_ ;
	wire _w86_ ;
	wire _w85_ ;
	wire _w84_ ;
	wire _w53_ ;
	wire _w52_ ;
	wire _w51_ ;
	wire _w50_ ;
	wire _w49_ ;
	wire _w48_ ;
	wire _w47_ ;
	wire _w46_ ;
	wire _w45_ ;
	wire _w44_ ;
	wire _w43_ ;
	wire _w42_ ;
	wire _w41_ ;
	wire _w40_ ;
	wire _w39_ ;
	wire _w38_ ;
	wire _w25_ ;
	wire _w26_ ;
	wire _w27_ ;
	wire _w28_ ;
	wire _w29_ ;
	wire _w30_ ;
	wire _w31_ ;
	wire _w32_ ;
	wire _w33_ ;
	wire _w34_ ;
	wire _w35_ ;
	wire _w36_ ;
	wire _w37_ ;
	wire _w54_ ;
	wire _w55_ ;
	wire _w56_ ;
	wire _w57_ ;
	wire _w58_ ;
	wire _w59_ ;
	wire _w60_ ;
	wire _w61_ ;
	wire _w62_ ;
	wire _w63_ ;
	wire _w64_ ;
	wire _w65_ ;
	wire _w66_ ;
	wire _w67_ ;
	wire _w68_ ;
	wire _w69_ ;
	wire _w70_ ;
	wire _w71_ ;
	wire _w72_ ;
	wire _w73_ ;
	wire _w74_ ;
	wire _w75_ ;
	wire _w76_ ;
	wire _w77_ ;
	wire _w78_ ;
	wire _w79_ ;
	wire _w80_ ;
	wire _w81_ ;
	wire _w82_ ;
	wire _w83_ ;
	LUT2 #(
		.INIT('h4)
	) name0 (
		\G14_reg/NET0131 ,
		\G15_reg/NET0131 ,
		_w25_
	);
	LUT2 #(
		.INIT('h2)
	) name1 (
		\G10_reg/NET0131 ,
		\G11_reg/NET0131 ,
		_w26_
	);
	LUT2 #(
		.INIT('h8)
	) name2 (
		_w25_,
		_w26_,
		_w27_
	);
	LUT2 #(
		.INIT('h1)
	) name3 (
		\G30_reg/NET0131 ,
		_w27_,
		_w28_
	);
	LUT2 #(
		.INIT('h2)
	) name4 (
		\G16_reg/NET0131 ,
		_w28_,
		_w29_
	);
	LUT2 #(
		.INIT('h8)
	) name5 (
		\G17_reg/NET0131 ,
		_w29_,
		_w30_
	);
	LUT2 #(
		.INIT('h1)
	) name6 (
		\G18_reg/NET0131 ,
		_w30_,
		_w31_
	);
	LUT2 #(
		.INIT('h8)
	) name7 (
		\G18_reg/NET0131 ,
		_w30_,
		_w32_
	);
	LUT2 #(
		.INIT('h1)
	) name8 (
		\G0_pad ,
		_w31_,
		_w33_
	);
	LUT2 #(
		.INIT('h4)
	) name9 (
		_w32_,
		_w33_,
		_w34_
	);
	LUT2 #(
		.INIT('h1)
	) name10 (
		\G17_reg/NET0131 ,
		\G18_reg/NET0131 ,
		_w35_
	);
	LUT2 #(
		.INIT('h8)
	) name11 (
		\G16_reg/NET0131 ,
		\G19_reg/NET0131 ,
		_w36_
	);
	LUT2 #(
		.INIT('h8)
	) name12 (
		_w35_,
		_w36_,
		_w37_
	);
	LUT2 #(
		.INIT('h4)
	) name13 (
		_w28_,
		_w37_,
		_w38_
	);
	LUT2 #(
		.INIT('h1)
	) name14 (
		\G20_reg/NET0131 ,
		_w38_,
		_w39_
	);
	LUT2 #(
		.INIT('h8)
	) name15 (
		\G20_reg/NET0131 ,
		_w38_,
		_w40_
	);
	LUT2 #(
		.INIT('h1)
	) name16 (
		\G0_pad ,
		_w40_,
		_w41_
	);
	LUT2 #(
		.INIT('h4)
	) name17 (
		_w39_,
		_w41_,
		_w42_
	);
	LUT2 #(
		.INIT('h2)
	) name18 (
		\G20_reg/NET0131 ,
		\G21_reg/NET0131 ,
		_w43_
	);
	LUT2 #(
		.INIT('h2)
	) name19 (
		\G12_reg/NET0131 ,
		\G13_reg/NET0131 ,
		_w44_
	);
	LUT2 #(
		.INIT('h4)
	) name20 (
		\G29_reg/NET0131 ,
		_w43_,
		_w45_
	);
	LUT2 #(
		.INIT('h8)
	) name21 (
		_w44_,
		_w45_,
		_w46_
	);
	LUT2 #(
		.INIT('h2)
	) name22 (
		\G22_reg/NET0131 ,
		_w46_,
		_w47_
	);
	LUT2 #(
		.INIT('h1)
	) name23 (
		\G20_reg/NET0131 ,
		\G21_reg/NET0131 ,
		_w48_
	);
	LUT2 #(
		.INIT('h8)
	) name24 (
		\G29_reg/NET0131 ,
		_w48_,
		_w49_
	);
	LUT2 #(
		.INIT('h8)
	) name25 (
		_w44_,
		_w49_,
		_w50_
	);
	LUT2 #(
		.INIT('h1)
	) name26 (
		_w47_,
		_w50_,
		_w51_
	);
	LUT2 #(
		.INIT('h1)
	) name27 (
		\G0_pad ,
		_w51_,
		_w52_
	);
	LUT2 #(
		.INIT('h4)
	) name28 (
		\G16_reg/NET0131 ,
		_w28_,
		_w53_
	);
	LUT2 #(
		.INIT('h1)
	) name29 (
		\G0_pad ,
		_w29_,
		_w54_
	);
	LUT2 #(
		.INIT('h4)
	) name30 (
		_w53_,
		_w54_,
		_w55_
	);
	LUT2 #(
		.INIT('h8)
	) name31 (
		\G10_reg/NET0131 ,
		\G11_reg/NET0131 ,
		_w56_
	);
	LUT2 #(
		.INIT('h8)
	) name32 (
		\G14_reg/NET0131 ,
		_w56_,
		_w57_
	);
	LUT2 #(
		.INIT('h1)
	) name33 (
		\G14_reg/NET0131 ,
		_w56_,
		_w58_
	);
	LUT2 #(
		.INIT('h1)
	) name34 (
		\G0_pad ,
		_w57_,
		_w59_
	);
	LUT2 #(
		.INIT('h4)
	) name35 (
		_w58_,
		_w59_,
		_w60_
	);
	LUT2 #(
		.INIT('h4)
	) name36 (
		\G14_reg/NET0131 ,
		_w26_,
		_w61_
	);
	LUT2 #(
		.INIT('h1)
	) name37 (
		\G15_reg/NET0131 ,
		_w57_,
		_w62_
	);
	LUT2 #(
		.INIT('h8)
	) name38 (
		\G15_reg/NET0131 ,
		_w57_,
		_w63_
	);
	LUT2 #(
		.INIT('h1)
	) name39 (
		\G0_pad ,
		_w61_,
		_w64_
	);
	LUT2 #(
		.INIT('h4)
	) name40 (
		_w62_,
		_w64_,
		_w65_
	);
	LUT2 #(
		.INIT('h4)
	) name41 (
		_w63_,
		_w65_,
		_w66_
	);
	LUT2 #(
		.INIT('h2)
	) name42 (
		\G10_reg/NET0131 ,
		_w25_,
		_w67_
	);
	LUT2 #(
		.INIT('h1)
	) name43 (
		\G11_reg/NET0131 ,
		_w67_,
		_w68_
	);
	LUT2 #(
		.INIT('h1)
	) name44 (
		\G0_pad ,
		_w56_,
		_w69_
	);
	LUT2 #(
		.INIT('h4)
	) name45 (
		_w68_,
		_w69_,
		_w70_
	);
	LUT2 #(
		.INIT('h2)
	) name46 (
		\G1_pad ,
		\G30_reg/NET0131 ,
		_w71_
	);
	LUT2 #(
		.INIT('h4)
	) name47 (
		\G1_pad ,
		\G30_reg/NET0131 ,
		_w72_
	);
	LUT2 #(
		.INIT('h1)
	) name48 (
		_w71_,
		_w72_,
		_w73_
	);
	LUT2 #(
		.INIT('h1)
	) name49 (
		\G0_pad ,
		_w73_,
		_w74_
	);
	LUT2 #(
		.INIT('h2)
	) name50 (
		\G29_reg/NET0131 ,
		\G2_pad ,
		_w75_
	);
	LUT2 #(
		.INIT('h4)
	) name51 (
		\G29_reg/NET0131 ,
		\G2_pad ,
		_w76_
	);
	LUT2 #(
		.INIT('h1)
	) name52 (
		_w75_,
		_w76_,
		_w77_
	);
	LUT2 #(
		.INIT('h1)
	) name53 (
		\G0_pad ,
		_w77_,
		_w78_
	);
	LUT2 #(
		.INIT('h1)
	) name54 (
		\G0_pad ,
		\G10_reg/NET0131 ,
		_w79_
	);
	LUT2 #(
		.INIT('h8)
	) name55 (
		\G12_reg/NET0131 ,
		\G21_reg/NET0131 ,
		_w80_
	);
	LUT2 #(
		.INIT('h1)
	) name56 (
		\G12_reg/NET0131 ,
		\G21_reg/NET0131 ,
		_w81_
	);
	LUT2 #(
		.INIT('h1)
	) name57 (
		_w80_,
		_w81_,
		_w82_
	);
	LUT2 #(
		.INIT('h2)
	) name58 (
		_w40_,
		_w82_,
		_w83_
	);
	LUT2 #(
		.INIT('h4)
	) name59 (
		\G0_pad ,
		\G13_reg/NET0131 ,
		_w84_
	);
	LUT2 #(
		.INIT('h4)
	) name60 (
		_w83_,
		_w84_,
		_w85_
	);
	LUT2 #(
		.INIT('h4)
	) name61 (
		\G0_pad ,
		\G12_reg/NET0131 ,
		_w86_
	);
	LUT2 #(
		.INIT('h4)
	) name62 (
		\G13_reg/NET0131 ,
		\G20_reg/NET0131 ,
		_w87_
	);
	LUT2 #(
		.INIT('h8)
	) name63 (
		\G21_reg/NET0131 ,
		_w87_,
		_w88_
	);
	LUT2 #(
		.INIT('h8)
	) name64 (
		_w86_,
		_w88_,
		_w89_
	);
	LUT2 #(
		.INIT('h8)
	) name65 (
		_w38_,
		_w89_,
		_w90_
	);
	LUT2 #(
		.INIT('h1)
	) name66 (
		_w85_,
		_w90_,
		_w91_
	);
	LUT2 #(
		.INIT('h1)
	) name67 (
		\G18_reg/NET0131 ,
		_w51_,
		_w92_
	);
	LUT2 #(
		.INIT('h8)
	) name68 (
		\G13_reg/NET0131 ,
		\G21_reg/NET0131 ,
		_w93_
	);
	LUT2 #(
		.INIT('h8)
	) name69 (
		\G199_pad ,
		_w93_,
		_w94_
	);
	LUT2 #(
		.INIT('h2)
	) name70 (
		\G13_reg/NET0131 ,
		\G20_reg/NET0131 ,
		_w95_
	);
	LUT2 #(
		.INIT('h4)
	) name71 (
		\G21_reg/NET0131 ,
		_w95_,
		_w96_
	);
	LUT2 #(
		.INIT('h1)
	) name72 (
		\G12_reg/NET0131 ,
		_w94_,
		_w97_
	);
	LUT2 #(
		.INIT('h4)
	) name73 (
		_w96_,
		_w97_,
		_w98_
	);
	LUT2 #(
		.INIT('h2)
	) name74 (
		_w51_,
		_w98_,
		_w99_
	);
	LUT2 #(
		.INIT('h1)
	) name75 (
		_w92_,
		_w99_,
		_w100_
	);
	LUT2 #(
		.INIT('h2)
	) name76 (
		\G13_reg/NET0131 ,
		\G22_reg/NET0131 ,
		_w101_
	);
	LUT2 #(
		.INIT('h2)
	) name77 (
		\G12_reg/NET0131 ,
		\G199_pad ,
		_w102_
	);
	LUT2 #(
		.INIT('h8)
	) name78 (
		_w101_,
		_w102_,
		_w103_
	);
	LUT2 #(
		.INIT('h1)
	) name79 (
		_w100_,
		_w103_,
		_w104_
	);
	LUT2 #(
		.INIT('h1)
	) name80 (
		\G12_reg/NET0131 ,
		_w93_,
		_w105_
	);
	LUT2 #(
		.INIT('h1)
	) name81 (
		\G148_pad ,
		_w105_,
		_w106_
	);
	LUT2 #(
		.INIT('h8)
	) name82 (
		_w81_,
		_w95_,
		_w107_
	);
	LUT2 #(
		.INIT('h1)
	) name83 (
		_w44_,
		_w107_,
		_w108_
	);
	LUT2 #(
		.INIT('h1)
	) name84 (
		_w88_,
		_w106_,
		_w109_
	);
	LUT2 #(
		.INIT('h8)
	) name85 (
		_w108_,
		_w109_,
		_w110_
	);
	LUT2 #(
		.INIT('h8)
	) name86 (
		_w51_,
		_w110_,
		_w111_
	);
	LUT2 #(
		.INIT('h1)
	) name87 (
		\G198_pad ,
		_w105_,
		_w112_
	);
	LUT2 #(
		.INIT('h2)
	) name88 (
		_w108_,
		_w112_,
		_w113_
	);
	LUT2 #(
		.INIT('h8)
	) name89 (
		_w51_,
		_w113_,
		_w114_
	);
	LUT2 #(
		.INIT('h8)
	) name90 (
		\G13_reg/NET0131 ,
		\G214_pad ,
		_w115_
	);
	LUT2 #(
		.INIT('h1)
	) name91 (
		_w87_,
		_w115_,
		_w116_
	);
	LUT2 #(
		.INIT('h1)
	) name92 (
		_w44_,
		_w81_,
		_w117_
	);
	LUT2 #(
		.INIT('h4)
	) name93 (
		_w116_,
		_w117_,
		_w118_
	);
	LUT2 #(
		.INIT('h8)
	) name94 (
		_w51_,
		_w118_,
		_w119_
	);
	LUT2 #(
		.INIT('h8)
	) name95 (
		\G21_reg/NET0131 ,
		_w41_,
		_w120_
	);
	LUT2 #(
		.INIT('h4)
	) name96 (
		\G12_reg/NET0131 ,
		\G13_reg/NET0131 ,
		_w121_
	);
	LUT2 #(
		.INIT('h4)
	) name97 (
		\G0_pad ,
		_w43_,
		_w122_
	);
	LUT2 #(
		.INIT('h4)
	) name98 (
		_w121_,
		_w122_,
		_w123_
	);
	LUT2 #(
		.INIT('h8)
	) name99 (
		_w38_,
		_w123_,
		_w124_
	);
	LUT2 #(
		.INIT('h1)
	) name100 (
		_w120_,
		_w124_,
		_w125_
	);
	LUT2 #(
		.INIT('h1)
	) name101 (
		\G213_pad ,
		_w81_,
		_w126_
	);
	LUT2 #(
		.INIT('h4)
	) name102 (
		\G12_reg/NET0131 ,
		_w43_,
		_w127_
	);
	LUT2 #(
		.INIT('h2)
	) name103 (
		_w101_,
		_w126_,
		_w128_
	);
	LUT2 #(
		.INIT('h4)
	) name104 (
		_w127_,
		_w128_,
		_w129_
	);
	LUT2 #(
		.INIT('h1)
	) name105 (
		_w92_,
		_w129_,
		_w130_
	);
	LUT2 #(
		.INIT('h8)
	) name106 (
		\G21_reg/NET0131 ,
		_w40_,
		_w131_
	);
	LUT2 #(
		.INIT('h2)
	) name107 (
		_w86_,
		_w131_,
		_w132_
	);
	LUT2 #(
		.INIT('h1)
	) name108 (
		\G0_pad ,
		\G12_reg/NET0131 ,
		_w133_
	);
	LUT2 #(
		.INIT('h8)
	) name109 (
		_w131_,
		_w133_,
		_w134_
	);
	LUT2 #(
		.INIT('h1)
	) name110 (
		_w132_,
		_w134_,
		_w135_
	);
	LUT2 #(
		.INIT('h1)
	) name111 (
		\G19_reg/NET0131 ,
		_w32_,
		_w136_
	);
	LUT2 #(
		.INIT('h8)
	) name112 (
		\G17_reg/NET0131 ,
		\G18_reg/NET0131 ,
		_w137_
	);
	LUT2 #(
		.INIT('h8)
	) name113 (
		\G19_reg/NET0131 ,
		_w137_,
		_w138_
	);
	LUT2 #(
		.INIT('h1)
	) name114 (
		_w35_,
		_w138_,
		_w139_
	);
	LUT2 #(
		.INIT('h2)
	) name115 (
		_w29_,
		_w139_,
		_w140_
	);
	LUT2 #(
		.INIT('h1)
	) name116 (
		\G0_pad ,
		_w140_,
		_w141_
	);
	LUT2 #(
		.INIT('h4)
	) name117 (
		_w136_,
		_w141_,
		_w142_
	);
	LUT2 #(
		.INIT('h2)
	) name118 (
		\G13_reg/NET0131 ,
		\G147_pad ,
		_w143_
	);
	LUT2 #(
		.INIT('h1)
	) name119 (
		_w105_,
		_w143_,
		_w144_
	);
	LUT2 #(
		.INIT('h8)
	) name120 (
		_w51_,
		_w144_,
		_w145_
	);
	LUT2 #(
		.INIT('h4)
	) name121 (
		\G18_reg/NET0131 ,
		\G19_reg/NET0131 ,
		_w146_
	);
	LUT2 #(
		.INIT('h2)
	) name122 (
		_w29_,
		_w146_,
		_w147_
	);
	LUT2 #(
		.INIT('h1)
	) name123 (
		\G17_reg/NET0131 ,
		_w147_,
		_w148_
	);
	LUT2 #(
		.INIT('h1)
	) name124 (
		\G0_pad ,
		_w30_,
		_w149_
	);
	LUT2 #(
		.INIT('h4)
	) name125 (
		_w148_,
		_w149_,
		_w150_
	);
	assign \_al_n0  = 1'b0;
	assign \_al_n1  = 1'b0;
	assign \g1001/_0_  = _w34_ ;
	assign \g1006/_0_  = _w42_ ;
	assign \g1008/_0_  = _w52_ ;
	assign \g1012/_0_  = _w55_ ;
	assign \g1020/_0_  = _w60_ ;
	assign \g1036/_0_  = _w66_ ;
	assign \g1056/_0_  = _w70_ ;
	assign \g1068/_0_  = _w74_ ;
	assign \g1070/_0_  = _w78_ ;
	assign \g1152/_0_  = _w79_ ;
	assign \g1298/_0_  = _w91_ ;
	assign \g1331/_2_  = _w104_ ;
	assign \g971/_2_  = _w111_ ;
	assign \g973/_2_  = _w114_ ;
	assign \g975/_2_  = _w119_ ;
	assign \g983/_0_  = _w125_ ;
	assign \g984/_0_  = _w130_ ;
	assign \g985/_0_  = _w135_ ;
	assign \g991/_2_  = _w142_ ;
	assign \g993/_0_  = _w145_ ;
	assign \g997/_0_  = _w150_ ;
endmodule;