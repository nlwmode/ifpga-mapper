module top( \a0_pad  , \a1_pad  , \a2_pad  , a_pad , \b0_pad  , \b1_pad  , \b2_pad  , b_pad , \c0_pad  , \c1_pad  , \c2_pad  , \d0_pad  , \d1_pad  , \d2_pad  , \e0_pad  , \e1_pad  , \e2_pad  , \f0_pad  , \f1_pad  , \f2_pad  , \g0_pad  , \g1_pad  , \g2_pad  , g_pad , \h0_pad  , \h1_pad  , \h2_pad  , h_pad , \i0_pad  , \i1_pad  , \i2_pad  , i_pad , \j1_pad  , \j2_pad  , \k0_pad  , \k1_pad  , \k2_pad  , k_pad , \l0_pad  , \l1_pad  , \l2_pad  , l_pad , \m0_pad  , \m1_pad  , \m2_pad  , m_pad , \n0_pad  , \n1_pad  , \n2_pad  , n_pad , \o0_pad  , \o1_pad  , \o2_pad  , o_pad , \p0_pad  , \p1_pad  , \p2_pad  , p_pad , \q0_pad  , \q1_pad  , \q2_pad  , q_pad , \r0_pad  , \r1_pad  , \r2_pad  , r_pad , \s0_pad  , \s1_pad  , \s2_pad  , s_pad , \t0_pad  , \t1_pad  , \t2_pad  , t_pad , \u0_pad  , \u1_pad  , \u2_pad  , u_pad , \v0_pad  , \v1_pad  , \v2_pad  , v_pad , \w0_pad  , \w1_pad  , w_pad , \x0_pad  , \x1_pad  , x_pad , \y0_pad  , \y1_pad  , y_pad , \z0_pad  , \z1_pad  , z_pad , \a3_pad  , \a4_pad  , \a5_pad  , \b3_pad  , \b4_pad  , \b5_pad  , \c3_pad  , \c4_pad  , \c5_pad  , \d3_pad  , \d4_pad  , \d5_pad  , \e3_pad  , \e4_pad  , \e5_pad  , \f3_pad  , \f4_pad  , \f5_pad  , \g3_pad  , \g4_pad  , \g5_pad  , \h3_pad  , \h4_pad  , \h5_pad  , \i3_pad  , \i4_pad  , \i5_pad  , \j3_pad  , \j4_pad  , \j5_pad  , \k3_pad  , \k4_pad  , \k5_pad  , \l3_pad  , \l4_pad  , \l5_pad  , \m3_pad  , \m4_pad  , \m5_pad  , \n3_pad  , \n4_pad  , \n5_pad  , \o3_pad  , \o4_pad  , \o5_pad  , \p3_pad  , \p4_pad  , \q3_pad  , \q4_pad  , \r3_pad  , \r4_pad  , \s3_pad  , \s4_pad  , \t3_pad  , \t4_pad  , \u3_pad  , \u4_pad  , \v3_pad  , \v4_pad  , \w2_pad  , \w3_pad  , \w4_pad  , \x2_pad  , \x3_pad  , \x4_pad  , \y2_pad  , \y3_pad  , \y4_pad  , \z2_pad  , \z3_pad  , \z4_pad  );
  input \a0_pad  ;
  input \a1_pad  ;
  input \a2_pad  ;
  input a_pad ;
  input \b0_pad  ;
  input \b1_pad  ;
  input \b2_pad  ;
  input b_pad ;
  input \c0_pad  ;
  input \c1_pad  ;
  input \c2_pad  ;
  input \d0_pad  ;
  input \d1_pad  ;
  input \d2_pad  ;
  input \e0_pad  ;
  input \e1_pad  ;
  input \e2_pad  ;
  input \f0_pad  ;
  input \f1_pad  ;
  input \f2_pad  ;
  input \g0_pad  ;
  input \g1_pad  ;
  input \g2_pad  ;
  input g_pad ;
  input \h0_pad  ;
  input \h1_pad  ;
  input \h2_pad  ;
  input h_pad ;
  input \i0_pad  ;
  input \i1_pad  ;
  input \i2_pad  ;
  input i_pad ;
  input \j1_pad  ;
  input \j2_pad  ;
  input \k0_pad  ;
  input \k1_pad  ;
  input \k2_pad  ;
  input k_pad ;
  input \l0_pad  ;
  input \l1_pad  ;
  input \l2_pad  ;
  input l_pad ;
  input \m0_pad  ;
  input \m1_pad  ;
  input \m2_pad  ;
  input m_pad ;
  input \n0_pad  ;
  input \n1_pad  ;
  input \n2_pad  ;
  input n_pad ;
  input \o0_pad  ;
  input \o1_pad  ;
  input \o2_pad  ;
  input o_pad ;
  input \p0_pad  ;
  input \p1_pad  ;
  input \p2_pad  ;
  input p_pad ;
  input \q0_pad  ;
  input \q1_pad  ;
  input \q2_pad  ;
  input q_pad ;
  input \r0_pad  ;
  input \r1_pad  ;
  input \r2_pad  ;
  input r_pad ;
  input \s0_pad  ;
  input \s1_pad  ;
  input \s2_pad  ;
  input s_pad ;
  input \t0_pad  ;
  input \t1_pad  ;
  input \t2_pad  ;
  input t_pad ;
  input \u0_pad  ;
  input \u1_pad  ;
  input \u2_pad  ;
  input u_pad ;
  input \v0_pad  ;
  input \v1_pad  ;
  input \v2_pad  ;
  input v_pad ;
  input \w0_pad  ;
  input \w1_pad  ;
  input w_pad ;
  input \x0_pad  ;
  input \x1_pad  ;
  input x_pad ;
  input \y0_pad  ;
  input \y1_pad  ;
  input y_pad ;
  input \z0_pad  ;
  input \z1_pad  ;
  input z_pad ;
  output \a3_pad  ;
  output \a4_pad  ;
  output \a5_pad  ;
  output \b3_pad  ;
  output \b4_pad  ;
  output \b5_pad  ;
  output \c3_pad  ;
  output \c4_pad  ;
  output \c5_pad  ;
  output \d3_pad  ;
  output \d4_pad  ;
  output \d5_pad  ;
  output \e3_pad  ;
  output \e4_pad  ;
  output \e5_pad  ;
  output \f3_pad  ;
  output \f4_pad  ;
  output \f5_pad  ;
  output \g3_pad  ;
  output \g4_pad  ;
  output \g5_pad  ;
  output \h3_pad  ;
  output \h4_pad  ;
  output \h5_pad  ;
  output \i3_pad  ;
  output \i4_pad  ;
  output \i5_pad  ;
  output \j3_pad  ;
  output \j4_pad  ;
  output \j5_pad  ;
  output \k3_pad  ;
  output \k4_pad  ;
  output \k5_pad  ;
  output \l3_pad  ;
  output \l4_pad  ;
  output \l5_pad  ;
  output \m3_pad  ;
  output \m4_pad  ;
  output \m5_pad  ;
  output \n3_pad  ;
  output \n4_pad  ;
  output \n5_pad  ;
  output \o3_pad  ;
  output \o4_pad  ;
  output \o5_pad  ;
  output \p3_pad  ;
  output \p4_pad  ;
  output \q3_pad  ;
  output \q4_pad  ;
  output \r3_pad  ;
  output \r4_pad  ;
  output \s3_pad  ;
  output \s4_pad  ;
  output \t3_pad  ;
  output \t4_pad  ;
  output \u3_pad  ;
  output \u4_pad  ;
  output \v3_pad  ;
  output \v4_pad  ;
  output \w2_pad  ;
  output \w3_pad  ;
  output \w4_pad  ;
  output \x2_pad  ;
  output \x3_pad  ;
  output \x4_pad  ;
  output \y2_pad  ;
  output \y3_pad  ;
  output \y4_pad  ;
  output \z2_pad  ;
  output \z3_pad  ;
  output \z4_pad  ;
  wire n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 ;
  assign n95 = ~\p2_pad  & ~\q2_pad  ;
  assign n96 = ~\r2_pad  & n95 ;
  assign n97 = \e1_pad  & ~\n2_pad  ;
  assign n98 = \o2_pad  & n97 ;
  assign n99 = n96 & n98 ;
  assign n100 = ~\h1_pad  & ~n99 ;
  assign n101 = ~\q0_pad  & ~\r2_pad  ;
  assign n102 = n95 & n101 ;
  assign n103 = n98 & n102 ;
  assign n104 = ~\c1_pad  & ~n103 ;
  assign n105 = ~n100 & n104 ;
  assign n106 = ~g_pad & ~h_pad ;
  assign n107 = \h0_pad  & ~i_pad ;
  assign n108 = n106 & n107 ;
  assign n109 = \g0_pad  & \v2_pad  ;
  assign n110 = \c0_pad  & \m1_pad  ;
  assign n111 = n109 & n110 ;
  assign n112 = ~n108 & n111 ;
  assign n113 = \m1_pad  & n109 ;
  assign n114 = ~n108 & n113 ;
  assign n115 = \e1_pad  & ~\m0_pad  ;
  assign n116 = ~\h2_pad  & ~n115 ;
  assign n117 = ~\i2_pad  & n115 ;
  assign n118 = ~n116 & ~n117 ;
  assign n119 = ~n114 & n118 ;
  assign n120 = ~n112 & ~n119 ;
  assign n121 = ~\i0_pad  & ~n120 ;
  assign n122 = ~\i1_pad  & ~n99 ;
  assign n123 = ~\r0_pad  & ~\r2_pad  ;
  assign n124 = n95 & n123 ;
  assign n125 = n98 & n124 ;
  assign n126 = ~\c1_pad  & ~n125 ;
  assign n127 = ~n122 & n126 ;
  assign n128 = \d0_pad  & \m1_pad  ;
  assign n129 = n109 & n128 ;
  assign n130 = ~n108 & n129 ;
  assign n131 = ~\i2_pad  & ~n115 ;
  assign n132 = ~\j2_pad  & n115 ;
  assign n133 = ~n131 & ~n132 ;
  assign n134 = ~n114 & n133 ;
  assign n135 = ~n130 & ~n134 ;
  assign n136 = ~\i0_pad  & ~n135 ;
  assign n137 = \e1_pad  & \n2_pad  ;
  assign n138 = ~\o2_pad  & n137 ;
  assign n139 = ~i_pad & ~\q2_pad  ;
  assign n140 = ~\p2_pad  & \r2_pad  ;
  assign n141 = ~n139 & n140 ;
  assign n142 = n138 & n141 ;
  assign n143 = \h0_pad  & ~\t2_pad  ;
  assign n144 = ~\h0_pad  & \t2_pad  ;
  assign n145 = ~n143 & ~n144 ;
  assign n146 = ~\i0_pad  & n145 ;
  assign n147 = n142 & n146 ;
  assign n148 = ~\i0_pad  & \s2_pad  ;
  assign n149 = ~n142 & n148 ;
  assign n150 = ~n147 & ~n149 ;
  assign n151 = ~\j1_pad  & ~n99 ;
  assign n152 = ~\r2_pad  & ~\s0_pad  ;
  assign n153 = n95 & n152 ;
  assign n154 = n98 & n153 ;
  assign n155 = ~\c1_pad  & ~n154 ;
  assign n156 = ~n151 & n155 ;
  assign n157 = ~\i0_pad  & \m1_pad  ;
  assign n158 = n109 & n157 ;
  assign n159 = ~n108 & n158 ;
  assign n160 = \e0_pad  & n159 ;
  assign n161 = \j2_pad  & ~n115 ;
  assign n162 = ~\i0_pad  & n161 ;
  assign n163 = ~n114 & n162 ;
  assign n164 = ~n160 & ~n163 ;
  assign n165 = \f0_pad  & \v2_pad  ;
  assign n166 = ~\k0_pad  & ~n165 ;
  assign n167 = ~\c1_pad  & ~n166 ;
  assign n168 = \m1_pad  & ~n108 ;
  assign n169 = ~\c1_pad  & n109 ;
  assign n170 = ~n168 & n169 ;
  assign n171 = ~n167 & ~n170 ;
  assign n172 = ~\k1_pad  & ~n99 ;
  assign n173 = ~\r2_pad  & ~\t0_pad  ;
  assign n174 = n95 & n173 ;
  assign n175 = n98 & n174 ;
  assign n176 = ~\c1_pad  & ~n175 ;
  assign n177 = ~n172 & n176 ;
  assign n178 = b_pad & ~\u0_pad  ;
  assign n179 = ~\k2_pad  & ~\u2_pad  ;
  assign n180 = ~n178 & n179 ;
  assign n181 = ~\c1_pad  & ~\k2_pad  ;
  assign n182 = ~\c1_pad  & ~\u2_pad  ;
  assign n183 = ~n178 & n182 ;
  assign n184 = ~n181 & ~n183 ;
  assign n185 = ~n180 & ~n184 ;
  assign n186 = n96 & n138 ;
  assign n187 = ~\l0_pad  & ~n186 ;
  assign n188 = ~\c1_pad  & ~n187 ;
  assign n189 = ~\l1_pad  & ~n186 ;
  assign n190 = ~\c1_pad  & ~n189 ;
  assign n191 = ~\u2_pad  & ~n178 ;
  assign n192 = \k2_pad  & \l2_pad  ;
  assign n193 = ~n191 & n192 ;
  assign n194 = ~\k2_pad  & \m2_pad  ;
  assign n195 = \l2_pad  & ~n194 ;
  assign n196 = ~\c1_pad  & n195 ;
  assign n197 = ~\c1_pad  & \k2_pad  ;
  assign n198 = ~n191 & n197 ;
  assign n199 = ~n196 & ~n198 ;
  assign n200 = ~n193 & ~n199 ;
  assign n201 = ~\i0_pad  & ~n109 ;
  assign n202 = ~n108 & n157 ;
  assign n203 = ~n201 & ~n202 ;
  assign n204 = \m0_pad  & ~n109 ;
  assign n205 = ~n203 & ~n204 ;
  assign n206 = ~\k2_pad  & \l2_pad  ;
  assign n207 = \m2_pad  & n206 ;
  assign n208 = n106 & n207 ;
  assign n209 = ~\m1_pad  & ~n208 ;
  assign n210 = n201 & ~n209 ;
  assign n211 = ~\l2_pad  & ~\m2_pad  ;
  assign n212 = ~\m2_pad  & ~\u2_pad  ;
  assign n213 = ~n178 & n212 ;
  assign n214 = ~n211 & ~n213 ;
  assign n215 = \l2_pad  & \m2_pad  ;
  assign n216 = ~n191 & n215 ;
  assign n217 = ~\c1_pad  & ~n206 ;
  assign n218 = ~n216 & n217 ;
  assign n219 = n214 & n218 ;
  assign n220 = ~\n0_pad  & ~n186 ;
  assign n221 = ~\c1_pad  & ~\i0_pad  ;
  assign n222 = ~n220 & n221 ;
  assign n223 = i_pad & \m1_pad  ;
  assign n224 = n109 & n223 ;
  assign n225 = \h0_pad  & n106 ;
  assign n226 = n113 & ~n225 ;
  assign n227 = ~\n1_pad  & ~n115 ;
  assign n228 = \o1_pad  & n115 ;
  assign n229 = ~n227 & ~n228 ;
  assign n230 = ~n226 & n229 ;
  assign n231 = ~n224 & ~n230 ;
  assign n232 = ~\i0_pad  & ~n231 ;
  assign n233 = ~\d1_pad  & ~\e1_pad  ;
  assign n234 = ~\n2_pad  & n233 ;
  assign n235 = ~n207 & n234 ;
  assign n236 = \n2_pad  & ~n233 ;
  assign n237 = \m2_pad  & \n2_pad  ;
  assign n238 = n206 & n237 ;
  assign n239 = ~n236 & ~n238 ;
  assign n240 = ~\c1_pad  & n239 ;
  assign n241 = ~n235 & n240 ;
  assign n242 = \o0_pad  & n221 ;
  assign n243 = ~\i0_pad  & ~n114 ;
  assign n244 = ~\p1_pad  & n115 ;
  assign n245 = \o1_pad  & ~n115 ;
  assign n246 = ~n244 & ~n245 ;
  assign n247 = n243 & n246 ;
  assign n248 = ~\c1_pad  & \o2_pad  ;
  assign n249 = n239 & n248 ;
  assign n250 = ~\c1_pad  & ~\o2_pad  ;
  assign n251 = ~n239 & n250 ;
  assign n252 = ~n249 & ~n251 ;
  assign n253 = \p0_pad  & n221 ;
  assign n254 = k_pad & n159 ;
  assign n255 = ~\p1_pad  & ~n115 ;
  assign n256 = ~\q1_pad  & n115 ;
  assign n257 = ~n255 & ~n256 ;
  assign n258 = n243 & n257 ;
  assign n259 = ~n254 & ~n258 ;
  assign n260 = \o2_pad  & ~n239 ;
  assign n261 = ~\p2_pad  & ~n260 ;
  assign n262 = \o2_pad  & \p2_pad  ;
  assign n263 = ~n239 & n262 ;
  assign n264 = ~\c1_pad  & ~n263 ;
  assign n265 = ~n261 & n264 ;
  assign n266 = \q0_pad  & n221 ;
  assign n267 = l_pad & \m1_pad  ;
  assign n268 = n109 & n267 ;
  assign n269 = ~n108 & n268 ;
  assign n270 = ~\q1_pad  & ~n115 ;
  assign n271 = ~\r1_pad  & n115 ;
  assign n272 = ~n270 & ~n271 ;
  assign n273 = ~n114 & n272 ;
  assign n274 = ~n269 & ~n273 ;
  assign n275 = ~\i0_pad  & ~n274 ;
  assign n276 = ~\q2_pad  & ~n263 ;
  assign n277 = \o2_pad  & \q2_pad  ;
  assign n278 = \p2_pad  & n277 ;
  assign n279 = ~n239 & n278 ;
  assign n280 = ~\c1_pad  & ~n279 ;
  assign n281 = ~n276 & n280 ;
  assign n282 = \r0_pad  & n221 ;
  assign n283 = \m1_pad  & m_pad ;
  assign n284 = n109 & n283 ;
  assign n285 = ~n108 & n284 ;
  assign n286 = ~\r1_pad  & ~n115 ;
  assign n287 = ~\s1_pad  & n115 ;
  assign n288 = ~n286 & ~n287 ;
  assign n289 = ~n114 & n288 ;
  assign n290 = ~n285 & ~n289 ;
  assign n291 = ~\i0_pad  & ~n290 ;
  assign n292 = ~\c1_pad  & \r2_pad  ;
  assign n293 = ~n279 & n292 ;
  assign n294 = ~\c1_pad  & ~\r2_pad  ;
  assign n295 = n279 & n294 ;
  assign n296 = ~n293 & ~n295 ;
  assign n297 = \s0_pad  & n221 ;
  assign n298 = \m1_pad  & n_pad ;
  assign n299 = n109 & n298 ;
  assign n300 = ~n108 & n299 ;
  assign n301 = ~\s1_pad  & ~n115 ;
  assign n302 = ~\t1_pad  & n115 ;
  assign n303 = ~n301 & ~n302 ;
  assign n304 = ~n114 & n303 ;
  assign n305 = ~n300 & ~n304 ;
  assign n306 = ~\i0_pad  & ~n305 ;
  assign n307 = \b1_pad  & ~\i0_pad  ;
  assign n308 = ~n115 & n307 ;
  assign n309 = ~\i0_pad  & \n1_pad  ;
  assign n310 = n115 & n309 ;
  assign n311 = ~n308 & ~n310 ;
  assign n312 = \t0_pad  & n221 ;
  assign n313 = \m1_pad  & o_pad ;
  assign n314 = n109 & n313 ;
  assign n315 = ~n108 & n314 ;
  assign n316 = ~\t1_pad  & ~n115 ;
  assign n317 = ~\u1_pad  & n115 ;
  assign n318 = ~n316 & ~n317 ;
  assign n319 = ~n114 & n318 ;
  assign n320 = ~n315 & ~n319 ;
  assign n321 = ~\i0_pad  & ~n320 ;
  assign n322 = \l1_pad  & \s2_pad  ;
  assign n323 = ~\c1_pad  & \t2_pad  ;
  assign n324 = ~n322 & n323 ;
  assign n325 = ~\c1_pad  & ~\t2_pad  ;
  assign n326 = n322 & n325 ;
  assign n327 = ~n324 & ~n326 ;
  assign n328 = b_pad & ~\i0_pad  ;
  assign n329 = \m1_pad  & p_pad ;
  assign n330 = n109 & n329 ;
  assign n331 = ~n108 & n330 ;
  assign n332 = ~\u1_pad  & ~n115 ;
  assign n333 = ~\v1_pad  & n115 ;
  assign n334 = ~n332 & ~n333 ;
  assign n335 = ~n114 & n334 ;
  assign n336 = ~n331 & ~n335 ;
  assign n337 = ~\i0_pad  & ~n336 ;
  assign n338 = ~n178 & n207 ;
  assign n339 = ~\i0_pad  & ~n191 ;
  assign n340 = ~n338 & n339 ;
  assign n341 = a_pad & ~\i0_pad  ;
  assign n342 = \m1_pad  & q_pad ;
  assign n343 = n109 & n342 ;
  assign n344 = ~n108 & n343 ;
  assign n345 = ~\v1_pad  & ~n115 ;
  assign n346 = ~\w1_pad  & n115 ;
  assign n347 = ~n345 & ~n346 ;
  assign n348 = ~n114 & n347 ;
  assign n349 = ~n344 & ~n348 ;
  assign n350 = ~\i0_pad  & ~n349 ;
  assign n351 = ~\f0_pad  & \v2_pad  ;
  assign n352 = ~n142 & ~n351 ;
  assign n353 = n201 & ~n352 ;
  assign n354 = ~\i0_pad  & \v0_pad  ;
  assign n355 = \m1_pad  & r_pad ;
  assign n356 = n109 & n355 ;
  assign n357 = ~n108 & n356 ;
  assign n358 = ~\w1_pad  & ~n115 ;
  assign n359 = ~\x1_pad  & n115 ;
  assign n360 = ~n358 & ~n359 ;
  assign n361 = ~n114 & n360 ;
  assign n362 = ~n357 & ~n361 ;
  assign n363 = ~\i0_pad  & ~n362 ;
  assign n364 = ~\i0_pad  & \w0_pad  ;
  assign n365 = \m1_pad  & s_pad ;
  assign n366 = n109 & n365 ;
  assign n367 = ~n108 & n366 ;
  assign n368 = ~\x1_pad  & ~n115 ;
  assign n369 = ~\y1_pad  & n115 ;
  assign n370 = ~n368 & ~n369 ;
  assign n371 = ~n114 & n370 ;
  assign n372 = ~n367 & ~n371 ;
  assign n373 = ~\i0_pad  & ~n372 ;
  assign n374 = ~\i0_pad  & \x0_pad  ;
  assign n375 = \m1_pad  & t_pad ;
  assign n376 = n109 & n375 ;
  assign n377 = ~n108 & n376 ;
  assign n378 = ~\y1_pad  & ~n115 ;
  assign n379 = ~\z1_pad  & n115 ;
  assign n380 = ~n378 & ~n379 ;
  assign n381 = ~n114 & n380 ;
  assign n382 = ~n377 & ~n381 ;
  assign n383 = ~\i0_pad  & ~n382 ;
  assign n384 = ~\i0_pad  & \y0_pad  ;
  assign n385 = \m1_pad  & u_pad ;
  assign n386 = n109 & n385 ;
  assign n387 = ~n108 & n386 ;
  assign n388 = ~\z1_pad  & ~n115 ;
  assign n389 = ~\a2_pad  & n115 ;
  assign n390 = ~n388 & ~n389 ;
  assign n391 = ~n114 & n390 ;
  assign n392 = ~n387 & ~n391 ;
  assign n393 = ~\i0_pad  & ~n392 ;
  assign n394 = ~\i0_pad  & \z0_pad  ;
  assign n395 = \m1_pad  & v_pad ;
  assign n396 = n109 & n395 ;
  assign n397 = ~n108 & n396 ;
  assign n398 = ~\a2_pad  & ~n115 ;
  assign n399 = ~\b2_pad  & n115 ;
  assign n400 = ~n398 & ~n399 ;
  assign n401 = ~n114 & n400 ;
  assign n402 = ~n397 & ~n401 ;
  assign n403 = ~\i0_pad  & ~n402 ;
  assign n404 = \a1_pad  & ~\i0_pad  ;
  assign n405 = \m1_pad  & w_pad ;
  assign n406 = n109 & n405 ;
  assign n407 = ~n108 & n406 ;
  assign n408 = ~\b2_pad  & ~n115 ;
  assign n409 = ~\c2_pad  & n115 ;
  assign n410 = ~n408 & ~n409 ;
  assign n411 = ~n114 & n410 ;
  assign n412 = ~n407 & ~n411 ;
  assign n413 = ~\i0_pad  & ~n412 ;
  assign n414 = ~n142 & ~n165 ;
  assign n415 = ~n203 & n414 ;
  assign n416 = \m1_pad  & x_pad ;
  assign n417 = n109 & n416 ;
  assign n418 = ~n108 & n417 ;
  assign n419 = ~\c2_pad  & ~n115 ;
  assign n420 = ~\d2_pad  & n115 ;
  assign n421 = ~n419 & ~n420 ;
  assign n422 = ~n114 & n421 ;
  assign n423 = ~n418 & ~n422 ;
  assign n424 = ~\i0_pad  & ~n423 ;
  assign n425 = ~\g0_pad  & \i0_pad  ;
  assign n426 = ~\m1_pad  & \v2_pad  ;
  assign n427 = n425 & n426 ;
  assign n428 = ~n108 & n427 ;
  assign n429 = \m1_pad  & y_pad ;
  assign n430 = n109 & n429 ;
  assign n431 = ~n108 & n430 ;
  assign n432 = ~\d2_pad  & ~n115 ;
  assign n433 = ~\e2_pad  & n115 ;
  assign n434 = ~n432 & ~n433 ;
  assign n435 = ~n114 & n434 ;
  assign n436 = ~n431 & ~n435 ;
  assign n437 = ~\i0_pad  & ~n436 ;
  assign n438 = ~\c1_pad  & ~n233 ;
  assign n439 = ~\c1_pad  & \m2_pad  ;
  assign n440 = n206 & n439 ;
  assign n441 = ~n438 & ~n440 ;
  assign n442 = \m1_pad  & z_pad ;
  assign n443 = n109 & n442 ;
  assign n444 = ~n108 & n443 ;
  assign n445 = ~\e2_pad  & ~n115 ;
  assign n446 = ~\f2_pad  & n115 ;
  assign n447 = ~n445 & ~n446 ;
  assign n448 = ~n114 & n447 ;
  assign n449 = ~n444 & ~n448 ;
  assign n450 = ~\i0_pad  & ~n449 ;
  assign n451 = ~\f1_pad  & ~n99 ;
  assign n452 = ~\o0_pad  & ~\r2_pad  ;
  assign n453 = n95 & n452 ;
  assign n454 = n98 & n453 ;
  assign n455 = ~\c1_pad  & ~n454 ;
  assign n456 = ~n451 & n455 ;
  assign n457 = \a0_pad  & \m1_pad  ;
  assign n458 = n109 & n457 ;
  assign n459 = ~n108 & n458 ;
  assign n460 = ~\f2_pad  & ~n115 ;
  assign n461 = ~\g2_pad  & n115 ;
  assign n462 = ~n460 & ~n461 ;
  assign n463 = ~n114 & n462 ;
  assign n464 = ~n459 & ~n463 ;
  assign n465 = ~\i0_pad  & ~n464 ;
  assign n466 = ~\g1_pad  & ~n99 ;
  assign n467 = ~\p0_pad  & ~\r2_pad  ;
  assign n468 = n95 & n467 ;
  assign n469 = n98 & n468 ;
  assign n470 = ~\c1_pad  & ~n469 ;
  assign n471 = ~n466 & n470 ;
  assign n472 = \b0_pad  & \m1_pad  ;
  assign n473 = n109 & n472 ;
  assign n474 = ~n108 & n473 ;
  assign n475 = ~\g2_pad  & ~n115 ;
  assign n476 = ~\h2_pad  & n115 ;
  assign n477 = ~n475 & ~n476 ;
  assign n478 = ~n114 & n477 ;
  assign n479 = ~n474 & ~n478 ;
  assign n480 = ~\i0_pad  & ~n479 ;
  assign \a3_pad  = ~\j1_pad  ;
  assign \a4_pad  = n105 ;
  assign \a5_pad  = n121 ;
  assign \b3_pad  = ~\k1_pad  ;
  assign \b4_pad  = n127 ;
  assign \b5_pad  = n136 ;
  assign \c3_pad  = ~n150 ;
  assign \c4_pad  = n156 ;
  assign \c5_pad  = ~n164 ;
  assign \d3_pad  = ~n171 ;
  assign \d4_pad  = n177 ;
  assign \d5_pad  = n185 ;
  assign \e3_pad  = n188 ;
  assign \e4_pad  = n190 ;
  assign \e5_pad  = n200 ;
  assign \f3_pad  = ~n205 ;
  assign \f4_pad  = n210 ;
  assign \f5_pad  = n219 ;
  assign \g3_pad  = n222 ;
  assign \g4_pad  = n232 ;
  assign \g5_pad  = n241 ;
  assign \h3_pad  = n242 ;
  assign \h4_pad  = ~n247 ;
  assign \h5_pad  = ~n252 ;
  assign \i3_pad  = n253 ;
  assign \i4_pad  = ~n259 ;
  assign \i5_pad  = n265 ;
  assign \j3_pad  = n266 ;
  assign \j4_pad  = n275 ;
  assign \j5_pad  = n281 ;
  assign \k3_pad  = n282 ;
  assign \k4_pad  = n291 ;
  assign \k5_pad  = ~n296 ;
  assign \l3_pad  = n297 ;
  assign \l4_pad  = n306 ;
  assign \l5_pad  = ~n311 ;
  assign \m3_pad  = n312 ;
  assign \m4_pad  = n321 ;
  assign \m5_pad  = ~n327 ;
  assign \n3_pad  = n328 ;
  assign \n4_pad  = n337 ;
  assign \n5_pad  = n340 ;
  assign \o3_pad  = n341 ;
  assign \o4_pad  = n350 ;
  assign \o5_pad  = n353 ;
  assign \p3_pad  = n354 ;
  assign \p4_pad  = n363 ;
  assign \q3_pad  = n364 ;
  assign \q4_pad  = n373 ;
  assign \r3_pad  = n374 ;
  assign \r4_pad  = n383 ;
  assign \s3_pad  = n384 ;
  assign \s4_pad  = n393 ;
  assign \t3_pad  = n394 ;
  assign \t4_pad  = n403 ;
  assign \u3_pad  = n404 ;
  assign \u4_pad  = n413 ;
  assign \v3_pad  = ~n415 ;
  assign \v4_pad  = n424 ;
  assign \w2_pad  = ~\f1_pad  ;
  assign \w3_pad  = n428 ;
  assign \w4_pad  = n437 ;
  assign \x2_pad  = ~\g1_pad  ;
  assign \x3_pad  = ~n441 ;
  assign \x4_pad  = n450 ;
  assign \y2_pad  = ~\h1_pad  ;
  assign \y3_pad  = n456 ;
  assign \y4_pad  = n465 ;
  assign \z2_pad  = ~\i1_pad  ;
  assign \z3_pad  = n471 ;
  assign \z4_pad  = n480 ;
endmodule
