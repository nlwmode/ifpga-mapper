module top (\cnt10_pad , \cnt13_pad , \cnt21_pad , \cnt261_pad , \cnt272_pad , \cnt283_pad , \cnt284_pad , \cnt44_pad , \cnt45_pad , \cnt509_pad , \cnt511_pad , \cnt567_pad , \cnt591_pad , john_pad, \pcnt12_pad , \pcnt17_pad , \pcnt241_pad , \pcnt27_pad , \pcnt6_pad , \st_0_reg/NET0131 , \st_1_reg/NET0131 , \st_2_reg/NET0131 , \st_3_reg/NET0131 , \st_4_reg/NET0131 , \st_5_reg/NET0131 , \_al_n0 , \_al_n1 , cblank_pad, cclr_pad, csm_pad, csync_pad, \g1235/_0_ , \g1258/_0_ , \g1273/_0_ , \g52/_0_ , \g869/_0_ , \g886/_0_ , pc_pad, pclr_pad, vsync_pad);
	input \cnt10_pad  ;
	input \cnt13_pad  ;
	input \cnt21_pad  ;
	input \cnt261_pad  ;
	input \cnt272_pad  ;
	input \cnt283_pad  ;
	input \cnt284_pad  ;
	input \cnt44_pad  ;
	input \cnt45_pad  ;
	input \cnt509_pad  ;
	input \cnt511_pad  ;
	input \cnt567_pad  ;
	input \cnt591_pad  ;
	input john_pad ;
	input \pcnt12_pad  ;
	input \pcnt17_pad  ;
	input \pcnt241_pad  ;
	input \pcnt27_pad  ;
	input \pcnt6_pad  ;
	input \st_0_reg/NET0131  ;
	input \st_1_reg/NET0131  ;
	input \st_2_reg/NET0131  ;
	input \st_3_reg/NET0131  ;
	input \st_4_reg/NET0131  ;
	input \st_5_reg/NET0131  ;
	output \_al_n0  ;
	output \_al_n1  ;
	output cblank_pad ;
	output cclr_pad ;
	output csm_pad ;
	output csync_pad ;
	output \g1235/_0_  ;
	output \g1258/_0_  ;
	output \g1273/_0_  ;
	output \g52/_0_  ;
	output \g869/_0_  ;
	output \g886/_0_  ;
	output pc_pad ;
	output pclr_pad ;
	output vsync_pad ;
	wire _w233_ ;
	wire _w232_ ;
	wire _w231_ ;
	wire _w230_ ;
	wire _w229_ ;
	wire _w228_ ;
	wire _w227_ ;
	wire _w226_ ;
	wire _w225_ ;
	wire _w224_ ;
	wire _w223_ ;
	wire _w222_ ;
	wire _w221_ ;
	wire _w220_ ;
	wire _w219_ ;
	wire _w218_ ;
	wire _w217_ ;
	wire _w216_ ;
	wire _w215_ ;
	wire _w214_ ;
	wire _w213_ ;
	wire _w212_ ;
	wire _w211_ ;
	wire _w210_ ;
	wire _w209_ ;
	wire _w208_ ;
	wire _w207_ ;
	wire _w206_ ;
	wire _w205_ ;
	wire _w204_ ;
	wire _w203_ ;
	wire _w202_ ;
	wire _w201_ ;
	wire _w200_ ;
	wire _w199_ ;
	wire _w198_ ;
	wire _w197_ ;
	wire _w196_ ;
	wire _w195_ ;
	wire _w194_ ;
	wire _w193_ ;
	wire _w192_ ;
	wire _w191_ ;
	wire _w190_ ;
	wire _w189_ ;
	wire _w188_ ;
	wire _w187_ ;
	wire _w186_ ;
	wire _w185_ ;
	wire _w184_ ;
	wire _w183_ ;
	wire _w182_ ;
	wire _w181_ ;
	wire _w180_ ;
	wire _w179_ ;
	wire _w178_ ;
	wire _w177_ ;
	wire _w176_ ;
	wire _w175_ ;
	wire _w174_ ;
	wire _w173_ ;
	wire _w172_ ;
	wire _w171_ ;
	wire _w170_ ;
	wire _w169_ ;
	wire _w168_ ;
	wire _w167_ ;
	wire _w166_ ;
	wire _w165_ ;
	wire _w164_ ;
	wire _w163_ ;
	wire _w162_ ;
	wire _w161_ ;
	wire _w160_ ;
	wire _w159_ ;
	wire _w158_ ;
	wire _w157_ ;
	wire _w156_ ;
	wire _w155_ ;
	wire _w154_ ;
	wire _w153_ ;
	wire _w84_ ;
	wire _w83_ ;
	wire _w82_ ;
	wire _w81_ ;
	wire _w80_ ;
	wire _w79_ ;
	wire _w78_ ;
	wire _w77_ ;
	wire _w76_ ;
	wire _w75_ ;
	wire _w74_ ;
	wire _w73_ ;
	wire _w72_ ;
	wire _w71_ ;
	wire _w70_ ;
	wire _w69_ ;
	wire _w68_ ;
	wire _w67_ ;
	wire _w66_ ;
	wire _w65_ ;
	wire _w64_ ;
	wire _w63_ ;
	wire _w62_ ;
	wire _w61_ ;
	wire _w60_ ;
	wire _w59_ ;
	wire _w58_ ;
	wire _w57_ ;
	wire _w56_ ;
	wire _w55_ ;
	wire _w38_ ;
	wire _w37_ ;
	wire _w36_ ;
	wire _w35_ ;
	wire _w34_ ;
	wire _w33_ ;
	wire _w32_ ;
	wire _w31_ ;
	wire _w30_ ;
	wire _w29_ ;
	wire _w28_ ;
	wire _w27_ ;
	wire _w26_ ;
	wire _w39_ ;
	wire _w40_ ;
	wire _w41_ ;
	wire _w42_ ;
	wire _w43_ ;
	wire _w44_ ;
	wire _w45_ ;
	wire _w46_ ;
	wire _w47_ ;
	wire _w48_ ;
	wire _w49_ ;
	wire _w50_ ;
	wire _w51_ ;
	wire _w52_ ;
	wire _w53_ ;
	wire _w54_ ;
	wire _w85_ ;
	wire _w86_ ;
	wire _w87_ ;
	wire _w88_ ;
	wire _w89_ ;
	wire _w90_ ;
	wire _w91_ ;
	wire _w92_ ;
	wire _w93_ ;
	wire _w94_ ;
	wire _w95_ ;
	wire _w96_ ;
	wire _w97_ ;
	wire _w98_ ;
	wire _w99_ ;
	wire _w100_ ;
	wire _w101_ ;
	wire _w102_ ;
	wire _w103_ ;
	wire _w104_ ;
	wire _w105_ ;
	wire _w106_ ;
	wire _w107_ ;
	wire _w108_ ;
	wire _w109_ ;
	wire _w110_ ;
	wire _w111_ ;
	wire _w112_ ;
	wire _w113_ ;
	wire _w114_ ;
	wire _w115_ ;
	wire _w116_ ;
	wire _w117_ ;
	wire _w118_ ;
	wire _w119_ ;
	wire _w120_ ;
	wire _w121_ ;
	wire _w122_ ;
	wire _w123_ ;
	wire _w124_ ;
	wire _w125_ ;
	wire _w126_ ;
	wire _w127_ ;
	wire _w128_ ;
	wire _w129_ ;
	wire _w130_ ;
	wire _w131_ ;
	wire _w132_ ;
	wire _w133_ ;
	wire _w134_ ;
	wire _w135_ ;
	wire _w136_ ;
	wire _w137_ ;
	wire _w138_ ;
	wire _w139_ ;
	wire _w140_ ;
	wire _w141_ ;
	wire _w142_ ;
	wire _w143_ ;
	wire _w144_ ;
	wire _w145_ ;
	wire _w146_ ;
	wire _w147_ ;
	wire _w148_ ;
	wire _w149_ ;
	wire _w150_ ;
	wire _w151_ ;
	wire _w152_ ;
	LUT2 #(
		.INIT('h2)
	) name0 (
		\st_3_reg/NET0131 ,
		\st_4_reg/NET0131 ,
		_w26_
	);
	LUT2 #(
		.INIT('h8)
	) name1 (
		\st_2_reg/NET0131 ,
		_w26_,
		_w27_
	);
	LUT2 #(
		.INIT('h4)
	) name2 (
		\st_0_reg/NET0131 ,
		_w27_,
		_w28_
	);
	LUT2 #(
		.INIT('h8)
	) name3 (
		\st_3_reg/NET0131 ,
		\st_4_reg/NET0131 ,
		_w29_
	);
	LUT2 #(
		.INIT('h1)
	) name4 (
		\st_5_reg/NET0131 ,
		_w29_,
		_w30_
	);
	LUT2 #(
		.INIT('h2)
	) name5 (
		\st_0_reg/NET0131 ,
		\st_2_reg/NET0131 ,
		_w31_
	);
	LUT2 #(
		.INIT('h8)
	) name6 (
		\st_1_reg/NET0131 ,
		_w31_,
		_w32_
	);
	LUT2 #(
		.INIT('h4)
	) name7 (
		_w30_,
		_w32_,
		_w33_
	);
	LUT2 #(
		.INIT('h8)
	) name8 (
		\st_2_reg/NET0131 ,
		\st_5_reg/NET0131 ,
		_w34_
	);
	LUT2 #(
		.INIT('h8)
	) name9 (
		\st_3_reg/NET0131 ,
		_w34_,
		_w35_
	);
	LUT2 #(
		.INIT('h1)
	) name10 (
		_w28_,
		_w35_,
		_w36_
	);
	LUT2 #(
		.INIT('h4)
	) name11 (
		_w33_,
		_w36_,
		_w37_
	);
	LUT2 #(
		.INIT('h1)
	) name12 (
		\st_0_reg/NET0131 ,
		\st_1_reg/NET0131 ,
		_w38_
	);
	LUT2 #(
		.INIT('h2)
	) name13 (
		\st_2_reg/NET0131 ,
		\st_3_reg/NET0131 ,
		_w39_
	);
	LUT2 #(
		.INIT('h8)
	) name14 (
		_w38_,
		_w39_,
		_w40_
	);
	LUT2 #(
		.INIT('h8)
	) name15 (
		\st_5_reg/NET0131 ,
		_w40_,
		_w41_
	);
	LUT2 #(
		.INIT('h1)
	) name16 (
		\st_3_reg/NET0131 ,
		\st_5_reg/NET0131 ,
		_w42_
	);
	LUT2 #(
		.INIT('h1)
	) name17 (
		\st_1_reg/NET0131 ,
		\st_2_reg/NET0131 ,
		_w43_
	);
	LUT2 #(
		.INIT('h8)
	) name18 (
		_w42_,
		_w43_,
		_w44_
	);
	LUT2 #(
		.INIT('h4)
	) name19 (
		\st_4_reg/NET0131 ,
		_w44_,
		_w45_
	);
	LUT2 #(
		.INIT('h8)
	) name20 (
		\st_0_reg/NET0131 ,
		\st_1_reg/NET0131 ,
		_w46_
	);
	LUT2 #(
		.INIT('h4)
	) name21 (
		_w42_,
		_w46_,
		_w47_
	);
	LUT2 #(
		.INIT('h2)
	) name22 (
		\st_0_reg/NET0131 ,
		\st_5_reg/NET0131 ,
		_w48_
	);
	LUT2 #(
		.INIT('h4)
	) name23 (
		\st_1_reg/NET0131 ,
		_w48_,
		_w49_
	);
	LUT2 #(
		.INIT('h8)
	) name24 (
		\st_0_reg/NET0131 ,
		\st_4_reg/NET0131 ,
		_w50_
	);
	LUT2 #(
		.INIT('h1)
	) name25 (
		_w31_,
		_w50_,
		_w51_
	);
	LUT2 #(
		.INIT('h4)
	) name26 (
		_w47_,
		_w51_,
		_w52_
	);
	LUT2 #(
		.INIT('h4)
	) name27 (
		_w49_,
		_w52_,
		_w53_
	);
	LUT2 #(
		.INIT('h1)
	) name28 (
		_w41_,
		_w45_,
		_w54_
	);
	LUT2 #(
		.INIT('h8)
	) name29 (
		_w53_,
		_w54_,
		_w55_
	);
	LUT2 #(
		.INIT('h2)
	) name30 (
		_w35_,
		_w38_,
		_w56_
	);
	LUT2 #(
		.INIT('h1)
	) name31 (
		\st_4_reg/NET0131 ,
		\st_5_reg/NET0131 ,
		_w57_
	);
	LUT2 #(
		.INIT('h1)
	) name32 (
		\st_2_reg/NET0131 ,
		_w57_,
		_w58_
	);
	LUT2 #(
		.INIT('h8)
	) name33 (
		\st_0_reg/NET0131 ,
		_w58_,
		_w59_
	);
	LUT2 #(
		.INIT('h2)
	) name34 (
		\st_1_reg/NET0131 ,
		_w42_,
		_w60_
	);
	LUT2 #(
		.INIT('h8)
	) name35 (
		\st_1_reg/NET0131 ,
		\st_2_reg/NET0131 ,
		_w61_
	);
	LUT2 #(
		.INIT('h1)
	) name36 (
		_w43_,
		_w61_,
		_w62_
	);
	LUT2 #(
		.INIT('h4)
	) name37 (
		\st_4_reg/NET0131 ,
		_w62_,
		_w63_
	);
	LUT2 #(
		.INIT('h1)
	) name38 (
		_w60_,
		_w63_,
		_w64_
	);
	LUT2 #(
		.INIT('h1)
	) name39 (
		\st_0_reg/NET0131 ,
		_w64_,
		_w65_
	);
	LUT2 #(
		.INIT('h4)
	) name40 (
		\st_0_reg/NET0131 ,
		\st_3_reg/NET0131 ,
		_w66_
	);
	LUT2 #(
		.INIT('h4)
	) name41 (
		\st_5_reg/NET0131 ,
		_w66_,
		_w67_
	);
	LUT2 #(
		.INIT('h2)
	) name42 (
		\st_1_reg/NET0131 ,
		\st_5_reg/NET0131 ,
		_w68_
	);
	LUT2 #(
		.INIT('h8)
	) name43 (
		\st_0_reg/NET0131 ,
		\st_2_reg/NET0131 ,
		_w69_
	);
	LUT2 #(
		.INIT('h8)
	) name44 (
		_w68_,
		_w69_,
		_w70_
	);
	LUT2 #(
		.INIT('h1)
	) name45 (
		_w67_,
		_w70_,
		_w71_
	);
	LUT2 #(
		.INIT('h1)
	) name46 (
		\st_4_reg/NET0131 ,
		_w71_,
		_w72_
	);
	LUT2 #(
		.INIT('h4)
	) name47 (
		\st_1_reg/NET0131 ,
		_w50_,
		_w73_
	);
	LUT2 #(
		.INIT('h1)
	) name48 (
		_w27_,
		_w73_,
		_w74_
	);
	LUT2 #(
		.INIT('h4)
	) name49 (
		_w59_,
		_w74_,
		_w75_
	);
	LUT2 #(
		.INIT('h4)
	) name50 (
		_w72_,
		_w75_,
		_w76_
	);
	LUT2 #(
		.INIT('h4)
	) name51 (
		_w65_,
		_w76_,
		_w77_
	);
	LUT2 #(
		.INIT('h8)
	) name52 (
		\st_3_reg/NET0131 ,
		_w58_,
		_w78_
	);
	LUT2 #(
		.INIT('h4)
	) name53 (
		\st_4_reg/NET0131 ,
		_w31_,
		_w79_
	);
	LUT2 #(
		.INIT('h1)
	) name54 (
		\st_5_reg/NET0131 ,
		_w79_,
		_w80_
	);
	LUT2 #(
		.INIT('h2)
	) name55 (
		_w46_,
		_w80_,
		_w81_
	);
	LUT2 #(
		.INIT('h4)
	) name56 (
		\st_3_reg/NET0131 ,
		_w50_,
		_w82_
	);
	LUT2 #(
		.INIT('h1)
	) name57 (
		_w27_,
		_w82_,
		_w83_
	);
	LUT2 #(
		.INIT('h1)
	) name58 (
		\st_1_reg/NET0131 ,
		_w83_,
		_w84_
	);
	LUT2 #(
		.INIT('h1)
	) name59 (
		_w67_,
		_w78_,
		_w85_
	);
	LUT2 #(
		.INIT('h4)
	) name60 (
		_w81_,
		_w85_,
		_w86_
	);
	LUT2 #(
		.INIT('h4)
	) name61 (
		_w84_,
		_w86_,
		_w87_
	);
	LUT2 #(
		.INIT('h8)
	) name62 (
		\st_2_reg/NET0131 ,
		\st_3_reg/NET0131 ,
		_w88_
	);
	LUT2 #(
		.INIT('h8)
	) name63 (
		_w46_,
		_w88_,
		_w89_
	);
	LUT2 #(
		.INIT('h4)
	) name64 (
		\st_0_reg/NET0131 ,
		\st_1_reg/NET0131 ,
		_w90_
	);
	LUT2 #(
		.INIT('h2)
	) name65 (
		\st_3_reg/NET0131 ,
		_w90_,
		_w91_
	);
	LUT2 #(
		.INIT('h1)
	) name66 (
		\st_0_reg/NET0131 ,
		\st_2_reg/NET0131 ,
		_w92_
	);
	LUT2 #(
		.INIT('h1)
	) name67 (
		_w69_,
		_w92_,
		_w93_
	);
	LUT2 #(
		.INIT('h4)
	) name68 (
		_w91_,
		_w93_,
		_w94_
	);
	LUT2 #(
		.INIT('h2)
	) name69 (
		\st_5_reg/NET0131 ,
		_w94_,
		_w95_
	);
	LUT2 #(
		.INIT('h1)
	) name70 (
		\st_1_reg/NET0131 ,
		_w79_,
		_w96_
	);
	LUT2 #(
		.INIT('h1)
	) name71 (
		\st_3_reg/NET0131 ,
		_w46_,
		_w97_
	);
	LUT2 #(
		.INIT('h4)
	) name72 (
		_w68_,
		_w97_,
		_w98_
	);
	LUT2 #(
		.INIT('h4)
	) name73 (
		_w96_,
		_w98_,
		_w99_
	);
	LUT2 #(
		.INIT('h1)
	) name74 (
		_w89_,
		_w95_,
		_w100_
	);
	LUT2 #(
		.INIT('h4)
	) name75 (
		_w99_,
		_w100_,
		_w101_
	);
	LUT2 #(
		.INIT('h8)
	) name76 (
		\st_1_reg/NET0131 ,
		\st_3_reg/NET0131 ,
		_w102_
	);
	LUT2 #(
		.INIT('h2)
	) name77 (
		_w31_,
		_w102_,
		_w103_
	);
	LUT2 #(
		.INIT('h8)
	) name78 (
		\st_5_reg/NET0131 ,
		_w103_,
		_w104_
	);
	LUT2 #(
		.INIT('h4)
	) name79 (
		\st_2_reg/NET0131 ,
		_w90_,
		_w105_
	);
	LUT2 #(
		.INIT('h2)
	) name80 (
		\cnt567_pad ,
		\pcnt27_pad ,
		_w106_
	);
	LUT2 #(
		.INIT('h2)
	) name81 (
		_w105_,
		_w106_,
		_w107_
	);
	LUT2 #(
		.INIT('h1)
	) name82 (
		_w73_,
		_w107_,
		_w108_
	);
	LUT2 #(
		.INIT('h2)
	) name83 (
		\st_3_reg/NET0131 ,
		_w108_,
		_w109_
	);
	LUT2 #(
		.INIT('h4)
	) name84 (
		\st_3_reg/NET0131 ,
		_w34_,
		_w110_
	);
	LUT2 #(
		.INIT('h1)
	) name85 (
		_w45_,
		_w110_,
		_w111_
	);
	LUT2 #(
		.INIT('h1)
	) name86 (
		\st_0_reg/NET0131 ,
		_w111_,
		_w112_
	);
	LUT2 #(
		.INIT('h8)
	) name87 (
		\cnt284_pad ,
		\pcnt17_pad ,
		_w113_
	);
	LUT2 #(
		.INIT('h2)
	) name88 (
		_w70_,
		_w113_,
		_w114_
	);
	LUT2 #(
		.INIT('h2)
	) name89 (
		\cnt44_pad ,
		\pcnt12_pad ,
		_w115_
	);
	LUT2 #(
		.INIT('h2)
	) name90 (
		_w105_,
		_w115_,
		_w116_
	);
	LUT2 #(
		.INIT('h1)
	) name91 (
		_w114_,
		_w116_,
		_w117_
	);
	LUT2 #(
		.INIT('h1)
	) name92 (
		\st_3_reg/NET0131 ,
		_w117_,
		_w118_
	);
	LUT2 #(
		.INIT('h4)
	) name93 (
		\cnt13_pad ,
		_w39_,
		_w119_
	);
	LUT2 #(
		.INIT('h2)
	) name94 (
		_w57_,
		_w119_,
		_w120_
	);
	LUT2 #(
		.INIT('h2)
	) name95 (
		_w90_,
		_w120_,
		_w121_
	);
	LUT2 #(
		.INIT('h2)
	) name96 (
		\cnt511_pad ,
		\pcnt241_pad ,
		_w122_
	);
	LUT2 #(
		.INIT('h8)
	) name97 (
		_w88_,
		_w90_,
		_w123_
	);
	LUT2 #(
		.INIT('h4)
	) name98 (
		_w122_,
		_w123_,
		_w124_
	);
	LUT2 #(
		.INIT('h1)
	) name99 (
		\st_3_reg/NET0131 ,
		\st_4_reg/NET0131 ,
		_w125_
	);
	LUT2 #(
		.INIT('h4)
	) name100 (
		_w29_,
		_w69_,
		_w126_
	);
	LUT2 #(
		.INIT('h4)
	) name101 (
		_w125_,
		_w126_,
		_w127_
	);
	LUT2 #(
		.INIT('h1)
	) name102 (
		_w104_,
		_w124_,
		_w128_
	);
	LUT2 #(
		.INIT('h4)
	) name103 (
		_w127_,
		_w128_,
		_w129_
	);
	LUT2 #(
		.INIT('h4)
	) name104 (
		_w121_,
		_w129_,
		_w130_
	);
	LUT2 #(
		.INIT('h1)
	) name105 (
		_w109_,
		_w112_,
		_w131_
	);
	LUT2 #(
		.INIT('h4)
	) name106 (
		_w118_,
		_w131_,
		_w132_
	);
	LUT2 #(
		.INIT('h8)
	) name107 (
		_w130_,
		_w132_,
		_w133_
	);
	LUT2 #(
		.INIT('h8)
	) name108 (
		\cnt511_pad ,
		_w123_,
		_w134_
	);
	LUT2 #(
		.INIT('h8)
	) name109 (
		\cnt284_pad ,
		\pcnt6_pad ,
		_w135_
	);
	LUT2 #(
		.INIT('h8)
	) name110 (
		_w40_,
		_w135_,
		_w136_
	);
	LUT2 #(
		.INIT('h8)
	) name111 (
		\cnt567_pad ,
		\st_3_reg/NET0131 ,
		_w137_
	);
	LUT2 #(
		.INIT('h8)
	) name112 (
		_w105_,
		_w137_,
		_w138_
	);
	LUT2 #(
		.INIT('h1)
	) name113 (
		_w134_,
		_w136_,
		_w139_
	);
	LUT2 #(
		.INIT('h4)
	) name114 (
		_w138_,
		_w139_,
		_w140_
	);
	LUT2 #(
		.INIT('h2)
	) name115 (
		_w57_,
		_w140_,
		_w141_
	);
	LUT2 #(
		.INIT('h4)
	) name116 (
		\st_1_reg/NET0131 ,
		_w88_,
		_w142_
	);
	LUT2 #(
		.INIT('h8)
	) name117 (
		\cnt509_pad ,
		\st_5_reg/NET0131 ,
		_w143_
	);
	LUT2 #(
		.INIT('h8)
	) name118 (
		_w142_,
		_w143_,
		_w144_
	);
	LUT2 #(
		.INIT('h8)
	) name119 (
		\cnt45_pad ,
		_w43_,
		_w145_
	);
	LUT2 #(
		.INIT('h4)
	) name120 (
		_w30_,
		_w145_,
		_w146_
	);
	LUT2 #(
		.INIT('h1)
	) name121 (
		_w144_,
		_w146_,
		_w147_
	);
	LUT2 #(
		.INIT('h1)
	) name122 (
		\st_0_reg/NET0131 ,
		_w147_,
		_w148_
	);
	LUT2 #(
		.INIT('h8)
	) name123 (
		john_pad,
		\st_4_reg/NET0131 ,
		_w149_
	);
	LUT2 #(
		.INIT('h8)
	) name124 (
		\cnt10_pad ,
		\st_5_reg/NET0131 ,
		_w150_
	);
	LUT2 #(
		.INIT('h1)
	) name125 (
		_w149_,
		_w150_,
		_w151_
	);
	LUT2 #(
		.INIT('h8)
	) name126 (
		_w39_,
		_w90_,
		_w152_
	);
	LUT2 #(
		.INIT('h4)
	) name127 (
		_w151_,
		_w152_,
		_w153_
	);
	LUT2 #(
		.INIT('h4)
	) name128 (
		\cnt261_pad ,
		\st_0_reg/NET0131 ,
		_w154_
	);
	LUT2 #(
		.INIT('h4)
	) name129 (
		\st_1_reg/NET0131 ,
		_w154_,
		_w155_
	);
	LUT2 #(
		.INIT('h8)
	) name130 (
		_w110_,
		_w155_,
		_w156_
	);
	LUT2 #(
		.INIT('h8)
	) name131 (
		\st_0_reg/NET0131 ,
		_w42_,
		_w157_
	);
	LUT2 #(
		.INIT('h1)
	) name132 (
		\st_4_reg/NET0131 ,
		_w62_,
		_w158_
	);
	LUT2 #(
		.INIT('h8)
	) name133 (
		_w157_,
		_w158_,
		_w159_
	);
	LUT2 #(
		.INIT('h4)
	) name134 (
		\cnt272_pad ,
		\st_2_reg/NET0131 ,
		_w160_
	);
	LUT2 #(
		.INIT('h4)
	) name135 (
		\st_5_reg/NET0131 ,
		_w26_,
		_w161_
	);
	LUT2 #(
		.INIT('h1)
	) name136 (
		\cnt591_pad ,
		\st_2_reg/NET0131 ,
		_w162_
	);
	LUT2 #(
		.INIT('h2)
	) name137 (
		_w38_,
		_w160_,
		_w163_
	);
	LUT2 #(
		.INIT('h4)
	) name138 (
		_w162_,
		_w163_,
		_w164_
	);
	LUT2 #(
		.INIT('h8)
	) name139 (
		_w161_,
		_w164_,
		_w165_
	);
	LUT2 #(
		.INIT('h1)
	) name140 (
		\st_5_reg/NET0131 ,
		_w125_,
		_w166_
	);
	LUT2 #(
		.INIT('h8)
	) name141 (
		\cnt44_pad ,
		_w105_,
		_w167_
	);
	LUT2 #(
		.INIT('h4)
	) name142 (
		_w166_,
		_w167_,
		_w168_
	);
	LUT2 #(
		.INIT('h8)
	) name143 (
		\cnt45_pad ,
		_w40_,
		_w169_
	);
	LUT2 #(
		.INIT('h2)
	) name144 (
		\cnt21_pad ,
		\st_3_reg/NET0131 ,
		_w170_
	);
	LUT2 #(
		.INIT('h8)
	) name145 (
		\cnt283_pad ,
		_w102_,
		_w171_
	);
	LUT2 #(
		.INIT('h1)
	) name146 (
		_w170_,
		_w171_,
		_w172_
	);
	LUT2 #(
		.INIT('h2)
	) name147 (
		_w92_,
		_w172_,
		_w173_
	);
	LUT2 #(
		.INIT('h1)
	) name148 (
		\cnt21_pad ,
		\st_0_reg/NET0131 ,
		_w174_
	);
	LUT2 #(
		.INIT('h2)
	) name149 (
		_w142_,
		_w174_,
		_w175_
	);
	LUT2 #(
		.INIT('h8)
	) name150 (
		\cnt10_pad ,
		_w123_,
		_w176_
	);
	LUT2 #(
		.INIT('h1)
	) name151 (
		_w169_,
		_w175_,
		_w177_
	);
	LUT2 #(
		.INIT('h4)
	) name152 (
		_w176_,
		_w177_,
		_w178_
	);
	LUT2 #(
		.INIT('h4)
	) name153 (
		_w173_,
		_w178_,
		_w179_
	);
	LUT2 #(
		.INIT('h2)
	) name154 (
		\st_4_reg/NET0131 ,
		_w179_,
		_w180_
	);
	LUT2 #(
		.INIT('h1)
	) name155 (
		_w153_,
		_w156_,
		_w181_
	);
	LUT2 #(
		.INIT('h4)
	) name156 (
		_w159_,
		_w181_,
		_w182_
	);
	LUT2 #(
		.INIT('h1)
	) name157 (
		_w165_,
		_w168_,
		_w183_
	);
	LUT2 #(
		.INIT('h8)
	) name158 (
		_w182_,
		_w183_,
		_w184_
	);
	LUT2 #(
		.INIT('h4)
	) name159 (
		_w148_,
		_w184_,
		_w185_
	);
	LUT2 #(
		.INIT('h4)
	) name160 (
		_w141_,
		_w185_,
		_w186_
	);
	LUT2 #(
		.INIT('h4)
	) name161 (
		_w180_,
		_w186_,
		_w187_
	);
	LUT2 #(
		.INIT('h8)
	) name162 (
		\st_2_reg/NET0131 ,
		\st_4_reg/NET0131 ,
		_w188_
	);
	LUT2 #(
		.INIT('h4)
	) name163 (
		\st_1_reg/NET0131 ,
		\st_2_reg/NET0131 ,
		_w189_
	);
	LUT2 #(
		.INIT('h4)
	) name164 (
		\st_5_reg/NET0131 ,
		_w189_,
		_w190_
	);
	LUT2 #(
		.INIT('h4)
	) name165 (
		\cnt284_pad ,
		_w190_,
		_w191_
	);
	LUT2 #(
		.INIT('h1)
	) name166 (
		_w188_,
		_w191_,
		_w192_
	);
	LUT2 #(
		.INIT('h1)
	) name167 (
		\st_0_reg/NET0131 ,
		_w192_,
		_w193_
	);
	LUT2 #(
		.INIT('h4)
	) name168 (
		\st_2_reg/NET0131 ,
		_w49_,
		_w194_
	);
	LUT2 #(
		.INIT('h1)
	) name169 (
		_w88_,
		_w194_,
		_w195_
	);
	LUT2 #(
		.INIT('h1)
	) name170 (
		\st_4_reg/NET0131 ,
		_w195_,
		_w196_
	);
	LUT2 #(
		.INIT('h8)
	) name171 (
		\st_0_reg/NET0131 ,
		\st_5_reg/NET0131 ,
		_w197_
	);
	LUT2 #(
		.INIT('h8)
	) name172 (
		_w62_,
		_w197_,
		_w198_
	);
	LUT2 #(
		.INIT('h2)
	) name173 (
		\cnt13_pad ,
		\st_5_reg/NET0131 ,
		_w199_
	);
	LUT2 #(
		.INIT('h8)
	) name174 (
		\st_2_reg/NET0131 ,
		_w90_,
		_w200_
	);
	LUT2 #(
		.INIT('h4)
	) name175 (
		_w199_,
		_w200_,
		_w201_
	);
	LUT2 #(
		.INIT('h2)
	) name176 (
		\cnt284_pad ,
		\pcnt17_pad ,
		_w202_
	);
	LUT2 #(
		.INIT('h2)
	) name177 (
		_w157_,
		_w202_,
		_w203_
	);
	LUT2 #(
		.INIT('h4)
	) name178 (
		_w26_,
		_w31_,
		_w204_
	);
	LUT2 #(
		.INIT('h1)
	) name179 (
		_w82_,
		_w204_,
		_w205_
	);
	LUT2 #(
		.INIT('h4)
	) name180 (
		_w203_,
		_w205_,
		_w206_
	);
	LUT2 #(
		.INIT('h2)
	) name181 (
		\st_1_reg/NET0131 ,
		_w206_,
		_w207_
	);
	LUT2 #(
		.INIT('h1)
	) name182 (
		_w142_,
		_w198_,
		_w208_
	);
	LUT2 #(
		.INIT('h4)
	) name183 (
		_w201_,
		_w208_,
		_w209_
	);
	LUT2 #(
		.INIT('h4)
	) name184 (
		_w193_,
		_w209_,
		_w210_
	);
	LUT2 #(
		.INIT('h1)
	) name185 (
		_w196_,
		_w207_,
		_w211_
	);
	LUT2 #(
		.INIT('h8)
	) name186 (
		_w210_,
		_w211_,
		_w212_
	);
	LUT2 #(
		.INIT('h8)
	) name187 (
		_w48_,
		_w63_,
		_w213_
	);
	LUT2 #(
		.INIT('h1)
	) name188 (
		\st_4_reg/NET0131 ,
		_w44_,
		_w214_
	);
	LUT2 #(
		.INIT('h1)
	) name189 (
		\st_0_reg/NET0131 ,
		_w214_,
		_w215_
	);
	LUT2 #(
		.INIT('h8)
	) name190 (
		\st_1_reg/NET0131 ,
		_w34_,
		_w216_
	);
	LUT2 #(
		.INIT('h1)
	) name191 (
		_w194_,
		_w216_,
		_w217_
	);
	LUT2 #(
		.INIT('h2)
	) name192 (
		\st_3_reg/NET0131 ,
		_w217_,
		_w218_
	);
	LUT2 #(
		.INIT('h1)
	) name193 (
		_w213_,
		_w215_,
		_w219_
	);
	LUT2 #(
		.INIT('h4)
	) name194 (
		_w218_,
		_w219_,
		_w220_
	);
	LUT2 #(
		.INIT('h8)
	) name195 (
		_w57_,
		_w103_,
		_w221_
	);
	LUT2 #(
		.INIT('h8)
	) name196 (
		\st_4_reg/NET0131 ,
		_w89_,
		_w222_
	);
	LUT2 #(
		.INIT('h1)
	) name197 (
		_w45_,
		_w221_,
		_w223_
	);
	LUT2 #(
		.INIT('h4)
	) name198 (
		_w222_,
		_w223_,
		_w224_
	);
	LUT2 #(
		.INIT('h8)
	) name199 (
		_w61_,
		_w82_,
		_w225_
	);
	LUT2 #(
		.INIT('h8)
	) name200 (
		_w32_,
		_w161_,
		_w226_
	);
	LUT2 #(
		.INIT('h1)
	) name201 (
		_w225_,
		_w226_,
		_w227_
	);
	LUT2 #(
		.INIT('h4)
	) name202 (
		\st_4_reg/NET0131 ,
		_w61_,
		_w228_
	);
	LUT2 #(
		.INIT('h4)
	) name203 (
		\st_2_reg/NET0131 ,
		_w38_,
		_w229_
	);
	LUT2 #(
		.INIT('h4)
	) name204 (
		_w58_,
		_w97_,
		_w230_
	);
	LUT2 #(
		.INIT('h1)
	) name205 (
		_w190_,
		_w228_,
		_w231_
	);
	LUT2 #(
		.INIT('h4)
	) name206 (
		_w229_,
		_w231_,
		_w232_
	);
	LUT2 #(
		.INIT('h8)
	) name207 (
		_w230_,
		_w232_,
		_w233_
	);
	assign \_al_n0  = 1'b0;
	assign \_al_n1  = 1'b0;
	assign cblank_pad = _w37_ ;
	assign cclr_pad = _w55_ ;
	assign csm_pad = _w56_ ;
	assign csync_pad = _w77_ ;
	assign \g1235/_0_  = _w87_ ;
	assign \g1258/_0_  = _w101_ ;
	assign \g1273/_0_  = _w133_ ;
	assign \g52/_0_  = _w187_ ;
	assign \g869/_0_  = _w212_ ;
	assign \g886/_0_  = _w220_ ;
	assign pc_pad = _w224_ ;
	assign pclr_pad = _w227_ ;
	assign vsync_pad = _w233_ ;
endmodule;