module top( \a0_pad  , a_pad , b_pad , c_pad , d_pad , e_pad , f_pad , g_pad , h_pad , i_pad , j_pad , k_pad , l_pad , m_pad , n_pad , o_pad , p_pad , q_pad , r_pad , s_pad , t_pad , u_pad , v_pad , w_pad , x_pad , y_pad , z_pad , \b0_pad  , \c0_pad  , \d0_pad  , \e0_pad  , \f0_pad  , \g0_pad  , \h0_pad  , \i0_pad  , \j0_pad  , \k0_pad  , \l0_pad  , \m0_pad  , \n0_pad  , \o0_pad  , \p0_pad  , \q0_pad  , \r0_pad  );
  input \a0_pad  ;
  input a_pad ;
  input b_pad ;
  input c_pad ;
  input d_pad ;
  input e_pad ;
  input f_pad ;
  input g_pad ;
  input h_pad ;
  input i_pad ;
  input j_pad ;
  input k_pad ;
  input l_pad ;
  input m_pad ;
  input n_pad ;
  input o_pad ;
  input p_pad ;
  input q_pad ;
  input r_pad ;
  input s_pad ;
  input t_pad ;
  input u_pad ;
  input v_pad ;
  input w_pad ;
  input x_pad ;
  input y_pad ;
  input z_pad ;
  output \b0_pad  ;
  output \c0_pad  ;
  output \d0_pad  ;
  output \e0_pad  ;
  output \f0_pad  ;
  output \g0_pad  ;
  output \h0_pad  ;
  output \i0_pad  ;
  output \j0_pad  ;
  output \k0_pad  ;
  output \l0_pad  ;
  output \m0_pad  ;
  output \n0_pad  ;
  output \o0_pad  ;
  output \p0_pad  ;
  output \q0_pad  ;
  output \r0_pad  ;
  wire n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 ;
  assign n28 = t_pad & u_pad ;
  assign n29 = v_pad & w_pad ;
  assign n30 = n28 & n29 ;
  assign n31 = x_pad & z_pad ;
  assign n32 = y_pad & n31 ;
  assign n33 = n30 & n32 ;
  assign n34 = ~i_pad & j_pad ;
  assign n35 = ~k_pad & n34 ;
  assign n36 = \a0_pad  & n35 ;
  assign n37 = n33 & n36 ;
  assign n38 = a_pad & i_pad ;
  assign n39 = b_pad & i_pad ;
  assign n40 = c_pad & i_pad ;
  assign n41 = d_pad & i_pad ;
  assign n42 = e_pad & i_pad ;
  assign n43 = f_pad & i_pad ;
  assign n44 = g_pad & i_pad ;
  assign n45 = h_pad & i_pad ;
  assign n46 = \a0_pad  & l_pad ;
  assign n47 = n35 & n46 ;
  assign n48 = n33 & n47 ;
  assign n49 = ~k_pad & ~t_pad ;
  assign n50 = n34 & n49 ;
  assign n51 = ~n38 & ~n50 ;
  assign n52 = ~n48 & n51 ;
  assign n53 = ~t_pad & ~u_pad ;
  assign n54 = ~n28 & ~n53 ;
  assign n55 = m_pad & ~n54 ;
  assign n56 = n37 & n55 ;
  assign n57 = n35 & n54 ;
  assign n58 = ~n39 & ~n57 ;
  assign n59 = ~n56 & n58 ;
  assign n60 = n_pad & ~v_pad ;
  assign n61 = ~n28 & n60 ;
  assign n62 = n_pad & v_pad ;
  assign n63 = n28 & n62 ;
  assign n64 = ~n61 & ~n63 ;
  assign n65 = n37 & ~n64 ;
  assign n66 = v_pad & n28 ;
  assign n67 = ~v_pad & ~n28 ;
  assign n68 = ~n66 & ~n67 ;
  assign n69 = n35 & n68 ;
  assign n70 = ~n40 & ~n69 ;
  assign n71 = ~n65 & n70 ;
  assign n72 = o_pad & ~w_pad ;
  assign n73 = ~n66 & n72 ;
  assign n74 = o_pad & w_pad ;
  assign n75 = n66 & n74 ;
  assign n76 = ~n73 & ~n75 ;
  assign n77 = n37 & ~n76 ;
  assign n78 = ~w_pad & ~n66 ;
  assign n79 = ~n30 & n35 ;
  assign n80 = ~n78 & n79 ;
  assign n81 = ~n41 & ~n80 ;
  assign n82 = ~n77 & n81 ;
  assign n83 = p_pad & ~x_pad ;
  assign n84 = ~n30 & n83 ;
  assign n85 = p_pad & x_pad ;
  assign n86 = n30 & n85 ;
  assign n87 = ~n84 & ~n86 ;
  assign n88 = n37 & ~n87 ;
  assign n89 = ~k_pad & x_pad ;
  assign n90 = n34 & n89 ;
  assign n91 = ~n30 & n90 ;
  assign n92 = ~k_pad & ~x_pad ;
  assign n93 = n34 & n92 ;
  assign n94 = n30 & n93 ;
  assign n95 = ~n91 & ~n94 ;
  assign n96 = ~n42 & n95 ;
  assign n97 = ~n88 & n96 ;
  assign n98 = x_pad & n30 ;
  assign n99 = q_pad & ~y_pad ;
  assign n100 = ~n98 & n99 ;
  assign n101 = q_pad & y_pad ;
  assign n102 = n98 & n101 ;
  assign n103 = ~n100 & ~n102 ;
  assign n104 = n37 & ~n103 ;
  assign n105 = ~y_pad & ~n98 ;
  assign n106 = x_pad & y_pad ;
  assign n107 = n30 & n106 ;
  assign n108 = n35 & ~n107 ;
  assign n109 = ~n105 & n108 ;
  assign n110 = ~n43 & ~n109 ;
  assign n111 = ~n104 & n110 ;
  assign n112 = ~z_pad & ~n107 ;
  assign n113 = ~n33 & n35 ;
  assign n114 = ~n112 & n113 ;
  assign n115 = \a0_pad  & r_pad ;
  assign n116 = n35 & n115 ;
  assign n117 = n33 & n116 ;
  assign n118 = ~n44 & ~n117 ;
  assign n119 = ~n114 & n118 ;
  assign n120 = \a0_pad  & ~s_pad ;
  assign n121 = n33 & n120 ;
  assign n122 = ~\a0_pad  & ~n33 ;
  assign n123 = n35 & ~n122 ;
  assign n124 = ~n121 & n123 ;
  assign n125 = ~n45 & ~n124 ;
  assign \b0_pad  = n37 ;
  assign \c0_pad  = n38 ;
  assign \d0_pad  = n39 ;
  assign \e0_pad  = n40 ;
  assign \f0_pad  = n41 ;
  assign \g0_pad  = n42 ;
  assign \h0_pad  = n43 ;
  assign \i0_pad  = n44 ;
  assign \j0_pad  = n45 ;
  assign \k0_pad  = ~n52 ;
  assign \l0_pad  = ~n59 ;
  assign \m0_pad  = ~n71 ;
  assign \n0_pad  = ~n82 ;
  assign \o0_pad  = ~n97 ;
  assign \p0_pad  = ~n111 ;
  assign \q0_pad  = ~n119 ;
  assign \r0_pad  = ~n125 ;
endmodule
