module top( \a0_pad  , a_pad , \b0_pad  , \c0_pad  , c_pad , \d0_pad  , d_pad , \e0_pad  , e_pad , \f0_pad  , f_pad , \g0_pad  , g_pad , \h0_pad  , h_pad , \i0_pad  , i_pad , \j0_pad  , j_pad , \k0_pad  , k_pad , \l0_pad  , l_pad , \m0_pad  , m_pad , \n0_pad  , n_pad , \o0_pad  , o_pad , \p0_pad  , p_pad , \q0_pad  , q_pad , \r0_pad  , r_pad , \s0_pad  , s_pad , \t0_pad  , t_pad , \u0_pad  , u_pad , \v0_pad  , v_pad , w_pad , x_pad , y_pad , z_pad , \a1_pad  , \a2_pad  , \b1_pad  , \b2_pad  , \c1_pad  , \c2_pad  , \d1_pad  , \d2_pad  , \e1_pad  , \e2_pad  , \f1_pad  , \f2_pad  , \g1_pad  , \h1_pad  , \i1_pad  , \j1_pad  , \k1_pad  , \l1_pad  , \m1_pad  , \n1_pad  , \o1_pad  , \p1_pad  , \q1_pad  , \r1_pad  , \s1_pad  , \t1_pad  , \u1_pad  , \v1_pad  , \w0_pad  , \w1_pad  , \x0_pad  , \x1_pad  , \y0_pad  , \y1_pad  , \z0_pad  , \z1_pad  );
  input \a0_pad  ;
  input a_pad ;
  input \b0_pad  ;
  input \c0_pad  ;
  input c_pad ;
  input \d0_pad  ;
  input d_pad ;
  input \e0_pad  ;
  input e_pad ;
  input \f0_pad  ;
  input f_pad ;
  input \g0_pad  ;
  input g_pad ;
  input \h0_pad  ;
  input h_pad ;
  input \i0_pad  ;
  input i_pad ;
  input \j0_pad  ;
  input j_pad ;
  input \k0_pad  ;
  input k_pad ;
  input \l0_pad  ;
  input l_pad ;
  input \m0_pad  ;
  input m_pad ;
  input \n0_pad  ;
  input n_pad ;
  input \o0_pad  ;
  input o_pad ;
  input \p0_pad  ;
  input p_pad ;
  input \q0_pad  ;
  input q_pad ;
  input \r0_pad  ;
  input r_pad ;
  input \s0_pad  ;
  input s_pad ;
  input \t0_pad  ;
  input t_pad ;
  input \u0_pad  ;
  input u_pad ;
  input \v0_pad  ;
  input v_pad ;
  input w_pad ;
  input x_pad ;
  input y_pad ;
  input z_pad ;
  output \a1_pad  ;
  output \a2_pad  ;
  output \b1_pad  ;
  output \b2_pad  ;
  output \c1_pad  ;
  output \c2_pad  ;
  output \d1_pad  ;
  output \d2_pad  ;
  output \e1_pad  ;
  output \e2_pad  ;
  output \f1_pad  ;
  output \f2_pad  ;
  output \g1_pad  ;
  output \h1_pad  ;
  output \i1_pad  ;
  output \j1_pad  ;
  output \k1_pad  ;
  output \l1_pad  ;
  output \m1_pad  ;
  output \n1_pad  ;
  output \o1_pad  ;
  output \p1_pad  ;
  output \q1_pad  ;
  output \r1_pad  ;
  output \s1_pad  ;
  output \t1_pad  ;
  output \u1_pad  ;
  output \v1_pad  ;
  output \w0_pad  ;
  output \w1_pad  ;
  output \x0_pad  ;
  output \x1_pad  ;
  output \y0_pad  ;
  output \y1_pad  ;
  output \z0_pad  ;
  output \z1_pad  ;
  wire n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 ;
  assign n49 = ~d_pad & i_pad ;
  assign n48 = ~i_pad & ~q_pad ;
  assign n50 = ~l_pad & ~n48 ;
  assign n51 = ~n49 & n50 ;
  assign n52 = k_pad & ~p_pad ;
  assign n54 = ~\r0_pad  & n52 ;
  assign n53 = ~\q0_pad  & ~n52 ;
  assign n55 = ~l_pad & ~n53 ;
  assign n56 = ~n54 & n55 ;
  assign n58 = ~e_pad & i_pad ;
  assign n57 = ~i_pad & ~r_pad ;
  assign n59 = ~l_pad & ~n57 ;
  assign n60 = ~n58 & n59 ;
  assign n62 = ~\s0_pad  & n52 ;
  assign n61 = ~\r0_pad  & ~n52 ;
  assign n63 = ~l_pad & ~n61 ;
  assign n64 = ~n62 & n63 ;
  assign n66 = j_pad & ~t_pad ;
  assign n65 = ~j_pad & ~s_pad ;
  assign n67 = ~l_pad & ~n65 ;
  assign n68 = ~n66 & n67 ;
  assign n70 = ~\t0_pad  & n52 ;
  assign n69 = ~\s0_pad  & ~n52 ;
  assign n71 = ~l_pad & ~n69 ;
  assign n72 = ~n70 & n71 ;
  assign n74 = j_pad & ~u_pad ;
  assign n73 = ~j_pad & ~t_pad ;
  assign n75 = ~l_pad & ~n73 ;
  assign n76 = ~n74 & n75 ;
  assign n78 = ~\u0_pad  & n52 ;
  assign n77 = ~\t0_pad  & ~n52 ;
  assign n79 = ~l_pad & ~n77 ;
  assign n80 = ~n78 & n79 ;
  assign n82 = j_pad & ~v_pad ;
  assign n81 = ~j_pad & ~u_pad ;
  assign n83 = ~l_pad & ~n81 ;
  assign n84 = ~n82 & n83 ;
  assign n86 = ~\v0_pad  & n52 ;
  assign n85 = ~\u0_pad  & ~n52 ;
  assign n87 = ~l_pad & ~n85 ;
  assign n88 = ~n86 & n87 ;
  assign n90 = j_pad & ~w_pad ;
  assign n89 = ~j_pad & ~v_pad ;
  assign n91 = ~l_pad & ~n89 ;
  assign n92 = ~n90 & n91 ;
  assign n94 = ~a_pad & n52 ;
  assign n93 = ~\v0_pad  & ~n52 ;
  assign n95 = ~l_pad & ~n93 ;
  assign n96 = ~n94 & n95 ;
  assign n98 = j_pad & ~x_pad ;
  assign n97 = ~j_pad & ~w_pad ;
  assign n99 = ~l_pad & ~n97 ;
  assign n100 = ~n98 & n99 ;
  assign n102 = j_pad & ~y_pad ;
  assign n101 = ~j_pad & ~x_pad ;
  assign n103 = ~l_pad & ~n101 ;
  assign n104 = ~n102 & n103 ;
  assign n106 = j_pad & ~z_pad ;
  assign n105 = ~j_pad & ~y_pad ;
  assign n107 = ~l_pad & ~n105 ;
  assign n108 = ~n106 & n107 ;
  assign n110 = ~\a0_pad  & j_pad ;
  assign n109 = ~j_pad & ~z_pad ;
  assign n111 = ~l_pad & ~n109 ;
  assign n112 = ~n110 & n111 ;
  assign n114 = ~\b0_pad  & j_pad ;
  assign n113 = ~\a0_pad  & ~j_pad ;
  assign n115 = ~l_pad & ~n113 ;
  assign n116 = ~n114 & n115 ;
  assign n118 = ~\c0_pad  & j_pad ;
  assign n117 = ~\b0_pad  & ~j_pad ;
  assign n119 = ~l_pad & ~n117 ;
  assign n120 = ~n118 & n119 ;
  assign n122 = ~\d0_pad  & j_pad ;
  assign n121 = ~\c0_pad  & ~j_pad ;
  assign n123 = ~l_pad & ~n121 ;
  assign n124 = ~n122 & n123 ;
  assign n126 = ~\e0_pad  & j_pad ;
  assign n125 = ~\d0_pad  & ~j_pad ;
  assign n127 = ~l_pad & ~n125 ;
  assign n128 = ~n126 & n127 ;
  assign n130 = ~\f0_pad  & j_pad ;
  assign n129 = ~\e0_pad  & ~j_pad ;
  assign n131 = ~l_pad & ~n129 ;
  assign n132 = ~n130 & n131 ;
  assign n134 = ~a_pad & j_pad ;
  assign n133 = ~\f0_pad  & ~j_pad ;
  assign n135 = ~l_pad & ~n133 ;
  assign n136 = ~n134 & n135 ;
  assign n138 = ~\h0_pad  & k_pad ;
  assign n137 = ~\g0_pad  & ~k_pad ;
  assign n139 = ~l_pad & ~n137 ;
  assign n140 = ~n138 & n139 ;
  assign n142 = ~\i0_pad  & k_pad ;
  assign n141 = ~\h0_pad  & ~k_pad ;
  assign n143 = ~l_pad & ~n141 ;
  assign n144 = ~n142 & n143 ;
  assign n146 = ~\j0_pad  & k_pad ;
  assign n145 = ~\i0_pad  & ~k_pad ;
  assign n147 = ~l_pad & ~n145 ;
  assign n148 = ~n146 & n147 ;
  assign n150 = ~\k0_pad  & k_pad ;
  assign n149 = ~\j0_pad  & ~k_pad ;
  assign n151 = ~l_pad & ~n149 ;
  assign n152 = ~n150 & n151 ;
  assign n154 = k_pad & ~\l0_pad  ;
  assign n153 = ~\k0_pad  & ~k_pad ;
  assign n155 = ~l_pad & ~n153 ;
  assign n156 = ~n154 & n155 ;
  assign n158 = k_pad & ~\m0_pad  ;
  assign n157 = ~k_pad & ~\l0_pad  ;
  assign n159 = ~l_pad & ~n157 ;
  assign n160 = ~n158 & n159 ;
  assign n162 = ~f_pad & i_pad ;
  assign n161 = ~i_pad & ~m_pad ;
  assign n163 = ~l_pad & ~n161 ;
  assign n164 = ~n162 & n163 ;
  assign n166 = k_pad & ~\n0_pad  ;
  assign n165 = ~k_pad & ~\m0_pad  ;
  assign n167 = ~l_pad & ~n165 ;
  assign n168 = ~n166 & n167 ;
  assign n170 = ~g_pad & i_pad ;
  assign n169 = ~i_pad & ~n_pad ;
  assign n171 = ~l_pad & ~n169 ;
  assign n172 = ~n170 & n171 ;
  assign n175 = a_pad & p_pad ;
  assign n174 = \o0_pad  & ~p_pad ;
  assign n176 = k_pad & ~n174 ;
  assign n177 = ~n175 & n176 ;
  assign n173 = ~k_pad & ~\n0_pad  ;
  assign n178 = ~l_pad & ~n173 ;
  assign n179 = ~n177 & n178 ;
  assign n181 = ~h_pad & i_pad ;
  assign n180 = ~i_pad & ~o_pad ;
  assign n182 = ~l_pad & ~n180 ;
  assign n183 = ~n181 & n182 ;
  assign n185 = ~\p0_pad  & n52 ;
  assign n184 = ~\o0_pad  & ~n52 ;
  assign n186 = ~l_pad & ~n184 ;
  assign n187 = ~n185 & n186 ;
  assign n189 = ~c_pad & i_pad ;
  assign n188 = ~i_pad & ~p_pad ;
  assign n190 = ~l_pad & ~n188 ;
  assign n191 = ~n189 & n190 ;
  assign n193 = ~\q0_pad  & n52 ;
  assign n192 = ~\p0_pad  & ~n52 ;
  assign n194 = ~l_pad & ~n192 ;
  assign n195 = ~n193 & n194 ;
  assign \a1_pad  = n51 ;
  assign \a2_pad  = n56 ;
  assign \b1_pad  = n60 ;
  assign \b2_pad  = n64 ;
  assign \c1_pad  = n68 ;
  assign \c2_pad  = n72 ;
  assign \d1_pad  = n76 ;
  assign \d2_pad  = n80 ;
  assign \e1_pad  = n84 ;
  assign \e2_pad  = n88 ;
  assign \f1_pad  = n92 ;
  assign \f2_pad  = n96 ;
  assign \g1_pad  = n100 ;
  assign \h1_pad  = n104 ;
  assign \i1_pad  = n108 ;
  assign \j1_pad  = n112 ;
  assign \k1_pad  = n116 ;
  assign \l1_pad  = n120 ;
  assign \m1_pad  = n124 ;
  assign \n1_pad  = n128 ;
  assign \o1_pad  = n132 ;
  assign \p1_pad  = n136 ;
  assign \q1_pad  = n140 ;
  assign \r1_pad  = n144 ;
  assign \s1_pad  = n148 ;
  assign \t1_pad  = n152 ;
  assign \u1_pad  = n156 ;
  assign \v1_pad  = n160 ;
  assign \w0_pad  = n164 ;
  assign \w1_pad  = n168 ;
  assign \x0_pad  = n172 ;
  assign \x1_pad  = n179 ;
  assign \y0_pad  = n183 ;
  assign \y1_pad  = n187 ;
  assign \z0_pad  = n191 ;
  assign \z1_pad  = n195 ;
endmodule
