module top (CLR_pad, \v0_pad , \v10_reg/NET0131 , \v11_reg/NET0131 , \v12_reg/NET0131 , \v1_pad , \v2_pad , \v3_pad , \v4_pad , \v5_pad , \v6_pad , \v7_reg/NET0131 , \v8_reg/NET0131 , \v9_reg/NET0131 , \_al_n0 , \_al_n1 , \g1757/_0_ , \g1763/_1_ , \g1787/_3_ , \g1800/_3_ , \g1821/_2_ , \g1940/_1_ , \g25/_0_ , \g2783/_3_ , \g2823/_0_ , \g38/_1_ , \g40/_1_ , \v13_D_11_pad , \v13_D_12_pad , \v13_D_13_pad , \v13_D_14_pad , \v13_D_16_pad , \v13_D_18_pad , \v13_D_19_pad , \v13_D_21_pad , \v13_D_22_pad , \v13_D_23_pad , \v13_D_24_pad , \v13_D_7_pad , \v13_D_8_pad , \v13_D_9_pad );
	input CLR_pad ;
	input \v0_pad  ;
	input \v10_reg/NET0131  ;
	input \v11_reg/NET0131  ;
	input \v12_reg/NET0131  ;
	input \v1_pad  ;
	input \v2_pad  ;
	input \v3_pad  ;
	input \v4_pad  ;
	input \v5_pad  ;
	input \v6_pad  ;
	input \v7_reg/NET0131  ;
	input \v8_reg/NET0131  ;
	input \v9_reg/NET0131  ;
	output \_al_n0  ;
	output \_al_n1  ;
	output \g1757/_0_  ;
	output \g1763/_1_  ;
	output \g1787/_3_  ;
	output \g1800/_3_  ;
	output \g1821/_2_  ;
	output \g1940/_1_  ;
	output \g25/_0_  ;
	output \g2783/_3_  ;
	output \g2823/_0_  ;
	output \g38/_1_  ;
	output \g40/_1_  ;
	output \v13_D_11_pad  ;
	output \v13_D_12_pad  ;
	output \v13_D_13_pad  ;
	output \v13_D_14_pad  ;
	output \v13_D_16_pad  ;
	output \v13_D_18_pad  ;
	output \v13_D_19_pad  ;
	output \v13_D_21_pad  ;
	output \v13_D_22_pad  ;
	output \v13_D_23_pad  ;
	output \v13_D_24_pad  ;
	output \v13_D_7_pad  ;
	output \v13_D_8_pad  ;
	output \v13_D_9_pad  ;
	wire _w579_ ;
	wire _w578_ ;
	wire _w577_ ;
	wire _w576_ ;
	wire _w575_ ;
	wire _w574_ ;
	wire _w573_ ;
	wire _w572_ ;
	wire _w571_ ;
	wire _w570_ ;
	wire _w569_ ;
	wire _w568_ ;
	wire _w567_ ;
	wire _w566_ ;
	wire _w565_ ;
	wire _w564_ ;
	wire _w563_ ;
	wire _w562_ ;
	wire _w561_ ;
	wire _w560_ ;
	wire _w559_ ;
	wire _w558_ ;
	wire _w557_ ;
	wire _w556_ ;
	wire _w271_ ;
	wire _w270_ ;
	wire _w269_ ;
	wire _w268_ ;
	wire _w267_ ;
	wire _w266_ ;
	wire _w265_ ;
	wire _w264_ ;
	wire _w263_ ;
	wire _w262_ ;
	wire _w261_ ;
	wire _w260_ ;
	wire _w259_ ;
	wire _w258_ ;
	wire _w257_ ;
	wire _w256_ ;
	wire _w255_ ;
	wire _w254_ ;
	wire _w253_ ;
	wire _w252_ ;
	wire _w251_ ;
	wire _w250_ ;
	wire _w249_ ;
	wire _w248_ ;
	wire _w247_ ;
	wire _w246_ ;
	wire _w245_ ;
	wire _w244_ ;
	wire _w243_ ;
	wire _w242_ ;
	wire _w241_ ;
	wire _w240_ ;
	wire _w239_ ;
	wire _w238_ ;
	wire _w237_ ;
	wire _w236_ ;
	wire _w235_ ;
	wire _w234_ ;
	wire _w233_ ;
	wire _w232_ ;
	wire _w231_ ;
	wire _w230_ ;
	wire _w229_ ;
	wire _w228_ ;
	wire _w227_ ;
	wire _w226_ ;
	wire _w225_ ;
	wire _w224_ ;
	wire _w223_ ;
	wire _w222_ ;
	wire _w221_ ;
	wire _w220_ ;
	wire _w219_ ;
	wire _w218_ ;
	wire _w217_ ;
	wire _w216_ ;
	wire _w215_ ;
	wire _w214_ ;
	wire _w213_ ;
	wire _w212_ ;
	wire _w211_ ;
	wire _w210_ ;
	wire _w209_ ;
	wire _w208_ ;
	wire _w207_ ;
	wire _w206_ ;
	wire _w205_ ;
	wire _w204_ ;
	wire _w203_ ;
	wire _w202_ ;
	wire _w201_ ;
	wire _w200_ ;
	wire _w199_ ;
	wire _w198_ ;
	wire _w197_ ;
	wire _w196_ ;
	wire _w195_ ;
	wire _w194_ ;
	wire _w193_ ;
	wire _w192_ ;
	wire _w191_ ;
	wire _w190_ ;
	wire _w189_ ;
	wire _w188_ ;
	wire _w187_ ;
	wire _w186_ ;
	wire _w185_ ;
	wire _w184_ ;
	wire _w183_ ;
	wire _w182_ ;
	wire _w181_ ;
	wire _w180_ ;
	wire _w179_ ;
	wire _w178_ ;
	wire _w177_ ;
	wire _w176_ ;
	wire _w175_ ;
	wire _w174_ ;
	wire _w173_ ;
	wire _w172_ ;
	wire _w171_ ;
	wire _w170_ ;
	wire _w169_ ;
	wire _w168_ ;
	wire _w167_ ;
	wire _w166_ ;
	wire _w165_ ;
	wire _w164_ ;
	wire _w163_ ;
	wire _w162_ ;
	wire _w161_ ;
	wire _w160_ ;
	wire _w159_ ;
	wire _w158_ ;
	wire _w157_ ;
	wire _w156_ ;
	wire _w155_ ;
	wire _w154_ ;
	wire _w153_ ;
	wire _w152_ ;
	wire _w151_ ;
	wire _w150_ ;
	wire _w149_ ;
	wire _w148_ ;
	wire _w147_ ;
	wire _w146_ ;
	wire _w145_ ;
	wire _w144_ ;
	wire _w143_ ;
	wire _w142_ ;
	wire _w73_ ;
	wire _w72_ ;
	wire _w71_ ;
	wire _w70_ ;
	wire _w69_ ;
	wire _w68_ ;
	wire _w67_ ;
	wire _w66_ ;
	wire _w65_ ;
	wire _w64_ ;
	wire _w63_ ;
	wire _w62_ ;
	wire _w61_ ;
	wire _w60_ ;
	wire _w59_ ;
	wire _w58_ ;
	wire _w57_ ;
	wire _w56_ ;
	wire _w55_ ;
	wire _w54_ ;
	wire _w53_ ;
	wire _w52_ ;
	wire _w51_ ;
	wire _w50_ ;
	wire _w49_ ;
	wire _w48_ ;
	wire _w47_ ;
	wire _w46_ ;
	wire _w45_ ;
	wire _w44_ ;
	wire _w27_ ;
	wire _w26_ ;
	wire _w25_ ;
	wire _w24_ ;
	wire _w23_ ;
	wire _w22_ ;
	wire _w21_ ;
	wire _w20_ ;
	wire _w19_ ;
	wire _w18_ ;
	wire _w17_ ;
	wire _w16_ ;
	wire _w15_ ;
	wire _w28_ ;
	wire _w29_ ;
	wire _w30_ ;
	wire _w31_ ;
	wire _w32_ ;
	wire _w33_ ;
	wire _w34_ ;
	wire _w35_ ;
	wire _w36_ ;
	wire _w37_ ;
	wire _w38_ ;
	wire _w39_ ;
	wire _w40_ ;
	wire _w41_ ;
	wire _w42_ ;
	wire _w43_ ;
	wire _w74_ ;
	wire _w75_ ;
	wire _w76_ ;
	wire _w77_ ;
	wire _w78_ ;
	wire _w79_ ;
	wire _w80_ ;
	wire _w81_ ;
	wire _w82_ ;
	wire _w83_ ;
	wire _w84_ ;
	wire _w85_ ;
	wire _w86_ ;
	wire _w87_ ;
	wire _w88_ ;
	wire _w89_ ;
	wire _w90_ ;
	wire _w91_ ;
	wire _w92_ ;
	wire _w93_ ;
	wire _w94_ ;
	wire _w95_ ;
	wire _w96_ ;
	wire _w97_ ;
	wire _w98_ ;
	wire _w99_ ;
	wire _w100_ ;
	wire _w101_ ;
	wire _w102_ ;
	wire _w103_ ;
	wire _w104_ ;
	wire _w105_ ;
	wire _w106_ ;
	wire _w107_ ;
	wire _w108_ ;
	wire _w109_ ;
	wire _w110_ ;
	wire _w111_ ;
	wire _w112_ ;
	wire _w113_ ;
	wire _w114_ ;
	wire _w115_ ;
	wire _w116_ ;
	wire _w117_ ;
	wire _w118_ ;
	wire _w119_ ;
	wire _w120_ ;
	wire _w121_ ;
	wire _w122_ ;
	wire _w123_ ;
	wire _w124_ ;
	wire _w125_ ;
	wire _w126_ ;
	wire _w127_ ;
	wire _w128_ ;
	wire _w129_ ;
	wire _w130_ ;
	wire _w131_ ;
	wire _w132_ ;
	wire _w133_ ;
	wire _w134_ ;
	wire _w135_ ;
	wire _w136_ ;
	wire _w137_ ;
	wire _w138_ ;
	wire _w139_ ;
	wire _w140_ ;
	wire _w141_ ;
	wire _w272_ ;
	wire _w273_ ;
	wire _w274_ ;
	wire _w275_ ;
	wire _w276_ ;
	wire _w277_ ;
	wire _w278_ ;
	wire _w279_ ;
	wire _w280_ ;
	wire _w281_ ;
	wire _w282_ ;
	wire _w283_ ;
	wire _w284_ ;
	wire _w285_ ;
	wire _w286_ ;
	wire _w287_ ;
	wire _w288_ ;
	wire _w289_ ;
	wire _w290_ ;
	wire _w291_ ;
	wire _w292_ ;
	wire _w293_ ;
	wire _w294_ ;
	wire _w295_ ;
	wire _w296_ ;
	wire _w297_ ;
	wire _w298_ ;
	wire _w299_ ;
	wire _w300_ ;
	wire _w301_ ;
	wire _w302_ ;
	wire _w303_ ;
	wire _w304_ ;
	wire _w305_ ;
	wire _w306_ ;
	wire _w307_ ;
	wire _w308_ ;
	wire _w309_ ;
	wire _w310_ ;
	wire _w311_ ;
	wire _w312_ ;
	wire _w313_ ;
	wire _w314_ ;
	wire _w315_ ;
	wire _w316_ ;
	wire _w317_ ;
	wire _w318_ ;
	wire _w319_ ;
	wire _w320_ ;
	wire _w321_ ;
	wire _w322_ ;
	wire _w323_ ;
	wire _w324_ ;
	wire _w325_ ;
	wire _w326_ ;
	wire _w327_ ;
	wire _w328_ ;
	wire _w329_ ;
	wire _w330_ ;
	wire _w331_ ;
	wire _w332_ ;
	wire _w333_ ;
	wire _w334_ ;
	wire _w335_ ;
	wire _w336_ ;
	wire _w337_ ;
	wire _w338_ ;
	wire _w339_ ;
	wire _w340_ ;
	wire _w341_ ;
	wire _w342_ ;
	wire _w343_ ;
	wire _w344_ ;
	wire _w345_ ;
	wire _w346_ ;
	wire _w347_ ;
	wire _w348_ ;
	wire _w349_ ;
	wire _w350_ ;
	wire _w351_ ;
	wire _w352_ ;
	wire _w353_ ;
	wire _w354_ ;
	wire _w355_ ;
	wire _w356_ ;
	wire _w357_ ;
	wire _w358_ ;
	wire _w359_ ;
	wire _w360_ ;
	wire _w361_ ;
	wire _w362_ ;
	wire _w363_ ;
	wire _w364_ ;
	wire _w365_ ;
	wire _w366_ ;
	wire _w367_ ;
	wire _w368_ ;
	wire _w369_ ;
	wire _w370_ ;
	wire _w371_ ;
	wire _w372_ ;
	wire _w373_ ;
	wire _w374_ ;
	wire _w375_ ;
	wire _w376_ ;
	wire _w377_ ;
	wire _w378_ ;
	wire _w379_ ;
	wire _w380_ ;
	wire _w381_ ;
	wire _w382_ ;
	wire _w383_ ;
	wire _w384_ ;
	wire _w385_ ;
	wire _w386_ ;
	wire _w387_ ;
	wire _w388_ ;
	wire _w389_ ;
	wire _w390_ ;
	wire _w391_ ;
	wire _w392_ ;
	wire _w393_ ;
	wire _w394_ ;
	wire _w395_ ;
	wire _w396_ ;
	wire _w397_ ;
	wire _w398_ ;
	wire _w399_ ;
	wire _w400_ ;
	wire _w401_ ;
	wire _w402_ ;
	wire _w403_ ;
	wire _w404_ ;
	wire _w405_ ;
	wire _w406_ ;
	wire _w407_ ;
	wire _w408_ ;
	wire _w409_ ;
	wire _w410_ ;
	wire _w411_ ;
	wire _w412_ ;
	wire _w413_ ;
	wire _w414_ ;
	wire _w415_ ;
	wire _w416_ ;
	wire _w417_ ;
	wire _w418_ ;
	wire _w419_ ;
	wire _w420_ ;
	wire _w421_ ;
	wire _w422_ ;
	wire _w423_ ;
	wire _w424_ ;
	wire _w425_ ;
	wire _w426_ ;
	wire _w427_ ;
	wire _w428_ ;
	wire _w429_ ;
	wire _w430_ ;
	wire _w431_ ;
	wire _w432_ ;
	wire _w433_ ;
	wire _w434_ ;
	wire _w435_ ;
	wire _w436_ ;
	wire _w437_ ;
	wire _w438_ ;
	wire _w439_ ;
	wire _w440_ ;
	wire _w441_ ;
	wire _w442_ ;
	wire _w443_ ;
	wire _w444_ ;
	wire _w445_ ;
	wire _w446_ ;
	wire _w447_ ;
	wire _w448_ ;
	wire _w449_ ;
	wire _w450_ ;
	wire _w451_ ;
	wire _w452_ ;
	wire _w453_ ;
	wire _w454_ ;
	wire _w455_ ;
	wire _w456_ ;
	wire _w457_ ;
	wire _w458_ ;
	wire _w459_ ;
	wire _w460_ ;
	wire _w461_ ;
	wire _w462_ ;
	wire _w463_ ;
	wire _w464_ ;
	wire _w465_ ;
	wire _w466_ ;
	wire _w467_ ;
	wire _w468_ ;
	wire _w469_ ;
	wire _w470_ ;
	wire _w471_ ;
	wire _w472_ ;
	wire _w473_ ;
	wire _w474_ ;
	wire _w475_ ;
	wire _w476_ ;
	wire _w477_ ;
	wire _w478_ ;
	wire _w479_ ;
	wire _w480_ ;
	wire _w481_ ;
	wire _w482_ ;
	wire _w483_ ;
	wire _w484_ ;
	wire _w485_ ;
	wire _w486_ ;
	wire _w487_ ;
	wire _w488_ ;
	wire _w489_ ;
	wire _w490_ ;
	wire _w491_ ;
	wire _w492_ ;
	wire _w493_ ;
	wire _w494_ ;
	wire _w495_ ;
	wire _w496_ ;
	wire _w497_ ;
	wire _w498_ ;
	wire _w499_ ;
	wire _w500_ ;
	wire _w501_ ;
	wire _w502_ ;
	wire _w503_ ;
	wire _w504_ ;
	wire _w505_ ;
	wire _w506_ ;
	wire _w507_ ;
	wire _w508_ ;
	wire _w509_ ;
	wire _w510_ ;
	wire _w511_ ;
	wire _w512_ ;
	wire _w513_ ;
	wire _w514_ ;
	wire _w515_ ;
	wire _w516_ ;
	wire _w517_ ;
	wire _w518_ ;
	wire _w519_ ;
	wire _w520_ ;
	wire _w521_ ;
	wire _w522_ ;
	wire _w523_ ;
	wire _w524_ ;
	wire _w525_ ;
	wire _w526_ ;
	wire _w527_ ;
	wire _w528_ ;
	wire _w529_ ;
	wire _w530_ ;
	wire _w531_ ;
	wire _w532_ ;
	wire _w533_ ;
	wire _w534_ ;
	wire _w535_ ;
	wire _w536_ ;
	wire _w537_ ;
	wire _w538_ ;
	wire _w539_ ;
	wire _w540_ ;
	wire _w541_ ;
	wire _w542_ ;
	wire _w543_ ;
	wire _w544_ ;
	wire _w545_ ;
	wire _w546_ ;
	wire _w547_ ;
	wire _w548_ ;
	wire _w549_ ;
	wire _w550_ ;
	wire _w551_ ;
	wire _w552_ ;
	wire _w553_ ;
	wire _w554_ ;
	wire _w555_ ;
	LUT2 #(
		.INIT('h2)
	) name0 (
		\v10_reg/NET0131 ,
		\v12_reg/NET0131 ,
		_w15_
	);
	LUT2 #(
		.INIT('h4)
	) name1 (
		\v11_reg/NET0131 ,
		_w15_,
		_w16_
	);
	LUT2 #(
		.INIT('h2)
	) name2 (
		\v9_reg/NET0131 ,
		_w16_,
		_w17_
	);
	LUT2 #(
		.INIT('h8)
	) name3 (
		\v10_reg/NET0131 ,
		\v11_reg/NET0131 ,
		_w18_
	);
	LUT2 #(
		.INIT('h4)
	) name4 (
		\v0_pad ,
		_w18_,
		_w19_
	);
	LUT2 #(
		.INIT('h1)
	) name5 (
		\v10_reg/NET0131 ,
		\v11_reg/NET0131 ,
		_w20_
	);
	LUT2 #(
		.INIT('h1)
	) name6 (
		_w19_,
		_w20_,
		_w21_
	);
	LUT2 #(
		.INIT('h8)
	) name7 (
		\v4_pad ,
		\v5_pad ,
		_w22_
	);
	LUT2 #(
		.INIT('h4)
	) name8 (
		\v12_reg/NET0131 ,
		_w22_,
		_w23_
	);
	LUT2 #(
		.INIT('h4)
	) name9 (
		_w21_,
		_w23_,
		_w24_
	);
	LUT2 #(
		.INIT('h4)
	) name10 (
		\v10_reg/NET0131 ,
		\v11_reg/NET0131 ,
		_w25_
	);
	LUT2 #(
		.INIT('h2)
	) name11 (
		\v10_reg/NET0131 ,
		\v11_reg/NET0131 ,
		_w26_
	);
	LUT2 #(
		.INIT('h1)
	) name12 (
		_w25_,
		_w26_,
		_w27_
	);
	LUT2 #(
		.INIT('h1)
	) name13 (
		\v10_reg/NET0131 ,
		\v3_pad ,
		_w28_
	);
	LUT2 #(
		.INIT('h4)
	) name14 (
		\v6_pad ,
		_w28_,
		_w29_
	);
	LUT2 #(
		.INIT('h2)
	) name15 (
		_w27_,
		_w29_,
		_w30_
	);
	LUT2 #(
		.INIT('h2)
	) name16 (
		\v12_reg/NET0131 ,
		_w30_,
		_w31_
	);
	LUT2 #(
		.INIT('h1)
	) name17 (
		_w17_,
		_w24_,
		_w32_
	);
	LUT2 #(
		.INIT('h4)
	) name18 (
		_w31_,
		_w32_,
		_w33_
	);
	LUT2 #(
		.INIT('h1)
	) name19 (
		\v8_reg/NET0131 ,
		_w33_,
		_w34_
	);
	LUT2 #(
		.INIT('h2)
	) name20 (
		\v12_reg/NET0131 ,
		\v3_pad ,
		_w35_
	);
	LUT2 #(
		.INIT('h2)
	) name21 (
		\v10_reg/NET0131 ,
		\v8_reg/NET0131 ,
		_w36_
	);
	LUT2 #(
		.INIT('h8)
	) name22 (
		_w35_,
		_w36_,
		_w37_
	);
	LUT2 #(
		.INIT('h4)
	) name23 (
		\v8_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w38_
	);
	LUT2 #(
		.INIT('h8)
	) name24 (
		\v11_reg/NET0131 ,
		\v12_reg/NET0131 ,
		_w39_
	);
	LUT2 #(
		.INIT('h1)
	) name25 (
		\v10_reg/NET0131 ,
		\v1_pad ,
		_w40_
	);
	LUT2 #(
		.INIT('h8)
	) name26 (
		_w39_,
		_w40_,
		_w41_
	);
	LUT2 #(
		.INIT('h1)
	) name27 (
		_w37_,
		_w38_,
		_w42_
	);
	LUT2 #(
		.INIT('h4)
	) name28 (
		_w41_,
		_w42_,
		_w43_
	);
	LUT2 #(
		.INIT('h2)
	) name29 (
		\v2_pad ,
		_w43_,
		_w44_
	);
	LUT2 #(
		.INIT('h8)
	) name30 (
		\v9_reg/NET0131 ,
		_w39_,
		_w45_
	);
	LUT2 #(
		.INIT('h4)
	) name31 (
		\v10_reg/NET0131 ,
		\v8_reg/NET0131 ,
		_w46_
	);
	LUT2 #(
		.INIT('h1)
	) name32 (
		\v12_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w47_
	);
	LUT2 #(
		.INIT('h8)
	) name33 (
		_w46_,
		_w47_,
		_w48_
	);
	LUT2 #(
		.INIT('h1)
	) name34 (
		_w45_,
		_w48_,
		_w49_
	);
	LUT2 #(
		.INIT('h4)
	) name35 (
		_w44_,
		_w49_,
		_w50_
	);
	LUT2 #(
		.INIT('h4)
	) name36 (
		_w34_,
		_w50_,
		_w51_
	);
	LUT2 #(
		.INIT('h1)
	) name37 (
		\v7_reg/NET0131 ,
		_w51_,
		_w52_
	);
	LUT2 #(
		.INIT('h4)
	) name38 (
		\v2_pad ,
		\v8_reg/NET0131 ,
		_w53_
	);
	LUT2 #(
		.INIT('h2)
	) name39 (
		\v12_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w54_
	);
	LUT2 #(
		.INIT('h8)
	) name40 (
		\v7_reg/NET0131 ,
		_w54_,
		_w55_
	);
	LUT2 #(
		.INIT('h8)
	) name41 (
		\v11_reg/NET0131 ,
		_w15_,
		_w56_
	);
	LUT2 #(
		.INIT('h1)
	) name42 (
		_w55_,
		_w56_,
		_w57_
	);
	LUT2 #(
		.INIT('h2)
	) name43 (
		_w53_,
		_w57_,
		_w58_
	);
	LUT2 #(
		.INIT('h1)
	) name44 (
		\v10_reg/NET0131 ,
		\v12_reg/NET0131 ,
		_w59_
	);
	LUT2 #(
		.INIT('h8)
	) name45 (
		\v3_pad ,
		_w59_,
		_w60_
	);
	LUT2 #(
		.INIT('h1)
	) name46 (
		_w54_,
		_w60_,
		_w61_
	);
	LUT2 #(
		.INIT('h4)
	) name47 (
		\v11_reg/NET0131 ,
		\v8_reg/NET0131 ,
		_w62_
	);
	LUT2 #(
		.INIT('h4)
	) name48 (
		_w61_,
		_w62_,
		_w63_
	);
	LUT2 #(
		.INIT('h8)
	) name49 (
		\v12_reg/NET0131 ,
		\v1_pad ,
		_w64_
	);
	LUT2 #(
		.INIT('h4)
	) name50 (
		\v10_reg/NET0131 ,
		_w64_,
		_w65_
	);
	LUT2 #(
		.INIT('h8)
	) name51 (
		\v8_reg/NET0131 ,
		_w23_,
		_w66_
	);
	LUT2 #(
		.INIT('h1)
	) name52 (
		_w65_,
		_w66_,
		_w67_
	);
	LUT2 #(
		.INIT('h2)
	) name53 (
		\v11_reg/NET0131 ,
		\v2_pad ,
		_w68_
	);
	LUT2 #(
		.INIT('h4)
	) name54 (
		\v7_reg/NET0131 ,
		_w68_,
		_w69_
	);
	LUT2 #(
		.INIT('h4)
	) name55 (
		_w67_,
		_w69_,
		_w70_
	);
	LUT2 #(
		.INIT('h4)
	) name56 (
		\v12_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w71_
	);
	LUT2 #(
		.INIT('h8)
	) name57 (
		_w18_,
		_w71_,
		_w72_
	);
	LUT2 #(
		.INIT('h2)
	) name58 (
		\v11_reg/NET0131 ,
		_w54_,
		_w73_
	);
	LUT2 #(
		.INIT('h2)
	) name59 (
		_w46_,
		_w73_,
		_w74_
	);
	LUT2 #(
		.INIT('h2)
	) name60 (
		\v11_reg/NET0131 ,
		_w46_,
		_w75_
	);
	LUT2 #(
		.INIT('h1)
	) name61 (
		\v12_reg/NET0131 ,
		_w36_,
		_w76_
	);
	LUT2 #(
		.INIT('h8)
	) name62 (
		_w75_,
		_w76_,
		_w77_
	);
	LUT2 #(
		.INIT('h1)
	) name63 (
		_w72_,
		_w74_,
		_w78_
	);
	LUT2 #(
		.INIT('h4)
	) name64 (
		_w77_,
		_w78_,
		_w79_
	);
	LUT2 #(
		.INIT('h2)
	) name65 (
		\v7_reg/NET0131 ,
		_w79_,
		_w80_
	);
	LUT2 #(
		.INIT('h1)
	) name66 (
		_w58_,
		_w63_,
		_w81_
	);
	LUT2 #(
		.INIT('h4)
	) name67 (
		_w70_,
		_w81_,
		_w82_
	);
	LUT2 #(
		.INIT('h4)
	) name68 (
		_w80_,
		_w82_,
		_w83_
	);
	LUT2 #(
		.INIT('h4)
	) name69 (
		_w52_,
		_w83_,
		_w84_
	);
	LUT2 #(
		.INIT('h2)
	) name70 (
		CLR_pad,
		_w84_,
		_w85_
	);
	LUT2 #(
		.INIT('h1)
	) name71 (
		\v9_reg/NET0131 ,
		_w64_,
		_w86_
	);
	LUT2 #(
		.INIT('h8)
	) name72 (
		\v11_reg/NET0131 ,
		_w46_,
		_w87_
	);
	LUT2 #(
		.INIT('h4)
	) name73 (
		_w86_,
		_w87_,
		_w88_
	);
	LUT2 #(
		.INIT('h1)
	) name74 (
		\v11_reg/NET0131 ,
		\v8_reg/NET0131 ,
		_w89_
	);
	LUT2 #(
		.INIT('h8)
	) name75 (
		_w71_,
		_w89_,
		_w90_
	);
	LUT2 #(
		.INIT('h4)
	) name76 (
		\v10_reg/NET0131 ,
		_w90_,
		_w91_
	);
	LUT2 #(
		.INIT('h1)
	) name77 (
		_w88_,
		_w91_,
		_w92_
	);
	LUT2 #(
		.INIT('h2)
	) name78 (
		\v2_pad ,
		_w92_,
		_w93_
	);
	LUT2 #(
		.INIT('h8)
	) name79 (
		\v2_pad ,
		_w26_,
		_w94_
	);
	LUT2 #(
		.INIT('h4)
	) name80 (
		_w22_,
		_w36_,
		_w95_
	);
	LUT2 #(
		.INIT('h1)
	) name81 (
		_w94_,
		_w95_,
		_w96_
	);
	LUT2 #(
		.INIT('h2)
	) name82 (
		_w47_,
		_w96_,
		_w97_
	);
	LUT2 #(
		.INIT('h8)
	) name83 (
		\v12_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w98_
	);
	LUT2 #(
		.INIT('h8)
	) name84 (
		_w26_,
		_w98_,
		_w99_
	);
	LUT2 #(
		.INIT('h4)
	) name85 (
		\v11_reg/NET0131 ,
		\v3_pad ,
		_w100_
	);
	LUT2 #(
		.INIT('h4)
	) name86 (
		\v12_reg/NET0131 ,
		_w46_,
		_w101_
	);
	LUT2 #(
		.INIT('h8)
	) name87 (
		_w100_,
		_w101_,
		_w102_
	);
	LUT2 #(
		.INIT('h1)
	) name88 (
		\v11_reg/NET0131 ,
		\v6_pad ,
		_w103_
	);
	LUT2 #(
		.INIT('h1)
	) name89 (
		\v10_reg/NET0131 ,
		\v8_reg/NET0131 ,
		_w104_
	);
	LUT2 #(
		.INIT('h8)
	) name90 (
		_w71_,
		_w104_,
		_w105_
	);
	LUT2 #(
		.INIT('h8)
	) name91 (
		_w103_,
		_w105_,
		_w106_
	);
	LUT2 #(
		.INIT('h2)
	) name92 (
		\v9_reg/NET0131 ,
		_w22_,
		_w107_
	);
	LUT2 #(
		.INIT('h8)
	) name93 (
		_w87_,
		_w107_,
		_w108_
	);
	LUT2 #(
		.INIT('h8)
	) name94 (
		\v8_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w109_
	);
	LUT2 #(
		.INIT('h2)
	) name95 (
		\v12_reg/NET0131 ,
		_w18_,
		_w110_
	);
	LUT2 #(
		.INIT('h8)
	) name96 (
		_w109_,
		_w110_,
		_w111_
	);
	LUT2 #(
		.INIT('h1)
	) name97 (
		\v10_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w112_
	);
	LUT2 #(
		.INIT('h8)
	) name98 (
		_w23_,
		_w112_,
		_w113_
	);
	LUT2 #(
		.INIT('h4)
	) name99 (
		\v11_reg/NET0131 ,
		_w113_,
		_w114_
	);
	LUT2 #(
		.INIT('h8)
	) name100 (
		_w39_,
		_w53_,
		_w115_
	);
	LUT2 #(
		.INIT('h1)
	) name101 (
		_w90_,
		_w115_,
		_w116_
	);
	LUT2 #(
		.INIT('h2)
	) name102 (
		_w40_,
		_w116_,
		_w117_
	);
	LUT2 #(
		.INIT('h1)
	) name103 (
		\v8_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w118_
	);
	LUT2 #(
		.INIT('h8)
	) name104 (
		\v12_reg/NET0131 ,
		_w25_,
		_w119_
	);
	LUT2 #(
		.INIT('h4)
	) name105 (
		\v0_pad ,
		\v11_reg/NET0131 ,
		_w120_
	);
	LUT2 #(
		.INIT('h2)
	) name106 (
		_w15_,
		_w120_,
		_w121_
	);
	LUT2 #(
		.INIT('h1)
	) name107 (
		_w119_,
		_w121_,
		_w122_
	);
	LUT2 #(
		.INIT('h2)
	) name108 (
		_w118_,
		_w122_,
		_w123_
	);
	LUT2 #(
		.INIT('h1)
	) name109 (
		\v7_reg/NET0131 ,
		_w99_,
		_w124_
	);
	LUT2 #(
		.INIT('h4)
	) name110 (
		_w102_,
		_w124_,
		_w125_
	);
	LUT2 #(
		.INIT('h1)
	) name111 (
		_w106_,
		_w108_,
		_w126_
	);
	LUT2 #(
		.INIT('h4)
	) name112 (
		_w111_,
		_w126_,
		_w127_
	);
	LUT2 #(
		.INIT('h4)
	) name113 (
		_w97_,
		_w125_,
		_w128_
	);
	LUT2 #(
		.INIT('h1)
	) name114 (
		_w114_,
		_w117_,
		_w129_
	);
	LUT2 #(
		.INIT('h4)
	) name115 (
		_w123_,
		_w129_,
		_w130_
	);
	LUT2 #(
		.INIT('h8)
	) name116 (
		_w127_,
		_w128_,
		_w131_
	);
	LUT2 #(
		.INIT('h4)
	) name117 (
		_w93_,
		_w131_,
		_w132_
	);
	LUT2 #(
		.INIT('h8)
	) name118 (
		_w130_,
		_w132_,
		_w133_
	);
	LUT2 #(
		.INIT('h2)
	) name119 (
		\v11_reg/NET0131 ,
		\v12_reg/NET0131 ,
		_w134_
	);
	LUT2 #(
		.INIT('h2)
	) name120 (
		\v10_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w135_
	);
	LUT2 #(
		.INIT('h2)
	) name121 (
		_w134_,
		_w135_,
		_w136_
	);
	LUT2 #(
		.INIT('h2)
	) name122 (
		\v12_reg/NET0131 ,
		_w68_,
		_w137_
	);
	LUT2 #(
		.INIT('h8)
	) name123 (
		_w27_,
		_w137_,
		_w138_
	);
	LUT2 #(
		.INIT('h1)
	) name124 (
		\v12_reg/NET0131 ,
		_w20_,
		_w139_
	);
	LUT2 #(
		.INIT('h2)
	) name125 (
		\v9_reg/NET0131 ,
		_w139_,
		_w140_
	);
	LUT2 #(
		.INIT('h2)
	) name126 (
		\v8_reg/NET0131 ,
		_w138_,
		_w141_
	);
	LUT2 #(
		.INIT('h4)
	) name127 (
		_w140_,
		_w141_,
		_w142_
	);
	LUT2 #(
		.INIT('h2)
	) name128 (
		\v7_reg/NET0131 ,
		_w136_,
		_w143_
	);
	LUT2 #(
		.INIT('h4)
	) name129 (
		_w142_,
		_w143_,
		_w144_
	);
	LUT2 #(
		.INIT('h1)
	) name130 (
		_w133_,
		_w144_,
		_w145_
	);
	LUT2 #(
		.INIT('h8)
	) name131 (
		\v11_reg/NET0131 ,
		\v3_pad ,
		_w146_
	);
	LUT2 #(
		.INIT('h2)
	) name132 (
		_w48_,
		_w146_,
		_w147_
	);
	LUT2 #(
		.INIT('h4)
	) name133 (
		\v6_pad ,
		_w104_,
		_w148_
	);
	LUT2 #(
		.INIT('h1)
	) name134 (
		\v7_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w149_
	);
	LUT2 #(
		.INIT('h8)
	) name135 (
		_w35_,
		_w149_,
		_w150_
	);
	LUT2 #(
		.INIT('h8)
	) name136 (
		_w148_,
		_w150_,
		_w151_
	);
	LUT2 #(
		.INIT('h1)
	) name137 (
		_w147_,
		_w151_,
		_w152_
	);
	LUT2 #(
		.INIT('h4)
	) name138 (
		_w145_,
		_w152_,
		_w153_
	);
	LUT2 #(
		.INIT('h2)
	) name139 (
		CLR_pad,
		_w153_,
		_w154_
	);
	LUT2 #(
		.INIT('h1)
	) name140 (
		\v7_reg/NET0131 ,
		\v8_reg/NET0131 ,
		_w155_
	);
	LUT2 #(
		.INIT('h8)
	) name141 (
		_w114_,
		_w155_,
		_w156_
	);
	LUT2 #(
		.INIT('h8)
	) name142 (
		\v11_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w157_
	);
	LUT2 #(
		.INIT('h8)
	) name143 (
		\v0_pad ,
		\v11_reg/NET0131 ,
		_w158_
	);
	LUT2 #(
		.INIT('h2)
	) name144 (
		_w149_,
		_w158_,
		_w159_
	);
	LUT2 #(
		.INIT('h1)
	) name145 (
		_w157_,
		_w159_,
		_w160_
	);
	LUT2 #(
		.INIT('h2)
	) name146 (
		\v10_reg/NET0131 ,
		_w160_,
		_w161_
	);
	LUT2 #(
		.INIT('h2)
	) name147 (
		\v8_reg/NET0131 ,
		_w112_,
		_w162_
	);
	LUT2 #(
		.INIT('h8)
	) name148 (
		\v11_reg/NET0131 ,
		_w162_,
		_w163_
	);
	LUT2 #(
		.INIT('h1)
	) name149 (
		_w161_,
		_w163_,
		_w164_
	);
	LUT2 #(
		.INIT('h1)
	) name150 (
		\v12_reg/NET0131 ,
		_w164_,
		_w165_
	);
	LUT2 #(
		.INIT('h1)
	) name151 (
		\v8_reg/NET0131 ,
		_w25_,
		_w166_
	);
	LUT2 #(
		.INIT('h1)
	) name152 (
		\v12_reg/NET0131 ,
		_w166_,
		_w167_
	);
	LUT2 #(
		.INIT('h8)
	) name153 (
		\v11_reg/NET0131 ,
		_w135_,
		_w168_
	);
	LUT2 #(
		.INIT('h8)
	) name154 (
		\v8_reg/NET0131 ,
		_w168_,
		_w169_
	);
	LUT2 #(
		.INIT('h1)
	) name155 (
		_w167_,
		_w169_,
		_w170_
	);
	LUT2 #(
		.INIT('h2)
	) name156 (
		\v7_reg/NET0131 ,
		_w170_,
		_w171_
	);
	LUT2 #(
		.INIT('h1)
	) name157 (
		_w165_,
		_w171_,
		_w172_
	);
	LUT2 #(
		.INIT('h2)
	) name158 (
		\v2_pad ,
		_w172_,
		_w173_
	);
	LUT2 #(
		.INIT('h1)
	) name159 (
		_w156_,
		_w173_,
		_w174_
	);
	LUT2 #(
		.INIT('h4)
	) name160 (
		\v2_pad ,
		\v9_reg/NET0131 ,
		_w175_
	);
	LUT2 #(
		.INIT('h8)
	) name161 (
		\v11_reg/NET0131 ,
		_w175_,
		_w176_
	);
	LUT2 #(
		.INIT('h1)
	) name162 (
		_w94_,
		_w176_,
		_w177_
	);
	LUT2 #(
		.INIT('h1)
	) name163 (
		\v12_reg/NET0131 ,
		_w177_,
		_w178_
	);
	LUT2 #(
		.INIT('h2)
	) name164 (
		\v8_reg/NET0131 ,
		_w178_,
		_w179_
	);
	LUT2 #(
		.INIT('h2)
	) name165 (
		\v11_reg/NET0131 ,
		_w104_,
		_w180_
	);
	LUT2 #(
		.INIT('h4)
	) name166 (
		\v4_pad ,
		\v5_pad ,
		_w181_
	);
	LUT2 #(
		.INIT('h1)
	) name167 (
		\v10_reg/NET0131 ,
		_w181_,
		_w182_
	);
	LUT2 #(
		.INIT('h1)
	) name168 (
		\v9_reg/NET0131 ,
		_w182_,
		_w183_
	);
	LUT2 #(
		.INIT('h1)
	) name169 (
		_w180_,
		_w183_,
		_w184_
	);
	LUT2 #(
		.INIT('h1)
	) name170 (
		\v12_reg/NET0131 ,
		_w184_,
		_w185_
	);
	LUT2 #(
		.INIT('h8)
	) name171 (
		\v11_reg/NET0131 ,
		_w112_,
		_w186_
	);
	LUT2 #(
		.INIT('h1)
	) name172 (
		_w185_,
		_w186_,
		_w187_
	);
	LUT2 #(
		.INIT('h1)
	) name173 (
		_w179_,
		_w187_,
		_w188_
	);
	LUT2 #(
		.INIT('h1)
	) name174 (
		\v7_reg/NET0131 ,
		_w188_,
		_w189_
	);
	LUT2 #(
		.INIT('h4)
	) name175 (
		\v10_reg/NET0131 ,
		_w54_,
		_w190_
	);
	LUT2 #(
		.INIT('h4)
	) name176 (
		\v11_reg/NET0131 ,
		_w190_,
		_w191_
	);
	LUT2 #(
		.INIT('h2)
	) name177 (
		\v9_reg/NET0131 ,
		_w20_,
		_w192_
	);
	LUT2 #(
		.INIT('h2)
	) name178 (
		\v8_reg/NET0131 ,
		_w192_,
		_w193_
	);
	LUT2 #(
		.INIT('h8)
	) name179 (
		\v7_reg/NET0131 ,
		_w112_,
		_w194_
	);
	LUT2 #(
		.INIT('h1)
	) name180 (
		\v12_reg/NET0131 ,
		_w194_,
		_w195_
	);
	LUT2 #(
		.INIT('h4)
	) name181 (
		_w191_,
		_w193_,
		_w196_
	);
	LUT2 #(
		.INIT('h4)
	) name182 (
		_w195_,
		_w196_,
		_w197_
	);
	LUT2 #(
		.INIT('h1)
	) name183 (
		_w189_,
		_w197_,
		_w198_
	);
	LUT2 #(
		.INIT('h4)
	) name184 (
		_w21_,
		_w118_,
		_w199_
	);
	LUT2 #(
		.INIT('h8)
	) name185 (
		\v11_reg/NET0131 ,
		\v8_reg/NET0131 ,
		_w200_
	);
	LUT2 #(
		.INIT('h8)
	) name186 (
		_w175_,
		_w200_,
		_w201_
	);
	LUT2 #(
		.INIT('h1)
	) name187 (
		_w199_,
		_w201_,
		_w202_
	);
	LUT2 #(
		.INIT('h1)
	) name188 (
		\v12_reg/NET0131 ,
		\v7_reg/NET0131 ,
		_w203_
	);
	LUT2 #(
		.INIT('h2)
	) name189 (
		\v4_pad ,
		\v5_pad ,
		_w204_
	);
	LUT2 #(
		.INIT('h8)
	) name190 (
		_w203_,
		_w204_,
		_w205_
	);
	LUT2 #(
		.INIT('h4)
	) name191 (
		_w202_,
		_w205_,
		_w206_
	);
	LUT2 #(
		.INIT('h4)
	) name192 (
		\v1_pad ,
		\v6_pad ,
		_w207_
	);
	LUT2 #(
		.INIT('h2)
	) name193 (
		\v8_reg/NET0131 ,
		_w207_,
		_w208_
	);
	LUT2 #(
		.INIT('h2)
	) name194 (
		\v10_reg/NET0131 ,
		\v7_reg/NET0131 ,
		_w209_
	);
	LUT2 #(
		.INIT('h8)
	) name195 (
		_w98_,
		_w146_,
		_w210_
	);
	LUT2 #(
		.INIT('h8)
	) name196 (
		_w209_,
		_w210_,
		_w211_
	);
	LUT2 #(
		.INIT('h8)
	) name197 (
		_w208_,
		_w211_,
		_w212_
	);
	LUT2 #(
		.INIT('h2)
	) name198 (
		\v10_reg/NET0131 ,
		\v2_pad ,
		_w213_
	);
	LUT2 #(
		.INIT('h4)
	) name199 (
		_w22_,
		_w213_,
		_w214_
	);
	LUT2 #(
		.INIT('h2)
	) name200 (
		_w134_,
		_w214_,
		_w215_
	);
	LUT2 #(
		.INIT('h2)
	) name201 (
		\v9_reg/NET0131 ,
		_w215_,
		_w216_
	);
	LUT2 #(
		.INIT('h2)
	) name202 (
		_w162_,
		_w216_,
		_w217_
	);
	LUT2 #(
		.INIT('h8)
	) name203 (
		\v12_reg/NET0131 ,
		\v3_pad ,
		_w218_
	);
	LUT2 #(
		.INIT('h8)
	) name204 (
		_w20_,
		_w118_,
		_w219_
	);
	LUT2 #(
		.INIT('h8)
	) name205 (
		\v10_reg/NET0131 ,
		_w158_,
		_w220_
	);
	LUT2 #(
		.INIT('h8)
	) name206 (
		_w208_,
		_w220_,
		_w221_
	);
	LUT2 #(
		.INIT('h1)
	) name207 (
		_w219_,
		_w221_,
		_w222_
	);
	LUT2 #(
		.INIT('h2)
	) name208 (
		_w218_,
		_w222_,
		_w223_
	);
	LUT2 #(
		.INIT('h1)
	) name209 (
		\v11_reg/NET0131 ,
		_w47_,
		_w224_
	);
	LUT2 #(
		.INIT('h2)
	) name210 (
		\v11_reg/NET0131 ,
		_w38_,
		_w225_
	);
	LUT2 #(
		.INIT('h1)
	) name211 (
		_w224_,
		_w225_,
		_w226_
	);
	LUT2 #(
		.INIT('h4)
	) name212 (
		\v9_reg/NET0131 ,
		_w22_,
		_w227_
	);
	LUT2 #(
		.INIT('h1)
	) name213 (
		\v0_pad ,
		\v12_reg/NET0131 ,
		_w228_
	);
	LUT2 #(
		.INIT('h8)
	) name214 (
		_w227_,
		_w228_,
		_w229_
	);
	LUT2 #(
		.INIT('h1)
	) name215 (
		_w226_,
		_w229_,
		_w230_
	);
	LUT2 #(
		.INIT('h2)
	) name216 (
		\v10_reg/NET0131 ,
		_w230_,
		_w231_
	);
	LUT2 #(
		.INIT('h8)
	) name217 (
		\v6_pad ,
		_w20_,
		_w232_
	);
	LUT2 #(
		.INIT('h8)
	) name218 (
		\v12_reg/NET0131 ,
		_w232_,
		_w233_
	);
	LUT2 #(
		.INIT('h8)
	) name219 (
		_w118_,
		_w233_,
		_w234_
	);
	LUT2 #(
		.INIT('h4)
	) name220 (
		\v0_pad ,
		\v10_reg/NET0131 ,
		_w235_
	);
	LUT2 #(
		.INIT('h8)
	) name221 (
		_w200_,
		_w207_,
		_w236_
	);
	LUT2 #(
		.INIT('h8)
	) name222 (
		_w218_,
		_w235_,
		_w237_
	);
	LUT2 #(
		.INIT('h8)
	) name223 (
		_w236_,
		_w237_,
		_w238_
	);
	LUT2 #(
		.INIT('h1)
	) name224 (
		_w234_,
		_w238_,
		_w239_
	);
	LUT2 #(
		.INIT('h4)
	) name225 (
		_w217_,
		_w239_,
		_w240_
	);
	LUT2 #(
		.INIT('h1)
	) name226 (
		_w223_,
		_w231_,
		_w241_
	);
	LUT2 #(
		.INIT('h8)
	) name227 (
		_w240_,
		_w241_,
		_w242_
	);
	LUT2 #(
		.INIT('h1)
	) name228 (
		\v7_reg/NET0131 ,
		_w242_,
		_w243_
	);
	LUT2 #(
		.INIT('h8)
	) name229 (
		\v8_reg/NET0131 ,
		_w135_,
		_w244_
	);
	LUT2 #(
		.INIT('h4)
	) name230 (
		_w137_,
		_w244_,
		_w245_
	);
	LUT2 #(
		.INIT('h1)
	) name231 (
		\v12_reg/NET0131 ,
		\v8_reg/NET0131 ,
		_w246_
	);
	LUT2 #(
		.INIT('h1)
	) name232 (
		_w224_,
		_w246_,
		_w247_
	);
	LUT2 #(
		.INIT('h1)
	) name233 (
		\v10_reg/NET0131 ,
		_w89_,
		_w248_
	);
	LUT2 #(
		.INIT('h4)
	) name234 (
		_w247_,
		_w248_,
		_w249_
	);
	LUT2 #(
		.INIT('h1)
	) name235 (
		_w72_,
		_w249_,
		_w250_
	);
	LUT2 #(
		.INIT('h2)
	) name236 (
		\v7_reg/NET0131 ,
		_w250_,
		_w251_
	);
	LUT2 #(
		.INIT('h1)
	) name237 (
		\v12_reg/NET0131 ,
		\v2_pad ,
		_w252_
	);
	LUT2 #(
		.INIT('h2)
	) name238 (
		\v1_pad ,
		\v7_reg/NET0131 ,
		_w253_
	);
	LUT2 #(
		.INIT('h8)
	) name239 (
		_w38_,
		_w253_,
		_w254_
	);
	LUT2 #(
		.INIT('h8)
	) name240 (
		_w252_,
		_w254_,
		_w255_
	);
	LUT2 #(
		.INIT('h8)
	) name241 (
		_w232_,
		_w255_,
		_w256_
	);
	LUT2 #(
		.INIT('h1)
	) name242 (
		_w245_,
		_w256_,
		_w257_
	);
	LUT2 #(
		.INIT('h4)
	) name243 (
		_w251_,
		_w257_,
		_w258_
	);
	LUT2 #(
		.INIT('h4)
	) name244 (
		_w243_,
		_w258_,
		_w259_
	);
	LUT2 #(
		.INIT('h2)
	) name245 (
		CLR_pad,
		_w259_,
		_w260_
	);
	LUT2 #(
		.INIT('h4)
	) name246 (
		\v8_reg/NET0131 ,
		_w158_,
		_w261_
	);
	LUT2 #(
		.INIT('h2)
	) name247 (
		_w26_,
		_w53_,
		_w262_
	);
	LUT2 #(
		.INIT('h1)
	) name248 (
		_w261_,
		_w262_,
		_w263_
	);
	LUT2 #(
		.INIT('h2)
	) name249 (
		_w149_,
		_w263_,
		_w264_
	);
	LUT2 #(
		.INIT('h2)
	) name250 (
		\v11_reg/NET0131 ,
		_w135_,
		_w265_
	);
	LUT2 #(
		.INIT('h4)
	) name251 (
		\v10_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w266_
	);
	LUT2 #(
		.INIT('h1)
	) name252 (
		\v8_reg/NET0131 ,
		_w266_,
		_w267_
	);
	LUT2 #(
		.INIT('h8)
	) name253 (
		_w265_,
		_w267_,
		_w268_
	);
	LUT2 #(
		.INIT('h2)
	) name254 (
		\v8_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w269_
	);
	LUT2 #(
		.INIT('h1)
	) name255 (
		_w149_,
		_w200_,
		_w270_
	);
	LUT2 #(
		.INIT('h2)
	) name256 (
		_w22_,
		_w269_,
		_w271_
	);
	LUT2 #(
		.INIT('h4)
	) name257 (
		_w270_,
		_w271_,
		_w272_
	);
	LUT2 #(
		.INIT('h1)
	) name258 (
		_w268_,
		_w272_,
		_w273_
	);
	LUT2 #(
		.INIT('h4)
	) name259 (
		_w264_,
		_w273_,
		_w274_
	);
	LUT2 #(
		.INIT('h1)
	) name260 (
		\v12_reg/NET0131 ,
		_w274_,
		_w275_
	);
	LUT2 #(
		.INIT('h2)
	) name261 (
		\v11_reg/NET0131 ,
		_w252_,
		_w276_
	);
	LUT2 #(
		.INIT('h1)
	) name262 (
		\v7_reg/NET0131 ,
		_w276_,
		_w277_
	);
	LUT2 #(
		.INIT('h2)
	) name263 (
		_w26_,
		_w47_,
		_w278_
	);
	LUT2 #(
		.INIT('h2)
	) name264 (
		\v8_reg/NET0131 ,
		_w98_,
		_w279_
	);
	LUT2 #(
		.INIT('h4)
	) name265 (
		_w186_,
		_w279_,
		_w280_
	);
	LUT2 #(
		.INIT('h4)
	) name266 (
		_w278_,
		_w280_,
		_w281_
	);
	LUT2 #(
		.INIT('h4)
	) name267 (
		_w277_,
		_w281_,
		_w282_
	);
	LUT2 #(
		.INIT('h1)
	) name268 (
		_w275_,
		_w282_,
		_w283_
	);
	LUT2 #(
		.INIT('h8)
	) name269 (
		_w71_,
		_w103_,
		_w284_
	);
	LUT2 #(
		.INIT('h4)
	) name270 (
		_w15_,
		_w157_,
		_w285_
	);
	LUT2 #(
		.INIT('h8)
	) name271 (
		_w26_,
		_w71_,
		_w286_
	);
	LUT2 #(
		.INIT('h1)
	) name272 (
		_w284_,
		_w285_,
		_w287_
	);
	LUT2 #(
		.INIT('h4)
	) name273 (
		_w286_,
		_w287_,
		_w288_
	);
	LUT2 #(
		.INIT('h1)
	) name274 (
		\v8_reg/NET0131 ,
		_w288_,
		_w289_
	);
	LUT2 #(
		.INIT('h4)
	) name275 (
		\v12_reg/NET0131 ,
		\v1_pad ,
		_w290_
	);
	LUT2 #(
		.INIT('h2)
	) name276 (
		_w18_,
		_w207_,
		_w291_
	);
	LUT2 #(
		.INIT('h1)
	) name277 (
		_w290_,
		_w291_,
		_w292_
	);
	LUT2 #(
		.INIT('h2)
	) name278 (
		\v3_pad ,
		_w292_,
		_w293_
	);
	LUT2 #(
		.INIT('h1)
	) name279 (
		\v12_reg/NET0131 ,
		_w89_,
		_w294_
	);
	LUT2 #(
		.INIT('h2)
	) name280 (
		\v12_reg/NET0131 ,
		\v8_reg/NET0131 ,
		_w295_
	);
	LUT2 #(
		.INIT('h8)
	) name281 (
		_w26_,
		_w295_,
		_w296_
	);
	LUT2 #(
		.INIT('h2)
	) name282 (
		\v9_reg/NET0131 ,
		_w294_,
		_w297_
	);
	LUT2 #(
		.INIT('h4)
	) name283 (
		_w296_,
		_w297_,
		_w298_
	);
	LUT2 #(
		.INIT('h4)
	) name284 (
		_w293_,
		_w298_,
		_w299_
	);
	LUT2 #(
		.INIT('h8)
	) name285 (
		_w118_,
		_w235_,
		_w300_
	);
	LUT2 #(
		.INIT('h8)
	) name286 (
		_w22_,
		_w134_,
		_w301_
	);
	LUT2 #(
		.INIT('h8)
	) name287 (
		_w300_,
		_w301_,
		_w302_
	);
	LUT2 #(
		.INIT('h1)
	) name288 (
		_w289_,
		_w302_,
		_w303_
	);
	LUT2 #(
		.INIT('h4)
	) name289 (
		_w299_,
		_w303_,
		_w304_
	);
	LUT2 #(
		.INIT('h1)
	) name290 (
		\v7_reg/NET0131 ,
		_w304_,
		_w305_
	);
	LUT2 #(
		.INIT('h8)
	) name291 (
		_w22_,
		_w200_,
		_w306_
	);
	LUT2 #(
		.INIT('h1)
	) name292 (
		_w89_,
		_w306_,
		_w307_
	);
	LUT2 #(
		.INIT('h4)
	) name293 (
		\v7_reg/NET0131 ,
		_w71_,
		_w308_
	);
	LUT2 #(
		.INIT('h4)
	) name294 (
		_w307_,
		_w308_,
		_w309_
	);
	LUT2 #(
		.INIT('h8)
	) name295 (
		\v7_reg/NET0131 ,
		\v8_reg/NET0131 ,
		_w310_
	);
	LUT2 #(
		.INIT('h8)
	) name296 (
		_w54_,
		_w310_,
		_w311_
	);
	LUT2 #(
		.INIT('h1)
	) name297 (
		_w309_,
		_w311_,
		_w312_
	);
	LUT2 #(
		.INIT('h1)
	) name298 (
		\v2_pad ,
		_w312_,
		_w313_
	);
	LUT2 #(
		.INIT('h2)
	) name299 (
		\v7_reg/NET0131 ,
		_w18_,
		_w314_
	);
	LUT2 #(
		.INIT('h4)
	) name300 (
		_w47_,
		_w314_,
		_w315_
	);
	LUT2 #(
		.INIT('h8)
	) name301 (
		_w193_,
		_w315_,
		_w316_
	);
	LUT2 #(
		.INIT('h1)
	) name302 (
		_w313_,
		_w316_,
		_w317_
	);
	LUT2 #(
		.INIT('h4)
	) name303 (
		_w305_,
		_w317_,
		_w318_
	);
	LUT2 #(
		.INIT('h2)
	) name304 (
		CLR_pad,
		_w318_,
		_w319_
	);
	LUT2 #(
		.INIT('h8)
	) name305 (
		\v0_pad ,
		_w207_,
		_w320_
	);
	LUT2 #(
		.INIT('h8)
	) name306 (
		\v3_pad ,
		_w98_,
		_w321_
	);
	LUT2 #(
		.INIT('h4)
	) name307 (
		_w320_,
		_w321_,
		_w322_
	);
	LUT2 #(
		.INIT('h1)
	) name308 (
		\v3_pad ,
		\v9_reg/NET0131 ,
		_w323_
	);
	LUT2 #(
		.INIT('h2)
	) name309 (
		_w134_,
		_w323_,
		_w324_
	);
	LUT2 #(
		.INIT('h1)
	) name310 (
		\v10_reg/NET0131 ,
		_w324_,
		_w325_
	);
	LUT2 #(
		.INIT('h1)
	) name311 (
		\v12_reg/NET0131 ,
		_w112_,
		_w326_
	);
	LUT2 #(
		.INIT('h1)
	) name312 (
		\v2_pad ,
		_w107_,
		_w327_
	);
	LUT2 #(
		.INIT('h8)
	) name313 (
		_w326_,
		_w327_,
		_w328_
	);
	LUT2 #(
		.INIT('h1)
	) name314 (
		_w224_,
		_w322_,
		_w329_
	);
	LUT2 #(
		.INIT('h4)
	) name315 (
		_w325_,
		_w329_,
		_w330_
	);
	LUT2 #(
		.INIT('h4)
	) name316 (
		_w328_,
		_w330_,
		_w331_
	);
	LUT2 #(
		.INIT('h2)
	) name317 (
		\v8_reg/NET0131 ,
		_w331_,
		_w332_
	);
	LUT2 #(
		.INIT('h4)
	) name318 (
		\v10_reg/NET0131 ,
		_w45_,
		_w333_
	);
	LUT2 #(
		.INIT('h4)
	) name319 (
		\v11_reg/NET0131 ,
		_w54_,
		_w334_
	);
	LUT2 #(
		.INIT('h1)
	) name320 (
		_w105_,
		_w334_,
		_w335_
	);
	LUT2 #(
		.INIT('h1)
	) name321 (
		\v6_pad ,
		_w335_,
		_w336_
	);
	LUT2 #(
		.INIT('h4)
	) name322 (
		\v1_pad ,
		_w266_,
		_w337_
	);
	LUT2 #(
		.INIT('h1)
	) name323 (
		_w168_,
		_w337_,
		_w338_
	);
	LUT2 #(
		.INIT('h2)
	) name324 (
		_w246_,
		_w338_,
		_w339_
	);
	LUT2 #(
		.INIT('h1)
	) name325 (
		_w278_,
		_w333_,
		_w340_
	);
	LUT2 #(
		.INIT('h4)
	) name326 (
		_w336_,
		_w340_,
		_w341_
	);
	LUT2 #(
		.INIT('h4)
	) name327 (
		_w339_,
		_w341_,
		_w342_
	);
	LUT2 #(
		.INIT('h4)
	) name328 (
		_w332_,
		_w342_,
		_w343_
	);
	LUT2 #(
		.INIT('h1)
	) name329 (
		\v7_reg/NET0131 ,
		_w343_,
		_w344_
	);
	LUT2 #(
		.INIT('h1)
	) name330 (
		\v10_reg/NET0131 ,
		_w200_,
		_w345_
	);
	LUT2 #(
		.INIT('h1)
	) name331 (
		\v11_reg/NET0131 ,
		\v12_reg/NET0131 ,
		_w346_
	);
	LUT2 #(
		.INIT('h1)
	) name332 (
		\v8_reg/NET0131 ,
		_w71_,
		_w347_
	);
	LUT2 #(
		.INIT('h2)
	) name333 (
		_w345_,
		_w346_,
		_w348_
	);
	LUT2 #(
		.INIT('h4)
	) name334 (
		_w347_,
		_w348_,
		_w349_
	);
	LUT2 #(
		.INIT('h8)
	) name335 (
		\v10_reg/NET0131 ,
		\v8_reg/NET0131 ,
		_w350_
	);
	LUT2 #(
		.INIT('h8)
	) name336 (
		\v11_reg/NET0131 ,
		\v2_pad ,
		_w351_
	);
	LUT2 #(
		.INIT('h8)
	) name337 (
		_w55_,
		_w351_,
		_w352_
	);
	LUT2 #(
		.INIT('h8)
	) name338 (
		_w350_,
		_w352_,
		_w353_
	);
	LUT2 #(
		.INIT('h4)
	) name339 (
		\v12_reg/NET0131 ,
		\v2_pad ,
		_w354_
	);
	LUT2 #(
		.INIT('h4)
	) name340 (
		\v7_reg/NET0131 ,
		_w266_,
		_w355_
	);
	LUT2 #(
		.INIT('h8)
	) name341 (
		_w354_,
		_w355_,
		_w356_
	);
	LUT2 #(
		.INIT('h1)
	) name342 (
		\v11_reg/NET0131 ,
		_w244_,
		_w357_
	);
	LUT2 #(
		.INIT('h4)
	) name343 (
		\v12_reg/NET0131 ,
		\v7_reg/NET0131 ,
		_w358_
	);
	LUT2 #(
		.INIT('h4)
	) name344 (
		_w180_,
		_w358_,
		_w359_
	);
	LUT2 #(
		.INIT('h4)
	) name345 (
		_w357_,
		_w359_,
		_w360_
	);
	LUT2 #(
		.INIT('h1)
	) name346 (
		_w349_,
		_w356_,
		_w361_
	);
	LUT2 #(
		.INIT('h1)
	) name347 (
		_w353_,
		_w360_,
		_w362_
	);
	LUT2 #(
		.INIT('h8)
	) name348 (
		_w361_,
		_w362_,
		_w363_
	);
	LUT2 #(
		.INIT('h4)
	) name349 (
		_w344_,
		_w363_,
		_w364_
	);
	LUT2 #(
		.INIT('h2)
	) name350 (
		CLR_pad,
		_w364_,
		_w365_
	);
	LUT2 #(
		.INIT('h1)
	) name351 (
		_w71_,
		_w104_,
		_w366_
	);
	LUT2 #(
		.INIT('h1)
	) name352 (
		\v3_pad ,
		_w246_,
		_w367_
	);
	LUT2 #(
		.INIT('h4)
	) name353 (
		_w366_,
		_w367_,
		_w368_
	);
	LUT2 #(
		.INIT('h1)
	) name354 (
		_w113_,
		_w368_,
		_w369_
	);
	LUT2 #(
		.INIT('h1)
	) name355 (
		\v11_reg/NET0131 ,
		_w369_,
		_w370_
	);
	LUT2 #(
		.INIT('h1)
	) name356 (
		\v11_reg/NET0131 ,
		_w354_,
		_w371_
	);
	LUT2 #(
		.INIT('h1)
	) name357 (
		_w59_,
		_w371_,
		_w372_
	);
	LUT2 #(
		.INIT('h2)
	) name358 (
		_w269_,
		_w372_,
		_w373_
	);
	LUT2 #(
		.INIT('h2)
	) name359 (
		\v10_reg/NET0131 ,
		_w38_,
		_w374_
	);
	LUT2 #(
		.INIT('h4)
	) name360 (
		_w104_,
		_w354_,
		_w375_
	);
	LUT2 #(
		.INIT('h4)
	) name361 (
		_w374_,
		_w375_,
		_w376_
	);
	LUT2 #(
		.INIT('h1)
	) name362 (
		_w168_,
		_w266_,
		_w377_
	);
	LUT2 #(
		.INIT('h4)
	) name363 (
		_w232_,
		_w377_,
		_w378_
	);
	LUT2 #(
		.INIT('h2)
	) name364 (
		_w295_,
		_w378_,
		_w379_
	);
	LUT2 #(
		.INIT('h8)
	) name365 (
		\v11_reg/NET0131 ,
		_w322_,
		_w380_
	);
	LUT2 #(
		.INIT('h4)
	) name366 (
		_w22_,
		_w59_,
		_w381_
	);
	LUT2 #(
		.INIT('h1)
	) name367 (
		_w119_,
		_w284_,
		_w382_
	);
	LUT2 #(
		.INIT('h4)
	) name368 (
		_w381_,
		_w382_,
		_w383_
	);
	LUT2 #(
		.INIT('h4)
	) name369 (
		_w380_,
		_w383_,
		_w384_
	);
	LUT2 #(
		.INIT('h2)
	) name370 (
		\v8_reg/NET0131 ,
		_w384_,
		_w385_
	);
	LUT2 #(
		.INIT('h1)
	) name371 (
		_w373_,
		_w376_,
		_w386_
	);
	LUT2 #(
		.INIT('h4)
	) name372 (
		_w370_,
		_w386_,
		_w387_
	);
	LUT2 #(
		.INIT('h4)
	) name373 (
		_w379_,
		_w387_,
		_w388_
	);
	LUT2 #(
		.INIT('h4)
	) name374 (
		_w385_,
		_w388_,
		_w389_
	);
	LUT2 #(
		.INIT('h1)
	) name375 (
		\v7_reg/NET0131 ,
		_w389_,
		_w390_
	);
	LUT2 #(
		.INIT('h2)
	) name376 (
		\v10_reg/NET0131 ,
		_w54_,
		_w391_
	);
	LUT2 #(
		.INIT('h2)
	) name377 (
		_w62_,
		_w190_,
		_w392_
	);
	LUT2 #(
		.INIT('h4)
	) name378 (
		_w391_,
		_w392_,
		_w393_
	);
	LUT2 #(
		.INIT('h1)
	) name379 (
		\v11_reg/NET0131 ,
		_w46_,
		_w394_
	);
	LUT2 #(
		.INIT('h8)
	) name380 (
		\v9_reg/NET0131 ,
		_w358_,
		_w395_
	);
	LUT2 #(
		.INIT('h4)
	) name381 (
		_w394_,
		_w395_,
		_w396_
	);
	LUT2 #(
		.INIT('h1)
	) name382 (
		_w393_,
		_w396_,
		_w397_
	);
	LUT2 #(
		.INIT('h4)
	) name383 (
		_w390_,
		_w397_,
		_w398_
	);
	LUT2 #(
		.INIT('h2)
	) name384 (
		CLR_pad,
		_w398_,
		_w399_
	);
	LUT2 #(
		.INIT('h8)
	) name385 (
		_w104_,
		_w134_,
		_w400_
	);
	LUT2 #(
		.INIT('h2)
	) name386 (
		_w22_,
		_w62_,
		_w401_
	);
	LUT2 #(
		.INIT('h1)
	) name387 (
		\v9_reg/NET0131 ,
		_w26_,
		_w402_
	);
	LUT2 #(
		.INIT('h4)
	) name388 (
		_w158_,
		_w402_,
		_w403_
	);
	LUT2 #(
		.INIT('h1)
	) name389 (
		\v8_reg/NET0131 ,
		_w403_,
		_w404_
	);
	LUT2 #(
		.INIT('h2)
	) name390 (
		\v8_reg/NET0131 ,
		_w68_,
		_w405_
	);
	LUT2 #(
		.INIT('h8)
	) name391 (
		\v6_pad ,
		_w100_,
		_w406_
	);
	LUT2 #(
		.INIT('h2)
	) name392 (
		_w405_,
		_w406_,
		_w407_
	);
	LUT2 #(
		.INIT('h1)
	) name393 (
		\v12_reg/NET0131 ,
		_w401_,
		_w408_
	);
	LUT2 #(
		.INIT('h4)
	) name394 (
		_w407_,
		_w408_,
		_w409_
	);
	LUT2 #(
		.INIT('h4)
	) name395 (
		_w404_,
		_w409_,
		_w410_
	);
	LUT2 #(
		.INIT('h1)
	) name396 (
		\v7_reg/NET0131 ,
		_w410_,
		_w411_
	);
	LUT2 #(
		.INIT('h1)
	) name397 (
		_w193_,
		_w400_,
		_w412_
	);
	LUT2 #(
		.INIT('h4)
	) name398 (
		_w411_,
		_w412_,
		_w413_
	);
	LUT2 #(
		.INIT('h2)
	) name399 (
		\v12_reg/NET0131 ,
		_w26_,
		_w414_
	);
	LUT2 #(
		.INIT('h4)
	) name400 (
		\v10_reg/NET0131 ,
		_w22_,
		_w415_
	);
	LUT2 #(
		.INIT('h1)
	) name401 (
		\v12_reg/NET0131 ,
		_w158_,
		_w416_
	);
	LUT2 #(
		.INIT('h4)
	) name402 (
		_w415_,
		_w416_,
		_w417_
	);
	LUT2 #(
		.INIT('h1)
	) name403 (
		\v9_reg/NET0131 ,
		_w414_,
		_w418_
	);
	LUT2 #(
		.INIT('h4)
	) name404 (
		_w417_,
		_w418_,
		_w419_
	);
	LUT2 #(
		.INIT('h1)
	) name405 (
		_w72_,
		_w419_,
		_w420_
	);
	LUT2 #(
		.INIT('h1)
	) name406 (
		\v7_reg/NET0131 ,
		_w420_,
		_w421_
	);
	LUT2 #(
		.INIT('h4)
	) name407 (
		\v12_reg/NET0131 ,
		_w186_,
		_w422_
	);
	LUT2 #(
		.INIT('h1)
	) name408 (
		_w421_,
		_w422_,
		_w423_
	);
	LUT2 #(
		.INIT('h1)
	) name409 (
		\v8_reg/NET0131 ,
		_w423_,
		_w424_
	);
	LUT2 #(
		.INIT('h1)
	) name410 (
		_w98_,
		_w112_,
		_w425_
	);
	LUT2 #(
		.INIT('h8)
	) name411 (
		_w276_,
		_w425_,
		_w426_
	);
	LUT2 #(
		.INIT('h1)
	) name412 (
		_w358_,
		_w426_,
		_w427_
	);
	LUT2 #(
		.INIT('h2)
	) name413 (
		\v8_reg/NET0131 ,
		_w427_,
		_w428_
	);
	LUT2 #(
		.INIT('h1)
	) name414 (
		_w424_,
		_w428_,
		_w429_
	);
	LUT2 #(
		.INIT('h2)
	) name415 (
		\v11_reg/NET0131 ,
		_w235_,
		_w430_
	);
	LUT2 #(
		.INIT('h1)
	) name416 (
		\v9_reg/NET0131 ,
		_w430_,
		_w431_
	);
	LUT2 #(
		.INIT('h4)
	) name417 (
		\v8_reg/NET0131 ,
		_w431_,
		_w432_
	);
	LUT2 #(
		.INIT('h1)
	) name418 (
		_w201_,
		_w432_,
		_w433_
	);
	LUT2 #(
		.INIT('h2)
	) name419 (
		_w22_,
		_w433_,
		_w434_
	);
	LUT2 #(
		.INIT('h8)
	) name420 (
		_w162_,
		_w351_,
		_w435_
	);
	LUT2 #(
		.INIT('h1)
	) name421 (
		_w434_,
		_w435_,
		_w436_
	);
	LUT2 #(
		.INIT('h1)
	) name422 (
		\v12_reg/NET0131 ,
		_w436_,
		_w437_
	);
	LUT2 #(
		.INIT('h1)
	) name423 (
		_w15_,
		_w295_,
		_w438_
	);
	LUT2 #(
		.INIT('h1)
	) name424 (
		\v9_reg/NET0131 ,
		_w27_,
		_w439_
	);
	LUT2 #(
		.INIT('h4)
	) name425 (
		_w438_,
		_w439_,
		_w440_
	);
	LUT2 #(
		.INIT('h1)
	) name426 (
		_w437_,
		_w440_,
		_w441_
	);
	LUT2 #(
		.INIT('h1)
	) name427 (
		\v7_reg/NET0131 ,
		_w441_,
		_w442_
	);
	LUT2 #(
		.INIT('h4)
	) name428 (
		_w39_,
		_w112_,
		_w443_
	);
	LUT2 #(
		.INIT('h1)
	) name429 (
		_w286_,
		_w443_,
		_w444_
	);
	LUT2 #(
		.INIT('h2)
	) name430 (
		\v8_reg/NET0131 ,
		_w444_,
		_w445_
	);
	LUT2 #(
		.INIT('h1)
	) name431 (
		_w400_,
		_w445_,
		_w446_
	);
	LUT2 #(
		.INIT('h2)
	) name432 (
		\v7_reg/NET0131 ,
		_w446_,
		_w447_
	);
	LUT2 #(
		.INIT('h1)
	) name433 (
		_w200_,
		_w203_,
		_w448_
	);
	LUT2 #(
		.INIT('h1)
	) name434 (
		\v9_reg/NET0131 ,
		_w448_,
		_w449_
	);
	LUT2 #(
		.INIT('h1)
	) name435 (
		_w290_,
		_w449_,
		_w450_
	);
	LUT2 #(
		.INIT('h4)
	) name436 (
		_w157_,
		_w290_,
		_w451_
	);
	LUT2 #(
		.INIT('h2)
	) name437 (
		\v10_reg/NET0131 ,
		_w451_,
		_w452_
	);
	LUT2 #(
		.INIT('h4)
	) name438 (
		_w450_,
		_w452_,
		_w453_
	);
	LUT2 #(
		.INIT('h1)
	) name439 (
		_w447_,
		_w453_,
		_w454_
	);
	LUT2 #(
		.INIT('h4)
	) name440 (
		_w442_,
		_w454_,
		_w455_
	);
	LUT2 #(
		.INIT('h1)
	) name441 (
		\v8_reg/NET0131 ,
		_w265_,
		_w456_
	);
	LUT2 #(
		.INIT('h2)
	) name442 (
		_w358_,
		_w456_,
		_w457_
	);
	LUT2 #(
		.INIT('h1)
	) name443 (
		\v8_reg/NET0131 ,
		_w431_,
		_w458_
	);
	LUT2 #(
		.INIT('h1)
	) name444 (
		\v4_pad ,
		\v5_pad ,
		_w459_
	);
	LUT2 #(
		.INIT('h1)
	) name445 (
		\v12_reg/NET0131 ,
		_w22_,
		_w460_
	);
	LUT2 #(
		.INIT('h1)
	) name446 (
		_w26_,
		_w459_,
		_w461_
	);
	LUT2 #(
		.INIT('h8)
	) name447 (
		_w460_,
		_w461_,
		_w462_
	);
	LUT2 #(
		.INIT('h4)
	) name448 (
		_w405_,
		_w462_,
		_w463_
	);
	LUT2 #(
		.INIT('h4)
	) name449 (
		_w458_,
		_w463_,
		_w464_
	);
	LUT2 #(
		.INIT('h1)
	) name450 (
		\v7_reg/NET0131 ,
		_w464_,
		_w465_
	);
	LUT2 #(
		.INIT('h1)
	) name451 (
		_w193_,
		_w457_,
		_w466_
	);
	LUT2 #(
		.INIT('h4)
	) name452 (
		_w465_,
		_w466_,
		_w467_
	);
	LUT2 #(
		.INIT('h8)
	) name453 (
		_w308_,
		_w406_,
		_w468_
	);
	LUT2 #(
		.INIT('h1)
	) name454 (
		_w352_,
		_w468_,
		_w469_
	);
	LUT2 #(
		.INIT('h2)
	) name455 (
		_w350_,
		_w469_,
		_w470_
	);
	LUT2 #(
		.INIT('h8)
	) name456 (
		_w22_,
		_w219_,
		_w471_
	);
	LUT2 #(
		.INIT('h8)
	) name457 (
		\v8_reg/NET0131 ,
		_w175_,
		_w472_
	);
	LUT2 #(
		.INIT('h1)
	) name458 (
		_w300_,
		_w472_,
		_w473_
	);
	LUT2 #(
		.INIT('h2)
	) name459 (
		\v11_reg/NET0131 ,
		_w459_,
		_w474_
	);
	LUT2 #(
		.INIT('h4)
	) name460 (
		_w473_,
		_w474_,
		_w475_
	);
	LUT2 #(
		.INIT('h1)
	) name461 (
		_w471_,
		_w475_,
		_w476_
	);
	LUT2 #(
		.INIT('h2)
	) name462 (
		_w203_,
		_w476_,
		_w477_
	);
	LUT2 #(
		.INIT('h8)
	) name463 (
		_w54_,
		_w148_,
		_w478_
	);
	LUT2 #(
		.INIT('h8)
	) name464 (
		\v6_pad ,
		_w15_,
		_w479_
	);
	LUT2 #(
		.INIT('h8)
	) name465 (
		_w109_,
		_w479_,
		_w480_
	);
	LUT2 #(
		.INIT('h1)
	) name466 (
		_w478_,
		_w480_,
		_w481_
	);
	LUT2 #(
		.INIT('h4)
	) name467 (
		\v7_reg/NET0131 ,
		_w100_,
		_w482_
	);
	LUT2 #(
		.INIT('h4)
	) name468 (
		_w481_,
		_w482_,
		_w483_
	);
	LUT2 #(
		.INIT('h1)
	) name469 (
		_w353_,
		_w483_,
		_w484_
	);
	LUT2 #(
		.INIT('h8)
	) name470 (
		_w89_,
		_w227_,
		_w485_
	);
	LUT2 #(
		.INIT('h8)
	) name471 (
		\v2_pad ,
		_w109_,
		_w486_
	);
	LUT2 #(
		.INIT('h1)
	) name472 (
		_w485_,
		_w486_,
		_w487_
	);
	LUT2 #(
		.INIT('h4)
	) name473 (
		\v10_reg/NET0131 ,
		_w203_,
		_w488_
	);
	LUT2 #(
		.INIT('h4)
	) name474 (
		_w487_,
		_w488_,
		_w489_
	);
	LUT2 #(
		.INIT('h8)
	) name475 (
		_w286_,
		_w310_,
		_w490_
	);
	LUT2 #(
		.INIT('h8)
	) name476 (
		_w62_,
		_w252_,
		_w491_
	);
	LUT2 #(
		.INIT('h8)
	) name477 (
		\v12_reg/NET0131 ,
		_w38_,
		_w492_
	);
	LUT2 #(
		.INIT('h1)
	) name478 (
		_w491_,
		_w492_,
		_w493_
	);
	LUT2 #(
		.INIT('h1)
	) name479 (
		\v10_reg/NET0131 ,
		\v7_reg/NET0131 ,
		_w494_
	);
	LUT2 #(
		.INIT('h4)
	) name480 (
		_w493_,
		_w494_,
		_w495_
	);
	LUT2 #(
		.INIT('h1)
	) name481 (
		_w490_,
		_w495_,
		_w496_
	);
	LUT2 #(
		.INIT('h8)
	) name482 (
		\v0_pad ,
		_w56_,
		_w497_
	);
	LUT2 #(
		.INIT('h1)
	) name483 (
		_w233_,
		_w497_,
		_w498_
	);
	LUT2 #(
		.INIT('h1)
	) name484 (
		\v9_reg/NET0131 ,
		_w498_,
		_w499_
	);
	LUT2 #(
		.INIT('h8)
	) name485 (
		\v10_reg/NET0131 ,
		_w45_,
		_w500_
	);
	LUT2 #(
		.INIT('h1)
	) name486 (
		_w499_,
		_w500_,
		_w501_
	);
	LUT2 #(
		.INIT('h2)
	) name487 (
		_w155_,
		_w501_,
		_w502_
	);
	LUT2 #(
		.INIT('h8)
	) name488 (
		_w100_,
		_w480_,
		_w503_
	);
	LUT2 #(
		.INIT('h1)
	) name489 (
		\v12_reg/NET0131 ,
		\v5_pad ,
		_w504_
	);
	LUT2 #(
		.INIT('h2)
	) name490 (
		_w27_,
		_w504_,
		_w505_
	);
	LUT2 #(
		.INIT('h2)
	) name491 (
		_w118_,
		_w139_,
		_w506_
	);
	LUT2 #(
		.INIT('h4)
	) name492 (
		_w505_,
		_w506_,
		_w507_
	);
	LUT2 #(
		.INIT('h1)
	) name493 (
		_w503_,
		_w507_,
		_w508_
	);
	LUT2 #(
		.INIT('h1)
	) name494 (
		\v7_reg/NET0131 ,
		_w508_,
		_w509_
	);
	LUT2 #(
		.INIT('h2)
	) name495 (
		\v10_reg/NET0131 ,
		_w109_,
		_w510_
	);
	LUT2 #(
		.INIT('h4)
	) name496 (
		\v10_reg/NET0131 ,
		_w109_,
		_w511_
	);
	LUT2 #(
		.INIT('h2)
	) name497 (
		_w358_,
		_w510_,
		_w512_
	);
	LUT2 #(
		.INIT('h4)
	) name498 (
		_w511_,
		_w512_,
		_w513_
	);
	LUT2 #(
		.INIT('h4)
	) name499 (
		\v10_reg/NET0131 ,
		\v7_reg/NET0131 ,
		_w514_
	);
	LUT2 #(
		.INIT('h8)
	) name500 (
		\v9_reg/NET0131 ,
		_w504_,
		_w515_
	);
	LUT2 #(
		.INIT('h1)
	) name501 (
		_w55_,
		_w515_,
		_w516_
	);
	LUT2 #(
		.INIT('h2)
	) name502 (
		_w53_,
		_w514_,
		_w517_
	);
	LUT2 #(
		.INIT('h4)
	) name503 (
		_w516_,
		_w517_,
		_w518_
	);
	LUT2 #(
		.INIT('h1)
	) name504 (
		_w513_,
		_w518_,
		_w519_
	);
	LUT2 #(
		.INIT('h2)
	) name505 (
		\v11_reg/NET0131 ,
		_w519_,
		_w520_
	);
	LUT2 #(
		.INIT('h8)
	) name506 (
		_w53_,
		_w514_,
		_w521_
	);
	LUT2 #(
		.INIT('h4)
	) name507 (
		\v5_pad ,
		_w18_,
		_w522_
	);
	LUT2 #(
		.INIT('h8)
	) name508 (
		_w155_,
		_w522_,
		_w523_
	);
	LUT2 #(
		.INIT('h1)
	) name509 (
		_w521_,
		_w523_,
		_w524_
	);
	LUT2 #(
		.INIT('h4)
	) name510 (
		\v0_pad ,
		_w47_,
		_w525_
	);
	LUT2 #(
		.INIT('h4)
	) name511 (
		_w524_,
		_w525_,
		_w526_
	);
	LUT2 #(
		.INIT('h1)
	) name512 (
		_w509_,
		_w526_,
		_w527_
	);
	LUT2 #(
		.INIT('h4)
	) name513 (
		_w520_,
		_w527_,
		_w528_
	);
	LUT2 #(
		.INIT('h1)
	) name514 (
		_w190_,
		_w326_,
		_w529_
	);
	LUT2 #(
		.INIT('h2)
	) name515 (
		_w62_,
		_w529_,
		_w530_
	);
	LUT2 #(
		.INIT('h8)
	) name516 (
		_w71_,
		_w75_,
		_w531_
	);
	LUT2 #(
		.INIT('h1)
	) name517 (
		_w530_,
		_w531_,
		_w532_
	);
	LUT2 #(
		.INIT('h2)
	) name518 (
		\v7_reg/NET0131 ,
		_w532_,
		_w533_
	);
	LUT2 #(
		.INIT('h1)
	) name519 (
		_w16_,
		_w119_,
		_w534_
	);
	LUT2 #(
		.INIT('h1)
	) name520 (
		\v8_reg/NET0131 ,
		_w534_,
		_w535_
	);
	LUT2 #(
		.INIT('h4)
	) name521 (
		\v12_reg/NET0131 ,
		_w94_,
		_w536_
	);
	LUT2 #(
		.INIT('h1)
	) name522 (
		_w535_,
		_w536_,
		_w537_
	);
	LUT2 #(
		.INIT('h1)
	) name523 (
		\v9_reg/NET0131 ,
		_w537_,
		_w538_
	);
	LUT2 #(
		.INIT('h1)
	) name524 (
		_w201_,
		_w300_,
		_w539_
	);
	LUT2 #(
		.INIT('h1)
	) name525 (
		\v12_reg/NET0131 ,
		_w181_,
		_w540_
	);
	LUT2 #(
		.INIT('h4)
	) name526 (
		_w539_,
		_w540_,
		_w541_
	);
	LUT2 #(
		.INIT('h1)
	) name527 (
		_w538_,
		_w541_,
		_w542_
	);
	LUT2 #(
		.INIT('h1)
	) name528 (
		\v7_reg/NET0131 ,
		_w542_,
		_w543_
	);
	LUT2 #(
		.INIT('h1)
	) name529 (
		_w533_,
		_w543_,
		_w544_
	);
	LUT2 #(
		.INIT('h2)
	) name530 (
		\v11_reg/NET0131 ,
		\v8_reg/NET0131 ,
		_w545_
	);
	LUT2 #(
		.INIT('h1)
	) name531 (
		_w175_,
		_w545_,
		_w546_
	);
	LUT2 #(
		.INIT('h1)
	) name532 (
		_w181_,
		_w546_,
		_w547_
	);
	LUT2 #(
		.INIT('h1)
	) name533 (
		\v8_reg/NET0131 ,
		_w15_,
		_w548_
	);
	LUT2 #(
		.INIT('h8)
	) name534 (
		\v10_reg/NET0131 ,
		_w252_,
		_w549_
	);
	LUT2 #(
		.INIT('h1)
	) name535 (
		_w548_,
		_w549_,
		_w550_
	);
	LUT2 #(
		.INIT('h1)
	) name536 (
		\v9_reg/NET0131 ,
		_w550_,
		_w551_
	);
	LUT2 #(
		.INIT('h1)
	) name537 (
		\v11_reg/NET0131 ,
		_w551_,
		_w552_
	);
	LUT2 #(
		.INIT('h2)
	) name538 (
		\v11_reg/NET0131 ,
		_w228_,
		_w553_
	);
	LUT2 #(
		.INIT('h1)
	) name539 (
		\v9_reg/NET0131 ,
		_w16_,
		_w554_
	);
	LUT2 #(
		.INIT('h4)
	) name540 (
		_w553_,
		_w554_,
		_w555_
	);
	LUT2 #(
		.INIT('h1)
	) name541 (
		\v8_reg/NET0131 ,
		_w555_,
		_w556_
	);
	LUT2 #(
		.INIT('h2)
	) name542 (
		_w112_,
		_w346_,
		_w557_
	);
	LUT2 #(
		.INIT('h1)
	) name543 (
		\v7_reg/NET0131 ,
		_w98_,
		_w558_
	);
	LUT2 #(
		.INIT('h4)
	) name544 (
		_w557_,
		_w558_,
		_w559_
	);
	LUT2 #(
		.INIT('h4)
	) name545 (
		_w547_,
		_w559_,
		_w560_
	);
	LUT2 #(
		.INIT('h4)
	) name546 (
		_w552_,
		_w560_,
		_w561_
	);
	LUT2 #(
		.INIT('h4)
	) name547 (
		_w556_,
		_w561_,
		_w562_
	);
	LUT2 #(
		.INIT('h2)
	) name548 (
		\v9_reg/NET0131 ,
		_w346_,
		_w563_
	);
	LUT2 #(
		.INIT('h4)
	) name549 (
		_w39_,
		_w350_,
		_w564_
	);
	LUT2 #(
		.INIT('h4)
	) name550 (
		_w563_,
		_w564_,
		_w565_
	);
	LUT2 #(
		.INIT('h2)
	) name551 (
		\v7_reg/NET0131 ,
		_w400_,
		_w566_
	);
	LUT2 #(
		.INIT('h4)
	) name552 (
		_w565_,
		_w566_,
		_w567_
	);
	LUT2 #(
		.INIT('h1)
	) name553 (
		_w562_,
		_w567_,
		_w568_
	);
	LUT2 #(
		.INIT('h2)
	) name554 (
		_w46_,
		_w47_,
		_w569_
	);
	LUT2 #(
		.INIT('h4)
	) name555 (
		_w157_,
		_w569_,
		_w570_
	);
	LUT2 #(
		.INIT('h1)
	) name556 (
		_w568_,
		_w570_,
		_w571_
	);
	LUT2 #(
		.INIT('h4)
	) name557 (
		\v9_reg/NET0131 ,
		_w53_,
		_w572_
	);
	LUT2 #(
		.INIT('h1)
	) name558 (
		_w261_,
		_w572_,
		_w573_
	);
	LUT2 #(
		.INIT('h2)
	) name559 (
		_w209_,
		_w573_,
		_w574_
	);
	LUT2 #(
		.INIT('h1)
	) name560 (
		_w310_,
		_w545_,
		_w575_
	);
	LUT2 #(
		.INIT('h2)
	) name561 (
		\v9_reg/NET0131 ,
		_w345_,
		_w576_
	);
	LUT2 #(
		.INIT('h4)
	) name562 (
		_w575_,
		_w576_,
		_w577_
	);
	LUT2 #(
		.INIT('h1)
	) name563 (
		_w574_,
		_w577_,
		_w578_
	);
	LUT2 #(
		.INIT('h1)
	) name564 (
		\v12_reg/NET0131 ,
		_w578_,
		_w579_
	);
	assign \_al_n0  = 1'b0;
	assign \_al_n1  = 1'b0;
	assign \g1757/_0_  = _w85_ ;
	assign \g1763/_1_  = _w154_ ;
	assign \g1787/_3_  = _w174_ ;
	assign \g1800/_3_  = _w198_ ;
	assign \g1821/_2_  = _w206_ ;
	assign \g1940/_1_  = _w212_ ;
	assign \g25/_0_  = _w260_ ;
	assign \g2783/_3_  = _w283_ ;
	assign \g2823/_0_  = _w319_ ;
	assign \g38/_1_  = _w365_ ;
	assign \g40/_1_  = _w399_ ;
	assign \v13_D_11_pad  = _w413_ ;
	assign \v13_D_12_pad  = _w429_ ;
	assign \v13_D_13_pad  = _w455_ ;
	assign \v13_D_14_pad  = _w467_ ;
	assign \v13_D_16_pad  = _w470_ ;
	assign \v13_D_18_pad  = _w477_ ;
	assign \v13_D_19_pad  = _w484_ ;
	assign \v13_D_21_pad  = _w489_ ;
	assign \v13_D_22_pad  = _w496_ ;
	assign \v13_D_23_pad  = _w502_ ;
	assign \v13_D_24_pad  = _w528_ ;
	assign \v13_D_7_pad  = _w544_ ;
	assign \v13_D_8_pad  = _w571_ ;
	assign \v13_D_9_pad  = _w579_ ;
endmodule;