module top (\a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] , \a[17] , \a[18] , \a[19] , \a[20] , \a[21] , \a[22] , \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[30] , \a[31] , \a[32] , \a[33] , \a[34] , \a[35] , \a[36] , \a[37] , \a[38] , \a[39] , \a[40] , \a[41] , \a[42] , \a[43] , \a[44] , \a[45] , \a[46] , \a[47] , \a[48] , \a[49] , \a[50] , \a[51] , \a[52] , \a[53] , \a[54] , \a[55] , \a[56] , \a[57] , \a[58] , \a[59] , \a[60] , \a[61] , \a[62] , \a[63] , \a[64] , \a[65] , \a[66] , \a[67] , \a[68] , \a[69] , \a[70] , \a[71] , \a[72] , \a[73] , \a[74] , \a[75] , \a[76] , \a[77] , \a[78] , \a[79] , \a[80] , \a[81] , \a[82] , \a[83] , \a[84] , \a[85] , \a[86] , \a[87] , \a[88] , \a[89] , \a[90] , \a[91] , \a[92] , \a[93] , \a[94] , \a[95] , \a[96] , \a[97] , \a[98] , \a[99] , \a[100] , \a[101] , \a[102] , \a[103] , \a[104] , \a[105] , \a[106] , \a[107] , \a[108] , \a[109] , \a[110] , \a[111] , \a[112] , \a[113] , \a[114] , \a[115] , \a[116] , \a[117] , \a[118] , \a[119] , \a[120] , \a[121] , \a[122] , \a[123] , \a[124] , \a[125] , \a[126] , \a[127] , \b[0] , \b[1] , \b[2] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] , \b[17] , \b[18] , \b[19] , \b[20] , \b[21] , \b[22] , \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[30] , \b[31] , \b[32] , \b[33] , \b[34] , \b[35] , \b[36] , \b[37] , \b[38] , \b[39] , \b[40] , \b[41] , \b[42] , \b[43] , \b[44] , \b[45] , \b[46] , \b[47] , \b[48] , \b[49] , \b[50] , \b[51] , \b[52] , \b[53] , \b[54] , \b[55] , \b[56] , \b[57] , \b[58] , \b[59] , \b[60] , \b[61] , \b[62] , \b[63] , \b[64] , \b[65] , \b[66] , \b[67] , \b[68] , \b[69] , \b[70] , \b[71] , \b[72] , \b[73] , \b[74] , \b[75] , \b[76] , \b[77] , \b[78] , \b[79] , \b[80] , \b[81] , \b[82] , \b[83] , \b[84] , \b[85] , \b[86] , \b[87] , \b[88] , \b[89] , \b[90] , \b[91] , \b[92] , \b[93] , \b[94] , \b[95] , \b[96] , \b[97] , \b[98] , \b[99] , \b[100] , \b[101] , \b[102] , \b[103] , \b[104] , \b[105] , \b[106] , \b[107] , \b[108] , \b[109] , \b[110] , \b[111] , \b[112] , \b[113] , \b[114] , \b[115] , \b[116] , \b[117] , \b[118] , \b[119] , \b[120] , \b[121] , \b[122] , \b[123] , \b[124] , \b[125] , \b[126] , \b[127] , \f[0] , \f[1] , \f[2] , \f[3] , \f[4] , \f[5] , \f[6] , \f[7] , \f[8] , \f[9] , \f[10] , \f[11] , \f[12] , \f[13] , \f[14] , \f[15] , \f[16] , \f[17] , \f[18] , \f[19] , \f[20] , \f[21] , \f[22] , \f[23] , \f[24] , \f[25] , \f[26] , \f[27] , \f[28] , \f[29] , \f[30] , \f[31] , \f[32] , \f[33] , \f[34] , \f[35] , \f[36] , \f[37] , \f[38] , \f[39] , \f[40] , \f[41] , \f[42] , \f[43] , \f[44] , \f[45] , \f[46] , \f[47] , \f[48] , \f[49] , \f[50] , \f[51] , \f[52] , \f[53] , \f[54] , \f[55] , \f[56] , \f[57] , \f[58] , \f[59] , \f[60] , \f[61] , \f[62] , \f[63] , \f[64] , \f[65] , \f[66] , \f[67] , \f[68] , \f[69] , \f[70] , \f[71] , \f[72] , \f[73] , \f[74] , \f[75] , \f[76] , \f[77] , \f[78] , \f[79] , \f[80] , \f[81] , \f[82] , \f[83] , \f[84] , \f[85] , \f[86] , \f[87] , \f[88] , \f[89] , \f[90] , \f[91] , \f[92] , \f[93] , \f[94] , \f[95] , \f[96] , \f[97] , \f[98] , \f[99] , \f[100] , \f[101] , \f[102] , \f[103] , \f[104] , \f[105] , \f[106] , \f[107] , \f[108] , \f[109] , \f[110] , \f[111] , \f[112] , \f[113] , \f[114] , \f[115] , \f[116] , \f[117] , \f[118] , \f[119] , \f[120] , \f[121] , \f[122] , \f[123] , \f[124] , \f[125] , \f[126] , \f[127] , cOut);
	input \a[0]  ;
	input \a[1]  ;
	input \a[2]  ;
	input \a[3]  ;
	input \a[4]  ;
	input \a[5]  ;
	input \a[6]  ;
	input \a[7]  ;
	input \a[8]  ;
	input \a[9]  ;
	input \a[10]  ;
	input \a[11]  ;
	input \a[12]  ;
	input \a[13]  ;
	input \a[14]  ;
	input \a[15]  ;
	input \a[16]  ;
	input \a[17]  ;
	input \a[18]  ;
	input \a[19]  ;
	input \a[20]  ;
	input \a[21]  ;
	input \a[22]  ;
	input \a[23]  ;
	input \a[24]  ;
	input \a[25]  ;
	input \a[26]  ;
	input \a[27]  ;
	input \a[28]  ;
	input \a[29]  ;
	input \a[30]  ;
	input \a[31]  ;
	input \a[32]  ;
	input \a[33]  ;
	input \a[34]  ;
	input \a[35]  ;
	input \a[36]  ;
	input \a[37]  ;
	input \a[38]  ;
	input \a[39]  ;
	input \a[40]  ;
	input \a[41]  ;
	input \a[42]  ;
	input \a[43]  ;
	input \a[44]  ;
	input \a[45]  ;
	input \a[46]  ;
	input \a[47]  ;
	input \a[48]  ;
	input \a[49]  ;
	input \a[50]  ;
	input \a[51]  ;
	input \a[52]  ;
	input \a[53]  ;
	input \a[54]  ;
	input \a[55]  ;
	input \a[56]  ;
	input \a[57]  ;
	input \a[58]  ;
	input \a[59]  ;
	input \a[60]  ;
	input \a[61]  ;
	input \a[62]  ;
	input \a[63]  ;
	input \a[64]  ;
	input \a[65]  ;
	input \a[66]  ;
	input \a[67]  ;
	input \a[68]  ;
	input \a[69]  ;
	input \a[70]  ;
	input \a[71]  ;
	input \a[72]  ;
	input \a[73]  ;
	input \a[74]  ;
	input \a[75]  ;
	input \a[76]  ;
	input \a[77]  ;
	input \a[78]  ;
	input \a[79]  ;
	input \a[80]  ;
	input \a[81]  ;
	input \a[82]  ;
	input \a[83]  ;
	input \a[84]  ;
	input \a[85]  ;
	input \a[86]  ;
	input \a[87]  ;
	input \a[88]  ;
	input \a[89]  ;
	input \a[90]  ;
	input \a[91]  ;
	input \a[92]  ;
	input \a[93]  ;
	input \a[94]  ;
	input \a[95]  ;
	input \a[96]  ;
	input \a[97]  ;
	input \a[98]  ;
	input \a[99]  ;
	input \a[100]  ;
	input \a[101]  ;
	input \a[102]  ;
	input \a[103]  ;
	input \a[104]  ;
	input \a[105]  ;
	input \a[106]  ;
	input \a[107]  ;
	input \a[108]  ;
	input \a[109]  ;
	input \a[110]  ;
	input \a[111]  ;
	input \a[112]  ;
	input \a[113]  ;
	input \a[114]  ;
	input \a[115]  ;
	input \a[116]  ;
	input \a[117]  ;
	input \a[118]  ;
	input \a[119]  ;
	input \a[120]  ;
	input \a[121]  ;
	input \a[122]  ;
	input \a[123]  ;
	input \a[124]  ;
	input \a[125]  ;
	input \a[126]  ;
	input \a[127]  ;
	input \b[0]  ;
	input \b[1]  ;
	input \b[2]  ;
	input \b[3]  ;
	input \b[4]  ;
	input \b[5]  ;
	input \b[6]  ;
	input \b[7]  ;
	input \b[8]  ;
	input \b[9]  ;
	input \b[10]  ;
	input \b[11]  ;
	input \b[12]  ;
	input \b[13]  ;
	input \b[14]  ;
	input \b[15]  ;
	input \b[16]  ;
	input \b[17]  ;
	input \b[18]  ;
	input \b[19]  ;
	input \b[20]  ;
	input \b[21]  ;
	input \b[22]  ;
	input \b[23]  ;
	input \b[24]  ;
	input \b[25]  ;
	input \b[26]  ;
	input \b[27]  ;
	input \b[28]  ;
	input \b[29]  ;
	input \b[30]  ;
	input \b[31]  ;
	input \b[32]  ;
	input \b[33]  ;
	input \b[34]  ;
	input \b[35]  ;
	input \b[36]  ;
	input \b[37]  ;
	input \b[38]  ;
	input \b[39]  ;
	input \b[40]  ;
	input \b[41]  ;
	input \b[42]  ;
	input \b[43]  ;
	input \b[44]  ;
	input \b[45]  ;
	input \b[46]  ;
	input \b[47]  ;
	input \b[48]  ;
	input \b[49]  ;
	input \b[50]  ;
	input \b[51]  ;
	input \b[52]  ;
	input \b[53]  ;
	input \b[54]  ;
	input \b[55]  ;
	input \b[56]  ;
	input \b[57]  ;
	input \b[58]  ;
	input \b[59]  ;
	input \b[60]  ;
	input \b[61]  ;
	input \b[62]  ;
	input \b[63]  ;
	input \b[64]  ;
	input \b[65]  ;
	input \b[66]  ;
	input \b[67]  ;
	input \b[68]  ;
	input \b[69]  ;
	input \b[70]  ;
	input \b[71]  ;
	input \b[72]  ;
	input \b[73]  ;
	input \b[74]  ;
	input \b[75]  ;
	input \b[76]  ;
	input \b[77]  ;
	input \b[78]  ;
	input \b[79]  ;
	input \b[80]  ;
	input \b[81]  ;
	input \b[82]  ;
	input \b[83]  ;
	input \b[84]  ;
	input \b[85]  ;
	input \b[86]  ;
	input \b[87]  ;
	input \b[88]  ;
	input \b[89]  ;
	input \b[90]  ;
	input \b[91]  ;
	input \b[92]  ;
	input \b[93]  ;
	input \b[94]  ;
	input \b[95]  ;
	input \b[96]  ;
	input \b[97]  ;
	input \b[98]  ;
	input \b[99]  ;
	input \b[100]  ;
	input \b[101]  ;
	input \b[102]  ;
	input \b[103]  ;
	input \b[104]  ;
	input \b[105]  ;
	input \b[106]  ;
	input \b[107]  ;
	input \b[108]  ;
	input \b[109]  ;
	input \b[110]  ;
	input \b[111]  ;
	input \b[112]  ;
	input \b[113]  ;
	input \b[114]  ;
	input \b[115]  ;
	input \b[116]  ;
	input \b[117]  ;
	input \b[118]  ;
	input \b[119]  ;
	input \b[120]  ;
	input \b[121]  ;
	input \b[122]  ;
	input \b[123]  ;
	input \b[124]  ;
	input \b[125]  ;
	input \b[126]  ;
	input \b[127]  ;
	output \f[0]  ;
	output \f[1]  ;
	output \f[2]  ;
	output \f[3]  ;
	output \f[4]  ;
	output \f[5]  ;
	output \f[6]  ;
	output \f[7]  ;
	output \f[8]  ;
	output \f[9]  ;
	output \f[10]  ;
	output \f[11]  ;
	output \f[12]  ;
	output \f[13]  ;
	output \f[14]  ;
	output \f[15]  ;
	output \f[16]  ;
	output \f[17]  ;
	output \f[18]  ;
	output \f[19]  ;
	output \f[20]  ;
	output \f[21]  ;
	output \f[22]  ;
	output \f[23]  ;
	output \f[24]  ;
	output \f[25]  ;
	output \f[26]  ;
	output \f[27]  ;
	output \f[28]  ;
	output \f[29]  ;
	output \f[30]  ;
	output \f[31]  ;
	output \f[32]  ;
	output \f[33]  ;
	output \f[34]  ;
	output \f[35]  ;
	output \f[36]  ;
	output \f[37]  ;
	output \f[38]  ;
	output \f[39]  ;
	output \f[40]  ;
	output \f[41]  ;
	output \f[42]  ;
	output \f[43]  ;
	output \f[44]  ;
	output \f[45]  ;
	output \f[46]  ;
	output \f[47]  ;
	output \f[48]  ;
	output \f[49]  ;
	output \f[50]  ;
	output \f[51]  ;
	output \f[52]  ;
	output \f[53]  ;
	output \f[54]  ;
	output \f[55]  ;
	output \f[56]  ;
	output \f[57]  ;
	output \f[58]  ;
	output \f[59]  ;
	output \f[60]  ;
	output \f[61]  ;
	output \f[62]  ;
	output \f[63]  ;
	output \f[64]  ;
	output \f[65]  ;
	output \f[66]  ;
	output \f[67]  ;
	output \f[68]  ;
	output \f[69]  ;
	output \f[70]  ;
	output \f[71]  ;
	output \f[72]  ;
	output \f[73]  ;
	output \f[74]  ;
	output \f[75]  ;
	output \f[76]  ;
	output \f[77]  ;
	output \f[78]  ;
	output \f[79]  ;
	output \f[80]  ;
	output \f[81]  ;
	output \f[82]  ;
	output \f[83]  ;
	output \f[84]  ;
	output \f[85]  ;
	output \f[86]  ;
	output \f[87]  ;
	output \f[88]  ;
	output \f[89]  ;
	output \f[90]  ;
	output \f[91]  ;
	output \f[92]  ;
	output \f[93]  ;
	output \f[94]  ;
	output \f[95]  ;
	output \f[96]  ;
	output \f[97]  ;
	output \f[98]  ;
	output \f[99]  ;
	output \f[100]  ;
	output \f[101]  ;
	output \f[102]  ;
	output \f[103]  ;
	output \f[104]  ;
	output \f[105]  ;
	output \f[106]  ;
	output \f[107]  ;
	output \f[108]  ;
	output \f[109]  ;
	output \f[110]  ;
	output \f[111]  ;
	output \f[112]  ;
	output \f[113]  ;
	output \f[114]  ;
	output \f[115]  ;
	output \f[116]  ;
	output \f[117]  ;
	output \f[118]  ;
	output \f[119]  ;
	output \f[120]  ;
	output \f[121]  ;
	output \f[122]  ;
	output \f[123]  ;
	output \f[124]  ;
	output \f[125]  ;
	output \f[126]  ;
	output \f[127]  ;
	output cOut ;
	wire _w1136_ ;
	wire _w1135_ ;
	wire _w1134_ ;
	wire _w1133_ ;
	wire _w1132_ ;
	wire _w1131_ ;
	wire _w1130_ ;
	wire _w1129_ ;
	wire _w1128_ ;
	wire _w1127_ ;
	wire _w1126_ ;
	wire _w1125_ ;
	wire _w1124_ ;
	wire _w1123_ ;
	wire _w1122_ ;
	wire _w1121_ ;
	wire _w1120_ ;
	wire _w1119_ ;
	wire _w1118_ ;
	wire _w1117_ ;
	wire _w1116_ ;
	wire _w1115_ ;
	wire _w1114_ ;
	wire _w1113_ ;
	wire _w1112_ ;
	wire _w1111_ ;
	wire _w1110_ ;
	wire _w1109_ ;
	wire _w1108_ ;
	wire _w1107_ ;
	wire _w1106_ ;
	wire _w1105_ ;
	wire _w1104_ ;
	wire _w1103_ ;
	wire _w1102_ ;
	wire _w1101_ ;
	wire _w1100_ ;
	wire _w1099_ ;
	wire _w1098_ ;
	wire _w1097_ ;
	wire _w1096_ ;
	wire _w1095_ ;
	wire _w1094_ ;
	wire _w1093_ ;
	wire _w1092_ ;
	wire _w1091_ ;
	wire _w1090_ ;
	wire _w1089_ ;
	wire _w1088_ ;
	wire _w1087_ ;
	wire _w1086_ ;
	wire _w1085_ ;
	wire _w1084_ ;
	wire _w1083_ ;
	wire _w1082_ ;
	wire _w1081_ ;
	wire _w1080_ ;
	wire _w1079_ ;
	wire _w1078_ ;
	wire _w1077_ ;
	wire _w1076_ ;
	wire _w1075_ ;
	wire _w1074_ ;
	wire _w1073_ ;
	wire _w1072_ ;
	wire _w1071_ ;
	wire _w1070_ ;
	wire _w1069_ ;
	wire _w1068_ ;
	wire _w1067_ ;
	wire _w1066_ ;
	wire _w1065_ ;
	wire _w1064_ ;
	wire _w1063_ ;
	wire _w1062_ ;
	wire _w1061_ ;
	wire _w1060_ ;
	wire _w1059_ ;
	wire _w1058_ ;
	wire _w1057_ ;
	wire _w1056_ ;
	wire _w1055_ ;
	wire _w1054_ ;
	wire _w1053_ ;
	wire _w1052_ ;
	wire _w1051_ ;
	wire _w1050_ ;
	wire _w1049_ ;
	wire _w1048_ ;
	wire _w1047_ ;
	wire _w1046_ ;
	wire _w1045_ ;
	wire _w1044_ ;
	wire _w1043_ ;
	wire _w1042_ ;
	wire _w1041_ ;
	wire _w1040_ ;
	wire _w1039_ ;
	wire _w1038_ ;
	wire _w1037_ ;
	wire _w1036_ ;
	wire _w1035_ ;
	wire _w1034_ ;
	wire _w1033_ ;
	wire _w1032_ ;
	wire _w1031_ ;
	wire _w1030_ ;
	wire _w1029_ ;
	wire _w1028_ ;
	wire _w1027_ ;
	wire _w1026_ ;
	wire _w1025_ ;
	wire _w1024_ ;
	wire _w1023_ ;
	wire _w1022_ ;
	wire _w1021_ ;
	wire _w1020_ ;
	wire _w1019_ ;
	wire _w1018_ ;
	wire _w1017_ ;
	wire _w1016_ ;
	wire _w1015_ ;
	wire _w1014_ ;
	wire _w1013_ ;
	wire _w1012_ ;
	wire _w1011_ ;
	wire _w1010_ ;
	wire _w1009_ ;
	wire _w1008_ ;
	wire _w1007_ ;
	wire _w1006_ ;
	wire _w1005_ ;
	wire _w1004_ ;
	wire _w1003_ ;
	wire _w1002_ ;
	wire _w1001_ ;
	wire _w1000_ ;
	wire _w999_ ;
	wire _w998_ ;
	wire _w997_ ;
	wire _w996_ ;
	wire _w995_ ;
	wire _w994_ ;
	wire _w993_ ;
	wire _w992_ ;
	wire _w991_ ;
	wire _w990_ ;
	wire _w989_ ;
	wire _w988_ ;
	wire _w987_ ;
	wire _w986_ ;
	wire _w985_ ;
	wire _w984_ ;
	wire _w983_ ;
	wire _w982_ ;
	wire _w981_ ;
	wire _w980_ ;
	wire _w979_ ;
	wire _w978_ ;
	wire _w977_ ;
	wire _w976_ ;
	wire _w975_ ;
	wire _w974_ ;
	wire _w973_ ;
	wire _w972_ ;
	wire _w971_ ;
	wire _w970_ ;
	wire _w969_ ;
	wire _w968_ ;
	wire _w967_ ;
	wire _w966_ ;
	wire _w965_ ;
	wire _w964_ ;
	wire _w963_ ;
	wire _w962_ ;
	wire _w961_ ;
	wire _w960_ ;
	wire _w959_ ;
	wire _w958_ ;
	wire _w957_ ;
	wire _w956_ ;
	wire _w955_ ;
	wire _w954_ ;
	wire _w953_ ;
	wire _w952_ ;
	wire _w951_ ;
	wire _w950_ ;
	wire _w949_ ;
	wire _w948_ ;
	wire _w947_ ;
	wire _w946_ ;
	wire _w945_ ;
	wire _w944_ ;
	wire _w943_ ;
	wire _w942_ ;
	wire _w941_ ;
	wire _w940_ ;
	wire _w939_ ;
	wire _w938_ ;
	wire _w937_ ;
	wire _w936_ ;
	wire _w935_ ;
	wire _w934_ ;
	wire _w933_ ;
	wire _w932_ ;
	wire _w931_ ;
	wire _w930_ ;
	wire _w929_ ;
	wire _w928_ ;
	wire _w927_ ;
	wire _w926_ ;
	wire _w925_ ;
	wire _w924_ ;
	wire _w923_ ;
	wire _w922_ ;
	wire _w921_ ;
	wire _w920_ ;
	wire _w919_ ;
	wire _w918_ ;
	wire _w917_ ;
	wire _w916_ ;
	wire _w915_ ;
	wire _w914_ ;
	wire _w913_ ;
	wire _w912_ ;
	wire _w911_ ;
	wire _w910_ ;
	wire _w909_ ;
	wire _w908_ ;
	wire _w907_ ;
	wire _w906_ ;
	wire _w905_ ;
	wire _w904_ ;
	wire _w903_ ;
	wire _w902_ ;
	wire _w901_ ;
	wire _w900_ ;
	wire _w899_ ;
	wire _w898_ ;
	wire _w897_ ;
	wire _w896_ ;
	wire _w895_ ;
	wire _w894_ ;
	wire _w893_ ;
	wire _w892_ ;
	wire _w891_ ;
	wire _w890_ ;
	wire _w889_ ;
	wire _w888_ ;
	wire _w887_ ;
	wire _w886_ ;
	wire _w885_ ;
	wire _w884_ ;
	wire _w883_ ;
	wire _w882_ ;
	wire _w881_ ;
	wire _w880_ ;
	wire _w879_ ;
	wire _w878_ ;
	wire _w877_ ;
	wire _w876_ ;
	wire _w875_ ;
	wire _w874_ ;
	wire _w873_ ;
	wire _w872_ ;
	wire _w871_ ;
	wire _w870_ ;
	wire _w869_ ;
	wire _w868_ ;
	wire _w867_ ;
	wire _w866_ ;
	wire _w865_ ;
	wire _w864_ ;
	wire _w863_ ;
	wire _w862_ ;
	wire _w861_ ;
	wire _w860_ ;
	wire _w859_ ;
	wire _w858_ ;
	wire _w857_ ;
	wire _w856_ ;
	wire _w855_ ;
	wire _w854_ ;
	wire _w853_ ;
	wire _w852_ ;
	wire _w851_ ;
	wire _w850_ ;
	wire _w849_ ;
	wire _w848_ ;
	wire _w847_ ;
	wire _w846_ ;
	wire _w845_ ;
	wire _w844_ ;
	wire _w843_ ;
	wire _w842_ ;
	wire _w841_ ;
	wire _w840_ ;
	wire _w839_ ;
	wire _w838_ ;
	wire _w837_ ;
	wire _w836_ ;
	wire _w835_ ;
	wire _w834_ ;
	wire _w833_ ;
	wire _w832_ ;
	wire _w831_ ;
	wire _w830_ ;
	wire _w829_ ;
	wire _w828_ ;
	wire _w827_ ;
	wire _w826_ ;
	wire _w825_ ;
	wire _w824_ ;
	wire _w823_ ;
	wire _w822_ ;
	wire _w821_ ;
	wire _w820_ ;
	wire _w819_ ;
	wire _w818_ ;
	wire _w817_ ;
	wire _w816_ ;
	wire _w815_ ;
	wire _w814_ ;
	wire _w813_ ;
	wire _w812_ ;
	wire _w811_ ;
	wire _w810_ ;
	wire _w809_ ;
	wire _w808_ ;
	wire _w807_ ;
	wire _w806_ ;
	wire _w805_ ;
	wire _w804_ ;
	wire _w803_ ;
	wire _w802_ ;
	wire _w801_ ;
	wire _w800_ ;
	wire _w799_ ;
	wire _w514_ ;
	wire _w513_ ;
	wire _w512_ ;
	wire _w511_ ;
	wire _w510_ ;
	wire _w509_ ;
	wire _w508_ ;
	wire _w507_ ;
	wire _w506_ ;
	wire _w505_ ;
	wire _w504_ ;
	wire _w503_ ;
	wire _w502_ ;
	wire _w501_ ;
	wire _w500_ ;
	wire _w499_ ;
	wire _w498_ ;
	wire _w497_ ;
	wire _w496_ ;
	wire _w495_ ;
	wire _w494_ ;
	wire _w493_ ;
	wire _w492_ ;
	wire _w491_ ;
	wire _w490_ ;
	wire _w489_ ;
	wire _w488_ ;
	wire _w487_ ;
	wire _w486_ ;
	wire _w485_ ;
	wire _w484_ ;
	wire _w483_ ;
	wire _w482_ ;
	wire _w481_ ;
	wire _w480_ ;
	wire _w479_ ;
	wire _w478_ ;
	wire _w477_ ;
	wire _w476_ ;
	wire _w475_ ;
	wire _w474_ ;
	wire _w473_ ;
	wire _w472_ ;
	wire _w471_ ;
	wire _w470_ ;
	wire _w469_ ;
	wire _w468_ ;
	wire _w467_ ;
	wire _w466_ ;
	wire _w465_ ;
	wire _w464_ ;
	wire _w463_ ;
	wire _w462_ ;
	wire _w461_ ;
	wire _w460_ ;
	wire _w459_ ;
	wire _w458_ ;
	wire _w457_ ;
	wire _w456_ ;
	wire _w455_ ;
	wire _w454_ ;
	wire _w453_ ;
	wire _w452_ ;
	wire _w451_ ;
	wire _w450_ ;
	wire _w449_ ;
	wire _w448_ ;
	wire _w447_ ;
	wire _w446_ ;
	wire _w445_ ;
	wire _w444_ ;
	wire _w443_ ;
	wire _w442_ ;
	wire _w441_ ;
	wire _w440_ ;
	wire _w439_ ;
	wire _w438_ ;
	wire _w437_ ;
	wire _w436_ ;
	wire _w435_ ;
	wire _w434_ ;
	wire _w433_ ;
	wire _w432_ ;
	wire _w431_ ;
	wire _w430_ ;
	wire _w429_ ;
	wire _w428_ ;
	wire _w427_ ;
	wire _w426_ ;
	wire _w425_ ;
	wire _w424_ ;
	wire _w423_ ;
	wire _w422_ ;
	wire _w421_ ;
	wire _w420_ ;
	wire _w419_ ;
	wire _w418_ ;
	wire _w417_ ;
	wire _w416_ ;
	wire _w415_ ;
	wire _w414_ ;
	wire _w413_ ;
	wire _w412_ ;
	wire _w411_ ;
	wire _w410_ ;
	wire _w409_ ;
	wire _w408_ ;
	wire _w407_ ;
	wire _w406_ ;
	wire _w405_ ;
	wire _w404_ ;
	wire _w403_ ;
	wire _w402_ ;
	wire _w401_ ;
	wire _w400_ ;
	wire _w399_ ;
	wire _w398_ ;
	wire _w397_ ;
	wire _w396_ ;
	wire _w395_ ;
	wire _w394_ ;
	wire _w393_ ;
	wire _w392_ ;
	wire _w391_ ;
	wire _w390_ ;
	wire _w389_ ;
	wire _w388_ ;
	wire _w387_ ;
	wire _w386_ ;
	wire _w385_ ;
	wire _w316_ ;
	wire _w315_ ;
	wire _w314_ ;
	wire _w313_ ;
	wire _w312_ ;
	wire _w311_ ;
	wire _w310_ ;
	wire _w309_ ;
	wire _w308_ ;
	wire _w307_ ;
	wire _w306_ ;
	wire _w305_ ;
	wire _w304_ ;
	wire _w303_ ;
	wire _w302_ ;
	wire _w301_ ;
	wire _w300_ ;
	wire _w299_ ;
	wire _w298_ ;
	wire _w297_ ;
	wire _w296_ ;
	wire _w295_ ;
	wire _w294_ ;
	wire _w293_ ;
	wire _w292_ ;
	wire _w291_ ;
	wire _w290_ ;
	wire _w289_ ;
	wire _w288_ ;
	wire _w287_ ;
	wire _w270_ ;
	wire _w269_ ;
	wire _w268_ ;
	wire _w267_ ;
	wire _w266_ ;
	wire _w265_ ;
	wire _w264_ ;
	wire _w263_ ;
	wire _w262_ ;
	wire _w261_ ;
	wire _w260_ ;
	wire _w259_ ;
	wire _w258_ ;
	wire _w271_ ;
	wire _w272_ ;
	wire _w273_ ;
	wire _w274_ ;
	wire _w275_ ;
	wire _w276_ ;
	wire _w277_ ;
	wire _w278_ ;
	wire _w279_ ;
	wire _w280_ ;
	wire _w281_ ;
	wire _w282_ ;
	wire _w283_ ;
	wire _w284_ ;
	wire _w285_ ;
	wire _w286_ ;
	wire _w317_ ;
	wire _w318_ ;
	wire _w319_ ;
	wire _w320_ ;
	wire _w321_ ;
	wire _w322_ ;
	wire _w323_ ;
	wire _w324_ ;
	wire _w325_ ;
	wire _w326_ ;
	wire _w327_ ;
	wire _w328_ ;
	wire _w329_ ;
	wire _w330_ ;
	wire _w331_ ;
	wire _w332_ ;
	wire _w333_ ;
	wire _w334_ ;
	wire _w335_ ;
	wire _w336_ ;
	wire _w337_ ;
	wire _w338_ ;
	wire _w339_ ;
	wire _w340_ ;
	wire _w341_ ;
	wire _w342_ ;
	wire _w343_ ;
	wire _w344_ ;
	wire _w345_ ;
	wire _w346_ ;
	wire _w347_ ;
	wire _w348_ ;
	wire _w349_ ;
	wire _w350_ ;
	wire _w351_ ;
	wire _w352_ ;
	wire _w353_ ;
	wire _w354_ ;
	wire _w355_ ;
	wire _w356_ ;
	wire _w357_ ;
	wire _w358_ ;
	wire _w359_ ;
	wire _w360_ ;
	wire _w361_ ;
	wire _w362_ ;
	wire _w363_ ;
	wire _w364_ ;
	wire _w365_ ;
	wire _w366_ ;
	wire _w367_ ;
	wire _w368_ ;
	wire _w369_ ;
	wire _w370_ ;
	wire _w371_ ;
	wire _w372_ ;
	wire _w373_ ;
	wire _w374_ ;
	wire _w375_ ;
	wire _w376_ ;
	wire _w377_ ;
	wire _w378_ ;
	wire _w379_ ;
	wire _w380_ ;
	wire _w381_ ;
	wire _w382_ ;
	wire _w383_ ;
	wire _w384_ ;
	wire _w515_ ;
	wire _w516_ ;
	wire _w517_ ;
	wire _w518_ ;
	wire _w519_ ;
	wire _w520_ ;
	wire _w521_ ;
	wire _w522_ ;
	wire _w523_ ;
	wire _w524_ ;
	wire _w525_ ;
	wire _w526_ ;
	wire _w527_ ;
	wire _w528_ ;
	wire _w529_ ;
	wire _w530_ ;
	wire _w531_ ;
	wire _w532_ ;
	wire _w533_ ;
	wire _w534_ ;
	wire _w535_ ;
	wire _w536_ ;
	wire _w537_ ;
	wire _w538_ ;
	wire _w539_ ;
	wire _w540_ ;
	wire _w541_ ;
	wire _w542_ ;
	wire _w543_ ;
	wire _w544_ ;
	wire _w545_ ;
	wire _w546_ ;
	wire _w547_ ;
	wire _w548_ ;
	wire _w549_ ;
	wire _w550_ ;
	wire _w551_ ;
	wire _w552_ ;
	wire _w553_ ;
	wire _w554_ ;
	wire _w555_ ;
	wire _w556_ ;
	wire _w557_ ;
	wire _w558_ ;
	wire _w559_ ;
	wire _w560_ ;
	wire _w561_ ;
	wire _w562_ ;
	wire _w563_ ;
	wire _w564_ ;
	wire _w565_ ;
	wire _w566_ ;
	wire _w567_ ;
	wire _w568_ ;
	wire _w569_ ;
	wire _w570_ ;
	wire _w571_ ;
	wire _w572_ ;
	wire _w573_ ;
	wire _w574_ ;
	wire _w575_ ;
	wire _w576_ ;
	wire _w577_ ;
	wire _w578_ ;
	wire _w579_ ;
	wire _w580_ ;
	wire _w581_ ;
	wire _w582_ ;
	wire _w583_ ;
	wire _w584_ ;
	wire _w585_ ;
	wire _w586_ ;
	wire _w587_ ;
	wire _w588_ ;
	wire _w589_ ;
	wire _w590_ ;
	wire _w591_ ;
	wire _w592_ ;
	wire _w593_ ;
	wire _w594_ ;
	wire _w595_ ;
	wire _w596_ ;
	wire _w597_ ;
	wire _w598_ ;
	wire _w599_ ;
	wire _w600_ ;
	wire _w601_ ;
	wire _w602_ ;
	wire _w603_ ;
	wire _w604_ ;
	wire _w605_ ;
	wire _w606_ ;
	wire _w607_ ;
	wire _w608_ ;
	wire _w609_ ;
	wire _w610_ ;
	wire _w611_ ;
	wire _w612_ ;
	wire _w613_ ;
	wire _w614_ ;
	wire _w615_ ;
	wire _w616_ ;
	wire _w617_ ;
	wire _w618_ ;
	wire _w619_ ;
	wire _w620_ ;
	wire _w621_ ;
	wire _w622_ ;
	wire _w623_ ;
	wire _w624_ ;
	wire _w625_ ;
	wire _w626_ ;
	wire _w627_ ;
	wire _w628_ ;
	wire _w629_ ;
	wire _w630_ ;
	wire _w631_ ;
	wire _w632_ ;
	wire _w633_ ;
	wire _w634_ ;
	wire _w635_ ;
	wire _w636_ ;
	wire _w637_ ;
	wire _w638_ ;
	wire _w639_ ;
	wire _w640_ ;
	wire _w641_ ;
	wire _w642_ ;
	wire _w643_ ;
	wire _w644_ ;
	wire _w645_ ;
	wire _w646_ ;
	wire _w647_ ;
	wire _w648_ ;
	wire _w649_ ;
	wire _w650_ ;
	wire _w651_ ;
	wire _w652_ ;
	wire _w653_ ;
	wire _w654_ ;
	wire _w655_ ;
	wire _w656_ ;
	wire _w657_ ;
	wire _w658_ ;
	wire _w659_ ;
	wire _w660_ ;
	wire _w661_ ;
	wire _w662_ ;
	wire _w663_ ;
	wire _w664_ ;
	wire _w665_ ;
	wire _w666_ ;
	wire _w667_ ;
	wire _w668_ ;
	wire _w669_ ;
	wire _w670_ ;
	wire _w671_ ;
	wire _w672_ ;
	wire _w673_ ;
	wire _w674_ ;
	wire _w675_ ;
	wire _w676_ ;
	wire _w677_ ;
	wire _w678_ ;
	wire _w679_ ;
	wire _w680_ ;
	wire _w681_ ;
	wire _w682_ ;
	wire _w683_ ;
	wire _w684_ ;
	wire _w685_ ;
	wire _w686_ ;
	wire _w687_ ;
	wire _w688_ ;
	wire _w689_ ;
	wire _w690_ ;
	wire _w691_ ;
	wire _w692_ ;
	wire _w693_ ;
	wire _w694_ ;
	wire _w695_ ;
	wire _w696_ ;
	wire _w697_ ;
	wire _w698_ ;
	wire _w699_ ;
	wire _w700_ ;
	wire _w701_ ;
	wire _w702_ ;
	wire _w703_ ;
	wire _w704_ ;
	wire _w705_ ;
	wire _w706_ ;
	wire _w707_ ;
	wire _w708_ ;
	wire _w709_ ;
	wire _w710_ ;
	wire _w711_ ;
	wire _w712_ ;
	wire _w713_ ;
	wire _w714_ ;
	wire _w715_ ;
	wire _w716_ ;
	wire _w717_ ;
	wire _w718_ ;
	wire _w719_ ;
	wire _w720_ ;
	wire _w721_ ;
	wire _w722_ ;
	wire _w723_ ;
	wire _w724_ ;
	wire _w725_ ;
	wire _w726_ ;
	wire _w727_ ;
	wire _w728_ ;
	wire _w729_ ;
	wire _w730_ ;
	wire _w731_ ;
	wire _w732_ ;
	wire _w733_ ;
	wire _w734_ ;
	wire _w735_ ;
	wire _w736_ ;
	wire _w737_ ;
	wire _w738_ ;
	wire _w739_ ;
	wire _w740_ ;
	wire _w741_ ;
	wire _w742_ ;
	wire _w743_ ;
	wire _w744_ ;
	wire _w745_ ;
	wire _w746_ ;
	wire _w747_ ;
	wire _w748_ ;
	wire _w749_ ;
	wire _w750_ ;
	wire _w751_ ;
	wire _w752_ ;
	wire _w753_ ;
	wire _w754_ ;
	wire _w755_ ;
	wire _w756_ ;
	wire _w757_ ;
	wire _w758_ ;
	wire _w759_ ;
	wire _w760_ ;
	wire _w761_ ;
	wire _w762_ ;
	wire _w763_ ;
	wire _w764_ ;
	wire _w765_ ;
	wire _w766_ ;
	wire _w767_ ;
	wire _w768_ ;
	wire _w769_ ;
	wire _w770_ ;
	wire _w771_ ;
	wire _w772_ ;
	wire _w773_ ;
	wire _w774_ ;
	wire _w775_ ;
	wire _w776_ ;
	wire _w777_ ;
	wire _w778_ ;
	wire _w779_ ;
	wire _w780_ ;
	wire _w781_ ;
	wire _w782_ ;
	wire _w783_ ;
	wire _w784_ ;
	wire _w785_ ;
	wire _w786_ ;
	wire _w787_ ;
	wire _w788_ ;
	wire _w789_ ;
	wire _w790_ ;
	wire _w791_ ;
	wire _w792_ ;
	wire _w793_ ;
	wire _w794_ ;
	wire _w795_ ;
	wire _w796_ ;
	wire _w797_ ;
	wire _w798_ ;
	LUT2 #(
		.INIT('h6)
	) name0 (
		\a[0] ,
		\b[0] ,
		_w258_
	);
	LUT4 #(
		.INIT('h936c)
	) name1 (
		\a[0] ,
		\a[1] ,
		\b[0] ,
		\b[1] ,
		_w259_
	);
	LUT2 #(
		.INIT('h8)
	) name2 (
		\a[2] ,
		\b[2] ,
		_w260_
	);
	LUT2 #(
		.INIT('h6)
	) name3 (
		\a[2] ,
		\b[2] ,
		_w261_
	);
	LUT4 #(
		.INIT('h135f)
	) name4 (
		\a[0] ,
		\a[1] ,
		\b[0] ,
		\b[1] ,
		_w262_
	);
	LUT4 #(
		.INIT('hec80)
	) name5 (
		\a[0] ,
		\a[1] ,
		\b[0] ,
		\b[1] ,
		_w263_
	);
	LUT2 #(
		.INIT('h6)
	) name6 (
		_w261_,
		_w263_,
		_w264_
	);
	LUT2 #(
		.INIT('h6)
	) name7 (
		\a[3] ,
		\b[3] ,
		_w265_
	);
	LUT4 #(
		.INIT('hfac8)
	) name8 (
		\a[1] ,
		\a[2] ,
		\b[1] ,
		\b[2] ,
		_w266_
	);
	LUT4 #(
		.INIT('h4b5a)
	) name9 (
		_w260_,
		_w262_,
		_w265_,
		_w266_,
		_w267_
	);
	LUT4 #(
		.INIT('h135f)
	) name10 (
		\a[2] ,
		\a[3] ,
		\b[2] ,
		\b[3] ,
		_w268_
	);
	LUT2 #(
		.INIT('h1)
	) name11 (
		\a[4] ,
		\b[4] ,
		_w269_
	);
	LUT2 #(
		.INIT('h8)
	) name12 (
		\a[4] ,
		\b[4] ,
		_w270_
	);
	LUT2 #(
		.INIT('h6)
	) name13 (
		\a[4] ,
		\b[4] ,
		_w271_
	);
	LUT4 #(
		.INIT('hc832)
	) name14 (
		\a[3] ,
		\a[4] ,
		\b[3] ,
		\b[4] ,
		_w272_
	);
	LUT4 #(
		.INIT('h4f00)
	) name15 (
		_w262_,
		_w266_,
		_w268_,
		_w272_,
		_w273_
	);
	LUT4 #(
		.INIT('h0104)
	) name16 (
		\a[3] ,
		\a[4] ,
		\b[3] ,
		\b[4] ,
		_w274_
	);
	LUT4 #(
		.INIT('hb000)
	) name17 (
		_w262_,
		_w266_,
		_w268_,
		_w271_,
		_w275_
	);
	LUT3 #(
		.INIT('hfe)
	) name18 (
		_w273_,
		_w274_,
		_w275_,
		_w276_
	);
	LUT4 #(
		.INIT('h00b0)
	) name19 (
		_w262_,
		_w266_,
		_w268_,
		_w270_,
		_w277_
	);
	LUT4 #(
		.INIT('h0105)
	) name20 (
		\a[3] ,
		\a[4] ,
		\b[3] ,
		\b[4] ,
		_w278_
	);
	LUT2 #(
		.INIT('h8)
	) name21 (
		\a[5] ,
		\b[5] ,
		_w279_
	);
	LUT2 #(
		.INIT('h6)
	) name22 (
		\a[5] ,
		\b[5] ,
		_w280_
	);
	LUT4 #(
		.INIT('hfe01)
	) name23 (
		_w269_,
		_w277_,
		_w278_,
		_w280_,
		_w281_
	);
	LUT2 #(
		.INIT('h6)
	) name24 (
		\a[6] ,
		\b[6] ,
		_w282_
	);
	LUT4 #(
		.INIT('hfac8)
	) name25 (
		\a[4] ,
		\a[5] ,
		\b[4] ,
		\b[5] ,
		_w283_
	);
	LUT2 #(
		.INIT('h4)
	) name26 (
		_w278_,
		_w283_,
		_w284_
	);
	LUT4 #(
		.INIT('h2d3c)
	) name27 (
		_w277_,
		_w279_,
		_w282_,
		_w284_,
		_w285_
	);
	LUT4 #(
		.INIT('h135f)
	) name28 (
		\a[5] ,
		\a[6] ,
		\b[5] ,
		\b[6] ,
		_w286_
	);
	LUT2 #(
		.INIT('h8)
	) name29 (
		\a[7] ,
		\b[7] ,
		_w287_
	);
	LUT2 #(
		.INIT('h6)
	) name30 (
		\a[7] ,
		\b[7] ,
		_w288_
	);
	LUT4 #(
		.INIT('hc832)
	) name31 (
		\a[6] ,
		\a[7] ,
		\b[6] ,
		\b[7] ,
		_w289_
	);
	LUT4 #(
		.INIT('h4f00)
	) name32 (
		_w277_,
		_w284_,
		_w286_,
		_w289_,
		_w290_
	);
	LUT4 #(
		.INIT('h0104)
	) name33 (
		\a[6] ,
		\a[7] ,
		\b[6] ,
		\b[7] ,
		_w291_
	);
	LUT2 #(
		.INIT('h8)
	) name34 (
		_w286_,
		_w288_,
		_w292_
	);
	LUT4 #(
		.INIT('h040f)
	) name35 (
		_w277_,
		_w284_,
		_w291_,
		_w292_,
		_w293_
	);
	LUT2 #(
		.INIT('hb)
	) name36 (
		_w290_,
		_w293_,
		_w294_
	);
	LUT2 #(
		.INIT('h2)
	) name37 (
		_w286_,
		_w287_,
		_w295_
	);
	LUT4 #(
		.INIT('h0105)
	) name38 (
		\a[6] ,
		\a[7] ,
		\b[6] ,
		\b[7] ,
		_w296_
	);
	LUT2 #(
		.INIT('h8)
	) name39 (
		\a[8] ,
		\b[8] ,
		_w297_
	);
	LUT2 #(
		.INIT('h6)
	) name40 (
		\a[8] ,
		\b[8] ,
		_w298_
	);
	LUT4 #(
		.INIT('hc832)
	) name41 (
		\a[7] ,
		\a[8] ,
		\b[7] ,
		\b[8] ,
		_w299_
	);
	LUT2 #(
		.INIT('h4)
	) name42 (
		_w296_,
		_w299_,
		_w300_
	);
	LUT4 #(
		.INIT('h4f00)
	) name43 (
		_w277_,
		_w284_,
		_w295_,
		_w300_,
		_w301_
	);
	LUT4 #(
		.INIT('hfec8)
	) name44 (
		\a[6] ,
		\a[7] ,
		\b[6] ,
		\b[7] ,
		_w302_
	);
	LUT4 #(
		.INIT('h4f00)
	) name45 (
		_w277_,
		_w284_,
		_w295_,
		_w302_,
		_w303_
	);
	LUT3 #(
		.INIT('hce)
	) name46 (
		_w298_,
		_w301_,
		_w303_,
		_w304_
	);
	LUT2 #(
		.INIT('h1)
	) name47 (
		\a[9] ,
		\b[9] ,
		_w305_
	);
	LUT2 #(
		.INIT('h6)
	) name48 (
		\a[9] ,
		\b[9] ,
		_w306_
	);
	LUT4 #(
		.INIT('hfac8)
	) name49 (
		\a[7] ,
		\a[8] ,
		\b[7] ,
		\b[8] ,
		_w307_
	);
	LUT2 #(
		.INIT('h4)
	) name50 (
		_w296_,
		_w307_,
		_w308_
	);
	LUT4 #(
		.INIT('h4f00)
	) name51 (
		_w277_,
		_w284_,
		_w295_,
		_w308_,
		_w309_
	);
	LUT3 #(
		.INIT('h36)
	) name52 (
		_w297_,
		_w306_,
		_w309_,
		_w310_
	);
	LUT4 #(
		.INIT('h135f)
	) name53 (
		\a[8] ,
		\a[9] ,
		\b[8] ,
		\b[9] ,
		_w311_
	);
	LUT2 #(
		.INIT('h8)
	) name54 (
		\a[10] ,
		\b[10] ,
		_w312_
	);
	LUT2 #(
		.INIT('h6)
	) name55 (
		\a[10] ,
		\b[10] ,
		_w313_
	);
	LUT4 #(
		.INIT('hba45)
	) name56 (
		_w305_,
		_w309_,
		_w311_,
		_w313_,
		_w314_
	);
	LUT2 #(
		.INIT('h2)
	) name57 (
		_w311_,
		_w312_,
		_w315_
	);
	LUT4 #(
		.INIT('h0105)
	) name58 (
		\a[9] ,
		\a[10] ,
		\b[9] ,
		\b[10] ,
		_w316_
	);
	LUT2 #(
		.INIT('h8)
	) name59 (
		\a[11] ,
		\b[11] ,
		_w317_
	);
	LUT2 #(
		.INIT('h6)
	) name60 (
		\a[11] ,
		\b[11] ,
		_w318_
	);
	LUT4 #(
		.INIT('hc832)
	) name61 (
		\a[10] ,
		\a[11] ,
		\b[10] ,
		\b[11] ,
		_w319_
	);
	LUT2 #(
		.INIT('h4)
	) name62 (
		_w316_,
		_w319_,
		_w320_
	);
	LUT3 #(
		.INIT('hb0)
	) name63 (
		_w309_,
		_w315_,
		_w320_,
		_w321_
	);
	LUT4 #(
		.INIT('hfec8)
	) name64 (
		\a[9] ,
		\a[10] ,
		\b[9] ,
		\b[10] ,
		_w322_
	);
	LUT4 #(
		.INIT('h40f0)
	) name65 (
		_w309_,
		_w315_,
		_w318_,
		_w322_,
		_w323_
	);
	LUT2 #(
		.INIT('he)
	) name66 (
		_w321_,
		_w323_,
		_w324_
	);
	LUT2 #(
		.INIT('h1)
	) name67 (
		\a[12] ,
		\b[12] ,
		_w325_
	);
	LUT2 #(
		.INIT('h6)
	) name68 (
		\a[12] ,
		\b[12] ,
		_w326_
	);
	LUT4 #(
		.INIT('hfac8)
	) name69 (
		\a[10] ,
		\a[11] ,
		\b[10] ,
		\b[11] ,
		_w327_
	);
	LUT2 #(
		.INIT('h4)
	) name70 (
		_w316_,
		_w327_,
		_w328_
	);
	LUT3 #(
		.INIT('hb0)
	) name71 (
		_w309_,
		_w315_,
		_w328_,
		_w329_
	);
	LUT3 #(
		.INIT('h36)
	) name72 (
		_w317_,
		_w326_,
		_w329_,
		_w330_
	);
	LUT4 #(
		.INIT('h135f)
	) name73 (
		\a[11] ,
		\a[12] ,
		\b[11] ,
		\b[12] ,
		_w331_
	);
	LUT4 #(
		.INIT('h4f00)
	) name74 (
		_w309_,
		_w315_,
		_w328_,
		_w331_,
		_w332_
	);
	LUT2 #(
		.INIT('h1)
	) name75 (
		\a[13] ,
		\b[13] ,
		_w333_
	);
	LUT2 #(
		.INIT('h8)
	) name76 (
		\a[13] ,
		\b[13] ,
		_w334_
	);
	LUT2 #(
		.INIT('h6)
	) name77 (
		\a[13] ,
		\b[13] ,
		_w335_
	);
	LUT2 #(
		.INIT('h8)
	) name78 (
		_w331_,
		_w335_,
		_w336_
	);
	LUT4 #(
		.INIT('h4f00)
	) name79 (
		_w309_,
		_w315_,
		_w328_,
		_w336_,
		_w337_
	);
	LUT4 #(
		.INIT('hffa1)
	) name80 (
		_w325_,
		_w332_,
		_w335_,
		_w337_,
		_w338_
	);
	LUT2 #(
		.INIT('h2)
	) name81 (
		_w331_,
		_w334_,
		_w339_
	);
	LUT4 #(
		.INIT('h4f00)
	) name82 (
		_w309_,
		_w315_,
		_w328_,
		_w339_,
		_w340_
	);
	LUT4 #(
		.INIT('h0105)
	) name83 (
		\a[12] ,
		\a[13] ,
		\b[12] ,
		\b[13] ,
		_w341_
	);
	LUT2 #(
		.INIT('h8)
	) name84 (
		\a[14] ,
		\b[14] ,
		_w342_
	);
	LUT2 #(
		.INIT('h6)
	) name85 (
		\a[14] ,
		\b[14] ,
		_w343_
	);
	LUT4 #(
		.INIT('hfe01)
	) name86 (
		_w333_,
		_w340_,
		_w341_,
		_w343_,
		_w344_
	);
	LUT2 #(
		.INIT('h6)
	) name87 (
		\a[15] ,
		\b[15] ,
		_w345_
	);
	LUT4 #(
		.INIT('hfac8)
	) name88 (
		\a[13] ,
		\a[14] ,
		\b[13] ,
		\b[14] ,
		_w346_
	);
	LUT2 #(
		.INIT('h4)
	) name89 (
		_w341_,
		_w346_,
		_w347_
	);
	LUT4 #(
		.INIT('h2d3c)
	) name90 (
		_w340_,
		_w342_,
		_w345_,
		_w347_,
		_w348_
	);
	LUT4 #(
		.INIT('h135f)
	) name91 (
		\a[14] ,
		\a[15] ,
		\b[14] ,
		\b[15] ,
		_w349_
	);
	LUT2 #(
		.INIT('h8)
	) name92 (
		\a[16] ,
		\b[16] ,
		_w350_
	);
	LUT2 #(
		.INIT('h6)
	) name93 (
		\a[16] ,
		\b[16] ,
		_w351_
	);
	LUT4 #(
		.INIT('hc832)
	) name94 (
		\a[15] ,
		\a[16] ,
		\b[15] ,
		\b[16] ,
		_w352_
	);
	LUT4 #(
		.INIT('h4f00)
	) name95 (
		_w340_,
		_w347_,
		_w349_,
		_w352_,
		_w353_
	);
	LUT4 #(
		.INIT('h0104)
	) name96 (
		\a[15] ,
		\a[16] ,
		\b[15] ,
		\b[16] ,
		_w354_
	);
	LUT2 #(
		.INIT('h8)
	) name97 (
		_w349_,
		_w351_,
		_w355_
	);
	LUT4 #(
		.INIT('h040f)
	) name98 (
		_w340_,
		_w347_,
		_w354_,
		_w355_,
		_w356_
	);
	LUT2 #(
		.INIT('hb)
	) name99 (
		_w353_,
		_w356_,
		_w357_
	);
	LUT2 #(
		.INIT('h2)
	) name100 (
		_w349_,
		_w350_,
		_w358_
	);
	LUT4 #(
		.INIT('h0105)
	) name101 (
		\a[15] ,
		\a[16] ,
		\b[15] ,
		\b[16] ,
		_w359_
	);
	LUT2 #(
		.INIT('h8)
	) name102 (
		\a[17] ,
		\b[17] ,
		_w360_
	);
	LUT2 #(
		.INIT('h6)
	) name103 (
		\a[17] ,
		\b[17] ,
		_w361_
	);
	LUT4 #(
		.INIT('hc832)
	) name104 (
		\a[16] ,
		\a[17] ,
		\b[16] ,
		\b[17] ,
		_w362_
	);
	LUT2 #(
		.INIT('h4)
	) name105 (
		_w359_,
		_w362_,
		_w363_
	);
	LUT4 #(
		.INIT('h4f00)
	) name106 (
		_w340_,
		_w347_,
		_w358_,
		_w363_,
		_w364_
	);
	LUT4 #(
		.INIT('hfec8)
	) name107 (
		\a[15] ,
		\a[16] ,
		\b[15] ,
		\b[16] ,
		_w365_
	);
	LUT4 #(
		.INIT('h4f00)
	) name108 (
		_w340_,
		_w347_,
		_w358_,
		_w365_,
		_w366_
	);
	LUT3 #(
		.INIT('hce)
	) name109 (
		_w361_,
		_w364_,
		_w366_,
		_w367_
	);
	LUT2 #(
		.INIT('h1)
	) name110 (
		\a[18] ,
		\b[18] ,
		_w368_
	);
	LUT2 #(
		.INIT('h6)
	) name111 (
		\a[18] ,
		\b[18] ,
		_w369_
	);
	LUT4 #(
		.INIT('hfac8)
	) name112 (
		\a[16] ,
		\a[17] ,
		\b[16] ,
		\b[17] ,
		_w370_
	);
	LUT2 #(
		.INIT('h4)
	) name113 (
		_w359_,
		_w370_,
		_w371_
	);
	LUT4 #(
		.INIT('h4f00)
	) name114 (
		_w340_,
		_w347_,
		_w358_,
		_w371_,
		_w372_
	);
	LUT3 #(
		.INIT('h36)
	) name115 (
		_w360_,
		_w369_,
		_w372_,
		_w373_
	);
	LUT4 #(
		.INIT('h135f)
	) name116 (
		\a[17] ,
		\a[18] ,
		\b[17] ,
		\b[18] ,
		_w374_
	);
	LUT2 #(
		.INIT('h8)
	) name117 (
		\a[19] ,
		\b[19] ,
		_w375_
	);
	LUT2 #(
		.INIT('h6)
	) name118 (
		\a[19] ,
		\b[19] ,
		_w376_
	);
	LUT4 #(
		.INIT('hba45)
	) name119 (
		_w368_,
		_w372_,
		_w374_,
		_w376_,
		_w377_
	);
	LUT2 #(
		.INIT('h2)
	) name120 (
		_w374_,
		_w375_,
		_w378_
	);
	LUT4 #(
		.INIT('h0105)
	) name121 (
		\a[18] ,
		\a[19] ,
		\b[18] ,
		\b[19] ,
		_w379_
	);
	LUT2 #(
		.INIT('h8)
	) name122 (
		\a[20] ,
		\b[20] ,
		_w380_
	);
	LUT2 #(
		.INIT('h6)
	) name123 (
		\a[20] ,
		\b[20] ,
		_w381_
	);
	LUT4 #(
		.INIT('hc832)
	) name124 (
		\a[19] ,
		\a[20] ,
		\b[19] ,
		\b[20] ,
		_w382_
	);
	LUT2 #(
		.INIT('h4)
	) name125 (
		_w379_,
		_w382_,
		_w383_
	);
	LUT3 #(
		.INIT('hb0)
	) name126 (
		_w372_,
		_w378_,
		_w383_,
		_w384_
	);
	LUT4 #(
		.INIT('hfec8)
	) name127 (
		\a[18] ,
		\a[19] ,
		\b[18] ,
		\b[19] ,
		_w385_
	);
	LUT4 #(
		.INIT('h40f0)
	) name128 (
		_w372_,
		_w378_,
		_w381_,
		_w385_,
		_w386_
	);
	LUT2 #(
		.INIT('he)
	) name129 (
		_w384_,
		_w386_,
		_w387_
	);
	LUT2 #(
		.INIT('h1)
	) name130 (
		\a[21] ,
		\b[21] ,
		_w388_
	);
	LUT2 #(
		.INIT('h6)
	) name131 (
		\a[21] ,
		\b[21] ,
		_w389_
	);
	LUT4 #(
		.INIT('hfac8)
	) name132 (
		\a[19] ,
		\a[20] ,
		\b[19] ,
		\b[20] ,
		_w390_
	);
	LUT2 #(
		.INIT('h4)
	) name133 (
		_w379_,
		_w390_,
		_w391_
	);
	LUT3 #(
		.INIT('hb0)
	) name134 (
		_w372_,
		_w378_,
		_w391_,
		_w392_
	);
	LUT3 #(
		.INIT('h36)
	) name135 (
		_w380_,
		_w389_,
		_w392_,
		_w393_
	);
	LUT4 #(
		.INIT('h135f)
	) name136 (
		\a[20] ,
		\a[21] ,
		\b[20] ,
		\b[21] ,
		_w394_
	);
	LUT4 #(
		.INIT('h4f00)
	) name137 (
		_w372_,
		_w378_,
		_w391_,
		_w394_,
		_w395_
	);
	LUT2 #(
		.INIT('h1)
	) name138 (
		\a[22] ,
		\b[22] ,
		_w396_
	);
	LUT2 #(
		.INIT('h8)
	) name139 (
		\a[22] ,
		\b[22] ,
		_w397_
	);
	LUT2 #(
		.INIT('h6)
	) name140 (
		\a[22] ,
		\b[22] ,
		_w398_
	);
	LUT2 #(
		.INIT('h8)
	) name141 (
		_w394_,
		_w398_,
		_w399_
	);
	LUT4 #(
		.INIT('h4f00)
	) name142 (
		_w372_,
		_w378_,
		_w391_,
		_w399_,
		_w400_
	);
	LUT4 #(
		.INIT('hffa1)
	) name143 (
		_w388_,
		_w395_,
		_w398_,
		_w400_,
		_w401_
	);
	LUT2 #(
		.INIT('h2)
	) name144 (
		_w394_,
		_w397_,
		_w402_
	);
	LUT4 #(
		.INIT('h4f00)
	) name145 (
		_w372_,
		_w378_,
		_w391_,
		_w402_,
		_w403_
	);
	LUT4 #(
		.INIT('h0105)
	) name146 (
		\a[21] ,
		\a[22] ,
		\b[21] ,
		\b[22] ,
		_w404_
	);
	LUT2 #(
		.INIT('h8)
	) name147 (
		\a[23] ,
		\b[23] ,
		_w405_
	);
	LUT2 #(
		.INIT('h6)
	) name148 (
		\a[23] ,
		\b[23] ,
		_w406_
	);
	LUT4 #(
		.INIT('hfe01)
	) name149 (
		_w396_,
		_w403_,
		_w404_,
		_w406_,
		_w407_
	);
	LUT2 #(
		.INIT('h6)
	) name150 (
		\a[24] ,
		\b[24] ,
		_w408_
	);
	LUT4 #(
		.INIT('hfac8)
	) name151 (
		\a[22] ,
		\a[23] ,
		\b[22] ,
		\b[23] ,
		_w409_
	);
	LUT2 #(
		.INIT('h4)
	) name152 (
		_w404_,
		_w409_,
		_w410_
	);
	LUT4 #(
		.INIT('h2d3c)
	) name153 (
		_w403_,
		_w405_,
		_w408_,
		_w410_,
		_w411_
	);
	LUT4 #(
		.INIT('h135f)
	) name154 (
		\a[23] ,
		\a[24] ,
		\b[23] ,
		\b[24] ,
		_w412_
	);
	LUT2 #(
		.INIT('h8)
	) name155 (
		\a[25] ,
		\b[25] ,
		_w413_
	);
	LUT2 #(
		.INIT('h6)
	) name156 (
		\a[25] ,
		\b[25] ,
		_w414_
	);
	LUT4 #(
		.INIT('hc832)
	) name157 (
		\a[24] ,
		\a[25] ,
		\b[24] ,
		\b[25] ,
		_w415_
	);
	LUT4 #(
		.INIT('h4f00)
	) name158 (
		_w403_,
		_w410_,
		_w412_,
		_w415_,
		_w416_
	);
	LUT4 #(
		.INIT('h0104)
	) name159 (
		\a[24] ,
		\a[25] ,
		\b[24] ,
		\b[25] ,
		_w417_
	);
	LUT2 #(
		.INIT('h8)
	) name160 (
		_w412_,
		_w414_,
		_w418_
	);
	LUT4 #(
		.INIT('h040f)
	) name161 (
		_w403_,
		_w410_,
		_w417_,
		_w418_,
		_w419_
	);
	LUT2 #(
		.INIT('hb)
	) name162 (
		_w416_,
		_w419_,
		_w420_
	);
	LUT2 #(
		.INIT('h2)
	) name163 (
		_w412_,
		_w413_,
		_w421_
	);
	LUT4 #(
		.INIT('h0105)
	) name164 (
		\a[24] ,
		\a[25] ,
		\b[24] ,
		\b[25] ,
		_w422_
	);
	LUT2 #(
		.INIT('h8)
	) name165 (
		\a[26] ,
		\b[26] ,
		_w423_
	);
	LUT2 #(
		.INIT('h6)
	) name166 (
		\a[26] ,
		\b[26] ,
		_w424_
	);
	LUT4 #(
		.INIT('hc832)
	) name167 (
		\a[25] ,
		\a[26] ,
		\b[25] ,
		\b[26] ,
		_w425_
	);
	LUT2 #(
		.INIT('h4)
	) name168 (
		_w422_,
		_w425_,
		_w426_
	);
	LUT4 #(
		.INIT('h4f00)
	) name169 (
		_w403_,
		_w410_,
		_w421_,
		_w426_,
		_w427_
	);
	LUT4 #(
		.INIT('hfec8)
	) name170 (
		\a[24] ,
		\a[25] ,
		\b[24] ,
		\b[25] ,
		_w428_
	);
	LUT4 #(
		.INIT('h4f00)
	) name171 (
		_w403_,
		_w410_,
		_w421_,
		_w428_,
		_w429_
	);
	LUT3 #(
		.INIT('hce)
	) name172 (
		_w424_,
		_w427_,
		_w429_,
		_w430_
	);
	LUT2 #(
		.INIT('h1)
	) name173 (
		\a[27] ,
		\b[27] ,
		_w431_
	);
	LUT2 #(
		.INIT('h6)
	) name174 (
		\a[27] ,
		\b[27] ,
		_w432_
	);
	LUT4 #(
		.INIT('hfac8)
	) name175 (
		\a[25] ,
		\a[26] ,
		\b[25] ,
		\b[26] ,
		_w433_
	);
	LUT2 #(
		.INIT('h4)
	) name176 (
		_w422_,
		_w433_,
		_w434_
	);
	LUT4 #(
		.INIT('h4f00)
	) name177 (
		_w403_,
		_w410_,
		_w421_,
		_w434_,
		_w435_
	);
	LUT3 #(
		.INIT('h36)
	) name178 (
		_w423_,
		_w432_,
		_w435_,
		_w436_
	);
	LUT4 #(
		.INIT('h135f)
	) name179 (
		\a[26] ,
		\a[27] ,
		\b[26] ,
		\b[27] ,
		_w437_
	);
	LUT2 #(
		.INIT('h8)
	) name180 (
		\a[28] ,
		\b[28] ,
		_w438_
	);
	LUT2 #(
		.INIT('h6)
	) name181 (
		\a[28] ,
		\b[28] ,
		_w439_
	);
	LUT4 #(
		.INIT('hba45)
	) name182 (
		_w431_,
		_w435_,
		_w437_,
		_w439_,
		_w440_
	);
	LUT2 #(
		.INIT('h2)
	) name183 (
		_w437_,
		_w438_,
		_w441_
	);
	LUT4 #(
		.INIT('h0105)
	) name184 (
		\a[27] ,
		\a[28] ,
		\b[27] ,
		\b[28] ,
		_w442_
	);
	LUT2 #(
		.INIT('h8)
	) name185 (
		\a[29] ,
		\b[29] ,
		_w443_
	);
	LUT2 #(
		.INIT('h6)
	) name186 (
		\a[29] ,
		\b[29] ,
		_w444_
	);
	LUT4 #(
		.INIT('hc832)
	) name187 (
		\a[28] ,
		\a[29] ,
		\b[28] ,
		\b[29] ,
		_w445_
	);
	LUT2 #(
		.INIT('h4)
	) name188 (
		_w442_,
		_w445_,
		_w446_
	);
	LUT3 #(
		.INIT('hb0)
	) name189 (
		_w435_,
		_w441_,
		_w446_,
		_w447_
	);
	LUT4 #(
		.INIT('hfec8)
	) name190 (
		\a[27] ,
		\a[28] ,
		\b[27] ,
		\b[28] ,
		_w448_
	);
	LUT4 #(
		.INIT('h40f0)
	) name191 (
		_w435_,
		_w441_,
		_w444_,
		_w448_,
		_w449_
	);
	LUT2 #(
		.INIT('he)
	) name192 (
		_w447_,
		_w449_,
		_w450_
	);
	LUT2 #(
		.INIT('h1)
	) name193 (
		\a[30] ,
		\b[30] ,
		_w451_
	);
	LUT2 #(
		.INIT('h6)
	) name194 (
		\a[30] ,
		\b[30] ,
		_w452_
	);
	LUT4 #(
		.INIT('hfac8)
	) name195 (
		\a[28] ,
		\a[29] ,
		\b[28] ,
		\b[29] ,
		_w453_
	);
	LUT2 #(
		.INIT('h4)
	) name196 (
		_w442_,
		_w453_,
		_w454_
	);
	LUT3 #(
		.INIT('hb0)
	) name197 (
		_w435_,
		_w441_,
		_w454_,
		_w455_
	);
	LUT3 #(
		.INIT('h36)
	) name198 (
		_w443_,
		_w452_,
		_w455_,
		_w456_
	);
	LUT4 #(
		.INIT('h135f)
	) name199 (
		\a[29] ,
		\a[30] ,
		\b[29] ,
		\b[30] ,
		_w457_
	);
	LUT4 #(
		.INIT('h4f00)
	) name200 (
		_w435_,
		_w441_,
		_w454_,
		_w457_,
		_w458_
	);
	LUT2 #(
		.INIT('h1)
	) name201 (
		\a[31] ,
		\b[31] ,
		_w459_
	);
	LUT2 #(
		.INIT('h8)
	) name202 (
		\a[31] ,
		\b[31] ,
		_w460_
	);
	LUT2 #(
		.INIT('h6)
	) name203 (
		\a[31] ,
		\b[31] ,
		_w461_
	);
	LUT2 #(
		.INIT('h8)
	) name204 (
		_w457_,
		_w461_,
		_w462_
	);
	LUT4 #(
		.INIT('h4f00)
	) name205 (
		_w435_,
		_w441_,
		_w454_,
		_w462_,
		_w463_
	);
	LUT4 #(
		.INIT('hffa1)
	) name206 (
		_w451_,
		_w458_,
		_w461_,
		_w463_,
		_w464_
	);
	LUT2 #(
		.INIT('h2)
	) name207 (
		_w457_,
		_w460_,
		_w465_
	);
	LUT4 #(
		.INIT('h4f00)
	) name208 (
		_w435_,
		_w441_,
		_w454_,
		_w465_,
		_w466_
	);
	LUT4 #(
		.INIT('h0105)
	) name209 (
		\a[30] ,
		\a[31] ,
		\b[30] ,
		\b[31] ,
		_w467_
	);
	LUT2 #(
		.INIT('h8)
	) name210 (
		\a[32] ,
		\b[32] ,
		_w468_
	);
	LUT2 #(
		.INIT('h6)
	) name211 (
		\a[32] ,
		\b[32] ,
		_w469_
	);
	LUT4 #(
		.INIT('hfe01)
	) name212 (
		_w459_,
		_w466_,
		_w467_,
		_w469_,
		_w470_
	);
	LUT2 #(
		.INIT('h6)
	) name213 (
		\a[33] ,
		\b[33] ,
		_w471_
	);
	LUT4 #(
		.INIT('hfac8)
	) name214 (
		\a[31] ,
		\a[32] ,
		\b[31] ,
		\b[32] ,
		_w472_
	);
	LUT2 #(
		.INIT('h4)
	) name215 (
		_w467_,
		_w472_,
		_w473_
	);
	LUT4 #(
		.INIT('h2d3c)
	) name216 (
		_w466_,
		_w468_,
		_w471_,
		_w473_,
		_w474_
	);
	LUT4 #(
		.INIT('h135f)
	) name217 (
		\a[32] ,
		\a[33] ,
		\b[32] ,
		\b[33] ,
		_w475_
	);
	LUT2 #(
		.INIT('h8)
	) name218 (
		\a[34] ,
		\b[34] ,
		_w476_
	);
	LUT2 #(
		.INIT('h6)
	) name219 (
		\a[34] ,
		\b[34] ,
		_w477_
	);
	LUT4 #(
		.INIT('hc832)
	) name220 (
		\a[33] ,
		\a[34] ,
		\b[33] ,
		\b[34] ,
		_w478_
	);
	LUT4 #(
		.INIT('h4f00)
	) name221 (
		_w466_,
		_w473_,
		_w475_,
		_w478_,
		_w479_
	);
	LUT4 #(
		.INIT('h0104)
	) name222 (
		\a[33] ,
		\a[34] ,
		\b[33] ,
		\b[34] ,
		_w480_
	);
	LUT2 #(
		.INIT('h8)
	) name223 (
		_w475_,
		_w477_,
		_w481_
	);
	LUT4 #(
		.INIT('h040f)
	) name224 (
		_w466_,
		_w473_,
		_w480_,
		_w481_,
		_w482_
	);
	LUT2 #(
		.INIT('hb)
	) name225 (
		_w479_,
		_w482_,
		_w483_
	);
	LUT2 #(
		.INIT('h2)
	) name226 (
		_w475_,
		_w476_,
		_w484_
	);
	LUT4 #(
		.INIT('h0105)
	) name227 (
		\a[33] ,
		\a[34] ,
		\b[33] ,
		\b[34] ,
		_w485_
	);
	LUT2 #(
		.INIT('h8)
	) name228 (
		\a[35] ,
		\b[35] ,
		_w486_
	);
	LUT2 #(
		.INIT('h6)
	) name229 (
		\a[35] ,
		\b[35] ,
		_w487_
	);
	LUT4 #(
		.INIT('hc832)
	) name230 (
		\a[34] ,
		\a[35] ,
		\b[34] ,
		\b[35] ,
		_w488_
	);
	LUT2 #(
		.INIT('h4)
	) name231 (
		_w485_,
		_w488_,
		_w489_
	);
	LUT4 #(
		.INIT('h4f00)
	) name232 (
		_w466_,
		_w473_,
		_w484_,
		_w489_,
		_w490_
	);
	LUT4 #(
		.INIT('hfec8)
	) name233 (
		\a[33] ,
		\a[34] ,
		\b[33] ,
		\b[34] ,
		_w491_
	);
	LUT4 #(
		.INIT('h4f00)
	) name234 (
		_w466_,
		_w473_,
		_w484_,
		_w491_,
		_w492_
	);
	LUT3 #(
		.INIT('hce)
	) name235 (
		_w487_,
		_w490_,
		_w492_,
		_w493_
	);
	LUT2 #(
		.INIT('h1)
	) name236 (
		\a[36] ,
		\b[36] ,
		_w494_
	);
	LUT2 #(
		.INIT('h6)
	) name237 (
		\a[36] ,
		\b[36] ,
		_w495_
	);
	LUT4 #(
		.INIT('hfac8)
	) name238 (
		\a[34] ,
		\a[35] ,
		\b[34] ,
		\b[35] ,
		_w496_
	);
	LUT2 #(
		.INIT('h4)
	) name239 (
		_w485_,
		_w496_,
		_w497_
	);
	LUT4 #(
		.INIT('h4f00)
	) name240 (
		_w466_,
		_w473_,
		_w484_,
		_w497_,
		_w498_
	);
	LUT3 #(
		.INIT('h36)
	) name241 (
		_w486_,
		_w495_,
		_w498_,
		_w499_
	);
	LUT4 #(
		.INIT('h135f)
	) name242 (
		\a[35] ,
		\a[36] ,
		\b[35] ,
		\b[36] ,
		_w500_
	);
	LUT2 #(
		.INIT('h8)
	) name243 (
		\a[37] ,
		\b[37] ,
		_w501_
	);
	LUT2 #(
		.INIT('h6)
	) name244 (
		\a[37] ,
		\b[37] ,
		_w502_
	);
	LUT4 #(
		.INIT('hba45)
	) name245 (
		_w494_,
		_w498_,
		_w500_,
		_w502_,
		_w503_
	);
	LUT2 #(
		.INIT('h2)
	) name246 (
		_w500_,
		_w501_,
		_w504_
	);
	LUT4 #(
		.INIT('h0105)
	) name247 (
		\a[36] ,
		\a[37] ,
		\b[36] ,
		\b[37] ,
		_w505_
	);
	LUT2 #(
		.INIT('h8)
	) name248 (
		\a[38] ,
		\b[38] ,
		_w506_
	);
	LUT2 #(
		.INIT('h6)
	) name249 (
		\a[38] ,
		\b[38] ,
		_w507_
	);
	LUT4 #(
		.INIT('hc832)
	) name250 (
		\a[37] ,
		\a[38] ,
		\b[37] ,
		\b[38] ,
		_w508_
	);
	LUT2 #(
		.INIT('h4)
	) name251 (
		_w505_,
		_w508_,
		_w509_
	);
	LUT3 #(
		.INIT('hb0)
	) name252 (
		_w498_,
		_w504_,
		_w509_,
		_w510_
	);
	LUT4 #(
		.INIT('hfec8)
	) name253 (
		\a[36] ,
		\a[37] ,
		\b[36] ,
		\b[37] ,
		_w511_
	);
	LUT4 #(
		.INIT('h40f0)
	) name254 (
		_w498_,
		_w504_,
		_w507_,
		_w511_,
		_w512_
	);
	LUT2 #(
		.INIT('he)
	) name255 (
		_w510_,
		_w512_,
		_w513_
	);
	LUT2 #(
		.INIT('h1)
	) name256 (
		\a[39] ,
		\b[39] ,
		_w514_
	);
	LUT2 #(
		.INIT('h6)
	) name257 (
		\a[39] ,
		\b[39] ,
		_w515_
	);
	LUT4 #(
		.INIT('hfac8)
	) name258 (
		\a[37] ,
		\a[38] ,
		\b[37] ,
		\b[38] ,
		_w516_
	);
	LUT2 #(
		.INIT('h4)
	) name259 (
		_w505_,
		_w516_,
		_w517_
	);
	LUT3 #(
		.INIT('hb0)
	) name260 (
		_w498_,
		_w504_,
		_w517_,
		_w518_
	);
	LUT3 #(
		.INIT('h36)
	) name261 (
		_w506_,
		_w515_,
		_w518_,
		_w519_
	);
	LUT4 #(
		.INIT('h135f)
	) name262 (
		\a[38] ,
		\a[39] ,
		\b[38] ,
		\b[39] ,
		_w520_
	);
	LUT4 #(
		.INIT('h4f00)
	) name263 (
		_w498_,
		_w504_,
		_w517_,
		_w520_,
		_w521_
	);
	LUT2 #(
		.INIT('h1)
	) name264 (
		\a[40] ,
		\b[40] ,
		_w522_
	);
	LUT2 #(
		.INIT('h8)
	) name265 (
		\a[40] ,
		\b[40] ,
		_w523_
	);
	LUT2 #(
		.INIT('h6)
	) name266 (
		\a[40] ,
		\b[40] ,
		_w524_
	);
	LUT2 #(
		.INIT('h8)
	) name267 (
		_w520_,
		_w524_,
		_w525_
	);
	LUT4 #(
		.INIT('h4f00)
	) name268 (
		_w498_,
		_w504_,
		_w517_,
		_w525_,
		_w526_
	);
	LUT4 #(
		.INIT('hffa1)
	) name269 (
		_w514_,
		_w521_,
		_w524_,
		_w526_,
		_w527_
	);
	LUT2 #(
		.INIT('h2)
	) name270 (
		_w520_,
		_w523_,
		_w528_
	);
	LUT4 #(
		.INIT('h4f00)
	) name271 (
		_w498_,
		_w504_,
		_w517_,
		_w528_,
		_w529_
	);
	LUT4 #(
		.INIT('h0105)
	) name272 (
		\a[39] ,
		\a[40] ,
		\b[39] ,
		\b[40] ,
		_w530_
	);
	LUT2 #(
		.INIT('h8)
	) name273 (
		\a[41] ,
		\b[41] ,
		_w531_
	);
	LUT2 #(
		.INIT('h6)
	) name274 (
		\a[41] ,
		\b[41] ,
		_w532_
	);
	LUT4 #(
		.INIT('hfe01)
	) name275 (
		_w522_,
		_w529_,
		_w530_,
		_w532_,
		_w533_
	);
	LUT2 #(
		.INIT('h6)
	) name276 (
		\a[42] ,
		\b[42] ,
		_w534_
	);
	LUT4 #(
		.INIT('hfac8)
	) name277 (
		\a[40] ,
		\a[41] ,
		\b[40] ,
		\b[41] ,
		_w535_
	);
	LUT2 #(
		.INIT('h4)
	) name278 (
		_w530_,
		_w535_,
		_w536_
	);
	LUT4 #(
		.INIT('h2d3c)
	) name279 (
		_w529_,
		_w531_,
		_w534_,
		_w536_,
		_w537_
	);
	LUT4 #(
		.INIT('h135f)
	) name280 (
		\a[41] ,
		\a[42] ,
		\b[41] ,
		\b[42] ,
		_w538_
	);
	LUT2 #(
		.INIT('h8)
	) name281 (
		\a[43] ,
		\b[43] ,
		_w539_
	);
	LUT2 #(
		.INIT('h6)
	) name282 (
		\a[43] ,
		\b[43] ,
		_w540_
	);
	LUT4 #(
		.INIT('hc832)
	) name283 (
		\a[42] ,
		\a[43] ,
		\b[42] ,
		\b[43] ,
		_w541_
	);
	LUT4 #(
		.INIT('h4f00)
	) name284 (
		_w529_,
		_w536_,
		_w538_,
		_w541_,
		_w542_
	);
	LUT4 #(
		.INIT('h0104)
	) name285 (
		\a[42] ,
		\a[43] ,
		\b[42] ,
		\b[43] ,
		_w543_
	);
	LUT2 #(
		.INIT('h8)
	) name286 (
		_w538_,
		_w540_,
		_w544_
	);
	LUT4 #(
		.INIT('h040f)
	) name287 (
		_w529_,
		_w536_,
		_w543_,
		_w544_,
		_w545_
	);
	LUT2 #(
		.INIT('hb)
	) name288 (
		_w542_,
		_w545_,
		_w546_
	);
	LUT2 #(
		.INIT('h2)
	) name289 (
		_w538_,
		_w539_,
		_w547_
	);
	LUT4 #(
		.INIT('h0105)
	) name290 (
		\a[42] ,
		\a[43] ,
		\b[42] ,
		\b[43] ,
		_w548_
	);
	LUT2 #(
		.INIT('h8)
	) name291 (
		\a[44] ,
		\b[44] ,
		_w549_
	);
	LUT2 #(
		.INIT('h6)
	) name292 (
		\a[44] ,
		\b[44] ,
		_w550_
	);
	LUT4 #(
		.INIT('hc832)
	) name293 (
		\a[43] ,
		\a[44] ,
		\b[43] ,
		\b[44] ,
		_w551_
	);
	LUT2 #(
		.INIT('h4)
	) name294 (
		_w548_,
		_w551_,
		_w552_
	);
	LUT4 #(
		.INIT('h4f00)
	) name295 (
		_w529_,
		_w536_,
		_w547_,
		_w552_,
		_w553_
	);
	LUT4 #(
		.INIT('hfec8)
	) name296 (
		\a[42] ,
		\a[43] ,
		\b[42] ,
		\b[43] ,
		_w554_
	);
	LUT4 #(
		.INIT('h4f00)
	) name297 (
		_w529_,
		_w536_,
		_w547_,
		_w554_,
		_w555_
	);
	LUT3 #(
		.INIT('hce)
	) name298 (
		_w550_,
		_w553_,
		_w555_,
		_w556_
	);
	LUT2 #(
		.INIT('h1)
	) name299 (
		\a[45] ,
		\b[45] ,
		_w557_
	);
	LUT2 #(
		.INIT('h6)
	) name300 (
		\a[45] ,
		\b[45] ,
		_w558_
	);
	LUT4 #(
		.INIT('hfac8)
	) name301 (
		\a[43] ,
		\a[44] ,
		\b[43] ,
		\b[44] ,
		_w559_
	);
	LUT2 #(
		.INIT('h4)
	) name302 (
		_w548_,
		_w559_,
		_w560_
	);
	LUT4 #(
		.INIT('h4f00)
	) name303 (
		_w529_,
		_w536_,
		_w547_,
		_w560_,
		_w561_
	);
	LUT3 #(
		.INIT('h36)
	) name304 (
		_w549_,
		_w558_,
		_w561_,
		_w562_
	);
	LUT4 #(
		.INIT('h135f)
	) name305 (
		\a[44] ,
		\a[45] ,
		\b[44] ,
		\b[45] ,
		_w563_
	);
	LUT2 #(
		.INIT('h8)
	) name306 (
		\a[46] ,
		\b[46] ,
		_w564_
	);
	LUT2 #(
		.INIT('h6)
	) name307 (
		\a[46] ,
		\b[46] ,
		_w565_
	);
	LUT4 #(
		.INIT('hba45)
	) name308 (
		_w557_,
		_w561_,
		_w563_,
		_w565_,
		_w566_
	);
	LUT2 #(
		.INIT('h2)
	) name309 (
		_w563_,
		_w564_,
		_w567_
	);
	LUT4 #(
		.INIT('h0105)
	) name310 (
		\a[45] ,
		\a[46] ,
		\b[45] ,
		\b[46] ,
		_w568_
	);
	LUT2 #(
		.INIT('h8)
	) name311 (
		\a[47] ,
		\b[47] ,
		_w569_
	);
	LUT2 #(
		.INIT('h6)
	) name312 (
		\a[47] ,
		\b[47] ,
		_w570_
	);
	LUT4 #(
		.INIT('hc832)
	) name313 (
		\a[46] ,
		\a[47] ,
		\b[46] ,
		\b[47] ,
		_w571_
	);
	LUT2 #(
		.INIT('h4)
	) name314 (
		_w568_,
		_w571_,
		_w572_
	);
	LUT3 #(
		.INIT('hb0)
	) name315 (
		_w561_,
		_w567_,
		_w572_,
		_w573_
	);
	LUT4 #(
		.INIT('hfec8)
	) name316 (
		\a[45] ,
		\a[46] ,
		\b[45] ,
		\b[46] ,
		_w574_
	);
	LUT4 #(
		.INIT('h40f0)
	) name317 (
		_w561_,
		_w567_,
		_w570_,
		_w574_,
		_w575_
	);
	LUT2 #(
		.INIT('he)
	) name318 (
		_w573_,
		_w575_,
		_w576_
	);
	LUT2 #(
		.INIT('h1)
	) name319 (
		\a[48] ,
		\b[48] ,
		_w577_
	);
	LUT2 #(
		.INIT('h6)
	) name320 (
		\a[48] ,
		\b[48] ,
		_w578_
	);
	LUT4 #(
		.INIT('hfac8)
	) name321 (
		\a[46] ,
		\a[47] ,
		\b[46] ,
		\b[47] ,
		_w579_
	);
	LUT2 #(
		.INIT('h4)
	) name322 (
		_w568_,
		_w579_,
		_w580_
	);
	LUT3 #(
		.INIT('hb0)
	) name323 (
		_w561_,
		_w567_,
		_w580_,
		_w581_
	);
	LUT3 #(
		.INIT('h36)
	) name324 (
		_w569_,
		_w578_,
		_w581_,
		_w582_
	);
	LUT4 #(
		.INIT('h135f)
	) name325 (
		\a[47] ,
		\a[48] ,
		\b[47] ,
		\b[48] ,
		_w583_
	);
	LUT4 #(
		.INIT('h4f00)
	) name326 (
		_w561_,
		_w567_,
		_w580_,
		_w583_,
		_w584_
	);
	LUT2 #(
		.INIT('h1)
	) name327 (
		\a[49] ,
		\b[49] ,
		_w585_
	);
	LUT2 #(
		.INIT('h8)
	) name328 (
		\a[49] ,
		\b[49] ,
		_w586_
	);
	LUT2 #(
		.INIT('h6)
	) name329 (
		\a[49] ,
		\b[49] ,
		_w587_
	);
	LUT2 #(
		.INIT('h8)
	) name330 (
		_w583_,
		_w587_,
		_w588_
	);
	LUT4 #(
		.INIT('h4f00)
	) name331 (
		_w561_,
		_w567_,
		_w580_,
		_w588_,
		_w589_
	);
	LUT4 #(
		.INIT('hffa1)
	) name332 (
		_w577_,
		_w584_,
		_w587_,
		_w589_,
		_w590_
	);
	LUT2 #(
		.INIT('h2)
	) name333 (
		_w583_,
		_w586_,
		_w591_
	);
	LUT4 #(
		.INIT('h4f00)
	) name334 (
		_w561_,
		_w567_,
		_w580_,
		_w591_,
		_w592_
	);
	LUT4 #(
		.INIT('h0105)
	) name335 (
		\a[48] ,
		\a[49] ,
		\b[48] ,
		\b[49] ,
		_w593_
	);
	LUT2 #(
		.INIT('h8)
	) name336 (
		\a[50] ,
		\b[50] ,
		_w594_
	);
	LUT2 #(
		.INIT('h6)
	) name337 (
		\a[50] ,
		\b[50] ,
		_w595_
	);
	LUT4 #(
		.INIT('hfe01)
	) name338 (
		_w585_,
		_w592_,
		_w593_,
		_w595_,
		_w596_
	);
	LUT2 #(
		.INIT('h6)
	) name339 (
		\a[51] ,
		\b[51] ,
		_w597_
	);
	LUT4 #(
		.INIT('hfac8)
	) name340 (
		\a[49] ,
		\a[50] ,
		\b[49] ,
		\b[50] ,
		_w598_
	);
	LUT2 #(
		.INIT('h4)
	) name341 (
		_w593_,
		_w598_,
		_w599_
	);
	LUT4 #(
		.INIT('h2d3c)
	) name342 (
		_w592_,
		_w594_,
		_w597_,
		_w599_,
		_w600_
	);
	LUT4 #(
		.INIT('h135f)
	) name343 (
		\a[50] ,
		\a[51] ,
		\b[50] ,
		\b[51] ,
		_w601_
	);
	LUT2 #(
		.INIT('h8)
	) name344 (
		\a[52] ,
		\b[52] ,
		_w602_
	);
	LUT2 #(
		.INIT('h6)
	) name345 (
		\a[52] ,
		\b[52] ,
		_w603_
	);
	LUT4 #(
		.INIT('hc832)
	) name346 (
		\a[51] ,
		\a[52] ,
		\b[51] ,
		\b[52] ,
		_w604_
	);
	LUT4 #(
		.INIT('h4f00)
	) name347 (
		_w592_,
		_w599_,
		_w601_,
		_w604_,
		_w605_
	);
	LUT4 #(
		.INIT('h0104)
	) name348 (
		\a[51] ,
		\a[52] ,
		\b[51] ,
		\b[52] ,
		_w606_
	);
	LUT2 #(
		.INIT('h8)
	) name349 (
		_w601_,
		_w603_,
		_w607_
	);
	LUT4 #(
		.INIT('h040f)
	) name350 (
		_w592_,
		_w599_,
		_w606_,
		_w607_,
		_w608_
	);
	LUT2 #(
		.INIT('hb)
	) name351 (
		_w605_,
		_w608_,
		_w609_
	);
	LUT2 #(
		.INIT('h2)
	) name352 (
		_w601_,
		_w602_,
		_w610_
	);
	LUT4 #(
		.INIT('h0105)
	) name353 (
		\a[51] ,
		\a[52] ,
		\b[51] ,
		\b[52] ,
		_w611_
	);
	LUT2 #(
		.INIT('h8)
	) name354 (
		\a[53] ,
		\b[53] ,
		_w612_
	);
	LUT2 #(
		.INIT('h6)
	) name355 (
		\a[53] ,
		\b[53] ,
		_w613_
	);
	LUT4 #(
		.INIT('hc832)
	) name356 (
		\a[52] ,
		\a[53] ,
		\b[52] ,
		\b[53] ,
		_w614_
	);
	LUT2 #(
		.INIT('h4)
	) name357 (
		_w611_,
		_w614_,
		_w615_
	);
	LUT4 #(
		.INIT('h4f00)
	) name358 (
		_w592_,
		_w599_,
		_w610_,
		_w615_,
		_w616_
	);
	LUT4 #(
		.INIT('hfec8)
	) name359 (
		\a[51] ,
		\a[52] ,
		\b[51] ,
		\b[52] ,
		_w617_
	);
	LUT4 #(
		.INIT('h4f00)
	) name360 (
		_w592_,
		_w599_,
		_w610_,
		_w617_,
		_w618_
	);
	LUT3 #(
		.INIT('hce)
	) name361 (
		_w613_,
		_w616_,
		_w618_,
		_w619_
	);
	LUT2 #(
		.INIT('h1)
	) name362 (
		\a[54] ,
		\b[54] ,
		_w620_
	);
	LUT2 #(
		.INIT('h6)
	) name363 (
		\a[54] ,
		\b[54] ,
		_w621_
	);
	LUT4 #(
		.INIT('hfac8)
	) name364 (
		\a[52] ,
		\a[53] ,
		\b[52] ,
		\b[53] ,
		_w622_
	);
	LUT2 #(
		.INIT('h4)
	) name365 (
		_w611_,
		_w622_,
		_w623_
	);
	LUT4 #(
		.INIT('h4f00)
	) name366 (
		_w592_,
		_w599_,
		_w610_,
		_w623_,
		_w624_
	);
	LUT3 #(
		.INIT('h36)
	) name367 (
		_w612_,
		_w621_,
		_w624_,
		_w625_
	);
	LUT4 #(
		.INIT('h135f)
	) name368 (
		\a[53] ,
		\a[54] ,
		\b[53] ,
		\b[54] ,
		_w626_
	);
	LUT2 #(
		.INIT('h8)
	) name369 (
		\a[55] ,
		\b[55] ,
		_w627_
	);
	LUT2 #(
		.INIT('h6)
	) name370 (
		\a[55] ,
		\b[55] ,
		_w628_
	);
	LUT4 #(
		.INIT('hba45)
	) name371 (
		_w620_,
		_w624_,
		_w626_,
		_w628_,
		_w629_
	);
	LUT2 #(
		.INIT('h2)
	) name372 (
		_w626_,
		_w627_,
		_w630_
	);
	LUT4 #(
		.INIT('h0105)
	) name373 (
		\a[54] ,
		\a[55] ,
		\b[54] ,
		\b[55] ,
		_w631_
	);
	LUT2 #(
		.INIT('h8)
	) name374 (
		\a[56] ,
		\b[56] ,
		_w632_
	);
	LUT2 #(
		.INIT('h6)
	) name375 (
		\a[56] ,
		\b[56] ,
		_w633_
	);
	LUT4 #(
		.INIT('hc832)
	) name376 (
		\a[55] ,
		\a[56] ,
		\b[55] ,
		\b[56] ,
		_w634_
	);
	LUT2 #(
		.INIT('h4)
	) name377 (
		_w631_,
		_w634_,
		_w635_
	);
	LUT3 #(
		.INIT('hb0)
	) name378 (
		_w624_,
		_w630_,
		_w635_,
		_w636_
	);
	LUT4 #(
		.INIT('hfec8)
	) name379 (
		\a[54] ,
		\a[55] ,
		\b[54] ,
		\b[55] ,
		_w637_
	);
	LUT4 #(
		.INIT('h40f0)
	) name380 (
		_w624_,
		_w630_,
		_w633_,
		_w637_,
		_w638_
	);
	LUT2 #(
		.INIT('he)
	) name381 (
		_w636_,
		_w638_,
		_w639_
	);
	LUT2 #(
		.INIT('h1)
	) name382 (
		\a[57] ,
		\b[57] ,
		_w640_
	);
	LUT2 #(
		.INIT('h6)
	) name383 (
		\a[57] ,
		\b[57] ,
		_w641_
	);
	LUT4 #(
		.INIT('hfac8)
	) name384 (
		\a[55] ,
		\a[56] ,
		\b[55] ,
		\b[56] ,
		_w642_
	);
	LUT2 #(
		.INIT('h4)
	) name385 (
		_w631_,
		_w642_,
		_w643_
	);
	LUT3 #(
		.INIT('hb0)
	) name386 (
		_w624_,
		_w630_,
		_w643_,
		_w644_
	);
	LUT3 #(
		.INIT('h36)
	) name387 (
		_w632_,
		_w641_,
		_w644_,
		_w645_
	);
	LUT4 #(
		.INIT('h135f)
	) name388 (
		\a[56] ,
		\a[57] ,
		\b[56] ,
		\b[57] ,
		_w646_
	);
	LUT4 #(
		.INIT('h4f00)
	) name389 (
		_w624_,
		_w630_,
		_w643_,
		_w646_,
		_w647_
	);
	LUT2 #(
		.INIT('h1)
	) name390 (
		\a[58] ,
		\b[58] ,
		_w648_
	);
	LUT2 #(
		.INIT('h8)
	) name391 (
		\a[58] ,
		\b[58] ,
		_w649_
	);
	LUT2 #(
		.INIT('h6)
	) name392 (
		\a[58] ,
		\b[58] ,
		_w650_
	);
	LUT2 #(
		.INIT('h8)
	) name393 (
		_w646_,
		_w650_,
		_w651_
	);
	LUT4 #(
		.INIT('h4f00)
	) name394 (
		_w624_,
		_w630_,
		_w643_,
		_w651_,
		_w652_
	);
	LUT4 #(
		.INIT('hffa1)
	) name395 (
		_w640_,
		_w647_,
		_w650_,
		_w652_,
		_w653_
	);
	LUT2 #(
		.INIT('h2)
	) name396 (
		_w646_,
		_w649_,
		_w654_
	);
	LUT4 #(
		.INIT('h4f00)
	) name397 (
		_w624_,
		_w630_,
		_w643_,
		_w654_,
		_w655_
	);
	LUT4 #(
		.INIT('h0105)
	) name398 (
		\a[57] ,
		\a[58] ,
		\b[57] ,
		\b[58] ,
		_w656_
	);
	LUT2 #(
		.INIT('h8)
	) name399 (
		\a[59] ,
		\b[59] ,
		_w657_
	);
	LUT2 #(
		.INIT('h6)
	) name400 (
		\a[59] ,
		\b[59] ,
		_w658_
	);
	LUT4 #(
		.INIT('hfe01)
	) name401 (
		_w648_,
		_w655_,
		_w656_,
		_w658_,
		_w659_
	);
	LUT2 #(
		.INIT('h6)
	) name402 (
		\a[60] ,
		\b[60] ,
		_w660_
	);
	LUT4 #(
		.INIT('hfac8)
	) name403 (
		\a[58] ,
		\a[59] ,
		\b[58] ,
		\b[59] ,
		_w661_
	);
	LUT2 #(
		.INIT('h4)
	) name404 (
		_w656_,
		_w661_,
		_w662_
	);
	LUT4 #(
		.INIT('h2d3c)
	) name405 (
		_w655_,
		_w657_,
		_w660_,
		_w662_,
		_w663_
	);
	LUT4 #(
		.INIT('h135f)
	) name406 (
		\a[59] ,
		\a[60] ,
		\b[59] ,
		\b[60] ,
		_w664_
	);
	LUT2 #(
		.INIT('h8)
	) name407 (
		\a[61] ,
		\b[61] ,
		_w665_
	);
	LUT2 #(
		.INIT('h6)
	) name408 (
		\a[61] ,
		\b[61] ,
		_w666_
	);
	LUT4 #(
		.INIT('hc832)
	) name409 (
		\a[60] ,
		\a[61] ,
		\b[60] ,
		\b[61] ,
		_w667_
	);
	LUT4 #(
		.INIT('h4f00)
	) name410 (
		_w655_,
		_w662_,
		_w664_,
		_w667_,
		_w668_
	);
	LUT4 #(
		.INIT('h0104)
	) name411 (
		\a[60] ,
		\a[61] ,
		\b[60] ,
		\b[61] ,
		_w669_
	);
	LUT2 #(
		.INIT('h8)
	) name412 (
		_w664_,
		_w666_,
		_w670_
	);
	LUT4 #(
		.INIT('h040f)
	) name413 (
		_w655_,
		_w662_,
		_w669_,
		_w670_,
		_w671_
	);
	LUT2 #(
		.INIT('hb)
	) name414 (
		_w668_,
		_w671_,
		_w672_
	);
	LUT2 #(
		.INIT('h2)
	) name415 (
		_w664_,
		_w665_,
		_w673_
	);
	LUT4 #(
		.INIT('h0105)
	) name416 (
		\a[60] ,
		\a[61] ,
		\b[60] ,
		\b[61] ,
		_w674_
	);
	LUT2 #(
		.INIT('h8)
	) name417 (
		\a[62] ,
		\b[62] ,
		_w675_
	);
	LUT2 #(
		.INIT('h6)
	) name418 (
		\a[62] ,
		\b[62] ,
		_w676_
	);
	LUT4 #(
		.INIT('hc832)
	) name419 (
		\a[61] ,
		\a[62] ,
		\b[61] ,
		\b[62] ,
		_w677_
	);
	LUT2 #(
		.INIT('h4)
	) name420 (
		_w674_,
		_w677_,
		_w678_
	);
	LUT4 #(
		.INIT('h4f00)
	) name421 (
		_w655_,
		_w662_,
		_w673_,
		_w678_,
		_w679_
	);
	LUT4 #(
		.INIT('hfec8)
	) name422 (
		\a[60] ,
		\a[61] ,
		\b[60] ,
		\b[61] ,
		_w680_
	);
	LUT4 #(
		.INIT('h4f00)
	) name423 (
		_w655_,
		_w662_,
		_w673_,
		_w680_,
		_w681_
	);
	LUT3 #(
		.INIT('hce)
	) name424 (
		_w676_,
		_w679_,
		_w681_,
		_w682_
	);
	LUT2 #(
		.INIT('h1)
	) name425 (
		\a[63] ,
		\b[63] ,
		_w683_
	);
	LUT2 #(
		.INIT('h6)
	) name426 (
		\a[63] ,
		\b[63] ,
		_w684_
	);
	LUT4 #(
		.INIT('hfac8)
	) name427 (
		\a[61] ,
		\a[62] ,
		\b[61] ,
		\b[62] ,
		_w685_
	);
	LUT2 #(
		.INIT('h4)
	) name428 (
		_w674_,
		_w685_,
		_w686_
	);
	LUT4 #(
		.INIT('h4f00)
	) name429 (
		_w655_,
		_w662_,
		_w673_,
		_w686_,
		_w687_
	);
	LUT3 #(
		.INIT('h36)
	) name430 (
		_w675_,
		_w684_,
		_w687_,
		_w688_
	);
	LUT4 #(
		.INIT('h135f)
	) name431 (
		\a[62] ,
		\a[63] ,
		\b[62] ,
		\b[63] ,
		_w689_
	);
	LUT2 #(
		.INIT('h8)
	) name432 (
		\a[64] ,
		\b[64] ,
		_w690_
	);
	LUT2 #(
		.INIT('h6)
	) name433 (
		\a[64] ,
		\b[64] ,
		_w691_
	);
	LUT4 #(
		.INIT('hba45)
	) name434 (
		_w683_,
		_w687_,
		_w689_,
		_w691_,
		_w692_
	);
	LUT2 #(
		.INIT('h2)
	) name435 (
		_w689_,
		_w690_,
		_w693_
	);
	LUT4 #(
		.INIT('h0105)
	) name436 (
		\a[63] ,
		\a[64] ,
		\b[63] ,
		\b[64] ,
		_w694_
	);
	LUT2 #(
		.INIT('h8)
	) name437 (
		\a[65] ,
		\b[65] ,
		_w695_
	);
	LUT2 #(
		.INIT('h6)
	) name438 (
		\a[65] ,
		\b[65] ,
		_w696_
	);
	LUT4 #(
		.INIT('hc832)
	) name439 (
		\a[64] ,
		\a[65] ,
		\b[64] ,
		\b[65] ,
		_w697_
	);
	LUT2 #(
		.INIT('h4)
	) name440 (
		_w694_,
		_w697_,
		_w698_
	);
	LUT3 #(
		.INIT('hb0)
	) name441 (
		_w687_,
		_w693_,
		_w698_,
		_w699_
	);
	LUT4 #(
		.INIT('hfec8)
	) name442 (
		\a[63] ,
		\a[64] ,
		\b[63] ,
		\b[64] ,
		_w700_
	);
	LUT4 #(
		.INIT('h40f0)
	) name443 (
		_w687_,
		_w693_,
		_w696_,
		_w700_,
		_w701_
	);
	LUT2 #(
		.INIT('he)
	) name444 (
		_w699_,
		_w701_,
		_w702_
	);
	LUT2 #(
		.INIT('h1)
	) name445 (
		\a[66] ,
		\b[66] ,
		_w703_
	);
	LUT2 #(
		.INIT('h6)
	) name446 (
		\a[66] ,
		\b[66] ,
		_w704_
	);
	LUT4 #(
		.INIT('hfac8)
	) name447 (
		\a[64] ,
		\a[65] ,
		\b[64] ,
		\b[65] ,
		_w705_
	);
	LUT2 #(
		.INIT('h4)
	) name448 (
		_w694_,
		_w705_,
		_w706_
	);
	LUT3 #(
		.INIT('hb0)
	) name449 (
		_w687_,
		_w693_,
		_w706_,
		_w707_
	);
	LUT3 #(
		.INIT('h36)
	) name450 (
		_w695_,
		_w704_,
		_w707_,
		_w708_
	);
	LUT4 #(
		.INIT('h135f)
	) name451 (
		\a[65] ,
		\a[66] ,
		\b[65] ,
		\b[66] ,
		_w709_
	);
	LUT4 #(
		.INIT('h4f00)
	) name452 (
		_w687_,
		_w693_,
		_w706_,
		_w709_,
		_w710_
	);
	LUT2 #(
		.INIT('h1)
	) name453 (
		\a[67] ,
		\b[67] ,
		_w711_
	);
	LUT2 #(
		.INIT('h8)
	) name454 (
		\a[67] ,
		\b[67] ,
		_w712_
	);
	LUT2 #(
		.INIT('h6)
	) name455 (
		\a[67] ,
		\b[67] ,
		_w713_
	);
	LUT2 #(
		.INIT('h8)
	) name456 (
		_w709_,
		_w713_,
		_w714_
	);
	LUT4 #(
		.INIT('h4f00)
	) name457 (
		_w687_,
		_w693_,
		_w706_,
		_w714_,
		_w715_
	);
	LUT4 #(
		.INIT('hffa1)
	) name458 (
		_w703_,
		_w710_,
		_w713_,
		_w715_,
		_w716_
	);
	LUT2 #(
		.INIT('h2)
	) name459 (
		_w709_,
		_w712_,
		_w717_
	);
	LUT4 #(
		.INIT('h4f00)
	) name460 (
		_w687_,
		_w693_,
		_w706_,
		_w717_,
		_w718_
	);
	LUT4 #(
		.INIT('h0105)
	) name461 (
		\a[66] ,
		\a[67] ,
		\b[66] ,
		\b[67] ,
		_w719_
	);
	LUT2 #(
		.INIT('h8)
	) name462 (
		\a[68] ,
		\b[68] ,
		_w720_
	);
	LUT2 #(
		.INIT('h6)
	) name463 (
		\a[68] ,
		\b[68] ,
		_w721_
	);
	LUT4 #(
		.INIT('hfe01)
	) name464 (
		_w711_,
		_w718_,
		_w719_,
		_w721_,
		_w722_
	);
	LUT2 #(
		.INIT('h6)
	) name465 (
		\a[69] ,
		\b[69] ,
		_w723_
	);
	LUT4 #(
		.INIT('hfac8)
	) name466 (
		\a[67] ,
		\a[68] ,
		\b[67] ,
		\b[68] ,
		_w724_
	);
	LUT2 #(
		.INIT('h4)
	) name467 (
		_w719_,
		_w724_,
		_w725_
	);
	LUT4 #(
		.INIT('h2d3c)
	) name468 (
		_w718_,
		_w720_,
		_w723_,
		_w725_,
		_w726_
	);
	LUT4 #(
		.INIT('h135f)
	) name469 (
		\a[68] ,
		\a[69] ,
		\b[68] ,
		\b[69] ,
		_w727_
	);
	LUT2 #(
		.INIT('h8)
	) name470 (
		\a[70] ,
		\b[70] ,
		_w728_
	);
	LUT2 #(
		.INIT('h6)
	) name471 (
		\a[70] ,
		\b[70] ,
		_w729_
	);
	LUT4 #(
		.INIT('hc832)
	) name472 (
		\a[69] ,
		\a[70] ,
		\b[69] ,
		\b[70] ,
		_w730_
	);
	LUT4 #(
		.INIT('h4f00)
	) name473 (
		_w718_,
		_w725_,
		_w727_,
		_w730_,
		_w731_
	);
	LUT4 #(
		.INIT('h0104)
	) name474 (
		\a[69] ,
		\a[70] ,
		\b[69] ,
		\b[70] ,
		_w732_
	);
	LUT2 #(
		.INIT('h8)
	) name475 (
		_w727_,
		_w729_,
		_w733_
	);
	LUT4 #(
		.INIT('h040f)
	) name476 (
		_w718_,
		_w725_,
		_w732_,
		_w733_,
		_w734_
	);
	LUT2 #(
		.INIT('hb)
	) name477 (
		_w731_,
		_w734_,
		_w735_
	);
	LUT2 #(
		.INIT('h2)
	) name478 (
		_w727_,
		_w728_,
		_w736_
	);
	LUT4 #(
		.INIT('h0105)
	) name479 (
		\a[69] ,
		\a[70] ,
		\b[69] ,
		\b[70] ,
		_w737_
	);
	LUT2 #(
		.INIT('h8)
	) name480 (
		\a[71] ,
		\b[71] ,
		_w738_
	);
	LUT2 #(
		.INIT('h6)
	) name481 (
		\a[71] ,
		\b[71] ,
		_w739_
	);
	LUT4 #(
		.INIT('hc832)
	) name482 (
		\a[70] ,
		\a[71] ,
		\b[70] ,
		\b[71] ,
		_w740_
	);
	LUT2 #(
		.INIT('h4)
	) name483 (
		_w737_,
		_w740_,
		_w741_
	);
	LUT4 #(
		.INIT('h4f00)
	) name484 (
		_w718_,
		_w725_,
		_w736_,
		_w741_,
		_w742_
	);
	LUT4 #(
		.INIT('hfec8)
	) name485 (
		\a[69] ,
		\a[70] ,
		\b[69] ,
		\b[70] ,
		_w743_
	);
	LUT4 #(
		.INIT('h4f00)
	) name486 (
		_w718_,
		_w725_,
		_w736_,
		_w743_,
		_w744_
	);
	LUT3 #(
		.INIT('hce)
	) name487 (
		_w739_,
		_w742_,
		_w744_,
		_w745_
	);
	LUT2 #(
		.INIT('h1)
	) name488 (
		\a[72] ,
		\b[72] ,
		_w746_
	);
	LUT2 #(
		.INIT('h6)
	) name489 (
		\a[72] ,
		\b[72] ,
		_w747_
	);
	LUT4 #(
		.INIT('hfac8)
	) name490 (
		\a[70] ,
		\a[71] ,
		\b[70] ,
		\b[71] ,
		_w748_
	);
	LUT2 #(
		.INIT('h4)
	) name491 (
		_w737_,
		_w748_,
		_w749_
	);
	LUT4 #(
		.INIT('h4f00)
	) name492 (
		_w718_,
		_w725_,
		_w736_,
		_w749_,
		_w750_
	);
	LUT3 #(
		.INIT('h36)
	) name493 (
		_w738_,
		_w747_,
		_w750_,
		_w751_
	);
	LUT4 #(
		.INIT('h135f)
	) name494 (
		\a[71] ,
		\a[72] ,
		\b[71] ,
		\b[72] ,
		_w752_
	);
	LUT2 #(
		.INIT('h8)
	) name495 (
		\a[73] ,
		\b[73] ,
		_w753_
	);
	LUT2 #(
		.INIT('h6)
	) name496 (
		\a[73] ,
		\b[73] ,
		_w754_
	);
	LUT4 #(
		.INIT('hba45)
	) name497 (
		_w746_,
		_w750_,
		_w752_,
		_w754_,
		_w755_
	);
	LUT2 #(
		.INIT('h2)
	) name498 (
		_w752_,
		_w753_,
		_w756_
	);
	LUT4 #(
		.INIT('h0105)
	) name499 (
		\a[72] ,
		\a[73] ,
		\b[72] ,
		\b[73] ,
		_w757_
	);
	LUT2 #(
		.INIT('h8)
	) name500 (
		\a[74] ,
		\b[74] ,
		_w758_
	);
	LUT2 #(
		.INIT('h6)
	) name501 (
		\a[74] ,
		\b[74] ,
		_w759_
	);
	LUT4 #(
		.INIT('hc832)
	) name502 (
		\a[73] ,
		\a[74] ,
		\b[73] ,
		\b[74] ,
		_w760_
	);
	LUT2 #(
		.INIT('h4)
	) name503 (
		_w757_,
		_w760_,
		_w761_
	);
	LUT3 #(
		.INIT('hb0)
	) name504 (
		_w750_,
		_w756_,
		_w761_,
		_w762_
	);
	LUT4 #(
		.INIT('hfec8)
	) name505 (
		\a[72] ,
		\a[73] ,
		\b[72] ,
		\b[73] ,
		_w763_
	);
	LUT4 #(
		.INIT('h40f0)
	) name506 (
		_w750_,
		_w756_,
		_w759_,
		_w763_,
		_w764_
	);
	LUT2 #(
		.INIT('he)
	) name507 (
		_w762_,
		_w764_,
		_w765_
	);
	LUT2 #(
		.INIT('h1)
	) name508 (
		\a[75] ,
		\b[75] ,
		_w766_
	);
	LUT2 #(
		.INIT('h6)
	) name509 (
		\a[75] ,
		\b[75] ,
		_w767_
	);
	LUT4 #(
		.INIT('hfac8)
	) name510 (
		\a[73] ,
		\a[74] ,
		\b[73] ,
		\b[74] ,
		_w768_
	);
	LUT2 #(
		.INIT('h4)
	) name511 (
		_w757_,
		_w768_,
		_w769_
	);
	LUT3 #(
		.INIT('hb0)
	) name512 (
		_w750_,
		_w756_,
		_w769_,
		_w770_
	);
	LUT3 #(
		.INIT('h36)
	) name513 (
		_w758_,
		_w767_,
		_w770_,
		_w771_
	);
	LUT4 #(
		.INIT('h135f)
	) name514 (
		\a[74] ,
		\a[75] ,
		\b[74] ,
		\b[75] ,
		_w772_
	);
	LUT4 #(
		.INIT('h4f00)
	) name515 (
		_w750_,
		_w756_,
		_w769_,
		_w772_,
		_w773_
	);
	LUT2 #(
		.INIT('h1)
	) name516 (
		\a[76] ,
		\b[76] ,
		_w774_
	);
	LUT2 #(
		.INIT('h8)
	) name517 (
		\a[76] ,
		\b[76] ,
		_w775_
	);
	LUT2 #(
		.INIT('h6)
	) name518 (
		\a[76] ,
		\b[76] ,
		_w776_
	);
	LUT2 #(
		.INIT('h8)
	) name519 (
		_w772_,
		_w776_,
		_w777_
	);
	LUT4 #(
		.INIT('h4f00)
	) name520 (
		_w750_,
		_w756_,
		_w769_,
		_w777_,
		_w778_
	);
	LUT4 #(
		.INIT('hffa1)
	) name521 (
		_w766_,
		_w773_,
		_w776_,
		_w778_,
		_w779_
	);
	LUT2 #(
		.INIT('h2)
	) name522 (
		_w772_,
		_w775_,
		_w780_
	);
	LUT4 #(
		.INIT('h4f00)
	) name523 (
		_w750_,
		_w756_,
		_w769_,
		_w780_,
		_w781_
	);
	LUT4 #(
		.INIT('h0105)
	) name524 (
		\a[75] ,
		\a[76] ,
		\b[75] ,
		\b[76] ,
		_w782_
	);
	LUT2 #(
		.INIT('h8)
	) name525 (
		\a[77] ,
		\b[77] ,
		_w783_
	);
	LUT2 #(
		.INIT('h6)
	) name526 (
		\a[77] ,
		\b[77] ,
		_w784_
	);
	LUT4 #(
		.INIT('hfe01)
	) name527 (
		_w774_,
		_w781_,
		_w782_,
		_w784_,
		_w785_
	);
	LUT2 #(
		.INIT('h6)
	) name528 (
		\a[78] ,
		\b[78] ,
		_w786_
	);
	LUT4 #(
		.INIT('hfac8)
	) name529 (
		\a[76] ,
		\a[77] ,
		\b[76] ,
		\b[77] ,
		_w787_
	);
	LUT2 #(
		.INIT('h4)
	) name530 (
		_w782_,
		_w787_,
		_w788_
	);
	LUT4 #(
		.INIT('h2d3c)
	) name531 (
		_w781_,
		_w783_,
		_w786_,
		_w788_,
		_w789_
	);
	LUT4 #(
		.INIT('h135f)
	) name532 (
		\a[77] ,
		\a[78] ,
		\b[77] ,
		\b[78] ,
		_w790_
	);
	LUT2 #(
		.INIT('h8)
	) name533 (
		\a[79] ,
		\b[79] ,
		_w791_
	);
	LUT2 #(
		.INIT('h6)
	) name534 (
		\a[79] ,
		\b[79] ,
		_w792_
	);
	LUT4 #(
		.INIT('hc832)
	) name535 (
		\a[78] ,
		\a[79] ,
		\b[78] ,
		\b[79] ,
		_w793_
	);
	LUT4 #(
		.INIT('h4f00)
	) name536 (
		_w781_,
		_w788_,
		_w790_,
		_w793_,
		_w794_
	);
	LUT4 #(
		.INIT('h0104)
	) name537 (
		\a[78] ,
		\a[79] ,
		\b[78] ,
		\b[79] ,
		_w795_
	);
	LUT2 #(
		.INIT('h8)
	) name538 (
		_w790_,
		_w792_,
		_w796_
	);
	LUT4 #(
		.INIT('h040f)
	) name539 (
		_w781_,
		_w788_,
		_w795_,
		_w796_,
		_w797_
	);
	LUT2 #(
		.INIT('hb)
	) name540 (
		_w794_,
		_w797_,
		_w798_
	);
	LUT2 #(
		.INIT('h2)
	) name541 (
		_w790_,
		_w791_,
		_w799_
	);
	LUT4 #(
		.INIT('h0105)
	) name542 (
		\a[78] ,
		\a[79] ,
		\b[78] ,
		\b[79] ,
		_w800_
	);
	LUT2 #(
		.INIT('h8)
	) name543 (
		\a[80] ,
		\b[80] ,
		_w801_
	);
	LUT2 #(
		.INIT('h6)
	) name544 (
		\a[80] ,
		\b[80] ,
		_w802_
	);
	LUT4 #(
		.INIT('hc832)
	) name545 (
		\a[79] ,
		\a[80] ,
		\b[79] ,
		\b[80] ,
		_w803_
	);
	LUT2 #(
		.INIT('h4)
	) name546 (
		_w800_,
		_w803_,
		_w804_
	);
	LUT4 #(
		.INIT('h4f00)
	) name547 (
		_w781_,
		_w788_,
		_w799_,
		_w804_,
		_w805_
	);
	LUT4 #(
		.INIT('hfec8)
	) name548 (
		\a[78] ,
		\a[79] ,
		\b[78] ,
		\b[79] ,
		_w806_
	);
	LUT4 #(
		.INIT('h4f00)
	) name549 (
		_w781_,
		_w788_,
		_w799_,
		_w806_,
		_w807_
	);
	LUT3 #(
		.INIT('hce)
	) name550 (
		_w802_,
		_w805_,
		_w807_,
		_w808_
	);
	LUT2 #(
		.INIT('h1)
	) name551 (
		\a[81] ,
		\b[81] ,
		_w809_
	);
	LUT2 #(
		.INIT('h6)
	) name552 (
		\a[81] ,
		\b[81] ,
		_w810_
	);
	LUT4 #(
		.INIT('hfac8)
	) name553 (
		\a[79] ,
		\a[80] ,
		\b[79] ,
		\b[80] ,
		_w811_
	);
	LUT2 #(
		.INIT('h4)
	) name554 (
		_w800_,
		_w811_,
		_w812_
	);
	LUT4 #(
		.INIT('h4f00)
	) name555 (
		_w781_,
		_w788_,
		_w799_,
		_w812_,
		_w813_
	);
	LUT3 #(
		.INIT('h36)
	) name556 (
		_w801_,
		_w810_,
		_w813_,
		_w814_
	);
	LUT4 #(
		.INIT('h135f)
	) name557 (
		\a[80] ,
		\a[81] ,
		\b[80] ,
		\b[81] ,
		_w815_
	);
	LUT2 #(
		.INIT('h8)
	) name558 (
		\a[82] ,
		\b[82] ,
		_w816_
	);
	LUT2 #(
		.INIT('h6)
	) name559 (
		\a[82] ,
		\b[82] ,
		_w817_
	);
	LUT4 #(
		.INIT('hba45)
	) name560 (
		_w809_,
		_w813_,
		_w815_,
		_w817_,
		_w818_
	);
	LUT2 #(
		.INIT('h2)
	) name561 (
		_w815_,
		_w816_,
		_w819_
	);
	LUT4 #(
		.INIT('h0105)
	) name562 (
		\a[81] ,
		\a[82] ,
		\b[81] ,
		\b[82] ,
		_w820_
	);
	LUT2 #(
		.INIT('h8)
	) name563 (
		\a[83] ,
		\b[83] ,
		_w821_
	);
	LUT2 #(
		.INIT('h6)
	) name564 (
		\a[83] ,
		\b[83] ,
		_w822_
	);
	LUT4 #(
		.INIT('hc832)
	) name565 (
		\a[82] ,
		\a[83] ,
		\b[82] ,
		\b[83] ,
		_w823_
	);
	LUT2 #(
		.INIT('h4)
	) name566 (
		_w820_,
		_w823_,
		_w824_
	);
	LUT3 #(
		.INIT('hb0)
	) name567 (
		_w813_,
		_w819_,
		_w824_,
		_w825_
	);
	LUT4 #(
		.INIT('hfec8)
	) name568 (
		\a[81] ,
		\a[82] ,
		\b[81] ,
		\b[82] ,
		_w826_
	);
	LUT4 #(
		.INIT('h40f0)
	) name569 (
		_w813_,
		_w819_,
		_w822_,
		_w826_,
		_w827_
	);
	LUT2 #(
		.INIT('he)
	) name570 (
		_w825_,
		_w827_,
		_w828_
	);
	LUT2 #(
		.INIT('h1)
	) name571 (
		\a[84] ,
		\b[84] ,
		_w829_
	);
	LUT2 #(
		.INIT('h6)
	) name572 (
		\a[84] ,
		\b[84] ,
		_w830_
	);
	LUT4 #(
		.INIT('hfac8)
	) name573 (
		\a[82] ,
		\a[83] ,
		\b[82] ,
		\b[83] ,
		_w831_
	);
	LUT2 #(
		.INIT('h4)
	) name574 (
		_w820_,
		_w831_,
		_w832_
	);
	LUT3 #(
		.INIT('hb0)
	) name575 (
		_w813_,
		_w819_,
		_w832_,
		_w833_
	);
	LUT3 #(
		.INIT('h36)
	) name576 (
		_w821_,
		_w830_,
		_w833_,
		_w834_
	);
	LUT4 #(
		.INIT('h135f)
	) name577 (
		\a[83] ,
		\a[84] ,
		\b[83] ,
		\b[84] ,
		_w835_
	);
	LUT4 #(
		.INIT('h4f00)
	) name578 (
		_w813_,
		_w819_,
		_w832_,
		_w835_,
		_w836_
	);
	LUT2 #(
		.INIT('h1)
	) name579 (
		\a[85] ,
		\b[85] ,
		_w837_
	);
	LUT2 #(
		.INIT('h8)
	) name580 (
		\a[85] ,
		\b[85] ,
		_w838_
	);
	LUT2 #(
		.INIT('h6)
	) name581 (
		\a[85] ,
		\b[85] ,
		_w839_
	);
	LUT2 #(
		.INIT('h8)
	) name582 (
		_w835_,
		_w839_,
		_w840_
	);
	LUT4 #(
		.INIT('h4f00)
	) name583 (
		_w813_,
		_w819_,
		_w832_,
		_w840_,
		_w841_
	);
	LUT4 #(
		.INIT('hffa1)
	) name584 (
		_w829_,
		_w836_,
		_w839_,
		_w841_,
		_w842_
	);
	LUT2 #(
		.INIT('h2)
	) name585 (
		_w835_,
		_w838_,
		_w843_
	);
	LUT4 #(
		.INIT('h4f00)
	) name586 (
		_w813_,
		_w819_,
		_w832_,
		_w843_,
		_w844_
	);
	LUT4 #(
		.INIT('h0105)
	) name587 (
		\a[84] ,
		\a[85] ,
		\b[84] ,
		\b[85] ,
		_w845_
	);
	LUT2 #(
		.INIT('h8)
	) name588 (
		\a[86] ,
		\b[86] ,
		_w846_
	);
	LUT2 #(
		.INIT('h6)
	) name589 (
		\a[86] ,
		\b[86] ,
		_w847_
	);
	LUT4 #(
		.INIT('hfe01)
	) name590 (
		_w837_,
		_w844_,
		_w845_,
		_w847_,
		_w848_
	);
	LUT2 #(
		.INIT('h6)
	) name591 (
		\a[87] ,
		\b[87] ,
		_w849_
	);
	LUT4 #(
		.INIT('hfac8)
	) name592 (
		\a[85] ,
		\a[86] ,
		\b[85] ,
		\b[86] ,
		_w850_
	);
	LUT2 #(
		.INIT('h4)
	) name593 (
		_w845_,
		_w850_,
		_w851_
	);
	LUT4 #(
		.INIT('h2d3c)
	) name594 (
		_w844_,
		_w846_,
		_w849_,
		_w851_,
		_w852_
	);
	LUT4 #(
		.INIT('h135f)
	) name595 (
		\a[86] ,
		\a[87] ,
		\b[86] ,
		\b[87] ,
		_w853_
	);
	LUT2 #(
		.INIT('h8)
	) name596 (
		\a[88] ,
		\b[88] ,
		_w854_
	);
	LUT2 #(
		.INIT('h6)
	) name597 (
		\a[88] ,
		\b[88] ,
		_w855_
	);
	LUT4 #(
		.INIT('hc832)
	) name598 (
		\a[87] ,
		\a[88] ,
		\b[87] ,
		\b[88] ,
		_w856_
	);
	LUT4 #(
		.INIT('h4f00)
	) name599 (
		_w844_,
		_w851_,
		_w853_,
		_w856_,
		_w857_
	);
	LUT4 #(
		.INIT('h0104)
	) name600 (
		\a[87] ,
		\a[88] ,
		\b[87] ,
		\b[88] ,
		_w858_
	);
	LUT2 #(
		.INIT('h8)
	) name601 (
		_w853_,
		_w855_,
		_w859_
	);
	LUT4 #(
		.INIT('h040f)
	) name602 (
		_w844_,
		_w851_,
		_w858_,
		_w859_,
		_w860_
	);
	LUT2 #(
		.INIT('hb)
	) name603 (
		_w857_,
		_w860_,
		_w861_
	);
	LUT2 #(
		.INIT('h2)
	) name604 (
		_w853_,
		_w854_,
		_w862_
	);
	LUT4 #(
		.INIT('h0105)
	) name605 (
		\a[87] ,
		\a[88] ,
		\b[87] ,
		\b[88] ,
		_w863_
	);
	LUT2 #(
		.INIT('h8)
	) name606 (
		\a[89] ,
		\b[89] ,
		_w864_
	);
	LUT2 #(
		.INIT('h6)
	) name607 (
		\a[89] ,
		\b[89] ,
		_w865_
	);
	LUT4 #(
		.INIT('hc832)
	) name608 (
		\a[88] ,
		\a[89] ,
		\b[88] ,
		\b[89] ,
		_w866_
	);
	LUT2 #(
		.INIT('h4)
	) name609 (
		_w863_,
		_w866_,
		_w867_
	);
	LUT4 #(
		.INIT('h4f00)
	) name610 (
		_w844_,
		_w851_,
		_w862_,
		_w867_,
		_w868_
	);
	LUT4 #(
		.INIT('hfec8)
	) name611 (
		\a[87] ,
		\a[88] ,
		\b[87] ,
		\b[88] ,
		_w869_
	);
	LUT4 #(
		.INIT('h4f00)
	) name612 (
		_w844_,
		_w851_,
		_w862_,
		_w869_,
		_w870_
	);
	LUT3 #(
		.INIT('hce)
	) name613 (
		_w865_,
		_w868_,
		_w870_,
		_w871_
	);
	LUT2 #(
		.INIT('h1)
	) name614 (
		\a[90] ,
		\b[90] ,
		_w872_
	);
	LUT2 #(
		.INIT('h6)
	) name615 (
		\a[90] ,
		\b[90] ,
		_w873_
	);
	LUT4 #(
		.INIT('hfac8)
	) name616 (
		\a[88] ,
		\a[89] ,
		\b[88] ,
		\b[89] ,
		_w874_
	);
	LUT2 #(
		.INIT('h4)
	) name617 (
		_w863_,
		_w874_,
		_w875_
	);
	LUT4 #(
		.INIT('h4f00)
	) name618 (
		_w844_,
		_w851_,
		_w862_,
		_w875_,
		_w876_
	);
	LUT3 #(
		.INIT('h36)
	) name619 (
		_w864_,
		_w873_,
		_w876_,
		_w877_
	);
	LUT4 #(
		.INIT('h135f)
	) name620 (
		\a[89] ,
		\a[90] ,
		\b[89] ,
		\b[90] ,
		_w878_
	);
	LUT2 #(
		.INIT('h8)
	) name621 (
		\a[91] ,
		\b[91] ,
		_w879_
	);
	LUT2 #(
		.INIT('h6)
	) name622 (
		\a[91] ,
		\b[91] ,
		_w880_
	);
	LUT4 #(
		.INIT('hba45)
	) name623 (
		_w872_,
		_w876_,
		_w878_,
		_w880_,
		_w881_
	);
	LUT2 #(
		.INIT('h2)
	) name624 (
		_w878_,
		_w879_,
		_w882_
	);
	LUT4 #(
		.INIT('h0105)
	) name625 (
		\a[90] ,
		\a[91] ,
		\b[90] ,
		\b[91] ,
		_w883_
	);
	LUT2 #(
		.INIT('h8)
	) name626 (
		\a[92] ,
		\b[92] ,
		_w884_
	);
	LUT2 #(
		.INIT('h6)
	) name627 (
		\a[92] ,
		\b[92] ,
		_w885_
	);
	LUT4 #(
		.INIT('hc832)
	) name628 (
		\a[91] ,
		\a[92] ,
		\b[91] ,
		\b[92] ,
		_w886_
	);
	LUT2 #(
		.INIT('h4)
	) name629 (
		_w883_,
		_w886_,
		_w887_
	);
	LUT3 #(
		.INIT('hb0)
	) name630 (
		_w876_,
		_w882_,
		_w887_,
		_w888_
	);
	LUT4 #(
		.INIT('hfec8)
	) name631 (
		\a[90] ,
		\a[91] ,
		\b[90] ,
		\b[91] ,
		_w889_
	);
	LUT4 #(
		.INIT('h40f0)
	) name632 (
		_w876_,
		_w882_,
		_w885_,
		_w889_,
		_w890_
	);
	LUT2 #(
		.INIT('he)
	) name633 (
		_w888_,
		_w890_,
		_w891_
	);
	LUT2 #(
		.INIT('h1)
	) name634 (
		\a[93] ,
		\b[93] ,
		_w892_
	);
	LUT2 #(
		.INIT('h6)
	) name635 (
		\a[93] ,
		\b[93] ,
		_w893_
	);
	LUT4 #(
		.INIT('hfac8)
	) name636 (
		\a[91] ,
		\a[92] ,
		\b[91] ,
		\b[92] ,
		_w894_
	);
	LUT2 #(
		.INIT('h4)
	) name637 (
		_w883_,
		_w894_,
		_w895_
	);
	LUT3 #(
		.INIT('hb0)
	) name638 (
		_w876_,
		_w882_,
		_w895_,
		_w896_
	);
	LUT3 #(
		.INIT('h36)
	) name639 (
		_w884_,
		_w893_,
		_w896_,
		_w897_
	);
	LUT4 #(
		.INIT('h135f)
	) name640 (
		\a[92] ,
		\a[93] ,
		\b[92] ,
		\b[93] ,
		_w898_
	);
	LUT4 #(
		.INIT('h4f00)
	) name641 (
		_w876_,
		_w882_,
		_w895_,
		_w898_,
		_w899_
	);
	LUT2 #(
		.INIT('h1)
	) name642 (
		\a[94] ,
		\b[94] ,
		_w900_
	);
	LUT2 #(
		.INIT('h8)
	) name643 (
		\a[94] ,
		\b[94] ,
		_w901_
	);
	LUT2 #(
		.INIT('h6)
	) name644 (
		\a[94] ,
		\b[94] ,
		_w902_
	);
	LUT2 #(
		.INIT('h8)
	) name645 (
		_w898_,
		_w902_,
		_w903_
	);
	LUT4 #(
		.INIT('h4f00)
	) name646 (
		_w876_,
		_w882_,
		_w895_,
		_w903_,
		_w904_
	);
	LUT4 #(
		.INIT('hffa1)
	) name647 (
		_w892_,
		_w899_,
		_w902_,
		_w904_,
		_w905_
	);
	LUT2 #(
		.INIT('h2)
	) name648 (
		_w898_,
		_w901_,
		_w906_
	);
	LUT4 #(
		.INIT('h4f00)
	) name649 (
		_w876_,
		_w882_,
		_w895_,
		_w906_,
		_w907_
	);
	LUT4 #(
		.INIT('h0105)
	) name650 (
		\a[93] ,
		\a[94] ,
		\b[93] ,
		\b[94] ,
		_w908_
	);
	LUT2 #(
		.INIT('h8)
	) name651 (
		\a[95] ,
		\b[95] ,
		_w909_
	);
	LUT2 #(
		.INIT('h6)
	) name652 (
		\a[95] ,
		\b[95] ,
		_w910_
	);
	LUT4 #(
		.INIT('hfe01)
	) name653 (
		_w900_,
		_w907_,
		_w908_,
		_w910_,
		_w911_
	);
	LUT2 #(
		.INIT('h6)
	) name654 (
		\a[96] ,
		\b[96] ,
		_w912_
	);
	LUT4 #(
		.INIT('hfac8)
	) name655 (
		\a[94] ,
		\a[95] ,
		\b[94] ,
		\b[95] ,
		_w913_
	);
	LUT2 #(
		.INIT('h4)
	) name656 (
		_w908_,
		_w913_,
		_w914_
	);
	LUT4 #(
		.INIT('h2d3c)
	) name657 (
		_w907_,
		_w909_,
		_w912_,
		_w914_,
		_w915_
	);
	LUT4 #(
		.INIT('h135f)
	) name658 (
		\a[95] ,
		\a[96] ,
		\b[95] ,
		\b[96] ,
		_w916_
	);
	LUT2 #(
		.INIT('h8)
	) name659 (
		\a[97] ,
		\b[97] ,
		_w917_
	);
	LUT2 #(
		.INIT('h6)
	) name660 (
		\a[97] ,
		\b[97] ,
		_w918_
	);
	LUT4 #(
		.INIT('hc832)
	) name661 (
		\a[96] ,
		\a[97] ,
		\b[96] ,
		\b[97] ,
		_w919_
	);
	LUT4 #(
		.INIT('h4f00)
	) name662 (
		_w907_,
		_w914_,
		_w916_,
		_w919_,
		_w920_
	);
	LUT4 #(
		.INIT('h0104)
	) name663 (
		\a[96] ,
		\a[97] ,
		\b[96] ,
		\b[97] ,
		_w921_
	);
	LUT2 #(
		.INIT('h8)
	) name664 (
		_w916_,
		_w918_,
		_w922_
	);
	LUT4 #(
		.INIT('h040f)
	) name665 (
		_w907_,
		_w914_,
		_w921_,
		_w922_,
		_w923_
	);
	LUT2 #(
		.INIT('hb)
	) name666 (
		_w920_,
		_w923_,
		_w924_
	);
	LUT2 #(
		.INIT('h2)
	) name667 (
		_w916_,
		_w917_,
		_w925_
	);
	LUT4 #(
		.INIT('h0105)
	) name668 (
		\a[96] ,
		\a[97] ,
		\b[96] ,
		\b[97] ,
		_w926_
	);
	LUT2 #(
		.INIT('h8)
	) name669 (
		\a[98] ,
		\b[98] ,
		_w927_
	);
	LUT2 #(
		.INIT('h6)
	) name670 (
		\a[98] ,
		\b[98] ,
		_w928_
	);
	LUT4 #(
		.INIT('hc832)
	) name671 (
		\a[97] ,
		\a[98] ,
		\b[97] ,
		\b[98] ,
		_w929_
	);
	LUT2 #(
		.INIT('h4)
	) name672 (
		_w926_,
		_w929_,
		_w930_
	);
	LUT4 #(
		.INIT('h4f00)
	) name673 (
		_w907_,
		_w914_,
		_w925_,
		_w930_,
		_w931_
	);
	LUT4 #(
		.INIT('hfec8)
	) name674 (
		\a[96] ,
		\a[97] ,
		\b[96] ,
		\b[97] ,
		_w932_
	);
	LUT4 #(
		.INIT('h4f00)
	) name675 (
		_w907_,
		_w914_,
		_w925_,
		_w932_,
		_w933_
	);
	LUT3 #(
		.INIT('hce)
	) name676 (
		_w928_,
		_w931_,
		_w933_,
		_w934_
	);
	LUT2 #(
		.INIT('h1)
	) name677 (
		\a[99] ,
		\b[99] ,
		_w935_
	);
	LUT2 #(
		.INIT('h6)
	) name678 (
		\a[99] ,
		\b[99] ,
		_w936_
	);
	LUT4 #(
		.INIT('hfac8)
	) name679 (
		\a[97] ,
		\a[98] ,
		\b[97] ,
		\b[98] ,
		_w937_
	);
	LUT2 #(
		.INIT('h4)
	) name680 (
		_w926_,
		_w937_,
		_w938_
	);
	LUT4 #(
		.INIT('h4f00)
	) name681 (
		_w907_,
		_w914_,
		_w925_,
		_w938_,
		_w939_
	);
	LUT3 #(
		.INIT('h36)
	) name682 (
		_w927_,
		_w936_,
		_w939_,
		_w940_
	);
	LUT4 #(
		.INIT('h135f)
	) name683 (
		\a[98] ,
		\a[99] ,
		\b[98] ,
		\b[99] ,
		_w941_
	);
	LUT2 #(
		.INIT('h8)
	) name684 (
		\a[100] ,
		\b[100] ,
		_w942_
	);
	LUT2 #(
		.INIT('h6)
	) name685 (
		\a[100] ,
		\b[100] ,
		_w943_
	);
	LUT4 #(
		.INIT('hba45)
	) name686 (
		_w935_,
		_w939_,
		_w941_,
		_w943_,
		_w944_
	);
	LUT2 #(
		.INIT('h2)
	) name687 (
		_w941_,
		_w942_,
		_w945_
	);
	LUT4 #(
		.INIT('h0105)
	) name688 (
		\a[99] ,
		\a[100] ,
		\b[99] ,
		\b[100] ,
		_w946_
	);
	LUT2 #(
		.INIT('h8)
	) name689 (
		\a[101] ,
		\b[101] ,
		_w947_
	);
	LUT2 #(
		.INIT('h6)
	) name690 (
		\a[101] ,
		\b[101] ,
		_w948_
	);
	LUT4 #(
		.INIT('hc832)
	) name691 (
		\a[100] ,
		\a[101] ,
		\b[100] ,
		\b[101] ,
		_w949_
	);
	LUT2 #(
		.INIT('h4)
	) name692 (
		_w946_,
		_w949_,
		_w950_
	);
	LUT3 #(
		.INIT('hb0)
	) name693 (
		_w939_,
		_w945_,
		_w950_,
		_w951_
	);
	LUT4 #(
		.INIT('hfec8)
	) name694 (
		\a[99] ,
		\a[100] ,
		\b[99] ,
		\b[100] ,
		_w952_
	);
	LUT4 #(
		.INIT('h40f0)
	) name695 (
		_w939_,
		_w945_,
		_w948_,
		_w952_,
		_w953_
	);
	LUT2 #(
		.INIT('he)
	) name696 (
		_w951_,
		_w953_,
		_w954_
	);
	LUT2 #(
		.INIT('h1)
	) name697 (
		\a[102] ,
		\b[102] ,
		_w955_
	);
	LUT2 #(
		.INIT('h6)
	) name698 (
		\a[102] ,
		\b[102] ,
		_w956_
	);
	LUT4 #(
		.INIT('hfac8)
	) name699 (
		\a[100] ,
		\a[101] ,
		\b[100] ,
		\b[101] ,
		_w957_
	);
	LUT2 #(
		.INIT('h4)
	) name700 (
		_w946_,
		_w957_,
		_w958_
	);
	LUT3 #(
		.INIT('hb0)
	) name701 (
		_w939_,
		_w945_,
		_w958_,
		_w959_
	);
	LUT3 #(
		.INIT('h36)
	) name702 (
		_w947_,
		_w956_,
		_w959_,
		_w960_
	);
	LUT4 #(
		.INIT('h135f)
	) name703 (
		\a[101] ,
		\a[102] ,
		\b[101] ,
		\b[102] ,
		_w961_
	);
	LUT4 #(
		.INIT('h4f00)
	) name704 (
		_w939_,
		_w945_,
		_w958_,
		_w961_,
		_w962_
	);
	LUT2 #(
		.INIT('h1)
	) name705 (
		\a[103] ,
		\b[103] ,
		_w963_
	);
	LUT2 #(
		.INIT('h8)
	) name706 (
		\a[103] ,
		\b[103] ,
		_w964_
	);
	LUT2 #(
		.INIT('h6)
	) name707 (
		\a[103] ,
		\b[103] ,
		_w965_
	);
	LUT2 #(
		.INIT('h8)
	) name708 (
		_w961_,
		_w965_,
		_w966_
	);
	LUT4 #(
		.INIT('h4f00)
	) name709 (
		_w939_,
		_w945_,
		_w958_,
		_w966_,
		_w967_
	);
	LUT4 #(
		.INIT('hffa1)
	) name710 (
		_w955_,
		_w962_,
		_w965_,
		_w967_,
		_w968_
	);
	LUT2 #(
		.INIT('h2)
	) name711 (
		_w961_,
		_w964_,
		_w969_
	);
	LUT4 #(
		.INIT('h4f00)
	) name712 (
		_w939_,
		_w945_,
		_w958_,
		_w969_,
		_w970_
	);
	LUT4 #(
		.INIT('h0105)
	) name713 (
		\a[102] ,
		\a[103] ,
		\b[102] ,
		\b[103] ,
		_w971_
	);
	LUT2 #(
		.INIT('h8)
	) name714 (
		\a[104] ,
		\b[104] ,
		_w972_
	);
	LUT2 #(
		.INIT('h6)
	) name715 (
		\a[104] ,
		\b[104] ,
		_w973_
	);
	LUT4 #(
		.INIT('hfe01)
	) name716 (
		_w963_,
		_w970_,
		_w971_,
		_w973_,
		_w974_
	);
	LUT2 #(
		.INIT('h6)
	) name717 (
		\a[105] ,
		\b[105] ,
		_w975_
	);
	LUT4 #(
		.INIT('hfac8)
	) name718 (
		\a[103] ,
		\a[104] ,
		\b[103] ,
		\b[104] ,
		_w976_
	);
	LUT2 #(
		.INIT('h4)
	) name719 (
		_w971_,
		_w976_,
		_w977_
	);
	LUT4 #(
		.INIT('h2d3c)
	) name720 (
		_w970_,
		_w972_,
		_w975_,
		_w977_,
		_w978_
	);
	LUT4 #(
		.INIT('h135f)
	) name721 (
		\a[104] ,
		\a[105] ,
		\b[104] ,
		\b[105] ,
		_w979_
	);
	LUT2 #(
		.INIT('h8)
	) name722 (
		\a[106] ,
		\b[106] ,
		_w980_
	);
	LUT2 #(
		.INIT('h6)
	) name723 (
		\a[106] ,
		\b[106] ,
		_w981_
	);
	LUT4 #(
		.INIT('hc832)
	) name724 (
		\a[105] ,
		\a[106] ,
		\b[105] ,
		\b[106] ,
		_w982_
	);
	LUT4 #(
		.INIT('h4f00)
	) name725 (
		_w970_,
		_w977_,
		_w979_,
		_w982_,
		_w983_
	);
	LUT4 #(
		.INIT('h0104)
	) name726 (
		\a[105] ,
		\a[106] ,
		\b[105] ,
		\b[106] ,
		_w984_
	);
	LUT2 #(
		.INIT('h8)
	) name727 (
		_w979_,
		_w981_,
		_w985_
	);
	LUT4 #(
		.INIT('h040f)
	) name728 (
		_w970_,
		_w977_,
		_w984_,
		_w985_,
		_w986_
	);
	LUT2 #(
		.INIT('hb)
	) name729 (
		_w983_,
		_w986_,
		_w987_
	);
	LUT2 #(
		.INIT('h2)
	) name730 (
		_w979_,
		_w980_,
		_w988_
	);
	LUT4 #(
		.INIT('h0105)
	) name731 (
		\a[105] ,
		\a[106] ,
		\b[105] ,
		\b[106] ,
		_w989_
	);
	LUT2 #(
		.INIT('h8)
	) name732 (
		\a[107] ,
		\b[107] ,
		_w990_
	);
	LUT2 #(
		.INIT('h6)
	) name733 (
		\a[107] ,
		\b[107] ,
		_w991_
	);
	LUT4 #(
		.INIT('hc832)
	) name734 (
		\a[106] ,
		\a[107] ,
		\b[106] ,
		\b[107] ,
		_w992_
	);
	LUT2 #(
		.INIT('h4)
	) name735 (
		_w989_,
		_w992_,
		_w993_
	);
	LUT4 #(
		.INIT('h4f00)
	) name736 (
		_w970_,
		_w977_,
		_w988_,
		_w993_,
		_w994_
	);
	LUT4 #(
		.INIT('hfec8)
	) name737 (
		\a[105] ,
		\a[106] ,
		\b[105] ,
		\b[106] ,
		_w995_
	);
	LUT4 #(
		.INIT('h4f00)
	) name738 (
		_w970_,
		_w977_,
		_w988_,
		_w995_,
		_w996_
	);
	LUT3 #(
		.INIT('hce)
	) name739 (
		_w991_,
		_w994_,
		_w996_,
		_w997_
	);
	LUT2 #(
		.INIT('h1)
	) name740 (
		\a[108] ,
		\b[108] ,
		_w998_
	);
	LUT2 #(
		.INIT('h6)
	) name741 (
		\a[108] ,
		\b[108] ,
		_w999_
	);
	LUT4 #(
		.INIT('hfac8)
	) name742 (
		\a[106] ,
		\a[107] ,
		\b[106] ,
		\b[107] ,
		_w1000_
	);
	LUT2 #(
		.INIT('h4)
	) name743 (
		_w989_,
		_w1000_,
		_w1001_
	);
	LUT4 #(
		.INIT('h4f00)
	) name744 (
		_w970_,
		_w977_,
		_w988_,
		_w1001_,
		_w1002_
	);
	LUT3 #(
		.INIT('h36)
	) name745 (
		_w990_,
		_w999_,
		_w1002_,
		_w1003_
	);
	LUT4 #(
		.INIT('h135f)
	) name746 (
		\a[107] ,
		\a[108] ,
		\b[107] ,
		\b[108] ,
		_w1004_
	);
	LUT2 #(
		.INIT('h8)
	) name747 (
		\a[109] ,
		\b[109] ,
		_w1005_
	);
	LUT2 #(
		.INIT('h6)
	) name748 (
		\a[109] ,
		\b[109] ,
		_w1006_
	);
	LUT4 #(
		.INIT('hba45)
	) name749 (
		_w998_,
		_w1002_,
		_w1004_,
		_w1006_,
		_w1007_
	);
	LUT2 #(
		.INIT('h2)
	) name750 (
		_w1004_,
		_w1005_,
		_w1008_
	);
	LUT4 #(
		.INIT('h0105)
	) name751 (
		\a[108] ,
		\a[109] ,
		\b[108] ,
		\b[109] ,
		_w1009_
	);
	LUT2 #(
		.INIT('h8)
	) name752 (
		\a[110] ,
		\b[110] ,
		_w1010_
	);
	LUT2 #(
		.INIT('h6)
	) name753 (
		\a[110] ,
		\b[110] ,
		_w1011_
	);
	LUT4 #(
		.INIT('hc832)
	) name754 (
		\a[109] ,
		\a[110] ,
		\b[109] ,
		\b[110] ,
		_w1012_
	);
	LUT2 #(
		.INIT('h4)
	) name755 (
		_w1009_,
		_w1012_,
		_w1013_
	);
	LUT3 #(
		.INIT('hb0)
	) name756 (
		_w1002_,
		_w1008_,
		_w1013_,
		_w1014_
	);
	LUT4 #(
		.INIT('hfec8)
	) name757 (
		\a[108] ,
		\a[109] ,
		\b[108] ,
		\b[109] ,
		_w1015_
	);
	LUT4 #(
		.INIT('h40f0)
	) name758 (
		_w1002_,
		_w1008_,
		_w1011_,
		_w1015_,
		_w1016_
	);
	LUT2 #(
		.INIT('he)
	) name759 (
		_w1014_,
		_w1016_,
		_w1017_
	);
	LUT2 #(
		.INIT('h1)
	) name760 (
		\a[111] ,
		\b[111] ,
		_w1018_
	);
	LUT2 #(
		.INIT('h6)
	) name761 (
		\a[111] ,
		\b[111] ,
		_w1019_
	);
	LUT4 #(
		.INIT('hfac8)
	) name762 (
		\a[109] ,
		\a[110] ,
		\b[109] ,
		\b[110] ,
		_w1020_
	);
	LUT2 #(
		.INIT('h4)
	) name763 (
		_w1009_,
		_w1020_,
		_w1021_
	);
	LUT3 #(
		.INIT('hb0)
	) name764 (
		_w1002_,
		_w1008_,
		_w1021_,
		_w1022_
	);
	LUT3 #(
		.INIT('h36)
	) name765 (
		_w1010_,
		_w1019_,
		_w1022_,
		_w1023_
	);
	LUT4 #(
		.INIT('h135f)
	) name766 (
		\a[110] ,
		\a[111] ,
		\b[110] ,
		\b[111] ,
		_w1024_
	);
	LUT4 #(
		.INIT('h4f00)
	) name767 (
		_w1002_,
		_w1008_,
		_w1021_,
		_w1024_,
		_w1025_
	);
	LUT2 #(
		.INIT('h1)
	) name768 (
		\a[112] ,
		\b[112] ,
		_w1026_
	);
	LUT2 #(
		.INIT('h8)
	) name769 (
		\a[112] ,
		\b[112] ,
		_w1027_
	);
	LUT2 #(
		.INIT('h6)
	) name770 (
		\a[112] ,
		\b[112] ,
		_w1028_
	);
	LUT2 #(
		.INIT('h8)
	) name771 (
		_w1024_,
		_w1028_,
		_w1029_
	);
	LUT4 #(
		.INIT('h4f00)
	) name772 (
		_w1002_,
		_w1008_,
		_w1021_,
		_w1029_,
		_w1030_
	);
	LUT4 #(
		.INIT('hffa1)
	) name773 (
		_w1018_,
		_w1025_,
		_w1028_,
		_w1030_,
		_w1031_
	);
	LUT2 #(
		.INIT('h2)
	) name774 (
		_w1024_,
		_w1027_,
		_w1032_
	);
	LUT4 #(
		.INIT('h4f00)
	) name775 (
		_w1002_,
		_w1008_,
		_w1021_,
		_w1032_,
		_w1033_
	);
	LUT4 #(
		.INIT('h0105)
	) name776 (
		\a[111] ,
		\a[112] ,
		\b[111] ,
		\b[112] ,
		_w1034_
	);
	LUT2 #(
		.INIT('h8)
	) name777 (
		\a[113] ,
		\b[113] ,
		_w1035_
	);
	LUT2 #(
		.INIT('h6)
	) name778 (
		\a[113] ,
		\b[113] ,
		_w1036_
	);
	LUT4 #(
		.INIT('hfe01)
	) name779 (
		_w1026_,
		_w1033_,
		_w1034_,
		_w1036_,
		_w1037_
	);
	LUT2 #(
		.INIT('h6)
	) name780 (
		\a[114] ,
		\b[114] ,
		_w1038_
	);
	LUT4 #(
		.INIT('hfac8)
	) name781 (
		\a[112] ,
		\a[113] ,
		\b[112] ,
		\b[113] ,
		_w1039_
	);
	LUT2 #(
		.INIT('h4)
	) name782 (
		_w1034_,
		_w1039_,
		_w1040_
	);
	LUT4 #(
		.INIT('h2d3c)
	) name783 (
		_w1033_,
		_w1035_,
		_w1038_,
		_w1040_,
		_w1041_
	);
	LUT4 #(
		.INIT('h135f)
	) name784 (
		\a[113] ,
		\a[114] ,
		\b[113] ,
		\b[114] ,
		_w1042_
	);
	LUT2 #(
		.INIT('h8)
	) name785 (
		\a[115] ,
		\b[115] ,
		_w1043_
	);
	LUT2 #(
		.INIT('h6)
	) name786 (
		\a[115] ,
		\b[115] ,
		_w1044_
	);
	LUT4 #(
		.INIT('hc832)
	) name787 (
		\a[114] ,
		\a[115] ,
		\b[114] ,
		\b[115] ,
		_w1045_
	);
	LUT4 #(
		.INIT('h4f00)
	) name788 (
		_w1033_,
		_w1040_,
		_w1042_,
		_w1045_,
		_w1046_
	);
	LUT4 #(
		.INIT('h0104)
	) name789 (
		\a[114] ,
		\a[115] ,
		\b[114] ,
		\b[115] ,
		_w1047_
	);
	LUT2 #(
		.INIT('h8)
	) name790 (
		_w1042_,
		_w1044_,
		_w1048_
	);
	LUT4 #(
		.INIT('h040f)
	) name791 (
		_w1033_,
		_w1040_,
		_w1047_,
		_w1048_,
		_w1049_
	);
	LUT2 #(
		.INIT('hb)
	) name792 (
		_w1046_,
		_w1049_,
		_w1050_
	);
	LUT2 #(
		.INIT('h2)
	) name793 (
		_w1042_,
		_w1043_,
		_w1051_
	);
	LUT4 #(
		.INIT('h0105)
	) name794 (
		\a[114] ,
		\a[115] ,
		\b[114] ,
		\b[115] ,
		_w1052_
	);
	LUT2 #(
		.INIT('h8)
	) name795 (
		\a[116] ,
		\b[116] ,
		_w1053_
	);
	LUT2 #(
		.INIT('h6)
	) name796 (
		\a[116] ,
		\b[116] ,
		_w1054_
	);
	LUT4 #(
		.INIT('hc832)
	) name797 (
		\a[115] ,
		\a[116] ,
		\b[115] ,
		\b[116] ,
		_w1055_
	);
	LUT2 #(
		.INIT('h4)
	) name798 (
		_w1052_,
		_w1055_,
		_w1056_
	);
	LUT4 #(
		.INIT('h4f00)
	) name799 (
		_w1033_,
		_w1040_,
		_w1051_,
		_w1056_,
		_w1057_
	);
	LUT4 #(
		.INIT('hfec8)
	) name800 (
		\a[114] ,
		\a[115] ,
		\b[114] ,
		\b[115] ,
		_w1058_
	);
	LUT4 #(
		.INIT('h4f00)
	) name801 (
		_w1033_,
		_w1040_,
		_w1051_,
		_w1058_,
		_w1059_
	);
	LUT3 #(
		.INIT('hce)
	) name802 (
		_w1054_,
		_w1057_,
		_w1059_,
		_w1060_
	);
	LUT2 #(
		.INIT('h1)
	) name803 (
		\a[117] ,
		\b[117] ,
		_w1061_
	);
	LUT2 #(
		.INIT('h6)
	) name804 (
		\a[117] ,
		\b[117] ,
		_w1062_
	);
	LUT4 #(
		.INIT('hfac8)
	) name805 (
		\a[115] ,
		\a[116] ,
		\b[115] ,
		\b[116] ,
		_w1063_
	);
	LUT2 #(
		.INIT('h4)
	) name806 (
		_w1052_,
		_w1063_,
		_w1064_
	);
	LUT4 #(
		.INIT('h4f00)
	) name807 (
		_w1033_,
		_w1040_,
		_w1051_,
		_w1064_,
		_w1065_
	);
	LUT3 #(
		.INIT('h36)
	) name808 (
		_w1053_,
		_w1062_,
		_w1065_,
		_w1066_
	);
	LUT4 #(
		.INIT('h135f)
	) name809 (
		\a[116] ,
		\a[117] ,
		\b[116] ,
		\b[117] ,
		_w1067_
	);
	LUT2 #(
		.INIT('h8)
	) name810 (
		\a[118] ,
		\b[118] ,
		_w1068_
	);
	LUT2 #(
		.INIT('h6)
	) name811 (
		\a[118] ,
		\b[118] ,
		_w1069_
	);
	LUT4 #(
		.INIT('hba45)
	) name812 (
		_w1061_,
		_w1065_,
		_w1067_,
		_w1069_,
		_w1070_
	);
	LUT2 #(
		.INIT('h2)
	) name813 (
		_w1067_,
		_w1068_,
		_w1071_
	);
	LUT4 #(
		.INIT('h0105)
	) name814 (
		\a[117] ,
		\a[118] ,
		\b[117] ,
		\b[118] ,
		_w1072_
	);
	LUT2 #(
		.INIT('h8)
	) name815 (
		\a[119] ,
		\b[119] ,
		_w1073_
	);
	LUT2 #(
		.INIT('h6)
	) name816 (
		\a[119] ,
		\b[119] ,
		_w1074_
	);
	LUT4 #(
		.INIT('hc832)
	) name817 (
		\a[118] ,
		\a[119] ,
		\b[118] ,
		\b[119] ,
		_w1075_
	);
	LUT2 #(
		.INIT('h4)
	) name818 (
		_w1072_,
		_w1075_,
		_w1076_
	);
	LUT3 #(
		.INIT('hb0)
	) name819 (
		_w1065_,
		_w1071_,
		_w1076_,
		_w1077_
	);
	LUT4 #(
		.INIT('hfec8)
	) name820 (
		\a[117] ,
		\a[118] ,
		\b[117] ,
		\b[118] ,
		_w1078_
	);
	LUT4 #(
		.INIT('h40f0)
	) name821 (
		_w1065_,
		_w1071_,
		_w1074_,
		_w1078_,
		_w1079_
	);
	LUT2 #(
		.INIT('he)
	) name822 (
		_w1077_,
		_w1079_,
		_w1080_
	);
	LUT2 #(
		.INIT('h1)
	) name823 (
		\a[120] ,
		\b[120] ,
		_w1081_
	);
	LUT2 #(
		.INIT('h6)
	) name824 (
		\a[120] ,
		\b[120] ,
		_w1082_
	);
	LUT4 #(
		.INIT('hfac8)
	) name825 (
		\a[118] ,
		\a[119] ,
		\b[118] ,
		\b[119] ,
		_w1083_
	);
	LUT2 #(
		.INIT('h4)
	) name826 (
		_w1072_,
		_w1083_,
		_w1084_
	);
	LUT3 #(
		.INIT('hb0)
	) name827 (
		_w1065_,
		_w1071_,
		_w1084_,
		_w1085_
	);
	LUT3 #(
		.INIT('h36)
	) name828 (
		_w1073_,
		_w1082_,
		_w1085_,
		_w1086_
	);
	LUT4 #(
		.INIT('h135f)
	) name829 (
		\a[119] ,
		\a[120] ,
		\b[119] ,
		\b[120] ,
		_w1087_
	);
	LUT4 #(
		.INIT('h4f00)
	) name830 (
		_w1065_,
		_w1071_,
		_w1084_,
		_w1087_,
		_w1088_
	);
	LUT2 #(
		.INIT('h1)
	) name831 (
		\a[121] ,
		\b[121] ,
		_w1089_
	);
	LUT2 #(
		.INIT('h8)
	) name832 (
		\a[121] ,
		\b[121] ,
		_w1090_
	);
	LUT2 #(
		.INIT('h6)
	) name833 (
		\a[121] ,
		\b[121] ,
		_w1091_
	);
	LUT2 #(
		.INIT('h8)
	) name834 (
		_w1087_,
		_w1091_,
		_w1092_
	);
	LUT4 #(
		.INIT('h4f00)
	) name835 (
		_w1065_,
		_w1071_,
		_w1084_,
		_w1092_,
		_w1093_
	);
	LUT4 #(
		.INIT('hffa1)
	) name836 (
		_w1081_,
		_w1088_,
		_w1091_,
		_w1093_,
		_w1094_
	);
	LUT2 #(
		.INIT('h2)
	) name837 (
		_w1087_,
		_w1090_,
		_w1095_
	);
	LUT4 #(
		.INIT('h4f00)
	) name838 (
		_w1065_,
		_w1071_,
		_w1084_,
		_w1095_,
		_w1096_
	);
	LUT4 #(
		.INIT('h0105)
	) name839 (
		\a[120] ,
		\a[121] ,
		\b[120] ,
		\b[121] ,
		_w1097_
	);
	LUT2 #(
		.INIT('h8)
	) name840 (
		\a[122] ,
		\b[122] ,
		_w1098_
	);
	LUT2 #(
		.INIT('h6)
	) name841 (
		\a[122] ,
		\b[122] ,
		_w1099_
	);
	LUT4 #(
		.INIT('hfe01)
	) name842 (
		_w1089_,
		_w1096_,
		_w1097_,
		_w1099_,
		_w1100_
	);
	LUT2 #(
		.INIT('h6)
	) name843 (
		\a[123] ,
		\b[123] ,
		_w1101_
	);
	LUT4 #(
		.INIT('hfac8)
	) name844 (
		\a[121] ,
		\a[122] ,
		\b[121] ,
		\b[122] ,
		_w1102_
	);
	LUT2 #(
		.INIT('h4)
	) name845 (
		_w1097_,
		_w1102_,
		_w1103_
	);
	LUT4 #(
		.INIT('h2d3c)
	) name846 (
		_w1096_,
		_w1098_,
		_w1101_,
		_w1103_,
		_w1104_
	);
	LUT4 #(
		.INIT('h135f)
	) name847 (
		\a[122] ,
		\a[123] ,
		\b[122] ,
		\b[123] ,
		_w1105_
	);
	LUT2 #(
		.INIT('h8)
	) name848 (
		\a[124] ,
		\b[124] ,
		_w1106_
	);
	LUT2 #(
		.INIT('h6)
	) name849 (
		\a[124] ,
		\b[124] ,
		_w1107_
	);
	LUT4 #(
		.INIT('hc832)
	) name850 (
		\a[123] ,
		\a[124] ,
		\b[123] ,
		\b[124] ,
		_w1108_
	);
	LUT4 #(
		.INIT('h4f00)
	) name851 (
		_w1096_,
		_w1103_,
		_w1105_,
		_w1108_,
		_w1109_
	);
	LUT4 #(
		.INIT('h0104)
	) name852 (
		\a[123] ,
		\a[124] ,
		\b[123] ,
		\b[124] ,
		_w1110_
	);
	LUT2 #(
		.INIT('h8)
	) name853 (
		_w1105_,
		_w1107_,
		_w1111_
	);
	LUT4 #(
		.INIT('h040f)
	) name854 (
		_w1096_,
		_w1103_,
		_w1110_,
		_w1111_,
		_w1112_
	);
	LUT2 #(
		.INIT('hb)
	) name855 (
		_w1109_,
		_w1112_,
		_w1113_
	);
	LUT2 #(
		.INIT('h2)
	) name856 (
		_w1105_,
		_w1106_,
		_w1114_
	);
	LUT4 #(
		.INIT('h0105)
	) name857 (
		\a[123] ,
		\a[124] ,
		\b[123] ,
		\b[124] ,
		_w1115_
	);
	LUT2 #(
		.INIT('h8)
	) name858 (
		\a[125] ,
		\b[125] ,
		_w1116_
	);
	LUT2 #(
		.INIT('h6)
	) name859 (
		\a[125] ,
		\b[125] ,
		_w1117_
	);
	LUT4 #(
		.INIT('hc832)
	) name860 (
		\a[124] ,
		\a[125] ,
		\b[124] ,
		\b[125] ,
		_w1118_
	);
	LUT2 #(
		.INIT('h4)
	) name861 (
		_w1115_,
		_w1118_,
		_w1119_
	);
	LUT4 #(
		.INIT('h4f00)
	) name862 (
		_w1096_,
		_w1103_,
		_w1114_,
		_w1119_,
		_w1120_
	);
	LUT4 #(
		.INIT('hfec8)
	) name863 (
		\a[123] ,
		\a[124] ,
		\b[123] ,
		\b[124] ,
		_w1121_
	);
	LUT4 #(
		.INIT('h4f00)
	) name864 (
		_w1096_,
		_w1103_,
		_w1114_,
		_w1121_,
		_w1122_
	);
	LUT3 #(
		.INIT('hce)
	) name865 (
		_w1117_,
		_w1120_,
		_w1122_,
		_w1123_
	);
	LUT2 #(
		.INIT('h1)
	) name866 (
		\a[126] ,
		\b[126] ,
		_w1124_
	);
	LUT2 #(
		.INIT('h6)
	) name867 (
		\a[126] ,
		\b[126] ,
		_w1125_
	);
	LUT4 #(
		.INIT('hfac8)
	) name868 (
		\a[124] ,
		\a[125] ,
		\b[124] ,
		\b[125] ,
		_w1126_
	);
	LUT2 #(
		.INIT('h4)
	) name869 (
		_w1115_,
		_w1126_,
		_w1127_
	);
	LUT4 #(
		.INIT('h4f00)
	) name870 (
		_w1096_,
		_w1103_,
		_w1114_,
		_w1127_,
		_w1128_
	);
	LUT3 #(
		.INIT('h36)
	) name871 (
		_w1116_,
		_w1125_,
		_w1128_,
		_w1129_
	);
	LUT4 #(
		.INIT('h135f)
	) name872 (
		\a[125] ,
		\a[126] ,
		\b[125] ,
		\b[126] ,
		_w1130_
	);
	LUT2 #(
		.INIT('h8)
	) name873 (
		\a[127] ,
		\b[127] ,
		_w1131_
	);
	LUT2 #(
		.INIT('h6)
	) name874 (
		\a[127] ,
		\b[127] ,
		_w1132_
	);
	LUT4 #(
		.INIT('hba45)
	) name875 (
		_w1124_,
		_w1128_,
		_w1130_,
		_w1132_,
		_w1133_
	);
	LUT2 #(
		.INIT('h2)
	) name876 (
		_w1130_,
		_w1131_,
		_w1134_
	);
	LUT4 #(
		.INIT('hfec8)
	) name877 (
		\a[126] ,
		\a[127] ,
		\b[126] ,
		\b[127] ,
		_w1135_
	);
	LUT3 #(
		.INIT('hb0)
	) name878 (
		_w1128_,
		_w1134_,
		_w1135_,
		_w1136_
	);
	assign \f[0]  = _w258_ ;
	assign \f[1]  = _w259_ ;
	assign \f[2]  = _w264_ ;
	assign \f[3]  = _w267_ ;
	assign \f[4]  = _w276_ ;
	assign \f[5]  = _w281_ ;
	assign \f[6]  = _w285_ ;
	assign \f[7]  = _w294_ ;
	assign \f[8]  = _w304_ ;
	assign \f[9]  = _w310_ ;
	assign \f[10]  = _w314_ ;
	assign \f[11]  = _w324_ ;
	assign \f[12]  = _w330_ ;
	assign \f[13]  = _w338_ ;
	assign \f[14]  = _w344_ ;
	assign \f[15]  = _w348_ ;
	assign \f[16]  = _w357_ ;
	assign \f[17]  = _w367_ ;
	assign \f[18]  = _w373_ ;
	assign \f[19]  = _w377_ ;
	assign \f[20]  = _w387_ ;
	assign \f[21]  = _w393_ ;
	assign \f[22]  = _w401_ ;
	assign \f[23]  = _w407_ ;
	assign \f[24]  = _w411_ ;
	assign \f[25]  = _w420_ ;
	assign \f[26]  = _w430_ ;
	assign \f[27]  = _w436_ ;
	assign \f[28]  = _w440_ ;
	assign \f[29]  = _w450_ ;
	assign \f[30]  = _w456_ ;
	assign \f[31]  = _w464_ ;
	assign \f[32]  = _w470_ ;
	assign \f[33]  = _w474_ ;
	assign \f[34]  = _w483_ ;
	assign \f[35]  = _w493_ ;
	assign \f[36]  = _w499_ ;
	assign \f[37]  = _w503_ ;
	assign \f[38]  = _w513_ ;
	assign \f[39]  = _w519_ ;
	assign \f[40]  = _w527_ ;
	assign \f[41]  = _w533_ ;
	assign \f[42]  = _w537_ ;
	assign \f[43]  = _w546_ ;
	assign \f[44]  = _w556_ ;
	assign \f[45]  = _w562_ ;
	assign \f[46]  = _w566_ ;
	assign \f[47]  = _w576_ ;
	assign \f[48]  = _w582_ ;
	assign \f[49]  = _w590_ ;
	assign \f[50]  = _w596_ ;
	assign \f[51]  = _w600_ ;
	assign \f[52]  = _w609_ ;
	assign \f[53]  = _w619_ ;
	assign \f[54]  = _w625_ ;
	assign \f[55]  = _w629_ ;
	assign \f[56]  = _w639_ ;
	assign \f[57]  = _w645_ ;
	assign \f[58]  = _w653_ ;
	assign \f[59]  = _w659_ ;
	assign \f[60]  = _w663_ ;
	assign \f[61]  = _w672_ ;
	assign \f[62]  = _w682_ ;
	assign \f[63]  = _w688_ ;
	assign \f[64]  = _w692_ ;
	assign \f[65]  = _w702_ ;
	assign \f[66]  = _w708_ ;
	assign \f[67]  = _w716_ ;
	assign \f[68]  = _w722_ ;
	assign \f[69]  = _w726_ ;
	assign \f[70]  = _w735_ ;
	assign \f[71]  = _w745_ ;
	assign \f[72]  = _w751_ ;
	assign \f[73]  = _w755_ ;
	assign \f[74]  = _w765_ ;
	assign \f[75]  = _w771_ ;
	assign \f[76]  = _w779_ ;
	assign \f[77]  = _w785_ ;
	assign \f[78]  = _w789_ ;
	assign \f[79]  = _w798_ ;
	assign \f[80]  = _w808_ ;
	assign \f[81]  = _w814_ ;
	assign \f[82]  = _w818_ ;
	assign \f[83]  = _w828_ ;
	assign \f[84]  = _w834_ ;
	assign \f[85]  = _w842_ ;
	assign \f[86]  = _w848_ ;
	assign \f[87]  = _w852_ ;
	assign \f[88]  = _w861_ ;
	assign \f[89]  = _w871_ ;
	assign \f[90]  = _w877_ ;
	assign \f[91]  = _w881_ ;
	assign \f[92]  = _w891_ ;
	assign \f[93]  = _w897_ ;
	assign \f[94]  = _w905_ ;
	assign \f[95]  = _w911_ ;
	assign \f[96]  = _w915_ ;
	assign \f[97]  = _w924_ ;
	assign \f[98]  = _w934_ ;
	assign \f[99]  = _w940_ ;
	assign \f[100]  = _w944_ ;
	assign \f[101]  = _w954_ ;
	assign \f[102]  = _w960_ ;
	assign \f[103]  = _w968_ ;
	assign \f[104]  = _w974_ ;
	assign \f[105]  = _w978_ ;
	assign \f[106]  = _w987_ ;
	assign \f[107]  = _w997_ ;
	assign \f[108]  = _w1003_ ;
	assign \f[109]  = _w1007_ ;
	assign \f[110]  = _w1017_ ;
	assign \f[111]  = _w1023_ ;
	assign \f[112]  = _w1031_ ;
	assign \f[113]  = _w1037_ ;
	assign \f[114]  = _w1041_ ;
	assign \f[115]  = _w1050_ ;
	assign \f[116]  = _w1060_ ;
	assign \f[117]  = _w1066_ ;
	assign \f[118]  = _w1070_ ;
	assign \f[119]  = _w1080_ ;
	assign \f[120]  = _w1086_ ;
	assign \f[121]  = _w1094_ ;
	assign \f[122]  = _w1100_ ;
	assign \f[123]  = _w1104_ ;
	assign \f[124]  = _w1113_ ;
	assign \f[125]  = _w1123_ ;
	assign \f[126]  = _w1129_ ;
	assign \f[127]  = _w1133_ ;
	assign cOut = _w1136_ ;
endmodule;