module top (\coda0_reg[0]/NET0131 , \coda0_reg[1]/NET0131 , \coda0_reg[2]/NET0131 , \coda1_reg[0]/NET0131 , \coda1_reg[1]/NET0131 , \coda1_reg[2]/NET0131 , \coda2_reg[0]/NET0131 , \coda2_reg[1]/NET0131 , \coda2_reg[2]/NET0131 , \coda3_reg[0]/NET0131 , \coda3_reg[1]/NET0131 , \coda3_reg[2]/NET0131 , \fu1_reg/NET0131 , \fu2_reg/NET0131 , \fu3_reg/NET0131 , \fu4_reg/NET0131 , \grant_o[0]_pad , \grant_o[1]_pad , \grant_o[2]_pad , \grant_o[3]_pad , \grant_reg[0]/NET0131 , \grant_reg[1]/NET0131 , \grant_reg[2]/NET0131 , \grant_reg[3]/NET0131 , \request1_pad , \request2_pad , \request3_pad , \request4_pad , \ru1_reg/NET0131 , \ru2_reg/NET0131 , \ru3_reg/NET0131 , \ru4_reg/NET0131 , \stato_reg[0]/NET0131 , \stato_reg[1]/NET0131 , \_al_n0 , \_al_n1 , \g1143/_0_ , \g1144/_0_ , \g1145/_0_ , \g1146/_0_ , \g1147/_0_ , \g1148/_0_ , \g1149/_0_ , \g1150/_0_ , \g1151/_0_ , \g1152/_0_ , \g1153/_0_ , \g1154/_0_ , \g1174/_0_ , \g1175/_0_ , \g1176/_0_ , \g1177/_0_ , \g1238/_0_ , \g1239/_0_ , \g1240/_0_ , \g1241/_0_ , \g1242/_0_ , \g1243/_0_ , \g1244/_0_ , \g1245/_0_ , \g1247/_0_ , \g1248/_0_ , \g1249/_0_ , \g1250/_0_ , \g1520/_0_ );
	input \coda0_reg[0]/NET0131  ;
	input \coda0_reg[1]/NET0131  ;
	input \coda0_reg[2]/NET0131  ;
	input \coda1_reg[0]/NET0131  ;
	input \coda1_reg[1]/NET0131  ;
	input \coda1_reg[2]/NET0131  ;
	input \coda2_reg[0]/NET0131  ;
	input \coda2_reg[1]/NET0131  ;
	input \coda2_reg[2]/NET0131  ;
	input \coda3_reg[0]/NET0131  ;
	input \coda3_reg[1]/NET0131  ;
	input \coda3_reg[2]/NET0131  ;
	input \fu1_reg/NET0131  ;
	input \fu2_reg/NET0131  ;
	input \fu3_reg/NET0131  ;
	input \fu4_reg/NET0131  ;
	input \grant_o[0]_pad  ;
	input \grant_o[1]_pad  ;
	input \grant_o[2]_pad  ;
	input \grant_o[3]_pad  ;
	input \grant_reg[0]/NET0131  ;
	input \grant_reg[1]/NET0131  ;
	input \grant_reg[2]/NET0131  ;
	input \grant_reg[3]/NET0131  ;
	input \request1_pad  ;
	input \request2_pad  ;
	input \request3_pad  ;
	input \request4_pad  ;
	input \ru1_reg/NET0131  ;
	input \ru2_reg/NET0131  ;
	input \ru3_reg/NET0131  ;
	input \ru4_reg/NET0131  ;
	input \stato_reg[0]/NET0131  ;
	input \stato_reg[1]/NET0131  ;
	output \_al_n0  ;
	output \_al_n1  ;
	output \g1143/_0_  ;
	output \g1144/_0_  ;
	output \g1145/_0_  ;
	output \g1146/_0_  ;
	output \g1147/_0_  ;
	output \g1148/_0_  ;
	output \g1149/_0_  ;
	output \g1150/_0_  ;
	output \g1151/_0_  ;
	output \g1152/_0_  ;
	output \g1153/_0_  ;
	output \g1154/_0_  ;
	output \g1174/_0_  ;
	output \g1175/_0_  ;
	output \g1176/_0_  ;
	output \g1177/_0_  ;
	output \g1238/_0_  ;
	output \g1239/_0_  ;
	output \g1240/_0_  ;
	output \g1241/_0_  ;
	output \g1242/_0_  ;
	output \g1243/_0_  ;
	output \g1244/_0_  ;
	output \g1245/_0_  ;
	output \g1247/_0_  ;
	output \g1248/_0_  ;
	output \g1249/_0_  ;
	output \g1250/_0_  ;
	output \g1520/_0_  ;
	wire _w203_ ;
	wire _w202_ ;
	wire _w201_ ;
	wire _w200_ ;
	wire _w199_ ;
	wire _w198_ ;
	wire _w197_ ;
	wire _w196_ ;
	wire _w195_ ;
	wire _w194_ ;
	wire _w193_ ;
	wire _w192_ ;
	wire _w191_ ;
	wire _w190_ ;
	wire _w189_ ;
	wire _w188_ ;
	wire _w187_ ;
	wire _w186_ ;
	wire _w185_ ;
	wire _w184_ ;
	wire _w183_ ;
	wire _w182_ ;
	wire _w181_ ;
	wire _w180_ ;
	wire _w179_ ;
	wire _w178_ ;
	wire _w177_ ;
	wire _w176_ ;
	wire _w175_ ;
	wire _w174_ ;
	wire _w173_ ;
	wire _w172_ ;
	wire _w171_ ;
	wire _w170_ ;
	wire _w169_ ;
	wire _w168_ ;
	wire _w167_ ;
	wire _w166_ ;
	wire _w165_ ;
	wire _w164_ ;
	wire _w163_ ;
	wire _w93_ ;
	wire _w92_ ;
	wire _w91_ ;
	wire _w90_ ;
	wire _w89_ ;
	wire _w88_ ;
	wire _w87_ ;
	wire _w86_ ;
	wire _w85_ ;
	wire _w84_ ;
	wire _w83_ ;
	wire _w82_ ;
	wire _w81_ ;
	wire _w80_ ;
	wire _w79_ ;
	wire _w78_ ;
	wire _w77_ ;
	wire _w76_ ;
	wire _w75_ ;
	wire _w74_ ;
	wire _w73_ ;
	wire _w72_ ;
	wire _w71_ ;
	wire _w70_ ;
	wire _w69_ ;
	wire _w68_ ;
	wire _w67_ ;
	wire _w66_ ;
	wire _w65_ ;
	wire _w47_ ;
	wire _w46_ ;
	wire _w45_ ;
	wire _w44_ ;
	wire _w43_ ;
	wire _w42_ ;
	wire _w41_ ;
	wire _w40_ ;
	wire _w39_ ;
	wire _w38_ ;
	wire _w37_ ;
	wire _w48_ ;
	wire _w94_ ;
	wire _w35_ ;
	wire _w162_ ;
	wire _w64_ ;
	wire _w49_ ;
	wire _w50_ ;
	wire _w51_ ;
	wire _w52_ ;
	wire _w53_ ;
	wire _w54_ ;
	wire _w55_ ;
	wire _w56_ ;
	wire _w57_ ;
	wire _w58_ ;
	wire _w59_ ;
	wire _w60_ ;
	wire _w61_ ;
	wire _w62_ ;
	wire _w63_ ;
	wire _w95_ ;
	wire _w96_ ;
	wire _w97_ ;
	wire _w98_ ;
	wire _w99_ ;
	wire _w100_ ;
	wire _w101_ ;
	wire _w102_ ;
	wire _w103_ ;
	wire _w104_ ;
	wire _w105_ ;
	wire _w106_ ;
	wire _w107_ ;
	wire _w108_ ;
	wire _w109_ ;
	wire _w110_ ;
	wire _w111_ ;
	wire _w112_ ;
	wire _w113_ ;
	wire _w114_ ;
	wire _w115_ ;
	wire _w116_ ;
	wire _w117_ ;
	wire _w118_ ;
	wire _w119_ ;
	wire _w120_ ;
	wire _w121_ ;
	wire _w122_ ;
	wire _w123_ ;
	wire _w124_ ;
	wire _w125_ ;
	wire _w126_ ;
	wire _w127_ ;
	wire _w128_ ;
	wire _w129_ ;
	wire _w130_ ;
	wire _w131_ ;
	wire _w132_ ;
	wire _w133_ ;
	wire _w134_ ;
	wire _w135_ ;
	wire _w136_ ;
	wire _w137_ ;
	wire _w138_ ;
	wire _w139_ ;
	wire _w140_ ;
	wire _w141_ ;
	wire _w142_ ;
	wire _w143_ ;
	wire _w144_ ;
	wire _w145_ ;
	wire _w146_ ;
	wire _w147_ ;
	wire _w148_ ;
	wire _w149_ ;
	wire _w150_ ;
	wire _w151_ ;
	wire _w152_ ;
	wire _w153_ ;
	wire _w154_ ;
	wire _w155_ ;
	wire _w156_ ;
	wire _w157_ ;
	wire _w158_ ;
	wire _w159_ ;
	wire _w160_ ;
	wire _w161_ ;
	LUT1 #(
		.INIT('h1)
	) name0 (
		\stato_reg[0]/NET0131 ,
		_w35_
	);
	LUT3 #(
		.INIT('h10)
	) name1 (
		\fu4_reg/NET0131 ,
		\ru3_reg/NET0131 ,
		\ru4_reg/NET0131 ,
		_w37_
	);
	LUT3 #(
		.INIT('h8a)
	) name2 (
		\coda0_reg[2]/NET0131 ,
		\fu3_reg/NET0131 ,
		\ru3_reg/NET0131 ,
		_w38_
	);
	LUT4 #(
		.INIT('h070f)
	) name3 (
		\coda0_reg[2]/NET0131 ,
		\fu2_reg/NET0131 ,
		\ru1_reg/NET0131 ,
		\ru2_reg/NET0131 ,
		_w39_
	);
	LUT4 #(
		.INIT('hab00)
	) name4 (
		\ru2_reg/NET0131 ,
		_w37_,
		_w38_,
		_w39_,
		_w40_
	);
	LUT3 #(
		.INIT('h40)
	) name5 (
		\coda0_reg[2]/NET0131 ,
		\fu1_reg/NET0131 ,
		\ru1_reg/NET0131 ,
		_w41_
	);
	LUT2 #(
		.INIT('h2)
	) name6 (
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		_w42_
	);
	LUT2 #(
		.INIT('h4)
	) name7 (
		_w41_,
		_w42_,
		_w43_
	);
	LUT4 #(
		.INIT('h0001)
	) name8 (
		\fu1_reg/NET0131 ,
		\fu2_reg/NET0131 ,
		\fu3_reg/NET0131 ,
		\fu4_reg/NET0131 ,
		_w44_
	);
	LUT2 #(
		.INIT('h4)
	) name9 (
		\coda1_reg[2]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		_w45_
	);
	LUT2 #(
		.INIT('h2)
	) name10 (
		\coda0_reg[2]/NET0131 ,
		\stato_reg[0]/NET0131 ,
		_w46_
	);
	LUT2 #(
		.INIT('h4)
	) name11 (
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		_w47_
	);
	LUT4 #(
		.INIT('hb1b0)
	) name12 (
		_w44_,
		_w45_,
		_w46_,
		_w47_,
		_w48_
	);
	LUT3 #(
		.INIT('hf4)
	) name13 (
		_w40_,
		_w43_,
		_w48_,
		_w49_
	);
	LUT3 #(
		.INIT('h80)
	) name14 (
		\coda0_reg[0]/NET0131 ,
		\fu1_reg/NET0131 ,
		\ru1_reg/NET0131 ,
		_w50_
	);
	LUT3 #(
		.INIT('h70)
	) name15 (
		\coda0_reg[0]/NET0131 ,
		\fu1_reg/NET0131 ,
		\ru1_reg/NET0131 ,
		_w51_
	);
	LUT4 #(
		.INIT('h0100)
	) name16 (
		\fu4_reg/NET0131 ,
		\ru2_reg/NET0131 ,
		\ru3_reg/NET0131 ,
		\ru4_reg/NET0131 ,
		_w52_
	);
	LUT3 #(
		.INIT('h10)
	) name17 (
		\fu3_reg/NET0131 ,
		\ru2_reg/NET0131 ,
		\ru3_reg/NET0131 ,
		_w53_
	);
	LUT3 #(
		.INIT('h8a)
	) name18 (
		\coda0_reg[0]/NET0131 ,
		\fu2_reg/NET0131 ,
		\ru2_reg/NET0131 ,
		_w54_
	);
	LUT4 #(
		.INIT('h0001)
	) name19 (
		_w50_,
		_w52_,
		_w53_,
		_w54_,
		_w55_
	);
	LUT2 #(
		.INIT('h4)
	) name20 (
		\coda1_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		_w56_
	);
	LUT2 #(
		.INIT('h2)
	) name21 (
		\coda0_reg[0]/NET0131 ,
		\stato_reg[0]/NET0131 ,
		_w57_
	);
	LUT4 #(
		.INIT('haf04)
	) name22 (
		_w44_,
		_w47_,
		_w56_,
		_w57_,
		_w58_
	);
	LUT4 #(
		.INIT('hff02)
	) name23 (
		_w42_,
		_w51_,
		_w55_,
		_w58_,
		_w59_
	);
	LUT3 #(
		.INIT('h80)
	) name24 (
		\coda0_reg[1]/NET0131 ,
		\fu1_reg/NET0131 ,
		\ru1_reg/NET0131 ,
		_w60_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name25 (
		\coda0_reg[1]/NET0131 ,
		\fu2_reg/NET0131 ,
		\ru1_reg/NET0131 ,
		\ru2_reg/NET0131 ,
		_w61_
	);
	LUT4 #(
		.INIT('h3233)
	) name26 (
		\fu4_reg/NET0131 ,
		\ru2_reg/NET0131 ,
		\ru3_reg/NET0131 ,
		\ru4_reg/NET0131 ,
		_w62_
	);
	LUT3 #(
		.INIT('h8a)
	) name27 (
		\coda0_reg[1]/NET0131 ,
		\fu3_reg/NET0131 ,
		\ru3_reg/NET0131 ,
		_w63_
	);
	LUT4 #(
		.INIT('heeae)
	) name28 (
		_w60_,
		_w61_,
		_w62_,
		_w63_,
		_w64_
	);
	LUT2 #(
		.INIT('h4)
	) name29 (
		\coda1_reg[1]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		_w65_
	);
	LUT2 #(
		.INIT('h2)
	) name30 (
		\coda0_reg[1]/NET0131 ,
		\stato_reg[0]/NET0131 ,
		_w66_
	);
	LUT4 #(
		.INIT('haf04)
	) name31 (
		_w44_,
		_w47_,
		_w65_,
		_w66_,
		_w67_
	);
	LUT3 #(
		.INIT('hf8)
	) name32 (
		_w42_,
		_w64_,
		_w67_,
		_w68_
	);
	LUT3 #(
		.INIT('h04)
	) name33 (
		\ru1_reg/NET0131 ,
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		_w69_
	);
	LUT4 #(
		.INIT('hca00)
	) name34 (
		\coda0_reg[1]/NET0131 ,
		\coda1_reg[1]/NET0131 ,
		\fu2_reg/NET0131 ,
		\ru2_reg/NET0131 ,
		_w70_
	);
	LUT2 #(
		.INIT('h8)
	) name35 (
		_w69_,
		_w70_,
		_w71_
	);
	LUT4 #(
		.INIT('hca00)
	) name36 (
		\coda0_reg[1]/NET0131 ,
		\coda1_reg[1]/NET0131 ,
		\fu3_reg/NET0131 ,
		\ru3_reg/NET0131 ,
		_w72_
	);
	LUT4 #(
		.INIT('h080a)
	) name37 (
		\coda1_reg[1]/NET0131 ,
		\fu4_reg/NET0131 ,
		\ru3_reg/NET0131 ,
		\ru4_reg/NET0131 ,
		_w73_
	);
	LUT4 #(
		.INIT('h0200)
	) name38 (
		\coda0_reg[1]/NET0131 ,
		\fu4_reg/NET0131 ,
		\ru3_reg/NET0131 ,
		\ru4_reg/NET0131 ,
		_w74_
	);
	LUT4 #(
		.INIT('h0010)
	) name39 (
		\ru1_reg/NET0131 ,
		\ru2_reg/NET0131 ,
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		_w75_
	);
	LUT4 #(
		.INIT('hfe00)
	) name40 (
		_w72_,
		_w73_,
		_w74_,
		_w75_,
		_w76_
	);
	LUT4 #(
		.INIT('hff70)
	) name41 (
		\fu1_reg/NET0131 ,
		\ru1_reg/NET0131 ,
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		_w77_
	);
	LUT4 #(
		.INIT('h20aa)
	) name42 (
		\coda1_reg[1]/NET0131 ,
		\stato_reg[0]/NET0131 ,
		_w44_,
		_w77_,
		_w78_
	);
	LUT3 #(
		.INIT('h20)
	) name43 (
		\coda2_reg[1]/NET0131 ,
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		_w79_
	);
	LUT4 #(
		.INIT('h0040)
	) name44 (
		\fu1_reg/NET0131 ,
		\ru1_reg/NET0131 ,
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		_w80_
	);
	LUT4 #(
		.INIT('h45cf)
	) name45 (
		\coda0_reg[1]/NET0131 ,
		_w44_,
		_w79_,
		_w80_,
		_w81_
	);
	LUT4 #(
		.INIT('hfeff)
	) name46 (
		_w71_,
		_w76_,
		_w78_,
		_w81_,
		_w82_
	);
	LUT4 #(
		.INIT('hca00)
	) name47 (
		\coda1_reg[2]/NET0131 ,
		\coda2_reg[2]/NET0131 ,
		\fu2_reg/NET0131 ,
		\ru2_reg/NET0131 ,
		_w83_
	);
	LUT2 #(
		.INIT('h8)
	) name48 (
		_w69_,
		_w83_,
		_w84_
	);
	LUT4 #(
		.INIT('hca00)
	) name49 (
		\coda1_reg[2]/NET0131 ,
		\coda2_reg[2]/NET0131 ,
		\fu3_reg/NET0131 ,
		\ru3_reg/NET0131 ,
		_w85_
	);
	LUT4 #(
		.INIT('h080a)
	) name50 (
		\coda2_reg[2]/NET0131 ,
		\fu4_reg/NET0131 ,
		\ru3_reg/NET0131 ,
		\ru4_reg/NET0131 ,
		_w86_
	);
	LUT4 #(
		.INIT('h0200)
	) name51 (
		\coda1_reg[2]/NET0131 ,
		\fu4_reg/NET0131 ,
		\ru3_reg/NET0131 ,
		\ru4_reg/NET0131 ,
		_w87_
	);
	LUT4 #(
		.INIT('haaa8)
	) name52 (
		_w75_,
		_w85_,
		_w86_,
		_w87_,
		_w88_
	);
	LUT4 #(
		.INIT('h20aa)
	) name53 (
		\coda2_reg[2]/NET0131 ,
		\stato_reg[0]/NET0131 ,
		_w44_,
		_w77_,
		_w89_
	);
	LUT3 #(
		.INIT('h20)
	) name54 (
		\coda3_reg[2]/NET0131 ,
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		_w90_
	);
	LUT4 #(
		.INIT('h4c5f)
	) name55 (
		\coda1_reg[2]/NET0131 ,
		_w44_,
		_w80_,
		_w90_,
		_w91_
	);
	LUT4 #(
		.INIT('hfeff)
	) name56 (
		_w84_,
		_w88_,
		_w89_,
		_w91_,
		_w92_
	);
	LUT4 #(
		.INIT('hca00)
	) name57 (
		\coda0_reg[2]/NET0131 ,
		\coda1_reg[2]/NET0131 ,
		\fu2_reg/NET0131 ,
		\ru2_reg/NET0131 ,
		_w93_
	);
	LUT2 #(
		.INIT('h8)
	) name58 (
		_w69_,
		_w93_,
		_w94_
	);
	LUT4 #(
		.INIT('hca00)
	) name59 (
		\coda0_reg[2]/NET0131 ,
		\coda1_reg[2]/NET0131 ,
		\fu3_reg/NET0131 ,
		\ru3_reg/NET0131 ,
		_w95_
	);
	LUT4 #(
		.INIT('h080a)
	) name60 (
		\coda1_reg[2]/NET0131 ,
		\fu4_reg/NET0131 ,
		\ru3_reg/NET0131 ,
		\ru4_reg/NET0131 ,
		_w96_
	);
	LUT4 #(
		.INIT('h0200)
	) name61 (
		\coda0_reg[2]/NET0131 ,
		\fu4_reg/NET0131 ,
		\ru3_reg/NET0131 ,
		\ru4_reg/NET0131 ,
		_w97_
	);
	LUT4 #(
		.INIT('haaa8)
	) name62 (
		_w75_,
		_w95_,
		_w96_,
		_w97_,
		_w98_
	);
	LUT4 #(
		.INIT('h20aa)
	) name63 (
		\coda1_reg[2]/NET0131 ,
		\stato_reg[0]/NET0131 ,
		_w44_,
		_w77_,
		_w99_
	);
	LUT3 #(
		.INIT('h20)
	) name64 (
		\coda2_reg[2]/NET0131 ,
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		_w100_
	);
	LUT4 #(
		.INIT('h4c5f)
	) name65 (
		\coda0_reg[2]/NET0131 ,
		_w44_,
		_w80_,
		_w100_,
		_w101_
	);
	LUT4 #(
		.INIT('hfeff)
	) name66 (
		_w94_,
		_w98_,
		_w99_,
		_w101_,
		_w102_
	);
	LUT4 #(
		.INIT('hca00)
	) name67 (
		\coda0_reg[0]/NET0131 ,
		\coda1_reg[0]/NET0131 ,
		\fu2_reg/NET0131 ,
		\ru2_reg/NET0131 ,
		_w103_
	);
	LUT2 #(
		.INIT('h8)
	) name68 (
		_w69_,
		_w103_,
		_w104_
	);
	LUT4 #(
		.INIT('hca00)
	) name69 (
		\coda0_reg[0]/NET0131 ,
		\coda1_reg[0]/NET0131 ,
		\fu3_reg/NET0131 ,
		\ru3_reg/NET0131 ,
		_w105_
	);
	LUT4 #(
		.INIT('h080a)
	) name70 (
		\coda1_reg[0]/NET0131 ,
		\fu4_reg/NET0131 ,
		\ru3_reg/NET0131 ,
		\ru4_reg/NET0131 ,
		_w106_
	);
	LUT4 #(
		.INIT('h0200)
	) name71 (
		\coda0_reg[0]/NET0131 ,
		\fu4_reg/NET0131 ,
		\ru3_reg/NET0131 ,
		\ru4_reg/NET0131 ,
		_w107_
	);
	LUT4 #(
		.INIT('haaa8)
	) name72 (
		_w75_,
		_w105_,
		_w106_,
		_w107_,
		_w108_
	);
	LUT4 #(
		.INIT('h20aa)
	) name73 (
		\coda1_reg[0]/NET0131 ,
		\stato_reg[0]/NET0131 ,
		_w44_,
		_w77_,
		_w109_
	);
	LUT3 #(
		.INIT('h20)
	) name74 (
		\coda2_reg[0]/NET0131 ,
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		_w110_
	);
	LUT4 #(
		.INIT('h4c5f)
	) name75 (
		\coda0_reg[0]/NET0131 ,
		_w44_,
		_w80_,
		_w110_,
		_w111_
	);
	LUT4 #(
		.INIT('hfeff)
	) name76 (
		_w104_,
		_w108_,
		_w109_,
		_w111_,
		_w112_
	);
	LUT4 #(
		.INIT('hca00)
	) name77 (
		\coda1_reg[0]/NET0131 ,
		\coda2_reg[0]/NET0131 ,
		\fu2_reg/NET0131 ,
		\ru2_reg/NET0131 ,
		_w113_
	);
	LUT2 #(
		.INIT('h8)
	) name78 (
		_w69_,
		_w113_,
		_w114_
	);
	LUT4 #(
		.INIT('hca00)
	) name79 (
		\coda1_reg[0]/NET0131 ,
		\coda2_reg[0]/NET0131 ,
		\fu3_reg/NET0131 ,
		\ru3_reg/NET0131 ,
		_w115_
	);
	LUT4 #(
		.INIT('h080a)
	) name80 (
		\coda2_reg[0]/NET0131 ,
		\fu4_reg/NET0131 ,
		\ru3_reg/NET0131 ,
		\ru4_reg/NET0131 ,
		_w116_
	);
	LUT4 #(
		.INIT('h0200)
	) name81 (
		\coda1_reg[0]/NET0131 ,
		\fu4_reg/NET0131 ,
		\ru3_reg/NET0131 ,
		\ru4_reg/NET0131 ,
		_w117_
	);
	LUT4 #(
		.INIT('haaa8)
	) name82 (
		_w75_,
		_w115_,
		_w116_,
		_w117_,
		_w118_
	);
	LUT4 #(
		.INIT('h20aa)
	) name83 (
		\coda2_reg[0]/NET0131 ,
		\stato_reg[0]/NET0131 ,
		_w44_,
		_w77_,
		_w119_
	);
	LUT3 #(
		.INIT('h20)
	) name84 (
		\coda3_reg[0]/NET0131 ,
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		_w120_
	);
	LUT4 #(
		.INIT('h4c5f)
	) name85 (
		\coda1_reg[0]/NET0131 ,
		_w44_,
		_w80_,
		_w120_,
		_w121_
	);
	LUT4 #(
		.INIT('hfeff)
	) name86 (
		_w114_,
		_w118_,
		_w119_,
		_w121_,
		_w122_
	);
	LUT4 #(
		.INIT('hca00)
	) name87 (
		\coda1_reg[1]/NET0131 ,
		\coda2_reg[1]/NET0131 ,
		\fu2_reg/NET0131 ,
		\ru2_reg/NET0131 ,
		_w123_
	);
	LUT2 #(
		.INIT('h8)
	) name88 (
		_w69_,
		_w123_,
		_w124_
	);
	LUT4 #(
		.INIT('hca00)
	) name89 (
		\coda1_reg[1]/NET0131 ,
		\coda2_reg[1]/NET0131 ,
		\fu3_reg/NET0131 ,
		\ru3_reg/NET0131 ,
		_w125_
	);
	LUT4 #(
		.INIT('h080a)
	) name90 (
		\coda2_reg[1]/NET0131 ,
		\fu4_reg/NET0131 ,
		\ru3_reg/NET0131 ,
		\ru4_reg/NET0131 ,
		_w126_
	);
	LUT4 #(
		.INIT('h0200)
	) name91 (
		\coda1_reg[1]/NET0131 ,
		\fu4_reg/NET0131 ,
		\ru3_reg/NET0131 ,
		\ru4_reg/NET0131 ,
		_w127_
	);
	LUT4 #(
		.INIT('haaa8)
	) name92 (
		_w75_,
		_w125_,
		_w126_,
		_w127_,
		_w128_
	);
	LUT3 #(
		.INIT('h08)
	) name93 (
		\ru1_reg/NET0131 ,
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		_w129_
	);
	LUT3 #(
		.INIT('hca)
	) name94 (
		\coda1_reg[1]/NET0131 ,
		\coda2_reg[1]/NET0131 ,
		\fu1_reg/NET0131 ,
		_w130_
	);
	LUT2 #(
		.INIT('h8)
	) name95 (
		_w129_,
		_w130_,
		_w131_
	);
	LUT2 #(
		.INIT('h4)
	) name96 (
		\coda3_reg[1]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		_w132_
	);
	LUT2 #(
		.INIT('h2)
	) name97 (
		\coda2_reg[1]/NET0131 ,
		\stato_reg[0]/NET0131 ,
		_w133_
	);
	LUT4 #(
		.INIT('haf04)
	) name98 (
		_w44_,
		_w47_,
		_w132_,
		_w133_,
		_w134_
	);
	LUT4 #(
		.INIT('hfffe)
	) name99 (
		_w124_,
		_w128_,
		_w131_,
		_w134_,
		_w135_
	);
	LUT2 #(
		.INIT('h4)
	) name100 (
		\coda3_reg[0]/NET0131 ,
		\fu2_reg/NET0131 ,
		_w136_
	);
	LUT4 #(
		.INIT('h0e00)
	) name101 (
		\coda2_reg[0]/NET0131 ,
		\fu2_reg/NET0131 ,
		\ru1_reg/NET0131 ,
		\ru2_reg/NET0131 ,
		_w137_
	);
	LUT3 #(
		.INIT('h20)
	) name102 (
		_w42_,
		_w136_,
		_w137_,
		_w138_
	);
	LUT4 #(
		.INIT('hca00)
	) name103 (
		\coda2_reg[0]/NET0131 ,
		\coda3_reg[0]/NET0131 ,
		\fu3_reg/NET0131 ,
		\ru3_reg/NET0131 ,
		_w139_
	);
	LUT4 #(
		.INIT('h080a)
	) name104 (
		\coda3_reg[0]/NET0131 ,
		\fu4_reg/NET0131 ,
		\ru3_reg/NET0131 ,
		\ru4_reg/NET0131 ,
		_w140_
	);
	LUT4 #(
		.INIT('h0200)
	) name105 (
		\coda2_reg[0]/NET0131 ,
		\fu4_reg/NET0131 ,
		\ru3_reg/NET0131 ,
		\ru4_reg/NET0131 ,
		_w141_
	);
	LUT4 #(
		.INIT('hfe00)
	) name106 (
		_w139_,
		_w140_,
		_w141_,
		_w75_,
		_w142_
	);
	LUT4 #(
		.INIT('h20aa)
	) name107 (
		\coda3_reg[0]/NET0131 ,
		\stato_reg[0]/NET0131 ,
		_w44_,
		_w77_,
		_w143_
	);
	LUT2 #(
		.INIT('h8)
	) name108 (
		\coda2_reg[0]/NET0131 ,
		_w80_,
		_w144_
	);
	LUT4 #(
		.INIT('hfffe)
	) name109 (
		_w138_,
		_w142_,
		_w143_,
		_w144_,
		_w145_
	);
	LUT2 #(
		.INIT('h4)
	) name110 (
		\coda3_reg[1]/NET0131 ,
		\fu2_reg/NET0131 ,
		_w146_
	);
	LUT4 #(
		.INIT('h0e00)
	) name111 (
		\coda2_reg[1]/NET0131 ,
		\fu2_reg/NET0131 ,
		\ru1_reg/NET0131 ,
		\ru2_reg/NET0131 ,
		_w147_
	);
	LUT3 #(
		.INIT('h20)
	) name112 (
		_w42_,
		_w146_,
		_w147_,
		_w148_
	);
	LUT4 #(
		.INIT('hca00)
	) name113 (
		\coda2_reg[1]/NET0131 ,
		\coda3_reg[1]/NET0131 ,
		\fu3_reg/NET0131 ,
		\ru3_reg/NET0131 ,
		_w149_
	);
	LUT4 #(
		.INIT('h080a)
	) name114 (
		\coda3_reg[1]/NET0131 ,
		\fu4_reg/NET0131 ,
		\ru3_reg/NET0131 ,
		\ru4_reg/NET0131 ,
		_w150_
	);
	LUT4 #(
		.INIT('h0200)
	) name115 (
		\coda2_reg[1]/NET0131 ,
		\fu4_reg/NET0131 ,
		\ru3_reg/NET0131 ,
		\ru4_reg/NET0131 ,
		_w151_
	);
	LUT4 #(
		.INIT('haaa8)
	) name116 (
		_w75_,
		_w149_,
		_w150_,
		_w151_,
		_w152_
	);
	LUT2 #(
		.INIT('h8)
	) name117 (
		\coda2_reg[1]/NET0131 ,
		_w80_,
		_w153_
	);
	LUT4 #(
		.INIT('h20aa)
	) name118 (
		\coda3_reg[1]/NET0131 ,
		\stato_reg[0]/NET0131 ,
		_w44_,
		_w77_,
		_w154_
	);
	LUT4 #(
		.INIT('hfffe)
	) name119 (
		_w148_,
		_w152_,
		_w153_,
		_w154_,
		_w155_
	);
	LUT2 #(
		.INIT('h4)
	) name120 (
		\coda3_reg[2]/NET0131 ,
		\fu2_reg/NET0131 ,
		_w156_
	);
	LUT4 #(
		.INIT('h0e00)
	) name121 (
		\coda2_reg[2]/NET0131 ,
		\fu2_reg/NET0131 ,
		\ru1_reg/NET0131 ,
		\ru2_reg/NET0131 ,
		_w157_
	);
	LUT3 #(
		.INIT('h20)
	) name122 (
		_w42_,
		_w156_,
		_w157_,
		_w158_
	);
	LUT4 #(
		.INIT('hca00)
	) name123 (
		\coda2_reg[2]/NET0131 ,
		\coda3_reg[2]/NET0131 ,
		\fu3_reg/NET0131 ,
		\ru3_reg/NET0131 ,
		_w159_
	);
	LUT4 #(
		.INIT('h080a)
	) name124 (
		\coda3_reg[2]/NET0131 ,
		\fu4_reg/NET0131 ,
		\ru3_reg/NET0131 ,
		\ru4_reg/NET0131 ,
		_w160_
	);
	LUT4 #(
		.INIT('h0200)
	) name125 (
		\coda2_reg[2]/NET0131 ,
		\fu4_reg/NET0131 ,
		\ru3_reg/NET0131 ,
		\ru4_reg/NET0131 ,
		_w161_
	);
	LUT4 #(
		.INIT('haaa8)
	) name126 (
		_w75_,
		_w159_,
		_w160_,
		_w161_,
		_w162_
	);
	LUT2 #(
		.INIT('h8)
	) name127 (
		\coda2_reg[2]/NET0131 ,
		_w80_,
		_w163_
	);
	LUT4 #(
		.INIT('h20aa)
	) name128 (
		\coda3_reg[2]/NET0131 ,
		\stato_reg[0]/NET0131 ,
		_w44_,
		_w77_,
		_w164_
	);
	LUT4 #(
		.INIT('hfffe)
	) name129 (
		_w158_,
		_w162_,
		_w163_,
		_w164_,
		_w165_
	);
	LUT2 #(
		.INIT('h2)
	) name130 (
		\grant_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		_w166_
	);
	LUT2 #(
		.INIT('h2)
	) name131 (
		\grant_reg[0]/NET0131 ,
		\stato_reg[0]/NET0131 ,
		_w167_
	);
	LUT3 #(
		.INIT('h13)
	) name132 (
		_w44_,
		_w166_,
		_w167_,
		_w168_
	);
	LUT3 #(
		.INIT('h20)
	) name133 (
		\coda0_reg[1]/NET0131 ,
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		_w169_
	);
	LUT2 #(
		.INIT('h8)
	) name134 (
		\coda0_reg[0]/NET0131 ,
		\coda0_reg[2]/NET0131 ,
		_w170_
	);
	LUT3 #(
		.INIT('h40)
	) name135 (
		_w44_,
		_w169_,
		_w170_,
		_w171_
	);
	LUT2 #(
		.INIT('hd)
	) name136 (
		_w168_,
		_w171_,
		_w172_
	);
	LUT2 #(
		.INIT('h2)
	) name137 (
		\grant_reg[1]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		_w173_
	);
	LUT2 #(
		.INIT('h2)
	) name138 (
		\grant_reg[1]/NET0131 ,
		\stato_reg[0]/NET0131 ,
		_w174_
	);
	LUT3 #(
		.INIT('h13)
	) name139 (
		_w44_,
		_w173_,
		_w174_,
		_w175_
	);
	LUT3 #(
		.INIT('h10)
	) name140 (
		\coda0_reg[1]/NET0131 ,
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		_w176_
	);
	LUT2 #(
		.INIT('h2)
	) name141 (
		\coda0_reg[0]/NET0131 ,
		\coda0_reg[2]/NET0131 ,
		_w177_
	);
	LUT3 #(
		.INIT('h40)
	) name142 (
		_w44_,
		_w176_,
		_w177_,
		_w178_
	);
	LUT2 #(
		.INIT('hd)
	) name143 (
		_w175_,
		_w178_,
		_w179_
	);
	LUT2 #(
		.INIT('h2)
	) name144 (
		\grant_reg[2]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		_w180_
	);
	LUT2 #(
		.INIT('h2)
	) name145 (
		\grant_reg[2]/NET0131 ,
		\stato_reg[0]/NET0131 ,
		_w181_
	);
	LUT3 #(
		.INIT('h13)
	) name146 (
		_w44_,
		_w180_,
		_w181_,
		_w182_
	);
	LUT2 #(
		.INIT('h1)
	) name147 (
		\coda0_reg[0]/NET0131 ,
		\coda0_reg[2]/NET0131 ,
		_w183_
	);
	LUT3 #(
		.INIT('h40)
	) name148 (
		_w44_,
		_w169_,
		_w183_,
		_w184_
	);
	LUT2 #(
		.INIT('hd)
	) name149 (
		_w182_,
		_w184_,
		_w185_
	);
	LUT2 #(
		.INIT('h2)
	) name150 (
		\grant_reg[3]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		_w186_
	);
	LUT2 #(
		.INIT('h2)
	) name151 (
		\grant_reg[3]/NET0131 ,
		\stato_reg[0]/NET0131 ,
		_w187_
	);
	LUT3 #(
		.INIT('h13)
	) name152 (
		_w44_,
		_w186_,
		_w187_,
		_w188_
	);
	LUT2 #(
		.INIT('h4)
	) name153 (
		\coda0_reg[0]/NET0131 ,
		\coda0_reg[2]/NET0131 ,
		_w189_
	);
	LUT3 #(
		.INIT('h40)
	) name154 (
		_w44_,
		_w176_,
		_w189_,
		_w190_
	);
	LUT2 #(
		.INIT('hd)
	) name155 (
		_w188_,
		_w190_,
		_w191_
	);
	LUT4 #(
		.INIT('h0aca)
	) name156 (
		\fu1_reg/NET0131 ,
		\ru1_reg/NET0131 ,
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		_w192_
	);
	LUT4 #(
		.INIT('h0aca)
	) name157 (
		\fu2_reg/NET0131 ,
		\ru2_reg/NET0131 ,
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		_w193_
	);
	LUT4 #(
		.INIT('h0aca)
	) name158 (
		\fu3_reg/NET0131 ,
		\ru3_reg/NET0131 ,
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		_w194_
	);
	LUT4 #(
		.INIT('h0aca)
	) name159 (
		\fu4_reg/NET0131 ,
		\ru4_reg/NET0131 ,
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		_w195_
	);
	LUT4 #(
		.INIT('h0aca)
	) name160 (
		\grant_o[0]_pad ,
		\grant_reg[0]/NET0131 ,
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		_w196_
	);
	LUT4 #(
		.INIT('h0aca)
	) name161 (
		\grant_o[1]_pad ,
		\grant_reg[1]/NET0131 ,
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		_w197_
	);
	LUT4 #(
		.INIT('h0aca)
	) name162 (
		\grant_o[2]_pad ,
		\grant_reg[2]/NET0131 ,
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		_w198_
	);
	LUT4 #(
		.INIT('h0aca)
	) name163 (
		\grant_o[3]_pad ,
		\grant_reg[3]/NET0131 ,
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		_w199_
	);
	LUT4 #(
		.INIT('h0aca)
	) name164 (
		\request1_pad ,
		\ru1_reg/NET0131 ,
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		_w200_
	);
	LUT4 #(
		.INIT('h0aca)
	) name165 (
		\request2_pad ,
		\ru2_reg/NET0131 ,
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		_w201_
	);
	LUT4 #(
		.INIT('h0aca)
	) name166 (
		\request3_pad ,
		\ru3_reg/NET0131 ,
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		_w202_
	);
	LUT4 #(
		.INIT('h0aca)
	) name167 (
		\request4_pad ,
		\ru4_reg/NET0131 ,
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		_w203_
	);
	assign \_al_n0  = 1'b0;
	assign \_al_n1  = 1'b1;
	assign \g1143/_0_  = _w49_ ;
	assign \g1144/_0_  = _w59_ ;
	assign \g1145/_0_  = _w68_ ;
	assign \g1146/_0_  = _w82_ ;
	assign \g1147/_0_  = _w92_ ;
	assign \g1148/_0_  = _w102_ ;
	assign \g1149/_0_  = _w112_ ;
	assign \g1150/_0_  = _w122_ ;
	assign \g1151/_0_  = _w135_ ;
	assign \g1152/_0_  = _w145_ ;
	assign \g1153/_0_  = _w155_ ;
	assign \g1154/_0_  = _w165_ ;
	assign \g1174/_0_  = _w172_ ;
	assign \g1175/_0_  = _w179_ ;
	assign \g1176/_0_  = _w185_ ;
	assign \g1177/_0_  = _w191_ ;
	assign \g1238/_0_  = _w192_ ;
	assign \g1239/_0_  = _w193_ ;
	assign \g1240/_0_  = _w194_ ;
	assign \g1241/_0_  = _w195_ ;
	assign \g1242/_0_  = _w196_ ;
	assign \g1243/_0_  = _w197_ ;
	assign \g1244/_0_  = _w198_ ;
	assign \g1245/_0_  = _w199_ ;
	assign \g1247/_0_  = _w200_ ;
	assign \g1248/_0_  = _w201_ ;
	assign \g1249/_0_  = _w202_ ;
	assign \g1250/_0_  = _w203_ ;
	assign \g1520/_0_  = _w35_ ;
endmodule;