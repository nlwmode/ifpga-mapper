module top (\a0_pad , a_pad, \b0_pad , b_pad, \c0_pad , c_pad, \d0_pad , d_pad, \e0_pad , e_pad, \f0_pad , f_pad, \g0_pad , g_pad, h_pad, i_pad, j_pad, k_pad, l_pad, m_pad, n_pad, o_pad, p_pad, q_pad, r_pad, s_pad, t_pad, u_pad, v_pad, w_pad, x_pad, y_pad, z_pad, \h0_pad , \i0_pad , \j0_pad , \k0_pad , \l0_pad , \m0_pad , \n0_pad , \o0_pad , \p0_pad , \q0_pad , \r0_pad , \s0_pad , \t0_pad , \u0_pad , \v0_pad , \w0_pad , \x0_pad );
	input \a0_pad  ;
	input a_pad ;
	input \b0_pad  ;
	input b_pad ;
	input \c0_pad  ;
	input c_pad ;
	input \d0_pad  ;
	input d_pad ;
	input \e0_pad  ;
	input e_pad ;
	input \f0_pad  ;
	input f_pad ;
	input \g0_pad  ;
	input g_pad ;
	input h_pad ;
	input i_pad ;
	input j_pad ;
	input k_pad ;
	input l_pad ;
	input m_pad ;
	input n_pad ;
	input o_pad ;
	input p_pad ;
	input q_pad ;
	input r_pad ;
	input s_pad ;
	input t_pad ;
	input u_pad ;
	input v_pad ;
	input w_pad ;
	input x_pad ;
	input y_pad ;
	input z_pad ;
	output \h0_pad  ;
	output \i0_pad  ;
	output \j0_pad  ;
	output \k0_pad  ;
	output \l0_pad  ;
	output \m0_pad  ;
	output \n0_pad  ;
	output \o0_pad  ;
	output \p0_pad  ;
	output \q0_pad  ;
	output \r0_pad  ;
	output \s0_pad  ;
	output \t0_pad  ;
	output \u0_pad  ;
	output \v0_pad  ;
	output \w0_pad  ;
	output \x0_pad  ;
	wire _w136_ ;
	wire _w135_ ;
	wire _w134_ ;
	wire _w133_ ;
	wire _w132_ ;
	wire _w131_ ;
	wire _w130_ ;
	wire _w129_ ;
	wire _w128_ ;
	wire _w127_ ;
	wire _w126_ ;
	wire _w125_ ;
	wire _w124_ ;
	wire _w123_ ;
	wire _w122_ ;
	wire _w121_ ;
	wire _w120_ ;
	wire _w119_ ;
	wire _w118_ ;
	wire _w117_ ;
	wire _w116_ ;
	wire _w115_ ;
	wire _w114_ ;
	wire _w113_ ;
	wire _w112_ ;
	wire _w111_ ;
	wire _w110_ ;
	wire _w109_ ;
	wire _w108_ ;
	wire _w107_ ;
	wire _w106_ ;
	wire _w105_ ;
	wire _w104_ ;
	wire _w103_ ;
	wire _w102_ ;
	wire _w101_ ;
	wire _w100_ ;
	wire _w99_ ;
	wire _w98_ ;
	wire _w97_ ;
	wire _w96_ ;
	wire _w95_ ;
	wire _w94_ ;
	wire _w63_ ;
	wire _w62_ ;
	wire _w61_ ;
	wire _w60_ ;
	wire _w59_ ;
	wire _w58_ ;
	wire _w57_ ;
	wire _w56_ ;
	wire _w55_ ;
	wire _w54_ ;
	wire _w53_ ;
	wire _w52_ ;
	wire _w51_ ;
	wire _w50_ ;
	wire _w49_ ;
	wire _w48_ ;
	wire _w35_ ;
	wire _w36_ ;
	wire _w37_ ;
	wire _w38_ ;
	wire _w39_ ;
	wire _w40_ ;
	wire _w41_ ;
	wire _w42_ ;
	wire _w43_ ;
	wire _w44_ ;
	wire _w45_ ;
	wire _w46_ ;
	wire _w47_ ;
	wire _w64_ ;
	wire _w65_ ;
	wire _w66_ ;
	wire _w67_ ;
	wire _w68_ ;
	wire _w69_ ;
	wire _w70_ ;
	wire _w71_ ;
	wire _w72_ ;
	wire _w73_ ;
	wire _w74_ ;
	wire _w75_ ;
	wire _w76_ ;
	wire _w77_ ;
	wire _w78_ ;
	wire _w79_ ;
	wire _w80_ ;
	wire _w81_ ;
	wire _w82_ ;
	wire _w83_ ;
	wire _w84_ ;
	wire _w85_ ;
	wire _w86_ ;
	wire _w87_ ;
	wire _w88_ ;
	wire _w89_ ;
	wire _w90_ ;
	wire _w91_ ;
	wire _w92_ ;
	wire _w93_ ;
	LUT2 #(
		.INIT('h1)
	) name0 (
		c_pad,
		s_pad,
		_w35_
	);
	LUT2 #(
		.INIT('h8)
	) name1 (
		d_pad,
		t_pad,
		_w36_
	);
	LUT4 #(
		.INIT('he8a0)
	) name2 (
		c_pad,
		d_pad,
		s_pad,
		t_pad,
		_w37_
	);
	LUT2 #(
		.INIT('h8)
	) name3 (
		e_pad,
		u_pad,
		_w38_
	);
	LUT2 #(
		.INIT('h1)
	) name4 (
		f_pad,
		v_pad,
		_w39_
	);
	LUT4 #(
		.INIT('h0013)
	) name5 (
		e_pad,
		f_pad,
		u_pad,
		v_pad,
		_w40_
	);
	LUT4 #(
		.INIT('hfac8)
	) name6 (
		g_pad,
		h_pad,
		w_pad,
		x_pad,
		_w41_
	);
	LUT2 #(
		.INIT('h8)
	) name7 (
		h_pad,
		x_pad,
		_w42_
	);
	LUT4 #(
		.INIT('hc800)
	) name8 (
		g_pad,
		h_pad,
		w_pad,
		x_pad,
		_w43_
	);
	LUT4 #(
		.INIT('hfac8)
	) name9 (
		\c0_pad ,
		\d0_pad ,
		m_pad,
		n_pad,
		_w44_
	);
	LUT2 #(
		.INIT('h8)
	) name10 (
		\d0_pad ,
		n_pad,
		_w45_
	);
	LUT4 #(
		.INIT('hc800)
	) name11 (
		\c0_pad ,
		\d0_pad ,
		m_pad,
		n_pad,
		_w46_
	);
	LUT3 #(
		.INIT('hc8)
	) name12 (
		\f0_pad ,
		\g0_pad ,
		p_pad,
		_w47_
	);
	LUT4 #(
		.INIT('h135f)
	) name13 (
		\e0_pad ,
		\f0_pad ,
		o_pad,
		p_pad,
		_w48_
	);
	LUT2 #(
		.INIT('h1)
	) name14 (
		\e0_pad ,
		o_pad,
		_w49_
	);
	LUT4 #(
		.INIT('h008a)
	) name15 (
		_w44_,
		_w47_,
		_w48_,
		_w49_,
		_w50_
	);
	LUT2 #(
		.INIT('h8)
	) name16 (
		\c0_pad ,
		m_pad,
		_w51_
	);
	LUT4 #(
		.INIT('h135f)
	) name17 (
		\b0_pad ,
		\c0_pad ,
		l_pad,
		m_pad,
		_w52_
	);
	LUT2 #(
		.INIT('h1)
	) name18 (
		\b0_pad ,
		l_pad,
		_w53_
	);
	LUT4 #(
		.INIT('hfac8)
	) name19 (
		\a0_pad ,
		j_pad,
		k_pad,
		z_pad,
		_w54_
	);
	LUT2 #(
		.INIT('h4)
	) name20 (
		_w53_,
		_w54_,
		_w55_
	);
	LUT4 #(
		.INIT('hef00)
	) name21 (
		_w46_,
		_w50_,
		_w52_,
		_w55_,
		_w56_
	);
	LUT2 #(
		.INIT('h8)
	) name22 (
		\a0_pad ,
		k_pad,
		_w57_
	);
	LUT4 #(
		.INIT('ha080)
	) name23 (
		\a0_pad ,
		j_pad,
		k_pad,
		z_pad,
		_w58_
	);
	LUT4 #(
		.INIT('h135f)
	) name24 (
		i_pad,
		j_pad,
		y_pad,
		z_pad,
		_w59_
	);
	LUT2 #(
		.INIT('h4)
	) name25 (
		_w58_,
		_w59_,
		_w60_
	);
	LUT2 #(
		.INIT('h1)
	) name26 (
		i_pad,
		y_pad,
		_w61_
	);
	LUT2 #(
		.INIT('h2)
	) name27 (
		_w41_,
		_w61_,
		_w62_
	);
	LUT4 #(
		.INIT('h1055)
	) name28 (
		_w43_,
		_w56_,
		_w60_,
		_w62_,
		_w63_
	);
	LUT2 #(
		.INIT('h8)
	) name29 (
		g_pad,
		w_pad,
		_w64_
	);
	LUT4 #(
		.INIT('h135f)
	) name30 (
		f_pad,
		g_pad,
		v_pad,
		w_pad,
		_w65_
	);
	LUT2 #(
		.INIT('h4)
	) name31 (
		_w38_,
		_w65_,
		_w66_
	);
	LUT4 #(
		.INIT('hfac8)
	) name32 (
		d_pad,
		e_pad,
		t_pad,
		u_pad,
		_w67_
	);
	LUT2 #(
		.INIT('h4)
	) name33 (
		_w35_,
		_w67_,
		_w68_
	);
	LUT4 #(
		.INIT('h1500)
	) name34 (
		_w40_,
		_w63_,
		_w66_,
		_w68_,
		_w69_
	);
	LUT2 #(
		.INIT('h1)
	) name35 (
		b_pad,
		r_pad,
		_w70_
	);
	LUT4 #(
		.INIT('h21a5)
	) name36 (
		a_pad,
		b_pad,
		q_pad,
		r_pad,
		_w71_
	);
	LUT4 #(
		.INIT('hf100)
	) name37 (
		_w37_,
		_w69_,
		_w70_,
		_w71_,
		_w72_
	);
	LUT4 #(
		.INIT('h5a48)
	) name38 (
		a_pad,
		b_pad,
		q_pad,
		r_pad,
		_w73_
	);
	LUT4 #(
		.INIT('h4800)
	) name39 (
		a_pad,
		b_pad,
		q_pad,
		r_pad,
		_w74_
	);
	LUT4 #(
		.INIT('h001f)
	) name40 (
		_w37_,
		_w69_,
		_w73_,
		_w74_,
		_w75_
	);
	LUT2 #(
		.INIT('h4)
	) name41 (
		_w72_,
		_w75_,
		_w76_
	);
	LUT2 #(
		.INIT('h6)
	) name42 (
		b_pad,
		r_pad,
		_w77_
	);
	LUT3 #(
		.INIT('h1e)
	) name43 (
		_w37_,
		_w69_,
		_w77_,
		_w78_
	);
	LUT2 #(
		.INIT('h6)
	) name44 (
		c_pad,
		s_pad,
		_w79_
	);
	LUT2 #(
		.INIT('h2)
	) name45 (
		_w67_,
		_w79_,
		_w80_
	);
	LUT4 #(
		.INIT('h1500)
	) name46 (
		_w40_,
		_w63_,
		_w66_,
		_w80_,
		_w81_
	);
	LUT4 #(
		.INIT('h1500)
	) name47 (
		_w40_,
		_w63_,
		_w66_,
		_w67_,
		_w82_
	);
	LUT4 #(
		.INIT('hf2f6)
	) name48 (
		_w36_,
		_w79_,
		_w81_,
		_w82_,
		_w83_
	);
	LUT4 #(
		.INIT('h5a48)
	) name49 (
		d_pad,
		e_pad,
		t_pad,
		u_pad,
		_w84_
	);
	LUT4 #(
		.INIT('h1500)
	) name50 (
		_w40_,
		_w63_,
		_w66_,
		_w84_,
		_w85_
	);
	LUT4 #(
		.INIT('hfac8)
	) name51 (
		e_pad,
		f_pad,
		u_pad,
		v_pad,
		_w86_
	);
	LUT4 #(
		.INIT('h21a5)
	) name52 (
		d_pad,
		e_pad,
		t_pad,
		u_pad,
		_w87_
	);
	LUT4 #(
		.INIT('h8f00)
	) name53 (
		_w63_,
		_w65_,
		_w86_,
		_w87_,
		_w88_
	);
	LUT2 #(
		.INIT('h1)
	) name54 (
		_w85_,
		_w88_,
		_w89_
	);
	LUT2 #(
		.INIT('h6)
	) name55 (
		e_pad,
		u_pad,
		_w90_
	);
	LUT4 #(
		.INIT('hea15)
	) name56 (
		_w39_,
		_w63_,
		_w65_,
		_w90_,
		_w91_
	);
	LUT2 #(
		.INIT('h6)
	) name57 (
		f_pad,
		v_pad,
		_w92_
	);
	LUT3 #(
		.INIT('h2d)
	) name58 (
		_w63_,
		_w64_,
		_w92_,
		_w93_
	);
	LUT4 #(
		.INIT('h5510)
	) name59 (
		_w42_,
		_w56_,
		_w60_,
		_w61_,
		_w94_
	);
	LUT4 #(
		.INIT('h5a48)
	) name60 (
		g_pad,
		h_pad,
		w_pad,
		x_pad,
		_w95_
	);
	LUT4 #(
		.INIT('hfac8)
	) name61 (
		h_pad,
		i_pad,
		x_pad,
		y_pad,
		_w96_
	);
	LUT4 #(
		.INIT('h21a5)
	) name62 (
		g_pad,
		h_pad,
		w_pad,
		x_pad,
		_w97_
	);
	LUT4 #(
		.INIT('h4f00)
	) name63 (
		_w56_,
		_w60_,
		_w96_,
		_w97_,
		_w98_
	);
	LUT3 #(
		.INIT('h0b)
	) name64 (
		_w94_,
		_w95_,
		_w98_,
		_w99_
	);
	LUT2 #(
		.INIT('h6)
	) name65 (
		h_pad,
		x_pad,
		_w100_
	);
	LUT4 #(
		.INIT('hf40b)
	) name66 (
		_w56_,
		_w60_,
		_w61_,
		_w100_,
		_w101_
	);
	LUT4 #(
		.INIT('h137f)
	) name67 (
		\a0_pad ,
		j_pad,
		k_pad,
		z_pad,
		_w102_
	);
	LUT2 #(
		.INIT('h6)
	) name68 (
		i_pad,
		y_pad,
		_w103_
	);
	LUT3 #(
		.INIT('h4b)
	) name69 (
		_w56_,
		_w102_,
		_w103_,
		_w104_
	);
	LUT4 #(
		.INIT('h32c8)
	) name70 (
		\a0_pad ,
		j_pad,
		k_pad,
		z_pad,
		_w105_
	);
	LUT4 #(
		.INIT('h0013)
	) name71 (
		\a0_pad ,
		\b0_pad ,
		k_pad,
		l_pad,
		_w106_
	);
	LUT2 #(
		.INIT('h2)
	) name72 (
		_w52_,
		_w57_,
		_w107_
	);
	LUT4 #(
		.INIT('h0e0f)
	) name73 (
		_w46_,
		_w50_,
		_w106_,
		_w107_,
		_w108_
	);
	LUT4 #(
		.INIT('hfac8)
	) name74 (
		\a0_pad ,
		\b0_pad ,
		k_pad,
		l_pad,
		_w109_
	);
	LUT4 #(
		.INIT('hef00)
	) name75 (
		_w46_,
		_w50_,
		_w52_,
		_w109_,
		_w110_
	);
	LUT4 #(
		.INIT('h4c13)
	) name76 (
		\a0_pad ,
		j_pad,
		k_pad,
		z_pad,
		_w111_
	);
	LUT4 #(
		.INIT('h7077)
	) name77 (
		_w105_,
		_w108_,
		_w110_,
		_w111_,
		_w112_
	);
	LUT2 #(
		.INIT('h6)
	) name78 (
		\a0_pad ,
		k_pad,
		_w113_
	);
	LUT4 #(
		.INIT('h5a48)
	) name79 (
		\a0_pad ,
		\b0_pad ,
		k_pad,
		l_pad,
		_w114_
	);
	LUT4 #(
		.INIT('hef00)
	) name80 (
		_w46_,
		_w50_,
		_w52_,
		_w114_,
		_w115_
	);
	LUT4 #(
		.INIT('h0021)
	) name81 (
		\a0_pad ,
		\b0_pad ,
		k_pad,
		l_pad,
		_w116_
	);
	LUT2 #(
		.INIT('h2)
	) name82 (
		_w52_,
		_w113_,
		_w117_
	);
	LUT4 #(
		.INIT('h0e0f)
	) name83 (
		_w46_,
		_w50_,
		_w116_,
		_w117_,
		_w118_
	);
	LUT2 #(
		.INIT('h4)
	) name84 (
		_w115_,
		_w118_,
		_w119_
	);
	LUT2 #(
		.INIT('h6)
	) name85 (
		\b0_pad ,
		l_pad,
		_w120_
	);
	LUT4 #(
		.INIT('h01fe)
	) name86 (
		_w46_,
		_w50_,
		_w51_,
		_w120_,
		_w121_
	);
	LUT4 #(
		.INIT('h5510)
	) name87 (
		_w45_,
		_w47_,
		_w48_,
		_w49_,
		_w122_
	);
	LUT4 #(
		.INIT('h5a48)
	) name88 (
		\c0_pad ,
		\d0_pad ,
		m_pad,
		n_pad,
		_w123_
	);
	LUT4 #(
		.INIT('hfac8)
	) name89 (
		\d0_pad ,
		\e0_pad ,
		n_pad,
		o_pad,
		_w124_
	);
	LUT4 #(
		.INIT('h21a5)
	) name90 (
		\c0_pad ,
		\d0_pad ,
		m_pad,
		n_pad,
		_w125_
	);
	LUT4 #(
		.INIT('h4f00)
	) name91 (
		_w47_,
		_w48_,
		_w124_,
		_w125_,
		_w126_
	);
	LUT3 #(
		.INIT('h0b)
	) name92 (
		_w122_,
		_w123_,
		_w126_,
		_w127_
	);
	LUT2 #(
		.INIT('h6)
	) name93 (
		\d0_pad ,
		n_pad,
		_w128_
	);
	LUT4 #(
		.INIT('hf40b)
	) name94 (
		_w47_,
		_w48_,
		_w49_,
		_w128_,
		_w129_
	);
	LUT3 #(
		.INIT('h17)
	) name95 (
		\f0_pad ,
		\g0_pad ,
		p_pad,
		_w130_
	);
	LUT2 #(
		.INIT('h6)
	) name96 (
		\e0_pad ,
		o_pad,
		_w131_
	);
	LUT2 #(
		.INIT('h9)
	) name97 (
		_w130_,
		_w131_,
		_w132_
	);
	LUT3 #(
		.INIT('h96)
	) name98 (
		\f0_pad ,
		\g0_pad ,
		p_pad,
		_w133_
	);
	LUT4 #(
		.INIT('h0517)
	) name99 (
		a_pad,
		b_pad,
		q_pad,
		r_pad,
		_w134_
	);
	LUT4 #(
		.INIT('h135f)
	) name100 (
		a_pad,
		b_pad,
		q_pad,
		r_pad,
		_w135_
	);
	LUT4 #(
		.INIT('h0e0f)
	) name101 (
		_w37_,
		_w69_,
		_w134_,
		_w135_,
		_w136_
	);
	assign \h0_pad  = _w76_ ;
	assign \i0_pad  = _w78_ ;
	assign \j0_pad  = _w83_ ;
	assign \k0_pad  = _w89_ ;
	assign \l0_pad  = _w91_ ;
	assign \m0_pad  = _w93_ ;
	assign \n0_pad  = _w99_ ;
	assign \o0_pad  = _w101_ ;
	assign \p0_pad  = _w104_ ;
	assign \q0_pad  = _w112_ ;
	assign \r0_pad  = _w119_ ;
	assign \s0_pad  = _w121_ ;
	assign \t0_pad  = _w127_ ;
	assign \u0_pad  = _w129_ ;
	assign \v0_pad  = _w132_ ;
	assign \w0_pad  = _w133_ ;
	assign \x0_pad  = _w136_ ;
endmodule;