module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , x255 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , x255 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 ;
  wire n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 ;
  assign n257 = x0 & ~x128 ;
  assign n258 = ~x0 & x128 ;
  assign n259 = ~n257 & ~n258 ;
  assign n260 = x0 & x128 ;
  assign n261 = ~x1 & ~x129 ;
  assign n262 = x1 & x129 ;
  assign n263 = ~n261 & ~n262 ;
  assign n264 = n260 & ~n263 ;
  assign n265 = ~n260 & n263 ;
  assign n266 = ~n264 & ~n265 ;
  assign n267 = n260 & ~n261 ;
  assign n268 = ~n262 & ~n267 ;
  assign n269 = ~x2 & ~x130 ;
  assign n270 = x2 & x130 ;
  assign n271 = ~n269 & ~n270 ;
  assign n272 = n268 & ~n271 ;
  assign n273 = ~n268 & n271 ;
  assign n274 = ~n272 & ~n273 ;
  assign n275 = ~n268 & ~n269 ;
  assign n276 = ~n270 & ~n275 ;
  assign n277 = ~x3 & ~x131 ;
  assign n278 = x3 & x131 ;
  assign n279 = ~n277 & ~n278 ;
  assign n280 = n276 & ~n279 ;
  assign n281 = ~n276 & n279 ;
  assign n282 = ~n280 & ~n281 ;
  assign n283 = ~n276 & ~n277 ;
  assign n284 = ~n278 & ~n283 ;
  assign n285 = ~x4 & ~x132 ;
  assign n286 = x4 & x132 ;
  assign n287 = ~n285 & ~n286 ;
  assign n288 = n284 & ~n287 ;
  assign n289 = ~n284 & n287 ;
  assign n290 = ~n288 & ~n289 ;
  assign n291 = ~n284 & ~n285 ;
  assign n292 = ~n286 & ~n291 ;
  assign n293 = ~x5 & ~x133 ;
  assign n294 = x5 & x133 ;
  assign n295 = ~n293 & ~n294 ;
  assign n296 = n292 & ~n295 ;
  assign n297 = ~n292 & n295 ;
  assign n298 = ~n296 & ~n297 ;
  assign n299 = ~n292 & ~n293 ;
  assign n300 = ~n294 & ~n299 ;
  assign n301 = ~x6 & ~x134 ;
  assign n302 = x6 & x134 ;
  assign n303 = ~n301 & ~n302 ;
  assign n304 = n300 & ~n303 ;
  assign n305 = ~n300 & n303 ;
  assign n306 = ~n304 & ~n305 ;
  assign n307 = ~n300 & ~n301 ;
  assign n308 = ~n302 & ~n307 ;
  assign n309 = ~x7 & ~x135 ;
  assign n310 = x7 & x135 ;
  assign n311 = ~n309 & ~n310 ;
  assign n312 = n308 & ~n311 ;
  assign n313 = ~n308 & n311 ;
  assign n314 = ~n312 & ~n313 ;
  assign n315 = ~n308 & ~n309 ;
  assign n316 = ~n310 & ~n315 ;
  assign n317 = ~x8 & ~x136 ;
  assign n318 = x8 & x136 ;
  assign n319 = ~n317 & ~n318 ;
  assign n320 = n316 & ~n319 ;
  assign n321 = ~n316 & n319 ;
  assign n322 = ~n320 & ~n321 ;
  assign n323 = ~n316 & ~n317 ;
  assign n324 = ~n318 & ~n323 ;
  assign n325 = ~x9 & ~x137 ;
  assign n326 = x9 & x137 ;
  assign n327 = ~n325 & ~n326 ;
  assign n328 = n324 & ~n327 ;
  assign n329 = ~n324 & n327 ;
  assign n330 = ~n328 & ~n329 ;
  assign n331 = ~n324 & ~n325 ;
  assign n332 = ~n326 & ~n331 ;
  assign n333 = ~x10 & ~x138 ;
  assign n334 = x10 & x138 ;
  assign n335 = ~n333 & ~n334 ;
  assign n336 = n332 & ~n335 ;
  assign n337 = ~n332 & n335 ;
  assign n338 = ~n336 & ~n337 ;
  assign n339 = ~n332 & ~n333 ;
  assign n340 = ~n334 & ~n339 ;
  assign n341 = ~x11 & ~x139 ;
  assign n342 = x11 & x139 ;
  assign n343 = ~n341 & ~n342 ;
  assign n344 = n340 & ~n343 ;
  assign n345 = ~n340 & n343 ;
  assign n346 = ~n344 & ~n345 ;
  assign n347 = ~n340 & ~n341 ;
  assign n348 = ~n342 & ~n347 ;
  assign n349 = ~x12 & ~x140 ;
  assign n350 = x12 & x140 ;
  assign n351 = ~n349 & ~n350 ;
  assign n352 = n348 & ~n351 ;
  assign n353 = ~n348 & n351 ;
  assign n354 = ~n352 & ~n353 ;
  assign n355 = ~n348 & ~n349 ;
  assign n356 = ~n350 & ~n355 ;
  assign n357 = ~x13 & ~x141 ;
  assign n358 = x13 & x141 ;
  assign n359 = ~n357 & ~n358 ;
  assign n360 = n356 & ~n359 ;
  assign n361 = ~n356 & n359 ;
  assign n362 = ~n360 & ~n361 ;
  assign n363 = ~n356 & ~n357 ;
  assign n364 = ~n358 & ~n363 ;
  assign n365 = ~x14 & ~x142 ;
  assign n366 = x14 & x142 ;
  assign n367 = ~n365 & ~n366 ;
  assign n368 = n364 & ~n367 ;
  assign n369 = ~n364 & n367 ;
  assign n370 = ~n368 & ~n369 ;
  assign n371 = ~n364 & ~n365 ;
  assign n372 = ~n366 & ~n371 ;
  assign n373 = ~x15 & ~x143 ;
  assign n374 = x15 & x143 ;
  assign n375 = ~n373 & ~n374 ;
  assign n376 = n372 & ~n375 ;
  assign n377 = ~n372 & n375 ;
  assign n378 = ~n376 & ~n377 ;
  assign n379 = ~n372 & ~n373 ;
  assign n380 = ~n374 & ~n379 ;
  assign n381 = ~x16 & ~x144 ;
  assign n382 = x16 & x144 ;
  assign n383 = ~n381 & ~n382 ;
  assign n384 = n380 & ~n383 ;
  assign n385 = ~n380 & n383 ;
  assign n386 = ~n384 & ~n385 ;
  assign n387 = ~n380 & ~n381 ;
  assign n388 = ~n382 & ~n387 ;
  assign n389 = ~x17 & ~x145 ;
  assign n390 = x17 & x145 ;
  assign n391 = ~n389 & ~n390 ;
  assign n392 = n388 & ~n391 ;
  assign n393 = ~n388 & n391 ;
  assign n394 = ~n392 & ~n393 ;
  assign n395 = ~n388 & ~n389 ;
  assign n396 = ~n390 & ~n395 ;
  assign n397 = ~x18 & ~x146 ;
  assign n398 = x18 & x146 ;
  assign n399 = ~n397 & ~n398 ;
  assign n400 = n396 & ~n399 ;
  assign n401 = ~n396 & n399 ;
  assign n402 = ~n400 & ~n401 ;
  assign n403 = ~n396 & ~n397 ;
  assign n404 = ~n398 & ~n403 ;
  assign n405 = ~x19 & ~x147 ;
  assign n406 = x19 & x147 ;
  assign n407 = ~n405 & ~n406 ;
  assign n408 = n404 & ~n407 ;
  assign n409 = ~n404 & n407 ;
  assign n410 = ~n408 & ~n409 ;
  assign n411 = ~n404 & ~n405 ;
  assign n412 = ~n406 & ~n411 ;
  assign n413 = ~x20 & ~x148 ;
  assign n414 = x20 & x148 ;
  assign n415 = ~n413 & ~n414 ;
  assign n416 = n412 & ~n415 ;
  assign n417 = ~n412 & n415 ;
  assign n418 = ~n416 & ~n417 ;
  assign n419 = ~n412 & ~n413 ;
  assign n420 = ~n414 & ~n419 ;
  assign n421 = ~x21 & ~x149 ;
  assign n422 = x21 & x149 ;
  assign n423 = ~n421 & ~n422 ;
  assign n424 = n420 & ~n423 ;
  assign n425 = ~n420 & n423 ;
  assign n426 = ~n424 & ~n425 ;
  assign n427 = ~n420 & ~n421 ;
  assign n428 = ~n422 & ~n427 ;
  assign n429 = ~x22 & ~x150 ;
  assign n430 = x22 & x150 ;
  assign n431 = ~n429 & ~n430 ;
  assign n432 = n428 & ~n431 ;
  assign n433 = ~n428 & n431 ;
  assign n434 = ~n432 & ~n433 ;
  assign n435 = ~n428 & ~n429 ;
  assign n436 = ~n430 & ~n435 ;
  assign n437 = ~x23 & ~x151 ;
  assign n438 = x23 & x151 ;
  assign n439 = ~n437 & ~n438 ;
  assign n440 = n436 & ~n439 ;
  assign n441 = ~n436 & n439 ;
  assign n442 = ~n440 & ~n441 ;
  assign n443 = ~n436 & ~n437 ;
  assign n444 = ~n438 & ~n443 ;
  assign n445 = ~x24 & ~x152 ;
  assign n446 = x24 & x152 ;
  assign n447 = ~n445 & ~n446 ;
  assign n448 = n444 & ~n447 ;
  assign n449 = ~n444 & n447 ;
  assign n450 = ~n448 & ~n449 ;
  assign n451 = ~n444 & ~n445 ;
  assign n452 = ~n446 & ~n451 ;
  assign n453 = ~x25 & ~x153 ;
  assign n454 = x25 & x153 ;
  assign n455 = ~n453 & ~n454 ;
  assign n456 = n452 & ~n455 ;
  assign n457 = ~n452 & n455 ;
  assign n458 = ~n456 & ~n457 ;
  assign n459 = ~n452 & ~n453 ;
  assign n460 = ~n454 & ~n459 ;
  assign n461 = ~x26 & ~x154 ;
  assign n462 = x26 & x154 ;
  assign n463 = ~n461 & ~n462 ;
  assign n464 = n460 & ~n463 ;
  assign n465 = ~n460 & n463 ;
  assign n466 = ~n464 & ~n465 ;
  assign n467 = ~n460 & ~n461 ;
  assign n468 = ~n462 & ~n467 ;
  assign n469 = ~x27 & ~x155 ;
  assign n470 = x27 & x155 ;
  assign n471 = ~n469 & ~n470 ;
  assign n472 = n468 & ~n471 ;
  assign n473 = ~n468 & n471 ;
  assign n474 = ~n472 & ~n473 ;
  assign n475 = ~n468 & ~n469 ;
  assign n476 = ~n470 & ~n475 ;
  assign n477 = ~x28 & ~x156 ;
  assign n478 = x28 & x156 ;
  assign n479 = ~n477 & ~n478 ;
  assign n480 = n476 & ~n479 ;
  assign n481 = ~n476 & n479 ;
  assign n482 = ~n480 & ~n481 ;
  assign n483 = ~n476 & ~n477 ;
  assign n484 = ~n478 & ~n483 ;
  assign n485 = ~x29 & ~x157 ;
  assign n486 = x29 & x157 ;
  assign n487 = ~n485 & ~n486 ;
  assign n488 = n484 & ~n487 ;
  assign n489 = ~n484 & n487 ;
  assign n490 = ~n488 & ~n489 ;
  assign n491 = ~n484 & ~n485 ;
  assign n492 = ~n486 & ~n491 ;
  assign n493 = ~x30 & ~x158 ;
  assign n494 = x30 & x158 ;
  assign n495 = ~n493 & ~n494 ;
  assign n496 = n492 & ~n495 ;
  assign n497 = ~n492 & n495 ;
  assign n498 = ~n496 & ~n497 ;
  assign n499 = ~n492 & ~n493 ;
  assign n500 = ~n494 & ~n499 ;
  assign n501 = ~x31 & ~x159 ;
  assign n502 = x31 & x159 ;
  assign n503 = ~n501 & ~n502 ;
  assign n504 = n500 & ~n503 ;
  assign n505 = ~n500 & n503 ;
  assign n506 = ~n504 & ~n505 ;
  assign n507 = ~n500 & ~n501 ;
  assign n508 = ~n502 & ~n507 ;
  assign n509 = ~x32 & ~x160 ;
  assign n510 = x32 & x160 ;
  assign n511 = ~n509 & ~n510 ;
  assign n512 = n508 & ~n511 ;
  assign n513 = ~n508 & n511 ;
  assign n514 = ~n512 & ~n513 ;
  assign n515 = ~n508 & ~n509 ;
  assign n516 = ~n510 & ~n515 ;
  assign n517 = ~x33 & ~x161 ;
  assign n518 = x33 & x161 ;
  assign n519 = ~n517 & ~n518 ;
  assign n520 = n516 & ~n519 ;
  assign n521 = ~n516 & n519 ;
  assign n522 = ~n520 & ~n521 ;
  assign n523 = ~n516 & ~n517 ;
  assign n524 = ~n518 & ~n523 ;
  assign n525 = ~x34 & ~x162 ;
  assign n526 = x34 & x162 ;
  assign n527 = ~n525 & ~n526 ;
  assign n528 = n524 & ~n527 ;
  assign n529 = ~n524 & n527 ;
  assign n530 = ~n528 & ~n529 ;
  assign n531 = ~n524 & ~n525 ;
  assign n532 = ~n526 & ~n531 ;
  assign n533 = ~x35 & ~x163 ;
  assign n534 = x35 & x163 ;
  assign n535 = ~n533 & ~n534 ;
  assign n536 = n532 & ~n535 ;
  assign n537 = ~n532 & n535 ;
  assign n538 = ~n536 & ~n537 ;
  assign n539 = ~n532 & ~n533 ;
  assign n540 = ~n534 & ~n539 ;
  assign n541 = ~x36 & ~x164 ;
  assign n542 = x36 & x164 ;
  assign n543 = ~n541 & ~n542 ;
  assign n544 = n540 & ~n543 ;
  assign n545 = ~n540 & n543 ;
  assign n546 = ~n544 & ~n545 ;
  assign n547 = ~n540 & ~n541 ;
  assign n548 = ~n542 & ~n547 ;
  assign n549 = ~x37 & ~x165 ;
  assign n550 = x37 & x165 ;
  assign n551 = ~n549 & ~n550 ;
  assign n552 = n548 & ~n551 ;
  assign n553 = ~n548 & n551 ;
  assign n554 = ~n552 & ~n553 ;
  assign n555 = ~n548 & ~n549 ;
  assign n556 = ~n550 & ~n555 ;
  assign n557 = ~x38 & ~x166 ;
  assign n558 = x38 & x166 ;
  assign n559 = ~n557 & ~n558 ;
  assign n560 = n556 & ~n559 ;
  assign n561 = ~n556 & n559 ;
  assign n562 = ~n560 & ~n561 ;
  assign n563 = ~n556 & ~n557 ;
  assign n564 = ~n558 & ~n563 ;
  assign n565 = ~x39 & ~x167 ;
  assign n566 = x39 & x167 ;
  assign n567 = ~n565 & ~n566 ;
  assign n568 = n564 & ~n567 ;
  assign n569 = ~n564 & n567 ;
  assign n570 = ~n568 & ~n569 ;
  assign n571 = ~n564 & ~n565 ;
  assign n572 = ~n566 & ~n571 ;
  assign n573 = ~x40 & ~x168 ;
  assign n574 = x40 & x168 ;
  assign n575 = ~n573 & ~n574 ;
  assign n576 = n572 & ~n575 ;
  assign n577 = ~n572 & n575 ;
  assign n578 = ~n576 & ~n577 ;
  assign n579 = ~n572 & ~n573 ;
  assign n580 = ~n574 & ~n579 ;
  assign n581 = ~x41 & ~x169 ;
  assign n582 = x41 & x169 ;
  assign n583 = ~n581 & ~n582 ;
  assign n584 = n580 & ~n583 ;
  assign n585 = ~n580 & n583 ;
  assign n586 = ~n584 & ~n585 ;
  assign n587 = ~n580 & ~n581 ;
  assign n588 = ~n582 & ~n587 ;
  assign n589 = ~x42 & ~x170 ;
  assign n590 = x42 & x170 ;
  assign n591 = ~n589 & ~n590 ;
  assign n592 = n588 & ~n591 ;
  assign n593 = ~n588 & n591 ;
  assign n594 = ~n592 & ~n593 ;
  assign n595 = ~n588 & ~n589 ;
  assign n596 = ~n590 & ~n595 ;
  assign n597 = ~x43 & ~x171 ;
  assign n598 = x43 & x171 ;
  assign n599 = ~n597 & ~n598 ;
  assign n600 = n596 & ~n599 ;
  assign n601 = ~n596 & n599 ;
  assign n602 = ~n600 & ~n601 ;
  assign n603 = ~n596 & ~n597 ;
  assign n604 = ~n598 & ~n603 ;
  assign n605 = ~x44 & ~x172 ;
  assign n606 = x44 & x172 ;
  assign n607 = ~n605 & ~n606 ;
  assign n608 = n604 & ~n607 ;
  assign n609 = ~n604 & n607 ;
  assign n610 = ~n608 & ~n609 ;
  assign n611 = ~n604 & ~n605 ;
  assign n612 = ~n606 & ~n611 ;
  assign n613 = ~x45 & ~x173 ;
  assign n614 = x45 & x173 ;
  assign n615 = ~n613 & ~n614 ;
  assign n616 = n612 & ~n615 ;
  assign n617 = ~n612 & n615 ;
  assign n618 = ~n616 & ~n617 ;
  assign n619 = ~n612 & ~n613 ;
  assign n620 = ~n614 & ~n619 ;
  assign n621 = ~x46 & ~x174 ;
  assign n622 = x46 & x174 ;
  assign n623 = ~n621 & ~n622 ;
  assign n624 = n620 & ~n623 ;
  assign n625 = ~n620 & n623 ;
  assign n626 = ~n624 & ~n625 ;
  assign n627 = ~n620 & ~n621 ;
  assign n628 = ~n622 & ~n627 ;
  assign n629 = ~x47 & ~x175 ;
  assign n630 = x47 & x175 ;
  assign n631 = ~n629 & ~n630 ;
  assign n632 = n628 & ~n631 ;
  assign n633 = ~n628 & n631 ;
  assign n634 = ~n632 & ~n633 ;
  assign n635 = ~n628 & ~n629 ;
  assign n636 = ~n630 & ~n635 ;
  assign n637 = ~x48 & ~x176 ;
  assign n638 = x48 & x176 ;
  assign n639 = ~n637 & ~n638 ;
  assign n640 = n636 & ~n639 ;
  assign n641 = ~n636 & n639 ;
  assign n642 = ~n640 & ~n641 ;
  assign n643 = ~n636 & ~n637 ;
  assign n644 = ~n638 & ~n643 ;
  assign n645 = ~x49 & ~x177 ;
  assign n646 = x49 & x177 ;
  assign n647 = ~n645 & ~n646 ;
  assign n648 = n644 & ~n647 ;
  assign n649 = ~n644 & n647 ;
  assign n650 = ~n648 & ~n649 ;
  assign n651 = ~n644 & ~n645 ;
  assign n652 = ~n646 & ~n651 ;
  assign n653 = ~x50 & ~x178 ;
  assign n654 = x50 & x178 ;
  assign n655 = ~n653 & ~n654 ;
  assign n656 = n652 & ~n655 ;
  assign n657 = ~n652 & n655 ;
  assign n658 = ~n656 & ~n657 ;
  assign n659 = ~n652 & ~n653 ;
  assign n660 = ~n654 & ~n659 ;
  assign n661 = ~x51 & ~x179 ;
  assign n662 = x51 & x179 ;
  assign n663 = ~n661 & ~n662 ;
  assign n664 = n660 & ~n663 ;
  assign n665 = ~n660 & n663 ;
  assign n666 = ~n664 & ~n665 ;
  assign n667 = ~n660 & ~n661 ;
  assign n668 = ~n662 & ~n667 ;
  assign n669 = ~x52 & ~x180 ;
  assign n670 = x52 & x180 ;
  assign n671 = ~n669 & ~n670 ;
  assign n672 = n668 & ~n671 ;
  assign n673 = ~n668 & n671 ;
  assign n674 = ~n672 & ~n673 ;
  assign n675 = ~n668 & ~n669 ;
  assign n676 = ~n670 & ~n675 ;
  assign n677 = ~x53 & ~x181 ;
  assign n678 = x53 & x181 ;
  assign n679 = ~n677 & ~n678 ;
  assign n680 = n676 & ~n679 ;
  assign n681 = ~n676 & n679 ;
  assign n682 = ~n680 & ~n681 ;
  assign n683 = ~n676 & ~n677 ;
  assign n684 = ~n678 & ~n683 ;
  assign n685 = ~x54 & ~x182 ;
  assign n686 = x54 & x182 ;
  assign n687 = ~n685 & ~n686 ;
  assign n688 = n684 & ~n687 ;
  assign n689 = ~n684 & n687 ;
  assign n690 = ~n688 & ~n689 ;
  assign n691 = ~n684 & ~n685 ;
  assign n692 = ~n686 & ~n691 ;
  assign n693 = ~x55 & ~x183 ;
  assign n694 = x55 & x183 ;
  assign n695 = ~n693 & ~n694 ;
  assign n696 = n692 & ~n695 ;
  assign n697 = ~n692 & n695 ;
  assign n698 = ~n696 & ~n697 ;
  assign n699 = ~n692 & ~n693 ;
  assign n700 = ~n694 & ~n699 ;
  assign n701 = ~x56 & ~x184 ;
  assign n702 = x56 & x184 ;
  assign n703 = ~n701 & ~n702 ;
  assign n704 = n700 & ~n703 ;
  assign n705 = ~n700 & n703 ;
  assign n706 = ~n704 & ~n705 ;
  assign n707 = ~n700 & ~n701 ;
  assign n708 = ~n702 & ~n707 ;
  assign n709 = ~x57 & ~x185 ;
  assign n710 = x57 & x185 ;
  assign n711 = ~n709 & ~n710 ;
  assign n712 = n708 & ~n711 ;
  assign n713 = ~n708 & n711 ;
  assign n714 = ~n712 & ~n713 ;
  assign n715 = ~n708 & ~n709 ;
  assign n716 = ~n710 & ~n715 ;
  assign n717 = ~x58 & ~x186 ;
  assign n718 = x58 & x186 ;
  assign n719 = ~n717 & ~n718 ;
  assign n720 = n716 & ~n719 ;
  assign n721 = ~n716 & n719 ;
  assign n722 = ~n720 & ~n721 ;
  assign n723 = ~n716 & ~n717 ;
  assign n724 = ~n718 & ~n723 ;
  assign n725 = ~x59 & ~x187 ;
  assign n726 = x59 & x187 ;
  assign n727 = ~n725 & ~n726 ;
  assign n728 = n724 & ~n727 ;
  assign n729 = ~n724 & n727 ;
  assign n730 = ~n728 & ~n729 ;
  assign n731 = ~n724 & ~n725 ;
  assign n732 = ~n726 & ~n731 ;
  assign n733 = ~x60 & ~x188 ;
  assign n734 = x60 & x188 ;
  assign n735 = ~n733 & ~n734 ;
  assign n736 = n732 & ~n735 ;
  assign n737 = ~n732 & n735 ;
  assign n738 = ~n736 & ~n737 ;
  assign n739 = ~n732 & ~n733 ;
  assign n740 = ~n734 & ~n739 ;
  assign n741 = ~x61 & ~x189 ;
  assign n742 = x61 & x189 ;
  assign n743 = ~n741 & ~n742 ;
  assign n744 = n740 & ~n743 ;
  assign n745 = ~n740 & n743 ;
  assign n746 = ~n744 & ~n745 ;
  assign n747 = ~n740 & ~n741 ;
  assign n748 = ~n742 & ~n747 ;
  assign n749 = ~x62 & ~x190 ;
  assign n750 = x62 & x190 ;
  assign n751 = ~n749 & ~n750 ;
  assign n752 = n748 & ~n751 ;
  assign n753 = ~n748 & n751 ;
  assign n754 = ~n752 & ~n753 ;
  assign n755 = ~n748 & ~n749 ;
  assign n756 = ~n750 & ~n755 ;
  assign n757 = ~x63 & ~x191 ;
  assign n758 = x63 & x191 ;
  assign n759 = ~n757 & ~n758 ;
  assign n760 = n756 & ~n759 ;
  assign n761 = ~n756 & n759 ;
  assign n762 = ~n760 & ~n761 ;
  assign n763 = ~n756 & ~n757 ;
  assign n764 = ~n758 & ~n763 ;
  assign n765 = ~x64 & ~x192 ;
  assign n766 = x64 & x192 ;
  assign n767 = ~n765 & ~n766 ;
  assign n768 = n764 & ~n767 ;
  assign n769 = ~n764 & n767 ;
  assign n770 = ~n768 & ~n769 ;
  assign n771 = ~n764 & ~n765 ;
  assign n772 = ~n766 & ~n771 ;
  assign n773 = ~x65 & ~x193 ;
  assign n774 = x65 & x193 ;
  assign n775 = ~n773 & ~n774 ;
  assign n776 = n772 & ~n775 ;
  assign n777 = ~n772 & n775 ;
  assign n778 = ~n776 & ~n777 ;
  assign n779 = ~n772 & ~n773 ;
  assign n780 = ~n774 & ~n779 ;
  assign n781 = ~x66 & ~x194 ;
  assign n782 = x66 & x194 ;
  assign n783 = ~n781 & ~n782 ;
  assign n784 = n780 & ~n783 ;
  assign n785 = ~n780 & n783 ;
  assign n786 = ~n784 & ~n785 ;
  assign n787 = ~n780 & ~n781 ;
  assign n788 = ~n782 & ~n787 ;
  assign n789 = ~x67 & ~x195 ;
  assign n790 = x67 & x195 ;
  assign n791 = ~n789 & ~n790 ;
  assign n792 = n788 & ~n791 ;
  assign n793 = ~n788 & n791 ;
  assign n794 = ~n792 & ~n793 ;
  assign n795 = ~n788 & ~n789 ;
  assign n796 = ~n790 & ~n795 ;
  assign n797 = ~x68 & ~x196 ;
  assign n798 = x68 & x196 ;
  assign n799 = ~n797 & ~n798 ;
  assign n800 = n796 & ~n799 ;
  assign n801 = ~n796 & n799 ;
  assign n802 = ~n800 & ~n801 ;
  assign n803 = ~n796 & ~n797 ;
  assign n804 = ~n798 & ~n803 ;
  assign n805 = ~x69 & ~x197 ;
  assign n806 = x69 & x197 ;
  assign n807 = ~n805 & ~n806 ;
  assign n808 = n804 & ~n807 ;
  assign n809 = ~n804 & n807 ;
  assign n810 = ~n808 & ~n809 ;
  assign n811 = ~n804 & ~n805 ;
  assign n812 = ~n806 & ~n811 ;
  assign n813 = ~x70 & ~x198 ;
  assign n814 = x70 & x198 ;
  assign n815 = ~n813 & ~n814 ;
  assign n816 = n812 & ~n815 ;
  assign n817 = ~n812 & n815 ;
  assign n818 = ~n816 & ~n817 ;
  assign n819 = ~n812 & ~n813 ;
  assign n820 = ~n814 & ~n819 ;
  assign n821 = ~x71 & ~x199 ;
  assign n822 = x71 & x199 ;
  assign n823 = ~n821 & ~n822 ;
  assign n824 = n820 & ~n823 ;
  assign n825 = ~n820 & n823 ;
  assign n826 = ~n824 & ~n825 ;
  assign n827 = ~n820 & ~n821 ;
  assign n828 = ~n822 & ~n827 ;
  assign n829 = ~x72 & ~x200 ;
  assign n830 = x72 & x200 ;
  assign n831 = ~n829 & ~n830 ;
  assign n832 = n828 & ~n831 ;
  assign n833 = ~n828 & n831 ;
  assign n834 = ~n832 & ~n833 ;
  assign n835 = ~n828 & ~n829 ;
  assign n836 = ~n830 & ~n835 ;
  assign n837 = ~x73 & ~x201 ;
  assign n838 = x73 & x201 ;
  assign n839 = ~n837 & ~n838 ;
  assign n840 = n836 & ~n839 ;
  assign n841 = ~n836 & n839 ;
  assign n842 = ~n840 & ~n841 ;
  assign n843 = ~n836 & ~n837 ;
  assign n844 = ~n838 & ~n843 ;
  assign n845 = ~x74 & ~x202 ;
  assign n846 = x74 & x202 ;
  assign n847 = ~n845 & ~n846 ;
  assign n848 = n844 & ~n847 ;
  assign n849 = ~n844 & n847 ;
  assign n850 = ~n848 & ~n849 ;
  assign n851 = ~n844 & ~n845 ;
  assign n852 = ~n846 & ~n851 ;
  assign n853 = ~x75 & ~x203 ;
  assign n854 = x75 & x203 ;
  assign n855 = ~n853 & ~n854 ;
  assign n856 = n852 & ~n855 ;
  assign n857 = ~n852 & n855 ;
  assign n858 = ~n856 & ~n857 ;
  assign n859 = ~n852 & ~n853 ;
  assign n860 = ~n854 & ~n859 ;
  assign n861 = ~x76 & ~x204 ;
  assign n862 = x76 & x204 ;
  assign n863 = ~n861 & ~n862 ;
  assign n864 = n860 & ~n863 ;
  assign n865 = ~n860 & n863 ;
  assign n866 = ~n864 & ~n865 ;
  assign n867 = ~n860 & ~n861 ;
  assign n868 = ~n862 & ~n867 ;
  assign n869 = ~x77 & ~x205 ;
  assign n870 = x77 & x205 ;
  assign n871 = ~n869 & ~n870 ;
  assign n872 = n868 & ~n871 ;
  assign n873 = ~n868 & n871 ;
  assign n874 = ~n872 & ~n873 ;
  assign n875 = ~n868 & ~n869 ;
  assign n876 = ~n870 & ~n875 ;
  assign n877 = ~x78 & ~x206 ;
  assign n878 = x78 & x206 ;
  assign n879 = ~n877 & ~n878 ;
  assign n880 = n876 & ~n879 ;
  assign n881 = ~n876 & n879 ;
  assign n882 = ~n880 & ~n881 ;
  assign n883 = ~n876 & ~n877 ;
  assign n884 = ~n878 & ~n883 ;
  assign n885 = ~x79 & ~x207 ;
  assign n886 = x79 & x207 ;
  assign n887 = ~n885 & ~n886 ;
  assign n888 = n884 & ~n887 ;
  assign n889 = ~n884 & n887 ;
  assign n890 = ~n888 & ~n889 ;
  assign n891 = ~n884 & ~n885 ;
  assign n892 = ~n886 & ~n891 ;
  assign n893 = ~x80 & ~x208 ;
  assign n894 = x80 & x208 ;
  assign n895 = ~n893 & ~n894 ;
  assign n896 = n892 & ~n895 ;
  assign n897 = ~n892 & n895 ;
  assign n898 = ~n896 & ~n897 ;
  assign n899 = ~n892 & ~n893 ;
  assign n900 = ~n894 & ~n899 ;
  assign n901 = ~x81 & ~x209 ;
  assign n902 = x81 & x209 ;
  assign n903 = ~n901 & ~n902 ;
  assign n904 = n900 & ~n903 ;
  assign n905 = ~n900 & n903 ;
  assign n906 = ~n904 & ~n905 ;
  assign n907 = ~n900 & ~n901 ;
  assign n908 = ~n902 & ~n907 ;
  assign n909 = ~x82 & ~x210 ;
  assign n910 = x82 & x210 ;
  assign n911 = ~n909 & ~n910 ;
  assign n912 = n908 & ~n911 ;
  assign n913 = ~n908 & n911 ;
  assign n914 = ~n912 & ~n913 ;
  assign n915 = ~n908 & ~n909 ;
  assign n916 = ~n910 & ~n915 ;
  assign n917 = ~x83 & ~x211 ;
  assign n918 = x83 & x211 ;
  assign n919 = ~n917 & ~n918 ;
  assign n920 = n916 & ~n919 ;
  assign n921 = ~n916 & n919 ;
  assign n922 = ~n920 & ~n921 ;
  assign n923 = ~n916 & ~n917 ;
  assign n924 = ~n918 & ~n923 ;
  assign n925 = ~x84 & ~x212 ;
  assign n926 = x84 & x212 ;
  assign n927 = ~n925 & ~n926 ;
  assign n928 = n924 & ~n927 ;
  assign n929 = ~n924 & n927 ;
  assign n930 = ~n928 & ~n929 ;
  assign n931 = ~n924 & ~n925 ;
  assign n932 = ~n926 & ~n931 ;
  assign n933 = ~x85 & ~x213 ;
  assign n934 = x85 & x213 ;
  assign n935 = ~n933 & ~n934 ;
  assign n936 = n932 & ~n935 ;
  assign n937 = ~n932 & n935 ;
  assign n938 = ~n936 & ~n937 ;
  assign n939 = ~n932 & ~n933 ;
  assign n940 = ~n934 & ~n939 ;
  assign n941 = ~x86 & ~x214 ;
  assign n942 = x86 & x214 ;
  assign n943 = ~n941 & ~n942 ;
  assign n944 = n940 & ~n943 ;
  assign n945 = ~n940 & n943 ;
  assign n946 = ~n944 & ~n945 ;
  assign n947 = ~n940 & ~n941 ;
  assign n948 = ~n942 & ~n947 ;
  assign n949 = ~x87 & ~x215 ;
  assign n950 = x87 & x215 ;
  assign n951 = ~n949 & ~n950 ;
  assign n952 = n948 & ~n951 ;
  assign n953 = ~n948 & n951 ;
  assign n954 = ~n952 & ~n953 ;
  assign n955 = ~n948 & ~n949 ;
  assign n956 = ~n950 & ~n955 ;
  assign n957 = ~x88 & ~x216 ;
  assign n958 = x88 & x216 ;
  assign n959 = ~n957 & ~n958 ;
  assign n960 = n956 & ~n959 ;
  assign n961 = ~n956 & n959 ;
  assign n962 = ~n960 & ~n961 ;
  assign n963 = ~n956 & ~n957 ;
  assign n964 = ~n958 & ~n963 ;
  assign n965 = ~x89 & ~x217 ;
  assign n966 = x89 & x217 ;
  assign n967 = ~n965 & ~n966 ;
  assign n968 = n964 & ~n967 ;
  assign n969 = ~n964 & n967 ;
  assign n970 = ~n968 & ~n969 ;
  assign n971 = ~n964 & ~n965 ;
  assign n972 = ~n966 & ~n971 ;
  assign n973 = ~x90 & ~x218 ;
  assign n974 = x90 & x218 ;
  assign n975 = ~n973 & ~n974 ;
  assign n976 = n972 & ~n975 ;
  assign n977 = ~n972 & n975 ;
  assign n978 = ~n976 & ~n977 ;
  assign n979 = ~n972 & ~n973 ;
  assign n980 = ~n974 & ~n979 ;
  assign n981 = ~x91 & ~x219 ;
  assign n982 = x91 & x219 ;
  assign n983 = ~n981 & ~n982 ;
  assign n984 = n980 & ~n983 ;
  assign n985 = ~n980 & n983 ;
  assign n986 = ~n984 & ~n985 ;
  assign n987 = ~n980 & ~n981 ;
  assign n988 = ~n982 & ~n987 ;
  assign n989 = ~x92 & ~x220 ;
  assign n990 = x92 & x220 ;
  assign n991 = ~n989 & ~n990 ;
  assign n992 = n988 & ~n991 ;
  assign n993 = ~n988 & n991 ;
  assign n994 = ~n992 & ~n993 ;
  assign n995 = ~n988 & ~n989 ;
  assign n996 = ~n990 & ~n995 ;
  assign n997 = ~x93 & ~x221 ;
  assign n998 = x93 & x221 ;
  assign n999 = ~n997 & ~n998 ;
  assign n1000 = n996 & ~n999 ;
  assign n1001 = ~n996 & n999 ;
  assign n1002 = ~n1000 & ~n1001 ;
  assign n1003 = ~n996 & ~n997 ;
  assign n1004 = ~n998 & ~n1003 ;
  assign n1005 = ~x94 & ~x222 ;
  assign n1006 = x94 & x222 ;
  assign n1007 = ~n1005 & ~n1006 ;
  assign n1008 = n1004 & ~n1007 ;
  assign n1009 = ~n1004 & n1007 ;
  assign n1010 = ~n1008 & ~n1009 ;
  assign n1011 = ~n1004 & ~n1005 ;
  assign n1012 = ~n1006 & ~n1011 ;
  assign n1013 = ~x95 & ~x223 ;
  assign n1014 = x95 & x223 ;
  assign n1015 = ~n1013 & ~n1014 ;
  assign n1016 = n1012 & ~n1015 ;
  assign n1017 = ~n1012 & n1015 ;
  assign n1018 = ~n1016 & ~n1017 ;
  assign n1019 = ~n1012 & ~n1013 ;
  assign n1020 = ~n1014 & ~n1019 ;
  assign n1021 = ~x96 & ~x224 ;
  assign n1022 = x96 & x224 ;
  assign n1023 = ~n1021 & ~n1022 ;
  assign n1024 = n1020 & ~n1023 ;
  assign n1025 = ~n1020 & n1023 ;
  assign n1026 = ~n1024 & ~n1025 ;
  assign n1027 = ~n1020 & ~n1021 ;
  assign n1028 = ~n1022 & ~n1027 ;
  assign n1029 = ~x97 & ~x225 ;
  assign n1030 = x97 & x225 ;
  assign n1031 = ~n1029 & ~n1030 ;
  assign n1032 = n1028 & ~n1031 ;
  assign n1033 = ~n1028 & n1031 ;
  assign n1034 = ~n1032 & ~n1033 ;
  assign n1035 = ~n1028 & ~n1029 ;
  assign n1036 = ~n1030 & ~n1035 ;
  assign n1037 = ~x98 & ~x226 ;
  assign n1038 = x98 & x226 ;
  assign n1039 = ~n1037 & ~n1038 ;
  assign n1040 = n1036 & ~n1039 ;
  assign n1041 = ~n1036 & n1039 ;
  assign n1042 = ~n1040 & ~n1041 ;
  assign n1043 = ~n1036 & ~n1037 ;
  assign n1044 = ~n1038 & ~n1043 ;
  assign n1045 = ~x99 & ~x227 ;
  assign n1046 = x99 & x227 ;
  assign n1047 = ~n1045 & ~n1046 ;
  assign n1048 = n1044 & ~n1047 ;
  assign n1049 = ~n1044 & n1047 ;
  assign n1050 = ~n1048 & ~n1049 ;
  assign n1051 = ~n1044 & ~n1045 ;
  assign n1052 = ~n1046 & ~n1051 ;
  assign n1053 = ~x100 & ~x228 ;
  assign n1054 = x100 & x228 ;
  assign n1055 = ~n1053 & ~n1054 ;
  assign n1056 = n1052 & ~n1055 ;
  assign n1057 = ~n1052 & n1055 ;
  assign n1058 = ~n1056 & ~n1057 ;
  assign n1059 = ~n1052 & ~n1053 ;
  assign n1060 = ~n1054 & ~n1059 ;
  assign n1061 = ~x101 & ~x229 ;
  assign n1062 = x101 & x229 ;
  assign n1063 = ~n1061 & ~n1062 ;
  assign n1064 = n1060 & ~n1063 ;
  assign n1065 = ~n1060 & n1063 ;
  assign n1066 = ~n1064 & ~n1065 ;
  assign n1067 = ~n1060 & ~n1061 ;
  assign n1068 = ~n1062 & ~n1067 ;
  assign n1069 = ~x102 & ~x230 ;
  assign n1070 = x102 & x230 ;
  assign n1071 = ~n1069 & ~n1070 ;
  assign n1072 = n1068 & ~n1071 ;
  assign n1073 = ~n1068 & n1071 ;
  assign n1074 = ~n1072 & ~n1073 ;
  assign n1075 = ~n1068 & ~n1069 ;
  assign n1076 = ~n1070 & ~n1075 ;
  assign n1077 = ~x103 & ~x231 ;
  assign n1078 = x103 & x231 ;
  assign n1079 = ~n1077 & ~n1078 ;
  assign n1080 = n1076 & ~n1079 ;
  assign n1081 = ~n1076 & n1079 ;
  assign n1082 = ~n1080 & ~n1081 ;
  assign n1083 = ~n1076 & ~n1077 ;
  assign n1084 = ~n1078 & ~n1083 ;
  assign n1085 = ~x104 & ~x232 ;
  assign n1086 = x104 & x232 ;
  assign n1087 = ~n1085 & ~n1086 ;
  assign n1088 = n1084 & ~n1087 ;
  assign n1089 = ~n1084 & n1087 ;
  assign n1090 = ~n1088 & ~n1089 ;
  assign n1091 = ~n1084 & ~n1085 ;
  assign n1092 = ~n1086 & ~n1091 ;
  assign n1093 = ~x105 & ~x233 ;
  assign n1094 = x105 & x233 ;
  assign n1095 = ~n1093 & ~n1094 ;
  assign n1096 = n1092 & ~n1095 ;
  assign n1097 = ~n1092 & n1095 ;
  assign n1098 = ~n1096 & ~n1097 ;
  assign n1099 = ~n1092 & ~n1093 ;
  assign n1100 = ~n1094 & ~n1099 ;
  assign n1101 = ~x106 & ~x234 ;
  assign n1102 = x106 & x234 ;
  assign n1103 = ~n1101 & ~n1102 ;
  assign n1104 = n1100 & ~n1103 ;
  assign n1105 = ~n1100 & n1103 ;
  assign n1106 = ~n1104 & ~n1105 ;
  assign n1107 = ~n1100 & ~n1101 ;
  assign n1108 = ~n1102 & ~n1107 ;
  assign n1109 = ~x107 & ~x235 ;
  assign n1110 = x107 & x235 ;
  assign n1111 = ~n1109 & ~n1110 ;
  assign n1112 = n1108 & ~n1111 ;
  assign n1113 = ~n1108 & n1111 ;
  assign n1114 = ~n1112 & ~n1113 ;
  assign n1115 = ~n1108 & ~n1109 ;
  assign n1116 = ~n1110 & ~n1115 ;
  assign n1117 = ~x108 & ~x236 ;
  assign n1118 = x108 & x236 ;
  assign n1119 = ~n1117 & ~n1118 ;
  assign n1120 = n1116 & ~n1119 ;
  assign n1121 = ~n1116 & n1119 ;
  assign n1122 = ~n1120 & ~n1121 ;
  assign n1123 = ~n1116 & ~n1117 ;
  assign n1124 = ~n1118 & ~n1123 ;
  assign n1125 = ~x109 & ~x237 ;
  assign n1126 = x109 & x237 ;
  assign n1127 = ~n1125 & ~n1126 ;
  assign n1128 = n1124 & ~n1127 ;
  assign n1129 = ~n1124 & n1127 ;
  assign n1130 = ~n1128 & ~n1129 ;
  assign n1131 = ~n1124 & ~n1125 ;
  assign n1132 = ~n1126 & ~n1131 ;
  assign n1133 = ~x110 & ~x238 ;
  assign n1134 = x110 & x238 ;
  assign n1135 = ~n1133 & ~n1134 ;
  assign n1136 = n1132 & ~n1135 ;
  assign n1137 = ~n1132 & n1135 ;
  assign n1138 = ~n1136 & ~n1137 ;
  assign n1139 = ~n1132 & ~n1133 ;
  assign n1140 = ~n1134 & ~n1139 ;
  assign n1141 = ~x111 & ~x239 ;
  assign n1142 = x111 & x239 ;
  assign n1143 = ~n1141 & ~n1142 ;
  assign n1144 = n1140 & ~n1143 ;
  assign n1145 = ~n1140 & n1143 ;
  assign n1146 = ~n1144 & ~n1145 ;
  assign n1147 = ~n1140 & ~n1141 ;
  assign n1148 = ~n1142 & ~n1147 ;
  assign n1149 = ~x112 & ~x240 ;
  assign n1150 = x112 & x240 ;
  assign n1151 = ~n1149 & ~n1150 ;
  assign n1152 = n1148 & ~n1151 ;
  assign n1153 = ~n1148 & n1151 ;
  assign n1154 = ~n1152 & ~n1153 ;
  assign n1155 = ~n1148 & ~n1149 ;
  assign n1156 = ~n1150 & ~n1155 ;
  assign n1157 = ~x113 & ~x241 ;
  assign n1158 = x113 & x241 ;
  assign n1159 = ~n1157 & ~n1158 ;
  assign n1160 = n1156 & ~n1159 ;
  assign n1161 = ~n1156 & n1159 ;
  assign n1162 = ~n1160 & ~n1161 ;
  assign n1163 = ~n1156 & ~n1157 ;
  assign n1164 = ~n1158 & ~n1163 ;
  assign n1165 = ~x114 & ~x242 ;
  assign n1166 = x114 & x242 ;
  assign n1167 = ~n1165 & ~n1166 ;
  assign n1168 = n1164 & ~n1167 ;
  assign n1169 = ~n1164 & n1167 ;
  assign n1170 = ~n1168 & ~n1169 ;
  assign n1171 = ~n1164 & ~n1165 ;
  assign n1172 = ~n1166 & ~n1171 ;
  assign n1173 = ~x115 & ~x243 ;
  assign n1174 = x115 & x243 ;
  assign n1175 = ~n1173 & ~n1174 ;
  assign n1176 = n1172 & ~n1175 ;
  assign n1177 = ~n1172 & n1175 ;
  assign n1178 = ~n1176 & ~n1177 ;
  assign n1179 = ~n1172 & ~n1173 ;
  assign n1180 = ~n1174 & ~n1179 ;
  assign n1181 = ~x116 & ~x244 ;
  assign n1182 = x116 & x244 ;
  assign n1183 = ~n1181 & ~n1182 ;
  assign n1184 = n1180 & ~n1183 ;
  assign n1185 = ~n1180 & n1183 ;
  assign n1186 = ~n1184 & ~n1185 ;
  assign n1187 = ~n1180 & ~n1181 ;
  assign n1188 = ~n1182 & ~n1187 ;
  assign n1189 = ~x117 & ~x245 ;
  assign n1190 = x117 & x245 ;
  assign n1191 = ~n1189 & ~n1190 ;
  assign n1192 = n1188 & ~n1191 ;
  assign n1193 = ~n1188 & n1191 ;
  assign n1194 = ~n1192 & ~n1193 ;
  assign n1195 = ~n1188 & ~n1189 ;
  assign n1196 = ~n1190 & ~n1195 ;
  assign n1197 = ~x118 & ~x246 ;
  assign n1198 = x118 & x246 ;
  assign n1199 = ~n1197 & ~n1198 ;
  assign n1200 = n1196 & ~n1199 ;
  assign n1201 = ~n1196 & n1199 ;
  assign n1202 = ~n1200 & ~n1201 ;
  assign n1203 = ~n1196 & ~n1197 ;
  assign n1204 = ~n1198 & ~n1203 ;
  assign n1205 = ~x119 & ~x247 ;
  assign n1206 = x119 & x247 ;
  assign n1207 = ~n1205 & ~n1206 ;
  assign n1208 = n1204 & ~n1207 ;
  assign n1209 = ~n1204 & n1207 ;
  assign n1210 = ~n1208 & ~n1209 ;
  assign n1211 = ~n1204 & ~n1205 ;
  assign n1212 = ~n1206 & ~n1211 ;
  assign n1213 = ~x120 & ~x248 ;
  assign n1214 = x120 & x248 ;
  assign n1215 = ~n1213 & ~n1214 ;
  assign n1216 = n1212 & ~n1215 ;
  assign n1217 = ~n1212 & n1215 ;
  assign n1218 = ~n1216 & ~n1217 ;
  assign n1219 = ~n1212 & ~n1213 ;
  assign n1220 = ~n1214 & ~n1219 ;
  assign n1221 = ~x121 & ~x249 ;
  assign n1222 = x121 & x249 ;
  assign n1223 = ~n1221 & ~n1222 ;
  assign n1224 = n1220 & ~n1223 ;
  assign n1225 = ~n1220 & n1223 ;
  assign n1226 = ~n1224 & ~n1225 ;
  assign n1227 = ~n1220 & ~n1221 ;
  assign n1228 = ~n1222 & ~n1227 ;
  assign n1229 = ~x122 & ~x250 ;
  assign n1230 = x122 & x250 ;
  assign n1231 = ~n1229 & ~n1230 ;
  assign n1232 = n1228 & ~n1231 ;
  assign n1233 = ~n1228 & n1231 ;
  assign n1234 = ~n1232 & ~n1233 ;
  assign n1235 = ~n1228 & ~n1229 ;
  assign n1236 = ~n1230 & ~n1235 ;
  assign n1237 = ~x123 & ~x251 ;
  assign n1238 = x123 & x251 ;
  assign n1239 = ~n1237 & ~n1238 ;
  assign n1240 = n1236 & ~n1239 ;
  assign n1241 = ~n1236 & n1239 ;
  assign n1242 = ~n1240 & ~n1241 ;
  assign n1243 = ~n1236 & ~n1237 ;
  assign n1244 = ~n1238 & ~n1243 ;
  assign n1245 = ~x124 & ~x252 ;
  assign n1246 = x124 & x252 ;
  assign n1247 = ~n1245 & ~n1246 ;
  assign n1248 = n1244 & ~n1247 ;
  assign n1249 = ~n1244 & n1247 ;
  assign n1250 = ~n1248 & ~n1249 ;
  assign n1251 = ~n1244 & ~n1245 ;
  assign n1252 = ~n1246 & ~n1251 ;
  assign n1253 = ~x125 & ~x253 ;
  assign n1254 = x125 & x253 ;
  assign n1255 = ~n1253 & ~n1254 ;
  assign n1256 = n1252 & ~n1255 ;
  assign n1257 = ~n1252 & n1255 ;
  assign n1258 = ~n1256 & ~n1257 ;
  assign n1259 = ~n1252 & ~n1253 ;
  assign n1260 = ~n1254 & ~n1259 ;
  assign n1261 = ~x126 & ~x254 ;
  assign n1262 = x126 & x254 ;
  assign n1263 = ~n1261 & ~n1262 ;
  assign n1264 = n1260 & ~n1263 ;
  assign n1265 = ~n1260 & n1263 ;
  assign n1266 = ~n1264 & ~n1265 ;
  assign n1267 = ~n1260 & ~n1261 ;
  assign n1268 = ~n1262 & ~n1267 ;
  assign n1269 = ~x127 & ~x255 ;
  assign n1270 = x127 & x255 ;
  assign n1271 = ~n1269 & ~n1270 ;
  assign n1272 = n1268 & ~n1271 ;
  assign n1273 = ~n1268 & n1271 ;
  assign n1274 = ~n1272 & ~n1273 ;
  assign n1275 = ~n1268 & ~n1269 ;
  assign n1276 = ~n1270 & ~n1275 ;
  assign y0 = ~n259 ;
  assign y1 = ~n266 ;
  assign y2 = n274 ;
  assign y3 = n282 ;
  assign y4 = n290 ;
  assign y5 = n298 ;
  assign y6 = n306 ;
  assign y7 = n314 ;
  assign y8 = n322 ;
  assign y9 = n330 ;
  assign y10 = n338 ;
  assign y11 = n346 ;
  assign y12 = n354 ;
  assign y13 = n362 ;
  assign y14 = n370 ;
  assign y15 = n378 ;
  assign y16 = n386 ;
  assign y17 = n394 ;
  assign y18 = n402 ;
  assign y19 = n410 ;
  assign y20 = n418 ;
  assign y21 = n426 ;
  assign y22 = n434 ;
  assign y23 = n442 ;
  assign y24 = n450 ;
  assign y25 = n458 ;
  assign y26 = n466 ;
  assign y27 = n474 ;
  assign y28 = n482 ;
  assign y29 = n490 ;
  assign y30 = n498 ;
  assign y31 = n506 ;
  assign y32 = n514 ;
  assign y33 = n522 ;
  assign y34 = n530 ;
  assign y35 = n538 ;
  assign y36 = n546 ;
  assign y37 = n554 ;
  assign y38 = n562 ;
  assign y39 = n570 ;
  assign y40 = n578 ;
  assign y41 = n586 ;
  assign y42 = n594 ;
  assign y43 = n602 ;
  assign y44 = n610 ;
  assign y45 = n618 ;
  assign y46 = n626 ;
  assign y47 = n634 ;
  assign y48 = n642 ;
  assign y49 = n650 ;
  assign y50 = n658 ;
  assign y51 = n666 ;
  assign y52 = n674 ;
  assign y53 = n682 ;
  assign y54 = n690 ;
  assign y55 = n698 ;
  assign y56 = n706 ;
  assign y57 = n714 ;
  assign y58 = n722 ;
  assign y59 = n730 ;
  assign y60 = n738 ;
  assign y61 = n746 ;
  assign y62 = n754 ;
  assign y63 = n762 ;
  assign y64 = n770 ;
  assign y65 = n778 ;
  assign y66 = n786 ;
  assign y67 = n794 ;
  assign y68 = n802 ;
  assign y69 = n810 ;
  assign y70 = n818 ;
  assign y71 = n826 ;
  assign y72 = n834 ;
  assign y73 = n842 ;
  assign y74 = n850 ;
  assign y75 = n858 ;
  assign y76 = n866 ;
  assign y77 = n874 ;
  assign y78 = n882 ;
  assign y79 = n890 ;
  assign y80 = n898 ;
  assign y81 = n906 ;
  assign y82 = n914 ;
  assign y83 = n922 ;
  assign y84 = n930 ;
  assign y85 = n938 ;
  assign y86 = n946 ;
  assign y87 = n954 ;
  assign y88 = n962 ;
  assign y89 = n970 ;
  assign y90 = n978 ;
  assign y91 = n986 ;
  assign y92 = n994 ;
  assign y93 = n1002 ;
  assign y94 = n1010 ;
  assign y95 = n1018 ;
  assign y96 = n1026 ;
  assign y97 = n1034 ;
  assign y98 = n1042 ;
  assign y99 = n1050 ;
  assign y100 = n1058 ;
  assign y101 = n1066 ;
  assign y102 = n1074 ;
  assign y103 = n1082 ;
  assign y104 = n1090 ;
  assign y105 = n1098 ;
  assign y106 = n1106 ;
  assign y107 = n1114 ;
  assign y108 = n1122 ;
  assign y109 = n1130 ;
  assign y110 = n1138 ;
  assign y111 = n1146 ;
  assign y112 = n1154 ;
  assign y113 = n1162 ;
  assign y114 = n1170 ;
  assign y115 = n1178 ;
  assign y116 = n1186 ;
  assign y117 = n1194 ;
  assign y118 = n1202 ;
  assign y119 = n1210 ;
  assign y120 = n1218 ;
  assign y121 = n1226 ;
  assign y122 = n1234 ;
  assign y123 = n1242 ;
  assign y124 = n1250 ;
  assign y125 = n1258 ;
  assign y126 = n1266 ;
  assign y127 = n1274 ;
  assign y128 = ~n1276 ;
endmodule
