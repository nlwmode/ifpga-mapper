module top( \G0_pad  , \G10_reg/NET0131  , \G11_reg/NET0131  , \G12_reg/NET0131  , \G13_reg/NET0131  , \G147_pad  , \G148_pad  , \G14_reg/NET0131  , \G15_reg/NET0131  , \G16_reg/NET0131  , \G17_reg/NET0131  , \G18_reg/NET0131  , \G198_pad  , \G199_pad  , \G19_reg/NET0131  , \G1_pad  , \G20_reg/NET0131  , \G213_pad  , \G214_pad  , \G21_reg/NET0131  , \G22_reg/NET0131  , \G29_reg/NET0131  , \G2_pad  , \G30_reg/NET0131  , \_al_n0  , \_al_n1  , \g1001/_0_  , \g1003/_0_  , \g1008/_0_  , \g1014/_0_  , \g1031/_0_  , \g1051/_0_  , \g1066/_0_  , \g1067/_0_  , \g1148/_0_  , \g1278/_0_  , \g1306/_3_  , \g1318/_2_  , \g1323/_3_  , \g1400/_0_  , \g1427/_2_  , \g1451/_0_  , \g22/_0_  , \g979/_0_  , \g982/_0_  , \g992/_0_  , \g995/_0_  );
  input \G0_pad  ;
  input \G10_reg/NET0131  ;
  input \G11_reg/NET0131  ;
  input \G12_reg/NET0131  ;
  input \G13_reg/NET0131  ;
  input \G147_pad  ;
  input \G148_pad  ;
  input \G14_reg/NET0131  ;
  input \G15_reg/NET0131  ;
  input \G16_reg/NET0131  ;
  input \G17_reg/NET0131  ;
  input \G18_reg/NET0131  ;
  input \G198_pad  ;
  input \G199_pad  ;
  input \G19_reg/NET0131  ;
  input \G1_pad  ;
  input \G20_reg/NET0131  ;
  input \G213_pad  ;
  input \G214_pad  ;
  input \G21_reg/NET0131  ;
  input \G22_reg/NET0131  ;
  input \G29_reg/NET0131  ;
  input \G2_pad  ;
  input \G30_reg/NET0131  ;
  output \_al_n0  ;
  output \_al_n1  ;
  output \g1001/_0_  ;
  output \g1003/_0_  ;
  output \g1008/_0_  ;
  output \g1014/_0_  ;
  output \g1031/_0_  ;
  output \g1051/_0_  ;
  output \g1066/_0_  ;
  output \g1067/_0_  ;
  output \g1148/_0_  ;
  output \g1278/_0_  ;
  output \g1306/_3_  ;
  output \g1318/_2_  ;
  output \g1323/_3_  ;
  output \g1400/_0_  ;
  output \g1427/_2_  ;
  output \g1451/_0_  ;
  output \g22/_0_  ;
  output \g979/_0_  ;
  output \g982/_0_  ;
  output \g992/_0_  ;
  output \g995/_0_  ;
  wire n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 ;
  assign n25 = ~\G14_reg/NET0131  & \G15_reg/NET0131  ;
  assign n26 = \G10_reg/NET0131  & ~\G11_reg/NET0131  ;
  assign n27 = n25 & n26 ;
  assign n28 = ~\G30_reg/NET0131  & ~n27 ;
  assign n29 = ~\G17_reg/NET0131  & ~\G18_reg/NET0131  ;
  assign n30 = \G16_reg/NET0131  & \G19_reg/NET0131  ;
  assign n31 = n29 & n30 ;
  assign n32 = ~n28 & n31 ;
  assign n33 = ~\G20_reg/NET0131  & ~n32 ;
  assign n34 = \G20_reg/NET0131  & n31 ;
  assign n35 = ~n28 & n34 ;
  assign n36 = ~\G0_pad  & ~n35 ;
  assign n37 = ~n33 & n36 ;
  assign n39 = \G20_reg/NET0131  & ~\G21_reg/NET0131  ;
  assign n38 = \G12_reg/NET0131  & ~\G13_reg/NET0131  ;
  assign n40 = ~\G29_reg/NET0131  & n38 ;
  assign n41 = n39 & n40 ;
  assign n42 = \G22_reg/NET0131  & ~n41 ;
  assign n43 = ~\G20_reg/NET0131  & ~\G21_reg/NET0131  ;
  assign n44 = \G29_reg/NET0131  & n38 ;
  assign n45 = n43 & n44 ;
  assign n46 = ~n42 & ~n45 ;
  assign n47 = ~\G0_pad  & ~n46 ;
  assign n49 = ~\G16_reg/NET0131  & n28 ;
  assign n48 = \G16_reg/NET0131  & ~n28 ;
  assign n50 = ~\G0_pad  & ~n48 ;
  assign n51 = ~n49 & n50 ;
  assign n52 = \G10_reg/NET0131  & \G11_reg/NET0131  ;
  assign n54 = ~\G14_reg/NET0131  & ~n52 ;
  assign n53 = \G14_reg/NET0131  & n52 ;
  assign n55 = ~\G0_pad  & ~n53 ;
  assign n56 = ~n54 & n55 ;
  assign n59 = \G15_reg/NET0131  & n53 ;
  assign n58 = ~\G15_reg/NET0131  & ~n53 ;
  assign n57 = ~\G14_reg/NET0131  & n26 ;
  assign n60 = ~\G0_pad  & ~n57 ;
  assign n61 = ~n58 & n60 ;
  assign n62 = ~n59 & n61 ;
  assign n63 = \G10_reg/NET0131  & ~n25 ;
  assign n64 = ~\G11_reg/NET0131  & ~n63 ;
  assign n65 = ~\G0_pad  & ~n52 ;
  assign n66 = ~n64 & n65 ;
  assign n67 = \G29_reg/NET0131  & ~\G2_pad  ;
  assign n68 = ~\G29_reg/NET0131  & \G2_pad  ;
  assign n69 = ~n67 & ~n68 ;
  assign n70 = ~\G0_pad  & ~n69 ;
  assign n71 = \G1_pad  & ~\G30_reg/NET0131  ;
  assign n72 = ~\G1_pad  & \G30_reg/NET0131  ;
  assign n73 = ~n71 & ~n72 ;
  assign n74 = ~\G0_pad  & ~n73 ;
  assign n75 = ~\G0_pad  & ~\G10_reg/NET0131  ;
  assign n76 = \G18_reg/NET0131  & ~n46 ;
  assign n77 = ~\G12_reg/NET0131  & ~\G21_reg/NET0131  ;
  assign n79 = \G20_reg/NET0131  & n77 ;
  assign n78 = ~\G213_pad  & ~n77 ;
  assign n80 = \G13_reg/NET0131  & ~n78 ;
  assign n81 = ~n79 & n80 ;
  assign n82 = n46 & ~n81 ;
  assign n83 = ~n76 & ~n82 ;
  assign n84 = \G13_reg/NET0131  & \G21_reg/NET0131  ;
  assign n85 = ~\G12_reg/NET0131  & ~n84 ;
  assign n86 = ~\G198_pad  & ~n85 ;
  assign n87 = \G12_reg/NET0131  & \G13_reg/NET0131  ;
  assign n88 = \G13_reg/NET0131  & n43 ;
  assign n89 = ~\G12_reg/NET0131  & ~n88 ;
  assign n90 = ~n87 & ~n89 ;
  assign n91 = n46 & ~n90 ;
  assign n92 = ~n86 & n91 ;
  assign n93 = ~\G13_reg/NET0131  & \G20_reg/NET0131  ;
  assign n94 = \G13_reg/NET0131  & \G214_pad  ;
  assign n95 = ~n93 & ~n94 ;
  assign n96 = ~n38 & ~n77 ;
  assign n97 = ~n95 & n96 ;
  assign n98 = n46 & n97 ;
  assign n99 = ~\G148_pad  & ~n85 ;
  assign n100 = \G21_reg/NET0131  & n93 ;
  assign n101 = ~n99 & ~n100 ;
  assign n102 = n91 & n101 ;
  assign n103 = ~\G0_pad  & \G19_reg/NET0131  ;
  assign n104 = \G17_reg/NET0131  & \G18_reg/NET0131  ;
  assign n105 = ~\G0_pad  & n104 ;
  assign n106 = n48 & n105 ;
  assign n107 = ~n103 & ~n106 ;
  assign n108 = ~n29 & ~n104 ;
  assign n109 = n48 & ~n108 ;
  assign n110 = \G19_reg/NET0131  & n109 ;
  assign n111 = ~n107 & ~n110 ;
  assign n112 = \G199_pad  & n84 ;
  assign n113 = ~\G199_pad  & n87 ;
  assign n114 = ~n89 & ~n113 ;
  assign n115 = ~n112 & ~n114 ;
  assign n116 = n46 & n115 ;
  assign n117 = ~n76 & ~n116 ;
  assign n121 = ~\G17_reg/NET0131  & ~n48 ;
  assign n118 = ~\G18_reg/NET0131  & \G19_reg/NET0131  ;
  assign n119 = ~\G17_reg/NET0131  & ~n118 ;
  assign n120 = n48 & ~n119 ;
  assign n122 = ~\G0_pad  & ~n120 ;
  assign n123 = ~n121 & n122 ;
  assign n124 = \G13_reg/NET0131  & ~\G147_pad  ;
  assign n125 = ~n85 & ~n124 ;
  assign n126 = n46 & n125 ;
  assign n127 = \G21_reg/NET0131  & n36 ;
  assign n128 = ~\G12_reg/NET0131  & \G13_reg/NET0131  ;
  assign n129 = ~\G0_pad  & n39 ;
  assign n130 = ~n128 & n129 ;
  assign n131 = n32 & n130 ;
  assign n132 = ~n127 & ~n131 ;
  assign n133 = \G21_reg/NET0131  & n35 ;
  assign n134 = ~\G0_pad  & \G12_reg/NET0131  ;
  assign n135 = ~n133 & n134 ;
  assign n136 = ~\G0_pad  & ~\G12_reg/NET0131  ;
  assign n137 = n133 & n136 ;
  assign n138 = ~n135 & ~n137 ;
  assign n139 = \G12_reg/NET0131  & \G21_reg/NET0131  ;
  assign n140 = ~n77 & ~n139 ;
  assign n141 = n35 & ~n140 ;
  assign n142 = ~\G0_pad  & \G13_reg/NET0131  ;
  assign n143 = ~n141 & n142 ;
  assign n144 = ~\G13_reg/NET0131  & n134 ;
  assign n145 = n133 & n144 ;
  assign n146 = ~n143 & ~n145 ;
  assign n147 = ~\G18_reg/NET0131  & ~n48 ;
  assign n148 = ~\G0_pad  & ~n109 ;
  assign n149 = ~n147 & n148 ;
  assign \_al_n0  = 1'b0 ;
  assign \_al_n1  = ~1'b0 ;
  assign \g1001/_0_  = n37 ;
  assign \g1003/_0_  = n47 ;
  assign \g1008/_0_  = n51 ;
  assign \g1014/_0_  = n56 ;
  assign \g1031/_0_  = n62 ;
  assign \g1051/_0_  = n66 ;
  assign \g1066/_0_  = n70 ;
  assign \g1067/_0_  = n74 ;
  assign \g1148/_0_  = n75 ;
  assign \g1278/_0_  = n83 ;
  assign \g1306/_3_  = n92 ;
  assign \g1318/_2_  = n98 ;
  assign \g1323/_3_  = n102 ;
  assign \g1400/_0_  = n111 ;
  assign \g1427/_2_  = n117 ;
  assign \g1451/_0_  = n123 ;
  assign \g22/_0_  = n126 ;
  assign \g979/_0_  = ~n132 ;
  assign \g982/_0_  = ~n138 ;
  assign \g992/_0_  = ~n146 ;
  assign \g995/_0_  = n149 ;
endmodule
