module top (\1_pad , \2_pad , \3_pad , \4_pad , \5_pad , \6_pad , \7_pad , \8_pad , \44_pad , \45_pad , \46_pad , \47_pad , \48_pad , \49_pad , \50_pad , \51_pad );
	input \1_pad  ;
	input \2_pad  ;
	input \3_pad  ;
	input \4_pad  ;
	input \5_pad  ;
	input \6_pad  ;
	input \7_pad  ;
	input \8_pad  ;
	output \44_pad  ;
	output \45_pad  ;
	output \46_pad  ;
	output \47_pad  ;
	output \48_pad  ;
	output \49_pad  ;
	output \50_pad  ;
	output \51_pad  ;
	wire _w134_ ;
	wire _w133_ ;
	wire _w132_ ;
	wire _w131_ ;
	wire _w130_ ;
	wire _w129_ ;
	wire _w128_ ;
	wire _w127_ ;
	wire _w126_ ;
	wire _w125_ ;
	wire _w124_ ;
	wire _w123_ ;
	wire _w122_ ;
	wire _w121_ ;
	wire _w120_ ;
	wire _w119_ ;
	wire _w118_ ;
	wire _w117_ ;
	wire _w116_ ;
	wire _w115_ ;
	wire _w114_ ;
	wire _w113_ ;
	wire _w112_ ;
	wire _w111_ ;
	wire _w110_ ;
	wire _w109_ ;
	wire _w108_ ;
	wire _w107_ ;
	wire _w106_ ;
	wire _w105_ ;
	wire _w104_ ;
	wire _w103_ ;
	wire _w102_ ;
	wire _w101_ ;
	wire _w100_ ;
	wire _w99_ ;
	wire _w98_ ;
	wire _w97_ ;
	wire _w96_ ;
	wire _w95_ ;
	wire _w94_ ;
	wire _w93_ ;
	wire _w92_ ;
	wire _w91_ ;
	wire _w90_ ;
	wire _w89_ ;
	wire _w88_ ;
	wire _w87_ ;
	wire _w86_ ;
	wire _w85_ ;
	wire _w84_ ;
	wire _w83_ ;
	wire _w82_ ;
	wire _w81_ ;
	wire _w80_ ;
	wire _w79_ ;
	wire _w78_ ;
	wire _w77_ ;
	wire _w76_ ;
	wire _w75_ ;
	wire _w74_ ;
	wire _w73_ ;
	wire _w72_ ;
	wire _w71_ ;
	wire _w70_ ;
	wire _w69_ ;
	wire _w68_ ;
	wire _w37_ ;
	wire _w36_ ;
	wire _w35_ ;
	wire _w34_ ;
	wire _w33_ ;
	wire _w32_ ;
	wire _w31_ ;
	wire _w30_ ;
	wire _w29_ ;
	wire _w28_ ;
	wire _w27_ ;
	wire _w26_ ;
	wire _w25_ ;
	wire _w24_ ;
	wire _w23_ ;
	wire _w22_ ;
	wire _w9_ ;
	wire _w10_ ;
	wire _w11_ ;
	wire _w12_ ;
	wire _w13_ ;
	wire _w14_ ;
	wire _w15_ ;
	wire _w16_ ;
	wire _w17_ ;
	wire _w18_ ;
	wire _w19_ ;
	wire _w20_ ;
	wire _w21_ ;
	wire _w38_ ;
	wire _w39_ ;
	wire _w40_ ;
	wire _w41_ ;
	wire _w42_ ;
	wire _w43_ ;
	wire _w44_ ;
	wire _w45_ ;
	wire _w46_ ;
	wire _w47_ ;
	wire _w48_ ;
	wire _w49_ ;
	wire _w50_ ;
	wire _w51_ ;
	wire _w52_ ;
	wire _w53_ ;
	wire _w54_ ;
	wire _w55_ ;
	wire _w56_ ;
	wire _w57_ ;
	wire _w58_ ;
	wire _w59_ ;
	wire _w60_ ;
	wire _w61_ ;
	wire _w62_ ;
	wire _w63_ ;
	wire _w64_ ;
	wire _w65_ ;
	wire _w66_ ;
	wire _w67_ ;
	LUT2 #(
		.INIT('h8)
	) name0 (
		\7_pad ,
		\8_pad ,
		_w9_
	);
	LUT2 #(
		.INIT('h4)
	) name1 (
		\1_pad ,
		\3_pad ,
		_w10_
	);
	LUT2 #(
		.INIT('h2)
	) name2 (
		\1_pad ,
		\3_pad ,
		_w11_
	);
	LUT2 #(
		.INIT('h1)
	) name3 (
		_w10_,
		_w11_,
		_w12_
	);
	LUT2 #(
		.INIT('h1)
	) name4 (
		\4_pad ,
		_w12_,
		_w13_
	);
	LUT2 #(
		.INIT('h2)
	) name5 (
		_w9_,
		_w13_,
		_w14_
	);
	LUT2 #(
		.INIT('h1)
	) name6 (
		\6_pad ,
		_w14_,
		_w15_
	);
	LUT2 #(
		.INIT('h1)
	) name7 (
		_w9_,
		_w13_,
		_w16_
	);
	LUT2 #(
		.INIT('h1)
	) name8 (
		\1_pad ,
		\2_pad ,
		_w17_
	);
	LUT2 #(
		.INIT('h8)
	) name9 (
		\1_pad ,
		\2_pad ,
		_w18_
	);
	LUT2 #(
		.INIT('h1)
	) name10 (
		_w17_,
		_w18_,
		_w19_
	);
	LUT2 #(
		.INIT('h8)
	) name11 (
		\3_pad ,
		_w19_,
		_w20_
	);
	LUT2 #(
		.INIT('h1)
	) name12 (
		\1_pad ,
		\3_pad ,
		_w21_
	);
	LUT2 #(
		.INIT('h1)
	) name13 (
		\4_pad ,
		_w21_,
		_w22_
	);
	LUT2 #(
		.INIT('h4)
	) name14 (
		_w20_,
		_w22_,
		_w23_
	);
	LUT2 #(
		.INIT('h8)
	) name15 (
		\6_pad ,
		_w23_,
		_w24_
	);
	LUT2 #(
		.INIT('h2)
	) name16 (
		_w9_,
		_w24_,
		_w25_
	);
	LUT2 #(
		.INIT('h1)
	) name17 (
		_w16_,
		_w25_,
		_w26_
	);
	LUT2 #(
		.INIT('h1)
	) name18 (
		\3_pad ,
		_w19_,
		_w27_
	);
	LUT2 #(
		.INIT('h2)
	) name19 (
		\4_pad ,
		_w10_,
		_w28_
	);
	LUT2 #(
		.INIT('h4)
	) name20 (
		_w27_,
		_w28_,
		_w29_
	);
	LUT2 #(
		.INIT('h1)
	) name21 (
		_w15_,
		_w29_,
		_w30_
	);
	LUT2 #(
		.INIT('h4)
	) name22 (
		_w26_,
		_w30_,
		_w31_
	);
	LUT2 #(
		.INIT('h1)
	) name23 (
		_w20_,
		_w27_,
		_w32_
	);
	LUT2 #(
		.INIT('h8)
	) name24 (
		\4_pad ,
		_w32_,
		_w33_
	);
	LUT2 #(
		.INIT('h4)
	) name25 (
		\6_pad ,
		_w16_,
		_w34_
	);
	LUT2 #(
		.INIT('h4)
	) name26 (
		_w33_,
		_w34_,
		_w35_
	);
	LUT2 #(
		.INIT('h1)
	) name27 (
		_w31_,
		_w35_,
		_w36_
	);
	LUT2 #(
		.INIT('h1)
	) name28 (
		\5_pad ,
		_w36_,
		_w37_
	);
	LUT2 #(
		.INIT('h8)
	) name29 (
		\4_pad ,
		_w12_,
		_w38_
	);
	LUT2 #(
		.INIT('h1)
	) name30 (
		\7_pad ,
		_w23_,
		_w39_
	);
	LUT2 #(
		.INIT('h1)
	) name31 (
		\8_pad ,
		_w39_,
		_w40_
	);
	LUT2 #(
		.INIT('h4)
	) name32 (
		\4_pad ,
		_w32_,
		_w41_
	);
	LUT2 #(
		.INIT('h8)
	) name33 (
		\8_pad ,
		_w41_,
		_w42_
	);
	LUT2 #(
		.INIT('h2)
	) name34 (
		\6_pad ,
		_w40_,
		_w43_
	);
	LUT2 #(
		.INIT('h4)
	) name35 (
		_w42_,
		_w43_,
		_w44_
	);
	LUT2 #(
		.INIT('h4)
	) name36 (
		\6_pad ,
		_w23_,
		_w45_
	);
	LUT2 #(
		.INIT('h8)
	) name37 (
		\6_pad ,
		_w41_,
		_w46_
	);
	LUT2 #(
		.INIT('h2)
	) name38 (
		\7_pad ,
		_w45_,
		_w47_
	);
	LUT2 #(
		.INIT('h4)
	) name39 (
		_w46_,
		_w47_,
		_w48_
	);
	LUT2 #(
		.INIT('h1)
	) name40 (
		_w44_,
		_w48_,
		_w49_
	);
	LUT2 #(
		.INIT('h1)
	) name41 (
		_w38_,
		_w49_,
		_w50_
	);
	LUT2 #(
		.INIT('h1)
	) name42 (
		\6_pad ,
		_w29_,
		_w51_
	);
	LUT2 #(
		.INIT('h8)
	) name43 (
		_w39_,
		_w51_,
		_w52_
	);
	LUT2 #(
		.INIT('h1)
	) name44 (
		_w50_,
		_w52_,
		_w53_
	);
	LUT2 #(
		.INIT('h2)
	) name45 (
		\5_pad ,
		_w53_,
		_w54_
	);
	LUT2 #(
		.INIT('h1)
	) name46 (
		_w37_,
		_w54_,
		_w55_
	);
	LUT2 #(
		.INIT('h1)
	) name47 (
		\3_pad ,
		\5_pad ,
		_w56_
	);
	LUT2 #(
		.INIT('h8)
	) name48 (
		\3_pad ,
		\5_pad ,
		_w57_
	);
	LUT2 #(
		.INIT('h1)
	) name49 (
		\6_pad ,
		_w57_,
		_w58_
	);
	LUT2 #(
		.INIT('h1)
	) name50 (
		_w56_,
		_w58_,
		_w59_
	);
	LUT2 #(
		.INIT('h8)
	) name51 (
		\3_pad ,
		\8_pad ,
		_w60_
	);
	LUT2 #(
		.INIT('h1)
	) name52 (
		\5_pad ,
		_w60_,
		_w61_
	);
	LUT2 #(
		.INIT('h2)
	) name53 (
		\7_pad ,
		_w61_,
		_w62_
	);
	LUT2 #(
		.INIT('h2)
	) name54 (
		\2_pad ,
		_w62_,
		_w63_
	);
	LUT2 #(
		.INIT('h2)
	) name55 (
		\4_pad ,
		_w63_,
		_w64_
	);
	LUT2 #(
		.INIT('h2)
	) name56 (
		\2_pad ,
		\4_pad ,
		_w65_
	);
	LUT2 #(
		.INIT('h1)
	) name57 (
		_w59_,
		_w65_,
		_w66_
	);
	LUT2 #(
		.INIT('h4)
	) name58 (
		_w64_,
		_w66_,
		_w67_
	);
	LUT2 #(
		.INIT('h1)
	) name59 (
		_w57_,
		_w62_,
		_w68_
	);
	LUT2 #(
		.INIT('h2)
	) name60 (
		\4_pad ,
		_w68_,
		_w69_
	);
	LUT2 #(
		.INIT('h8)
	) name61 (
		\4_pad ,
		\5_pad ,
		_w70_
	);
	LUT2 #(
		.INIT('h2)
	) name62 (
		\3_pad ,
		\5_pad ,
		_w71_
	);
	LUT2 #(
		.INIT('h4)
	) name63 (
		\7_pad ,
		_w71_,
		_w72_
	);
	LUT2 #(
		.INIT('h4)
	) name64 (
		\3_pad ,
		\7_pad ,
		_w73_
	);
	LUT2 #(
		.INIT('h1)
	) name65 (
		\8_pad ,
		_w56_,
		_w74_
	);
	LUT2 #(
		.INIT('h1)
	) name66 (
		_w57_,
		_w73_,
		_w75_
	);
	LUT2 #(
		.INIT('h8)
	) name67 (
		_w74_,
		_w75_,
		_w76_
	);
	LUT2 #(
		.INIT('h1)
	) name68 (
		_w70_,
		_w72_,
		_w77_
	);
	LUT2 #(
		.INIT('h4)
	) name69 (
		_w76_,
		_w77_,
		_w78_
	);
	LUT2 #(
		.INIT('h2)
	) name70 (
		\6_pad ,
		_w78_,
		_w79_
	);
	LUT2 #(
		.INIT('h1)
	) name71 (
		_w69_,
		_w79_,
		_w80_
	);
	LUT2 #(
		.INIT('h1)
	) name72 (
		\2_pad ,
		_w80_,
		_w81_
	);
	LUT2 #(
		.INIT('h1)
	) name73 (
		\3_pad ,
		\8_pad ,
		_w82_
	);
	LUT2 #(
		.INIT('h2)
	) name74 (
		\5_pad ,
		_w82_,
		_w83_
	);
	LUT2 #(
		.INIT('h1)
	) name75 (
		_w62_,
		_w83_,
		_w84_
	);
	LUT2 #(
		.INIT('h4)
	) name76 (
		_w58_,
		_w65_,
		_w85_
	);
	LUT2 #(
		.INIT('h4)
	) name77 (
		_w84_,
		_w85_,
		_w86_
	);
	LUT2 #(
		.INIT('h1)
	) name78 (
		_w67_,
		_w86_,
		_w87_
	);
	LUT2 #(
		.INIT('h4)
	) name79 (
		_w81_,
		_w87_,
		_w88_
	);
	LUT2 #(
		.INIT('h1)
	) name80 (
		\4_pad ,
		\8_pad ,
		_w89_
	);
	LUT2 #(
		.INIT('h2)
	) name81 (
		\6_pad ,
		_w89_,
		_w90_
	);
	LUT2 #(
		.INIT('h8)
	) name82 (
		\4_pad ,
		_w9_,
		_w91_
	);
	LUT2 #(
		.INIT('h2)
	) name83 (
		_w56_,
		_w91_,
		_w92_
	);
	LUT2 #(
		.INIT('h1)
	) name84 (
		\4_pad ,
		\6_pad ,
		_w93_
	);
	LUT2 #(
		.INIT('h2)
	) name85 (
		\7_pad ,
		_w93_,
		_w94_
	);
	LUT2 #(
		.INIT('h2)
	) name86 (
		_w57_,
		_w94_,
		_w95_
	);
	LUT2 #(
		.INIT('h1)
	) name87 (
		_w92_,
		_w95_,
		_w96_
	);
	LUT2 #(
		.INIT('h1)
	) name88 (
		_w90_,
		_w96_,
		_w97_
	);
	LUT2 #(
		.INIT('h4)
	) name89 (
		\7_pad ,
		\8_pad ,
		_w98_
	);
	LUT2 #(
		.INIT('h4)
	) name90 (
		\4_pad ,
		_w98_,
		_w99_
	);
	LUT2 #(
		.INIT('h1)
	) name91 (
		_w70_,
		_w99_,
		_w100_
	);
	LUT2 #(
		.INIT('h1)
	) name92 (
		\3_pad ,
		_w100_,
		_w101_
	);
	LUT2 #(
		.INIT('h8)
	) name93 (
		\4_pad ,
		_w71_,
		_w102_
	);
	LUT2 #(
		.INIT('h1)
	) name94 (
		_w101_,
		_w102_,
		_w103_
	);
	LUT2 #(
		.INIT('h2)
	) name95 (
		\6_pad ,
		_w103_,
		_w104_
	);
	LUT2 #(
		.INIT('h1)
	) name96 (
		_w57_,
		_w93_,
		_w105_
	);
	LUT2 #(
		.INIT('h8)
	) name97 (
		_w62_,
		_w105_,
		_w106_
	);
	LUT2 #(
		.INIT('h1)
	) name98 (
		_w97_,
		_w106_,
		_w107_
	);
	LUT2 #(
		.INIT('h4)
	) name99 (
		_w104_,
		_w107_,
		_w108_
	);
	LUT2 #(
		.INIT('h8)
	) name100 (
		\4_pad ,
		\6_pad ,
		_w109_
	);
	LUT2 #(
		.INIT('h1)
	) name101 (
		\7_pad ,
		_w93_,
		_w110_
	);
	LUT2 #(
		.INIT('h4)
	) name102 (
		_w109_,
		_w110_,
		_w111_
	);
	LUT2 #(
		.INIT('h1)
	) name103 (
		\4_pad ,
		\5_pad ,
		_w112_
	);
	LUT2 #(
		.INIT('h1)
	) name104 (
		_w70_,
		_w112_,
		_w113_
	);
	LUT2 #(
		.INIT('h8)
	) name105 (
		\6_pad ,
		_w113_,
		_w114_
	);
	LUT2 #(
		.INIT('h1)
	) name106 (
		\6_pad ,
		_w113_,
		_w115_
	);
	LUT2 #(
		.INIT('h2)
	) name107 (
		\7_pad ,
		_w114_,
		_w116_
	);
	LUT2 #(
		.INIT('h4)
	) name108 (
		_w115_,
		_w116_,
		_w117_
	);
	LUT2 #(
		.INIT('h1)
	) name109 (
		_w111_,
		_w117_,
		_w118_
	);
	LUT2 #(
		.INIT('h1)
	) name110 (
		\8_pad ,
		_w118_,
		_w119_
	);
	LUT2 #(
		.INIT('h1)
	) name111 (
		_w93_,
		_w109_,
		_w120_
	);
	LUT2 #(
		.INIT('h2)
	) name112 (
		\7_pad ,
		_w120_,
		_w121_
	);
	LUT2 #(
		.INIT('h2)
	) name113 (
		_w110_,
		_w114_,
		_w122_
	);
	LUT2 #(
		.INIT('h1)
	) name114 (
		_w121_,
		_w122_,
		_w123_
	);
	LUT2 #(
		.INIT('h2)
	) name115 (
		\8_pad ,
		_w123_,
		_w124_
	);
	LUT2 #(
		.INIT('h1)
	) name116 (
		_w119_,
		_w124_,
		_w125_
	);
	LUT2 #(
		.INIT('h2)
	) name117 (
		\7_pad ,
		\8_pad ,
		_w126_
	);
	LUT2 #(
		.INIT('h8)
	) name118 (
		\6_pad ,
		_w98_,
		_w127_
	);
	LUT2 #(
		.INIT('h1)
	) name119 (
		_w126_,
		_w127_,
		_w128_
	);
	LUT2 #(
		.INIT('h2)
	) name120 (
		\5_pad ,
		_w128_,
		_w129_
	);
	LUT2 #(
		.INIT('h4)
	) name121 (
		\5_pad ,
		_w128_,
		_w130_
	);
	LUT2 #(
		.INIT('h1)
	) name122 (
		_w129_,
		_w130_,
		_w131_
	);
	LUT2 #(
		.INIT('h1)
	) name123 (
		\6_pad ,
		_w98_,
		_w132_
	);
	LUT2 #(
		.INIT('h1)
	) name124 (
		_w127_,
		_w132_,
		_w133_
	);
	LUT2 #(
		.INIT('h1)
	) name125 (
		_w98_,
		_w126_,
		_w134_
	);
	assign \44_pad  = _w55_ ;
	assign \45_pad  = _w88_ ;
	assign \46_pad  = _w108_ ;
	assign \47_pad  = _w125_ ;
	assign \48_pad  = _w131_ ;
	assign \49_pad  = _w133_ ;
	assign \50_pad  = _w134_ ;
	assign \51_pad  = \8_pad ;
endmodule;