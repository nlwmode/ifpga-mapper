module top (\a0_pad , a_pad, \b0_pad , \c0_pad , c_pad, \d0_pad , d_pad, \e0_pad , e_pad, \f0_pad , f_pad, \g0_pad , g_pad, \h0_pad , h_pad, \i0_pad , i_pad, \j0_pad , j_pad, \k0_pad , k_pad, \l0_pad , l_pad, \m0_pad , m_pad, \n0_pad , n_pad, \o0_pad , o_pad, \p0_pad , p_pad, \q0_pad , q_pad, \r0_pad , r_pad, \s0_pad , s_pad, \t0_pad , t_pad, \u0_pad , u_pad, \v0_pad , v_pad, w_pad, x_pad, y_pad, z_pad, \a1_pad , \a2_pad , \b1_pad , \b2_pad , \c1_pad , \c2_pad , \d1_pad , \d2_pad , \e1_pad , \e2_pad , \f1_pad , \f2_pad , \g1_pad , \h1_pad , \i1_pad , \j1_pad , \k1_pad , \l1_pad , \m1_pad , \n1_pad , \o1_pad , \p1_pad , \q1_pad , \r1_pad , \s1_pad , \t1_pad , \u1_pad , \v1_pad , \w0_pad , \w1_pad , \x0_pad , \x1_pad , \y0_pad , \y1_pad , \z0_pad , \z1_pad );
	input \a0_pad  ;
	input a_pad ;
	input \b0_pad  ;
	input \c0_pad  ;
	input c_pad ;
	input \d0_pad  ;
	input d_pad ;
	input \e0_pad  ;
	input e_pad ;
	input \f0_pad  ;
	input f_pad ;
	input \g0_pad  ;
	input g_pad ;
	input \h0_pad  ;
	input h_pad ;
	input \i0_pad  ;
	input i_pad ;
	input \j0_pad  ;
	input j_pad ;
	input \k0_pad  ;
	input k_pad ;
	input \l0_pad  ;
	input l_pad ;
	input \m0_pad  ;
	input m_pad ;
	input \n0_pad  ;
	input n_pad ;
	input \o0_pad  ;
	input o_pad ;
	input \p0_pad  ;
	input p_pad ;
	input \q0_pad  ;
	input q_pad ;
	input \r0_pad  ;
	input r_pad ;
	input \s0_pad  ;
	input s_pad ;
	input \t0_pad  ;
	input t_pad ;
	input \u0_pad  ;
	input u_pad ;
	input \v0_pad  ;
	input v_pad ;
	input w_pad ;
	input x_pad ;
	input y_pad ;
	input z_pad ;
	output \a1_pad  ;
	output \a2_pad  ;
	output \b1_pad  ;
	output \b2_pad  ;
	output \c1_pad  ;
	output \c2_pad  ;
	output \d1_pad  ;
	output \d2_pad  ;
	output \e1_pad  ;
	output \e2_pad  ;
	output \f1_pad  ;
	output \f2_pad  ;
	output \g1_pad  ;
	output \h1_pad  ;
	output \i1_pad  ;
	output \j1_pad  ;
	output \k1_pad  ;
	output \l1_pad  ;
	output \m1_pad  ;
	output \n1_pad  ;
	output \o1_pad  ;
	output \p1_pad  ;
	output \q1_pad  ;
	output \r1_pad  ;
	output \s1_pad  ;
	output \t1_pad  ;
	output \u1_pad  ;
	output \v1_pad  ;
	output \w0_pad  ;
	output \w1_pad  ;
	output \x0_pad  ;
	output \x1_pad  ;
	output \y0_pad  ;
	output \y1_pad  ;
	output \z0_pad  ;
	output \z1_pad  ;
	wire _w195_ ;
	wire _w194_ ;
	wire _w193_ ;
	wire _w192_ ;
	wire _w191_ ;
	wire _w190_ ;
	wire _w189_ ;
	wire _w188_ ;
	wire _w187_ ;
	wire _w186_ ;
	wire _w185_ ;
	wire _w184_ ;
	wire _w183_ ;
	wire _w182_ ;
	wire _w181_ ;
	wire _w180_ ;
	wire _w179_ ;
	wire _w178_ ;
	wire _w177_ ;
	wire _w176_ ;
	wire _w175_ ;
	wire _w106_ ;
	wire _w105_ ;
	wire _w104_ ;
	wire _w103_ ;
	wire _w102_ ;
	wire _w101_ ;
	wire _w100_ ;
	wire _w99_ ;
	wire _w98_ ;
	wire _w97_ ;
	wire _w96_ ;
	wire _w95_ ;
	wire _w94_ ;
	wire _w93_ ;
	wire _w92_ ;
	wire _w91_ ;
	wire _w90_ ;
	wire _w89_ ;
	wire _w88_ ;
	wire _w87_ ;
	wire _w86_ ;
	wire _w85_ ;
	wire _w84_ ;
	wire _w83_ ;
	wire _w82_ ;
	wire _w81_ ;
	wire _w80_ ;
	wire _w79_ ;
	wire _w78_ ;
	wire _w77_ ;
	wire _w60_ ;
	wire _w59_ ;
	wire _w58_ ;
	wire _w57_ ;
	wire _w56_ ;
	wire _w55_ ;
	wire _w54_ ;
	wire _w53_ ;
	wire _w52_ ;
	wire _w51_ ;
	wire _w50_ ;
	wire _w49_ ;
	wire _w48_ ;
	wire _w61_ ;
	wire _w62_ ;
	wire _w63_ ;
	wire _w64_ ;
	wire _w65_ ;
	wire _w66_ ;
	wire _w67_ ;
	wire _w68_ ;
	wire _w69_ ;
	wire _w70_ ;
	wire _w71_ ;
	wire _w72_ ;
	wire _w73_ ;
	wire _w74_ ;
	wire _w75_ ;
	wire _w76_ ;
	wire _w107_ ;
	wire _w108_ ;
	wire _w109_ ;
	wire _w110_ ;
	wire _w111_ ;
	wire _w112_ ;
	wire _w113_ ;
	wire _w114_ ;
	wire _w115_ ;
	wire _w116_ ;
	wire _w117_ ;
	wire _w118_ ;
	wire _w119_ ;
	wire _w120_ ;
	wire _w121_ ;
	wire _w122_ ;
	wire _w123_ ;
	wire _w124_ ;
	wire _w125_ ;
	wire _w126_ ;
	wire _w127_ ;
	wire _w128_ ;
	wire _w129_ ;
	wire _w130_ ;
	wire _w131_ ;
	wire _w132_ ;
	wire _w133_ ;
	wire _w134_ ;
	wire _w135_ ;
	wire _w136_ ;
	wire _w137_ ;
	wire _w138_ ;
	wire _w139_ ;
	wire _w140_ ;
	wire _w141_ ;
	wire _w142_ ;
	wire _w143_ ;
	wire _w144_ ;
	wire _w145_ ;
	wire _w146_ ;
	wire _w147_ ;
	wire _w148_ ;
	wire _w149_ ;
	wire _w150_ ;
	wire _w151_ ;
	wire _w152_ ;
	wire _w153_ ;
	wire _w154_ ;
	wire _w155_ ;
	wire _w156_ ;
	wire _w157_ ;
	wire _w158_ ;
	wire _w159_ ;
	wire _w160_ ;
	wire _w161_ ;
	wire _w162_ ;
	wire _w163_ ;
	wire _w164_ ;
	wire _w165_ ;
	wire _w166_ ;
	wire _w167_ ;
	wire _w168_ ;
	wire _w169_ ;
	wire _w170_ ;
	wire _w171_ ;
	wire _w172_ ;
	wire _w173_ ;
	wire _w174_ ;
	LUT2 #(
		.INIT('h1)
	) name0 (
		i_pad,
		q_pad,
		_w48_
	);
	LUT2 #(
		.INIT('h4)
	) name1 (
		d_pad,
		i_pad,
		_w49_
	);
	LUT2 #(
		.INIT('h1)
	) name2 (
		l_pad,
		_w48_,
		_w50_
	);
	LUT2 #(
		.INIT('h4)
	) name3 (
		_w49_,
		_w50_,
		_w51_
	);
	LUT2 #(
		.INIT('h2)
	) name4 (
		k_pad,
		p_pad,
		_w52_
	);
	LUT2 #(
		.INIT('h1)
	) name5 (
		\q0_pad ,
		_w52_,
		_w53_
	);
	LUT2 #(
		.INIT('h4)
	) name6 (
		\r0_pad ,
		_w52_,
		_w54_
	);
	LUT2 #(
		.INIT('h1)
	) name7 (
		l_pad,
		_w53_,
		_w55_
	);
	LUT2 #(
		.INIT('h4)
	) name8 (
		_w54_,
		_w55_,
		_w56_
	);
	LUT2 #(
		.INIT('h1)
	) name9 (
		i_pad,
		r_pad,
		_w57_
	);
	LUT2 #(
		.INIT('h4)
	) name10 (
		e_pad,
		i_pad,
		_w58_
	);
	LUT2 #(
		.INIT('h1)
	) name11 (
		l_pad,
		_w57_,
		_w59_
	);
	LUT2 #(
		.INIT('h4)
	) name12 (
		_w58_,
		_w59_,
		_w60_
	);
	LUT2 #(
		.INIT('h1)
	) name13 (
		\r0_pad ,
		_w52_,
		_w61_
	);
	LUT2 #(
		.INIT('h4)
	) name14 (
		\s0_pad ,
		_w52_,
		_w62_
	);
	LUT2 #(
		.INIT('h1)
	) name15 (
		l_pad,
		_w61_,
		_w63_
	);
	LUT2 #(
		.INIT('h4)
	) name16 (
		_w62_,
		_w63_,
		_w64_
	);
	LUT2 #(
		.INIT('h1)
	) name17 (
		j_pad,
		s_pad,
		_w65_
	);
	LUT2 #(
		.INIT('h2)
	) name18 (
		j_pad,
		t_pad,
		_w66_
	);
	LUT2 #(
		.INIT('h1)
	) name19 (
		l_pad,
		_w65_,
		_w67_
	);
	LUT2 #(
		.INIT('h4)
	) name20 (
		_w66_,
		_w67_,
		_w68_
	);
	LUT2 #(
		.INIT('h1)
	) name21 (
		\s0_pad ,
		_w52_,
		_w69_
	);
	LUT2 #(
		.INIT('h4)
	) name22 (
		\t0_pad ,
		_w52_,
		_w70_
	);
	LUT2 #(
		.INIT('h1)
	) name23 (
		l_pad,
		_w69_,
		_w71_
	);
	LUT2 #(
		.INIT('h4)
	) name24 (
		_w70_,
		_w71_,
		_w72_
	);
	LUT2 #(
		.INIT('h1)
	) name25 (
		j_pad,
		t_pad,
		_w73_
	);
	LUT2 #(
		.INIT('h2)
	) name26 (
		j_pad,
		u_pad,
		_w74_
	);
	LUT2 #(
		.INIT('h1)
	) name27 (
		l_pad,
		_w73_,
		_w75_
	);
	LUT2 #(
		.INIT('h4)
	) name28 (
		_w74_,
		_w75_,
		_w76_
	);
	LUT2 #(
		.INIT('h1)
	) name29 (
		\t0_pad ,
		_w52_,
		_w77_
	);
	LUT2 #(
		.INIT('h4)
	) name30 (
		\u0_pad ,
		_w52_,
		_w78_
	);
	LUT2 #(
		.INIT('h1)
	) name31 (
		l_pad,
		_w77_,
		_w79_
	);
	LUT2 #(
		.INIT('h4)
	) name32 (
		_w78_,
		_w79_,
		_w80_
	);
	LUT2 #(
		.INIT('h1)
	) name33 (
		j_pad,
		u_pad,
		_w81_
	);
	LUT2 #(
		.INIT('h2)
	) name34 (
		j_pad,
		v_pad,
		_w82_
	);
	LUT2 #(
		.INIT('h1)
	) name35 (
		l_pad,
		_w81_,
		_w83_
	);
	LUT2 #(
		.INIT('h4)
	) name36 (
		_w82_,
		_w83_,
		_w84_
	);
	LUT2 #(
		.INIT('h1)
	) name37 (
		\u0_pad ,
		_w52_,
		_w85_
	);
	LUT2 #(
		.INIT('h4)
	) name38 (
		\v0_pad ,
		_w52_,
		_w86_
	);
	LUT2 #(
		.INIT('h1)
	) name39 (
		l_pad,
		_w85_,
		_w87_
	);
	LUT2 #(
		.INIT('h4)
	) name40 (
		_w86_,
		_w87_,
		_w88_
	);
	LUT2 #(
		.INIT('h1)
	) name41 (
		j_pad,
		v_pad,
		_w89_
	);
	LUT2 #(
		.INIT('h2)
	) name42 (
		j_pad,
		w_pad,
		_w90_
	);
	LUT2 #(
		.INIT('h1)
	) name43 (
		l_pad,
		_w89_,
		_w91_
	);
	LUT2 #(
		.INIT('h4)
	) name44 (
		_w90_,
		_w91_,
		_w92_
	);
	LUT2 #(
		.INIT('h1)
	) name45 (
		\v0_pad ,
		_w52_,
		_w93_
	);
	LUT2 #(
		.INIT('h4)
	) name46 (
		a_pad,
		_w52_,
		_w94_
	);
	LUT2 #(
		.INIT('h1)
	) name47 (
		l_pad,
		_w93_,
		_w95_
	);
	LUT2 #(
		.INIT('h4)
	) name48 (
		_w94_,
		_w95_,
		_w96_
	);
	LUT2 #(
		.INIT('h1)
	) name49 (
		j_pad,
		w_pad,
		_w97_
	);
	LUT2 #(
		.INIT('h2)
	) name50 (
		j_pad,
		x_pad,
		_w98_
	);
	LUT2 #(
		.INIT('h1)
	) name51 (
		l_pad,
		_w97_,
		_w99_
	);
	LUT2 #(
		.INIT('h4)
	) name52 (
		_w98_,
		_w99_,
		_w100_
	);
	LUT2 #(
		.INIT('h1)
	) name53 (
		j_pad,
		x_pad,
		_w101_
	);
	LUT2 #(
		.INIT('h2)
	) name54 (
		j_pad,
		y_pad,
		_w102_
	);
	LUT2 #(
		.INIT('h1)
	) name55 (
		l_pad,
		_w101_,
		_w103_
	);
	LUT2 #(
		.INIT('h4)
	) name56 (
		_w102_,
		_w103_,
		_w104_
	);
	LUT2 #(
		.INIT('h1)
	) name57 (
		j_pad,
		y_pad,
		_w105_
	);
	LUT2 #(
		.INIT('h2)
	) name58 (
		j_pad,
		z_pad,
		_w106_
	);
	LUT2 #(
		.INIT('h1)
	) name59 (
		l_pad,
		_w105_,
		_w107_
	);
	LUT2 #(
		.INIT('h4)
	) name60 (
		_w106_,
		_w107_,
		_w108_
	);
	LUT2 #(
		.INIT('h1)
	) name61 (
		j_pad,
		z_pad,
		_w109_
	);
	LUT2 #(
		.INIT('h4)
	) name62 (
		\a0_pad ,
		j_pad,
		_w110_
	);
	LUT2 #(
		.INIT('h1)
	) name63 (
		l_pad,
		_w109_,
		_w111_
	);
	LUT2 #(
		.INIT('h4)
	) name64 (
		_w110_,
		_w111_,
		_w112_
	);
	LUT2 #(
		.INIT('h1)
	) name65 (
		\a0_pad ,
		j_pad,
		_w113_
	);
	LUT2 #(
		.INIT('h4)
	) name66 (
		\b0_pad ,
		j_pad,
		_w114_
	);
	LUT2 #(
		.INIT('h1)
	) name67 (
		l_pad,
		_w113_,
		_w115_
	);
	LUT2 #(
		.INIT('h4)
	) name68 (
		_w114_,
		_w115_,
		_w116_
	);
	LUT2 #(
		.INIT('h1)
	) name69 (
		\b0_pad ,
		j_pad,
		_w117_
	);
	LUT2 #(
		.INIT('h4)
	) name70 (
		\c0_pad ,
		j_pad,
		_w118_
	);
	LUT2 #(
		.INIT('h1)
	) name71 (
		l_pad,
		_w117_,
		_w119_
	);
	LUT2 #(
		.INIT('h4)
	) name72 (
		_w118_,
		_w119_,
		_w120_
	);
	LUT2 #(
		.INIT('h1)
	) name73 (
		\c0_pad ,
		j_pad,
		_w121_
	);
	LUT2 #(
		.INIT('h4)
	) name74 (
		\d0_pad ,
		j_pad,
		_w122_
	);
	LUT2 #(
		.INIT('h1)
	) name75 (
		l_pad,
		_w121_,
		_w123_
	);
	LUT2 #(
		.INIT('h4)
	) name76 (
		_w122_,
		_w123_,
		_w124_
	);
	LUT2 #(
		.INIT('h1)
	) name77 (
		\d0_pad ,
		j_pad,
		_w125_
	);
	LUT2 #(
		.INIT('h4)
	) name78 (
		\e0_pad ,
		j_pad,
		_w126_
	);
	LUT2 #(
		.INIT('h1)
	) name79 (
		l_pad,
		_w125_,
		_w127_
	);
	LUT2 #(
		.INIT('h4)
	) name80 (
		_w126_,
		_w127_,
		_w128_
	);
	LUT2 #(
		.INIT('h1)
	) name81 (
		\e0_pad ,
		j_pad,
		_w129_
	);
	LUT2 #(
		.INIT('h4)
	) name82 (
		\f0_pad ,
		j_pad,
		_w130_
	);
	LUT2 #(
		.INIT('h1)
	) name83 (
		l_pad,
		_w129_,
		_w131_
	);
	LUT2 #(
		.INIT('h4)
	) name84 (
		_w130_,
		_w131_,
		_w132_
	);
	LUT2 #(
		.INIT('h1)
	) name85 (
		\f0_pad ,
		j_pad,
		_w133_
	);
	LUT2 #(
		.INIT('h4)
	) name86 (
		a_pad,
		j_pad,
		_w134_
	);
	LUT2 #(
		.INIT('h1)
	) name87 (
		l_pad,
		_w133_,
		_w135_
	);
	LUT2 #(
		.INIT('h4)
	) name88 (
		_w134_,
		_w135_,
		_w136_
	);
	LUT2 #(
		.INIT('h1)
	) name89 (
		\g0_pad ,
		k_pad,
		_w137_
	);
	LUT2 #(
		.INIT('h4)
	) name90 (
		\h0_pad ,
		k_pad,
		_w138_
	);
	LUT2 #(
		.INIT('h1)
	) name91 (
		l_pad,
		_w137_,
		_w139_
	);
	LUT2 #(
		.INIT('h4)
	) name92 (
		_w138_,
		_w139_,
		_w140_
	);
	LUT2 #(
		.INIT('h1)
	) name93 (
		\h0_pad ,
		k_pad,
		_w141_
	);
	LUT2 #(
		.INIT('h4)
	) name94 (
		\i0_pad ,
		k_pad,
		_w142_
	);
	LUT2 #(
		.INIT('h1)
	) name95 (
		l_pad,
		_w141_,
		_w143_
	);
	LUT2 #(
		.INIT('h4)
	) name96 (
		_w142_,
		_w143_,
		_w144_
	);
	LUT2 #(
		.INIT('h1)
	) name97 (
		\i0_pad ,
		k_pad,
		_w145_
	);
	LUT2 #(
		.INIT('h4)
	) name98 (
		\j0_pad ,
		k_pad,
		_w146_
	);
	LUT2 #(
		.INIT('h1)
	) name99 (
		l_pad,
		_w145_,
		_w147_
	);
	LUT2 #(
		.INIT('h4)
	) name100 (
		_w146_,
		_w147_,
		_w148_
	);
	LUT2 #(
		.INIT('h1)
	) name101 (
		\j0_pad ,
		k_pad,
		_w149_
	);
	LUT2 #(
		.INIT('h4)
	) name102 (
		\k0_pad ,
		k_pad,
		_w150_
	);
	LUT2 #(
		.INIT('h1)
	) name103 (
		l_pad,
		_w149_,
		_w151_
	);
	LUT2 #(
		.INIT('h4)
	) name104 (
		_w150_,
		_w151_,
		_w152_
	);
	LUT2 #(
		.INIT('h1)
	) name105 (
		\k0_pad ,
		k_pad,
		_w153_
	);
	LUT2 #(
		.INIT('h2)
	) name106 (
		k_pad,
		\l0_pad ,
		_w154_
	);
	LUT2 #(
		.INIT('h1)
	) name107 (
		l_pad,
		_w153_,
		_w155_
	);
	LUT2 #(
		.INIT('h4)
	) name108 (
		_w154_,
		_w155_,
		_w156_
	);
	LUT2 #(
		.INIT('h1)
	) name109 (
		k_pad,
		\l0_pad ,
		_w157_
	);
	LUT2 #(
		.INIT('h2)
	) name110 (
		k_pad,
		\m0_pad ,
		_w158_
	);
	LUT2 #(
		.INIT('h1)
	) name111 (
		l_pad,
		_w157_,
		_w159_
	);
	LUT2 #(
		.INIT('h4)
	) name112 (
		_w158_,
		_w159_,
		_w160_
	);
	LUT2 #(
		.INIT('h1)
	) name113 (
		i_pad,
		m_pad,
		_w161_
	);
	LUT2 #(
		.INIT('h4)
	) name114 (
		f_pad,
		i_pad,
		_w162_
	);
	LUT2 #(
		.INIT('h1)
	) name115 (
		l_pad,
		_w161_,
		_w163_
	);
	LUT2 #(
		.INIT('h4)
	) name116 (
		_w162_,
		_w163_,
		_w164_
	);
	LUT2 #(
		.INIT('h1)
	) name117 (
		k_pad,
		\m0_pad ,
		_w165_
	);
	LUT2 #(
		.INIT('h2)
	) name118 (
		k_pad,
		\n0_pad ,
		_w166_
	);
	LUT2 #(
		.INIT('h1)
	) name119 (
		l_pad,
		_w165_,
		_w167_
	);
	LUT2 #(
		.INIT('h4)
	) name120 (
		_w166_,
		_w167_,
		_w168_
	);
	LUT2 #(
		.INIT('h1)
	) name121 (
		i_pad,
		n_pad,
		_w169_
	);
	LUT2 #(
		.INIT('h4)
	) name122 (
		g_pad,
		i_pad,
		_w170_
	);
	LUT2 #(
		.INIT('h1)
	) name123 (
		l_pad,
		_w169_,
		_w171_
	);
	LUT2 #(
		.INIT('h4)
	) name124 (
		_w170_,
		_w171_,
		_w172_
	);
	LUT2 #(
		.INIT('h1)
	) name125 (
		k_pad,
		\n0_pad ,
		_w173_
	);
	LUT2 #(
		.INIT('h2)
	) name126 (
		\o0_pad ,
		p_pad,
		_w174_
	);
	LUT2 #(
		.INIT('h8)
	) name127 (
		a_pad,
		p_pad,
		_w175_
	);
	LUT2 #(
		.INIT('h2)
	) name128 (
		k_pad,
		_w174_,
		_w176_
	);
	LUT2 #(
		.INIT('h4)
	) name129 (
		_w175_,
		_w176_,
		_w177_
	);
	LUT2 #(
		.INIT('h1)
	) name130 (
		l_pad,
		_w173_,
		_w178_
	);
	LUT2 #(
		.INIT('h4)
	) name131 (
		_w177_,
		_w178_,
		_w179_
	);
	LUT2 #(
		.INIT('h1)
	) name132 (
		i_pad,
		o_pad,
		_w180_
	);
	LUT2 #(
		.INIT('h4)
	) name133 (
		h_pad,
		i_pad,
		_w181_
	);
	LUT2 #(
		.INIT('h1)
	) name134 (
		l_pad,
		_w180_,
		_w182_
	);
	LUT2 #(
		.INIT('h4)
	) name135 (
		_w181_,
		_w182_,
		_w183_
	);
	LUT2 #(
		.INIT('h1)
	) name136 (
		\o0_pad ,
		_w52_,
		_w184_
	);
	LUT2 #(
		.INIT('h4)
	) name137 (
		\p0_pad ,
		_w52_,
		_w185_
	);
	LUT2 #(
		.INIT('h1)
	) name138 (
		l_pad,
		_w184_,
		_w186_
	);
	LUT2 #(
		.INIT('h4)
	) name139 (
		_w185_,
		_w186_,
		_w187_
	);
	LUT2 #(
		.INIT('h1)
	) name140 (
		i_pad,
		p_pad,
		_w188_
	);
	LUT2 #(
		.INIT('h4)
	) name141 (
		c_pad,
		i_pad,
		_w189_
	);
	LUT2 #(
		.INIT('h1)
	) name142 (
		l_pad,
		_w188_,
		_w190_
	);
	LUT2 #(
		.INIT('h4)
	) name143 (
		_w189_,
		_w190_,
		_w191_
	);
	LUT2 #(
		.INIT('h1)
	) name144 (
		\p0_pad ,
		_w52_,
		_w192_
	);
	LUT2 #(
		.INIT('h4)
	) name145 (
		\q0_pad ,
		_w52_,
		_w193_
	);
	LUT2 #(
		.INIT('h1)
	) name146 (
		l_pad,
		_w192_,
		_w194_
	);
	LUT2 #(
		.INIT('h4)
	) name147 (
		_w193_,
		_w194_,
		_w195_
	);
	assign \a1_pad  = _w51_ ;
	assign \a2_pad  = _w56_ ;
	assign \b1_pad  = _w60_ ;
	assign \b2_pad  = _w64_ ;
	assign \c1_pad  = _w68_ ;
	assign \c2_pad  = _w72_ ;
	assign \d1_pad  = _w76_ ;
	assign \d2_pad  = _w80_ ;
	assign \e1_pad  = _w84_ ;
	assign \e2_pad  = _w88_ ;
	assign \f1_pad  = _w92_ ;
	assign \f2_pad  = _w96_ ;
	assign \g1_pad  = _w100_ ;
	assign \h1_pad  = _w104_ ;
	assign \i1_pad  = _w108_ ;
	assign \j1_pad  = _w112_ ;
	assign \k1_pad  = _w116_ ;
	assign \l1_pad  = _w120_ ;
	assign \m1_pad  = _w124_ ;
	assign \n1_pad  = _w128_ ;
	assign \o1_pad  = _w132_ ;
	assign \p1_pad  = _w136_ ;
	assign \q1_pad  = _w140_ ;
	assign \r1_pad  = _w144_ ;
	assign \s1_pad  = _w148_ ;
	assign \t1_pad  = _w152_ ;
	assign \u1_pad  = _w156_ ;
	assign \v1_pad  = _w160_ ;
	assign \w0_pad  = _w164_ ;
	assign \w1_pad  = _w168_ ;
	assign \x0_pad  = _w172_ ;
	assign \x1_pad  = _w179_ ;
	assign \y0_pad  = _w183_ ;
	assign \y1_pad  = _w187_ ;
	assign \z0_pad  = _w191_ ;
	assign \z1_pad  = _w195_ ;
endmodule;