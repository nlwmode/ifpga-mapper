module top (\100(51)_pad , \103(52)_pad , \109(54)_pad , \110(55)_pad , \111(56)_pad , \112(57)_pad , \113(58)_pad , \114(59)_pad , \115(60)_pad , \118(61)_pad , \1197(165)_pad , \12(3)_pad , \121(62)_pad , \124(63)_pad , \127(64)_pad , \130(65)_pad , \133(66)_pad , \134(67)_pad , \135(68)_pad , \138(69)_pad , \141(70)_pad , \144(71)_pad , \1455(166)_pad , \147(72)_pad , \15(4)_pad , \150(73)_pad , \151(74)_pad , \152(75)_pad , \153(76)_pad , \154(77)_pad , \155(78)_pad , \156(79)_pad , \157(80)_pad , \158(81)_pad , \159(82)_pad , \160(83)_pad , \161(84)_pad , \162(85)_pad , \163(86)_pad , \164(87)_pad , \165(88)_pad , \166(89)_pad , \167(90)_pad , \168(91)_pad , \169(92)_pad , \170(93)_pad , \171(94)_pad , \172(95)_pad , \173(96)_pad , \174(97)_pad , \175(98)_pad , \176(99)_pad , \177(100)_pad , \178(101)_pad , \179(102)_pad , \18(5)_pad , \180(103)_pad , \181(104)_pad , \182(105)_pad , \183(106)_pad , \184(107)_pad , \185(108)_pad , \186(109)_pad , \187(110)_pad , \188(111)_pad , \189(112)_pad , \190(113)_pad , \191(114)_pad , \192(115)_pad , \193(116)_pad , \194(117)_pad , \195(118)_pad , \196(119)_pad , \197(120)_pad , \198(121)_pad , \199(122)_pad , \200(123)_pad , \201(124)_pad , \202(125)_pad , \203(126)_pad , \204(127)_pad , \205(128)_pad , \206(129)_pad , \207(130)_pad , \208(131)_pad , \209(132)_pad , \210(133)_pad , \211(134)_pad , \212(135)_pad , \213(136)_pad , \214(137)_pad , \215(138)_pad , \216(139)_pad , \217(140)_pad , \218(141)_pad , \219(142)_pad , \220(143)_pad , \2204(174)_pad , \221(144)_pad , \222(145)_pad , \223(146)_pad , \224(147)_pad , \225(148)_pad , \226(149)_pad , \227(150)_pad , \228(151)_pad , \229(152)_pad , \23(6)_pad , \230(153)_pad , \231(154)_pad , \232(155)_pad , \233(156)_pad , \234(157)_pad , \235(158)_pad , \236(159)_pad , \237(160)_pad , \238(161)_pad , \239(162)_pad , \240(163)_pad , \26(7)_pad , \29(8)_pad , \32(9)_pad , \35(10)_pad , \38(11)_pad , \41(12)_pad , \436(286)_pad , \438(274)_pad , \44(13)_pad , \440(277)_pad , \442(280)_pad , \444(282)_pad , \446(393)_pad , \448(284)_pad , \450(288)_pad , \4526(205)_pad , \4528(206)_pad , \453(596)_pad , \47(14)_pad , \478(269)_pad , \480(250)_pad , \482(253)_pad , \484(256)_pad , \486(258)_pad , \488(260)_pad , \490(263)_pad , \492(265)_pad , \494(267)_pad , \496(271)_pad , \5(1)_pad , \50(15)_pad , \522(226)_pad , \524(210)_pad , \526(212)_pad , \528(214)_pad , \53(16)_pad , \530(216)_pad , \532(218)_pad , \534(220)_pad , \536(222)_pad , \538(224)_pad , \54(17)_pad , \540(227)_pad , \542(246)_pad , \544(230)_pad , \546(232)_pad , \548(234)_pad , \55(18)_pad , \550(236)_pad , \552(238)_pad , \554(240)_pad , \556(242)_pad , \558(244)_pad , \56(19)_pad , \560(248)_pad , \57(20)_pad , \58(21)_pad , \59(22)_pad , \60(23)_pad , \61(24)_pad , \62(25)_pad , \63(26)_pad , \64(27)_pad , \65(28)_pad , \66(29)_pad , \69(30)_pad , \70(31)_pad , \73(32)_pad , \74(33)_pad , \75(34)_pad , \76(35)_pad , \77(36)_pad , \78(37)_pad , \79(38)_pad , \80(39)_pad , \81(40)_pad , \82(41)_pad , \83(42)_pad , \84(43)_pad , \85(44)_pad , \86(45)_pad , \87(46)_pad , \88(47)_pad , \89(48)_pad , \9(2)_pad , \94(49)_pad , \97(50)_pad , \252(3450)_pad , \258(3122)_pad , \270(3109)_pad , \278(536)_pad , \281(547)_pad , \284(384)_pad , \286(419)_pad , \292(392)_pad , \295(3352)_pad , \298(3387)_pad , \301(3388)_pad , \304(3390)_pad , \307(3389)_pad , \310(3393)_pad , \313(3396)_pad , \316(3397)_pad , \319(3398)_pad , \321(3715)_pad , \324(3363)_pad , \327(3408)_pad , \330(3411)_pad , \333(3416)_pad , \336(3412)_pad , \338(3716)_pad , \344(3382)_pad , \347(3420)_pad , \350(3421)_pad , \353(3425)_pad , \356(3424)_pad , \359(3426)_pad , \362(3429)_pad , \365(3430)_pad , \368(3431)_pad , \370(3718)_pad , \373(2994)_pad , \376(3206)_pad , \379(3207)_pad , \382(3148)_pad , \385(3151)_pad , \388(3093)_pad , \391(3094)_pad , \394(3095)_pad , \397(3097)_pad , \399(3717)_pad , \402(395)_pad , \404(390)_pad , \406(388)_pad , \408(385)_pad , \410(387)_pad , \412(3369)_pad , \414(3338)_pad , \416(3368)_pad , \418(3449)_pad , \419(3444)_pad , \422(3451)_pad );
	input \100(51)_pad  ;
	input \103(52)_pad  ;
	input \109(54)_pad  ;
	input \110(55)_pad  ;
	input \111(56)_pad  ;
	input \112(57)_pad  ;
	input \113(58)_pad  ;
	input \114(59)_pad  ;
	input \115(60)_pad  ;
	input \118(61)_pad  ;
	input \1197(165)_pad  ;
	input \12(3)_pad  ;
	input \121(62)_pad  ;
	input \124(63)_pad  ;
	input \127(64)_pad  ;
	input \130(65)_pad  ;
	input \133(66)_pad  ;
	input \134(67)_pad  ;
	input \135(68)_pad  ;
	input \138(69)_pad  ;
	input \141(70)_pad  ;
	input \144(71)_pad  ;
	input \1455(166)_pad  ;
	input \147(72)_pad  ;
	input \15(4)_pad  ;
	input \150(73)_pad  ;
	input \151(74)_pad  ;
	input \152(75)_pad  ;
	input \153(76)_pad  ;
	input \154(77)_pad  ;
	input \155(78)_pad  ;
	input \156(79)_pad  ;
	input \157(80)_pad  ;
	input \158(81)_pad  ;
	input \159(82)_pad  ;
	input \160(83)_pad  ;
	input \161(84)_pad  ;
	input \162(85)_pad  ;
	input \163(86)_pad  ;
	input \164(87)_pad  ;
	input \165(88)_pad  ;
	input \166(89)_pad  ;
	input \167(90)_pad  ;
	input \168(91)_pad  ;
	input \169(92)_pad  ;
	input \170(93)_pad  ;
	input \171(94)_pad  ;
	input \172(95)_pad  ;
	input \173(96)_pad  ;
	input \174(97)_pad  ;
	input \175(98)_pad  ;
	input \176(99)_pad  ;
	input \177(100)_pad  ;
	input \178(101)_pad  ;
	input \179(102)_pad  ;
	input \18(5)_pad  ;
	input \180(103)_pad  ;
	input \181(104)_pad  ;
	input \182(105)_pad  ;
	input \183(106)_pad  ;
	input \184(107)_pad  ;
	input \185(108)_pad  ;
	input \186(109)_pad  ;
	input \187(110)_pad  ;
	input \188(111)_pad  ;
	input \189(112)_pad  ;
	input \190(113)_pad  ;
	input \191(114)_pad  ;
	input \192(115)_pad  ;
	input \193(116)_pad  ;
	input \194(117)_pad  ;
	input \195(118)_pad  ;
	input \196(119)_pad  ;
	input \197(120)_pad  ;
	input \198(121)_pad  ;
	input \199(122)_pad  ;
	input \200(123)_pad  ;
	input \201(124)_pad  ;
	input \202(125)_pad  ;
	input \203(126)_pad  ;
	input \204(127)_pad  ;
	input \205(128)_pad  ;
	input \206(129)_pad  ;
	input \207(130)_pad  ;
	input \208(131)_pad  ;
	input \209(132)_pad  ;
	input \210(133)_pad  ;
	input \211(134)_pad  ;
	input \212(135)_pad  ;
	input \213(136)_pad  ;
	input \214(137)_pad  ;
	input \215(138)_pad  ;
	input \216(139)_pad  ;
	input \217(140)_pad  ;
	input \218(141)_pad  ;
	input \219(142)_pad  ;
	input \220(143)_pad  ;
	input \2204(174)_pad  ;
	input \221(144)_pad  ;
	input \222(145)_pad  ;
	input \223(146)_pad  ;
	input \224(147)_pad  ;
	input \225(148)_pad  ;
	input \226(149)_pad  ;
	input \227(150)_pad  ;
	input \228(151)_pad  ;
	input \229(152)_pad  ;
	input \23(6)_pad  ;
	input \230(153)_pad  ;
	input \231(154)_pad  ;
	input \232(155)_pad  ;
	input \233(156)_pad  ;
	input \234(157)_pad  ;
	input \235(158)_pad  ;
	input \236(159)_pad  ;
	input \237(160)_pad  ;
	input \238(161)_pad  ;
	input \239(162)_pad  ;
	input \240(163)_pad  ;
	input \26(7)_pad  ;
	input \29(8)_pad  ;
	input \32(9)_pad  ;
	input \35(10)_pad  ;
	input \38(11)_pad  ;
	input \41(12)_pad  ;
	input \436(286)_pad  ;
	input \438(274)_pad  ;
	input \44(13)_pad  ;
	input \440(277)_pad  ;
	input \442(280)_pad  ;
	input \444(282)_pad  ;
	input \446(393)_pad  ;
	input \448(284)_pad  ;
	input \450(288)_pad  ;
	input \4526(205)_pad  ;
	input \4528(206)_pad  ;
	input \453(596)_pad  ;
	input \47(14)_pad  ;
	input \478(269)_pad  ;
	input \480(250)_pad  ;
	input \482(253)_pad  ;
	input \484(256)_pad  ;
	input \486(258)_pad  ;
	input \488(260)_pad  ;
	input \490(263)_pad  ;
	input \492(265)_pad  ;
	input \494(267)_pad  ;
	input \496(271)_pad  ;
	input \5(1)_pad  ;
	input \50(15)_pad  ;
	input \522(226)_pad  ;
	input \524(210)_pad  ;
	input \526(212)_pad  ;
	input \528(214)_pad  ;
	input \53(16)_pad  ;
	input \530(216)_pad  ;
	input \532(218)_pad  ;
	input \534(220)_pad  ;
	input \536(222)_pad  ;
	input \538(224)_pad  ;
	input \54(17)_pad  ;
	input \540(227)_pad  ;
	input \542(246)_pad  ;
	input \544(230)_pad  ;
	input \546(232)_pad  ;
	input \548(234)_pad  ;
	input \55(18)_pad  ;
	input \550(236)_pad  ;
	input \552(238)_pad  ;
	input \554(240)_pad  ;
	input \556(242)_pad  ;
	input \558(244)_pad  ;
	input \56(19)_pad  ;
	input \560(248)_pad  ;
	input \57(20)_pad  ;
	input \58(21)_pad  ;
	input \59(22)_pad  ;
	input \60(23)_pad  ;
	input \61(24)_pad  ;
	input \62(25)_pad  ;
	input \63(26)_pad  ;
	input \64(27)_pad  ;
	input \65(28)_pad  ;
	input \66(29)_pad  ;
	input \69(30)_pad  ;
	input \70(31)_pad  ;
	input \73(32)_pad  ;
	input \74(33)_pad  ;
	input \75(34)_pad  ;
	input \76(35)_pad  ;
	input \77(36)_pad  ;
	input \78(37)_pad  ;
	input \79(38)_pad  ;
	input \80(39)_pad  ;
	input \81(40)_pad  ;
	input \82(41)_pad  ;
	input \83(42)_pad  ;
	input \84(43)_pad  ;
	input \85(44)_pad  ;
	input \86(45)_pad  ;
	input \87(46)_pad  ;
	input \88(47)_pad  ;
	input \89(48)_pad  ;
	input \9(2)_pad  ;
	input \94(49)_pad  ;
	input \97(50)_pad  ;
	output \252(3450)_pad  ;
	output \258(3122)_pad  ;
	output \270(3109)_pad  ;
	output \278(536)_pad  ;
	output \281(547)_pad  ;
	output \284(384)_pad  ;
	output \286(419)_pad  ;
	output \292(392)_pad  ;
	output \295(3352)_pad  ;
	output \298(3387)_pad  ;
	output \301(3388)_pad  ;
	output \304(3390)_pad  ;
	output \307(3389)_pad  ;
	output \310(3393)_pad  ;
	output \313(3396)_pad  ;
	output \316(3397)_pad  ;
	output \319(3398)_pad  ;
	output \321(3715)_pad  ;
	output \324(3363)_pad  ;
	output \327(3408)_pad  ;
	output \330(3411)_pad  ;
	output \333(3416)_pad  ;
	output \336(3412)_pad  ;
	output \338(3716)_pad  ;
	output \344(3382)_pad  ;
	output \347(3420)_pad  ;
	output \350(3421)_pad  ;
	output \353(3425)_pad  ;
	output \356(3424)_pad  ;
	output \359(3426)_pad  ;
	output \362(3429)_pad  ;
	output \365(3430)_pad  ;
	output \368(3431)_pad  ;
	output \370(3718)_pad  ;
	output \373(2994)_pad  ;
	output \376(3206)_pad  ;
	output \379(3207)_pad  ;
	output \382(3148)_pad  ;
	output \385(3151)_pad  ;
	output \388(3093)_pad  ;
	output \391(3094)_pad  ;
	output \394(3095)_pad  ;
	output \397(3097)_pad  ;
	output \399(3717)_pad  ;
	output \402(395)_pad  ;
	output \404(390)_pad  ;
	output \406(388)_pad  ;
	output \408(385)_pad  ;
	output \410(387)_pad  ;
	output \412(3369)_pad  ;
	output \414(3338)_pad  ;
	output \416(3368)_pad  ;
	output \418(3449)_pad  ;
	output \419(3444)_pad  ;
	output \422(3451)_pad  ;
	wire _w932_ ;
	wire _w931_ ;
	wire _w930_ ;
	wire _w929_ ;
	wire _w928_ ;
	wire _w927_ ;
	wire _w926_ ;
	wire _w925_ ;
	wire _w924_ ;
	wire _w923_ ;
	wire _w922_ ;
	wire _w921_ ;
	wire _w920_ ;
	wire _w919_ ;
	wire _w918_ ;
	wire _w917_ ;
	wire _w916_ ;
	wire _w915_ ;
	wire _w914_ ;
	wire _w913_ ;
	wire _w912_ ;
	wire _w911_ ;
	wire _w910_ ;
	wire _w909_ ;
	wire _w908_ ;
	wire _w907_ ;
	wire _w906_ ;
	wire _w905_ ;
	wire _w904_ ;
	wire _w903_ ;
	wire _w902_ ;
	wire _w901_ ;
	wire _w900_ ;
	wire _w899_ ;
	wire _w898_ ;
	wire _w897_ ;
	wire _w896_ ;
	wire _w895_ ;
	wire _w894_ ;
	wire _w893_ ;
	wire _w892_ ;
	wire _w891_ ;
	wire _w890_ ;
	wire _w889_ ;
	wire _w888_ ;
	wire _w887_ ;
	wire _w886_ ;
	wire _w885_ ;
	wire _w884_ ;
	wire _w883_ ;
	wire _w882_ ;
	wire _w881_ ;
	wire _w880_ ;
	wire _w879_ ;
	wire _w878_ ;
	wire _w877_ ;
	wire _w876_ ;
	wire _w875_ ;
	wire _w874_ ;
	wire _w873_ ;
	wire _w872_ ;
	wire _w871_ ;
	wire _w870_ ;
	wire _w869_ ;
	wire _w868_ ;
	wire _w867_ ;
	wire _w866_ ;
	wire _w865_ ;
	wire _w864_ ;
	wire _w863_ ;
	wire _w862_ ;
	wire _w861_ ;
	wire _w860_ ;
	wire _w859_ ;
	wire _w858_ ;
	wire _w857_ ;
	wire _w856_ ;
	wire _w855_ ;
	wire _w854_ ;
	wire _w853_ ;
	wire _w852_ ;
	wire _w851_ ;
	wire _w850_ ;
	wire _w849_ ;
	wire _w848_ ;
	wire _w847_ ;
	wire _w846_ ;
	wire _w845_ ;
	wire _w844_ ;
	wire _w843_ ;
	wire _w842_ ;
	wire _w841_ ;
	wire _w840_ ;
	wire _w839_ ;
	wire _w838_ ;
	wire _w837_ ;
	wire _w836_ ;
	wire _w835_ ;
	wire _w834_ ;
	wire _w833_ ;
	wire _w832_ ;
	wire _w831_ ;
	wire _w830_ ;
	wire _w829_ ;
	wire _w828_ ;
	wire _w827_ ;
	wire _w826_ ;
	wire _w825_ ;
	wire _w824_ ;
	wire _w823_ ;
	wire _w822_ ;
	wire _w821_ ;
	wire _w820_ ;
	wire _w819_ ;
	wire _w818_ ;
	wire _w817_ ;
	wire _w816_ ;
	wire _w815_ ;
	wire _w814_ ;
	wire _w813_ ;
	wire _w812_ ;
	wire _w811_ ;
	wire _w810_ ;
	wire _w809_ ;
	wire _w808_ ;
	wire _w807_ ;
	wire _w806_ ;
	wire _w805_ ;
	wire _w804_ ;
	wire _w803_ ;
	wire _w802_ ;
	wire _w801_ ;
	wire _w800_ ;
	wire _w799_ ;
	wire _w798_ ;
	wire _w797_ ;
	wire _w796_ ;
	wire _w795_ ;
	wire _w794_ ;
	wire _w793_ ;
	wire _w792_ ;
	wire _w791_ ;
	wire _w790_ ;
	wire _w789_ ;
	wire _w788_ ;
	wire _w787_ ;
	wire _w786_ ;
	wire _w785_ ;
	wire _w784_ ;
	wire _w783_ ;
	wire _w782_ ;
	wire _w781_ ;
	wire _w780_ ;
	wire _w779_ ;
	wire _w778_ ;
	wire _w777_ ;
	wire _w776_ ;
	wire _w775_ ;
	wire _w774_ ;
	wire _w773_ ;
	wire _w772_ ;
	wire _w771_ ;
	wire _w770_ ;
	wire _w769_ ;
	wire _w768_ ;
	wire _w767_ ;
	wire _w766_ ;
	wire _w765_ ;
	wire _w764_ ;
	wire _w763_ ;
	wire _w762_ ;
	wire _w761_ ;
	wire _w760_ ;
	wire _w759_ ;
	wire _w758_ ;
	wire _w757_ ;
	wire _w756_ ;
	wire _w755_ ;
	wire _w754_ ;
	wire _w753_ ;
	wire _w752_ ;
	wire _w751_ ;
	wire _w750_ ;
	wire _w749_ ;
	wire _w464_ ;
	wire _w463_ ;
	wire _w462_ ;
	wire _w461_ ;
	wire _w460_ ;
	wire _w459_ ;
	wire _w458_ ;
	wire _w457_ ;
	wire _w456_ ;
	wire _w455_ ;
	wire _w454_ ;
	wire _w453_ ;
	wire _w452_ ;
	wire _w451_ ;
	wire _w450_ ;
	wire _w449_ ;
	wire _w448_ ;
	wire _w447_ ;
	wire _w446_ ;
	wire _w445_ ;
	wire _w444_ ;
	wire _w443_ ;
	wire _w442_ ;
	wire _w441_ ;
	wire _w440_ ;
	wire _w439_ ;
	wire _w438_ ;
	wire _w437_ ;
	wire _w436_ ;
	wire _w435_ ;
	wire _w434_ ;
	wire _w433_ ;
	wire _w432_ ;
	wire _w431_ ;
	wire _w430_ ;
	wire _w429_ ;
	wire _w428_ ;
	wire _w427_ ;
	wire _w426_ ;
	wire _w425_ ;
	wire _w424_ ;
	wire _w423_ ;
	wire _w422_ ;
	wire _w421_ ;
	wire _w420_ ;
	wire _w419_ ;
	wire _w418_ ;
	wire _w417_ ;
	wire _w416_ ;
	wire _w415_ ;
	wire _w414_ ;
	wire _w413_ ;
	wire _w412_ ;
	wire _w411_ ;
	wire _w410_ ;
	wire _w409_ ;
	wire _w408_ ;
	wire _w407_ ;
	wire _w406_ ;
	wire _w405_ ;
	wire _w404_ ;
	wire _w403_ ;
	wire _w402_ ;
	wire _w401_ ;
	wire _w400_ ;
	wire _w399_ ;
	wire _w398_ ;
	wire _w397_ ;
	wire _w396_ ;
	wire _w395_ ;
	wire _w394_ ;
	wire _w393_ ;
	wire _w392_ ;
	wire _w391_ ;
	wire _w390_ ;
	wire _w389_ ;
	wire _w388_ ;
	wire _w387_ ;
	wire _w386_ ;
	wire _w385_ ;
	wire _w384_ ;
	wire _w383_ ;
	wire _w382_ ;
	wire _w381_ ;
	wire _w380_ ;
	wire _w379_ ;
	wire _w378_ ;
	wire _w377_ ;
	wire _w376_ ;
	wire _w375_ ;
	wire _w374_ ;
	wire _w373_ ;
	wire _w372_ ;
	wire _w371_ ;
	wire _w370_ ;
	wire _w369_ ;
	wire _w368_ ;
	wire _w367_ ;
	wire _w366_ ;
	wire _w365_ ;
	wire _w364_ ;
	wire _w363_ ;
	wire _w362_ ;
	wire _w361_ ;
	wire _w360_ ;
	wire _w359_ ;
	wire _w358_ ;
	wire _w357_ ;
	wire _w356_ ;
	wire _w355_ ;
	wire _w354_ ;
	wire _w353_ ;
	wire _w352_ ;
	wire _w351_ ;
	wire _w350_ ;
	wire _w349_ ;
	wire _w348_ ;
	wire _w347_ ;
	wire _w346_ ;
	wire _w345_ ;
	wire _w344_ ;
	wire _w343_ ;
	wire _w342_ ;
	wire _w341_ ;
	wire _w340_ ;
	wire _w339_ ;
	wire _w338_ ;
	wire _w337_ ;
	wire _w336_ ;
	wire _w335_ ;
	wire _w266_ ;
	wire _w265_ ;
	wire _w264_ ;
	wire _w262_ ;
	wire _w261_ ;
	wire _w260_ ;
	wire _w259_ ;
	wire _w258_ ;
	wire _w257_ ;
	wire _w256_ ;
	wire _w255_ ;
	wire _w254_ ;
	wire _w253_ ;
	wire _w252_ ;
	wire _w251_ ;
	wire _w250_ ;
	wire _w249_ ;
	wire _w248_ ;
	wire _w247_ ;
	wire _w246_ ;
	wire _w245_ ;
	wire _w244_ ;
	wire _w243_ ;
	wire _w242_ ;
	wire _w241_ ;
	wire _w240_ ;
	wire _w239_ ;
	wire _w238_ ;
	wire _w237_ ;
	wire _w220_ ;
	wire _w219_ ;
	wire _w218_ ;
	wire _w217_ ;
	wire _w216_ ;
	wire _w215_ ;
	wire _w214_ ;
	wire _w213_ ;
	wire _w212_ ;
	wire _w211_ ;
	wire _w210_ ;
	wire _w209_ ;
	wire _w263_ ;
	wire _w281_ ;
	wire _w230_ ;
	wire _w221_ ;
	wire _w222_ ;
	wire _w223_ ;
	wire _w224_ ;
	wire _w225_ ;
	wire _w226_ ;
	wire _w227_ ;
	wire _w228_ ;
	wire _w229_ ;
	wire _w231_ ;
	wire _w232_ ;
	wire _w233_ ;
	wire _w234_ ;
	wire _w235_ ;
	wire _w236_ ;
	wire _w267_ ;
	wire _w268_ ;
	wire _w269_ ;
	wire _w270_ ;
	wire _w271_ ;
	wire _w272_ ;
	wire _w273_ ;
	wire _w274_ ;
	wire _w275_ ;
	wire _w276_ ;
	wire _w277_ ;
	wire _w278_ ;
	wire _w279_ ;
	wire _w280_ ;
	wire _w282_ ;
	wire _w283_ ;
	wire _w27_ ;
	wire _w568_ ;
	wire _w284_ ;
	wire _w285_ ;
	wire _w286_ ;
	wire _w287_ ;
	wire _w288_ ;
	wire _w289_ ;
	wire _w290_ ;
	wire _w291_ ;
	wire _w292_ ;
	wire _w293_ ;
	wire _w294_ ;
	wire _w295_ ;
	wire _w296_ ;
	wire _w297_ ;
	wire _w298_ ;
	wire _w299_ ;
	wire _w300_ ;
	wire _w301_ ;
	wire _w302_ ;
	wire _w303_ ;
	wire _w304_ ;
	wire _w305_ ;
	wire _w306_ ;
	wire _w307_ ;
	wire _w308_ ;
	wire _w309_ ;
	wire _w310_ ;
	wire _w311_ ;
	wire _w312_ ;
	wire _w313_ ;
	wire _w314_ ;
	wire _w315_ ;
	wire _w316_ ;
	wire _w317_ ;
	wire _w318_ ;
	wire _w319_ ;
	wire _w320_ ;
	wire _w321_ ;
	wire _w322_ ;
	wire _w323_ ;
	wire _w324_ ;
	wire _w325_ ;
	wire _w326_ ;
	wire _w327_ ;
	wire _w328_ ;
	wire _w329_ ;
	wire _w330_ ;
	wire _w331_ ;
	wire _w332_ ;
	wire _w333_ ;
	wire _w334_ ;
	wire _w465_ ;
	wire _w466_ ;
	wire _w467_ ;
	wire _w468_ ;
	wire _w469_ ;
	wire _w470_ ;
	wire _w471_ ;
	wire _w472_ ;
	wire _w473_ ;
	wire _w474_ ;
	wire _w475_ ;
	wire _w476_ ;
	wire _w477_ ;
	wire _w478_ ;
	wire _w479_ ;
	wire _w480_ ;
	wire _w481_ ;
	wire _w482_ ;
	wire _w483_ ;
	wire _w484_ ;
	wire _w485_ ;
	wire _w486_ ;
	wire _w487_ ;
	wire _w488_ ;
	wire _w489_ ;
	wire _w490_ ;
	wire _w491_ ;
	wire _w492_ ;
	wire _w493_ ;
	wire _w494_ ;
	wire _w495_ ;
	wire _w496_ ;
	wire _w497_ ;
	wire _w498_ ;
	wire _w499_ ;
	wire _w500_ ;
	wire _w501_ ;
	wire _w502_ ;
	wire _w503_ ;
	wire _w504_ ;
	wire _w505_ ;
	wire _w506_ ;
	wire _w507_ ;
	wire _w508_ ;
	wire _w509_ ;
	wire _w510_ ;
	wire _w511_ ;
	wire _w512_ ;
	wire _w513_ ;
	wire _w514_ ;
	wire _w515_ ;
	wire _w516_ ;
	wire _w517_ ;
	wire _w518_ ;
	wire _w519_ ;
	wire _w520_ ;
	wire _w521_ ;
	wire _w522_ ;
	wire _w523_ ;
	wire _w524_ ;
	wire _w525_ ;
	wire _w526_ ;
	wire _w527_ ;
	wire _w528_ ;
	wire _w529_ ;
	wire _w530_ ;
	wire _w531_ ;
	wire _w532_ ;
	wire _w533_ ;
	wire _w534_ ;
	wire _w535_ ;
	wire _w536_ ;
	wire _w537_ ;
	wire _w538_ ;
	wire _w539_ ;
	wire _w540_ ;
	wire _w541_ ;
	wire _w542_ ;
	wire _w543_ ;
	wire _w544_ ;
	wire _w545_ ;
	wire _w546_ ;
	wire _w547_ ;
	wire _w548_ ;
	wire _w549_ ;
	wire _w550_ ;
	wire _w551_ ;
	wire _w552_ ;
	wire _w553_ ;
	wire _w554_ ;
	wire _w555_ ;
	wire _w556_ ;
	wire _w557_ ;
	wire _w558_ ;
	wire _w559_ ;
	wire _w560_ ;
	wire _w561_ ;
	wire _w562_ ;
	wire _w563_ ;
	wire _w564_ ;
	wire _w565_ ;
	wire _w566_ ;
	wire _w567_ ;
	wire _w569_ ;
	wire _w570_ ;
	wire _w571_ ;
	wire _w572_ ;
	wire _w573_ ;
	wire _w574_ ;
	wire _w575_ ;
	wire _w576_ ;
	wire _w577_ ;
	wire _w578_ ;
	wire _w579_ ;
	wire _w580_ ;
	wire _w581_ ;
	wire _w582_ ;
	wire _w583_ ;
	wire _w584_ ;
	wire _w585_ ;
	wire _w586_ ;
	wire _w587_ ;
	wire _w588_ ;
	wire _w589_ ;
	wire _w590_ ;
	wire _w591_ ;
	wire _w592_ ;
	wire _w593_ ;
	wire _w594_ ;
	wire _w595_ ;
	wire _w596_ ;
	wire _w597_ ;
	wire _w598_ ;
	wire _w599_ ;
	wire _w600_ ;
	wire _w601_ ;
	wire _w602_ ;
	wire _w603_ ;
	wire _w604_ ;
	wire _w605_ ;
	wire _w606_ ;
	wire _w607_ ;
	wire _w608_ ;
	wire _w609_ ;
	wire _w610_ ;
	wire _w611_ ;
	wire _w612_ ;
	wire _w613_ ;
	wire _w614_ ;
	wire _w615_ ;
	wire _w616_ ;
	wire _w617_ ;
	wire _w618_ ;
	wire _w619_ ;
	wire _w620_ ;
	wire _w621_ ;
	wire _w622_ ;
	wire _w623_ ;
	wire _w624_ ;
	wire _w625_ ;
	wire _w626_ ;
	wire _w627_ ;
	wire _w628_ ;
	wire _w629_ ;
	wire _w630_ ;
	wire _w631_ ;
	wire _w632_ ;
	wire _w633_ ;
	wire _w634_ ;
	wire _w635_ ;
	wire _w636_ ;
	wire _w637_ ;
	wire _w638_ ;
	wire _w639_ ;
	wire _w640_ ;
	wire _w641_ ;
	wire _w642_ ;
	wire _w643_ ;
	wire _w644_ ;
	wire _w645_ ;
	wire _w646_ ;
	wire _w647_ ;
	wire _w648_ ;
	wire _w649_ ;
	wire _w650_ ;
	wire _w651_ ;
	wire _w652_ ;
	wire _w653_ ;
	wire _w654_ ;
	wire _w655_ ;
	wire _w656_ ;
	wire _w657_ ;
	wire _w658_ ;
	wire _w659_ ;
	wire _w660_ ;
	wire _w661_ ;
	wire _w662_ ;
	wire _w663_ ;
	wire _w664_ ;
	wire _w665_ ;
	wire _w666_ ;
	wire _w667_ ;
	wire _w668_ ;
	wire _w669_ ;
	wire _w670_ ;
	wire _w671_ ;
	wire _w672_ ;
	wire _w673_ ;
	wire _w674_ ;
	wire _w675_ ;
	wire _w676_ ;
	wire _w677_ ;
	wire _w678_ ;
	wire _w679_ ;
	wire _w680_ ;
	wire _w681_ ;
	wire _w682_ ;
	wire _w683_ ;
	wire _w684_ ;
	wire _w685_ ;
	wire _w686_ ;
	wire _w687_ ;
	wire _w688_ ;
	wire _w689_ ;
	wire _w690_ ;
	wire _w691_ ;
	wire _w692_ ;
	wire _w693_ ;
	wire _w694_ ;
	wire _w695_ ;
	wire _w696_ ;
	wire _w697_ ;
	wire _w698_ ;
	wire _w699_ ;
	wire _w700_ ;
	wire _w701_ ;
	wire _w702_ ;
	wire _w703_ ;
	wire _w704_ ;
	wire _w705_ ;
	wire _w706_ ;
	wire _w707_ ;
	wire _w708_ ;
	wire _w709_ ;
	wire _w710_ ;
	wire _w711_ ;
	wire _w712_ ;
	wire _w713_ ;
	wire _w714_ ;
	wire _w715_ ;
	wire _w716_ ;
	wire _w717_ ;
	wire _w718_ ;
	wire _w719_ ;
	wire _w720_ ;
	wire _w721_ ;
	wire _w722_ ;
	wire _w723_ ;
	wire _w724_ ;
	wire _w725_ ;
	wire _w726_ ;
	wire _w727_ ;
	wire _w728_ ;
	wire _w729_ ;
	wire _w730_ ;
	wire _w731_ ;
	wire _w732_ ;
	wire _w733_ ;
	wire _w734_ ;
	wire _w735_ ;
	wire _w736_ ;
	wire _w737_ ;
	wire _w738_ ;
	wire _w739_ ;
	wire _w740_ ;
	wire _w741_ ;
	wire _w742_ ;
	wire _w743_ ;
	wire _w744_ ;
	wire _w745_ ;
	wire _w746_ ;
	wire _w747_ ;
	wire _w748_ ;
	LUT1 #(
		.INIT('h1)
	) name0 (
		\15(4)_pad ,
		_w27_
	);
	LUT3 #(
		.INIT('h27)
	) name1 (
		\18(5)_pad ,
		\195(118)_pad ,
		\94(49)_pad ,
		_w209_
	);
	LUT3 #(
		.INIT('h8d)
	) name2 (
		\18(5)_pad ,
		\536(222)_pad ,
		\59(22)_pad ,
		_w210_
	);
	LUT3 #(
		.INIT('h27)
	) name3 (
		\18(5)_pad ,
		\196(119)_pad ,
		\97(50)_pad ,
		_w211_
	);
	LUT3 #(
		.INIT('h8d)
	) name4 (
		\18(5)_pad ,
		\538(224)_pad ,
		\78(37)_pad ,
		_w212_
	);
	LUT4 #(
		.INIT('h0777)
	) name5 (
		_w209_,
		_w210_,
		_w211_,
		_w212_,
		_w213_
	);
	LUT3 #(
		.INIT('h27)
	) name6 (
		\18(5)_pad ,
		\193(116)_pad ,
		\47(14)_pad ,
		_w214_
	);
	LUT3 #(
		.INIT('h8d)
	) name7 (
		\18(5)_pad ,
		\532(218)_pad ,
		\80(39)_pad ,
		_w215_
	);
	LUT2 #(
		.INIT('h1)
	) name8 (
		_w214_,
		_w215_,
		_w216_
	);
	LUT3 #(
		.INIT('h1d)
	) name9 (
		\121(62)_pad ,
		\18(5)_pad ,
		\194(117)_pad ,
		_w217_
	);
	LUT3 #(
		.INIT('h8d)
	) name10 (
		\18(5)_pad ,
		\534(220)_pad ,
		\81(40)_pad ,
		_w218_
	);
	LUT4 #(
		.INIT('heee0)
	) name11 (
		_w209_,
		_w210_,
		_w217_,
		_w218_,
		_w219_
	);
	LUT3 #(
		.INIT('h10)
	) name12 (
		_w213_,
		_w216_,
		_w219_,
		_w220_
	);
	LUT3 #(
		.INIT('h27)
	) name13 (
		\18(5)_pad ,
		\205(128)_pad ,
		\23(6)_pad ,
		_w221_
	);
	LUT3 #(
		.INIT('h8d)
	) name14 (
		\18(5)_pad ,
		\554(240)_pad ,
		\75(34)_pad ,
		_w222_
	);
	LUT3 #(
		.INIT('h1d)
	) name15 (
		\103(52)_pad ,
		\18(5)_pad ,
		\204(127)_pad ,
		_w223_
	);
	LUT3 #(
		.INIT('h8d)
	) name16 (
		\18(5)_pad ,
		\552(238)_pad ,
		\73(32)_pad ,
		_w224_
	);
	LUT4 #(
		.INIT('h0777)
	) name17 (
		_w221_,
		_w222_,
		_w223_,
		_w224_,
		_w225_
	);
	LUT3 #(
		.INIT('h27)
	) name18 (
		\18(5)_pad ,
		\206(129)_pad ,
		\26(7)_pad ,
		_w226_
	);
	LUT3 #(
		.INIT('h8d)
	) name19 (
		\18(5)_pad ,
		\556(242)_pad ,
		\76(35)_pad ,
		_w227_
	);
	LUT4 #(
		.INIT('heee0)
	) name20 (
		_w221_,
		_w222_,
		_w226_,
		_w227_,
		_w228_
	);
	LUT3 #(
		.INIT('h40)
	) name21 (
		\18(5)_pad ,
		\41(12)_pad ,
		\70(31)_pad ,
		_w229_
	);
	LUT4 #(
		.INIT('hfe00)
	) name22 (
		\18(5)_pad ,
		\41(12)_pad ,
		\70(31)_pad ,
		\89(48)_pad ,
		_w230_
	);
	LUT3 #(
		.INIT('h27)
	) name23 (
		\18(5)_pad ,
		\207(130)_pad ,
		\29(8)_pad ,
		_w231_
	);
	LUT3 #(
		.INIT('h8d)
	) name24 (
		\18(5)_pad ,
		\558(244)_pad ,
		\74(33)_pad ,
		_w232_
	);
	LUT4 #(
		.INIT('h1110)
	) name25 (
		_w229_,
		_w230_,
		_w231_,
		_w232_,
		_w233_
	);
	LUT4 #(
		.INIT('h0777)
	) name26 (
		_w226_,
		_w227_,
		_w231_,
		_w232_,
		_w234_
	);
	LUT4 #(
		.INIT('hd5dd)
	) name27 (
		_w225_,
		_w228_,
		_w233_,
		_w234_,
		_w235_
	);
	LUT3 #(
		.INIT('h1d)
	) name28 (
		\124(63)_pad ,
		\18(5)_pad ,
		\201(124)_pad ,
		_w236_
	);
	LUT3 #(
		.INIT('h8d)
	) name29 (
		\18(5)_pad ,
		\546(232)_pad ,
		\55(18)_pad ,
		_w237_
	);
	LUT3 #(
		.INIT('h1d)
	) name30 (
		\127(64)_pad ,
		\18(5)_pad ,
		\202(125)_pad ,
		_w238_
	);
	LUT3 #(
		.INIT('hb1)
	) name31 (
		\18(5)_pad ,
		\54(17)_pad ,
		\548(234)_pad ,
		_w239_
	);
	LUT4 #(
		.INIT('h0007)
	) name32 (
		_w236_,
		_w237_,
		_w238_,
		_w239_,
		_w240_
	);
	LUT3 #(
		.INIT('h1d)
	) name33 (
		\100(51)_pad ,
		\18(5)_pad ,
		\200(123)_pad ,
		_w241_
	);
	LUT3 #(
		.INIT('h8d)
	) name34 (
		\18(5)_pad ,
		\544(230)_pad ,
		\56(19)_pad ,
		_w242_
	);
	LUT4 #(
		.INIT('heee0)
	) name35 (
		_w236_,
		_w237_,
		_w241_,
		_w242_,
		_w243_
	);
	LUT3 #(
		.INIT('h1d)
	) name36 (
		\130(65)_pad ,
		\18(5)_pad ,
		\203(126)_pad ,
		_w244_
	);
	LUT3 #(
		.INIT('hb1)
	) name37 (
		\18(5)_pad ,
		\53(16)_pad ,
		\550(236)_pad ,
		_w245_
	);
	LUT4 #(
		.INIT('heee0)
	) name38 (
		_w223_,
		_w224_,
		_w244_,
		_w245_,
		_w246_
	);
	LUT3 #(
		.INIT('h40)
	) name39 (
		_w240_,
		_w243_,
		_w246_,
		_w247_
	);
	LUT4 #(
		.INIT('h0777)
	) name40 (
		_w236_,
		_w237_,
		_w238_,
		_w239_,
		_w248_
	);
	LUT4 #(
		.INIT('h0eee)
	) name41 (
		_w238_,
		_w239_,
		_w244_,
		_w245_,
		_w249_
	);
	LUT4 #(
		.INIT('h0444)
	) name42 (
		_w240_,
		_w243_,
		_w248_,
		_w249_,
		_w250_
	);
	LUT3 #(
		.INIT('h1d)
	) name43 (
		\118(61)_pad ,
		\18(5)_pad ,
		\187(110)_pad ,
		_w251_
	);
	LUT3 #(
		.INIT('h8d)
	) name44 (
		\18(5)_pad ,
		\522(226)_pad ,
		\77(36)_pad ,
		_w252_
	);
	LUT4 #(
		.INIT('h0777)
	) name45 (
		_w241_,
		_w242_,
		_w251_,
		_w252_,
		_w253_
	);
	LUT4 #(
		.INIT('h0700)
	) name46 (
		_w235_,
		_w247_,
		_w250_,
		_w253_,
		_w254_
	);
	LUT4 #(
		.INIT('heee0)
	) name47 (
		_w211_,
		_w212_,
		_w251_,
		_w252_,
		_w255_
	);
	LUT3 #(
		.INIT('h40)
	) name48 (
		_w216_,
		_w219_,
		_w255_,
		_w256_
	);
	LUT3 #(
		.INIT('h45)
	) name49 (
		_w220_,
		_w254_,
		_w256_,
		_w257_
	);
	LUT4 #(
		.INIT('he888)
	) name50 (
		_w214_,
		_w215_,
		_w217_,
		_w218_,
		_w258_
	);
	LUT3 #(
		.INIT('h27)
	) name51 (
		\18(5)_pad ,
		\189(112)_pad ,
		\66(29)_pad ,
		_w259_
	);
	LUT3 #(
		.INIT('h8d)
	) name52 (
		\18(5)_pad ,
		\524(210)_pad ,
		\62(25)_pad ,
		_w260_
	);
	LUT2 #(
		.INIT('h8)
	) name53 (
		_w259_,
		_w260_,
		_w261_
	);
	LUT3 #(
		.INIT('h27)
	) name54 (
		\18(5)_pad ,
		\191(114)_pad ,
		\32(9)_pad ,
		_w262_
	);
	LUT3 #(
		.INIT('h8d)
	) name55 (
		\18(5)_pad ,
		\528(214)_pad ,
		\60(23)_pad ,
		_w263_
	);
	LUT4 #(
		.INIT('h0777)
	) name56 (
		_w259_,
		_w260_,
		_w262_,
		_w263_,
		_w264_
	);
	LUT3 #(
		.INIT('h27)
	) name57 (
		\18(5)_pad ,
		\190(113)_pad ,
		\50(15)_pad ,
		_w265_
	);
	LUT3 #(
		.INIT('h8d)
	) name58 (
		\18(5)_pad ,
		\526(212)_pad ,
		\61(24)_pad ,
		_w266_
	);
	LUT4 #(
		.INIT('h0eee)
	) name59 (
		_w262_,
		_w263_,
		_w265_,
		_w266_,
		_w267_
	);
	LUT4 #(
		.INIT('heee0)
	) name60 (
		_w259_,
		_w260_,
		_w265_,
		_w266_,
		_w268_
	);
	LUT3 #(
		.INIT('h27)
	) name61 (
		\18(5)_pad ,
		\192(115)_pad ,
		\35(10)_pad ,
		_w269_
	);
	LUT3 #(
		.INIT('h8d)
	) name62 (
		\18(5)_pad ,
		\530(216)_pad ,
		\79(38)_pad ,
		_w270_
	);
	LUT2 #(
		.INIT('h1)
	) name63 (
		_w269_,
		_w270_,
		_w271_
	);
	LUT2 #(
		.INIT('h6)
	) name64 (
		_w269_,
		_w270_,
		_w272_
	);
	LUT4 #(
		.INIT('h8000)
	) name65 (
		_w264_,
		_w267_,
		_w268_,
		_w272_,
		_w273_
	);
	LUT2 #(
		.INIT('h4)
	) name66 (
		_w258_,
		_w273_,
		_w274_
	);
	LUT4 #(
		.INIT('h4500)
	) name67 (
		_w220_,
		_w254_,
		_w256_,
		_w274_,
		_w275_
	);
	LUT4 #(
		.INIT('h8000)
	) name68 (
		_w264_,
		_w267_,
		_w268_,
		_w271_,
		_w276_
	);
	LUT4 #(
		.INIT('h0111)
	) name69 (
		_w262_,
		_w263_,
		_w265_,
		_w266_,
		_w277_
	);
	LUT3 #(
		.INIT('h51)
	) name70 (
		_w261_,
		_w268_,
		_w277_,
		_w278_
	);
	LUT2 #(
		.INIT('h1)
	) name71 (
		_w276_,
		_w278_,
		_w279_
	);
	LUT2 #(
		.INIT('hb)
	) name72 (
		_w275_,
		_w279_,
		_w280_
	);
	LUT2 #(
		.INIT('h8)
	) name73 (
		\12(3)_pad ,
		\9(2)_pad ,
		_w281_
	);
	LUT4 #(
		.INIT('h45cf)
	) name74 (
		\12(3)_pad ,
		\167(90)_pad ,
		\18(5)_pad ,
		\9(2)_pad ,
		_w282_
	);
	LUT3 #(
		.INIT('hd1)
	) name75 (
		\112(57)_pad ,
		\18(5)_pad ,
		\444(282)_pad ,
		_w283_
	);
	LUT4 #(
		.INIT('h45cf)
	) name76 (
		\12(3)_pad ,
		\168(91)_pad ,
		\18(5)_pad ,
		\9(2)_pad ,
		_w284_
	);
	LUT3 #(
		.INIT('h8d)
	) name77 (
		\18(5)_pad ,
		\446(393)_pad ,
		\87(46)_pad ,
		_w285_
	);
	LUT4 #(
		.INIT('h9009)
	) name78 (
		_w282_,
		_w283_,
		_w284_,
		_w285_,
		_w286_
	);
	LUT2 #(
		.INIT('h4)
	) name79 (
		\169(92)_pad ,
		\18(5)_pad ,
		_w287_
	);
	LUT4 #(
		.INIT('h45cf)
	) name80 (
		\12(3)_pad ,
		\169(92)_pad ,
		\18(5)_pad ,
		\9(2)_pad ,
		_w288_
	);
	LUT3 #(
		.INIT('hd1)
	) name81 (
		\111(56)_pad ,
		\18(5)_pad ,
		\448(284)_pad ,
		_w289_
	);
	LUT2 #(
		.INIT('h2)
	) name82 (
		_w288_,
		_w289_,
		_w290_
	);
	LUT2 #(
		.INIT('h9)
	) name83 (
		_w288_,
		_w289_,
		_w291_
	);
	LUT4 #(
		.INIT('h0700)
	) name84 (
		\1455(166)_pad ,
		\2204(174)_pad ,
		\38(11)_pad ,
		\4528(206)_pad ,
		_w292_
	);
	LUT2 #(
		.INIT('h4)
	) name85 (
		\166(89)_pad ,
		\18(5)_pad ,
		_w293_
	);
	LUT4 #(
		.INIT('h45cf)
	) name86 (
		\12(3)_pad ,
		\166(89)_pad ,
		\18(5)_pad ,
		\9(2)_pad ,
		_w294_
	);
	LUT3 #(
		.INIT('h8d)
	) name87 (
		\18(5)_pad ,
		\442(280)_pad ,
		\88(47)_pad ,
		_w295_
	);
	LUT4 #(
		.INIT('he0f0)
	) name88 (
		\1455(166)_pad ,
		\2204(174)_pad ,
		\38(11)_pad ,
		\4528(206)_pad ,
		_w296_
	);
	LUT4 #(
		.INIT('h0045)
	) name89 (
		_w292_,
		_w294_,
		_w295_,
		_w296_,
		_w297_
	);
	LUT2 #(
		.INIT('h2)
	) name90 (
		_w294_,
		_w295_,
		_w298_
	);
	LUT3 #(
		.INIT('hd1)
	) name91 (
		\113(58)_pad ,
		\18(5)_pad ,
		\436(286)_pad ,
		_w299_
	);
	LUT4 #(
		.INIT('h54aa)
	) name92 (
		_w281_,
		_w293_,
		_w295_,
		_w299_,
		_w300_
	);
	LUT4 #(
		.INIT('h8000)
	) name93 (
		_w286_,
		_w291_,
		_w297_,
		_w300_,
		_w301_
	);
	LUT4 #(
		.INIT('h00fb)
	) name94 (
		_w294_,
		_w295_,
		_w296_,
		_w292_,
		_w302_
	);
	LUT4 #(
		.INIT('h22b2)
	) name95 (
		_w282_,
		_w283_,
		_w284_,
		_w285_,
		_w303_
	);
	LUT4 #(
		.INIT('h0007)
	) name96 (
		_w286_,
		_w290_,
		_w298_,
		_w303_,
		_w304_
	);
	LUT4 #(
		.INIT('h0014)
	) name97 (
		_w281_,
		_w287_,
		_w289_,
		_w299_,
		_w305_
	);
	LUT3 #(
		.INIT('h13)
	) name98 (
		_w286_,
		_w296_,
		_w305_,
		_w306_
	);
	LUT3 #(
		.INIT('h2a)
	) name99 (
		_w302_,
		_w304_,
		_w306_,
		_w307_
	);
	LUT4 #(
		.INIT('h5111)
	) name100 (
		_w301_,
		_w302_,
		_w304_,
		_w306_,
		_w308_
	);
	LUT4 #(
		.INIT('h45cf)
	) name101 (
		\12(3)_pad ,
		\177(100)_pad ,
		\18(5)_pad ,
		\9(2)_pad ,
		_w309_
	);
	LUT3 #(
		.INIT('h8d)
	) name102 (
		\18(5)_pad ,
		\488(260)_pad ,
		\64(27)_pad ,
		_w310_
	);
	LUT3 #(
		.INIT('h35)
	) name103 (
		\135(68)_pad ,
		\178(101)_pad ,
		\18(5)_pad ,
		_w311_
	);
	LUT3 #(
		.INIT('h8d)
	) name104 (
		\18(5)_pad ,
		\490(263)_pad ,
		\85(44)_pad ,
		_w312_
	);
	LUT4 #(
		.INIT('hddd0)
	) name105 (
		_w309_,
		_w310_,
		_w311_,
		_w312_,
		_w313_
	);
	LUT4 #(
		.INIT('h45cf)
	) name106 (
		\12(3)_pad ,
		\175(98)_pad ,
		\18(5)_pad ,
		\9(2)_pad ,
		_w314_
	);
	LUT3 #(
		.INIT('h8d)
	) name107 (
		\18(5)_pad ,
		\484(256)_pad ,
		\86(45)_pad ,
		_w315_
	);
	LUT2 #(
		.INIT('h4)
	) name108 (
		_w314_,
		_w315_,
		_w316_
	);
	LUT4 #(
		.INIT('h45cf)
	) name109 (
		\12(3)_pad ,
		\176(99)_pad ,
		\18(5)_pad ,
		\9(2)_pad ,
		_w317_
	);
	LUT3 #(
		.INIT('h8d)
	) name110 (
		\18(5)_pad ,
		\486(258)_pad ,
		\63(26)_pad ,
		_w318_
	);
	LUT2 #(
		.INIT('h2)
	) name111 (
		_w317_,
		_w318_,
		_w319_
	);
	LUT4 #(
		.INIT('hbb0b)
	) name112 (
		_w314_,
		_w315_,
		_w317_,
		_w318_,
		_w320_
	);
	LUT3 #(
		.INIT('h35)
	) name113 (
		\144(71)_pad ,
		\179(102)_pad ,
		\18(5)_pad ,
		_w321_
	);
	LUT3 #(
		.INIT('h8d)
	) name114 (
		\18(5)_pad ,
		\492(265)_pad ,
		\84(43)_pad ,
		_w322_
	);
	LUT4 #(
		.INIT('h0777)
	) name115 (
		_w311_,
		_w312_,
		_w321_,
		_w322_,
		_w323_
	);
	LUT3 #(
		.INIT('h80)
	) name116 (
		_w313_,
		_w320_,
		_w323_,
		_w324_
	);
	LUT4 #(
		.INIT('h45cf)
	) name117 (
		\12(3)_pad ,
		\174(97)_pad ,
		\18(5)_pad ,
		\9(2)_pad ,
		_w325_
	);
	LUT3 #(
		.INIT('hd1)
	) name118 (
		\109(54)_pad ,
		\18(5)_pad ,
		\482(253)_pad ,
		_w326_
	);
	LUT4 #(
		.INIT('h45cf)
	) name119 (
		\12(3)_pad ,
		\173(96)_pad ,
		\18(5)_pad ,
		\9(2)_pad ,
		_w327_
	);
	LUT3 #(
		.INIT('hd1)
	) name120 (
		\110(55)_pad ,
		\18(5)_pad ,
		\480(250)_pad ,
		_w328_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name121 (
		_w325_,
		_w326_,
		_w327_,
		_w328_,
		_w329_
	);
	LUT2 #(
		.INIT('h2)
	) name122 (
		_w327_,
		_w328_,
		_w330_
	);
	LUT3 #(
		.INIT('h1d)
	) name123 (
		\138(69)_pad ,
		\18(5)_pad ,
		\180(103)_pad ,
		_w331_
	);
	LUT3 #(
		.INIT('h8d)
	) name124 (
		\18(5)_pad ,
		\494(267)_pad ,
		\83(42)_pad ,
		_w332_
	);
	LUT3 #(
		.INIT('h35)
	) name125 (
		\147(72)_pad ,
		\171(94)_pad ,
		\18(5)_pad ,
		_w333_
	);
	LUT3 #(
		.INIT('h8d)
	) name126 (
		\18(5)_pad ,
		\478(269)_pad ,
		\65(28)_pad ,
		_w334_
	);
	LUT4 #(
		.INIT('h0777)
	) name127 (
		_w331_,
		_w332_,
		_w333_,
		_w334_,
		_w335_
	);
	LUT3 #(
		.INIT('h20)
	) name128 (
		_w329_,
		_w330_,
		_w335_,
		_w336_
	);
	LUT2 #(
		.INIT('h1)
	) name129 (
		_w331_,
		_w332_,
		_w337_
	);
	LUT4 #(
		.INIT('heee0)
	) name130 (
		_w321_,
		_w322_,
		_w333_,
		_w334_,
		_w338_
	);
	LUT4 #(
		.INIT('hdd0d)
	) name131 (
		_w314_,
		_w315_,
		_w325_,
		_w326_,
		_w339_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name132 (
		_w309_,
		_w310_,
		_w317_,
		_w318_,
		_w340_
	);
	LUT4 #(
		.INIT('h4000)
	) name133 (
		_w337_,
		_w338_,
		_w339_,
		_w340_,
		_w341_
	);
	LUT4 #(
		.INIT('h8000)
	) name134 (
		_w273_,
		_w324_,
		_w336_,
		_w341_,
		_w342_
	);
	LUT2 #(
		.INIT('h4)
	) name135 (
		_w258_,
		_w342_,
		_w343_
	);
	LUT3 #(
		.INIT('h80)
	) name136 (
		_w324_,
		_w336_,
		_w341_,
		_w344_
	);
	LUT2 #(
		.INIT('h4)
	) name137 (
		_w279_,
		_w344_,
		_w345_
	);
	LUT4 #(
		.INIT('h4f04)
	) name138 (
		_w325_,
		_w326_,
		_w327_,
		_w328_,
		_w346_
	);
	LUT4 #(
		.INIT('he000)
	) name139 (
		_w321_,
		_w322_,
		_w331_,
		_w332_,
		_w347_
	);
	LUT4 #(
		.INIT('h008a)
	) name140 (
		_w323_,
		_w337_,
		_w338_,
		_w347_,
		_w348_
	);
	LUT2 #(
		.INIT('h2)
	) name141 (
		_w313_,
		_w319_,
		_w349_
	);
	LUT4 #(
		.INIT('h4f04)
	) name142 (
		_w309_,
		_w310_,
		_w317_,
		_w318_,
		_w350_
	);
	LUT2 #(
		.INIT('h1)
	) name143 (
		_w316_,
		_w350_,
		_w351_
	);
	LUT2 #(
		.INIT('h4)
	) name144 (
		_w330_,
		_w339_,
		_w352_
	);
	LUT4 #(
		.INIT('h4f00)
	) name145 (
		_w348_,
		_w349_,
		_w351_,
		_w352_,
		_w353_
	);
	LUT3 #(
		.INIT('h54)
	) name146 (
		_w307_,
		_w346_,
		_w353_,
		_w354_
	);
	LUT4 #(
		.INIT('h0700)
	) name147 (
		_w257_,
		_w343_,
		_w345_,
		_w354_,
		_w355_
	);
	LUT2 #(
		.INIT('h1)
	) name148 (
		_w308_,
		_w355_,
		_w356_
	);
	LUT4 #(
		.INIT('h45cf)
	) name149 (
		\12(3)_pad ,
		\155(78)_pad ,
		\18(5)_pad ,
		\9(2)_pad ,
		_w357_
	);
	LUT2 #(
		.INIT('h2)
	) name150 (
		\484(256)_pad ,
		_w357_,
		_w358_
	);
	LUT4 #(
		.INIT('h45cf)
	) name151 (
		\12(3)_pad ,
		\156(79)_pad ,
		\18(5)_pad ,
		\9(2)_pad ,
		_w359_
	);
	LUT2 #(
		.INIT('h9)
	) name152 (
		\486(258)_pad ,
		_w359_,
		_w360_
	);
	LUT4 #(
		.INIT('h8421)
	) name153 (
		\484(256)_pad ,
		\486(258)_pad ,
		_w357_,
		_w359_,
		_w361_
	);
	LUT3 #(
		.INIT('h35)
	) name154 (
		\147(72)_pad ,
		\151(74)_pad ,
		\18(5)_pad ,
		_w362_
	);
	LUT4 #(
		.INIT('h00ca)
	) name155 (
		\147(72)_pad ,
		\151(74)_pad ,
		\18(5)_pad ,
		\478(269)_pad ,
		_w363_
	);
	LUT4 #(
		.INIT('h3500)
	) name156 (
		\147(72)_pad ,
		\151(74)_pad ,
		\18(5)_pad ,
		\478(269)_pad ,
		_w364_
	);
	LUT4 #(
		.INIT('hca35)
	) name157 (
		\147(72)_pad ,
		\151(74)_pad ,
		\18(5)_pad ,
		\478(269)_pad ,
		_w365_
	);
	LUT3 #(
		.INIT('h35)
	) name158 (
		\144(71)_pad ,
		\159(82)_pad ,
		\18(5)_pad ,
		_w366_
	);
	LUT4 #(
		.INIT('h00ca)
	) name159 (
		\144(71)_pad ,
		\159(82)_pad ,
		\18(5)_pad ,
		\492(265)_pad ,
		_w367_
	);
	LUT4 #(
		.INIT('h3500)
	) name160 (
		\144(71)_pad ,
		\159(82)_pad ,
		\18(5)_pad ,
		\492(265)_pad ,
		_w368_
	);
	LUT4 #(
		.INIT('hca35)
	) name161 (
		\144(71)_pad ,
		\159(82)_pad ,
		\18(5)_pad ,
		\492(265)_pad ,
		_w369_
	);
	LUT3 #(
		.INIT('h35)
	) name162 (
		\138(69)_pad ,
		\160(83)_pad ,
		\18(5)_pad ,
		_w370_
	);
	LUT4 #(
		.INIT('h00ca)
	) name163 (
		\138(69)_pad ,
		\160(83)_pad ,
		\18(5)_pad ,
		\494(267)_pad ,
		_w371_
	);
	LUT4 #(
		.INIT('h3500)
	) name164 (
		\138(69)_pad ,
		\160(83)_pad ,
		\18(5)_pad ,
		\494(267)_pad ,
		_w372_
	);
	LUT4 #(
		.INIT('hca35)
	) name165 (
		\138(69)_pad ,
		\160(83)_pad ,
		\18(5)_pad ,
		\494(267)_pad ,
		_w373_
	);
	LUT3 #(
		.INIT('h80)
	) name166 (
		_w365_,
		_w369_,
		_w373_,
		_w374_
	);
	LUT3 #(
		.INIT('h35)
	) name167 (
		\135(68)_pad ,
		\158(81)_pad ,
		\18(5)_pad ,
		_w375_
	);
	LUT4 #(
		.INIT('h00ca)
	) name168 (
		\135(68)_pad ,
		\158(81)_pad ,
		\18(5)_pad ,
		\490(263)_pad ,
		_w376_
	);
	LUT4 #(
		.INIT('h3500)
	) name169 (
		\135(68)_pad ,
		\158(81)_pad ,
		\18(5)_pad ,
		\490(263)_pad ,
		_w377_
	);
	LUT4 #(
		.INIT('hca35)
	) name170 (
		\135(68)_pad ,
		\158(81)_pad ,
		\18(5)_pad ,
		\490(263)_pad ,
		_w378_
	);
	LUT4 #(
		.INIT('h45cf)
	) name171 (
		\12(3)_pad ,
		\157(80)_pad ,
		\18(5)_pad ,
		\9(2)_pad ,
		_w379_
	);
	LUT2 #(
		.INIT('h9)
	) name172 (
		\488(260)_pad ,
		_w379_,
		_w380_
	);
	LUT3 #(
		.INIT('h84)
	) name173 (
		\488(260)_pad ,
		_w378_,
		_w379_,
		_w381_
	);
	LUT4 #(
		.INIT('h45cf)
	) name174 (
		\12(3)_pad ,
		\154(77)_pad ,
		\18(5)_pad ,
		\9(2)_pad ,
		_w382_
	);
	LUT2 #(
		.INIT('h4)
	) name175 (
		\482(253)_pad ,
		_w382_,
		_w383_
	);
	LUT2 #(
		.INIT('h2)
	) name176 (
		\482(253)_pad ,
		_w382_,
		_w384_
	);
	LUT2 #(
		.INIT('h9)
	) name177 (
		\482(253)_pad ,
		_w382_,
		_w385_
	);
	LUT4 #(
		.INIT('h45cf)
	) name178 (
		\12(3)_pad ,
		\153(76)_pad ,
		\18(5)_pad ,
		\9(2)_pad ,
		_w386_
	);
	LUT2 #(
		.INIT('h2)
	) name179 (
		\480(250)_pad ,
		_w386_,
		_w387_
	);
	LUT2 #(
		.INIT('h9)
	) name180 (
		\480(250)_pad ,
		_w386_,
		_w388_
	);
	LUT4 #(
		.INIT('h8241)
	) name181 (
		\480(250)_pad ,
		\482(253)_pad ,
		_w382_,
		_w386_,
		_w389_
	);
	LUT4 #(
		.INIT('h8000)
	) name182 (
		_w361_,
		_w374_,
		_w381_,
		_w389_,
		_w390_
	);
	LUT4 #(
		.INIT('h0b02)
	) name183 (
		\494(267)_pad ,
		_w363_,
		_w367_,
		_w370_,
		_w391_
	);
	LUT4 #(
		.INIT('h0301)
	) name184 (
		\488(260)_pad ,
		_w368_,
		_w377_,
		_w379_,
		_w392_
	);
	LUT3 #(
		.INIT('h2b)
	) name185 (
		\488(260)_pad ,
		_w376_,
		_w379_,
		_w393_
	);
	LUT3 #(
		.INIT('hb0)
	) name186 (
		_w391_,
		_w392_,
		_w393_,
		_w394_
	);
	LUT4 #(
		.INIT('hc341)
	) name187 (
		\480(250)_pad ,
		\482(253)_pad ,
		_w382_,
		_w386_,
		_w395_
	);
	LUT2 #(
		.INIT('h8)
	) name188 (
		_w361_,
		_w395_,
		_w396_
	);
	LUT4 #(
		.INIT('h51f3)
	) name189 (
		\12(3)_pad ,
		\18(5)_pad ,
		\216(139)_pad ,
		\9(2)_pad ,
		_w397_
	);
	LUT2 #(
		.INIT('h4)
	) name190 (
		\448(284)_pad ,
		_w397_,
		_w398_
	);
	LUT4 #(
		.INIT('h51f3)
	) name191 (
		\12(3)_pad ,
		\18(5)_pad ,
		\209(132)_pad ,
		\9(2)_pad ,
		_w399_
	);
	LUT2 #(
		.INIT('h4)
	) name192 (
		\436(286)_pad ,
		_w399_,
		_w400_
	);
	LUT4 #(
		.INIT('h8acf)
	) name193 (
		\436(286)_pad ,
		\448(284)_pad ,
		_w397_,
		_w399_,
		_w401_
	);
	LUT4 #(
		.INIT('h51f3)
	) name194 (
		\12(3)_pad ,
		\18(5)_pad ,
		\215(138)_pad ,
		\9(2)_pad ,
		_w402_
	);
	LUT4 #(
		.INIT('hf351)
	) name195 (
		\446(393)_pad ,
		\448(284)_pad ,
		_w397_,
		_w402_,
		_w403_
	);
	LUT2 #(
		.INIT('h4)
	) name196 (
		\446(393)_pad ,
		_w402_,
		_w404_
	);
	LUT4 #(
		.INIT('h51f3)
	) name197 (
		\12(3)_pad ,
		\18(5)_pad ,
		\214(137)_pad ,
		\9(2)_pad ,
		_w405_
	);
	LUT4 #(
		.INIT('h8acf)
	) name198 (
		\444(282)_pad ,
		\446(393)_pad ,
		_w402_,
		_w405_,
		_w406_
	);
	LUT3 #(
		.INIT('hb0)
	) name199 (
		_w401_,
		_w403_,
		_w406_,
		_w407_
	);
	LUT4 #(
		.INIT('h8caf)
	) name200 (
		\484(256)_pad ,
		\486(258)_pad ,
		_w357_,
		_w359_,
		_w408_
	);
	LUT4 #(
		.INIT('hf351)
	) name201 (
		\482(253)_pad ,
		\484(256)_pad ,
		_w357_,
		_w382_,
		_w409_
	);
	LUT4 #(
		.INIT('h8acf)
	) name202 (
		\480(250)_pad ,
		\482(253)_pad ,
		_w382_,
		_w386_,
		_w410_
	);
	LUT4 #(
		.INIT('h1055)
	) name203 (
		_w387_,
		_w408_,
		_w409_,
		_w410_,
		_w411_
	);
	LUT4 #(
		.INIT('h00b0)
	) name204 (
		_w394_,
		_w396_,
		_w407_,
		_w411_,
		_w412_
	);
	LUT2 #(
		.INIT('h4)
	) name205 (
		_w390_,
		_w412_,
		_w413_
	);
	LUT3 #(
		.INIT('h1d)
	) name206 (
		\100(51)_pad ,
		\18(5)_pad ,
		\231(154)_pad ,
		_w414_
	);
	LUT4 #(
		.INIT('h1d00)
	) name207 (
		\100(51)_pad ,
		\18(5)_pad ,
		\231(154)_pad ,
		\544(230)_pad ,
		_w415_
	);
	LUT3 #(
		.INIT('h1d)
	) name208 (
		\127(64)_pad ,
		\18(5)_pad ,
		\233(156)_pad ,
		_w416_
	);
	LUT3 #(
		.INIT('h1d)
	) name209 (
		\130(65)_pad ,
		\18(5)_pad ,
		\234(157)_pad ,
		_w417_
	);
	LUT4 #(
		.INIT('h00e2)
	) name210 (
		\130(65)_pad ,
		\18(5)_pad ,
		\234(157)_pad ,
		\550(236)_pad ,
		_w418_
	);
	LUT3 #(
		.INIT('h1d)
	) name211 (
		\124(63)_pad ,
		\18(5)_pad ,
		\232(155)_pad ,
		_w419_
	);
	LUT4 #(
		.INIT('h1d00)
	) name212 (
		\124(63)_pad ,
		\18(5)_pad ,
		\232(155)_pad ,
		\546(232)_pad ,
		_w420_
	);
	LUT4 #(
		.INIT('h0071)
	) name213 (
		\548(234)_pad ,
		_w416_,
		_w418_,
		_w420_,
		_w421_
	);
	LUT4 #(
		.INIT('h00e2)
	) name214 (
		\124(63)_pad ,
		\18(5)_pad ,
		\232(155)_pad ,
		\546(232)_pad ,
		_w422_
	);
	LUT4 #(
		.INIT('h00e2)
	) name215 (
		\100(51)_pad ,
		\18(5)_pad ,
		\231(154)_pad ,
		\544(230)_pad ,
		_w423_
	);
	LUT2 #(
		.INIT('h1)
	) name216 (
		_w422_,
		_w423_,
		_w424_
	);
	LUT3 #(
		.INIT('h45)
	) name217 (
		_w415_,
		_w421_,
		_w424_,
		_w425_
	);
	LUT3 #(
		.INIT('h27)
	) name218 (
		\18(5)_pad ,
		\220(143)_pad ,
		\50(15)_pad ,
		_w426_
	);
	LUT4 #(
		.INIT('h00d8)
	) name219 (
		\18(5)_pad ,
		\220(143)_pad ,
		\50(15)_pad ,
		\526(212)_pad ,
		_w427_
	);
	LUT4 #(
		.INIT('h2700)
	) name220 (
		\18(5)_pad ,
		\220(143)_pad ,
		\50(15)_pad ,
		\526(212)_pad ,
		_w428_
	);
	LUT4 #(
		.INIT('hd827)
	) name221 (
		\18(5)_pad ,
		\220(143)_pad ,
		\50(15)_pad ,
		\526(212)_pad ,
		_w429_
	);
	LUT3 #(
		.INIT('h27)
	) name222 (
		\18(5)_pad ,
		\221(144)_pad ,
		\32(9)_pad ,
		_w430_
	);
	LUT4 #(
		.INIT('hd827)
	) name223 (
		\18(5)_pad ,
		\221(144)_pad ,
		\32(9)_pad ,
		\528(214)_pad ,
		_w431_
	);
	LUT3 #(
		.INIT('h27)
	) name224 (
		\18(5)_pad ,
		\222(145)_pad ,
		\35(10)_pad ,
		_w432_
	);
	LUT4 #(
		.INIT('h00d8)
	) name225 (
		\18(5)_pad ,
		\222(145)_pad ,
		\35(10)_pad ,
		\530(216)_pad ,
		_w433_
	);
	LUT4 #(
		.INIT('h2700)
	) name226 (
		\18(5)_pad ,
		\222(145)_pad ,
		\35(10)_pad ,
		\530(216)_pad ,
		_w434_
	);
	LUT4 #(
		.INIT('hd827)
	) name227 (
		\18(5)_pad ,
		\222(145)_pad ,
		\35(10)_pad ,
		\530(216)_pad ,
		_w435_
	);
	LUT2 #(
		.INIT('h8)
	) name228 (
		_w431_,
		_w435_,
		_w436_
	);
	LUT3 #(
		.INIT('h80)
	) name229 (
		_w429_,
		_w431_,
		_w435_,
		_w437_
	);
	LUT3 #(
		.INIT('h1d)
	) name230 (
		\118(61)_pad ,
		\18(5)_pad ,
		\217(140)_pad ,
		_w438_
	);
	LUT4 #(
		.INIT('h00e2)
	) name231 (
		\118(61)_pad ,
		\18(5)_pad ,
		\217(140)_pad ,
		\522(226)_pad ,
		_w439_
	);
	LUT4 #(
		.INIT('h1d00)
	) name232 (
		\118(61)_pad ,
		\18(5)_pad ,
		\217(140)_pad ,
		\522(226)_pad ,
		_w440_
	);
	LUT4 #(
		.INIT('he21d)
	) name233 (
		\118(61)_pad ,
		\18(5)_pad ,
		\217(140)_pad ,
		\522(226)_pad ,
		_w441_
	);
	LUT3 #(
		.INIT('h27)
	) name234 (
		\18(5)_pad ,
		\226(149)_pad ,
		\97(50)_pad ,
		_w442_
	);
	LUT4 #(
		.INIT('h2070)
	) name235 (
		\18(5)_pad ,
		\226(149)_pad ,
		\538(224)_pad ,
		\97(50)_pad ,
		_w443_
	);
	LUT4 #(
		.INIT('h0d08)
	) name236 (
		\18(5)_pad ,
		\226(149)_pad ,
		\538(224)_pad ,
		\97(50)_pad ,
		_w444_
	);
	LUT4 #(
		.INIT('hd287)
	) name237 (
		\18(5)_pad ,
		\226(149)_pad ,
		\538(224)_pad ,
		\97(50)_pad ,
		_w445_
	);
	LUT3 #(
		.INIT('h27)
	) name238 (
		\18(5)_pad ,
		\225(148)_pad ,
		\94(49)_pad ,
		_w446_
	);
	LUT4 #(
		.INIT('h0d08)
	) name239 (
		\18(5)_pad ,
		\225(148)_pad ,
		\536(222)_pad ,
		\94(49)_pad ,
		_w447_
	);
	LUT4 #(
		.INIT('h2070)
	) name240 (
		\18(5)_pad ,
		\225(148)_pad ,
		\536(222)_pad ,
		\94(49)_pad ,
		_w448_
	);
	LUT4 #(
		.INIT('hd287)
	) name241 (
		\18(5)_pad ,
		\225(148)_pad ,
		\536(222)_pad ,
		\94(49)_pad ,
		_w449_
	);
	LUT3 #(
		.INIT('h80)
	) name242 (
		_w441_,
		_w445_,
		_w449_,
		_w450_
	);
	LUT3 #(
		.INIT('h1d)
	) name243 (
		\121(62)_pad ,
		\18(5)_pad ,
		\224(147)_pad ,
		_w451_
	);
	LUT4 #(
		.INIT('h1d00)
	) name244 (
		\121(62)_pad ,
		\18(5)_pad ,
		\224(147)_pad ,
		\534(220)_pad ,
		_w452_
	);
	LUT4 #(
		.INIT('h00e2)
	) name245 (
		\121(62)_pad ,
		\18(5)_pad ,
		\224(147)_pad ,
		\534(220)_pad ,
		_w453_
	);
	LUT4 #(
		.INIT('he21d)
	) name246 (
		\121(62)_pad ,
		\18(5)_pad ,
		\224(147)_pad ,
		\534(220)_pad ,
		_w454_
	);
	LUT3 #(
		.INIT('h27)
	) name247 (
		\18(5)_pad ,
		\223(146)_pad ,
		\47(14)_pad ,
		_w455_
	);
	LUT4 #(
		.INIT('h00d8)
	) name248 (
		\18(5)_pad ,
		\223(146)_pad ,
		\47(14)_pad ,
		\532(218)_pad ,
		_w456_
	);
	LUT4 #(
		.INIT('h2700)
	) name249 (
		\18(5)_pad ,
		\223(146)_pad ,
		\47(14)_pad ,
		\532(218)_pad ,
		_w457_
	);
	LUT4 #(
		.INIT('hd827)
	) name250 (
		\18(5)_pad ,
		\223(146)_pad ,
		\47(14)_pad ,
		\532(218)_pad ,
		_w458_
	);
	LUT2 #(
		.INIT('h8)
	) name251 (
		_w454_,
		_w458_,
		_w459_
	);
	LUT3 #(
		.INIT('h27)
	) name252 (
		\18(5)_pad ,
		\219(142)_pad ,
		\66(29)_pad ,
		_w460_
	);
	LUT4 #(
		.INIT('h2070)
	) name253 (
		\18(5)_pad ,
		\219(142)_pad ,
		\524(210)_pad ,
		\66(29)_pad ,
		_w461_
	);
	LUT4 #(
		.INIT('h0d08)
	) name254 (
		\18(5)_pad ,
		\219(142)_pad ,
		\524(210)_pad ,
		\66(29)_pad ,
		_w462_
	);
	LUT4 #(
		.INIT('hd287)
	) name255 (
		\18(5)_pad ,
		\219(142)_pad ,
		\524(210)_pad ,
		\66(29)_pad ,
		_w463_
	);
	LUT3 #(
		.INIT('h80)
	) name256 (
		_w454_,
		_w458_,
		_w463_,
		_w464_
	);
	LUT3 #(
		.INIT('h80)
	) name257 (
		_w437_,
		_w450_,
		_w464_,
		_w465_
	);
	LUT2 #(
		.INIT('h8)
	) name258 (
		_w425_,
		_w465_,
		_w466_
	);
	LUT3 #(
		.INIT('h1b)
	) name259 (
		\18(5)_pad ,
		\23(6)_pad ,
		\236(159)_pad ,
		_w467_
	);
	LUT4 #(
		.INIT('h00e4)
	) name260 (
		\18(5)_pad ,
		\23(6)_pad ,
		\236(159)_pad ,
		\554(240)_pad ,
		_w468_
	);
	LUT4 #(
		.INIT('h1b00)
	) name261 (
		\18(5)_pad ,
		\23(6)_pad ,
		\236(159)_pad ,
		\554(240)_pad ,
		_w469_
	);
	LUT3 #(
		.INIT('h1d)
	) name262 (
		\103(52)_pad ,
		\18(5)_pad ,
		\235(158)_pad ,
		_w470_
	);
	LUT4 #(
		.INIT('h1d00)
	) name263 (
		\103(52)_pad ,
		\18(5)_pad ,
		\235(158)_pad ,
		\552(238)_pad ,
		_w471_
	);
	LUT3 #(
		.INIT('h01)
	) name264 (
		\554(240)_pad ,
		_w467_,
		_w471_,
		_w472_
	);
	LUT3 #(
		.INIT('h27)
	) name265 (
		\18(5)_pad ,
		\238(161)_pad ,
		\29(8)_pad ,
		_w473_
	);
	LUT3 #(
		.INIT('h04)
	) name266 (
		\18(5)_pad ,
		\41(12)_pad ,
		\542(246)_pad ,
		_w474_
	);
	LUT3 #(
		.INIT('h27)
	) name267 (
		\18(5)_pad ,
		\237(160)_pad ,
		\26(7)_pad ,
		_w475_
	);
	LUT4 #(
		.INIT('h00d8)
	) name268 (
		\18(5)_pad ,
		\237(160)_pad ,
		\26(7)_pad ,
		\556(242)_pad ,
		_w476_
	);
	LUT4 #(
		.INIT('h008e)
	) name269 (
		\558(244)_pad ,
		_w473_,
		_w474_,
		_w476_,
		_w477_
	);
	LUT4 #(
		.INIT('h2700)
	) name270 (
		\18(5)_pad ,
		\237(160)_pad ,
		\26(7)_pad ,
		\556(242)_pad ,
		_w478_
	);
	LUT3 #(
		.INIT('h01)
	) name271 (
		_w469_,
		_w471_,
		_w478_,
		_w479_
	);
	LUT3 #(
		.INIT('h45)
	) name272 (
		_w472_,
		_w477_,
		_w479_,
		_w480_
	);
	LUT4 #(
		.INIT('h00e2)
	) name273 (
		\103(52)_pad ,
		\18(5)_pad ,
		\235(158)_pad ,
		\552(238)_pad ,
		_w481_
	);
	LUT4 #(
		.INIT('hd827)
	) name274 (
		\18(5)_pad ,
		\237(160)_pad ,
		\26(7)_pad ,
		\556(242)_pad ,
		_w482_
	);
	LUT3 #(
		.INIT('h10)
	) name275 (
		\18(5)_pad ,
		\41(12)_pad ,
		\542(246)_pad ,
		_w483_
	);
	LUT3 #(
		.INIT('heb)
	) name276 (
		\18(5)_pad ,
		\41(12)_pad ,
		\542(246)_pad ,
		_w484_
	);
	LUT4 #(
		.INIT('hd827)
	) name277 (
		\18(5)_pad ,
		\238(161)_pad ,
		\29(8)_pad ,
		\558(244)_pad ,
		_w485_
	);
	LUT2 #(
		.INIT('h8)
	) name278 (
		_w484_,
		_w485_,
		_w486_
	);
	LUT4 #(
		.INIT('h0028)
	) name279 (
		\4526(205)_pad ,
		\554(240)_pad ,
		_w467_,
		_w471_,
		_w487_
	);
	LUT3 #(
		.INIT('h80)
	) name280 (
		_w482_,
		_w486_,
		_w487_,
		_w488_
	);
	LUT4 #(
		.INIT('h1555)
	) name281 (
		_w481_,
		_w482_,
		_w486_,
		_w487_,
		_w489_
	);
	LUT4 #(
		.INIT('he21d)
	) name282 (
		\127(64)_pad ,
		\18(5)_pad ,
		\233(156)_pad ,
		\548(234)_pad ,
		_w490_
	);
	LUT4 #(
		.INIT('h1d00)
	) name283 (
		\130(65)_pad ,
		\18(5)_pad ,
		\234(157)_pad ,
		\550(236)_pad ,
		_w491_
	);
	LUT4 #(
		.INIT('he21d)
	) name284 (
		\130(65)_pad ,
		\18(5)_pad ,
		\234(157)_pad ,
		\550(236)_pad ,
		_w492_
	);
	LUT2 #(
		.INIT('h8)
	) name285 (
		_w490_,
		_w492_,
		_w493_
	);
	LUT4 #(
		.INIT('he21d)
	) name286 (
		\124(63)_pad ,
		\18(5)_pad ,
		\232(155)_pad ,
		\546(232)_pad ,
		_w494_
	);
	LUT4 #(
		.INIT('he21d)
	) name287 (
		\100(51)_pad ,
		\18(5)_pad ,
		\231(154)_pad ,
		\544(230)_pad ,
		_w495_
	);
	LUT4 #(
		.INIT('h8000)
	) name288 (
		_w490_,
		_w492_,
		_w494_,
		_w495_,
		_w496_
	);
	LUT4 #(
		.INIT('h8000)
	) name289 (
		_w437_,
		_w450_,
		_w464_,
		_w496_,
		_w497_
	);
	LUT3 #(
		.INIT('h70)
	) name290 (
		_w480_,
		_w489_,
		_w497_,
		_w498_
	);
	LUT2 #(
		.INIT('h1)
	) name291 (
		_w427_,
		_w462_,
		_w499_
	);
	LUT4 #(
		.INIT('h0080)
	) name292 (
		_w429_,
		_w431_,
		_w435_,
		_w457_,
		_w500_
	);
	LUT4 #(
		.INIT('h1301)
	) name293 (
		\528(214)_pad ,
		_w428_,
		_w430_,
		_w433_,
		_w501_
	);
	LUT2 #(
		.INIT('h1)
	) name294 (
		_w500_,
		_w501_,
		_w502_
	);
	LUT4 #(
		.INIT('h00b2)
	) name295 (
		\538(224)_pad ,
		_w439_,
		_w442_,
		_w447_,
		_w503_
	);
	LUT2 #(
		.INIT('h1)
	) name296 (
		_w448_,
		_w452_,
		_w504_
	);
	LUT2 #(
		.INIT('h4)
	) name297 (
		_w503_,
		_w504_,
		_w505_
	);
	LUT2 #(
		.INIT('h1)
	) name298 (
		_w453_,
		_w456_,
		_w506_
	);
	LUT4 #(
		.INIT('h4500)
	) name299 (
		_w501_,
		_w503_,
		_w504_,
		_w506_,
		_w507_
	);
	LUT4 #(
		.INIT('h1115)
	) name300 (
		_w461_,
		_w499_,
		_w502_,
		_w507_,
		_w508_
	);
	LUT4 #(
		.INIT('h0002)
	) name301 (
		_w412_,
		_w466_,
		_w498_,
		_w508_,
		_w509_
	);
	LUT2 #(
		.INIT('h9)
	) name302 (
		\446(393)_pad ,
		_w402_,
		_w510_
	);
	LUT4 #(
		.INIT('h8241)
	) name303 (
		\446(393)_pad ,
		\448(284)_pad ,
		_w397_,
		_w402_,
		_w511_
	);
	LUT2 #(
		.INIT('h9)
	) name304 (
		\436(286)_pad ,
		_w399_,
		_w512_
	);
	LUT2 #(
		.INIT('h8)
	) name305 (
		_w511_,
		_w512_,
		_w513_
	);
	LUT2 #(
		.INIT('h2)
	) name306 (
		_w407_,
		_w513_,
		_w514_
	);
	LUT4 #(
		.INIT('h51f3)
	) name307 (
		\12(3)_pad ,
		\18(5)_pad ,
		\213(136)_pad ,
		\9(2)_pad ,
		_w515_
	);
	LUT2 #(
		.INIT('h4)
	) name308 (
		\442(280)_pad ,
		_w515_,
		_w516_
	);
	LUT2 #(
		.INIT('h9)
	) name309 (
		\442(280)_pad ,
		_w515_,
		_w517_
	);
	LUT2 #(
		.INIT('h2)
	) name310 (
		\444(282)_pad ,
		_w405_,
		_w518_
	);
	LUT4 #(
		.INIT('ha251)
	) name311 (
		\442(280)_pad ,
		\444(282)_pad ,
		_w405_,
		_w515_,
		_w519_
	);
	LUT3 #(
		.INIT('hd0)
	) name312 (
		_w407_,
		_w513_,
		_w519_,
		_w520_
	);
	LUT3 #(
		.INIT('h10)
	) name313 (
		_w413_,
		_w509_,
		_w520_,
		_w521_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name314 (
		\38(11)_pad ,
		\438(274)_pad ,
		\440(277)_pad ,
		\4528(206)_pad ,
		_w522_
	);
	LUT3 #(
		.INIT('h0b)
	) name315 (
		\442(280)_pad ,
		_w515_,
		_w522_,
		_w523_
	);
	LUT4 #(
		.INIT('hef00)
	) name316 (
		_w413_,
		_w509_,
		_w520_,
		_w523_,
		_w524_
	);
	LUT4 #(
		.INIT('h5400)
	) name317 (
		\38(11)_pad ,
		\438(274)_pad ,
		\440(277)_pad ,
		\4528(206)_pad ,
		_w525_
	);
	LUT2 #(
		.INIT('h1)
	) name318 (
		_w524_,
		_w525_,
		_w526_
	);
	LUT2 #(
		.INIT('h8)
	) name319 (
		\163(86)_pad ,
		\453(596)_pad ,
		_w527_
	);
	LUT3 #(
		.INIT('hf7)
	) name320 (
		\133(66)_pad ,
		\134(67)_pad ,
		\5(1)_pad ,
		_w528_
	);
	LUT2 #(
		.INIT('hd)
	) name321 (
		\1197(165)_pad ,
		\5(1)_pad ,
		_w529_
	);
	LUT3 #(
		.INIT('h01)
	) name322 (
		_w466_,
		_w498_,
		_w508_,
		_w530_
	);
	LUT4 #(
		.INIT('h5556)
	) name323 (
		_w365_,
		_w466_,
		_w498_,
		_w508_,
		_w531_
	);
	LUT2 #(
		.INIT('h8)
	) name324 (
		_w361_,
		_w385_,
		_w532_
	);
	LUT2 #(
		.INIT('h8)
	) name325 (
		_w374_,
		_w381_,
		_w533_
	);
	LUT2 #(
		.INIT('h2)
	) name326 (
		_w394_,
		_w533_,
		_w534_
	);
	LUT4 #(
		.INIT('h0002)
	) name327 (
		_w394_,
		_w466_,
		_w498_,
		_w508_,
		_w535_
	);
	LUT3 #(
		.INIT('h45)
	) name328 (
		_w383_,
		_w408_,
		_w409_,
		_w536_
	);
	LUT4 #(
		.INIT('h1011)
	) name329 (
		_w383_,
		_w388_,
		_w408_,
		_w409_,
		_w537_
	);
	LUT4 #(
		.INIT('hfd00)
	) name330 (
		_w532_,
		_w534_,
		_w535_,
		_w537_,
		_w538_
	);
	LUT2 #(
		.INIT('h8)
	) name331 (
		_w361_,
		_w389_,
		_w539_
	);
	LUT4 #(
		.INIT('h8c88)
	) name332 (
		_w383_,
		_w388_,
		_w408_,
		_w409_,
		_w540_
	);
	LUT4 #(
		.INIT('h00ef)
	) name333 (
		_w534_,
		_w535_,
		_w539_,
		_w540_,
		_w541_
	);
	LUT2 #(
		.INIT('h4)
	) name334 (
		_w538_,
		_w541_,
		_w542_
	);
	LUT4 #(
		.INIT('h7150)
	) name335 (
		\484(256)_pad ,
		\486(258)_pad ,
		_w357_,
		_w359_,
		_w543_
	);
	LUT4 #(
		.INIT('hf571)
	) name336 (
		\484(256)_pad ,
		\486(258)_pad ,
		_w357_,
		_w359_,
		_w544_
	);
	LUT2 #(
		.INIT('h4)
	) name337 (
		_w385_,
		_w544_,
		_w545_
	);
	LUT4 #(
		.INIT('hf100)
	) name338 (
		_w534_,
		_w535_,
		_w543_,
		_w545_,
		_w546_
	);
	LUT2 #(
		.INIT('h2)
	) name339 (
		_w385_,
		_w544_,
		_w547_
	);
	LUT2 #(
		.INIT('h2)
	) name340 (
		_w385_,
		_w543_,
		_w548_
	);
	LUT4 #(
		.INIT('h010f)
	) name341 (
		_w534_,
		_w535_,
		_w547_,
		_w548_,
		_w549_
	);
	LUT2 #(
		.INIT('hb)
	) name342 (
		_w546_,
		_w549_,
		_w550_
	);
	LUT4 #(
		.INIT('ha569)
	) name343 (
		\484(256)_pad ,
		\486(258)_pad ,
		_w357_,
		_w359_,
		_w551_
	);
	LUT4 #(
		.INIT('h0057)
	) name344 (
		_w360_,
		_w534_,
		_w535_,
		_w551_,
		_w552_
	);
	LUT3 #(
		.INIT('ha8)
	) name345 (
		_w361_,
		_w534_,
		_w535_,
		_w553_
	);
	LUT2 #(
		.INIT('he)
	) name346 (
		_w552_,
		_w553_,
		_w554_
	);
	LUT3 #(
		.INIT('ha9)
	) name347 (
		_w360_,
		_w534_,
		_w535_,
		_w555_
	);
	LUT4 #(
		.INIT('h0001)
	) name348 (
		_w363_,
		_w466_,
		_w498_,
		_w508_,
		_w556_
	);
	LUT3 #(
		.INIT('h04)
	) name349 (
		_w364_,
		_w369_,
		_w372_,
		_w557_
	);
	LUT2 #(
		.INIT('h8)
	) name350 (
		_w369_,
		_w371_,
		_w558_
	);
	LUT4 #(
		.INIT('h008e)
	) name351 (
		\492(265)_pad ,
		_w366_,
		_w371_,
		_w376_,
		_w559_
	);
	LUT3 #(
		.INIT('h21)
	) name352 (
		\488(260)_pad ,
		_w377_,
		_w379_,
		_w560_
	);
	LUT4 #(
		.INIT('h4f00)
	) name353 (
		_w556_,
		_w557_,
		_w559_,
		_w560_,
		_w561_
	);
	LUT4 #(
		.INIT('h1055)
	) name354 (
		_w377_,
		_w556_,
		_w557_,
		_w559_,
		_w562_
	);
	LUT3 #(
		.INIT('h32)
	) name355 (
		_w380_,
		_w561_,
		_w562_,
		_w563_
	);
	LUT3 #(
		.INIT('h8e)
	) name356 (
		\492(265)_pad ,
		_w366_,
		_w371_,
		_w564_
	);
	LUT4 #(
		.INIT('h1055)
	) name357 (
		_w378_,
		_w556_,
		_w557_,
		_w564_,
		_w565_
	);
	LUT4 #(
		.INIT('h8e00)
	) name358 (
		\492(265)_pad ,
		_w366_,
		_w371_,
		_w378_,
		_w566_
	);
	LUT3 #(
		.INIT('hb0)
	) name359 (
		_w556_,
		_w557_,
		_w566_,
		_w567_
	);
	LUT2 #(
		.INIT('he)
	) name360 (
		_w565_,
		_w567_,
		_w568_
	);
	LUT3 #(
		.INIT('h0b)
	) name361 (
		_w556_,
		_w557_,
		_w558_,
		_w569_
	);
	LUT2 #(
		.INIT('h1)
	) name362 (
		_w364_,
		_w372_,
		_w570_
	);
	LUT2 #(
		.INIT('h1)
	) name363 (
		_w369_,
		_w371_,
		_w571_
	);
	LUT3 #(
		.INIT('hb0)
	) name364 (
		_w556_,
		_w570_,
		_w571_,
		_w572_
	);
	LUT2 #(
		.INIT('h2)
	) name365 (
		_w569_,
		_w572_,
		_w573_
	);
	LUT3 #(
		.INIT('hc9)
	) name366 (
		_w364_,
		_w373_,
		_w556_,
		_w574_
	);
	LUT2 #(
		.INIT('h6)
	) name367 (
		_w369_,
		_w373_,
		_w575_
	);
	LUT3 #(
		.INIT('h81)
	) name368 (
		\494(267)_pad ,
		_w363_,
		_w370_,
		_w576_
	);
	LUT2 #(
		.INIT('h1)
	) name369 (
		_w368_,
		_w377_,
		_w577_
	);
	LUT2 #(
		.INIT('h4)
	) name370 (
		_w391_,
		_w577_,
		_w578_
	);
	LUT2 #(
		.INIT('h1)
	) name371 (
		_w368_,
		_w391_,
		_w579_
	);
	LUT3 #(
		.INIT('h32)
	) name372 (
		_w368_,
		_w376_,
		_w391_,
		_w580_
	);
	LUT4 #(
		.INIT('h3c39)
	) name373 (
		_w376_,
		_w576_,
		_w578_,
		_w579_,
		_w581_
	);
	LUT2 #(
		.INIT('h6)
	) name374 (
		_w365_,
		_w581_,
		_w582_
	);
	LUT4 #(
		.INIT('h0080)
	) name375 (
		_w365_,
		_w369_,
		_w373_,
		_w377_,
		_w583_
	);
	LUT3 #(
		.INIT('h0b)
	) name376 (
		_w391_,
		_w577_,
		_w583_,
		_w584_
	);
	LUT3 #(
		.INIT('h24)
	) name377 (
		\494(267)_pad ,
		_w364_,
		_w370_,
		_w585_
	);
	LUT4 #(
		.INIT('hb04f)
	) name378 (
		_w374_,
		_w580_,
		_w584_,
		_w585_,
		_w586_
	);
	LUT3 #(
		.INIT('h4e)
	) name379 (
		_w365_,
		_w581_,
		_w586_,
		_w587_
	);
	LUT4 #(
		.INIT('h93c6)
	) name380 (
		_w530_,
		_w575_,
		_w582_,
		_w587_,
		_w588_
	);
	LUT3 #(
		.INIT('h69)
	) name381 (
		\488(260)_pad ,
		_w378_,
		_w379_,
		_w589_
	);
	LUT4 #(
		.INIT('h6996)
	) name382 (
		\480(250)_pad ,
		\482(253)_pad ,
		_w382_,
		_w386_,
		_w590_
	);
	LUT2 #(
		.INIT('h6)
	) name383 (
		_w589_,
		_w590_,
		_w591_
	);
	LUT3 #(
		.INIT('h70)
	) name384 (
		_w361_,
		_w385_,
		_w544_,
		_w592_
	);
	LUT4 #(
		.INIT('h96a5)
	) name385 (
		\484(256)_pad ,
		\486(258)_pad ,
		_w357_,
		_w359_,
		_w593_
	);
	LUT2 #(
		.INIT('h2)
	) name386 (
		_w383_,
		_w544_,
		_w594_
	);
	LUT4 #(
		.INIT('h0f78)
	) name387 (
		_w536_,
		_w592_,
		_w593_,
		_w594_,
		_w595_
	);
	LUT4 #(
		.INIT('hccd8)
	) name388 (
		_w358_,
		_w383_,
		_w384_,
		_w408_,
		_w596_
	);
	LUT2 #(
		.INIT('h9)
	) name389 (
		_w551_,
		_w596_,
		_w597_
	);
	LUT4 #(
		.INIT('hef01)
	) name390 (
		_w534_,
		_w535_,
		_w595_,
		_w597_,
		_w598_
	);
	LUT3 #(
		.INIT('h69)
	) name391 (
		_w588_,
		_w591_,
		_w598_,
		_w599_
	);
	LUT3 #(
		.INIT('h0b)
	) name392 (
		_w394_,
		_w396_,
		_w411_,
		_w600_
	);
	LUT4 #(
		.INIT('h0045)
	) name393 (
		_w390_,
		_w394_,
		_w396_,
		_w411_,
		_w601_
	);
	LUT4 #(
		.INIT('h0100)
	) name394 (
		_w466_,
		_w498_,
		_w508_,
		_w600_,
		_w602_
	);
	LUT2 #(
		.INIT('h1)
	) name395 (
		_w601_,
		_w602_,
		_w603_
	);
	LUT3 #(
		.INIT('ha9)
	) name396 (
		_w512_,
		_w601_,
		_w602_,
		_w604_
	);
	LUT3 #(
		.INIT('h0d)
	) name397 (
		_w407_,
		_w513_,
		_w518_,
		_w605_
	);
	LUT4 #(
		.INIT('h0e0f)
	) name398 (
		_w413_,
		_w509_,
		_w517_,
		_w605_,
		_w606_
	);
	LUT2 #(
		.INIT('h1)
	) name399 (
		_w521_,
		_w606_,
		_w607_
	);
	LUT2 #(
		.INIT('h9)
	) name400 (
		\444(282)_pad ,
		_w405_,
		_w608_
	);
	LUT3 #(
		.INIT('h0b)
	) name401 (
		_w401_,
		_w403_,
		_w404_,
		_w609_
	);
	LUT3 #(
		.INIT('h10)
	) name402 (
		_w513_,
		_w608_,
		_w609_,
		_w610_
	);
	LUT4 #(
		.INIT('h000b)
	) name403 (
		_w401_,
		_w403_,
		_w404_,
		_w608_,
		_w611_
	);
	LUT4 #(
		.INIT('h010f)
	) name404 (
		_w601_,
		_w602_,
		_w610_,
		_w611_,
		_w612_
	);
	LUT3 #(
		.INIT('h8c)
	) name405 (
		_w513_,
		_w608_,
		_w609_,
		_w613_
	);
	LUT4 #(
		.INIT('h1f00)
	) name406 (
		_w601_,
		_w602_,
		_w609_,
		_w613_,
		_w614_
	);
	LUT2 #(
		.INIT('h2)
	) name407 (
		_w612_,
		_w614_,
		_w615_
	);
	LUT4 #(
		.INIT('hf351)
	) name408 (
		\436(286)_pad ,
		\448(284)_pad ,
		_w397_,
		_w399_,
		_w616_
	);
	LUT4 #(
		.INIT('hab00)
	) name409 (
		_w400_,
		_w601_,
		_w602_,
		_w616_,
		_w617_
	);
	LUT2 #(
		.INIT('h8)
	) name410 (
		_w510_,
		_w616_,
		_w618_
	);
	LUT4 #(
		.INIT('hab00)
	) name411 (
		_w400_,
		_w601_,
		_w602_,
		_w618_,
		_w619_
	);
	LUT4 #(
		.INIT('h0076)
	) name412 (
		_w398_,
		_w510_,
		_w617_,
		_w619_,
		_w620_
	);
	LUT4 #(
		.INIT('h3c14)
	) name413 (
		\436(286)_pad ,
		\448(284)_pad ,
		_w397_,
		_w399_,
		_w621_
	);
	LUT4 #(
		.INIT('hab00)
	) name414 (
		_w400_,
		_w601_,
		_w602_,
		_w621_,
		_w622_
	);
	LUT4 #(
		.INIT('h0082)
	) name415 (
		\436(286)_pad ,
		\448(284)_pad ,
		_w397_,
		_w399_,
		_w623_
	);
	LUT4 #(
		.INIT('h82c3)
	) name416 (
		\436(286)_pad ,
		\448(284)_pad ,
		_w397_,
		_w399_,
		_w624_
	);
	LUT4 #(
		.INIT('h010f)
	) name417 (
		_w601_,
		_w602_,
		_w623_,
		_w624_,
		_w625_
	);
	LUT2 #(
		.INIT('hb)
	) name418 (
		_w622_,
		_w625_,
		_w626_
	);
	LUT4 #(
		.INIT('h6996)
	) name419 (
		\446(393)_pad ,
		\448(284)_pad ,
		_w397_,
		_w402_,
		_w627_
	);
	LUT2 #(
		.INIT('h6)
	) name420 (
		_w517_,
		_w627_,
		_w628_
	);
	LUT4 #(
		.INIT('h2430)
	) name421 (
		\436(286)_pad ,
		\448(284)_pad ,
		_w397_,
		_w399_,
		_w629_
	);
	LUT4 #(
		.INIT('hb000)
	) name422 (
		_w401_,
		_w403_,
		_w406_,
		_w629_,
		_w630_
	);
	LUT2 #(
		.INIT('h4)
	) name423 (
		_w518_,
		_w629_,
		_w631_
	);
	LUT3 #(
		.INIT('h23)
	) name424 (
		_w609_,
		_w630_,
		_w631_,
		_w632_
	);
	LUT4 #(
		.INIT('h00f4)
	) name425 (
		_w401_,
		_w403_,
		_w404_,
		_w518_,
		_w633_
	);
	LUT4 #(
		.INIT('h004f)
	) name426 (
		_w401_,
		_w403_,
		_w406_,
		_w629_,
		_w634_
	);
	LUT2 #(
		.INIT('h4)
	) name427 (
		_w633_,
		_w634_,
		_w635_
	);
	LUT4 #(
		.INIT('h8421)
	) name428 (
		\436(286)_pad ,
		\444(282)_pad ,
		_w399_,
		_w405_,
		_w636_
	);
	LUT4 #(
		.INIT('h6696)
	) name429 (
		_w512_,
		_w608_,
		_w632_,
		_w635_,
		_w637_
	);
	LUT3 #(
		.INIT('h0e)
	) name430 (
		_w601_,
		_w602_,
		_w637_,
		_w638_
	);
	LUT3 #(
		.INIT('h51)
	) name431 (
		_w512_,
		_w632_,
		_w635_,
		_w639_
	);
	LUT3 #(
		.INIT('h23)
	) name432 (
		_w513_,
		_w518_,
		_w609_,
		_w640_
	);
	LUT4 #(
		.INIT('h0c24)
	) name433 (
		\436(286)_pad ,
		\448(284)_pad ,
		_w397_,
		_w399_,
		_w641_
	);
	LUT4 #(
		.INIT('h02a8)
	) name434 (
		_w512_,
		_w514_,
		_w640_,
		_w641_,
		_w642_
	);
	LUT3 #(
		.INIT('ha9)
	) name435 (
		_w608_,
		_w639_,
		_w642_,
		_w643_
	);
	LUT4 #(
		.INIT('hc9c3)
	) name436 (
		_w603_,
		_w628_,
		_w638_,
		_w643_,
		_w644_
	);
	LUT3 #(
		.INIT('h80)
	) name437 (
		_w511_,
		_w517_,
		_w636_,
		_w645_
	);
	LUT4 #(
		.INIT('hf351)
	) name438 (
		\442(280)_pad ,
		\444(282)_pad ,
		_w405_,
		_w515_,
		_w646_
	);
	LUT4 #(
		.INIT('h4f00)
	) name439 (
		_w401_,
		_w403_,
		_w406_,
		_w646_,
		_w647_
	);
	LUT4 #(
		.INIT('hc955)
	) name440 (
		\38(11)_pad ,
		\438(274)_pad ,
		\440(277)_pad ,
		\4528(206)_pad ,
		_w648_
	);
	LUT3 #(
		.INIT('hb0)
	) name441 (
		\442(280)_pad ,
		_w515_,
		_w648_,
		_w649_
	);
	LUT2 #(
		.INIT('h4)
	) name442 (
		_w647_,
		_w649_,
		_w650_
	);
	LUT4 #(
		.INIT('hef00)
	) name443 (
		_w601_,
		_w602_,
		_w645_,
		_w650_,
		_w651_
	);
	LUT2 #(
		.INIT('h1)
	) name444 (
		_w516_,
		_w647_,
		_w652_
	);
	LUT4 #(
		.INIT('hef00)
	) name445 (
		_w601_,
		_w602_,
		_w645_,
		_w652_,
		_w653_
	);
	LUT4 #(
		.INIT('h6c00)
	) name446 (
		\38(11)_pad ,
		\438(274)_pad ,
		\440(277)_pad ,
		\4528(206)_pad ,
		_w654_
	);
	LUT3 #(
		.INIT('h54)
	) name447 (
		_w651_,
		_w653_,
		_w654_,
		_w655_
	);
	LUT2 #(
		.INIT('h6)
	) name448 (
		_w644_,
		_w655_,
		_w656_
	);
	LUT2 #(
		.INIT('h4)
	) name449 (
		_w415_,
		_w441_,
		_w657_
	);
	LUT3 #(
		.INIT('hb0)
	) name450 (
		_w421_,
		_w424_,
		_w657_,
		_w658_
	);
	LUT2 #(
		.INIT('h8)
	) name451 (
		_w441_,
		_w496_,
		_w659_
	);
	LUT4 #(
		.INIT('hf7f0)
	) name452 (
		_w480_,
		_w489_,
		_w658_,
		_w659_,
		_w660_
	);
	LUT2 #(
		.INIT('h2)
	) name453 (
		_w415_,
		_w441_,
		_w661_
	);
	LUT3 #(
		.INIT('h01)
	) name454 (
		_w422_,
		_w423_,
		_w441_,
		_w662_
	);
	LUT3 #(
		.INIT('h23)
	) name455 (
		_w421_,
		_w661_,
		_w662_,
		_w663_
	);
	LUT4 #(
		.INIT('h3130)
	) name456 (
		_w421_,
		_w496_,
		_w661_,
		_w662_,
		_w664_
	);
	LUT4 #(
		.INIT('h00f7)
	) name457 (
		_w480_,
		_w489_,
		_w663_,
		_w664_,
		_w665_
	);
	LUT2 #(
		.INIT('h4)
	) name458 (
		_w660_,
		_w665_,
		_w666_
	);
	LUT2 #(
		.INIT('h1)
	) name459 (
		_w427_,
		_w501_,
		_w667_
	);
	LUT3 #(
		.INIT('h01)
	) name460 (
		_w427_,
		_w437_,
		_w501_,
		_w668_
	);
	LUT3 #(
		.INIT('h4d)
	) name461 (
		\532(218)_pad ,
		_w453_,
		_w455_,
		_w669_
	);
	LUT3 #(
		.INIT('h01)
	) name462 (
		_w448_,
		_w452_,
		_w457_,
		_w670_
	);
	LUT3 #(
		.INIT('h23)
	) name463 (
		_w503_,
		_w669_,
		_w670_,
		_w671_
	);
	LUT3 #(
		.INIT('h13)
	) name464 (
		_w667_,
		_w668_,
		_w671_,
		_w672_
	);
	LUT4 #(
		.INIT('h00ba)
	) name465 (
		_w415_,
		_w421_,
		_w424_,
		_w496_,
		_w673_
	);
	LUT4 #(
		.INIT('h00bf)
	) name466 (
		_w425_,
		_w480_,
		_w489_,
		_w673_,
		_w674_
	);
	LUT2 #(
		.INIT('h8)
	) name467 (
		_w450_,
		_w459_,
		_w675_
	);
	LUT2 #(
		.INIT('h4)
	) name468 (
		_w668_,
		_w675_,
		_w676_
	);
	LUT4 #(
		.INIT('h5666)
	) name469 (
		_w463_,
		_w672_,
		_w674_,
		_w676_,
		_w677_
	);
	LUT3 #(
		.INIT('h71)
	) name470 (
		\528(214)_pad ,
		_w430_,
		_w433_,
		_w678_
	);
	LUT4 #(
		.INIT('h0023)
	) name471 (
		_w503_,
		_w669_,
		_w670_,
		_w678_,
		_w679_
	);
	LUT3 #(
		.INIT('h17)
	) name472 (
		\528(214)_pad ,
		_w430_,
		_w434_,
		_w680_
	);
	LUT4 #(
		.INIT('h0113)
	) name473 (
		\528(214)_pad ,
		_w429_,
		_w430_,
		_w434_,
		_w681_
	);
	LUT4 #(
		.INIT('h8f00)
	) name474 (
		_w674_,
		_w675_,
		_w679_,
		_w681_,
		_w682_
	);
	LUT4 #(
		.INIT('h8f00)
	) name475 (
		_w674_,
		_w675_,
		_w679_,
		_w680_,
		_w683_
	);
	LUT3 #(
		.INIT('hce)
	) name476 (
		_w429_,
		_w682_,
		_w683_,
		_w684_
	);
	LUT4 #(
		.INIT('h080a)
	) name477 (
		_w435_,
		_w503_,
		_w669_,
		_w670_,
		_w685_
	);
	LUT2 #(
		.INIT('h6)
	) name478 (
		_w431_,
		_w434_,
		_w686_
	);
	LUT4 #(
		.INIT('h008f)
	) name479 (
		_w674_,
		_w675_,
		_w685_,
		_w686_,
		_w687_
	);
	LUT4 #(
		.INIT('h080a)
	) name480 (
		_w436_,
		_w503_,
		_w669_,
		_w670_,
		_w688_
	);
	LUT3 #(
		.INIT('h70)
	) name481 (
		_w674_,
		_w675_,
		_w688_,
		_w689_
	);
	LUT2 #(
		.INIT('he)
	) name482 (
		_w687_,
		_w689_,
		_w690_
	);
	LUT4 #(
		.INIT('h5999)
	) name483 (
		_w435_,
		_w671_,
		_w674_,
		_w675_,
		_w691_
	);
	LUT2 #(
		.INIT('h1)
	) name484 (
		_w448_,
		_w503_,
		_w692_
	);
	LUT4 #(
		.INIT('h0517)
	) name485 (
		\534(220)_pad ,
		_w448_,
		_w451_,
		_w503_,
		_w693_
	);
	LUT4 #(
		.INIT('h0080)
	) name486 (
		_w441_,
		_w445_,
		_w449_,
		_w452_,
		_w694_
	);
	LUT4 #(
		.INIT('h565a)
	) name487 (
		_w458_,
		_w674_,
		_w693_,
		_w694_,
		_w695_
	);
	LUT4 #(
		.INIT('h336c)
	) name488 (
		_w450_,
		_w454_,
		_w674_,
		_w692_,
		_w696_
	);
	LUT2 #(
		.INIT('h1)
	) name489 (
		_w439_,
		_w444_,
		_w697_
	);
	LUT4 #(
		.INIT('h9c99)
	) name490 (
		_w443_,
		_w449_,
		_w660_,
		_w697_,
		_w698_
	);
	LUT3 #(
		.INIT('h36)
	) name491 (
		_w439_,
		_w445_,
		_w660_,
		_w699_
	);
	LUT2 #(
		.INIT('h6)
	) name492 (
		_w445_,
		_w449_,
		_w700_
	);
	LUT3 #(
		.INIT('h81)
	) name493 (
		\538(224)_pad ,
		_w439_,
		_w442_,
		_w701_
	);
	LUT4 #(
		.INIT('h32cd)
	) name494 (
		_w453_,
		_w505_,
		_w692_,
		_w701_,
		_w702_
	);
	LUT3 #(
		.INIT('h04)
	) name495 (
		_w660_,
		_w665_,
		_w702_,
		_w703_
	);
	LUT3 #(
		.INIT('h32)
	) name496 (
		_w448_,
		_w450_,
		_w503_,
		_w704_
	);
	LUT3 #(
		.INIT('hdb)
	) name497 (
		\538(224)_pad ,
		_w440_,
		_w442_,
		_w705_
	);
	LUT4 #(
		.INIT('he718)
	) name498 (
		\534(220)_pad ,
		_w451_,
		_w704_,
		_w705_,
		_w706_
	);
	LUT4 #(
		.INIT('h45cf)
	) name499 (
		_w660_,
		_w665_,
		_w702_,
		_w706_,
		_w707_
	);
	LUT4 #(
		.INIT('h41cb)
	) name500 (
		_w660_,
		_w665_,
		_w702_,
		_w706_,
		_w708_
	);
	LUT2 #(
		.INIT('h2)
	) name501 (
		_w700_,
		_w708_,
		_w709_
	);
	LUT4 #(
		.INIT('h9669)
	) name502 (
		_w429_,
		_w454_,
		_w458_,
		_w463_,
		_w710_
	);
	LUT4 #(
		.INIT('h00ef)
	) name503 (
		_w700_,
		_w703_,
		_w707_,
		_w710_,
		_w711_
	);
	LUT4 #(
		.INIT('h2032)
	) name504 (
		\528(214)_pad ,
		_w427_,
		_w430_,
		_w433_,
		_w712_
	);
	LUT3 #(
		.INIT('h36)
	) name505 (
		_w501_,
		_w686_,
		_w712_,
		_w713_
	);
	LUT2 #(
		.INIT('h8)
	) name506 (
		_w671_,
		_w713_,
		_w714_
	);
	LUT3 #(
		.INIT('h70)
	) name507 (
		_w674_,
		_w675_,
		_w714_,
		_w715_
	);
	LUT4 #(
		.INIT('h0100)
	) name508 (
		_w427_,
		_w437_,
		_w501_,
		_w680_,
		_w716_
	);
	LUT2 #(
		.INIT('h6)
	) name509 (
		_w431_,
		_w433_,
		_w717_
	);
	LUT4 #(
		.INIT('h175f)
	) name510 (
		\528(214)_pad ,
		\530(216)_pad ,
		_w430_,
		_w432_,
		_w718_
	);
	LUT3 #(
		.INIT('hc4)
	) name511 (
		_w427_,
		_w717_,
		_w718_,
		_w719_
	);
	LUT2 #(
		.INIT('h4)
	) name512 (
		_w716_,
		_w719_,
		_w720_
	);
	LUT3 #(
		.INIT('h02)
	) name513 (
		_w427_,
		_w717_,
		_w718_,
		_w721_
	);
	LUT4 #(
		.INIT('h0516)
	) name514 (
		\528(214)_pad ,
		\530(216)_pad ,
		_w430_,
		_w432_,
		_w722_
	);
	LUT4 #(
		.INIT('h0100)
	) name515 (
		_w427_,
		_w437_,
		_w501_,
		_w722_,
		_w723_
	);
	LUT3 #(
		.INIT('h01)
	) name516 (
		_w671_,
		_w721_,
		_w723_,
		_w724_
	);
	LUT3 #(
		.INIT('h02)
	) name517 (
		_w675_,
		_w721_,
		_w723_,
		_w725_
	);
	LUT4 #(
		.INIT('h3230)
	) name518 (
		_w674_,
		_w720_,
		_w724_,
		_w725_,
		_w726_
	);
	LUT2 #(
		.INIT('h1)
	) name519 (
		_w715_,
		_w726_,
		_w727_
	);
	LUT3 #(
		.INIT('h9f)
	) name520 (
		_w700_,
		_w708_,
		_w710_,
		_w728_
	);
	LUT4 #(
		.INIT('hb40f)
	) name521 (
		_w709_,
		_w711_,
		_w727_,
		_w728_,
		_w729_
	);
	LUT4 #(
		.INIT('he0b0)
	) name522 (
		\18(5)_pad ,
		\41(12)_pad ,
		\4526(205)_pad ,
		\542(246)_pad ,
		_w730_
	);
	LUT4 #(
		.INIT('hfefb)
	) name523 (
		\18(5)_pad ,
		\41(12)_pad ,
		\4526(205)_pad ,
		\542(246)_pad ,
		_w731_
	);
	LUT4 #(
		.INIT('h1e4b)
	) name524 (
		\18(5)_pad ,
		\41(12)_pad ,
		\4526(205)_pad ,
		\542(246)_pad ,
		_w732_
	);
	LUT2 #(
		.INIT('h1)
	) name525 (
		_w421_,
		_w422_,
		_w733_
	);
	LUT3 #(
		.INIT('h80)
	) name526 (
		_w490_,
		_w492_,
		_w494_,
		_w734_
	);
	LUT4 #(
		.INIT('h0f0e)
	) name527 (
		_w421_,
		_w422_,
		_w495_,
		_w734_,
		_w735_
	);
	LUT4 #(
		.INIT('h7f00)
	) name528 (
		_w480_,
		_w489_,
		_w733_,
		_w735_,
		_w736_
	);
	LUT3 #(
		.INIT('h10)
	) name529 (
		_w421_,
		_w422_,
		_w495_,
		_w737_
	);
	LUT2 #(
		.INIT('h4)
	) name530 (
		_w422_,
		_w495_,
		_w738_
	);
	LUT3 #(
		.INIT('h10)
	) name531 (
		_w421_,
		_w734_,
		_w738_,
		_w739_
	);
	LUT4 #(
		.INIT('h007f)
	) name532 (
		_w480_,
		_w489_,
		_w737_,
		_w739_,
		_w740_
	);
	LUT2 #(
		.INIT('hb)
	) name533 (
		_w736_,
		_w740_,
		_w741_
	);
	LUT3 #(
		.INIT('h71)
	) name534 (
		\548(234)_pad ,
		_w416_,
		_w418_,
		_w742_
	);
	LUT4 #(
		.INIT('h0045)
	) name535 (
		_w472_,
		_w477_,
		_w479_,
		_w742_,
		_w743_
	);
	LUT3 #(
		.INIT('h17)
	) name536 (
		\548(234)_pad ,
		_w416_,
		_w491_,
		_w744_
	);
	LUT4 #(
		.INIT('h0017)
	) name537 (
		\548(234)_pad ,
		_w416_,
		_w491_,
		_w494_,
		_w745_
	);
	LUT3 #(
		.INIT('h70)
	) name538 (
		_w489_,
		_w743_,
		_w745_,
		_w746_
	);
	LUT4 #(
		.INIT('he800)
	) name539 (
		\548(234)_pad ,
		_w416_,
		_w491_,
		_w494_,
		_w747_
	);
	LUT4 #(
		.INIT('h8e00)
	) name540 (
		\548(234)_pad ,
		_w416_,
		_w418_,
		_w494_,
		_w748_
	);
	LUT4 #(
		.INIT('h4500)
	) name541 (
		_w472_,
		_w477_,
		_w479_,
		_w748_,
		_w749_
	);
	LUT3 #(
		.INIT('h13)
	) name542 (
		_w489_,
		_w747_,
		_w749_,
		_w750_
	);
	LUT2 #(
		.INIT('hb)
	) name543 (
		_w746_,
		_w750_,
		_w751_
	);
	LUT2 #(
		.INIT('h4)
	) name544 (
		_w481_,
		_w492_,
		_w752_
	);
	LUT4 #(
		.INIT('h7f00)
	) name545 (
		_w482_,
		_w486_,
		_w487_,
		_w752_,
		_w753_
	);
	LUT2 #(
		.INIT('h9)
	) name546 (
		_w490_,
		_w491_,
		_w754_
	);
	LUT3 #(
		.INIT('h70)
	) name547 (
		_w480_,
		_w753_,
		_w754_,
		_w755_
	);
	LUT4 #(
		.INIT('h4500)
	) name548 (
		_w472_,
		_w477_,
		_w479_,
		_w493_,
		_w756_
	);
	LUT2 #(
		.INIT('h8)
	) name549 (
		_w489_,
		_w756_,
		_w757_
	);
	LUT2 #(
		.INIT('he)
	) name550 (
		_w755_,
		_w757_,
		_w758_
	);
	LUT4 #(
		.INIT('h02fd)
	) name551 (
		_w480_,
		_w481_,
		_w488_,
		_w492_,
		_w759_
	);
	LUT4 #(
		.INIT('he21d)
	) name552 (
		\103(52)_pad ,
		\18(5)_pad ,
		\235(158)_pad ,
		\552(238)_pad ,
		_w760_
	);
	LUT3 #(
		.INIT('h8e)
	) name553 (
		\558(244)_pad ,
		_w473_,
		_w474_,
		_w761_
	);
	LUT4 #(
		.INIT('h888e)
	) name554 (
		\558(244)_pad ,
		_w473_,
		_w474_,
		_w730_,
		_w762_
	);
	LUT4 #(
		.INIT('he41b)
	) name555 (
		\18(5)_pad ,
		\23(6)_pad ,
		\236(159)_pad ,
		\554(240)_pad ,
		_w763_
	);
	LUT2 #(
		.INIT('h8)
	) name556 (
		_w482_,
		_w763_,
		_w764_
	);
	LUT3 #(
		.INIT('h8e)
	) name557 (
		\554(240)_pad ,
		_w467_,
		_w476_,
		_w765_
	);
	LUT4 #(
		.INIT('h1055)
	) name558 (
		_w760_,
		_w762_,
		_w764_,
		_w765_,
		_w766_
	);
	LUT4 #(
		.INIT('h8e00)
	) name559 (
		\554(240)_pad ,
		_w467_,
		_w476_,
		_w760_,
		_w767_
	);
	LUT3 #(
		.INIT('hb0)
	) name560 (
		_w762_,
		_w764_,
		_w767_,
		_w768_
	);
	LUT2 #(
		.INIT('he)
	) name561 (
		_w766_,
		_w768_,
		_w769_
	);
	LUT4 #(
		.INIT('he817)
	) name562 (
		\556(242)_pad ,
		_w475_,
		_w762_,
		_w763_,
		_w770_
	);
	LUT2 #(
		.INIT('h9)
	) name563 (
		_w482_,
		_w762_,
		_w771_
	);
	LUT4 #(
		.INIT('he0f4)
	) name564 (
		\18(5)_pad ,
		\41(12)_pad ,
		\4526(205)_pad ,
		\542(246)_pad ,
		_w772_
	);
	LUT2 #(
		.INIT('h6)
	) name565 (
		_w485_,
		_w772_,
		_w773_
	);
	LUT4 #(
		.INIT('h008e)
	) name566 (
		\548(234)_pad ,
		_w416_,
		_w418_,
		_w422_,
		_w774_
	);
	LUT3 #(
		.INIT('hc9)
	) name567 (
		_w421_,
		_w754_,
		_w774_,
		_w775_
	);
	LUT3 #(
		.INIT('h80)
	) name568 (
		_w480_,
		_w489_,
		_w775_,
		_w776_
	);
	LUT2 #(
		.INIT('h6)
	) name569 (
		_w418_,
		_w490_,
		_w777_
	);
	LUT3 #(
		.INIT('h2a)
	) name570 (
		_w422_,
		_w490_,
		_w492_,
		_w778_
	);
	LUT3 #(
		.INIT('h10)
	) name571 (
		_w742_,
		_w777_,
		_w778_,
		_w779_
	);
	LUT4 #(
		.INIT('h0516)
	) name572 (
		\548(234)_pad ,
		\550(236)_pad ,
		_w416_,
		_w417_,
		_w780_
	);
	LUT4 #(
		.INIT('h0100)
	) name573 (
		_w421_,
		_w422_,
		_w734_,
		_w780_,
		_w781_
	);
	LUT2 #(
		.INIT('h1)
	) name574 (
		_w779_,
		_w781_,
		_w782_
	);
	LUT4 #(
		.INIT('h0100)
	) name575 (
		_w421_,
		_w422_,
		_w734_,
		_w744_,
		_w783_
	);
	LUT3 #(
		.INIT('h8c)
	) name576 (
		_w742_,
		_w777_,
		_w778_,
		_w784_
	);
	LUT4 #(
		.INIT('h7077)
	) name577 (
		_w480_,
		_w489_,
		_w783_,
		_w784_,
		_w785_
	);
	LUT3 #(
		.INIT('h15)
	) name578 (
		_w776_,
		_w782_,
		_w785_,
		_w786_
	);
	LUT3 #(
		.INIT('h80)
	) name579 (
		_w482_,
		_w484_,
		_w485_,
		_w787_
	);
	LUT4 #(
		.INIT('h5501)
	) name580 (
		_w469_,
		_w477_,
		_w478_,
		_w787_,
		_w788_
	);
	LUT4 #(
		.INIT('h0054)
	) name581 (
		_w468_,
		_w477_,
		_w478_,
		_w787_,
		_w789_
	);
	LUT4 #(
		.INIT('h88fe)
	) name582 (
		\558(244)_pad ,
		_w473_,
		_w483_,
		_w474_,
		_w790_
	);
	LUT3 #(
		.INIT('h23)
	) name583 (
		_w474_,
		_w483_,
		_w485_,
		_w791_
	);
	LUT3 #(
		.INIT('hc4)
	) name584 (
		_w761_,
		_w790_,
		_w791_,
		_w792_
	);
	LUT4 #(
		.INIT('hfd57)
	) name585 (
		_w730_,
		_w788_,
		_w789_,
		_w792_,
		_w793_
	);
	LUT4 #(
		.INIT('h4cc8)
	) name586 (
		\558(244)_pad ,
		_w469_,
		_w473_,
		_w474_,
		_w794_
	);
	LUT4 #(
		.INIT('h4cc8)
	) name587 (
		\558(244)_pad ,
		_w468_,
		_w473_,
		_w474_,
		_w795_
	);
	LUT4 #(
		.INIT('h01ef)
	) name588 (
		_w477_,
		_w478_,
		_w794_,
		_w795_,
		_w796_
	);
	LUT4 #(
		.INIT('h2001)
	) name589 (
		\558(244)_pad ,
		_w468_,
		_w473_,
		_w474_,
		_w797_
	);
	LUT4 #(
		.INIT('h2001)
	) name590 (
		\558(244)_pad ,
		_w469_,
		_w473_,
		_w474_,
		_w798_
	);
	LUT4 #(
		.INIT('h0e1f)
	) name591 (
		_w477_,
		_w478_,
		_w797_,
		_w798_,
		_w799_
	);
	LUT4 #(
		.INIT('hcbbb)
	) name592 (
		_w730_,
		_w731_,
		_w796_,
		_w799_,
		_w800_
	);
	LUT2 #(
		.INIT('h8)
	) name593 (
		_w793_,
		_w800_,
		_w801_
	);
	LUT4 #(
		.INIT('h6996)
	) name594 (
		_w482_,
		_w495_,
		_w760_,
		_w763_,
		_w802_
	);
	LUT2 #(
		.INIT('h9)
	) name595 (
		_w485_,
		_w494_,
		_w803_
	);
	LUT4 #(
		.INIT('h9669)
	) name596 (
		_w786_,
		_w801_,
		_w802_,
		_w803_,
		_w804_
	);
	LUT2 #(
		.INIT('he)
	) name597 (
		\5(1)_pad ,
		\57(20)_pad ,
		_w805_
	);
	LUT4 #(
		.INIT('h8000)
	) name598 (
		\150(73)_pad ,
		\184(107)_pad ,
		\228(151)_pad ,
		\240(163)_pad ,
		_w806_
	);
	LUT4 #(
		.INIT('h7fff)
	) name599 (
		\150(73)_pad ,
		\184(107)_pad ,
		\228(151)_pad ,
		\240(163)_pad ,
		_w807_
	);
	LUT4 #(
		.INIT('h8000)
	) name600 (
		\152(75)_pad ,
		\210(133)_pad ,
		\218(141)_pad ,
		\230(153)_pad ,
		_w808_
	);
	LUT4 #(
		.INIT('h7fff)
	) name601 (
		\152(75)_pad ,
		\210(133)_pad ,
		\218(141)_pad ,
		\230(153)_pad ,
		_w809_
	);
	LUT4 #(
		.INIT('h8000)
	) name602 (
		\182(105)_pad ,
		\183(106)_pad ,
		\185(108)_pad ,
		\186(109)_pad ,
		_w810_
	);
	LUT4 #(
		.INIT('h7fff)
	) name603 (
		\182(105)_pad ,
		\183(106)_pad ,
		\185(108)_pad ,
		\186(109)_pad ,
		_w811_
	);
	LUT4 #(
		.INIT('h8000)
	) name604 (
		\162(85)_pad ,
		\172(95)_pad ,
		\188(111)_pad ,
		\199(122)_pad ,
		_w812_
	);
	LUT4 #(
		.INIT('h7fff)
	) name605 (
		\162(85)_pad ,
		\172(95)_pad ,
		\188(111)_pad ,
		\199(122)_pad ,
		_w813_
	);
	LUT4 #(
		.INIT('h9669)
	) name606 (
		_w426_,
		_w430_,
		_w442_,
		_w446_,
		_w814_
	);
	LUT2 #(
		.INIT('h6)
	) name607 (
		_w451_,
		_w814_,
		_w815_
	);
	LUT3 #(
		.INIT('h1d)
	) name608 (
		\115(60)_pad ,
		\18(5)_pad ,
		\227(150)_pad ,
		_w816_
	);
	LUT2 #(
		.INIT('h6)
	) name609 (
		_w455_,
		_w816_,
		_w817_
	);
	LUT4 #(
		.INIT('h6996)
	) name610 (
		_w432_,
		_w438_,
		_w460_,
		_w817_,
		_w818_
	);
	LUT2 #(
		.INIT('h9)
	) name611 (
		\211(134)_pad ,
		\212(135)_pad ,
		_w819_
	);
	LUT3 #(
		.INIT('h4c)
	) name612 (
		\12(3)_pad ,
		\18(5)_pad ,
		\9(2)_pad ,
		_w820_
	);
	LUT3 #(
		.INIT('h60)
	) name613 (
		\209(132)_pad ,
		_w819_,
		_w820_,
		_w821_
	);
	LUT2 #(
		.INIT('h6)
	) name614 (
		\215(138)_pad ,
		\216(139)_pad ,
		_w822_
	);
	LUT2 #(
		.INIT('h8)
	) name615 (
		_w820_,
		_w822_,
		_w823_
	);
	LUT2 #(
		.INIT('h6)
	) name616 (
		\213(136)_pad ,
		\214(137)_pad ,
		_w824_
	);
	LUT3 #(
		.INIT('h57)
	) name617 (
		_w820_,
		_w822_,
		_w824_,
		_w825_
	);
	LUT3 #(
		.INIT('h20)
	) name618 (
		_w820_,
		_w822_,
		_w824_,
		_w826_
	);
	LUT3 #(
		.INIT('h1b)
	) name619 (
		_w821_,
		_w825_,
		_w826_,
		_w827_
	);
	LUT4 #(
		.INIT('h0f9f)
	) name620 (
		\209(132)_pad ,
		_w819_,
		_w820_,
		_w824_,
		_w828_
	);
	LUT4 #(
		.INIT('h6000)
	) name621 (
		\209(132)_pad ,
		_w819_,
		_w820_,
		_w824_,
		_w829_
	);
	LUT3 #(
		.INIT('h02)
	) name622 (
		_w823_,
		_w828_,
		_w829_,
		_w830_
	);
	LUT4 #(
		.INIT('hbb0b)
	) name623 (
		_w815_,
		_w818_,
		_w827_,
		_w830_,
		_w831_
	);
	LUT4 #(
		.INIT('h9909)
	) name624 (
		_w815_,
		_w818_,
		_w827_,
		_w830_,
		_w832_
	);
	LUT4 #(
		.INIT('h6996)
	) name625 (
		_w414_,
		_w417_,
		_w419_,
		_w470_,
		_w833_
	);
	LUT3 #(
		.INIT('h69)
	) name626 (
		_w416_,
		_w467_,
		_w475_,
		_w834_
	);
	LUT3 #(
		.INIT('h27)
	) name627 (
		\18(5)_pad ,
		\239(162)_pad ,
		\44(13)_pad ,
		_w835_
	);
	LUT3 #(
		.INIT('h27)
	) name628 (
		\18(5)_pad ,
		\229(152)_pad ,
		\41(12)_pad ,
		_w836_
	);
	LUT2 #(
		.INIT('h6)
	) name629 (
		_w473_,
		_w836_,
		_w837_
	);
	LUT4 #(
		.INIT('h6996)
	) name630 (
		_w833_,
		_w834_,
		_w835_,
		_w837_,
		_w838_
	);
	LUT3 #(
		.INIT('h69)
	) name631 (
		_w366_,
		_w370_,
		_w375_,
		_w839_
	);
	LUT3 #(
		.INIT('he0)
	) name632 (
		\153(76)_pad ,
		\154(77)_pad ,
		\18(5)_pad ,
		_w840_
	);
	LUT4 #(
		.INIT('h153f)
	) name633 (
		\12(3)_pad ,
		\153(76)_pad ,
		\154(77)_pad ,
		\9(2)_pad ,
		_w841_
	);
	LUT3 #(
		.INIT('h6a)
	) name634 (
		_w362_,
		_w840_,
		_w841_,
		_w842_
	);
	LUT3 #(
		.INIT('h35)
	) name635 (
		\141(70)_pad ,
		\161(84)_pad ,
		\18(5)_pad ,
		_w843_
	);
	LUT2 #(
		.INIT('h6)
	) name636 (
		_w379_,
		_w843_,
		_w844_
	);
	LUT3 #(
		.INIT('he0)
	) name637 (
		\155(78)_pad ,
		\156(79)_pad ,
		\18(5)_pad ,
		_w845_
	);
	LUT4 #(
		.INIT('h153f)
	) name638 (
		\12(3)_pad ,
		\155(78)_pad ,
		\156(79)_pad ,
		\9(2)_pad ,
		_w846_
	);
	LUT2 #(
		.INIT('h8)
	) name639 (
		_w845_,
		_w846_,
		_w847_
	);
	LUT4 #(
		.INIT('h6996)
	) name640 (
		_w839_,
		_w842_,
		_w844_,
		_w847_,
		_w848_
	);
	LUT2 #(
		.INIT('h4)
	) name641 (
		_w838_,
		_w848_,
		_w849_
	);
	LUT2 #(
		.INIT('h7)
	) name642 (
		_w832_,
		_w849_,
		_w850_
	);
	LUT3 #(
		.INIT('h69)
	) name643 (
		_w283_,
		_w285_,
		_w289_,
		_w851_
	);
	LUT3 #(
		.INIT('h82)
	) name644 (
		\18(5)_pad ,
		\438(274)_pad ,
		\440(277)_pad ,
		_w852_
	);
	LUT3 #(
		.INIT('h21)
	) name645 (
		\1455(166)_pad ,
		\18(5)_pad ,
		\2204(174)_pad ,
		_w853_
	);
	LUT2 #(
		.INIT('h1)
	) name646 (
		_w852_,
		_w853_,
		_w854_
	);
	LUT3 #(
		.INIT('hd1)
	) name647 (
		\114(59)_pad ,
		\18(5)_pad ,
		\450(288)_pad ,
		_w855_
	);
	LUT3 #(
		.INIT('h69)
	) name648 (
		_w295_,
		_w299_,
		_w855_,
		_w856_
	);
	LUT3 #(
		.INIT('h69)
	) name649 (
		_w851_,
		_w854_,
		_w856_,
		_w857_
	);
	LUT2 #(
		.INIT('h6)
	) name650 (
		_w227_,
		_w245_,
		_w858_
	);
	LUT4 #(
		.INIT('h6996)
	) name651 (
		_w224_,
		_w232_,
		_w237_,
		_w858_,
		_w859_
	);
	LUT3 #(
		.INIT('h72)
	) name652 (
		\18(5)_pad ,
		\560(248)_pad ,
		\69(30)_pad ,
		_w860_
	);
	LUT2 #(
		.INIT('h6)
	) name653 (
		_w222_,
		_w860_,
		_w861_
	);
	LUT3 #(
		.INIT('h72)
	) name654 (
		\18(5)_pad ,
		\542(246)_pad ,
		\70(31)_pad ,
		_w862_
	);
	LUT4 #(
		.INIT('h6996)
	) name655 (
		_w239_,
		_w242_,
		_w861_,
		_w862_,
		_w863_
	);
	LUT3 #(
		.INIT('h14)
	) name656 (
		_w857_,
		_w859_,
		_w863_,
		_w864_
	);
	LUT4 #(
		.INIT('h6996)
	) name657 (
		_w310_,
		_w318_,
		_w328_,
		_w334_,
		_w865_
	);
	LUT3 #(
		.INIT('h69)
	) name658 (
		_w322_,
		_w326_,
		_w332_,
		_w866_
	);
	LUT3 #(
		.INIT('h72)
	) name659 (
		\18(5)_pad ,
		\496(271)_pad ,
		\82(41)_pad ,
		_w867_
	);
	LUT2 #(
		.INIT('h6)
	) name660 (
		_w315_,
		_w867_,
		_w868_
	);
	LUT4 #(
		.INIT('h9669)
	) name661 (
		_w312_,
		_w865_,
		_w866_,
		_w868_,
		_w869_
	);
	LUT3 #(
		.INIT('h8d)
	) name662 (
		\18(5)_pad ,
		\540(227)_pad ,
		\58(21)_pad ,
		_w870_
	);
	LUT2 #(
		.INIT('h6)
	) name663 (
		_w266_,
		_w870_,
		_w871_
	);
	LUT4 #(
		.INIT('h9669)
	) name664 (
		_w218_,
		_w252_,
		_w260_,
		_w871_,
		_w872_
	);
	LUT2 #(
		.INIT('h9)
	) name665 (
		_w210_,
		_w215_,
		_w873_
	);
	LUT3 #(
		.INIT('h69)
	) name666 (
		_w212_,
		_w263_,
		_w270_,
		_w874_
	);
	LUT4 #(
		.INIT('h1441)
	) name667 (
		_w869_,
		_w872_,
		_w873_,
		_w874_,
		_w875_
	);
	LUT2 #(
		.INIT('h8)
	) name668 (
		_w864_,
		_w875_,
		_w876_
	);
	LUT2 #(
		.INIT('h7)
	) name669 (
		_w864_,
		_w875_,
		_w877_
	);
	LUT4 #(
		.INIT('h6996)
	) name670 (
		_w223_,
		_w236_,
		_w238_,
		_w244_,
		_w878_
	);
	LUT3 #(
		.INIT('h69)
	) name671 (
		_w221_,
		_w226_,
		_w231_,
		_w879_
	);
	LUT3 #(
		.INIT('h27)
	) name672 (
		\18(5)_pad ,
		\208(131)_pad ,
		\44(13)_pad ,
		_w880_
	);
	LUT3 #(
		.INIT('h27)
	) name673 (
		\18(5)_pad ,
		\198(121)_pad ,
		\41(12)_pad ,
		_w881_
	);
	LUT2 #(
		.INIT('h6)
	) name674 (
		_w241_,
		_w881_,
		_w882_
	);
	LUT4 #(
		.INIT('h6996)
	) name675 (
		_w878_,
		_w879_,
		_w880_,
		_w882_,
		_w883_
	);
	LUT4 #(
		.INIT('h9669)
	) name676 (
		_w209_,
		_w217_,
		_w259_,
		_w262_,
		_w884_
	);
	LUT2 #(
		.INIT('h6)
	) name677 (
		_w265_,
		_w884_,
		_w885_
	);
	LUT3 #(
		.INIT('h1d)
	) name678 (
		\115(60)_pad ,
		\18(5)_pad ,
		\197(120)_pad ,
		_w886_
	);
	LUT2 #(
		.INIT('h6)
	) name679 (
		_w251_,
		_w886_,
		_w887_
	);
	LUT4 #(
		.INIT('h6996)
	) name680 (
		_w211_,
		_w214_,
		_w269_,
		_w887_,
		_w888_
	);
	LUT2 #(
		.INIT('h2)
	) name681 (
		_w885_,
		_w888_,
		_w889_
	);
	LUT2 #(
		.INIT('h4)
	) name682 (
		_w885_,
		_w888_,
		_w890_
	);
	LUT2 #(
		.INIT('h9)
	) name683 (
		\164(87)_pad ,
		\165(88)_pad ,
		_w891_
	);
	LUT3 #(
		.INIT('h90)
	) name684 (
		\164(87)_pad ,
		\165(88)_pad ,
		\170(93)_pad ,
		_w892_
	);
	LUT3 #(
		.INIT('h06)
	) name685 (
		\164(87)_pad ,
		\165(88)_pad ,
		\170(93)_pad ,
		_w893_
	);
	LUT2 #(
		.INIT('h2)
	) name686 (
		_w820_,
		_w893_,
		_w894_
	);
	LUT3 #(
		.INIT('h48)
	) name687 (
		\170(93)_pad ,
		_w820_,
		_w891_,
		_w895_
	);
	LUT3 #(
		.INIT('he0)
	) name688 (
		\166(89)_pad ,
		\167(90)_pad ,
		\18(5)_pad ,
		_w896_
	);
	LUT4 #(
		.INIT('h153f)
	) name689 (
		\12(3)_pad ,
		\166(89)_pad ,
		\167(90)_pad ,
		\9(2)_pad ,
		_w897_
	);
	LUT2 #(
		.INIT('h8)
	) name690 (
		_w896_,
		_w897_,
		_w898_
	);
	LUT3 #(
		.INIT('he0)
	) name691 (
		\168(91)_pad ,
		\169(92)_pad ,
		\18(5)_pad ,
		_w899_
	);
	LUT4 #(
		.INIT('h153f)
	) name692 (
		\12(3)_pad ,
		\168(91)_pad ,
		\169(92)_pad ,
		\9(2)_pad ,
		_w900_
	);
	LUT2 #(
		.INIT('h8)
	) name693 (
		_w899_,
		_w900_,
		_w901_
	);
	LUT3 #(
		.INIT('hde)
	) name694 (
		_w895_,
		_w898_,
		_w901_,
		_w902_
	);
	LUT2 #(
		.INIT('h1)
	) name695 (
		_w895_,
		_w901_,
		_w903_
	);
	LUT3 #(
		.INIT('h40)
	) name696 (
		_w892_,
		_w899_,
		_w900_,
		_w904_
	);
	LUT3 #(
		.INIT('h4c)
	) name697 (
		_w894_,
		_w898_,
		_w904_,
		_w905_
	);
	LUT3 #(
		.INIT('h8a)
	) name698 (
		_w902_,
		_w903_,
		_w905_,
		_w906_
	);
	LUT3 #(
		.INIT('h01)
	) name699 (
		_w889_,
		_w890_,
		_w906_,
		_w907_
	);
	LUT3 #(
		.INIT('h69)
	) name700 (
		_w311_,
		_w321_,
		_w331_,
		_w908_
	);
	LUT3 #(
		.INIT('he0)
	) name701 (
		\173(96)_pad ,
		\174(97)_pad ,
		\18(5)_pad ,
		_w909_
	);
	LUT4 #(
		.INIT('h153f)
	) name702 (
		\12(3)_pad ,
		\173(96)_pad ,
		\174(97)_pad ,
		\9(2)_pad ,
		_w910_
	);
	LUT3 #(
		.INIT('h6a)
	) name703 (
		_w309_,
		_w909_,
		_w910_,
		_w911_
	);
	LUT3 #(
		.INIT('h1d)
	) name704 (
		\141(70)_pad ,
		\18(5)_pad ,
		\181(104)_pad ,
		_w912_
	);
	LUT2 #(
		.INIT('h6)
	) name705 (
		_w333_,
		_w912_,
		_w913_
	);
	LUT3 #(
		.INIT('he0)
	) name706 (
		\175(98)_pad ,
		\176(99)_pad ,
		\18(5)_pad ,
		_w914_
	);
	LUT4 #(
		.INIT('h153f)
	) name707 (
		\12(3)_pad ,
		\175(98)_pad ,
		\176(99)_pad ,
		\9(2)_pad ,
		_w915_
	);
	LUT2 #(
		.INIT('h8)
	) name708 (
		_w914_,
		_w915_,
		_w916_
	);
	LUT4 #(
		.INIT('h6996)
	) name709 (
		_w908_,
		_w911_,
		_w913_,
		_w916_,
		_w917_
	);
	LUT4 #(
		.INIT('h0900)
	) name710 (
		_w885_,
		_w888_,
		_w906_,
		_w917_,
		_w918_
	);
	LUT2 #(
		.INIT('hb)
	) name711 (
		_w883_,
		_w918_,
		_w919_
	);
	LUT2 #(
		.INIT('h4)
	) name712 (
		_w883_,
		_w917_,
		_w920_
	);
	LUT4 #(
		.INIT('h8000)
	) name713 (
		_w806_,
		_w808_,
		_w810_,
		_w812_,
		_w921_
	);
	LUT3 #(
		.INIT('hd0)
	) name714 (
		_w815_,
		_w818_,
		_w921_,
		_w922_
	);
	LUT4 #(
		.INIT('h8000)
	) name715 (
		_w831_,
		_w849_,
		_w920_,
		_w922_,
		_w923_
	);
	LUT3 #(
		.INIT('h7f)
	) name716 (
		_w876_,
		_w907_,
		_w923_,
		_w924_
	);
	LUT3 #(
		.INIT('h6a)
	) name717 (
		\38(11)_pad ,
		\440(277)_pad ,
		\4528(206)_pad ,
		_w925_
	);
	LUT3 #(
		.INIT('h0b)
	) name718 (
		\442(280)_pad ,
		_w515_,
		_w925_,
		_w926_
	);
	LUT4 #(
		.INIT('hef00)
	) name719 (
		_w413_,
		_w509_,
		_w520_,
		_w926_,
		_w927_
	);
	LUT4 #(
		.INIT('h0e0f)
	) name720 (
		_w413_,
		_w509_,
		_w516_,
		_w520_,
		_w928_
	);
	LUT3 #(
		.INIT('hce)
	) name721 (
		_w925_,
		_w927_,
		_w928_,
		_w929_
	);
	LUT3 #(
		.INIT('h0b)
	) name722 (
		\442(280)_pad ,
		_w515_,
		_w654_,
		_w930_
	);
	LUT4 #(
		.INIT('hef00)
	) name723 (
		_w413_,
		_w509_,
		_w520_,
		_w930_,
		_w931_
	);
	LUT3 #(
		.INIT('hf1)
	) name724 (
		_w648_,
		_w928_,
		_w931_,
		_w932_
	);
	assign \252(3450)_pad  = _w280_ ;
	assign \258(3122)_pad  = _w356_ ;
	assign \270(3109)_pad  = _w526_ ;
	assign \278(536)_pad  = _w527_ ;
	assign \281(547)_pad  = _w528_ ;
	assign \284(384)_pad  = _w529_ ;
	assign \286(419)_pad  = _w27_ ;
	assign \292(392)_pad  = _w528_ ;
	assign \295(3352)_pad  = _w531_ ;
	assign \298(3387)_pad  = _w542_ ;
	assign \301(3388)_pad  = _w550_ ;
	assign \304(3390)_pad  = _w554_ ;
	assign \307(3389)_pad  = _w555_ ;
	assign \310(3393)_pad  = _w563_ ;
	assign \313(3396)_pad  = _w568_ ;
	assign \316(3397)_pad  = _w573_ ;
	assign \319(3398)_pad  = _w574_ ;
	assign \321(3715)_pad  = _w599_ ;
	assign \324(3363)_pad  = _w604_ ;
	assign \327(3408)_pad  = _w607_ ;
	assign \330(3411)_pad  = _w615_ ;
	assign \333(3416)_pad  = _w620_ ;
	assign \336(3412)_pad  = _w626_ ;
	assign \338(3716)_pad  = _w656_ ;
	assign \344(3382)_pad  = _w666_ ;
	assign \347(3420)_pad  = _w677_ ;
	assign \350(3421)_pad  = _w684_ ;
	assign \353(3425)_pad  = _w690_ ;
	assign \356(3424)_pad  = _w691_ ;
	assign \359(3426)_pad  = _w695_ ;
	assign \362(3429)_pad  = _w696_ ;
	assign \365(3430)_pad  = _w698_ ;
	assign \368(3431)_pad  = _w699_ ;
	assign \370(3718)_pad  = _w729_ ;
	assign \373(2994)_pad  = _w732_ ;
	assign \376(3206)_pad  = _w741_ ;
	assign \379(3207)_pad  = _w751_ ;
	assign \382(3148)_pad  = _w758_ ;
	assign \385(3151)_pad  = _w759_ ;
	assign \388(3093)_pad  = _w769_ ;
	assign \391(3094)_pad  = _w770_ ;
	assign \394(3095)_pad  = _w771_ ;
	assign \397(3097)_pad  = _w773_ ;
	assign \399(3717)_pad  = _w804_ ;
	assign \402(395)_pad  = _w805_ ;
	assign \404(390)_pad  = _w807_ ;
	assign \406(388)_pad  = _w809_ ;
	assign \408(385)_pad  = _w811_ ;
	assign \410(387)_pad  = _w813_ ;
	assign \412(3369)_pad  = _w850_ ;
	assign \414(3338)_pad  = _w877_ ;
	assign \416(3368)_pad  = _w919_ ;
	assign \418(3449)_pad  = _w924_ ;
	assign \419(3444)_pad  = _w929_ ;
	assign \422(3451)_pad  = _w932_ ;
endmodule;