module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 ;
  wire n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 ;
  assign n8 = x0 & ~x1 ;
  assign n9 = x3 & x4 ;
  assign n10 = n8 & n9 ;
  assign n11 = x1 & x3 ;
  assign n12 = x4 & n11 ;
  assign n13 = ~n10 & ~n12 ;
  assign n14 = ~x2 & ~n13 ;
  assign n15 = ~x1 & x3 ;
  assign n16 = x4 & n15 ;
  assign n17 = ~x3 & ~x4 ;
  assign n18 = ~n9 & ~n17 ;
  assign n19 = x1 & ~n18 ;
  assign n20 = ~n16 & ~n19 ;
  assign n21 = x2 & ~n20 ;
  assign n22 = ~n14 & ~n21 ;
  assign n23 = ~x0 & ~n9 ;
  assign n24 = ~x0 & ~n23 ;
  assign n25 = ~x1 & ~n24 ;
  assign n26 = ~x3 & ~n17 ;
  assign n27 = x1 & ~n26 ;
  assign n28 = ~n25 & ~n27 ;
  assign n29 = ~x2 & ~n28 ;
  assign n30 = ~x3 & x4 ;
  assign n31 = ~x3 & ~n30 ;
  assign n32 = x1 & ~n31 ;
  assign n33 = x1 & ~n32 ;
  assign n34 = x2 & ~n33 ;
  assign n35 = ~n29 & ~n34 ;
  assign n36 = ~x0 & ~n18 ;
  assign n37 = x3 & ~n9 ;
  assign n38 = x0 & ~n37 ;
  assign n39 = ~n36 & ~n38 ;
  assign n40 = x1 & ~n39 ;
  assign n41 = ~n25 & ~n40 ;
  assign n42 = ~x2 & ~n41 ;
  assign n43 = ~x2 & ~n42 ;
  assign n44 = ~x0 & ~x3 ;
  assign n45 = ~n30 & n44 ;
  assign n46 = x0 & ~n18 ;
  assign n47 = ~n45 & ~n46 ;
  assign n48 = ~x1 & ~n47 ;
  assign n49 = ~n27 & ~n48 ;
  assign n50 = ~x2 & ~n49 ;
  assign n51 = x2 & ~n26 ;
  assign n52 = ~n50 & ~n51 ;
  assign n53 = ~x0 & x3 ;
  assign n54 = x4 & x5 ;
  assign n55 = n53 & n54 ;
  assign n56 = x3 & ~x6 ;
  assign n57 = ~n9 & n56 ;
  assign n58 = x3 & ~x5 ;
  assign n59 = ~n9 & n58 ;
  assign n60 = x3 & x5 ;
  assign n61 = ~n59 & ~n60 ;
  assign n62 = x6 & ~n61 ;
  assign n63 = ~n57 & ~n62 ;
  assign n64 = x0 & ~n63 ;
  assign n65 = ~n55 & ~n64 ;
  assign n66 = x1 & ~n65 ;
  assign n67 = ~x2 & ~n66 ;
  assign n68 = x0 & ~n26 ;
  assign n69 = x0 & ~n68 ;
  assign n70 = x2 & ~n69 ;
  assign n71 = ~n67 & ~n70 ;
  assign n72 = x3 & x6 ;
  assign n73 = ~n57 & ~n72 ;
  assign n74 = x1 & ~n73 ;
  assign n75 = ~x2 & ~n74 ;
  assign n76 = x1 & ~n27 ;
  assign n77 = x2 & ~n76 ;
  assign n78 = ~n75 & ~n77 ;
  assign n79 = ~x1 & ~n9 ;
  assign n80 = ~n17 & n79 ;
  assign n81 = ~n17 & n23 ;
  assign n82 = x0 & ~n31 ;
  assign n83 = ~n81 & ~n82 ;
  assign n84 = x1 & ~n83 ;
  assign n85 = ~n80 & ~n84 ;
  assign n86 = ~x2 & ~n85 ;
  assign n87 = x2 & x3 ;
  assign n88 = x4 & n87 ;
  assign n89 = ~n86 & ~n88 ;
  assign n90 = ~x1 & ~x2 ;
  assign n91 = ~n25 & n90 ;
  assign n92 = x1 & ~n47 ;
  assign n93 = ~n10 & ~n92 ;
  assign n94 = x2 & ~n93 ;
  assign n95 = ~n91 & ~n94 ;
  assign n96 = ~x0 & ~n26 ;
  assign n97 = ~x0 & ~n96 ;
  assign n98 = x1 & ~n97 ;
  assign n99 = x1 & ~x2 ;
  assign n100 = ~n98 & n99 ;
  assign n101 = x1 & x2 ;
  assign n102 = ~n18 & n101 ;
  assign n103 = ~n100 & ~n102 ;
  assign n104 = ~n79 & ~n98 ;
  assign n105 = ~x2 & ~n104 ;
  assign n106 = ~n34 & ~n105 ;
  assign n107 = ~n53 & ~n82 ;
  assign n108 = x1 & ~n107 ;
  assign n109 = ~x2 & ~n80 ;
  assign n110 = ~n108 & n109 ;
  assign n111 = ~n51 & ~n110 ;
  assign n112 = ~x0 & ~n31 ;
  assign n113 = ~x0 & ~n112 ;
  assign n114 = ~x1 & ~n113 ;
  assign n115 = ~x1 & ~n114 ;
  assign n116 = ~x2 & ~n115 ;
  assign n117 = ~x2 & ~n116 ;
  assign n118 = ~x1 & ~n107 ;
  assign n119 = ~n32 & ~n118 ;
  assign n120 = ~x2 & ~n119 ;
  assign n121 = ~x1 & x4 ;
  assign n122 = x1 & ~n37 ;
  assign n123 = ~n121 & ~n122 ;
  assign n124 = x2 & ~n123 ;
  assign n125 = ~n120 & ~n124 ;
  assign n126 = x0 & ~n82 ;
  assign n127 = x2 & ~n126 ;
  assign n128 = x2 & ~n127 ;
  assign n129 = x2 & ~n113 ;
  assign n130 = x2 & ~n129 ;
  assign n131 = ~x0 & ~n37 ;
  assign n132 = ~x0 & ~n131 ;
  assign n133 = ~x1 & ~n132 ;
  assign n134 = ~x1 & ~n133 ;
  assign n135 = x2 & ~n134 ;
  assign n136 = x2 & ~n135 ;
  assign n137 = x0 & ~n38 ;
  assign n138 = ~x1 & ~n137 ;
  assign n139 = ~x1 & ~n138 ;
  assign n140 = x2 & ~n139 ;
  assign n141 = x2 & ~n140 ;
  assign n142 = x1 & ~n137 ;
  assign n143 = x1 & ~n142 ;
  assign n144 = x2 & ~n143 ;
  assign n145 = x2 & ~n144 ;
  assign n146 = x1 & ~n132 ;
  assign n147 = x1 & ~n146 ;
  assign n148 = x2 & ~n147 ;
  assign n149 = x2 & ~n148 ;
  assign n150 = x2 & ~n31 ;
  assign n151 = x2 & ~n150 ;
  assign n152 = x0 & x1 ;
  assign n153 = ~n61 & n152 ;
  assign n154 = n8 & ~n38 ;
  assign n155 = ~x2 & ~n154 ;
  assign n156 = ~n153 & n155 ;
  assign n157 = x1 & ~n24 ;
  assign n158 = ~n79 & ~n157 ;
  assign n159 = x2 & ~n158 ;
  assign n160 = ~n156 & ~n159 ;
  assign n161 = x5 & n9 ;
  assign n162 = ~x6 & ~n161 ;
  assign n163 = ~x6 & ~n162 ;
  assign n164 = x0 & ~n163 ;
  assign n165 = x0 & ~n164 ;
  assign n166 = x1 & ~n165 ;
  assign n167 = ~n138 & ~n166 ;
  assign n168 = ~x2 & ~n167 ;
  assign n169 = ~x2 & ~n168 ;
  assign n170 = ~n63 & n152 ;
  assign n171 = ~x2 & ~n170 ;
  assign n172 = ~n159 & ~n171 ;
  assign n173 = ~x1 & ~n97 ;
  assign n174 = x1 & ~n69 ;
  assign n175 = ~n173 & ~n174 ;
  assign n176 = ~x2 & ~n175 ;
  assign n177 = ~x2 & ~n176 ;
  assign n178 = ~x1 & ~n69 ;
  assign n179 = ~x1 & ~n178 ;
  assign n180 = ~x2 & ~n179 ;
  assign n181 = ~x2 & ~n180 ;
  assign y0 = ~n22 ;
  assign y1 = n35 ;
  assign y2 = n43 ;
  assign y3 = n52 ;
  assign y4 = n71 ;
  assign y5 = n78 ;
  assign y6 = ~n89 ;
  assign y7 = ~n95 ;
  assign y8 = ~n103 ;
  assign y9 = n106 ;
  assign y10 = n111 ;
  assign y11 = n117 ;
  assign y12 = ~n125 ;
  assign y13 = n128 ;
  assign y14 = n130 ;
  assign y15 = n136 ;
  assign y16 = n141 ;
  assign y17 = n145 ;
  assign y18 = n149 ;
  assign y19 = n151 ;
  assign y20 = n160 ;
  assign y21 = n169 ;
  assign y22 = n172 ;
  assign y23 = ~1'b0 ;
  assign y24 = n177 ;
  assign y25 = n181 ;
endmodule
