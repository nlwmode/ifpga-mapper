module top( a_pad , b_pad , c_pad , d_pad , e_pad , f_pad , g_pad , i_pad , j_pad , k_pad , l_pad , m_pad , n_pad , o_pad , p_pad , q_pad , r_pad , s_pad , t_pad , u_pad , v_pad , w_pad , x_pad , y_pad , z_pad );
  input a_pad ;
  input b_pad ;
  input c_pad ;
  input d_pad ;
  input e_pad ;
  input f_pad ;
  input g_pad ;
  input i_pad ;
  input j_pad ;
  input k_pad ;
  input l_pad ;
  input m_pad ;
  input n_pad ;
  input o_pad ;
  output p_pad ;
  output q_pad ;
  output r_pad ;
  output s_pad ;
  output t_pad ;
  output u_pad ;
  output v_pad ;
  output w_pad ;
  output x_pad ;
  output y_pad ;
  output z_pad ;
  wire n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 ;
  assign n16 = ~c_pad & f_pad ;
  assign n17 = c_pad & e_pad ;
  assign n18 = ~n16 & ~n17 ;
  assign n15 = e_pad & f_pad ;
  assign n19 = ~d_pad & ~n15 ;
  assign n20 = ~n18 & n19 ;
  assign n21 = ~a_pad & ~b_pad ;
  assign n22 = ~d_pad & ~e_pad ;
  assign n23 = ~o_pad & n22 ;
  assign n24 = n16 & n23 ;
  assign n25 = n21 & n24 ;
  assign n26 = a_pad & n24 ;
  assign n27 = ~b_pad & n26 ;
  assign n28 = ~a_pad & b_pad ;
  assign n29 = n24 & n28 ;
  assign n30 = b_pad & n26 ;
  assign n34 = b_pad & ~m_pad ;
  assign n39 = a_pad & n34 ;
  assign n35 = ~b_pad & ~k_pad ;
  assign n40 = l_pad & ~n21 ;
  assign n41 = ~n35 & n40 ;
  assign n42 = ~n39 & n41 ;
  assign n36 = a_pad & ~l_pad ;
  assign n37 = ~n34 & n36 ;
  assign n38 = ~n35 & n37 ;
  assign n32 = f_pad & ~n_pad ;
  assign n33 = o_pad & n32 ;
  assign n31 = j_pad & n21 ;
  assign n43 = ~i_pad & ~n31 ;
  assign n44 = n33 & n43 ;
  assign n45 = ~n38 & n44 ;
  assign n46 = ~n42 & n45 ;
  assign n47 = ~c_pad & ~n46 ;
  assign n48 = ~f_pad & ~o_pad ;
  assign n49 = c_pad & ~n48 ;
  assign n50 = ~d_pad & e_pad ;
  assign n51 = ~n49 & n50 ;
  assign n52 = ~n47 & n51 ;
  assign n53 = ~c_pad & ~n33 ;
  assign n54 = n51 & ~n53 ;
  assign n55 = g_pad & o_pad ;
  assign n56 = c_pad & f_pad ;
  assign n57 = ~d_pad & g_pad ;
  assign n58 = ~n56 & n57 ;
  assign p_pad = ~n20 ;
  assign q_pad = n20 ;
  assign r_pad = n25 ;
  assign s_pad = n27 ;
  assign t_pad = n29 ;
  assign u_pad = n30 ;
  assign v_pad = n52 ;
  assign w_pad = n24 ;
  assign x_pad = n54 ;
  assign y_pad = n55 ;
  assign z_pad = n58 ;
endmodule
