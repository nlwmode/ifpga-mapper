module top( \1(0)_pad  , \107(12)_pad  , \116(13)_pad  , \124(14)_pad  , \125(15)_pad  , \128(16)_pad  , \13(1)_pad  , \132(17)_pad  , \137(18)_pad  , \143(19)_pad  , \150(20)_pad  , \159(21)_pad  , \169(22)_pad  , \1698(48)_pad  , \179(23)_pad  , \190(24)_pad  , \20(2)_pad  , \200(25)_pad  , \213(26)_pad  , \222(27)_pad  , \223(28)_pad  , \226(29)_pad  , \232(30)_pad  , \238(31)_pad  , \244(32)_pad  , \250(33)_pad  , \257(34)_pad  , \264(35)_pad  , \270(36)_pad  , \274(37)_pad  , \283(38)_pad  , \2897(49)_pad  , \294(39)_pad  , \303(40)_pad  , \311(41)_pad  , \317(42)_pad  , \322(43)_pad  , \326(44)_pad  , \329(45)_pad  , \33(3)_pad  , \330(46)_pad  , \343(47)_pad  , \41(4)_pad  , \45(5)_pad  , \50(6)_pad  , \58(7)_pad  , \68(8)_pad  , \77(9)_pad  , \87(10)_pad  , \97(11)_pad  , \2690(1611)  , \2709(1587)  , \353(405)_pad  , \355(399)_pad  , \358(1161)_pad  , \361(940)_pad  , \364(1484)_pad  , \367(1585)_pad  , \369(1321)_pad  , \372(1243)_pad  , \381(1626)_pad  , \384(1553)_pad  , \387(1616)_pad  , \390(1603)_pad  , \393(1605)_pad  , \396(1504)_pad  , \399(1428)_pad  , \402(1718)_pad  , \404(1714)  , \407(1657)_pad  , \409(1670)_pad  , \605(1186)  );
  input \1(0)_pad  ;
  input \107(12)_pad  ;
  input \116(13)_pad  ;
  input \124(14)_pad  ;
  input \125(15)_pad  ;
  input \128(16)_pad  ;
  input \13(1)_pad  ;
  input \132(17)_pad  ;
  input \137(18)_pad  ;
  input \143(19)_pad  ;
  input \150(20)_pad  ;
  input \159(21)_pad  ;
  input \169(22)_pad  ;
  input \1698(48)_pad  ;
  input \179(23)_pad  ;
  input \190(24)_pad  ;
  input \20(2)_pad  ;
  input \200(25)_pad  ;
  input \213(26)_pad  ;
  input \222(27)_pad  ;
  input \223(28)_pad  ;
  input \226(29)_pad  ;
  input \232(30)_pad  ;
  input \238(31)_pad  ;
  input \244(32)_pad  ;
  input \250(33)_pad  ;
  input \257(34)_pad  ;
  input \264(35)_pad  ;
  input \270(36)_pad  ;
  input \274(37)_pad  ;
  input \283(38)_pad  ;
  input \2897(49)_pad  ;
  input \294(39)_pad  ;
  input \303(40)_pad  ;
  input \311(41)_pad  ;
  input \317(42)_pad  ;
  input \322(43)_pad  ;
  input \326(44)_pad  ;
  input \329(45)_pad  ;
  input \33(3)_pad  ;
  input \330(46)_pad  ;
  input \343(47)_pad  ;
  input \41(4)_pad  ;
  input \45(5)_pad  ;
  input \50(6)_pad  ;
  input \58(7)_pad  ;
  input \68(8)_pad  ;
  input \77(9)_pad  ;
  input \87(10)_pad  ;
  input \97(11)_pad  ;
  output \2690(1611)  ;
  output \2709(1587)  ;
  output \353(405)_pad  ;
  output \355(399)_pad  ;
  output \358(1161)_pad  ;
  output \361(940)_pad  ;
  output \364(1484)_pad  ;
  output \367(1585)_pad  ;
  output \369(1321)_pad  ;
  output \372(1243)_pad  ;
  output \381(1626)_pad  ;
  output \384(1553)_pad  ;
  output \387(1616)_pad  ;
  output \390(1603)_pad  ;
  output \393(1605)_pad  ;
  output \396(1504)_pad  ;
  output \399(1428)_pad  ;
  output \402(1718)_pad  ;
  output \404(1714)  ;
  output \407(1657)_pad  ;
  output \409(1670)_pad  ;
  output \605(1186)  ;
  wire n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 ;
  assign n51 = \13(1)_pad  & ~\20(2)_pad  ;
  assign n52 = ~\1(0)_pad  & \213(26)_pad  ;
  assign n53 = n51 & n52 ;
  assign n100 = \343(47)_pad  & n53 ;
  assign n190 = ~\33(3)_pad  & \97(11)_pad  ;
  assign n189 = \283(38)_pad  & \33(3)_pad  ;
  assign n191 = ~\20(2)_pad  & ~n189 ;
  assign n192 = ~n190 & n191 ;
  assign n54 = \1(0)_pad  & \13(1)_pad  ;
  assign n55 = \1(0)_pad  & \20(2)_pad  ;
  assign n56 = \33(3)_pad  & n55 ;
  assign n57 = ~n54 & ~n56 ;
  assign n188 = ~\116(13)_pad  & \20(2)_pad  ;
  assign n193 = ~n57 & ~n188 ;
  assign n194 = ~n192 & n193 ;
  assign n69 = \13(1)_pad  & \20(2)_pad  ;
  assign n70 = ~\1(0)_pad  & n69 ;
  assign n186 = ~\116(13)_pad  & n70 ;
  assign n172 = ~\33(3)_pad  & ~n69 ;
  assign n173 = ~\1(0)_pad  & ~n172 ;
  assign n174 = n57 & ~n173 ;
  assign n187 = \116(13)_pad  & n174 ;
  assign n195 = ~n186 & ~n187 ;
  assign n196 = ~n194 & n195 ;
  assign n77 = \33(3)_pad  & \41(4)_pad  ;
  assign n78 = n54 & ~n77 ;
  assign n83 = \274(37)_pad  & ~n78 ;
  assign n162 = ~\1(0)_pad  & \45(5)_pad  ;
  assign n197 = ~\41(4)_pad  & n162 ;
  assign n198 = n83 & n197 ;
  assign n85 = ~\1698(48)_pad  & ~\33(3)_pad  ;
  assign n200 = \257(34)_pad  & n85 ;
  assign n87 = \1698(48)_pad  & ~\33(3)_pad  ;
  assign n199 = \264(35)_pad  & n87 ;
  assign n201 = \303(40)_pad  & \33(3)_pad  ;
  assign n202 = ~n199 & ~n201 ;
  assign n203 = ~n200 & n202 ;
  assign n204 = n78 & ~n203 ;
  assign n205 = ~n78 & ~n197 ;
  assign n206 = \270(36)_pad  & n205 ;
  assign n207 = ~n204 & ~n206 ;
  assign n208 = ~n198 & n207 ;
  assign n209 = \169(22)_pad  & ~n208 ;
  assign n210 = \179(23)_pad  & n208 ;
  assign n211 = ~n209 & ~n210 ;
  assign n212 = ~n196 & ~n211 ;
  assign n331 = \190(24)_pad  & n208 ;
  assign n330 = \200(25)_pad  & ~n208 ;
  assign n332 = n196 & ~n330 ;
  assign n333 = ~n331 & n332 ;
  assign n334 = ~n212 & ~n333 ;
  assign n157 = \244(32)_pad  & n87 ;
  assign n156 = \238(31)_pad  & n85 ;
  assign n158 = \116(13)_pad  & \33(3)_pad  ;
  assign n159 = ~n156 & ~n158 ;
  assign n160 = ~n157 & n159 ;
  assign n161 = n78 & ~n160 ;
  assign n164 = ~\274(37)_pad  & n162 ;
  assign n163 = ~\250(33)_pad  & ~n162 ;
  assign n165 = ~n78 & ~n163 ;
  assign n166 = ~n164 & n165 ;
  assign n167 = ~n161 & ~n166 ;
  assign n168 = \179(23)_pad  & n167 ;
  assign n169 = \169(22)_pad  & ~n167 ;
  assign n170 = ~n168 & ~n169 ;
  assign n176 = ~\107(12)_pad  & ~\87(10)_pad  ;
  assign n177 = ~\97(11)_pad  & n176 ;
  assign n178 = \20(2)_pad  & ~n177 ;
  assign n115 = \33(3)_pad  & \97(11)_pad  ;
  assign n64 = ~\20(2)_pad  & ~\33(3)_pad  ;
  assign n179 = \68(8)_pad  & n64 ;
  assign n180 = ~n115 & ~n179 ;
  assign n181 = ~n178 & n180 ;
  assign n182 = ~n57 & ~n181 ;
  assign n171 = ~\87(10)_pad  & n70 ;
  assign n175 = \87(10)_pad  & n174 ;
  assign n183 = ~n171 & ~n175 ;
  assign n184 = ~n182 & n183 ;
  assign n185 = ~n170 & ~n184 ;
  assign n272 = \200(25)_pad  & ~n167 ;
  assign n271 = \190(24)_pad  & n167 ;
  assign n273 = n184 & ~n271 ;
  assign n274 = ~n272 & n273 ;
  assign n335 = ~n185 & ~n274 ;
  assign n223 = \250(33)_pad  & n85 ;
  assign n222 = \257(34)_pad  & n87 ;
  assign n224 = \294(39)_pad  & \33(3)_pad  ;
  assign n225 = ~n222 & ~n224 ;
  assign n226 = ~n223 & n225 ;
  assign n227 = n78 & ~n226 ;
  assign n221 = \264(35)_pad  & n205 ;
  assign n228 = ~n198 & ~n221 ;
  assign n229 = ~n227 & n228 ;
  assign n236 = \200(25)_pad  & ~n229 ;
  assign n214 = \107(12)_pad  & n174 ;
  assign n101 = ~\13(1)_pad  & ~\33(3)_pad  ;
  assign n102 = n55 & ~n101 ;
  assign n103 = ~n70 & ~n102 ;
  assign n213 = ~\107(12)_pad  & ~n103 ;
  assign n215 = ~\33(3)_pad  & \87(10)_pad  ;
  assign n216 = ~n158 & ~n215 ;
  assign n217 = ~\20(2)_pad  & ~n216 ;
  assign n218 = ~n57 & n217 ;
  assign n219 = ~n213 & ~n218 ;
  assign n220 = ~n214 & n219 ;
  assign n235 = \190(24)_pad  & n229 ;
  assign n237 = n220 & ~n235 ;
  assign n238 = ~n236 & n237 ;
  assign n241 = \250(33)_pad  & n87 ;
  assign n240 = \244(32)_pad  & n85 ;
  assign n242 = ~n189 & ~n240 ;
  assign n243 = ~n241 & n242 ;
  assign n244 = n78 & ~n243 ;
  assign n239 = \257(34)_pad  & n205 ;
  assign n245 = ~n198 & ~n239 ;
  assign n246 = ~n244 & n245 ;
  assign n261 = \200(25)_pad  & ~n246 ;
  assign n247 = \190(24)_pad  & n246 ;
  assign n253 = ~\107(12)_pad  & ~\97(11)_pad  ;
  assign n254 = \107(12)_pad  & \97(11)_pad  ;
  assign n255 = ~n253 & ~n254 ;
  assign n256 = \20(2)_pad  & n255 ;
  assign n250 = ~\33(3)_pad  & \77(9)_pad  ;
  assign n145 = \107(12)_pad  & \33(3)_pad  ;
  assign n251 = ~\20(2)_pad  & ~n145 ;
  assign n252 = ~n250 & n251 ;
  assign n257 = ~n57 & ~n252 ;
  assign n258 = ~n256 & n257 ;
  assign n248 = ~\97(11)_pad  & n70 ;
  assign n249 = \97(11)_pad  & n174 ;
  assign n259 = ~n248 & ~n249 ;
  assign n260 = ~n258 & n259 ;
  assign n262 = ~n247 & n260 ;
  assign n263 = ~n261 & n262 ;
  assign n264 = ~n238 & ~n263 ;
  assign n231 = ~\179(23)_pad  & n229 ;
  assign n230 = ~\169(22)_pad  & ~n229 ;
  assign n232 = ~n220 & ~n230 ;
  assign n233 = ~n231 & n232 ;
  assign n267 = ~\179(23)_pad  & n246 ;
  assign n266 = ~\169(22)_pad  & ~n246 ;
  assign n268 = ~n260 & ~n266 ;
  assign n269 = ~n267 & n268 ;
  assign n336 = ~n233 & ~n269 ;
  assign n337 = n264 & n336 ;
  assign n338 = n335 & n337 ;
  assign n339 = n334 & n338 ;
  assign n340 = ~n100 & ~n339 ;
  assign n344 = ~\179(23)_pad  & ~n167 ;
  assign n345 = ~n229 & ~n246 ;
  assign n346 = n344 & n345 ;
  assign n347 = ~n208 & n346 ;
  assign n341 = n207 & n229 ;
  assign n342 = n246 & n341 ;
  assign n343 = n168 & n342 ;
  assign n348 = n100 & ~n343 ;
  assign n349 = ~n347 & n348 ;
  assign n350 = \330(46)_pad  & ~n349 ;
  assign n351 = ~n340 & n350 ;
  assign n234 = ~n212 & ~n233 ;
  assign n265 = ~n234 & n264 ;
  assign n270 = ~n265 & ~n269 ;
  assign n275 = ~n270 & ~n274 ;
  assign n276 = ~n185 & ~n275 ;
  assign n433 = ~n100 & ~n276 ;
  assign n434 = ~n351 & ~n433 ;
  assign n116 = \232(30)_pad  & n87 ;
  assign n114 = \226(29)_pad  & n85 ;
  assign n117 = ~n114 & ~n115 ;
  assign n118 = ~n116 & n117 ;
  assign n119 = n78 & ~n118 ;
  assign n79 = ~\41(4)_pad  & ~\45(5)_pad  ;
  assign n80 = ~\1(0)_pad  & ~n79 ;
  assign n84 = n80 & n83 ;
  assign n81 = ~n78 & ~n80 ;
  assign n113 = \238(31)_pad  & n81 ;
  assign n120 = ~n84 & ~n113 ;
  assign n121 = ~n119 & n120 ;
  assign n123 = ~\179(23)_pad  & n121 ;
  assign n72 = ~\1(0)_pad  & \20(2)_pad  ;
  assign n73 = n57 & ~n72 ;
  assign n105 = \68(8)_pad  & n73 ;
  assign n104 = ~\68(8)_pad  & ~n103 ;
  assign n106 = \33(3)_pad  & \77(9)_pad  ;
  assign n107 = ~\33(3)_pad  & \50(6)_pad  ;
  assign n108 = ~n106 & ~n107 ;
  assign n109 = ~\20(2)_pad  & ~n108 ;
  assign n110 = ~n57 & n109 ;
  assign n111 = ~n104 & ~n110 ;
  assign n112 = ~n105 & n111 ;
  assign n122 = ~\169(22)_pad  & ~n121 ;
  assign n124 = ~n112 & ~n122 ;
  assign n125 = ~n123 & n124 ;
  assign n127 = \200(25)_pad  & ~n121 ;
  assign n126 = \190(24)_pad  & n121 ;
  assign n128 = n112 & ~n126 ;
  assign n129 = ~n127 & n128 ;
  assign n130 = ~n125 & ~n129 ;
  assign n88 = \226(29)_pad  & n87 ;
  assign n86 = \223(28)_pad  & n85 ;
  assign n89 = \33(3)_pad  & \87(10)_pad  ;
  assign n90 = ~n86 & ~n89 ;
  assign n91 = ~n88 & n90 ;
  assign n92 = n78 & ~n91 ;
  assign n82 = \232(30)_pad  & n81 ;
  assign n93 = ~n82 & ~n84 ;
  assign n94 = ~n92 & n93 ;
  assign n96 = ~\179(23)_pad  & n94 ;
  assign n74 = \58(7)_pad  & n73 ;
  assign n60 = ~\58(7)_pad  & ~\68(8)_pad  ;
  assign n61 = \58(7)_pad  & \68(8)_pad  ;
  assign n62 = ~n60 & ~n61 ;
  assign n63 = \20(2)_pad  & ~n62 ;
  assign n58 = ~\20(2)_pad  & \33(3)_pad  ;
  assign n59 = \68(8)_pad  & n58 ;
  assign n65 = \159(21)_pad  & n64 ;
  assign n66 = ~n59 & ~n65 ;
  assign n67 = ~n63 & n66 ;
  assign n68 = ~n57 & ~n67 ;
  assign n71 = ~\58(7)_pad  & n70 ;
  assign n75 = ~n68 & ~n71 ;
  assign n76 = ~n74 & n75 ;
  assign n95 = ~\169(22)_pad  & ~n94 ;
  assign n97 = ~n76 & ~n95 ;
  assign n98 = ~n96 & n97 ;
  assign n291 = \200(25)_pad  & ~n94 ;
  assign n290 = \190(24)_pad  & n94 ;
  assign n292 = n76 & ~n290 ;
  assign n293 = ~n291 & n292 ;
  assign n435 = ~n98 & ~n293 ;
  assign n436 = n130 & n435 ;
  assign n146 = \238(31)_pad  & n87 ;
  assign n144 = \232(30)_pad  & n85 ;
  assign n147 = ~n144 & ~n145 ;
  assign n148 = ~n146 & n147 ;
  assign n149 = n78 & ~n148 ;
  assign n143 = \244(32)_pad  & n81 ;
  assign n150 = ~n84 & ~n143 ;
  assign n151 = ~n149 & n150 ;
  assign n153 = ~\179(23)_pad  & n151 ;
  assign n136 = ~\33(3)_pad  & \58(7)_pad  ;
  assign n137 = ~\20(2)_pad  & ~n89 ;
  assign n138 = ~n136 & n137 ;
  assign n135 = \20(2)_pad  & ~\77(9)_pad  ;
  assign n139 = ~n57 & ~n135 ;
  assign n140 = ~n138 & n139 ;
  assign n133 = ~\77(9)_pad  & n70 ;
  assign n134 = \77(9)_pad  & n73 ;
  assign n141 = ~n133 & ~n134 ;
  assign n142 = ~n140 & n141 ;
  assign n152 = ~\169(22)_pad  & ~n151 ;
  assign n154 = ~n142 & ~n152 ;
  assign n155 = ~n153 & n154 ;
  assign n279 = \190(24)_pad  & n151 ;
  assign n278 = \200(25)_pad  & ~n151 ;
  assign n280 = n142 & ~n278 ;
  assign n281 = ~n279 & n280 ;
  assign n282 = ~n155 & ~n281 ;
  assign n311 = \223(28)_pad  & n87 ;
  assign n310 = \222(27)_pad  & n85 ;
  assign n312 = ~n106 & ~n310 ;
  assign n313 = ~n311 & n312 ;
  assign n314 = n78 & ~n313 ;
  assign n309 = \226(29)_pad  & n81 ;
  assign n315 = ~n84 & ~n309 ;
  assign n316 = ~n314 & n315 ;
  assign n318 = ~\179(23)_pad  & n316 ;
  assign n306 = \50(6)_pad  & n73 ;
  assign n299 = ~\50(6)_pad  & n60 ;
  assign n300 = \20(2)_pad  & ~n299 ;
  assign n298 = \58(7)_pad  & n58 ;
  assign n301 = \150(20)_pad  & n64 ;
  assign n302 = ~n298 & ~n301 ;
  assign n303 = ~n300 & n302 ;
  assign n304 = ~n57 & ~n303 ;
  assign n305 = ~\50(6)_pad  & n70 ;
  assign n307 = ~n304 & ~n305 ;
  assign n308 = ~n306 & n307 ;
  assign n317 = ~\169(22)_pad  & ~n316 ;
  assign n319 = ~n308 & ~n317 ;
  assign n320 = ~n318 & n319 ;
  assign n322 = \200(25)_pad  & ~n316 ;
  assign n321 = \190(24)_pad  & n316 ;
  assign n323 = n308 & ~n321 ;
  assign n324 = ~n322 & n323 ;
  assign n325 = ~n320 & ~n324 ;
  assign n437 = n282 & n325 ;
  assign n438 = n436 & n437 ;
  assign n439 = ~n434 & n438 ;
  assign n440 = ~n129 & n155 ;
  assign n441 = ~n125 & ~n440 ;
  assign n442 = ~n293 & ~n441 ;
  assign n443 = ~n98 & ~n442 ;
  assign n444 = ~n324 & ~n443 ;
  assign n445 = ~n320 & ~n444 ;
  assign n446 = ~n439 & n445 ;
  assign n131 = n100 & ~n112 ;
  assign n132 = n130 & ~n131 ;
  assign n355 = n100 & n125 ;
  assign n356 = ~n132 & ~n355 ;
  assign n277 = n100 & ~n142 ;
  assign n283 = ~n277 & n282 ;
  assign n353 = n100 & n155 ;
  assign n354 = ~n283 & ~n353 ;
  assign n447 = n351 & ~n354 ;
  assign n448 = n356 & ~n447 ;
  assign n357 = ~n354 & ~n356 ;
  assign n449 = n351 & n357 ;
  assign n450 = ~n448 & ~n449 ;
  assign n284 = ~n276 & n283 ;
  assign n285 = ~n155 & ~n284 ;
  assign n451 = ~n100 & ~n285 ;
  assign n452 = ~n450 & n451 ;
  assign n453 = n450 & ~n451 ;
  assign n454 = ~n452 & ~n453 ;
  assign n455 = n446 & ~n454 ;
  assign n286 = n132 & ~n285 ;
  assign n287 = ~n125 & ~n286 ;
  assign n288 = ~n100 & ~n287 ;
  assign n99 = ~n53 & n98 ;
  assign n289 = n53 & ~n76 ;
  assign n294 = ~n289 & ~n293 ;
  assign n295 = ~n98 & ~n294 ;
  assign n352 = ~n99 & ~n295 ;
  assign n358 = n352 & n357 ;
  assign n359 = n351 & n358 ;
  assign n456 = ~n352 & ~n449 ;
  assign n457 = ~n359 & ~n456 ;
  assign n458 = ~n288 & n457 ;
  assign n459 = n288 & ~n457 ;
  assign n460 = ~n458 & ~n459 ;
  assign n461 = n455 & ~n460 ;
  assign n462 = n446 & ~n461 ;
  assign n296 = n288 & ~n295 ;
  assign n297 = ~n99 & ~n296 ;
  assign n326 = n53 & ~n308 ;
  assign n327 = n325 & ~n326 ;
  assign n328 = n53 & n320 ;
  assign n329 = ~n327 & ~n328 ;
  assign n360 = ~n329 & n359 ;
  assign n361 = n329 & ~n359 ;
  assign n362 = ~n360 & ~n361 ;
  assign n363 = n297 & n362 ;
  assign n364 = ~n297 & ~n362 ;
  assign n365 = ~n363 & ~n364 ;
  assign n369 = ~\13(1)_pad  & n55 ;
  assign n370 = ~\41(4)_pad  & n369 ;
  assign n463 = ~n365 & n370 ;
  assign n464 = ~n462 & n463 ;
  assign n366 = \45(5)_pad  & n51 ;
  assign n367 = \1(0)_pad  & ~n366 ;
  assign n368 = ~n365 & ~n367 ;
  assign n427 = n101 & n329 ;
  assign n372 = ~\169(22)_pad  & \20(2)_pad  ;
  assign n373 = n54 & ~n372 ;
  assign n375 = \179(23)_pad  & \20(2)_pad  ;
  assign n384 = ~\200(25)_pad  & n375 ;
  assign n389 = ~\190(24)_pad  & n384 ;
  assign n414 = \87(10)_pad  & n389 ;
  assign n376 = \200(25)_pad  & n375 ;
  assign n377 = \190(24)_pad  & n376 ;
  assign n412 = \116(13)_pad  & n377 ;
  assign n379 = \20(2)_pad  & \200(25)_pad  ;
  assign n380 = ~n375 & ~n379 ;
  assign n381 = ~\190(24)_pad  & \20(2)_pad  ;
  assign n382 = n380 & ~n381 ;
  assign n413 = \68(8)_pad  & n382 ;
  assign n419 = ~n412 & ~n413 ;
  assign n420 = ~n414 & n419 ;
  assign n393 = ~n375 & n379 ;
  assign n396 = ~\190(24)_pad  & n393 ;
  assign n407 = \58(7)_pad  & n396 ;
  assign n415 = \33(3)_pad  & ~\41(4)_pad  ;
  assign n416 = ~n407 & n415 ;
  assign n387 = n380 & n381 ;
  assign n408 = \283(38)_pad  & n387 ;
  assign n394 = \190(24)_pad  & n393 ;
  assign n409 = \77(9)_pad  & n394 ;
  assign n417 = ~n408 & ~n409 ;
  assign n391 = ~\190(24)_pad  & n376 ;
  assign n410 = \97(11)_pad  & n391 ;
  assign n385 = \190(24)_pad  & n384 ;
  assign n411 = \107(12)_pad  & n385 ;
  assign n418 = ~n410 & ~n411 ;
  assign n421 = n417 & n418 ;
  assign n422 = n416 & n421 ;
  assign n423 = n420 & n422 ;
  assign n374 = \41(4)_pad  & ~\50(6)_pad  ;
  assign n397 = \159(21)_pad  & n396 ;
  assign n392 = \132(17)_pad  & n391 ;
  assign n395 = \143(19)_pad  & n394 ;
  assign n402 = ~n392 & ~n395 ;
  assign n403 = ~n397 & n402 ;
  assign n378 = \125(15)_pad  & n377 ;
  assign n398 = ~\33(3)_pad  & ~\41(4)_pad  ;
  assign n399 = ~n378 & n398 ;
  assign n383 = \150(20)_pad  & n382 ;
  assign n386 = \128(16)_pad  & n385 ;
  assign n400 = ~n383 & ~n386 ;
  assign n388 = \124(14)_pad  & n387 ;
  assign n390 = \137(18)_pad  & n389 ;
  assign n401 = ~n388 & ~n390 ;
  assign n404 = n400 & n401 ;
  assign n405 = n399 & n404 ;
  assign n406 = n403 & n405 ;
  assign n424 = ~n374 & ~n406 ;
  assign n425 = ~n423 & n424 ;
  assign n426 = n373 & ~n425 ;
  assign n371 = n367 & ~n370 ;
  assign n428 = ~n101 & ~n373 ;
  assign n429 = ~\50(6)_pad  & n428 ;
  assign n430 = n371 & ~n429 ;
  assign n431 = ~n426 & n430 ;
  assign n432 = ~n427 & n431 ;
  assign n465 = ~n368 & ~n432 ;
  assign n466 = ~n464 & n465 ;
  assign n507 = ~n455 & n460 ;
  assign n508 = n370 & ~n461 ;
  assign n509 = ~n507 & n508 ;
  assign n467 = ~n367 & ~n460 ;
  assign n502 = n101 & ~n352 ;
  assign n475 = \159(21)_pad  & n382 ;
  assign n473 = \150(20)_pad  & n394 ;
  assign n474 = \128(16)_pad  & n377 ;
  assign n479 = ~n473 & ~n474 ;
  assign n480 = ~n475 & n479 ;
  assign n468 = \137(18)_pad  & n391 ;
  assign n476 = ~\33(3)_pad  & ~n468 ;
  assign n469 = \50(6)_pad  & n396 ;
  assign n470 = \132(17)_pad  & n385 ;
  assign n477 = ~n469 & ~n470 ;
  assign n471 = \143(19)_pad  & n389 ;
  assign n472 = \125(15)_pad  & n387 ;
  assign n478 = ~n471 & ~n472 ;
  assign n481 = n477 & n478 ;
  assign n482 = n476 & n481 ;
  assign n483 = n480 & n482 ;
  assign n491 = \283(38)_pad  & n377 ;
  assign n489 = \77(9)_pad  & n382 ;
  assign n490 = \107(12)_pad  & n391 ;
  assign n495 = ~n489 & ~n490 ;
  assign n496 = ~n491 & n495 ;
  assign n484 = \68(8)_pad  & n396 ;
  assign n492 = \33(3)_pad  & ~n484 ;
  assign n485 = \87(10)_pad  & n394 ;
  assign n486 = \294(39)_pad  & n387 ;
  assign n493 = ~n485 & ~n486 ;
  assign n487 = \97(11)_pad  & n389 ;
  assign n488 = \116(13)_pad  & n385 ;
  assign n494 = ~n487 & ~n488 ;
  assign n497 = n493 & n494 ;
  assign n498 = n492 & n497 ;
  assign n499 = n496 & n498 ;
  assign n500 = ~n483 & ~n499 ;
  assign n501 = n373 & ~n500 ;
  assign n503 = ~\58(7)_pad  & n428 ;
  assign n504 = n371 & ~n503 ;
  assign n505 = ~n501 & n504 ;
  assign n506 = ~n502 & n505 ;
  assign n510 = ~n467 & ~n506 ;
  assign n511 = ~n509 & n510 ;
  assign n512 = ~\50(6)_pad  & ~\77(9)_pad  ;
  assign n513 = n60 & n512 ;
  assign n514 = \87(10)_pad  & ~n253 ;
  assign n515 = ~\257(34)_pad  & ~\264(35)_pad  ;
  assign n516 = \257(34)_pad  & \264(35)_pad  ;
  assign n517 = ~n515 & ~n516 ;
  assign n518 = \250(33)_pad  & ~\270(36)_pad  ;
  assign n519 = ~\250(33)_pad  & \270(36)_pad  ;
  assign n520 = ~n518 & ~n519 ;
  assign n521 = n517 & n520 ;
  assign n522 = ~n517 & ~n520 ;
  assign n523 = ~n521 & ~n522 ;
  assign n524 = \226(29)_pad  & ~\232(30)_pad  ;
  assign n525 = ~\226(29)_pad  & \232(30)_pad  ;
  assign n526 = ~n524 & ~n525 ;
  assign n527 = \238(31)_pad  & ~\244(32)_pad  ;
  assign n528 = ~\238(31)_pad  & \244(32)_pad  ;
  assign n529 = ~n527 & ~n528 ;
  assign n530 = n526 & n529 ;
  assign n531 = ~n526 & ~n529 ;
  assign n532 = ~n530 & ~n531 ;
  assign n533 = n523 & n532 ;
  assign n534 = ~n523 & ~n532 ;
  assign n535 = ~n533 & ~n534 ;
  assign n540 = \116(13)_pad  & \270(36)_pad  ;
  assign n541 = \107(12)_pad  & \264(35)_pad  ;
  assign n546 = ~n540 & ~n541 ;
  assign n542 = \238(31)_pad  & \68(8)_pad  ;
  assign n543 = \257(34)_pad  & \97(11)_pad  ;
  assign n547 = ~n542 & ~n543 ;
  assign n548 = n546 & n547 ;
  assign n536 = \232(30)_pad  & \58(7)_pad  ;
  assign n537 = \226(29)_pad  & \50(6)_pad  ;
  assign n544 = ~n536 & ~n537 ;
  assign n538 = \250(33)_pad  & \87(10)_pad  ;
  assign n539 = \244(32)_pad  & \77(9)_pad  ;
  assign n545 = ~n538 & ~n539 ;
  assign n549 = n544 & n545 ;
  assign n550 = n548 & n549 ;
  assign n551 = ~n55 & ~n550 ;
  assign n552 = \50(6)_pad  & ~n60 ;
  assign n553 = \1(0)_pad  & n69 ;
  assign n554 = n552 & n553 ;
  assign n555 = \250(33)_pad  & ~n515 ;
  assign n556 = n369 & n555 ;
  assign n557 = ~n554 & ~n556 ;
  assign n558 = ~n551 & n557 ;
  assign n560 = ~\1(0)_pad  & ~n434 ;
  assign n559 = n370 & n552 ;
  assign n561 = ~\116(13)_pad  & n177 ;
  assign n562 = \1(0)_pad  & ~n370 ;
  assign n563 = n561 & n562 ;
  assign n564 = ~n559 & ~n563 ;
  assign n565 = ~n560 & n564 ;
  assign n566 = ~\50(6)_pad  & \68(8)_pad  ;
  assign n567 = \50(6)_pad  & \77(9)_pad  ;
  assign n568 = n62 & n567 ;
  assign n569 = ~n566 & ~n568 ;
  assign n570 = ~\13(1)_pad  & ~n569 ;
  assign n571 = \116(13)_pad  & n255 ;
  assign n572 = n69 & n571 ;
  assign n573 = ~n570 & ~n572 ;
  assign n574 = \1(0)_pad  & ~n573 ;
  assign n577 = n358 & n438 ;
  assign n576 = ~n358 & ~n438 ;
  assign n578 = n351 & ~n576 ;
  assign n579 = ~n577 & n578 ;
  assign n580 = ~n297 & n579 ;
  assign n581 = n297 & ~n579 ;
  assign n582 = ~n580 & ~n581 ;
  assign n583 = n433 & n438 ;
  assign n584 = n445 & ~n583 ;
  assign n586 = ~n582 & n584 ;
  assign n575 = \1(0)_pad  & ~n51 ;
  assign n585 = n582 & ~n584 ;
  assign n587 = ~n575 & ~n585 ;
  assign n588 = ~n586 & n587 ;
  assign n589 = ~n574 & ~n588 ;
  assign n590 = ~n276 & n438 ;
  assign n591 = n445 & ~n590 ;
  assign n592 = n339 & n438 ;
  assign n632 = ~n446 & n454 ;
  assign n633 = n370 & ~n455 ;
  assign n634 = ~n632 & n633 ;
  assign n593 = ~n367 & ~n454 ;
  assign n627 = n101 & n356 ;
  assign n601 = \303(40)_pad  & n387 ;
  assign n599 = \116(13)_pad  & n391 ;
  assign n600 = \283(38)_pad  & n385 ;
  assign n605 = ~n599 & ~n600 ;
  assign n606 = ~n601 & n605 ;
  assign n594 = \87(10)_pad  & n382 ;
  assign n602 = \33(3)_pad  & ~n594 ;
  assign n595 = \97(11)_pad  & n394 ;
  assign n596 = \77(9)_pad  & n396 ;
  assign n603 = ~n595 & ~n596 ;
  assign n597 = \294(39)_pad  & n377 ;
  assign n598 = \107(12)_pad  & n389 ;
  assign n604 = ~n597 & ~n598 ;
  assign n607 = n603 & n604 ;
  assign n608 = n602 & n607 ;
  assign n609 = n606 & n608 ;
  assign n616 = \150(20)_pad  & n389 ;
  assign n614 = \50(6)_pad  & n382 ;
  assign n615 = \143(19)_pad  & n391 ;
  assign n620 = ~n614 & ~n615 ;
  assign n621 = ~n616 & n620 ;
  assign n617 = ~\33(3)_pad  & ~n407 ;
  assign n610 = \132(17)_pad  & n377 ;
  assign n611 = \159(21)_pad  & n394 ;
  assign n618 = ~n610 & ~n611 ;
  assign n612 = \137(18)_pad  & n385 ;
  assign n613 = \128(16)_pad  & n387 ;
  assign n619 = ~n612 & ~n613 ;
  assign n622 = n618 & n619 ;
  assign n623 = n617 & n622 ;
  assign n624 = n621 & n623 ;
  assign n625 = ~n609 & ~n624 ;
  assign n626 = n373 & ~n625 ;
  assign n628 = ~\68(8)_pad  & n428 ;
  assign n629 = n371 & ~n628 ;
  assign n630 = ~n626 & n629 ;
  assign n631 = ~n627 & n630 ;
  assign n635 = ~n593 & ~n631 ;
  assign n636 = ~n634 & n635 ;
  assign n637 = ~n351 & n354 ;
  assign n638 = ~n447 & ~n637 ;
  assign n640 = ~n433 & ~n638 ;
  assign n639 = n433 & n638 ;
  assign n641 = ~n371 & ~n639 ;
  assign n642 = ~n640 & n641 ;
  assign n676 = n101 & n354 ;
  assign n650 = \311(41)_pad  & n387 ;
  assign n648 = \283(38)_pad  & n391 ;
  assign n649 = \294(39)_pad  & n385 ;
  assign n654 = ~n648 & ~n649 ;
  assign n655 = ~n650 & n654 ;
  assign n643 = \97(11)_pad  & n382 ;
  assign n651 = \33(3)_pad  & ~n643 ;
  assign n644 = \107(12)_pad  & n394 ;
  assign n645 = \87(10)_pad  & n396 ;
  assign n652 = ~n644 & ~n645 ;
  assign n646 = \303(40)_pad  & n377 ;
  assign n647 = \116(13)_pad  & n389 ;
  assign n653 = ~n646 & ~n647 ;
  assign n656 = n652 & n653 ;
  assign n657 = n651 & n656 ;
  assign n658 = n655 & n657 ;
  assign n665 = \159(21)_pad  & n389 ;
  assign n663 = \58(7)_pad  & n382 ;
  assign n664 = \150(20)_pad  & n391 ;
  assign n669 = ~n663 & ~n664 ;
  assign n670 = ~n665 & n669 ;
  assign n666 = ~\33(3)_pad  & ~n484 ;
  assign n659 = \137(18)_pad  & n377 ;
  assign n660 = \50(6)_pad  & n394 ;
  assign n667 = ~n659 & ~n660 ;
  assign n661 = \143(19)_pad  & n385 ;
  assign n662 = \132(17)_pad  & n387 ;
  assign n668 = ~n661 & ~n662 ;
  assign n671 = n667 & n668 ;
  assign n672 = n666 & n671 ;
  assign n673 = n670 & n672 ;
  assign n674 = ~n658 & ~n673 ;
  assign n675 = n373 & ~n674 ;
  assign n677 = ~\77(9)_pad  & n428 ;
  assign n678 = n371 & ~n677 ;
  assign n679 = ~n675 & n678 ;
  assign n680 = ~n676 & n679 ;
  assign n681 = ~n642 & ~n680 ;
  assign n682 = ~\13(1)_pad  & n64 ;
  assign n683 = n100 & ~n184 ;
  assign n684 = n335 & ~n683 ;
  assign n685 = n100 & n185 ;
  assign n686 = ~n684 & ~n685 ;
  assign n687 = n682 & n686 ;
  assign n693 = \50(6)_pad  & n389 ;
  assign n691 = \58(7)_pad  & n394 ;
  assign n692 = \150(20)_pad  & n385 ;
  assign n697 = ~n691 & ~n692 ;
  assign n698 = ~n693 & n697 ;
  assign n694 = ~\33(3)_pad  & ~n413 ;
  assign n688 = \159(21)_pad  & n391 ;
  assign n695 = ~n596 & ~n688 ;
  assign n689 = \137(18)_pad  & n387 ;
  assign n690 = \143(19)_pad  & n377 ;
  assign n696 = ~n689 & ~n690 ;
  assign n699 = n695 & n696 ;
  assign n700 = n694 & n699 ;
  assign n701 = n698 & n700 ;
  assign n709 = \107(12)_pad  & n382 ;
  assign n707 = \116(13)_pad  & n394 ;
  assign n708 = \283(38)_pad  & n389 ;
  assign n713 = ~n707 & ~n708 ;
  assign n714 = ~n709 & n713 ;
  assign n702 = \294(39)_pad  & n391 ;
  assign n710 = \33(3)_pad  & ~n702 ;
  assign n703 = \97(11)_pad  & n396 ;
  assign n704 = \311(41)_pad  & n377 ;
  assign n711 = ~n703 & ~n704 ;
  assign n705 = \303(40)_pad  & n385 ;
  assign n706 = \317(42)_pad  & n387 ;
  assign n712 = ~n705 & ~n706 ;
  assign n715 = n711 & n712 ;
  assign n716 = n710 & n715 ;
  assign n717 = n714 & n716 ;
  assign n718 = ~n701 & ~n717 ;
  assign n719 = n373 & ~n718 ;
  assign n721 = ~\13(1)_pad  & n56 ;
  assign n722 = n523 & n721 ;
  assign n720 = ~n373 & ~n682 ;
  assign n723 = \87(10)_pad  & ~n369 ;
  assign n724 = n720 & ~n723 ;
  assign n725 = ~n722 & n724 ;
  assign n726 = n371 & ~n725 ;
  assign n727 = ~n719 & n726 ;
  assign n728 = ~n687 & n727 ;
  assign n729 = n100 & ~n196 ;
  assign n730 = n334 & ~n729 ;
  assign n731 = ~n211 & n729 ;
  assign n732 = ~n730 & ~n731 ;
  assign n733 = \330(46)_pad  & ~n732 ;
  assign n734 = ~n100 & n212 ;
  assign n735 = ~n100 & n233 ;
  assign n736 = n100 & ~n220 ;
  assign n737 = ~n238 & ~n736 ;
  assign n738 = ~n233 & ~n737 ;
  assign n739 = ~n735 & ~n738 ;
  assign n740 = ~n734 & ~n739 ;
  assign n741 = ~n233 & ~n238 ;
  assign n742 = n734 & n741 ;
  assign n743 = ~n740 & ~n742 ;
  assign n744 = ~n733 & n743 ;
  assign n745 = n733 & ~n743 ;
  assign n746 = ~n744 & ~n745 ;
  assign n747 = n434 & ~n746 ;
  assign n748 = ~n100 & n269 ;
  assign n749 = n100 & ~n260 ;
  assign n750 = ~n263 & ~n749 ;
  assign n751 = ~n269 & ~n750 ;
  assign n752 = ~n748 & ~n751 ;
  assign n753 = n733 & ~n738 ;
  assign n754 = ~n735 & ~n753 ;
  assign n755 = ~n742 & n754 ;
  assign n756 = n742 & ~n754 ;
  assign n757 = ~n755 & ~n756 ;
  assign n758 = n752 & ~n757 ;
  assign n759 = ~n752 & n757 ;
  assign n760 = ~n758 & ~n759 ;
  assign n761 = n747 & ~n760 ;
  assign n762 = n434 & ~n761 ;
  assign n763 = n370 & ~n762 ;
  assign n764 = n367 & ~n763 ;
  assign n765 = ~n751 & n757 ;
  assign n766 = ~n748 & ~n765 ;
  assign n767 = ~n686 & ~n766 ;
  assign n768 = n686 & n766 ;
  assign n769 = ~n767 & ~n768 ;
  assign n770 = ~n764 & n769 ;
  assign n771 = ~n728 & ~n770 ;
  assign n818 = ~n747 & n760 ;
  assign n819 = n370 & ~n761 ;
  assign n820 = ~n818 & n819 ;
  assign n772 = ~n367 & ~n760 ;
  assign n814 = n682 & ~n752 ;
  assign n789 = \303(40)_pad  & n391 ;
  assign n787 = \317(42)_pad  & n377 ;
  assign n788 = \311(41)_pad  & n385 ;
  assign n793 = ~n787 & ~n788 ;
  assign n794 = ~n789 & n793 ;
  assign n782 = \116(13)_pad  & n382 ;
  assign n790 = \33(3)_pad  & ~n782 ;
  assign n783 = \294(39)_pad  & n389 ;
  assign n784 = \322(43)_pad  & n387 ;
  assign n791 = ~n783 & ~n784 ;
  assign n785 = \283(38)_pad  & n394 ;
  assign n786 = \107(12)_pad  & n396 ;
  assign n792 = ~n785 & ~n786 ;
  assign n795 = n791 & n792 ;
  assign n796 = n790 & n795 ;
  assign n797 = n794 & n796 ;
  assign n803 = \58(7)_pad  & n389 ;
  assign n801 = \68(8)_pad  & n394 ;
  assign n802 = \159(21)_pad  & n385 ;
  assign n807 = ~n801 & ~n802 ;
  assign n808 = ~n803 & n807 ;
  assign n804 = ~\33(3)_pad  & ~n489 ;
  assign n798 = \50(6)_pad  & n391 ;
  assign n805 = ~n645 & ~n798 ;
  assign n799 = \143(19)_pad  & n387 ;
  assign n800 = \150(20)_pad  & n377 ;
  assign n806 = ~n799 & ~n800 ;
  assign n809 = n805 & n806 ;
  assign n810 = n804 & n809 ;
  assign n811 = n808 & n810 ;
  assign n812 = ~n797 & ~n811 ;
  assign n813 = n373 & ~n812 ;
  assign n774 = ~\116(13)_pad  & ~n255 ;
  assign n775 = ~n571 & ~n774 ;
  assign n776 = \87(10)_pad  & n775 ;
  assign n777 = ~\87(10)_pad  & ~n775 ;
  assign n778 = ~n776 & ~n777 ;
  assign n779 = n721 & ~n778 ;
  assign n773 = \97(11)_pad  & ~n369 ;
  assign n780 = n720 & ~n773 ;
  assign n781 = ~n779 & n780 ;
  assign n815 = n371 & ~n781 ;
  assign n816 = ~n813 & n815 ;
  assign n817 = ~n814 & n816 ;
  assign n821 = ~n772 & ~n817 ;
  assign n822 = ~n820 & n821 ;
  assign n873 = ~n434 & n746 ;
  assign n874 = n370 & ~n747 ;
  assign n875 = ~n873 & n874 ;
  assign n823 = ~n367 & ~n746 ;
  assign n824 = n682 & ~n739 ;
  assign n843 = \159(21)_pad  & n377 ;
  assign n841 = \68(8)_pad  & n389 ;
  assign n842 = \58(7)_pad  & n391 ;
  assign n847 = ~n841 & ~n842 ;
  assign n848 = ~n843 & n847 ;
  assign n844 = ~\33(3)_pad  & ~n409 ;
  assign n845 = ~n594 & ~n703 ;
  assign n839 = \150(20)_pad  & n387 ;
  assign n840 = \50(6)_pad  & n385 ;
  assign n846 = ~n839 & ~n840 ;
  assign n849 = n845 & n846 ;
  assign n850 = n844 & n849 ;
  assign n851 = n848 & n850 ;
  assign n859 = \311(41)_pad  & n391 ;
  assign n857 = \294(39)_pad  & n394 ;
  assign n858 = \322(43)_pad  & n377 ;
  assign n863 = ~n857 & ~n858 ;
  assign n864 = ~n859 & n863 ;
  assign n852 = \303(40)_pad  & n389 ;
  assign n860 = \33(3)_pad  & ~n852 ;
  assign n853 = \116(13)_pad  & n396 ;
  assign n854 = \317(42)_pad  & n385 ;
  assign n861 = ~n853 & ~n854 ;
  assign n855 = \326(44)_pad  & n387 ;
  assign n856 = \283(38)_pad  & n382 ;
  assign n862 = ~n855 & ~n856 ;
  assign n865 = n861 & n862 ;
  assign n866 = n860 & n865 ;
  assign n867 = n864 & n866 ;
  assign n868 = ~n851 & ~n867 ;
  assign n869 = n373 & ~n868 ;
  assign n828 = \45(5)_pad  & ~n532 ;
  assign n829 = \68(8)_pad  & \77(9)_pad  ;
  assign n830 = ~\45(5)_pad  & ~\50(6)_pad  ;
  assign n831 = \58(7)_pad  & n830 ;
  assign n832 = ~n829 & n831 ;
  assign n833 = n561 & n832 ;
  assign n834 = n721 & ~n833 ;
  assign n835 = ~n828 & n834 ;
  assign n825 = ~\107(12)_pad  & ~n369 ;
  assign n826 = ~\33(3)_pad  & n369 ;
  assign n827 = ~n561 & n826 ;
  assign n836 = ~n825 & ~n827 ;
  assign n837 = ~n835 & n836 ;
  assign n838 = n720 & ~n837 ;
  assign n870 = n371 & ~n838 ;
  assign n871 = ~n869 & n870 ;
  assign n872 = ~n824 & n871 ;
  assign n876 = ~n823 & ~n872 ;
  assign n877 = ~n875 & n876 ;
  assign n878 = ~\330(46)_pad  & n732 ;
  assign n879 = ~n371 & ~n733 ;
  assign n880 = ~n878 & n879 ;
  assign n881 = n682 & n732 ;
  assign n889 = \283(38)_pad  & n396 ;
  assign n887 = \303(40)_pad  & n394 ;
  assign n888 = \326(44)_pad  & n377 ;
  assign n893 = ~n887 & ~n888 ;
  assign n894 = ~n889 & n893 ;
  assign n882 = \322(43)_pad  & n385 ;
  assign n890 = \33(3)_pad  & ~n882 ;
  assign n883 = \294(39)_pad  & n382 ;
  assign n884 = \329(45)_pad  & n387 ;
  assign n891 = ~n883 & ~n884 ;
  assign n885 = \317(42)_pad  & n391 ;
  assign n886 = \311(41)_pad  & n389 ;
  assign n892 = ~n885 & ~n886 ;
  assign n895 = n891 & n892 ;
  assign n896 = n890 & n895 ;
  assign n897 = n894 & n896 ;
  assign n902 = \50(6)_pad  & n377 ;
  assign n900 = \58(7)_pad  & n385 ;
  assign n901 = \77(9)_pad  & n389 ;
  assign n906 = ~n900 & ~n901 ;
  assign n907 = ~n902 & n906 ;
  assign n903 = ~\33(3)_pad  & ~n485 ;
  assign n904 = ~n643 & ~n786 ;
  assign n898 = \159(21)_pad  & n387 ;
  assign n899 = \68(8)_pad  & n391 ;
  assign n905 = ~n898 & ~n899 ;
  assign n908 = n904 & n905 ;
  assign n909 = n903 & n908 ;
  assign n910 = n907 & n909 ;
  assign n911 = ~n897 & ~n910 ;
  assign n912 = n373 & ~n911 ;
  assign n916 = ~n512 & ~n567 ;
  assign n917 = n62 & ~n916 ;
  assign n918 = ~n62 & n916 ;
  assign n919 = ~n917 & ~n918 ;
  assign n920 = \45(5)_pad  & n919 ;
  assign n915 = ~\45(5)_pad  & n552 ;
  assign n921 = n721 & ~n915 ;
  assign n922 = ~n920 & n921 ;
  assign n913 = ~\116(13)_pad  & ~n369 ;
  assign n914 = ~n514 & n826 ;
  assign n923 = ~n913 & ~n914 ;
  assign n924 = ~n922 & n923 ;
  assign n925 = n720 & ~n924 ;
  assign n926 = n371 & ~n925 ;
  assign n927 = ~n912 & n926 ;
  assign n928 = ~n881 & n927 ;
  assign n929 = ~n880 & ~n928 ;
  assign n930 = ~n466 & ~n511 ;
  assign n931 = n466 & n511 ;
  assign n932 = ~n930 & ~n931 ;
  assign n933 = n877 & ~n929 ;
  assign n934 = ~n877 & n929 ;
  assign n935 = ~n933 & ~n934 ;
  assign n936 = n771 & n935 ;
  assign n937 = ~n771 & ~n935 ;
  assign n938 = ~n936 & ~n937 ;
  assign n939 = ~n636 & n681 ;
  assign n940 = n636 & ~n681 ;
  assign n941 = ~n939 & ~n940 ;
  assign n942 = n822 & ~n941 ;
  assign n943 = ~n822 & n941 ;
  assign n944 = ~n942 & ~n943 ;
  assign n945 = n938 & n944 ;
  assign n946 = ~n938 & ~n944 ;
  assign n947 = ~n945 & ~n946 ;
  assign n948 = n932 & n947 ;
  assign n949 = ~n932 & ~n947 ;
  assign n950 = ~n948 & ~n949 ;
  assign n951 = \213(26)_pad  & ~\343(47)_pad  ;
  assign n952 = ~n932 & ~n951 ;
  assign n953 = ~\2897(49)_pad  & n951 ;
  assign n954 = ~n952 & ~n953 ;
  assign n955 = n947 & n954 ;
  assign n956 = ~n947 & ~n954 ;
  assign n957 = ~n955 & ~n956 ;
  assign n958 = n681 & n929 ;
  assign n959 = n877 & n958 ;
  assign n960 = n636 & n959 ;
  assign n961 = n822 & n960 ;
  assign n962 = n771 & n961 ;
  assign n963 = n931 & n962 ;
  assign n964 = n931 & n951 ;
  assign n965 = \213(26)_pad  & ~n963 ;
  assign n966 = ~n964 & n965 ;
  assign n967 = n778 & n919 ;
  assign n968 = ~n778 & ~n919 ;
  assign n969 = ~n967 & ~n968 ;
  assign \2690(1611)  = ~n466 ;
  assign \2709(1587)  = ~n511 ;
  assign \353(405)_pad  = n513 ;
  assign \355(399)_pad  = ~n514 ;
  assign \358(1161)_pad  = n535 ;
  assign \361(940)_pad  = n558 ;
  assign \364(1484)_pad  = ~n565 ;
  assign \367(1585)_pad  = ~n589 ;
  assign \369(1321)_pad  = ~n591 ;
  assign \372(1243)_pad  = n592 ;
  assign \381(1626)_pad  = ~n636 ;
  assign \384(1553)_pad  = ~n681 ;
  assign \387(1616)_pad  = ~n771 ;
  assign \390(1603)_pad  = ~n822 ;
  assign \393(1605)_pad  = ~n877 ;
  assign \396(1504)_pad  = ~n929 ;
  assign \399(1428)_pad  = ~n755 ;
  assign \402(1718)_pad  = n950 ;
  assign \404(1714)  = n957 ;
  assign \407(1657)_pad  = ~n963 ;
  assign \409(1670)_pad  = ~n966 ;
  assign \605(1186)  = n969 ;
endmodule
