module top( \dcnt_reg[0]/P0001  , \dcnt_reg[1]/P0001  , \dcnt_reg[2]/P0001  , \dcnt_reg[3]/P0001  , \key[0]_pad  , \key[100]_pad  , \key[101]_pad  , \key[102]_pad  , \key[103]_pad  , \key[104]_pad  , \key[105]_pad  , \key[106]_pad  , \key[107]_pad  , \key[108]_pad  , \key[109]_pad  , \key[10]_pad  , \key[110]_pad  , \key[111]_pad  , \key[112]_pad  , \key[113]_pad  , \key[114]_pad  , \key[115]_pad  , \key[116]_pad  , \key[117]_pad  , \key[118]_pad  , \key[119]_pad  , \key[11]_pad  , \key[120]_pad  , \key[121]_pad  , \key[122]_pad  , \key[123]_pad  , \key[124]_pad  , \key[125]_pad  , \key[126]_pad  , \key[127]_pad  , \key[12]_pad  , \key[13]_pad  , \key[14]_pad  , \key[15]_pad  , \key[16]_pad  , \key[17]_pad  , \key[18]_pad  , \key[19]_pad  , \key[1]_pad  , \key[20]_pad  , \key[21]_pad  , \key[22]_pad  , \key[23]_pad  , \key[24]_pad  , \key[25]_pad  , \key[26]_pad  , \key[27]_pad  , \key[28]_pad  , \key[29]_pad  , \key[2]_pad  , \key[30]_pad  , \key[31]_pad  , \key[32]_pad  , \key[33]_pad  , \key[34]_pad  , \key[35]_pad  , \key[36]_pad  , \key[37]_pad  , \key[38]_pad  , \key[39]_pad  , \key[3]_pad  , \key[40]_pad  , \key[41]_pad  , \key[42]_pad  , \key[43]_pad  , \key[44]_pad  , \key[45]_pad  , \key[46]_pad  , \key[47]_pad  , \key[48]_pad  , \key[49]_pad  , \key[4]_pad  , \key[50]_pad  , \key[51]_pad  , \key[52]_pad  , \key[53]_pad  , \key[54]_pad  , \key[55]_pad  , \key[56]_pad  , \key[57]_pad  , \key[58]_pad  , \key[59]_pad  , \key[5]_pad  , \key[60]_pad  , \key[61]_pad  , \key[62]_pad  , \key[63]_pad  , \key[64]_pad  , \key[65]_pad  , \key[66]_pad  , \key[67]_pad  , \key[68]_pad  , \key[69]_pad  , \key[6]_pad  , \key[70]_pad  , \key[71]_pad  , \key[72]_pad  , \key[73]_pad  , \key[74]_pad  , \key[75]_pad  , \key[76]_pad  , \key[77]_pad  , \key[78]_pad  , \key[79]_pad  , \key[7]_pad  , \key[80]_pad  , \key[81]_pad  , \key[82]_pad  , \key[83]_pad  , \key[84]_pad  , \key[85]_pad  , \key[86]_pad  , \key[87]_pad  , \key[88]_pad  , \key[89]_pad  , \key[8]_pad  , \key[90]_pad  , \key[91]_pad  , \key[92]_pad  , \key[93]_pad  , \key[94]_pad  , \key[95]_pad  , \key[96]_pad  , \key[97]_pad  , \key[98]_pad  , \key[99]_pad  , \key[9]_pad  , ld_pad , \ld_r_reg/P0001  , rst_pad , \sa00_reg[0]/P0001  , \sa00_reg[1]/P0001  , \sa00_reg[2]/P0001  , \sa00_reg[3]/P0001  , \sa00_reg[4]/P0001  , \sa00_reg[5]/P0001  , \sa00_reg[6]/NET0131  , \sa00_reg[7]/NET0131  , \sa01_reg[0]/P0001  , \sa01_reg[1]/P0001  , \sa01_reg[2]/P0001  , \sa01_reg[3]/P0001  , \sa01_reg[4]/P0001  , \sa01_reg[5]/P0001  , \sa01_reg[6]/NET0131  , \sa01_reg[7]/NET0131  , \sa02_reg[0]/P0001  , \sa02_reg[1]/P0001  , \sa02_reg[2]/P0001  , \sa02_reg[3]/P0001  , \sa02_reg[4]/P0001  , \sa02_reg[5]/P0001  , \sa02_reg[6]/NET0131  , \sa02_reg[7]/NET0131  , \sa03_reg[0]/P0001  , \sa03_reg[1]/P0001  , \sa03_reg[2]/P0001  , \sa03_reg[3]/P0001  , \sa03_reg[4]/P0001  , \sa03_reg[5]/P0001  , \sa03_reg[6]/NET0131  , \sa03_reg[7]/NET0131  , \sa10_reg[0]/P0001  , \sa10_reg[1]/P0001  , \sa10_reg[2]/P0001  , \sa10_reg[3]/P0001  , \sa10_reg[4]/P0001  , \sa10_reg[5]/P0001  , \sa10_reg[6]/NET0131  , \sa10_reg[7]/NET0131  , \sa11_reg[0]/P0001  , \sa11_reg[1]/P0001  , \sa11_reg[2]/P0001  , \sa11_reg[3]/P0001  , \sa11_reg[4]/P0001  , \sa11_reg[5]/P0001  , \sa11_reg[6]/NET0131  , \sa11_reg[7]/NET0131  , \sa12_reg[0]/P0001  , \sa12_reg[1]/P0001  , \sa12_reg[2]/P0001  , \sa12_reg[3]/P0001  , \sa12_reg[4]/P0001  , \sa12_reg[5]/P0001  , \sa12_reg[6]/NET0131  , \sa12_reg[7]/NET0131  , \sa13_reg[0]/P0001  , \sa13_reg[1]/P0001  , \sa13_reg[2]/P0001  , \sa13_reg[3]/P0001  , \sa13_reg[4]/P0001  , \sa13_reg[5]/P0001  , \sa13_reg[6]/NET0131  , \sa13_reg[7]/NET0131  , \sa20_reg[0]/P0001  , \sa20_reg[1]/P0001  , \sa20_reg[2]/P0001  , \sa20_reg[3]/P0001  , \sa20_reg[4]/P0001  , \sa20_reg[5]/P0001  , \sa20_reg[6]/NET0131  , \sa20_reg[7]/NET0131  , \sa21_reg[0]/P0001  , \sa21_reg[1]/P0001  , \sa21_reg[2]/P0001  , \sa21_reg[3]/P0001  , \sa21_reg[4]/P0001  , \sa21_reg[5]/P0001  , \sa21_reg[6]/NET0131  , \sa21_reg[7]/P0001  , \sa22_reg[0]/P0001  , \sa22_reg[1]/P0001  , \sa22_reg[2]/P0001  , \sa22_reg[3]/P0001  , \sa22_reg[4]/P0001  , \sa22_reg[5]/P0001  , \sa22_reg[6]/NET0131  , \sa22_reg[7]/NET0131  , \sa23_reg[0]/P0001  , \sa23_reg[1]/P0001  , \sa23_reg[2]/P0001  , \sa23_reg[3]/P0001  , \sa23_reg[4]/P0001  , \sa23_reg[5]/P0001  , \sa23_reg[6]/NET0131  , \sa23_reg[7]/NET0131  , \sa30_reg[0]/P0002  , \sa30_reg[1]/P0001  , \sa30_reg[2]/P0001  , \sa30_reg[3]/P0001  , \sa30_reg[4]/P0001  , \sa30_reg[5]/P0001  , \sa30_reg[6]/NET0131  , \sa30_reg[7]/P0001  , \sa31_reg[0]/P0002  , \sa31_reg[1]/P0001  , \sa31_reg[2]/P0001  , \sa31_reg[3]/P0001  , \sa31_reg[4]/P0001  , \sa31_reg[5]/P0001  , \sa31_reg[6]/NET0131  , \sa31_reg[7]/P0001  , \sa32_reg[0]/P0002  , \sa32_reg[1]/P0001  , \sa32_reg[2]/P0001  , \sa32_reg[3]/P0001  , \sa32_reg[4]/P0001  , \sa32_reg[5]/P0001  , \sa32_reg[6]/NET0131  , \sa32_reg[7]/P0001  , \sa33_reg[0]/P0001  , \sa33_reg[1]/P0001  , \sa33_reg[2]/P0001  , \sa33_reg[3]/P0001  , \sa33_reg[4]/P0001  , \sa33_reg[5]/P0001  , \sa33_reg[6]/P0001  , \sa33_reg[7]/NET0131  , \text_in_r_reg[0]/P0001  , \text_in_r_reg[100]/P0001  , \text_in_r_reg[101]/P0001  , \text_in_r_reg[102]/P0001  , \text_in_r_reg[103]/P0001  , \text_in_r_reg[104]/P0001  , \text_in_r_reg[105]/P0001  , \text_in_r_reg[106]/P0001  , \text_in_r_reg[107]/P0001  , \text_in_r_reg[108]/P0001  , \text_in_r_reg[109]/P0001  , \text_in_r_reg[10]/P0001  , \text_in_r_reg[110]/P0001  , \text_in_r_reg[111]/P0001  , \text_in_r_reg[112]/P0001  , \text_in_r_reg[113]/P0001  , \text_in_r_reg[114]/P0001  , \text_in_r_reg[115]/P0001  , \text_in_r_reg[116]/P0001  , \text_in_r_reg[117]/P0001  , \text_in_r_reg[118]/P0001  , \text_in_r_reg[119]/P0001  , \text_in_r_reg[11]/P0001  , \text_in_r_reg[120]/P0001  , \text_in_r_reg[121]/P0001  , \text_in_r_reg[122]/P0001  , \text_in_r_reg[123]/P0001  , \text_in_r_reg[124]/P0001  , \text_in_r_reg[125]/P0001  , \text_in_r_reg[126]/P0001  , \text_in_r_reg[127]/P0001  , \text_in_r_reg[12]/P0001  , \text_in_r_reg[13]/P0001  , \text_in_r_reg[14]/P0001  , \text_in_r_reg[15]/P0001  , \text_in_r_reg[16]/P0001  , \text_in_r_reg[17]/P0001  , \text_in_r_reg[18]/P0001  , \text_in_r_reg[19]/P0001  , \text_in_r_reg[1]/P0001  , \text_in_r_reg[20]/P0001  , \text_in_r_reg[21]/P0001  , \text_in_r_reg[22]/P0001  , \text_in_r_reg[23]/P0001  , \text_in_r_reg[24]/P0001  , \text_in_r_reg[25]/P0001  , \text_in_r_reg[26]/P0001  , \text_in_r_reg[27]/P0001  , \text_in_r_reg[28]/P0001  , \text_in_r_reg[29]/P0001  , \text_in_r_reg[2]/P0001  , \text_in_r_reg[30]/P0001  , \text_in_r_reg[31]/P0001  , \text_in_r_reg[32]/P0001  , \text_in_r_reg[33]/P0001  , \text_in_r_reg[34]/P0001  , \text_in_r_reg[35]/P0001  , \text_in_r_reg[36]/P0001  , \text_in_r_reg[37]/P0001  , \text_in_r_reg[38]/P0001  , \text_in_r_reg[39]/P0001  , \text_in_r_reg[3]/P0001  , \text_in_r_reg[40]/P0001  , \text_in_r_reg[41]/P0001  , \text_in_r_reg[42]/P0001  , \text_in_r_reg[43]/P0001  , \text_in_r_reg[44]/P0001  , \text_in_r_reg[45]/P0001  , \text_in_r_reg[46]/P0001  , \text_in_r_reg[47]/P0001  , \text_in_r_reg[48]/P0001  , \text_in_r_reg[49]/P0001  , \text_in_r_reg[4]/P0001  , \text_in_r_reg[50]/P0001  , \text_in_r_reg[51]/P0001  , \text_in_r_reg[52]/P0001  , \text_in_r_reg[53]/P0001  , \text_in_r_reg[54]/P0001  , \text_in_r_reg[55]/P0001  , \text_in_r_reg[56]/P0001  , \text_in_r_reg[57]/P0001  , \text_in_r_reg[58]/P0001  , \text_in_r_reg[59]/P0001  , \text_in_r_reg[5]/P0001  , \text_in_r_reg[60]/P0001  , \text_in_r_reg[61]/P0001  , \text_in_r_reg[62]/P0001  , \text_in_r_reg[63]/P0001  , \text_in_r_reg[64]/P0001  , \text_in_r_reg[65]/P0001  , \text_in_r_reg[66]/P0001  , \text_in_r_reg[67]/P0001  , \text_in_r_reg[68]/P0001  , \text_in_r_reg[69]/P0001  , \text_in_r_reg[6]/P0001  , \text_in_r_reg[70]/P0001  , \text_in_r_reg[71]/P0001  , \text_in_r_reg[72]/P0001  , \text_in_r_reg[73]/P0001  , \text_in_r_reg[74]/P0001  , \text_in_r_reg[75]/P0001  , \text_in_r_reg[76]/P0001  , \text_in_r_reg[77]/P0001  , \text_in_r_reg[78]/P0001  , \text_in_r_reg[79]/P0001  , \text_in_r_reg[7]/P0001  , \text_in_r_reg[80]/P0001  , \text_in_r_reg[81]/P0001  , \text_in_r_reg[82]/P0001  , \text_in_r_reg[83]/P0001  , \text_in_r_reg[84]/P0001  , \text_in_r_reg[85]/P0001  , \text_in_r_reg[86]/P0001  , \text_in_r_reg[87]/P0001  , \text_in_r_reg[88]/P0001  , \text_in_r_reg[89]/P0001  , \text_in_r_reg[8]/P0001  , \text_in_r_reg[90]/P0001  , \text_in_r_reg[91]/P0001  , \text_in_r_reg[92]/P0001  , \text_in_r_reg[93]/P0001  , \text_in_r_reg[94]/P0001  , \text_in_r_reg[95]/P0001  , \text_in_r_reg[96]/P0001  , \text_in_r_reg[97]/P0001  , \text_in_r_reg[98]/P0001  , \text_in_r_reg[99]/P0001  , \text_in_r_reg[9]/P0001  , \u0_r0_out_reg[24]/P0001  , \u0_r0_out_reg[25]/P0001  , \u0_r0_out_reg[26]/P0001  , \u0_r0_out_reg[27]/P0001  , \u0_r0_out_reg[28]/P0001  , \u0_r0_out_reg[29]/P0001  , \u0_r0_out_reg[30]/P0001  , \u0_r0_out_reg[31]/P0001  , \u0_r0_rcnt_reg[0]/P0001  , \u0_r0_rcnt_reg[1]/P0001  , \u0_r0_rcnt_reg[2]/P0001  , \u0_r0_rcnt_reg[3]/P0001  , \u0_w_reg[0][0]/P0001  , \u0_w_reg[0][10]/P0001  , \u0_w_reg[0][11]/P0001  , \u0_w_reg[0][12]/P0001  , \u0_w_reg[0][13]/P0001  , \u0_w_reg[0][14]/P0001  , \u0_w_reg[0][15]/P0001  , \u0_w_reg[0][16]/P0001  , \u0_w_reg[0][17]/P0001  , \u0_w_reg[0][18]/P0001  , \u0_w_reg[0][19]/P0001  , \u0_w_reg[0][1]/P0001  , \u0_w_reg[0][20]/P0001  , \u0_w_reg[0][21]/P0001  , \u0_w_reg[0][22]/P0001  , \u0_w_reg[0][23]/P0001  , \u0_w_reg[0][24]/P0001  , \u0_w_reg[0][25]/P0001  , \u0_w_reg[0][26]/P0001  , \u0_w_reg[0][27]/P0001  , \u0_w_reg[0][28]/P0001  , \u0_w_reg[0][29]/P0001  , \u0_w_reg[0][2]/P0001  , \u0_w_reg[0][30]/P0001  , \u0_w_reg[0][31]/P0001  , \u0_w_reg[0][3]/P0001  , \u0_w_reg[0][4]/P0001  , \u0_w_reg[0][5]/P0001  , \u0_w_reg[0][6]/P0001  , \u0_w_reg[0][7]/P0001  , \u0_w_reg[0][8]/P0001  , \u0_w_reg[0][9]/P0001  , \u0_w_reg[1][0]/P0001  , \u0_w_reg[1][10]/P0001  , \u0_w_reg[1][11]/P0001  , \u0_w_reg[1][12]/P0001  , \u0_w_reg[1][13]/P0001  , \u0_w_reg[1][14]/P0001  , \u0_w_reg[1][15]/P0001  , \u0_w_reg[1][16]/P0001  , \u0_w_reg[1][17]/P0001  , \u0_w_reg[1][18]/P0001  , \u0_w_reg[1][19]/P0001  , \u0_w_reg[1][1]/P0001  , \u0_w_reg[1][20]/P0001  , \u0_w_reg[1][21]/P0001  , \u0_w_reg[1][22]/P0001  , \u0_w_reg[1][23]/P0001  , \u0_w_reg[1][24]/P0002  , \u0_w_reg[1][25]/P0001  , \u0_w_reg[1][26]/P0001  , \u0_w_reg[1][27]/P0001  , \u0_w_reg[1][28]/P0001  , \u0_w_reg[1][29]/P0002  , \u0_w_reg[1][2]/P0001  , \u0_w_reg[1][30]/P0001  , \u0_w_reg[1][31]/P0001  , \u0_w_reg[1][3]/P0001  , \u0_w_reg[1][4]/P0001  , \u0_w_reg[1][5]/P0001  , \u0_w_reg[1][6]/P0001  , \u0_w_reg[1][7]/P0001  , \u0_w_reg[1][8]/P0001  , \u0_w_reg[1][9]/P0001  , \u0_w_reg[2][0]/P0001  , \u0_w_reg[2][10]/P0001  , \u0_w_reg[2][11]/P0001  , \u0_w_reg[2][12]/P0001  , \u0_w_reg[2][13]/P0001  , \u0_w_reg[2][14]/P0001  , \u0_w_reg[2][15]/P0001  , \u0_w_reg[2][16]/P0001  , \u0_w_reg[2][17]/P0001  , \u0_w_reg[2][18]/P0001  , \u0_w_reg[2][19]/P0001  , \u0_w_reg[2][1]/P0001  , \u0_w_reg[2][20]/P0001  , \u0_w_reg[2][21]/P0001  , \u0_w_reg[2][22]/P0001  , \u0_w_reg[2][23]/P0001  , \u0_w_reg[2][24]/P0001  , \u0_w_reg[2][25]/P0001  , \u0_w_reg[2][26]/P0001  , \u0_w_reg[2][27]/P0001  , \u0_w_reg[2][28]/P0001  , \u0_w_reg[2][29]/P0001  , \u0_w_reg[2][2]/P0001  , \u0_w_reg[2][30]/P0001  , \u0_w_reg[2][31]/P0001  , \u0_w_reg[2][3]/P0001  , \u0_w_reg[2][4]/P0001  , \u0_w_reg[2][5]/P0001  , \u0_w_reg[2][6]/P0001  , \u0_w_reg[2][7]/P0001  , \u0_w_reg[2][8]/P0001  , \u0_w_reg[2][9]/P0001  , \u0_w_reg[3][0]/P0001  , \u0_w_reg[3][10]/P0001  , \u0_w_reg[3][11]/P0001  , \u0_w_reg[3][12]/P0001  , \u0_w_reg[3][13]/P0001  , \u0_w_reg[3][14]/P0001  , \u0_w_reg[3][15]/P0001  , \u0_w_reg[3][16]/P0001  , \u0_w_reg[3][17]/P0001  , \u0_w_reg[3][18]/P0001  , \u0_w_reg[3][19]/P0001  , \u0_w_reg[3][1]/P0001  , \u0_w_reg[3][20]/P0001  , \u0_w_reg[3][21]/P0001  , \u0_w_reg[3][22]/P0001  , \u0_w_reg[3][23]/P0001  , \u0_w_reg[3][24]/P0001  , \u0_w_reg[3][25]/P0001  , \u0_w_reg[3][26]/P0001  , \u0_w_reg[3][27]/P0001  , \u0_w_reg[3][28]/P0001  , \u0_w_reg[3][29]/P0001  , \u0_w_reg[3][2]/P0001  , \u0_w_reg[3][30]/P0001  , \u0_w_reg[3][31]/P0001  , \u0_w_reg[3][3]/P0001  , \u0_w_reg[3][4]/P0001  , \u0_w_reg[3][5]/P0001  , \u0_w_reg[3][6]/P0001  , \u0_w_reg[3][7]/P0001  , \u0_w_reg[3][8]/P0001  , \u0_w_reg[3][9]/P0001  , \_al_n0  , \_al_n1  , \g21/_0_  , \g56610/_0_  , \g56611/_0_  , \g56612/_0_  , \g56613/_0_  , \g56614/_0_  , \g56615/_0_  , \g56616/_0_  , \g56617/_0_  , \g56630/_0_  , \g56631/_0_  , \g56632/_0_  , \g56633/_0_  , \g56634/_0_  , \g56635/_0_  , \g56645/_0_  , \g56646/_0_  , \g56647/_0_  , \g56648/_0_  , \g56649/_0_  , \g56650/_0_  , \g56651/_0_  , \g56652/_0_  , \g56666/_0_  , \g56667/_0_  , \g56668/_0_  , \g56669/_0_  , \g56670/_0_  , \g56671/_0_  , \g56672/_0_  , \g56674/_0_  , \g56675/_0_  , \g56704/_0_  , \g56739/_0_  , \g56743/_0_  , \g56763/_0_  , \g56776/_0_  , \g56812/_0_  , \g56818/_0_  , \g56861/_0_  , \g56874/_0_  , \g56919/_0_  , \g56920/_0_  , \g56921/_0_  , \g56923/_0_  , \g56924/_0_  , \g56925/_0_  , \g56926/_0_  , \g56956/_0_  , \g56957/_0_  , \g56958/_0_  , \g56959/_0_  , \g56960/_0_  , \g56961/_0_  , \g56972/_0_  , \g56973/_0_  , \g56974/_0_  , \g56976/_0_  , \g56977/_0_  , \g56978/_0_  , \g56979/_0_  , \g56980/_0_  , \g57008/_0_  , \g57010/_0_  , \g57011/_0_  , \g57012/_0_  , \g57013/_0_  , \g57014/_0_  , \g57015/_0_  , \g57016/_0_  , \g57017/_0_  , \g57086/_0_  , \g57091/_0_  , \g57114/_0_  , \g57129/_0_  , \g57163/_0_  , \g57171/_0_  , \g57204/_0_  , \g57218/_0_  , \g57262/_0_  , \g57263/_0_  , \g57264/_0_  , \g57265/_0_  , \g57266/_0_  , \g57267/_0_  , \g57268/_0_  , \g57269/_0_  , \g57300/_0_  , \g57301/_0_  , \g57302/_0_  , \g57303/_0_  , \g57304/_0_  , \g57316/_0_  , \g57317/_0_  , \g57319/_0_  , \g57320/_0_  , \g57321/_0_  , \g57322/_0_  , \g57323/_0_  , \g57324/_0_  , \g57350/_0_  , \g57353/_0_  , \g57354/_0_  , \g57355/_0_  , \g57356/_0_  , \g57357/_0_  , \g57358/_0_  , \g57359/_0_  , \g57360/_0_  , \g57427/_0_  , \g57432/_0_  , \g57456/_0_  , \g57471/_0_  , \g57506/_0_  , \g57512/_0_  , \g57540/_0_  , \g57547/_0_  , \g57654/_0_  , \g57655/_0_  , \g57656/_0_  , \g57657/_0_  , \g57658/_0_  , \g57676/_0_  , \g57677/_0_  , \g57678/_0_  , \g57679/_0_  , \g57680/_0_  , \g57681/_0_  , \g57682/_0_  , \g57683/_0_  , \g57684/_0_  , \g57685/_0_  , \g57686/_0_  , \g57687/_0_  , \g57688/_0_  , \g57689/_0_  , \g57690/_0_  , \g57691/_0_  , \g57700/_0_  , \g57701/_0_  , \g57702/_0_  , \g57703/_0_  , \g57704/_0_  , \g57705/_0_  , \g57706/_0_  , \g57707/_0_  , \g57708/_0_  , \g57709/_3_  , \g57710/_3_  , \g57711/_0_  , \g57712/_3_  , \g57715/_3_  , \g57716/_3_  , \g57767/_0_  , \g57768/_3_  , \g57769/_3_  , \g57770/_3_  , \g57771/_3_  , \g57777/_3_  , \g57779/_3_  , \g57804/_3_  , \g57805/_3_  , \g57806/_3_  , \g57807/_3_  , \g57808/_3_  , \g57809/_3_  , \g57810/_3_  , \g57811/_3_  , \g57812/_3_  , \g57813/_3_  , \g57814/_3_  , \g57815/_3_  , \g57816/_0_  , \g57817/_3_  , \g57818/_3_  , \g57819/_3_  , \g57822/_3_  , \g57823/_3_  , \g57824/_3_  , \g57830/_3_  , \g57835/_3_  , \g57836/_3_  , \g57837/_3_  , \g57841/_3_  , \g57842/_3_  , \g57843/_3_  , \g57854/_3_  , \g57855/_3_  , \g57856/_3_  , \g57857/_3_  , \g57858/_3_  , \g57859/_3_  , \g57860/_3_  , \g57861/_3_  , \g57871/_3_  , \g57872/_3_  , \g57874/_3_  , \g57968/_3_  , \g57969/_3_  , \g57970/_3_  , \g57971/_3_  , \g57980/_3_  , \g57983/_3_  , \g57984/_3_  , \g57985/_3_  , \g58012/_3_  , \g58013/_3_  , \g58015/_3_  , \g58057/_3_  , \g58058/_3_  , \g58059/_3_  , \g58189/_3_  , \g58190/_3_  , \g58191/_3_  , \g58192/_3_  , \g58193/_3_  , \g58194/_3_  , \g58195/_3_  , \g58196/_3_  , \g58197/_3_  , \g58224/_3_  , \g58226/_3_  , \g58229/_3_  , \g58255/_3_  , \g58256/_3_  , \g58257/_3_  , \g58258/_3_  , \g58259/_3_  , \g58260/_3_  , \g58261/_3_  , \g58262/_3_  , \g58263/_3_  , \g58264/_3_  , \g58265/_3_  , \g58266/_3_  , \g58267/_3_  , \g58268/_3_  , \g58269/_3_  , \g58270/_0_  , \g58271/_3_  , \g58272/_3_  , \g58273/_3_  , \g58274/_3_  , \g58275/_3_  , \g58276/_3_  , \g58277/_3_  , \g58278/_3_  , \g58279/_3_  , \g58285/_3_  , \g58286/_3_  , \g58288/_3_  , \g58289/_3_  , \g58290/_3_  , \g58292/_3_  , \g58294/_3_  , \g58295/_3_  , \g58297/_3_  , \g58330/_0_  , \g58331/_0_  , \g58332/_0_  , \g58333/_0_  , \g58444/_3_  , \g58445/_3_  , \g58446/_3_  , \g58462/_0_  , \g58506/_0_  , \g58507/_0_  , \g58508/_0_  , \g58509/_0_  , \g58531/_0_  , \g58532/_0_  , \g58533/_0_  , \g58550/_0_  , \g58551/_0_  , \g58552/_0_  , \g58553/_0_  , \g58554/_0_  , \g58555/_0_  , \g58556/_0_  , \g58557/_0_  , \g58558/_0_  , \g58559/_0_  , \g58560/_0_  , \g58600/_3_  , \g58601/_3_  , \g58602/_3_  , \g58603/_3_  , \g58604/_3_  , \g58605/_3_  , \g58606/_3_  , \g58607/_3_  , \g58608/_3_  , \g58611/_0_  , \g58612/_0_  , \g58613/_0_  , \g58614/_0_  , \g58617/_0_  , \g58618/_0_  , \g58619/_0_  , \g58634/_0_  , \g58635/_0_  , \g58636/_0_  , \g58637/_0_  , \g58638/_0_  , \g58639/_0_  , \g58640/_0_  , \g58641/_0_  , \g58829/_3_  , \g58830/_3_  , \g58831/_3_  , \g58832/_3_  , \g58833/_3_  , \g58834/_3_  , \g58835/_0_  , \g58844/_0_  , \g58902/_0_  , \g58903/_0_  , \g58904/_0_  , \g58905/_0_  , \g58910/_0_  , \g58913/_0_  , \g58934/_0_  , \g58935/_0_  , \g58936/_0_  , \g58937/_0_  , \g58938/_0_  , \g58970/_0_  , \g58972/_0_  , \g58994/_0_  , \g58995/_0_  , \g58996/_0_  , \g58997/_0_  , \g58998/_0_  , \g58999/_0_  , \g59000/_0_  , \g59002/_0_  , \g59003/_0_  , \g59004/_0_  , \g59254/_0_  , \g59257/_0_  , \g59258/_0_  , \g59259/_0_  , \g59276/_0_  , \g59277/_0_  , \g59278/_0_  , \g59279/_0_  , \g59280/_0_  , \g59291/_0_  , \g59292/_0_  , \g59293/_0_  , \g59294/_0_  , \g59295/_0_  , \g59308/_0_  , \g59309/_0_  , \g59310/_0_  , \g59311/_0_  , \g59330/_0_  , \g59331/_0_  , \g59332/_0_  , \g59333/_0_  , \g59334/_0_  , \g59335/_0_  , \g59336/_0_  , \g59337/_0_  , \g59338/_0_  , \g59339/_0_  , \g59596/_0_  , \g59597/_0_  , \g59598/_0_  , \g59599/_0_  , \g59625/_0_  , \g59626/_0_  , \g59627/_0_  , \g59628/_0_  , \g59837/_0_  , \g59838/_0_  , \g59839/_0_  , \g59840/_0_  , \g60090/_0_  , \g60320/_0_  , \g60321/_0_  , \g60409/_0_  , \g60539/_0_  , \g60860/_0_  , \g60977/_0_  , \g61012/_0_  , \g61185/_0_  , \g61524/_2_  , \g61776/_0_  , \g61895/_0_  , \g61897/_0_  , \g62220/_0_  , \g65958/_0_  , \g72347/_3_  , \g77848/_0_  , \g85056/_0_  , \sa30_reg[0]/_05_  , \sa31_reg[0]/_05_  , \sa32_reg[0]/_05_  , \u0_w_reg[1][24]/_05_  , \u0_w_reg[1][29]/_05_  );
  input \dcnt_reg[0]/P0001  ;
  input \dcnt_reg[1]/P0001  ;
  input \dcnt_reg[2]/P0001  ;
  input \dcnt_reg[3]/P0001  ;
  input \key[0]_pad  ;
  input \key[100]_pad  ;
  input \key[101]_pad  ;
  input \key[102]_pad  ;
  input \key[103]_pad  ;
  input \key[104]_pad  ;
  input \key[105]_pad  ;
  input \key[106]_pad  ;
  input \key[107]_pad  ;
  input \key[108]_pad  ;
  input \key[109]_pad  ;
  input \key[10]_pad  ;
  input \key[110]_pad  ;
  input \key[111]_pad  ;
  input \key[112]_pad  ;
  input \key[113]_pad  ;
  input \key[114]_pad  ;
  input \key[115]_pad  ;
  input \key[116]_pad  ;
  input \key[117]_pad  ;
  input \key[118]_pad  ;
  input \key[119]_pad  ;
  input \key[11]_pad  ;
  input \key[120]_pad  ;
  input \key[121]_pad  ;
  input \key[122]_pad  ;
  input \key[123]_pad  ;
  input \key[124]_pad  ;
  input \key[125]_pad  ;
  input \key[126]_pad  ;
  input \key[127]_pad  ;
  input \key[12]_pad  ;
  input \key[13]_pad  ;
  input \key[14]_pad  ;
  input \key[15]_pad  ;
  input \key[16]_pad  ;
  input \key[17]_pad  ;
  input \key[18]_pad  ;
  input \key[19]_pad  ;
  input \key[1]_pad  ;
  input \key[20]_pad  ;
  input \key[21]_pad  ;
  input \key[22]_pad  ;
  input \key[23]_pad  ;
  input \key[24]_pad  ;
  input \key[25]_pad  ;
  input \key[26]_pad  ;
  input \key[27]_pad  ;
  input \key[28]_pad  ;
  input \key[29]_pad  ;
  input \key[2]_pad  ;
  input \key[30]_pad  ;
  input \key[31]_pad  ;
  input \key[32]_pad  ;
  input \key[33]_pad  ;
  input \key[34]_pad  ;
  input \key[35]_pad  ;
  input \key[36]_pad  ;
  input \key[37]_pad  ;
  input \key[38]_pad  ;
  input \key[39]_pad  ;
  input \key[3]_pad  ;
  input \key[40]_pad  ;
  input \key[41]_pad  ;
  input \key[42]_pad  ;
  input \key[43]_pad  ;
  input \key[44]_pad  ;
  input \key[45]_pad  ;
  input \key[46]_pad  ;
  input \key[47]_pad  ;
  input \key[48]_pad  ;
  input \key[49]_pad  ;
  input \key[4]_pad  ;
  input \key[50]_pad  ;
  input \key[51]_pad  ;
  input \key[52]_pad  ;
  input \key[53]_pad  ;
  input \key[54]_pad  ;
  input \key[55]_pad  ;
  input \key[56]_pad  ;
  input \key[57]_pad  ;
  input \key[58]_pad  ;
  input \key[59]_pad  ;
  input \key[5]_pad  ;
  input \key[60]_pad  ;
  input \key[61]_pad  ;
  input \key[62]_pad  ;
  input \key[63]_pad  ;
  input \key[64]_pad  ;
  input \key[65]_pad  ;
  input \key[66]_pad  ;
  input \key[67]_pad  ;
  input \key[68]_pad  ;
  input \key[69]_pad  ;
  input \key[6]_pad  ;
  input \key[70]_pad  ;
  input \key[71]_pad  ;
  input \key[72]_pad  ;
  input \key[73]_pad  ;
  input \key[74]_pad  ;
  input \key[75]_pad  ;
  input \key[76]_pad  ;
  input \key[77]_pad  ;
  input \key[78]_pad  ;
  input \key[79]_pad  ;
  input \key[7]_pad  ;
  input \key[80]_pad  ;
  input \key[81]_pad  ;
  input \key[82]_pad  ;
  input \key[83]_pad  ;
  input \key[84]_pad  ;
  input \key[85]_pad  ;
  input \key[86]_pad  ;
  input \key[87]_pad  ;
  input \key[88]_pad  ;
  input \key[89]_pad  ;
  input \key[8]_pad  ;
  input \key[90]_pad  ;
  input \key[91]_pad  ;
  input \key[92]_pad  ;
  input \key[93]_pad  ;
  input \key[94]_pad  ;
  input \key[95]_pad  ;
  input \key[96]_pad  ;
  input \key[97]_pad  ;
  input \key[98]_pad  ;
  input \key[99]_pad  ;
  input \key[9]_pad  ;
  input ld_pad ;
  input \ld_r_reg/P0001  ;
  input rst_pad ;
  input \sa00_reg[0]/P0001  ;
  input \sa00_reg[1]/P0001  ;
  input \sa00_reg[2]/P0001  ;
  input \sa00_reg[3]/P0001  ;
  input \sa00_reg[4]/P0001  ;
  input \sa00_reg[5]/P0001  ;
  input \sa00_reg[6]/NET0131  ;
  input \sa00_reg[7]/NET0131  ;
  input \sa01_reg[0]/P0001  ;
  input \sa01_reg[1]/P0001  ;
  input \sa01_reg[2]/P0001  ;
  input \sa01_reg[3]/P0001  ;
  input \sa01_reg[4]/P0001  ;
  input \sa01_reg[5]/P0001  ;
  input \sa01_reg[6]/NET0131  ;
  input \sa01_reg[7]/NET0131  ;
  input \sa02_reg[0]/P0001  ;
  input \sa02_reg[1]/P0001  ;
  input \sa02_reg[2]/P0001  ;
  input \sa02_reg[3]/P0001  ;
  input \sa02_reg[4]/P0001  ;
  input \sa02_reg[5]/P0001  ;
  input \sa02_reg[6]/NET0131  ;
  input \sa02_reg[7]/NET0131  ;
  input \sa03_reg[0]/P0001  ;
  input \sa03_reg[1]/P0001  ;
  input \sa03_reg[2]/P0001  ;
  input \sa03_reg[3]/P0001  ;
  input \sa03_reg[4]/P0001  ;
  input \sa03_reg[5]/P0001  ;
  input \sa03_reg[6]/NET0131  ;
  input \sa03_reg[7]/NET0131  ;
  input \sa10_reg[0]/P0001  ;
  input \sa10_reg[1]/P0001  ;
  input \sa10_reg[2]/P0001  ;
  input \sa10_reg[3]/P0001  ;
  input \sa10_reg[4]/P0001  ;
  input \sa10_reg[5]/P0001  ;
  input \sa10_reg[6]/NET0131  ;
  input \sa10_reg[7]/NET0131  ;
  input \sa11_reg[0]/P0001  ;
  input \sa11_reg[1]/P0001  ;
  input \sa11_reg[2]/P0001  ;
  input \sa11_reg[3]/P0001  ;
  input \sa11_reg[4]/P0001  ;
  input \sa11_reg[5]/P0001  ;
  input \sa11_reg[6]/NET0131  ;
  input \sa11_reg[7]/NET0131  ;
  input \sa12_reg[0]/P0001  ;
  input \sa12_reg[1]/P0001  ;
  input \sa12_reg[2]/P0001  ;
  input \sa12_reg[3]/P0001  ;
  input \sa12_reg[4]/P0001  ;
  input \sa12_reg[5]/P0001  ;
  input \sa12_reg[6]/NET0131  ;
  input \sa12_reg[7]/NET0131  ;
  input \sa13_reg[0]/P0001  ;
  input \sa13_reg[1]/P0001  ;
  input \sa13_reg[2]/P0001  ;
  input \sa13_reg[3]/P0001  ;
  input \sa13_reg[4]/P0001  ;
  input \sa13_reg[5]/P0001  ;
  input \sa13_reg[6]/NET0131  ;
  input \sa13_reg[7]/NET0131  ;
  input \sa20_reg[0]/P0001  ;
  input \sa20_reg[1]/P0001  ;
  input \sa20_reg[2]/P0001  ;
  input \sa20_reg[3]/P0001  ;
  input \sa20_reg[4]/P0001  ;
  input \sa20_reg[5]/P0001  ;
  input \sa20_reg[6]/NET0131  ;
  input \sa20_reg[7]/NET0131  ;
  input \sa21_reg[0]/P0001  ;
  input \sa21_reg[1]/P0001  ;
  input \sa21_reg[2]/P0001  ;
  input \sa21_reg[3]/P0001  ;
  input \sa21_reg[4]/P0001  ;
  input \sa21_reg[5]/P0001  ;
  input \sa21_reg[6]/NET0131  ;
  input \sa21_reg[7]/P0001  ;
  input \sa22_reg[0]/P0001  ;
  input \sa22_reg[1]/P0001  ;
  input \sa22_reg[2]/P0001  ;
  input \sa22_reg[3]/P0001  ;
  input \sa22_reg[4]/P0001  ;
  input \sa22_reg[5]/P0001  ;
  input \sa22_reg[6]/NET0131  ;
  input \sa22_reg[7]/NET0131  ;
  input \sa23_reg[0]/P0001  ;
  input \sa23_reg[1]/P0001  ;
  input \sa23_reg[2]/P0001  ;
  input \sa23_reg[3]/P0001  ;
  input \sa23_reg[4]/P0001  ;
  input \sa23_reg[5]/P0001  ;
  input \sa23_reg[6]/NET0131  ;
  input \sa23_reg[7]/NET0131  ;
  input \sa30_reg[0]/P0002  ;
  input \sa30_reg[1]/P0001  ;
  input \sa30_reg[2]/P0001  ;
  input \sa30_reg[3]/P0001  ;
  input \sa30_reg[4]/P0001  ;
  input \sa30_reg[5]/P0001  ;
  input \sa30_reg[6]/NET0131  ;
  input \sa30_reg[7]/P0001  ;
  input \sa31_reg[0]/P0002  ;
  input \sa31_reg[1]/P0001  ;
  input \sa31_reg[2]/P0001  ;
  input \sa31_reg[3]/P0001  ;
  input \sa31_reg[4]/P0001  ;
  input \sa31_reg[5]/P0001  ;
  input \sa31_reg[6]/NET0131  ;
  input \sa31_reg[7]/P0001  ;
  input \sa32_reg[0]/P0002  ;
  input \sa32_reg[1]/P0001  ;
  input \sa32_reg[2]/P0001  ;
  input \sa32_reg[3]/P0001  ;
  input \sa32_reg[4]/P0001  ;
  input \sa32_reg[5]/P0001  ;
  input \sa32_reg[6]/NET0131  ;
  input \sa32_reg[7]/P0001  ;
  input \sa33_reg[0]/P0001  ;
  input \sa33_reg[1]/P0001  ;
  input \sa33_reg[2]/P0001  ;
  input \sa33_reg[3]/P0001  ;
  input \sa33_reg[4]/P0001  ;
  input \sa33_reg[5]/P0001  ;
  input \sa33_reg[6]/P0001  ;
  input \sa33_reg[7]/NET0131  ;
  input \text_in_r_reg[0]/P0001  ;
  input \text_in_r_reg[100]/P0001  ;
  input \text_in_r_reg[101]/P0001  ;
  input \text_in_r_reg[102]/P0001  ;
  input \text_in_r_reg[103]/P0001  ;
  input \text_in_r_reg[104]/P0001  ;
  input \text_in_r_reg[105]/P0001  ;
  input \text_in_r_reg[106]/P0001  ;
  input \text_in_r_reg[107]/P0001  ;
  input \text_in_r_reg[108]/P0001  ;
  input \text_in_r_reg[109]/P0001  ;
  input \text_in_r_reg[10]/P0001  ;
  input \text_in_r_reg[110]/P0001  ;
  input \text_in_r_reg[111]/P0001  ;
  input \text_in_r_reg[112]/P0001  ;
  input \text_in_r_reg[113]/P0001  ;
  input \text_in_r_reg[114]/P0001  ;
  input \text_in_r_reg[115]/P0001  ;
  input \text_in_r_reg[116]/P0001  ;
  input \text_in_r_reg[117]/P0001  ;
  input \text_in_r_reg[118]/P0001  ;
  input \text_in_r_reg[119]/P0001  ;
  input \text_in_r_reg[11]/P0001  ;
  input \text_in_r_reg[120]/P0001  ;
  input \text_in_r_reg[121]/P0001  ;
  input \text_in_r_reg[122]/P0001  ;
  input \text_in_r_reg[123]/P0001  ;
  input \text_in_r_reg[124]/P0001  ;
  input \text_in_r_reg[125]/P0001  ;
  input \text_in_r_reg[126]/P0001  ;
  input \text_in_r_reg[127]/P0001  ;
  input \text_in_r_reg[12]/P0001  ;
  input \text_in_r_reg[13]/P0001  ;
  input \text_in_r_reg[14]/P0001  ;
  input \text_in_r_reg[15]/P0001  ;
  input \text_in_r_reg[16]/P0001  ;
  input \text_in_r_reg[17]/P0001  ;
  input \text_in_r_reg[18]/P0001  ;
  input \text_in_r_reg[19]/P0001  ;
  input \text_in_r_reg[1]/P0001  ;
  input \text_in_r_reg[20]/P0001  ;
  input \text_in_r_reg[21]/P0001  ;
  input \text_in_r_reg[22]/P0001  ;
  input \text_in_r_reg[23]/P0001  ;
  input \text_in_r_reg[24]/P0001  ;
  input \text_in_r_reg[25]/P0001  ;
  input \text_in_r_reg[26]/P0001  ;
  input \text_in_r_reg[27]/P0001  ;
  input \text_in_r_reg[28]/P0001  ;
  input \text_in_r_reg[29]/P0001  ;
  input \text_in_r_reg[2]/P0001  ;
  input \text_in_r_reg[30]/P0001  ;
  input \text_in_r_reg[31]/P0001  ;
  input \text_in_r_reg[32]/P0001  ;
  input \text_in_r_reg[33]/P0001  ;
  input \text_in_r_reg[34]/P0001  ;
  input \text_in_r_reg[35]/P0001  ;
  input \text_in_r_reg[36]/P0001  ;
  input \text_in_r_reg[37]/P0001  ;
  input \text_in_r_reg[38]/P0001  ;
  input \text_in_r_reg[39]/P0001  ;
  input \text_in_r_reg[3]/P0001  ;
  input \text_in_r_reg[40]/P0001  ;
  input \text_in_r_reg[41]/P0001  ;
  input \text_in_r_reg[42]/P0001  ;
  input \text_in_r_reg[43]/P0001  ;
  input \text_in_r_reg[44]/P0001  ;
  input \text_in_r_reg[45]/P0001  ;
  input \text_in_r_reg[46]/P0001  ;
  input \text_in_r_reg[47]/P0001  ;
  input \text_in_r_reg[48]/P0001  ;
  input \text_in_r_reg[49]/P0001  ;
  input \text_in_r_reg[4]/P0001  ;
  input \text_in_r_reg[50]/P0001  ;
  input \text_in_r_reg[51]/P0001  ;
  input \text_in_r_reg[52]/P0001  ;
  input \text_in_r_reg[53]/P0001  ;
  input \text_in_r_reg[54]/P0001  ;
  input \text_in_r_reg[55]/P0001  ;
  input \text_in_r_reg[56]/P0001  ;
  input \text_in_r_reg[57]/P0001  ;
  input \text_in_r_reg[58]/P0001  ;
  input \text_in_r_reg[59]/P0001  ;
  input \text_in_r_reg[5]/P0001  ;
  input \text_in_r_reg[60]/P0001  ;
  input \text_in_r_reg[61]/P0001  ;
  input \text_in_r_reg[62]/P0001  ;
  input \text_in_r_reg[63]/P0001  ;
  input \text_in_r_reg[64]/P0001  ;
  input \text_in_r_reg[65]/P0001  ;
  input \text_in_r_reg[66]/P0001  ;
  input \text_in_r_reg[67]/P0001  ;
  input \text_in_r_reg[68]/P0001  ;
  input \text_in_r_reg[69]/P0001  ;
  input \text_in_r_reg[6]/P0001  ;
  input \text_in_r_reg[70]/P0001  ;
  input \text_in_r_reg[71]/P0001  ;
  input \text_in_r_reg[72]/P0001  ;
  input \text_in_r_reg[73]/P0001  ;
  input \text_in_r_reg[74]/P0001  ;
  input \text_in_r_reg[75]/P0001  ;
  input \text_in_r_reg[76]/P0001  ;
  input \text_in_r_reg[77]/P0001  ;
  input \text_in_r_reg[78]/P0001  ;
  input \text_in_r_reg[79]/P0001  ;
  input \text_in_r_reg[7]/P0001  ;
  input \text_in_r_reg[80]/P0001  ;
  input \text_in_r_reg[81]/P0001  ;
  input \text_in_r_reg[82]/P0001  ;
  input \text_in_r_reg[83]/P0001  ;
  input \text_in_r_reg[84]/P0001  ;
  input \text_in_r_reg[85]/P0001  ;
  input \text_in_r_reg[86]/P0001  ;
  input \text_in_r_reg[87]/P0001  ;
  input \text_in_r_reg[88]/P0001  ;
  input \text_in_r_reg[89]/P0001  ;
  input \text_in_r_reg[8]/P0001  ;
  input \text_in_r_reg[90]/P0001  ;
  input \text_in_r_reg[91]/P0001  ;
  input \text_in_r_reg[92]/P0001  ;
  input \text_in_r_reg[93]/P0001  ;
  input \text_in_r_reg[94]/P0001  ;
  input \text_in_r_reg[95]/P0001  ;
  input \text_in_r_reg[96]/P0001  ;
  input \text_in_r_reg[97]/P0001  ;
  input \text_in_r_reg[98]/P0001  ;
  input \text_in_r_reg[99]/P0001  ;
  input \text_in_r_reg[9]/P0001  ;
  input \u0_r0_out_reg[24]/P0001  ;
  input \u0_r0_out_reg[25]/P0001  ;
  input \u0_r0_out_reg[26]/P0001  ;
  input \u0_r0_out_reg[27]/P0001  ;
  input \u0_r0_out_reg[28]/P0001  ;
  input \u0_r0_out_reg[29]/P0001  ;
  input \u0_r0_out_reg[30]/P0001  ;
  input \u0_r0_out_reg[31]/P0001  ;
  input \u0_r0_rcnt_reg[0]/P0001  ;
  input \u0_r0_rcnt_reg[1]/P0001  ;
  input \u0_r0_rcnt_reg[2]/P0001  ;
  input \u0_r0_rcnt_reg[3]/P0001  ;
  input \u0_w_reg[0][0]/P0001  ;
  input \u0_w_reg[0][10]/P0001  ;
  input \u0_w_reg[0][11]/P0001  ;
  input \u0_w_reg[0][12]/P0001  ;
  input \u0_w_reg[0][13]/P0001  ;
  input \u0_w_reg[0][14]/P0001  ;
  input \u0_w_reg[0][15]/P0001  ;
  input \u0_w_reg[0][16]/P0001  ;
  input \u0_w_reg[0][17]/P0001  ;
  input \u0_w_reg[0][18]/P0001  ;
  input \u0_w_reg[0][19]/P0001  ;
  input \u0_w_reg[0][1]/P0001  ;
  input \u0_w_reg[0][20]/P0001  ;
  input \u0_w_reg[0][21]/P0001  ;
  input \u0_w_reg[0][22]/P0001  ;
  input \u0_w_reg[0][23]/P0001  ;
  input \u0_w_reg[0][24]/P0001  ;
  input \u0_w_reg[0][25]/P0001  ;
  input \u0_w_reg[0][26]/P0001  ;
  input \u0_w_reg[0][27]/P0001  ;
  input \u0_w_reg[0][28]/P0001  ;
  input \u0_w_reg[0][29]/P0001  ;
  input \u0_w_reg[0][2]/P0001  ;
  input \u0_w_reg[0][30]/P0001  ;
  input \u0_w_reg[0][31]/P0001  ;
  input \u0_w_reg[0][3]/P0001  ;
  input \u0_w_reg[0][4]/P0001  ;
  input \u0_w_reg[0][5]/P0001  ;
  input \u0_w_reg[0][6]/P0001  ;
  input \u0_w_reg[0][7]/P0001  ;
  input \u0_w_reg[0][8]/P0001  ;
  input \u0_w_reg[0][9]/P0001  ;
  input \u0_w_reg[1][0]/P0001  ;
  input \u0_w_reg[1][10]/P0001  ;
  input \u0_w_reg[1][11]/P0001  ;
  input \u0_w_reg[1][12]/P0001  ;
  input \u0_w_reg[1][13]/P0001  ;
  input \u0_w_reg[1][14]/P0001  ;
  input \u0_w_reg[1][15]/P0001  ;
  input \u0_w_reg[1][16]/P0001  ;
  input \u0_w_reg[1][17]/P0001  ;
  input \u0_w_reg[1][18]/P0001  ;
  input \u0_w_reg[1][19]/P0001  ;
  input \u0_w_reg[1][1]/P0001  ;
  input \u0_w_reg[1][20]/P0001  ;
  input \u0_w_reg[1][21]/P0001  ;
  input \u0_w_reg[1][22]/P0001  ;
  input \u0_w_reg[1][23]/P0001  ;
  input \u0_w_reg[1][24]/P0002  ;
  input \u0_w_reg[1][25]/P0001  ;
  input \u0_w_reg[1][26]/P0001  ;
  input \u0_w_reg[1][27]/P0001  ;
  input \u0_w_reg[1][28]/P0001  ;
  input \u0_w_reg[1][29]/P0002  ;
  input \u0_w_reg[1][2]/P0001  ;
  input \u0_w_reg[1][30]/P0001  ;
  input \u0_w_reg[1][31]/P0001  ;
  input \u0_w_reg[1][3]/P0001  ;
  input \u0_w_reg[1][4]/P0001  ;
  input \u0_w_reg[1][5]/P0001  ;
  input \u0_w_reg[1][6]/P0001  ;
  input \u0_w_reg[1][7]/P0001  ;
  input \u0_w_reg[1][8]/P0001  ;
  input \u0_w_reg[1][9]/P0001  ;
  input \u0_w_reg[2][0]/P0001  ;
  input \u0_w_reg[2][10]/P0001  ;
  input \u0_w_reg[2][11]/P0001  ;
  input \u0_w_reg[2][12]/P0001  ;
  input \u0_w_reg[2][13]/P0001  ;
  input \u0_w_reg[2][14]/P0001  ;
  input \u0_w_reg[2][15]/P0001  ;
  input \u0_w_reg[2][16]/P0001  ;
  input \u0_w_reg[2][17]/P0001  ;
  input \u0_w_reg[2][18]/P0001  ;
  input \u0_w_reg[2][19]/P0001  ;
  input \u0_w_reg[2][1]/P0001  ;
  input \u0_w_reg[2][20]/P0001  ;
  input \u0_w_reg[2][21]/P0001  ;
  input \u0_w_reg[2][22]/P0001  ;
  input \u0_w_reg[2][23]/P0001  ;
  input \u0_w_reg[2][24]/P0001  ;
  input \u0_w_reg[2][25]/P0001  ;
  input \u0_w_reg[2][26]/P0001  ;
  input \u0_w_reg[2][27]/P0001  ;
  input \u0_w_reg[2][28]/P0001  ;
  input \u0_w_reg[2][29]/P0001  ;
  input \u0_w_reg[2][2]/P0001  ;
  input \u0_w_reg[2][30]/P0001  ;
  input \u0_w_reg[2][31]/P0001  ;
  input \u0_w_reg[2][3]/P0001  ;
  input \u0_w_reg[2][4]/P0001  ;
  input \u0_w_reg[2][5]/P0001  ;
  input \u0_w_reg[2][6]/P0001  ;
  input \u0_w_reg[2][7]/P0001  ;
  input \u0_w_reg[2][8]/P0001  ;
  input \u0_w_reg[2][9]/P0001  ;
  input \u0_w_reg[3][0]/P0001  ;
  input \u0_w_reg[3][10]/P0001  ;
  input \u0_w_reg[3][11]/P0001  ;
  input \u0_w_reg[3][12]/P0001  ;
  input \u0_w_reg[3][13]/P0001  ;
  input \u0_w_reg[3][14]/P0001  ;
  input \u0_w_reg[3][15]/P0001  ;
  input \u0_w_reg[3][16]/P0001  ;
  input \u0_w_reg[3][17]/P0001  ;
  input \u0_w_reg[3][18]/P0001  ;
  input \u0_w_reg[3][19]/P0001  ;
  input \u0_w_reg[3][1]/P0001  ;
  input \u0_w_reg[3][20]/P0001  ;
  input \u0_w_reg[3][21]/P0001  ;
  input \u0_w_reg[3][22]/P0001  ;
  input \u0_w_reg[3][23]/P0001  ;
  input \u0_w_reg[3][24]/P0001  ;
  input \u0_w_reg[3][25]/P0001  ;
  input \u0_w_reg[3][26]/P0001  ;
  input \u0_w_reg[3][27]/P0001  ;
  input \u0_w_reg[3][28]/P0001  ;
  input \u0_w_reg[3][29]/P0001  ;
  input \u0_w_reg[3][2]/P0001  ;
  input \u0_w_reg[3][30]/P0001  ;
  input \u0_w_reg[3][31]/P0001  ;
  input \u0_w_reg[3][3]/P0001  ;
  input \u0_w_reg[3][4]/P0001  ;
  input \u0_w_reg[3][5]/P0001  ;
  input \u0_w_reg[3][6]/P0001  ;
  input \u0_w_reg[3][7]/P0001  ;
  input \u0_w_reg[3][8]/P0001  ;
  input \u0_w_reg[3][9]/P0001  ;
  output \_al_n0  ;
  output \_al_n1  ;
  output \g21/_0_  ;
  output \g56610/_0_  ;
  output \g56611/_0_  ;
  output \g56612/_0_  ;
  output \g56613/_0_  ;
  output \g56614/_0_  ;
  output \g56615/_0_  ;
  output \g56616/_0_  ;
  output \g56617/_0_  ;
  output \g56630/_0_  ;
  output \g56631/_0_  ;
  output \g56632/_0_  ;
  output \g56633/_0_  ;
  output \g56634/_0_  ;
  output \g56635/_0_  ;
  output \g56645/_0_  ;
  output \g56646/_0_  ;
  output \g56647/_0_  ;
  output \g56648/_0_  ;
  output \g56649/_0_  ;
  output \g56650/_0_  ;
  output \g56651/_0_  ;
  output \g56652/_0_  ;
  output \g56666/_0_  ;
  output \g56667/_0_  ;
  output \g56668/_0_  ;
  output \g56669/_0_  ;
  output \g56670/_0_  ;
  output \g56671/_0_  ;
  output \g56672/_0_  ;
  output \g56674/_0_  ;
  output \g56675/_0_  ;
  output \g56704/_0_  ;
  output \g56739/_0_  ;
  output \g56743/_0_  ;
  output \g56763/_0_  ;
  output \g56776/_0_  ;
  output \g56812/_0_  ;
  output \g56818/_0_  ;
  output \g56861/_0_  ;
  output \g56874/_0_  ;
  output \g56919/_0_  ;
  output \g56920/_0_  ;
  output \g56921/_0_  ;
  output \g56923/_0_  ;
  output \g56924/_0_  ;
  output \g56925/_0_  ;
  output \g56926/_0_  ;
  output \g56956/_0_  ;
  output \g56957/_0_  ;
  output \g56958/_0_  ;
  output \g56959/_0_  ;
  output \g56960/_0_  ;
  output \g56961/_0_  ;
  output \g56972/_0_  ;
  output \g56973/_0_  ;
  output \g56974/_0_  ;
  output \g56976/_0_  ;
  output \g56977/_0_  ;
  output \g56978/_0_  ;
  output \g56979/_0_  ;
  output \g56980/_0_  ;
  output \g57008/_0_  ;
  output \g57010/_0_  ;
  output \g57011/_0_  ;
  output \g57012/_0_  ;
  output \g57013/_0_  ;
  output \g57014/_0_  ;
  output \g57015/_0_  ;
  output \g57016/_0_  ;
  output \g57017/_0_  ;
  output \g57086/_0_  ;
  output \g57091/_0_  ;
  output \g57114/_0_  ;
  output \g57129/_0_  ;
  output \g57163/_0_  ;
  output \g57171/_0_  ;
  output \g57204/_0_  ;
  output \g57218/_0_  ;
  output \g57262/_0_  ;
  output \g57263/_0_  ;
  output \g57264/_0_  ;
  output \g57265/_0_  ;
  output \g57266/_0_  ;
  output \g57267/_0_  ;
  output \g57268/_0_  ;
  output \g57269/_0_  ;
  output \g57300/_0_  ;
  output \g57301/_0_  ;
  output \g57302/_0_  ;
  output \g57303/_0_  ;
  output \g57304/_0_  ;
  output \g57316/_0_  ;
  output \g57317/_0_  ;
  output \g57319/_0_  ;
  output \g57320/_0_  ;
  output \g57321/_0_  ;
  output \g57322/_0_  ;
  output \g57323/_0_  ;
  output \g57324/_0_  ;
  output \g57350/_0_  ;
  output \g57353/_0_  ;
  output \g57354/_0_  ;
  output \g57355/_0_  ;
  output \g57356/_0_  ;
  output \g57357/_0_  ;
  output \g57358/_0_  ;
  output \g57359/_0_  ;
  output \g57360/_0_  ;
  output \g57427/_0_  ;
  output \g57432/_0_  ;
  output \g57456/_0_  ;
  output \g57471/_0_  ;
  output \g57506/_0_  ;
  output \g57512/_0_  ;
  output \g57540/_0_  ;
  output \g57547/_0_  ;
  output \g57654/_0_  ;
  output \g57655/_0_  ;
  output \g57656/_0_  ;
  output \g57657/_0_  ;
  output \g57658/_0_  ;
  output \g57676/_0_  ;
  output \g57677/_0_  ;
  output \g57678/_0_  ;
  output \g57679/_0_  ;
  output \g57680/_0_  ;
  output \g57681/_0_  ;
  output \g57682/_0_  ;
  output \g57683/_0_  ;
  output \g57684/_0_  ;
  output \g57685/_0_  ;
  output \g57686/_0_  ;
  output \g57687/_0_  ;
  output \g57688/_0_  ;
  output \g57689/_0_  ;
  output \g57690/_0_  ;
  output \g57691/_0_  ;
  output \g57700/_0_  ;
  output \g57701/_0_  ;
  output \g57702/_0_  ;
  output \g57703/_0_  ;
  output \g57704/_0_  ;
  output \g57705/_0_  ;
  output \g57706/_0_  ;
  output \g57707/_0_  ;
  output \g57708/_0_  ;
  output \g57709/_3_  ;
  output \g57710/_3_  ;
  output \g57711/_0_  ;
  output \g57712/_3_  ;
  output \g57715/_3_  ;
  output \g57716/_3_  ;
  output \g57767/_0_  ;
  output \g57768/_3_  ;
  output \g57769/_3_  ;
  output \g57770/_3_  ;
  output \g57771/_3_  ;
  output \g57777/_3_  ;
  output \g57779/_3_  ;
  output \g57804/_3_  ;
  output \g57805/_3_  ;
  output \g57806/_3_  ;
  output \g57807/_3_  ;
  output \g57808/_3_  ;
  output \g57809/_3_  ;
  output \g57810/_3_  ;
  output \g57811/_3_  ;
  output \g57812/_3_  ;
  output \g57813/_3_  ;
  output \g57814/_3_  ;
  output \g57815/_3_  ;
  output \g57816/_0_  ;
  output \g57817/_3_  ;
  output \g57818/_3_  ;
  output \g57819/_3_  ;
  output \g57822/_3_  ;
  output \g57823/_3_  ;
  output \g57824/_3_  ;
  output \g57830/_3_  ;
  output \g57835/_3_  ;
  output \g57836/_3_  ;
  output \g57837/_3_  ;
  output \g57841/_3_  ;
  output \g57842/_3_  ;
  output \g57843/_3_  ;
  output \g57854/_3_  ;
  output \g57855/_3_  ;
  output \g57856/_3_  ;
  output \g57857/_3_  ;
  output \g57858/_3_  ;
  output \g57859/_3_  ;
  output \g57860/_3_  ;
  output \g57861/_3_  ;
  output \g57871/_3_  ;
  output \g57872/_3_  ;
  output \g57874/_3_  ;
  output \g57968/_3_  ;
  output \g57969/_3_  ;
  output \g57970/_3_  ;
  output \g57971/_3_  ;
  output \g57980/_3_  ;
  output \g57983/_3_  ;
  output \g57984/_3_  ;
  output \g57985/_3_  ;
  output \g58012/_3_  ;
  output \g58013/_3_  ;
  output \g58015/_3_  ;
  output \g58057/_3_  ;
  output \g58058/_3_  ;
  output \g58059/_3_  ;
  output \g58189/_3_  ;
  output \g58190/_3_  ;
  output \g58191/_3_  ;
  output \g58192/_3_  ;
  output \g58193/_3_  ;
  output \g58194/_3_  ;
  output \g58195/_3_  ;
  output \g58196/_3_  ;
  output \g58197/_3_  ;
  output \g58224/_3_  ;
  output \g58226/_3_  ;
  output \g58229/_3_  ;
  output \g58255/_3_  ;
  output \g58256/_3_  ;
  output \g58257/_3_  ;
  output \g58258/_3_  ;
  output \g58259/_3_  ;
  output \g58260/_3_  ;
  output \g58261/_3_  ;
  output \g58262/_3_  ;
  output \g58263/_3_  ;
  output \g58264/_3_  ;
  output \g58265/_3_  ;
  output \g58266/_3_  ;
  output \g58267/_3_  ;
  output \g58268/_3_  ;
  output \g58269/_3_  ;
  output \g58270/_0_  ;
  output \g58271/_3_  ;
  output \g58272/_3_  ;
  output \g58273/_3_  ;
  output \g58274/_3_  ;
  output \g58275/_3_  ;
  output \g58276/_3_  ;
  output \g58277/_3_  ;
  output \g58278/_3_  ;
  output \g58279/_3_  ;
  output \g58285/_3_  ;
  output \g58286/_3_  ;
  output \g58288/_3_  ;
  output \g58289/_3_  ;
  output \g58290/_3_  ;
  output \g58292/_3_  ;
  output \g58294/_3_  ;
  output \g58295/_3_  ;
  output \g58297/_3_  ;
  output \g58330/_0_  ;
  output \g58331/_0_  ;
  output \g58332/_0_  ;
  output \g58333/_0_  ;
  output \g58444/_3_  ;
  output \g58445/_3_  ;
  output \g58446/_3_  ;
  output \g58462/_0_  ;
  output \g58506/_0_  ;
  output \g58507/_0_  ;
  output \g58508/_0_  ;
  output \g58509/_0_  ;
  output \g58531/_0_  ;
  output \g58532/_0_  ;
  output \g58533/_0_  ;
  output \g58550/_0_  ;
  output \g58551/_0_  ;
  output \g58552/_0_  ;
  output \g58553/_0_  ;
  output \g58554/_0_  ;
  output \g58555/_0_  ;
  output \g58556/_0_  ;
  output \g58557/_0_  ;
  output \g58558/_0_  ;
  output \g58559/_0_  ;
  output \g58560/_0_  ;
  output \g58600/_3_  ;
  output \g58601/_3_  ;
  output \g58602/_3_  ;
  output \g58603/_3_  ;
  output \g58604/_3_  ;
  output \g58605/_3_  ;
  output \g58606/_3_  ;
  output \g58607/_3_  ;
  output \g58608/_3_  ;
  output \g58611/_0_  ;
  output \g58612/_0_  ;
  output \g58613/_0_  ;
  output \g58614/_0_  ;
  output \g58617/_0_  ;
  output \g58618/_0_  ;
  output \g58619/_0_  ;
  output \g58634/_0_  ;
  output \g58635/_0_  ;
  output \g58636/_0_  ;
  output \g58637/_0_  ;
  output \g58638/_0_  ;
  output \g58639/_0_  ;
  output \g58640/_0_  ;
  output \g58641/_0_  ;
  output \g58829/_3_  ;
  output \g58830/_3_  ;
  output \g58831/_3_  ;
  output \g58832/_3_  ;
  output \g58833/_3_  ;
  output \g58834/_3_  ;
  output \g58835/_0_  ;
  output \g58844/_0_  ;
  output \g58902/_0_  ;
  output \g58903/_0_  ;
  output \g58904/_0_  ;
  output \g58905/_0_  ;
  output \g58910/_0_  ;
  output \g58913/_0_  ;
  output \g58934/_0_  ;
  output \g58935/_0_  ;
  output \g58936/_0_  ;
  output \g58937/_0_  ;
  output \g58938/_0_  ;
  output \g58970/_0_  ;
  output \g58972/_0_  ;
  output \g58994/_0_  ;
  output \g58995/_0_  ;
  output \g58996/_0_  ;
  output \g58997/_0_  ;
  output \g58998/_0_  ;
  output \g58999/_0_  ;
  output \g59000/_0_  ;
  output \g59002/_0_  ;
  output \g59003/_0_  ;
  output \g59004/_0_  ;
  output \g59254/_0_  ;
  output \g59257/_0_  ;
  output \g59258/_0_  ;
  output \g59259/_0_  ;
  output \g59276/_0_  ;
  output \g59277/_0_  ;
  output \g59278/_0_  ;
  output \g59279/_0_  ;
  output \g59280/_0_  ;
  output \g59291/_0_  ;
  output \g59292/_0_  ;
  output \g59293/_0_  ;
  output \g59294/_0_  ;
  output \g59295/_0_  ;
  output \g59308/_0_  ;
  output \g59309/_0_  ;
  output \g59310/_0_  ;
  output \g59311/_0_  ;
  output \g59330/_0_  ;
  output \g59331/_0_  ;
  output \g59332/_0_  ;
  output \g59333/_0_  ;
  output \g59334/_0_  ;
  output \g59335/_0_  ;
  output \g59336/_0_  ;
  output \g59337/_0_  ;
  output \g59338/_0_  ;
  output \g59339/_0_  ;
  output \g59596/_0_  ;
  output \g59597/_0_  ;
  output \g59598/_0_  ;
  output \g59599/_0_  ;
  output \g59625/_0_  ;
  output \g59626/_0_  ;
  output \g59627/_0_  ;
  output \g59628/_0_  ;
  output \g59837/_0_  ;
  output \g59838/_0_  ;
  output \g59839/_0_  ;
  output \g59840/_0_  ;
  output \g60090/_0_  ;
  output \g60320/_0_  ;
  output \g60321/_0_  ;
  output \g60409/_0_  ;
  output \g60539/_0_  ;
  output \g60860/_0_  ;
  output \g60977/_0_  ;
  output \g61012/_0_  ;
  output \g61185/_0_  ;
  output \g61524/_2_  ;
  output \g61776/_0_  ;
  output \g61895/_0_  ;
  output \g61897/_0_  ;
  output \g62220/_0_  ;
  output \g65958/_0_  ;
  output \g72347/_3_  ;
  output \g77848/_0_  ;
  output \g85056/_0_  ;
  output \sa30_reg[0]/_05_  ;
  output \sa31_reg[0]/_05_  ;
  output \sa32_reg[0]/_05_  ;
  output \u0_w_reg[1][24]/_05_  ;
  output \u0_w_reg[1][29]/_05_  ;
  wire n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , n6000 , n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , n6089 , n6090 , n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , n6170 , n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , n6230 , n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , n6240 , n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , n6250 , n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , n6259 , n6260 , n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , n6300 , n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , n6310 , n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , n6320 , n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , n6340 , n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , n6349 , n6350 , n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , n6359 , n6360 , n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , n6367 , n6368 , n6369 , n6370 , n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , n6380 , n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , n6390 , n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , n6400 , n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , n6409 , n6410 , n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , n6420 , n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , n6429 , n6430 , n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , n6439 , n6440 , n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , n6449 , n6450 , n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , n6460 , n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , n6470 , n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , n6480 , n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , n6490 , n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , n6499 , n6500 , n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , n6509 , n6510 , n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , n6519 , n6520 , n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , n6529 , n6530 , n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , n6539 , n6540 , n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , n6549 , n6550 , n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , n6559 , n6560 , n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , n6569 , n6570 , n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , n6579 , n6580 , n6581 , n6582 , n6583 , n6584 , n6585 , n6586 , n6587 , n6588 , n6589 , n6590 , n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , n6599 , n6600 , n6601 , n6602 , n6603 , n6604 , n6605 , n6606 , n6607 , n6608 , n6609 , n6610 , n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , n6617 , n6618 , n6619 , n6620 , n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , n6627 , n6628 , n6629 , n6630 , n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , n6639 , n6640 , n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , n6647 , n6648 , n6649 , n6650 , n6651 , n6652 , n6653 , n6654 , n6655 , n6656 , n6657 , n6658 , n6659 , n6660 , n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , n6667 , n6668 , n6669 , n6670 , n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , n6679 , n6680 , n6681 , n6682 , n6683 , n6684 , n6685 , n6686 , n6687 , n6688 , n6689 , n6690 , n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , n6697 , n6698 , n6699 , n6700 , n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , n6707 , n6708 , n6709 , n6710 , n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , n6717 , n6718 , n6719 , n6720 , n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , n6729 , n6730 , n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , n6739 , n6740 , n6741 , n6742 , n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , n6749 , n6750 , n6751 , n6752 , n6753 , n6754 , n6755 , n6756 , n6757 , n6758 , n6759 , n6760 , n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , n6770 , n6771 , n6772 , n6773 , n6774 , n6775 , n6776 , n6777 , n6778 , n6779 , n6780 , n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , n6789 , n6790 , n6791 , n6792 , n6793 , n6794 , n6795 , n6796 , n6797 , n6798 , n6799 , n6800 , n6801 , n6802 , n6803 , n6804 , n6805 , n6806 , n6807 , n6808 , n6809 , n6810 , n6811 , n6812 , n6813 , n6814 , n6815 , n6816 , n6817 , n6818 , n6819 , n6820 , n6821 , n6822 , n6823 , n6824 , n6825 , n6826 , n6827 , n6828 , n6829 , n6830 , n6831 , n6832 , n6833 , n6834 , n6835 , n6836 , n6837 , n6838 , n6839 , n6840 , n6841 , n6842 , n6843 , n6844 , n6845 , n6846 , n6847 , n6848 , n6849 , n6850 , n6851 , n6852 , n6853 , n6854 , n6855 , n6856 , n6857 , n6858 , n6859 , n6860 , n6861 , n6862 , n6863 , n6864 , n6865 , n6866 , n6867 , n6868 , n6869 , n6870 , n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , n6877 , n6878 , n6879 , n6880 , n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , n6887 , n6888 , n6889 , n6890 , n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , n6897 , n6898 , n6899 , n6900 , n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , n6907 , n6908 , n6909 , n6910 , n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , n6919 , n6920 , n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , n6927 , n6928 , n6929 , n6930 , n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , n6937 , n6938 , n6939 , n6940 , n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , n6949 , n6950 , n6951 , n6952 , n6953 , n6954 , n6955 , n6956 , n6957 , n6958 , n6959 , n6960 , n6961 , n6962 , n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , n6969 , n6970 , n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , n6979 , n6980 , n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , n6987 , n6988 , n6989 , n6990 , n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , n6997 , n6998 , n6999 , n7000 , n7001 , n7002 , n7003 , n7004 , n7005 , n7006 , n7007 , n7008 , n7009 , n7010 , n7011 , n7012 , n7013 , n7014 , n7015 , n7016 , n7017 , n7018 , n7019 , n7020 , n7021 , n7022 , n7023 , n7024 , n7025 , n7026 , n7027 , n7028 , n7029 , n7030 , n7031 , n7032 , n7033 , n7034 , n7035 , n7036 , n7037 , n7038 , n7039 , n7040 , n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , n7047 , n7048 , n7049 , n7050 , n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , n7057 , n7058 , n7059 , n7060 , n7061 , n7062 , n7063 , n7064 , n7065 , n7066 , n7067 , n7068 , n7069 , n7070 , n7071 , n7072 , n7073 , n7074 , n7075 , n7076 , n7077 , n7078 , n7079 , n7080 , n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , n7087 , n7088 , n7089 , n7090 , n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , n7097 , n7098 , n7099 , n7100 , n7101 , n7102 , n7103 , n7104 , n7105 , n7106 , n7107 , n7108 , n7109 , n7110 , n7111 , n7112 , n7113 , n7114 , n7115 , n7116 , n7117 , n7118 , n7119 , n7120 , n7121 , n7122 , n7123 , n7124 , n7125 , n7126 , n7127 , n7128 , n7129 , n7130 , n7131 , n7132 , n7133 , n7134 , n7135 , n7136 , n7137 , n7138 , n7139 , n7140 , n7141 , n7142 , n7143 , n7144 , n7145 , n7146 , n7147 , n7148 , n7149 , n7150 , n7151 , n7152 , n7153 , n7154 , n7155 , n7156 , n7157 , n7158 , n7159 , n7160 , n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , n7167 , n7168 , n7169 , n7170 , n7171 , n7172 , n7173 , n7174 , n7175 , n7176 , n7177 , n7178 , n7179 , n7180 , n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , n7187 , n7188 , n7189 , n7190 , n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , n7197 , n7198 , n7199 , n7200 , n7201 , n7202 , n7203 , n7204 , n7205 , n7206 , n7207 , n7208 , n7209 , n7210 , n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , n7217 , n7218 , n7219 , n7220 , n7221 , n7222 , n7223 , n7224 , n7225 , n7226 , n7227 , n7228 , n7229 , n7230 , n7231 , n7232 , n7233 , n7234 , n7235 , n7236 , n7237 , n7238 , n7239 , n7240 , n7241 , n7242 , n7243 , n7244 , n7245 , n7246 , n7247 , n7248 , n7249 , n7250 , n7251 , n7252 , n7253 , n7254 , n7255 , n7256 , n7257 , n7258 , n7259 , n7260 , n7261 , n7262 , n7263 , n7264 , n7265 , n7266 , n7267 , n7268 , n7269 , n7270 , n7271 , n7272 , n7273 , n7274 , n7275 , n7276 , n7277 , n7278 , n7279 , n7280 , n7281 , n7282 , n7283 , n7284 , n7285 , n7286 , n7287 , n7288 , n7289 , n7290 , n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , n7297 , n7298 , n7299 , n7300 , n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , n7307 , n7308 , n7309 , n7310 , n7311 , n7312 , n7313 , n7314 , n7315 , n7316 , n7317 , n7318 , n7319 , n7320 , n7321 , n7322 , n7323 , n7324 , n7325 , n7326 , n7327 , n7328 , n7329 , n7330 , n7331 , n7332 , n7333 , n7334 , n7335 , n7336 , n7337 , n7338 , n7339 , n7340 , n7341 , n7342 , n7343 , n7344 , n7345 , n7346 , n7347 , n7348 , n7349 , n7350 , n7351 , n7352 , n7353 , n7354 , n7355 , n7356 , n7357 , n7358 , n7359 , n7360 , n7361 , n7362 , n7363 , n7364 , n7365 , n7366 , n7367 , n7368 , n7369 , n7370 , n7371 , n7372 , n7373 , n7374 , n7375 , n7376 , n7377 , n7378 , n7379 , n7380 , n7381 , n7382 , n7383 , n7384 , n7385 , n7386 , n7387 , n7388 , n7389 , n7390 , n7391 , n7392 , n7393 , n7394 , n7395 , n7396 , n7397 , n7398 , n7399 , n7400 , n7401 , n7402 , n7403 , n7404 , n7405 , n7406 , n7407 , n7408 , n7409 , n7410 , n7411 , n7412 , n7413 , n7414 , n7415 , n7416 , n7417 , n7418 , n7419 , n7420 , n7421 , n7422 , n7423 , n7424 , n7425 , n7426 , n7427 , n7428 , n7429 , n7430 , n7431 , n7432 , n7433 , n7434 , n7435 , n7436 , n7437 , n7438 , n7439 , n7440 , n7441 , n7442 , n7443 , n7444 , n7445 , n7446 , n7447 , n7448 , n7449 , n7450 , n7451 , n7452 , n7453 , n7454 , n7455 , n7456 , n7457 , n7458 , n7459 , n7460 , n7461 , n7462 , n7463 , n7464 , n7465 , n7466 , n7467 , n7468 , n7469 , n7470 , n7471 , n7472 , n7473 , n7474 , n7475 , n7476 , n7477 , n7478 , n7479 , n7480 , n7481 , n7482 , n7483 , n7484 , n7485 , n7486 , n7487 , n7488 , n7489 , n7490 , n7491 , n7492 , n7493 , n7494 , n7495 , n7496 , n7497 , n7498 , n7499 , n7500 , n7501 , n7502 , n7503 , n7504 , n7505 , n7506 , n7507 , n7508 , n7509 , n7510 , n7511 , n7512 , n7513 , n7514 , n7515 , n7516 , n7517 , n7518 , n7519 , n7520 , n7521 , n7522 , n7523 , n7524 , n7525 , n7526 , n7527 , n7528 , n7529 , n7530 , n7531 , n7532 , n7533 , n7534 , n7535 , n7536 , n7537 , n7538 , n7539 , n7540 , n7541 , n7542 , n7543 , n7544 , n7545 , n7546 , n7547 , n7548 , n7549 , n7550 , n7551 , n7552 , n7553 , n7554 , n7555 , n7556 , n7557 , n7558 , n7559 , n7560 , n7561 , n7562 , n7563 , n7564 , n7565 , n7566 , n7567 , n7568 , n7569 , n7570 , n7571 , n7572 , n7573 , n7574 , n7575 , n7576 , n7577 , n7578 , n7579 , n7580 , n7581 , n7582 , n7583 , n7584 , n7585 , n7586 , n7587 , n7588 , n7589 , n7590 , n7591 , n7592 , n7593 , n7594 , n7595 , n7596 , n7597 , n7598 , n7599 , n7600 , n7601 , n7602 , n7603 , n7604 , n7605 , n7606 , n7607 , n7608 , n7609 , n7610 , n7611 , n7612 , n7613 , n7614 , n7615 , n7616 , n7617 , n7618 , n7619 , n7620 , n7621 , n7622 , n7623 , n7624 , n7625 , n7626 , n7627 , n7628 , n7629 , n7630 , n7631 , n7632 , n7633 , n7634 , n7635 , n7636 , n7637 , n7638 , n7639 , n7640 , n7641 , n7642 , n7643 , n7644 , n7645 , n7646 , n7647 , n7648 , n7649 , n7650 , n7651 , n7652 , n7653 , n7654 , n7655 , n7656 , n7657 , n7658 , n7659 , n7660 , n7661 , n7662 , n7663 , n7664 , n7665 , n7666 , n7667 , n7668 , n7669 , n7670 , n7671 , n7672 , n7673 , n7674 , n7675 , n7676 , n7677 , n7678 , n7679 , n7680 , n7681 , n7682 , n7683 , n7684 , n7685 , n7686 , n7687 , n7688 , n7689 , n7690 , n7691 , n7692 , n7693 , n7694 , n7695 , n7696 , n7697 , n7698 , n7699 , n7700 , n7701 , n7702 , n7703 , n7704 , n7705 , n7706 , n7707 , n7708 , n7709 , n7710 , n7711 , n7712 , n7713 , n7714 , n7715 , n7716 , n7717 , n7718 , n7719 , n7720 , n7721 , n7722 , n7723 , n7724 , n7725 , n7726 , n7727 , n7728 , n7729 , n7730 , n7731 , n7732 , n7733 , n7734 , n7735 , n7736 , n7737 , n7738 , n7739 , n7740 , n7741 , n7742 , n7743 , n7744 , n7745 , n7746 , n7747 , n7748 , n7749 , n7750 , n7751 , n7752 , n7753 , n7754 , n7755 , n7756 , n7757 , n7758 , n7759 , n7760 , n7761 , n7762 , n7763 , n7764 , n7765 , n7766 , n7767 , n7768 , n7769 , n7770 , n7771 , n7772 , n7773 , n7774 , n7775 , n7776 , n7777 , n7778 , n7779 , n7780 , n7781 , n7782 , n7783 , n7784 , n7785 , n7786 , n7787 , n7788 , n7789 , n7790 , n7791 , n7792 , n7793 , n7794 , n7795 , n7796 , n7797 , n7798 , n7799 , n7800 , n7801 , n7802 , n7803 , n7804 , n7805 , n7806 , n7807 , n7808 , n7809 , n7810 , n7811 , n7812 , n7813 , n7814 , n7815 , n7816 , n7817 , n7818 , n7819 , n7820 , n7821 , n7822 , n7823 , n7824 , n7825 , n7826 , n7827 , n7828 , n7829 , n7830 , n7831 , n7832 , n7833 , n7834 , n7835 , n7836 , n7837 , n7838 , n7839 , n7840 , n7841 , n7842 , n7843 , n7844 , n7845 , n7846 , n7847 , n7848 , n7849 , n7850 , n7851 , n7852 , n7853 , n7854 , n7855 , n7856 , n7857 , n7858 , n7859 , n7860 , n7861 , n7862 , n7863 , n7864 , n7865 , n7866 , n7867 , n7868 , n7869 , n7870 , n7871 , n7872 , n7873 , n7874 , n7875 , n7876 , n7877 , n7878 , n7879 , n7880 , n7881 , n7882 , n7883 , n7884 , n7885 , n7886 , n7887 , n7888 , n7889 , n7890 , n7891 , n7892 , n7893 , n7894 , n7895 , n7896 , n7897 , n7898 , n7899 , n7900 , n7901 , n7902 , n7903 , n7904 , n7905 , n7906 , n7907 , n7908 , n7909 , n7910 , n7911 , n7912 , n7913 , n7914 , n7915 , n7916 , n7917 , n7918 , n7919 , n7920 , n7921 , n7922 , n7923 , n7924 , n7925 , n7926 , n7927 , n7928 , n7929 , n7930 , n7931 , n7932 , n7933 , n7934 , n7935 , n7936 , n7937 , n7938 , n7939 , n7940 , n7941 , n7942 , n7943 , n7944 , n7945 , n7946 , n7947 , n7948 , n7949 , n7950 , n7951 , n7952 , n7953 , n7954 , n7955 , n7956 , n7957 , n7958 , n7959 , n7960 , n7961 , n7962 , n7963 , n7964 , n7965 , n7966 , n7967 , n7968 , n7969 , n7970 , n7971 , n7972 , n7973 , n7974 , n7975 , n7976 , n7977 , n7978 , n7979 , n7980 , n7981 , n7982 , n7983 , n7984 , n7985 , n7986 , n7987 , n7988 , n7989 , n7990 , n7991 , n7992 , n7993 , n7994 , n7995 , n7996 , n7997 , n7998 , n7999 , n8000 , n8001 , n8002 , n8003 , n8004 , n8005 , n8006 , n8007 , n8008 , n8009 , n8010 , n8011 , n8012 , n8013 , n8014 , n8015 , n8016 , n8017 , n8018 , n8019 , n8020 , n8021 , n8022 , n8023 , n8024 , n8025 , n8026 , n8027 , n8028 , n8029 , n8030 , n8031 , n8032 , n8033 , n8034 , n8035 , n8036 , n8037 , n8038 , n8039 , n8040 , n8041 , n8042 , n8043 , n8044 , n8045 , n8046 , n8047 , n8048 , n8049 , n8050 , n8051 , n8052 , n8053 , n8054 , n8055 , n8056 , n8057 , n8058 , n8059 , n8060 , n8061 , n8062 , n8063 , n8064 , n8065 , n8066 , n8067 , n8068 , n8069 , n8070 , n8071 , n8072 , n8073 , n8074 , n8075 , n8076 , n8077 , n8078 , n8079 , n8080 , n8081 , n8082 , n8083 , n8084 , n8085 , n8086 , n8087 , n8088 , n8089 , n8090 , n8091 , n8092 , n8093 , n8094 , n8095 , n8096 , n8097 , n8098 , n8099 , n8100 , n8101 , n8102 , n8103 , n8104 , n8105 , n8106 , n8107 , n8108 , n8109 , n8110 , n8111 , n8112 , n8113 , n8114 , n8115 , n8116 , n8117 , n8118 , n8119 , n8120 , n8121 , n8122 , n8123 , n8124 , n8125 , n8126 , n8127 , n8128 , n8129 , n8130 , n8131 , n8132 , n8133 , n8134 , n8135 , n8136 , n8137 , n8138 , n8139 , n8140 , n8141 , n8142 , n8143 , n8144 , n8145 , n8146 , n8147 , n8148 , n8149 , n8150 , n8151 , n8152 , n8153 , n8154 , n8155 , n8156 , n8157 , n8158 , n8159 , n8160 , n8161 , n8162 , n8163 , n8164 , n8165 , n8166 , n8167 , n8168 , n8169 , n8170 , n8171 , n8172 , n8173 , n8174 , n8175 , n8176 , n8177 , n8178 , n8179 , n8180 , n8181 , n8182 , n8183 , n8184 , n8185 , n8186 , n8187 , n8188 , n8189 , n8190 , n8191 , n8192 , n8193 , n8194 , n8195 , n8196 , n8197 , n8198 , n8199 , n8200 , n8201 , n8202 , n8203 , n8204 , n8205 , n8206 , n8207 , n8208 , n8209 , n8210 , n8211 , n8212 , n8213 , n8214 , n8215 , n8216 , n8217 , n8218 , n8219 , n8220 , n8221 , n8222 , n8223 , n8224 , n8225 , n8226 , n8227 , n8228 , n8229 , n8230 , n8231 , n8232 , n8233 , n8234 , n8235 , n8236 , n8237 , n8238 , n8239 , n8240 , n8241 , n8242 , n8243 , n8244 , n8245 , n8246 , n8247 , n8248 , n8249 , n8250 , n8251 , n8252 , n8253 , n8254 , n8255 , n8256 , n8257 , n8258 , n8259 , n8260 , n8261 , n8262 , n8263 , n8264 , n8265 , n8266 , n8267 , n8268 , n8269 , n8270 , n8271 , n8272 , n8273 , n8274 , n8275 , n8276 , n8277 , n8278 , n8279 , n8280 , n8281 , n8282 , n8283 , n8284 , n8285 , n8286 , n8287 , n8288 , n8289 , n8290 , n8291 , n8292 , n8293 , n8294 , n8295 , n8296 , n8297 , n8298 , n8299 , n8300 , n8301 , n8302 , n8303 , n8304 , n8305 , n8306 , n8307 , n8308 , n8309 , n8310 , n8311 , n8312 , n8313 , n8314 , n8315 , n8316 , n8317 , n8318 , n8319 , n8320 , n8321 , n8322 , n8323 , n8324 , n8325 , n8326 , n8327 , n8328 , n8329 , n8330 , n8331 , n8332 , n8333 , n8334 , n8335 , n8336 , n8337 , n8338 , n8339 , n8340 , n8341 , n8342 , n8343 , n8344 , n8345 , n8346 , n8347 , n8348 , n8349 , n8350 , n8351 , n8352 , n8353 , n8354 , n8355 , n8356 , n8357 , n8358 , n8359 , n8360 , n8361 , n8362 , n8363 , n8364 , n8365 , n8366 , n8367 , n8368 , n8369 , n8370 , n8371 , n8372 , n8373 , n8374 , n8375 , n8376 , n8377 , n8378 , n8379 , n8380 , n8381 , n8382 , n8383 , n8384 , n8385 , n8386 , n8387 , n8388 , n8389 , n8390 , n8391 , n8392 , n8393 , n8394 , n8395 , n8396 , n8397 , n8398 , n8399 , n8400 , n8401 , n8402 , n8403 , n8404 , n8405 , n8406 , n8407 , n8408 , n8409 , n8410 , n8411 , n8412 , n8413 , n8414 , n8415 , n8416 , n8417 , n8418 , n8419 , n8420 , n8421 , n8422 , n8423 , n8424 , n8425 , n8426 , n8427 , n8428 , n8429 , n8430 , n8431 , n8432 , n8433 , n8434 , n8435 , n8436 , n8437 , n8438 , n8439 , n8440 , n8441 , n8442 , n8443 , n8444 , n8445 , n8446 , n8447 , n8448 , n8449 , n8450 , n8451 , n8452 , n8453 , n8454 , n8455 , n8456 , n8457 , n8458 , n8459 , n8460 , n8461 , n8462 , n8463 , n8464 , n8465 , n8466 , n8467 , n8468 , n8469 , n8470 , n8471 , n8472 , n8473 , n8474 , n8475 , n8476 , n8477 , n8478 , n8479 , n8480 , n8481 , n8482 , n8483 , n8484 , n8485 , n8486 , n8487 , n8488 , n8489 , n8490 , n8491 , n8492 , n8493 , n8494 , n8495 , n8496 , n8497 , n8498 , n8499 , n8500 , n8501 , n8502 , n8503 , n8504 , n8505 , n8506 , n8507 , n8508 , n8509 , n8510 , n8511 , n8512 , n8513 , n8514 , n8515 , n8516 , n8517 , n8518 , n8519 , n8520 , n8521 , n8522 , n8523 , n8524 , n8525 , n8526 , n8527 , n8528 , n8529 , n8530 , n8531 , n8532 , n8533 , n8534 , n8535 , n8536 , n8537 , n8538 , n8539 , n8540 , n8541 , n8542 , n8543 , n8544 , n8545 , n8546 , n8547 , n8548 , n8549 , n8550 , n8551 , n8552 , n8553 , n8554 , n8555 , n8556 , n8557 , n8558 , n8559 , n8560 , n8561 , n8562 , n8563 , n8564 , n8565 , n8566 , n8567 , n8568 , n8569 , n8570 , n8571 , n8572 , n8573 , n8574 , n8575 , n8576 , n8577 , n8578 , n8579 , n8580 , n8581 , n8582 , n8583 , n8584 , n8585 , n8586 , n8587 , n8588 , n8589 , n8590 , n8591 , n8592 , n8593 , n8594 , n8595 , n8596 , n8597 , n8598 , n8599 , n8600 , n8601 , n8602 , n8603 , n8604 , n8605 , n8606 , n8607 , n8608 , n8609 , n8610 , n8611 , n8612 , n8613 , n8614 , n8615 , n8616 , n8617 , n8618 , n8619 , n8620 , n8621 , n8622 , n8623 , n8624 , n8625 , n8626 , n8627 , n8628 , n8629 , n8630 , n8631 , n8632 , n8633 , n8634 , n8635 , n8636 , n8637 , n8638 , n8639 , n8640 , n8641 , n8642 , n8643 , n8644 , n8645 , n8646 , n8647 , n8648 , n8649 , n8650 , n8651 , n8652 , n8653 , n8654 , n8655 , n8656 , n8657 , n8658 , n8659 , n8660 , n8661 , n8662 , n8663 , n8664 , n8665 , n8666 , n8667 , n8668 , n8669 , n8670 , n8671 , n8672 , n8673 , n8674 , n8675 , n8676 , n8677 , n8678 , n8679 , n8680 , n8681 , n8682 , n8683 , n8684 , n8685 , n8686 , n8687 , n8688 , n8689 , n8690 , n8691 , n8692 , n8693 , n8694 , n8695 , n8696 , n8697 , n8698 , n8699 , n8700 , n8701 , n8702 , n8703 , n8704 , n8705 , n8706 , n8707 , n8708 , n8709 , n8710 , n8711 , n8712 , n8713 , n8714 , n8715 , n8716 , n8717 , n8718 , n8719 , n8720 , n8721 , n8722 , n8723 , n8724 , n8725 , n8726 , n8727 , n8728 , n8729 , n8730 , n8731 , n8732 , n8733 , n8734 , n8735 , n8736 , n8737 , n8738 , n8739 , n8740 , n8741 , n8742 , n8743 , n8744 , n8745 , n8746 , n8747 , n8748 , n8749 , n8750 , n8751 , n8752 , n8753 , n8754 , n8755 , n8756 , n8757 , n8758 , n8759 , n8760 , n8761 , n8762 , n8763 , n8764 , n8765 , n8766 , n8767 , n8768 , n8769 , n8770 , n8771 , n8772 , n8773 , n8774 , n8775 , n8776 , n8777 , n8778 , n8779 , n8780 , n8781 , n8782 , n8783 , n8784 , n8785 , n8786 , n8787 , n8788 , n8789 , n8790 , n8791 , n8792 , n8793 , n8794 , n8795 , n8796 , n8797 , n8798 , n8799 , n8800 , n8801 , n8802 , n8803 , n8804 , n8805 , n8806 , n8807 , n8808 , n8809 , n8810 , n8811 , n8812 , n8813 , n8814 , n8815 , n8816 , n8817 , n8818 , n8819 , n8820 , n8821 , n8822 , n8823 , n8824 , n8825 , n8826 , n8827 , n8828 , n8829 , n8830 , n8831 , n8832 , n8833 , n8834 , n8835 , n8836 , n8837 , n8838 , n8839 , n8840 , n8841 , n8842 , n8843 , n8844 , n8845 , n8846 , n8847 , n8848 , n8849 , n8850 , n8851 , n8852 , n8853 , n8854 , n8855 , n8856 , n8857 , n8858 , n8859 , n8860 , n8861 , n8862 , n8863 , n8864 , n8865 , n8866 , n8867 , n8868 , n8869 , n8870 , n8871 , n8872 , n8873 , n8874 , n8875 , n8876 , n8877 , n8878 , n8879 , n8880 , n8881 , n8882 , n8883 , n8884 , n8885 , n8886 , n8887 , n8888 , n8889 , n8890 , n8891 , n8892 , n8893 , n8894 , n8895 , n8896 , n8897 , n8898 , n8899 , n8900 , n8901 , n8902 , n8903 , n8904 , n8905 , n8906 , n8907 , n8908 , n8909 , n8910 , n8911 , n8912 , n8913 , n8914 , n8915 , n8916 , n8917 , n8918 , n8919 , n8920 , n8921 , n8922 , n8923 , n8924 , n8925 , n8926 , n8927 , n8928 , n8929 , n8930 , n8931 , n8932 , n8933 , n8934 , n8935 , n8936 , n8937 , n8938 , n8939 , n8940 , n8941 , n8942 , n8943 , n8944 , n8945 , n8946 , n8947 , n8948 , n8949 , n8950 , n8951 , n8952 , n8953 , n8954 , n8955 , n8956 , n8957 , n8958 , n8959 , n8960 , n8961 , n8962 , n8963 , n8964 , n8965 , n8966 , n8967 , n8968 , n8969 , n8970 , n8971 , n8972 , n8973 , n8974 , n8975 , n8976 , n8977 , n8978 , n8979 , n8980 , n8981 , n8982 , n8983 , n8984 , n8985 , n8986 , n8987 , n8988 , n8989 , n8990 , n8991 , n8992 , n8993 , n8994 , n8995 , n8996 , n8997 , n8998 , n8999 , n9000 , n9001 , n9002 , n9003 , n9004 , n9005 , n9006 , n9007 , n9008 , n9009 , n9010 , n9011 , n9012 , n9013 , n9014 , n9015 , n9016 , n9017 , n9018 , n9019 , n9020 , n9021 , n9022 , n9023 , n9024 , n9025 , n9026 , n9027 , n9028 , n9029 , n9030 , n9031 , n9032 , n9033 , n9034 , n9035 , n9036 , n9037 , n9038 , n9039 , n9040 , n9041 , n9042 , n9043 , n9044 , n9045 , n9046 , n9047 , n9048 , n9049 , n9050 , n9051 , n9052 , n9053 , n9054 , n9055 , n9056 , n9057 , n9058 , n9059 , n9060 , n9061 , n9062 , n9063 , n9064 , n9065 , n9066 , n9067 , n9068 , n9069 , n9070 , n9071 , n9072 , n9073 , n9074 , n9075 , n9076 , n9077 , n9078 , n9079 , n9080 , n9081 , n9082 , n9083 , n9084 , n9085 , n9086 , n9087 , n9088 , n9089 , n9090 , n9091 , n9092 , n9093 , n9094 , n9095 , n9096 , n9097 , n9098 , n9099 , n9100 , n9101 , n9102 , n9103 , n9104 , n9105 , n9106 , n9107 , n9108 , n9109 , n9110 , n9111 , n9112 , n9113 , n9114 , n9115 , n9116 , n9117 , n9118 , n9119 , n9120 , n9121 , n9122 , n9123 , n9124 , n9125 , n9126 , n9127 , n9128 , n9129 , n9130 , n9131 , n9132 , n9133 , n9134 , n9135 , n9136 , n9137 , n9138 , n9139 , n9140 , n9141 , n9142 , n9143 , n9144 , n9145 , n9146 , n9147 , n9148 , n9149 , n9150 , n9151 , n9152 , n9153 , n9154 , n9155 , n9156 , n9157 , n9158 , n9159 , n9160 , n9161 , n9162 , n9163 , n9164 , n9165 , n9166 , n9167 , n9168 , n9169 , n9170 , n9171 , n9172 , n9173 , n9174 , n9175 , n9176 , n9177 , n9178 , n9179 , n9180 , n9181 , n9182 , n9183 , n9184 , n9185 , n9186 , n9187 , n9188 , n9189 , n9190 , n9191 , n9192 , n9193 , n9194 , n9195 , n9196 , n9197 , n9198 , n9199 , n9200 , n9201 , n9202 , n9203 , n9204 , n9205 , n9206 , n9207 , n9208 , n9209 , n9210 , n9211 , n9212 , n9213 , n9214 , n9215 , n9216 , n9217 , n9218 , n9219 , n9220 , n9221 , n9222 , n9223 , n9224 , n9225 , n9226 , n9227 , n9228 , n9229 , n9230 , n9231 , n9232 , n9233 , n9234 , n9235 , n9236 , n9237 , n9238 , n9239 , n9240 , n9241 , n9242 , n9243 , n9244 , n9245 , n9246 , n9247 , n9248 , n9249 , n9250 , n9251 , n9252 , n9253 , n9254 , n9255 , n9256 , n9257 , n9258 , n9259 , n9260 , n9261 , n9262 , n9263 , n9264 , n9265 , n9266 , n9267 , n9268 , n9269 , n9270 , n9271 , n9272 , n9273 , n9274 , n9275 , n9276 , n9277 , n9278 , n9279 , n9280 , n9281 , n9282 , n9283 , n9284 , n9285 , n9286 , n9287 , n9288 , n9289 , n9290 , n9291 , n9292 , n9293 , n9294 , n9295 , n9296 , n9297 , n9298 , n9299 , n9300 , n9301 , n9302 , n9303 , n9304 , n9305 , n9306 , n9307 , n9308 , n9309 , n9310 , n9311 , n9312 , n9313 , n9314 , n9315 , n9316 , n9317 , n9318 , n9319 , n9320 , n9321 , n9322 , n9323 , n9324 , n9325 , n9326 , n9327 , n9328 , n9329 , n9330 , n9331 , n9332 , n9333 , n9334 , n9335 , n9336 , n9337 , n9338 , n9339 , n9340 , n9341 , n9342 , n9343 , n9344 , n9345 , n9346 , n9347 , n9348 , n9349 , n9350 , n9351 , n9352 , n9353 , n9354 , n9355 , n9356 , n9357 , n9358 , n9359 , n9360 , n9361 , n9362 , n9363 , n9364 , n9365 , n9366 , n9367 , n9368 , n9369 , n9370 , n9371 , n9372 , n9373 , n9374 , n9375 , n9376 , n9377 , n9378 , n9379 , n9380 , n9381 , n9382 , n9383 , n9384 , n9385 , n9386 , n9387 , n9388 , n9389 , n9390 , n9391 , n9392 , n9393 , n9394 , n9395 , n9396 , n9397 , n9398 , n9399 , n9400 , n9401 , n9402 , n9403 , n9404 , n9405 , n9406 , n9407 , n9408 , n9409 , n9410 , n9411 , n9412 , n9413 , n9414 , n9415 , n9416 , n9417 , n9418 , n9419 , n9420 , n9421 , n9422 , n9423 , n9424 , n9425 , n9426 , n9427 , n9428 , n9429 , n9430 , n9431 , n9432 , n9433 , n9434 , n9435 , n9436 , n9437 , n9438 , n9439 , n9440 , n9441 , n9442 , n9443 , n9444 , n9445 , n9446 , n9447 , n9448 , n9449 , n9450 , n9451 , n9452 , n9453 , n9454 , n9455 , n9456 , n9457 , n9458 , n9459 , n9460 , n9461 , n9462 , n9463 , n9464 , n9465 , n9466 , n9467 , n9468 , n9469 , n9470 , n9471 , n9472 , n9473 , n9474 , n9475 , n9476 , n9477 , n9478 , n9479 , n9480 , n9481 , n9482 , n9483 , n9484 , n9485 , n9486 , n9487 , n9488 , n9489 , n9490 , n9491 , n9492 , n9493 , n9494 , n9495 , n9496 , n9497 , n9498 , n9499 , n9500 , n9501 , n9502 , n9503 , n9504 , n9505 , n9506 , n9507 , n9508 , n9509 , n9510 , n9511 , n9512 , n9513 , n9514 , n9515 , n9516 , n9517 , n9518 , n9519 , n9520 , n9521 , n9522 , n9523 , n9524 , n9525 , n9526 , n9527 , n9528 , n9529 , n9530 , n9531 , n9532 , n9533 , n9534 , n9535 , n9536 , n9537 , n9538 , n9539 , n9540 , n9541 , n9542 , n9543 , n9544 , n9545 , n9546 , n9547 , n9548 , n9549 , n9550 , n9551 , n9552 , n9553 , n9554 , n9555 , n9556 , n9557 , n9558 , n9559 , n9560 , n9561 , n9562 , n9563 , n9564 , n9565 , n9566 , n9567 , n9568 , n9569 , n9570 , n9571 , n9572 , n9573 , n9574 , n9575 , n9576 , n9577 , n9578 , n9579 , n9580 , n9581 , n9582 , n9583 , n9584 , n9585 , n9586 , n9587 , n9588 , n9589 , n9590 , n9591 , n9592 , n9593 , n9594 , n9595 , n9596 , n9597 , n9598 , n9599 , n9600 , n9601 , n9602 , n9603 , n9604 , n9605 , n9606 , n9607 , n9608 , n9609 , n9610 , n9611 , n9612 , n9613 , n9614 , n9615 , n9616 , n9617 , n9618 , n9619 , n9620 , n9621 , n9622 , n9623 , n9624 , n9625 , n9626 , n9627 , n9628 , n9629 , n9630 , n9631 , n9632 , n9633 , n9634 , n9635 , n9636 , n9637 , n9638 , n9639 , n9640 , n9641 , n9642 , n9643 , n9644 , n9645 , n9646 , n9647 , n9648 , n9649 , n9650 , n9651 , n9652 , n9653 , n9654 , n9655 , n9656 , n9657 , n9658 , n9659 , n9660 , n9661 , n9662 , n9663 , n9664 , n9665 , n9666 , n9667 , n9668 , n9669 , n9670 , n9671 , n9672 , n9673 , n9674 , n9675 , n9676 , n9677 , n9678 , n9679 , n9680 , n9681 , n9682 , n9683 , n9684 , n9685 , n9686 , n9687 , n9688 , n9689 , n9690 , n9691 , n9692 , n9693 , n9694 , n9695 , n9696 , n9697 , n9698 , n9699 , n9700 , n9701 , n9702 , n9703 , n9704 , n9705 , n9706 , n9707 , n9708 , n9709 , n9710 , n9711 , n9712 , n9713 , n9714 , n9715 , n9716 , n9717 , n9718 , n9719 , n9720 , n9721 , n9722 , n9723 , n9724 , n9725 , n9726 , n9727 , n9728 , n9729 , n9730 , n9731 , n9732 , n9733 , n9734 , n9735 , n9736 , n9737 , n9738 , n9739 , n9740 , n9741 , n9742 , n9743 , n9744 , n9745 , n9746 , n9747 , n9748 , n9749 , n9750 , n9751 , n9752 , n9753 , n9754 , n9755 , n9756 , n9757 , n9758 , n9759 , n9760 , n9761 , n9762 , n9763 , n9764 , n9765 , n9766 , n9767 , n9768 , n9769 , n9770 , n9771 , n9772 , n9773 , n9774 , n9775 , n9776 , n9777 , n9778 , n9779 , n9780 , n9781 , n9782 , n9783 , n9784 , n9785 , n9786 , n9787 , n9788 , n9789 , n9790 , n9791 , n9792 , n9793 , n9794 , n9795 , n9796 , n9797 , n9798 , n9799 , n9800 , n9801 , n9802 , n9803 , n9804 , n9805 , n9806 , n9807 , n9808 , n9809 , n9810 , n9811 , n9812 , n9813 , n9814 , n9815 , n9816 , n9817 , n9818 , n9819 , n9820 , n9821 , n9822 , n9823 , n9824 , n9825 , n9826 , n9827 , n9828 , n9829 , n9830 , n9831 , n9832 , n9833 , n9834 , n9835 , n9836 , n9837 , n9838 , n9839 , n9840 , n9841 , n9842 , n9843 , n9844 , n9845 , n9846 , n9847 , n9848 , n9849 , n9850 , n9851 , n9852 , n9853 , n9854 , n9855 , n9856 , n9857 , n9858 , n9859 , n9860 , n9861 , n9862 , n9863 , n9864 , n9865 , n9866 , n9867 , n9868 , n9869 , n9870 , n9871 , n9872 , n9873 , n9874 , n9875 , n9876 , n9877 , n9878 , n9879 , n9880 , n9881 , n9882 , n9883 , n9884 , n9885 , n9886 , n9887 , n9888 , n9889 , n9890 , n9891 , n9892 , n9893 , n9894 , n9895 , n9896 , n9897 , n9898 , n9899 , n9900 , n9901 , n9902 , n9903 , n9904 , n9905 , n9906 , n9907 , n9908 , n9909 , n9910 , n9911 , n9912 , n9913 , n9914 , n9915 , n9916 , n9917 , n9918 , n9919 , n9920 , n9921 , n9922 , n9923 , n9924 , n9925 , n9926 , n9927 , n9928 , n9929 , n9930 , n9931 , n9932 , n9933 , n9934 , n9935 , n9936 , n9937 , n9938 , n9939 , n9940 , n9941 , n9942 , n9943 , n9944 , n9945 , n9946 , n9947 , n9948 , n9949 , n9950 , n9951 , n9952 , n9953 , n9954 , n9955 , n9956 , n9957 , n9958 , n9959 , n9960 , n9961 , n9962 , n9963 , n9964 , n9965 , n9966 , n9967 , n9968 , n9969 , n9970 , n9971 , n9972 , n9973 , n9974 , n9975 , n9976 , n9977 , n9978 , n9979 , n9980 , n9981 , n9982 , n9983 , n9984 , n9985 , n9986 , n9987 , n9988 , n9989 , n9990 , n9991 , n9992 , n9993 , n9994 , n9995 , n9996 , n9997 , n9998 , n9999 , n10000 , n10001 , n10002 , n10003 , n10004 , n10005 , n10006 , n10007 , n10008 , n10009 , n10010 , n10011 , n10012 , n10013 , n10014 , n10015 , n10016 , n10017 , n10018 , n10019 , n10020 , n10021 , n10022 , n10023 , n10024 , n10025 , n10026 , n10027 , n10028 , n10029 , n10030 , n10031 , n10032 , n10033 , n10034 , n10035 , n10036 , n10037 , n10038 , n10039 , n10040 , n10041 , n10042 , n10043 , n10044 , n10045 , n10046 , n10047 , n10048 , n10049 , n10050 , n10051 , n10052 , n10053 , n10054 , n10055 , n10056 , n10057 , n10058 , n10059 , n10060 , n10061 , n10062 , n10063 , n10064 , n10065 , n10066 , n10067 , n10068 , n10069 , n10070 , n10071 , n10072 , n10073 , n10074 , n10075 , n10076 , n10077 , n10078 , n10079 , n10080 , n10081 , n10082 , n10083 , n10084 , n10085 , n10086 , n10087 , n10088 , n10089 , n10090 , n10091 , n10092 , n10093 , n10094 , n10095 , n10096 , n10097 , n10098 , n10099 , n10100 , n10101 , n10102 , n10103 , n10104 , n10105 , n10106 , n10107 , n10108 , n10109 , n10110 , n10111 , n10112 , n10113 , n10114 , n10115 , n10116 , n10117 , n10118 , n10119 , n10120 , n10121 , n10122 , n10123 , n10124 , n10125 , n10126 , n10127 , n10128 , n10129 , n10130 , n10131 , n10132 , n10133 , n10134 , n10135 , n10136 , n10137 , n10138 , n10139 , n10140 , n10141 , n10142 , n10143 , n10144 , n10145 , n10146 , n10147 , n10148 , n10149 , n10150 , n10151 , n10152 , n10153 , n10154 , n10155 , n10156 , n10157 , n10158 , n10159 , n10160 , n10161 , n10162 , n10163 , n10164 , n10165 , n10166 , n10167 , n10168 , n10169 , n10170 , n10171 , n10172 , n10173 , n10174 , n10175 , n10176 , n10177 , n10178 , n10179 , n10180 , n10181 , n10182 , n10183 , n10184 , n10185 , n10186 , n10187 , n10188 , n10189 , n10190 , n10191 , n10192 , n10193 , n10194 , n10195 , n10196 , n10197 , n10198 , n10199 , n10200 , n10201 , n10202 , n10203 , n10204 , n10205 , n10206 , n10207 , n10208 , n10209 , n10210 , n10211 , n10212 , n10213 , n10214 , n10215 , n10216 , n10217 , n10218 , n10219 , n10220 , n10221 , n10222 , n10223 , n10224 , n10225 , n10226 , n10227 , n10228 , n10229 , n10230 , n10231 , n10232 , n10233 , n10234 , n10235 , n10236 , n10237 , n10238 , n10239 , n10240 , n10241 , n10242 , n10243 , n10244 , n10245 , n10246 , n10247 , n10248 , n10249 , n10250 , n10251 , n10252 , n10253 , n10254 , n10255 , n10256 , n10257 , n10258 , n10259 , n10260 , n10261 , n10262 , n10263 , n10264 , n10265 , n10266 , n10267 , n10268 , n10269 , n10270 , n10271 , n10272 , n10273 , n10274 , n10275 , n10276 , n10277 , n10278 , n10279 , n10280 , n10281 , n10282 , n10283 , n10284 , n10285 , n10286 , n10287 , n10288 , n10289 , n10290 , n10291 , n10292 , n10293 , n10294 , n10295 , n10296 , n10297 , n10298 , n10299 , n10300 , n10301 , n10302 , n10303 , n10304 , n10305 , n10306 , n10307 , n10308 , n10309 , n10310 , n10311 , n10312 , n10313 , n10314 , n10315 , n10316 , n10317 , n10318 , n10319 , n10320 , n10321 , n10322 , n10323 , n10324 , n10325 , n10326 , n10327 , n10328 , n10329 , n10330 , n10331 , n10332 , n10333 , n10334 , n10335 , n10336 , n10337 , n10338 , n10339 , n10340 , n10341 , n10342 , n10343 , n10344 , n10345 , n10346 , n10347 , n10348 , n10349 , n10350 , n10351 , n10352 , n10353 , n10354 , n10355 , n10356 , n10357 , n10358 , n10359 , n10360 , n10361 , n10362 , n10363 , n10364 , n10365 , n10366 , n10367 , n10368 , n10369 , n10370 , n10371 , n10372 , n10373 , n10374 , n10375 , n10376 , n10377 , n10378 , n10379 , n10380 , n10381 , n10382 , n10383 , n10384 , n10385 , n10386 , n10387 , n10388 , n10389 , n10390 , n10391 , n10392 , n10393 , n10394 , n10395 , n10396 , n10397 , n10398 , n10399 , n10400 , n10401 , n10402 , n10403 , n10404 , n10405 , n10406 , n10407 , n10408 , n10409 , n10410 , n10411 , n10412 , n10413 , n10414 , n10415 , n10416 , n10417 , n10418 , n10419 , n10420 , n10421 , n10422 , n10423 , n10424 , n10425 , n10426 , n10427 , n10428 , n10429 , n10430 , n10431 , n10432 , n10433 , n10434 , n10435 , n10436 , n10437 , n10438 , n10439 , n10440 , n10441 , n10442 , n10443 , n10444 , n10445 , n10446 , n10447 , n10448 , n10449 , n10450 , n10451 , n10452 , n10453 , n10454 , n10455 , n10456 , n10457 , n10458 , n10459 , n10460 , n10461 , n10462 , n10463 , n10464 , n10465 , n10466 , n10467 , n10468 , n10469 , n10470 , n10471 , n10472 , n10473 , n10474 , n10475 , n10476 , n10477 , n10478 , n10479 , n10480 , n10481 , n10482 , n10483 , n10484 , n10485 , n10486 , n10487 , n10488 , n10489 , n10490 , n10491 , n10492 , n10493 , n10494 , n10495 , n10496 , n10497 , n10498 , n10499 , n10500 , n10501 , n10502 , n10503 , n10504 , n10505 , n10506 , n10507 , n10508 , n10509 , n10510 , n10511 , n10512 , n10513 , n10514 , n10515 , n10516 , n10517 , n10518 , n10519 , n10520 , n10521 , n10522 , n10523 , n10524 , n10525 , n10526 , n10527 , n10528 , n10529 , n10530 , n10531 , n10532 , n10533 , n10534 , n10535 , n10536 , n10537 , n10538 , n10539 , n10540 , n10541 , n10542 , n10543 , n10544 , n10545 , n10546 , n10547 , n10548 , n10549 , n10550 , n10551 , n10552 , n10553 , n10554 , n10555 , n10556 , n10557 , n10558 , n10559 , n10560 , n10561 , n10562 , n10563 , n10564 , n10565 , n10566 , n10567 , n10568 , n10569 , n10570 , n10571 , n10572 , n10573 , n10574 , n10575 , n10576 , n10577 , n10578 , n10579 , n10580 , n10581 , n10582 , n10583 , n10584 , n10585 , n10586 , n10587 , n10588 , n10589 , n10590 , n10591 , n10592 , n10593 , n10594 , n10595 , n10596 , n10597 , n10598 , n10599 , n10600 , n10601 , n10602 , n10603 , n10604 , n10605 , n10606 , n10607 , n10608 , n10609 , n10610 , n10611 , n10612 , n10613 , n10614 , n10615 , n10616 , n10617 , n10618 , n10619 , n10620 , n10621 , n10622 , n10623 , n10624 , n10625 , n10626 , n10627 , n10628 , n10629 , n10630 , n10631 , n10632 , n10633 , n10634 , n10635 , n10636 , n10637 , n10638 , n10639 , n10640 , n10641 , n10642 , n10643 , n10644 , n10645 , n10646 , n10647 , n10648 , n10649 , n10650 , n10651 , n10652 , n10653 , n10654 , n10655 , n10656 , n10657 , n10658 , n10659 , n10660 , n10661 , n10662 , n10663 , n10664 , n10665 , n10666 , n10667 , n10668 , n10669 , n10670 , n10671 , n10672 , n10673 , n10674 , n10675 , n10676 , n10677 , n10678 , n10679 , n10680 , n10681 , n10682 , n10683 , n10684 , n10685 , n10686 , n10687 , n10688 , n10689 , n10690 , n10691 , n10692 , n10693 , n10694 , n10695 , n10696 , n10697 , n10698 , n10699 , n10700 , n10701 , n10702 , n10703 , n10704 , n10705 , n10706 , n10707 , n10708 , n10709 , n10710 , n10711 , n10712 , n10713 , n10714 , n10715 , n10716 , n10717 , n10718 , n10719 , n10720 , n10721 , n10722 , n10723 , n10724 , n10725 , n10726 , n10727 , n10728 , n10729 , n10730 , n10731 , n10732 , n10733 , n10734 , n10735 , n10736 , n10737 , n10738 , n10739 , n10740 , n10741 , n10742 , n10743 , n10744 , n10745 , n10746 , n10747 , n10748 , n10749 , n10750 , n10751 , n10752 , n10753 , n10754 , n10755 , n10756 , n10757 , n10758 , n10759 , n10760 , n10761 , n10762 , n10763 , n10764 , n10765 , n10766 , n10767 , n10768 , n10769 , n10770 , n10771 , n10772 , n10773 , n10774 , n10775 , n10776 , n10777 , n10778 , n10779 , n10780 , n10781 , n10782 , n10783 , n10784 , n10785 , n10786 , n10787 , n10788 , n10789 , n10790 , n10791 , n10792 , n10793 , n10794 , n10795 , n10796 , n10797 , n10798 , n10799 , n10800 , n10801 , n10802 , n10803 , n10804 , n10805 , n10806 , n10807 , n10808 , n10809 , n10810 , n10811 , n10812 , n10813 , n10814 , n10815 , n10816 , n10817 , n10818 , n10819 , n10820 , n10821 , n10822 , n10823 , n10824 , n10825 , n10826 , n10827 , n10828 , n10829 , n10830 , n10831 , n10832 , n10833 , n10834 , n10835 , n10836 , n10837 , n10838 , n10839 , n10840 , n10841 , n10842 , n10843 , n10844 , n10845 , n10846 , n10847 , n10848 , n10849 , n10850 , n10851 , n10852 , n10853 , n10854 , n10855 , n10856 , n10857 , n10858 , n10859 , n10860 , n10861 , n10862 , n10863 , n10864 , n10865 , n10866 , n10867 , n10868 , n10869 , n10870 , n10871 , n10872 , n10873 , n10874 , n10875 , n10876 , n10877 , n10878 , n10879 , n10880 , n10881 , n10882 , n10883 , n10884 , n10885 , n10886 , n10887 , n10888 , n10889 , n10890 , n10891 , n10892 , n10893 , n10894 , n10895 , n10896 , n10897 , n10898 , n10899 , n10900 , n10901 , n10902 , n10903 , n10904 , n10905 , n10906 , n10907 , n10908 , n10909 , n10910 , n10911 , n10912 , n10913 , n10914 , n10915 , n10916 , n10917 , n10918 , n10919 , n10920 , n10921 , n10922 , n10923 , n10924 , n10925 , n10926 , n10927 , n10928 , n10929 , n10930 , n10931 , n10932 , n10933 , n10934 , n10935 , n10936 , n10937 , n10938 , n10939 , n10940 , n10941 , n10942 , n10943 , n10944 , n10945 , n10946 , n10947 , n10948 , n10949 , n10950 , n10951 , n10952 , n10953 , n10954 , n10955 , n10956 , n10957 , n10958 , n10959 , n10960 , n10961 , n10962 , n10963 , n10964 , n10965 , n10966 , n10967 , n10968 , n10969 , n10970 , n10971 , n10972 , n10973 , n10974 , n10975 , n10976 , n10977 , n10978 , n10979 , n10980 , n10981 , n10982 , n10983 , n10984 , n10985 , n10986 , n10987 , n10988 , n10989 , n10990 , n10991 , n10992 , n10993 , n10994 , n10995 , n10996 , n10997 , n10998 , n10999 , n11000 , n11001 , n11002 , n11003 , n11004 , n11005 , n11006 , n11007 , n11008 , n11009 , n11010 , n11011 , n11012 , n11013 , n11014 , n11015 , n11016 , n11017 , n11018 , n11019 , n11020 , n11021 , n11022 , n11023 , n11024 , n11025 , n11026 , n11027 , n11028 , n11029 , n11030 , n11031 , n11032 , n11033 , n11034 , n11035 , n11036 , n11037 , n11038 , n11039 , n11040 , n11041 , n11042 , n11043 , n11044 , n11045 , n11046 , n11047 , n11048 , n11049 , n11050 , n11051 , n11052 , n11053 , n11054 , n11055 , n11056 , n11057 , n11058 , n11059 , n11060 , n11061 , n11062 , n11063 , n11064 , n11065 , n11066 , n11067 , n11068 , n11069 , n11070 , n11071 , n11072 , n11073 , n11074 , n11075 , n11076 , n11077 , n11078 , n11079 , n11080 , n11081 , n11082 , n11083 , n11084 , n11085 , n11086 , n11087 , n11088 , n11089 , n11090 , n11091 , n11092 , n11093 , n11094 , n11095 , n11096 , n11097 , n11098 , n11099 , n11100 , n11101 , n11102 , n11103 , n11104 , n11105 , n11106 , n11107 , n11108 , n11109 , n11110 , n11111 , n11112 , n11113 , n11114 , n11115 , n11116 , n11117 , n11118 , n11119 , n11120 , n11121 , n11122 , n11123 , n11124 , n11125 , n11126 , n11127 , n11128 , n11129 , n11130 , n11131 , n11132 , n11133 , n11134 , n11135 , n11136 , n11137 , n11138 , n11139 , n11140 , n11141 , n11142 , n11143 , n11144 , n11145 , n11146 , n11147 , n11148 , n11149 , n11150 , n11151 , n11152 , n11153 , n11154 , n11155 , n11156 , n11157 , n11158 , n11159 , n11160 , n11161 , n11162 , n11163 , n11164 , n11165 , n11166 , n11167 , n11168 , n11169 , n11170 , n11171 , n11172 , n11173 , n11174 , n11175 , n11176 , n11177 , n11178 , n11179 , n11180 , n11181 , n11182 , n11183 , n11184 , n11185 , n11186 , n11187 , n11188 , n11189 , n11190 , n11191 , n11192 , n11193 , n11194 , n11195 , n11196 , n11197 , n11198 , n11199 , n11200 , n11201 , n11202 , n11203 , n11204 , n11205 , n11206 , n11207 , n11208 , n11209 , n11210 , n11211 , n11212 , n11213 , n11214 , n11215 , n11216 , n11217 , n11218 , n11219 , n11220 , n11221 , n11222 , n11223 , n11224 , n11225 , n11226 , n11227 , n11228 , n11229 , n11230 , n11231 , n11232 , n11233 , n11234 , n11235 , n11236 , n11237 , n11238 , n11239 , n11240 , n11241 , n11242 , n11243 , n11244 , n11245 , n11246 , n11247 , n11248 , n11249 , n11250 , n11251 , n11252 , n11253 , n11254 , n11255 , n11256 , n11257 , n11258 , n11259 , n11260 , n11261 , n11262 , n11263 , n11264 , n11265 , n11266 , n11267 , n11268 , n11269 , n11270 , n11271 , n11272 , n11273 , n11274 , n11275 , n11276 , n11277 , n11278 , n11279 , n11280 , n11281 , n11282 , n11283 , n11284 , n11285 , n11286 , n11287 , n11288 , n11289 , n11290 , n11291 , n11292 , n11293 , n11294 , n11295 , n11296 , n11297 , n11298 , n11299 , n11300 , n11301 , n11302 , n11303 , n11304 , n11305 , n11306 , n11307 , n11308 , n11309 , n11310 , n11311 , n11312 , n11313 , n11314 , n11315 , n11316 , n11317 , n11318 , n11319 , n11320 , n11321 , n11322 , n11323 , n11324 , n11325 , n11326 , n11327 , n11328 , n11329 , n11330 , n11331 , n11332 , n11333 , n11334 , n11335 , n11336 , n11337 , n11338 , n11339 , n11340 , n11341 , n11342 , n11343 , n11344 , n11345 , n11346 , n11347 , n11348 , n11349 , n11350 , n11351 , n11352 , n11353 , n11354 , n11355 , n11356 , n11357 , n11358 , n11359 , n11360 , n11361 , n11362 , n11363 , n11364 , n11365 , n11366 , n11367 , n11368 , n11369 , n11370 , n11371 , n11372 , n11373 , n11374 , n11375 , n11376 , n11377 , n11378 , n11379 , n11380 , n11381 , n11382 , n11383 , n11384 , n11385 , n11386 , n11387 , n11388 , n11389 , n11390 , n11391 , n11392 , n11393 , n11394 , n11395 , n11396 , n11397 , n11398 , n11399 , n11400 , n11401 , n11402 , n11403 , n11404 , n11405 , n11406 , n11407 , n11408 , n11409 , n11410 , n11411 , n11412 , n11413 , n11414 , n11415 , n11416 , n11417 , n11418 , n11419 , n11420 , n11421 , n11422 , n11423 , n11424 , n11425 , n11426 , n11427 , n11428 , n11429 , n11430 , n11431 , n11432 , n11433 , n11434 , n11435 , n11436 , n11437 , n11438 , n11439 , n11440 , n11441 , n11442 , n11443 , n11444 , n11445 , n11446 , n11447 , n11448 , n11449 , n11450 , n11451 , n11452 , n11453 , n11454 , n11455 , n11456 , n11457 , n11458 , n11459 , n11460 , n11461 , n11462 , n11463 , n11464 , n11465 , n11466 , n11467 , n11468 , n11469 , n11470 , n11471 , n11472 , n11473 , n11474 , n11475 , n11476 , n11477 , n11478 , n11479 , n11480 , n11481 , n11482 , n11483 , n11484 , n11485 , n11486 , n11487 , n11488 , n11489 , n11490 , n11491 , n11492 , n11493 , n11494 , n11495 , n11496 , n11497 , n11498 , n11499 , n11500 , n11501 , n11502 , n11503 , n11504 , n11505 , n11506 , n11507 , n11508 , n11509 , n11510 , n11511 , n11512 , n11513 , n11514 , n11515 , n11516 , n11517 , n11518 , n11519 , n11520 , n11521 , n11522 , n11523 , n11524 , n11525 , n11526 , n11527 , n11528 , n11529 , n11530 , n11531 , n11532 , n11533 , n11534 , n11535 , n11536 , n11537 , n11538 , n11539 , n11540 , n11541 , n11542 , n11543 , n11544 , n11545 , n11546 , n11547 , n11548 , n11549 , n11550 , n11551 , n11552 , n11553 , n11554 , n11555 , n11556 , n11557 , n11558 , n11559 , n11560 , n11561 , n11562 , n11563 , n11564 , n11565 , n11566 , n11567 , n11568 , n11569 , n11570 , n11571 , n11572 , n11573 , n11574 , n11575 , n11576 , n11577 , n11578 , n11579 , n11580 , n11581 , n11582 , n11583 , n11584 , n11585 , n11586 , n11587 , n11588 , n11589 , n11590 , n11591 , n11592 , n11593 , n11594 , n11595 , n11596 , n11597 , n11598 , n11599 , n11600 , n11601 , n11602 , n11603 , n11604 , n11605 , n11606 , n11607 , n11608 , n11609 , n11610 , n11611 , n11612 , n11613 , n11614 , n11615 , n11616 , n11617 , n11618 , n11619 , n11620 , n11621 , n11622 , n11623 , n11624 , n11625 , n11626 , n11627 , n11628 , n11629 , n11630 , n11631 , n11632 , n11633 , n11634 , n11635 , n11636 , n11637 , n11638 , n11639 , n11640 , n11641 , n11642 , n11643 , n11644 , n11645 , n11646 , n11647 , n11648 , n11649 , n11650 , n11651 , n11652 , n11653 , n11654 , n11655 , n11656 , n11657 , n11658 , n11659 , n11660 , n11661 , n11662 , n11663 , n11664 , n11665 , n11666 , n11667 , n11668 , n11669 , n11670 , n11671 , n11672 , n11673 , n11674 , n11675 , n11676 , n11677 , n11678 , n11679 , n11680 , n11681 , n11682 , n11683 , n11684 , n11685 , n11686 , n11687 , n11688 , n11689 , n11690 , n11691 , n11692 , n11693 , n11694 , n11695 , n11696 , n11697 , n11698 , n11699 , n11700 , n11701 , n11702 , n11703 , n11704 , n11705 , n11706 , n11707 , n11708 , n11709 , n11710 , n11711 , n11712 , n11713 , n11714 , n11715 , n11716 , n11717 , n11718 , n11719 , n11720 , n11721 , n11722 , n11723 , n11724 , n11725 , n11726 , n11727 , n11728 , n11729 , n11730 , n11731 , n11732 , n11733 , n11734 , n11735 , n11736 , n11737 , n11738 , n11739 , n11740 , n11741 , n11742 , n11743 , n11744 , n11745 , n11746 , n11747 , n11748 , n11749 , n11750 , n11751 , n11752 , n11753 , n11754 , n11755 , n11756 , n11757 , n11758 , n11759 , n11760 , n11761 , n11762 , n11763 , n11764 , n11765 , n11766 , n11767 , n11768 , n11769 , n11770 , n11771 , n11772 , n11773 , n11774 , n11775 , n11776 , n11777 , n11778 , n11779 , n11780 , n11781 , n11782 , n11783 , n11784 , n11785 , n11786 , n11787 , n11788 , n11789 , n11790 , n11791 , n11792 , n11793 , n11794 , n11795 , n11796 , n11797 , n11798 , n11799 , n11800 , n11801 , n11802 , n11803 , n11804 , n11805 , n11806 , n11807 , n11808 , n11809 , n11810 , n11811 , n11812 , n11813 , n11814 , n11815 , n11816 , n11817 , n11818 , n11819 , n11820 , n11821 , n11822 , n11823 , n11824 , n11825 , n11826 , n11827 , n11828 , n11829 , n11830 , n11831 , n11832 , n11833 , n11834 , n11835 , n11836 , n11837 , n11838 , n11839 , n11840 , n11841 , n11842 , n11843 , n11844 , n11845 , n11846 , n11847 , n11848 , n11849 , n11850 , n11851 , n11852 , n11853 , n11854 , n11855 , n11856 , n11857 , n11858 , n11859 , n11860 , n11861 , n11862 , n11863 , n11864 , n11865 , n11866 , n11867 , n11868 , n11869 , n11870 , n11871 , n11872 , n11873 , n11874 , n11875 , n11876 , n11877 , n11878 , n11879 , n11880 , n11881 , n11882 , n11883 , n11884 , n11885 , n11886 , n11887 , n11888 , n11889 , n11890 , n11891 , n11892 , n11893 , n11894 , n11895 , n11896 , n11897 , n11898 , n11899 , n11900 , n11901 , n11902 , n11903 , n11904 , n11905 , n11906 , n11907 , n11908 , n11909 , n11910 , n11911 , n11912 , n11913 , n11914 , n11915 , n11916 , n11917 , n11918 , n11919 , n11920 , n11921 , n11922 , n11923 , n11924 , n11925 , n11926 , n11927 , n11928 , n11929 , n11930 , n11931 , n11932 , n11933 , n11934 , n11935 , n11936 , n11937 , n11938 , n11939 , n11940 , n11941 , n11942 , n11943 , n11944 , n11945 , n11946 , n11947 , n11948 , n11949 , n11950 , n11951 , n11952 , n11953 , n11954 , n11955 , n11956 , n11957 , n11958 , n11959 , n11960 , n11961 , n11962 , n11963 , n11964 , n11965 , n11966 , n11967 , n11968 , n11969 , n11970 , n11971 , n11972 , n11973 , n11974 , n11975 , n11976 , n11977 , n11978 , n11979 , n11980 , n11981 , n11982 , n11983 , n11984 , n11985 , n11986 , n11987 , n11988 , n11989 , n11990 , n11991 , n11992 , n11993 , n11994 , n11995 , n11996 , n11997 , n11998 , n11999 , n12000 , n12001 , n12002 , n12003 , n12004 , n12005 , n12006 , n12007 , n12008 , n12009 , n12010 , n12011 , n12012 , n12013 , n12014 , n12015 , n12016 , n12017 , n12018 , n12019 , n12020 , n12021 , n12022 , n12023 , n12024 , n12025 , n12026 , n12027 , n12028 , n12029 , n12030 , n12031 , n12032 , n12033 , n12034 , n12035 , n12036 , n12037 , n12038 , n12039 , n12040 , n12041 , n12042 , n12043 , n12044 , n12045 , n12046 , n12047 , n12048 , n12049 , n12050 , n12051 , n12052 , n12053 , n12054 , n12055 , n12056 , n12057 , n12058 , n12059 , n12060 , n12061 , n12062 , n12063 , n12064 , n12065 , n12066 , n12067 , n12068 , n12069 , n12070 , n12071 , n12072 , n12073 , n12074 , n12075 , n12076 , n12077 , n12078 , n12079 , n12080 , n12081 , n12082 , n12083 , n12084 , n12085 , n12086 , n12087 , n12088 , n12089 , n12090 , n12091 , n12092 , n12093 , n12094 , n12095 , n12096 , n12097 , n12098 , n12099 , n12100 , n12101 , n12102 , n12103 , n12104 , n12105 , n12106 , n12107 , n12108 , n12109 , n12110 , n12111 , n12112 , n12113 , n12114 , n12115 , n12116 , n12117 , n12118 , n12119 , n12120 , n12121 , n12122 , n12123 , n12124 , n12125 , n12126 , n12127 , n12128 , n12129 , n12130 , n12131 , n12132 , n12133 , n12134 , n12135 , n12136 , n12137 , n12138 , n12139 , n12140 , n12141 , n12142 , n12143 , n12144 , n12145 , n12146 , n12147 , n12148 , n12149 , n12150 , n12151 , n12152 , n12153 , n12154 , n12155 , n12156 , n12157 , n12158 , n12159 , n12160 , n12161 , n12162 , n12163 , n12164 , n12165 , n12166 , n12167 , n12168 , n12169 , n12170 , n12171 , n12172 , n12173 , n12174 , n12175 , n12176 , n12177 , n12178 , n12179 , n12180 , n12181 , n12182 , n12183 , n12184 , n12185 , n12186 , n12187 , n12188 , n12189 , n12190 , n12191 , n12192 , n12193 , n12194 , n12195 , n12196 , n12197 , n12198 , n12199 , n12200 , n12201 , n12202 , n12203 , n12204 , n12205 , n12206 , n12207 , n12208 , n12209 , n12210 , n12211 , n12212 , n12213 , n12214 , n12215 , n12216 , n12217 , n12218 , n12219 , n12220 , n12221 , n12222 , n12223 , n12224 , n12225 , n12226 , n12227 , n12228 , n12229 , n12230 , n12231 , n12232 , n12233 , n12234 , n12235 , n12236 , n12237 , n12238 , n12239 , n12240 , n12241 , n12242 , n12243 , n12244 , n12245 , n12246 , n12247 , n12248 , n12249 , n12250 , n12251 , n12252 , n12253 , n12254 , n12255 , n12256 , n12257 , n12258 , n12259 , n12260 , n12261 , n12262 , n12263 , n12264 , n12265 , n12266 , n12267 , n12268 , n12269 , n12270 , n12271 , n12272 , n12273 , n12274 , n12275 , n12276 , n12277 , n12278 , n12279 , n12280 , n12281 , n12282 , n12283 , n12284 , n12285 , n12286 , n12287 , n12288 , n12289 , n12290 , n12291 , n12292 , n12293 , n12294 , n12295 , n12296 , n12297 , n12298 , n12299 , n12300 , n12301 , n12302 , n12303 , n12304 , n12305 , n12306 , n12307 , n12308 , n12309 , n12310 , n12311 , n12312 , n12313 , n12314 , n12315 , n12316 , n12317 , n12318 , n12319 , n12320 , n12321 , n12322 , n12323 , n12324 , n12325 , n12326 , n12327 , n12328 , n12329 , n12330 , n12331 , n12332 , n12333 , n12334 , n12335 , n12336 , n12337 , n12338 , n12339 , n12340 , n12341 , n12342 , n12343 , n12344 , n12345 , n12346 , n12347 , n12348 , n12349 , n12350 , n12351 , n12352 , n12353 , n12354 , n12355 , n12356 , n12357 , n12358 , n12359 , n12360 , n12361 , n12362 , n12363 , n12364 , n12365 , n12366 , n12367 , n12368 , n12369 , n12370 , n12371 , n12372 , n12373 , n12374 , n12375 , n12376 , n12377 , n12378 , n12379 , n12380 , n12381 , n12382 , n12383 , n12384 , n12385 , n12386 , n12387 , n12388 , n12389 , n12390 , n12391 , n12392 , n12393 , n12394 , n12395 , n12396 , n12397 , n12398 , n12399 , n12400 , n12401 , n12402 , n12403 , n12404 , n12405 , n12406 , n12407 , n12408 , n12409 , n12410 , n12411 , n12412 , n12413 , n12414 , n12415 , n12416 , n12417 , n12418 , n12419 , n12420 , n12421 , n12422 , n12423 , n12424 , n12425 , n12426 , n12427 , n12428 , n12429 , n12430 , n12431 , n12432 , n12433 , n12434 , n12435 , n12436 , n12437 , n12438 , n12439 , n12440 , n12441 , n12442 , n12443 , n12444 , n12445 , n12446 , n12447 , n12448 , n12449 , n12450 , n12451 , n12452 , n12453 , n12454 , n12455 , n12456 , n12457 , n12458 , n12459 , n12460 , n12461 , n12462 , n12463 , n12464 , n12465 , n12466 , n12467 , n12468 , n12469 , n12470 , n12471 , n12472 , n12473 , n12474 , n12475 , n12476 , n12477 , n12478 , n12479 , n12480 , n12481 , n12482 , n12483 , n12484 , n12485 , n12486 , n12487 , n12488 , n12489 , n12490 , n12491 , n12492 , n12493 , n12494 , n12495 , n12496 , n12497 , n12498 , n12499 , n12500 , n12501 , n12502 , n12503 , n12504 , n12505 , n12506 , n12507 , n12508 , n12509 , n12510 , n12511 , n12512 , n12513 , n12514 , n12515 , n12516 , n12517 , n12518 , n12519 , n12520 , n12521 , n12522 , n12523 , n12524 , n12525 , n12526 , n12527 , n12528 , n12529 , n12530 , n12531 , n12532 , n12533 , n12534 , n12535 , n12536 , n12537 , n12538 , n12539 , n12540 , n12541 , n12542 , n12543 , n12544 , n12545 , n12546 , n12547 , n12548 , n12549 , n12550 , n12551 , n12552 , n12553 , n12554 , n12555 , n12556 , n12557 , n12558 , n12559 , n12560 , n12561 , n12562 , n12563 , n12564 , n12565 , n12566 , n12567 , n12568 , n12569 , n12570 , n12571 , n12572 , n12573 , n12574 , n12575 , n12576 , n12577 , n12578 , n12579 , n12580 , n12581 , n12582 , n12583 , n12584 , n12585 , n12586 , n12587 , n12588 , n12589 , n12590 , n12591 , n12592 , n12593 , n12594 , n12595 , n12596 , n12597 , n12598 , n12599 , n12600 , n12601 , n12602 , n12603 , n12604 , n12605 , n12606 , n12607 , n12608 , n12609 , n12610 , n12611 , n12612 , n12613 , n12614 , n12615 , n12616 , n12617 , n12618 , n12619 , n12620 , n12621 , n12622 , n12623 , n12624 , n12625 , n12626 , n12627 , n12628 , n12629 , n12630 , n12631 , n12632 , n12633 , n12634 , n12635 , n12636 , n12637 , n12638 , n12639 , n12640 , n12641 , n12642 , n12643 , n12644 , n12645 , n12646 , n12647 , n12648 , n12649 , n12650 , n12651 , n12652 , n12653 , n12654 , n12655 , n12656 , n12657 , n12658 , n12659 , n12660 , n12661 , n12662 , n12663 , n12664 , n12665 , n12666 , n12667 , n12668 , n12669 , n12670 , n12671 , n12672 , n12673 , n12674 , n12675 , n12676 , n12677 , n12678 , n12679 , n12680 , n12681 , n12682 , n12683 , n12684 , n12685 , n12686 , n12687 , n12688 , n12689 , n12690 , n12691 , n12692 , n12693 , n12694 , n12695 , n12696 , n12697 , n12698 , n12699 , n12700 , n12701 , n12702 , n12703 , n12704 , n12705 , n12706 , n12707 , n12708 , n12709 , n12710 , n12711 , n12712 , n12713 , n12714 , n12715 , n12716 , n12717 , n12718 , n12719 , n12720 , n12721 , n12722 , n12723 , n12724 , n12725 , n12726 , n12727 , n12728 , n12729 , n12730 , n12731 , n12732 , n12733 , n12734 , n12735 , n12736 , n12737 , n12738 , n12739 , n12740 , n12741 , n12742 , n12743 , n12744 , n12745 , n12746 , n12747 , n12748 , n12749 , n12750 , n12751 , n12752 , n12753 , n12754 , n12755 , n12756 , n12757 , n12758 , n12759 , n12760 , n12761 , n12762 , n12763 , n12764 , n12765 , n12766 , n12767 , n12768 , n12769 , n12770 , n12771 , n12772 , n12773 , n12774 , n12775 , n12776 , n12777 , n12778 , n12779 , n12780 , n12781 , n12782 , n12783 , n12784 , n12785 , n12786 , n12787 , n12788 , n12789 , n12790 , n12791 , n12792 , n12793 , n12794 , n12795 , n12796 , n12797 , n12798 , n12799 , n12800 , n12801 , n12802 , n12803 , n12804 , n12805 , n12806 , n12807 , n12808 , n12809 , n12810 , n12811 , n12812 , n12813 , n12814 , n12815 , n12816 , n12817 , n12818 , n12819 , n12820 , n12821 , n12822 , n12823 , n12824 , n12825 , n12826 , n12827 , n12828 , n12829 , n12830 , n12831 , n12832 , n12833 , n12834 , n12835 , n12836 , n12837 , n12838 , n12839 , n12840 , n12841 , n12842 , n12843 , n12844 , n12845 , n12846 , n12847 , n12848 , n12849 , n12850 , n12851 , n12852 , n12853 , n12854 , n12855 , n12856 , n12857 , n12858 , n12859 , n12860 , n12861 , n12862 , n12863 , n12864 , n12865 , n12866 , n12867 , n12868 , n12869 , n12870 , n12871 , n12872 , n12873 , n12874 , n12875 , n12876 , n12877 , n12878 , n12879 , n12880 , n12881 , n12882 , n12883 , n12884 , n12885 , n12886 , n12887 , n12888 , n12889 , n12890 , n12891 , n12892 , n12893 , n12894 , n12895 , n12896 , n12897 , n12898 , n12899 , n12900 , n12901 , n12902 , n12903 , n12904 , n12905 , n12906 , n12907 , n12908 , n12909 , n12910 , n12911 , n12912 , n12913 , n12914 , n12915 , n12916 , n12917 , n12918 , n12919 , n12920 , n12921 , n12922 , n12923 , n12924 , n12925 , n12926 , n12927 , n12928 , n12929 , n12930 , n12931 , n12932 , n12933 , n12934 , n12935 , n12936 , n12937 , n12938 , n12939 , n12940 , n12941 , n12942 , n12943 , n12944 , n12945 , n12946 , n12947 , n12948 , n12949 , n12950 , n12951 , n12952 , n12953 , n12954 , n12955 , n12956 , n12957 , n12958 , n12959 , n12960 , n12961 , n12962 , n12963 , n12964 , n12965 , n12966 , n12967 , n12968 , n12969 , n12970 , n12971 , n12972 , n12973 , n12974 , n12975 , n12976 , n12977 , n12978 , n12979 , n12980 , n12981 , n12982 , n12983 , n12984 , n12985 , n12986 , n12987 , n12988 , n12989 , n12990 , n12991 , n12992 , n12993 , n12994 , n12995 , n12996 , n12997 , n12998 , n12999 , n13000 , n13001 , n13002 , n13003 , n13004 , n13005 , n13006 , n13007 , n13008 , n13009 , n13010 , n13011 , n13012 , n13013 , n13014 , n13015 , n13016 , n13017 , n13018 , n13019 , n13020 , n13021 , n13022 , n13023 , n13024 , n13025 , n13026 , n13027 , n13028 , n13029 , n13030 , n13031 , n13032 , n13033 , n13034 , n13035 , n13036 , n13037 , n13038 , n13039 , n13040 , n13041 , n13042 , n13043 , n13044 , n13045 , n13046 , n13047 , n13048 , n13049 , n13050 , n13051 , n13052 , n13053 , n13054 , n13055 , n13056 , n13057 , n13058 , n13059 , n13060 , n13061 , n13062 , n13063 , n13064 , n13065 , n13066 , n13067 , n13068 , n13069 , n13070 , n13071 , n13072 , n13073 , n13074 , n13075 , n13076 , n13077 , n13078 , n13079 , n13080 , n13081 , n13082 , n13083 , n13084 , n13085 , n13086 , n13087 , n13088 , n13089 , n13090 , n13091 , n13092 , n13093 , n13094 , n13095 , n13096 , n13097 , n13098 , n13099 , n13100 , n13101 , n13102 , n13103 , n13104 , n13105 , n13106 , n13107 , n13108 , n13109 , n13110 , n13111 , n13112 , n13113 , n13114 , n13115 , n13116 , n13117 , n13118 , n13119 , n13120 , n13121 , n13122 , n13123 , n13124 , n13125 , n13126 , n13127 , n13128 , n13129 , n13130 , n13131 , n13132 , n13133 , n13134 , n13135 , n13136 , n13137 , n13138 , n13139 , n13140 , n13141 , n13142 , n13143 , n13144 , n13145 , n13146 , n13147 , n13148 , n13149 , n13150 , n13151 , n13152 , n13153 , n13154 , n13155 , n13156 , n13157 , n13158 , n13159 , n13160 , n13161 , n13162 , n13163 , n13164 , n13165 , n13166 , n13167 , n13168 , n13169 , n13170 , n13171 , n13172 , n13173 , n13174 , n13175 , n13176 , n13177 , n13178 , n13179 , n13180 , n13181 , n13182 , n13183 , n13184 , n13185 , n13186 , n13187 , n13188 , n13189 , n13190 , n13191 , n13192 , n13193 , n13194 , n13195 , n13196 , n13197 , n13198 , n13199 , n13200 , n13201 , n13202 , n13203 , n13204 , n13205 , n13206 , n13207 , n13208 , n13209 , n13210 , n13211 , n13212 , n13213 , n13214 , n13215 , n13216 , n13217 , n13218 , n13219 , n13220 , n13221 , n13222 , n13223 , n13224 , n13225 , n13226 , n13227 , n13228 , n13229 , n13230 , n13231 , n13232 , n13233 , n13234 , n13235 , n13236 , n13237 , n13238 , n13239 , n13240 , n13241 , n13242 , n13243 , n13244 , n13245 , n13246 , n13247 , n13248 , n13249 , n13250 , n13251 , n13252 , n13253 , n13254 , n13255 , n13256 , n13257 , n13258 , n13259 , n13260 , n13261 , n13262 , n13263 , n13264 , n13265 , n13266 , n13267 , n13268 , n13269 , n13270 , n13271 , n13272 , n13273 , n13274 , n13275 , n13276 , n13277 , n13278 , n13279 , n13280 , n13281 , n13282 , n13283 , n13284 , n13285 , n13286 , n13287 , n13288 , n13289 , n13290 , n13291 , n13292 , n13293 , n13294 , n13295 , n13296 , n13297 , n13298 , n13299 , n13300 , n13301 , n13302 , n13303 , n13304 , n13305 , n13306 , n13307 , n13308 , n13309 , n13310 , n13311 , n13312 , n13313 , n13314 , n13315 , n13316 , n13317 , n13318 , n13319 , n13320 , n13321 , n13322 , n13323 , n13324 , n13325 , n13326 , n13327 , n13328 , n13329 , n13330 , n13331 , n13332 , n13333 , n13334 , n13335 , n13336 , n13337 , n13338 , n13339 , n13340 , n13341 , n13342 , n13343 , n13344 , n13345 , n13346 , n13347 , n13348 , n13349 , n13350 , n13351 , n13352 , n13353 , n13354 , n13355 , n13356 , n13357 , n13358 , n13359 , n13360 , n13361 , n13362 , n13363 , n13364 , n13365 , n13366 , n13367 , n13368 , n13369 , n13370 , n13371 , n13372 , n13373 , n13374 , n13375 , n13376 , n13377 , n13378 , n13379 , n13380 , n13381 , n13382 , n13383 , n13384 , n13385 , n13386 , n13387 , n13388 , n13389 , n13390 , n13391 , n13392 , n13393 , n13394 , n13395 , n13396 , n13397 , n13398 , n13399 , n13400 , n13401 , n13402 , n13403 , n13404 , n13405 , n13406 , n13407 , n13408 , n13409 , n13410 , n13411 , n13412 , n13413 , n13414 , n13415 , n13416 , n13417 , n13418 , n13419 , n13420 , n13421 , n13422 , n13423 , n13424 , n13425 , n13426 , n13427 , n13428 , n13429 , n13430 , n13431 , n13432 , n13433 , n13434 , n13435 , n13436 , n13437 , n13438 , n13439 , n13440 , n13441 , n13442 , n13443 , n13444 , n13445 , n13446 , n13447 , n13448 , n13449 , n13450 , n13451 , n13452 , n13453 , n13454 , n13455 , n13456 , n13457 , n13458 , n13459 , n13460 , n13461 , n13462 , n13463 , n13464 , n13465 , n13466 , n13467 , n13468 , n13469 , n13470 , n13471 , n13472 , n13473 , n13474 , n13475 , n13476 , n13477 , n13478 , n13479 , n13480 , n13481 , n13482 , n13483 , n13484 , n13485 , n13486 , n13487 , n13488 , n13489 , n13490 , n13491 , n13492 , n13493 , n13494 , n13495 , n13496 , n13497 , n13498 , n13499 , n13500 , n13501 , n13502 , n13503 , n13504 , n13505 , n13506 , n13507 , n13508 , n13509 , n13510 , n13511 , n13512 , n13513 , n13514 , n13515 , n13516 , n13517 , n13518 , n13519 , n13520 , n13521 , n13522 , n13523 , n13524 , n13525 , n13526 , n13527 , n13528 , n13529 , n13530 , n13531 , n13532 , n13533 , n13534 , n13535 , n13536 , n13537 , n13538 , n13539 , n13540 , n13541 , n13542 , n13543 , n13544 , n13545 , n13546 , n13547 , n13548 , n13549 , n13550 , n13551 , n13552 , n13553 , n13554 , n13555 , n13556 , n13557 , n13558 , n13559 , n13560 , n13561 , n13562 , n13563 , n13564 , n13565 , n13566 , n13567 , n13568 , n13569 , n13570 , n13571 , n13572 , n13573 , n13574 , n13575 , n13576 , n13577 , n13578 , n13579 , n13580 , n13581 , n13582 , n13583 , n13584 , n13585 , n13586 , n13587 , n13588 , n13589 , n13590 , n13591 , n13592 , n13593 , n13594 , n13595 , n13596 , n13597 , n13598 , n13599 , n13600 , n13601 , n13602 , n13603 , n13604 , n13605 , n13606 , n13607 , n13608 , n13609 , n13610 , n13611 , n13612 , n13613 , n13614 , n13615 , n13616 , n13617 , n13618 , n13619 , n13620 , n13621 , n13622 , n13623 , n13624 , n13625 , n13626 , n13627 , n13628 , n13629 , n13630 , n13631 , n13632 , n13633 , n13634 , n13635 , n13636 , n13637 , n13638 , n13639 , n13640 , n13641 , n13642 , n13643 , n13644 , n13645 , n13646 , n13647 , n13648 , n13649 , n13650 , n13651 , n13652 , n13653 , n13654 , n13655 , n13656 , n13657 , n13658 , n13659 , n13660 , n13661 , n13662 , n13663 , n13664 , n13665 , n13666 , n13667 , n13668 , n13669 , n13670 , n13671 , n13672 , n13673 , n13674 , n13675 , n13676 , n13677 , n13678 , n13679 , n13680 , n13681 , n13682 , n13683 , n13684 , n13685 , n13686 , n13687 , n13688 , n13689 , n13690 , n13691 , n13692 , n13693 , n13694 , n13695 , n13696 , n13697 , n13698 , n13699 , n13700 , n13701 , n13702 , n13703 , n13704 , n13705 , n13706 , n13707 , n13708 , n13709 , n13710 , n13711 , n13712 , n13713 , n13714 , n13715 , n13716 , n13717 , n13718 , n13719 , n13720 , n13721 , n13722 , n13723 , n13724 , n13725 , n13726 , n13727 , n13728 , n13729 , n13730 , n13731 , n13732 , n13733 , n13734 , n13735 , n13736 , n13737 , n13738 , n13739 , n13740 , n13741 , n13742 , n13743 , n13744 , n13745 , n13746 , n13747 , n13748 , n13749 , n13750 , n13751 , n13752 , n13753 , n13754 , n13755 , n13756 , n13757 , n13758 , n13759 , n13760 , n13761 , n13762 , n13763 , n13764 , n13765 , n13766 , n13767 , n13768 , n13769 , n13770 , n13771 , n13772 , n13773 , n13774 , n13775 , n13776 , n13777 , n13778 , n13779 , n13780 , n13781 , n13782 , n13783 , n13784 , n13785 , n13786 , n13787 , n13788 , n13789 , n13790 , n13791 , n13792 , n13793 , n13794 , n13795 , n13796 , n13797 , n13798 , n13799 , n13800 , n13801 , n13802 , n13803 , n13804 , n13805 , n13806 , n13807 , n13808 , n13809 , n13810 , n13811 , n13812 , n13813 , n13814 , n13815 , n13816 , n13817 , n13818 , n13819 , n13820 , n13821 , n13822 , n13823 , n13824 , n13825 , n13826 , n13827 , n13828 , n13829 , n13830 , n13831 , n13832 , n13833 , n13834 , n13835 , n13836 , n13837 , n13838 , n13839 , n13840 , n13841 , n13842 , n13843 , n13844 , n13845 , n13846 , n13847 , n13848 , n13849 , n13850 , n13851 , n13852 , n13853 , n13854 , n13855 , n13856 , n13857 , n13858 , n13859 , n13860 , n13861 , n13862 , n13863 , n13864 , n13865 , n13866 , n13867 , n13868 , n13869 , n13870 , n13871 , n13872 , n13873 , n13874 , n13875 , n13876 , n13877 , n13878 , n13879 , n13880 , n13881 , n13882 , n13883 , n13884 , n13885 , n13886 , n13887 , n13888 , n13889 , n13890 , n13891 , n13892 , n13893 , n13894 , n13895 , n13896 , n13897 , n13898 , n13899 , n13900 , n13901 , n13902 , n13903 , n13904 , n13905 , n13906 , n13907 , n13908 , n13909 , n13910 , n13911 , n13912 , n13913 , n13914 , n13915 , n13916 , n13917 , n13918 , n13919 , n13920 , n13921 , n13922 , n13923 , n13924 , n13925 , n13926 , n13927 , n13928 , n13929 , n13930 , n13931 , n13932 , n13933 , n13934 , n13935 , n13936 , n13937 , n13938 , n13939 , n13940 , n13941 , n13942 , n13943 , n13944 , n13945 , n13946 , n13947 , n13948 , n13949 , n13950 , n13951 , n13952 , n13953 , n13954 , n13955 , n13956 , n13957 , n13958 , n13959 , n13960 , n13961 , n13962 , n13963 , n13964 , n13965 , n13966 , n13967 , n13968 , n13969 , n13970 , n13971 , n13972 , n13973 , n13974 , n13975 , n13976 , n13977 , n13978 , n13979 , n13980 , n13981 , n13982 , n13983 , n13984 , n13985 , n13986 , n13987 , n13988 , n13989 , n13990 , n13991 , n13992 , n13993 , n13994 , n13995 , n13996 , n13997 , n13998 , n13999 , n14000 , n14001 , n14002 , n14003 , n14004 , n14005 , n14006 , n14007 , n14008 , n14009 , n14010 , n14011 , n14012 , n14013 , n14014 , n14015 , n14016 , n14017 , n14018 , n14019 , n14020 , n14021 , n14022 , n14023 , n14024 , n14025 , n14026 , n14027 , n14028 , n14029 , n14030 , n14031 , n14032 , n14033 , n14034 , n14035 , n14036 , n14037 , n14038 , n14039 , n14040 , n14041 , n14042 , n14043 , n14044 , n14045 , n14046 , n14047 , n14048 , n14049 , n14050 , n14051 , n14052 , n14053 , n14054 , n14055 , n14056 , n14057 , n14058 , n14059 , n14060 , n14061 , n14062 , n14063 , n14064 , n14065 , n14066 , n14067 , n14068 , n14069 , n14070 , n14071 , n14072 , n14073 , n14074 , n14075 , n14076 , n14077 , n14078 , n14079 , n14080 , n14081 , n14082 , n14083 , n14084 , n14085 , n14086 , n14087 , n14088 , n14089 , n14090 , n14091 , n14092 , n14093 , n14094 , n14095 , n14096 , n14097 , n14098 , n14099 , n14100 , n14101 , n14102 , n14103 , n14104 , n14105 , n14106 , n14107 , n14108 , n14109 , n14110 , n14111 , n14112 , n14113 , n14114 , n14115 , n14116 , n14117 , n14118 , n14119 , n14120 , n14121 , n14122 , n14123 , n14124 , n14125 , n14126 , n14127 , n14128 , n14129 , n14130 , n14131 , n14132 , n14133 , n14134 , n14135 , n14136 , n14137 , n14138 , n14139 , n14140 , n14141 , n14142 , n14143 , n14144 , n14145 , n14146 , n14147 , n14148 , n14149 , n14150 , n14151 , n14152 , n14153 , n14154 , n14155 , n14156 , n14157 , n14158 , n14159 , n14160 , n14161 , n14162 , n14163 , n14164 , n14165 , n14166 , n14167 , n14168 , n14169 , n14170 , n14171 , n14172 , n14173 , n14174 , n14175 , n14176 , n14177 , n14178 , n14179 , n14180 , n14181 , n14182 , n14183 , n14184 , n14185 , n14186 , n14187 , n14188 , n14189 , n14190 , n14191 , n14192 , n14193 , n14194 , n14195 , n14196 , n14197 , n14198 , n14199 , n14200 , n14201 , n14202 , n14203 , n14204 , n14205 , n14206 , n14207 , n14208 , n14209 , n14210 , n14211 , n14212 , n14213 , n14214 , n14215 , n14216 , n14217 , n14218 , n14219 , n14220 , n14221 , n14222 , n14223 , n14224 , n14225 , n14226 , n14227 , n14228 , n14229 , n14230 , n14231 , n14232 , n14233 , n14234 , n14235 , n14236 , n14237 , n14238 , n14239 , n14240 , n14241 , n14242 , n14243 , n14244 , n14245 , n14246 , n14247 , n14248 , n14249 , n14250 , n14251 , n14252 , n14253 , n14254 , n14255 , n14256 , n14257 , n14258 , n14259 , n14260 , n14261 , n14262 , n14263 , n14264 , n14265 , n14266 , n14267 , n14268 , n14269 , n14270 , n14271 , n14272 , n14273 , n14274 , n14275 , n14276 , n14277 , n14278 , n14279 , n14280 , n14281 , n14282 , n14283 , n14284 , n14285 , n14286 , n14287 , n14288 , n14289 , n14290 , n14291 , n14292 , n14293 , n14294 , n14295 , n14296 , n14297 , n14298 , n14299 , n14300 , n14301 , n14302 , n14303 , n14304 , n14305 , n14306 , n14307 , n14308 , n14309 , n14310 , n14311 , n14312 , n14313 , n14314 , n14315 , n14316 , n14317 , n14318 , n14319 , n14320 , n14321 , n14322 , n14323 , n14324 , n14325 , n14326 , n14327 , n14328 , n14329 , n14330 , n14331 , n14332 , n14333 , n14334 , n14335 , n14336 , n14337 , n14338 , n14339 , n14340 , n14341 , n14342 , n14343 , n14344 , n14345 , n14346 , n14347 , n14348 , n14349 , n14350 , n14351 , n14352 , n14353 , n14354 , n14355 , n14356 , n14357 , n14358 , n14359 , n14360 , n14361 , n14362 , n14363 , n14364 , n14365 , n14366 , n14367 , n14368 , n14369 , n14370 , n14371 , n14372 , n14373 , n14374 , n14375 , n14376 , n14377 , n14378 , n14379 , n14380 , n14381 , n14382 , n14383 , n14384 , n14385 , n14386 , n14387 , n14388 , n14389 , n14390 , n14391 , n14392 , n14393 , n14394 , n14395 , n14396 , n14397 , n14398 , n14399 , n14400 , n14401 , n14402 , n14403 , n14404 , n14405 , n14406 , n14407 , n14408 , n14409 , n14410 , n14411 , n14412 , n14413 , n14414 , n14415 , n14416 , n14417 , n14418 , n14419 , n14420 , n14421 , n14422 , n14423 , n14424 , n14425 , n14426 , n14427 , n14428 , n14429 , n14430 , n14431 , n14432 , n14433 , n14434 , n14435 , n14436 , n14437 , n14438 , n14439 , n14440 , n14441 , n14442 , n14443 , n14444 , n14445 , n14446 , n14447 , n14448 , n14449 , n14450 , n14451 , n14452 , n14453 , n14454 , n14455 , n14456 , n14457 , n14458 , n14459 , n14460 , n14461 , n14462 , n14463 , n14464 , n14465 , n14466 , n14467 , n14468 , n14469 , n14470 , n14471 , n14472 , n14473 , n14474 , n14475 , n14476 , n14477 , n14478 , n14479 , n14480 , n14481 , n14482 , n14483 , n14484 , n14485 , n14486 , n14487 , n14488 , n14489 , n14490 , n14491 , n14492 , n14493 , n14494 , n14495 , n14496 , n14497 , n14498 , n14499 , n14500 , n14501 , n14502 , n14503 , n14504 , n14505 , n14506 , n14507 , n14508 , n14509 , n14510 , n14511 , n14512 , n14513 , n14514 , n14515 , n14516 , n14517 , n14518 , n14519 , n14520 , n14521 , n14522 , n14523 , n14524 , n14525 , n14526 , n14527 , n14528 , n14529 , n14530 , n14531 , n14532 , n14533 , n14534 , n14535 , n14536 , n14537 , n14538 , n14539 , n14540 , n14541 , n14542 , n14543 , n14544 , n14545 , n14546 , n14547 , n14548 , n14549 , n14550 , n14551 , n14552 , n14553 , n14554 , n14555 , n14556 , n14557 , n14558 , n14559 , n14560 , n14561 , n14562 , n14563 , n14564 , n14565 , n14566 , n14567 , n14568 , n14569 , n14570 , n14571 , n14572 , n14573 , n14574 , n14575 , n14576 , n14577 , n14578 , n14579 , n14580 , n14581 , n14582 , n14583 , n14584 , n14585 , n14586 , n14587 , n14588 , n14589 , n14590 , n14591 , n14592 , n14593 , n14594 , n14595 , n14596 , n14597 , n14598 , n14599 , n14600 , n14601 , n14602 , n14603 , n14604 , n14605 , n14606 , n14607 , n14608 , n14609 , n14610 , n14611 , n14612 , n14613 , n14614 , n14615 , n14616 , n14617 , n14618 , n14619 , n14620 , n14621 , n14622 , n14623 , n14624 , n14625 , n14626 , n14627 , n14628 , n14629 , n14630 , n14631 , n14632 , n14633 , n14634 , n14635 , n14636 , n14637 , n14638 , n14639 , n14640 , n14641 , n14642 , n14643 , n14644 , n14645 , n14646 , n14647 , n14648 , n14649 , n14650 , n14651 , n14652 , n14653 , n14654 , n14655 , n14656 , n14657 , n14658 , n14659 , n14660 , n14661 , n14662 , n14663 , n14664 , n14665 , n14666 , n14667 , n14668 , n14669 , n14670 , n14671 , n14672 , n14673 , n14674 , n14675 , n14676 , n14677 , n14678 , n14679 , n14680 , n14681 , n14682 , n14683 , n14684 , n14685 , n14686 , n14687 , n14688 , n14689 , n14690 , n14691 , n14692 , n14693 , n14694 , n14695 , n14696 , n14697 , n14698 , n14699 , n14700 , n14701 , n14702 , n14703 , n14704 , n14705 , n14706 , n14707 , n14708 , n14709 , n14710 , n14711 , n14712 , n14713 , n14714 , n14715 , n14716 , n14717 , n14718 , n14719 , n14720 , n14721 , n14722 , n14723 , n14724 , n14725 , n14726 , n14727 , n14728 , n14729 , n14730 , n14731 , n14732 , n14733 , n14734 , n14735 , n14736 , n14737 , n14738 , n14739 , n14740 , n14741 , n14742 , n14743 , n14744 , n14745 , n14746 , n14747 , n14748 , n14749 , n14750 , n14751 , n14752 , n14753 , n14754 , n14755 , n14756 , n14757 , n14758 , n14759 , n14760 , n14761 , n14762 , n14763 , n14764 , n14765 , n14766 , n14767 , n14768 , n14769 , n14770 , n14771 , n14772 , n14773 , n14774 , n14775 , n14776 , n14777 , n14778 , n14779 , n14780 , n14781 , n14782 , n14783 , n14784 , n14785 , n14786 , n14787 , n14788 , n14789 , n14790 , n14791 , n14792 , n14793 , n14794 , n14795 , n14796 , n14797 , n14798 , n14799 , n14800 , n14801 , n14802 , n14803 , n14804 , n14805 , n14806 , n14807 , n14808 , n14809 , n14810 , n14811 , n14812 , n14813 , n14814 , n14815 , n14816 , n14817 , n14818 , n14819 , n14820 , n14821 , n14822 , n14823 , n14824 , n14825 , n14826 , n14827 , n14828 , n14829 , n14830 , n14831 , n14832 , n14833 , n14834 , n14835 , n14836 , n14837 , n14838 , n14839 , n14840 , n14841 , n14842 , n14843 , n14844 , n14845 , n14846 , n14847 , n14848 , n14849 , n14850 , n14851 , n14852 , n14853 , n14854 , n14855 , n14856 , n14857 , n14858 , n14859 , n14860 , n14861 , n14862 , n14863 , n14864 , n14865 , n14866 , n14867 , n14868 , n14869 , n14870 , n14871 , n14872 , n14873 , n14874 , n14875 , n14876 , n14877 , n14878 , n14879 , n14880 , n14881 , n14882 , n14883 , n14884 , n14885 , n14886 , n14887 , n14888 , n14889 , n14890 , n14891 , n14892 , n14893 , n14894 , n14895 , n14896 , n14897 , n14898 , n14899 , n14900 , n14901 , n14902 , n14903 , n14904 , n14905 , n14906 , n14907 , n14908 , n14909 , n14910 , n14911 , n14912 , n14913 , n14914 , n14915 , n14916 , n14917 , n14918 , n14919 , n14920 , n14921 , n14922 , n14923 , n14924 , n14925 , n14926 , n14927 , n14928 , n14929 , n14930 , n14931 , n14932 , n14933 , n14934 , n14935 , n14936 , n14937 , n14938 , n14939 , n14940 , n14941 , n14942 , n14943 , n14944 , n14945 , n14946 , n14947 , n14948 , n14949 , n14950 , n14951 , n14952 , n14953 , n14954 , n14955 , n14956 , n14957 , n14958 , n14959 , n14960 , n14961 , n14962 , n14963 , n14964 , n14965 , n14966 , n14967 , n14968 , n14969 , n14970 , n14971 , n14972 , n14973 , n14974 , n14975 , n14976 , n14977 , n14978 , n14979 , n14980 , n14981 , n14982 , n14983 , n14984 , n14985 , n14986 , n14987 , n14988 , n14989 , n14990 , n14991 , n14992 , n14993 , n14994 , n14995 , n14996 , n14997 , n14998 , n14999 , n15000 , n15001 , n15002 , n15003 , n15004 , n15005 , n15006 , n15007 , n15008 , n15009 , n15010 , n15011 , n15012 , n15013 , n15014 , n15015 , n15016 , n15017 , n15018 , n15019 , n15020 , n15021 , n15022 , n15023 , n15024 , n15025 , n15026 , n15027 , n15028 , n15029 , n15030 , n15031 , n15032 , n15033 , n15034 , n15035 , n15036 , n15037 , n15038 , n15039 , n15040 , n15041 , n15042 , n15043 , n15044 , n15045 , n15046 , n15047 , n15048 , n15049 , n15050 , n15051 , n15052 , n15053 , n15054 , n15055 , n15056 , n15057 , n15058 , n15059 , n15060 , n15061 , n15062 , n15063 , n15064 , n15065 , n15066 , n15067 , n15068 , n15069 , n15070 , n15071 , n15072 , n15073 , n15074 , n15075 , n15076 , n15077 , n15078 , n15079 , n15080 , n15081 , n15082 , n15083 , n15084 , n15085 , n15086 , n15087 , n15088 , n15089 , n15090 , n15091 , n15092 , n15093 , n15094 , n15095 , n15096 , n15097 , n15098 , n15099 , n15100 , n15101 , n15102 , n15103 , n15104 , n15105 , n15106 , n15107 , n15108 , n15109 , n15110 , n15111 , n15112 , n15113 , n15114 , n15115 , n15116 , n15117 , n15118 , n15119 , n15120 , n15121 , n15122 , n15123 , n15124 , n15125 , n15126 , n15127 , n15128 , n15129 , n15130 , n15131 , n15132 , n15133 , n15134 , n15135 , n15136 , n15137 , n15138 , n15139 , n15140 , n15141 , n15142 , n15143 , n15144 , n15145 , n15146 , n15147 , n15148 , n15149 , n15150 , n15151 , n15152 , n15153 , n15154 , n15155 , n15156 , n15157 , n15158 , n15159 , n15160 , n15161 , n15162 , n15163 , n15164 , n15165 , n15166 , n15167 , n15168 , n15169 , n15170 , n15171 , n15172 , n15173 , n15174 , n15175 , n15176 , n15177 , n15178 , n15179 , n15180 , n15181 , n15182 , n15183 , n15184 , n15185 , n15186 , n15187 , n15188 , n15189 , n15190 , n15191 , n15192 , n15193 , n15194 , n15195 , n15196 , n15197 , n15198 , n15199 , n15200 , n15201 , n15202 , n15203 , n15204 , n15205 , n15206 , n15207 , n15208 , n15209 , n15210 , n15211 , n15212 , n15213 , n15214 , n15215 , n15216 , n15217 , n15218 , n15219 , n15220 , n15221 , n15222 , n15223 , n15224 , n15225 , n15226 , n15227 , n15228 , n15229 , n15230 , n15231 , n15232 , n15233 , n15234 , n15235 , n15236 , n15237 , n15238 , n15239 , n15240 , n15241 , n15242 , n15243 , n15244 , n15245 , n15246 , n15247 , n15248 , n15249 , n15250 , n15251 , n15252 , n15253 , n15254 , n15255 , n15256 , n15257 , n15258 , n15259 , n15260 , n15261 , n15262 , n15263 , n15264 , n15265 , n15266 , n15267 , n15268 , n15269 , n15270 , n15271 , n15272 , n15273 , n15274 , n15275 , n15276 , n15277 , n15278 , n15279 , n15280 , n15281 , n15282 , n15283 , n15284 , n15285 , n15286 , n15287 , n15288 , n15289 , n15290 , n15291 , n15292 , n15293 , n15294 , n15295 , n15296 , n15297 , n15298 , n15299 , n15300 , n15301 , n15302 , n15303 , n15304 , n15305 , n15306 , n15307 , n15308 , n15309 , n15310 , n15311 , n15312 , n15313 , n15314 , n15315 , n15316 , n15317 , n15318 , n15319 , n15320 , n15321 , n15322 , n15323 , n15324 , n15325 , n15326 , n15327 , n15328 , n15329 , n15330 , n15331 , n15332 , n15333 , n15334 , n15335 , n15336 , n15337 , n15338 , n15339 , n15340 , n15341 , n15342 , n15343 , n15344 , n15345 , n15346 , n15347 , n15348 , n15349 , n15350 , n15351 , n15352 , n15353 , n15354 , n15355 , n15356 , n15357 , n15358 , n15359 , n15360 , n15361 , n15362 , n15363 , n15364 , n15365 , n15366 , n15367 , n15368 , n15369 , n15370 , n15371 , n15372 , n15373 , n15374 , n15375 , n15376 , n15377 , n15378 , n15379 , n15380 , n15381 , n15382 , n15383 , n15384 , n15385 , n15386 , n15387 , n15388 , n15389 , n15390 , n15391 , n15392 , n15393 , n15394 , n15395 , n15396 , n15397 , n15398 , n15399 , n15400 , n15401 , n15402 , n15403 , n15404 , n15405 , n15406 , n15407 , n15408 , n15409 , n15410 , n15411 , n15412 , n15413 , n15414 , n15415 , n15416 , n15417 , n15418 , n15419 , n15420 , n15421 , n15422 , n15423 , n15424 , n15425 , n15426 , n15427 , n15428 , n15429 , n15430 , n15431 , n15432 , n15433 , n15434 , n15435 , n15436 , n15437 , n15438 , n15439 , n15440 , n15441 , n15442 , n15443 , n15444 , n15445 , n15446 , n15447 , n15448 , n15449 , n15450 , n15451 , n15452 , n15453 , n15454 , n15455 , n15456 , n15457 , n15458 , n15459 , n15460 , n15461 , n15462 , n15463 , n15464 , n15465 , n15466 , n15467 , n15468 , n15469 , n15470 , n15471 , n15472 , n15473 , n15474 , n15475 , n15476 , n15477 , n15478 , n15479 , n15480 , n15481 , n15482 , n15483 , n15484 , n15485 , n15486 , n15487 , n15488 , n15489 , n15490 , n15491 , n15492 , n15493 , n15494 , n15495 , n15496 , n15497 , n15498 , n15499 , n15500 , n15501 , n15502 , n15503 , n15504 , n15505 , n15506 , n15507 , n15508 , n15509 , n15510 , n15511 , n15512 , n15513 , n15514 , n15515 , n15516 , n15517 , n15518 , n15519 , n15520 , n15521 , n15522 , n15523 , n15524 , n15525 , n15526 , n15527 , n15528 , n15529 , n15530 , n15531 , n15532 , n15533 , n15534 , n15535 , n15536 , n15537 , n15538 , n15539 , n15540 , n15541 , n15542 , n15543 , n15544 , n15545 , n15546 , n15547 , n15548 , n15549 , n15550 , n15551 , n15552 , n15553 , n15554 , n15555 , n15556 , n15557 , n15558 , n15559 , n15560 , n15561 , n15562 , n15563 , n15564 , n15565 , n15566 , n15567 , n15568 , n15569 , n15570 , n15571 , n15572 , n15573 , n15574 , n15575 , n15576 , n15577 , n15578 , n15579 , n15580 , n15581 , n15582 , n15583 , n15584 , n15585 , n15586 , n15587 , n15588 , n15589 , n15590 , n15591 , n15592 , n15593 , n15594 , n15595 , n15596 , n15597 , n15598 , n15599 , n15600 , n15601 , n15602 , n15603 , n15604 , n15605 , n15606 , n15607 , n15608 , n15609 , n15610 , n15611 , n15612 , n15613 , n15614 , n15615 , n15616 , n15617 , n15618 , n15619 , n15620 , n15621 , n15622 , n15623 , n15624 , n15625 , n15626 , n15627 , n15628 , n15629 , n15630 , n15631 , n15632 , n15633 , n15634 , n15635 , n15636 , n15637 , n15638 , n15639 , n15640 , n15641 , n15642 , n15643 , n15644 , n15645 , n15646 , n15647 , n15648 , n15649 , n15650 , n15651 , n15652 , n15653 , n15654 , n15655 , n15656 , n15657 , n15658 , n15659 , n15660 , n15661 , n15662 , n15663 , n15664 , n15665 , n15666 , n15667 , n15668 , n15669 , n15670 , n15671 , n15672 , n15673 , n15674 , n15675 , n15676 , n15677 , n15678 , n15679 , n15680 , n15681 , n15682 , n15683 , n15684 , n15685 , n15686 , n15687 , n15688 , n15689 , n15690 , n15691 , n15692 , n15693 , n15694 , n15695 , n15696 , n15697 , n15698 , n15699 , n15700 , n15701 , n15702 , n15703 , n15704 , n15705 , n15706 , n15707 , n15708 , n15709 , n15710 , n15711 , n15712 , n15713 , n15714 , n15715 , n15716 , n15717 , n15718 , n15719 , n15720 , n15721 , n15722 , n15723 , n15724 , n15725 , n15726 , n15727 , n15728 , n15729 , n15730 , n15731 , n15732 , n15733 , n15734 , n15735 , n15736 , n15737 , n15738 , n15739 , n15740 , n15741 , n15742 , n15743 , n15744 , n15745 , n15746 , n15747 , n15748 , n15749 , n15750 , n15751 , n15752 , n15753 , n15754 , n15755 , n15756 , n15757 , n15758 , n15759 , n15760 , n15761 , n15762 , n15763 , n15764 , n15765 , n15766 , n15767 , n15768 , n15769 , n15770 , n15771 , n15772 , n15773 , n15774 , n15775 , n15776 , n15777 , n15778 , n15779 , n15780 , n15781 , n15782 , n15783 , n15784 , n15785 , n15786 , n15787 , n15788 , n15789 , n15790 , n15791 , n15792 , n15793 , n15794 , n15795 , n15796 , n15797 , n15798 , n15799 , n15800 , n15801 , n15802 , n15803 , n15804 , n15805 , n15806 , n15807 , n15808 , n15809 , n15810 , n15811 , n15812 , n15813 , n15814 , n15815 , n15816 , n15817 , n15818 , n15819 , n15820 , n15821 , n15822 , n15823 , n15824 , n15825 , n15826 , n15827 , n15828 , n15829 , n15830 , n15831 , n15832 , n15833 , n15834 , n15835 , n15836 , n15837 , n15838 , n15839 , n15840 , n15841 , n15842 , n15843 , n15844 , n15845 , n15846 , n15847 , n15848 , n15849 , n15850 , n15851 , n15852 , n15853 , n15854 , n15855 , n15856 , n15857 , n15858 , n15859 , n15860 , n15861 , n15862 , n15863 , n15864 , n15865 , n15866 , n15867 , n15868 , n15869 , n15870 , n15871 , n15872 , n15873 , n15874 , n15875 , n15876 , n15877 , n15878 , n15879 , n15880 , n15881 , n15882 , n15883 , n15884 , n15885 , n15886 , n15887 , n15888 , n15889 , n15890 , n15891 , n15892 , n15893 , n15894 , n15895 , n15896 , n15897 , n15898 , n15899 , n15900 , n15901 , n15902 , n15903 , n15904 , n15905 , n15906 , n15907 , n15908 , n15909 , n15910 , n15911 , n15912 , n15913 , n15914 , n15915 , n15916 , n15917 , n15918 , n15919 , n15920 , n15921 , n15922 , n15923 , n15924 , n15925 , n15926 , n15927 , n15928 , n15929 , n15930 , n15931 , n15932 , n15933 , n15934 , n15935 , n15936 , n15937 , n15938 , n15939 , n15940 , n15941 , n15942 , n15943 , n15944 , n15945 , n15946 , n15947 , n15948 , n15949 , n15950 , n15951 , n15952 , n15953 , n15954 , n15955 , n15956 , n15957 , n15958 , n15959 , n15960 , n15961 , n15962 , n15963 , n15964 , n15965 , n15966 , n15967 , n15968 , n15969 , n15970 , n15971 , n15972 , n15973 , n15974 , n15975 , n15976 , n15977 , n15978 , n15979 , n15980 , n15981 , n15982 , n15983 , n15984 , n15985 , n15986 , n15987 , n15988 , n15989 , n15990 , n15991 , n15992 , n15993 , n15994 , n15995 , n15996 , n15997 , n15998 , n15999 , n16000 , n16001 , n16002 , n16003 , n16004 , n16005 , n16006 , n16007 , n16008 , n16009 , n16010 , n16011 , n16012 , n16013 , n16014 , n16015 , n16016 , n16017 , n16018 , n16019 , n16020 , n16021 , n16022 , n16023 , n16024 , n16025 , n16026 , n16027 , n16028 , n16029 , n16030 , n16031 , n16032 , n16033 , n16034 , n16035 , n16036 , n16037 , n16038 , n16039 , n16040 , n16041 , n16042 , n16043 , n16044 , n16045 , n16046 , n16047 , n16048 , n16049 , n16050 , n16051 , n16052 , n16053 , n16054 , n16055 , n16056 , n16057 , n16058 , n16059 , n16060 , n16061 , n16062 , n16063 , n16064 , n16065 , n16066 , n16067 , n16068 , n16069 , n16070 , n16071 , n16072 , n16073 , n16074 , n16075 , n16076 , n16077 , n16078 , n16079 , n16080 , n16081 , n16082 , n16083 , n16084 , n16085 , n16086 , n16087 , n16088 , n16089 , n16090 , n16091 , n16092 , n16093 , n16094 , n16095 , n16096 , n16097 , n16098 , n16099 , n16100 , n16101 , n16102 , n16103 , n16104 , n16105 , n16106 , n16107 , n16108 , n16109 , n16110 , n16111 , n16112 , n16113 , n16114 , n16115 , n16116 , n16117 , n16118 , n16119 , n16120 , n16121 , n16122 , n16123 , n16124 , n16125 , n16126 , n16127 , n16128 , n16129 , n16130 , n16131 , n16132 , n16133 , n16134 , n16135 , n16136 , n16137 , n16138 , n16139 , n16140 , n16141 , n16142 , n16143 , n16144 , n16145 , n16146 , n16147 , n16148 , n16149 , n16150 , n16151 , n16152 , n16153 , n16154 , n16155 , n16156 , n16157 , n16158 , n16159 , n16160 , n16161 , n16162 , n16163 , n16164 , n16165 , n16166 , n16167 , n16168 , n16169 , n16170 , n16171 , n16172 , n16173 , n16174 , n16175 , n16176 , n16177 , n16178 , n16179 , n16180 , n16181 , n16182 , n16183 , n16184 , n16185 , n16186 , n16187 , n16188 , n16189 , n16190 , n16191 , n16192 , n16193 , n16194 , n16195 , n16196 , n16197 , n16198 , n16199 , n16200 , n16201 , n16202 , n16203 , n16204 , n16205 , n16206 , n16207 , n16208 , n16209 , n16210 , n16211 , n16212 , n16213 , n16214 , n16215 , n16216 , n16217 , n16218 , n16219 , n16220 , n16221 , n16222 , n16223 , n16224 , n16225 , n16226 , n16227 , n16228 , n16229 , n16230 , n16231 , n16232 , n16233 , n16234 , n16235 , n16236 , n16237 , n16238 , n16239 , n16240 , n16241 , n16242 , n16243 , n16244 , n16245 , n16246 , n16247 , n16248 , n16249 , n16250 , n16251 , n16252 , n16253 , n16254 , n16255 , n16256 , n16257 , n16258 , n16259 , n16260 , n16261 , n16262 , n16263 , n16264 , n16265 , n16266 , n16267 , n16268 , n16269 , n16270 , n16271 , n16272 , n16273 , n16274 , n16275 , n16276 , n16277 , n16278 , n16279 , n16280 , n16281 , n16282 , n16283 , n16284 , n16285 , n16286 , n16287 , n16288 , n16289 , n16290 , n16291 , n16292 , n16293 , n16294 , n16295 , n16296 , n16297 , n16298 , n16299 , n16300 , n16301 , n16302 , n16303 , n16304 , n16305 , n16306 , n16307 , n16308 , n16309 , n16310 , n16311 , n16312 , n16313 , n16314 , n16315 , n16316 , n16317 , n16318 , n16319 , n16320 , n16321 , n16322 , n16323 , n16324 , n16325 , n16326 , n16327 , n16328 , n16329 , n16330 , n16331 , n16332 , n16333 , n16334 , n16335 , n16336 , n16337 , n16338 , n16339 , n16340 , n16341 , n16342 , n16343 , n16344 , n16345 , n16346 , n16347 , n16348 , n16349 , n16350 , n16351 , n16352 , n16353 , n16354 , n16355 , n16356 , n16357 , n16358 , n16359 , n16360 , n16361 , n16362 , n16363 , n16364 , n16365 , n16366 , n16367 , n16368 , n16369 , n16370 , n16371 , n16372 , n16373 , n16374 , n16375 , n16376 , n16377 , n16378 , n16379 , n16380 , n16381 , n16382 , n16383 , n16384 , n16385 , n16386 , n16387 , n16388 , n16389 , n16390 , n16391 , n16392 , n16393 , n16394 , n16395 , n16396 , n16397 , n16398 , n16399 , n16400 , n16401 , n16402 , n16403 , n16404 , n16405 , n16406 , n16407 , n16408 , n16409 , n16410 , n16411 , n16412 , n16413 , n16414 , n16415 , n16416 , n16417 , n16418 , n16419 , n16420 , n16421 , n16422 , n16423 , n16424 , n16425 , n16426 , n16427 , n16428 , n16429 , n16430 , n16431 , n16432 , n16433 , n16434 , n16435 , n16436 , n16437 , n16438 , n16439 , n16440 , n16441 , n16442 , n16443 , n16444 , n16445 , n16446 , n16447 , n16448 , n16449 , n16450 , n16451 , n16452 , n16453 , n16454 , n16455 , n16456 , n16457 , n16458 , n16459 , n16460 , n16461 , n16462 , n16463 , n16464 , n16465 , n16466 , n16467 , n16468 , n16469 , n16470 , n16471 , n16472 , n16473 , n16474 , n16475 , n16476 , n16477 , n16478 , n16479 , n16480 , n16481 , n16482 , n16483 , n16484 , n16485 , n16486 , n16487 , n16488 , n16489 , n16490 , n16491 , n16492 , n16493 , n16494 , n16495 , n16496 , n16497 , n16498 , n16499 , n16500 , n16501 , n16502 , n16503 , n16504 , n16505 , n16506 , n16507 , n16508 , n16509 , n16510 , n16511 , n16512 , n16513 , n16514 , n16515 , n16516 , n16517 , n16518 , n16519 , n16520 , n16521 , n16522 , n16523 , n16524 , n16525 , n16526 , n16527 , n16528 , n16529 , n16530 , n16531 , n16532 , n16533 , n16534 , n16535 , n16536 , n16537 , n16538 , n16539 , n16540 , n16541 , n16542 , n16543 , n16544 , n16545 , n16546 , n16547 , n16548 , n16549 , n16550 , n16551 , n16552 , n16553 , n16554 , n16555 , n16556 , n16557 , n16558 , n16559 , n16560 , n16561 , n16562 , n16563 , n16564 , n16565 , n16566 , n16567 , n16568 , n16569 , n16570 , n16571 , n16572 , n16573 , n16574 , n16575 , n16576 , n16577 , n16578 , n16579 , n16580 , n16581 , n16582 , n16583 , n16584 , n16585 , n16586 , n16587 , n16588 , n16589 , n16590 , n16591 , n16592 , n16593 , n16594 , n16595 , n16596 , n16597 , n16598 , n16599 , n16600 , n16601 , n16602 , n16603 , n16604 , n16605 , n16606 , n16607 , n16608 , n16609 , n16610 , n16611 , n16612 , n16613 , n16614 , n16615 , n16616 , n16617 , n16618 , n16619 , n16620 , n16621 , n16622 , n16623 , n16624 , n16625 , n16626 , n16627 , n16628 , n16629 , n16630 , n16631 , n16632 , n16633 , n16634 , n16635 , n16636 , n16637 , n16638 , n16639 , n16640 , n16641 , n16642 , n16643 , n16644 , n16645 , n16646 , n16647 , n16648 , n16649 , n16650 , n16651 , n16652 , n16653 , n16654 , n16655 , n16656 , n16657 , n16658 , n16659 , n16660 , n16661 , n16662 , n16663 , n16664 , n16665 , n16666 , n16667 , n16668 , n16669 , n16670 , n16671 , n16672 , n16673 , n16674 , n16675 , n16676 , n16677 , n16678 , n16679 , n16680 , n16681 , n16682 , n16683 , n16684 , n16685 , n16686 , n16687 , n16688 , n16689 , n16690 , n16691 , n16692 , n16693 , n16694 , n16695 , n16696 , n16697 , n16698 , n16699 , n16700 , n16701 , n16702 , n16703 , n16704 , n16705 , n16706 , n16707 , n16708 , n16709 , n16710 , n16711 , n16712 , n16713 , n16714 , n16715 , n16716 , n16717 , n16718 , n16719 , n16720 , n16721 , n16722 , n16723 , n16724 , n16725 , n16726 , n16727 , n16728 , n16729 , n16730 , n16731 , n16732 , n16733 , n16734 , n16735 , n16736 , n16737 , n16738 , n16739 , n16740 , n16741 , n16742 , n16743 , n16744 , n16745 , n16746 , n16747 , n16748 , n16749 , n16750 , n16751 , n16752 , n16753 , n16754 , n16755 , n16756 , n16757 , n16758 , n16759 , n16760 , n16761 , n16762 , n16763 , n16764 , n16765 , n16766 , n16767 , n16768 , n16769 , n16770 , n16771 , n16772 , n16773 , n16774 , n16775 , n16776 , n16777 , n16778 , n16779 , n16780 , n16781 , n16782 , n16783 , n16784 , n16785 , n16786 , n16787 , n16788 , n16789 , n16790 , n16791 , n16792 , n16793 , n16794 , n16795 , n16796 , n16797 , n16798 , n16799 , n16800 , n16801 , n16802 , n16803 , n16804 , n16805 , n16806 , n16807 , n16808 , n16809 , n16810 , n16811 , n16812 , n16813 , n16814 , n16815 , n16816 , n16817 , n16818 , n16819 , n16820 , n16821 , n16822 , n16823 , n16824 , n16825 , n16826 , n16827 , n16828 , n16829 , n16830 , n16831 , n16832 , n16833 , n16834 , n16835 , n16836 , n16837 , n16838 , n16839 , n16840 , n16841 , n16842 , n16843 , n16844 , n16845 , n16846 , n16847 , n16848 , n16849 , n16850 , n16851 , n16852 , n16853 , n16854 , n16855 , n16856 , n16857 , n16858 , n16859 , n16860 , n16861 , n16862 , n16863 , n16864 , n16865 , n16866 , n16867 , n16868 , n16869 , n16870 , n16871 , n16872 , n16873 , n16874 , n16875 , n16876 , n16877 , n16878 , n16879 , n16880 , n16881 , n16882 , n16883 , n16884 , n16885 , n16886 , n16887 , n16888 , n16889 , n16890 , n16891 , n16892 , n16893 , n16894 , n16895 , n16896 , n16897 , n16898 , n16899 , n16900 , n16901 , n16902 , n16903 , n16904 , n16905 , n16906 , n16907 , n16908 , n16909 , n16910 , n16911 , n16912 , n16913 , n16914 , n16915 , n16916 , n16917 , n16918 , n16919 , n16920 , n16921 , n16922 , n16923 , n16924 , n16925 , n16926 , n16927 , n16928 , n16929 , n16930 , n16931 , n16932 , n16933 , n16934 , n16935 , n16936 , n16937 , n16938 , n16939 , n16940 , n16941 , n16942 , n16943 , n16944 , n16945 , n16946 , n16947 , n16948 , n16949 , n16950 , n16951 , n16952 , n16953 , n16954 , n16955 , n16956 , n16957 , n16958 , n16959 , n16960 , n16961 , n16962 , n16963 , n16964 , n16965 , n16966 , n16967 , n16968 , n16969 , n16970 , n16971 , n16972 , n16973 , n16974 , n16975 , n16976 , n16977 , n16978 , n16979 , n16980 , n16981 , n16982 , n16983 , n16984 , n16985 , n16986 , n16987 , n16988 , n16989 , n16990 , n16991 , n16992 , n16993 , n16994 , n16995 , n16996 , n16997 , n16998 , n16999 , n17000 , n17001 , n17002 , n17003 , n17004 , n17005 , n17006 , n17007 , n17008 , n17009 , n17010 , n17011 , n17012 , n17013 , n17014 , n17015 , n17016 , n17017 , n17018 , n17019 , n17020 , n17021 , n17022 , n17023 , n17024 , n17025 , n17026 , n17027 , n17028 , n17029 , n17030 , n17031 , n17032 , n17033 , n17034 , n17035 , n17036 , n17037 , n17038 , n17039 , n17040 , n17041 , n17042 , n17043 , n17044 , n17045 , n17046 , n17047 , n17048 , n17049 , n17050 , n17051 , n17052 , n17053 , n17054 , n17055 , n17056 , n17057 , n17058 , n17059 , n17060 , n17061 , n17062 , n17063 , n17064 , n17065 , n17066 , n17067 , n17068 , n17069 , n17070 , n17071 , n17072 , n17073 , n17074 , n17075 , n17076 , n17077 , n17078 , n17079 , n17080 , n17081 , n17082 , n17083 , n17084 , n17085 , n17086 , n17087 , n17088 , n17089 , n17090 , n17091 , n17092 , n17093 , n17094 , n17095 , n17096 , n17097 , n17098 , n17099 , n17100 , n17101 , n17102 , n17103 , n17104 , n17105 , n17106 , n17107 , n17108 , n17109 , n17110 , n17111 , n17112 , n17113 , n17114 , n17115 , n17116 , n17117 , n17118 , n17119 , n17120 , n17121 , n17122 , n17123 , n17124 , n17125 , n17126 , n17127 , n17128 , n17129 , n17130 , n17131 , n17132 , n17133 , n17134 , n17135 , n17136 , n17137 , n17138 , n17139 , n17140 , n17141 , n17142 , n17143 , n17144 , n17145 , n17146 , n17147 , n17148 , n17149 , n17150 , n17151 , n17152 , n17153 , n17154 , n17155 , n17156 , n17157 , n17158 , n17159 , n17160 , n17161 , n17162 , n17163 , n17164 , n17165 , n17166 , n17167 , n17168 , n17169 , n17170 , n17171 , n17172 , n17173 , n17174 , n17175 , n17176 , n17177 , n17178 , n17179 , n17180 , n17181 , n17182 , n17183 , n17184 , n17185 , n17186 , n17187 , n17188 , n17189 , n17190 , n17191 , n17192 , n17193 , n17194 , n17195 , n17196 , n17197 , n17198 , n17199 , n17200 , n17201 , n17202 , n17203 , n17204 , n17205 , n17206 , n17207 , n17208 , n17209 , n17210 , n17211 , n17212 , n17213 , n17214 , n17215 , n17216 , n17217 , n17218 , n17219 , n17220 , n17221 , n17222 , n17223 , n17224 , n17225 , n17226 , n17227 , n17228 , n17229 , n17230 , n17231 , n17232 , n17233 , n17234 , n17235 , n17236 , n17237 , n17238 , n17239 , n17240 , n17241 , n17242 , n17243 , n17244 , n17245 , n17246 , n17247 , n17248 , n17249 , n17250 , n17251 , n17252 , n17253 , n17254 , n17255 , n17256 , n17257 , n17258 , n17259 , n17260 , n17261 , n17262 , n17263 , n17264 , n17265 , n17266 , n17267 , n17268 , n17269 , n17270 , n17271 , n17272 , n17273 , n17274 , n17275 , n17276 , n17277 , n17278 , n17279 , n17280 , n17281 , n17282 , n17283 , n17284 , n17285 , n17286 , n17287 , n17288 , n17289 , n17290 , n17291 , n17292 , n17293 , n17294 , n17295 , n17296 , n17297 , n17298 , n17299 , n17300 , n17301 , n17302 , n17303 , n17304 , n17305 , n17306 , n17307 , n17308 , n17309 , n17310 , n17311 , n17312 , n17313 , n17314 , n17315 , n17316 , n17317 , n17318 , n17319 , n17320 , n17321 , n17322 , n17323 , n17324 , n17325 , n17326 , n17327 , n17328 , n17329 , n17330 , n17331 , n17332 , n17333 , n17334 , n17335 , n17336 , n17337 , n17338 , n17339 , n17340 , n17341 , n17342 , n17343 , n17344 , n17345 , n17346 , n17347 , n17348 , n17349 , n17350 , n17351 , n17352 , n17353 , n17354 , n17355 , n17356 , n17357 , n17358 , n17359 , n17360 , n17361 , n17362 , n17363 , n17364 , n17365 , n17366 , n17367 , n17368 , n17369 , n17370 , n17371 , n17372 , n17373 , n17374 , n17375 , n17376 , n17377 , n17378 , n17379 , n17380 , n17381 , n17382 , n17383 , n17384 , n17385 , n17386 , n17387 , n17388 , n17389 , n17390 , n17391 , n17392 , n17393 , n17394 , n17395 , n17396 , n17397 , n17398 , n17399 , n17400 , n17401 , n17402 , n17403 , n17404 , n17405 , n17406 , n17407 , n17408 , n17409 , n17410 , n17411 , n17412 , n17413 , n17414 , n17415 , n17416 , n17417 , n17418 , n17419 , n17420 , n17421 , n17422 , n17423 , n17424 , n17425 , n17426 , n17427 , n17428 , n17429 , n17430 , n17431 , n17432 , n17433 , n17434 , n17435 , n17436 , n17437 , n17438 , n17439 , n17440 , n17441 , n17442 , n17443 , n17444 , n17445 , n17446 , n17447 , n17448 , n17449 , n17450 , n17451 , n17452 , n17453 , n17454 , n17455 , n17456 , n17457 , n17458 , n17459 , n17460 , n17461 , n17462 , n17463 , n17464 , n17465 , n17466 , n17467 , n17468 , n17469 , n17470 , n17471 , n17472 , n17473 , n17474 , n17475 , n17476 , n17477 , n17478 , n17479 , n17480 , n17481 , n17482 , n17483 , n17484 , n17485 , n17486 , n17487 , n17488 , n17489 , n17490 , n17491 , n17492 , n17493 , n17494 , n17495 , n17496 , n17497 , n17498 , n17499 , n17500 , n17501 , n17502 , n17503 , n17504 , n17505 , n17506 , n17507 , n17508 , n17509 , n17510 , n17511 , n17512 , n17513 , n17514 , n17515 , n17516 , n17517 , n17518 , n17519 , n17520 , n17521 , n17522 , n17523 , n17524 , n17525 , n17526 , n17527 , n17528 , n17529 , n17530 , n17531 , n17532 , n17533 , n17534 , n17535 , n17536 , n17537 , n17538 , n17539 , n17540 , n17541 , n17542 , n17543 , n17544 , n17545 , n17546 , n17547 , n17548 , n17549 , n17550 , n17551 , n17552 , n17553 , n17554 , n17555 , n17556 , n17557 , n17558 , n17559 , n17560 , n17561 , n17562 , n17563 , n17564 , n17565 , n17566 , n17567 , n17568 , n17569 , n17570 , n17571 , n17572 , n17573 , n17574 , n17575 , n17576 , n17577 , n17578 , n17579 , n17580 , n17581 , n17582 , n17583 , n17584 , n17585 , n17586 , n17587 , n17588 , n17589 , n17590 , n17591 , n17592 , n17593 , n17594 , n17595 , n17596 , n17597 , n17598 , n17599 , n17600 , n17601 , n17602 , n17603 , n17604 , n17605 , n17606 , n17607 , n17608 , n17609 , n17610 , n17611 , n17612 , n17613 , n17614 , n17615 , n17616 , n17617 , n17618 , n17619 , n17620 , n17621 , n17622 , n17623 , n17624 , n17625 , n17626 , n17627 , n17628 , n17629 , n17630 , n17631 , n17632 , n17633 , n17634 , n17635 , n17636 , n17637 , n17638 , n17639 , n17640 , n17641 , n17642 , n17643 , n17644 , n17645 , n17646 , n17647 , n17648 , n17649 , n17650 , n17651 , n17652 , n17653 , n17654 , n17655 , n17656 , n17657 , n17658 , n17659 , n17660 , n17661 , n17662 , n17663 , n17664 , n17665 , n17666 , n17667 , n17668 , n17669 , n17670 , n17671 , n17672 , n17673 , n17674 , n17675 , n17676 , n17677 , n17678 , n17679 , n17680 , n17681 , n17682 , n17683 , n17684 , n17685 , n17686 , n17687 , n17688 , n17689 , n17690 , n17691 , n17692 , n17693 , n17694 , n17695 , n17696 , n17697 , n17698 , n17699 , n17700 , n17701 , n17702 , n17703 , n17704 , n17705 , n17706 , n17707 , n17708 , n17709 , n17710 , n17711 , n17712 , n17713 , n17714 , n17715 , n17716 , n17717 , n17718 , n17719 , n17720 , n17721 , n17722 , n17723 , n17724 , n17725 , n17726 , n17727 , n17728 , n17729 , n17730 , n17731 , n17732 , n17733 , n17734 , n17735 , n17736 , n17737 , n17738 , n17739 , n17740 , n17741 , n17742 , n17743 , n17744 , n17745 , n17746 , n17747 , n17748 , n17749 , n17750 , n17751 , n17752 , n17753 , n17754 , n17755 , n17756 , n17757 , n17758 , n17759 , n17760 , n17761 , n17762 , n17763 , n17764 , n17765 , n17766 , n17767 , n17768 , n17769 , n17770 , n17771 , n17772 , n17773 , n17774 , n17775 , n17776 , n17777 , n17778 , n17779 , n17780 , n17781 , n17782 , n17783 , n17784 , n17785 , n17786 , n17787 , n17788 , n17789 , n17790 , n17791 , n17792 , n17793 , n17794 , n17795 , n17796 , n17797 , n17798 , n17799 , n17800 , n17801 , n17802 , n17803 , n17804 , n17805 , n17806 , n17807 , n17808 , n17809 , n17810 , n17811 , n17812 , n17813 , n17814 , n17815 , n17816 , n17817 , n17818 , n17819 , n17820 , n17821 , n17822 , n17823 , n17824 , n17825 , n17826 , n17827 , n17828 , n17829 , n17830 , n17831 , n17832 , n17833 , n17834 , n17835 , n17836 , n17837 , n17838 , n17839 , n17840 , n17841 , n17842 , n17843 , n17844 , n17845 , n17846 , n17847 , n17848 , n17849 , n17850 , n17851 , n17852 , n17853 , n17854 , n17855 , n17856 , n17857 , n17858 , n17859 , n17860 , n17861 , n17862 , n17863 , n17864 , n17865 , n17866 , n17867 , n17868 , n17869 , n17870 , n17871 , n17872 , n17873 , n17874 , n17875 , n17876 , n17877 , n17878 , n17879 , n17880 , n17881 , n17882 , n17883 , n17884 , n17885 , n17886 , n17887 , n17888 , n17889 , n17890 , n17891 , n17892 , n17893 , n17894 , n17895 , n17896 , n17897 , n17898 , n17899 , n17900 , n17901 , n17902 , n17903 , n17904 , n17905 , n17906 , n17907 , n17908 , n17909 , n17910 , n17911 , n17912 , n17913 , n17914 , n17915 , n17916 , n17917 , n17918 , n17919 , n17920 , n17921 , n17922 , n17923 , n17924 , n17925 , n17926 , n17927 , n17928 , n17929 , n17930 , n17931 , n17932 , n17933 , n17934 , n17935 , n17936 , n17937 , n17938 , n17939 , n17940 , n17941 , n17942 , n17943 , n17944 , n17945 , n17946 , n17947 , n17948 , n17949 , n17950 , n17951 , n17952 , n17953 , n17954 , n17955 , n17956 , n17957 , n17958 , n17959 , n17960 , n17961 , n17962 , n17963 , n17964 , n17965 , n17966 , n17967 , n17968 , n17969 , n17970 , n17971 , n17972 , n17973 , n17974 , n17975 , n17976 , n17977 , n17978 , n17979 , n17980 , n17981 , n17982 , n17983 , n17984 , n17985 , n17986 , n17987 , n17988 , n17989 , n17990 , n17991 , n17992 , n17993 , n17994 , n17995 , n17996 , n17997 , n17998 , n17999 , n18000 , n18001 , n18002 , n18003 , n18004 , n18005 , n18006 , n18007 , n18008 , n18009 , n18010 , n18011 , n18012 , n18013 , n18014 , n18015 , n18016 , n18017 , n18018 , n18019 , n18020 , n18021 , n18022 , n18023 , n18024 , n18025 , n18026 , n18027 , n18028 , n18029 , n18030 , n18031 , n18032 , n18033 , n18034 , n18035 , n18036 , n18037 , n18038 , n18039 , n18040 , n18041 , n18042 , n18043 , n18044 , n18045 , n18046 , n18047 , n18048 , n18049 , n18050 , n18051 , n18052 , n18053 , n18054 , n18055 , n18056 , n18057 , n18058 , n18059 , n18060 , n18061 , n18062 , n18063 , n18064 , n18065 , n18066 , n18067 , n18068 , n18069 , n18070 , n18071 , n18072 , n18073 , n18074 , n18075 , n18076 , n18077 , n18078 , n18079 , n18080 , n18081 , n18082 , n18083 , n18084 , n18085 , n18086 , n18087 , n18088 , n18089 , n18090 , n18091 , n18092 , n18093 , n18094 , n18095 , n18096 , n18097 , n18098 , n18099 , n18100 , n18101 , n18102 , n18103 , n18104 , n18105 , n18106 , n18107 , n18108 , n18109 , n18110 , n18111 , n18112 , n18113 , n18114 , n18115 , n18116 , n18117 , n18118 , n18119 , n18120 , n18121 , n18122 , n18123 , n18124 , n18125 , n18126 , n18127 , n18128 , n18129 , n18130 , n18131 , n18132 , n18133 , n18134 , n18135 , n18136 , n18137 , n18138 , n18139 , n18140 , n18141 , n18142 , n18143 , n18144 , n18145 , n18146 , n18147 , n18148 , n18149 , n18150 , n18151 , n18152 , n18153 , n18154 , n18155 , n18156 , n18157 , n18158 , n18159 , n18160 , n18161 , n18162 , n18163 , n18164 , n18165 , n18166 , n18167 , n18168 , n18169 , n18170 , n18171 , n18172 , n18173 , n18174 , n18175 , n18176 , n18177 , n18178 , n18179 , n18180 , n18181 , n18182 , n18183 , n18184 , n18185 , n18186 , n18187 , n18188 , n18189 , n18190 , n18191 , n18192 , n18193 , n18194 , n18195 , n18196 , n18197 , n18198 , n18199 , n18200 , n18201 , n18202 , n18203 , n18204 , n18205 , n18206 , n18207 , n18208 , n18209 , n18210 , n18211 , n18212 , n18213 , n18214 , n18215 , n18216 , n18217 , n18218 , n18219 , n18220 , n18221 , n18222 , n18223 , n18224 , n18225 , n18226 , n18227 , n18228 , n18229 , n18230 , n18231 , n18232 , n18233 , n18234 , n18235 , n18236 , n18237 , n18238 , n18239 , n18240 , n18241 , n18242 , n18243 , n18244 , n18245 , n18246 , n18247 , n18248 , n18249 , n18250 , n18251 , n18252 , n18253 , n18254 , n18255 , n18256 , n18257 , n18258 , n18259 , n18260 , n18261 , n18262 , n18263 , n18264 , n18265 , n18266 , n18267 , n18268 , n18269 , n18270 , n18271 , n18272 , n18273 , n18274 , n18275 , n18276 , n18277 , n18278 , n18279 , n18280 , n18281 , n18282 , n18283 , n18284 , n18285 , n18286 , n18287 , n18288 , n18289 , n18290 , n18291 , n18292 , n18293 , n18294 , n18295 , n18296 , n18297 , n18298 , n18299 , n18300 , n18301 , n18302 , n18303 , n18304 , n18305 , n18306 , n18307 , n18308 , n18309 , n18310 , n18311 , n18312 , n18313 , n18314 , n18315 , n18316 , n18317 , n18318 , n18319 , n18320 , n18321 , n18322 , n18323 , n18324 , n18325 , n18326 , n18327 , n18328 , n18329 , n18330 , n18331 , n18332 , n18333 , n18334 , n18335 , n18336 , n18337 , n18338 , n18339 , n18340 , n18341 , n18342 , n18343 , n18344 , n18345 , n18346 , n18347 , n18348 , n18349 , n18350 , n18351 , n18352 , n18353 , n18354 , n18355 , n18356 , n18357 , n18358 , n18359 , n18360 , n18361 , n18362 , n18363 , n18364 , n18365 , n18366 , n18367 , n18368 , n18369 , n18370 , n18371 , n18372 , n18373 , n18374 , n18375 , n18376 , n18377 , n18378 , n18379 , n18380 , n18381 , n18382 , n18383 , n18384 , n18385 , n18386 , n18387 , n18388 , n18389 , n18390 , n18391 , n18392 , n18393 , n18394 , n18395 , n18396 , n18397 , n18398 , n18399 , n18400 , n18401 , n18402 , n18403 , n18404 , n18405 , n18406 , n18407 , n18408 , n18409 , n18410 , n18411 , n18412 , n18413 , n18414 , n18415 , n18416 , n18417 , n18418 , n18419 , n18420 , n18421 , n18422 , n18423 , n18424 , n18425 , n18426 , n18427 , n18428 , n18429 , n18430 , n18431 , n18432 , n18433 , n18434 , n18435 , n18436 , n18437 , n18438 , n18439 , n18440 , n18441 , n18442 , n18443 , n18444 , n18445 , n18446 , n18447 , n18448 , n18449 , n18450 , n18451 , n18452 , n18453 , n18454 , n18455 , n18456 , n18457 , n18458 , n18459 , n18460 , n18461 , n18462 , n18463 , n18464 , n18465 , n18466 , n18467 , n18468 , n18469 , n18470 , n18471 , n18472 , n18473 , n18474 , n18475 , n18476 , n18477 , n18478 , n18479 , n18480 , n18481 , n18482 , n18483 , n18484 , n18485 , n18486 , n18487 , n18488 , n18489 , n18490 , n18491 , n18492 , n18493 , n18494 , n18495 , n18496 , n18497 , n18498 , n18499 , n18500 , n18501 , n18502 , n18503 , n18504 , n18505 , n18506 , n18507 , n18508 , n18509 , n18510 , n18511 , n18512 , n18513 , n18514 , n18515 , n18516 , n18517 , n18518 , n18519 , n18520 , n18521 , n18522 , n18523 , n18524 , n18525 , n18526 , n18527 , n18528 , n18529 , n18530 , n18531 , n18532 , n18533 , n18534 , n18535 , n18536 , n18537 , n18538 , n18539 , n18540 , n18541 , n18542 , n18543 , n18544 , n18545 , n18546 , n18547 , n18548 , n18549 , n18550 , n18551 , n18552 , n18553 , n18554 , n18555 , n18556 , n18557 , n18558 , n18559 , n18560 , n18561 , n18562 , n18563 , n18564 , n18565 , n18566 , n18567 , n18568 , n18569 , n18570 , n18571 , n18572 , n18573 , n18574 , n18575 , n18576 , n18577 , n18578 , n18579 , n18580 , n18581 , n18582 , n18583 , n18584 , n18585 , n18586 , n18587 , n18588 , n18589 , n18590 , n18591 , n18592 , n18593 , n18594 , n18595 , n18596 , n18597 , n18598 , n18599 , n18600 , n18601 , n18602 , n18603 , n18604 , n18605 , n18606 , n18607 , n18608 , n18609 , n18610 , n18611 , n18612 , n18613 , n18614 , n18615 , n18616 , n18617 , n18618 , n18619 , n18620 , n18621 , n18622 , n18623 , n18624 , n18625 , n18626 , n18627 , n18628 , n18629 , n18630 , n18631 , n18632 , n18633 , n18634 , n18635 , n18636 , n18637 , n18638 , n18639 , n18640 , n18641 , n18642 , n18643 , n18644 , n18645 , n18646 , n18647 , n18648 , n18649 , n18650 , n18651 , n18652 , n18653 , n18654 , n18655 , n18656 , n18657 , n18658 , n18659 , n18660 , n18661 , n18662 , n18663 , n18664 , n18665 , n18666 , n18667 , n18668 , n18669 , n18670 , n18671 , n18672 , n18673 , n18674 , n18675 , n18676 , n18677 , n18678 , n18679 , n18680 , n18681 , n18682 , n18683 , n18684 , n18685 , n18686 , n18687 , n18688 , n18689 , n18690 , n18691 , n18692 , n18693 , n18694 , n18695 , n18696 , n18697 , n18698 , n18699 , n18700 , n18701 , n18702 , n18703 , n18704 , n18705 , n18706 , n18707 , n18708 , n18709 , n18710 , n18711 , n18712 , n18713 , n18714 , n18715 , n18716 , n18717 , n18718 , n18719 , n18720 , n18721 , n18722 , n18723 , n18724 , n18725 , n18726 , n18727 , n18728 , n18729 , n18730 , n18731 , n18732 , n18733 , n18734 , n18735 , n18736 , n18737 , n18738 , n18739 , n18740 , n18741 , n18742 , n18743 , n18744 , n18745 , n18746 , n18747 , n18748 , n18749 , n18750 , n18751 , n18752 , n18753 , n18754 , n18755 , n18756 , n18757 , n18758 , n18759 , n18760 , n18761 , n18762 , n18763 , n18764 , n18765 , n18766 , n18767 , n18768 , n18769 , n18770 , n18771 , n18772 , n18773 , n18774 , n18775 , n18776 , n18777 , n18778 , n18779 , n18780 , n18781 , n18782 , n18783 , n18784 , n18785 , n18786 , n18787 , n18788 , n18789 , n18790 , n18791 , n18792 , n18793 , n18794 , n18795 , n18796 , n18797 , n18798 , n18799 , n18800 , n18801 , n18802 , n18803 , n18804 , n18805 , n18806 , n18807 , n18808 , n18809 , n18810 , n18811 , n18812 , n18813 , n18814 , n18815 , n18816 , n18817 , n18818 , n18819 , n18820 , n18821 , n18822 , n18823 , n18824 , n18825 , n18826 , n18827 , n18828 , n18829 , n18830 , n18831 , n18832 , n18833 , n18834 , n18835 , n18836 , n18837 , n18838 , n18839 , n18840 , n18841 , n18842 , n18843 , n18844 , n18845 , n18846 , n18847 , n18848 , n18849 , n18850 , n18851 , n18852 , n18853 , n18854 , n18855 , n18856 , n18857 , n18858 , n18859 , n18860 , n18861 , n18862 , n18863 , n18864 , n18865 , n18866 , n18867 , n18868 , n18869 , n18870 , n18871 , n18872 , n18873 , n18874 , n18875 , n18876 , n18877 , n18878 , n18879 , n18880 , n18881 , n18882 , n18883 , n18884 , n18885 , n18886 , n18887 , n18888 , n18889 , n18890 , n18891 , n18892 , n18893 , n18894 , n18895 , n18896 , n18897 , n18898 , n18899 , n18900 , n18901 , n18902 , n18903 , n18904 , n18905 , n18906 , n18907 , n18908 , n18909 , n18910 , n18911 , n18912 , n18913 , n18914 , n18915 , n18916 , n18917 , n18918 , n18919 , n18920 , n18921 , n18922 , n18923 , n18924 , n18925 , n18926 , n18927 , n18928 , n18929 , n18930 , n18931 , n18932 , n18933 , n18934 , n18935 , n18936 , n18937 , n18938 , n18939 , n18940 , n18941 , n18942 , n18943 , n18944 , n18945 , n18946 , n18947 , n18948 , n18949 , n18950 , n18951 , n18952 , n18953 , n18954 , n18955 , n18956 , n18957 , n18958 , n18959 , n18960 , n18961 , n18962 , n18963 , n18964 , n18965 , n18966 , n18967 , n18968 , n18969 , n18970 , n18971 , n18972 , n18973 , n18974 , n18975 , n18976 , n18977 , n18978 , n18979 , n18980 , n18981 , n18982 , n18983 , n18984 , n18985 , n18986 , n18987 , n18988 , n18989 , n18990 , n18991 , n18992 , n18993 , n18994 , n18995 , n18996 , n18997 , n18998 , n18999 , n19000 , n19001 , n19002 , n19003 , n19004 , n19005 , n19006 , n19007 , n19008 , n19009 , n19010 , n19011 , n19012 , n19013 , n19014 , n19015 , n19016 , n19017 , n19018 , n19019 , n19020 , n19021 , n19022 , n19023 , n19024 , n19025 , n19026 , n19027 , n19028 , n19029 , n19030 , n19031 , n19032 , n19033 , n19034 , n19035 , n19036 , n19037 , n19038 , n19039 , n19040 , n19041 , n19042 , n19043 , n19044 , n19045 , n19046 , n19047 , n19048 , n19049 , n19050 , n19051 , n19052 , n19053 , n19054 , n19055 , n19056 , n19057 , n19058 , n19059 , n19060 , n19061 , n19062 , n19063 , n19064 , n19065 , n19066 , n19067 , n19068 , n19069 , n19070 , n19071 , n19072 , n19073 , n19074 , n19075 , n19076 , n19077 , n19078 , n19079 , n19080 , n19081 , n19082 , n19083 , n19084 , n19085 , n19086 , n19087 , n19088 , n19089 , n19090 , n19091 , n19092 , n19093 , n19094 , n19095 , n19096 , n19097 , n19098 , n19099 , n19100 , n19101 , n19102 , n19103 , n19104 , n19105 , n19106 , n19107 , n19108 , n19109 , n19110 , n19111 , n19112 , n19113 , n19114 , n19115 , n19116 , n19117 , n19118 , n19119 , n19120 , n19121 , n19122 , n19123 , n19124 , n19125 , n19126 , n19127 , n19128 , n19129 , n19130 , n19131 , n19132 , n19133 , n19134 , n19135 , n19136 , n19137 , n19138 , n19139 , n19140 , n19141 , n19142 , n19143 , n19144 , n19145 , n19146 , n19147 , n19148 , n19149 , n19150 , n19151 , n19152 , n19153 , n19154 , n19155 , n19156 , n19157 , n19158 , n19159 , n19160 , n19161 , n19162 , n19163 , n19164 , n19165 , n19166 , n19167 , n19168 , n19169 , n19170 , n19171 , n19172 , n19173 , n19174 , n19175 , n19176 , n19177 , n19178 , n19179 , n19180 , n19181 , n19182 , n19183 , n19184 , n19185 , n19186 , n19187 , n19188 , n19189 , n19190 , n19191 , n19192 , n19193 , n19194 , n19195 , n19196 , n19197 , n19198 , n19199 , n19200 , n19201 , n19202 , n19203 , n19204 , n19205 , n19206 , n19207 , n19208 , n19209 , n19210 , n19211 , n19212 , n19213 , n19214 , n19215 , n19216 , n19217 , n19218 , n19219 , n19220 , n19221 , n19222 , n19223 , n19224 , n19225 , n19226 , n19227 , n19228 , n19229 , n19230 , n19231 , n19232 , n19233 , n19234 , n19235 , n19236 , n19237 , n19238 , n19239 , n19240 , n19241 , n19242 , n19243 , n19244 , n19245 , n19246 , n19247 , n19248 , n19249 , n19250 , n19251 , n19252 , n19253 , n19254 , n19255 , n19256 , n19257 , n19258 , n19259 , n19260 , n19261 , n19262 , n19263 , n19264 , n19265 , n19266 , n19267 , n19268 , n19269 , n19270 , n19271 , n19272 , n19273 , n19274 , n19275 , n19276 , n19277 , n19278 , n19279 , n19280 , n19281 , n19282 , n19283 , n19284 , n19285 , n19286 , n19287 , n19288 , n19289 , n19290 , n19291 , n19292 , n19293 , n19294 , n19295 , n19296 , n19297 , n19298 , n19299 , n19300 , n19301 , n19302 , n19303 , n19304 , n19305 , n19306 , n19307 , n19308 , n19309 , n19310 , n19311 , n19312 , n19313 , n19314 , n19315 , n19316 , n19317 , n19318 , n19319 , n19320 , n19321 , n19322 , n19323 , n19324 , n19325 , n19326 , n19327 , n19328 , n19329 , n19330 , n19331 , n19332 , n19333 , n19334 , n19335 , n19336 , n19337 , n19338 , n19339 , n19340 , n19341 , n19342 , n19343 , n19344 , n19345 , n19346 , n19347 , n19348 , n19349 , n19350 , n19351 , n19352 , n19353 , n19354 , n19355 , n19356 , n19357 , n19358 , n19359 , n19360 , n19361 , n19362 , n19363 , n19364 , n19365 , n19366 , n19367 , n19368 , n19369 , n19370 , n19371 , n19372 , n19373 , n19374 , n19375 , n19376 , n19377 , n19378 , n19379 , n19380 , n19381 , n19382 , n19383 , n19384 , n19385 , n19386 , n19387 , n19388 , n19389 , n19390 , n19391 , n19392 , n19393 , n19394 , n19395 , n19396 , n19397 , n19398 , n19399 , n19400 , n19401 , n19402 , n19403 , n19404 , n19405 , n19406 , n19407 , n19408 , n19409 , n19410 , n19411 , n19412 , n19413 , n19414 , n19415 , n19416 , n19417 , n19418 , n19419 , n19420 , n19421 , n19422 , n19423 , n19424 , n19425 , n19426 , n19427 , n19428 , n19429 , n19430 , n19431 , n19432 , n19433 , n19434 , n19435 , n19436 , n19437 , n19438 , n19439 , n19440 , n19441 , n19442 , n19443 , n19444 , n19445 , n19446 , n19447 , n19448 , n19449 , n19450 , n19451 , n19452 , n19453 , n19454 , n19455 , n19456 , n19457 , n19458 , n19459 , n19460 , n19461 , n19462 , n19463 , n19464 , n19465 , n19466 , n19467 , n19468 , n19469 , n19470 , n19471 , n19472 , n19473 , n19474 , n19475 , n19476 , n19477 , n19478 , n19479 , n19480 , n19481 , n19482 , n19483 , n19484 , n19485 , n19486 , n19487 , n19488 , n19489 , n19490 , n19491 , n19492 , n19493 , n19494 , n19495 , n19496 , n19497 , n19498 , n19499 , n19500 , n19501 , n19502 , n19503 , n19504 , n19505 , n19506 , n19507 , n19508 , n19509 , n19510 , n19511 , n19512 , n19513 , n19514 , n19515 , n19516 , n19517 , n19518 , n19519 , n19520 , n19521 , n19522 , n19523 , n19524 , n19525 , n19526 , n19527 , n19528 , n19529 , n19530 , n19531 , n19532 , n19533 , n19534 , n19535 , n19536 , n19537 , n19538 , n19539 , n19540 , n19541 , n19542 , n19543 , n19544 , n19545 , n19546 , n19547 , n19548 , n19549 , n19550 , n19551 , n19552 , n19553 , n19554 , n19555 , n19556 , n19557 , n19558 , n19559 , n19560 , n19561 , n19562 , n19563 , n19564 , n19565 , n19566 , n19567 , n19568 , n19569 , n19570 , n19571 , n19572 , n19573 , n19574 , n19575 , n19576 , n19577 , n19578 , n19579 , n19580 , n19581 , n19582 , n19583 , n19584 , n19585 , n19586 , n19587 , n19588 , n19589 , n19590 , n19591 , n19592 , n19593 , n19594 , n19595 , n19596 , n19597 , n19598 , n19599 , n19600 , n19601 , n19602 , n19603 , n19604 , n19605 , n19606 , n19607 , n19608 , n19609 , n19610 , n19611 , n19612 , n19613 , n19614 , n19615 , n19616 , n19617 , n19618 , n19619 , n19620 , n19621 , n19622 , n19623 , n19624 , n19625 , n19626 , n19627 , n19628 , n19629 , n19630 , n19631 , n19632 , n19633 , n19634 , n19635 , n19636 , n19637 , n19638 , n19639 , n19640 , n19641 , n19642 , n19643 , n19644 , n19645 , n19646 , n19647 , n19648 , n19649 , n19650 , n19651 , n19652 , n19653 , n19654 , n19655 , n19656 , n19657 , n19658 , n19659 , n19660 , n19661 , n19662 , n19663 , n19664 , n19665 , n19666 , n19667 , n19668 , n19669 , n19670 , n19671 , n19672 , n19673 , n19674 , n19675 , n19676 , n19677 , n19678 , n19679 , n19680 , n19681 , n19682 , n19683 , n19684 , n19685 , n19686 , n19687 , n19688 , n19689 , n19690 , n19691 , n19692 , n19693 , n19694 , n19695 , n19696 , n19697 , n19698 , n19699 , n19700 , n19701 , n19702 , n19703 , n19704 , n19705 , n19706 , n19707 , n19708 , n19709 , n19710 , n19711 , n19712 , n19713 , n19714 , n19715 , n19716 , n19717 , n19718 , n19719 , n19720 , n19721 , n19722 , n19723 , n19724 , n19725 , n19726 , n19727 , n19728 , n19729 , n19730 , n19731 , n19732 , n19733 , n19734 , n19735 , n19736 , n19737 , n19738 , n19739 , n19740 , n19741 , n19742 , n19743 , n19744 , n19745 , n19746 , n19747 , n19748 , n19749 , n19750 , n19751 , n19752 , n19753 , n19754 , n19755 , n19756 , n19757 , n19758 , n19759 , n19760 , n19761 , n19762 , n19763 , n19764 , n19765 , n19766 , n19767 , n19768 , n19769 , n19770 , n19771 , n19772 , n19773 , n19774 , n19775 , n19776 , n19777 , n19778 , n19779 , n19780 , n19781 , n19782 , n19783 , n19784 , n19785 , n19786 , n19787 , n19788 , n19789 , n19790 , n19791 , n19792 , n19793 , n19794 , n19795 , n19796 , n19797 , n19798 , n19799 , n19800 , n19801 , n19802 , n19803 , n19804 , n19805 , n19806 , n19807 , n19808 , n19809 , n19810 , n19811 , n19812 , n19813 , n19814 , n19815 , n19816 , n19817 , n19818 , n19819 , n19820 , n19821 , n19822 , n19823 , n19824 , n19825 , n19826 , n19827 , n19828 , n19829 , n19830 , n19831 , n19832 , n19833 , n19834 , n19835 , n19836 , n19837 , n19838 , n19839 , n19840 , n19841 , n19842 , n19843 , n19844 , n19845 , n19846 , n19847 , n19848 , n19849 , n19850 , n19851 , n19852 , n19853 , n19854 , n19855 , n19856 , n19857 , n19858 , n19859 , n19860 , n19861 , n19862 , n19863 , n19864 , n19865 , n19866 , n19867 , n19868 , n19869 , n19870 , n19871 , n19872 , n19873 , n19874 , n19875 , n19876 , n19877 , n19878 , n19879 , n19880 , n19881 , n19882 , n19883 , n19884 , n19885 , n19886 , n19887 , n19888 , n19889 , n19890 , n19891 , n19892 , n19893 , n19894 , n19895 , n19896 , n19897 , n19898 , n19899 , n19900 , n19901 , n19902 , n19903 , n19904 , n19905 , n19906 , n19907 , n19908 , n19909 , n19910 , n19911 , n19912 , n19913 , n19914 , n19915 , n19916 , n19917 , n19918 , n19919 , n19920 , n19921 , n19922 , n19923 , n19924 , n19925 , n19926 , n19927 , n19928 , n19929 , n19930 , n19931 , n19932 , n19933 , n19934 , n19935 , n19936 , n19937 , n19938 , n19939 , n19940 , n19941 , n19942 , n19943 , n19944 , n19945 , n19946 , n19947 , n19948 , n19949 , n19950 , n19951 , n19952 , n19953 , n19954 , n19955 , n19956 , n19957 , n19958 , n19959 , n19960 , n19961 , n19962 , n19963 , n19964 , n19965 , n19966 , n19967 ;
  assign n563 = ~\sa13_reg[4]/P0001  & \sa13_reg[6]/NET0131  ;
  assign n570 = ~\sa13_reg[5]/P0001  & \sa13_reg[7]/NET0131  ;
  assign n571 = n563 & n570 ;
  assign n572 = ~\sa13_reg[3]/P0001  & n571 ;
  assign n543 = \sa13_reg[6]/NET0131  & ~\sa13_reg[7]/NET0131  ;
  assign n567 = \sa13_reg[4]/P0001  & n543 ;
  assign n549 = ~\sa13_reg[6]/NET0131  & \sa13_reg[7]/NET0131  ;
  assign n568 = \sa13_reg[5]/P0001  & n549 ;
  assign n569 = ~\sa13_reg[4]/P0001  & n568 ;
  assign n573 = ~n567 & ~n569 ;
  assign n574 = ~n572 & n573 ;
  assign n575 = \sa13_reg[2]/P0001  & ~n574 ;
  assign n555 = \sa13_reg[3]/P0001  & \sa13_reg[4]/P0001  ;
  assign n556 = ~\sa13_reg[6]/NET0131  & ~\sa13_reg[7]/NET0131  ;
  assign n557 = \sa13_reg[5]/P0001  & n556 ;
  assign n558 = n555 & n557 ;
  assign n559 = \sa13_reg[5]/P0001  & \sa13_reg[7]/NET0131  ;
  assign n560 = \sa13_reg[3]/P0001  & n559 ;
  assign n561 = ~\sa13_reg[4]/P0001  & n560 ;
  assign n562 = ~n558 & ~n561 ;
  assign n564 = ~\sa13_reg[2]/P0001  & ~\sa13_reg[5]/P0001  ;
  assign n565 = ~\sa13_reg[3]/P0001  & n564 ;
  assign n566 = ~n563 & n565 ;
  assign n576 = n562 & ~n566 ;
  assign n577 = ~n575 & n576 ;
  assign n578 = \sa13_reg[1]/P0001  & ~n577 ;
  assign n589 = ~\sa13_reg[3]/P0001  & n557 ;
  assign n590 = ~\sa13_reg[2]/P0001  & ~n589 ;
  assign n592 = \sa13_reg[7]/NET0131  & n555 ;
  assign n591 = ~\sa13_reg[5]/P0001  & n543 ;
  assign n593 = \sa13_reg[2]/P0001  & ~n591 ;
  assign n594 = ~n592 & n593 ;
  assign n595 = ~n590 & ~n594 ;
  assign n579 = ~\sa13_reg[5]/P0001  & ~\sa13_reg[7]/NET0131  ;
  assign n580 = \sa13_reg[4]/P0001  & n579 ;
  assign n581 = ~\sa13_reg[2]/P0001  & \sa13_reg[3]/P0001  ;
  assign n582 = n580 & n581 ;
  assign n583 = \sa13_reg[6]/NET0131  & \sa13_reg[7]/NET0131  ;
  assign n584 = ~\sa13_reg[4]/P0001  & n583 ;
  assign n585 = n564 & n584 ;
  assign n586 = ~n582 & ~n585 ;
  assign n532 = \sa13_reg[5]/P0001  & ~\sa13_reg[6]/NET0131  ;
  assign n587 = \sa13_reg[4]/P0001  & \sa13_reg[7]/NET0131  ;
  assign n588 = n532 & n587 ;
  assign n596 = n586 & ~n588 ;
  assign n597 = ~n595 & n596 ;
  assign n598 = ~\sa13_reg[1]/P0001  & ~n597 ;
  assign n533 = ~\sa13_reg[3]/P0001  & \sa13_reg[4]/P0001  ;
  assign n534 = n532 & n533 ;
  assign n535 = \sa13_reg[5]/P0001  & \sa13_reg[6]/NET0131  ;
  assign n536 = ~\sa13_reg[4]/P0001  & ~\sa13_reg[7]/NET0131  ;
  assign n537 = n535 & n536 ;
  assign n538 = ~n534 & ~n537 ;
  assign n539 = ~\sa13_reg[2]/P0001  & ~n538 ;
  assign n540 = \sa13_reg[7]/NET0131  & n535 ;
  assign n541 = ~\sa13_reg[3]/P0001  & n540 ;
  assign n542 = \sa13_reg[4]/P0001  & n541 ;
  assign n544 = \sa13_reg[3]/P0001  & n543 ;
  assign n545 = \sa13_reg[4]/P0001  & n544 ;
  assign n546 = ~n542 & ~n545 ;
  assign n547 = ~\sa13_reg[5]/P0001  & ~\sa13_reg[6]/NET0131  ;
  assign n548 = n536 & n547 ;
  assign n550 = \sa13_reg[3]/P0001  & ~\sa13_reg[5]/P0001  ;
  assign n551 = n549 & n550 ;
  assign n552 = ~n548 & ~n551 ;
  assign n553 = n546 & n552 ;
  assign n554 = \sa13_reg[2]/P0001  & ~n553 ;
  assign n599 = ~n539 & ~n554 ;
  assign n600 = ~n598 & n599 ;
  assign n601 = ~n578 & n600 ;
  assign n602 = \sa13_reg[0]/P0001  & ~n601 ;
  assign n603 = \sa13_reg[2]/P0001  & ~\sa13_reg[3]/P0001  ;
  assign n604 = ~\sa13_reg[4]/P0001  & n579 ;
  assign n605 = \sa13_reg[4]/P0001  & n559 ;
  assign n606 = ~n604 & ~n605 ;
  assign n607 = n603 & ~n606 ;
  assign n610 = ~\sa13_reg[4]/P0001  & n547 ;
  assign n611 = ~\sa13_reg[2]/P0001  & ~\sa13_reg[7]/NET0131  ;
  assign n612 = n610 & n611 ;
  assign n608 = \sa13_reg[5]/P0001  & n555 ;
  assign n609 = n543 & n608 ;
  assign n613 = \sa13_reg[1]/P0001  & ~n609 ;
  assign n614 = ~n612 & n613 ;
  assign n615 = ~n607 & n614 ;
  assign n623 = \sa13_reg[2]/P0001  & \sa13_reg[3]/P0001  ;
  assign n624 = n557 & n623 ;
  assign n625 = n581 & n587 ;
  assign n626 = ~\sa13_reg[1]/P0001  & ~n537 ;
  assign n627 = ~n625 & n626 ;
  assign n628 = ~n624 & n627 ;
  assign n616 = \sa13_reg[3]/P0001  & n570 ;
  assign n617 = ~\sa13_reg[3]/P0001  & n549 ;
  assign n618 = ~n616 & ~n617 ;
  assign n619 = ~\sa13_reg[4]/P0001  & ~n618 ;
  assign n620 = \sa13_reg[6]/NET0131  & n533 ;
  assign n621 = ~\sa13_reg[5]/P0001  & n620 ;
  assign n622 = \sa13_reg[7]/NET0131  & n621 ;
  assign n629 = ~n619 & ~n622 ;
  assign n630 = n628 & n629 ;
  assign n631 = ~n615 & ~n630 ;
  assign n632 = \sa13_reg[4]/P0001  & n547 ;
  assign n633 = ~\sa13_reg[3]/P0001  & n632 ;
  assign n639 = ~\sa13_reg[2]/P0001  & ~n633 ;
  assign n634 = n550 & ~n556 ;
  assign n635 = \sa13_reg[4]/P0001  & ~n583 ;
  assign n636 = n634 & ~n635 ;
  assign n637 = ~\sa13_reg[7]/NET0131  & n533 ;
  assign n638 = n535 & n637 ;
  assign n640 = ~n636 & ~n638 ;
  assign n641 = n639 & n640 ;
  assign n642 = ~\sa13_reg[3]/P0001  & n610 ;
  assign n643 = \sa13_reg[2]/P0001  & ~n642 ;
  assign n644 = ~n622 & n643 ;
  assign n645 = ~n641 & ~n644 ;
  assign n646 = ~n631 & ~n645 ;
  assign n647 = ~\sa13_reg[0]/P0001  & ~n646 ;
  assign n655 = \sa13_reg[3]/P0001  & ~\sa13_reg[4]/P0001  ;
  assign n656 = \sa13_reg[5]/P0001  & n655 ;
  assign n657 = n549 & n656 ;
  assign n652 = ~\sa13_reg[6]/NET0131  & n580 ;
  assign n653 = ~\sa13_reg[3]/P0001  & ~\sa13_reg[4]/P0001  ;
  assign n654 = n556 & n653 ;
  assign n658 = ~n652 & ~n654 ;
  assign n659 = ~n657 & n658 ;
  assign n660 = \sa13_reg[1]/P0001  & ~n659 ;
  assign n648 = n543 & n550 ;
  assign n649 = \sa13_reg[4]/P0001  & n648 ;
  assign n650 = ~\sa13_reg[5]/P0001  & n556 ;
  assign n651 = ~\sa13_reg[3]/P0001  & n650 ;
  assign n661 = ~n649 & ~n651 ;
  assign n662 = ~n660 & n661 ;
  assign n663 = \sa13_reg[2]/P0001  & ~n662 ;
  assign n664 = n568 & ~n653 ;
  assign n665 = ~\sa13_reg[5]/P0001  & n567 ;
  assign n666 = ~n664 & ~n665 ;
  assign n667 = ~\sa13_reg[2]/P0001  & ~n666 ;
  assign n668 = n535 & n653 ;
  assign n669 = ~\sa13_reg[6]/NET0131  & n592 ;
  assign n674 = ~n668 & ~n669 ;
  assign n670 = \sa13_reg[2]/P0001  & ~\sa13_reg[4]/P0001  ;
  assign n671 = n540 & n670 ;
  assign n672 = ~\sa13_reg[4]/P0001  & n556 ;
  assign n673 = n623 & n672 ;
  assign n675 = ~n671 & ~n673 ;
  assign n676 = n674 & n675 ;
  assign n677 = ~n667 & n676 ;
  assign n678 = ~\sa13_reg[1]/P0001  & ~n677 ;
  assign n680 = \sa13_reg[1]/P0001  & ~\sa13_reg[2]/P0001  ;
  assign n681 = n557 & n655 ;
  assign n682 = n680 & n681 ;
  assign n679 = n581 & n588 ;
  assign n683 = ~\sa13_reg[5]/P0001  & n654 ;
  assign n684 = ~n679 & ~n683 ;
  assign n685 = ~n682 & n684 ;
  assign n686 = ~n678 & n685 ;
  assign n687 = ~n663 & n686 ;
  assign n688 = ~n647 & n687 ;
  assign n689 = ~n602 & n688 ;
  assign n735 = ~\sa20_reg[5]/P0001  & \sa20_reg[6]/NET0131  ;
  assign n736 = ~\sa20_reg[3]/P0001  & \sa20_reg[7]/NET0131  ;
  assign n737 = n735 & n736 ;
  assign n738 = ~\sa20_reg[4]/P0001  & n737 ;
  assign n693 = \sa20_reg[6]/NET0131  & ~\sa20_reg[7]/NET0131  ;
  assign n739 = \sa20_reg[4]/P0001  & n693 ;
  assign n694 = ~\sa20_reg[4]/P0001  & \sa20_reg[5]/P0001  ;
  assign n705 = ~\sa20_reg[6]/NET0131  & \sa20_reg[7]/NET0131  ;
  assign n740 = n694 & n705 ;
  assign n741 = ~n739 & ~n740 ;
  assign n742 = ~n738 & n741 ;
  assign n743 = \sa20_reg[2]/P0001  & ~n742 ;
  assign n716 = \sa20_reg[3]/P0001  & \sa20_reg[4]/P0001  ;
  assign n750 = ~\sa20_reg[6]/NET0131  & n716 ;
  assign n751 = \sa20_reg[5]/P0001  & n750 ;
  assign n752 = ~\sa20_reg[7]/NET0131  & n751 ;
  assign n744 = \sa20_reg[5]/P0001  & \sa20_reg[7]/NET0131  ;
  assign n745 = \sa20_reg[3]/P0001  & ~\sa20_reg[4]/P0001  ;
  assign n746 = n744 & n745 ;
  assign n747 = ~\sa20_reg[2]/P0001  & ~\sa20_reg[3]/P0001  ;
  assign n719 = ~\sa20_reg[4]/P0001  & \sa20_reg[6]/NET0131  ;
  assign n748 = ~\sa20_reg[5]/P0001  & ~n719 ;
  assign n749 = n747 & n748 ;
  assign n753 = ~n746 & ~n749 ;
  assign n754 = ~n752 & n753 ;
  assign n755 = ~n743 & n754 ;
  assign n756 = \sa20_reg[1]/P0001  & ~n755 ;
  assign n717 = ~\sa20_reg[5]/P0001  & ~\sa20_reg[7]/NET0131  ;
  assign n718 = n716 & n717 ;
  assign n720 = ~\sa20_reg[5]/P0001  & \sa20_reg[7]/NET0131  ;
  assign n721 = n719 & n720 ;
  assign n722 = ~n718 & ~n721 ;
  assign n723 = ~\sa20_reg[6]/NET0131  & ~\sa20_reg[7]/NET0131  ;
  assign n724 = \sa20_reg[5]/P0001  & n723 ;
  assign n725 = ~\sa20_reg[3]/P0001  & n724 ;
  assign n726 = n722 & ~n725 ;
  assign n727 = ~\sa20_reg[2]/P0001  & ~n726 ;
  assign n690 = \sa20_reg[5]/P0001  & ~\sa20_reg[6]/NET0131  ;
  assign n714 = \sa20_reg[4]/P0001  & \sa20_reg[7]/NET0131  ;
  assign n715 = n690 & n714 ;
  assign n728 = ~\sa20_reg[5]/P0001  & n693 ;
  assign n729 = \sa20_reg[3]/P0001  & n714 ;
  assign n730 = ~n728 & ~n729 ;
  assign n731 = \sa20_reg[2]/P0001  & ~n730 ;
  assign n732 = ~n715 & ~n731 ;
  assign n733 = ~n727 & n732 ;
  assign n734 = ~\sa20_reg[1]/P0001  & ~n733 ;
  assign n691 = ~\sa20_reg[3]/P0001  & \sa20_reg[4]/P0001  ;
  assign n692 = n690 & n691 ;
  assign n695 = n693 & n694 ;
  assign n696 = ~n692 & ~n695 ;
  assign n697 = ~\sa20_reg[2]/P0001  & ~n696 ;
  assign n698 = \sa20_reg[3]/P0001  & \sa20_reg[6]/NET0131  ;
  assign n699 = ~\sa20_reg[7]/NET0131  & n698 ;
  assign n700 = \sa20_reg[4]/P0001  & n699 ;
  assign n701 = \sa20_reg[5]/P0001  & \sa20_reg[6]/NET0131  ;
  assign n702 = n691 & n701 ;
  assign n703 = \sa20_reg[7]/NET0131  & n702 ;
  assign n704 = ~n700 & ~n703 ;
  assign n706 = \sa20_reg[3]/P0001  & ~\sa20_reg[5]/P0001  ;
  assign n707 = n705 & n706 ;
  assign n708 = ~\sa20_reg[5]/P0001  & ~\sa20_reg[6]/NET0131  ;
  assign n709 = ~\sa20_reg[4]/P0001  & ~\sa20_reg[7]/NET0131  ;
  assign n710 = n708 & n709 ;
  assign n711 = ~n707 & ~n710 ;
  assign n712 = n704 & n711 ;
  assign n713 = \sa20_reg[2]/P0001  & ~n712 ;
  assign n757 = ~n697 & ~n713 ;
  assign n758 = ~n734 & n757 ;
  assign n759 = ~n756 & n758 ;
  assign n760 = \sa20_reg[0]/P0001  & ~n759 ;
  assign n771 = ~\sa20_reg[1]/P0001  & ~n695 ;
  assign n763 = ~\sa20_reg[2]/P0001  & \sa20_reg[3]/P0001  ;
  assign n764 = n714 & n763 ;
  assign n765 = ~\sa20_reg[4]/P0001  & \sa20_reg[7]/NET0131  ;
  assign n766 = n706 & n765 ;
  assign n772 = ~n764 & ~n766 ;
  assign n773 = n771 & n772 ;
  assign n769 = ~\sa20_reg[6]/NET0131  & n736 ;
  assign n770 = ~\sa20_reg[4]/P0001  & n769 ;
  assign n761 = \sa20_reg[2]/P0001  & \sa20_reg[3]/P0001  ;
  assign n762 = n724 & n761 ;
  assign n767 = \sa20_reg[4]/P0001  & n735 ;
  assign n768 = n736 & n767 ;
  assign n774 = ~n762 & ~n768 ;
  assign n775 = ~n770 & n774 ;
  assign n776 = n773 & n775 ;
  assign n781 = \sa20_reg[4]/P0001  & n744 ;
  assign n782 = ~\sa20_reg[4]/P0001  & n717 ;
  assign n783 = ~n781 & ~n782 ;
  assign n780 = ~\sa20_reg[2]/P0001  & ~n710 ;
  assign n784 = ~n761 & ~n780 ;
  assign n785 = ~n783 & n784 ;
  assign n777 = \sa20_reg[5]/P0001  & ~\sa20_reg[7]/NET0131  ;
  assign n778 = n698 & n777 ;
  assign n779 = \sa20_reg[4]/P0001  & n778 ;
  assign n786 = \sa20_reg[1]/P0001  & ~n779 ;
  assign n787 = ~n785 & n786 ;
  assign n788 = ~n776 & ~n787 ;
  assign n791 = \sa20_reg[4]/P0001  & n708 ;
  assign n792 = n706 & ~n723 ;
  assign n793 = ~n791 & ~n792 ;
  assign n794 = ~n716 & ~n793 ;
  assign n789 = ~\sa20_reg[7]/NET0131  & n691 ;
  assign n790 = n701 & n789 ;
  assign n795 = n698 & n720 ;
  assign n796 = ~\sa20_reg[2]/P0001  & ~n795 ;
  assign n797 = ~n790 & n796 ;
  assign n798 = ~n794 & n797 ;
  assign n799 = ~\sa20_reg[3]/P0001  & ~\sa20_reg[4]/P0001  ;
  assign n800 = n708 & n799 ;
  assign n801 = \sa20_reg[2]/P0001  & ~n800 ;
  assign n802 = ~n768 & n801 ;
  assign n803 = ~n798 & ~n802 ;
  assign n804 = ~n788 & ~n803 ;
  assign n805 = ~\sa20_reg[0]/P0001  & ~n804 ;
  assign n826 = \sa20_reg[6]/NET0131  & \sa20_reg[7]/NET0131  ;
  assign n827 = n694 & n826 ;
  assign n828 = \sa20_reg[2]/P0001  & ~n827 ;
  assign n829 = n723 & n745 ;
  assign n830 = n828 & ~n829 ;
  assign n833 = \sa20_reg[3]/P0001  & n744 ;
  assign n834 = ~\sa20_reg[6]/NET0131  & n833 ;
  assign n831 = ~\sa20_reg[2]/P0001  & ~n715 ;
  assign n832 = ~\sa20_reg[5]/P0001  & n739 ;
  assign n835 = n831 & ~n832 ;
  assign n836 = ~n834 & n835 ;
  assign n837 = ~n830 & ~n836 ;
  assign n838 = n701 & n799 ;
  assign n839 = n705 & n716 ;
  assign n840 = ~n838 & ~n839 ;
  assign n841 = ~n837 & n840 ;
  assign n842 = ~\sa20_reg[1]/P0001  & ~n841 ;
  assign n806 = \sa20_reg[1]/P0001  & \sa20_reg[2]/P0001  ;
  assign n810 = \sa20_reg[5]/P0001  & n745 ;
  assign n811 = n705 & n810 ;
  assign n807 = \sa20_reg[4]/P0001  & n723 ;
  assign n808 = ~\sa20_reg[5]/P0001  & n807 ;
  assign n809 = n723 & n799 ;
  assign n812 = ~n808 & ~n809 ;
  assign n813 = ~n811 & n812 ;
  assign n814 = n806 & ~n813 ;
  assign n825 = n715 & n763 ;
  assign n819 = \sa20_reg[2]/P0001  & ~\sa20_reg[3]/P0001  ;
  assign n820 = ~\sa20_reg[5]/P0001  & n723 ;
  assign n821 = n819 & n820 ;
  assign n824 = ~\sa20_reg[7]/NET0131  & n800 ;
  assign n843 = ~n821 & ~n824 ;
  assign n844 = ~n825 & n843 ;
  assign n815 = \sa20_reg[1]/P0001  & ~\sa20_reg[2]/P0001  ;
  assign n816 = ~\sa20_reg[6]/NET0131  & n745 ;
  assign n817 = n777 & n816 ;
  assign n818 = n815 & n817 ;
  assign n822 = n716 & n728 ;
  assign n823 = \sa20_reg[2]/P0001  & n822 ;
  assign n845 = ~n818 & ~n823 ;
  assign n846 = n844 & n845 ;
  assign n847 = ~n814 & n846 ;
  assign n848 = ~n842 & n847 ;
  assign n849 = ~n805 & n848 ;
  assign n850 = ~n760 & n849 ;
  assign n851 = n689 & ~n850 ;
  assign n852 = ~n689 & n850 ;
  assign n853 = ~n851 & ~n852 ;
  assign n861 = \sa13_reg[5]/P0001  & n543 ;
  assign n862 = ~\sa13_reg[3]/P0001  & n861 ;
  assign n863 = ~\sa13_reg[4]/P0001  & n862 ;
  assign n854 = n550 & n556 ;
  assign n870 = ~n569 & ~n854 ;
  assign n855 = ~\sa13_reg[5]/P0001  & n583 ;
  assign n856 = ~\sa13_reg[3]/P0001  & n855 ;
  assign n857 = \sa13_reg[7]/NET0131  & n608 ;
  assign n871 = ~n856 & ~n857 ;
  assign n872 = n870 & n871 ;
  assign n873 = ~n863 & n872 ;
  assign n858 = \sa13_reg[5]/P0001  & n567 ;
  assign n859 = ~n560 & ~n858 ;
  assign n860 = \sa13_reg[2]/P0001  & ~n859 ;
  assign n865 = ~\sa13_reg[4]/P0001  & n543 ;
  assign n866 = ~\sa13_reg[3]/P0001  & n865 ;
  assign n864 = \sa13_reg[3]/P0001  & n549 ;
  assign n867 = ~n534 & ~n864 ;
  assign n868 = ~n866 & n867 ;
  assign n869 = ~\sa13_reg[2]/P0001  & ~n868 ;
  assign n874 = ~n860 & ~n869 ;
  assign n875 = n873 & n874 ;
  assign n876 = \sa13_reg[1]/P0001  & ~n875 ;
  assign n883 = \sa13_reg[2]/P0001  & n655 ;
  assign n884 = \sa13_reg[7]/NET0131  & n533 ;
  assign n885 = ~n883 & ~n884 ;
  assign n886 = n547 & ~n885 ;
  assign n887 = \sa13_reg[2]/P0001  & n650 ;
  assign n888 = n559 & n563 ;
  assign n889 = ~n887 & ~n888 ;
  assign n890 = ~\sa13_reg[3]/P0001  & ~n889 ;
  assign n891 = ~n886 & ~n890 ;
  assign n892 = ~\sa13_reg[1]/P0001  & ~n891 ;
  assign n877 = ~\sa13_reg[3]/P0001  & n591 ;
  assign n878 = ~n604 & ~n877 ;
  assign n879 = ~n653 & ~n878 ;
  assign n880 = ~n672 & ~n857 ;
  assign n881 = ~n879 & n880 ;
  assign n882 = \sa13_reg[2]/P0001  & ~n881 ;
  assign n893 = ~\sa13_reg[2]/P0001  & n588 ;
  assign n894 = ~n548 & ~n893 ;
  assign n895 = n586 & n894 ;
  assign n896 = ~n882 & n895 ;
  assign n897 = ~n892 & n896 ;
  assign n898 = ~n876 & n897 ;
  assign n899 = ~\sa13_reg[0]/P0001  & ~n898 ;
  assign n902 = \sa13_reg[3]/P0001  & n861 ;
  assign n932 = ~n542 & ~n902 ;
  assign n926 = ~n551 & ~n861 ;
  assign n927 = ~\sa13_reg[2]/P0001  & ~n926 ;
  assign n912 = ~\sa13_reg[5]/P0001  & \sa13_reg[6]/NET0131  ;
  assign n928 = ~\sa13_reg[4]/P0001  & n912 ;
  assign n929 = n555 & n556 ;
  assign n930 = ~n928 & ~n929 ;
  assign n931 = \sa13_reg[2]/P0001  & ~n930 ;
  assign n933 = ~n927 & ~n931 ;
  assign n934 = n932 & n933 ;
  assign n935 = ~\sa13_reg[1]/P0001  & ~n934 ;
  assign n918 = ~\sa13_reg[3]/P0001  & n652 ;
  assign n920 = ~\sa13_reg[3]/P0001  & n532 ;
  assign n921 = n587 & n920 ;
  assign n919 = ~\sa13_reg[4]/P0001  & n864 ;
  assign n922 = ~n558 & ~n919 ;
  assign n923 = ~n921 & n922 ;
  assign n924 = ~n918 & n923 ;
  assign n925 = \sa13_reg[1]/P0001  & ~n924 ;
  assign n900 = \sa13_reg[5]/P0001  & ~\sa13_reg[7]/NET0131  ;
  assign n901 = ~\sa13_reg[4]/P0001  & n900 ;
  assign n903 = ~\sa13_reg[4]/P0001  & n544 ;
  assign n904 = ~n902 & ~n903 ;
  assign n905 = ~n901 & n904 ;
  assign n906 = ~\sa13_reg[2]/P0001  & ~n905 ;
  assign n915 = ~n580 & ~n610 ;
  assign n916 = ~n656 & n915 ;
  assign n917 = n680 & ~n916 ;
  assign n907 = n535 & n587 ;
  assign n908 = n563 & n579 ;
  assign n909 = ~n907 & ~n908 ;
  assign n910 = n603 & ~n909 ;
  assign n911 = \sa13_reg[3]/P0001  & n537 ;
  assign n913 = n587 & n912 ;
  assign n914 = ~\sa13_reg[2]/P0001  & n913 ;
  assign n936 = ~n911 & ~n914 ;
  assign n937 = ~n910 & n936 ;
  assign n938 = ~n917 & n937 ;
  assign n939 = ~n906 & n938 ;
  assign n940 = ~n925 & n939 ;
  assign n941 = ~n935 & n940 ;
  assign n942 = \sa13_reg[0]/P0001  & ~n941 ;
  assign n943 = ~n543 & ~n549 ;
  assign n944 = ~\sa13_reg[5]/P0001  & ~n943 ;
  assign n945 = n533 & n944 ;
  assign n946 = ~\sa13_reg[6]/NET0131  & n555 ;
  assign n947 = \sa13_reg[5]/P0001  & n946 ;
  assign n948 = ~n542 & ~n947 ;
  assign n949 = ~n945 & n948 ;
  assign n950 = \sa13_reg[2]/P0001  & ~n949 ;
  assign n951 = ~n654 & ~n950 ;
  assign n952 = ~\sa13_reg[1]/P0001  & ~n951 ;
  assign n962 = ~\sa13_reg[1]/P0001  & ~\sa13_reg[2]/P0001  ;
  assign n963 = ~\sa13_reg[3]/P0001  & n559 ;
  assign n964 = ~\sa13_reg[4]/P0001  & n963 ;
  assign n965 = ~n609 & ~n913 ;
  assign n966 = ~n964 & n965 ;
  assign n967 = n962 & ~n966 ;
  assign n954 = n603 & n858 ;
  assign n955 = \sa13_reg[3]/P0001  & n547 ;
  assign n956 = n536 & n955 ;
  assign n957 = ~n893 & ~n956 ;
  assign n958 = ~n954 & n957 ;
  assign n959 = \sa13_reg[1]/P0001  & ~n958 ;
  assign n953 = \sa13_reg[4]/P0001  & n624 ;
  assign n960 = ~n681 & ~n856 ;
  assign n961 = ~\sa13_reg[2]/P0001  & ~n960 ;
  assign n968 = ~n953 & ~n961 ;
  assign n969 = ~n959 & n968 ;
  assign n970 = ~n967 & n969 ;
  assign n971 = ~n952 & n970 ;
  assign n972 = ~n942 & n971 ;
  assign n973 = ~n899 & n972 ;
  assign n1011 = ~\sa02_reg[5]/P0001  & \sa02_reg[6]/NET0131  ;
  assign n1090 = ~\sa02_reg[4]/P0001  & n1011 ;
  assign n979 = ~\sa02_reg[6]/NET0131  & ~\sa02_reg[7]/NET0131  ;
  assign n1038 = \sa02_reg[3]/P0001  & \sa02_reg[4]/P0001  ;
  assign n1091 = n979 & n1038 ;
  assign n1092 = ~n1090 & ~n1091 ;
  assign n1093 = \sa02_reg[2]/P0001  & ~n1092 ;
  assign n1023 = ~\sa02_reg[6]/NET0131  & \sa02_reg[7]/NET0131  ;
  assign n1094 = ~\sa02_reg[5]/P0001  & n1023 ;
  assign n1095 = ~\sa02_reg[2]/P0001  & \sa02_reg[3]/P0001  ;
  assign n1096 = n1094 & n1095 ;
  assign n975 = \sa02_reg[5]/P0001  & \sa02_reg[6]/NET0131  ;
  assign n976 = \sa02_reg[7]/NET0131  & n975 ;
  assign n986 = ~\sa02_reg[3]/P0001  & \sa02_reg[4]/P0001  ;
  assign n1071 = n976 & n986 ;
  assign n978 = \sa02_reg[2]/P0001  & ~\sa02_reg[3]/P0001  ;
  assign n1025 = \sa02_reg[6]/NET0131  & ~\sa02_reg[7]/NET0131  ;
  assign n1088 = \sa02_reg[5]/P0001  & n1025 ;
  assign n1089 = ~n978 & n1088 ;
  assign n1097 = ~n1071 & ~n1089 ;
  assign n1098 = ~n1096 & n1097 ;
  assign n1099 = ~n1093 & n1098 ;
  assign n1100 = ~\sa02_reg[1]/P0001  & ~n1099 ;
  assign n1059 = \sa02_reg[3]/P0001  & ~\sa02_reg[4]/P0001  ;
  assign n1078 = \sa02_reg[5]/P0001  & n1059 ;
  assign n982 = ~\sa02_reg[5]/P0001  & ~\sa02_reg[6]/NET0131  ;
  assign n983 = ~\sa02_reg[4]/P0001  & n982 ;
  assign n1006 = \sa02_reg[4]/P0001  & ~\sa02_reg[7]/NET0131  ;
  assign n1007 = ~\sa02_reg[5]/P0001  & n1006 ;
  assign n1079 = ~n983 & ~n1007 ;
  assign n1080 = ~n1078 & n1079 ;
  assign n1081 = \sa02_reg[1]/P0001  & ~n1080 ;
  assign n1015 = ~\sa02_reg[4]/P0001  & ~\sa02_reg[7]/NET0131  ;
  assign n1068 = \sa02_reg[3]/P0001  & \sa02_reg[6]/NET0131  ;
  assign n1069 = n1015 & n1068 ;
  assign n1056 = \sa02_reg[5]/P0001  & ~\sa02_reg[7]/NET0131  ;
  assign n1082 = n1056 & n1068 ;
  assign n1083 = ~n1069 & ~n1082 ;
  assign n1084 = ~\sa02_reg[4]/P0001  & n1056 ;
  assign n1085 = n1083 & ~n1084 ;
  assign n1086 = ~n1081 & n1085 ;
  assign n1087 = ~\sa02_reg[2]/P0001  & ~n1086 ;
  assign n1057 = n1038 & n1056 ;
  assign n1058 = ~\sa02_reg[6]/NET0131  & n1057 ;
  assign n1060 = n1023 & n1059 ;
  assign n1064 = ~n1058 & ~n1060 ;
  assign n987 = n982 & n986 ;
  assign n1061 = ~\sa02_reg[7]/NET0131  & n987 ;
  assign n1000 = \sa02_reg[4]/P0001  & \sa02_reg[7]/NET0131  ;
  assign n999 = \sa02_reg[5]/P0001  & ~\sa02_reg[6]/NET0131  ;
  assign n1062 = ~\sa02_reg[3]/P0001  & n999 ;
  assign n1063 = n1000 & n1062 ;
  assign n1065 = ~n1061 & ~n1063 ;
  assign n1066 = n1064 & n1065 ;
  assign n1067 = \sa02_reg[1]/P0001  & ~n1066 ;
  assign n995 = ~\sa02_reg[5]/P0001  & ~\sa02_reg[7]/NET0131  ;
  assign n1004 = ~\sa02_reg[4]/P0001  & \sa02_reg[6]/NET0131  ;
  assign n1072 = n995 & n1004 ;
  assign n1073 = ~\sa02_reg[3]/P0001  & n1072 ;
  assign n1074 = ~n1071 & ~n1073 ;
  assign n1075 = \sa02_reg[2]/P0001  & ~n1074 ;
  assign n1070 = \sa02_reg[5]/P0001  & n1069 ;
  assign n1076 = n1000 & n1011 ;
  assign n1077 = ~\sa02_reg[2]/P0001  & n1076 ;
  assign n1101 = ~n1070 & ~n1077 ;
  assign n1102 = ~n1075 & n1101 ;
  assign n1103 = ~n1067 & n1102 ;
  assign n1104 = ~n1087 & n1103 ;
  assign n1105 = ~n1100 & n1104 ;
  assign n1106 = \sa02_reg[0]/P0001  & ~n1105 ;
  assign n1022 = n986 & n999 ;
  assign n1027 = ~\sa02_reg[2]/P0001  & ~n1022 ;
  assign n1024 = \sa02_reg[3]/P0001  & n1023 ;
  assign n974 = ~\sa02_reg[3]/P0001  & ~\sa02_reg[4]/P0001  ;
  assign n1026 = n974 & n1025 ;
  assign n1028 = ~n1024 & ~n1026 ;
  assign n1029 = n1027 & n1028 ;
  assign n1031 = n975 & n1006 ;
  assign n993 = \sa02_reg[5]/P0001  & \sa02_reg[7]/NET0131  ;
  assign n1030 = \sa02_reg[3]/P0001  & n993 ;
  assign n1032 = \sa02_reg[2]/P0001  & ~n1030 ;
  assign n1033 = ~n1031 & n1032 ;
  assign n1034 = ~n1029 & ~n1033 ;
  assign n1039 = \sa02_reg[7]/NET0131  & n1038 ;
  assign n1040 = ~n1026 & ~n1039 ;
  assign n1041 = \sa02_reg[5]/P0001  & ~n1040 ;
  assign n1042 = \sa02_reg[5]/P0001  & n1023 ;
  assign n1043 = ~\sa02_reg[4]/P0001  & n1042 ;
  assign n1019 = \sa02_reg[6]/NET0131  & \sa02_reg[7]/NET0131  ;
  assign n1020 = ~\sa02_reg[5]/P0001  & n1019 ;
  assign n1021 = ~\sa02_reg[3]/P0001  & n1020 ;
  assign n1035 = \sa02_reg[3]/P0001  & ~\sa02_reg[5]/P0001  ;
  assign n1036 = ~\sa02_reg[6]/NET0131  & n1035 ;
  assign n1037 = ~\sa02_reg[7]/NET0131  & n1036 ;
  assign n1044 = ~n1021 & ~n1037 ;
  assign n1045 = ~n1043 & n1044 ;
  assign n1046 = ~n1041 & n1045 ;
  assign n1047 = ~n1034 & n1046 ;
  assign n1048 = \sa02_reg[1]/P0001  & ~n1047 ;
  assign n977 = n974 & n976 ;
  assign n980 = ~\sa02_reg[5]/P0001  & n979 ;
  assign n981 = n978 & n980 ;
  assign n989 = ~n977 & ~n981 ;
  assign n984 = \sa02_reg[2]/P0001  & \sa02_reg[3]/P0001  ;
  assign n985 = n983 & n984 ;
  assign n988 = \sa02_reg[7]/NET0131  & n987 ;
  assign n990 = ~n985 & ~n988 ;
  assign n991 = n989 & n990 ;
  assign n992 = ~\sa02_reg[1]/P0001  & ~n991 ;
  assign n1003 = ~\sa02_reg[5]/P0001  & \sa02_reg[7]/NET0131  ;
  assign n1005 = n1003 & n1004 ;
  assign n1008 = \sa02_reg[3]/P0001  & n1007 ;
  assign n1009 = ~n1005 & ~n1008 ;
  assign n1010 = ~\sa02_reg[2]/P0001  & ~n1009 ;
  assign n1012 = n986 & n1011 ;
  assign n1013 = \sa02_reg[2]/P0001  & n1012 ;
  assign n1014 = ~\sa02_reg[7]/NET0131  & n1013 ;
  assign n994 = \sa02_reg[4]/P0001  & n993 ;
  assign n996 = ~\sa02_reg[4]/P0001  & n995 ;
  assign n997 = ~n994 & ~n996 ;
  assign n998 = n984 & ~n997 ;
  assign n1001 = n999 & n1000 ;
  assign n1002 = ~\sa02_reg[2]/P0001  & n1001 ;
  assign n1016 = \sa02_reg[2]/P0001  & ~\sa02_reg[6]/NET0131  ;
  assign n1017 = ~n982 & ~n1016 ;
  assign n1018 = n1015 & ~n1017 ;
  assign n1049 = ~n1002 & ~n1018 ;
  assign n1050 = ~n998 & n1049 ;
  assign n1051 = ~n1014 & n1050 ;
  assign n1052 = ~n1010 & n1051 ;
  assign n1053 = ~n992 & n1052 ;
  assign n1054 = ~n1048 & n1053 ;
  assign n1055 = ~\sa02_reg[0]/P0001  & ~n1054 ;
  assign n1122 = \sa02_reg[7]/NET0131  & n974 ;
  assign n1123 = n1025 & n1038 ;
  assign n1124 = ~n1122 & ~n1123 ;
  assign n1125 = \sa02_reg[5]/P0001  & ~n1124 ;
  assign n1126 = ~n1076 & ~n1125 ;
  assign n1127 = ~\sa02_reg[2]/P0001  & ~n1126 ;
  assign n1121 = n974 & n979 ;
  assign n1130 = ~\sa02_reg[5]/P0001  & n1025 ;
  assign n1131 = ~n1094 & ~n1130 ;
  assign n1132 = ~\sa02_reg[3]/P0001  & ~n976 ;
  assign n1133 = n1131 & n1132 ;
  assign n1128 = \sa02_reg[2]/P0001  & \sa02_reg[4]/P0001  ;
  assign n1129 = \sa02_reg[3]/P0001  & ~n999 ;
  assign n1134 = n1128 & ~n1129 ;
  assign n1135 = ~n1133 & n1134 ;
  assign n1136 = ~n1121 & ~n1135 ;
  assign n1137 = ~n1127 & n1136 ;
  assign n1138 = ~\sa02_reg[1]/P0001  & ~n1137 ;
  assign n1107 = \sa02_reg[2]/P0001  & ~n1058 ;
  assign n1108 = ~\sa02_reg[2]/P0001  & ~n1021 ;
  assign n1109 = ~\sa02_reg[6]/NET0131  & n1059 ;
  assign n1110 = n1056 & n1109 ;
  assign n1111 = n1108 & ~n1110 ;
  assign n1112 = ~n1107 & ~n1111 ;
  assign n1113 = n978 & n1025 ;
  assign n1114 = \sa02_reg[4]/P0001  & n1113 ;
  assign n1115 = \sa02_reg[5]/P0001  & n1114 ;
  assign n1116 = n979 & n1059 ;
  assign n1117 = ~\sa02_reg[5]/P0001  & n1116 ;
  assign n1118 = ~n1002 & ~n1117 ;
  assign n1119 = ~n1115 & n1118 ;
  assign n1120 = \sa02_reg[1]/P0001  & ~n1119 ;
  assign n1139 = ~n1112 & ~n1120 ;
  assign n1140 = ~n1138 & n1139 ;
  assign n1141 = ~n1055 & n1140 ;
  assign n1142 = ~n1106 & n1141 ;
  assign n1143 = ~n973 & ~n1142 ;
  assign n1144 = n973 & n1142 ;
  assign n1145 = ~n1143 & ~n1144 ;
  assign n1151 = ~\sa31_reg[5]/P0001  & \sa31_reg[6]/NET0131  ;
  assign n1152 = ~\sa31_reg[3]/P0001  & ~\sa31_reg[4]/P0001  ;
  assign n1153 = \sa31_reg[7]/P0001  & n1152 ;
  assign n1154 = n1151 & n1153 ;
  assign n1146 = ~\sa31_reg[6]/NET0131  & \sa31_reg[7]/P0001  ;
  assign n1147 = \sa31_reg[5]/P0001  & n1146 ;
  assign n1148 = ~\sa31_reg[4]/P0001  & n1147 ;
  assign n1149 = \sa31_reg[6]/NET0131  & ~\sa31_reg[7]/P0001  ;
  assign n1150 = \sa31_reg[4]/P0001  & n1149 ;
  assign n1155 = ~n1148 & ~n1150 ;
  assign n1156 = ~n1154 & n1155 ;
  assign n1157 = \sa31_reg[2]/P0001  & ~n1156 ;
  assign n1166 = \sa31_reg[5]/P0001  & \sa31_reg[7]/P0001  ;
  assign n1167 = \sa31_reg[3]/P0001  & n1166 ;
  assign n1168 = ~\sa31_reg[4]/P0001  & n1167 ;
  assign n1158 = \sa31_reg[5]/P0001  & ~\sa31_reg[7]/P0001  ;
  assign n1159 = \sa31_reg[3]/P0001  & \sa31_reg[4]/P0001  ;
  assign n1160 = ~\sa31_reg[6]/NET0131  & n1159 ;
  assign n1161 = n1158 & n1160 ;
  assign n1162 = ~\sa31_reg[2]/P0001  & ~\sa31_reg[3]/P0001  ;
  assign n1163 = ~\sa31_reg[4]/P0001  & \sa31_reg[6]/NET0131  ;
  assign n1164 = ~\sa31_reg[5]/P0001  & ~n1163 ;
  assign n1165 = n1162 & n1164 ;
  assign n1169 = ~n1161 & ~n1165 ;
  assign n1170 = ~n1168 & n1169 ;
  assign n1171 = ~n1157 & n1170 ;
  assign n1172 = \sa31_reg[1]/P0001  & ~n1171 ;
  assign n1180 = ~\sa31_reg[5]/P0001  & ~\sa31_reg[7]/P0001  ;
  assign n1181 = n1159 & n1180 ;
  assign n1182 = ~\sa31_reg[5]/P0001  & \sa31_reg[7]/P0001  ;
  assign n1183 = n1163 & n1182 ;
  assign n1184 = ~n1181 & ~n1183 ;
  assign n1185 = ~\sa31_reg[2]/P0001  & ~n1184 ;
  assign n1173 = ~\sa31_reg[5]/P0001  & n1149 ;
  assign n1174 = \sa31_reg[4]/P0001  & \sa31_reg[7]/P0001  ;
  assign n1175 = \sa31_reg[3]/P0001  & n1174 ;
  assign n1176 = ~n1173 & ~n1175 ;
  assign n1177 = \sa31_reg[2]/P0001  & ~n1176 ;
  assign n1178 = \sa31_reg[5]/P0001  & ~\sa31_reg[6]/NET0131  ;
  assign n1179 = n1174 & n1178 ;
  assign n1186 = ~\sa31_reg[6]/NET0131  & ~\sa31_reg[7]/P0001  ;
  assign n1187 = \sa31_reg[5]/P0001  & n1186 ;
  assign n1188 = n1162 & n1187 ;
  assign n1189 = ~n1179 & ~n1188 ;
  assign n1190 = ~n1177 & n1189 ;
  assign n1191 = ~n1185 & n1190 ;
  assign n1192 = ~\sa31_reg[1]/P0001  & ~n1191 ;
  assign n1193 = \sa31_reg[5]/P0001  & \sa31_reg[6]/NET0131  ;
  assign n1194 = ~\sa31_reg[7]/P0001  & n1193 ;
  assign n1195 = ~\sa31_reg[4]/P0001  & n1194 ;
  assign n1196 = ~\sa31_reg[3]/P0001  & \sa31_reg[4]/P0001  ;
  assign n1197 = n1178 & n1196 ;
  assign n1198 = ~n1195 & ~n1197 ;
  assign n1199 = ~\sa31_reg[2]/P0001  & ~n1198 ;
  assign n1200 = \sa31_reg[3]/P0001  & n1150 ;
  assign n1201 = \sa31_reg[6]/NET0131  & n1166 ;
  assign n1202 = n1196 & n1201 ;
  assign n1203 = ~n1200 & ~n1202 ;
  assign n1204 = ~\sa31_reg[4]/P0001  & n1180 ;
  assign n1205 = ~\sa31_reg[6]/NET0131  & n1204 ;
  assign n1206 = \sa31_reg[3]/P0001  & n1146 ;
  assign n1207 = ~\sa31_reg[5]/P0001  & n1206 ;
  assign n1208 = ~n1205 & ~n1207 ;
  assign n1209 = n1203 & n1208 ;
  assign n1210 = \sa31_reg[2]/P0001  & ~n1209 ;
  assign n1211 = ~n1199 & ~n1210 ;
  assign n1212 = ~n1192 & n1211 ;
  assign n1213 = ~n1172 & n1212 ;
  assign n1214 = \sa31_reg[0]/P0002  & ~n1213 ;
  assign n1265 = \sa31_reg[2]/P0001  & \sa31_reg[3]/P0001  ;
  assign n1266 = n1187 & n1265 ;
  assign n1222 = ~\sa31_reg[2]/P0001  & n1175 ;
  assign n1272 = ~\sa31_reg[1]/P0001  & ~n1222 ;
  assign n1273 = ~n1266 & n1272 ;
  assign n1225 = \sa31_reg[3]/P0001  & ~\sa31_reg[4]/P0001  ;
  assign n1260 = \sa31_reg[6]/NET0131  & n1196 ;
  assign n1267 = ~n1225 & ~n1260 ;
  assign n1268 = n1182 & ~n1267 ;
  assign n1269 = ~\sa31_reg[3]/P0001  & n1146 ;
  assign n1270 = ~n1194 & ~n1269 ;
  assign n1271 = ~\sa31_reg[4]/P0001  & ~n1270 ;
  assign n1274 = ~n1268 & ~n1271 ;
  assign n1275 = n1273 & n1274 ;
  assign n1283 = ~\sa31_reg[2]/P0001  & n1205 ;
  assign n1279 = \sa31_reg[2]/P0001  & ~\sa31_reg[3]/P0001  ;
  assign n1280 = \sa31_reg[4]/P0001  & n1166 ;
  assign n1281 = ~n1204 & ~n1280 ;
  assign n1282 = n1279 & ~n1281 ;
  assign n1276 = \sa31_reg[3]/P0001  & ~\sa31_reg[7]/P0001  ;
  assign n1277 = \sa31_reg[4]/P0001  & n1193 ;
  assign n1278 = n1276 & n1277 ;
  assign n1284 = \sa31_reg[1]/P0001  & ~n1278 ;
  assign n1285 = ~n1282 & n1284 ;
  assign n1286 = ~n1283 & n1285 ;
  assign n1287 = ~n1275 & ~n1286 ;
  assign n1261 = n1158 & n1260 ;
  assign n1229 = ~\sa31_reg[5]/P0001  & ~\sa31_reg[6]/NET0131  ;
  assign n1255 = n1196 & n1229 ;
  assign n1256 = \sa31_reg[6]/NET0131  & \sa31_reg[7]/P0001  ;
  assign n1257 = \sa31_reg[4]/P0001  & ~n1256 ;
  assign n1216 = \sa31_reg[3]/P0001  & ~\sa31_reg[5]/P0001  ;
  assign n1258 = ~n1186 & n1216 ;
  assign n1259 = ~n1257 & n1258 ;
  assign n1262 = ~n1255 & ~n1259 ;
  assign n1263 = ~n1261 & n1262 ;
  assign n1264 = ~\sa31_reg[2]/P0001  & ~n1263 ;
  assign n1288 = n1164 & n1279 ;
  assign n1289 = ~n1257 & n1288 ;
  assign n1290 = ~n1264 & ~n1289 ;
  assign n1291 = ~n1287 & n1290 ;
  assign n1292 = ~\sa31_reg[0]/P0002  & ~n1291 ;
  assign n1240 = \sa31_reg[5]/P0001  & n1206 ;
  assign n1239 = ~\sa31_reg[5]/P0001  & n1150 ;
  assign n1241 = ~n1179 & ~n1239 ;
  assign n1242 = ~n1240 & n1241 ;
  assign n1243 = ~\sa31_reg[2]/P0001  & ~n1242 ;
  assign n1244 = \sa31_reg[2]/P0001  & ~\sa31_reg[4]/P0001  ;
  assign n1248 = \sa31_reg[3]/P0001  & n1244 ;
  assign n1249 = n1186 & n1248 ;
  assign n1245 = n1201 & n1244 ;
  assign n1246 = n1146 & n1159 ;
  assign n1247 = n1152 & n1193 ;
  assign n1250 = ~n1246 & ~n1247 ;
  assign n1251 = ~n1245 & n1250 ;
  assign n1252 = ~n1249 & n1251 ;
  assign n1253 = ~n1243 & n1252 ;
  assign n1254 = ~\sa31_reg[1]/P0001  & ~n1253 ;
  assign n1232 = \sa31_reg[1]/P0001  & \sa31_reg[2]/P0001  ;
  assign n1235 = \sa31_reg[3]/P0001  & n1148 ;
  assign n1219 = ~\sa31_reg[5]/P0001  & n1186 ;
  assign n1233 = \sa31_reg[4]/P0001  & n1219 ;
  assign n1234 = n1152 & n1186 ;
  assign n1236 = ~n1233 & ~n1234 ;
  assign n1237 = ~n1235 & n1236 ;
  assign n1238 = n1232 & ~n1237 ;
  assign n1220 = ~\sa31_reg[3]/P0001  & n1219 ;
  assign n1221 = \sa31_reg[2]/P0001  & n1220 ;
  assign n1215 = \sa31_reg[2]/P0001  & \sa31_reg[4]/P0001  ;
  assign n1217 = n1149 & n1216 ;
  assign n1218 = n1215 & n1217 ;
  assign n1230 = ~\sa31_reg[7]/P0001  & n1152 ;
  assign n1231 = n1229 & n1230 ;
  assign n1293 = ~n1218 & ~n1231 ;
  assign n1294 = ~n1221 & n1293 ;
  assign n1223 = n1178 & n1222 ;
  assign n1224 = \sa31_reg[1]/P0001  & ~\sa31_reg[2]/P0001  ;
  assign n1226 = ~\sa31_reg[6]/NET0131  & n1225 ;
  assign n1227 = n1158 & n1226 ;
  assign n1228 = n1224 & n1227 ;
  assign n1295 = ~n1223 & ~n1228 ;
  assign n1296 = n1294 & n1295 ;
  assign n1297 = ~n1238 & n1296 ;
  assign n1298 = ~n1254 & n1297 ;
  assign n1299 = ~n1292 & n1298 ;
  assign n1300 = ~n1214 & n1299 ;
  assign n1301 = \u0_w_reg[2][30]/P0001  & ~n1300 ;
  assign n1302 = ~\u0_w_reg[2][30]/P0001  & n1300 ;
  assign n1303 = ~n1301 & ~n1302 ;
  assign n1304 = n1145 & n1303 ;
  assign n1305 = ~n1145 & ~n1303 ;
  assign n1306 = ~n1304 & ~n1305 ;
  assign n1308 = n853 & n1306 ;
  assign n1307 = ~n853 & ~n1306 ;
  assign n1309 = ~\ld_r_reg/P0001  & ~n1307 ;
  assign n1310 = ~n1308 & n1309 ;
  assign n1312 = ~\text_in_r_reg[62]/P0001  & \u0_w_reg[2][30]/P0001  ;
  assign n1311 = \text_in_r_reg[62]/P0001  & ~\u0_w_reg[2][30]/P0001  ;
  assign n1313 = \ld_r_reg/P0001  & ~n1311 ;
  assign n1314 = ~n1312 & n1313 ;
  assign n1315 = ~n1310 & ~n1314 ;
  assign n1318 = \sa03_reg[6]/NET0131  & ~\sa03_reg[7]/NET0131  ;
  assign n1435 = \sa03_reg[5]/P0001  & n1318 ;
  assign n1446 = \sa03_reg[3]/P0001  & n1435 ;
  assign n1383 = ~\sa03_reg[4]/P0001  & ~\sa03_reg[7]/NET0131  ;
  assign n1398 = \sa03_reg[3]/P0001  & \sa03_reg[6]/NET0131  ;
  assign n1447 = n1383 & n1398 ;
  assign n1448 = ~n1446 & ~n1447 ;
  assign n1326 = ~\sa03_reg[5]/P0001  & \sa03_reg[6]/NET0131  ;
  assign n1396 = \sa03_reg[4]/P0001  & n1326 ;
  assign n1397 = \sa03_reg[7]/NET0131  & n1396 ;
  assign n1449 = \sa03_reg[5]/P0001  & ~\sa03_reg[7]/NET0131  ;
  assign n1450 = ~\sa03_reg[4]/P0001  & n1449 ;
  assign n1451 = ~n1397 & ~n1450 ;
  assign n1452 = n1448 & n1451 ;
  assign n1453 = ~\sa03_reg[2]/P0001  & ~n1452 ;
  assign n1334 = ~\sa03_reg[3]/P0001  & \sa03_reg[4]/P0001  ;
  assign n1342 = \sa03_reg[5]/P0001  & \sa03_reg[6]/NET0131  ;
  assign n1353 = \sa03_reg[7]/NET0131  & n1342 ;
  assign n1438 = n1334 & n1353 ;
  assign n1319 = ~\sa03_reg[4]/P0001  & n1318 ;
  assign n1320 = ~\sa03_reg[3]/P0001  & n1319 ;
  assign n1443 = ~\sa03_reg[5]/P0001  & n1320 ;
  assign n1444 = ~n1438 & ~n1443 ;
  assign n1445 = \sa03_reg[2]/P0001  & ~n1444 ;
  assign n1423 = \sa03_reg[3]/P0001  & ~\sa03_reg[4]/P0001  ;
  assign n1454 = \sa03_reg[5]/P0001  & n1423 ;
  assign n1469 = n1318 & n1454 ;
  assign n1470 = ~n1445 & ~n1469 ;
  assign n1471 = ~n1453 & n1470 ;
  assign n1431 = ~\sa03_reg[4]/P0001  & n1326 ;
  assign n1316 = \sa03_reg[3]/P0001  & \sa03_reg[4]/P0001  ;
  assign n1323 = ~\sa03_reg[6]/NET0131  & ~\sa03_reg[7]/NET0131  ;
  assign n1432 = n1316 & n1323 ;
  assign n1433 = ~n1431 & ~n1432 ;
  assign n1434 = \sa03_reg[2]/P0001  & ~n1433 ;
  assign n1332 = ~\sa03_reg[6]/NET0131  & \sa03_reg[7]/NET0131  ;
  assign n1404 = ~\sa03_reg[5]/P0001  & n1332 ;
  assign n1429 = ~\sa03_reg[2]/P0001  & \sa03_reg[3]/P0001  ;
  assign n1430 = n1404 & n1429 ;
  assign n1436 = \sa03_reg[2]/P0001  & ~\sa03_reg[3]/P0001  ;
  assign n1437 = n1435 & ~n1436 ;
  assign n1439 = ~n1430 & ~n1437 ;
  assign n1440 = ~n1438 & n1439 ;
  assign n1441 = ~n1434 & n1440 ;
  assign n1442 = ~\sa03_reg[1]/P0001  & ~n1441 ;
  assign n1355 = ~\sa03_reg[5]/P0001  & ~\sa03_reg[6]/NET0131  ;
  assign n1455 = ~\sa03_reg[4]/P0001  & n1355 ;
  assign n1341 = \sa03_reg[4]/P0001  & ~\sa03_reg[7]/NET0131  ;
  assign n1370 = ~\sa03_reg[5]/P0001  & n1341 ;
  assign n1456 = ~n1370 & ~n1454 ;
  assign n1457 = ~n1455 & n1456 ;
  assign n1458 = ~\sa03_reg[2]/P0001  & ~n1457 ;
  assign n1459 = \sa03_reg[5]/P0001  & n1432 ;
  assign n1463 = n1332 & n1423 ;
  assign n1464 = ~n1459 & ~n1463 ;
  assign n1460 = ~\sa03_reg[7]/NET0131  & n1355 ;
  assign n1461 = n1334 & n1460 ;
  assign n1339 = \sa03_reg[5]/P0001  & \sa03_reg[7]/NET0131  ;
  assign n1375 = \sa03_reg[4]/P0001  & n1339 ;
  assign n1408 = ~\sa03_reg[3]/P0001  & ~\sa03_reg[6]/NET0131  ;
  assign n1462 = n1375 & n1408 ;
  assign n1465 = ~n1461 & ~n1462 ;
  assign n1466 = n1464 & n1465 ;
  assign n1467 = ~n1458 & n1466 ;
  assign n1468 = \sa03_reg[1]/P0001  & ~n1467 ;
  assign n1472 = ~n1442 & ~n1468 ;
  assign n1473 = n1471 & n1472 ;
  assign n1474 = \sa03_reg[0]/P0001  & ~n1473 ;
  assign n1329 = \sa03_reg[5]/P0001  & ~\sa03_reg[6]/NET0131  ;
  assign n1335 = n1329 & n1334 ;
  assign n1333 = \sa03_reg[3]/P0001  & n1332 ;
  assign n1336 = ~\sa03_reg[2]/P0001  & ~n1333 ;
  assign n1337 = ~n1335 & n1336 ;
  assign n1338 = ~n1320 & n1337 ;
  assign n1343 = n1341 & n1342 ;
  assign n1340 = \sa03_reg[3]/P0001  & n1339 ;
  assign n1344 = \sa03_reg[2]/P0001  & ~n1340 ;
  assign n1345 = ~n1343 & n1344 ;
  assign n1346 = ~n1338 & ~n1345 ;
  assign n1317 = \sa03_reg[7]/NET0131  & n1316 ;
  assign n1321 = ~n1317 & ~n1320 ;
  assign n1322 = \sa03_reg[5]/P0001  & ~n1321 ;
  assign n1330 = ~\sa03_reg[4]/P0001  & \sa03_reg[7]/NET0131  ;
  assign n1331 = n1329 & n1330 ;
  assign n1324 = \sa03_reg[3]/P0001  & ~\sa03_reg[5]/P0001  ;
  assign n1325 = n1323 & n1324 ;
  assign n1327 = ~\sa03_reg[3]/P0001  & \sa03_reg[7]/NET0131  ;
  assign n1328 = n1326 & n1327 ;
  assign n1347 = ~n1325 & ~n1328 ;
  assign n1348 = ~n1331 & n1347 ;
  assign n1349 = ~n1322 & n1348 ;
  assign n1350 = ~n1346 & n1349 ;
  assign n1351 = \sa03_reg[1]/P0001  & ~n1350 ;
  assign n1359 = n1327 & n1355 ;
  assign n1360 = \sa03_reg[4]/P0001  & n1359 ;
  assign n1352 = ~\sa03_reg[3]/P0001  & ~\sa03_reg[4]/P0001  ;
  assign n1354 = n1352 & n1353 ;
  assign n1356 = \sa03_reg[2]/P0001  & ~n1316 ;
  assign n1357 = ~n1327 & n1355 ;
  assign n1358 = n1356 & n1357 ;
  assign n1361 = ~n1354 & ~n1358 ;
  assign n1362 = ~n1360 & n1361 ;
  assign n1363 = ~\sa03_reg[1]/P0001  & ~n1362 ;
  assign n1367 = ~\sa03_reg[5]/P0001  & \sa03_reg[7]/NET0131  ;
  assign n1368 = ~\sa03_reg[4]/P0001  & \sa03_reg[6]/NET0131  ;
  assign n1369 = n1367 & n1368 ;
  assign n1371 = \sa03_reg[3]/P0001  & n1370 ;
  assign n1372 = ~n1369 & ~n1371 ;
  assign n1373 = ~\sa03_reg[2]/P0001  & ~n1372 ;
  assign n1374 = \sa03_reg[2]/P0001  & \sa03_reg[3]/P0001  ;
  assign n1376 = ~\sa03_reg[5]/P0001  & ~\sa03_reg[7]/NET0131  ;
  assign n1377 = ~\sa03_reg[4]/P0001  & n1376 ;
  assign n1378 = ~n1375 & ~n1377 ;
  assign n1379 = n1374 & ~n1378 ;
  assign n1364 = \sa03_reg[4]/P0001  & n1329 ;
  assign n1365 = \sa03_reg[7]/NET0131  & n1364 ;
  assign n1366 = ~\sa03_reg[2]/P0001  & n1365 ;
  assign n1380 = ~\sa03_reg[5]/P0001  & n1318 ;
  assign n1381 = \sa03_reg[2]/P0001  & n1334 ;
  assign n1382 = n1380 & n1381 ;
  assign n1384 = \sa03_reg[2]/P0001  & ~\sa03_reg[6]/NET0131  ;
  assign n1385 = ~n1355 & ~n1384 ;
  assign n1386 = n1383 & ~n1385 ;
  assign n1387 = ~n1382 & ~n1386 ;
  assign n1388 = ~n1366 & n1387 ;
  assign n1389 = ~n1379 & n1388 ;
  assign n1390 = ~n1373 & n1389 ;
  assign n1391 = ~n1363 & n1390 ;
  assign n1392 = ~n1351 & n1391 ;
  assign n1393 = ~\sa03_reg[0]/P0001  & ~n1392 ;
  assign n1399 = n1341 & n1398 ;
  assign n1400 = \sa03_reg[5]/P0001  & n1399 ;
  assign n1395 = n1339 & n1352 ;
  assign n1401 = ~n1395 & ~n1397 ;
  assign n1402 = ~n1400 & n1401 ;
  assign n1403 = ~\sa03_reg[2]/P0001  & ~n1402 ;
  assign n1405 = ~n1380 & ~n1404 ;
  assign n1406 = ~n1353 & n1405 ;
  assign n1407 = n1381 & ~n1406 ;
  assign n1394 = n1364 & n1374 ;
  assign n1409 = n1383 & n1408 ;
  assign n1410 = ~n1394 & ~n1409 ;
  assign n1411 = ~n1407 & n1410 ;
  assign n1412 = ~n1403 & n1411 ;
  assign n1413 = ~\sa03_reg[1]/P0001  & ~n1412 ;
  assign n1420 = n1334 & n1342 ;
  assign n1421 = ~\sa03_reg[7]/NET0131  & n1420 ;
  assign n1422 = \sa03_reg[2]/P0001  & n1421 ;
  assign n1424 = ~\sa03_reg[6]/NET0131  & n1423 ;
  assign n1425 = n1376 & n1424 ;
  assign n1426 = ~n1366 & ~n1425 ;
  assign n1427 = ~n1422 & n1426 ;
  assign n1428 = \sa03_reg[1]/P0001  & ~n1427 ;
  assign n1414 = n1329 & n1341 ;
  assign n1415 = n1374 & n1414 ;
  assign n1416 = n1329 & n1383 ;
  assign n1417 = \sa03_reg[3]/P0001  & n1416 ;
  assign n1418 = ~n1328 & ~n1417 ;
  assign n1419 = ~\sa03_reg[2]/P0001  & ~n1418 ;
  assign n1475 = ~n1415 & ~n1419 ;
  assign n1476 = ~n1428 & n1475 ;
  assign n1477 = ~n1413 & n1476 ;
  assign n1478 = ~n1393 & n1477 ;
  assign n1479 = ~n1474 & n1478 ;
  assign n1504 = n1408 & n1449 ;
  assign n1505 = ~\sa03_reg[2]/P0001  & n1504 ;
  assign n1506 = ~n1365 & ~n1505 ;
  assign n1507 = ~n1373 & n1506 ;
  assign n1508 = ~\sa03_reg[1]/P0001  & ~n1507 ;
  assign n1480 = n1339 & n1423 ;
  assign n1481 = ~n1459 & ~n1480 ;
  assign n1483 = ~\sa03_reg[4]/P0001  & n1328 ;
  assign n1482 = \sa03_reg[4]/P0001  & n1318 ;
  assign n1484 = ~n1331 & ~n1482 ;
  assign n1485 = ~n1483 & n1484 ;
  assign n1486 = \sa03_reg[2]/P0001  & ~n1485 ;
  assign n1487 = n1481 & ~n1486 ;
  assign n1488 = \sa03_reg[1]/P0001  & ~n1487 ;
  assign n1489 = ~n1399 & ~n1438 ;
  assign n1490 = n1355 & n1383 ;
  assign n1491 = n1489 & ~n1490 ;
  assign n1492 = \sa03_reg[2]/P0001  & ~n1491 ;
  assign n1498 = \sa03_reg[1]/P0001  & ~\sa03_reg[3]/P0001  ;
  assign n1499 = ~\sa03_reg[5]/P0001  & n1498 ;
  assign n1500 = ~n1368 & n1499 ;
  assign n1497 = n1342 & n1383 ;
  assign n1501 = ~n1335 & ~n1497 ;
  assign n1502 = ~n1500 & n1501 ;
  assign n1503 = ~\sa03_reg[2]/P0001  & ~n1502 ;
  assign n1493 = ~n1317 & ~n1380 ;
  assign n1494 = ~\sa03_reg[1]/P0001  & \sa03_reg[2]/P0001  ;
  assign n1495 = ~n1493 & n1494 ;
  assign n1496 = n1374 & n1404 ;
  assign n1509 = ~n1495 & ~n1496 ;
  assign n1510 = ~n1503 & n1509 ;
  assign n1511 = ~n1492 & n1510 ;
  assign n1512 = ~n1488 & n1511 ;
  assign n1513 = ~n1508 & n1512 ;
  assign n1514 = \sa03_reg[0]/P0001  & ~n1513 ;
  assign n1517 = ~n1378 & n1436 ;
  assign n1515 = ~\sa03_reg[2]/P0001  & ~\sa03_reg[4]/P0001  ;
  assign n1516 = n1460 & n1515 ;
  assign n1518 = \sa03_reg[1]/P0001  & ~n1400 ;
  assign n1519 = ~n1516 & n1518 ;
  assign n1520 = ~n1517 & n1519 ;
  assign n1521 = \sa03_reg[3]/P0001  & n1384 ;
  assign n1522 = n1449 & n1521 ;
  assign n1527 = ~\sa03_reg[1]/P0001  & ~n1497 ;
  assign n1528 = ~n1522 & n1527 ;
  assign n1526 = \sa03_reg[4]/P0001  & n1328 ;
  assign n1523 = ~\sa03_reg[2]/P0001  & n1317 ;
  assign n1524 = ~n1324 & ~n1408 ;
  assign n1525 = n1330 & ~n1524 ;
  assign n1529 = ~n1523 & ~n1525 ;
  assign n1530 = ~n1526 & n1529 ;
  assign n1531 = n1528 & n1530 ;
  assign n1532 = ~n1520 & ~n1531 ;
  assign n1533 = \sa03_reg[4]/P0001  & n1355 ;
  assign n1534 = ~n1323 & n1324 ;
  assign n1535 = ~n1533 & ~n1534 ;
  assign n1536 = ~n1316 & ~n1535 ;
  assign n1537 = n1367 & n1398 ;
  assign n1538 = ~\sa03_reg[2]/P0001  & ~n1537 ;
  assign n1539 = ~n1421 & n1538 ;
  assign n1540 = ~n1536 & n1539 ;
  assign n1541 = n1352 & n1355 ;
  assign n1542 = \sa03_reg[2]/P0001  & ~n1541 ;
  assign n1543 = ~n1526 & n1542 ;
  assign n1544 = ~n1540 & ~n1543 ;
  assign n1545 = ~n1532 & ~n1544 ;
  assign n1546 = ~\sa03_reg[0]/P0001  & ~n1545 ;
  assign n1561 = n1339 & n1368 ;
  assign n1562 = \sa03_reg[2]/P0001  & ~n1561 ;
  assign n1563 = ~\sa03_reg[7]/NET0131  & n1424 ;
  assign n1564 = n1562 & ~n1563 ;
  assign n1567 = ~\sa03_reg[2]/P0001  & ~n1365 ;
  assign n1565 = ~\sa03_reg[6]/NET0131  & n1340 ;
  assign n1566 = ~\sa03_reg[7]/NET0131  & n1396 ;
  assign n1568 = ~n1565 & ~n1566 ;
  assign n1569 = n1567 & n1568 ;
  assign n1570 = ~n1564 & ~n1569 ;
  assign n1571 = n1342 & n1352 ;
  assign n1572 = ~\sa03_reg[6]/NET0131  & n1317 ;
  assign n1573 = ~n1571 & ~n1572 ;
  assign n1574 = ~n1570 & n1573 ;
  assign n1575 = ~\sa03_reg[1]/P0001  & ~n1574 ;
  assign n1548 = ~\sa03_reg[6]/NET0131  & n1480 ;
  assign n1547 = n1341 & n1355 ;
  assign n1549 = ~n1409 & ~n1547 ;
  assign n1550 = ~n1548 & n1549 ;
  assign n1551 = \sa03_reg[1]/P0001  & ~n1550 ;
  assign n1552 = n1316 & n1380 ;
  assign n1553 = ~n1551 & ~n1552 ;
  assign n1554 = \sa03_reg[2]/P0001  & ~n1553 ;
  assign n1560 = n1365 & n1429 ;
  assign n1555 = ~\sa03_reg[2]/P0001  & \sa03_reg[4]/P0001  ;
  assign n1556 = n1376 & n1408 ;
  assign n1557 = ~n1555 & n1556 ;
  assign n1558 = \sa03_reg[1]/P0001  & ~\sa03_reg[2]/P0001  ;
  assign n1559 = n1417 & n1558 ;
  assign n1576 = ~n1557 & ~n1559 ;
  assign n1577 = ~n1560 & n1576 ;
  assign n1578 = ~n1554 & n1577 ;
  assign n1579 = ~n1575 & n1578 ;
  assign n1580 = ~n1546 & n1579 ;
  assign n1581 = ~n1514 & n1580 ;
  assign n1607 = ~\sa10_reg[4]/P0001  & \sa10_reg[6]/NET0131  ;
  assign n1608 = ~\sa10_reg[5]/P0001  & \sa10_reg[7]/NET0131  ;
  assign n1609 = n1607 & n1608 ;
  assign n1639 = ~\sa10_reg[3]/P0001  & n1609 ;
  assign n1593 = \sa10_reg[6]/NET0131  & ~\sa10_reg[7]/NET0131  ;
  assign n1636 = \sa10_reg[4]/P0001  & n1593 ;
  assign n1582 = \sa10_reg[5]/P0001  & ~\sa10_reg[6]/NET0131  ;
  assign n1637 = ~\sa10_reg[4]/P0001  & \sa10_reg[7]/NET0131  ;
  assign n1638 = n1582 & n1637 ;
  assign n1640 = ~n1636 & ~n1638 ;
  assign n1641 = ~n1639 & n1640 ;
  assign n1642 = \sa10_reg[2]/P0001  & ~n1641 ;
  assign n1626 = \sa10_reg[5]/P0001  & \sa10_reg[7]/NET0131  ;
  assign n1627 = \sa10_reg[3]/P0001  & ~\sa10_reg[4]/P0001  ;
  assign n1628 = n1626 & n1627 ;
  assign n1629 = \sa10_reg[5]/P0001  & ~\sa10_reg[7]/NET0131  ;
  assign n1594 = \sa10_reg[3]/P0001  & \sa10_reg[4]/P0001  ;
  assign n1630 = ~\sa10_reg[6]/NET0131  & n1594 ;
  assign n1631 = n1629 & n1630 ;
  assign n1632 = ~n1628 & ~n1631 ;
  assign n1633 = ~\sa10_reg[2]/P0001  & ~\sa10_reg[3]/P0001  ;
  assign n1634 = ~\sa10_reg[5]/P0001  & ~n1607 ;
  assign n1635 = n1633 & n1634 ;
  assign n1643 = n1632 & ~n1635 ;
  assign n1644 = ~n1642 & n1643 ;
  assign n1645 = \sa10_reg[1]/P0001  & ~n1644 ;
  assign n1614 = ~\sa10_reg[6]/NET0131  & ~\sa10_reg[7]/NET0131  ;
  assign n1615 = \sa10_reg[5]/P0001  & n1614 ;
  assign n1616 = ~\sa10_reg[3]/P0001  & n1615 ;
  assign n1617 = ~\sa10_reg[2]/P0001  & ~n1616 ;
  assign n1619 = \sa10_reg[7]/NET0131  & n1594 ;
  assign n1618 = ~\sa10_reg[5]/P0001  & n1593 ;
  assign n1620 = \sa10_reg[2]/P0001  & ~n1618 ;
  assign n1621 = ~n1619 & n1620 ;
  assign n1622 = ~n1617 & ~n1621 ;
  assign n1600 = ~\sa10_reg[5]/P0001  & ~\sa10_reg[7]/NET0131  ;
  assign n1606 = n1594 & n1600 ;
  assign n1610 = ~n1606 & ~n1609 ;
  assign n1611 = ~\sa10_reg[2]/P0001  & ~n1610 ;
  assign n1612 = \sa10_reg[4]/P0001  & \sa10_reg[7]/NET0131  ;
  assign n1613 = n1582 & n1612 ;
  assign n1623 = ~n1611 & ~n1613 ;
  assign n1624 = ~n1622 & n1623 ;
  assign n1625 = ~\sa10_reg[1]/P0001  & ~n1624 ;
  assign n1583 = ~\sa10_reg[3]/P0001  & \sa10_reg[4]/P0001  ;
  assign n1584 = n1582 & n1583 ;
  assign n1585 = \sa10_reg[5]/P0001  & \sa10_reg[6]/NET0131  ;
  assign n1586 = ~\sa10_reg[4]/P0001  & ~\sa10_reg[7]/NET0131  ;
  assign n1587 = n1585 & n1586 ;
  assign n1588 = ~n1584 & ~n1587 ;
  assign n1589 = ~\sa10_reg[2]/P0001  & ~n1588 ;
  assign n1590 = ~\sa10_reg[3]/P0001  & \sa10_reg[7]/NET0131  ;
  assign n1591 = n1585 & n1590 ;
  assign n1592 = \sa10_reg[4]/P0001  & n1591 ;
  assign n1595 = n1593 & n1594 ;
  assign n1596 = ~n1592 & ~n1595 ;
  assign n1597 = ~\sa10_reg[6]/NET0131  & \sa10_reg[7]/NET0131  ;
  assign n1598 = \sa10_reg[3]/P0001  & ~\sa10_reg[5]/P0001  ;
  assign n1599 = n1597 & n1598 ;
  assign n1601 = ~\sa10_reg[4]/P0001  & n1600 ;
  assign n1602 = ~\sa10_reg[6]/NET0131  & n1601 ;
  assign n1603 = ~n1599 & ~n1602 ;
  assign n1604 = n1596 & n1603 ;
  assign n1605 = \sa10_reg[2]/P0001  & ~n1604 ;
  assign n1646 = ~n1589 & ~n1605 ;
  assign n1647 = ~n1625 & n1646 ;
  assign n1648 = ~n1645 & n1647 ;
  assign n1649 = \sa10_reg[0]/P0001  & ~n1648 ;
  assign n1675 = ~\sa10_reg[1]/P0001  & ~n1587 ;
  assign n1666 = ~\sa10_reg[2]/P0001  & \sa10_reg[3]/P0001  ;
  assign n1667 = n1612 & n1666 ;
  assign n1671 = n1608 & n1627 ;
  assign n1676 = ~n1667 & ~n1671 ;
  assign n1677 = n1675 & n1676 ;
  assign n1672 = ~\sa10_reg[5]/P0001  & \sa10_reg[6]/NET0131  ;
  assign n1673 = \sa10_reg[4]/P0001  & n1672 ;
  assign n1674 = n1590 & n1673 ;
  assign n1664 = \sa10_reg[2]/P0001  & \sa10_reg[3]/P0001  ;
  assign n1665 = n1615 & n1664 ;
  assign n1668 = ~\sa10_reg[3]/P0001  & ~\sa10_reg[4]/P0001  ;
  assign n1669 = \sa10_reg[7]/NET0131  & n1668 ;
  assign n1670 = ~\sa10_reg[6]/NET0131  & n1669 ;
  assign n1678 = ~n1665 & ~n1670 ;
  assign n1679 = ~n1674 & n1678 ;
  assign n1680 = n1677 & n1679 ;
  assign n1687 = ~\sa10_reg[5]/P0001  & n1614 ;
  assign n1688 = ~\sa10_reg[2]/P0001  & n1687 ;
  assign n1689 = ~\sa10_reg[4]/P0001  & n1688 ;
  assign n1661 = \sa10_reg[2]/P0001  & ~\sa10_reg[3]/P0001  ;
  assign n1684 = \sa10_reg[4]/P0001  & n1626 ;
  assign n1685 = ~n1601 & ~n1684 ;
  assign n1686 = n1661 & ~n1685 ;
  assign n1681 = \sa10_reg[3]/P0001  & \sa10_reg[6]/NET0131  ;
  assign n1682 = n1629 & n1681 ;
  assign n1683 = \sa10_reg[4]/P0001  & n1682 ;
  assign n1690 = \sa10_reg[1]/P0001  & ~n1683 ;
  assign n1691 = ~n1686 & n1690 ;
  assign n1692 = ~n1689 & n1691 ;
  assign n1693 = ~n1680 & ~n1692 ;
  assign n1656 = ~\sa10_reg[7]/NET0131  & n1583 ;
  assign n1657 = n1585 & n1656 ;
  assign n1650 = ~\sa10_reg[5]/P0001  & ~\sa10_reg[6]/NET0131  ;
  assign n1651 = n1583 & n1650 ;
  assign n1652 = \sa10_reg[6]/NET0131  & \sa10_reg[7]/NET0131  ;
  assign n1653 = \sa10_reg[4]/P0001  & ~n1652 ;
  assign n1654 = n1598 & ~n1614 ;
  assign n1655 = ~n1653 & n1654 ;
  assign n1658 = ~n1651 & ~n1655 ;
  assign n1659 = ~n1657 & n1658 ;
  assign n1660 = ~\sa10_reg[2]/P0001  & ~n1659 ;
  assign n1662 = n1634 & n1661 ;
  assign n1663 = ~n1653 & n1662 ;
  assign n1694 = ~n1660 & ~n1663 ;
  assign n1695 = ~n1693 & n1694 ;
  assign n1696 = ~\sa10_reg[0]/P0001  & ~n1695 ;
  assign n1699 = ~\sa10_reg[6]/NET0131  & n1626 ;
  assign n1707 = ~n1668 & n1699 ;
  assign n1708 = ~\sa10_reg[5]/P0001  & n1636 ;
  assign n1709 = ~n1707 & ~n1708 ;
  assign n1710 = ~\sa10_reg[2]/P0001  & ~n1709 ;
  assign n1711 = n1585 & n1668 ;
  assign n1712 = ~\sa10_reg[6]/NET0131  & n1619 ;
  assign n1717 = ~n1711 & ~n1712 ;
  assign n1713 = n1607 & n1626 ;
  assign n1714 = \sa10_reg[2]/P0001  & n1713 ;
  assign n1715 = \sa10_reg[2]/P0001  & n1627 ;
  assign n1716 = n1614 & n1715 ;
  assign n1718 = ~n1714 & ~n1716 ;
  assign n1719 = n1717 & n1718 ;
  assign n1720 = ~n1710 & n1719 ;
  assign n1721 = ~\sa10_reg[1]/P0001  & ~n1720 ;
  assign n1697 = \sa10_reg[1]/P0001  & \sa10_reg[2]/P0001  ;
  assign n1698 = ~\sa10_reg[3]/P0001  & n1614 ;
  assign n1700 = \sa10_reg[3]/P0001  & n1699 ;
  assign n1701 = ~n1698 & ~n1700 ;
  assign n1702 = ~\sa10_reg[4]/P0001  & ~n1701 ;
  assign n1703 = \sa10_reg[4]/P0001  & n1614 ;
  assign n1704 = ~\sa10_reg[5]/P0001  & n1703 ;
  assign n1705 = ~n1702 & ~n1704 ;
  assign n1706 = n1697 & ~n1705 ;
  assign n1726 = \sa10_reg[5]/P0001  & n1627 ;
  assign n1727 = n1614 & n1726 ;
  assign n1728 = ~\sa10_reg[2]/P0001  & n1727 ;
  assign n1729 = \sa10_reg[1]/P0001  & n1728 ;
  assign n1722 = \sa10_reg[2]/P0001  & ~\sa10_reg[5]/P0001  ;
  assign n1723 = ~n1595 & ~n1698 ;
  assign n1724 = n1722 & ~n1723 ;
  assign n1725 = n1613 & n1666 ;
  assign n1730 = n1614 & n1668 ;
  assign n1731 = ~\sa10_reg[5]/P0001  & n1730 ;
  assign n1732 = ~n1725 & ~n1731 ;
  assign n1733 = ~n1724 & n1732 ;
  assign n1734 = ~n1729 & n1733 ;
  assign n1735 = ~n1706 & n1734 ;
  assign n1736 = ~n1721 & n1735 ;
  assign n1737 = ~n1696 & n1736 ;
  assign n1738 = ~n1649 & n1737 ;
  assign n1739 = ~n1581 & ~n1738 ;
  assign n1740 = n1581 & n1738 ;
  assign n1741 = ~n1739 & ~n1740 ;
  assign n1742 = ~n1479 & ~n1741 ;
  assign n1743 = n1479 & n1741 ;
  assign n1744 = ~n1742 & ~n1743 ;
  assign n1772 = \sa21_reg[5]/P0001  & ~\sa21_reg[6]/NET0131  ;
  assign n1799 = ~\sa21_reg[3]/P0001  & ~\sa21_reg[7]/P0001  ;
  assign n1800 = n1772 & n1799 ;
  assign n1801 = ~\sa21_reg[2]/P0001  & ~n1800 ;
  assign n1761 = \sa21_reg[6]/NET0131  & ~\sa21_reg[7]/P0001  ;
  assign n1804 = ~\sa21_reg[5]/P0001  & n1761 ;
  assign n1802 = \sa21_reg[3]/P0001  & \sa21_reg[4]/P0001  ;
  assign n1803 = \sa21_reg[7]/P0001  & n1802 ;
  assign n1805 = \sa21_reg[2]/P0001  & ~n1803 ;
  assign n1806 = ~n1804 & n1805 ;
  assign n1807 = ~n1801 & ~n1806 ;
  assign n1763 = ~\sa21_reg[6]/NET0131  & \sa21_reg[7]/P0001  ;
  assign n1764 = \sa21_reg[5]/P0001  & n1763 ;
  assign n1792 = \sa21_reg[4]/P0001  & n1764 ;
  assign n1758 = ~\sa21_reg[5]/P0001  & \sa21_reg[6]/NET0131  ;
  assign n1793 = ~\sa21_reg[4]/P0001  & \sa21_reg[7]/P0001  ;
  assign n1794 = n1758 & n1793 ;
  assign n1784 = ~\sa21_reg[5]/P0001  & ~\sa21_reg[7]/P0001  ;
  assign n1795 = \sa21_reg[4]/P0001  & n1784 ;
  assign n1796 = \sa21_reg[3]/P0001  & n1795 ;
  assign n1797 = ~n1794 & ~n1796 ;
  assign n1798 = ~\sa21_reg[2]/P0001  & ~n1797 ;
  assign n1808 = ~n1792 & ~n1798 ;
  assign n1809 = ~n1807 & n1808 ;
  assign n1810 = ~\sa21_reg[1]/P0001  & ~n1809 ;
  assign n1765 = ~\sa21_reg[4]/P0001  & n1764 ;
  assign n1757 = ~\sa21_reg[3]/P0001  & \sa21_reg[7]/P0001  ;
  assign n1759 = ~\sa21_reg[4]/P0001  & n1758 ;
  assign n1760 = n1757 & n1759 ;
  assign n1762 = \sa21_reg[4]/P0001  & n1761 ;
  assign n1766 = ~n1760 & ~n1762 ;
  assign n1767 = ~n1765 & n1766 ;
  assign n1768 = \sa21_reg[2]/P0001  & ~n1767 ;
  assign n1745 = \sa21_reg[5]/P0001  & ~\sa21_reg[7]/P0001  ;
  assign n1746 = \sa21_reg[3]/P0001  & ~\sa21_reg[6]/NET0131  ;
  assign n1747 = \sa21_reg[4]/P0001  & n1746 ;
  assign n1748 = n1745 & n1747 ;
  assign n1749 = \sa21_reg[5]/P0001  & \sa21_reg[7]/P0001  ;
  assign n1750 = \sa21_reg[3]/P0001  & n1749 ;
  assign n1751 = ~\sa21_reg[4]/P0001  & n1750 ;
  assign n1752 = ~n1748 & ~n1751 ;
  assign n1753 = ~\sa21_reg[4]/P0001  & \sa21_reg[6]/NET0131  ;
  assign n1754 = ~\sa21_reg[2]/P0001  & ~\sa21_reg[3]/P0001  ;
  assign n1755 = ~\sa21_reg[5]/P0001  & n1754 ;
  assign n1756 = ~n1753 & n1755 ;
  assign n1769 = n1752 & ~n1756 ;
  assign n1770 = ~n1768 & n1769 ;
  assign n1771 = \sa21_reg[1]/P0001  & ~n1770 ;
  assign n1773 = ~\sa21_reg[3]/P0001  & \sa21_reg[4]/P0001  ;
  assign n1774 = n1772 & n1773 ;
  assign n1775 = ~\sa21_reg[4]/P0001  & n1761 ;
  assign n1776 = \sa21_reg[5]/P0001  & n1775 ;
  assign n1777 = ~n1774 & ~n1776 ;
  assign n1778 = ~\sa21_reg[2]/P0001  & ~n1777 ;
  assign n1779 = \sa21_reg[3]/P0001  & n1761 ;
  assign n1780 = \sa21_reg[4]/P0001  & n1779 ;
  assign n1781 = \sa21_reg[6]/NET0131  & n1749 ;
  assign n1782 = n1773 & n1781 ;
  assign n1783 = ~n1780 & ~n1782 ;
  assign n1785 = ~\sa21_reg[4]/P0001  & n1784 ;
  assign n1786 = ~\sa21_reg[6]/NET0131  & n1785 ;
  assign n1787 = \sa21_reg[3]/P0001  & ~\sa21_reg[5]/P0001  ;
  assign n1788 = n1763 & n1787 ;
  assign n1789 = ~n1786 & ~n1788 ;
  assign n1790 = n1783 & n1789 ;
  assign n1791 = \sa21_reg[2]/P0001  & ~n1790 ;
  assign n1811 = ~n1778 & ~n1791 ;
  assign n1812 = ~n1771 & n1811 ;
  assign n1813 = ~n1810 & n1812 ;
  assign n1814 = \sa21_reg[0]/P0001  & ~n1813 ;
  assign n1852 = ~\sa21_reg[2]/P0001  & n1786 ;
  assign n1831 = \sa21_reg[2]/P0001  & ~\sa21_reg[3]/P0001  ;
  assign n1849 = \sa21_reg[4]/P0001  & n1749 ;
  assign n1850 = ~n1785 & ~n1849 ;
  assign n1851 = n1831 & ~n1850 ;
  assign n1837 = \sa21_reg[5]/P0001  & \sa21_reg[6]/NET0131  ;
  assign n1853 = \sa21_reg[4]/P0001  & n1837 ;
  assign n1854 = \sa21_reg[3]/P0001  & ~\sa21_reg[7]/P0001  ;
  assign n1855 = n1853 & n1854 ;
  assign n1856 = ~n1851 & ~n1855 ;
  assign n1857 = ~n1852 & n1856 ;
  assign n1858 = \sa21_reg[1]/P0001  & ~n1857 ;
  assign n1818 = n1787 & n1793 ;
  assign n1825 = ~n1776 & ~n1818 ;
  assign n1815 = ~\sa21_reg[3]/P0001  & ~\sa21_reg[4]/P0001  ;
  assign n1816 = \sa21_reg[7]/P0001  & n1815 ;
  assign n1817 = ~\sa21_reg[6]/NET0131  & n1816 ;
  assign n1819 = \sa21_reg[2]/P0001  & n1745 ;
  assign n1820 = n1746 & n1819 ;
  assign n1826 = ~n1817 & ~n1820 ;
  assign n1821 = ~\sa21_reg[2]/P0001  & n1803 ;
  assign n1822 = \sa21_reg[6]/NET0131  & \sa21_reg[7]/P0001  ;
  assign n1823 = ~\sa21_reg[5]/P0001  & n1822 ;
  assign n1824 = n1773 & n1823 ;
  assign n1827 = ~n1821 & ~n1824 ;
  assign n1828 = n1826 & n1827 ;
  assign n1829 = n1825 & n1828 ;
  assign n1830 = ~\sa21_reg[1]/P0001  & ~n1829 ;
  assign n1832 = ~\sa21_reg[5]/P0001  & ~\sa21_reg[6]/NET0131  ;
  assign n1833 = ~\sa21_reg[4]/P0001  & n1832 ;
  assign n1834 = \sa21_reg[4]/P0001  & n1823 ;
  assign n1835 = ~n1833 & ~n1834 ;
  assign n1836 = n1831 & ~n1835 ;
  assign n1844 = \sa21_reg[4]/P0001  & n1832 ;
  assign n1845 = ~\sa21_reg[3]/P0001  & n1844 ;
  assign n1838 = n1799 & n1837 ;
  assign n1839 = \sa21_reg[4]/P0001  & n1838 ;
  assign n1840 = \sa21_reg[4]/P0001  & ~n1822 ;
  assign n1841 = ~\sa21_reg[6]/NET0131  & ~\sa21_reg[7]/P0001  ;
  assign n1842 = n1787 & ~n1841 ;
  assign n1843 = ~n1840 & n1842 ;
  assign n1846 = ~n1839 & ~n1843 ;
  assign n1847 = ~n1845 & n1846 ;
  assign n1848 = ~\sa21_reg[2]/P0001  & ~n1847 ;
  assign n1859 = ~n1836 & ~n1848 ;
  assign n1860 = ~n1830 & n1859 ;
  assign n1861 = ~n1858 & n1860 ;
  assign n1862 = ~\sa21_reg[0]/P0001  & ~n1861 ;
  assign n1885 = ~\sa21_reg[6]/NET0131  & n1750 ;
  assign n1884 = ~\sa21_reg[5]/P0001  & n1762 ;
  assign n1886 = ~n1792 & ~n1884 ;
  assign n1887 = ~n1885 & n1886 ;
  assign n1888 = ~\sa21_reg[2]/P0001  & ~n1887 ;
  assign n1889 = ~\sa21_reg[6]/NET0131  & n1803 ;
  assign n1890 = ~\sa21_reg[3]/P0001  & n1753 ;
  assign n1891 = \sa21_reg[5]/P0001  & n1890 ;
  assign n1897 = ~n1889 & ~n1891 ;
  assign n1892 = n1793 & n1837 ;
  assign n1893 = \sa21_reg[2]/P0001  & n1892 ;
  assign n1894 = \sa21_reg[2]/P0001  & \sa21_reg[3]/P0001  ;
  assign n1895 = ~\sa21_reg[4]/P0001  & n1894 ;
  assign n1896 = n1841 & n1895 ;
  assign n1898 = ~n1893 & ~n1896 ;
  assign n1899 = n1897 & n1898 ;
  assign n1900 = ~n1888 & n1899 ;
  assign n1901 = ~\sa21_reg[1]/P0001  & ~n1900 ;
  assign n1863 = \sa21_reg[1]/P0001  & \sa21_reg[2]/P0001  ;
  assign n1866 = \sa21_reg[3]/P0001  & ~\sa21_reg[4]/P0001  ;
  assign n1867 = \sa21_reg[5]/P0001  & n1866 ;
  assign n1868 = n1763 & n1867 ;
  assign n1864 = ~\sa21_reg[6]/NET0131  & n1795 ;
  assign n1865 = n1815 & n1841 ;
  assign n1869 = ~n1864 & ~n1865 ;
  assign n1870 = ~n1868 & n1869 ;
  assign n1871 = n1863 & ~n1870 ;
  assign n1877 = ~\sa21_reg[2]/P0001  & \sa21_reg[3]/P0001  ;
  assign n1879 = ~\sa21_reg[4]/P0001  & n1745 ;
  assign n1880 = ~\sa21_reg[6]/NET0131  & n1879 ;
  assign n1881 = n1877 & n1880 ;
  assign n1882 = \sa21_reg[1]/P0001  & n1881 ;
  assign n1872 = n1799 & n1832 ;
  assign n1873 = n1758 & n1802 ;
  assign n1874 = ~\sa21_reg[7]/P0001  & n1873 ;
  assign n1875 = ~n1872 & ~n1874 ;
  assign n1876 = \sa21_reg[2]/P0001  & ~n1875 ;
  assign n1878 = n1792 & n1877 ;
  assign n1883 = n1799 & n1833 ;
  assign n1902 = ~n1878 & ~n1883 ;
  assign n1903 = ~n1876 & n1902 ;
  assign n1904 = ~n1882 & n1903 ;
  assign n1905 = ~n1871 & n1904 ;
  assign n1906 = ~n1901 & n1905 ;
  assign n1907 = ~n1862 & n1906 ;
  assign n1908 = ~n1814 & n1907 ;
  assign n1981 = \sa32_reg[6]/NET0131  & ~\sa32_reg[7]/P0001  ;
  assign n1982 = ~\sa32_reg[3]/P0001  & n1981 ;
  assign n1983 = ~\sa32_reg[4]/P0001  & n1982 ;
  assign n1923 = ~\sa32_reg[6]/NET0131  & \sa32_reg[7]/P0001  ;
  assign n1932 = \sa32_reg[3]/P0001  & n1923 ;
  assign n1919 = ~\sa32_reg[3]/P0001  & \sa32_reg[4]/P0001  ;
  assign n1939 = \sa32_reg[5]/P0001  & ~\sa32_reg[6]/NET0131  ;
  assign n1940 = n1919 & n1939 ;
  assign n1984 = ~n1932 & ~n1940 ;
  assign n1985 = ~n1983 & n1984 ;
  assign n1986 = ~\sa32_reg[2]/P0001  & ~n1985 ;
  assign n1920 = \sa32_reg[5]/P0001  & \sa32_reg[7]/P0001  ;
  assign n1977 = \sa32_reg[3]/P0001  & n1920 ;
  assign n1909 = \sa32_reg[5]/P0001  & \sa32_reg[6]/NET0131  ;
  assign n1910 = ~\sa32_reg[7]/P0001  & n1909 ;
  assign n1978 = \sa32_reg[4]/P0001  & n1910 ;
  assign n1979 = ~n1977 & ~n1978 ;
  assign n1980 = \sa32_reg[2]/P0001  & ~n1979 ;
  assign n1987 = \sa32_reg[6]/NET0131  & \sa32_reg[7]/P0001  ;
  assign n1988 = ~\sa32_reg[5]/P0001  & n1987 ;
  assign n1989 = ~\sa32_reg[3]/P0001  & n1988 ;
  assign n1912 = \sa32_reg[3]/P0001  & \sa32_reg[4]/P0001  ;
  assign n1993 = n1912 & n1920 ;
  assign n1970 = ~\sa32_reg[4]/P0001  & \sa32_reg[5]/P0001  ;
  assign n1994 = n1923 & n1970 ;
  assign n1997 = ~n1993 & ~n1994 ;
  assign n1998 = ~n1989 & n1997 ;
  assign n1990 = ~\sa32_reg[5]/P0001  & ~\sa32_reg[6]/NET0131  ;
  assign n1991 = \sa32_reg[3]/P0001  & n1990 ;
  assign n1992 = ~\sa32_reg[7]/P0001  & n1991 ;
  assign n1995 = ~\sa32_reg[3]/P0001  & ~\sa32_reg[4]/P0001  ;
  assign n1996 = n1910 & n1995 ;
  assign n1999 = ~n1992 & ~n1996 ;
  assign n2000 = n1998 & n1999 ;
  assign n2001 = ~n1980 & n2000 ;
  assign n2002 = ~n1986 & n2001 ;
  assign n2003 = \sa32_reg[1]/P0001  & ~n2002 ;
  assign n1951 = \sa32_reg[3]/P0001  & ~\sa32_reg[4]/P0001  ;
  assign n2004 = ~\sa32_reg[6]/NET0131  & n1951 ;
  assign n2005 = \sa32_reg[2]/P0001  & n2004 ;
  assign n2006 = n1919 & n1923 ;
  assign n2007 = ~n2005 & ~n2006 ;
  assign n2008 = ~\sa32_reg[5]/P0001  & ~n2007 ;
  assign n1913 = ~\sa32_reg[6]/NET0131  & ~\sa32_reg[7]/P0001  ;
  assign n1937 = ~\sa32_reg[5]/P0001  & n1913 ;
  assign n2009 = ~\sa32_reg[3]/P0001  & n1937 ;
  assign n2010 = \sa32_reg[2]/P0001  & n2009 ;
  assign n2011 = \sa32_reg[7]/P0001  & n1909 ;
  assign n2012 = ~\sa32_reg[3]/P0001  & n2011 ;
  assign n2013 = ~\sa32_reg[4]/P0001  & n2012 ;
  assign n2014 = ~n2010 & ~n2013 ;
  assign n2015 = ~n2008 & n2014 ;
  assign n2016 = ~\sa32_reg[1]/P0001  & ~n2015 ;
  assign n2019 = ~\sa32_reg[5]/P0001  & n1981 ;
  assign n2020 = n1919 & n2019 ;
  assign n1948 = ~\sa32_reg[4]/P0001  & ~\sa32_reg[7]/P0001  ;
  assign n1924 = \sa32_reg[3]/P0001  & ~\sa32_reg[5]/P0001  ;
  assign n2017 = \sa32_reg[6]/NET0131  & ~n1924 ;
  assign n2018 = n1948 & ~n2017 ;
  assign n2021 = ~n1993 & ~n2018 ;
  assign n2022 = ~n2020 & n2021 ;
  assign n2023 = \sa32_reg[2]/P0001  & ~n2022 ;
  assign n2026 = ~\sa32_reg[2]/P0001  & \sa32_reg[3]/P0001  ;
  assign n2027 = ~\sa32_reg[5]/P0001  & ~\sa32_reg[7]/P0001  ;
  assign n2028 = \sa32_reg[4]/P0001  & n2027 ;
  assign n2029 = n2026 & n2028 ;
  assign n2030 = ~\sa32_reg[2]/P0001  & ~\sa32_reg[4]/P0001  ;
  assign n2031 = n1988 & n2030 ;
  assign n2032 = ~n2029 & ~n2031 ;
  assign n1953 = \sa32_reg[4]/P0001  & \sa32_reg[7]/P0001  ;
  assign n2024 = n1939 & n1953 ;
  assign n2025 = ~\sa32_reg[2]/P0001  & n2024 ;
  assign n2033 = n1948 & n1990 ;
  assign n2034 = ~n2025 & ~n2033 ;
  assign n2035 = n2032 & n2034 ;
  assign n2036 = ~n2023 & n2035 ;
  assign n2037 = ~n2016 & n2036 ;
  assign n2038 = ~n2003 & n2037 ;
  assign n2039 = ~\sa32_reg[0]/P0002  & ~n2038 ;
  assign n1952 = \sa32_reg[5]/P0001  & n1951 ;
  assign n1954 = ~\sa32_reg[4]/P0001  & \sa32_reg[6]/NET0131  ;
  assign n1955 = ~\sa32_reg[5]/P0001  & ~n1954 ;
  assign n1956 = ~n1953 & n1955 ;
  assign n1957 = ~n1952 & ~n1956 ;
  assign n1958 = \sa32_reg[1]/P0001  & ~n1957 ;
  assign n1911 = \sa32_reg[3]/P0001  & n1910 ;
  assign n1947 = \sa32_reg[3]/P0001  & \sa32_reg[6]/NET0131  ;
  assign n1949 = n1947 & n1948 ;
  assign n1950 = ~n1911 & ~n1949 ;
  assign n1934 = \sa32_reg[5]/P0001  & ~\sa32_reg[7]/P0001  ;
  assign n1959 = ~\sa32_reg[4]/P0001  & n1934 ;
  assign n1960 = n1950 & ~n1959 ;
  assign n1961 = ~n1958 & n1960 ;
  assign n1962 = ~\sa32_reg[2]/P0001  & ~n1961 ;
  assign n1921 = n1919 & n1920 ;
  assign n1922 = \sa32_reg[6]/NET0131  & n1921 ;
  assign n1928 = ~\sa32_reg[1]/P0001  & ~n1911 ;
  assign n1929 = ~n1922 & n1928 ;
  assign n1914 = n1912 & n1913 ;
  assign n1915 = ~\sa32_reg[5]/P0001  & \sa32_reg[6]/NET0131  ;
  assign n1916 = ~\sa32_reg[4]/P0001  & n1915 ;
  assign n1917 = ~n1914 & ~n1916 ;
  assign n1918 = \sa32_reg[2]/P0001  & ~n1917 ;
  assign n1925 = n1923 & n1924 ;
  assign n1926 = ~n1910 & ~n1925 ;
  assign n1927 = ~\sa32_reg[2]/P0001  & ~n1926 ;
  assign n1930 = ~n1918 & ~n1927 ;
  assign n1931 = n1929 & n1930 ;
  assign n1933 = ~\sa32_reg[4]/P0001  & n1932 ;
  assign n1942 = \sa32_reg[1]/P0001  & ~n1933 ;
  assign n1941 = \sa32_reg[7]/P0001  & n1940 ;
  assign n1935 = n1912 & n1934 ;
  assign n1936 = ~\sa32_reg[6]/NET0131  & n1935 ;
  assign n1938 = n1919 & n1937 ;
  assign n1943 = ~n1936 & ~n1938 ;
  assign n1944 = ~n1941 & n1943 ;
  assign n1945 = n1942 & n1944 ;
  assign n1946 = ~n1931 & ~n1945 ;
  assign n1965 = ~\sa32_reg[3]/P0001  & n1915 ;
  assign n1966 = n1948 & n1965 ;
  assign n1967 = ~n1922 & ~n1966 ;
  assign n1968 = \sa32_reg[2]/P0001  & ~n1967 ;
  assign n1963 = n1915 & n1953 ;
  assign n1964 = ~\sa32_reg[2]/P0001  & n1963 ;
  assign n1969 = ~\sa32_reg[7]/P0001  & n1947 ;
  assign n1971 = n1969 & n1970 ;
  assign n1972 = ~n1964 & ~n1971 ;
  assign n1973 = ~n1968 & n1972 ;
  assign n1974 = ~n1946 & n1973 ;
  assign n1975 = ~n1962 & n1974 ;
  assign n1976 = \sa32_reg[0]/P0002  & ~n1975 ;
  assign n2052 = \sa32_reg[6]/NET0131  & n1935 ;
  assign n2049 = ~\sa32_reg[4]/P0001  & \sa32_reg[7]/P0001  ;
  assign n2050 = ~\sa32_reg[3]/P0001  & n2049 ;
  assign n2051 = \sa32_reg[5]/P0001  & n2050 ;
  assign n2053 = ~n1963 & ~n2051 ;
  assign n2054 = ~n2052 & n2053 ;
  assign n2055 = ~\sa32_reg[2]/P0001  & ~n2054 ;
  assign n2040 = n1913 & n1995 ;
  assign n2041 = ~\sa32_reg[5]/P0001  & n1923 ;
  assign n2042 = ~n2019 & ~n2041 ;
  assign n2043 = ~\sa32_reg[3]/P0001  & ~n2011 ;
  assign n2044 = n2042 & n2043 ;
  assign n2045 = \sa32_reg[3]/P0001  & ~n1939 ;
  assign n2046 = \sa32_reg[2]/P0001  & \sa32_reg[4]/P0001  ;
  assign n2047 = ~n2045 & n2046 ;
  assign n2048 = ~n2044 & n2047 ;
  assign n2056 = ~n2040 & ~n2048 ;
  assign n2057 = ~n2055 & n2056 ;
  assign n2058 = ~\sa32_reg[1]/P0001  & ~n2057 ;
  assign n2067 = \sa32_reg[2]/P0001  & n1981 ;
  assign n2068 = \sa32_reg[5]/P0001  & n2067 ;
  assign n2069 = n1919 & n2068 ;
  assign n2066 = n1937 & n1951 ;
  assign n2070 = ~n2025 & ~n2066 ;
  assign n2071 = ~n2069 & n2070 ;
  assign n2072 = \sa32_reg[1]/P0001  & ~n2071 ;
  assign n2059 = \sa32_reg[2]/P0001  & \sa32_reg[3]/P0001  ;
  assign n2060 = \sa32_reg[5]/P0001  & n1913 ;
  assign n2061 = n2059 & n2060 ;
  assign n2062 = \sa32_reg[4]/P0001  & n2061 ;
  assign n2063 = n1934 & n2004 ;
  assign n2064 = ~n1989 & ~n2063 ;
  assign n2065 = ~\sa32_reg[2]/P0001  & ~n2064 ;
  assign n2073 = ~n2062 & ~n2065 ;
  assign n2074 = ~n2072 & n2073 ;
  assign n2075 = ~n2058 & n2074 ;
  assign n2076 = ~n1976 & n2075 ;
  assign n2077 = ~n2039 & n2076 ;
  assign n2078 = \u0_w_reg[3][6]/P0001  & ~n2077 ;
  assign n2079 = ~\u0_w_reg[3][6]/P0001  & n2077 ;
  assign n2080 = ~n2078 & ~n2079 ;
  assign n2081 = n1908 & n2080 ;
  assign n2082 = ~n1908 & ~n2080 ;
  assign n2083 = ~n2081 & ~n2082 ;
  assign n2085 = n1744 & ~n2083 ;
  assign n2084 = ~n1744 & n2083 ;
  assign n2086 = ~\ld_r_reg/P0001  & ~n2084 ;
  assign n2087 = ~n2085 & n2086 ;
  assign n2089 = ~\text_in_r_reg[6]/P0001  & \u0_w_reg[3][6]/P0001  ;
  assign n2088 = \text_in_r_reg[6]/P0001  & ~\u0_w_reg[3][6]/P0001  ;
  assign n2090 = \ld_r_reg/P0001  & ~n2088 ;
  assign n2091 = ~n2089 & n2090 ;
  assign n2092 = ~n2087 & ~n2091 ;
  assign n2128 = n1583 & n1672 ;
  assign n2129 = \sa10_reg[2]/P0001  & ~n2128 ;
  assign n2130 = n1593 & n1598 ;
  assign n2131 = ~\sa10_reg[2]/P0001  & ~n2130 ;
  assign n2132 = ~n1630 & n2131 ;
  assign n2133 = ~n2129 & ~n2132 ;
  assign n2134 = ~n1674 & ~n1700 ;
  assign n2135 = ~n2133 & n2134 ;
  assign n2136 = \sa10_reg[1]/P0001  & ~n2135 ;
  assign n2123 = n1629 & n1668 ;
  assign n2124 = ~n1591 & ~n2123 ;
  assign n2125 = ~n1683 & ~n1704 ;
  assign n2126 = n2124 & n2125 ;
  assign n2127 = ~\sa10_reg[2]/P0001  & ~n2126 ;
  assign n2110 = \sa10_reg[2]/P0001  & n1594 ;
  assign n2111 = n1608 & n2110 ;
  assign n2112 = \sa10_reg[2]/P0001  & ~\sa10_reg[6]/NET0131  ;
  assign n2113 = n1600 & n2112 ;
  assign n2109 = ~\sa10_reg[2]/P0001  & n1637 ;
  assign n2114 = ~n1628 & ~n2109 ;
  assign n2115 = ~n2113 & n2114 ;
  assign n2116 = ~n2111 & n2115 ;
  assign n2117 = ~\sa10_reg[1]/P0001  & ~n2116 ;
  assign n2119 = \sa10_reg[5]/P0001  & n1703 ;
  assign n2118 = n1585 & n1612 ;
  assign n2120 = ~n1602 & ~n2118 ;
  assign n2121 = ~n2119 & n2120 ;
  assign n2122 = n1664 & ~n2121 ;
  assign n2137 = ~n2117 & ~n2122 ;
  assign n2138 = ~n2127 & n2137 ;
  assign n2139 = ~n2136 & n2138 ;
  assign n2140 = ~\sa10_reg[0]/P0001  & ~n2139 ;
  assign n2093 = n1600 & n1607 ;
  assign n2094 = ~n1713 & ~n2093 ;
  assign n2095 = n1582 & ~n1637 ;
  assign n2096 = n2094 & ~n2095 ;
  assign n2097 = n1666 & ~n2096 ;
  assign n2098 = \sa10_reg[4]/P0001  & n1650 ;
  assign n2099 = ~n1607 & ~n2098 ;
  assign n2100 = \sa10_reg[7]/NET0131  & ~n2099 ;
  assign n2101 = n1582 & n1586 ;
  assign n2102 = ~n2100 & ~n2101 ;
  assign n2103 = ~\sa10_reg[3]/P0001  & ~n2102 ;
  assign n2104 = ~n1609 & ~n1682 ;
  assign n2105 = ~n2103 & n2104 ;
  assign n2106 = \sa10_reg[2]/P0001  & ~n2105 ;
  assign n2107 = ~n2097 & ~n2106 ;
  assign n2108 = \sa10_reg[1]/P0001  & ~n2107 ;
  assign n2142 = ~\sa10_reg[2]/P0001  & ~n1582 ;
  assign n2143 = \sa10_reg[5]/P0001  & ~n1637 ;
  assign n2144 = ~n1653 & ~n2143 ;
  assign n2145 = n2142 & ~n2144 ;
  assign n2148 = \sa10_reg[6]/NET0131  & n1656 ;
  assign n2141 = n1669 & n1722 ;
  assign n2146 = n1582 & n1627 ;
  assign n2147 = n1593 & n1633 ;
  assign n2149 = ~n2146 & ~n2147 ;
  assign n2150 = ~n2141 & n2149 ;
  assign n2151 = ~n2148 & n2150 ;
  assign n2152 = ~n2145 & n2151 ;
  assign n2153 = ~\sa10_reg[1]/P0001  & ~n2152 ;
  assign n2154 = n1608 & n1633 ;
  assign n2155 = ~\sa10_reg[6]/NET0131  & n2154 ;
  assign n2156 = n1619 & n1672 ;
  assign n2157 = ~n2155 & ~n2156 ;
  assign n2158 = \sa10_reg[1]/P0001  & ~n2157 ;
  assign n2161 = \sa10_reg[4]/P0001  & n2147 ;
  assign n2159 = n1672 & n1715 ;
  assign n2160 = \sa10_reg[5]/P0001  & n1656 ;
  assign n2172 = ~n2159 & ~n2160 ;
  assign n2173 = ~n2161 & n2172 ;
  assign n2174 = ~n2158 & n2173 ;
  assign n2162 = \sa10_reg[3]/P0001  & ~\sa10_reg[7]/NET0131  ;
  assign n2163 = \sa10_reg[6]/NET0131  & n2162 ;
  assign n2164 = ~n1698 & ~n2163 ;
  assign n2165 = n2099 & n2164 ;
  assign n2166 = n1697 & ~n2165 ;
  assign n2168 = \sa10_reg[5]/P0001  & n1636 ;
  assign n2167 = n1590 & n1607 ;
  assign n2169 = ~n1584 & ~n2167 ;
  assign n2170 = ~n2168 & n2169 ;
  assign n2171 = \sa10_reg[2]/P0001  & ~n2170 ;
  assign n2175 = ~n2166 & ~n2171 ;
  assign n2176 = n2174 & n2175 ;
  assign n2177 = ~n2153 & n2176 ;
  assign n2178 = \sa10_reg[0]/P0001  & ~n2177 ;
  assign n2189 = n1583 & n1626 ;
  assign n2191 = ~n1671 & ~n2189 ;
  assign n2192 = n2124 & n2191 ;
  assign n2190 = \sa10_reg[2]/P0001  & ~n2189 ;
  assign n2193 = ~\sa10_reg[1]/P0001  & ~n2190 ;
  assign n2194 = ~n2192 & n2193 ;
  assign n2179 = ~\sa10_reg[7]/NET0131  & n1711 ;
  assign n2180 = ~\sa10_reg[6]/NET0131  & n1606 ;
  assign n2181 = ~n2179 & ~n2180 ;
  assign n2182 = ~\sa10_reg[2]/P0001  & ~n2181 ;
  assign n2183 = ~\sa10_reg[1]/P0001  & \sa10_reg[2]/P0001  ;
  assign n2184 = n1583 & n1585 ;
  assign n2185 = n1598 & n1614 ;
  assign n2186 = ~n2184 & ~n2185 ;
  assign n2187 = ~n2156 & n2186 ;
  assign n2188 = n2183 & ~n2187 ;
  assign n2195 = ~n2182 & ~n2188 ;
  assign n2196 = ~n2194 & n2195 ;
  assign n2197 = ~n2178 & n2196 ;
  assign n2198 = ~n2108 & n2197 ;
  assign n2199 = ~n2140 & n2198 ;
  assign n2218 = ~\sa03_reg[6]/NET0131  & n1316 ;
  assign n2219 = n1376 & n1398 ;
  assign n2220 = ~n2218 & ~n2219 ;
  assign n2221 = ~\sa03_reg[2]/P0001  & ~n2220 ;
  assign n2215 = ~\sa03_reg[2]/P0001  & ~\sa03_reg[7]/NET0131  ;
  assign n2216 = n1326 & n1334 ;
  assign n2217 = ~n2215 & n2216 ;
  assign n2222 = ~n1565 & ~n2217 ;
  assign n2223 = ~n2221 & n2222 ;
  assign n2224 = \sa03_reg[1]/P0001  & ~n2223 ;
  assign n2229 = n1316 & n1367 ;
  assign n2230 = ~n1460 & ~n2229 ;
  assign n2231 = n1494 & ~n2230 ;
  assign n2226 = \sa03_reg[5]/P0001  & ~n1332 ;
  assign n2225 = ~\sa03_reg[2]/P0001  & ~\sa03_reg[3]/P0001  ;
  assign n2227 = ~n1341 & n2225 ;
  assign n2228 = n2226 & n2227 ;
  assign n2241 = ~\sa03_reg[0]/P0001  & ~n2228 ;
  assign n2242 = ~n2231 & n2241 ;
  assign n2232 = ~n1454 & ~n1515 ;
  assign n2233 = ~\sa03_reg[1]/P0001  & \sa03_reg[7]/NET0131  ;
  assign n2234 = ~n2232 & n2233 ;
  assign n2235 = \sa03_reg[2]/P0001  & n1425 ;
  assign n2243 = ~n2234 & ~n2235 ;
  assign n2244 = n2242 & n2243 ;
  assign n2236 = \sa03_reg[4]/P0001  & n1353 ;
  assign n2237 = ~n1414 & ~n2236 ;
  assign n2238 = n1374 & ~n2237 ;
  assign n2239 = ~n1400 & ~n1547 ;
  assign n2240 = ~\sa03_reg[2]/P0001  & ~n2239 ;
  assign n2245 = ~n2238 & ~n2240 ;
  assign n2246 = n2244 & n2245 ;
  assign n2247 = ~n2224 & n2246 ;
  assign n2260 = \sa03_reg[4]/P0001  & n1342 ;
  assign n2261 = ~n1482 & ~n1533 ;
  assign n2262 = ~n2260 & n2261 ;
  assign n2263 = ~\sa03_reg[2]/P0001  & ~n2262 ;
  assign n2267 = \sa03_reg[2]/P0001  & ~n1334 ;
  assign n2268 = n1318 & ~n1324 ;
  assign n2269 = ~n2267 & n2268 ;
  assign n2264 = ~\sa03_reg[4]/P0001  & n1367 ;
  assign n2265 = n1436 & n2264 ;
  assign n2266 = n1329 & n1423 ;
  assign n2270 = ~n2265 & ~n2266 ;
  assign n2271 = ~n2269 & n2270 ;
  assign n2272 = ~n2263 & n2271 ;
  assign n2273 = ~\sa03_reg[1]/P0001  & ~n2272 ;
  assign n2252 = ~n1398 & ~n1408 ;
  assign n2253 = ~\sa03_reg[7]/NET0131  & ~n2252 ;
  assign n2254 = ~n1368 & ~n1533 ;
  assign n2255 = ~n2253 & n2254 ;
  assign n2256 = \sa03_reg[2]/P0001  & ~n2255 ;
  assign n2248 = n1316 & n1326 ;
  assign n2249 = \sa03_reg[7]/NET0131  & n2248 ;
  assign n2250 = n1367 & n2225 ;
  assign n2251 = ~\sa03_reg[6]/NET0131  & n2250 ;
  assign n2257 = ~n2249 & ~n2251 ;
  assign n2258 = ~n2256 & n2257 ;
  assign n2259 = \sa03_reg[1]/P0001  & ~n2258 ;
  assign n2205 = \sa03_reg[7]/NET0131  & n1368 ;
  assign n2274 = ~n1364 & ~n2205 ;
  assign n2275 = ~\sa03_reg[3]/P0001  & ~n2274 ;
  assign n2276 = ~n1343 & ~n2275 ;
  assign n2277 = \sa03_reg[2]/P0001  & ~n2276 ;
  assign n2280 = n1482 & n2225 ;
  assign n2278 = n1374 & n1431 ;
  assign n2279 = n1334 & n1449 ;
  assign n2281 = \sa03_reg[0]/P0001  & ~n2279 ;
  assign n2282 = ~n2278 & n2281 ;
  assign n2283 = ~n2280 & n2282 ;
  assign n2284 = ~n2277 & n2283 ;
  assign n2285 = ~n2259 & n2284 ;
  assign n2286 = ~n2273 & n2285 ;
  assign n2287 = ~n2247 & ~n2286 ;
  assign n2200 = n1368 & n1376 ;
  assign n2201 = ~n1561 & ~n2200 ;
  assign n2202 = n1329 & ~n1330 ;
  assign n2203 = n2201 & ~n2202 ;
  assign n2204 = n1429 & ~n2203 ;
  assign n2206 = \sa03_reg[4]/P0001  & n1404 ;
  assign n2207 = ~n1416 & ~n2205 ;
  assign n2208 = ~n2206 & n2207 ;
  assign n2209 = ~\sa03_reg[3]/P0001  & ~n2208 ;
  assign n2210 = ~n1369 & ~n1446 ;
  assign n2211 = ~n2209 & n2210 ;
  assign n2212 = \sa03_reg[2]/P0001  & ~n2211 ;
  assign n2213 = ~n2204 & ~n2212 ;
  assign n2214 = \sa03_reg[1]/P0001  & ~n2213 ;
  assign n2288 = n1376 & n2218 ;
  assign n2289 = ~\sa03_reg[3]/P0001  & n1435 ;
  assign n2290 = ~\sa03_reg[4]/P0001  & n2289 ;
  assign n2291 = ~n2288 & ~n2290 ;
  assign n2292 = ~\sa03_reg[2]/P0001  & ~n2291 ;
  assign n2294 = ~n1325 & ~n1420 ;
  assign n2295 = ~n2249 & n2294 ;
  assign n2296 = \sa03_reg[2]/P0001  & ~n2295 ;
  assign n2297 = n1429 & n2264 ;
  assign n2293 = n1334 & n1339 ;
  assign n2298 = ~n2228 & ~n2293 ;
  assign n2299 = ~n2297 & n2298 ;
  assign n2300 = ~n2296 & n2299 ;
  assign n2301 = ~\sa03_reg[1]/P0001  & ~n2300 ;
  assign n2302 = ~n2292 & ~n2301 ;
  assign n2303 = ~n2214 & n2302 ;
  assign n2304 = ~n2287 & n2303 ;
  assign n2305 = n2199 & ~n2304 ;
  assign n2306 = ~n2199 & n2304 ;
  assign n2307 = ~n2305 & ~n2306 ;
  assign n2308 = ~n1581 & ~n2307 ;
  assign n2309 = n1581 & n2307 ;
  assign n2310 = ~n2308 & ~n2309 ;
  assign n2332 = ~\sa32_reg[3]/P0001  & n2060 ;
  assign n2333 = ~\sa32_reg[2]/P0001  & ~n2332 ;
  assign n2334 = \sa32_reg[7]/P0001  & n1912 ;
  assign n2335 = \sa32_reg[2]/P0001  & ~n2019 ;
  assign n2336 = ~n2334 & n2335 ;
  assign n2337 = ~n2333 & ~n2336 ;
  assign n2338 = ~n2024 & n2032 ;
  assign n2339 = ~n2337 & n2338 ;
  assign n2340 = ~\sa32_reg[1]/P0001  & ~n2339 ;
  assign n2316 = n1915 & n1995 ;
  assign n2317 = \sa32_reg[7]/P0001  & n2316 ;
  assign n2315 = \sa32_reg[4]/P0001  & n1981 ;
  assign n2318 = ~n1994 & ~n2315 ;
  assign n2319 = ~n2317 & n2318 ;
  assign n2320 = \sa32_reg[2]/P0001  & ~n2319 ;
  assign n2311 = n1920 & n1951 ;
  assign n2312 = ~n1936 & ~n2311 ;
  assign n2313 = ~\sa32_reg[2]/P0001  & ~\sa32_reg[3]/P0001  ;
  assign n2314 = n1955 & n2313 ;
  assign n2321 = n2312 & ~n2314 ;
  assign n2322 = ~n2320 & n2321 ;
  assign n2323 = \sa32_reg[1]/P0001  & ~n2322 ;
  assign n2324 = n1970 & n1981 ;
  assign n2325 = ~n1940 & ~n2324 ;
  assign n2326 = ~\sa32_reg[2]/P0001  & ~n2325 ;
  assign n2327 = \sa32_reg[4]/P0001  & n1969 ;
  assign n2328 = ~n1922 & ~n2327 ;
  assign n2329 = ~n1925 & ~n2033 ;
  assign n2330 = n2328 & n2329 ;
  assign n2331 = \sa32_reg[2]/P0001  & ~n2330 ;
  assign n2341 = ~n2326 & ~n2331 ;
  assign n2342 = ~n2323 & n2341 ;
  assign n2343 = ~n2340 & n2342 ;
  assign n2344 = \sa32_reg[0]/P0002  & ~n2343 ;
  assign n2378 = ~n1910 & ~n1990 ;
  assign n2379 = n1919 & ~n2378 ;
  assign n2375 = ~n1913 & n1924 ;
  assign n2376 = \sa32_reg[4]/P0001  & ~n1987 ;
  assign n2377 = n2375 & ~n2376 ;
  assign n2380 = ~\sa32_reg[2]/P0001  & ~n2377 ;
  assign n2381 = ~n2379 & n2380 ;
  assign n2383 = n1953 & n1965 ;
  assign n2382 = n1990 & n1995 ;
  assign n2384 = \sa32_reg[2]/P0001  & ~n2382 ;
  assign n2385 = ~n2383 & n2384 ;
  assign n2386 = ~n2381 & ~n2385 ;
  assign n2387 = ~\sa32_reg[5]/P0001  & \sa32_reg[7]/P0001  ;
  assign n2388 = n1951 & n2387 ;
  assign n2391 = ~\sa32_reg[1]/P0001  & ~n2324 ;
  assign n2392 = ~n2388 & n2391 ;
  assign n2364 = ~\sa32_reg[2]/P0001  & n2334 ;
  assign n2393 = ~n2061 & ~n2364 ;
  assign n2389 = ~\sa32_reg[3]/P0001  & n1923 ;
  assign n2390 = ~\sa32_reg[4]/P0001  & n2389 ;
  assign n2394 = ~n2383 & ~n2390 ;
  assign n2395 = n2393 & n2394 ;
  assign n2396 = n2392 & n2395 ;
  assign n2397 = \sa32_reg[2]/P0001  & ~\sa32_reg[3]/P0001  ;
  assign n2398 = \sa32_reg[4]/P0001  & n1920 ;
  assign n2399 = ~\sa32_reg[4]/P0001  & n2027 ;
  assign n2400 = ~n2398 & ~n2399 ;
  assign n2401 = n2397 & ~n2400 ;
  assign n2402 = ~\sa32_reg[2]/P0001  & n2033 ;
  assign n2403 = \sa32_reg[1]/P0001  & ~n2052 ;
  assign n2404 = ~n2402 & n2403 ;
  assign n2405 = ~n2401 & n2404 ;
  assign n2406 = ~n2396 & ~n2405 ;
  assign n2407 = ~n2386 & ~n2406 ;
  assign n2408 = ~\sa32_reg[0]/P0002  & ~n2407 ;
  assign n2352 = \sa32_reg[5]/P0001  & n1932 ;
  assign n2351 = ~\sa32_reg[5]/P0001  & n2315 ;
  assign n2353 = ~n2024 & ~n2351 ;
  assign n2354 = ~n2352 & n2353 ;
  assign n2355 = ~\sa32_reg[2]/P0001  & ~n2354 ;
  assign n2348 = \sa32_reg[2]/P0001  & ~\sa32_reg[4]/P0001  ;
  assign n2349 = n1913 & n2348 ;
  assign n2350 = \sa32_reg[3]/P0001  & n2349 ;
  assign n2346 = n1970 & n1987 ;
  assign n2347 = \sa32_reg[2]/P0001  & n2346 ;
  assign n2345 = n1909 & n1995 ;
  assign n2356 = n1912 & n1923 ;
  assign n2357 = ~n2345 & ~n2356 ;
  assign n2358 = ~n2347 & n2357 ;
  assign n2359 = ~n2350 & n2358 ;
  assign n2360 = ~n2355 & n2359 ;
  assign n2361 = ~\sa32_reg[1]/P0001  & ~n2360 ;
  assign n2365 = n1939 & n2364 ;
  assign n2362 = ~\sa32_reg[7]/P0001  & n1995 ;
  assign n2363 = n1990 & n2362 ;
  assign n2366 = n1924 & n1981 ;
  assign n2367 = n2046 & n2366 ;
  assign n2409 = ~n2363 & ~n2367 ;
  assign n2410 = ~n2010 & n2409 ;
  assign n2411 = ~n2365 & n2410 ;
  assign n2368 = ~\sa32_reg[2]/P0001  & n2063 ;
  assign n2369 = \sa32_reg[1]/P0001  & n2368 ;
  assign n2371 = ~n2028 & ~n2311 ;
  assign n2372 = ~n2362 & n2371 ;
  assign n2370 = \sa32_reg[1]/P0001  & \sa32_reg[2]/P0001  ;
  assign n2373 = ~\sa32_reg[6]/NET0131  & n2370 ;
  assign n2374 = ~n2372 & n2373 ;
  assign n2412 = ~n2369 & ~n2374 ;
  assign n2413 = n2411 & n2412 ;
  assign n2414 = ~n2361 & n2413 ;
  assign n2415 = ~n2408 & n2414 ;
  assign n2416 = ~n2344 & n2415 ;
  assign n2447 = ~\sa21_reg[6]/NET0131  & n1867 ;
  assign n2446 = n1754 & n1761 ;
  assign n2448 = ~\sa21_reg[2]/P0001  & ~\sa21_reg[7]/P0001  ;
  assign n2449 = n1837 & n2448 ;
  assign n2458 = ~n2446 & ~n2449 ;
  assign n2459 = ~n2447 & n2458 ;
  assign n2455 = ~\sa21_reg[2]/P0001  & \sa21_reg[4]/P0001  ;
  assign n2456 = ~n1772 & n2455 ;
  assign n2457 = ~n1823 & n2456 ;
  assign n2450 = \sa21_reg[6]/NET0131  & n1773 ;
  assign n2451 = ~\sa21_reg[7]/P0001  & n2450 ;
  assign n2452 = ~\sa21_reg[5]/P0001  & \sa21_reg[7]/P0001  ;
  assign n2453 = \sa21_reg[2]/P0001  & n1815 ;
  assign n2454 = n2452 & n2453 ;
  assign n2460 = ~n2451 & ~n2454 ;
  assign n2461 = ~n2457 & n2460 ;
  assign n2462 = n2459 & n2461 ;
  assign n2463 = ~\sa21_reg[1]/P0001  & ~n2462 ;
  assign n2437 = ~\sa21_reg[3]/P0001  & n1841 ;
  assign n2438 = ~n1779 & ~n2437 ;
  assign n2439 = ~n1753 & ~n1844 ;
  assign n2440 = n2438 & n2439 ;
  assign n2441 = \sa21_reg[1]/P0001  & ~n2440 ;
  assign n2436 = \sa21_reg[5]/P0001  & n1762 ;
  assign n2435 = \sa21_reg[7]/P0001  & n1890 ;
  assign n2442 = ~n1774 & ~n2435 ;
  assign n2443 = ~n2436 & n2442 ;
  assign n2444 = ~n2441 & n2443 ;
  assign n2445 = \sa21_reg[2]/P0001  & ~n2444 ;
  assign n2465 = n1802 & n1823 ;
  assign n2425 = ~\sa21_reg[5]/P0001  & n1763 ;
  assign n2466 = n1754 & n2425 ;
  assign n2467 = ~n2465 & ~n2466 ;
  assign n2468 = \sa21_reg[1]/P0001  & ~n2467 ;
  assign n2470 = n1754 & n1762 ;
  assign n2464 = n1759 & n1894 ;
  assign n2469 = n1745 & n1773 ;
  assign n2471 = ~n2464 & ~n2469 ;
  assign n2472 = ~n2470 & n2471 ;
  assign n2473 = ~n2468 & n2472 ;
  assign n2474 = ~n2445 & n2473 ;
  assign n2475 = ~n2463 & n2474 ;
  assign n2476 = \sa21_reg[0]/P0001  & ~n2475 ;
  assign n2417 = n1753 & n1784 ;
  assign n2418 = ~n1892 & ~n2417 ;
  assign n2419 = n1772 & ~n1793 ;
  assign n2420 = n2418 & ~n2419 ;
  assign n2421 = n1877 & ~n2420 ;
  assign n2422 = \sa21_reg[5]/P0001  & n1841 ;
  assign n2423 = ~n1822 & ~n2422 ;
  assign n2424 = ~\sa21_reg[4]/P0001  & ~n2423 ;
  assign n2426 = \sa21_reg[4]/P0001  & n2425 ;
  assign n2427 = ~n2424 & ~n2426 ;
  assign n2428 = ~\sa21_reg[3]/P0001  & ~n2427 ;
  assign n2429 = n1837 & n1854 ;
  assign n2430 = ~n1794 & ~n2429 ;
  assign n2431 = ~n2428 & n2430 ;
  assign n2432 = \sa21_reg[2]/P0001  & ~n2431 ;
  assign n2433 = ~n2421 & ~n2432 ;
  assign n2434 = \sa21_reg[1]/P0001  & ~n2433 ;
  assign n2492 = \sa21_reg[4]/P0001  & n1841 ;
  assign n2493 = \sa21_reg[5]/P0001  & n2492 ;
  assign n2489 = \sa21_reg[6]/NET0131  & n1849 ;
  assign n2490 = \sa21_reg[4]/P0001  & n2452 ;
  assign n2491 = ~\sa21_reg[1]/P0001  & n2490 ;
  assign n2494 = ~n2489 & ~n2491 ;
  assign n2495 = ~n2493 & n2494 ;
  assign n2496 = n1894 & ~n2495 ;
  assign n2477 = ~\sa21_reg[5]/P0001  & n1841 ;
  assign n2478 = \sa21_reg[2]/P0001  & n2477 ;
  assign n2479 = ~\sa21_reg[2]/P0001  & ~\sa21_reg[4]/P0001  ;
  assign n2480 = ~n1867 & ~n2479 ;
  assign n2481 = \sa21_reg[7]/P0001  & ~n2480 ;
  assign n2482 = ~n2478 & ~n2481 ;
  assign n2483 = ~\sa21_reg[1]/P0001  & ~n2482 ;
  assign n2487 = ~n1855 & ~n1864 ;
  assign n2488 = ~\sa21_reg[2]/P0001  & ~n2487 ;
  assign n2484 = ~n1781 & ~n1879 ;
  assign n2485 = n1754 & ~n2484 ;
  assign n2486 = n1786 & n1894 ;
  assign n2497 = ~n2485 & ~n2486 ;
  assign n2498 = ~n2488 & n2497 ;
  assign n2499 = ~n2483 & n2498 ;
  assign n2500 = ~n2496 & n2499 ;
  assign n2501 = ~\sa21_reg[0]/P0001  & ~n2500 ;
  assign n2503 = \sa21_reg[5]/P0001  & n2450 ;
  assign n2502 = n1832 & n1854 ;
  assign n2504 = ~n2465 & ~n2502 ;
  assign n2505 = ~n2503 & n2504 ;
  assign n2506 = \sa21_reg[2]/P0001  & ~n2505 ;
  assign n2507 = ~\sa21_reg[2]/P0001  & n1818 ;
  assign n2508 = n1749 & n1773 ;
  assign n2509 = ~n2507 & ~n2508 ;
  assign n2510 = ~n2485 & n2509 ;
  assign n2511 = ~n2506 & n2510 ;
  assign n2512 = ~\sa21_reg[1]/P0001  & ~n2511 ;
  assign n2516 = ~\sa21_reg[5]/P0001  & n2450 ;
  assign n2517 = ~n2448 & n2516 ;
  assign n2513 = n1761 & n1787 ;
  assign n2514 = ~n1747 & ~n2513 ;
  assign n2515 = ~\sa21_reg[2]/P0001  & ~n2514 ;
  assign n2518 = ~n1885 & ~n2515 ;
  assign n2519 = ~n2517 & n2518 ;
  assign n2520 = ~\sa21_reg[0]/P0001  & \sa21_reg[1]/P0001  ;
  assign n2521 = ~n2519 & n2520 ;
  assign n2522 = ~\sa21_reg[5]/P0001  & n1747 ;
  assign n2523 = ~n1891 & ~n2522 ;
  assign n2524 = n2448 & ~n2523 ;
  assign n2525 = ~n2521 & ~n2524 ;
  assign n2526 = ~n2512 & n2525 ;
  assign n2527 = ~n2501 & n2526 ;
  assign n2528 = ~n2434 & n2527 ;
  assign n2529 = ~n2476 & n2528 ;
  assign n2530 = \u0_w_reg[3][7]/P0001  & ~n2529 ;
  assign n2531 = ~\u0_w_reg[3][7]/P0001  & n2529 ;
  assign n2532 = ~n2530 & ~n2531 ;
  assign n2533 = n2416 & n2532 ;
  assign n2534 = ~n2416 & ~n2532 ;
  assign n2535 = ~n2533 & ~n2534 ;
  assign n2537 = n2310 & n2535 ;
  assign n2536 = ~n2310 & ~n2535 ;
  assign n2538 = ~\ld_r_reg/P0001  & ~n2536 ;
  assign n2539 = ~n2537 & n2538 ;
  assign n2541 = ~\text_in_r_reg[7]/P0001  & \u0_w_reg[3][7]/P0001  ;
  assign n2540 = \text_in_r_reg[7]/P0001  & ~\u0_w_reg[3][7]/P0001  ;
  assign n2542 = \ld_r_reg/P0001  & ~n2540 ;
  assign n2543 = ~n2541 & n2542 ;
  assign n2544 = ~n2539 & ~n2543 ;
  assign n2560 = \sa10_reg[2]/P0001  & ~n1682 ;
  assign n2561 = ~n2146 & n2560 ;
  assign n2559 = n1650 & n1669 ;
  assign n2558 = n1619 & n1650 ;
  assign n2562 = ~n1616 & ~n2558 ;
  assign n2563 = ~n2559 & n2562 ;
  assign n2564 = n2561 & n2563 ;
  assign n2566 = n1637 & n1681 ;
  assign n2567 = \sa10_reg[5]/P0001  & n2566 ;
  assign n2565 = n1590 & n1672 ;
  assign n2568 = ~\sa10_reg[2]/P0001  & ~n2128 ;
  assign n2569 = ~n2565 & n2568 ;
  assign n2570 = ~n2567 & n2569 ;
  assign n2571 = ~n2564 & ~n2570 ;
  assign n2572 = ~\sa10_reg[4]/P0001  & n1616 ;
  assign n2573 = ~\sa10_reg[1]/P0001  & ~n1683 ;
  assign n2574 = ~n2572 & n2573 ;
  assign n2575 = ~n2571 & n2574 ;
  assign n2576 = n1593 & n1661 ;
  assign n2577 = \sa10_reg[4]/P0001  & n2576 ;
  assign n2578 = \sa10_reg[1]/P0001  & ~n1665 ;
  assign n2579 = ~n2577 & n2578 ;
  assign n2580 = ~n2575 & ~n2579 ;
  assign n2545 = ~\sa10_reg[2]/P0001  & n2093 ;
  assign n2546 = \sa10_reg[4]/P0001  & n1585 ;
  assign n2547 = \sa10_reg[2]/P0001  & n2546 ;
  assign n2548 = ~n2545 & ~n2547 ;
  assign n2549 = \sa10_reg[3]/P0001  & ~n2548 ;
  assign n2550 = ~\sa10_reg[4]/P0001  & n1591 ;
  assign n2551 = ~n1654 & ~n1731 ;
  assign n2552 = ~n2550 & n2551 ;
  assign n2553 = ~\sa10_reg[2]/P0001  & ~n2552 ;
  assign n2554 = ~\sa10_reg[4]/P0001  & n1599 ;
  assign n2555 = ~n2156 & ~n2554 ;
  assign n2556 = ~n2553 & n2555 ;
  assign n2557 = \sa10_reg[1]/P0001  & ~n2556 ;
  assign n2644 = ~n2549 & ~n2557 ;
  assign n2645 = ~n2580 & n2644 ;
  assign n2582 = ~\sa10_reg[4]/P0001  & n1593 ;
  assign n2583 = \sa10_reg[7]/NET0131  & n2098 ;
  assign n2584 = ~n2582 & ~n2583 ;
  assign n2585 = ~\sa10_reg[2]/P0001  & ~n2584 ;
  assign n2581 = ~\sa10_reg[7]/NET0131  & n1651 ;
  assign n2586 = n1637 & n2112 ;
  assign n2587 = \sa10_reg[1]/P0001  & ~n2586 ;
  assign n2588 = ~n1727 & n2587 ;
  assign n2589 = ~n2581 & n2588 ;
  assign n2590 = ~n2585 & n2589 ;
  assign n2591 = n1666 & n1703 ;
  assign n2592 = ~\sa10_reg[1]/P0001  & ~n2591 ;
  assign n2594 = n1684 & n2112 ;
  assign n2595 = ~\sa10_reg[2]/P0001  & ~\sa10_reg[4]/P0001  ;
  assign n2596 = n1626 & n2595 ;
  assign n2593 = \sa10_reg[3]/P0001  & n1626 ;
  assign n2597 = ~n2566 & ~n2593 ;
  assign n2598 = ~n2596 & n2597 ;
  assign n2599 = ~n2594 & n2598 ;
  assign n2600 = n2592 & n2599 ;
  assign n2601 = ~n2590 & ~n2600 ;
  assign n2602 = \sa10_reg[2]/P0001  & ~n1599 ;
  assign n2603 = ~\sa10_reg[6]/NET0131  & n1627 ;
  assign n2604 = ~n1656 & ~n1713 ;
  assign n2605 = ~n2603 & n2604 ;
  assign n2606 = n2602 & n2605 ;
  assign n2608 = n1593 & n1627 ;
  assign n2607 = n1608 & n1681 ;
  assign n2609 = ~\sa10_reg[2]/P0001  & ~n2607 ;
  assign n2610 = ~n2608 & n2609 ;
  assign n2611 = ~n1731 & n2610 ;
  assign n2612 = ~n2606 & ~n2611 ;
  assign n2613 = ~n2601 & ~n2612 ;
  assign n2614 = \sa10_reg[0]/P0001  & ~n2613 ;
  assign n2618 = ~\sa10_reg[1]/P0001  & ~n2547 ;
  assign n2615 = \sa10_reg[5]/P0001  & n2147 ;
  assign n2616 = ~n1627 & ~n1722 ;
  assign n2617 = n1614 & ~n2616 ;
  assign n2619 = ~n2615 & ~n2617 ;
  assign n2620 = n2618 & n2619 ;
  assign n2625 = n1637 & n1650 ;
  assign n2626 = ~n1627 & n1699 ;
  assign n2627 = ~n2625 & ~n2626 ;
  assign n2628 = ~\sa10_reg[2]/P0001  & ~n2627 ;
  assign n2623 = \sa10_reg[4]/P0001  & n1608 ;
  assign n2624 = n1661 & n2623 ;
  assign n2621 = \sa10_reg[5]/P0001  & n1593 ;
  assign n2622 = \sa10_reg[2]/P0001  & n2621 ;
  assign n2629 = \sa10_reg[1]/P0001  & ~n1595 ;
  assign n2630 = ~n2622 & n2629 ;
  assign n2631 = ~n2624 & n2630 ;
  assign n2632 = ~n2628 & n2631 ;
  assign n2633 = ~n2620 & ~n2632 ;
  assign n2634 = n1612 & n1672 ;
  assign n2635 = ~\sa10_reg[2]/P0001  & n2634 ;
  assign n2636 = n1607 & n1722 ;
  assign n2637 = ~n2101 & ~n2636 ;
  assign n2638 = ~n2635 & n2637 ;
  assign n2639 = ~\sa10_reg[3]/P0001  & ~n2638 ;
  assign n2640 = \sa10_reg[2]/P0001  & n2180 ;
  assign n2641 = ~n2639 & ~n2640 ;
  assign n2642 = ~n2633 & n2641 ;
  assign n2643 = ~\sa10_reg[0]/P0001  & ~n2642 ;
  assign n2646 = ~n2614 & ~n2643 ;
  assign n2647 = n2645 & n2646 ;
  assign n2710 = \sa03_reg[5]/P0001  & n1332 ;
  assign n2711 = ~n1423 & n2710 ;
  assign n2712 = n1330 & n1355 ;
  assign n2713 = ~n2711 & ~n2712 ;
  assign n2714 = ~\sa03_reg[2]/P0001  & ~n2713 ;
  assign n2716 = n1367 & n1381 ;
  assign n2715 = \sa03_reg[2]/P0001  & n1435 ;
  assign n2717 = \sa03_reg[1]/P0001  & ~n1399 ;
  assign n2718 = ~n2715 & n2717 ;
  assign n2719 = ~n2716 & n2718 ;
  assign n2720 = ~n2714 & n2719 ;
  assign n2721 = ~\sa03_reg[2]/P0001  & ~n2289 ;
  assign n2722 = \sa03_reg[2]/P0001  & ~n2260 ;
  assign n2723 = ~n1460 & n2722 ;
  assign n2724 = ~n2721 & ~n2723 ;
  assign n2725 = ~\sa03_reg[1]/P0001  & ~n1563 ;
  assign n2726 = ~n2724 & n2725 ;
  assign n2727 = ~n2720 & ~n2726 ;
  assign n2704 = ~\sa03_reg[3]/P0001  & n1431 ;
  assign n2705 = ~n2288 & ~n2704 ;
  assign n2706 = \sa03_reg[2]/P0001  & ~n2705 ;
  assign n2707 = ~\sa03_reg[2]/P0001  & n1397 ;
  assign n2708 = ~n1416 & ~n2707 ;
  assign n2709 = ~\sa03_reg[3]/P0001  & ~n2708 ;
  assign n2728 = ~n2706 & ~n2709 ;
  assign n2729 = ~n2727 & n2728 ;
  assign n2730 = ~\sa03_reg[0]/P0001  & ~n2729 ;
  assign n2648 = ~n1319 & ~n2206 ;
  assign n2649 = ~\sa03_reg[2]/P0001  & ~n2648 ;
  assign n2650 = n1330 & n1384 ;
  assign n2651 = \sa03_reg[1]/P0001  & ~n2650 ;
  assign n2652 = ~n1417 & n2651 ;
  assign n2653 = ~n1461 & n2652 ;
  assign n2654 = ~n2649 & n2653 ;
  assign n2655 = n1330 & n1398 ;
  assign n2656 = ~\sa03_reg[1]/P0001  & ~n2655 ;
  assign n2657 = n2215 & n2218 ;
  assign n2661 = n2656 & ~n2657 ;
  assign n2658 = n1375 & n1384 ;
  assign n2659 = ~\sa03_reg[3]/P0001  & ~n1515 ;
  assign n2660 = n1339 & ~n2659 ;
  assign n2662 = ~n2658 & ~n2660 ;
  assign n2663 = n2661 & n2662 ;
  assign n2664 = ~n2654 & ~n2663 ;
  assign n2666 = ~\sa03_reg[3]/P0001  & n1341 ;
  assign n2665 = n1324 & n1332 ;
  assign n2667 = ~n1424 & ~n2665 ;
  assign n2668 = ~n2666 & n2667 ;
  assign n2669 = n1562 & n2668 ;
  assign n2670 = ~\sa03_reg[7]/NET0131  & n1541 ;
  assign n2671 = ~n1447 & n1538 ;
  assign n2672 = ~n2670 & n2671 ;
  assign n2673 = ~n2669 & ~n2672 ;
  assign n2674 = ~n2664 & ~n2673 ;
  assign n2675 = \sa03_reg[0]/P0001  & ~n2674 ;
  assign n2677 = n1449 & ~n2252 ;
  assign n2680 = \sa03_reg[2]/P0001  & ~n2266 ;
  assign n2681 = ~n2677 & n2680 ;
  assign n2678 = n1327 & n1455 ;
  assign n2679 = n1317 & n1355 ;
  assign n2682 = ~n2678 & ~n2679 ;
  assign n2683 = n2681 & n2682 ;
  assign n2684 = \sa03_reg[6]/NET0131  & \sa03_reg[7]/NET0131  ;
  assign n2685 = n1454 & n2684 ;
  assign n2686 = ~\sa03_reg[2]/P0001  & ~n1328 ;
  assign n2687 = ~n2216 & n2686 ;
  assign n2688 = ~n2685 & n2687 ;
  assign n2689 = ~n2683 & ~n2688 ;
  assign n2676 = ~\sa03_reg[3]/P0001  & n1416 ;
  assign n2690 = ~\sa03_reg[1]/P0001  & ~n1400 ;
  assign n2691 = ~n2676 & n2690 ;
  assign n2692 = ~n2689 & n2691 ;
  assign n2695 = ~n1354 & ~n1534 ;
  assign n2696 = ~n2670 & n2695 ;
  assign n2697 = ~\sa03_reg[2]/P0001  & ~n2696 ;
  assign n2698 = \sa03_reg[1]/P0001  & ~n1522 ;
  assign n2694 = n1436 & n1482 ;
  assign n2693 = n1367 & n1424 ;
  assign n2699 = ~n2249 & ~n2693 ;
  assign n2700 = ~n2694 & n2699 ;
  assign n2701 = n2698 & n2700 ;
  assign n2702 = ~n2697 & n2701 ;
  assign n2703 = ~n2692 & ~n2702 ;
  assign n2731 = ~\sa03_reg[2]/P0001  & ~n2200 ;
  assign n2732 = \sa03_reg[3]/P0001  & ~n2722 ;
  assign n2733 = ~n2731 & n2732 ;
  assign n2734 = ~n2703 & ~n2733 ;
  assign n2735 = ~n2675 & n2734 ;
  assign n2736 = ~n2730 & n2735 ;
  assign n2737 = n2647 & ~n2736 ;
  assign n2738 = ~n2647 & n2736 ;
  assign n2739 = ~n2737 & ~n2738 ;
  assign n2773 = ~n2168 & ~n2593 ;
  assign n2774 = \sa10_reg[2]/P0001  & ~n2773 ;
  assign n2754 = n1593 & n1668 ;
  assign n2775 = ~n1584 & ~n2754 ;
  assign n2776 = ~\sa10_reg[2]/P0001  & ~n2775 ;
  assign n2778 = n1597 & n1666 ;
  assign n2777 = n1594 & n1626 ;
  assign n2780 = ~n2565 & ~n2777 ;
  assign n2781 = ~n2778 & n2780 ;
  assign n2779 = ~n1638 & ~n2185 ;
  assign n2782 = ~n2179 & n2779 ;
  assign n2783 = n2781 & n2782 ;
  assign n2784 = ~n2776 & n2783 ;
  assign n2785 = ~n2774 & n2784 ;
  assign n2786 = \sa10_reg[1]/P0001  & ~n2785 ;
  assign n2787 = ~\sa10_reg[3]/P0001  & n1618 ;
  assign n2788 = ~n1601 & ~n2787 ;
  assign n2789 = ~n1668 & ~n2788 ;
  assign n2790 = ~\sa10_reg[4]/P0001  & n1614 ;
  assign n2791 = ~n2777 & ~n2790 ;
  assign n2792 = ~n2789 & n2791 ;
  assign n2793 = \sa10_reg[2]/P0001  & ~n2792 ;
  assign n2794 = ~n1651 & ~n1711 ;
  assign n2795 = \sa10_reg[7]/NET0131  & ~n2794 ;
  assign n2796 = ~n1698 & ~n2603 ;
  assign n2797 = n1722 & ~n2796 ;
  assign n2798 = ~n2795 & ~n2797 ;
  assign n2799 = ~\sa10_reg[1]/P0001  & ~n2798 ;
  assign n2800 = ~\sa10_reg[2]/P0001  & n1613 ;
  assign n2801 = ~n1602 & ~n2800 ;
  assign n2802 = ~n1611 & n2801 ;
  assign n2803 = ~n2799 & n2802 ;
  assign n2804 = ~n2793 & n2803 ;
  assign n2805 = ~n2786 & n2804 ;
  assign n2806 = ~\sa10_reg[0]/P0001  & ~n2805 ;
  assign n2759 = ~n1599 & ~n2621 ;
  assign n2760 = ~\sa10_reg[2]/P0001  & ~n2759 ;
  assign n2761 = n1664 & n1703 ;
  assign n2762 = ~n1682 & ~n2636 ;
  assign n2763 = ~n1592 & n2762 ;
  assign n2764 = ~n2761 & n2763 ;
  assign n2765 = ~n2760 & n2764 ;
  assign n2766 = ~\sa10_reg[1]/P0001  & ~n2765 ;
  assign n2741 = ~n1612 & n1634 ;
  assign n2742 = ~n1726 & ~n2741 ;
  assign n2743 = \sa10_reg[1]/P0001  & ~n2742 ;
  assign n2740 = ~\sa10_reg[4]/P0001  & n1629 ;
  assign n2744 = ~n1682 & ~n2608 ;
  assign n2745 = ~n2740 & n2744 ;
  assign n2746 = ~n2743 & n2745 ;
  assign n2747 = ~\sa10_reg[2]/P0001  & ~n2746 ;
  assign n2749 = n1597 & n1627 ;
  assign n2750 = ~n1631 & ~n2749 ;
  assign n2748 = \sa10_reg[7]/NET0131  & n1584 ;
  assign n2751 = ~n2581 & ~n2748 ;
  assign n2752 = n2750 & n2751 ;
  assign n2753 = \sa10_reg[1]/P0001  & ~n2752 ;
  assign n2755 = ~\sa10_reg[5]/P0001  & n2754 ;
  assign n2756 = ~n1592 & ~n2755 ;
  assign n2757 = \sa10_reg[2]/P0001  & ~n2756 ;
  assign n2758 = n1627 & n2621 ;
  assign n2767 = ~n2635 & ~n2758 ;
  assign n2768 = ~n2757 & n2767 ;
  assign n2769 = ~n2753 & n2768 ;
  assign n2770 = ~n2747 & n2769 ;
  assign n2771 = ~n2766 & n2770 ;
  assign n2772 = \sa10_reg[0]/P0001  & ~n2771 ;
  assign n2809 = \sa10_reg[6]/NET0131  & n1626 ;
  assign n2810 = ~n1593 & ~n1597 ;
  assign n2811 = ~\sa10_reg[5]/P0001  & ~n2810 ;
  assign n2812 = ~n2809 & ~n2811 ;
  assign n2813 = \sa10_reg[2]/P0001  & n1583 ;
  assign n2814 = ~n2812 & n2813 ;
  assign n2808 = n1582 & n2110 ;
  assign n2815 = ~n1730 & ~n2808 ;
  assign n2816 = ~n2814 & n2815 ;
  assign n2817 = ~\sa10_reg[1]/P0001  & ~n2816 ;
  assign n2818 = n1661 & n2168 ;
  assign n2819 = n1598 & n2790 ;
  assign n2820 = ~n2800 & ~n2819 ;
  assign n2821 = ~n2818 & n2820 ;
  assign n2822 = \sa10_reg[1]/P0001  & ~n2821 ;
  assign n2825 = ~\sa10_reg[1]/P0001  & ~\sa10_reg[2]/P0001  ;
  assign n2826 = n1626 & n1668 ;
  assign n2827 = ~n2634 & ~n2826 ;
  assign n2828 = ~n1683 & n2827 ;
  assign n2829 = n2825 & ~n2828 ;
  assign n2807 = \sa10_reg[5]/P0001  & n2761 ;
  assign n2823 = ~n1727 & ~n2565 ;
  assign n2824 = ~\sa10_reg[2]/P0001  & ~n2823 ;
  assign n2830 = ~n2807 & ~n2824 ;
  assign n2831 = ~n2829 & n2830 ;
  assign n2832 = ~n2822 & n2831 ;
  assign n2833 = ~n2817 & n2832 ;
  assign n2834 = ~n2772 & n2833 ;
  assign n2835 = ~n2806 & n2834 ;
  assign n2884 = \sa21_reg[3]/P0001  & n2492 ;
  assign n2885 = ~n1759 & ~n2884 ;
  assign n2886 = \sa21_reg[2]/P0001  & ~n2885 ;
  assign n2887 = n1877 & n2425 ;
  assign n2888 = ~n2429 & ~n2449 ;
  assign n2889 = ~n1782 & n2888 ;
  assign n2890 = ~n2887 & n2889 ;
  assign n2891 = ~n2886 & n2890 ;
  assign n2892 = ~\sa21_reg[1]/P0001  & ~n2891 ;
  assign n2878 = ~n1795 & ~n1833 ;
  assign n2879 = ~n1867 & n2878 ;
  assign n2880 = \sa21_reg[1]/P0001  & ~n2879 ;
  assign n2876 = n1753 & n1854 ;
  assign n2877 = ~n2429 & ~n2876 ;
  assign n2881 = ~n1879 & n2877 ;
  assign n2882 = ~n2880 & n2881 ;
  assign n2883 = ~\sa21_reg[2]/P0001  & ~n2882 ;
  assign n2893 = n1764 & n1773 ;
  assign n2896 = ~n1748 & ~n2893 ;
  assign n2894 = n1799 & n1844 ;
  assign n2842 = \sa21_reg[3]/P0001  & n1763 ;
  assign n2895 = ~\sa21_reg[4]/P0001  & n2842 ;
  assign n2897 = ~n2894 & ~n2895 ;
  assign n2898 = n2896 & n2897 ;
  assign n2899 = \sa21_reg[1]/P0001  & ~n2898 ;
  assign n2901 = n1758 & n1799 ;
  assign n2902 = ~\sa21_reg[4]/P0001  & n2901 ;
  assign n2903 = ~n1782 & ~n2902 ;
  assign n2904 = \sa21_reg[2]/P0001  & ~n2903 ;
  assign n2900 = n1823 & n2455 ;
  assign n2905 = ~\sa21_reg[4]/P0001  & n1854 ;
  assign n2906 = n1837 & n2905 ;
  assign n2907 = ~n2900 & ~n2906 ;
  assign n2908 = ~n2904 & n2907 ;
  assign n2909 = ~n2899 & n2908 ;
  assign n2910 = ~n2883 & n2909 ;
  assign n2911 = ~n2892 & n2910 ;
  assign n2912 = \sa21_reg[0]/P0001  & ~n2911 ;
  assign n2843 = ~\sa21_reg[3]/P0001  & n1775 ;
  assign n2844 = ~n1774 & ~n2842 ;
  assign n2845 = ~n2843 & n2844 ;
  assign n2846 = ~\sa21_reg[2]/P0001  & ~n2845 ;
  assign n2836 = ~n1750 & ~n2436 ;
  assign n2837 = \sa21_reg[2]/P0001  & ~n2836 ;
  assign n2840 = ~n1764 & ~n1838 ;
  assign n2841 = ~\sa21_reg[4]/P0001  & ~n2840 ;
  assign n2839 = \sa21_reg[4]/P0001  & n1750 ;
  assign n2838 = n1757 & n1758 ;
  assign n2847 = ~n2502 & ~n2838 ;
  assign n2848 = ~n2839 & n2847 ;
  assign n2849 = ~n2841 & n2848 ;
  assign n2850 = ~n2837 & n2849 ;
  assign n2851 = ~n2846 & n2850 ;
  assign n2852 = \sa21_reg[1]/P0001  & ~n2851 ;
  assign n2854 = ~n2426 & ~n2478 ;
  assign n2855 = ~\sa21_reg[3]/P0001  & ~n2854 ;
  assign n2853 = n1816 & n1837 ;
  assign n2856 = \sa21_reg[2]/P0001  & ~\sa21_reg[4]/P0001  ;
  assign n2857 = \sa21_reg[3]/P0001  & n1832 ;
  assign n2858 = n2856 & n2857 ;
  assign n2859 = ~n2853 & ~n2858 ;
  assign n2860 = ~n2855 & n2859 ;
  assign n2861 = ~\sa21_reg[1]/P0001  & ~n2860 ;
  assign n2863 = \sa21_reg[3]/P0001  & ~n1850 ;
  assign n2862 = ~\sa21_reg[4]/P0001  & n1841 ;
  assign n2864 = \sa21_reg[4]/P0001  & n1799 ;
  assign n2865 = n1758 & n2864 ;
  assign n2866 = ~n2862 & ~n2865 ;
  assign n2867 = ~n2863 & n2866 ;
  assign n2868 = \sa21_reg[2]/P0001  & ~n2867 ;
  assign n2869 = n1764 & n2455 ;
  assign n2870 = ~n1786 & ~n2869 ;
  assign n2871 = ~n1798 & n2870 ;
  assign n2872 = ~n2868 & n2871 ;
  assign n2873 = ~n2861 & n2872 ;
  assign n2874 = ~n2852 & n2873 ;
  assign n2875 = ~\sa21_reg[0]/P0001  & ~n2874 ;
  assign n2913 = ~n1780 & ~n1816 ;
  assign n2914 = \sa21_reg[5]/P0001  & ~n2913 ;
  assign n2915 = ~n1834 & ~n2914 ;
  assign n2916 = ~\sa21_reg[2]/P0001  & ~n2915 ;
  assign n2919 = ~n1804 & ~n2425 ;
  assign n2920 = ~\sa21_reg[3]/P0001  & ~n1781 ;
  assign n2921 = n2919 & n2920 ;
  assign n2917 = \sa21_reg[2]/P0001  & \sa21_reg[4]/P0001  ;
  assign n2918 = \sa21_reg[3]/P0001  & ~n1772 ;
  assign n2922 = n2917 & ~n2918 ;
  assign n2923 = ~n2921 & n2922 ;
  assign n2924 = ~n1865 & ~n2923 ;
  assign n2925 = ~n2916 & n2924 ;
  assign n2926 = ~\sa21_reg[1]/P0001  & ~n2925 ;
  assign n2930 = n1831 & n2436 ;
  assign n2929 = n1833 & n1854 ;
  assign n2931 = ~n2869 & ~n2929 ;
  assign n2932 = ~n2930 & n2931 ;
  assign n2933 = \sa21_reg[1]/P0001  & ~n2932 ;
  assign n2927 = n1755 & n1822 ;
  assign n2928 = n1747 & n1819 ;
  assign n2934 = ~n2927 & ~n2928 ;
  assign n2935 = ~n1881 & n2934 ;
  assign n2936 = ~n2933 & n2935 ;
  assign n2937 = ~n2926 & n2936 ;
  assign n2938 = ~n2875 & n2937 ;
  assign n2939 = ~n2912 & n2938 ;
  assign n2940 = n2835 & ~n2939 ;
  assign n2941 = ~n2835 & n2939 ;
  assign n2942 = ~n2940 & ~n2941 ;
  assign n2943 = \u0_w_reg[3][29]/P0001  & ~n2077 ;
  assign n2944 = ~\u0_w_reg[3][29]/P0001  & n2077 ;
  assign n2945 = ~n2943 & ~n2944 ;
  assign n2946 = n2942 & n2945 ;
  assign n2947 = ~n2942 & ~n2945 ;
  assign n2948 = ~n2946 & ~n2947 ;
  assign n2950 = n2739 & n2948 ;
  assign n2949 = ~n2739 & ~n2948 ;
  assign n2951 = ~\ld_r_reg/P0001  & ~n2949 ;
  assign n2952 = ~n2950 & n2951 ;
  assign n2954 = \text_in_r_reg[29]/P0001  & \u0_w_reg[3][29]/P0001  ;
  assign n2953 = ~\text_in_r_reg[29]/P0001  & ~\u0_w_reg[3][29]/P0001  ;
  assign n2955 = \ld_r_reg/P0001  & ~n2953 ;
  assign n2956 = ~n2954 & n2955 ;
  assign n2957 = ~n2952 & ~n2956 ;
  assign n2958 = n1738 & ~n1908 ;
  assign n2959 = ~n1738 & n1908 ;
  assign n2960 = ~n2958 & ~n2959 ;
  assign n2961 = ~n1479 & ~n2835 ;
  assign n2962 = n1479 & n2835 ;
  assign n2963 = ~n2961 & ~n2962 ;
  assign n2964 = \u0_w_reg[3][30]/P0001  & ~n2416 ;
  assign n2965 = ~\u0_w_reg[3][30]/P0001  & n2416 ;
  assign n2966 = ~n2964 & ~n2965 ;
  assign n2967 = n2963 & n2966 ;
  assign n2968 = ~n2963 & ~n2966 ;
  assign n2969 = ~n2967 & ~n2968 ;
  assign n2971 = n2960 & n2969 ;
  assign n2970 = ~n2960 & ~n2969 ;
  assign n2972 = ~\ld_r_reg/P0001  & ~n2970 ;
  assign n2973 = ~n2971 & n2972 ;
  assign n2975 = ~\text_in_r_reg[30]/P0001  & \u0_w_reg[3][30]/P0001  ;
  assign n2974 = \text_in_r_reg[30]/P0001  & ~\u0_w_reg[3][30]/P0001  ;
  assign n2976 = \ld_r_reg/P0001  & ~n2974 ;
  assign n2977 = ~n2975 & n2976 ;
  assign n2978 = ~n2973 & ~n2977 ;
  assign n3028 = ~\sa21_reg[2]/P0001  & n2884 ;
  assign n3030 = n1764 & n2917 ;
  assign n3026 = ~\sa21_reg[3]/P0001  & ~n2479 ;
  assign n3027 = n1749 & ~n3026 ;
  assign n3029 = n1822 & n1866 ;
  assign n3031 = ~n3027 & ~n3029 ;
  assign n3032 = ~n3030 & n3031 ;
  assign n3033 = ~n3028 & n3032 ;
  assign n3034 = ~\sa21_reg[1]/P0001  & ~n3033 ;
  assign n3018 = ~n1775 & ~n2426 ;
  assign n3019 = ~\sa21_reg[2]/P0001  & ~n3018 ;
  assign n3020 = n1841 & n1867 ;
  assign n3021 = n1763 & n2856 ;
  assign n3022 = ~n2894 & ~n3021 ;
  assign n3023 = ~n3020 & n3022 ;
  assign n3024 = ~n3019 & n3023 ;
  assign n3025 = \sa21_reg[1]/P0001  & ~n3024 ;
  assign n3035 = ~n1746 & ~n1781 ;
  assign n3036 = ~\sa21_reg[4]/P0001  & ~n3035 ;
  assign n3037 = \sa21_reg[2]/P0001  & ~n1788 ;
  assign n3038 = ~n2864 & n3037 ;
  assign n3039 = ~n3036 & n3038 ;
  assign n3040 = n1787 & n1822 ;
  assign n3041 = ~\sa21_reg[2]/P0001  & ~n2876 ;
  assign n3042 = ~n3040 & n3041 ;
  assign n3043 = ~n1883 & n3042 ;
  assign n3044 = ~n3039 & ~n3043 ;
  assign n3045 = ~n3025 & ~n3044 ;
  assign n3046 = ~n3034 & n3045 ;
  assign n3047 = \sa21_reg[0]/P0001  & ~n3046 ;
  assign n2992 = n1764 & ~n1866 ;
  assign n2993 = n1793 & n1832 ;
  assign n2994 = ~n2992 & ~n2993 ;
  assign n2995 = ~\sa21_reg[2]/P0001  & ~n2994 ;
  assign n2997 = \sa21_reg[6]/NET0131  & n1819 ;
  assign n2996 = n1831 & n2490 ;
  assign n2998 = ~n1780 & ~n2996 ;
  assign n2999 = ~n2997 & n2998 ;
  assign n3000 = ~n2995 & n2999 ;
  assign n3001 = \sa21_reg[1]/P0001  & ~n3000 ;
  assign n2988 = \sa21_reg[2]/P0001  & n1759 ;
  assign n2989 = ~n1880 & ~n2900 ;
  assign n2990 = ~n2988 & n2989 ;
  assign n2991 = ~\sa21_reg[3]/P0001  & ~n2990 ;
  assign n2979 = \sa21_reg[5]/P0001  & n2446 ;
  assign n2980 = \sa21_reg[3]/P0001  & n2862 ;
  assign n2981 = ~n2979 & ~n2980 ;
  assign n2982 = ~\sa21_reg[1]/P0001  & ~n2981 ;
  assign n2983 = ~n1853 & ~n2477 ;
  assign n2984 = ~\sa21_reg[1]/P0001  & ~n2983 ;
  assign n2985 = n1802 & n2477 ;
  assign n2986 = ~n2984 & ~n2985 ;
  assign n2987 = \sa21_reg[2]/P0001  & ~n2986 ;
  assign n3002 = ~n2982 & ~n2987 ;
  assign n3003 = ~n2991 & n3002 ;
  assign n3004 = ~n3001 & n3003 ;
  assign n3005 = ~\sa21_reg[0]/P0001  & ~n3004 ;
  assign n3054 = \sa21_reg[5]/P0001  & ~n2438 ;
  assign n3056 = n1802 & n2425 ;
  assign n3055 = n1757 & n1833 ;
  assign n3057 = ~n2447 & ~n3055 ;
  assign n3058 = ~n3056 & n3057 ;
  assign n3059 = ~n3054 & n3058 ;
  assign n3060 = \sa21_reg[2]/P0001  & ~n3059 ;
  assign n3050 = n1822 & n1867 ;
  assign n3051 = ~n2516 & ~n2838 ;
  assign n3052 = ~n3050 & n3051 ;
  assign n3053 = ~\sa21_reg[2]/P0001  & ~n3052 ;
  assign n3048 = ~\sa21_reg[7]/P0001  & n1815 ;
  assign n3049 = n1772 & n3048 ;
  assign n3061 = ~n1855 & ~n3049 ;
  assign n3062 = ~n3053 & n3061 ;
  assign n3063 = ~n3060 & n3062 ;
  assign n3064 = ~\sa21_reg[1]/P0001  & ~n3063 ;
  assign n3007 = ~n1842 & ~n1883 ;
  assign n3008 = ~n2853 & n3007 ;
  assign n3009 = ~\sa21_reg[2]/P0001  & ~n3008 ;
  assign n3010 = ~\sa21_reg[5]/P0001  & n2895 ;
  assign n3006 = n1762 & n1831 ;
  assign n3011 = ~n1820 & ~n2465 ;
  assign n3012 = ~n3006 & n3011 ;
  assign n3013 = ~n3010 & n3012 ;
  assign n3014 = ~n3009 & n3013 ;
  assign n3015 = \sa21_reg[1]/P0001  & ~n3014 ;
  assign n3016 = n1853 & n1894 ;
  assign n3017 = n1877 & n2417 ;
  assign n3065 = ~n3016 & ~n3017 ;
  assign n3066 = ~n3015 & n3065 ;
  assign n3067 = ~n3064 & n3066 ;
  assign n3068 = ~n3005 & n3067 ;
  assign n3069 = ~n3047 & n3068 ;
  assign n3070 = n2647 & ~n3069 ;
  assign n3071 = ~n2647 & n3069 ;
  assign n3072 = ~n3070 & ~n3071 ;
  assign n3073 = ~n1479 & ~n3072 ;
  assign n3074 = n1479 & n3072 ;
  assign n3075 = ~n3073 & ~n3074 ;
  assign n3076 = \u0_w_reg[3][21]/P0001  & ~n2077 ;
  assign n3077 = ~\u0_w_reg[3][21]/P0001  & n2077 ;
  assign n3078 = ~n3076 & ~n3077 ;
  assign n3079 = n2939 & n3078 ;
  assign n3080 = ~n2939 & ~n3078 ;
  assign n3081 = ~n3079 & ~n3080 ;
  assign n3083 = n3075 & n3081 ;
  assign n3082 = ~n3075 & ~n3081 ;
  assign n3084 = ~\ld_r_reg/P0001  & ~n3082 ;
  assign n3085 = ~n3083 & n3084 ;
  assign n3087 = ~\text_in_r_reg[21]/P0001  & \u0_w_reg[3][21]/P0001  ;
  assign n3086 = \text_in_r_reg[21]/P0001  & ~\u0_w_reg[3][21]/P0001  ;
  assign n3088 = \ld_r_reg/P0001  & ~n3086 ;
  assign n3089 = ~n3087 & n3088 ;
  assign n3090 = ~n3085 & ~n3089 ;
  assign n3091 = ~n1581 & ~n2942 ;
  assign n3092 = n1581 & n2942 ;
  assign n3093 = ~n3091 & ~n3092 ;
  assign n3094 = \u0_w_reg[3][22]/P0001  & ~n2416 ;
  assign n3095 = ~\u0_w_reg[3][22]/P0001  & n2416 ;
  assign n3096 = ~n3094 & ~n3095 ;
  assign n3097 = n1908 & n3096 ;
  assign n3098 = ~n1908 & ~n3096 ;
  assign n3099 = ~n3097 & ~n3098 ;
  assign n3101 = n3093 & n3099 ;
  assign n3100 = ~n3093 & ~n3099 ;
  assign n3102 = ~\ld_r_reg/P0001  & ~n3100 ;
  assign n3103 = ~n3101 & n3102 ;
  assign n3105 = ~\text_in_r_reg[22]/P0001  & \u0_w_reg[3][22]/P0001  ;
  assign n3104 = \text_in_r_reg[22]/P0001  & ~\u0_w_reg[3][22]/P0001  ;
  assign n3106 = \ld_r_reg/P0001  & ~n3104 ;
  assign n3107 = ~n3105 & n3106 ;
  assign n3108 = ~n3103 & ~n3107 ;
  assign n3109 = ~n2963 & ~n3069 ;
  assign n3110 = n2963 & n3069 ;
  assign n3111 = ~n3109 & ~n3110 ;
  assign n3129 = n1939 & n1951 ;
  assign n3130 = \sa32_reg[2]/P0001  & ~n3129 ;
  assign n3131 = ~n1911 & n3130 ;
  assign n3127 = ~n1919 & ~n1951 ;
  assign n3128 = n2041 & n3127 ;
  assign n3132 = ~n2332 & ~n3128 ;
  assign n3133 = n3131 & n3132 ;
  assign n3135 = ~n1948 & n1965 ;
  assign n3134 = n1951 & n2011 ;
  assign n3136 = ~\sa32_reg[2]/P0001  & ~n3134 ;
  assign n3137 = ~n3135 & n3136 ;
  assign n3138 = ~n3133 & ~n3137 ;
  assign n3126 = n1939 & n2362 ;
  assign n3139 = ~n2052 & ~n3126 ;
  assign n3140 = ~n3138 & n3139 ;
  assign n3141 = ~\sa32_reg[1]/P0001  & ~n3140 ;
  assign n3112 = ~n2363 & ~n2375 ;
  assign n3113 = ~n2013 & n3112 ;
  assign n3114 = ~\sa32_reg[2]/P0001  & ~n3113 ;
  assign n3116 = ~\sa32_reg[5]/P0001  & n1933 ;
  assign n3117 = \sa32_reg[3]/P0001  & n1963 ;
  assign n3115 = n2315 & n2397 ;
  assign n3118 = ~n2061 & ~n3115 ;
  assign n3119 = ~n3117 & n3118 ;
  assign n3120 = ~n3116 & n3119 ;
  assign n3121 = ~n3114 & n3120 ;
  assign n3122 = \sa32_reg[1]/P0001  & ~n3121 ;
  assign n3123 = n2030 & n2366 ;
  assign n3124 = \sa32_reg[4]/P0001  & n1909 ;
  assign n3125 = n2059 & n3124 ;
  assign n3201 = ~n3123 & ~n3125 ;
  assign n3202 = ~n3122 & n3201 ;
  assign n3203 = ~n3141 & n3202 ;
  assign n3143 = \sa32_reg[5]/P0001  & n1923 ;
  assign n3144 = ~n1951 & n3143 ;
  assign n3145 = ~\sa32_reg[5]/P0001  & n2049 ;
  assign n3146 = ~\sa32_reg[6]/NET0131  & n3145 ;
  assign n3147 = ~n3144 & ~n3146 ;
  assign n3148 = ~\sa32_reg[2]/P0001  & ~n3147 ;
  assign n3149 = \sa32_reg[4]/P0001  & n2387 ;
  assign n3150 = n2397 & n3149 ;
  assign n3151 = ~n2068 & ~n2327 ;
  assign n3152 = ~n3150 & n3151 ;
  assign n3153 = ~n3148 & n3152 ;
  assign n3154 = \sa32_reg[1]/P0001  & ~n3153 ;
  assign n3155 = n1909 & n2313 ;
  assign n3156 = ~n2004 & ~n3155 ;
  assign n3157 = ~\sa32_reg[7]/P0001  & ~n3156 ;
  assign n3158 = ~n1937 & ~n3124 ;
  assign n3159 = \sa32_reg[2]/P0001  & ~n3158 ;
  assign n3160 = ~n3157 & ~n3159 ;
  assign n3161 = ~\sa32_reg[1]/P0001  & ~n3160 ;
  assign n3162 = ~\sa32_reg[5]/P0001  & n1914 ;
  assign n3163 = ~n2316 & ~n3162 ;
  assign n3164 = \sa32_reg[2]/P0001  & ~n3163 ;
  assign n3142 = ~\sa32_reg[3]/P0001  & n1964 ;
  assign n3165 = ~n3126 & ~n3142 ;
  assign n3166 = ~n3164 & n3165 ;
  assign n3167 = ~n3161 & n3166 ;
  assign n3168 = ~n3154 & n3167 ;
  assign n3169 = ~\sa32_reg[0]/P0002  & ~n3168 ;
  assign n3170 = ~\sa32_reg[3]/P0001  & ~n2030 ;
  assign n3171 = n1920 & ~n3170 ;
  assign n3172 = n1947 & n2049 ;
  assign n3173 = ~\sa32_reg[1]/P0001  & ~n3172 ;
  assign n3176 = ~n3171 & n3173 ;
  assign n3174 = \sa32_reg[2]/P0001  & n2024 ;
  assign n3175 = ~\sa32_reg[2]/P0001  & n1914 ;
  assign n3177 = ~n3174 & ~n3175 ;
  assign n3178 = n3176 & n3177 ;
  assign n3180 = ~\sa32_reg[4]/P0001  & n1981 ;
  assign n3181 = n1953 & n1990 ;
  assign n3182 = ~n3180 & ~n3181 ;
  assign n3183 = ~\sa32_reg[2]/P0001  & ~n3182 ;
  assign n3179 = \sa32_reg[1]/P0001  & ~n2063 ;
  assign n3184 = n1923 & n2348 ;
  assign n3185 = ~n1938 & ~n3184 ;
  assign n3186 = n3179 & n3185 ;
  assign n3187 = ~n3183 & n3186 ;
  assign n3188 = ~n3178 & ~n3187 ;
  assign n3190 = \sa32_reg[2]/P0001  & ~n1925 ;
  assign n3189 = ~\sa32_reg[7]/P0001  & n1919 ;
  assign n3191 = ~n2004 & ~n2346 ;
  assign n3192 = ~n3189 & n3191 ;
  assign n3193 = n3190 & n3192 ;
  assign n3194 = n1924 & n1987 ;
  assign n3195 = ~\sa32_reg[2]/P0001  & ~n1949 ;
  assign n3196 = ~n3194 & n3195 ;
  assign n3197 = ~n2363 & n3196 ;
  assign n3198 = ~n3193 & ~n3197 ;
  assign n3199 = ~n3188 & ~n3198 ;
  assign n3200 = \sa32_reg[0]/P0002  & ~n3199 ;
  assign n3204 = ~n3169 & ~n3200 ;
  assign n3205 = n3203 & n3204 ;
  assign n3206 = \u0_w_reg[3][13]/P0001  & ~n3205 ;
  assign n3207 = ~\u0_w_reg[3][13]/P0001  & n3205 ;
  assign n3208 = ~n3206 & ~n3207 ;
  assign n3209 = n2077 & n3208 ;
  assign n3210 = ~n2077 & ~n3208 ;
  assign n3211 = ~n3209 & ~n3210 ;
  assign n3213 = n3111 & n3211 ;
  assign n3212 = ~n3111 & ~n3211 ;
  assign n3214 = ~\ld_r_reg/P0001  & ~n3212 ;
  assign n3215 = ~n3213 & n3214 ;
  assign n3217 = \text_in_r_reg[13]/P0001  & \u0_w_reg[3][13]/P0001  ;
  assign n3216 = ~\text_in_r_reg[13]/P0001  & ~\u0_w_reg[3][13]/P0001  ;
  assign n3218 = \ld_r_reg/P0001  & ~n3216 ;
  assign n3219 = ~n3217 & n3218 ;
  assign n3220 = ~n3215 & ~n3219 ;
  assign n3221 = ~n1741 & ~n2939 ;
  assign n3222 = n1741 & n2939 ;
  assign n3223 = ~n3221 & ~n3222 ;
  assign n3224 = \u0_w_reg[3][14]/P0001  & ~n2416 ;
  assign n3225 = ~\u0_w_reg[3][14]/P0001  & n2416 ;
  assign n3226 = ~n3224 & ~n3225 ;
  assign n3227 = n2077 & n3226 ;
  assign n3228 = ~n2077 & ~n3226 ;
  assign n3229 = ~n3227 & ~n3228 ;
  assign n3231 = n3223 & n3229 ;
  assign n3230 = ~n3223 & ~n3229 ;
  assign n3232 = ~\ld_r_reg/P0001  & ~n3230 ;
  assign n3233 = ~n3231 & n3232 ;
  assign n3235 = \text_in_r_reg[14]/P0001  & \u0_w_reg[3][14]/P0001  ;
  assign n3234 = ~\text_in_r_reg[14]/P0001  & ~\u0_w_reg[3][14]/P0001  ;
  assign n3236 = \ld_r_reg/P0001  & ~n3234 ;
  assign n3237 = ~n3235 & n3236 ;
  assign n3238 = ~n3233 & ~n3237 ;
  assign n3258 = ~n1963 & ~n1978 ;
  assign n3259 = ~n2009 & n3258 ;
  assign n3260 = \sa32_reg[2]/P0001  & ~n3259 ;
  assign n3253 = n2041 & n2313 ;
  assign n3254 = \sa32_reg[4]/P0001  & n3253 ;
  assign n3255 = \sa32_reg[5]/P0001  & ~n1923 ;
  assign n3256 = n1951 & ~n3255 ;
  assign n3257 = n1934 & n1995 ;
  assign n3261 = ~n3256 & ~n3257 ;
  assign n3262 = ~n3254 & n3261 ;
  assign n3263 = ~n3260 & n3262 ;
  assign n3264 = ~\sa32_reg[1]/P0001  & ~n3263 ;
  assign n3250 = ~n1941 & ~n3146 ;
  assign n3251 = n2312 & n3250 ;
  assign n3252 = \sa32_reg[2]/P0001  & ~n3251 ;
  assign n3239 = ~n1909 & ~n1937 ;
  assign n3240 = ~\sa32_reg[2]/P0001  & ~n3239 ;
  assign n3241 = ~n2351 & ~n3240 ;
  assign n3242 = \sa32_reg[1]/P0001  & ~n3241 ;
  assign n3245 = n1909 & n1953 ;
  assign n3246 = n1919 & n1934 ;
  assign n3247 = ~n3245 & ~n3246 ;
  assign n3248 = ~\sa32_reg[2]/P0001  & ~n3247 ;
  assign n3243 = ~n1915 & ~n1948 ;
  assign n3244 = n2026 & ~n3243 ;
  assign n3249 = ~\sa32_reg[3]/P0001  & n1910 ;
  assign n3265 = ~n3244 & ~n3249 ;
  assign n3266 = ~n3116 & n3265 ;
  assign n3267 = ~n3248 & n3266 ;
  assign n3268 = ~n3242 & n3267 ;
  assign n3269 = ~n3252 & n3268 ;
  assign n3270 = ~n3264 & n3269 ;
  assign n3271 = \sa32_reg[0]/P0002  & ~n3270 ;
  assign n3305 = ~n1970 & n1982 ;
  assign n3306 = ~n3126 & ~n3305 ;
  assign n3307 = ~\sa32_reg[2]/P0001  & ~n3306 ;
  assign n3302 = \sa32_reg[7]/P0001  & n2382 ;
  assign n3303 = ~n2345 & ~n3302 ;
  assign n3304 = \sa32_reg[2]/P0001  & ~n3303 ;
  assign n3308 = n1934 & n2026 ;
  assign n3309 = n1954 & n3308 ;
  assign n3310 = ~\sa32_reg[1]/P0001  & ~n3309 ;
  assign n3311 = ~n2062 & n3310 ;
  assign n3312 = ~n3304 & n3311 ;
  assign n3313 = ~n3307 & n3312 ;
  assign n3314 = ~n2040 & ~n3115 ;
  assign n3315 = ~\sa32_reg[5]/P0001  & ~n3314 ;
  assign n3316 = n2041 & n2059 ;
  assign n3317 = ~\sa32_reg[2]/P0001  & n1921 ;
  assign n3318 = ~n3316 & ~n3317 ;
  assign n3319 = n3179 & n3318 ;
  assign n3320 = ~n3315 & n3319 ;
  assign n3321 = ~n3313 & ~n3320 ;
  assign n3274 = ~n1915 & ~n2060 ;
  assign n3275 = n1951 & ~n3274 ;
  assign n3272 = ~\sa32_reg[1]/P0001  & n1920 ;
  assign n3273 = ~n1947 & n3272 ;
  assign n3276 = \sa32_reg[2]/P0001  & ~n3273 ;
  assign n3277 = ~n3275 & n3276 ;
  assign n3278 = \sa32_reg[7]/P0001  & n1947 ;
  assign n3279 = \sa32_reg[5]/P0001  & n3278 ;
  assign n3280 = ~n1941 & ~n3279 ;
  assign n3281 = ~\sa32_reg[2]/P0001  & ~n2382 ;
  assign n3282 = n3280 & n3281 ;
  assign n3283 = ~n3277 & ~n3282 ;
  assign n3286 = \sa32_reg[3]/P0001  & n2068 ;
  assign n3284 = n1947 & n1953 ;
  assign n3288 = \sa32_reg[1]/P0001  & ~n3284 ;
  assign n3285 = n2313 & n2387 ;
  assign n3287 = ~n1912 & n1913 ;
  assign n3289 = ~n3285 & ~n3287 ;
  assign n3290 = n3288 & n3289 ;
  assign n3291 = ~n3286 & n3290 ;
  assign n3292 = n1915 & n1948 ;
  assign n3293 = ~n2346 & ~n3292 ;
  assign n3294 = ~\sa32_reg[3]/P0001  & ~n3293 ;
  assign n3295 = ~\sa32_reg[1]/P0001  & ~n3175 ;
  assign n3296 = ~n3294 & n3295 ;
  assign n3297 = ~n3291 & ~n3296 ;
  assign n3298 = ~n3283 & ~n3297 ;
  assign n3299 = ~\sa32_reg[0]/P0002  & ~n3298 ;
  assign n3300 = n1995 & n2068 ;
  assign n3301 = ~\sa32_reg[2]/P0001  & n3284 ;
  assign n3322 = ~n3300 & ~n3301 ;
  assign n3323 = ~n3299 & n3322 ;
  assign n3324 = ~n3321 & n3323 ;
  assign n3325 = ~n3271 & n3324 ;
  assign n3374 = \sa32_reg[4]/P0001  & n1990 ;
  assign n3375 = ~n1954 & ~n3374 ;
  assign n3376 = ~\sa32_reg[3]/P0001  & n1913 ;
  assign n3377 = ~n1969 & ~n3376 ;
  assign n3378 = n3375 & n3377 ;
  assign n3379 = \sa32_reg[2]/P0001  & ~n3378 ;
  assign n3380 = ~n3117 & ~n3253 ;
  assign n3381 = ~n3379 & n3380 ;
  assign n3382 = \sa32_reg[1]/P0001  & ~n3381 ;
  assign n3363 = \sa32_reg[4]/P0001  & ~n1939 ;
  assign n3364 = ~n1988 & n3363 ;
  assign n3365 = ~n1910 & ~n3364 ;
  assign n3366 = ~\sa32_reg[2]/P0001  & ~n3365 ;
  assign n3367 = ~\sa32_reg[5]/P0001  & n2050 ;
  assign n3368 = \sa32_reg[2]/P0001  & n3367 ;
  assign n3369 = n1982 & ~n2348 ;
  assign n3370 = ~n3129 & ~n3369 ;
  assign n3371 = ~n3368 & n3370 ;
  assign n3372 = ~n3366 & n3371 ;
  assign n3373 = ~\sa32_reg[1]/P0001  & ~n3372 ;
  assign n3356 = ~\sa32_reg[5]/P0001  & n1951 ;
  assign n3357 = ~n2050 & ~n3356 ;
  assign n3358 = \sa32_reg[6]/NET0131  & ~n3357 ;
  assign n3359 = ~n1940 & ~n1978 ;
  assign n3360 = ~n3358 & n3359 ;
  assign n3361 = \sa32_reg[2]/P0001  & ~n3360 ;
  assign n3362 = n2313 & n2315 ;
  assign n3383 = ~n3246 & ~n3362 ;
  assign n3384 = ~n3361 & n3383 ;
  assign n3385 = ~n3373 & n3384 ;
  assign n3386 = ~n3382 & n3385 ;
  assign n3387 = \sa32_reg[0]/P0002  & ~n3386 ;
  assign n3342 = ~\sa32_reg[6]/NET0131  & n1912 ;
  assign n3343 = ~n2366 & ~n3342 ;
  assign n3344 = ~\sa32_reg[2]/P0001  & ~n3343 ;
  assign n3345 = \sa32_reg[4]/P0001  & n1915 ;
  assign n3346 = n2397 & n3345 ;
  assign n3347 = ~n2352 & ~n2383 ;
  assign n3348 = ~n3346 & n3347 ;
  assign n3349 = ~n3344 & n3348 ;
  assign n3350 = \sa32_reg[1]/P0001  & ~n3349 ;
  assign n3337 = ~n2012 & ~n3257 ;
  assign n3338 = ~\sa32_reg[6]/NET0131  & n2028 ;
  assign n3339 = ~n2052 & ~n3338 ;
  assign n3340 = n3337 & n3339 ;
  assign n3341 = ~\sa32_reg[2]/P0001  & ~n3340 ;
  assign n3326 = n2059 & n3149 ;
  assign n3327 = ~n1952 & ~n2030 ;
  assign n3328 = \sa32_reg[7]/P0001  & ~n3327 ;
  assign n3329 = ~n3326 & ~n3328 ;
  assign n3330 = ~\sa32_reg[1]/P0001  & ~n3329 ;
  assign n3331 = \sa32_reg[4]/P0001  & n2060 ;
  assign n3332 = ~n3245 & ~n3331 ;
  assign n3333 = n2059 & ~n3332 ;
  assign n3334 = \sa32_reg[1]/P0001  & ~n1951 ;
  assign n3335 = \sa32_reg[2]/P0001  & n1937 ;
  assign n3336 = ~n3334 & n3335 ;
  assign n3351 = ~n3333 & ~n3336 ;
  assign n3352 = ~n3330 & n3351 ;
  assign n3353 = ~n3341 & n3352 ;
  assign n3354 = ~n3350 & n3353 ;
  assign n3355 = ~\sa32_reg[0]/P0002  & ~n3354 ;
  assign n3404 = \sa32_reg[7]/P0001  & ~n3375 ;
  assign n3405 = n1913 & n1970 ;
  assign n3406 = ~n3404 & ~n3405 ;
  assign n3407 = ~\sa32_reg[3]/P0001  & ~n3406 ;
  assign n3408 = n1954 & n2387 ;
  assign n3409 = ~n1911 & ~n3408 ;
  assign n3410 = ~n3407 & n3409 ;
  assign n3411 = n2370 & ~n3410 ;
  assign n3388 = \sa32_reg[2]/P0001  & ~n1921 ;
  assign n3389 = ~n1921 & ~n2388 ;
  assign n3390 = n3337 & n3389 ;
  assign n3391 = ~n3388 & ~n3390 ;
  assign n3392 = ~\sa32_reg[3]/P0001  & n3124 ;
  assign n3393 = ~n1992 & ~n3117 ;
  assign n3394 = ~n3392 & n3393 ;
  assign n3395 = \sa32_reg[2]/P0001  & ~n3394 ;
  assign n3396 = ~n3391 & ~n3395 ;
  assign n3397 = ~\sa32_reg[1]/P0001  & ~n3396 ;
  assign n3398 = ~n1996 & ~n3162 ;
  assign n3399 = ~\sa32_reg[2]/P0001  & ~n3398 ;
  assign n3400 = n1939 & ~n2049 ;
  assign n3401 = n3293 & ~n3400 ;
  assign n3402 = \sa32_reg[1]/P0001  & n2026 ;
  assign n3403 = ~n3401 & n3402 ;
  assign n3412 = ~n3399 & ~n3403 ;
  assign n3413 = ~n3397 & n3412 ;
  assign n3414 = ~n3411 & n3413 ;
  assign n3415 = ~n3355 & n3414 ;
  assign n3416 = ~n3387 & n3415 ;
  assign n3417 = n3325 & ~n3416 ;
  assign n3418 = ~n3325 & n3416 ;
  assign n3419 = ~n3417 & ~n3418 ;
  assign n3438 = ~n2317 & ~n2351 ;
  assign n3439 = ~\sa32_reg[2]/P0001  & ~n3438 ;
  assign n3435 = ~n3194 & ~n3249 ;
  assign n3436 = \sa32_reg[2]/P0001  & ~n3435 ;
  assign n3437 = n1924 & n2315 ;
  assign n3440 = ~n3134 & ~n3437 ;
  assign n3441 = ~n3436 & n3440 ;
  assign n3442 = ~n3439 & n3441 ;
  assign n3443 = ~\sa32_reg[1]/P0001  & ~n3442 ;
  assign n3423 = \sa32_reg[3]/P0001  & n3345 ;
  assign n3422 = ~\sa32_reg[4]/P0001  & n1990 ;
  assign n3424 = ~n2389 & ~n3422 ;
  assign n3425 = ~n3423 & n3424 ;
  assign n3426 = ~\sa32_reg[2]/P0001  & ~n3425 ;
  assign n3420 = ~n2012 & ~n2398 ;
  assign n3421 = \sa32_reg[2]/P0001  & ~n3420 ;
  assign n3427 = n1950 & ~n1992 ;
  assign n3428 = ~n3421 & n3427 ;
  assign n3429 = ~n3426 & n3428 ;
  assign n3430 = \sa32_reg[1]/P0001  & ~n3429 ;
  assign n3433 = ~n1941 & ~n3134 ;
  assign n3434 = ~\sa32_reg[2]/P0001  & ~n3433 ;
  assign n3431 = ~n2009 & ~n2362 ;
  assign n3432 = \sa32_reg[2]/P0001  & ~n3431 ;
  assign n3444 = ~n2040 & ~n2062 ;
  assign n3445 = ~n3432 & n3444 ;
  assign n3446 = ~n3434 & n3445 ;
  assign n3447 = ~n3430 & n3446 ;
  assign n3448 = ~n3443 & n3447 ;
  assign n3449 = ~\sa32_reg[0]/P0002  & ~n3448 ;
  assign n3470 = ~\sa32_reg[1]/P0001  & n1994 ;
  assign n3469 = n1988 & ~n2030 ;
  assign n3471 = ~n3331 & ~n3469 ;
  assign n3472 = ~n3470 & n3471 ;
  assign n3473 = ~\sa32_reg[3]/P0001  & ~n3472 ;
  assign n3465 = ~n2352 & ~n3292 ;
  assign n3466 = ~n3249 & ~n3331 ;
  assign n3467 = n3465 & n3466 ;
  assign n3468 = ~\sa32_reg[2]/P0001  & ~n3467 ;
  assign n3474 = n1932 & ~n2348 ;
  assign n3475 = ~n1935 & ~n3292 ;
  assign n3476 = ~n3474 & n3475 ;
  assign n3477 = ~\sa32_reg[1]/P0001  & ~n3476 ;
  assign n3478 = ~n3468 & ~n3477 ;
  assign n3479 = ~n3473 & n3478 ;
  assign n3480 = \sa32_reg[0]/P0002  & ~n3479 ;
  assign n3450 = n1909 & n2334 ;
  assign n3451 = ~n3408 & ~n3450 ;
  assign n3452 = ~n3145 & ~n3278 ;
  assign n3453 = ~n3345 & n3452 ;
  assign n3454 = \sa32_reg[2]/P0001  & ~n3453 ;
  assign n3455 = n3451 & ~n3454 ;
  assign n3456 = \sa32_reg[0]/P0002  & ~n3455 ;
  assign n3457 = ~\sa32_reg[3]/P0001  & n1939 ;
  assign n3458 = ~n2033 & ~n3457 ;
  assign n3459 = ~n1953 & ~n3458 ;
  assign n3460 = ~n1992 & ~n2324 ;
  assign n3461 = ~n3459 & n3460 ;
  assign n3462 = ~\sa32_reg[2]/P0001  & ~n3461 ;
  assign n3463 = ~n3456 & ~n3462 ;
  assign n3464 = \sa32_reg[1]/P0001  & ~n3463 ;
  assign n3491 = ~\sa32_reg[3]/P0001  & n2041 ;
  assign n3492 = ~n1922 & ~n2040 ;
  assign n3493 = ~n3491 & n3492 ;
  assign n3494 = \sa32_reg[2]/P0001  & ~n3493 ;
  assign n3487 = ~n2311 & ~n2366 ;
  assign n3488 = ~n1938 & n3487 ;
  assign n3489 = ~\sa32_reg[2]/P0001  & ~n3488 ;
  assign n3490 = n1990 & n2334 ;
  assign n3495 = ~n1936 & ~n3490 ;
  assign n3496 = ~n3489 & n3495 ;
  assign n3497 = ~n3494 & n3496 ;
  assign n3498 = ~\sa32_reg[1]/P0001  & ~n3497 ;
  assign n3481 = n1988 & ~n3127 ;
  assign n3482 = \sa32_reg[3]/P0001  & n3124 ;
  assign n3483 = ~n3481 & ~n3482 ;
  assign n3484 = n2370 & ~n3483 ;
  assign n3485 = ~n2033 & ~n3181 ;
  assign n3486 = n2059 & ~n3485 ;
  assign n3499 = ~n3484 & ~n3486 ;
  assign n3500 = ~n3498 & n3499 ;
  assign n3501 = ~n3464 & n3500 ;
  assign n3502 = ~n3480 & n3501 ;
  assign n3503 = ~n3449 & n3502 ;
  assign n3504 = \u0_w_reg[3][9]/P0001  & ~n3503 ;
  assign n3505 = ~\u0_w_reg[3][9]/P0001  & n3503 ;
  assign n3506 = ~n3504 & ~n3505 ;
  assign n3507 = n3419 & n3506 ;
  assign n3508 = ~n3419 & ~n3506 ;
  assign n3509 = ~n3507 & ~n3508 ;
  assign n3537 = ~n1834 & ~n1872 ;
  assign n3538 = ~n2436 & n3537 ;
  assign n3539 = \sa21_reg[2]/P0001  & ~n3538 ;
  assign n3542 = ~\sa21_reg[6]/NET0131  & n1757 ;
  assign n3543 = ~\sa21_reg[5]/P0001  & n3542 ;
  assign n3544 = n2455 & n3543 ;
  assign n3540 = \sa21_reg[5]/P0001  & ~n1763 ;
  assign n3541 = n1866 & ~n3540 ;
  assign n3545 = n1745 & n1815 ;
  assign n3546 = ~n3541 & ~n3545 ;
  assign n3547 = ~n3544 & n3546 ;
  assign n3548 = ~n3539 & n3547 ;
  assign n3549 = ~\sa21_reg[1]/P0001  & ~n3548 ;
  assign n3554 = \sa21_reg[3]/P0001  & n1758 ;
  assign n3555 = ~\sa21_reg[2]/P0001  & ~n3554 ;
  assign n3556 = ~n2469 & ~n2905 ;
  assign n3557 = ~n2489 & n3556 ;
  assign n3558 = n3555 & n3557 ;
  assign n3559 = \sa21_reg[2]/P0001  & ~n2993 ;
  assign n3560 = ~n2893 & n3559 ;
  assign n3561 = n1752 & n3560 ;
  assign n3562 = ~n3558 & ~n3561 ;
  assign n3550 = ~n1837 & ~n2477 ;
  assign n3551 = ~\sa21_reg[2]/P0001  & ~n3550 ;
  assign n3552 = ~n1884 & ~n3551 ;
  assign n3553 = \sa21_reg[1]/P0001  & ~n3552 ;
  assign n3563 = ~n1838 & ~n3010 ;
  assign n3564 = ~n3553 & n3563 ;
  assign n3565 = ~n3562 & n3564 ;
  assign n3566 = ~n3549 & n3565 ;
  assign n3567 = \sa21_reg[0]/P0001  & ~n3566 ;
  assign n3510 = \sa21_reg[6]/NET0131  & n1750 ;
  assign n3511 = ~n2893 & ~n3510 ;
  assign n3512 = ~\sa21_reg[3]/P0001  & n1833 ;
  assign n3513 = n3511 & ~n3512 ;
  assign n3514 = ~\sa21_reg[2]/P0001  & ~n3513 ;
  assign n3526 = ~n1758 & ~n2422 ;
  assign n3527 = n1895 & ~n3526 ;
  assign n3528 = ~n1757 & ~n1763 ;
  assign n3529 = ~\sa21_reg[1]/P0001  & \sa21_reg[2]/P0001  ;
  assign n3530 = \sa21_reg[5]/P0001  & n3529 ;
  assign n3531 = ~n3528 & n3530 ;
  assign n3532 = ~n3527 & ~n3531 ;
  assign n3533 = ~n3514 & n3532 ;
  assign n3517 = ~n1802 & ~n1841 ;
  assign n3518 = \sa21_reg[3]/P0001  & n1840 ;
  assign n3519 = ~n3517 & ~n3518 ;
  assign n3515 = n1754 & n2452 ;
  assign n3516 = \sa21_reg[2]/P0001  & n2429 ;
  assign n3520 = ~n3515 & ~n3516 ;
  assign n3521 = ~n3519 & n3520 ;
  assign n3522 = \sa21_reg[1]/P0001  & ~n3521 ;
  assign n3523 = ~\sa21_reg[3]/P0001  & ~n2418 ;
  assign n3524 = ~n3028 & ~n3523 ;
  assign n3525 = ~\sa21_reg[1]/P0001  & ~n3524 ;
  assign n3534 = ~n3522 & ~n3525 ;
  assign n3535 = n3533 & n3534 ;
  assign n3536 = ~\sa21_reg[0]/P0001  & ~n3535 ;
  assign n3573 = ~\sa21_reg[2]/P0001  & ~n2901 ;
  assign n3574 = ~n2451 & n3573 ;
  assign n3575 = ~n3049 & n3574 ;
  assign n3576 = \sa21_reg[2]/P0001  & ~n1891 ;
  assign n3577 = ~n3055 & n3576 ;
  assign n3578 = ~n3575 & ~n3577 ;
  assign n3571 = n1745 & n1877 ;
  assign n3572 = n1753 & n3571 ;
  assign n3579 = ~n2928 & ~n3572 ;
  assign n3580 = ~n3578 & n3579 ;
  assign n3581 = ~\sa21_reg[1]/P0001  & ~n3580 ;
  assign n3568 = n1831 & n1879 ;
  assign n3569 = ~n1821 & ~n3568 ;
  assign n3570 = \sa21_reg[6]/NET0131  & ~n3569 ;
  assign n3582 = ~n1788 & ~n2865 ;
  assign n3583 = \sa21_reg[2]/P0001  & ~n3582 ;
  assign n3584 = n1754 & n1849 ;
  assign n3585 = ~n1883 & ~n3020 ;
  assign n3586 = ~n3584 & n3585 ;
  assign n3587 = ~n3583 & n3586 ;
  assign n3588 = \sa21_reg[1]/P0001  & ~n3587 ;
  assign n3589 = ~n3570 & ~n3588 ;
  assign n3590 = ~n3581 & n3589 ;
  assign n3591 = ~n3536 & n3590 ;
  assign n3592 = ~n3567 & n3591 ;
  assign n3593 = n2529 & ~n3592 ;
  assign n3594 = ~n2529 & n3592 ;
  assign n3595 = ~n3593 & ~n3594 ;
  assign n3613 = n1585 & n1619 ;
  assign n3614 = ~n1609 & ~n3613 ;
  assign n3616 = \sa10_reg[4]/P0001  & ~n1681 ;
  assign n3615 = \sa10_reg[5]/P0001  & ~n1681 ;
  assign n3617 = \sa10_reg[7]/NET0131  & ~n3615 ;
  assign n3618 = ~n3616 & n3617 ;
  assign n3619 = ~n1673 & ~n3618 ;
  assign n3620 = \sa10_reg[2]/P0001  & ~n3619 ;
  assign n3621 = n3614 & ~n3620 ;
  assign n3622 = \sa10_reg[1]/P0001  & ~n3621 ;
  assign n3630 = ~n1700 & ~n2093 ;
  assign n3599 = ~\sa10_reg[3]/P0001  & n2621 ;
  assign n3631 = ~n2119 & ~n3599 ;
  assign n3632 = n3630 & n3631 ;
  assign n3633 = ~\sa10_reg[2]/P0001  & ~n3632 ;
  assign n3624 = n1594 & ~n1652 ;
  assign n3625 = ~n1600 & n3624 ;
  assign n3623 = ~\sa10_reg[6]/NET0131  & n2826 ;
  assign n3626 = ~n2093 & ~n2778 ;
  assign n3627 = ~n3623 & n3626 ;
  assign n3628 = ~n3625 & n3627 ;
  assign n3629 = ~\sa10_reg[1]/P0001  & ~n3628 ;
  assign n3634 = n2565 & ~n2595 ;
  assign n3635 = \sa10_reg[4]/P0001  & n1616 ;
  assign n3636 = ~n3634 & ~n3635 ;
  assign n3637 = ~n3629 & n3636 ;
  assign n3638 = ~n3633 & n3637 ;
  assign n3639 = ~n3622 & n3638 ;
  assign n3640 = \sa10_reg[0]/P0001  & ~n3639 ;
  assign n3600 = ~n2607 & ~n3599 ;
  assign n3601 = \sa10_reg[2]/P0001  & ~n3600 ;
  assign n3596 = ~n1639 & ~n1708 ;
  assign n3597 = ~\sa10_reg[2]/P0001  & ~n3596 ;
  assign n3598 = n1598 & n1636 ;
  assign n3602 = ~n2567 & ~n3598 ;
  assign n3603 = ~n3597 & n3602 ;
  assign n3604 = ~n3601 & n3603 ;
  assign n3605 = ~\sa10_reg[0]/P0001  & ~n3604 ;
  assign n3606 = ~n1628 & ~n2130 ;
  assign n3607 = ~n2581 & n3606 ;
  assign n3608 = ~\sa10_reg[2]/P0001  & ~n3607 ;
  assign n3609 = ~n1631 & ~n2558 ;
  assign n3610 = ~n3608 & n3609 ;
  assign n3611 = ~n3605 & n3610 ;
  assign n3612 = ~\sa10_reg[1]/P0001  & ~n3611 ;
  assign n3641 = ~\sa10_reg[6]/NET0131  & n1590 ;
  assign n3642 = n1634 & ~n3616 ;
  assign n3643 = ~n3641 & ~n3642 ;
  assign n3644 = ~\sa10_reg[2]/P0001  & ~n3643 ;
  assign n3645 = ~n1591 & ~n1684 ;
  assign n3646 = \sa10_reg[2]/P0001  & ~n3645 ;
  assign n3647 = ~n2185 & n2744 ;
  assign n3648 = ~n3646 & n3647 ;
  assign n3649 = ~n3644 & n3648 ;
  assign n3650 = \sa10_reg[1]/P0001  & ~n3649 ;
  assign n3653 = ~n2567 & ~n2748 ;
  assign n3654 = ~\sa10_reg[2]/P0001  & ~n3653 ;
  assign n3651 = ~n1586 & ~n1687 ;
  assign n3652 = n1661 & ~n3651 ;
  assign n3655 = ~n1730 & ~n2807 ;
  assign n3656 = ~n3652 & n3655 ;
  assign n3657 = ~n3654 & n3656 ;
  assign n3658 = ~n3650 & n3657 ;
  assign n3659 = ~\sa10_reg[0]/P0001  & ~n3658 ;
  assign n3660 = n1582 & n1668 ;
  assign n3661 = ~n1587 & ~n2185 ;
  assign n3662 = ~n3660 & n3661 ;
  assign n3663 = ~n1602 & ~n1616 ;
  assign n3664 = n3662 & n3663 ;
  assign n3665 = \sa10_reg[1]/P0001  & ~n3664 ;
  assign n3666 = ~\sa10_reg[2]/P0001  & ~n3665 ;
  assign n3667 = ~\sa10_reg[5]/P0001  & n3641 ;
  assign n3668 = ~\sa10_reg[1]/P0001  & ~n1730 ;
  assign n3669 = ~n1592 & n3668 ;
  assign n3670 = ~n3667 & n3669 ;
  assign n3671 = ~n1609 & ~n2546 ;
  assign n3672 = \sa10_reg[3]/P0001  & ~n3671 ;
  assign n3673 = ~n1674 & n1697 ;
  assign n3674 = ~n3672 & n3673 ;
  assign n3675 = ~n3670 & ~n3674 ;
  assign n3676 = ~n2558 & ~n2819 ;
  assign n3677 = ~n3675 & n3676 ;
  assign n3678 = ~n3666 & ~n3677 ;
  assign n3679 = ~n3659 & ~n3678 ;
  assign n3680 = ~n3612 & n3679 ;
  assign n3681 = ~n3640 & n3680 ;
  assign n3699 = ~n1483 & ~n1566 ;
  assign n3700 = ~\sa03_reg[2]/P0001  & ~n3699 ;
  assign n3701 = ~n1552 & ~n2685 ;
  assign n3702 = ~n3700 & n3701 ;
  assign n3703 = ~\sa03_reg[1]/P0001  & ~n3702 ;
  assign n3692 = \sa03_reg[7]/NET0131  & n1408 ;
  assign n3693 = ~n1455 & ~n2248 ;
  assign n3694 = ~n3692 & n3693 ;
  assign n3695 = ~\sa03_reg[2]/P0001  & ~n3694 ;
  assign n3696 = ~n1325 & n1448 ;
  assign n3697 = ~n3695 & n3696 ;
  assign n3698 = \sa03_reg[1]/P0001  & ~n3697 ;
  assign n3690 = ~n1383 & ~n1460 ;
  assign n3691 = n1436 & ~n3690 ;
  assign n3686 = \sa03_reg[1]/P0001  & \sa03_reg[2]/P0001  ;
  assign n3687 = n1327 & n1342 ;
  assign n3688 = ~n1375 & ~n3687 ;
  assign n3689 = n3686 & ~n3688 ;
  assign n3704 = ~n1409 & ~n1415 ;
  assign n3705 = ~n3689 & n3704 ;
  assign n3706 = ~n3691 & n3705 ;
  assign n3682 = ~n1462 & ~n2685 ;
  assign n3683 = ~\sa03_reg[2]/P0001  & ~n3682 ;
  assign n3684 = ~n1537 & ~n2289 ;
  assign n3685 = n1494 & ~n3684 ;
  assign n3707 = ~n3683 & ~n3685 ;
  assign n3708 = n3706 & n3707 ;
  assign n3709 = ~n3698 & n3708 ;
  assign n3710 = ~n3703 & n3709 ;
  assign n3711 = ~\sa03_reg[0]/P0001  & ~n3710 ;
  assign n3712 = n1316 & n1353 ;
  assign n3713 = ~n1369 & ~n3712 ;
  assign n3714 = \sa03_reg[3]/P0001  & n2684 ;
  assign n3715 = ~n1396 & ~n2264 ;
  assign n3716 = ~n3714 & n3715 ;
  assign n3717 = \sa03_reg[2]/P0001  & ~n3716 ;
  assign n3718 = n3713 & ~n3717 ;
  assign n3719 = \sa03_reg[1]/P0001  & ~n3718 ;
  assign n3731 = ~n1414 & ~n1565 ;
  assign n3732 = ~n2289 & n3731 ;
  assign n3733 = ~\sa03_reg[2]/P0001  & ~n3732 ;
  assign n3720 = n1316 & ~n2684 ;
  assign n3721 = ~n1376 & n3720 ;
  assign n3722 = n1332 & n1429 ;
  assign n3723 = ~n3721 & ~n3722 ;
  assign n3724 = ~\sa03_reg[1]/P0001  & ~n3723 ;
  assign n3726 = ~\sa03_reg[3]/P0001  & n1329 ;
  assign n3727 = ~\sa03_reg[1]/P0001  & n1330 ;
  assign n3728 = ~n1341 & ~n3727 ;
  assign n3729 = n3726 & ~n3728 ;
  assign n3725 = n1328 & ~n1515 ;
  assign n3730 = n2200 & ~n3686 ;
  assign n3734 = ~n3725 & ~n3730 ;
  assign n3735 = ~n3729 & n3734 ;
  assign n3736 = ~n3724 & n3735 ;
  assign n3737 = ~n3733 & n3736 ;
  assign n3738 = ~n3719 & n3737 ;
  assign n3739 = \sa03_reg[0]/P0001  & ~n3738 ;
  assign n3740 = ~n1359 & ~n1409 ;
  assign n3741 = ~n1438 & n3740 ;
  assign n3742 = \sa03_reg[2]/P0001  & ~n3741 ;
  assign n3743 = ~n1459 & ~n2679 ;
  assign n3744 = ~n3742 & n3743 ;
  assign n3745 = ~\sa03_reg[1]/P0001  & ~n3744 ;
  assign n3757 = ~n1369 & ~n2260 ;
  assign n3758 = \sa03_reg[3]/P0001  & ~n3757 ;
  assign n3759 = ~n1526 & ~n3758 ;
  assign n3760 = n3686 & ~n3759 ;
  assign n3746 = ~n1334 & n1355 ;
  assign n3747 = ~n3726 & ~n3746 ;
  assign n3748 = ~\sa03_reg[7]/NET0131  & ~n3747 ;
  assign n3749 = ~\sa03_reg[4]/P0001  & n3726 ;
  assign n3750 = ~n1497 & ~n3749 ;
  assign n3751 = ~n3748 & n3750 ;
  assign n3752 = n1558 & ~n3751 ;
  assign n3753 = ~\sa03_reg[1]/P0001  & ~\sa03_reg[2]/P0001  ;
  assign n3754 = ~n1480 & ~n2219 ;
  assign n3755 = ~n1461 & n3754 ;
  assign n3756 = n3753 & ~n3755 ;
  assign n3761 = n1384 & n2229 ;
  assign n3762 = ~n2235 & ~n3761 ;
  assign n3763 = ~n3756 & n3762 ;
  assign n3764 = ~n3752 & n3763 ;
  assign n3765 = ~n3760 & n3764 ;
  assign n3766 = ~n3745 & n3765 ;
  assign n3767 = ~n3739 & n3766 ;
  assign n3768 = ~n3711 & n3767 ;
  assign n3769 = ~n3681 & ~n3768 ;
  assign n3770 = n3681 & n3768 ;
  assign n3771 = ~n3769 & ~n3770 ;
  assign n3772 = n3595 & n3771 ;
  assign n3773 = ~n3595 & ~n3771 ;
  assign n3774 = ~n3772 & ~n3773 ;
  assign n3776 = n3509 & n3774 ;
  assign n3775 = ~n3509 & ~n3774 ;
  assign n3777 = ~\ld_r_reg/P0001  & ~n3775 ;
  assign n3778 = ~n3776 & n3777 ;
  assign n3780 = \text_in_r_reg[9]/P0001  & \u0_w_reg[3][9]/P0001  ;
  assign n3779 = ~\text_in_r_reg[9]/P0001  & ~\u0_w_reg[3][9]/P0001  ;
  assign n3781 = \ld_r_reg/P0001  & ~n3779 ;
  assign n3782 = ~n3780 & n3781 ;
  assign n3783 = ~n3778 & ~n3782 ;
  assign n3784 = ~n2736 & ~n2963 ;
  assign n3785 = n2736 & n2963 ;
  assign n3786 = ~n3784 & ~n3785 ;
  assign n3787 = \u0_w_reg[3][5]/P0001  & ~n3205 ;
  assign n3788 = ~\u0_w_reg[3][5]/P0001  & n3205 ;
  assign n3789 = ~n3787 & ~n3788 ;
  assign n3790 = n2939 & n3789 ;
  assign n3791 = ~n2939 & ~n3789 ;
  assign n3792 = ~n3790 & ~n3791 ;
  assign n3794 = n3786 & n3792 ;
  assign n3793 = ~n3786 & ~n3792 ;
  assign n3795 = ~\ld_r_reg/P0001  & ~n3793 ;
  assign n3796 = ~n3794 & n3795 ;
  assign n3798 = \text_in_r_reg[5]/P0001  & \u0_w_reg[3][5]/P0001  ;
  assign n3797 = ~\text_in_r_reg[5]/P0001  & ~\u0_w_reg[3][5]/P0001  ;
  assign n3799 = \ld_r_reg/P0001  & ~n3797 ;
  assign n3800 = ~n3798 & n3799 ;
  assign n3801 = ~n3796 & ~n3800 ;
  assign n3802 = \u0_w_reg[3][28]/P0001  & ~n3205 ;
  assign n3803 = ~\u0_w_reg[3][28]/P0001  & n3205 ;
  assign n3804 = ~n3802 & ~n3803 ;
  assign n3805 = n3072 & n3804 ;
  assign n3806 = ~n3072 & ~n3804 ;
  assign n3807 = ~n3805 & ~n3806 ;
  assign n3818 = ~n1329 & ~n1398 ;
  assign n3819 = ~\sa03_reg[7]/NET0131  & n3818 ;
  assign n3820 = ~\sa03_reg[2]/P0001  & ~n3819 ;
  assign n3822 = \sa03_reg[2]/P0001  & ~n2710 ;
  assign n3821 = \sa03_reg[4]/P0001  & n1367 ;
  assign n3823 = ~n3726 & ~n3821 ;
  assign n3824 = n3822 & n3823 ;
  assign n3825 = ~n3820 & ~n3824 ;
  assign n3826 = ~n1537 & ~n2293 ;
  assign n3827 = ~n1365 & n3826 ;
  assign n3828 = ~n3825 & n3827 ;
  assign n3829 = \sa03_reg[1]/P0001  & ~n3828 ;
  assign n3810 = \sa03_reg[2]/P0001  & n1450 ;
  assign n3813 = ~n2679 & ~n2715 ;
  assign n3814 = ~n3810 & n3813 ;
  assign n3808 = ~n1328 & ~n2219 ;
  assign n3809 = ~\sa03_reg[2]/P0001  & ~n3808 ;
  assign n3811 = ~n1409 & ~n1571 ;
  assign n3812 = ~n1496 & n3811 ;
  assign n3815 = ~n3809 & n3812 ;
  assign n3816 = n3814 & n3815 ;
  assign n3817 = ~\sa03_reg[1]/P0001  & ~n3816 ;
  assign n3830 = ~\sa03_reg[3]/P0001  & n1330 ;
  assign n3831 = ~\sa03_reg[5]/P0001  & n3830 ;
  assign n3832 = \sa03_reg[6]/NET0131  & n1340 ;
  assign n3833 = ~n1462 & ~n3832 ;
  assign n3834 = ~n3831 & n3833 ;
  assign n3835 = ~\sa03_reg[2]/P0001  & ~n3834 ;
  assign n3836 = ~n1333 & n1405 ;
  assign n3837 = \sa03_reg[2]/P0001  & \sa03_reg[4]/P0001  ;
  assign n3838 = ~n3836 & n3837 ;
  assign n3839 = ~n1469 & ~n3838 ;
  assign n3840 = ~n3835 & n3839 ;
  assign n3841 = ~n3817 & n3840 ;
  assign n3842 = ~n3829 & n3841 ;
  assign n3843 = \sa03_reg[0]/P0001  & ~n3842 ;
  assign n3862 = ~n1377 & ~n1421 ;
  assign n3863 = \sa03_reg[2]/P0001  & ~n3862 ;
  assign n3865 = \sa03_reg[1]/P0001  & ~n2665 ;
  assign n3866 = ~n1354 & n3865 ;
  assign n3864 = ~\sa03_reg[2]/P0001  & n1331 ;
  assign n3867 = ~n3712 & ~n3864 ;
  assign n3868 = n3866 & n3867 ;
  assign n3869 = ~n3863 & n3868 ;
  assign n3873 = ~\sa03_reg[1]/P0001  & ~n3831 ;
  assign n3870 = n1341 & ~n1385 ;
  assign n3871 = \sa03_reg[2]/P0001  & ~n1355 ;
  assign n3872 = n1327 & n3871 ;
  assign n3874 = ~n3870 & ~n3872 ;
  assign n3875 = n3873 & n3874 ;
  assign n3876 = ~n1560 & n3875 ;
  assign n3877 = ~n3869 & ~n3876 ;
  assign n3858 = ~\sa03_reg[2]/P0001  & n1489 ;
  assign n3859 = n1324 & n1383 ;
  assign n3860 = n1562 & ~n3859 ;
  assign n3861 = ~n3858 & ~n3860 ;
  assign n3878 = ~n1443 & ~n3861 ;
  assign n3879 = ~n3877 & n3878 ;
  assign n3880 = ~\sa03_reg[0]/P0001  & ~n3879 ;
  assign n3846 = ~n1319 & ~n1331 ;
  assign n3847 = ~n1533 & n3846 ;
  assign n3848 = n2225 & ~n3847 ;
  assign n3845 = ~\sa03_reg[2]/P0001  & n2693 ;
  assign n3849 = ~n2658 & ~n3845 ;
  assign n3850 = ~n3848 & n3849 ;
  assign n3851 = \sa03_reg[1]/P0001  & ~n3850 ;
  assign n3855 = ~n1443 & ~n1461 ;
  assign n3856 = n1494 & ~n3855 ;
  assign n3852 = \sa03_reg[6]/NET0131  & n1454 ;
  assign n3853 = ~n1537 & ~n3852 ;
  assign n3854 = n3686 & ~n3853 ;
  assign n3881 = ~n1552 & ~n3761 ;
  assign n3844 = n1369 & n1374 ;
  assign n3857 = n2655 & n3753 ;
  assign n3882 = ~n3844 & ~n3857 ;
  assign n3883 = n3881 & n3882 ;
  assign n3884 = ~n3854 & n3883 ;
  assign n3885 = ~n3856 & n3884 ;
  assign n3886 = ~n3851 & n3885 ;
  assign n3887 = ~n3880 & n3886 ;
  assign n3888 = ~n3843 & n3887 ;
  assign n3947 = n2131 & ~n2565 ;
  assign n3948 = ~n2621 & ~n2740 ;
  assign n3949 = n2602 & n3948 ;
  assign n3950 = ~n3947 & ~n3949 ;
  assign n3951 = ~n1711 & ~n1730 ;
  assign n3952 = ~n2558 & n3951 ;
  assign n3953 = ~n3950 & n3952 ;
  assign n3954 = ~\sa10_reg[1]/P0001  & ~n3953 ;
  assign n3931 = n1582 & ~n2162 ;
  assign n3932 = ~n2623 & ~n3931 ;
  assign n3933 = \sa10_reg[2]/P0001  & ~n3932 ;
  assign n3930 = n1626 & n3616 ;
  assign n3934 = ~n2147 & ~n2607 ;
  assign n3935 = ~n1688 & n3934 ;
  assign n3936 = ~n3930 & n3935 ;
  assign n3937 = ~n3933 & n3936 ;
  assign n3938 = \sa10_reg[1]/P0001  & ~n3937 ;
  assign n3902 = n1608 & n1668 ;
  assign n3939 = \sa10_reg[6]/NET0131  & n2593 ;
  assign n3940 = ~n2748 & ~n3939 ;
  assign n3941 = ~n3902 & n3940 ;
  assign n3942 = ~\sa10_reg[2]/P0001  & ~n3941 ;
  assign n3943 = \sa10_reg[2]/P0001  & \sa10_reg[4]/P0001  ;
  assign n3944 = \sa10_reg[3]/P0001  & n1597 ;
  assign n3945 = ~n2811 & ~n3944 ;
  assign n3946 = n3943 & ~n3945 ;
  assign n3955 = ~n2758 & ~n3946 ;
  assign n3956 = ~n3942 & n3955 ;
  assign n3957 = ~n3938 & n3956 ;
  assign n3958 = ~n3954 & n3957 ;
  assign n3959 = \sa10_reg[0]/P0001  & ~n3958 ;
  assign n3899 = n1590 & ~n1650 ;
  assign n3900 = ~n1703 & ~n3899 ;
  assign n3901 = \sa10_reg[2]/P0001  & ~n3900 ;
  assign n3903 = ~n1704 & ~n3902 ;
  assign n3904 = ~n1725 & n3903 ;
  assign n3905 = ~n3901 & n3904 ;
  assign n3906 = ~\sa10_reg[1]/P0001  & ~n3905 ;
  assign n3889 = ~n1601 & ~n1657 ;
  assign n3890 = \sa10_reg[2]/P0001  & ~n3889 ;
  assign n3892 = ~n1599 & ~n2550 ;
  assign n3891 = n1582 & n2109 ;
  assign n3893 = ~n3613 & ~n3891 ;
  assign n3894 = n3892 & n3893 ;
  assign n3895 = ~n3890 & n3894 ;
  assign n3896 = \sa10_reg[1]/P0001  & ~n3895 ;
  assign n3898 = ~\sa10_reg[2]/P0001  & ~n1596 ;
  assign n3897 = n1601 & n1664 ;
  assign n3907 = ~n1714 & ~n2755 ;
  assign n3908 = ~n3897 & n3907 ;
  assign n3909 = ~n3898 & n3908 ;
  assign n3910 = ~n3896 & n3909 ;
  assign n3911 = ~n3906 & n3910 ;
  assign n3912 = ~\sa10_reg[0]/P0001  & ~n3911 ;
  assign n3919 = ~n1638 & ~n2098 ;
  assign n3920 = ~n2582 & n3919 ;
  assign n3921 = n1633 & ~n3920 ;
  assign n3922 = \sa10_reg[3]/P0001  & n1650 ;
  assign n3923 = n2109 & n3922 ;
  assign n3924 = ~n2594 & ~n3923 ;
  assign n3925 = ~n3921 & n3924 ;
  assign n3926 = \sa10_reg[1]/P0001  & ~n3925 ;
  assign n3914 = \sa10_reg[6]/NET0131  & n1726 ;
  assign n3915 = ~n2607 & ~n3914 ;
  assign n3916 = \sa10_reg[1]/P0001  & ~n3915 ;
  assign n3917 = ~n2558 & ~n3916 ;
  assign n3918 = \sa10_reg[2]/P0001  & ~n3917 ;
  assign n3927 = ~n2581 & ~n2755 ;
  assign n3928 = n2183 & ~n3927 ;
  assign n3929 = n2566 & n2825 ;
  assign n3913 = n1609 & n1664 ;
  assign n3960 = ~n3598 & ~n3913 ;
  assign n3961 = ~n3929 & n3960 ;
  assign n3962 = ~n3928 & n3961 ;
  assign n3963 = ~n3918 & n3962 ;
  assign n3964 = ~n3926 & n3963 ;
  assign n3965 = ~n3912 & n3964 ;
  assign n3966 = ~n3959 & n3965 ;
  assign n3967 = n3888 & ~n3966 ;
  assign n3968 = ~n3888 & n3966 ;
  assign n3969 = ~n3967 & ~n3968 ;
  assign n3970 = ~n2307 & n3969 ;
  assign n3971 = n2307 & ~n3969 ;
  assign n3972 = ~n3970 & ~n3971 ;
  assign n3974 = ~n3807 & n3972 ;
  assign n3973 = n3807 & ~n3972 ;
  assign n3975 = ~\ld_r_reg/P0001  & ~n3973 ;
  assign n3976 = ~n3974 & n3975 ;
  assign n3978 = ~\text_in_r_reg[28]/P0001  & \u0_w_reg[3][28]/P0001  ;
  assign n3977 = \text_in_r_reg[28]/P0001  & ~\u0_w_reg[3][28]/P0001  ;
  assign n3979 = \ld_r_reg/P0001  & ~n3977 ;
  assign n3980 = ~n3978 & n3979 ;
  assign n3981 = ~n3976 & ~n3980 ;
  assign n4033 = n1772 & ~n1854 ;
  assign n4034 = ~n2490 & ~n4033 ;
  assign n4035 = \sa21_reg[2]/P0001  & ~n4034 ;
  assign n4032 = n1832 & n2448 ;
  assign n4037 = ~n2508 & ~n3040 ;
  assign n4038 = ~n4032 & n4037 ;
  assign n4036 = \sa21_reg[1]/P0001  & ~n2446 ;
  assign n4039 = ~n1792 & n4036 ;
  assign n4040 = n4038 & n4039 ;
  assign n4041 = ~n4035 & n4040 ;
  assign n4046 = ~\sa21_reg[1]/P0001  & ~n1865 ;
  assign n4047 = ~n1891 & n4046 ;
  assign n4048 = ~n2997 & n4047 ;
  assign n4042 = ~n2513 & ~n2838 ;
  assign n4043 = ~\sa21_reg[2]/P0001  & ~n4042 ;
  assign n4044 = ~n1788 & ~n1879 ;
  assign n4045 = ~n2479 & ~n4044 ;
  assign n4049 = ~n4043 & ~n4045 ;
  assign n4050 = n4048 & n4049 ;
  assign n4051 = ~n4041 & ~n4050 ;
  assign n3994 = ~\sa21_reg[5]/P0001  & n1816 ;
  assign n4028 = n3511 & ~n3994 ;
  assign n4029 = ~\sa21_reg[2]/P0001  & ~n4028 ;
  assign n4030 = ~n2842 & n2919 ;
  assign n4031 = n2917 & ~n4030 ;
  assign n4052 = ~n2906 & ~n4031 ;
  assign n4053 = ~n4029 & n4052 ;
  assign n4054 = ~n4051 & n4053 ;
  assign n4055 = \sa21_reg[0]/P0001  & ~n4054 ;
  assign n3984 = ~n1785 & ~n1839 ;
  assign n3985 = \sa21_reg[2]/P0001  & ~n3984 ;
  assign n3986 = \sa21_reg[1]/P0001  & ~n1788 ;
  assign n3987 = ~n2853 & n3986 ;
  assign n3982 = n1781 & n1802 ;
  assign n3983 = n1764 & n2479 ;
  assign n3988 = ~n3982 & ~n3983 ;
  assign n3989 = n3987 & n3988 ;
  assign n3990 = ~n3985 & n3989 ;
  assign n3995 = ~\sa21_reg[1]/P0001  & ~n1864 ;
  assign n3996 = ~n3994 & n3995 ;
  assign n3991 = n1757 & ~n1832 ;
  assign n3992 = ~n2492 & ~n3991 ;
  assign n3993 = \sa21_reg[2]/P0001  & ~n3992 ;
  assign n3997 = ~n1878 & ~n3993 ;
  assign n3998 = n3996 & n3997 ;
  assign n3999 = ~n3990 & ~n3998 ;
  assign n4000 = ~\sa21_reg[2]/P0001  & ~n1783 ;
  assign n4001 = ~n1890 & ~n1895 ;
  assign n4002 = n1784 & ~n4001 ;
  assign n4003 = ~n1893 & ~n4002 ;
  assign n4004 = ~n4000 & n4003 ;
  assign n4005 = ~n3999 & n4004 ;
  assign n4006 = ~\sa21_reg[0]/P0001  & ~n4005 ;
  assign n4011 = \sa21_reg[6]/NET0131  & n1867 ;
  assign n4012 = ~n1792 & ~n4011 ;
  assign n4013 = \sa21_reg[2]/P0001  & ~n4012 ;
  assign n4008 = ~n1775 & ~n1844 ;
  assign n4009 = ~n1765 & n4008 ;
  assign n4010 = n1754 & ~n4009 ;
  assign n4014 = n1877 & n2993 ;
  assign n4007 = \sa21_reg[2]/P0001  & n3040 ;
  assign n4015 = \sa21_reg[1]/P0001  & ~n4007 ;
  assign n4016 = ~n4014 & n4015 ;
  assign n4017 = ~n4010 & n4016 ;
  assign n4018 = ~n4013 & n4017 ;
  assign n4021 = ~n1864 & ~n2417 ;
  assign n4022 = n1831 & ~n4021 ;
  assign n4019 = \sa21_reg[3]/P0001  & n1822 ;
  assign n4020 = n2479 & n4019 ;
  assign n4023 = ~\sa21_reg[1]/P0001  & ~n4020 ;
  assign n4024 = ~n4022 & n4023 ;
  assign n4025 = ~n4018 & ~n4024 ;
  assign n4026 = ~n1794 & ~n2426 ;
  assign n4027 = n1894 & ~n4026 ;
  assign n4056 = ~n1874 & ~n4027 ;
  assign n4057 = ~n4025 & n4056 ;
  assign n4058 = ~n4006 & n4057 ;
  assign n4059 = ~n4055 & n4058 ;
  assign n4060 = n3966 & ~n4059 ;
  assign n4061 = ~n3966 & n4059 ;
  assign n4062 = ~n4060 & ~n4061 ;
  assign n4063 = n2199 & ~n2736 ;
  assign n4064 = ~n2199 & n2736 ;
  assign n4065 = ~n4063 & ~n4064 ;
  assign n4066 = n4062 & n4065 ;
  assign n4067 = ~n4062 & ~n4065 ;
  assign n4068 = ~n4066 & ~n4067 ;
  assign n4069 = ~\u0_w_reg[3][20]/P0001  & ~n3205 ;
  assign n4070 = \u0_w_reg[3][20]/P0001  & n3205 ;
  assign n4071 = ~n4069 & ~n4070 ;
  assign n4072 = n2529 & ~n3069 ;
  assign n4073 = ~n2529 & n3069 ;
  assign n4074 = ~n4072 & ~n4073 ;
  assign n4075 = n4071 & n4074 ;
  assign n4076 = ~n4071 & ~n4074 ;
  assign n4077 = ~n4075 & ~n4076 ;
  assign n4079 = ~n4068 & n4077 ;
  assign n4078 = n4068 & ~n4077 ;
  assign n4080 = ~\ld_r_reg/P0001  & ~n4078 ;
  assign n4081 = ~n4079 & n4080 ;
  assign n4083 = ~\text_in_r_reg[20]/P0001  & \u0_w_reg[3][20]/P0001  ;
  assign n4082 = \text_in_r_reg[20]/P0001  & ~\u0_w_reg[3][20]/P0001  ;
  assign n4084 = \ld_r_reg/P0001  & ~n4082 ;
  assign n4085 = ~n4083 & n4084 ;
  assign n4086 = ~n4081 & ~n4085 ;
  assign n4103 = ~n1343 & ~n1556 ;
  assign n4104 = ~n1397 & n4103 ;
  assign n4105 = \sa03_reg[2]/P0001  & ~n4104 ;
  assign n4100 = n2206 & n2225 ;
  assign n4101 = n1423 & ~n2226 ;
  assign n4102 = n1352 & n1449 ;
  assign n4106 = ~n4101 & ~n4102 ;
  assign n4107 = ~n4100 & n4106 ;
  assign n4108 = ~n4105 & n4107 ;
  assign n4109 = ~\sa03_reg[1]/P0001  & ~n4108 ;
  assign n4090 = ~n1326 & ~n1383 ;
  assign n4091 = \sa03_reg[3]/P0001  & ~n4090 ;
  assign n4092 = ~n2236 & ~n2279 ;
  assign n4093 = ~n4091 & n4092 ;
  assign n4094 = ~\sa03_reg[2]/P0001  & ~n4093 ;
  assign n4087 = ~n1462 & ~n2712 ;
  assign n4088 = n1481 & n4087 ;
  assign n4089 = \sa03_reg[2]/P0001  & ~n4088 ;
  assign n4095 = ~n1326 & ~n1329 ;
  assign n4096 = ~\sa03_reg[2]/P0001  & ~n1332 ;
  assign n4097 = n4095 & n4096 ;
  assign n4098 = ~n1566 & ~n4097 ;
  assign n4099 = \sa03_reg[1]/P0001  & ~n4098 ;
  assign n4110 = ~n2289 & ~n2693 ;
  assign n4111 = ~n4099 & n4110 ;
  assign n4112 = ~n4089 & n4111 ;
  assign n4113 = ~n4094 & n4112 ;
  assign n4114 = ~n4109 & n4113 ;
  assign n4115 = \sa03_reg[0]/P0001  & ~n4114 ;
  assign n4116 = ~n1541 & n3833 ;
  assign n4117 = ~\sa03_reg[2]/P0001  & ~n4116 ;
  assign n4118 = \sa03_reg[5]/P0001  & ~n1323 ;
  assign n4119 = n1423 & n3871 ;
  assign n4120 = ~n4118 & n4119 ;
  assign n4121 = n1339 & ~n1398 ;
  assign n4122 = n1494 & n4121 ;
  assign n4132 = ~n4120 & ~n4122 ;
  assign n4133 = ~n4117 & n4132 ;
  assign n4123 = ~\sa03_reg[3]/P0001  & ~n2201 ;
  assign n4124 = ~n2657 & ~n4123 ;
  assign n4125 = ~\sa03_reg[1]/P0001  & ~n4124 ;
  assign n4128 = \sa03_reg[3]/P0001  & n2715 ;
  assign n4126 = ~n1316 & ~n1323 ;
  assign n4127 = ~n3720 & ~n4126 ;
  assign n4129 = ~n2250 & ~n4127 ;
  assign n4130 = ~n4128 & n4129 ;
  assign n4131 = \sa03_reg[1]/P0001  & ~n4130 ;
  assign n4134 = ~n4125 & ~n4131 ;
  assign n4135 = n4133 & n4134 ;
  assign n4136 = ~\sa03_reg[0]/P0001  & ~n4135 ;
  assign n4141 = ~n1380 & ~n1416 ;
  assign n4142 = ~n1482 & n4141 ;
  assign n4143 = n2225 & ~n4142 ;
  assign n4140 = n1446 & n1515 ;
  assign n4137 = \sa03_reg[2]/P0001  & n1352 ;
  assign n4138 = ~n1376 & n4137 ;
  assign n4139 = n4095 & n4138 ;
  assign n4144 = ~n1415 & ~n4139 ;
  assign n4145 = ~n4140 & n4144 ;
  assign n4146 = ~n4143 & n4145 ;
  assign n4147 = ~\sa03_reg[1]/P0001  & ~n4146 ;
  assign n4150 = n1436 & n1566 ;
  assign n4152 = ~n1417 & ~n1496 ;
  assign n4151 = ~\sa03_reg[2]/P0001  & n2293 ;
  assign n4153 = ~n2670 & ~n4151 ;
  assign n4154 = n4152 & n4153 ;
  assign n4155 = ~n4150 & n4154 ;
  assign n4156 = \sa03_reg[1]/P0001  & ~n4155 ;
  assign n4148 = n1435 & n4137 ;
  assign n4149 = \sa03_reg[6]/NET0131  & n1523 ;
  assign n4157 = ~n4148 & ~n4149 ;
  assign n4158 = ~n4156 & n4157 ;
  assign n4159 = ~n4147 & n4158 ;
  assign n4160 = ~n4136 & n4159 ;
  assign n4161 = ~n4115 & n4160 ;
  assign n4162 = ~n2304 & ~n4161 ;
  assign n4163 = n2304 & n4161 ;
  assign n4164 = ~n4162 & ~n4163 ;
  assign n4165 = n3771 & ~n4164 ;
  assign n4166 = ~n3771 & n4164 ;
  assign n4167 = ~n4165 & ~n4166 ;
  assign n4205 = ~n1784 & n3518 ;
  assign n4206 = n1772 & n1816 ;
  assign n4204 = ~\sa21_reg[2]/P0001  & n2842 ;
  assign n4207 = ~n2417 & ~n4204 ;
  assign n4208 = ~n4206 & n4207 ;
  assign n4209 = ~n4205 & n4208 ;
  assign n4210 = ~\sa21_reg[1]/P0001  & ~n4209 ;
  assign n4196 = ~n1794 & ~n3982 ;
  assign n4198 = ~\sa21_reg[5]/P0001  & n1793 ;
  assign n4197 = \sa21_reg[4]/P0001  & n1758 ;
  assign n4199 = ~n4019 & ~n4197 ;
  assign n4200 = ~n4198 & n4199 ;
  assign n4201 = \sa21_reg[2]/P0001  & ~n4200 ;
  assign n4202 = n4196 & ~n4201 ;
  assign n4203 = \sa21_reg[1]/P0001  & ~n4202 ;
  assign n4213 = ~n1838 & ~n2417 ;
  assign n4214 = ~n1885 & n4213 ;
  assign n4215 = ~\sa21_reg[2]/P0001  & ~n4214 ;
  assign n4211 = n1823 & n3026 ;
  assign n4212 = ~n1894 & n2493 ;
  assign n4216 = ~n4211 & ~n4212 ;
  assign n4217 = ~n4215 & n4216 ;
  assign n4218 = ~n4203 & n4217 ;
  assign n4219 = ~n4210 & n4218 ;
  assign n4220 = \sa21_reg[0]/P0001  & ~n4219 ;
  assign n4174 = ~n1760 & ~n1884 ;
  assign n4175 = ~\sa21_reg[2]/P0001  & ~n4174 ;
  assign n4177 = ~\sa21_reg[1]/P0001  & ~n1874 ;
  assign n4176 = \sa21_reg[2]/P0001  & n1838 ;
  assign n4178 = ~n3050 & ~n4007 ;
  assign n4179 = ~n4176 & n4178 ;
  assign n4180 = n4177 & n4179 ;
  assign n4181 = ~n4175 & n4180 ;
  assign n4182 = ~\sa21_reg[2]/P0001  & ~n1833 ;
  assign n4183 = ~n1873 & ~n3542 ;
  assign n4184 = n4182 & n4183 ;
  assign n4185 = ~\sa21_reg[3]/P0001  & n1781 ;
  assign n4186 = \sa21_reg[2]/P0001  & ~n1849 ;
  assign n4187 = ~n4185 & n4186 ;
  assign n4188 = ~n4184 & ~n4187 ;
  assign n4189 = \sa21_reg[1]/P0001  & ~n2502 ;
  assign n4190 = n2877 & n4189 ;
  assign n4191 = ~n4188 & n4190 ;
  assign n4192 = ~n4181 & ~n4191 ;
  assign n4168 = \sa21_reg[2]/P0001  & ~n1872 ;
  assign n4169 = ~n3048 & n4168 ;
  assign n4170 = ~\sa21_reg[2]/P0001  & ~n1865 ;
  assign n4171 = ~n2893 & n4170 ;
  assign n4172 = ~n3050 & n4171 ;
  assign n4173 = ~n4169 & ~n4172 ;
  assign n4193 = ~n2928 & ~n4173 ;
  assign n4194 = ~n4192 & n4193 ;
  assign n4195 = ~\sa21_reg[0]/P0001  & ~n4194 ;
  assign n4237 = ~n1751 & ~n2513 ;
  assign n4238 = ~n2894 & n4237 ;
  assign n4239 = ~\sa21_reg[2]/P0001  & ~n4238 ;
  assign n4240 = ~n1748 & ~n3056 ;
  assign n4241 = ~n4239 & n4240 ;
  assign n4242 = ~\sa21_reg[1]/P0001  & ~n4241 ;
  assign n4221 = ~n1794 & ~n1853 ;
  assign n4222 = \sa21_reg[3]/P0001  & ~n4221 ;
  assign n4223 = ~n1824 & ~n4222 ;
  assign n4224 = n1863 & ~n4223 ;
  assign n4225 = ~n1786 & ~n2426 ;
  assign n4226 = n1894 & ~n4225 ;
  assign n4243 = ~n4224 & ~n4226 ;
  assign n4227 = n1772 & n1815 ;
  assign n4228 = ~n1800 & ~n2502 ;
  assign n4229 = ~n4227 & n4228 ;
  assign n4230 = ~n1776 & ~n1786 ;
  assign n4231 = n4229 & n4230 ;
  assign n4232 = \sa21_reg[1]/P0001  & ~\sa21_reg[2]/P0001  ;
  assign n4233 = ~n4231 & n4232 ;
  assign n4234 = ~n1782 & ~n1865 ;
  assign n4235 = ~n3543 & n4234 ;
  assign n4236 = n3529 & ~n4235 ;
  assign n4244 = ~n4233 & ~n4236 ;
  assign n4245 = n4243 & n4244 ;
  assign n4246 = ~n4242 & n4245 ;
  assign n4247 = ~n4195 & n4246 ;
  assign n4248 = ~n4220 & n4247 ;
  assign n4249 = \u0_w_reg[3][1]/P0001  & ~n4248 ;
  assign n4250 = ~\u0_w_reg[3][1]/P0001  & n4248 ;
  assign n4251 = ~n4249 & ~n4250 ;
  assign n4252 = n3419 & n4251 ;
  assign n4253 = ~n3419 & ~n4251 ;
  assign n4254 = ~n4252 & ~n4253 ;
  assign n4256 = n4167 & n4254 ;
  assign n4255 = ~n4167 & ~n4254 ;
  assign n4257 = ~\ld_r_reg/P0001  & ~n4255 ;
  assign n4258 = ~n4256 & n4257 ;
  assign n4260 = \text_in_r_reg[1]/P0001  & \u0_w_reg[3][1]/P0001  ;
  assign n4259 = ~\text_in_r_reg[1]/P0001  & ~\u0_w_reg[3][1]/P0001  ;
  assign n4261 = \ld_r_reg/P0001  & ~n4259 ;
  assign n4262 = ~n4260 & n4261 ;
  assign n4263 = ~n4258 & ~n4262 ;
  assign n4293 = n1910 & n1919 ;
  assign n4294 = ~n2399 & ~n4293 ;
  assign n4295 = \sa32_reg[2]/P0001  & ~n4294 ;
  assign n4292 = ~\sa32_reg[2]/P0001  & n1994 ;
  assign n4296 = \sa32_reg[1]/P0001  & ~n1925 ;
  assign n4297 = ~n3450 & n4296 ;
  assign n4298 = ~n4292 & n4297 ;
  assign n4299 = ~n2013 & n4298 ;
  assign n4300 = ~n4295 & n4299 ;
  assign n4301 = n1913 & n2046 ;
  assign n4304 = ~\sa32_reg[1]/P0001  & ~n4301 ;
  assign n4305 = ~n3338 & n4304 ;
  assign n4302 = \sa32_reg[7]/P0001  & ~n1990 ;
  assign n4303 = n2397 & n4302 ;
  assign n4306 = ~n3367 & ~n4303 ;
  assign n4307 = n4305 & n4306 ;
  assign n4308 = ~n2365 & n4307 ;
  assign n4309 = ~n4300 & ~n4308 ;
  assign n4310 = ~\sa32_reg[2]/P0001  & ~n2328 ;
  assign n4311 = n2059 & n2399 ;
  assign n4312 = ~n1966 & ~n2347 ;
  assign n4313 = ~n4311 & n4312 ;
  assign n4314 = ~n4310 & n4313 ;
  assign n4315 = ~n4309 & n4314 ;
  assign n4316 = ~\sa32_reg[0]/P0002  & ~n4315 ;
  assign n4266 = n1926 & ~n1959 ;
  assign n4267 = \sa32_reg[2]/P0001  & ~n4266 ;
  assign n4264 = ~n1989 & ~n2366 ;
  assign n4265 = ~\sa32_reg[2]/P0001  & ~n4264 ;
  assign n4268 = ~n2040 & ~n2345 ;
  assign n4269 = ~n3490 & n4268 ;
  assign n4270 = ~n4265 & n4269 ;
  assign n4271 = ~n4267 & n4270 ;
  assign n4272 = ~\sa32_reg[1]/P0001  & ~n4271 ;
  assign n4278 = ~n3143 & ~n3149 ;
  assign n4279 = ~n3457 & n4278 ;
  assign n4280 = \sa32_reg[2]/P0001  & ~n4279 ;
  assign n4281 = ~n1937 & ~n1982 ;
  assign n4282 = ~\sa32_reg[2]/P0001  & ~n4281 ;
  assign n4277 = ~n2024 & ~n3194 ;
  assign n4283 = ~n1921 & n4277 ;
  assign n4284 = ~n4282 & n4283 ;
  assign n4285 = ~n4280 & n4284 ;
  assign n4286 = \sa32_reg[1]/P0001  & ~n4285 ;
  assign n4273 = n3280 & ~n3367 ;
  assign n4274 = ~\sa32_reg[2]/P0001  & ~n4273 ;
  assign n4275 = ~n1932 & n2042 ;
  assign n4276 = n2046 & ~n4275 ;
  assign n4287 = ~n1971 & ~n4276 ;
  assign n4288 = ~n4274 & n4287 ;
  assign n4289 = ~n4286 & n4288 ;
  assign n4290 = ~n4272 & n4289 ;
  assign n4291 = \sa32_reg[0]/P0002  & ~n4290 ;
  assign n4321 = ~n1994 & ~n3180 ;
  assign n4322 = ~n3374 & n4321 ;
  assign n4323 = n2313 & ~n4322 ;
  assign n4317 = n1925 & n2030 ;
  assign n4318 = \sa32_reg[6]/NET0131  & n1952 ;
  assign n4319 = n4277 & ~n4318 ;
  assign n4320 = \sa32_reg[2]/P0001  & ~n4319 ;
  assign n4324 = ~n4317 & ~n4320 ;
  assign n4325 = ~n4323 & n4324 ;
  assign n4326 = \sa32_reg[1]/P0001  & ~n4325 ;
  assign n4329 = \sa32_reg[2]/P0001  & ~n1938 ;
  assign n4330 = ~n1966 & n4329 ;
  assign n4331 = ~\sa32_reg[2]/P0001  & ~n3172 ;
  assign n4332 = ~\sa32_reg[1]/P0001  & ~n4331 ;
  assign n4333 = ~n4330 & n4332 ;
  assign n4327 = ~n3181 & ~n3408 ;
  assign n4328 = n2059 & ~n4327 ;
  assign n4334 = ~n3437 & ~n4328 ;
  assign n4335 = ~n4333 & n4334 ;
  assign n4336 = ~n4326 & n4335 ;
  assign n4337 = ~n4291 & n4336 ;
  assign n4338 = ~n4316 & n4337 ;
  assign n4339 = n3416 & ~n4338 ;
  assign n4340 = ~n3416 & n4338 ;
  assign n4341 = ~n4339 & ~n4340 ;
  assign n4342 = \u0_w_reg[3][12]/P0001  & ~n3205 ;
  assign n4343 = ~\u0_w_reg[3][12]/P0001  & n3205 ;
  assign n4344 = ~n4342 & ~n4343 ;
  assign n4345 = n4341 & n4344 ;
  assign n4346 = ~n4341 & ~n4344 ;
  assign n4347 = ~n4345 & ~n4346 ;
  assign n4348 = n2529 & ~n4059 ;
  assign n4349 = ~n2529 & n4059 ;
  assign n4350 = ~n4348 & ~n4349 ;
  assign n4351 = ~n2739 & n4350 ;
  assign n4352 = n2739 & ~n4350 ;
  assign n4353 = ~n4351 & ~n4352 ;
  assign n4355 = ~n4347 & n4353 ;
  assign n4354 = n4347 & ~n4353 ;
  assign n4356 = ~\ld_r_reg/P0001  & ~n4354 ;
  assign n4357 = ~n4355 & n4356 ;
  assign n4359 = ~\text_in_r_reg[12]/P0001  & \u0_w_reg[3][12]/P0001  ;
  assign n4358 = \text_in_r_reg[12]/P0001  & ~\u0_w_reg[3][12]/P0001  ;
  assign n4360 = \ld_r_reg/P0001  & ~n4358 ;
  assign n4361 = ~n4359 & n4360 ;
  assign n4362 = ~n4357 & ~n4361 ;
  assign n4364 = ~n2123 & ~n2566 ;
  assign n4365 = ~n2576 & ~n2586 ;
  assign n4366 = n4364 & n4365 ;
  assign n4367 = ~n1616 & ~n2622 ;
  assign n4363 = n1698 & n2595 ;
  assign n4368 = ~n2635 & ~n4363 ;
  assign n4369 = n4367 & n4368 ;
  assign n4370 = n4366 & n4369 ;
  assign n4371 = ~\sa10_reg[1]/P0001  & ~n4370 ;
  assign n4377 = n1629 & n1666 ;
  assign n4378 = n1607 & n4377 ;
  assign n4376 = n2142 & n3616 ;
  assign n4379 = n1586 & n2112 ;
  assign n4380 = ~n4376 & ~n4379 ;
  assign n4381 = ~n4378 & n4380 ;
  assign n4382 = \sa10_reg[1]/P0001  & ~n4381 ;
  assign n4373 = ~n1708 & ~n2809 ;
  assign n4374 = ~n2119 & n4373 ;
  assign n4375 = n1664 & ~n4374 ;
  assign n4372 = \sa10_reg[5]/P0001  & n2576 ;
  assign n4383 = ~n2559 & ~n4372 ;
  assign n4384 = ~n2572 & n4383 ;
  assign n4385 = ~n4375 & n4384 ;
  assign n4386 = ~n4382 & n4385 ;
  assign n4387 = ~n4371 & n4386 ;
  assign n4388 = \sa10_reg[0]/P0001  & ~n4387 ;
  assign n4417 = ~n1698 & ~n2608 ;
  assign n4418 = \sa10_reg[2]/P0001  & ~n4417 ;
  assign n4419 = ~n1586 & ~n1681 ;
  assign n4420 = ~\sa10_reg[2]/P0001  & ~n1629 ;
  assign n4421 = ~n4419 & n4420 ;
  assign n4422 = ~n1700 & ~n4421 ;
  assign n4423 = ~n4418 & n4422 ;
  assign n4424 = ~\sa10_reg[0]/P0001  & ~n4423 ;
  assign n4414 = \sa10_reg[4]/P0001  & n3641 ;
  assign n4415 = n3614 & ~n4414 ;
  assign n4416 = ~\sa10_reg[2]/P0001  & ~n4415 ;
  assign n4425 = ~n2565 & ~n4416 ;
  assign n4426 = ~n4424 & n4425 ;
  assign n4427 = \sa10_reg[1]/P0001  & ~n4426 ;
  assign n4389 = n2190 & ~n3922 ;
  assign n4390 = ~n2567 & n4389 ;
  assign n4391 = ~n1683 & ~n2101 ;
  assign n4392 = ~n1712 & n4391 ;
  assign n4393 = n1617 & n4392 ;
  assign n4394 = ~n4390 & ~n4393 ;
  assign n4395 = ~n1583 & ~n1586 ;
  assign n4396 = n1650 & n4395 ;
  assign n4397 = ~n4394 & ~n4396 ;
  assign n4398 = ~\sa10_reg[1]/P0001  & ~n4397 ;
  assign n4405 = ~n2189 & ~n4377 ;
  assign n4406 = ~\sa10_reg[1]/P0001  & ~n4405 ;
  assign n4407 = n2607 & n3943 ;
  assign n4408 = ~n1613 & ~n4407 ;
  assign n4409 = ~n1728 & n4408 ;
  assign n4410 = ~n4406 & n4409 ;
  assign n4411 = ~\sa10_reg[0]/P0001  & ~n4410 ;
  assign n4399 = ~n1608 & ~n1615 ;
  assign n4400 = n1668 & ~n4399 ;
  assign n4401 = ~n1669 & ~n2634 ;
  assign n4402 = \sa10_reg[1]/P0001  & ~n4401 ;
  assign n4403 = ~n4400 & ~n4402 ;
  assign n4404 = \sa10_reg[2]/P0001  & ~n4403 ;
  assign n4412 = \sa10_reg[1]/P0001  & n1664 ;
  assign n4413 = n2093 & n4412 ;
  assign n4428 = ~n3923 & ~n4413 ;
  assign n4429 = ~n4404 & n4428 ;
  assign n4430 = ~n4411 & n4429 ;
  assign n4431 = ~n4398 & n4430 ;
  assign n4432 = ~n4427 & n4431 ;
  assign n4433 = ~n4388 & n4432 ;
  assign n4460 = ~\sa03_reg[7]/NET0131  & n1408 ;
  assign n4461 = ~n1447 & ~n4460 ;
  assign n4462 = \sa03_reg[2]/P0001  & ~n4461 ;
  assign n4457 = ~n1383 & ~n1398 ;
  assign n4458 = ~\sa03_reg[2]/P0001  & ~n1449 ;
  assign n4459 = ~n4457 & n4458 ;
  assign n4463 = \sa03_reg[1]/P0001  & ~n1565 ;
  assign n4464 = ~n4459 & n4463 ;
  assign n4465 = ~n4462 & n4464 ;
  assign n4466 = n1429 & n1449 ;
  assign n4467 = ~\sa03_reg[1]/P0001  & ~n2293 ;
  assign n4468 = ~n4466 & n4467 ;
  assign n4469 = ~n4465 & ~n4468 ;
  assign n4471 = \sa03_reg[2]/P0001  & n2249 ;
  assign n4470 = ~\sa03_reg[2]/P0001  & n1417 ;
  assign n4472 = ~\sa03_reg[0]/P0001  & ~n1365 ;
  assign n4473 = ~n4470 & n4472 ;
  assign n4474 = ~n4471 & n4473 ;
  assign n4475 = ~n4469 & n4474 ;
  assign n4476 = ~\sa03_reg[2]/P0001  & n1409 ;
  assign n4481 = n2656 & ~n2715 ;
  assign n4482 = ~n4476 & n4481 ;
  assign n4478 = ~n1504 & ~n2650 ;
  assign n4477 = n1318 & n1436 ;
  assign n4479 = ~n4102 & ~n4477 ;
  assign n4480 = n4478 & n4479 ;
  assign n4483 = ~n2707 & n4480 ;
  assign n4484 = n4482 & n4483 ;
  assign n4486 = n1555 & n3818 ;
  assign n4485 = n1383 & n1384 ;
  assign n4487 = \sa03_reg[1]/P0001  & ~n4485 ;
  assign n4488 = ~n4486 & n4487 ;
  assign n4489 = ~n4140 & n4488 ;
  assign n4490 = ~n4484 & ~n4489 ;
  assign n4492 = ~n1353 & ~n1414 ;
  assign n4493 = ~n1566 & n4492 ;
  assign n4494 = n1374 & ~n4493 ;
  assign n4495 = \sa03_reg[0]/P0001  & ~n2676 ;
  assign n4491 = n1435 & n1436 ;
  assign n4496 = ~n2678 & ~n4491 ;
  assign n4497 = n4495 & n4496 ;
  assign n4498 = ~n4494 & n4497 ;
  assign n4499 = ~n4490 & n4498 ;
  assign n4500 = ~n4475 & ~n4499 ;
  assign n4451 = \sa03_reg[4]/P0001  & n3692 ;
  assign n4452 = n3713 & ~n4451 ;
  assign n4453 = ~\sa03_reg[2]/P0001  & ~n4452 ;
  assign n4449 = ~n1397 & ~n3830 ;
  assign n4450 = \sa03_reg[2]/P0001  & ~n4449 ;
  assign n4454 = ~n1328 & ~n4450 ;
  assign n4455 = ~n4453 & n4454 ;
  assign n4456 = \sa03_reg[1]/P0001  & ~n4455 ;
  assign n4434 = ~n1383 & n3746 ;
  assign n4435 = ~\sa03_reg[6]/NET0131  & n1324 ;
  assign n4436 = \sa03_reg[2]/P0001  & ~n2293 ;
  assign n4437 = ~n4435 & n4436 ;
  assign n4438 = ~n2685 & n4437 ;
  assign n4439 = ~\sa03_reg[2]/P0001  & ~n1416 ;
  assign n4440 = ~n1504 & n4439 ;
  assign n4441 = ~n1400 & ~n1572 ;
  assign n4442 = n4440 & n4441 ;
  assign n4443 = ~n4438 & ~n4442 ;
  assign n4444 = ~n4434 & ~n4443 ;
  assign n4445 = ~\sa03_reg[1]/P0001  & ~n4444 ;
  assign n4448 = ~n4118 & n4138 ;
  assign n4446 = \sa03_reg[1]/P0001  & n1374 ;
  assign n4447 = n2200 & n4446 ;
  assign n4501 = ~n3845 & ~n4447 ;
  assign n4502 = ~n4448 & n4501 ;
  assign n4503 = ~n4445 & n4502 ;
  assign n4504 = ~n4456 & n4503 ;
  assign n4505 = ~n4500 & n4504 ;
  assign n4506 = n4433 & ~n4505 ;
  assign n4507 = ~n4433 & n4505 ;
  assign n4508 = ~n4506 & ~n4507 ;
  assign n4509 = ~n3768 & ~n4508 ;
  assign n4510 = n3768 & n4508 ;
  assign n4511 = ~n4509 & ~n4510 ;
  assign n4541 = ~n3021 & ~n3029 ;
  assign n4538 = n1761 & n1831 ;
  assign n4542 = ~n3545 & ~n4538 ;
  assign n4543 = n4541 & n4542 ;
  assign n4540 = ~\sa21_reg[1]/P0001  & ~n1800 ;
  assign n4544 = ~n2900 & n4540 ;
  assign n4539 = n2437 & n2479 ;
  assign n4545 = ~n2997 & ~n4539 ;
  assign n4546 = n4544 & n4545 ;
  assign n4547 = n4543 & n4546 ;
  assign n4549 = ~n1844 & ~n2450 ;
  assign n4550 = ~\sa21_reg[2]/P0001  & ~n4549 ;
  assign n4548 = \sa21_reg[2]/P0001  & n2862 ;
  assign n4551 = \sa21_reg[1]/P0001  & ~n3572 ;
  assign n4552 = ~n4548 & n4551 ;
  assign n4553 = ~n4550 & n4552 ;
  assign n4554 = ~n4547 & ~n4553 ;
  assign n4535 = ~n1781 & ~n1884 ;
  assign n4536 = ~n2493 & n4535 ;
  assign n4537 = n1894 & ~n4536 ;
  assign n4555 = \sa21_reg[0]/P0001  & ~n3049 ;
  assign n4556 = ~n3055 & ~n4176 ;
  assign n4557 = n4555 & n4556 ;
  assign n4558 = ~n4537 & n4557 ;
  assign n4559 = ~n4554 & n4558 ;
  assign n4560 = ~\sa21_reg[1]/P0001  & ~n2508 ;
  assign n4561 = ~n3571 & n4560 ;
  assign n4562 = ~n1785 & ~n4019 ;
  assign n4563 = n3555 & n4562 ;
  assign n4564 = \sa21_reg[2]/P0001  & ~n2437 ;
  assign n4565 = ~n2876 & n4564 ;
  assign n4566 = ~n4563 & ~n4565 ;
  assign n4567 = \sa21_reg[1]/P0001  & ~n1885 ;
  assign n4568 = ~n4566 & n4567 ;
  assign n4569 = ~n4561 & ~n4568 ;
  assign n4570 = \sa21_reg[2]/P0001  & n2465 ;
  assign n4571 = ~\sa21_reg[0]/P0001  & ~n1792 ;
  assign n4572 = ~n1881 & n4571 ;
  assign n4573 = ~n4570 & n4572 ;
  assign n4574 = ~n4569 & n4573 ;
  assign n4575 = ~n4559 & ~n4574 ;
  assign n4514 = n1801 & ~n1855 ;
  assign n4515 = ~n1880 & ~n1889 ;
  assign n4516 = n4514 & n4515 ;
  assign n4517 = \sa21_reg[2]/P0001  & ~n2508 ;
  assign n4518 = ~n2857 & n4517 ;
  assign n4519 = ~n3050 & n4518 ;
  assign n4520 = ~n4516 & ~n4519 ;
  assign n4521 = ~\sa21_reg[1]/P0001  & ~n2993 ;
  assign n4522 = ~n2522 & n4521 ;
  assign n4523 = ~n4520 & n4522 ;
  assign n4524 = n1759 & n1854 ;
  assign n4525 = \sa21_reg[2]/P0001  & ~n1816 ;
  assign n4526 = ~n1834 & n4525 ;
  assign n4527 = ~n4524 & n4526 ;
  assign n4528 = \sa21_reg[4]/P0001  & n3542 ;
  assign n4529 = ~\sa21_reg[2]/P0001  & ~n4528 ;
  assign n4530 = n4196 & n4529 ;
  assign n4531 = ~n4527 & ~n4530 ;
  assign n4532 = \sa21_reg[1]/P0001  & ~n2838 ;
  assign n4533 = ~n4531 & n4532 ;
  assign n4534 = ~n4523 & ~n4533 ;
  assign n4512 = ~n2422 & ~n2452 ;
  assign n4513 = n2453 & ~n4512 ;
  assign n4576 = ~n4014 & ~n4513 ;
  assign n4577 = ~n4534 & n4576 ;
  assign n4578 = ~n4575 & n4577 ;
  assign n4579 = \u0_w_reg[3][2]/P0001  & ~n4578 ;
  assign n4580 = ~\u0_w_reg[3][2]/P0001  & n4578 ;
  assign n4581 = ~n4579 & ~n4580 ;
  assign n4582 = n3503 & n4581 ;
  assign n4583 = ~n3503 & ~n4581 ;
  assign n4584 = ~n4582 & ~n4583 ;
  assign n4586 = n4511 & ~n4584 ;
  assign n4585 = ~n4511 & n4584 ;
  assign n4587 = ~\ld_r_reg/P0001  & ~n4585 ;
  assign n4588 = ~n4586 & n4587 ;
  assign n4590 = \text_in_r_reg[2]/P0001  & \u0_w_reg[3][2]/P0001  ;
  assign n4589 = ~\text_in_r_reg[2]/P0001  & ~\u0_w_reg[3][2]/P0001  ;
  assign n4591 = \ld_r_reg/P0001  & ~n4589 ;
  assign n4592 = ~n4590 & n4591 ;
  assign n4593 = ~n4588 & ~n4592 ;
  assign n4594 = n3681 & ~n4248 ;
  assign n4595 = ~n3681 & n4248 ;
  assign n4596 = ~n4594 & ~n4595 ;
  assign n4597 = \u0_w_reg[3][25]/P0001  & ~n3503 ;
  assign n4598 = ~\u0_w_reg[3][25]/P0001  & n3503 ;
  assign n4599 = ~n4597 & ~n4598 ;
  assign n4600 = n4596 & n4599 ;
  assign n4601 = ~n4596 & ~n4599 ;
  assign n4602 = ~n4600 & ~n4601 ;
  assign n4616 = ~n2168 & ~n2634 ;
  assign n4617 = \sa10_reg[2]/P0001  & ~n4616 ;
  assign n4618 = ~n2113 & ~n2740 ;
  assign n4619 = ~\sa10_reg[3]/P0001  & ~n4618 ;
  assign n4615 = \sa10_reg[4]/P0001  & n2155 ;
  assign n4620 = \sa10_reg[5]/P0001  & ~n1597 ;
  assign n4621 = n1627 & ~n4620 ;
  assign n4622 = ~n4615 & ~n4621 ;
  assign n4623 = ~n4619 & n4622 ;
  assign n4624 = ~n4617 & n4623 ;
  assign n4625 = ~\sa10_reg[1]/P0001  & ~n4624 ;
  assign n4612 = ~n2625 & ~n2748 ;
  assign n4613 = n1632 & n4612 ;
  assign n4614 = \sa10_reg[2]/P0001  & ~n4613 ;
  assign n4607 = ~n1586 & ~n1672 ;
  assign n4608 = \sa10_reg[3]/P0001  & ~n4607 ;
  assign n4609 = ~n2118 & ~n2160 ;
  assign n4610 = ~n4608 & n4609 ;
  assign n4611 = ~\sa10_reg[2]/P0001  & ~n4610 ;
  assign n4603 = ~\sa10_reg[5]/P0001  & ~n1614 ;
  assign n4604 = n2142 & ~n4603 ;
  assign n4605 = ~n1708 & ~n4604 ;
  assign n4606 = \sa10_reg[1]/P0001  & ~n4605 ;
  assign n4626 = ~n2554 & ~n3599 ;
  assign n4627 = ~n4606 & n4626 ;
  assign n4628 = ~n4611 & n4627 ;
  assign n4629 = ~n4614 & n4628 ;
  assign n4630 = ~n4625 & n4629 ;
  assign n4631 = \sa10_reg[0]/P0001  & ~n4630 ;
  assign n4641 = n1650 & n1668 ;
  assign n4642 = n3940 & ~n4641 ;
  assign n4643 = ~\sa10_reg[2]/P0001  & ~n4642 ;
  assign n4632 = ~\sa10_reg[3]/P0001  & ~n2094 ;
  assign n4633 = n2592 & ~n4632 ;
  assign n4635 = ~n1594 & ~n1614 ;
  assign n4636 = ~n3624 & ~n4635 ;
  assign n4634 = n1664 & n2621 ;
  assign n4637 = \sa10_reg[1]/P0001  & ~n2154 ;
  assign n4638 = ~n4634 & n4637 ;
  assign n4639 = ~n4636 & n4638 ;
  assign n4640 = ~n4633 & ~n4639 ;
  assign n4644 = ~n1615 & ~n1672 ;
  assign n4645 = n1715 & ~n4644 ;
  assign n4646 = \sa10_reg[7]/NET0131  & n2183 ;
  assign n4647 = n3615 & n4646 ;
  assign n4648 = ~n4645 & ~n4647 ;
  assign n4649 = ~n4640 & n4648 ;
  assign n4650 = ~n4643 & n4649 ;
  assign n4651 = ~\sa10_reg[0]/P0001  & ~n4650 ;
  assign n4652 = ~n2148 & ~n2787 ;
  assign n4653 = ~n2572 & n4652 ;
  assign n4654 = ~\sa10_reg[2]/P0001  & ~n4653 ;
  assign n4655 = ~n2807 & ~n4378 ;
  assign n4656 = ~n4654 & n4655 ;
  assign n4657 = ~\sa10_reg[1]/P0001  & ~n4656 ;
  assign n4659 = ~n1730 & ~n2577 ;
  assign n4660 = ~\sa10_reg[5]/P0001  & ~n4659 ;
  assign n4661 = ~\sa10_reg[2]/P0001  & ~n2189 ;
  assign n4662 = ~n2602 & ~n4661 ;
  assign n4663 = ~n1727 & ~n4662 ;
  assign n4664 = ~n4660 & n4663 ;
  assign n4665 = \sa10_reg[1]/P0001  & ~n4664 ;
  assign n4658 = \sa10_reg[6]/NET0131  & n1667 ;
  assign n4667 = \sa10_reg[1]/P0001  & ~n2179 ;
  assign n4666 = ~n1711 & ~n2559 ;
  assign n4668 = \sa10_reg[2]/P0001  & ~n4666 ;
  assign n4669 = ~n4667 & n4668 ;
  assign n4670 = ~n4658 & ~n4669 ;
  assign n4671 = ~n4665 & n4670 ;
  assign n4672 = ~n4657 & n4671 ;
  assign n4673 = ~n4651 & n4672 ;
  assign n4674 = ~n4631 & n4673 ;
  assign n4675 = n4161 & ~n4674 ;
  assign n4676 = ~n4161 & n4674 ;
  assign n4677 = ~n4675 & ~n4676 ;
  assign n4678 = ~n2307 & n4677 ;
  assign n4679 = n2307 & ~n4677 ;
  assign n4680 = ~n4678 & ~n4679 ;
  assign n4682 = n4602 & n4680 ;
  assign n4681 = ~n4602 & ~n4680 ;
  assign n4683 = ~\ld_r_reg/P0001  & ~n4681 ;
  assign n4684 = ~n4682 & n4683 ;
  assign n4686 = \text_in_r_reg[25]/P0001  & \u0_w_reg[3][25]/P0001  ;
  assign n4685 = ~\text_in_r_reg[25]/P0001  & ~\u0_w_reg[3][25]/P0001  ;
  assign n4687 = \ld_r_reg/P0001  & ~n4685 ;
  assign n4688 = ~n4686 & n4687 ;
  assign n4689 = ~n4684 & ~n4688 ;
  assign n4690 = ~n1908 & ~n2307 ;
  assign n4691 = n1908 & n2307 ;
  assign n4692 = ~n4690 & ~n4691 ;
  assign n4693 = \u0_w_reg[3][15]/P0001  & ~n3416 ;
  assign n4694 = ~\u0_w_reg[3][15]/P0001  & n3416 ;
  assign n4695 = ~n4693 & ~n4694 ;
  assign n4696 = n2416 & n4695 ;
  assign n4697 = ~n2416 & ~n4695 ;
  assign n4698 = ~n4696 & ~n4697 ;
  assign n4700 = n4692 & n4698 ;
  assign n4699 = ~n4692 & ~n4698 ;
  assign n4701 = ~\ld_r_reg/P0001  & ~n4699 ;
  assign n4702 = ~n4700 & n4701 ;
  assign n4704 = ~\text_in_r_reg[15]/P0001  & \u0_w_reg[3][15]/P0001  ;
  assign n4703 = \text_in_r_reg[15]/P0001  & ~\u0_w_reg[3][15]/P0001  ;
  assign n4705 = \ld_r_reg/P0001  & ~n4703 ;
  assign n4706 = ~n4704 & n4705 ;
  assign n4707 = ~n4702 & ~n4706 ;
  assign n4708 = n2304 & ~n3888 ;
  assign n4709 = ~n2304 & n3888 ;
  assign n4710 = ~n4708 & ~n4709 ;
  assign n4711 = n2739 & n4710 ;
  assign n4712 = ~n2739 & ~n4710 ;
  assign n4713 = ~n4711 & ~n4712 ;
  assign n4714 = \u0_w_reg[3][4]/P0001  & ~n3069 ;
  assign n4715 = ~\u0_w_reg[3][4]/P0001  & n3069 ;
  assign n4716 = ~n4714 & ~n4715 ;
  assign n4717 = n4341 & n4716 ;
  assign n4718 = ~n4341 & ~n4716 ;
  assign n4719 = ~n4717 & ~n4718 ;
  assign n4721 = n4713 & n4719 ;
  assign n4720 = ~n4713 & ~n4719 ;
  assign n4722 = ~\ld_r_reg/P0001  & ~n4720 ;
  assign n4723 = ~n4721 & n4722 ;
  assign n4725 = ~\text_in_r_reg[4]/P0001  & \u0_w_reg[3][4]/P0001  ;
  assign n4724 = \text_in_r_reg[4]/P0001  & ~\u0_w_reg[3][4]/P0001  ;
  assign n4726 = \ld_r_reg/P0001  & ~n4724 ;
  assign n4727 = ~n4725 & n4726 ;
  assign n4728 = ~n4723 & ~n4727 ;
  assign n4729 = \u0_w_reg[3][27]/P0001  & ~n4338 ;
  assign n4730 = ~\u0_w_reg[3][27]/P0001  & n4338 ;
  assign n4731 = ~n4729 & ~n4730 ;
  assign n4732 = n4062 & n4731 ;
  assign n4733 = ~n4062 & ~n4731 ;
  assign n4734 = ~n4732 & ~n4733 ;
  assign n4735 = ~n2307 & n4508 ;
  assign n4736 = n2307 & ~n4508 ;
  assign n4737 = ~n4735 & ~n4736 ;
  assign n4739 = ~n4734 & n4737 ;
  assign n4738 = n4734 & ~n4737 ;
  assign n4740 = ~\ld_r_reg/P0001  & ~n4738 ;
  assign n4741 = ~n4739 & n4740 ;
  assign n4743 = ~\text_in_r_reg[27]/P0001  & \u0_w_reg[3][27]/P0001  ;
  assign n4742 = \text_in_r_reg[27]/P0001  & ~\u0_w_reg[3][27]/P0001  ;
  assign n4744 = \ld_r_reg/P0001  & ~n4742 ;
  assign n4745 = ~n4743 & n4744 ;
  assign n4746 = ~n4741 & ~n4745 ;
  assign n4747 = \u0_w_reg[3][19]/P0001  & ~n4338 ;
  assign n4748 = ~\u0_w_reg[3][19]/P0001  & n4338 ;
  assign n4749 = ~n4747 & ~n4748 ;
  assign n4750 = n4350 & n4749 ;
  assign n4751 = ~n4350 & ~n4749 ;
  assign n4752 = ~n4750 & ~n4751 ;
  assign n4753 = n4433 & ~n4578 ;
  assign n4754 = ~n4433 & n4578 ;
  assign n4755 = ~n4753 & ~n4754 ;
  assign n4756 = n2199 & ~n3888 ;
  assign n4757 = ~n2199 & n3888 ;
  assign n4758 = ~n4756 & ~n4757 ;
  assign n4759 = n4755 & n4758 ;
  assign n4760 = ~n4755 & ~n4758 ;
  assign n4761 = ~n4759 & ~n4760 ;
  assign n4763 = n4752 & n4761 ;
  assign n4762 = ~n4752 & ~n4761 ;
  assign n4764 = ~\ld_r_reg/P0001  & ~n4762 ;
  assign n4765 = ~n4763 & n4764 ;
  assign n4767 = ~\text_in_r_reg[19]/P0001  & \u0_w_reg[3][19]/P0001  ;
  assign n4766 = \text_in_r_reg[19]/P0001  & ~\u0_w_reg[3][19]/P0001  ;
  assign n4768 = \ld_r_reg/P0001  & ~n4766 ;
  assign n4769 = ~n4767 & n4768 ;
  assign n4770 = ~n4765 & ~n4769 ;
  assign n4771 = n3592 & ~n4674 ;
  assign n4772 = ~n3592 & n4674 ;
  assign n4773 = ~n4771 & ~n4772 ;
  assign n4774 = n2199 & ~n3768 ;
  assign n4775 = ~n2199 & n3768 ;
  assign n4776 = ~n4774 & ~n4775 ;
  assign n4777 = n4773 & n4776 ;
  assign n4778 = ~n4773 & ~n4776 ;
  assign n4779 = ~n4777 & ~n4778 ;
  assign n4780 = ~n2529 & ~n3503 ;
  assign n4781 = n2529 & n3503 ;
  assign n4782 = ~n4780 & ~n4781 ;
  assign n4783 = \u0_w_reg[3][17]/P0001  & ~n4248 ;
  assign n4784 = ~\u0_w_reg[3][17]/P0001  & n4248 ;
  assign n4785 = ~n4783 & ~n4784 ;
  assign n4786 = n4782 & n4785 ;
  assign n4787 = ~n4782 & ~n4785 ;
  assign n4788 = ~n4786 & ~n4787 ;
  assign n4790 = n4779 & n4788 ;
  assign n4789 = ~n4779 & ~n4788 ;
  assign n4791 = ~\ld_r_reg/P0001  & ~n4789 ;
  assign n4792 = ~n4790 & n4791 ;
  assign n4794 = \text_in_r_reg[17]/P0001  & \u0_w_reg[3][17]/P0001  ;
  assign n4793 = ~\text_in_r_reg[17]/P0001  & ~\u0_w_reg[3][17]/P0001  ;
  assign n4795 = \ld_r_reg/P0001  & ~n4793 ;
  assign n4796 = ~n4794 & n4795 ;
  assign n4797 = ~n4792 & ~n4796 ;
  assign n4798 = n2529 & ~n4578 ;
  assign n4799 = ~n2529 & n4578 ;
  assign n4800 = ~n4798 & ~n4799 ;
  assign n4801 = n3969 & n4800 ;
  assign n4802 = ~n3969 & ~n4800 ;
  assign n4803 = ~n4801 & ~n4802 ;
  assign n4832 = ~n3184 & ~n3257 ;
  assign n4833 = ~n1964 & n4832 ;
  assign n4834 = ~n2332 & n3173 ;
  assign n4830 = ~n1924 & n2067 ;
  assign n4831 = ~\sa32_reg[2]/P0001  & n2040 ;
  assign n4835 = ~n4830 & ~n4831 ;
  assign n4836 = n4834 & n4835 ;
  assign n4837 = n4833 & n4836 ;
  assign n4838 = ~\sa32_reg[2]/P0001  & ~n1947 ;
  assign n4839 = n3363 & n4838 ;
  assign n4840 = \sa32_reg[1]/P0001  & ~n2349 ;
  assign n4841 = ~n3309 & n4840 ;
  assign n4842 = ~n4839 & n4841 ;
  assign n4843 = ~n4837 & ~n4842 ;
  assign n4827 = ~n2011 & ~n2351 ;
  assign n4828 = ~n3331 & n4827 ;
  assign n4829 = n2059 & ~n4828 ;
  assign n4844 = ~n2068 & ~n3146 ;
  assign n4845 = ~\sa32_reg[3]/P0001  & ~n4844 ;
  assign n4846 = \sa32_reg[0]/P0002  & ~n3126 ;
  assign n4847 = ~n4845 & n4846 ;
  assign n4848 = ~n4829 & n4847 ;
  assign n4849 = ~n4843 & n4848 ;
  assign n4853 = ~n1949 & ~n3376 ;
  assign n4854 = \sa32_reg[2]/P0001  & ~n4853 ;
  assign n4850 = ~n1947 & ~n1948 ;
  assign n4851 = ~\sa32_reg[2]/P0001  & ~n1934 ;
  assign n4852 = ~n4850 & n4851 ;
  assign n4855 = \sa32_reg[1]/P0001  & ~n2352 ;
  assign n4856 = ~n4852 & n4855 ;
  assign n4857 = ~n4854 & n4856 ;
  assign n4858 = ~\sa32_reg[1]/P0001  & ~n1921 ;
  assign n4859 = ~n3308 & n4858 ;
  assign n4860 = ~n4857 & ~n4859 ;
  assign n4861 = \sa32_reg[6]/NET0131  & n3326 ;
  assign n4862 = ~\sa32_reg[0]/P0002  & ~n2024 ;
  assign n4863 = ~n2368 & n4862 ;
  assign n4864 = ~n4861 & n4863 ;
  assign n4865 = ~n4860 & n4864 ;
  assign n4866 = ~n4849 & ~n4865 ;
  assign n4808 = ~n2006 & n3451 ;
  assign n4809 = ~\sa32_reg[2]/P0001  & ~n4808 ;
  assign n4804 = ~\sa32_reg[4]/P0001  & n2366 ;
  assign n4805 = ~n1963 & ~n2050 ;
  assign n4806 = ~n4804 & n4805 ;
  assign n4807 = \sa32_reg[2]/P0001  & ~n4806 ;
  assign n4810 = \sa32_reg[1]/P0001  & ~n1989 ;
  assign n4811 = ~n4807 & n4810 ;
  assign n4812 = ~n4809 & n4811 ;
  assign n4815 = ~n2356 & ~n3405 ;
  assign n4816 = ~n2052 & n4815 ;
  assign n4817 = n2333 & n4816 ;
  assign n4818 = ~n1991 & ~n3134 ;
  assign n4819 = n3388 & n4818 ;
  assign n4820 = ~n4817 & ~n4819 ;
  assign n4813 = ~n1919 & ~n1948 ;
  assign n4814 = n1990 & n4813 ;
  assign n4821 = ~\sa32_reg[1]/P0001  & ~n4814 ;
  assign n4822 = ~n4820 & n4821 ;
  assign n4823 = ~n4812 & ~n4822 ;
  assign n4824 = ~n2060 & ~n2387 ;
  assign n4825 = ~\sa32_reg[3]/P0001  & n2348 ;
  assign n4826 = ~n4824 & n4825 ;
  assign n4867 = ~n4317 & ~n4826 ;
  assign n4868 = ~n4823 & n4867 ;
  assign n4869 = ~n4866 & n4868 ;
  assign n4870 = \u0_w_reg[3][11]/P0001  & ~n4869 ;
  assign n4871 = ~\u0_w_reg[3][11]/P0001  & n4869 ;
  assign n4872 = ~n4870 & ~n4871 ;
  assign n4873 = n4341 & n4872 ;
  assign n4874 = ~n4341 & ~n4872 ;
  assign n4875 = ~n4873 & ~n4874 ;
  assign n4877 = n4803 & n4875 ;
  assign n4876 = ~n4803 & ~n4875 ;
  assign n4878 = ~\ld_r_reg/P0001  & ~n4876 ;
  assign n4879 = ~n4877 & n4878 ;
  assign n4881 = ~\text_in_r_reg[11]/P0001  & \u0_w_reg[3][11]/P0001  ;
  assign n4880 = \text_in_r_reg[11]/P0001  & ~\u0_w_reg[3][11]/P0001  ;
  assign n4882 = \ld_r_reg/P0001  & ~n4880 ;
  assign n4883 = ~n4881 & n4882 ;
  assign n4884 = ~n4879 & ~n4883 ;
  assign n4885 = \u0_w_reg[3][26]/P0001  & ~n4869 ;
  assign n4886 = ~\u0_w_reg[3][26]/P0001  & n4869 ;
  assign n4887 = ~n4885 & ~n4886 ;
  assign n4888 = n4755 & n4887 ;
  assign n4889 = ~n4755 & ~n4887 ;
  assign n4890 = ~n4888 & ~n4889 ;
  assign n4892 = n3771 & n4890 ;
  assign n4891 = ~n3771 & ~n4890 ;
  assign n4893 = ~\ld_r_reg/P0001  & ~n4891 ;
  assign n4894 = ~n4892 & n4893 ;
  assign n4896 = ~\text_in_r_reg[26]/P0001  & \u0_w_reg[3][26]/P0001  ;
  assign n4895 = \text_in_r_reg[26]/P0001  & ~\u0_w_reg[3][26]/P0001  ;
  assign n4897 = \ld_r_reg/P0001  & ~n4895 ;
  assign n4898 = ~n4896 & n4897 ;
  assign n4899 = ~n4894 & ~n4898 ;
  assign n4900 = n2304 & ~n4505 ;
  assign n4901 = ~n2304 & n4505 ;
  assign n4902 = ~n4900 & ~n4901 ;
  assign n4903 = n3969 & n4902 ;
  assign n4904 = ~n3969 & ~n4902 ;
  assign n4905 = ~n4903 & ~n4904 ;
  assign n4906 = ~n3416 & ~n4059 ;
  assign n4907 = n3416 & n4059 ;
  assign n4908 = ~n4906 & ~n4907 ;
  assign n4909 = \u0_w_reg[3][3]/P0001  & ~n4869 ;
  assign n4910 = ~\u0_w_reg[3][3]/P0001  & n4869 ;
  assign n4911 = ~n4909 & ~n4910 ;
  assign n4912 = n4908 & n4911 ;
  assign n4913 = ~n4908 & ~n4911 ;
  assign n4914 = ~n4912 & ~n4913 ;
  assign n4916 = ~n4905 & n4914 ;
  assign n4915 = n4905 & ~n4914 ;
  assign n4917 = ~\ld_r_reg/P0001  & ~n4915 ;
  assign n4918 = ~n4916 & n4917 ;
  assign n4920 = ~\text_in_r_reg[3]/P0001  & \u0_w_reg[3][3]/P0001  ;
  assign n4919 = \text_in_r_reg[3]/P0001  & ~\u0_w_reg[3][3]/P0001  ;
  assign n4921 = \ld_r_reg/P0001  & ~n4919 ;
  assign n4922 = ~n4920 & n4921 ;
  assign n4923 = ~n4918 & ~n4922 ;
  assign n4924 = ~\u0_w_reg[3][24]/P0001  & ~n3325 ;
  assign n4925 = \u0_w_reg[3][24]/P0001  & n3325 ;
  assign n4926 = ~n4924 & ~n4925 ;
  assign n4927 = ~n2307 & n4773 ;
  assign n4928 = n2307 & ~n4773 ;
  assign n4929 = ~n4927 & ~n4928 ;
  assign n4931 = n4926 & n4929 ;
  assign n4930 = ~n4926 & ~n4929 ;
  assign n4932 = ~\ld_r_reg/P0001  & ~n4930 ;
  assign n4933 = ~n4931 & n4932 ;
  assign n4935 = \text_in_r_reg[24]/P0001  & \u0_w_reg[3][24]/P0001  ;
  assign n4934 = ~\text_in_r_reg[24]/P0001  & ~\u0_w_reg[3][24]/P0001  ;
  assign n4936 = \ld_r_reg/P0001  & ~n4934 ;
  assign n4937 = ~n4935 & n4936 ;
  assign n4938 = ~n4933 & ~n4937 ;
  assign n4939 = n2529 & ~n3416 ;
  assign n4940 = ~n2529 & n3416 ;
  assign n4941 = ~n4939 & ~n4940 ;
  assign n4942 = \u0_w_reg[3][31]/P0001  & ~n2199 ;
  assign n4943 = ~\u0_w_reg[3][31]/P0001  & n2199 ;
  assign n4944 = ~n4942 & ~n4943 ;
  assign n4945 = n4941 & n4944 ;
  assign n4946 = ~n4941 & ~n4944 ;
  assign n4947 = ~n4945 & ~n4946 ;
  assign n4949 = n1741 & ~n4947 ;
  assign n4948 = ~n1741 & n4947 ;
  assign n4950 = ~\ld_r_reg/P0001  & ~n4948 ;
  assign n4951 = ~n4949 & n4950 ;
  assign n4953 = \text_in_r_reg[31]/P0001  & \u0_w_reg[3][31]/P0001  ;
  assign n4952 = ~\text_in_r_reg[31]/P0001  & ~\u0_w_reg[3][31]/P0001  ;
  assign n4954 = \ld_r_reg/P0001  & ~n4952 ;
  assign n4955 = ~n4953 & n4954 ;
  assign n4956 = ~n4951 & ~n4955 ;
  assign n4957 = ~\u0_w_reg[3][16]/P0001  & ~n3325 ;
  assign n4958 = \u0_w_reg[3][16]/P0001  & n3325 ;
  assign n4959 = ~n4957 & ~n4958 ;
  assign n4960 = n2199 & ~n4161 ;
  assign n4961 = ~n2199 & n4161 ;
  assign n4962 = ~n4960 & ~n4961 ;
  assign n4963 = n3595 & n4962 ;
  assign n4964 = ~n3595 & ~n4962 ;
  assign n4965 = ~n4963 & ~n4964 ;
  assign n4967 = n4959 & ~n4965 ;
  assign n4966 = ~n4959 & n4965 ;
  assign n4968 = ~\ld_r_reg/P0001  & ~n4966 ;
  assign n4969 = ~n4967 & n4968 ;
  assign n4971 = \text_in_r_reg[16]/P0001  & \u0_w_reg[3][16]/P0001  ;
  assign n4970 = ~\text_in_r_reg[16]/P0001  & ~\u0_w_reg[3][16]/P0001  ;
  assign n4972 = \ld_r_reg/P0001  & ~n4970 ;
  assign n4973 = ~n4971 & n4972 ;
  assign n4974 = ~n4969 & ~n4973 ;
  assign n4975 = ~n4505 & ~n4596 ;
  assign n4976 = n4505 & n4596 ;
  assign n4977 = ~n4975 & ~n4976 ;
  assign n4978 = \u0_w_reg[3][18]/P0001  & ~n4869 ;
  assign n4979 = ~\u0_w_reg[3][18]/P0001  & n4869 ;
  assign n4980 = ~n4978 & ~n4979 ;
  assign n4981 = n4578 & n4980 ;
  assign n4982 = ~n4578 & ~n4980 ;
  assign n4983 = ~n4981 & ~n4982 ;
  assign n4985 = n4977 & n4983 ;
  assign n4984 = ~n4977 & ~n4983 ;
  assign n4986 = ~\ld_r_reg/P0001  & ~n4984 ;
  assign n4987 = ~n4985 & n4986 ;
  assign n4989 = ~\text_in_r_reg[18]/P0001  & \u0_w_reg[3][18]/P0001  ;
  assign n4988 = \text_in_r_reg[18]/P0001  & ~\u0_w_reg[3][18]/P0001  ;
  assign n4990 = \ld_r_reg/P0001  & ~n4988 ;
  assign n4991 = ~n4989 & n4990 ;
  assign n4992 = ~n4987 & ~n4991 ;
  assign n4993 = ~n2304 & ~n2960 ;
  assign n4994 = n2304 & n2960 ;
  assign n4995 = ~n4993 & ~n4994 ;
  assign n4996 = ~\u0_w_reg[3][23]/P0001  & ~n4941 ;
  assign n4997 = \u0_w_reg[3][23]/P0001  & n4941 ;
  assign n4998 = ~n4996 & ~n4997 ;
  assign n5000 = n4995 & n4998 ;
  assign n4999 = ~n4995 & ~n4998 ;
  assign n5001 = ~\ld_r_reg/P0001  & ~n4999 ;
  assign n5002 = ~n5000 & n5001 ;
  assign n5004 = ~\text_in_r_reg[23]/P0001  & \u0_w_reg[3][23]/P0001  ;
  assign n5003 = \text_in_r_reg[23]/P0001  & ~\u0_w_reg[3][23]/P0001  ;
  assign n5005 = \ld_r_reg/P0001  & ~n5003 ;
  assign n5006 = ~n5004 & n5005 ;
  assign n5007 = ~n5002 & ~n5006 ;
  assign n5008 = ~n4248 & ~n4508 ;
  assign n5009 = n4248 & n4508 ;
  assign n5010 = ~n5008 & ~n5009 ;
  assign n5011 = \u0_w_reg[3][10]/P0001  & ~n4869 ;
  assign n5012 = ~\u0_w_reg[3][10]/P0001  & n4869 ;
  assign n5013 = ~n5011 & ~n5012 ;
  assign n5014 = n3503 & n5013 ;
  assign n5015 = ~n3503 & ~n5013 ;
  assign n5016 = ~n5014 & ~n5015 ;
  assign n5018 = n5010 & n5016 ;
  assign n5017 = ~n5010 & ~n5016 ;
  assign n5019 = ~\ld_r_reg/P0001  & ~n5017 ;
  assign n5020 = ~n5018 & n5019 ;
  assign n5022 = ~\text_in_r_reg[10]/P0001  & \u0_w_reg[3][10]/P0001  ;
  assign n5021 = \text_in_r_reg[10]/P0001  & ~\u0_w_reg[3][10]/P0001  ;
  assign n5023 = \ld_r_reg/P0001  & ~n5021 ;
  assign n5024 = ~n5022 & n5023 ;
  assign n5025 = ~n5020 & ~n5024 ;
  assign n5026 = ~\u0_w_reg[3][8]/P0001  & ~n3325 ;
  assign n5027 = \u0_w_reg[3][8]/P0001  & n3325 ;
  assign n5028 = ~n5026 & ~n5027 ;
  assign n5029 = n4677 & ~n4941 ;
  assign n5030 = ~n4677 & n4941 ;
  assign n5031 = ~n5029 & ~n5030 ;
  assign n5033 = n5028 & ~n5031 ;
  assign n5032 = ~n5028 & n5031 ;
  assign n5034 = ~\ld_r_reg/P0001  & ~n5032 ;
  assign n5035 = ~n5033 & n5034 ;
  assign n5037 = ~\text_in_r_reg[8]/P0001  & \u0_w_reg[3][8]/P0001  ;
  assign n5036 = \text_in_r_reg[8]/P0001  & ~\u0_w_reg[3][8]/P0001  ;
  assign n5038 = \ld_r_reg/P0001  & ~n5036 ;
  assign n5039 = ~n5037 & n5038 ;
  assign n5040 = ~n5035 & ~n5039 ;
  assign n5041 = ~\u0_w_reg[3][0]/P0001  & ~n3416 ;
  assign n5042 = \u0_w_reg[3][0]/P0001  & n3416 ;
  assign n5043 = ~n5041 & ~n5042 ;
  assign n5044 = n4164 & n4773 ;
  assign n5045 = ~n4164 & ~n4773 ;
  assign n5046 = ~n5044 & ~n5045 ;
  assign n5048 = n5043 & n5046 ;
  assign n5047 = ~n5043 & ~n5046 ;
  assign n5049 = ~\ld_r_reg/P0001  & ~n5047 ;
  assign n5050 = ~n5048 & n5049 ;
  assign n5052 = \text_in_r_reg[0]/P0001  & \u0_w_reg[3][0]/P0001  ;
  assign n5051 = ~\text_in_r_reg[0]/P0001  & ~\u0_w_reg[3][0]/P0001  ;
  assign n5053 = \ld_r_reg/P0001  & ~n5051 ;
  assign n5054 = ~n5052 & n5053 ;
  assign n5055 = ~n5050 & ~n5054 ;
  assign n5056 = ~\u0_w_reg[3][5]/P0001  & ~n2077 ;
  assign n5057 = \u0_w_reg[3][5]/P0001  & n2077 ;
  assign n5058 = ~n5056 & ~n5057 ;
  assign n5059 = ~\u0_w_reg[3][6]/P0001  & ~n2416 ;
  assign n5060 = \u0_w_reg[3][6]/P0001  & n2416 ;
  assign n5061 = ~n5059 & ~n5060 ;
  assign n5062 = ~\u0_w_reg[3][4]/P0001  & ~n3205 ;
  assign n5063 = \u0_w_reg[3][4]/P0001  & n3205 ;
  assign n5064 = ~n5062 & ~n5063 ;
  assign n5065 = ~\u0_w_reg[3][0]/P0001  & ~n3325 ;
  assign n5066 = \u0_w_reg[3][0]/P0001  & n3325 ;
  assign n5067 = ~n5065 & ~n5066 ;
  assign n5068 = ~\u0_w_reg[3][3]/P0001  & ~n4338 ;
  assign n5069 = \u0_w_reg[3][3]/P0001  & n4338 ;
  assign n5070 = ~n5068 & ~n5069 ;
  assign n5071 = ~\u0_w_reg[3][1]/P0001  & ~n3503 ;
  assign n5072 = \u0_w_reg[3][1]/P0001  & n3503 ;
  assign n5073 = ~n5071 & ~n5072 ;
  assign n5074 = ~\u0_w_reg[3][2]/P0001  & ~n4869 ;
  assign n5075 = \u0_w_reg[3][2]/P0001  & n4869 ;
  assign n5076 = ~n5074 & ~n5075 ;
  assign n5077 = ~\u0_w_reg[3][7]/P0001  & ~n3416 ;
  assign n5078 = \u0_w_reg[3][7]/P0001  & n3416 ;
  assign n5079 = ~n5077 & ~n5078 ;
  assign n5091 = \sa02_reg[5]/P0001  & n979 ;
  assign n5092 = ~\sa02_reg[3]/P0001  & n5091 ;
  assign n5093 = n1009 & ~n5092 ;
  assign n5094 = ~\sa02_reg[2]/P0001  & ~n5093 ;
  assign n5095 = ~n1001 & ~n5094 ;
  assign n5096 = ~\sa02_reg[1]/P0001  & ~n5095 ;
  assign n5083 = ~\sa02_reg[3]/P0001  & n1090 ;
  assign n5084 = \sa02_reg[7]/NET0131  & n5083 ;
  assign n5082 = \sa02_reg[4]/P0001  & n1025 ;
  assign n5085 = ~n1043 & ~n5082 ;
  assign n5086 = ~n5084 & n5085 ;
  assign n5087 = \sa02_reg[1]/P0001  & ~n5086 ;
  assign n5080 = ~n1071 & ~n1123 ;
  assign n5081 = n982 & n1015 ;
  assign n5088 = n5080 & ~n5081 ;
  assign n5089 = ~n5087 & n5088 ;
  assign n5090 = \sa02_reg[2]/P0001  & ~n5089 ;
  assign n5102 = n993 & n1059 ;
  assign n5103 = ~n1058 & ~n5102 ;
  assign n5104 = \sa02_reg[1]/P0001  & ~n5103 ;
  assign n5105 = ~n1039 & ~n1130 ;
  assign n5106 = ~\sa02_reg[1]/P0001  & \sa02_reg[2]/P0001  ;
  assign n5107 = ~n5105 & n5106 ;
  assign n5099 = n975 & n1015 ;
  assign n5100 = ~n1022 & ~n5099 ;
  assign n5101 = ~\sa02_reg[2]/P0001  & ~n5100 ;
  assign n5097 = \sa02_reg[2]/P0001  & ~\sa02_reg[5]/P0001  ;
  assign n5098 = n1024 & n5097 ;
  assign n5108 = ~\sa02_reg[2]/P0001  & ~\sa02_reg[3]/P0001  ;
  assign n5109 = \sa02_reg[1]/P0001  & ~\sa02_reg[5]/P0001  ;
  assign n5110 = ~n1004 & n5109 ;
  assign n5111 = n5108 & n5110 ;
  assign n5112 = ~n5098 & ~n5111 ;
  assign n5113 = ~n5101 & n5112 ;
  assign n5114 = ~n5107 & n5113 ;
  assign n5115 = ~n5104 & n5114 ;
  assign n5116 = ~n5090 & n5115 ;
  assign n5117 = ~n5096 & n5116 ;
  assign n5118 = \sa02_reg[0]/P0001  & ~n5117 ;
  assign n5121 = n978 & ~n997 ;
  assign n5119 = ~\sa02_reg[2]/P0001  & n980 ;
  assign n5120 = ~\sa02_reg[4]/P0001  & n5119 ;
  assign n5122 = \sa02_reg[6]/NET0131  & n1057 ;
  assign n5123 = \sa02_reg[1]/P0001  & ~n5122 ;
  assign n5124 = ~n5120 & n5123 ;
  assign n5125 = ~n5121 & n5124 ;
  assign n5126 = \sa02_reg[4]/P0001  & n1021 ;
  assign n5132 = n1000 & n1095 ;
  assign n5129 = n974 & n1023 ;
  assign n5130 = ~\sa02_reg[4]/P0001  & \sa02_reg[7]/NET0131  ;
  assign n5131 = n1035 & n5130 ;
  assign n5134 = ~n5129 & ~n5131 ;
  assign n5135 = ~n5132 & n5134 ;
  assign n5127 = \sa02_reg[3]/P0001  & n1056 ;
  assign n5128 = n1016 & n5127 ;
  assign n5133 = ~\sa02_reg[1]/P0001  & ~n5099 ;
  assign n5136 = ~n5128 & n5133 ;
  assign n5137 = n5135 & n5136 ;
  assign n5138 = ~n5126 & n5137 ;
  assign n5139 = ~n5125 & ~n5138 ;
  assign n5142 = ~n979 & n1035 ;
  assign n5143 = \sa02_reg[4]/P0001  & ~n1019 ;
  assign n5144 = n5142 & ~n5143 ;
  assign n5140 = n975 & n986 ;
  assign n5141 = ~\sa02_reg[7]/NET0131  & n5140 ;
  assign n5145 = ~\sa02_reg[2]/P0001  & ~n987 ;
  assign n5146 = ~n5141 & n5145 ;
  assign n5147 = ~n5144 & n5146 ;
  assign n5148 = n974 & n982 ;
  assign n5149 = \sa02_reg[2]/P0001  & ~n5148 ;
  assign n5150 = ~n5126 & n5149 ;
  assign n5151 = ~n5147 & ~n5150 ;
  assign n5152 = ~n5139 & ~n5151 ;
  assign n5153 = ~\sa02_reg[0]/P0001  & ~n5152 ;
  assign n5163 = \sa02_reg[6]/NET0131  & n1007 ;
  assign n5156 = ~\sa02_reg[6]/NET0131  & n1030 ;
  assign n5164 = ~n1001 & ~n5156 ;
  assign n5165 = ~n5163 & n5164 ;
  assign n5166 = ~\sa02_reg[2]/P0001  & ~n5165 ;
  assign n5172 = n993 & n1004 ;
  assign n5173 = \sa02_reg[2]/P0001  & n5172 ;
  assign n5168 = \sa02_reg[2]/P0001  & ~\sa02_reg[4]/P0001  ;
  assign n5169 = n979 & n5168 ;
  assign n5170 = \sa02_reg[3]/P0001  & n5169 ;
  assign n5167 = n1023 & n1038 ;
  assign n5171 = n974 & n975 ;
  assign n5174 = ~n5167 & ~n5171 ;
  assign n5175 = ~n5170 & n5174 ;
  assign n5176 = ~n5173 & n5175 ;
  assign n5177 = ~n5166 & n5176 ;
  assign n5178 = ~\sa02_reg[1]/P0001  & ~n5177 ;
  assign n5154 = \sa02_reg[1]/P0001  & \sa02_reg[2]/P0001  ;
  assign n5155 = ~\sa02_reg[3]/P0001  & n979 ;
  assign n5157 = ~n5155 & ~n5156 ;
  assign n5158 = ~\sa02_reg[4]/P0001  & ~n5157 ;
  assign n5159 = \sa02_reg[4]/P0001  & ~\sa02_reg[6]/NET0131  ;
  assign n5160 = n995 & n5159 ;
  assign n5161 = ~n5158 & ~n5160 ;
  assign n5162 = n5154 & ~n5161 ;
  assign n5182 = n1001 & n1095 ;
  assign n5181 = ~\sa02_reg[7]/NET0131  & n5148 ;
  assign n5184 = ~n981 & ~n5181 ;
  assign n5185 = ~n5182 & n5184 ;
  assign n5179 = \sa02_reg[1]/P0001  & ~\sa02_reg[2]/P0001  ;
  assign n5180 = n1110 & n5179 ;
  assign n5183 = n984 & n5163 ;
  assign n5186 = ~n5180 & ~n5183 ;
  assign n5187 = n5185 & n5186 ;
  assign n5188 = ~n5162 & n5187 ;
  assign n5189 = ~n5178 & n5188 ;
  assign n5190 = ~n5153 & n5189 ;
  assign n5191 = ~n5118 & n5190 ;
  assign n5192 = n689 & ~n5191 ;
  assign n5193 = ~n689 & n5191 ;
  assign n5194 = ~n5192 & ~n5193 ;
  assign n5195 = ~n1142 & ~n5194 ;
  assign n5196 = n1142 & n5194 ;
  assign n5197 = ~n5195 & ~n5196 ;
  assign n5198 = \sa31_reg[4]/P0001  & n1178 ;
  assign n5199 = ~\sa31_reg[4]/P0001  & n1149 ;
  assign n5200 = ~n5198 & ~n5199 ;
  assign n5201 = ~\sa31_reg[3]/P0001  & ~n5200 ;
  assign n5202 = ~n1206 & ~n5201 ;
  assign n5203 = ~\sa31_reg[2]/P0001  & ~n5202 ;
  assign n5209 = \sa31_reg[4]/P0001  & n1194 ;
  assign n5210 = ~n1167 & ~n5209 ;
  assign n5211 = \sa31_reg[2]/P0001  & ~n5210 ;
  assign n5204 = n1186 & n1216 ;
  assign n5212 = ~n1148 & ~n5204 ;
  assign n5208 = \sa31_reg[4]/P0001  & n1167 ;
  assign n5205 = ~\sa31_reg[5]/P0001  & n1256 ;
  assign n5206 = ~\sa31_reg[3]/P0001  & n5205 ;
  assign n5207 = n1152 & n1194 ;
  assign n5213 = ~n5206 & ~n5207 ;
  assign n5214 = ~n5208 & n5213 ;
  assign n5215 = n5212 & n5214 ;
  assign n5216 = ~n5211 & n5215 ;
  assign n5217 = ~n5203 & n5216 ;
  assign n5218 = \sa31_reg[1]/P0001  & ~n5217 ;
  assign n5225 = ~n1247 & ~n1255 ;
  assign n5226 = \sa31_reg[7]/P0001  & ~n5225 ;
  assign n5227 = n1229 & n1248 ;
  assign n5228 = ~n1221 & ~n5227 ;
  assign n5229 = ~n5226 & n5228 ;
  assign n5230 = ~\sa31_reg[1]/P0001  & ~n5229 ;
  assign n5221 = ~\sa31_reg[3]/P0001  & n1239 ;
  assign n5219 = \sa31_reg[3]/P0001  & ~n1281 ;
  assign n5220 = ~\sa31_reg[4]/P0001  & n1186 ;
  assign n5222 = ~n5219 & ~n5220 ;
  assign n5223 = ~n5221 & n5222 ;
  assign n5224 = \sa31_reg[2]/P0001  & ~n5223 ;
  assign n5231 = ~\sa31_reg[2]/P0001  & n1179 ;
  assign n5232 = ~n1205 & ~n5231 ;
  assign n5233 = ~n1185 & n5232 ;
  assign n5234 = ~n5224 & n5233 ;
  assign n5235 = ~n5230 & n5234 ;
  assign n5236 = ~n5218 & n5235 ;
  assign n5237 = ~\sa31_reg[0]/P0002  & ~n5236 ;
  assign n5263 = \sa31_reg[5]/P0001  & n1225 ;
  assign n5265 = n1164 & ~n1174 ;
  assign n5266 = ~n5263 & ~n5265 ;
  assign n5267 = \sa31_reg[1]/P0001  & ~n5266 ;
  assign n5268 = ~\sa31_reg[4]/P0001  & n1158 ;
  assign n5269 = \sa31_reg[3]/P0001  & \sa31_reg[6]/NET0131  ;
  assign n5270 = n1158 & n5269 ;
  assign n5271 = n1149 & n1225 ;
  assign n5272 = ~n5270 & ~n5271 ;
  assign n5273 = ~n5268 & n5272 ;
  assign n5274 = ~n5267 & n5273 ;
  assign n5275 = ~\sa31_reg[2]/P0001  & ~n5274 ;
  assign n5241 = ~\sa31_reg[4]/P0001  & n1151 ;
  assign n5242 = n1159 & n1186 ;
  assign n5243 = ~n5241 & ~n5242 ;
  assign n5244 = \sa31_reg[2]/P0001  & ~n5243 ;
  assign n5245 = n1194 & ~n1279 ;
  assign n5238 = ~\sa31_reg[2]/P0001  & \sa31_reg[3]/P0001  ;
  assign n5239 = ~\sa31_reg[5]/P0001  & n1146 ;
  assign n5240 = n5238 & n5239 ;
  assign n5246 = ~n1202 & ~n5240 ;
  assign n5247 = ~n5245 & n5246 ;
  assign n5248 = ~n5244 & n5247 ;
  assign n5249 = ~\sa31_reg[1]/P0001  & ~n5248 ;
  assign n5250 = \sa31_reg[7]/P0001  & n1197 ;
  assign n5251 = ~n1161 & ~n5250 ;
  assign n5252 = ~\sa31_reg[7]/P0001  & n1196 ;
  assign n5253 = n1229 & n5252 ;
  assign n5254 = ~\sa31_reg[4]/P0001  & n1206 ;
  assign n5255 = ~n5253 & ~n5254 ;
  assign n5256 = n5251 & n5255 ;
  assign n5257 = \sa31_reg[1]/P0001  & ~n5256 ;
  assign n5258 = n1151 & n1230 ;
  assign n5259 = ~n1202 & ~n5258 ;
  assign n5260 = \sa31_reg[2]/P0001  & ~n5259 ;
  assign n5261 = n1151 & n1174 ;
  assign n5262 = ~\sa31_reg[2]/P0001  & n5261 ;
  assign n5264 = n1149 & n5263 ;
  assign n5276 = ~n5262 & ~n5264 ;
  assign n5277 = ~n5260 & n5276 ;
  assign n5278 = ~n5257 & n5277 ;
  assign n5279 = ~n5249 & n5278 ;
  assign n5280 = ~n5275 & n5279 ;
  assign n5281 = \sa31_reg[0]/P0002  & ~n5280 ;
  assign n5282 = ~n1153 & ~n1200 ;
  assign n5283 = \sa31_reg[5]/P0001  & ~n5282 ;
  assign n5284 = ~n5261 & ~n5283 ;
  assign n5285 = ~\sa31_reg[2]/P0001  & ~n5284 ;
  assign n5287 = ~n1173 & ~n5239 ;
  assign n5288 = ~\sa31_reg[3]/P0001  & ~n1201 ;
  assign n5289 = n5287 & n5288 ;
  assign n5286 = \sa31_reg[3]/P0001  & ~n1178 ;
  assign n5290 = n1215 & ~n5286 ;
  assign n5291 = ~n5289 & n5290 ;
  assign n5292 = ~n1234 & ~n5291 ;
  assign n5293 = ~n5285 & n5292 ;
  assign n5294 = ~\sa31_reg[1]/P0001  & ~n5293 ;
  assign n5298 = \sa31_reg[2]/P0001  & n1261 ;
  assign n5299 = ~\sa31_reg[4]/P0001  & n5204 ;
  assign n5300 = ~n5231 & ~n5299 ;
  assign n5301 = ~n5298 & n5300 ;
  assign n5302 = \sa31_reg[1]/P0001  & ~n5301 ;
  assign n5295 = \sa31_reg[4]/P0001  & n1266 ;
  assign n5296 = ~n1227 & ~n5206 ;
  assign n5297 = ~\sa31_reg[2]/P0001  & ~n5296 ;
  assign n5303 = ~n5295 & ~n5297 ;
  assign n5304 = ~n5302 & n5303 ;
  assign n5305 = ~n5294 & n5304 ;
  assign n5306 = ~n5281 & n5305 ;
  assign n5307 = ~n5237 & n5306 ;
  assign n5308 = \u0_w_reg[2][6]/P0001  & ~n5307 ;
  assign n5309 = ~\u0_w_reg[2][6]/P0001  & n5307 ;
  assign n5310 = ~n5308 & ~n5309 ;
  assign n5311 = n850 & n5310 ;
  assign n5312 = ~n850 & ~n5310 ;
  assign n5313 = ~n5311 & ~n5312 ;
  assign n5315 = n5197 & ~n5313 ;
  assign n5314 = ~n5197 & n5313 ;
  assign n5316 = ~\ld_r_reg/P0001  & ~n5314 ;
  assign n5317 = ~n5315 & n5316 ;
  assign n5319 = \text_in_r_reg[38]/P0001  & \u0_w_reg[2][6]/P0001  ;
  assign n5318 = ~\text_in_r_reg[38]/P0001  & ~\u0_w_reg[2][6]/P0001  ;
  assign n5320 = \ld_r_reg/P0001  & ~n5318 ;
  assign n5321 = ~n5319 & n5320 ;
  assign n5322 = ~n5317 & ~n5321 ;
  assign n5389 = ~n1072 & ~n5172 ;
  assign n5390 = n999 & ~n5130 ;
  assign n5391 = n5389 & ~n5390 ;
  assign n5392 = n1095 & ~n5391 ;
  assign n5323 = \sa02_reg[4]/P0001  & n982 ;
  assign n5324 = ~n1004 & ~n5323 ;
  assign n5393 = \sa02_reg[7]/NET0131  & ~n5324 ;
  assign n5394 = ~\sa02_reg[6]/NET0131  & n1084 ;
  assign n5395 = ~n5393 & ~n5394 ;
  assign n5396 = ~\sa02_reg[3]/P0001  & ~n5395 ;
  assign n5397 = ~n1005 & ~n1082 ;
  assign n5398 = ~n5396 & n5397 ;
  assign n5399 = \sa02_reg[2]/P0001  & ~n5398 ;
  assign n5400 = ~n5392 & ~n5399 ;
  assign n5401 = \sa02_reg[1]/P0001  & ~n5400 ;
  assign n5348 = \sa02_reg[4]/P0001  & ~n999 ;
  assign n5349 = ~\sa02_reg[2]/P0001  & ~n1020 ;
  assign n5350 = n5348 & n5349 ;
  assign n5344 = \sa02_reg[2]/P0001  & ~n986 ;
  assign n5345 = n1025 & ~n1035 ;
  assign n5346 = ~n5344 & n5345 ;
  assign n5342 = \sa02_reg[2]/P0001  & n974 ;
  assign n5343 = n1003 & n5342 ;
  assign n5347 = n999 & n1059 ;
  assign n5351 = ~n5343 & ~n5347 ;
  assign n5352 = ~n5346 & n5351 ;
  assign n5353 = ~n5350 & n5352 ;
  assign n5354 = ~\sa02_reg[1]/P0001  & ~n5353 ;
  assign n5325 = \sa02_reg[3]/P0001  & n1025 ;
  assign n5326 = ~n5155 & ~n5325 ;
  assign n5327 = n5324 & n5326 ;
  assign n5328 = \sa02_reg[1]/P0001  & ~n5327 ;
  assign n5329 = n974 & n1019 ;
  assign n5330 = ~n1022 & ~n1031 ;
  assign n5331 = ~n5329 & n5330 ;
  assign n5332 = ~n5328 & n5331 ;
  assign n5333 = \sa02_reg[2]/P0001  & ~n5332 ;
  assign n5338 = n1011 & n1039 ;
  assign n5339 = n1094 & n5108 ;
  assign n5340 = ~n5338 & ~n5339 ;
  assign n5341 = \sa02_reg[1]/P0001  & ~n5340 ;
  assign n5335 = ~\sa02_reg[2]/P0001  & n1025 ;
  assign n5336 = ~n1056 & ~n5335 ;
  assign n5337 = n986 & ~n5336 ;
  assign n5334 = n984 & n1090 ;
  assign n5355 = \sa02_reg[0]/P0001  & ~n5334 ;
  assign n5356 = ~n5337 & n5355 ;
  assign n5357 = ~n5341 & n5356 ;
  assign n5358 = ~n5333 & n5357 ;
  assign n5359 = ~n5354 & n5358 ;
  assign n5370 = ~n979 & ~n1039 ;
  assign n5371 = n5097 & ~n5370 ;
  assign n5372 = ~\sa02_reg[2]/P0001  & n5130 ;
  assign n5373 = ~\sa02_reg[1]/P0001  & ~n5102 ;
  assign n5374 = ~n5372 & n5373 ;
  assign n5375 = ~n5371 & n5374 ;
  assign n5378 = \sa02_reg[1]/P0001  & ~n1013 ;
  assign n5379 = ~n5156 & n5378 ;
  assign n5376 = ~n1130 & ~n5159 ;
  assign n5377 = n1095 & ~n5376 ;
  assign n5380 = ~n5126 & ~n5377 ;
  assign n5381 = n5379 & n5380 ;
  assign n5382 = ~n5375 & ~n5381 ;
  assign n5360 = ~n5122 & ~n5160 ;
  assign n5361 = ~\sa02_reg[2]/P0001  & ~n5360 ;
  assign n5363 = n1056 & n5159 ;
  assign n5364 = n975 & n1000 ;
  assign n5365 = ~n5363 & ~n5364 ;
  assign n5366 = n984 & ~n5365 ;
  assign n5362 = n1037 & n5168 ;
  assign n5367 = \sa02_reg[5]/P0001  & ~n1023 ;
  assign n5368 = ~n1006 & n5108 ;
  assign n5369 = n5367 & n5368 ;
  assign n5383 = ~\sa02_reg[0]/P0001  & ~n5369 ;
  assign n5384 = ~n5362 & n5383 ;
  assign n5385 = ~n5366 & n5384 ;
  assign n5386 = ~n5361 & n5385 ;
  assign n5387 = ~n5382 & n5386 ;
  assign n5388 = ~n5359 & ~n5387 ;
  assign n5402 = ~\sa02_reg[7]/NET0131  & n5171 ;
  assign n5403 = ~\sa02_reg[5]/P0001  & n1091 ;
  assign n5404 = ~n5402 & ~n5403 ;
  assign n5405 = ~\sa02_reg[2]/P0001  & ~n5404 ;
  assign n5406 = ~n1037 & ~n5140 ;
  assign n5407 = ~n5338 & n5406 ;
  assign n5408 = \sa02_reg[2]/P0001  & ~n5407 ;
  assign n5410 = n1035 & n5372 ;
  assign n5409 = n986 & n993 ;
  assign n5411 = ~n5369 & ~n5409 ;
  assign n5412 = ~n5410 & n5411 ;
  assign n5413 = ~n5408 & n5412 ;
  assign n5414 = ~\sa02_reg[1]/P0001  & ~n5413 ;
  assign n5415 = ~n5405 & ~n5414 ;
  assign n5416 = ~n5388 & n5415 ;
  assign n5417 = ~n5401 & n5416 ;
  assign n5487 = ~n888 & ~n908 ;
  assign n5458 = ~\sa13_reg[4]/P0001  & \sa13_reg[7]/NET0131  ;
  assign n5488 = n532 & ~n5458 ;
  assign n5489 = n5487 & ~n5488 ;
  assign n5490 = n581 & ~n5489 ;
  assign n5441 = ~n563 & ~n632 ;
  assign n5491 = \sa13_reg[7]/NET0131  & ~n5441 ;
  assign n5492 = ~\sa13_reg[6]/NET0131  & n901 ;
  assign n5493 = ~n5491 & ~n5492 ;
  assign n5494 = ~\sa13_reg[3]/P0001  & ~n5493 ;
  assign n5495 = ~n571 & ~n902 ;
  assign n5496 = ~n5494 & n5495 ;
  assign n5497 = \sa13_reg[2]/P0001  & ~n5496 ;
  assign n5498 = ~n5490 & ~n5497 ;
  assign n5499 = \sa13_reg[1]/P0001  & ~n5498 ;
  assign n5442 = ~\sa13_reg[3]/P0001  & n556 ;
  assign n5443 = ~n544 & ~n5442 ;
  assign n5444 = n5441 & n5443 ;
  assign n5445 = \sa13_reg[2]/P0001  & ~n5444 ;
  assign n5440 = \sa13_reg[3]/P0001  & n913 ;
  assign n5446 = n549 & n565 ;
  assign n5447 = ~n5440 & ~n5446 ;
  assign n5448 = ~n5445 & n5447 ;
  assign n5449 = \sa13_reg[1]/P0001  & ~n5448 ;
  assign n5418 = \sa13_reg[4]/P0001  & ~n532 ;
  assign n5419 = ~n855 & n5418 ;
  assign n5420 = ~n861 & ~n5419 ;
  assign n5421 = ~\sa13_reg[2]/P0001  & ~n5420 ;
  assign n5426 = n570 & n653 ;
  assign n5427 = \sa13_reg[2]/P0001  & n5426 ;
  assign n5422 = ~\sa13_reg[7]/NET0131  & n620 ;
  assign n5423 = n532 & n655 ;
  assign n5424 = ~\sa13_reg[2]/P0001  & ~\sa13_reg[3]/P0001  ;
  assign n5425 = n543 & n5424 ;
  assign n5428 = ~n5423 & ~n5425 ;
  assign n5429 = ~n5422 & n5428 ;
  assign n5430 = ~n5427 & n5429 ;
  assign n5431 = ~n5421 & n5430 ;
  assign n5432 = ~\sa13_reg[1]/P0001  & ~n5431 ;
  assign n5434 = ~\sa13_reg[3]/P0001  & n584 ;
  assign n5435 = ~n534 & ~n858 ;
  assign n5436 = ~n5434 & n5435 ;
  assign n5437 = \sa13_reg[2]/P0001  & ~n5436 ;
  assign n5433 = ~\sa13_reg[2]/P0001  & n5422 ;
  assign n5439 = n623 & n928 ;
  assign n5438 = n533 & n900 ;
  assign n5450 = \sa13_reg[0]/P0001  & ~n5438 ;
  assign n5451 = ~n5439 & n5450 ;
  assign n5452 = ~n5433 & n5451 ;
  assign n5453 = ~n5437 & n5452 ;
  assign n5454 = ~n5432 & n5453 ;
  assign n5455 = ~n5449 & n5454 ;
  assign n5474 = ~n648 & ~n946 ;
  assign n5475 = ~\sa13_reg[2]/P0001  & ~n5474 ;
  assign n5473 = ~n611 & n621 ;
  assign n5476 = \sa13_reg[5]/P0001  & n864 ;
  assign n5477 = ~n5473 & ~n5476 ;
  assign n5478 = ~n5475 & n5477 ;
  assign n5479 = \sa13_reg[1]/P0001  & ~n5478 ;
  assign n5459 = ~\sa13_reg[2]/P0001  & n5458 ;
  assign n5460 = ~n561 & ~n5459 ;
  assign n5456 = \sa13_reg[4]/P0001  & n570 ;
  assign n5457 = n623 & n5456 ;
  assign n5461 = ~n887 & ~n5457 ;
  assign n5462 = n5460 & n5461 ;
  assign n5463 = ~\sa13_reg[1]/P0001  & ~n5462 ;
  assign n5469 = ~n540 & ~n901 ;
  assign n5470 = n5424 & ~n5469 ;
  assign n5464 = n604 & n623 ;
  assign n5465 = ~\sa13_reg[6]/NET0131  & n5464 ;
  assign n5480 = ~\sa13_reg[0]/P0001  & ~n5465 ;
  assign n5481 = ~n5470 & n5480 ;
  assign n5466 = \sa13_reg[4]/P0001  & n557 ;
  assign n5467 = ~n907 & ~n5466 ;
  assign n5468 = n623 & ~n5467 ;
  assign n5471 = ~n609 & ~n652 ;
  assign n5472 = ~\sa13_reg[2]/P0001  & ~n5471 ;
  assign n5482 = ~n5468 & ~n5472 ;
  assign n5483 = n5481 & n5482 ;
  assign n5484 = ~n5463 & n5483 ;
  assign n5485 = ~n5479 & n5484 ;
  assign n5486 = ~n5455 & ~n5485 ;
  assign n5500 = n579 & n946 ;
  assign n5501 = ~n863 & ~n5500 ;
  assign n5502 = ~\sa13_reg[2]/P0001  & ~n5501 ;
  assign n5505 = \sa13_reg[4]/P0001  & n535 ;
  assign n5506 = ~\sa13_reg[3]/P0001  & n5505 ;
  assign n5507 = ~n854 & ~n5440 ;
  assign n5508 = ~n5506 & n5507 ;
  assign n5509 = \sa13_reg[2]/P0001  & ~n5508 ;
  assign n5503 = n550 & n5459 ;
  assign n5504 = n533 & n559 ;
  assign n5510 = ~n5503 & ~n5504 ;
  assign n5511 = ~n5470 & n5510 ;
  assign n5512 = ~n5509 & n5511 ;
  assign n5513 = ~\sa13_reg[1]/P0001  & ~n5512 ;
  assign n5514 = ~n5502 & ~n5513 ;
  assign n5515 = ~n5486 & n5514 ;
  assign n5516 = ~n5499 & n5515 ;
  assign n5517 = n5417 & ~n5516 ;
  assign n5518 = ~n5417 & n5516 ;
  assign n5519 = ~n5517 & ~n5518 ;
  assign n5520 = ~n5191 & ~n5519 ;
  assign n5521 = n5191 & n5519 ;
  assign n5522 = ~n5520 & ~n5521 ;
  assign n5567 = n717 & n719 ;
  assign n5568 = ~n827 & ~n5567 ;
  assign n5569 = n690 & ~n765 ;
  assign n5570 = n5568 & ~n5569 ;
  assign n5571 = n763 & ~n5570 ;
  assign n5551 = ~n719 & ~n791 ;
  assign n5572 = \sa20_reg[7]/NET0131  & ~n5551 ;
  assign n5573 = n694 & n723 ;
  assign n5574 = ~n5572 & ~n5573 ;
  assign n5575 = ~\sa20_reg[3]/P0001  & ~n5574 ;
  assign n5576 = ~n721 & ~n778 ;
  assign n5577 = ~n5575 & n5576 ;
  assign n5578 = \sa20_reg[2]/P0001  & ~n5577 ;
  assign n5579 = ~n5571 & ~n5578 ;
  assign n5580 = \sa20_reg[1]/P0001  & ~n5579 ;
  assign n5552 = ~\sa20_reg[3]/P0001  & n723 ;
  assign n5553 = ~n699 & ~n5552 ;
  assign n5554 = n5551 & n5553 ;
  assign n5555 = \sa20_reg[1]/P0001  & ~n5554 ;
  assign n5556 = \sa20_reg[5]/P0001  & n739 ;
  assign n5550 = n719 & n736 ;
  assign n5557 = ~n692 & ~n5550 ;
  assign n5558 = ~n5556 & n5557 ;
  assign n5559 = ~n5555 & n5558 ;
  assign n5560 = \sa20_reg[2]/P0001  & ~n5559 ;
  assign n5529 = ~\sa20_reg[4]/P0001  & n720 ;
  assign n5530 = ~\sa20_reg[3]/P0001  & n5529 ;
  assign n5531 = \sa20_reg[2]/P0001  & ~n5530 ;
  assign n5533 = ~\sa20_reg[2]/P0001  & ~n739 ;
  assign n5532 = \sa20_reg[4]/P0001  & n701 ;
  assign n5534 = ~n791 & ~n5532 ;
  assign n5535 = n5533 & n5534 ;
  assign n5536 = ~n5531 & ~n5535 ;
  assign n5526 = \sa20_reg[2]/P0001  & ~\sa20_reg[4]/P0001  ;
  assign n5527 = ~\sa20_reg[3]/P0001  & n693 ;
  assign n5528 = ~n5526 & n5527 ;
  assign n5523 = ~\sa20_reg[2]/P0001  & \sa20_reg[6]/NET0131  ;
  assign n5524 = n777 & n5523 ;
  assign n5525 = n690 & n745 ;
  assign n5537 = ~n5524 & ~n5525 ;
  assign n5538 = ~n5528 & n5537 ;
  assign n5539 = ~n5536 & n5538 ;
  assign n5540 = ~\sa20_reg[1]/P0001  & ~n5539 ;
  assign n5543 = \sa20_reg[4]/P0001  & n795 ;
  assign n5544 = ~\sa20_reg[5]/P0001  & n705 ;
  assign n5545 = n747 & n5544 ;
  assign n5546 = ~n5543 & ~n5545 ;
  assign n5547 = \sa20_reg[1]/P0001  & ~n5546 ;
  assign n5548 = n739 & n747 ;
  assign n5541 = n735 & n5526 ;
  assign n5542 = \sa20_reg[3]/P0001  & n5541 ;
  assign n5549 = n691 & n777 ;
  assign n5561 = ~n5542 & ~n5549 ;
  assign n5562 = ~n5548 & n5561 ;
  assign n5563 = ~n5547 & n5562 ;
  assign n5564 = ~n5540 & n5563 ;
  assign n5565 = ~n5560 & n5564 ;
  assign n5566 = \sa20_reg[0]/P0001  & ~n5565 ;
  assign n5582 = ~\sa20_reg[2]/P0001  & ~\sa20_reg[4]/P0001  ;
  assign n5583 = ~n810 & ~n5582 ;
  assign n5584 = \sa20_reg[7]/NET0131  & ~n5583 ;
  assign n5585 = \sa20_reg[4]/P0001  & n720 ;
  assign n5586 = n761 & n5585 ;
  assign n5581 = \sa20_reg[2]/P0001  & n820 ;
  assign n5587 = ~\sa20_reg[1]/P0001  & ~n5581 ;
  assign n5588 = ~n5586 & n5587 ;
  assign n5589 = ~n5584 & n5588 ;
  assign n5591 = n693 & n706 ;
  assign n5592 = ~n750 & ~n5591 ;
  assign n5593 = ~\sa20_reg[2]/P0001  & ~n5592 ;
  assign n5590 = \sa20_reg[1]/P0001  & ~n834 ;
  assign n5594 = ~n736 & ~n819 ;
  assign n5595 = n767 & ~n5594 ;
  assign n5596 = n5590 & ~n5595 ;
  assign n5597 = ~n5593 & n5596 ;
  assign n5598 = ~n5589 & ~n5597 ;
  assign n5599 = n701 & n736 ;
  assign n5600 = n777 & n799 ;
  assign n5601 = ~n5599 & ~n5600 ;
  assign n5602 = ~n779 & ~n808 ;
  assign n5603 = n5601 & n5602 ;
  assign n5604 = ~\sa20_reg[2]/P0001  & ~n5603 ;
  assign n5606 = \sa20_reg[4]/P0001  & n724 ;
  assign n5605 = n701 & n714 ;
  assign n5607 = ~n710 & ~n5605 ;
  assign n5608 = ~n5606 & n5607 ;
  assign n5609 = n761 & ~n5608 ;
  assign n5610 = ~n5604 & ~n5609 ;
  assign n5611 = ~n5598 & n5610 ;
  assign n5612 = ~\sa20_reg[0]/P0001  & ~n5611 ;
  assign n5613 = n694 & n5527 ;
  assign n5614 = ~\sa20_reg[6]/NET0131  & n718 ;
  assign n5615 = ~n5613 & ~n5614 ;
  assign n5616 = ~\sa20_reg[2]/P0001  & ~n5615 ;
  assign n5617 = n691 & n744 ;
  assign n5618 = \sa20_reg[2]/P0001  & ~n5543 ;
  assign n5619 = \sa20_reg[3]/P0001  & n708 ;
  assign n5620 = ~\sa20_reg[7]/NET0131  & n5619 ;
  assign n5621 = ~n702 & ~n5620 ;
  assign n5622 = n5618 & n5621 ;
  assign n5623 = ~\sa20_reg[2]/P0001  & ~n766 ;
  assign n5624 = n5601 & n5623 ;
  assign n5625 = ~n5622 & ~n5624 ;
  assign n5626 = ~n5617 & ~n5625 ;
  assign n5627 = ~\sa20_reg[1]/P0001  & ~n5626 ;
  assign n5628 = ~n5616 & ~n5627 ;
  assign n5629 = ~n5612 & n5628 ;
  assign n5630 = ~n5566 & n5629 ;
  assign n5631 = ~n5580 & n5630 ;
  assign n5632 = \u0_w_reg[2][7]/P0001  & ~n5631 ;
  assign n5633 = ~\u0_w_reg[2][7]/P0001  & n5631 ;
  assign n5634 = ~n5632 & ~n5633 ;
  assign n5635 = n1300 & n5634 ;
  assign n5636 = ~n1300 & ~n5634 ;
  assign n5637 = ~n5635 & ~n5636 ;
  assign n5639 = n5522 & n5637 ;
  assign n5638 = ~n5522 & ~n5637 ;
  assign n5640 = ~\ld_r_reg/P0001  & ~n5638 ;
  assign n5641 = ~n5639 & n5640 ;
  assign n5643 = ~\text_in_r_reg[39]/P0001  & \u0_w_reg[2][7]/P0001  ;
  assign n5642 = \text_in_r_reg[39]/P0001  & ~\u0_w_reg[2][7]/P0001  ;
  assign n5644 = \ld_r_reg/P0001  & ~n5642 ;
  assign n5645 = ~n5643 & n5644 ;
  assign n5646 = ~n5641 & ~n5645 ;
  assign n5647 = \sa13_reg[2]/P0001  & n588 ;
  assign n5652 = ~\sa13_reg[1]/P0001  & ~n560 ;
  assign n5653 = ~n5647 & n5652 ;
  assign n5650 = \sa13_reg[3]/P0001  & n583 ;
  assign n5651 = ~\sa13_reg[4]/P0001  & n5650 ;
  assign n5648 = \sa13_reg[5]/P0001  & n5459 ;
  assign n5649 = n611 & n946 ;
  assign n5654 = ~n5648 & ~n5649 ;
  assign n5655 = ~n5651 & n5654 ;
  assign n5656 = n5653 & n5655 ;
  assign n5658 = \sa13_reg[7]/NET0131  & n632 ;
  assign n5659 = ~n865 & ~n5658 ;
  assign n5660 = ~\sa13_reg[2]/P0001  & ~n5659 ;
  assign n5657 = \sa13_reg[1]/P0001  & ~n681 ;
  assign n5661 = n549 & n670 ;
  assign n5662 = ~n918 & ~n5661 ;
  assign n5663 = n5657 & n5662 ;
  assign n5664 = ~n5660 & n5663 ;
  assign n5665 = ~n5656 & ~n5664 ;
  assign n5666 = ~n616 & ~n655 ;
  assign n5667 = ~\sa13_reg[6]/NET0131  & ~n5666 ;
  assign n5668 = \sa13_reg[2]/P0001  & ~n637 ;
  assign n5669 = ~n888 & n5668 ;
  assign n5670 = ~n5667 & n5669 ;
  assign n5671 = n550 & n583 ;
  assign n5672 = ~\sa13_reg[2]/P0001  & ~n5671 ;
  assign n5673 = ~n683 & n5672 ;
  assign n5674 = ~n903 & n5673 ;
  assign n5675 = ~n5670 & ~n5674 ;
  assign n5676 = ~n5665 & ~n5675 ;
  assign n5677 = \sa13_reg[0]/P0001  & ~n5676 ;
  assign n5679 = n547 & n5458 ;
  assign n5721 = n568 & ~n655 ;
  assign n5722 = ~n5679 & ~n5721 ;
  assign n5723 = ~\sa13_reg[2]/P0001  & ~n5722 ;
  assign n5725 = \sa13_reg[2]/P0001  & n861 ;
  assign n5724 = n603 & n5456 ;
  assign n5726 = ~n545 & ~n5724 ;
  assign n5727 = ~n5725 & n5726 ;
  assign n5728 = ~n5723 & n5727 ;
  assign n5729 = \sa13_reg[1]/P0001  & ~n5728 ;
  assign n5696 = \sa13_reg[2]/P0001  & n5505 ;
  assign n5717 = ~n887 & ~n5696 ;
  assign n5715 = \sa13_reg[3]/P0001  & n672 ;
  assign n5716 = n861 & n5424 ;
  assign n5718 = ~n5715 & ~n5716 ;
  assign n5719 = n5717 & n5718 ;
  assign n5720 = ~\sa13_reg[1]/P0001  & ~n5719 ;
  assign n5710 = ~n914 & ~n5492 ;
  assign n5711 = ~\sa13_reg[3]/P0001  & ~n5710 ;
  assign n5712 = n653 & n912 ;
  assign n5713 = ~n5500 & ~n5712 ;
  assign n5714 = \sa13_reg[2]/P0001  & ~n5713 ;
  assign n5730 = ~n5711 & ~n5714 ;
  assign n5731 = ~n5720 & n5730 ;
  assign n5732 = ~n5729 & n5731 ;
  assign n5733 = ~\sa13_reg[0]/P0001  & ~n5732 ;
  assign n5681 = \sa13_reg[5]/P0001  & ~n5443 ;
  assign n5682 = n547 & n592 ;
  assign n5680 = ~\sa13_reg[3]/P0001  & n5679 ;
  assign n5683 = \sa13_reg[2]/P0001  & ~n5423 ;
  assign n5684 = ~n5680 & n5683 ;
  assign n5685 = ~n5682 & n5684 ;
  assign n5686 = ~n5681 & n5685 ;
  assign n5687 = \sa13_reg[5]/P0001  & n5651 ;
  assign n5688 = ~\sa13_reg[2]/P0001  & ~n621 ;
  assign n5689 = ~n856 & n5688 ;
  assign n5690 = ~n5687 & n5689 ;
  assign n5691 = ~n5686 & ~n5690 ;
  assign n5678 = n557 & n653 ;
  assign n5692 = ~n609 & ~n5678 ;
  assign n5693 = ~n5691 & n5692 ;
  assign n5694 = ~\sa13_reg[1]/P0001  & ~n5693 ;
  assign n5695 = ~\sa13_reg[2]/P0001  & n908 ;
  assign n5697 = ~n5695 & ~n5696 ;
  assign n5698 = \sa13_reg[3]/P0001  & ~n5697 ;
  assign n5699 = \sa13_reg[7]/NET0131  & n668 ;
  assign n5700 = ~n634 & ~n683 ;
  assign n5701 = ~n5699 & n5700 ;
  assign n5702 = ~\sa13_reg[2]/P0001  & ~n5701 ;
  assign n5705 = ~n624 & ~n5440 ;
  assign n5703 = n567 & n603 ;
  assign n5704 = n955 & n5458 ;
  assign n5706 = ~n5703 & ~n5704 ;
  assign n5707 = n5705 & n5706 ;
  assign n5708 = ~n5702 & n5707 ;
  assign n5709 = \sa13_reg[1]/P0001  & ~n5708 ;
  assign n5734 = ~n5698 & ~n5709 ;
  assign n5735 = ~n5694 & n5734 ;
  assign n5736 = ~n5733 & n5735 ;
  assign n5737 = ~n5677 & n5736 ;
  assign n5749 = n1042 & ~n1059 ;
  assign n5750 = n982 & n5130 ;
  assign n5751 = ~n5749 & ~n5750 ;
  assign n5752 = ~\sa02_reg[2]/P0001  & ~n5751 ;
  assign n5755 = \sa02_reg[4]/P0001  & n1003 ;
  assign n5756 = n978 & n5755 ;
  assign n5753 = \sa02_reg[2]/P0001  & n1056 ;
  assign n5754 = \sa02_reg[6]/NET0131  & n5753 ;
  assign n5757 = ~n1123 & ~n5754 ;
  assign n5758 = ~n5756 & n5757 ;
  assign n5759 = ~n5752 & n5758 ;
  assign n5760 = \sa02_reg[1]/P0001  & ~n5759 ;
  assign n5738 = ~\sa02_reg[3]/P0001  & n1088 ;
  assign n5739 = ~\sa02_reg[2]/P0001  & n5738 ;
  assign n5740 = ~n1116 & ~n5739 ;
  assign n5741 = ~\sa02_reg[1]/P0001  & ~n5740 ;
  assign n5747 = ~n1077 & ~n5394 ;
  assign n5748 = ~\sa02_reg[3]/P0001  & ~n5747 ;
  assign n5742 = ~n5083 & ~n5403 ;
  assign n5743 = \sa02_reg[2]/P0001  & ~n5742 ;
  assign n5744 = \sa02_reg[4]/P0001  & n975 ;
  assign n5745 = ~n980 & ~n5744 ;
  assign n5746 = n5106 & ~n5745 ;
  assign n5761 = ~n5743 & ~n5746 ;
  assign n5762 = ~n5748 & n5761 ;
  assign n5763 = ~n5741 & n5762 ;
  assign n5764 = ~n5760 & n5763 ;
  assign n5765 = ~\sa02_reg[0]/P0001  & ~n5764 ;
  assign n5767 = ~\sa02_reg[4]/P0001  & n1025 ;
  assign n5768 = n982 & n1000 ;
  assign n5769 = ~n5767 & ~n5768 ;
  assign n5770 = ~\sa02_reg[2]/P0001  & ~n5769 ;
  assign n5766 = n1016 & n5130 ;
  assign n5771 = \sa02_reg[1]/P0001  & ~n5766 ;
  assign n5772 = ~n1061 & n5771 ;
  assign n5773 = ~n1110 & n5772 ;
  assign n5774 = ~n5770 & n5773 ;
  assign n5775 = \sa02_reg[2]/P0001  & n1001 ;
  assign n5780 = n1068 & n5130 ;
  assign n5781 = ~\sa02_reg[1]/P0001  & ~n5780 ;
  assign n5782 = ~n5775 & n5781 ;
  assign n5776 = ~\sa02_reg[2]/P0001  & n1091 ;
  assign n5777 = ~\sa02_reg[2]/P0001  & ~\sa02_reg[4]/P0001  ;
  assign n5778 = ~\sa02_reg[3]/P0001  & ~n5777 ;
  assign n5779 = n993 & ~n5778 ;
  assign n5783 = ~n5776 & ~n5779 ;
  assign n5784 = n5782 & n5783 ;
  assign n5785 = ~n5774 & ~n5784 ;
  assign n5788 = \sa02_reg[2]/P0001  & ~n1109 ;
  assign n5787 = n1023 & n1035 ;
  assign n5786 = ~\sa02_reg[7]/NET0131  & n986 ;
  assign n5789 = ~n5172 & ~n5786 ;
  assign n5790 = ~n5787 & n5789 ;
  assign n5791 = n5788 & n5790 ;
  assign n5792 = n1019 & n1035 ;
  assign n5793 = ~\sa02_reg[2]/P0001  & ~n1069 ;
  assign n5794 = ~n5792 & n5793 ;
  assign n5795 = ~n5181 & n5794 ;
  assign n5796 = ~n5791 & ~n5795 ;
  assign n5797 = ~n5785 & ~n5796 ;
  assign n5798 = \sa02_reg[0]/P0001  & ~n5797 ;
  assign n5819 = ~n977 & ~n5142 ;
  assign n5820 = ~n5181 & n5819 ;
  assign n5821 = ~\sa02_reg[2]/P0001  & ~n5820 ;
  assign n5822 = ~n1114 & ~n5128 ;
  assign n5818 = n1059 & n1094 ;
  assign n5823 = ~n5338 & ~n5818 ;
  assign n5824 = n5822 & n5823 ;
  assign n5825 = ~n5821 & n5824 ;
  assign n5826 = \sa02_reg[1]/P0001  & ~n5825 ;
  assign n5799 = \sa02_reg[5]/P0001  & ~n5326 ;
  assign n5800 = ~n986 & ~n1059 ;
  assign n5801 = n1094 & n5800 ;
  assign n5802 = \sa02_reg[2]/P0001  & ~n5347 ;
  assign n5803 = ~n5801 & n5802 ;
  assign n5804 = ~n5799 & n5803 ;
  assign n5805 = n1004 & n1030 ;
  assign n5806 = ~n1012 & ~n5805 ;
  assign n5807 = n1108 & n5806 ;
  assign n5808 = ~n5804 & ~n5807 ;
  assign n5809 = ~\sa02_reg[3]/P0001  & n1084 ;
  assign n5810 = ~\sa02_reg[6]/NET0131  & n5809 ;
  assign n5811 = ~n5122 & ~n5810 ;
  assign n5812 = ~n5808 & n5811 ;
  assign n5813 = ~\sa02_reg[1]/P0001  & ~n5812 ;
  assign n5815 = \sa02_reg[2]/P0001  & ~n5744 ;
  assign n5814 = ~\sa02_reg[2]/P0001  & ~n1072 ;
  assign n5816 = \sa02_reg[3]/P0001  & ~n5814 ;
  assign n5817 = ~n5815 & n5816 ;
  assign n5827 = ~n5813 & ~n5817 ;
  assign n5828 = ~n5826 & n5827 ;
  assign n5829 = ~n5798 & n5828 ;
  assign n5830 = ~n5765 & n5829 ;
  assign n5831 = n5737 & ~n5830 ;
  assign n5832 = ~n5737 & n5830 ;
  assign n5833 = ~n5831 & ~n5832 ;
  assign n5844 = n693 & n799 ;
  assign n5845 = ~\sa20_reg[2]/P0001  & ~n692 ;
  assign n5846 = ~n5844 & n5845 ;
  assign n5847 = \sa20_reg[2]/P0001  & ~n833 ;
  assign n5848 = ~n5556 & n5847 ;
  assign n5849 = ~n5846 & ~n5848 ;
  assign n5843 = n705 & n763 ;
  assign n5839 = n716 & n744 ;
  assign n5851 = ~n740 & ~n5839 ;
  assign n5852 = ~n5843 & n5851 ;
  assign n5850 = \sa20_reg[1]/P0001  & ~n737 ;
  assign n5853 = ~n5613 & n5850 ;
  assign n5854 = ~n5620 & n5853 ;
  assign n5855 = n5852 & n5854 ;
  assign n5856 = ~n5849 & n5855 ;
  assign n5861 = ~\sa20_reg[1]/P0001  & ~n821 ;
  assign n5860 = n5526 & n5619 ;
  assign n5857 = n736 & n791 ;
  assign n5858 = \sa20_reg[6]/NET0131  & n744 ;
  assign n5859 = n799 & n5858 ;
  assign n5862 = ~n5857 & ~n5859 ;
  assign n5863 = ~n5860 & n5862 ;
  assign n5864 = n5861 & n5863 ;
  assign n5865 = ~n5856 & ~n5864 ;
  assign n5834 = n722 & n831 ;
  assign n5835 = n691 & n728 ;
  assign n5836 = \sa20_reg[2]/P0001  & ~n5835 ;
  assign n5837 = \sa20_reg[6]/NET0131  & ~n706 ;
  assign n5838 = n709 & ~n5837 ;
  assign n5840 = ~n5838 & ~n5839 ;
  assign n5841 = n5836 & n5840 ;
  assign n5842 = ~n5834 & ~n5841 ;
  assign n5866 = ~\sa20_reg[0]/P0001  & ~n710 ;
  assign n5867 = ~n5842 & n5866 ;
  assign n5868 = ~n5865 & n5867 ;
  assign n5883 = ~\sa20_reg[4]/P0001  & n735 ;
  assign n5884 = n716 & n723 ;
  assign n5885 = ~n5883 & ~n5884 ;
  assign n5886 = \sa20_reg[2]/P0001  & ~n5885 ;
  assign n5887 = ~\sa20_reg[1]/P0001  & ~n778 ;
  assign n5888 = ~n5524 & n5887 ;
  assign n5882 = n763 & n5544 ;
  assign n5889 = ~n703 & ~n5882 ;
  assign n5890 = n5888 & n5889 ;
  assign n5891 = ~n5886 & n5890 ;
  assign n5892 = ~\sa20_reg[3]/P0001  & n715 ;
  assign n5893 = ~n752 & ~n5892 ;
  assign n5894 = n691 & n820 ;
  assign n5895 = n705 & n745 ;
  assign n5896 = \sa20_reg[1]/P0001  & ~n5895 ;
  assign n5897 = ~n5894 & n5896 ;
  assign n5898 = n5893 & n5897 ;
  assign n5899 = ~n5891 & ~n5898 ;
  assign n5869 = ~n714 & n748 ;
  assign n5870 = ~n810 & ~n5869 ;
  assign n5871 = \sa20_reg[1]/P0001  & ~n5870 ;
  assign n5872 = n693 & n745 ;
  assign n5873 = ~n778 & ~n5872 ;
  assign n5874 = ~\sa20_reg[4]/P0001  & n777 ;
  assign n5875 = ~\sa20_reg[2]/P0001  & ~n5874 ;
  assign n5876 = n5873 & n5875 ;
  assign n5877 = ~n5871 & n5876 ;
  assign n5878 = n728 & n799 ;
  assign n5879 = \sa20_reg[2]/P0001  & ~n703 ;
  assign n5880 = ~n5878 & n5879 ;
  assign n5881 = ~n5877 & ~n5880 ;
  assign n5901 = n694 & n699 ;
  assign n5900 = n5523 & n5585 ;
  assign n5902 = \sa20_reg[0]/P0001  & ~n5900 ;
  assign n5903 = ~n5901 & n5902 ;
  assign n5904 = ~n5881 & n5903 ;
  assign n5905 = ~n5899 & n5904 ;
  assign n5906 = ~n5868 & ~n5905 ;
  assign n5916 = \sa20_reg[2]/P0001  & ~n790 ;
  assign n5917 = ~n831 & ~n5916 ;
  assign n5915 = \sa20_reg[3]/P0001  & n710 ;
  assign n5918 = \sa20_reg[1]/P0001  & ~n5915 ;
  assign n5919 = ~n5917 & n5918 ;
  assign n5920 = ~n728 & ~n5544 ;
  assign n5921 = ~n5858 & n5920 ;
  assign n5922 = n691 & ~n5921 ;
  assign n5923 = ~n751 & ~n5922 ;
  assign n5924 = \sa20_reg[2]/P0001  & ~n5923 ;
  assign n5925 = ~\sa20_reg[1]/P0001  & ~n809 ;
  assign n5926 = ~n5924 & n5925 ;
  assign n5927 = ~n5919 & ~n5926 ;
  assign n5907 = n714 & n735 ;
  assign n5908 = n694 & n736 ;
  assign n5909 = ~n5907 & ~n5908 ;
  assign n5910 = ~n779 & n5909 ;
  assign n5911 = ~\sa20_reg[1]/P0001  & ~n5910 ;
  assign n5912 = ~n737 & ~n817 ;
  assign n5913 = ~n5911 & n5912 ;
  assign n5914 = ~\sa20_reg[2]/P0001  & ~n5913 ;
  assign n5928 = n761 & n5606 ;
  assign n5929 = ~n5914 & ~n5928 ;
  assign n5930 = ~n5927 & n5929 ;
  assign n5931 = ~n5906 & n5930 ;
  assign n5932 = n973 & ~n5931 ;
  assign n5933 = ~n973 & n5931 ;
  assign n5934 = ~n5932 & ~n5933 ;
  assign n5935 = \u0_w_reg[2][29]/P0001  & ~n5307 ;
  assign n5936 = ~\u0_w_reg[2][29]/P0001  & n5307 ;
  assign n5937 = ~n5935 & ~n5936 ;
  assign n5938 = n5934 & n5937 ;
  assign n5939 = ~n5934 & ~n5937 ;
  assign n5940 = ~n5938 & ~n5939 ;
  assign n5942 = n5833 & ~n5940 ;
  assign n5941 = ~n5833 & n5940 ;
  assign n5943 = ~\ld_r_reg/P0001  & ~n5941 ;
  assign n5944 = ~n5942 & n5943 ;
  assign n5946 = ~\text_in_r_reg[61]/P0001  & \u0_w_reg[2][29]/P0001  ;
  assign n5945 = \text_in_r_reg[61]/P0001  & ~\u0_w_reg[2][29]/P0001  ;
  assign n5947 = \ld_r_reg/P0001  & ~n5945 ;
  assign n5948 = ~n5946 & n5947 ;
  assign n5949 = ~n5944 & ~n5948 ;
  assign n5950 = ~n5191 & ~n5934 ;
  assign n5951 = n5191 & n5934 ;
  assign n5952 = ~n5950 & ~n5951 ;
  assign n5953 = \u0_w_reg[2][22]/P0001  & ~n1300 ;
  assign n5954 = ~\u0_w_reg[2][22]/P0001  & n1300 ;
  assign n5955 = ~n5953 & ~n5954 ;
  assign n5956 = n850 & n5955 ;
  assign n5957 = ~n850 & ~n5955 ;
  assign n5958 = ~n5956 & ~n5957 ;
  assign n5960 = n5952 & n5958 ;
  assign n5959 = ~n5952 & ~n5958 ;
  assign n5961 = ~\ld_r_reg/P0001  & ~n5959 ;
  assign n5962 = ~n5960 & n5961 ;
  assign n5964 = ~\text_in_r_reg[54]/P0001  & \u0_w_reg[2][22]/P0001  ;
  assign n5963 = \text_in_r_reg[54]/P0001  & ~\u0_w_reg[2][22]/P0001  ;
  assign n5965 = \ld_r_reg/P0001  & ~n5963 ;
  assign n5966 = ~n5964 & n5965 ;
  assign n5967 = ~n5962 & ~n5966 ;
  assign n5979 = \sa20_reg[5]/P0001  & n705 ;
  assign n5980 = ~n745 & n5979 ;
  assign n5981 = n708 & n765 ;
  assign n5982 = ~n5980 & ~n5981 ;
  assign n5983 = ~\sa20_reg[2]/P0001  & ~n5982 ;
  assign n5986 = n819 & n5585 ;
  assign n5984 = \sa20_reg[2]/P0001  & ~\sa20_reg[7]/NET0131  ;
  assign n5985 = n701 & n5984 ;
  assign n5987 = ~n700 & ~n5985 ;
  assign n5988 = ~n5986 & n5987 ;
  assign n5989 = ~n5983 & n5988 ;
  assign n5990 = \sa20_reg[1]/P0001  & ~n5989 ;
  assign n5973 = \sa20_reg[5]/P0001  & n5527 ;
  assign n5974 = ~\sa20_reg[2]/P0001  & n5973 ;
  assign n5972 = \sa20_reg[2]/P0001  & n5532 ;
  assign n5975 = ~n829 & ~n5581 ;
  assign n5976 = ~n5972 & n5975 ;
  assign n5977 = ~n5974 & n5976 ;
  assign n5978 = ~\sa20_reg[1]/P0001  & ~n5977 ;
  assign n5969 = ~n5541 & ~n5900 ;
  assign n5970 = ~\sa20_reg[3]/P0001  & ~n5969 ;
  assign n5968 = n724 & n799 ;
  assign n5971 = n716 & n5581 ;
  assign n5991 = ~n5968 & ~n5971 ;
  assign n5992 = ~n5970 & n5991 ;
  assign n5993 = ~n5978 & n5992 ;
  assign n5994 = ~n5990 & n5993 ;
  assign n5995 = ~\sa20_reg[0]/P0001  & ~n5994 ;
  assign n6038 = \sa20_reg[2]/P0001  & ~n778 ;
  assign n6039 = ~n5525 & n6038 ;
  assign n6037 = \sa20_reg[7]/NET0131  & n800 ;
  assign n6036 = n714 & n5619 ;
  assign n6040 = ~n725 & ~n6036 ;
  assign n6041 = ~n6037 & n6040 ;
  assign n6042 = n6039 & n6041 ;
  assign n6046 = ~\sa20_reg[2]/P0001  & ~n779 ;
  assign n6043 = n810 & n826 ;
  assign n6044 = ~\sa20_reg[3]/P0001  & ~n709 ;
  assign n6045 = n735 & n6044 ;
  assign n6047 = ~n6043 & ~n6045 ;
  assign n6048 = n6046 & n6047 ;
  assign n6049 = ~n6042 & ~n6048 ;
  assign n6050 = ~n5968 & ~n6049 ;
  assign n6051 = ~\sa20_reg[1]/P0001  & ~n6050 ;
  assign n5997 = ~\sa20_reg[4]/P0001  & n693 ;
  assign n5998 = n708 & n714 ;
  assign n5999 = ~n5997 & ~n5998 ;
  assign n6000 = ~\sa20_reg[2]/P0001  & ~n5999 ;
  assign n5996 = \sa20_reg[1]/P0001  & ~n817 ;
  assign n6001 = n705 & n5526 ;
  assign n6002 = ~n5894 & ~n6001 ;
  assign n6003 = n5996 & n6002 ;
  assign n6004 = ~n6000 & n6003 ;
  assign n6005 = n745 & n826 ;
  assign n6006 = ~\sa20_reg[1]/P0001  & ~n6005 ;
  assign n6007 = n763 & n807 ;
  assign n6011 = n6006 & ~n6007 ;
  assign n6008 = \sa20_reg[2]/P0001  & n715 ;
  assign n6009 = ~\sa20_reg[3]/P0001  & ~n5582 ;
  assign n6010 = n744 & ~n6009 ;
  assign n6012 = ~n6008 & ~n6010 ;
  assign n6013 = n6011 & n6012 ;
  assign n6014 = ~n6004 & ~n6013 ;
  assign n6015 = n796 & ~n5872 ;
  assign n6016 = ~n824 & n6015 ;
  assign n6017 = ~n707 & ~n789 ;
  assign n6018 = ~n816 & n6017 ;
  assign n6019 = n828 & n6018 ;
  assign n6020 = ~n6016 & ~n6019 ;
  assign n6021 = ~n6014 & ~n6020 ;
  assign n6022 = \sa20_reg[0]/P0001  & ~n6021 ;
  assign n6023 = n782 & n5523 ;
  assign n6024 = ~n5972 & ~n6023 ;
  assign n6025 = \sa20_reg[3]/P0001  & ~n6024 ;
  assign n6026 = ~n792 & ~n824 ;
  assign n6027 = ~n5859 & n6026 ;
  assign n6028 = ~\sa20_reg[2]/P0001  & ~n6027 ;
  assign n6031 = ~n762 & ~n5543 ;
  assign n6029 = ~\sa20_reg[5]/P0001  & n5895 ;
  assign n6030 = n739 & n819 ;
  assign n6032 = ~n6029 & ~n6030 ;
  assign n6033 = n6031 & n6032 ;
  assign n6034 = ~n6028 & n6033 ;
  assign n6035 = \sa20_reg[1]/P0001  & ~n6034 ;
  assign n6052 = ~n6025 & ~n6035 ;
  assign n6053 = ~n6022 & n6052 ;
  assign n6054 = ~n6051 & n6053 ;
  assign n6055 = ~n5995 & n6054 ;
  assign n6056 = n5737 & ~n6055 ;
  assign n6057 = ~n5737 & n6055 ;
  assign n6058 = ~n6056 & ~n6057 ;
  assign n6059 = ~n1142 & ~n6058 ;
  assign n6060 = n1142 & n6058 ;
  assign n6061 = ~n6059 & ~n6060 ;
  assign n6062 = \u0_w_reg[2][21]/P0001  & ~n5307 ;
  assign n6063 = ~\u0_w_reg[2][21]/P0001  & n5307 ;
  assign n6064 = ~n6062 & ~n6063 ;
  assign n6065 = n5931 & n6064 ;
  assign n6066 = ~n5931 & ~n6064 ;
  assign n6067 = ~n6065 & ~n6066 ;
  assign n6069 = n6061 & n6067 ;
  assign n6068 = ~n6061 & ~n6067 ;
  assign n6070 = ~\ld_r_reg/P0001  & ~n6068 ;
  assign n6071 = ~n6069 & n6070 ;
  assign n6073 = ~\text_in_r_reg[53]/P0001  & \u0_w_reg[2][21]/P0001  ;
  assign n6072 = \text_in_r_reg[53]/P0001  & ~\u0_w_reg[2][21]/P0001  ;
  assign n6074 = \ld_r_reg/P0001  & ~n6072 ;
  assign n6075 = ~n6073 & n6074 ;
  assign n6076 = ~n6071 & ~n6075 ;
  assign n6077 = ~n1145 & ~n6055 ;
  assign n6078 = n1145 & n6055 ;
  assign n6079 = ~n6077 & ~n6078 ;
  assign n6114 = \sa31_reg[2]/P0001  & ~n1207 ;
  assign n6115 = n1163 & n1166 ;
  assign n6116 = ~n1226 & ~n5252 ;
  assign n6117 = ~n6115 & n6116 ;
  assign n6118 = n6114 & n6117 ;
  assign n6119 = n1182 & n5269 ;
  assign n6120 = ~\sa31_reg[2]/P0001  & ~n5271 ;
  assign n6121 = ~n6119 & n6120 ;
  assign n6122 = ~n1231 & n6121 ;
  assign n6123 = ~n6118 & ~n6122 ;
  assign n6092 = \sa31_reg[4]/P0001  & n1182 ;
  assign n6124 = ~\sa31_reg[6]/NET0131  & n6092 ;
  assign n6125 = ~n5199 & ~n6124 ;
  assign n6126 = ~\sa31_reg[2]/P0001  & ~n6125 ;
  assign n6127 = n1146 & n1244 ;
  assign n6128 = \sa31_reg[1]/P0001  & ~n6127 ;
  assign n6129 = ~n1227 & n6128 ;
  assign n6130 = ~n5253 & n6129 ;
  assign n6131 = ~n6126 & n6130 ;
  assign n6132 = ~\sa31_reg[2]/P0001  & n5242 ;
  assign n6133 = ~\sa31_reg[1]/P0001  & ~n6132 ;
  assign n6136 = ~\sa31_reg[2]/P0001  & ~\sa31_reg[4]/P0001  ;
  assign n6137 = ~\sa31_reg[3]/P0001  & ~n6136 ;
  assign n6138 = n1166 & ~n6137 ;
  assign n6134 = n1225 & n1256 ;
  assign n6135 = \sa31_reg[2]/P0001  & n1179 ;
  assign n6139 = ~n6134 & ~n6135 ;
  assign n6140 = ~n6138 & n6139 ;
  assign n6141 = n6133 & n6140 ;
  assign n6142 = ~n6131 & ~n6141 ;
  assign n6143 = ~n6123 & ~n6142 ;
  assign n6144 = \sa31_reg[0]/P0002  & ~n6143 ;
  assign n6088 = n1147 & ~n1225 ;
  assign n6089 = ~\sa31_reg[4]/P0001  & n5239 ;
  assign n6090 = ~n6088 & ~n6089 ;
  assign n6091 = ~\sa31_reg[2]/P0001  & ~n6090 ;
  assign n6094 = \sa31_reg[1]/P0001  & ~n1200 ;
  assign n6087 = \sa31_reg[2]/P0001  & n1194 ;
  assign n6093 = n1279 & n6092 ;
  assign n6095 = ~n6087 & ~n6093 ;
  assign n6096 = n6094 & n6095 ;
  assign n6097 = ~n6091 & n6096 ;
  assign n6100 = n1162 & n1193 ;
  assign n6101 = ~n1226 & ~n6100 ;
  assign n6102 = ~\sa31_reg[7]/P0001  & ~n6101 ;
  assign n6098 = \sa31_reg[2]/P0001  & n1219 ;
  assign n6099 = ~\sa31_reg[1]/P0001  & ~n6098 ;
  assign n6103 = \sa31_reg[2]/P0001  & n1277 ;
  assign n6104 = n6099 & ~n6103 ;
  assign n6105 = ~n6102 & n6104 ;
  assign n6106 = ~n6097 & ~n6105 ;
  assign n6080 = ~\sa31_reg[6]/NET0131  & n1181 ;
  assign n6081 = ~\sa31_reg[3]/P0001  & n5241 ;
  assign n6082 = ~n6080 & ~n6081 ;
  assign n6083 = \sa31_reg[2]/P0001  & ~n6082 ;
  assign n6084 = ~\sa31_reg[6]/NET0131  & n5268 ;
  assign n6085 = ~n5262 & ~n6084 ;
  assign n6086 = ~\sa31_reg[3]/P0001  & ~n6085 ;
  assign n6107 = ~n6083 & ~n6086 ;
  assign n6108 = ~n6106 & n6107 ;
  assign n6109 = ~\sa31_reg[0]/P0002  & ~n6108 ;
  assign n6110 = n1163 & n1180 ;
  assign n6111 = ~\sa31_reg[2]/P0001  & n6110 ;
  assign n6112 = ~n6103 & ~n6111 ;
  assign n6113 = \sa31_reg[3]/P0001  & ~n6112 ;
  assign n6148 = \sa31_reg[7]/P0001  & n1247 ;
  assign n6149 = ~n1231 & ~n1258 ;
  assign n6150 = ~n6148 & n6149 ;
  assign n6151 = ~\sa31_reg[2]/P0001  & ~n6150 ;
  assign n6154 = \sa31_reg[1]/P0001  & ~n1266 ;
  assign n6152 = n1159 & n1256 ;
  assign n6153 = ~\sa31_reg[5]/P0001  & n6152 ;
  assign n6145 = n1225 & n5239 ;
  assign n6146 = n1149 & n1279 ;
  assign n6147 = \sa31_reg[4]/P0001  & n6146 ;
  assign n6155 = ~n6145 & ~n6147 ;
  assign n6156 = ~n6153 & n6155 ;
  assign n6157 = n6154 & n6156 ;
  assign n6158 = ~n6151 & n6157 ;
  assign n6160 = n1256 & n5263 ;
  assign n6161 = ~\sa31_reg[2]/P0001  & ~n6160 ;
  assign n6162 = ~\sa31_reg[5]/P0001  & n1260 ;
  assign n6163 = ~n5206 & ~n6162 ;
  assign n6164 = n6161 & n6163 ;
  assign n6165 = ~n1196 & ~n1225 ;
  assign n6166 = n5239 & n6165 ;
  assign n6169 = \sa31_reg[2]/P0001  & ~n5270 ;
  assign n6170 = ~n6166 & n6169 ;
  assign n6167 = ~\sa31_reg[6]/NET0131  & n5263 ;
  assign n6168 = ~\sa31_reg[3]/P0001  & n1187 ;
  assign n6171 = ~n6167 & ~n6168 ;
  assign n6172 = n6170 & n6171 ;
  assign n6173 = ~n6164 & ~n6172 ;
  assign n6159 = n1178 & n1230 ;
  assign n6174 = ~\sa31_reg[1]/P0001  & ~n1278 ;
  assign n6175 = ~n6159 & n6174 ;
  assign n6176 = ~n6173 & n6175 ;
  assign n6177 = ~n6158 & ~n6176 ;
  assign n6178 = ~n6113 & ~n6177 ;
  assign n6179 = ~n6109 & n6178 ;
  assign n6180 = ~n6144 & n6179 ;
  assign n6181 = \u0_w_reg[2][13]/P0001  & ~n6180 ;
  assign n6182 = ~\u0_w_reg[2][13]/P0001  & n6180 ;
  assign n6183 = ~n6181 & ~n6182 ;
  assign n6184 = n5307 & n6183 ;
  assign n6185 = ~n5307 & ~n6183 ;
  assign n6186 = ~n6184 & ~n6185 ;
  assign n6188 = n6079 & n6186 ;
  assign n6187 = ~n6079 & ~n6186 ;
  assign n6189 = ~\ld_r_reg/P0001  & ~n6187 ;
  assign n6190 = ~n6188 & n6189 ;
  assign n6192 = \text_in_r_reg[45]/P0001  & \u0_w_reg[2][13]/P0001  ;
  assign n6191 = ~\text_in_r_reg[45]/P0001  & ~\u0_w_reg[2][13]/P0001  ;
  assign n6193 = \ld_r_reg/P0001  & ~n6191 ;
  assign n6194 = ~n6192 & n6193 ;
  assign n6195 = ~n6190 & ~n6194 ;
  assign n6196 = ~n5194 & ~n5931 ;
  assign n6197 = n5194 & n5931 ;
  assign n6198 = ~n6196 & ~n6197 ;
  assign n6199 = \u0_w_reg[2][14]/P0001  & ~n1300 ;
  assign n6200 = ~\u0_w_reg[2][14]/P0001  & n1300 ;
  assign n6201 = ~n6199 & ~n6200 ;
  assign n6202 = n5307 & n6201 ;
  assign n6203 = ~n5307 & ~n6201 ;
  assign n6204 = ~n6202 & ~n6203 ;
  assign n6206 = n6198 & n6204 ;
  assign n6205 = ~n6198 & ~n6204 ;
  assign n6207 = ~\ld_r_reg/P0001  & ~n6205 ;
  assign n6208 = ~n6206 & n6207 ;
  assign n6210 = ~\text_in_r_reg[46]/P0001  & \u0_w_reg[2][14]/P0001  ;
  assign n6209 = \text_in_r_reg[46]/P0001  & ~\u0_w_reg[2][14]/P0001  ;
  assign n6211 = \ld_r_reg/P0001  & ~n6209 ;
  assign n6212 = ~n6210 & n6211 ;
  assign n6213 = ~n6208 & ~n6212 ;
  assign n6229 = ~\sa13_reg[2]/P0001  & ~n572 ;
  assign n6230 = ~n665 & n6229 ;
  assign n6231 = \sa13_reg[2]/P0001  & ~n5671 ;
  assign n6232 = ~n862 & n6231 ;
  assign n6233 = ~n6230 & ~n6232 ;
  assign n6234 = ~n649 & ~n5687 ;
  assign n6235 = ~n6233 & n6234 ;
  assign n6236 = ~\sa13_reg[1]/P0001  & ~n6235 ;
  assign n6216 = \sa13_reg[6]/NET0131  & n550 ;
  assign n6217 = \sa13_reg[4]/P0001  & n6216 ;
  assign n6218 = ~n610 & ~n617 ;
  assign n6219 = ~n6217 & n6218 ;
  assign n6220 = ~\sa13_reg[2]/P0001  & ~n6219 ;
  assign n6214 = ~n541 & ~n605 ;
  assign n6215 = \sa13_reg[2]/P0001  & ~n6214 ;
  assign n6221 = ~n854 & n904 ;
  assign n6222 = ~n6215 & n6221 ;
  assign n6223 = ~n6220 & n6222 ;
  assign n6224 = \sa13_reg[1]/P0001  & ~n6223 ;
  assign n6227 = ~n921 & ~n5687 ;
  assign n6228 = ~\sa13_reg[2]/P0001  & ~n6227 ;
  assign n6225 = ~n536 & ~n650 ;
  assign n6226 = n603 & ~n6225 ;
  assign n6237 = ~n654 & ~n953 ;
  assign n6238 = ~n6226 & n6237 ;
  assign n6239 = ~n6228 & n6238 ;
  assign n6240 = ~n6224 & n6239 ;
  assign n6241 = ~n6236 & n6240 ;
  assign n6242 = ~\sa13_reg[0]/P0001  & ~n6241 ;
  assign n6243 = n540 & n555 ;
  assign n6244 = ~n571 & ~n6243 ;
  assign n6246 = ~\sa13_reg[5]/P0001  & n5458 ;
  assign n6245 = \sa13_reg[4]/P0001  & n912 ;
  assign n6247 = ~n5650 & ~n6245 ;
  assign n6248 = ~n6246 & n6247 ;
  assign n6249 = \sa13_reg[2]/P0001  & ~n6248 ;
  assign n6250 = n6244 & ~n6249 ;
  assign n6251 = \sa13_reg[1]/P0001  & ~n6250 ;
  assign n6264 = \sa13_reg[2]/P0001  & n855 ;
  assign n6265 = ~n913 & ~n5466 ;
  assign n6266 = ~n6264 & n6265 ;
  assign n6267 = ~\sa13_reg[3]/P0001  & ~n6266 ;
  assign n6254 = ~n608 & ~n928 ;
  assign n6255 = ~\sa13_reg[7]/NET0131  & ~n6254 ;
  assign n6252 = ~\sa13_reg[3]/P0001  & n5458 ;
  assign n6253 = n532 & n6252 ;
  assign n6256 = ~n670 & n864 ;
  assign n6257 = ~n6253 & ~n6256 ;
  assign n6258 = ~n6255 & n6257 ;
  assign n6259 = ~\sa13_reg[1]/P0001  & ~n6258 ;
  assign n6260 = ~n862 & ~n908 ;
  assign n6261 = ~n5466 & ~n5476 ;
  assign n6262 = n6260 & n6261 ;
  assign n6263 = ~\sa13_reg[2]/P0001  & ~n6262 ;
  assign n6268 = ~n6259 & ~n6263 ;
  assign n6269 = ~n6267 & n6268 ;
  assign n6270 = ~n6251 & n6269 ;
  assign n6271 = \sa13_reg[0]/P0001  & ~n6270 ;
  assign n6291 = ~n561 & ~n648 ;
  assign n6292 = ~n918 & n6291 ;
  assign n6293 = ~\sa13_reg[2]/P0001  & ~n6292 ;
  assign n6294 = ~n558 & ~n5682 ;
  assign n6295 = ~n6293 & n6294 ;
  assign n6296 = ~\sa13_reg[1]/P0001  & ~n6295 ;
  assign n6286 = \sa13_reg[1]/P0001  & \sa13_reg[2]/P0001  ;
  assign n6287 = ~n571 & ~n5505 ;
  assign n6288 = \sa13_reg[3]/P0001  & ~n6287 ;
  assign n6289 = ~n622 & ~n6288 ;
  assign n6290 = n6286 & ~n6289 ;
  assign n6272 = ~\sa13_reg[1]/P0001  & \sa13_reg[2]/P0001  ;
  assign n6273 = ~\sa13_reg[5]/P0001  & n617 ;
  assign n6274 = ~n654 & ~n6273 ;
  assign n6275 = ~n542 & n6274 ;
  assign n6276 = n6272 & ~n6275 ;
  assign n6277 = ~n587 & n920 ;
  assign n6278 = ~n537 & ~n548 ;
  assign n6279 = ~n6277 & n6278 ;
  assign n6280 = n680 & ~n6279 ;
  assign n6281 = \sa13_reg[2]/P0001  & \sa13_reg[4]/P0001  ;
  assign n6282 = n551 & n6281 ;
  assign n6283 = \sa13_reg[1]/P0001  & \sa13_reg[3]/P0001  ;
  assign n6284 = n547 & n611 ;
  assign n6285 = n6283 & n6284 ;
  assign n6297 = ~n6282 & ~n6285 ;
  assign n6298 = ~n5465 & n6297 ;
  assign n6299 = ~n6280 & n6298 ;
  assign n6300 = ~n6276 & n6299 ;
  assign n6301 = ~n6290 & n6300 ;
  assign n6302 = ~n6296 & n6301 ;
  assign n6303 = ~n6271 & n6302 ;
  assign n6304 = ~n6242 & n6303 ;
  assign n6337 = n976 & n1038 ;
  assign n6338 = ~n1005 & ~n6337 ;
  assign n6339 = ~\sa02_reg[5]/P0001  & ~n1015 ;
  assign n6340 = ~n5159 & n6339 ;
  assign n6341 = \sa02_reg[7]/NET0131  & n1068 ;
  assign n6342 = ~n6340 & ~n6341 ;
  assign n6343 = \sa02_reg[2]/P0001  & ~n6342 ;
  assign n6344 = n6338 & ~n6343 ;
  assign n6345 = \sa02_reg[1]/P0001  & ~n6344 ;
  assign n6354 = n1024 & ~n5168 ;
  assign n6353 = n999 & n1122 ;
  assign n6355 = ~n1057 & ~n1072 ;
  assign n6356 = ~n6353 & n6355 ;
  assign n6357 = ~n6354 & n6356 ;
  assign n6358 = ~\sa02_reg[1]/P0001  & ~n6357 ;
  assign n6346 = n1020 & ~n5777 ;
  assign n6347 = ~n5363 & ~n6346 ;
  assign n6348 = ~\sa02_reg[3]/P0001  & ~n6347 ;
  assign n6349 = ~n1072 & ~n5363 ;
  assign n6350 = ~n5156 & n6349 ;
  assign n6351 = ~n5738 & n6350 ;
  assign n6352 = ~\sa02_reg[2]/P0001  & ~n6351 ;
  assign n6359 = ~n6348 & ~n6352 ;
  assign n6360 = ~n6358 & n6359 ;
  assign n6361 = ~n6345 & n6360 ;
  assign n6362 = \sa02_reg[0]/P0001  & ~n6361 ;
  assign n6306 = ~n5084 & ~n5163 ;
  assign n6307 = ~\sa02_reg[2]/P0001  & ~n6306 ;
  assign n6305 = n1035 & n5082 ;
  assign n6308 = ~\sa02_reg[1]/P0001  & ~n5805 ;
  assign n6309 = ~n6305 & n6308 ;
  assign n6310 = ~n6307 & n6309 ;
  assign n6312 = ~\sa02_reg[3]/P0001  & n1023 ;
  assign n6311 = n1011 & n1038 ;
  assign n6313 = ~n983 & ~n6311 ;
  assign n6314 = ~n6312 & n6313 ;
  assign n6315 = ~\sa02_reg[2]/P0001  & ~n6314 ;
  assign n6316 = \sa02_reg[1]/P0001  & ~n1037 ;
  assign n6317 = n1083 & n6316 ;
  assign n6318 = ~n6315 & n6317 ;
  assign n6319 = ~n6310 & ~n6318 ;
  assign n6328 = ~n980 & ~n1015 ;
  assign n6329 = n978 & ~n6328 ;
  assign n6320 = \sa02_reg[2]/P0001  & n1058 ;
  assign n6330 = ~n1121 & ~n6320 ;
  assign n6331 = ~n6329 & n6330 ;
  assign n6325 = ~\sa02_reg[3]/P0001  & n976 ;
  assign n6326 = ~n994 & ~n6325 ;
  assign n6327 = n5154 & ~n6326 ;
  assign n6321 = ~n5738 & ~n5792 ;
  assign n6322 = n5106 & ~n6321 ;
  assign n6323 = ~n1063 & ~n5805 ;
  assign n6324 = ~\sa02_reg[2]/P0001  & ~n6323 ;
  assign n6332 = ~n6322 & ~n6324 ;
  assign n6333 = ~n6327 & n6332 ;
  assign n6334 = n6331 & n6333 ;
  assign n6335 = ~n6319 & n6334 ;
  assign n6336 = ~\sa02_reg[0]/P0001  & ~n6335 ;
  assign n6381 = ~\sa02_reg[3]/P0001  & n1094 ;
  assign n6382 = ~n1071 & ~n1121 ;
  assign n6383 = ~n6381 & n6382 ;
  assign n6384 = \sa02_reg[2]/P0001  & ~n6383 ;
  assign n6377 = n1038 & n1094 ;
  assign n6385 = ~n1058 & ~n6377 ;
  assign n6386 = ~n6384 & n6385 ;
  assign n6387 = ~\sa02_reg[1]/P0001  & ~n6386 ;
  assign n6373 = n1020 & ~n5800 ;
  assign n6374 = \sa02_reg[3]/P0001  & n5744 ;
  assign n6375 = ~n6373 & ~n6374 ;
  assign n6376 = \sa02_reg[1]/P0001  & ~n6375 ;
  assign n6378 = ~n1117 & ~n6377 ;
  assign n6379 = ~n6376 & n6378 ;
  assign n6380 = \sa02_reg[2]/P0001  & ~n6379 ;
  assign n6363 = ~\sa02_reg[1]/P0001  & ~\sa02_reg[2]/P0001  ;
  assign n6364 = n1025 & n1035 ;
  assign n6365 = ~n5102 & ~n6364 ;
  assign n6366 = ~n1061 & n6365 ;
  assign n6367 = n6363 & ~n6366 ;
  assign n6368 = ~n1000 & n1062 ;
  assign n6369 = ~n5081 & ~n5099 ;
  assign n6370 = ~n1037 & n6369 ;
  assign n6371 = ~n6368 & n6370 ;
  assign n6372 = n5179 & ~n6371 ;
  assign n6388 = ~n6367 & ~n6372 ;
  assign n6389 = ~n6380 & n6388 ;
  assign n6390 = ~n6387 & n6389 ;
  assign n6391 = ~n6336 & n6390 ;
  assign n6392 = ~n6362 & n6391 ;
  assign n6393 = ~n6304 & ~n6392 ;
  assign n6394 = n6304 & n6392 ;
  assign n6395 = ~n6393 & ~n6394 ;
  assign n6399 = ~\sa02_reg[5]/P0001  & n5155 ;
  assign n6400 = ~n1031 & ~n1076 ;
  assign n6401 = ~n6399 & n6400 ;
  assign n6402 = \sa02_reg[2]/P0001  & ~n6401 ;
  assign n6398 = n1059 & ~n5367 ;
  assign n6396 = n1003 & n5108 ;
  assign n6397 = n5159 & n6396 ;
  assign n6403 = ~n5809 & ~n6397 ;
  assign n6404 = ~n6398 & n6403 ;
  assign n6405 = ~n6402 & n6404 ;
  assign n6406 = \sa02_reg[0]/P0001  & ~n6405 ;
  assign n6407 = ~n975 & ~n1094 ;
  assign n6408 = n974 & ~n6407 ;
  assign n6409 = n1107 & ~n6408 ;
  assign n6410 = ~n1130 & ~n5082 ;
  assign n6411 = ~n5394 & n6410 ;
  assign n6412 = ~\sa02_reg[3]/P0001  & ~n6411 ;
  assign n6413 = ~\sa02_reg[2]/P0001  & ~n1070 ;
  assign n6414 = ~n6412 & n6413 ;
  assign n6415 = ~n6409 & ~n6414 ;
  assign n6416 = ~n6406 & ~n6415 ;
  assign n6417 = ~\sa02_reg[1]/P0001  & ~n6416 ;
  assign n6445 = ~n1110 & ~n5098 ;
  assign n6444 = n994 & n5108 ;
  assign n6446 = ~n5181 & ~n6444 ;
  assign n6447 = n6445 & n6446 ;
  assign n6448 = ~n1014 & n6447 ;
  assign n6449 = \sa02_reg[1]/P0001  & ~n6448 ;
  assign n6442 = \sa02_reg[6]/NET0131  & n5132 ;
  assign n6443 = n5168 & n5738 ;
  assign n6468 = ~n6442 & ~n6443 ;
  assign n6469 = ~n6449 & n6468 ;
  assign n6470 = ~n6417 & n6469 ;
  assign n6418 = \sa02_reg[6]/NET0131  & n1030 ;
  assign n6419 = ~n1063 & ~n6418 ;
  assign n6420 = ~n5148 & n6419 ;
  assign n6421 = ~\sa02_reg[2]/P0001  & ~n6420 ;
  assign n6424 = n1068 & n5753 ;
  assign n6422 = \sa02_reg[4]/P0001  & n6341 ;
  assign n6423 = n979 & ~n1038 ;
  assign n6425 = ~n6396 & ~n6423 ;
  assign n6426 = ~n6422 & n6425 ;
  assign n6427 = ~n6424 & n6426 ;
  assign n6428 = \sa02_reg[1]/P0001  & ~n6427 ;
  assign n6438 = ~n6421 & ~n6428 ;
  assign n6429 = ~\sa02_reg[3]/P0001  & ~n5389 ;
  assign n6430 = ~n5776 & ~n6429 ;
  assign n6431 = ~\sa02_reg[1]/P0001  & ~n6430 ;
  assign n6432 = ~n1011 & ~n5091 ;
  assign n6433 = n1059 & ~n6432 ;
  assign n6434 = ~\sa02_reg[1]/P0001  & n993 ;
  assign n6435 = ~n1068 & n6434 ;
  assign n6436 = ~n6433 & ~n6435 ;
  assign n6437 = \sa02_reg[2]/P0001  & ~n6436 ;
  assign n6439 = ~n6431 & ~n6437 ;
  assign n6440 = n6438 & n6439 ;
  assign n6441 = ~\sa02_reg[0]/P0001  & ~n6440 ;
  assign n6458 = ~n975 & ~n980 ;
  assign n6459 = ~\sa02_reg[2]/P0001  & ~n6458 ;
  assign n6460 = ~n5163 & ~n6459 ;
  assign n6461 = \sa02_reg[1]/P0001  & ~n6460 ;
  assign n6450 = ~n1063 & ~n5750 ;
  assign n6451 = n5103 & n6450 ;
  assign n6452 = \sa02_reg[2]/P0001  & ~n6451 ;
  assign n6453 = \sa02_reg[5]/P0001  & n5786 ;
  assign n6454 = ~n5364 & ~n6453 ;
  assign n6455 = ~\sa02_reg[2]/P0001  & ~n6454 ;
  assign n6456 = ~n1011 & ~n1015 ;
  assign n6457 = n1095 & ~n6456 ;
  assign n6462 = ~n5738 & ~n5818 ;
  assign n6463 = ~n6457 & n6462 ;
  assign n6464 = ~n6455 & n6463 ;
  assign n6465 = ~n6452 & n6464 ;
  assign n6466 = ~n6461 & n6465 ;
  assign n6467 = \sa02_reg[0]/P0001  & ~n6466 ;
  assign n6471 = ~n6441 & ~n6467 ;
  assign n6472 = n6470 & n6471 ;
  assign n6473 = ~n5417 & ~n6472 ;
  assign n6474 = n5417 & n6472 ;
  assign n6475 = ~n6473 & ~n6474 ;
  assign n6476 = n6395 & ~n6475 ;
  assign n6477 = ~n6395 & n6475 ;
  assign n6478 = ~n6476 & ~n6477 ;
  assign n6500 = ~n1220 & ~n5261 ;
  assign n6501 = ~n5209 & n6500 ;
  assign n6502 = \sa31_reg[2]/P0001  & ~n6501 ;
  assign n6495 = n1162 & n5239 ;
  assign n6496 = \sa31_reg[4]/P0001  & n6495 ;
  assign n6497 = \sa31_reg[5]/P0001  & ~n1146 ;
  assign n6498 = n1225 & ~n6497 ;
  assign n6499 = n1152 & n1158 ;
  assign n6503 = ~n6498 & ~n6499 ;
  assign n6504 = ~n6496 & n6503 ;
  assign n6505 = ~n6502 & n6504 ;
  assign n6506 = ~\sa31_reg[1]/P0001  & ~n6505 ;
  assign n6492 = ~n1168 & ~n6089 ;
  assign n6493 = n5251 & n6492 ;
  assign n6494 = \sa31_reg[2]/P0001  & ~n6493 ;
  assign n6479 = ~n1193 & ~n1219 ;
  assign n6480 = ~\sa31_reg[2]/P0001  & ~n6479 ;
  assign n6481 = ~n1239 & ~n6480 ;
  assign n6482 = \sa31_reg[1]/P0001  & ~n6481 ;
  assign n6487 = n1158 & n1196 ;
  assign n6488 = \sa31_reg[7]/P0001  & n1277 ;
  assign n6489 = ~n6487 & ~n6488 ;
  assign n6490 = ~\sa31_reg[2]/P0001  & ~n6489 ;
  assign n6483 = \sa31_reg[3]/P0001  & n1151 ;
  assign n6484 = ~\sa31_reg[4]/P0001  & n1276 ;
  assign n6485 = ~n6483 & ~n6484 ;
  assign n6486 = ~\sa31_reg[2]/P0001  & ~n6485 ;
  assign n6491 = ~\sa31_reg[3]/P0001  & n1194 ;
  assign n6507 = ~n6145 & ~n6491 ;
  assign n6508 = ~n6486 & n6507 ;
  assign n6509 = ~n6490 & n6508 ;
  assign n6510 = ~n6482 & n6509 ;
  assign n6511 = ~n6494 & n6510 ;
  assign n6512 = ~n6506 & n6511 ;
  assign n6513 = \sa31_reg[0]/P0002  & ~n6512 ;
  assign n6543 = n1152 & n1178 ;
  assign n6544 = ~n1260 & ~n6543 ;
  assign n6545 = ~\sa31_reg[7]/P0001  & ~n6544 ;
  assign n6546 = ~\sa31_reg[3]/P0001  & n1173 ;
  assign n6547 = ~n5264 & ~n6546 ;
  assign n6548 = ~n6545 & n6547 ;
  assign n6549 = ~\sa31_reg[2]/P0001  & ~n6548 ;
  assign n6530 = ~\sa31_reg[4]/P0001  & n1229 ;
  assign n6531 = ~\sa31_reg[3]/P0001  & n6530 ;
  assign n6540 = \sa31_reg[7]/P0001  & n6531 ;
  assign n6541 = ~n1247 & ~n6540 ;
  assign n6542 = \sa31_reg[2]/P0001  & ~n6541 ;
  assign n6550 = ~n5295 & ~n6542 ;
  assign n6551 = ~n6549 & n6550 ;
  assign n6552 = ~\sa31_reg[1]/P0001  & ~n6551 ;
  assign n6528 = n1166 & n5269 ;
  assign n6529 = ~n5250 & ~n6528 ;
  assign n6532 = n6529 & ~n6531 ;
  assign n6533 = ~\sa31_reg[2]/P0001  & ~n6532 ;
  assign n6517 = ~n6110 & ~n6115 ;
  assign n6518 = ~\sa31_reg[3]/P0001  & ~n6517 ;
  assign n6519 = n6133 & ~n6518 ;
  assign n6520 = n1194 & n1265 ;
  assign n6523 = \sa31_reg[1]/P0001  & ~n6152 ;
  assign n6521 = ~n1159 & n1186 ;
  assign n6522 = n1162 & n1182 ;
  assign n6524 = ~n6521 & ~n6522 ;
  assign n6525 = n6523 & n6524 ;
  assign n6526 = ~n6520 & n6525 ;
  assign n6527 = ~n6519 & ~n6526 ;
  assign n6514 = ~\sa31_reg[1]/P0001  & \sa31_reg[2]/P0001  ;
  assign n6515 = n1166 & ~n5269 ;
  assign n6516 = n6514 & n6515 ;
  assign n6534 = ~n1151 & ~n1187 ;
  assign n6535 = n1248 & ~n6534 ;
  assign n6536 = ~n6516 & ~n6535 ;
  assign n6537 = ~n6527 & n6536 ;
  assign n6538 = ~n6533 & n6537 ;
  assign n6539 = ~\sa31_reg[0]/P0002  & ~n6538 ;
  assign n6553 = \sa31_reg[2]/P0001  & n6162 ;
  assign n6554 = ~n6167 & ~n6553 ;
  assign n6555 = ~\sa31_reg[7]/P0001  & ~n6554 ;
  assign n6556 = n1166 & n1196 ;
  assign n6557 = ~\sa31_reg[2]/P0001  & ~n6556 ;
  assign n6558 = ~n6114 & ~n6557 ;
  assign n6559 = ~n1231 & ~n6558 ;
  assign n6560 = ~n6555 & n6559 ;
  assign n6561 = \sa31_reg[1]/P0001  & ~n6560 ;
  assign n6562 = \sa31_reg[6]/NET0131  & n1222 ;
  assign n6563 = n1152 & n6087 ;
  assign n6564 = ~n6562 & ~n6563 ;
  assign n6565 = ~n6561 & n6564 ;
  assign n6566 = ~n6539 & n6565 ;
  assign n6567 = ~n6552 & n6566 ;
  assign n6568 = ~n6513 & n6567 ;
  assign n6635 = \sa31_reg[1]/P0001  & ~n1240 ;
  assign n6639 = ~n6553 & n6635 ;
  assign n6636 = \sa31_reg[7]/P0001  & n6162 ;
  assign n6637 = ~n1160 & ~n1217 ;
  assign n6638 = ~\sa31_reg[2]/P0001  & ~n6637 ;
  assign n6640 = ~n6636 & ~n6638 ;
  assign n6641 = n6639 & n6640 ;
  assign n6642 = ~n5263 & ~n6136 ;
  assign n6643 = \sa31_reg[7]/P0001  & ~n6642 ;
  assign n6644 = n1265 & n6092 ;
  assign n6645 = n6099 & ~n6644 ;
  assign n6646 = ~n6643 & n6645 ;
  assign n6647 = ~n6641 & ~n6646 ;
  assign n6627 = \sa31_reg[4]/P0001  & n1187 ;
  assign n6628 = ~n6488 & ~n6627 ;
  assign n6629 = \sa31_reg[3]/P0001  & ~n6628 ;
  assign n6630 = \sa31_reg[2]/P0001  & ~n6629 ;
  assign n6631 = ~\sa31_reg[2]/P0001  & ~n1278 ;
  assign n6581 = ~\sa31_reg[3]/P0001  & n1201 ;
  assign n6582 = ~n6499 & ~n6581 ;
  assign n6632 = ~n1233 & n6582 ;
  assign n6633 = n6631 & n6632 ;
  assign n6634 = ~n6630 & ~n6633 ;
  assign n6648 = n1225 & n6098 ;
  assign n6649 = ~n6634 & ~n6648 ;
  assign n6650 = ~n6647 & n6649 ;
  assign n6651 = ~\sa31_reg[0]/P0002  & ~n6650 ;
  assign n6589 = ~\sa31_reg[4]/P0001  & n1256 ;
  assign n6590 = ~n5198 & ~n6589 ;
  assign n6591 = ~\sa31_reg[3]/P0001  & ~n6590 ;
  assign n6592 = ~n5209 & ~n6591 ;
  assign n6593 = \sa31_reg[2]/P0001  & ~n6592 ;
  assign n6596 = \sa31_reg[4]/P0001  & ~n1276 ;
  assign n6597 = \sa31_reg[6]/NET0131  & ~n6596 ;
  assign n6598 = \sa31_reg[4]/P0001  & n1229 ;
  assign n6599 = ~\sa31_reg[3]/P0001  & n1186 ;
  assign n6600 = ~n6598 & ~n6599 ;
  assign n6601 = ~n6597 & n6600 ;
  assign n6602 = n1232 & ~n6601 ;
  assign n6594 = ~n6153 & ~n6495 ;
  assign n6595 = \sa31_reg[1]/P0001  & ~n6594 ;
  assign n6604 = n1150 & n1162 ;
  assign n6603 = n1151 & n1248 ;
  assign n6605 = ~n6487 & ~n6603 ;
  assign n6606 = ~n6604 & n6605 ;
  assign n6607 = ~n6595 & n6606 ;
  assign n6608 = ~n6602 & n6607 ;
  assign n6609 = ~n6593 & n6608 ;
  assign n6610 = \sa31_reg[0]/P0002  & ~n6609 ;
  assign n6573 = \sa31_reg[4]/P0001  & ~n1178 ;
  assign n6574 = ~n5205 & n6573 ;
  assign n6575 = ~n1194 & ~n6574 ;
  assign n6576 = ~\sa31_reg[2]/P0001  & ~n6575 ;
  assign n6571 = ~\sa31_reg[4]/P0001  & n1182 ;
  assign n6572 = n1279 & n6571 ;
  assign n6569 = ~\sa31_reg[3]/P0001  & n1149 ;
  assign n6570 = ~n1244 & n6569 ;
  assign n6577 = ~n6167 & ~n6570 ;
  assign n6578 = ~n6572 & n6577 ;
  assign n6579 = ~n6576 & n6578 ;
  assign n6580 = \sa31_reg[0]/P0002  & ~n6579 ;
  assign n6583 = ~\sa31_reg[2]/P0001  & ~n6582 ;
  assign n6584 = n5238 & n6571 ;
  assign n6585 = ~n6556 & ~n6584 ;
  assign n6586 = ~n6583 & n6585 ;
  assign n6587 = ~n6580 & n6586 ;
  assign n6588 = ~\sa31_reg[1]/P0001  & ~n6587 ;
  assign n6611 = ~n6084 & ~n6589 ;
  assign n6612 = ~n6124 & n6611 ;
  assign n6613 = ~\sa31_reg[3]/P0001  & ~n6612 ;
  assign n6614 = ~n1183 & ~n5270 ;
  assign n6615 = ~n6613 & n6614 ;
  assign n6616 = n1232 & ~n6615 ;
  assign n6623 = \sa31_reg[5]/P0001  & n1260 ;
  assign n6624 = ~n5204 & ~n6153 ;
  assign n6625 = ~n6623 & n6624 ;
  assign n6626 = n6514 & ~n6625 ;
  assign n6617 = ~n5207 & ~n6080 ;
  assign n6618 = ~\sa31_reg[2]/P0001  & ~n6617 ;
  assign n6619 = ~n1187 & ~n5198 ;
  assign n6620 = n6517 & n6619 ;
  assign n6621 = \sa31_reg[1]/P0001  & n5238 ;
  assign n6622 = ~n6620 & n6621 ;
  assign n6652 = ~n6618 & ~n6622 ;
  assign n6653 = ~n6626 & n6652 ;
  assign n6654 = ~n6616 & n6653 ;
  assign n6655 = ~n6588 & n6654 ;
  assign n6656 = ~n6610 & n6655 ;
  assign n6657 = ~n6651 & n6656 ;
  assign n6658 = n6568 & ~n6657 ;
  assign n6659 = ~n6568 & n6657 ;
  assign n6660 = ~n6658 & ~n6659 ;
  assign n6689 = n716 & n5858 ;
  assign n6690 = ~n721 & ~n6689 ;
  assign n6691 = \sa20_reg[7]/NET0131  & n698 ;
  assign n6692 = ~n767 & ~n5529 ;
  assign n6693 = ~n6691 & n6692 ;
  assign n6694 = \sa20_reg[2]/P0001  & ~n6693 ;
  assign n6695 = n6690 & ~n6694 ;
  assign n6696 = \sa20_reg[1]/P0001  & ~n6695 ;
  assign n6706 = ~n834 & ~n5567 ;
  assign n6707 = ~n5606 & ~n5973 ;
  assign n6708 = n6706 & n6707 ;
  assign n6709 = ~\sa20_reg[2]/P0001  & ~n6708 ;
  assign n6699 = ~\sa20_reg[6]/NET0131  & n5908 ;
  assign n6697 = n716 & ~n826 ;
  assign n6698 = ~n717 & n6697 ;
  assign n6700 = ~n5567 & ~n5843 ;
  assign n6701 = ~n6698 & n6700 ;
  assign n6702 = ~n6699 & n6701 ;
  assign n6703 = ~\sa20_reg[1]/P0001  & ~n6702 ;
  assign n6704 = n737 & ~n5582 ;
  assign n6705 = \sa20_reg[4]/P0001  & n725 ;
  assign n6710 = ~n6704 & ~n6705 ;
  assign n6711 = ~n6703 & n6710 ;
  assign n6712 = ~n6709 & n6711 ;
  assign n6713 = ~n6696 & n6712 ;
  assign n6714 = \sa20_reg[0]/P0001  & ~n6713 ;
  assign n6673 = ~n738 & ~n832 ;
  assign n6674 = ~\sa20_reg[2]/P0001  & ~n6673 ;
  assign n6671 = ~n795 & ~n5973 ;
  assign n6672 = \sa20_reg[2]/P0001  & ~n6671 ;
  assign n6675 = ~n822 & ~n6043 ;
  assign n6676 = ~n6672 & n6675 ;
  assign n6677 = ~n6674 & n6676 ;
  assign n6678 = ~\sa20_reg[1]/P0001  & ~n6677 ;
  assign n6663 = \sa20_reg[4]/P0001  & ~n698 ;
  assign n6664 = n748 & ~n6663 ;
  assign n6665 = ~n769 & ~n6664 ;
  assign n6666 = ~\sa20_reg[2]/P0001  & ~n6665 ;
  assign n6661 = ~n781 & ~n5599 ;
  assign n6662 = \sa20_reg[2]/P0001  & ~n6661 ;
  assign n6667 = ~n5620 & n5873 ;
  assign n6668 = ~n6662 & n6667 ;
  assign n6669 = ~n6666 & n6668 ;
  assign n6670 = \sa20_reg[1]/P0001  & ~n6669 ;
  assign n6679 = ~n5892 & ~n6043 ;
  assign n6680 = ~\sa20_reg[2]/P0001  & ~n6679 ;
  assign n6681 = ~n709 & ~n820 ;
  assign n6682 = n819 & ~n6681 ;
  assign n6683 = ~n809 & ~n5928 ;
  assign n6684 = ~n6682 & n6683 ;
  assign n6685 = ~n6680 & n6684 ;
  assign n6686 = ~n6670 & n6685 ;
  assign n6687 = ~n6678 & n6686 ;
  assign n6688 = ~\sa20_reg[0]/P0001  & ~n6687 ;
  assign n6732 = ~n746 & ~n5591 ;
  assign n6733 = ~n5894 & n6732 ;
  assign n6734 = ~\sa20_reg[2]/P0001  & ~n6733 ;
  assign n6735 = ~n752 & ~n6036 ;
  assign n6736 = ~n6734 & n6735 ;
  assign n6737 = ~\sa20_reg[1]/P0001  & ~n6736 ;
  assign n6715 = ~\sa20_reg[3]/P0001  & n690 ;
  assign n6716 = ~n710 & ~n6715 ;
  assign n6717 = ~n5620 & n6716 ;
  assign n6718 = ~n714 & ~n6717 ;
  assign n6719 = ~n695 & ~n6718 ;
  assign n6720 = n815 & ~n6719 ;
  assign n6721 = ~n721 & ~n5532 ;
  assign n6722 = \sa20_reg[3]/P0001  & ~n6721 ;
  assign n6723 = ~n768 & ~n6722 ;
  assign n6724 = n806 & ~n6723 ;
  assign n6725 = ~n710 & ~n5998 ;
  assign n6726 = n761 & ~n6725 ;
  assign n6727 = ~\sa20_reg[1]/P0001  & \sa20_reg[2]/P0001  ;
  assign n6728 = n708 & n736 ;
  assign n6729 = ~n809 & ~n6728 ;
  assign n6730 = ~n703 & n6729 ;
  assign n6731 = n6727 & ~n6730 ;
  assign n6738 = ~n6726 & ~n6731 ;
  assign n6739 = ~n6724 & n6738 ;
  assign n6740 = ~n6720 & n6739 ;
  assign n6741 = ~n6737 & n6740 ;
  assign n6742 = ~n6688 & n6741 ;
  assign n6743 = ~n6714 & n6742 ;
  assign n6744 = \u0_w_reg[2][1]/P0001  & ~n6743 ;
  assign n6745 = ~\u0_w_reg[2][1]/P0001  & n6743 ;
  assign n6746 = ~n6744 & ~n6745 ;
  assign n6747 = n6660 & n6746 ;
  assign n6748 = ~n6660 & ~n6746 ;
  assign n6749 = ~n6747 & ~n6748 ;
  assign n6751 = n6478 & n6749 ;
  assign n6750 = ~n6478 & ~n6749 ;
  assign n6752 = ~\ld_r_reg/P0001  & ~n6750 ;
  assign n6753 = ~n6751 & n6752 ;
  assign n6755 = \text_in_r_reg[33]/P0001  & \u0_w_reg[2][1]/P0001  ;
  assign n6754 = ~\text_in_r_reg[33]/P0001  & ~\u0_w_reg[2][1]/P0001  ;
  assign n6756 = \ld_r_reg/P0001  & ~n6754 ;
  assign n6757 = ~n6755 & n6756 ;
  assign n6758 = ~n6753 & ~n6757 ;
  assign n6787 = \sa31_reg[3]/P0001  & n6488 ;
  assign n6788 = ~n1183 & ~n6787 ;
  assign n6790 = \sa31_reg[7]/P0001  & n5269 ;
  assign n6789 = \sa31_reg[4]/P0001  & n1151 ;
  assign n6791 = ~n6571 & ~n6789 ;
  assign n6792 = ~n6790 & n6791 ;
  assign n6793 = \sa31_reg[2]/P0001  & ~n6792 ;
  assign n6794 = n6788 & ~n6793 ;
  assign n6795 = \sa31_reg[1]/P0001  & ~n6794 ;
  assign n6805 = n1153 & n1178 ;
  assign n6803 = n1159 & ~n1180 ;
  assign n6804 = ~n1256 & n6803 ;
  assign n6806 = n1146 & n5238 ;
  assign n6807 = ~n6110 & ~n6806 ;
  assign n6808 = ~n6804 & n6807 ;
  assign n6809 = ~n6805 & n6808 ;
  assign n6810 = ~\sa31_reg[1]/P0001  & ~n6809 ;
  assign n6796 = n5205 & ~n6136 ;
  assign n6797 = ~n6627 & ~n6796 ;
  assign n6798 = ~\sa31_reg[3]/P0001  & ~n6797 ;
  assign n6799 = ~n1240 & ~n6110 ;
  assign n6800 = ~n6491 & ~n6627 ;
  assign n6801 = n6799 & n6800 ;
  assign n6802 = ~\sa31_reg[2]/P0001  & ~n6801 ;
  assign n6811 = ~n6798 & ~n6802 ;
  assign n6812 = ~n6810 & n6811 ;
  assign n6813 = ~n6795 & n6812 ;
  assign n6814 = \sa31_reg[0]/P0002  & ~n6813 ;
  assign n6763 = ~n1280 & ~n6581 ;
  assign n6764 = \sa31_reg[2]/P0001  & ~n6763 ;
  assign n6759 = \sa31_reg[4]/P0001  & n6483 ;
  assign n6760 = ~n1269 & ~n6530 ;
  assign n6761 = ~n6759 & n6760 ;
  assign n6762 = ~\sa31_reg[2]/P0001  & ~n6761 ;
  assign n6765 = \sa31_reg[1]/P0001  & ~n5204 ;
  assign n6766 = n5272 & n6765 ;
  assign n6767 = ~n6762 & n6766 ;
  assign n6768 = ~n6764 & n6767 ;
  assign n6772 = ~n1154 & ~n1239 ;
  assign n6773 = ~\sa31_reg[2]/P0001  & ~n6772 ;
  assign n6770 = ~n6119 & ~n6491 ;
  assign n6771 = \sa31_reg[2]/P0001  & ~n6770 ;
  assign n6769 = \sa31_reg[6]/NET0131  & n1181 ;
  assign n6774 = ~\sa31_reg[1]/P0001  & ~n6160 ;
  assign n6775 = ~n6769 & n6774 ;
  assign n6776 = ~n6771 & n6775 ;
  assign n6777 = ~n6773 & n6776 ;
  assign n6778 = ~n6768 & ~n6777 ;
  assign n6779 = ~n5250 & n6161 ;
  assign n6780 = \sa31_reg[2]/P0001  & ~n1230 ;
  assign n6781 = ~n1220 & n6780 ;
  assign n6782 = ~n6779 & ~n6781 ;
  assign n6783 = ~n1234 & ~n5295 ;
  assign n6784 = ~n6782 & n6783 ;
  assign n6785 = ~n6778 & n6784 ;
  assign n6786 = ~\sa31_reg[0]/P0002  & ~n6785 ;
  assign n6829 = ~n1168 & ~n1217 ;
  assign n6830 = ~n5253 & n6829 ;
  assign n6831 = ~\sa31_reg[2]/P0001  & ~n6830 ;
  assign n6832 = n1160 & n1182 ;
  assign n6833 = ~n1161 & ~n6832 ;
  assign n6834 = ~n6831 & n6833 ;
  assign n6835 = ~\sa31_reg[1]/P0001  & ~n6834 ;
  assign n6815 = ~\sa31_reg[5]/P0001  & n1269 ;
  assign n6816 = ~n1202 & ~n1234 ;
  assign n6817 = ~n6815 & n6816 ;
  assign n6818 = n6514 & ~n6817 ;
  assign n6824 = ~\sa31_reg[6]/NET0131  & n6644 ;
  assign n6836 = ~n6648 & ~n6824 ;
  assign n6837 = ~n6818 & n6836 ;
  assign n6819 = ~n5204 & ~n6543 ;
  assign n6820 = ~n1195 & n6819 ;
  assign n6821 = ~n1205 & ~n6168 ;
  assign n6822 = n6820 & n6821 ;
  assign n6823 = n1224 & ~n6822 ;
  assign n6825 = ~n1183 & ~n1277 ;
  assign n6826 = \sa31_reg[3]/P0001  & ~n6825 ;
  assign n6827 = ~n6636 & ~n6826 ;
  assign n6828 = n1232 & ~n6827 ;
  assign n6838 = ~n6823 & ~n6828 ;
  assign n6839 = n6837 & n6838 ;
  assign n6840 = ~n6835 & n6839 ;
  assign n6841 = ~n6786 & n6840 ;
  assign n6842 = ~n6814 & n6841 ;
  assign n6843 = \u0_w_reg[2][9]/P0001  & ~n6842 ;
  assign n6844 = ~\u0_w_reg[2][9]/P0001  & n6842 ;
  assign n6845 = ~n6843 & ~n6844 ;
  assign n6846 = n6660 & n6845 ;
  assign n6847 = ~n6660 & ~n6845 ;
  assign n6848 = ~n6846 & ~n6847 ;
  assign n6851 = ~\sa20_reg[3]/P0001  & n820 ;
  assign n6852 = ~n5556 & ~n5907 ;
  assign n6853 = ~n6851 & n6852 ;
  assign n6854 = \sa20_reg[2]/P0001  & ~n6853 ;
  assign n6850 = ~\sa20_reg[2]/P0001  & n5857 ;
  assign n6849 = ~\sa20_reg[4]/P0001  & n706 ;
  assign n6855 = ~n5600 & ~n5895 ;
  assign n6856 = ~n6849 & n6855 ;
  assign n6857 = ~n6850 & n6856 ;
  assign n6858 = ~n6854 & n6857 ;
  assign n6859 = ~\sa20_reg[1]/P0001  & ~n6858 ;
  assign n6860 = ~n746 & ~n5981 ;
  assign n6861 = n5893 & n6860 ;
  assign n6862 = \sa20_reg[2]/P0001  & ~n6861 ;
  assign n6867 = ~\sa20_reg[2]/P0001  & ~n690 ;
  assign n6868 = ~\sa20_reg[5]/P0001  & ~n723 ;
  assign n6869 = n6867 & ~n6868 ;
  assign n6870 = ~n832 & ~n6869 ;
  assign n6871 = \sa20_reg[1]/P0001  & ~n6870 ;
  assign n6863 = ~n5549 & ~n5605 ;
  assign n6864 = ~\sa20_reg[2]/P0001  & ~n6863 ;
  assign n6865 = ~n709 & ~n735 ;
  assign n6866 = n763 & ~n6865 ;
  assign n6872 = ~n5973 & ~n6029 ;
  assign n6873 = ~n6866 & n6872 ;
  assign n6874 = ~n6864 & n6873 ;
  assign n6875 = ~n6871 & n6874 ;
  assign n6876 = ~n6862 & n6875 ;
  assign n6877 = ~n6859 & n6876 ;
  assign n6878 = \sa20_reg[0]/P0001  & ~n6877 ;
  assign n6879 = \sa20_reg[6]/NET0131  & n833 ;
  assign n6880 = ~n5892 & ~n6879 ;
  assign n6881 = ~n800 & n6880 ;
  assign n6882 = ~\sa20_reg[2]/P0001  & ~n6881 ;
  assign n6883 = ~n724 & ~n735 ;
  assign n6884 = \sa20_reg[2]/P0001  & n745 ;
  assign n6885 = ~n6883 & n6884 ;
  assign n6886 = ~n698 & n744 ;
  assign n6887 = n6727 & n6886 ;
  assign n6899 = ~n6885 & ~n6887 ;
  assign n6900 = ~n6882 & n6899 ;
  assign n6888 = ~\sa20_reg[3]/P0001  & ~n5568 ;
  assign n6889 = ~n6007 & ~n6888 ;
  assign n6890 = ~\sa20_reg[1]/P0001  & ~n6889 ;
  assign n6894 = \sa20_reg[2]/P0001  & n698 ;
  assign n6895 = n777 & n6894 ;
  assign n6891 = n720 & n747 ;
  assign n6892 = ~n716 & ~n723 ;
  assign n6893 = ~n6697 & ~n6892 ;
  assign n6896 = ~n6891 & ~n6893 ;
  assign n6897 = ~n6895 & n6896 ;
  assign n6898 = \sa20_reg[1]/P0001  & ~n6897 ;
  assign n6901 = ~n6890 & ~n6898 ;
  assign n6902 = n6900 & n6901 ;
  assign n6903 = ~\sa20_reg[0]/P0001  & ~n6902 ;
  assign n6910 = ~n694 & n5527 ;
  assign n6911 = ~n5968 & ~n6910 ;
  assign n6912 = ~\sa20_reg[2]/P0001  & ~n6911 ;
  assign n6906 = \sa20_reg[2]/P0001  & n799 ;
  assign n6907 = ~n701 & ~n5544 ;
  assign n6908 = n6906 & ~n6907 ;
  assign n6909 = n695 & n763 ;
  assign n6913 = ~\sa20_reg[1]/P0001  & ~n6909 ;
  assign n6914 = ~n5928 & n6913 ;
  assign n6915 = ~n6908 & n6914 ;
  assign n6916 = ~n6912 & n6915 ;
  assign n6918 = ~\sa20_reg[2]/P0001  & ~n5617 ;
  assign n6919 = ~n5836 & ~n6918 ;
  assign n6917 = \sa20_reg[2]/P0001  & n707 ;
  assign n6920 = ~n824 & ~n6917 ;
  assign n6921 = n5996 & n6920 ;
  assign n6922 = ~n6919 & n6921 ;
  assign n6923 = ~n6916 & ~n6922 ;
  assign n6904 = n729 & n5523 ;
  assign n6905 = n5526 & n5973 ;
  assign n6924 = ~n6904 & ~n6905 ;
  assign n6925 = ~n6923 & n6924 ;
  assign n6926 = ~n6903 & n6925 ;
  assign n6927 = ~n6878 & n6926 ;
  assign n6928 = n5631 & ~n6927 ;
  assign n6929 = ~n5631 & n6927 ;
  assign n6930 = ~n6928 & ~n6929 ;
  assign n6931 = n6395 & n6930 ;
  assign n6932 = ~n6395 & ~n6930 ;
  assign n6933 = ~n6931 & ~n6932 ;
  assign n6935 = n6848 & n6933 ;
  assign n6934 = ~n6848 & ~n6933 ;
  assign n6936 = ~\ld_r_reg/P0001  & ~n6934 ;
  assign n6937 = ~n6935 & n6936 ;
  assign n6939 = \text_in_r_reg[41]/P0001  & \u0_w_reg[2][9]/P0001  ;
  assign n6938 = ~\text_in_r_reg[41]/P0001  & ~\u0_w_reg[2][9]/P0001  ;
  assign n6940 = \ld_r_reg/P0001  & ~n6938 ;
  assign n6941 = ~n6939 & n6940 ;
  assign n6942 = ~n6937 & ~n6941 ;
  assign n6943 = ~n1145 & ~n5830 ;
  assign n6944 = n1145 & n5830 ;
  assign n6945 = ~n6943 & ~n6944 ;
  assign n6946 = \u0_w_reg[2][5]/P0001  & ~n6180 ;
  assign n6947 = ~\u0_w_reg[2][5]/P0001  & n6180 ;
  assign n6948 = ~n6946 & ~n6947 ;
  assign n6949 = n5931 & n6948 ;
  assign n6950 = ~n5931 & ~n6948 ;
  assign n6951 = ~n6949 & ~n6950 ;
  assign n6953 = n6945 & n6951 ;
  assign n6952 = ~n6945 & ~n6951 ;
  assign n6954 = ~\ld_r_reg/P0001  & ~n6952 ;
  assign n6955 = ~n6953 & n6954 ;
  assign n6957 = \text_in_r_reg[37]/P0001  & \u0_w_reg[2][5]/P0001  ;
  assign n6956 = ~\text_in_r_reg[37]/P0001  & ~\u0_w_reg[2][5]/P0001  ;
  assign n6958 = \ld_r_reg/P0001  & ~n6956 ;
  assign n6959 = ~n6957 & n6958 ;
  assign n6960 = ~n6955 & ~n6959 ;
  assign n6961 = \u0_w_reg[2][28]/P0001  & ~n6180 ;
  assign n6962 = ~\u0_w_reg[2][28]/P0001  & n6180 ;
  assign n6963 = ~n6961 & ~n6962 ;
  assign n6964 = n6058 & n6963 ;
  assign n6965 = ~n6058 & ~n6963 ;
  assign n6966 = ~n6964 & ~n6965 ;
  assign n7000 = ~n1042 & ~n1062 ;
  assign n7001 = ~n5755 & n7000 ;
  assign n7002 = \sa02_reg[2]/P0001  & ~n7001 ;
  assign n7003 = n994 & ~n1068 ;
  assign n7004 = n1025 & n5108 ;
  assign n7005 = ~n5792 & ~n7004 ;
  assign n7006 = ~n5119 & n7005 ;
  assign n7007 = ~n7003 & n7006 ;
  assign n7008 = ~n7002 & n7007 ;
  assign n7009 = \sa02_reg[1]/P0001  & ~n7008 ;
  assign n6991 = ~n1021 & ~n6364 ;
  assign n6992 = ~\sa02_reg[2]/P0001  & ~n6991 ;
  assign n6994 = ~n1121 & ~n5171 ;
  assign n6995 = ~n5098 & n6994 ;
  assign n6993 = ~n5159 & n5753 ;
  assign n6996 = ~n6377 & ~n6993 ;
  assign n6997 = n6995 & n6996 ;
  assign n6998 = ~n6992 & n6997 ;
  assign n6999 = ~\sa02_reg[1]/P0001  & ~n6998 ;
  assign n6976 = n974 & n1003 ;
  assign n7010 = n6419 & ~n6976 ;
  assign n7011 = ~\sa02_reg[2]/P0001  & ~n7010 ;
  assign n7012 = ~n1024 & n1131 ;
  assign n7013 = n1128 & ~n7012 ;
  assign n7014 = ~n1070 & ~n7013 ;
  assign n7015 = ~n7011 & n7014 ;
  assign n7016 = ~n6999 & n7015 ;
  assign n7017 = ~n7009 & n7016 ;
  assign n7018 = \sa02_reg[0]/P0001  & ~n7017 ;
  assign n6968 = ~n996 & ~n5141 ;
  assign n6969 = \sa02_reg[2]/P0001  & ~n6968 ;
  assign n6967 = ~\sa02_reg[2]/P0001  & n1043 ;
  assign n6970 = ~n977 & ~n5787 ;
  assign n6971 = ~n6337 & n6970 ;
  assign n6972 = ~n6967 & n6971 ;
  assign n6973 = ~n6969 & n6972 ;
  assign n6974 = \sa02_reg[1]/P0001  & ~n6973 ;
  assign n6979 = ~n5182 & ~n6976 ;
  assign n6975 = n1006 & ~n1017 ;
  assign n6977 = \sa02_reg[7]/NET0131  & n978 ;
  assign n6978 = ~n982 & n6977 ;
  assign n6980 = ~n6975 & ~n6978 ;
  assign n6981 = n6979 & n6980 ;
  assign n6982 = ~\sa02_reg[1]/P0001  & ~n6981 ;
  assign n6983 = ~\sa02_reg[2]/P0001  & ~n5080 ;
  assign n6984 = n984 & n996 ;
  assign n6985 = ~n1073 & ~n5173 ;
  assign n6986 = ~n6984 & n6985 ;
  assign n6987 = ~n6983 & n6986 ;
  assign n6988 = ~n6982 & n6987 ;
  assign n6989 = ~n6974 & n6988 ;
  assign n6990 = ~\sa02_reg[0]/P0001  & ~n6989 ;
  assign n7020 = ~n5323 & ~n5767 ;
  assign n7021 = ~n1043 & n7020 ;
  assign n7022 = n5108 & ~n7021 ;
  assign n7019 = ~\sa02_reg[2]/P0001  & n5818 ;
  assign n7023 = ~n5775 & ~n7019 ;
  assign n7024 = ~n7022 & n7023 ;
  assign n7025 = \sa02_reg[1]/P0001  & ~n7024 ;
  assign n7028 = \sa02_reg[6]/NET0131  & n1078 ;
  assign n7029 = ~n5792 & ~n7028 ;
  assign n7030 = n5154 & ~n7029 ;
  assign n7026 = ~n1061 & ~n1073 ;
  assign n7027 = n5106 & ~n7026 ;
  assign n7032 = ~n1005 & ~n5768 ;
  assign n7033 = n984 & ~n7032 ;
  assign n7031 = n5780 & n6363 ;
  assign n7034 = ~n6305 & ~n7031 ;
  assign n7035 = ~n7033 & n7034 ;
  assign n7036 = ~n7027 & n7035 ;
  assign n7037 = ~n7030 & n7036 ;
  assign n7038 = ~n7025 & n7037 ;
  assign n7039 = ~n6990 & n7038 ;
  assign n7040 = ~n7018 & n7039 ;
  assign n7067 = ~n648 & ~n856 ;
  assign n7068 = ~\sa13_reg[2]/P0001  & ~n7067 ;
  assign n7065 = ~n901 & n926 ;
  assign n7066 = \sa13_reg[2]/P0001  & ~n7065 ;
  assign n7069 = ~n654 & ~n668 ;
  assign n7070 = ~n5682 & n7069 ;
  assign n7071 = ~n7066 & n7070 ;
  assign n7072 = ~n7068 & n7071 ;
  assign n7073 = ~\sa13_reg[1]/P0001  & ~n7072 ;
  assign n7074 = ~n568 & ~n920 ;
  assign n7075 = ~n5456 & n7074 ;
  assign n7076 = \sa13_reg[2]/P0001  & ~n7075 ;
  assign n7077 = ~n588 & ~n5425 ;
  assign n7078 = ~n5504 & ~n5671 ;
  assign n7079 = ~n6284 & n7078 ;
  assign n7080 = n7077 & n7079 ;
  assign n7081 = ~n7076 & n7080 ;
  assign n7082 = \sa13_reg[1]/P0001  & ~n7081 ;
  assign n7083 = \sa13_reg[3]/P0001  & n540 ;
  assign n7084 = ~n921 & ~n7083 ;
  assign n7085 = ~n5426 & n7084 ;
  assign n7086 = ~\sa13_reg[2]/P0001  & ~n7085 ;
  assign n7087 = ~n864 & ~n944 ;
  assign n7088 = n6281 & ~n7087 ;
  assign n7089 = ~n911 & ~n7088 ;
  assign n7090 = ~n7086 & n7089 ;
  assign n7091 = ~n7082 & n7090 ;
  assign n7092 = ~n7073 & n7091 ;
  assign n7093 = \sa13_reg[0]/P0001  & ~n7092 ;
  assign n7042 = ~n604 & ~n638 ;
  assign n7043 = \sa13_reg[2]/P0001  & ~n7042 ;
  assign n7044 = ~n551 & ~n5699 ;
  assign n7041 = n532 & n5459 ;
  assign n7045 = ~n6243 & ~n7041 ;
  assign n7046 = n7044 & n7045 ;
  assign n7047 = ~n7043 & n7046 ;
  assign n7048 = \sa13_reg[1]/P0001  & ~n7047 ;
  assign n7053 = n556 & n6281 ;
  assign n7054 = ~n5426 & ~n7053 ;
  assign n7055 = ~n652 & n7054 ;
  assign n7051 = \sa13_reg[7]/NET0131  & ~n547 ;
  assign n7052 = n603 & n7051 ;
  assign n7056 = ~n679 & ~n7052 ;
  assign n7057 = n7055 & n7056 ;
  assign n7058 = ~\sa13_reg[1]/P0001  & ~n7057 ;
  assign n7049 = ~\sa13_reg[2]/P0001  & ~n546 ;
  assign n7050 = n591 & n653 ;
  assign n7059 = ~n671 & ~n5464 ;
  assign n7060 = ~n7050 & n7059 ;
  assign n7061 = ~n7049 & n7060 ;
  assign n7062 = ~n7058 & n7061 ;
  assign n7063 = ~n7048 & n7062 ;
  assign n7064 = ~\sa13_reg[0]/P0001  & ~n7063 ;
  assign n7095 = ~n632 & ~n865 ;
  assign n7096 = ~n569 & n7095 ;
  assign n7097 = n5424 & ~n7096 ;
  assign n7098 = n955 & n5459 ;
  assign n7099 = ~n5647 & ~n7098 ;
  assign n7100 = ~n7097 & n7099 ;
  assign n7101 = \sa13_reg[1]/P0001  & ~n7100 ;
  assign n7102 = ~n918 & ~n7050 ;
  assign n7103 = n6272 & ~n7102 ;
  assign n7104 = \sa13_reg[6]/NET0131  & n656 ;
  assign n7105 = ~n5671 & ~n7104 ;
  assign n7106 = n6286 & ~n7105 ;
  assign n7107 = n962 & n5651 ;
  assign n7094 = n571 & n623 ;
  assign n7108 = ~n649 & ~n6282 ;
  assign n7109 = ~n7094 & n7108 ;
  assign n7110 = ~n7107 & n7109 ;
  assign n7111 = ~n7106 & n7110 ;
  assign n7112 = ~n7103 & n7111 ;
  assign n7113 = ~n7101 & n7112 ;
  assign n7114 = ~n7064 & n7113 ;
  assign n7115 = ~n7093 & n7114 ;
  assign n7116 = n7040 & ~n7115 ;
  assign n7117 = ~n7040 & n7115 ;
  assign n7118 = ~n7116 & ~n7117 ;
  assign n7119 = ~n5519 & n7118 ;
  assign n7120 = n5519 & ~n7118 ;
  assign n7121 = ~n7119 & ~n7120 ;
  assign n7123 = ~n6966 & n7121 ;
  assign n7122 = n6966 & ~n7121 ;
  assign n7124 = ~\ld_r_reg/P0001  & ~n7122 ;
  assign n7125 = ~n7123 & n7124 ;
  assign n7127 = ~\text_in_r_reg[60]/P0001  & \u0_w_reg[2][28]/P0001  ;
  assign n7126 = \text_in_r_reg[60]/P0001  & ~\u0_w_reg[2][28]/P0001  ;
  assign n7128 = \ld_r_reg/P0001  & ~n7126 ;
  assign n7129 = ~n7127 & n7128 ;
  assign n7130 = ~n7125 & ~n7129 ;
  assign n7174 = ~n708 & n736 ;
  assign n7175 = ~n807 & ~n7174 ;
  assign n7176 = \sa20_reg[2]/P0001  & ~n7175 ;
  assign n7177 = ~n808 & ~n825 ;
  assign n7178 = ~n5530 & n7177 ;
  assign n7179 = ~n7176 & n7178 ;
  assign n7180 = ~\sa20_reg[1]/P0001  & ~n7179 ;
  assign n7162 = ~n782 & ~n790 ;
  assign n7163 = \sa20_reg[2]/P0001  & ~n7162 ;
  assign n7165 = ~n707 & ~n5859 ;
  assign n7164 = ~\sa20_reg[2]/P0001  & n740 ;
  assign n7166 = ~n6689 & ~n7164 ;
  assign n7167 = n7165 & n7166 ;
  assign n7168 = ~n7163 & n7167 ;
  assign n7169 = \sa20_reg[1]/P0001  & ~n7168 ;
  assign n7170 = ~\sa20_reg[2]/P0001  & n704 ;
  assign n7171 = ~\sa20_reg[7]/NET0131  & n6849 ;
  assign n7172 = n828 & ~n7171 ;
  assign n7173 = ~n7170 & ~n7172 ;
  assign n7181 = ~n5878 & ~n7173 ;
  assign n7182 = ~n7169 & n7181 ;
  assign n7183 = ~n7180 & n7182 ;
  assign n7184 = ~\sa20_reg[0]/P0001  & ~n7183 ;
  assign n7133 = ~n820 & ~n5527 ;
  assign n7134 = ~\sa20_reg[2]/P0001  & ~n7133 ;
  assign n7135 = ~n715 & ~n795 ;
  assign n7136 = ~n5617 & n7135 ;
  assign n7137 = ~n7134 & n7136 ;
  assign n7138 = \sa20_reg[1]/P0001  & ~n7137 ;
  assign n7131 = ~n5530 & n6880 ;
  assign n7132 = ~\sa20_reg[2]/P0001  & ~n7131 ;
  assign n7157 = ~n5901 & ~n7132 ;
  assign n7158 = ~n7138 & n7157 ;
  assign n7139 = ~n737 & ~n5591 ;
  assign n7140 = ~\sa20_reg[2]/P0001  & ~n7139 ;
  assign n7143 = ~n809 & ~n838 ;
  assign n7144 = ~n6036 & n7143 ;
  assign n7141 = ~n694 & ~n701 ;
  assign n7142 = n5984 & ~n7141 ;
  assign n7145 = ~n6917 & ~n7142 ;
  assign n7146 = n7144 & n7145 ;
  assign n7147 = ~n7140 & n7146 ;
  assign n7148 = ~\sa20_reg[1]/P0001  & ~n7147 ;
  assign n7149 = \sa20_reg[3]/P0001  & n705 ;
  assign n7150 = n5920 & ~n7149 ;
  assign n7151 = \sa20_reg[4]/P0001  & ~n7150 ;
  assign n7152 = ~n5585 & ~n5979 ;
  assign n7153 = ~n6715 & n7152 ;
  assign n7154 = \sa20_reg[1]/P0001  & ~n7153 ;
  assign n7155 = ~n7151 & ~n7154 ;
  assign n7156 = \sa20_reg[2]/P0001  & ~n7155 ;
  assign n7159 = ~n7148 & ~n7156 ;
  assign n7160 = n7158 & n7159 ;
  assign n7161 = \sa20_reg[0]/P0001  & ~n7160 ;
  assign n7188 = ~n740 & ~n791 ;
  assign n7189 = ~n5997 & n7188 ;
  assign n7190 = n747 & ~n7189 ;
  assign n7186 = ~n694 & ~n720 ;
  assign n7187 = n6894 & ~n7186 ;
  assign n7185 = n763 & n5981 ;
  assign n7191 = ~n6008 & ~n7185 ;
  assign n7192 = ~n7187 & n7191 ;
  assign n7193 = ~n7190 & n7192 ;
  assign n7194 = \sa20_reg[1]/P0001  & ~n7193 ;
  assign n7198 = \sa20_reg[2]/P0001  & ~n5878 ;
  assign n7199 = ~n5894 & n7198 ;
  assign n7197 = ~\sa20_reg[2]/P0001  & ~n6005 ;
  assign n7200 = ~\sa20_reg[1]/P0001  & ~n7197 ;
  assign n7201 = ~n7199 & n7200 ;
  assign n7195 = ~n721 & ~n5998 ;
  assign n7196 = n761 & ~n7195 ;
  assign n7202 = ~n822 & ~n7196 ;
  assign n7203 = ~n7201 & n7202 ;
  assign n7204 = ~n7194 & n7203 ;
  assign n7205 = ~n7161 & n7204 ;
  assign n7206 = ~n7184 & n7205 ;
  assign n7207 = n7115 & ~n7206 ;
  assign n7208 = ~n7115 & n7206 ;
  assign n7209 = ~n7207 & ~n7208 ;
  assign n7210 = n5516 & ~n5830 ;
  assign n7211 = ~n5516 & n5830 ;
  assign n7212 = ~n7210 & ~n7211 ;
  assign n7213 = n7209 & n7212 ;
  assign n7214 = ~n7209 & ~n7212 ;
  assign n7215 = ~n7213 & ~n7214 ;
  assign n7216 = ~n5631 & ~n6055 ;
  assign n7217 = n5631 & n6055 ;
  assign n7218 = ~n7216 & ~n7217 ;
  assign n7219 = \u0_w_reg[2][20]/P0001  & ~n6180 ;
  assign n7220 = ~\u0_w_reg[2][20]/P0001  & n6180 ;
  assign n7221 = ~n7219 & ~n7220 ;
  assign n7222 = n7218 & n7221 ;
  assign n7223 = ~n7218 & ~n7221 ;
  assign n7224 = ~n7222 & ~n7223 ;
  assign n7226 = ~n7215 & n7224 ;
  assign n7225 = n7215 & ~n7224 ;
  assign n7227 = ~\ld_r_reg/P0001  & ~n7225 ;
  assign n7228 = ~n7226 & n7227 ;
  assign n7230 = ~\text_in_r_reg[52]/P0001  & \u0_w_reg[2][20]/P0001  ;
  assign n7229 = \text_in_r_reg[52]/P0001  & ~\u0_w_reg[2][20]/P0001  ;
  assign n7231 = \ld_r_reg/P0001  & ~n7229 ;
  assign n7232 = ~n7230 & n7231 ;
  assign n7233 = ~n7228 & ~n7232 ;
  assign n7234 = ~n6180 & ~n6657 ;
  assign n7235 = n6180 & n6657 ;
  assign n7236 = ~n7234 & ~n7235 ;
  assign n7268 = ~n1204 & ~n1261 ;
  assign n7269 = \sa31_reg[2]/P0001  & ~n7268 ;
  assign n7267 = n1147 & n6136 ;
  assign n7270 = ~n1207 & ~n6148 ;
  assign n7271 = ~n7267 & n7270 ;
  assign n7272 = ~n6787 & n7271 ;
  assign n7273 = ~n7269 & n7272 ;
  assign n7274 = \sa31_reg[1]/P0001  & ~n7273 ;
  assign n7276 = \sa31_reg[7]/P0001  & ~n1229 ;
  assign n7277 = n1279 & n7276 ;
  assign n7257 = n1152 & n1182 ;
  assign n7275 = n1186 & n1215 ;
  assign n7278 = ~n7257 & ~n7275 ;
  assign n7279 = ~n1233 & n7278 ;
  assign n7280 = ~n7277 & n7279 ;
  assign n7281 = ~n1223 & n7280 ;
  assign n7282 = ~\sa31_reg[1]/P0001  & ~n7281 ;
  assign n7283 = ~\sa31_reg[2]/P0001  & ~n1203 ;
  assign n7284 = n1204 & n1265 ;
  assign n7285 = ~n1245 & ~n5258 ;
  assign n7286 = ~n7284 & n7285 ;
  assign n7287 = ~n7283 & n7286 ;
  assign n7288 = ~n7282 & n7287 ;
  assign n7289 = ~n7274 & n7288 ;
  assign n7290 = ~\sa31_reg[0]/P0002  & ~n7289 ;
  assign n7239 = ~n1194 & ~n5268 ;
  assign n7240 = ~n1207 & n7239 ;
  assign n7241 = \sa31_reg[2]/P0001  & ~n7240 ;
  assign n7237 = ~n1217 & ~n5206 ;
  assign n7238 = ~\sa31_reg[2]/P0001  & ~n7237 ;
  assign n7242 = ~n1234 & ~n1247 ;
  assign n7243 = ~n6832 & n7242 ;
  assign n7244 = ~n7238 & n7243 ;
  assign n7245 = ~n7241 & n7244 ;
  assign n7246 = ~\sa31_reg[1]/P0001  & ~n7245 ;
  assign n7251 = ~n1219 & ~n6569 ;
  assign n7252 = ~\sa31_reg[2]/P0001  & ~n7251 ;
  assign n7248 = n1178 & ~n1276 ;
  assign n7249 = ~n6092 & ~n7248 ;
  assign n7250 = \sa31_reg[2]/P0001  & ~n7249 ;
  assign n7247 = \sa31_reg[4]/P0001  & n6515 ;
  assign n7253 = ~n6119 & ~n7247 ;
  assign n7254 = ~n7250 & n7253 ;
  assign n7255 = ~n7252 & n7254 ;
  assign n7256 = \sa31_reg[1]/P0001  & ~n7255 ;
  assign n7258 = n6529 & ~n7257 ;
  assign n7259 = ~\sa31_reg[2]/P0001  & ~n7258 ;
  assign n7260 = ~n1206 & n5287 ;
  assign n7261 = n1215 & ~n7260 ;
  assign n7262 = ~n5264 & ~n7261 ;
  assign n7263 = ~n7259 & n7262 ;
  assign n7264 = ~n7256 & n7263 ;
  assign n7265 = ~n7246 & n7264 ;
  assign n7266 = \sa31_reg[0]/P0002  & ~n7265 ;
  assign n7294 = \sa31_reg[6]/NET0131  & n5263 ;
  assign n7295 = ~n6119 & ~n7294 ;
  assign n7296 = \sa31_reg[2]/P0001  & ~n7295 ;
  assign n7291 = ~n5199 & ~n6598 ;
  assign n7292 = ~n1148 & n7291 ;
  assign n7293 = n1162 & ~n7292 ;
  assign n7297 = ~\sa31_reg[6]/NET0131  & n6584 ;
  assign n7298 = ~n6135 & ~n7297 ;
  assign n7299 = ~n7293 & n7298 ;
  assign n7300 = ~n7296 & n7299 ;
  assign n7301 = \sa31_reg[1]/P0001  & ~n7300 ;
  assign n7302 = ~n1233 & ~n6110 ;
  assign n7303 = n1279 & ~n7302 ;
  assign n7304 = n6136 & n6790 ;
  assign n7305 = ~n7303 & ~n7304 ;
  assign n7306 = ~\sa31_reg[1]/P0001  & ~n7305 ;
  assign n7307 = ~n1183 & ~n6124 ;
  assign n7308 = n1265 & ~n7307 ;
  assign n7309 = ~n6769 & ~n7308 ;
  assign n7310 = ~n7306 & n7309 ;
  assign n7311 = ~n7301 & n7310 ;
  assign n7312 = ~n7266 & n7311 ;
  assign n7313 = ~n7290 & n7312 ;
  assign n7314 = \u0_w_reg[2][12]/P0001  & ~n7313 ;
  assign n7315 = ~\u0_w_reg[2][12]/P0001  & n7313 ;
  assign n7316 = ~n7314 & ~n7315 ;
  assign n7317 = n7236 & n7316 ;
  assign n7318 = ~n7236 & ~n7316 ;
  assign n7319 = ~n7317 & ~n7318 ;
  assign n7320 = n5631 & ~n7206 ;
  assign n7321 = ~n5631 & n7206 ;
  assign n7322 = ~n7320 & ~n7321 ;
  assign n7323 = ~n5833 & n7322 ;
  assign n7324 = n5833 & ~n7322 ;
  assign n7325 = ~n7323 & ~n7324 ;
  assign n7327 = n7319 & n7325 ;
  assign n7326 = ~n7319 & ~n7325 ;
  assign n7328 = ~\ld_r_reg/P0001  & ~n7326 ;
  assign n7329 = ~n7327 & n7328 ;
  assign n7331 = ~\text_in_r_reg[44]/P0001  & \u0_w_reg[2][12]/P0001  ;
  assign n7330 = \text_in_r_reg[44]/P0001  & ~\u0_w_reg[2][12]/P0001  ;
  assign n7332 = \ld_r_reg/P0001  & ~n7330 ;
  assign n7333 = ~n7331 & n7332 ;
  assign n7334 = ~n7329 & ~n7333 ;
  assign n7339 = ~n651 & ~n913 ;
  assign n7340 = ~n858 & n7339 ;
  assign n7341 = \sa13_reg[2]/P0001  & ~n7340 ;
  assign n7337 = \sa13_reg[4]/P0001  & n5446 ;
  assign n7335 = \sa13_reg[5]/P0001  & ~n549 ;
  assign n7336 = n655 & ~n7335 ;
  assign n7338 = n653 & n900 ;
  assign n7342 = ~n7336 & ~n7338 ;
  assign n7343 = ~n7337 & n7342 ;
  assign n7344 = ~n7341 & n7343 ;
  assign n7345 = ~\sa13_reg[1]/P0001  & ~n7344 ;
  assign n7353 = ~n535 & ~n650 ;
  assign n7354 = ~\sa13_reg[2]/P0001  & ~n7353 ;
  assign n7355 = ~n665 & ~n7354 ;
  assign n7356 = \sa13_reg[1]/P0001  & ~n7355 ;
  assign n7346 = ~n921 & ~n5679 ;
  assign n7347 = n562 & n7346 ;
  assign n7348 = \sa13_reg[2]/P0001  & ~n7347 ;
  assign n7349 = ~n907 & ~n5438 ;
  assign n7350 = ~\sa13_reg[2]/P0001  & ~n7349 ;
  assign n7351 = ~n536 & ~n912 ;
  assign n7352 = n581 & ~n7351 ;
  assign n7357 = ~n862 & ~n5704 ;
  assign n7358 = ~n7352 & n7357 ;
  assign n7359 = ~n7350 & n7358 ;
  assign n7360 = ~n7348 & n7359 ;
  assign n7361 = ~n7356 & n7360 ;
  assign n7362 = ~n7345 & n7361 ;
  assign n7363 = \sa13_reg[0]/P0001  & ~n7362 ;
  assign n7373 = n570 & n5424 ;
  assign n7374 = \sa13_reg[1]/P0001  & ~n5442 ;
  assign n7375 = ~n7373 & n7374 ;
  assign n7370 = ~n555 & ~n556 ;
  assign n7371 = ~n635 & ~n7370 ;
  assign n7372 = n623 & n861 ;
  assign n7376 = ~n7371 & ~n7372 ;
  assign n7377 = n7375 & n7376 ;
  assign n7378 = ~\sa13_reg[3]/P0001  & ~n5487 ;
  assign n7379 = ~\sa13_reg[1]/P0001  & ~n5649 ;
  assign n7380 = ~n7378 & n7379 ;
  assign n7381 = ~n7377 & ~n7380 ;
  assign n7364 = ~n642 & n7084 ;
  assign n7365 = ~\sa13_reg[2]/P0001  & ~n7364 ;
  assign n7366 = ~n557 & ~n912 ;
  assign n7367 = n883 & ~n7366 ;
  assign n7368 = ~n568 & ~n963 ;
  assign n7369 = n6272 & ~n7368 ;
  assign n7382 = ~n7367 & ~n7369 ;
  assign n7383 = ~n7365 & n7382 ;
  assign n7384 = ~n7381 & n7383 ;
  assign n7385 = ~\sa13_reg[0]/P0001  & ~n7384 ;
  assign n7392 = \sa13_reg[4]/P0001  & n877 ;
  assign n7393 = ~n551 & ~n7392 ;
  assign n7394 = \sa13_reg[2]/P0001  & ~n7393 ;
  assign n7391 = ~\sa13_reg[2]/P0001  & n5504 ;
  assign n7395 = ~n683 & ~n7391 ;
  assign n7396 = n5657 & n7395 ;
  assign n7397 = ~n7394 & n7396 ;
  assign n7398 = ~n877 & ~n911 ;
  assign n7399 = ~n5422 & ~n5678 ;
  assign n7400 = n7398 & n7399 ;
  assign n7401 = ~\sa13_reg[2]/P0001  & ~n7400 ;
  assign n7402 = ~\sa13_reg[1]/P0001  & ~n953 ;
  assign n7403 = ~n7401 & n7402 ;
  assign n7404 = ~n7397 & ~n7403 ;
  assign n7386 = ~n668 & ~n5680 ;
  assign n7387 = n6272 & ~n7386 ;
  assign n7388 = n603 & n901 ;
  assign n7389 = ~n625 & ~n7388 ;
  assign n7390 = \sa13_reg[6]/NET0131  & ~n7389 ;
  assign n7405 = ~n7387 & ~n7390 ;
  assign n7406 = ~n7404 & n7405 ;
  assign n7407 = ~n7385 & n7406 ;
  assign n7408 = ~n7363 & n7407 ;
  assign n7409 = n5516 & ~n7408 ;
  assign n7410 = ~n5516 & n7408 ;
  assign n7411 = ~n7409 & ~n7410 ;
  assign n7412 = n6392 & ~n6927 ;
  assign n7413 = ~n6392 & n6927 ;
  assign n7414 = ~n7412 & ~n7413 ;
  assign n7415 = n7411 & n7414 ;
  assign n7416 = ~n7411 & ~n7414 ;
  assign n7417 = ~n7415 & ~n7416 ;
  assign n7418 = ~\u0_w_reg[2][17]/P0001  & ~n6842 ;
  assign n7419 = \u0_w_reg[2][17]/P0001  & n6842 ;
  assign n7420 = ~n7418 & ~n7419 ;
  assign n7421 = n5631 & ~n6743 ;
  assign n7422 = ~n5631 & n6743 ;
  assign n7423 = ~n7421 & ~n7422 ;
  assign n7424 = n7420 & n7423 ;
  assign n7425 = ~n7420 & ~n7423 ;
  assign n7426 = ~n7424 & ~n7425 ;
  assign n7428 = n7417 & n7426 ;
  assign n7427 = ~n7417 & ~n7426 ;
  assign n7429 = ~\ld_r_reg/P0001  & ~n7427 ;
  assign n7430 = ~n7428 & n7429 ;
  assign n7432 = \text_in_r_reg[49]/P0001  & \u0_w_reg[2][17]/P0001  ;
  assign n7431 = ~\text_in_r_reg[49]/P0001  & ~\u0_w_reg[2][17]/P0001  ;
  assign n7433 = \ld_r_reg/P0001  & ~n7431 ;
  assign n7434 = ~n7432 & n7433 ;
  assign n7435 = ~n7430 & ~n7434 ;
  assign n7447 = ~n540 & ~n665 ;
  assign n7448 = ~n5466 & n7447 ;
  assign n7449 = \sa13_reg[3]/P0001  & ~n7448 ;
  assign n7446 = \sa13_reg[1]/P0001  & n672 ;
  assign n7450 = ~n862 & ~n7446 ;
  assign n7451 = ~n7449 & n7450 ;
  assign n7452 = \sa13_reg[2]/P0001  & ~n7451 ;
  assign n7441 = ~n589 & ~n5651 ;
  assign n7442 = ~n5725 & n7441 ;
  assign n7436 = ~n654 & ~n913 ;
  assign n7437 = ~\sa13_reg[2]/P0001  & ~n7436 ;
  assign n7438 = n543 & n603 ;
  assign n7439 = ~n5661 & ~n7338 ;
  assign n7440 = ~n7438 & n7439 ;
  assign n7443 = ~n7437 & n7440 ;
  assign n7444 = n7442 & n7443 ;
  assign n7445 = ~\sa13_reg[1]/P0001  & ~n7444 ;
  assign n7453 = ~n620 & ~n632 ;
  assign n7454 = ~n911 & n7453 ;
  assign n7455 = n680 & ~n7454 ;
  assign n7456 = ~n5678 & ~n5680 ;
  assign n7457 = ~n7455 & n7456 ;
  assign n7458 = ~n7445 & n7457 ;
  assign n7459 = ~n7452 & n7458 ;
  assign n7460 = \sa13_reg[0]/P0001  & ~n7459 ;
  assign n7485 = \sa13_reg[2]/P0001  & ~n5442 ;
  assign n7486 = ~n903 & n7485 ;
  assign n7487 = ~\sa13_reg[2]/P0001  & ~n604 ;
  assign n7488 = ~n5650 & ~n6216 ;
  assign n7489 = n7487 & n7488 ;
  assign n7490 = ~n7486 & ~n7489 ;
  assign n7491 = ~n5476 & ~n7490 ;
  assign n7492 = \sa13_reg[1]/P0001  & ~n7491 ;
  assign n7493 = ~\sa13_reg[1]/P0001  & n900 ;
  assign n7494 = ~n5492 & ~n7493 ;
  assign n7495 = n581 & ~n7494 ;
  assign n7497 = ~\sa13_reg[1]/P0001  & n5504 ;
  assign n7496 = n5671 & n6281 ;
  assign n7498 = ~n588 & ~n7496 ;
  assign n7499 = ~n7497 & n7498 ;
  assign n7500 = ~n7495 & n7499 ;
  assign n7501 = ~n7492 & n7500 ;
  assign n7502 = ~\sa13_reg[0]/P0001  & ~n7501 ;
  assign n7461 = ~n609 & ~n669 ;
  assign n7462 = ~n5492 & n7461 ;
  assign n7463 = n590 & n7462 ;
  assign n7464 = \sa13_reg[2]/P0001  & ~n955 ;
  assign n7465 = ~n5504 & n7464 ;
  assign n7466 = ~n5687 & n7465 ;
  assign n7467 = ~n7463 & ~n7466 ;
  assign n7468 = ~n533 & ~n536 ;
  assign n7469 = n547 & n7468 ;
  assign n7470 = ~n7467 & ~n7469 ;
  assign n7471 = ~\sa13_reg[1]/P0001  & ~n7470 ;
  assign n7472 = ~\sa13_reg[6]/NET0131  & n884 ;
  assign n7473 = n6244 & ~n7472 ;
  assign n7474 = ~\sa13_reg[2]/P0001  & ~n7473 ;
  assign n7475 = ~n856 & ~n7474 ;
  assign n7476 = \sa13_reg[1]/P0001  & ~n7475 ;
  assign n7479 = ~n557 & ~n570 ;
  assign n7480 = n653 & ~n7479 ;
  assign n7481 = ~n913 & ~n6252 ;
  assign n7482 = \sa13_reg[1]/P0001  & ~n7481 ;
  assign n7483 = ~n7480 & ~n7482 ;
  assign n7484 = \sa13_reg[2]/P0001  & ~n7483 ;
  assign n7477 = \sa13_reg[2]/P0001  & n6283 ;
  assign n7478 = n908 & n7477 ;
  assign n7503 = ~n7098 & ~n7478 ;
  assign n7504 = ~n7484 & n7503 ;
  assign n7505 = ~n7476 & n7504 ;
  assign n7506 = ~n7471 & n7505 ;
  assign n7507 = ~n7502 & n7506 ;
  assign n7508 = ~n7460 & n7507 ;
  assign n7524 = ~n5092 & ~n5754 ;
  assign n7525 = ~n5809 & n7524 ;
  assign n7520 = ~n1076 & ~n1121 ;
  assign n7521 = ~\sa02_reg[2]/P0001  & ~n7520 ;
  assign n7522 = ~n1113 & ~n5766 ;
  assign n7523 = ~n5780 & n7522 ;
  assign n7526 = ~n7521 & n7523 ;
  assign n7527 = n7525 & n7526 ;
  assign n7528 = ~\sa02_reg[1]/P0001  & ~n7527 ;
  assign n7509 = ~n1068 & n5348 ;
  assign n7510 = ~n1070 & ~n7509 ;
  assign n7511 = ~\sa02_reg[2]/P0001  & ~n7510 ;
  assign n7512 = ~n5169 & ~n7511 ;
  assign n7513 = \sa02_reg[1]/P0001  & ~n7512 ;
  assign n7514 = ~n976 & ~n5363 ;
  assign n7515 = ~n5163 & n7514 ;
  assign n7516 = n984 & ~n7515 ;
  assign n7517 = ~n5394 & ~n5750 ;
  assign n7518 = ~n5754 & n7517 ;
  assign n7519 = ~\sa02_reg[3]/P0001  & ~n7518 ;
  assign n7529 = ~n7516 & ~n7519 ;
  assign n7530 = ~n7513 & n7529 ;
  assign n7531 = ~n7528 & n7530 ;
  assign n7532 = \sa02_reg[0]/P0001  & ~n7531 ;
  assign n7559 = ~\sa02_reg[2]/P0001  & ~n5167 ;
  assign n7560 = ~n5092 & n7559 ;
  assign n7561 = ~n5122 & ~n5394 ;
  assign n7562 = n7560 & n7561 ;
  assign n7563 = \sa02_reg[2]/P0001  & ~n1036 ;
  assign n7564 = ~n5409 & n7563 ;
  assign n7565 = ~n5805 & n7564 ;
  assign n7566 = ~n7562 & ~n7565 ;
  assign n7557 = ~\sa02_reg[6]/NET0131  & ~n986 ;
  assign n7558 = n6339 & n7557 ;
  assign n7567 = ~\sa02_reg[1]/P0001  & ~n7558 ;
  assign n7568 = ~n7566 & n7567 ;
  assign n7569 = \sa02_reg[4]/P0001  & n6312 ;
  assign n7570 = n6338 & ~n7569 ;
  assign n7571 = ~\sa02_reg[2]/P0001  & ~n7570 ;
  assign n7572 = \sa02_reg[1]/P0001  & ~n1021 ;
  assign n7573 = ~n7571 & n7572 ;
  assign n7574 = ~n7568 & ~n7573 ;
  assign n7533 = ~n1069 & ~n5155 ;
  assign n7534 = \sa02_reg[2]/P0001  & ~n7533 ;
  assign n7535 = ~n1015 & ~n1068 ;
  assign n7536 = ~\sa02_reg[2]/P0001  & ~n1056 ;
  assign n7537 = ~n7535 & n7536 ;
  assign n7538 = ~n5156 & ~n7537 ;
  assign n7539 = ~n7534 & n7538 ;
  assign n7540 = \sa02_reg[1]/P0001  & ~n7539 ;
  assign n7542 = ~\sa02_reg[1]/P0001  & n5127 ;
  assign n7543 = ~n1110 & ~n7542 ;
  assign n7544 = ~\sa02_reg[2]/P0001  & ~n7543 ;
  assign n7545 = \sa02_reg[2]/P0001  & n5338 ;
  assign n7541 = n986 & n6434 ;
  assign n7546 = ~n1001 & ~n7541 ;
  assign n7547 = ~n7545 & n7546 ;
  assign n7548 = ~n7544 & n7547 ;
  assign n7549 = ~n7540 & n7548 ;
  assign n7550 = ~\sa02_reg[0]/P0001  & ~n7549 ;
  assign n7553 = \sa02_reg[1]/P0001  & n984 ;
  assign n7554 = n1072 & n7553 ;
  assign n7575 = ~n7019 & ~n7554 ;
  assign n7551 = ~n1076 & ~n1122 ;
  assign n7552 = n5154 & ~n7551 ;
  assign n7555 = ~n1003 & ~n5091 ;
  assign n7556 = n5342 & ~n7555 ;
  assign n7576 = ~n7552 & ~n7556 ;
  assign n7577 = n7575 & n7576 ;
  assign n7578 = ~n7550 & n7577 ;
  assign n7579 = ~n7574 & n7578 ;
  assign n7580 = ~n7532 & n7579 ;
  assign n7581 = n7508 & ~n7580 ;
  assign n7582 = ~n7508 & n7580 ;
  assign n7583 = ~n7581 & ~n7582 ;
  assign n7584 = ~n6392 & ~n7583 ;
  assign n7585 = n6392 & n7583 ;
  assign n7586 = ~n7584 & ~n7585 ;
  assign n7613 = ~n809 & ~n5907 ;
  assign n7614 = ~\sa20_reg[2]/P0001  & ~n7613 ;
  assign n7616 = ~n5600 & ~n5985 ;
  assign n7615 = n693 & n819 ;
  assign n7617 = ~n6001 & ~n7615 ;
  assign n7618 = n7616 & n7617 ;
  assign n7619 = ~n725 & n6006 ;
  assign n7620 = n7618 & n7619 ;
  assign n7621 = ~n7614 & n7620 ;
  assign n7623 = n6663 & n6867 ;
  assign n7622 = n723 & n5526 ;
  assign n7624 = \sa20_reg[1]/P0001  & ~n7622 ;
  assign n7625 = ~n6909 & n7624 ;
  assign n7626 = ~n7623 & n7625 ;
  assign n7627 = ~n7621 & ~n7626 ;
  assign n7610 = ~n832 & ~n5858 ;
  assign n7611 = ~n5606 & n7610 ;
  assign n7612 = n761 & ~n7611 ;
  assign n7628 = ~n809 & ~n7615 ;
  assign n7629 = \sa20_reg[5]/P0001  & ~n7628 ;
  assign n7630 = \sa20_reg[0]/P0001  & ~n6037 ;
  assign n7631 = ~n7629 & n7630 ;
  assign n7632 = ~n7612 & n7631 ;
  assign n7633 = ~n7627 & n7632 ;
  assign n7640 = ~n5552 & ~n5872 ;
  assign n7641 = \sa20_reg[2]/P0001  & ~n7640 ;
  assign n7642 = n5590 & ~n7641 ;
  assign n7643 = n763 & n777 ;
  assign n7644 = ~\sa20_reg[1]/P0001  & ~n5617 ;
  assign n7645 = ~n7643 & n7644 ;
  assign n7646 = ~n7642 & ~n7645 ;
  assign n7634 = ~n698 & ~n709 ;
  assign n7635 = \sa20_reg[1]/P0001  & ~n777 ;
  assign n7636 = ~\sa20_reg[2]/P0001  & ~n7635 ;
  assign n7637 = ~n7634 & ~n7636 ;
  assign n7638 = ~n817 & ~n7637 ;
  assign n7639 = ~n5618 & ~n7638 ;
  assign n7647 = ~\sa20_reg[0]/P0001  & ~n715 ;
  assign n7648 = ~n7639 & n7647 ;
  assign n7649 = ~n7646 & n7648 ;
  assign n7650 = ~n7633 & ~n7649 ;
  assign n7592 = ~\sa20_reg[2]/P0001  & ~n839 ;
  assign n7593 = ~n5573 & n7592 ;
  assign n7594 = ~n725 & ~n779 ;
  assign n7595 = n7593 & n7594 ;
  assign n7596 = \sa20_reg[2]/P0001  & ~n5617 ;
  assign n7597 = ~n5619 & n7596 ;
  assign n7598 = ~n6043 & n7597 ;
  assign n7599 = ~n7595 & ~n7598 ;
  assign n7600 = ~n691 & n708 ;
  assign n7601 = ~n709 & n7600 ;
  assign n7602 = ~n7599 & ~n7601 ;
  assign n7603 = ~\sa20_reg[1]/P0001  & ~n7602 ;
  assign n7587 = \sa20_reg[4]/P0001  & n769 ;
  assign n7588 = n6690 & ~n7587 ;
  assign n7589 = ~\sa20_reg[2]/P0001  & ~n7588 ;
  assign n7590 = ~n737 & ~n7589 ;
  assign n7591 = \sa20_reg[1]/P0001  & ~n7590 ;
  assign n7604 = ~n736 & ~n5591 ;
  assign n7605 = ~\sa20_reg[4]/P0001  & ~n7604 ;
  assign n7606 = ~n5907 & ~n7605 ;
  assign n7607 = n806 & ~n7606 ;
  assign n7608 = ~n720 & ~n724 ;
  assign n7609 = n6906 & ~n7608 ;
  assign n7651 = ~n7185 & ~n7609 ;
  assign n7652 = ~n7607 & n7651 ;
  assign n7653 = ~n7591 & n7652 ;
  assign n7654 = ~n7603 & n7653 ;
  assign n7655 = ~n7650 & n7654 ;
  assign n7656 = \u0_w_reg[2][2]/P0001  & ~n7655 ;
  assign n7657 = ~\u0_w_reg[2][2]/P0001  & n7655 ;
  assign n7658 = ~n7656 & ~n7657 ;
  assign n7659 = n6842 & n7658 ;
  assign n7660 = ~n6842 & ~n7658 ;
  assign n7661 = ~n7659 & ~n7660 ;
  assign n7663 = n7586 & ~n7661 ;
  assign n7662 = ~n7586 & n7661 ;
  assign n7664 = ~\ld_r_reg/P0001  & ~n7662 ;
  assign n7665 = ~n7663 & n7664 ;
  assign n7667 = \text_in_r_reg[34]/P0001  & \u0_w_reg[2][2]/P0001  ;
  assign n7666 = ~\text_in_r_reg[34]/P0001  & ~\u0_w_reg[2][2]/P0001  ;
  assign n7668 = \ld_r_reg/P0001  & ~n7666 ;
  assign n7669 = ~n7667 & n7668 ;
  assign n7670 = ~n7665 & ~n7669 ;
  assign n7671 = ~n6304 & n6743 ;
  assign n7672 = n6304 & ~n6743 ;
  assign n7673 = ~n7671 & ~n7672 ;
  assign n7674 = \u0_w_reg[2][25]/P0001  & ~n6842 ;
  assign n7675 = ~\u0_w_reg[2][25]/P0001  & n6842 ;
  assign n7676 = ~n7674 & ~n7675 ;
  assign n7677 = n7673 & n7676 ;
  assign n7678 = ~n7673 & ~n7676 ;
  assign n7679 = ~n7677 & ~n7678 ;
  assign n7680 = n6475 & n7411 ;
  assign n7681 = ~n6475 & ~n7411 ;
  assign n7682 = ~n7680 & ~n7681 ;
  assign n7684 = n7679 & n7682 ;
  assign n7683 = ~n7679 & ~n7682 ;
  assign n7685 = ~\ld_r_reg/P0001  & ~n7683 ;
  assign n7686 = ~n7684 & n7685 ;
  assign n7688 = \text_in_r_reg[57]/P0001  & \u0_w_reg[2][25]/P0001  ;
  assign n7687 = ~\text_in_r_reg[57]/P0001  & ~\u0_w_reg[2][25]/P0001  ;
  assign n7689 = \ld_r_reg/P0001  & ~n7687 ;
  assign n7690 = ~n7688 & n7689 ;
  assign n7691 = ~n7686 & ~n7690 ;
  assign n7692 = ~n850 & ~n5519 ;
  assign n7693 = n850 & n5519 ;
  assign n7694 = ~n7692 & ~n7693 ;
  assign n7695 = \u0_w_reg[2][15]/P0001  & ~n6657 ;
  assign n7696 = ~\u0_w_reg[2][15]/P0001  & n6657 ;
  assign n7697 = ~n7695 & ~n7696 ;
  assign n7698 = n1300 & n7697 ;
  assign n7699 = ~n1300 & ~n7697 ;
  assign n7700 = ~n7698 & ~n7699 ;
  assign n7702 = n7694 & n7700 ;
  assign n7701 = ~n7694 & ~n7700 ;
  assign n7703 = ~\ld_r_reg/P0001  & ~n7701 ;
  assign n7704 = ~n7702 & n7703 ;
  assign n7706 = ~\text_in_r_reg[47]/P0001  & \u0_w_reg[2][15]/P0001  ;
  assign n7705 = \text_in_r_reg[47]/P0001  & ~\u0_w_reg[2][15]/P0001  ;
  assign n7707 = \ld_r_reg/P0001  & ~n7705 ;
  assign n7708 = ~n7706 & n7707 ;
  assign n7709 = ~n7704 & ~n7708 ;
  assign n7710 = n5417 & ~n7040 ;
  assign n7711 = ~n5417 & n7040 ;
  assign n7712 = ~n7710 & ~n7711 ;
  assign n7713 = n5833 & n7712 ;
  assign n7714 = ~n5833 & ~n7712 ;
  assign n7715 = ~n7713 & ~n7714 ;
  assign n7716 = ~n6055 & ~n6657 ;
  assign n7717 = n6055 & n6657 ;
  assign n7718 = ~n7716 & ~n7717 ;
  assign n7719 = \u0_w_reg[2][4]/P0001  & ~n7313 ;
  assign n7720 = ~\u0_w_reg[2][4]/P0001  & n7313 ;
  assign n7721 = ~n7719 & ~n7720 ;
  assign n7722 = n7718 & n7721 ;
  assign n7723 = ~n7718 & ~n7721 ;
  assign n7724 = ~n7722 & ~n7723 ;
  assign n7726 = ~n7715 & n7724 ;
  assign n7725 = n7715 & ~n7724 ;
  assign n7727 = ~\ld_r_reg/P0001  & ~n7725 ;
  assign n7728 = ~n7726 & n7727 ;
  assign n7730 = ~\text_in_r_reg[36]/P0001  & \u0_w_reg[2][4]/P0001  ;
  assign n7729 = \text_in_r_reg[36]/P0001  & ~\u0_w_reg[2][4]/P0001  ;
  assign n7731 = \ld_r_reg/P0001  & ~n7729 ;
  assign n7732 = ~n7730 & n7731 ;
  assign n7733 = ~n7728 & ~n7732 ;
  assign n7734 = \u0_w_reg[2][27]/P0001  & ~n7313 ;
  assign n7735 = ~\u0_w_reg[2][27]/P0001  & n7313 ;
  assign n7736 = ~n7734 & ~n7735 ;
  assign n7737 = n7209 & n7736 ;
  assign n7738 = ~n7209 & ~n7736 ;
  assign n7739 = ~n7737 & ~n7738 ;
  assign n7740 = ~n5519 & n7583 ;
  assign n7741 = n5519 & ~n7583 ;
  assign n7742 = ~n7740 & ~n7741 ;
  assign n7744 = ~n7739 & n7742 ;
  assign n7743 = n7739 & ~n7742 ;
  assign n7745 = ~\ld_r_reg/P0001  & ~n7743 ;
  assign n7746 = ~n7744 & n7745 ;
  assign n7748 = ~\text_in_r_reg[59]/P0001  & \u0_w_reg[2][27]/P0001  ;
  assign n7747 = \text_in_r_reg[59]/P0001  & ~\u0_w_reg[2][27]/P0001  ;
  assign n7749 = \ld_r_reg/P0001  & ~n7747 ;
  assign n7750 = ~n7748 & n7749 ;
  assign n7751 = ~n7746 & ~n7750 ;
  assign n7752 = \u0_w_reg[2][19]/P0001  & ~n7313 ;
  assign n7753 = ~\u0_w_reg[2][19]/P0001  & n7313 ;
  assign n7754 = ~n7752 & ~n7753 ;
  assign n7755 = n7322 & n7754 ;
  assign n7756 = ~n7322 & ~n7754 ;
  assign n7757 = ~n7755 & ~n7756 ;
  assign n7758 = n7508 & ~n7655 ;
  assign n7759 = ~n7508 & n7655 ;
  assign n7760 = ~n7758 & ~n7759 ;
  assign n7761 = n5516 & ~n7040 ;
  assign n7762 = ~n5516 & n7040 ;
  assign n7763 = ~n7761 & ~n7762 ;
  assign n7764 = n7760 & n7763 ;
  assign n7765 = ~n7760 & ~n7763 ;
  assign n7766 = ~n7764 & ~n7765 ;
  assign n7768 = n7757 & n7766 ;
  assign n7767 = ~n7757 & ~n7766 ;
  assign n7769 = ~\ld_r_reg/P0001  & ~n7767 ;
  assign n7770 = ~n7768 & n7769 ;
  assign n7772 = ~\text_in_r_reg[51]/P0001  & \u0_w_reg[2][19]/P0001  ;
  assign n7771 = \text_in_r_reg[51]/P0001  & ~\u0_w_reg[2][19]/P0001  ;
  assign n7773 = \ld_r_reg/P0001  & ~n7771 ;
  assign n7774 = ~n7772 & n7773 ;
  assign n7775 = ~n7770 & ~n7774 ;
  assign n7776 = n5631 & ~n7655 ;
  assign n7777 = ~n5631 & n7655 ;
  assign n7778 = ~n7776 & ~n7777 ;
  assign n7779 = n7118 & n7778 ;
  assign n7780 = ~n7118 & ~n7778 ;
  assign n7781 = ~n7779 & ~n7780 ;
  assign n7811 = n6136 & n6599 ;
  assign n7816 = ~n6087 & ~n6168 ;
  assign n7817 = ~n7811 & n7816 ;
  assign n7813 = ~n6134 & ~n6146 ;
  assign n7814 = ~n6499 & n7813 ;
  assign n7812 = ~\sa31_reg[1]/P0001  & ~n6127 ;
  assign n7815 = ~n5262 & n7812 ;
  assign n7818 = n7814 & n7815 ;
  assign n7819 = n7817 & n7818 ;
  assign n7821 = ~n5269 & n6573 ;
  assign n7822 = ~n5264 & ~n7821 ;
  assign n7823 = ~\sa31_reg[2]/P0001  & ~n7822 ;
  assign n7820 = \sa31_reg[2]/P0001  & n5220 ;
  assign n7824 = \sa31_reg[1]/P0001  & ~n7820 ;
  assign n7825 = ~n7823 & n7824 ;
  assign n7826 = ~n7819 & ~n7825 ;
  assign n7808 = ~n1201 & ~n1239 ;
  assign n7809 = ~n6627 & n7808 ;
  assign n7810 = n1265 & ~n7809 ;
  assign n7827 = n1194 & n1279 ;
  assign n7828 = \sa31_reg[0]/P0002  & ~n6159 ;
  assign n7829 = ~n7827 & n7828 ;
  assign n7830 = ~n6540 & n7829 ;
  assign n7831 = ~n7810 & n7830 ;
  assign n7832 = ~n7826 & n7831 ;
  assign n7833 = \sa31_reg[2]/P0001  & ~n5271 ;
  assign n7834 = ~n6599 & n7833 ;
  assign n7835 = ~n1158 & n5269 ;
  assign n7836 = ~\sa31_reg[2]/P0001  & ~n1204 ;
  assign n7837 = ~n7835 & n7836 ;
  assign n7838 = ~n7834 & ~n7837 ;
  assign n7839 = n6635 & ~n7838 ;
  assign n7840 = n1158 & n5238 ;
  assign n7841 = ~\sa31_reg[1]/P0001  & ~n6556 ;
  assign n7842 = ~n7840 & n7841 ;
  assign n7843 = ~n7839 & ~n7842 ;
  assign n7845 = ~\sa31_reg[2]/P0001  & n1227 ;
  assign n7844 = \sa31_reg[2]/P0001  & n6153 ;
  assign n7846 = ~\sa31_reg[0]/P0002  & ~n1179 ;
  assign n7847 = ~n7844 & n7846 ;
  assign n7848 = ~n7845 & n7847 ;
  assign n7849 = ~n7843 & n7848 ;
  assign n7850 = ~n7832 & ~n7849 ;
  assign n7786 = ~n1246 & ~n6084 ;
  assign n7787 = ~n6168 & n7786 ;
  assign n7788 = n6631 & n7787 ;
  assign n7789 = ~\sa31_reg[6]/NET0131  & n1216 ;
  assign n7790 = \sa31_reg[2]/P0001  & ~n6556 ;
  assign n7791 = ~n7789 & n7790 ;
  assign n7792 = ~n6160 & n7791 ;
  assign n7793 = ~n7788 & ~n7792 ;
  assign n7785 = ~\sa31_reg[5]/P0001  & n1160 ;
  assign n7794 = ~\sa31_reg[1]/P0001  & ~n6089 ;
  assign n7795 = ~n7785 & n7794 ;
  assign n7796 = ~n7793 & n7795 ;
  assign n7797 = \sa31_reg[4]/P0001  & n1269 ;
  assign n7798 = ~\sa31_reg[2]/P0001  & ~n7797 ;
  assign n7799 = n6788 & n7798 ;
  assign n7800 = n1276 & n5241 ;
  assign n7801 = \sa31_reg[2]/P0001  & ~n1153 ;
  assign n7802 = ~n5261 & n7801 ;
  assign n7803 = ~n7800 & n7802 ;
  assign n7804 = ~n7799 & ~n7803 ;
  assign n7805 = \sa31_reg[1]/P0001  & ~n5206 ;
  assign n7806 = ~n7804 & n7805 ;
  assign n7807 = ~n7796 & ~n7806 ;
  assign n7782 = ~n1182 & ~n1187 ;
  assign n7783 = ~\sa31_reg[3]/P0001  & n1244 ;
  assign n7784 = ~n7782 & n7783 ;
  assign n7851 = ~n7297 & ~n7784 ;
  assign n7852 = ~n7807 & n7851 ;
  assign n7853 = ~n7850 & n7852 ;
  assign n7854 = n6657 & ~n7853 ;
  assign n7855 = ~n6657 & n7853 ;
  assign n7856 = ~n7854 & ~n7855 ;
  assign n7857 = \u0_w_reg[2][11]/P0001  & ~n7313 ;
  assign n7858 = ~\u0_w_reg[2][11]/P0001  & n7313 ;
  assign n7859 = ~n7857 & ~n7858 ;
  assign n7860 = n7856 & n7859 ;
  assign n7861 = ~n7856 & ~n7859 ;
  assign n7862 = ~n7860 & ~n7861 ;
  assign n7864 = n7781 & n7862 ;
  assign n7863 = ~n7781 & ~n7862 ;
  assign n7865 = ~\ld_r_reg/P0001  & ~n7863 ;
  assign n7866 = ~n7864 & n7865 ;
  assign n7868 = ~\text_in_r_reg[43]/P0001  & \u0_w_reg[2][11]/P0001  ;
  assign n7867 = \text_in_r_reg[43]/P0001  & ~\u0_w_reg[2][11]/P0001  ;
  assign n7869 = \ld_r_reg/P0001  & ~n7867 ;
  assign n7870 = ~n7868 & n7869 ;
  assign n7871 = ~n7866 & ~n7870 ;
  assign n7872 = \u0_w_reg[2][26]/P0001  & ~n7853 ;
  assign n7873 = ~\u0_w_reg[2][26]/P0001  & n7853 ;
  assign n7874 = ~n7872 & ~n7873 ;
  assign n7875 = n7760 & n7874 ;
  assign n7876 = ~n7760 & ~n7874 ;
  assign n7877 = ~n7875 & ~n7876 ;
  assign n7879 = n6395 & ~n7877 ;
  assign n7878 = ~n6395 & n7877 ;
  assign n7880 = ~\ld_r_reg/P0001  & ~n7878 ;
  assign n7881 = ~n7879 & n7880 ;
  assign n7883 = \text_in_r_reg[58]/P0001  & \u0_w_reg[2][26]/P0001  ;
  assign n7882 = ~\text_in_r_reg[58]/P0001  & ~\u0_w_reg[2][26]/P0001  ;
  assign n7884 = \ld_r_reg/P0001  & ~n7882 ;
  assign n7885 = ~n7883 & n7884 ;
  assign n7886 = ~n7881 & ~n7885 ;
  assign n7887 = n5417 & ~n7580 ;
  assign n7888 = ~n5417 & n7580 ;
  assign n7889 = ~n7887 & ~n7888 ;
  assign n7890 = n7118 & n7889 ;
  assign n7891 = ~n7118 & ~n7889 ;
  assign n7892 = ~n7890 & ~n7891 ;
  assign n7893 = \u0_w_reg[2][3]/P0001  & ~n7206 ;
  assign n7894 = ~\u0_w_reg[2][3]/P0001  & n7206 ;
  assign n7895 = ~n7893 & ~n7894 ;
  assign n7896 = n7856 & n7895 ;
  assign n7897 = ~n7856 & ~n7895 ;
  assign n7898 = ~n7896 & ~n7897 ;
  assign n7900 = n7892 & n7898 ;
  assign n7899 = ~n7892 & ~n7898 ;
  assign n7901 = ~\ld_r_reg/P0001  & ~n7899 ;
  assign n7902 = ~n7900 & n7901 ;
  assign n7904 = ~\text_in_r_reg[35]/P0001  & \u0_w_reg[2][3]/P0001  ;
  assign n7903 = \text_in_r_reg[35]/P0001  & ~\u0_w_reg[2][3]/P0001  ;
  assign n7905 = \ld_r_reg/P0001  & ~n7903 ;
  assign n7906 = ~n7904 & n7905 ;
  assign n7907 = ~n7902 & ~n7906 ;
  assign n7908 = \u0_w_reg[2][31]/P0001  & ~n5516 ;
  assign n7909 = ~\u0_w_reg[2][31]/P0001  & n5516 ;
  assign n7910 = ~n7908 & ~n7909 ;
  assign n7911 = n5631 & ~n6657 ;
  assign n7912 = ~n5631 & n6657 ;
  assign n7913 = ~n7911 & ~n7912 ;
  assign n7914 = n5194 & n7913 ;
  assign n7915 = ~n5194 & ~n7913 ;
  assign n7916 = ~n7914 & ~n7915 ;
  assign n7918 = n7910 & ~n7916 ;
  assign n7917 = ~n7910 & n7916 ;
  assign n7919 = ~\ld_r_reg/P0001  & ~n7917 ;
  assign n7920 = ~n7918 & n7919 ;
  assign n7922 = ~\text_in_r_reg[63]/P0001  & \u0_w_reg[2][31]/P0001  ;
  assign n7921 = \text_in_r_reg[63]/P0001  & ~\u0_w_reg[2][31]/P0001  ;
  assign n7923 = \ld_r_reg/P0001  & ~n7921 ;
  assign n7924 = ~n7922 & n7923 ;
  assign n7925 = ~n7920 & ~n7924 ;
  assign n7926 = ~\u0_w_reg[2][24]/P0001  & ~n6568 ;
  assign n7927 = \u0_w_reg[2][24]/P0001  & n6568 ;
  assign n7928 = ~n7926 & ~n7927 ;
  assign n7929 = n6927 & ~n7408 ;
  assign n7930 = ~n6927 & n7408 ;
  assign n7931 = ~n7929 & ~n7930 ;
  assign n7932 = ~n5519 & n7931 ;
  assign n7933 = n5519 & ~n7931 ;
  assign n7934 = ~n7932 & ~n7933 ;
  assign n7936 = n7928 & n7934 ;
  assign n7935 = ~n7928 & ~n7934 ;
  assign n7937 = ~\ld_r_reg/P0001  & ~n7935 ;
  assign n7938 = ~n7936 & n7937 ;
  assign n7940 = \text_in_r_reg[56]/P0001  & \u0_w_reg[2][24]/P0001  ;
  assign n7939 = ~\text_in_r_reg[56]/P0001  & ~\u0_w_reg[2][24]/P0001  ;
  assign n7941 = \ld_r_reg/P0001  & ~n7939 ;
  assign n7942 = ~n7940 & n7941 ;
  assign n7943 = ~n7938 & ~n7942 ;
  assign n7944 = ~\u0_w_reg[2][16]/P0001  & ~n6568 ;
  assign n7945 = \u0_w_reg[2][16]/P0001  & n6568 ;
  assign n7946 = ~n7944 & ~n7945 ;
  assign n7947 = n5516 & ~n6472 ;
  assign n7948 = ~n5516 & n6472 ;
  assign n7949 = ~n7947 & ~n7948 ;
  assign n7950 = n6930 & n7949 ;
  assign n7951 = ~n6930 & ~n7949 ;
  assign n7952 = ~n7950 & ~n7951 ;
  assign n7954 = n7946 & ~n7952 ;
  assign n7953 = ~n7946 & n7952 ;
  assign n7955 = ~\ld_r_reg/P0001  & ~n7953 ;
  assign n7956 = ~n7954 & n7955 ;
  assign n7958 = \text_in_r_reg[48]/P0001  & \u0_w_reg[2][16]/P0001  ;
  assign n7957 = ~\text_in_r_reg[48]/P0001  & ~\u0_w_reg[2][16]/P0001  ;
  assign n7959 = \ld_r_reg/P0001  & ~n7957 ;
  assign n7960 = ~n7958 & n7959 ;
  assign n7961 = ~n7956 & ~n7960 ;
  assign n7962 = ~n7580 & ~n7673 ;
  assign n7963 = n7580 & n7673 ;
  assign n7964 = ~n7962 & ~n7963 ;
  assign n7965 = \u0_w_reg[2][18]/P0001  & ~n7853 ;
  assign n7966 = ~\u0_w_reg[2][18]/P0001  & n7853 ;
  assign n7967 = ~n7965 & ~n7966 ;
  assign n7968 = n7655 & n7967 ;
  assign n7969 = ~n7655 & ~n7967 ;
  assign n7970 = ~n7968 & ~n7969 ;
  assign n7972 = n7964 & n7970 ;
  assign n7971 = ~n7964 & ~n7970 ;
  assign n7973 = ~\ld_r_reg/P0001  & ~n7971 ;
  assign n7974 = ~n7972 & n7973 ;
  assign n7976 = ~\text_in_r_reg[50]/P0001  & \u0_w_reg[2][18]/P0001  ;
  assign n7975 = \text_in_r_reg[50]/P0001  & ~\u0_w_reg[2][18]/P0001  ;
  assign n7977 = \ld_r_reg/P0001  & ~n7975 ;
  assign n7978 = ~n7976 & n7977 ;
  assign n7979 = ~n7974 & ~n7978 ;
  assign n7980 = ~n853 & ~n5417 ;
  assign n7981 = n853 & n5417 ;
  assign n7982 = ~n7980 & ~n7981 ;
  assign n7983 = ~\u0_w_reg[2][23]/P0001  & ~n7913 ;
  assign n7984 = \u0_w_reg[2][23]/P0001  & n7913 ;
  assign n7985 = ~n7983 & ~n7984 ;
  assign n7987 = n7982 & n7985 ;
  assign n7986 = ~n7982 & ~n7985 ;
  assign n7988 = ~\ld_r_reg/P0001  & ~n7986 ;
  assign n7989 = ~n7987 & n7988 ;
  assign n7991 = ~\text_in_r_reg[55]/P0001  & \u0_w_reg[2][23]/P0001  ;
  assign n7990 = \text_in_r_reg[55]/P0001  & ~\u0_w_reg[2][23]/P0001  ;
  assign n7992 = \ld_r_reg/P0001  & ~n7990 ;
  assign n7993 = ~n7991 & n7992 ;
  assign n7994 = ~n7989 & ~n7993 ;
  assign n7995 = ~\u0_w_reg[2][8]/P0001  & ~n6568 ;
  assign n7996 = \u0_w_reg[2][8]/P0001  & n6568 ;
  assign n7997 = ~n7995 & ~n7996 ;
  assign n7998 = n6472 & ~n7408 ;
  assign n7999 = ~n6472 & n7408 ;
  assign n8000 = ~n7998 & ~n7999 ;
  assign n8001 = n7913 & n8000 ;
  assign n8002 = ~n7913 & ~n8000 ;
  assign n8003 = ~n8001 & ~n8002 ;
  assign n8005 = n7997 & n8003 ;
  assign n8004 = ~n7997 & ~n8003 ;
  assign n8006 = ~\ld_r_reg/P0001  & ~n8004 ;
  assign n8007 = ~n8005 & n8006 ;
  assign n8009 = ~\text_in_r_reg[40]/P0001  & \u0_w_reg[2][8]/P0001  ;
  assign n8008 = \text_in_r_reg[40]/P0001  & ~\u0_w_reg[2][8]/P0001  ;
  assign n8010 = \ld_r_reg/P0001  & ~n8008 ;
  assign n8011 = ~n8009 & n8010 ;
  assign n8012 = ~n8007 & ~n8011 ;
  assign n8013 = ~n6743 & ~n7583 ;
  assign n8014 = n6743 & n7583 ;
  assign n8015 = ~n8013 & ~n8014 ;
  assign n8016 = \u0_w_reg[2][10]/P0001  & ~n7853 ;
  assign n8017 = ~\u0_w_reg[2][10]/P0001  & n7853 ;
  assign n8018 = ~n8016 & ~n8017 ;
  assign n8019 = n6842 & n8018 ;
  assign n8020 = ~n6842 & ~n8018 ;
  assign n8021 = ~n8019 & ~n8020 ;
  assign n8023 = n8015 & n8021 ;
  assign n8022 = ~n8015 & ~n8021 ;
  assign n8024 = ~\ld_r_reg/P0001  & ~n8022 ;
  assign n8025 = ~n8023 & n8024 ;
  assign n8027 = ~\text_in_r_reg[42]/P0001  & \u0_w_reg[2][10]/P0001  ;
  assign n8026 = \text_in_r_reg[42]/P0001  & ~\u0_w_reg[2][10]/P0001  ;
  assign n8028 = \ld_r_reg/P0001  & ~n8026 ;
  assign n8029 = ~n8027 & n8028 ;
  assign n8030 = ~n8025 & ~n8029 ;
  assign n8031 = ~\u0_w_reg[2][5]/P0001  & ~n5307 ;
  assign n8032 = \u0_w_reg[2][5]/P0001  & n5307 ;
  assign n8033 = ~n8031 & ~n8032 ;
  assign n8034 = ~\u0_w_reg[2][6]/P0001  & ~n1300 ;
  assign n8035 = \u0_w_reg[2][6]/P0001  & n1300 ;
  assign n8036 = ~n8034 & ~n8035 ;
  assign n8037 = ~\u0_w_reg[2][4]/P0001  & ~n6180 ;
  assign n8038 = \u0_w_reg[2][4]/P0001  & n6180 ;
  assign n8039 = ~n8037 & ~n8038 ;
  assign n8040 = ~\u0_w_reg[2][0]/P0001  & ~n6568 ;
  assign n8041 = \u0_w_reg[2][0]/P0001  & n6568 ;
  assign n8042 = ~n8040 & ~n8041 ;
  assign n8043 = ~\u0_w_reg[2][3]/P0001  & ~n7313 ;
  assign n8044 = \u0_w_reg[2][3]/P0001  & n7313 ;
  assign n8045 = ~n8043 & ~n8044 ;
  assign n8046 = ~\u0_w_reg[2][1]/P0001  & ~n6842 ;
  assign n8047 = \u0_w_reg[2][1]/P0001  & n6842 ;
  assign n8048 = ~n8046 & ~n8047 ;
  assign n8049 = ~\u0_w_reg[2][2]/P0001  & ~n7853 ;
  assign n8050 = \u0_w_reg[2][2]/P0001  & n7853 ;
  assign n8051 = ~n8049 & ~n8050 ;
  assign n8052 = ~\u0_w_reg[2][7]/P0001  & ~n6657 ;
  assign n8053 = \u0_w_reg[2][7]/P0001  & n6657 ;
  assign n8054 = ~n8052 & ~n8053 ;
  assign n8060 = \sa12_reg[6]/NET0131  & ~\sa12_reg[7]/NET0131  ;
  assign n8146 = ~\sa12_reg[4]/P0001  & n8060 ;
  assign n8080 = \sa12_reg[4]/P0001  & \sa12_reg[7]/NET0131  ;
  assign n8082 = ~\sa12_reg[5]/P0001  & ~\sa12_reg[6]/NET0131  ;
  assign n8147 = n8080 & n8082 ;
  assign n8148 = ~n8146 & ~n8147 ;
  assign n8149 = ~\sa12_reg[2]/P0001  & ~n8148 ;
  assign n8074 = \sa12_reg[5]/P0001  & ~\sa12_reg[7]/NET0131  ;
  assign n8078 = \sa12_reg[3]/P0001  & ~\sa12_reg[4]/P0001  ;
  assign n8129 = ~\sa12_reg[6]/NET0131  & n8078 ;
  assign n8150 = n8074 & n8129 ;
  assign n8094 = ~\sa12_reg[3]/P0001  & \sa12_reg[4]/P0001  ;
  assign n8142 = ~\sa12_reg[7]/NET0131  & n8082 ;
  assign n8143 = n8094 & n8142 ;
  assign n8126 = ~\sa12_reg[6]/NET0131  & \sa12_reg[7]/NET0131  ;
  assign n8144 = \sa12_reg[2]/P0001  & ~\sa12_reg[4]/P0001  ;
  assign n8145 = n8126 & n8144 ;
  assign n8151 = \sa12_reg[1]/P0001  & ~n8145 ;
  assign n8152 = ~n8143 & n8151 ;
  assign n8153 = ~n8150 & n8152 ;
  assign n8154 = ~n8149 & n8153 ;
  assign n8161 = \sa12_reg[5]/P0001  & \sa12_reg[7]/NET0131  ;
  assign n8165 = \sa12_reg[4]/P0001  & n8161 ;
  assign n8166 = ~\sa12_reg[6]/NET0131  & n8165 ;
  assign n8167 = \sa12_reg[2]/P0001  & n8166 ;
  assign n8155 = ~\sa12_reg[2]/P0001  & \sa12_reg[3]/P0001  ;
  assign n8055 = ~\sa12_reg[6]/NET0131  & ~\sa12_reg[7]/NET0131  ;
  assign n8156 = \sa12_reg[4]/P0001  & n8055 ;
  assign n8157 = n8155 & n8156 ;
  assign n8158 = ~\sa12_reg[1]/P0001  & ~n8157 ;
  assign n8075 = \sa12_reg[3]/P0001  & \sa12_reg[6]/NET0131  ;
  assign n8159 = \sa12_reg[7]/NET0131  & n8075 ;
  assign n8160 = ~\sa12_reg[4]/P0001  & n8159 ;
  assign n8162 = ~\sa12_reg[2]/P0001  & ~\sa12_reg[4]/P0001  ;
  assign n8163 = ~\sa12_reg[3]/P0001  & ~n8162 ;
  assign n8164 = n8161 & ~n8163 ;
  assign n8168 = ~n8160 & ~n8164 ;
  assign n8169 = n8158 & n8168 ;
  assign n8170 = ~n8167 & n8169 ;
  assign n8171 = ~n8154 & ~n8170 ;
  assign n8065 = \sa12_reg[5]/P0001  & \sa12_reg[6]/NET0131  ;
  assign n8130 = \sa12_reg[7]/NET0131  & n8065 ;
  assign n8131 = ~n8094 & ~n8130 ;
  assign n8132 = ~n8080 & ~n8131 ;
  assign n8110 = \sa12_reg[3]/P0001  & ~\sa12_reg[5]/P0001  ;
  assign n8127 = n8110 & n8126 ;
  assign n8128 = \sa12_reg[2]/P0001  & ~n8127 ;
  assign n8133 = n8128 & ~n8129 ;
  assign n8134 = ~n8132 & n8133 ;
  assign n8135 = ~\sa12_reg[5]/P0001  & \sa12_reg[7]/NET0131  ;
  assign n8136 = n8075 & n8135 ;
  assign n8137 = ~\sa12_reg[2]/P0001  & ~n8136 ;
  assign n8104 = ~\sa12_reg[3]/P0001  & ~\sa12_reg[4]/P0001  ;
  assign n8117 = n8082 & n8104 ;
  assign n8118 = ~\sa12_reg[7]/NET0131  & n8117 ;
  assign n8138 = n8060 & n8078 ;
  assign n8139 = ~n8118 & ~n8138 ;
  assign n8140 = n8137 & n8139 ;
  assign n8141 = ~n8134 & ~n8140 ;
  assign n8172 = \sa12_reg[0]/P0001  & ~n8141 ;
  assign n8173 = ~n8171 & n8172 ;
  assign n8111 = ~\sa12_reg[4]/P0001  & \sa12_reg[7]/NET0131  ;
  assign n8184 = n8082 & n8111 ;
  assign n8185 = \sa12_reg[5]/P0001  & n8126 ;
  assign n8186 = ~n8078 & n8185 ;
  assign n8187 = ~n8184 & ~n8186 ;
  assign n8188 = ~\sa12_reg[2]/P0001  & ~n8187 ;
  assign n8174 = \sa12_reg[5]/P0001  & n8060 ;
  assign n8189 = \sa12_reg[2]/P0001  & n8174 ;
  assign n8059 = \sa12_reg[2]/P0001  & ~\sa12_reg[3]/P0001  ;
  assign n8182 = \sa12_reg[4]/P0001  & n8135 ;
  assign n8183 = n8059 & n8182 ;
  assign n8180 = \sa12_reg[3]/P0001  & \sa12_reg[4]/P0001  ;
  assign n8181 = n8060 & n8180 ;
  assign n8190 = \sa12_reg[1]/P0001  & ~n8181 ;
  assign n8191 = ~n8183 & n8190 ;
  assign n8192 = ~n8189 & n8191 ;
  assign n8193 = ~n8188 & n8192 ;
  assign n8195 = ~\sa12_reg[7]/NET0131  & n8129 ;
  assign n8194 = \sa12_reg[2]/P0001  & n8142 ;
  assign n8066 = \sa12_reg[2]/P0001  & \sa12_reg[4]/P0001  ;
  assign n8067 = n8065 & n8066 ;
  assign n8196 = ~\sa12_reg[1]/P0001  & ~n8067 ;
  assign n8197 = ~n8194 & n8196 ;
  assign n8198 = ~n8195 & n8197 ;
  assign n8199 = ~n8193 & ~n8198 ;
  assign n8175 = ~\sa12_reg[3]/P0001  & n8174 ;
  assign n8176 = ~\sa12_reg[1]/P0001  & n8175 ;
  assign n8093 = ~\sa12_reg[5]/P0001  & \sa12_reg[6]/NET0131  ;
  assign n8095 = n8093 & n8094 ;
  assign n8177 = \sa12_reg[7]/NET0131  & n8095 ;
  assign n8178 = ~n8176 & ~n8177 ;
  assign n8179 = ~\sa12_reg[2]/P0001  & ~n8178 ;
  assign n8069 = ~\sa12_reg[5]/P0001  & ~\sa12_reg[7]/NET0131  ;
  assign n8200 = n8069 & n8180 ;
  assign n8201 = ~\sa12_reg[6]/NET0131  & n8200 ;
  assign n8202 = ~\sa12_reg[4]/P0001  & n8093 ;
  assign n8203 = ~\sa12_reg[3]/P0001  & n8202 ;
  assign n8204 = ~n8201 & ~n8203 ;
  assign n8205 = \sa12_reg[2]/P0001  & ~n8204 ;
  assign n8056 = \sa12_reg[5]/P0001  & n8055 ;
  assign n8105 = n8056 & n8104 ;
  assign n8206 = ~\sa12_reg[0]/P0001  & ~n8105 ;
  assign n8207 = ~n8205 & n8206 ;
  assign n8208 = ~n8179 & n8207 ;
  assign n8209 = ~n8199 & n8208 ;
  assign n8210 = ~n8173 & ~n8209 ;
  assign n8077 = \sa12_reg[5]/P0001  & ~\sa12_reg[6]/NET0131  ;
  assign n8079 = n8077 & n8078 ;
  assign n8076 = n8074 & n8075 ;
  assign n8088 = \sa12_reg[2]/P0001  & ~n8076 ;
  assign n8089 = ~n8079 & n8088 ;
  assign n8087 = ~\sa12_reg[3]/P0001  & n8056 ;
  assign n8081 = \sa12_reg[3]/P0001  & n8080 ;
  assign n8083 = n8081 & n8082 ;
  assign n8084 = ~\sa12_reg[3]/P0001  & \sa12_reg[7]/NET0131  ;
  assign n8085 = ~\sa12_reg[4]/P0001  & n8084 ;
  assign n8086 = n8082 & n8085 ;
  assign n8090 = ~n8083 & ~n8086 ;
  assign n8091 = ~n8087 & n8090 ;
  assign n8092 = n8089 & n8091 ;
  assign n8097 = n8065 & n8078 ;
  assign n8098 = \sa12_reg[7]/NET0131  & n8097 ;
  assign n8096 = n8084 & n8093 ;
  assign n8099 = ~\sa12_reg[2]/P0001  & ~n8095 ;
  assign n8100 = ~n8096 & n8099 ;
  assign n8101 = ~n8098 & n8100 ;
  assign n8102 = ~n8092 & ~n8101 ;
  assign n8103 = \sa12_reg[4]/P0001  & n8076 ;
  assign n8106 = ~\sa12_reg[1]/P0001  & ~n8103 ;
  assign n8107 = ~n8105 & n8106 ;
  assign n8108 = ~n8102 & n8107 ;
  assign n8114 = n8065 & n8084 ;
  assign n8115 = ~\sa12_reg[4]/P0001  & n8114 ;
  assign n8116 = ~n8055 & n8110 ;
  assign n8119 = ~n8115 & ~n8116 ;
  assign n8120 = ~n8118 & n8119 ;
  assign n8121 = ~\sa12_reg[2]/P0001  & ~n8120 ;
  assign n8112 = n8110 & n8111 ;
  assign n8113 = ~\sa12_reg[6]/NET0131  & n8112 ;
  assign n8109 = n8081 & n8093 ;
  assign n8122 = \sa12_reg[1]/P0001  & ~n8109 ;
  assign n8123 = ~n8113 & n8122 ;
  assign n8124 = ~n8121 & n8123 ;
  assign n8125 = ~n8108 & ~n8124 ;
  assign n8057 = \sa12_reg[2]/P0001  & \sa12_reg[3]/P0001  ;
  assign n8058 = n8056 & n8057 ;
  assign n8061 = \sa12_reg[4]/P0001  & n8060 ;
  assign n8062 = n8059 & n8061 ;
  assign n8063 = ~n8058 & ~n8062 ;
  assign n8064 = \sa12_reg[1]/P0001  & ~n8063 ;
  assign n8068 = ~\sa12_reg[4]/P0001  & \sa12_reg[6]/NET0131  ;
  assign n8070 = n8068 & n8069 ;
  assign n8071 = ~\sa12_reg[2]/P0001  & n8070 ;
  assign n8072 = ~n8067 & ~n8071 ;
  assign n8073 = \sa12_reg[3]/P0001  & ~n8072 ;
  assign n8211 = ~n8064 & ~n8073 ;
  assign n8212 = ~n8125 & n8211 ;
  assign n8213 = ~n8210 & n8212 ;
  assign n8218 = \sa01_reg[3]/P0001  & ~\sa01_reg[4]/P0001  ;
  assign n8221 = ~\sa01_reg[6]/NET0131  & \sa01_reg[7]/NET0131  ;
  assign n8279 = \sa01_reg[5]/P0001  & n8221 ;
  assign n8280 = ~n8218 & n8279 ;
  assign n8281 = ~\sa01_reg[4]/P0001  & \sa01_reg[7]/NET0131  ;
  assign n8282 = ~\sa01_reg[5]/P0001  & n8281 ;
  assign n8283 = ~\sa01_reg[6]/NET0131  & n8282 ;
  assign n8284 = ~n8280 & ~n8283 ;
  assign n8285 = ~\sa01_reg[2]/P0001  & ~n8284 ;
  assign n8254 = ~\sa01_reg[5]/P0001  & \sa01_reg[7]/NET0131  ;
  assign n8214 = ~\sa01_reg[3]/P0001  & \sa01_reg[4]/P0001  ;
  assign n8287 = \sa01_reg[2]/P0001  & n8214 ;
  assign n8288 = n8254 & n8287 ;
  assign n8276 = \sa01_reg[6]/NET0131  & ~\sa01_reg[7]/NET0131  ;
  assign n8277 = \sa01_reg[5]/P0001  & n8276 ;
  assign n8278 = \sa01_reg[2]/P0001  & n8277 ;
  assign n8238 = \sa01_reg[3]/P0001  & \sa01_reg[4]/P0001  ;
  assign n8286 = n8238 & n8276 ;
  assign n8289 = \sa01_reg[1]/P0001  & ~n8286 ;
  assign n8290 = ~n8278 & n8289 ;
  assign n8291 = ~n8288 & n8290 ;
  assign n8292 = ~n8285 & n8291 ;
  assign n8215 = ~\sa01_reg[6]/NET0131  & ~\sa01_reg[7]/NET0131  ;
  assign n8216 = ~\sa01_reg[5]/P0001  & n8215 ;
  assign n8257 = \sa01_reg[5]/P0001  & \sa01_reg[6]/NET0131  ;
  assign n8295 = \sa01_reg[4]/P0001  & n8257 ;
  assign n8296 = ~n8216 & ~n8295 ;
  assign n8297 = \sa01_reg[2]/P0001  & ~n8296 ;
  assign n8293 = ~\sa01_reg[3]/P0001  & n8277 ;
  assign n8294 = ~\sa01_reg[2]/P0001  & n8293 ;
  assign n8298 = n8215 & n8218 ;
  assign n8299 = ~\sa01_reg[1]/P0001  & ~n8298 ;
  assign n8300 = ~n8294 & n8299 ;
  assign n8301 = ~n8297 & n8300 ;
  assign n8302 = ~n8292 & ~n8301 ;
  assign n8303 = \sa01_reg[2]/P0001  & ~\sa01_reg[5]/P0001  ;
  assign n8267 = ~\sa01_reg[3]/P0001  & ~\sa01_reg[4]/P0001  ;
  assign n8304 = \sa01_reg[6]/NET0131  & n8267 ;
  assign n8305 = n8215 & n8238 ;
  assign n8306 = ~n8304 & ~n8305 ;
  assign n8307 = n8303 & ~n8306 ;
  assign n8308 = ~\sa01_reg[4]/P0001  & \sa01_reg[5]/P0001  ;
  assign n8309 = n8215 & n8308 ;
  assign n8310 = ~\sa01_reg[5]/P0001  & \sa01_reg[6]/NET0131  ;
  assign n8224 = \sa01_reg[4]/P0001  & \sa01_reg[7]/NET0131  ;
  assign n8311 = ~\sa01_reg[2]/P0001  & n8224 ;
  assign n8312 = n8310 & n8311 ;
  assign n8313 = ~n8309 & ~n8312 ;
  assign n8314 = ~\sa01_reg[3]/P0001  & ~n8313 ;
  assign n8315 = ~n8307 & ~n8314 ;
  assign n8316 = ~n8302 & n8315 ;
  assign n8317 = ~\sa01_reg[0]/P0001  & ~n8316 ;
  assign n8227 = ~\sa01_reg[5]/P0001  & ~\sa01_reg[6]/NET0131  ;
  assign n8228 = \sa01_reg[7]/NET0131  & ~n8227 ;
  assign n8225 = ~\sa01_reg[4]/P0001  & \sa01_reg[6]/NET0131  ;
  assign n8226 = ~n8224 & ~n8225 ;
  assign n8229 = ~\sa01_reg[2]/P0001  & ~n8226 ;
  assign n8230 = ~n8228 & n8229 ;
  assign n8219 = \sa01_reg[5]/P0001  & n8215 ;
  assign n8220 = n8218 & n8219 ;
  assign n8217 = n8214 & n8216 ;
  assign n8222 = \sa01_reg[2]/P0001  & ~\sa01_reg[4]/P0001  ;
  assign n8223 = n8221 & n8222 ;
  assign n8231 = \sa01_reg[1]/P0001  & ~n8223 ;
  assign n8232 = ~n8217 & n8231 ;
  assign n8233 = ~n8220 & n8232 ;
  assign n8234 = ~n8230 & n8233 ;
  assign n8235 = \sa01_reg[6]/NET0131  & \sa01_reg[7]/NET0131  ;
  assign n8236 = n8218 & n8235 ;
  assign n8237 = ~\sa01_reg[1]/P0001  & ~n8236 ;
  assign n8239 = ~\sa01_reg[6]/NET0131  & n8238 ;
  assign n8240 = ~\sa01_reg[2]/P0001  & ~\sa01_reg[7]/NET0131  ;
  assign n8241 = n8239 & n8240 ;
  assign n8249 = n8237 & ~n8241 ;
  assign n8242 = \sa01_reg[5]/P0001  & ~\sa01_reg[6]/NET0131  ;
  assign n8243 = n8224 & n8242 ;
  assign n8244 = \sa01_reg[2]/P0001  & n8243 ;
  assign n8245 = \sa01_reg[5]/P0001  & \sa01_reg[7]/NET0131  ;
  assign n8246 = ~\sa01_reg[2]/P0001  & ~\sa01_reg[4]/P0001  ;
  assign n8247 = ~\sa01_reg[3]/P0001  & ~n8246 ;
  assign n8248 = n8245 & ~n8247 ;
  assign n8250 = ~n8244 & ~n8248 ;
  assign n8251 = n8249 & n8250 ;
  assign n8252 = ~n8234 & ~n8251 ;
  assign n8258 = \sa01_reg[7]/NET0131  & n8257 ;
  assign n8253 = \sa01_reg[3]/P0001  & ~\sa01_reg[6]/NET0131  ;
  assign n8256 = ~\sa01_reg[4]/P0001  & n8253 ;
  assign n8259 = ~n8214 & ~n8256 ;
  assign n8260 = ~n8258 & n8259 ;
  assign n8261 = ~n8224 & ~n8260 ;
  assign n8255 = n8253 & n8254 ;
  assign n8262 = \sa01_reg[2]/P0001  & ~n8255 ;
  assign n8263 = ~n8261 & n8262 ;
  assign n8268 = n8216 & n8267 ;
  assign n8264 = \sa01_reg[3]/P0001  & \sa01_reg[6]/NET0131  ;
  assign n8269 = n8254 & n8264 ;
  assign n8265 = ~\sa01_reg[4]/P0001  & ~\sa01_reg[7]/NET0131  ;
  assign n8266 = n8264 & n8265 ;
  assign n8270 = ~\sa01_reg[2]/P0001  & ~n8266 ;
  assign n8271 = ~n8269 & n8270 ;
  assign n8272 = ~n8268 & n8271 ;
  assign n8273 = ~n8263 & ~n8272 ;
  assign n8274 = ~n8252 & ~n8273 ;
  assign n8275 = \sa01_reg[0]/P0001  & ~n8274 ;
  assign n8320 = \sa01_reg[7]/NET0131  & n8267 ;
  assign n8321 = \sa01_reg[5]/P0001  & n8320 ;
  assign n8322 = \sa01_reg[6]/NET0131  & n8321 ;
  assign n8318 = \sa01_reg[3]/P0001  & ~\sa01_reg[5]/P0001  ;
  assign n8319 = ~n8215 & n8318 ;
  assign n8323 = ~n8268 & ~n8319 ;
  assign n8324 = ~n8322 & n8323 ;
  assign n8325 = ~\sa01_reg[2]/P0001  & ~n8324 ;
  assign n8326 = ~\sa01_reg[3]/P0001  & n8276 ;
  assign n8327 = \sa01_reg[2]/P0001  & \sa01_reg[4]/P0001  ;
  assign n8328 = n8326 & n8327 ;
  assign n8334 = \sa01_reg[1]/P0001  & ~n8328 ;
  assign n8333 = n8254 & n8256 ;
  assign n8329 = \sa01_reg[2]/P0001  & \sa01_reg[3]/P0001  ;
  assign n8330 = n8219 & n8329 ;
  assign n8331 = ~\sa01_reg[5]/P0001  & n8224 ;
  assign n8332 = n8264 & n8331 ;
  assign n8335 = ~n8330 & ~n8332 ;
  assign n8336 = ~n8333 & n8335 ;
  assign n8337 = n8334 & n8336 ;
  assign n8338 = ~n8325 & n8337 ;
  assign n8342 = \sa01_reg[5]/P0001  & ~\sa01_reg[7]/NET0131  ;
  assign n8343 = n8264 & n8342 ;
  assign n8341 = n8253 & n8308 ;
  assign n8347 = \sa01_reg[2]/P0001  & ~n8341 ;
  assign n8348 = ~n8343 & n8347 ;
  assign n8339 = ~\sa01_reg[3]/P0001  & n8215 ;
  assign n8340 = \sa01_reg[5]/P0001  & n8339 ;
  assign n8344 = ~\sa01_reg[5]/P0001  & n8221 ;
  assign n8345 = ~n8214 & ~n8218 ;
  assign n8346 = n8344 & n8345 ;
  assign n8349 = ~n8340 & ~n8346 ;
  assign n8350 = n8348 & n8349 ;
  assign n8354 = \sa01_reg[3]/P0001  & n8308 ;
  assign n8355 = n8235 & n8354 ;
  assign n8351 = ~\sa01_reg[3]/P0001  & ~\sa01_reg[5]/P0001  ;
  assign n8352 = n8235 & n8351 ;
  assign n8353 = ~\sa01_reg[2]/P0001  & ~n8352 ;
  assign n8356 = n8214 & n8310 ;
  assign n8357 = n8353 & ~n8356 ;
  assign n8358 = ~n8355 & n8357 ;
  assign n8359 = ~n8350 & ~n8358 ;
  assign n8362 = n8215 & n8267 ;
  assign n8363 = \sa01_reg[5]/P0001  & n8362 ;
  assign n8360 = n8238 & n8342 ;
  assign n8361 = \sa01_reg[6]/NET0131  & n8360 ;
  assign n8364 = ~\sa01_reg[1]/P0001  & ~n8361 ;
  assign n8365 = ~n8363 & n8364 ;
  assign n8366 = ~n8359 & n8365 ;
  assign n8367 = ~n8338 & ~n8366 ;
  assign n8371 = \sa01_reg[2]/P0001  & ~n8295 ;
  assign n8368 = ~\sa01_reg[5]/P0001  & ~\sa01_reg[7]/NET0131  ;
  assign n8369 = n8225 & n8368 ;
  assign n8370 = ~\sa01_reg[2]/P0001  & ~n8369 ;
  assign n8372 = \sa01_reg[3]/P0001  & ~n8370 ;
  assign n8373 = ~n8371 & n8372 ;
  assign n8374 = ~n8367 & ~n8373 ;
  assign n8375 = ~n8275 & n8374 ;
  assign n8376 = ~n8317 & n8375 ;
  assign n8377 = n8213 & ~n8376 ;
  assign n8378 = ~n8213 & n8376 ;
  assign n8379 = ~n8377 & ~n8378 ;
  assign n8382 = ~\sa12_reg[3]/P0001  & n8146 ;
  assign n8380 = n8077 & n8094 ;
  assign n8381 = \sa12_reg[3]/P0001  & n8126 ;
  assign n8383 = ~n8380 & ~n8381 ;
  assign n8384 = ~n8382 & n8383 ;
  assign n8385 = ~\sa12_reg[2]/P0001  & ~n8384 ;
  assign n8389 = \sa12_reg[3]/P0001  & n8161 ;
  assign n8390 = \sa12_reg[4]/P0001  & \sa12_reg[6]/NET0131  ;
  assign n8391 = n8074 & n8390 ;
  assign n8392 = ~n8389 & ~n8391 ;
  assign n8393 = \sa12_reg[2]/P0001  & ~n8392 ;
  assign n8394 = n8065 & n8104 ;
  assign n8395 = ~\sa12_reg[7]/NET0131  & n8394 ;
  assign n8386 = n8161 & n8180 ;
  assign n8396 = ~n8096 & ~n8386 ;
  assign n8387 = n8055 & n8110 ;
  assign n8388 = n8077 & n8111 ;
  assign n8397 = ~n8387 & ~n8388 ;
  assign n8398 = n8396 & n8397 ;
  assign n8399 = ~n8395 & n8398 ;
  assign n8400 = ~n8393 & n8399 ;
  assign n8401 = ~n8385 & n8400 ;
  assign n8402 = \sa12_reg[1]/P0001  & ~n8401 ;
  assign n8412 = ~\sa12_reg[5]/P0001  & n8060 ;
  assign n8413 = ~\sa12_reg[3]/P0001  & n8412 ;
  assign n8414 = ~\sa12_reg[4]/P0001  & n8069 ;
  assign n8415 = ~n8413 & ~n8414 ;
  assign n8416 = ~n8104 & ~n8415 ;
  assign n8417 = ~\sa12_reg[4]/P0001  & n8055 ;
  assign n8418 = ~n8386 & ~n8417 ;
  assign n8419 = ~n8416 & n8418 ;
  assign n8420 = \sa12_reg[2]/P0001  & ~n8419 ;
  assign n8403 = \sa12_reg[2]/P0001  & n8129 ;
  assign n8404 = ~\sa12_reg[6]/NET0131  & n8084 ;
  assign n8405 = \sa12_reg[4]/P0001  & n8404 ;
  assign n8406 = ~n8403 & ~n8405 ;
  assign n8407 = ~\sa12_reg[5]/P0001  & ~n8406 ;
  assign n8408 = ~\sa12_reg[3]/P0001  & n8194 ;
  assign n8409 = ~n8115 & ~n8408 ;
  assign n8410 = ~n8407 & n8409 ;
  assign n8411 = ~\sa12_reg[1]/P0001  & ~n8410 ;
  assign n8422 = n8068 & n8135 ;
  assign n8423 = ~n8200 & ~n8422 ;
  assign n8424 = ~\sa12_reg[2]/P0001  & ~n8423 ;
  assign n8421 = ~\sa12_reg[2]/P0001  & n8166 ;
  assign n8425 = ~\sa12_reg[4]/P0001  & n8142 ;
  assign n8426 = ~n8421 & ~n8425 ;
  assign n8427 = ~n8424 & n8426 ;
  assign n8428 = ~n8411 & n8427 ;
  assign n8429 = ~n8420 & n8428 ;
  assign n8430 = ~n8402 & n8429 ;
  assign n8431 = ~\sa12_reg[0]/P0001  & ~n8430 ;
  assign n8434 = n8055 & n8180 ;
  assign n8435 = \sa12_reg[2]/P0001  & ~n8202 ;
  assign n8436 = ~n8434 & n8435 ;
  assign n8437 = ~\sa12_reg[2]/P0001  & ~n8127 ;
  assign n8438 = ~n8174 & n8437 ;
  assign n8439 = ~n8436 & ~n8438 ;
  assign n8432 = n8065 & n8080 ;
  assign n8433 = ~\sa12_reg[3]/P0001  & n8432 ;
  assign n8440 = ~n8076 & ~n8433 ;
  assign n8441 = ~n8439 & n8440 ;
  assign n8442 = ~\sa12_reg[1]/P0001  & ~n8441 ;
  assign n8459 = ~\sa12_reg[6]/NET0131  & n8180 ;
  assign n8460 = n8074 & n8459 ;
  assign n8461 = \sa12_reg[7]/NET0131  & n8380 ;
  assign n8462 = ~n8460 & ~n8461 ;
  assign n8463 = n8078 & n8126 ;
  assign n8464 = ~n8143 & ~n8463 ;
  assign n8465 = n8462 & n8464 ;
  assign n8466 = \sa12_reg[1]/P0001  & ~n8465 ;
  assign n8443 = ~\sa12_reg[4]/P0001  & n8074 ;
  assign n8444 = ~n8076 & ~n8138 ;
  assign n8445 = ~n8443 & n8444 ;
  assign n8446 = ~\sa12_reg[2]/P0001  & ~n8445 ;
  assign n8454 = \sa12_reg[5]/P0001  & ~n8078 ;
  assign n8455 = \sa12_reg[1]/P0001  & ~\sa12_reg[2]/P0001  ;
  assign n8456 = ~n8080 & n8455 ;
  assign n8457 = ~n8202 & n8456 ;
  assign n8458 = ~n8454 & n8457 ;
  assign n8447 = \sa12_reg[2]/P0001  & n8104 ;
  assign n8448 = n8412 & n8447 ;
  assign n8449 = ~\sa12_reg[7]/NET0131  & n8097 ;
  assign n8467 = ~n8448 & ~n8449 ;
  assign n8450 = \sa12_reg[2]/P0001  & n8094 ;
  assign n8451 = n8130 & n8450 ;
  assign n8452 = n8080 & n8093 ;
  assign n8453 = ~\sa12_reg[2]/P0001  & n8452 ;
  assign n8468 = ~n8451 & ~n8453 ;
  assign n8469 = n8467 & n8468 ;
  assign n8470 = ~n8458 & n8469 ;
  assign n8471 = ~n8446 & n8470 ;
  assign n8472 = ~n8466 & n8471 ;
  assign n8473 = ~n8442 & n8472 ;
  assign n8474 = \sa12_reg[0]/P0001  & ~n8473 ;
  assign n8475 = ~n8085 & ~n8181 ;
  assign n8476 = \sa12_reg[5]/P0001  & ~n8475 ;
  assign n8477 = ~n8452 & ~n8476 ;
  assign n8478 = ~\sa12_reg[2]/P0001  & ~n8477 ;
  assign n8481 = ~\sa12_reg[5]/P0001  & n8126 ;
  assign n8482 = ~n8412 & ~n8481 ;
  assign n8483 = ~n8130 & n8482 ;
  assign n8484 = n8450 & ~n8483 ;
  assign n8479 = \sa12_reg[2]/P0001  & n8180 ;
  assign n8480 = n8077 & n8479 ;
  assign n8485 = n8055 & n8104 ;
  assign n8486 = ~n8480 & ~n8485 ;
  assign n8487 = ~n8484 & n8486 ;
  assign n8488 = ~n8478 & n8487 ;
  assign n8489 = ~\sa12_reg[1]/P0001  & ~n8488 ;
  assign n8494 = n8074 & n8094 ;
  assign n8495 = \sa12_reg[6]/NET0131  & n8494 ;
  assign n8496 = \sa12_reg[2]/P0001  & n8495 ;
  assign n8497 = ~\sa12_reg[6]/NET0131  & n8110 ;
  assign n8498 = ~\sa12_reg[4]/P0001  & ~\sa12_reg[7]/NET0131  ;
  assign n8499 = n8497 & n8498 ;
  assign n8500 = ~n8421 & ~n8499 ;
  assign n8501 = ~n8496 & n8500 ;
  assign n8502 = \sa12_reg[1]/P0001  & ~n8501 ;
  assign n8490 = \sa12_reg[5]/P0001  & n8156 ;
  assign n8491 = n8057 & n8490 ;
  assign n8492 = ~n8096 & ~n8150 ;
  assign n8493 = ~\sa12_reg[2]/P0001  & ~n8492 ;
  assign n8503 = ~n8491 & ~n8493 ;
  assign n8504 = ~n8502 & n8503 ;
  assign n8505 = ~n8489 & n8504 ;
  assign n8506 = ~n8474 & n8505 ;
  assign n8507 = ~n8431 & n8506 ;
  assign n8513 = \sa23_reg[6]/NET0131  & ~\sa23_reg[7]/NET0131  ;
  assign n8514 = ~\sa23_reg[4]/P0001  & n8513 ;
  assign n8515 = ~\sa23_reg[3]/P0001  & n8514 ;
  assign n8508 = \sa23_reg[5]/P0001  & ~\sa23_reg[6]/NET0131  ;
  assign n8509 = ~\sa23_reg[3]/P0001  & n8508 ;
  assign n8510 = \sa23_reg[4]/P0001  & n8509 ;
  assign n8511 = ~\sa23_reg[6]/NET0131  & \sa23_reg[7]/NET0131  ;
  assign n8512 = \sa23_reg[3]/P0001  & n8511 ;
  assign n8516 = ~n8510 & ~n8512 ;
  assign n8517 = ~n8515 & n8516 ;
  assign n8518 = ~\sa23_reg[2]/P0001  & ~n8517 ;
  assign n8531 = \sa23_reg[5]/P0001  & \sa23_reg[7]/NET0131  ;
  assign n8532 = \sa23_reg[3]/P0001  & n8531 ;
  assign n8521 = \sa23_reg[5]/P0001  & \sa23_reg[6]/NET0131  ;
  assign n8533 = \sa23_reg[4]/P0001  & n8521 ;
  assign n8534 = ~\sa23_reg[7]/NET0131  & n8533 ;
  assign n8535 = ~n8532 & ~n8534 ;
  assign n8536 = \sa23_reg[2]/P0001  & ~n8535 ;
  assign n8522 = ~\sa23_reg[3]/P0001  & ~\sa23_reg[4]/P0001  ;
  assign n8523 = ~\sa23_reg[7]/NET0131  & n8522 ;
  assign n8524 = n8521 & n8523 ;
  assign n8519 = ~\sa23_reg[4]/P0001  & \sa23_reg[7]/NET0131  ;
  assign n8520 = n8508 & n8519 ;
  assign n8525 = ~\sa23_reg[5]/P0001  & \sa23_reg[6]/NET0131  ;
  assign n8526 = ~\sa23_reg[3]/P0001  & \sa23_reg[7]/NET0131  ;
  assign n8527 = n8525 & n8526 ;
  assign n8539 = ~n8520 & ~n8527 ;
  assign n8528 = ~\sa23_reg[6]/NET0131  & ~\sa23_reg[7]/NET0131  ;
  assign n8529 = \sa23_reg[3]/P0001  & ~\sa23_reg[5]/P0001  ;
  assign n8530 = n8528 & n8529 ;
  assign n8537 = \sa23_reg[3]/P0001  & \sa23_reg[4]/P0001  ;
  assign n8538 = n8531 & n8537 ;
  assign n8540 = ~n8530 & ~n8538 ;
  assign n8541 = n8539 & n8540 ;
  assign n8542 = ~n8524 & n8541 ;
  assign n8543 = ~n8536 & n8542 ;
  assign n8544 = ~n8518 & n8543 ;
  assign n8545 = \sa23_reg[1]/P0001  & ~n8544 ;
  assign n8550 = ~\sa23_reg[6]/NET0131  & n8526 ;
  assign n8551 = \sa23_reg[4]/P0001  & n8550 ;
  assign n8552 = ~\sa23_reg[3]/P0001  & n8528 ;
  assign n8553 = \sa23_reg[2]/P0001  & n8552 ;
  assign n8554 = ~n8551 & ~n8553 ;
  assign n8555 = ~\sa23_reg[5]/P0001  & ~n8554 ;
  assign n8546 = \sa23_reg[2]/P0001  & \sa23_reg[3]/P0001  ;
  assign n8547 = ~\sa23_reg[5]/P0001  & ~\sa23_reg[6]/NET0131  ;
  assign n8548 = ~\sa23_reg[4]/P0001  & n8547 ;
  assign n8549 = n8546 & n8548 ;
  assign n8556 = ~\sa23_reg[4]/P0001  & \sa23_reg[6]/NET0131  ;
  assign n8557 = n8531 & n8556 ;
  assign n8558 = ~\sa23_reg[3]/P0001  & n8557 ;
  assign n8559 = ~n8549 & ~n8558 ;
  assign n8560 = ~n8555 & n8559 ;
  assign n8561 = ~\sa23_reg[1]/P0001  & ~n8560 ;
  assign n8564 = ~\sa23_reg[5]/P0001  & ~\sa23_reg[7]/NET0131  ;
  assign n8572 = \sa23_reg[3]/P0001  & ~\sa23_reg[4]/P0001  ;
  assign n8573 = ~\sa23_reg[3]/P0001  & \sa23_reg[4]/P0001  ;
  assign n8574 = \sa23_reg[6]/NET0131  & n8573 ;
  assign n8575 = ~n8572 & ~n8574 ;
  assign n8576 = n8564 & ~n8575 ;
  assign n8577 = ~\sa23_reg[4]/P0001  & ~\sa23_reg[7]/NET0131  ;
  assign n8578 = ~\sa23_reg[6]/NET0131  & n8577 ;
  assign n8579 = ~n8538 & ~n8578 ;
  assign n8580 = ~n8576 & n8579 ;
  assign n8581 = \sa23_reg[2]/P0001  & ~n8580 ;
  assign n8562 = ~\sa23_reg[5]/P0001  & \sa23_reg[7]/NET0131  ;
  assign n8563 = n8556 & n8562 ;
  assign n8565 = n8537 & n8564 ;
  assign n8566 = ~n8563 & ~n8565 ;
  assign n8567 = ~\sa23_reg[2]/P0001  & ~n8566 ;
  assign n8568 = ~\sa23_reg[7]/NET0131  & n8548 ;
  assign n8569 = \sa23_reg[4]/P0001  & \sa23_reg[7]/NET0131  ;
  assign n8570 = n8508 & n8569 ;
  assign n8571 = ~\sa23_reg[2]/P0001  & n8570 ;
  assign n8582 = ~n8568 & ~n8571 ;
  assign n8583 = ~n8567 & n8582 ;
  assign n8584 = ~n8581 & n8583 ;
  assign n8585 = ~n8561 & n8584 ;
  assign n8586 = ~n8545 & n8585 ;
  assign n8587 = ~\sa23_reg[0]/P0001  & ~n8586 ;
  assign n8622 = ~\sa23_reg[4]/P0001  & n8525 ;
  assign n8623 = \sa23_reg[4]/P0001  & ~\sa23_reg[7]/NET0131  ;
  assign n8624 = \sa23_reg[3]/P0001  & ~\sa23_reg[6]/NET0131  ;
  assign n8625 = n8623 & n8624 ;
  assign n8626 = ~n8622 & ~n8625 ;
  assign n8627 = \sa23_reg[2]/P0001  & ~n8626 ;
  assign n8614 = \sa23_reg[5]/P0001  & n8513 ;
  assign n8615 = n8511 & n8529 ;
  assign n8616 = ~n8614 & ~n8615 ;
  assign n8617 = ~\sa23_reg[2]/P0001  & ~n8616 ;
  assign n8589 = \sa23_reg[5]/P0001  & ~\sa23_reg[7]/NET0131  ;
  assign n8618 = \sa23_reg[3]/P0001  & n8589 ;
  assign n8619 = n8531 & n8573 ;
  assign n8620 = ~n8618 & ~n8619 ;
  assign n8621 = \sa23_reg[6]/NET0131  & ~n8620 ;
  assign n8628 = ~n8617 & ~n8621 ;
  assign n8629 = ~n8627 & n8628 ;
  assign n8630 = ~\sa23_reg[1]/P0001  & ~n8629 ;
  assign n8631 = \sa23_reg[5]/P0001  & n8528 ;
  assign n8632 = n8537 & n8631 ;
  assign n8633 = n8509 & n8569 ;
  assign n8634 = ~n8632 & ~n8633 ;
  assign n8635 = ~\sa23_reg[7]/NET0131  & n8573 ;
  assign n8636 = n8547 & n8635 ;
  assign n8637 = ~\sa23_reg[4]/P0001  & n8512 ;
  assign n8638 = ~n8636 & ~n8637 ;
  assign n8639 = n8634 & n8638 ;
  assign n8640 = \sa23_reg[1]/P0001  & ~n8639 ;
  assign n8641 = n8531 & n8574 ;
  assign n8642 = ~\sa23_reg[3]/P0001  & n8525 ;
  assign n8643 = n8577 & n8642 ;
  assign n8644 = ~n8641 & ~n8643 ;
  assign n8645 = \sa23_reg[2]/P0001  & ~n8644 ;
  assign n8602 = n8525 & n8569 ;
  assign n8646 = ~\sa23_reg[2]/P0001  & n8602 ;
  assign n8647 = n8572 & n8614 ;
  assign n8648 = ~n8646 & ~n8647 ;
  assign n8649 = ~n8645 & n8648 ;
  assign n8650 = ~n8640 & n8649 ;
  assign n8651 = ~n8630 & n8650 ;
  assign n8652 = \sa23_reg[0]/P0001  & ~n8651 ;
  assign n8593 = \sa23_reg[5]/P0001  & n8572 ;
  assign n8594 = ~\sa23_reg[5]/P0001  & ~n8556 ;
  assign n8595 = ~n8569 & n8594 ;
  assign n8596 = ~n8593 & ~n8595 ;
  assign n8597 = \sa23_reg[1]/P0001  & ~n8596 ;
  assign n8588 = \sa23_reg[3]/P0001  & \sa23_reg[6]/NET0131  ;
  assign n8590 = n8588 & n8589 ;
  assign n8591 = n8513 & n8572 ;
  assign n8592 = ~n8590 & ~n8591 ;
  assign n8598 = ~\sa23_reg[4]/P0001  & n8589 ;
  assign n8599 = n8592 & ~n8598 ;
  assign n8600 = ~n8597 & n8599 ;
  assign n8601 = \sa23_reg[0]/P0001  & ~n8600 ;
  assign n8603 = ~\sa23_reg[3]/P0001  & n8519 ;
  assign n8604 = n8513 & n8537 ;
  assign n8605 = ~n8603 & ~n8604 ;
  assign n8606 = \sa23_reg[5]/P0001  & ~n8605 ;
  assign n8607 = ~n8602 & ~n8606 ;
  assign n8608 = ~\sa23_reg[1]/P0001  & ~n8607 ;
  assign n8609 = n8528 & n8593 ;
  assign n8610 = ~n8527 & ~n8609 ;
  assign n8611 = ~n8608 & n8610 ;
  assign n8612 = ~n8601 & n8611 ;
  assign n8613 = ~\sa23_reg[2]/P0001  & ~n8612 ;
  assign n8653 = \sa23_reg[6]/NET0131  & n8531 ;
  assign n8654 = ~\sa23_reg[5]/P0001  & n8511 ;
  assign n8655 = ~\sa23_reg[5]/P0001  & n8513 ;
  assign n8656 = ~n8654 & ~n8655 ;
  assign n8657 = ~n8653 & n8656 ;
  assign n8658 = \sa23_reg[2]/P0001  & n8573 ;
  assign n8659 = ~n8657 & n8658 ;
  assign n8660 = \sa23_reg[2]/P0001  & ~\sa23_reg[6]/NET0131  ;
  assign n8661 = \sa23_reg[5]/P0001  & n8537 ;
  assign n8662 = n8660 & n8661 ;
  assign n8663 = n8522 & n8528 ;
  assign n8664 = ~n8662 & ~n8663 ;
  assign n8665 = ~n8659 & n8664 ;
  assign n8666 = ~\sa23_reg[1]/P0001  & ~n8665 ;
  assign n8667 = n8508 & n8623 ;
  assign n8668 = n8546 & n8667 ;
  assign n8670 = n8529 & n8578 ;
  assign n8669 = n8614 & n8658 ;
  assign n8671 = ~n8571 & ~n8669 ;
  assign n8672 = ~n8670 & n8671 ;
  assign n8673 = \sa23_reg[1]/P0001  & ~n8672 ;
  assign n8674 = ~n8668 & ~n8673 ;
  assign n8675 = ~n8666 & n8674 ;
  assign n8676 = ~n8613 & n8675 ;
  assign n8677 = ~n8652 & n8676 ;
  assign n8678 = ~n8587 & n8677 ;
  assign n8679 = n8507 & ~n8678 ;
  assign n8680 = ~n8507 & n8678 ;
  assign n8681 = ~n8679 & ~n8680 ;
  assign n8697 = \sa30_reg[5]/P0001  & \sa30_reg[6]/NET0131  ;
  assign n8705 = ~\sa30_reg[7]/P0001  & n8697 ;
  assign n8682 = ~\sa30_reg[6]/NET0131  & \sa30_reg[7]/P0001  ;
  assign n8702 = \sa30_reg[3]/P0001  & ~\sa30_reg[5]/P0001  ;
  assign n8796 = n8682 & n8702 ;
  assign n8797 = ~n8705 & ~n8796 ;
  assign n8798 = ~\sa30_reg[2]/P0001  & ~n8797 ;
  assign n8695 = \sa30_reg[3]/P0001  & \sa30_reg[4]/P0001  ;
  assign n8701 = ~\sa30_reg[6]/NET0131  & ~\sa30_reg[7]/P0001  ;
  assign n8791 = n8695 & n8701 ;
  assign n8792 = ~\sa30_reg[5]/P0001  & \sa30_reg[6]/NET0131  ;
  assign n8793 = ~\sa30_reg[4]/P0001  & n8792 ;
  assign n8794 = ~n8791 & ~n8793 ;
  assign n8795 = \sa30_reg[2]/P0001  & ~n8794 ;
  assign n8756 = \sa30_reg[5]/P0001  & ~\sa30_reg[7]/P0001  ;
  assign n8758 = \sa30_reg[3]/P0001  & \sa30_reg[6]/NET0131  ;
  assign n8759 = n8756 & n8758 ;
  assign n8694 = \sa30_reg[5]/P0001  & \sa30_reg[7]/P0001  ;
  assign n8721 = ~\sa30_reg[3]/P0001  & \sa30_reg[4]/P0001  ;
  assign n8735 = \sa30_reg[6]/NET0131  & n8721 ;
  assign n8769 = n8694 & n8735 ;
  assign n8799 = ~n8759 & ~n8769 ;
  assign n8800 = ~n8795 & n8799 ;
  assign n8801 = ~n8798 & n8800 ;
  assign n8802 = ~\sa30_reg[1]/P0001  & ~n8801 ;
  assign n8780 = n8695 & n8756 ;
  assign n8781 = ~\sa30_reg[6]/NET0131  & n8780 ;
  assign n8683 = \sa30_reg[3]/P0001  & n8682 ;
  assign n8782 = ~\sa30_reg[4]/P0001  & n8683 ;
  assign n8787 = ~n8781 & ~n8782 ;
  assign n8775 = ~\sa30_reg[5]/P0001  & ~\sa30_reg[6]/NET0131  ;
  assign n8783 = ~\sa30_reg[7]/P0001  & n8721 ;
  assign n8784 = n8775 & n8783 ;
  assign n8785 = n8694 & n8721 ;
  assign n8786 = ~\sa30_reg[6]/NET0131  & n8785 ;
  assign n8788 = ~n8784 & ~n8786 ;
  assign n8789 = n8787 & n8788 ;
  assign n8790 = \sa30_reg[1]/P0001  & ~n8789 ;
  assign n8757 = ~\sa30_reg[4]/P0001  & n8756 ;
  assign n8686 = \sa30_reg[6]/NET0131  & ~\sa30_reg[7]/P0001  ;
  assign n8725 = \sa30_reg[3]/P0001  & ~\sa30_reg[4]/P0001  ;
  assign n8760 = n8686 & n8725 ;
  assign n8761 = ~n8759 & ~n8760 ;
  assign n8762 = ~n8757 & n8761 ;
  assign n8763 = ~\sa30_reg[2]/P0001  & ~n8762 ;
  assign n8764 = n8705 & n8725 ;
  assign n8709 = \sa30_reg[6]/NET0131  & \sa30_reg[7]/P0001  ;
  assign n8710 = ~\sa30_reg[5]/P0001  & n8709 ;
  assign n8741 = ~\sa30_reg[2]/P0001  & \sa30_reg[4]/P0001  ;
  assign n8765 = n8710 & n8741 ;
  assign n8803 = ~n8764 & ~n8765 ;
  assign n8804 = ~n8763 & n8803 ;
  assign n8734 = ~\sa30_reg[5]/P0001  & ~\sa30_reg[7]/P0001  ;
  assign n8766 = ~\sa30_reg[4]/P0001  & \sa30_reg[6]/NET0131  ;
  assign n8767 = n8734 & n8766 ;
  assign n8768 = ~\sa30_reg[3]/P0001  & n8767 ;
  assign n8770 = ~n8768 & ~n8769 ;
  assign n8771 = \sa30_reg[2]/P0001  & ~n8770 ;
  assign n8772 = \sa30_reg[1]/P0001  & ~\sa30_reg[2]/P0001  ;
  assign n8776 = ~\sa30_reg[4]/P0001  & n8775 ;
  assign n8773 = \sa30_reg[5]/P0001  & n8725 ;
  assign n8774 = \sa30_reg[4]/P0001  & n8734 ;
  assign n8777 = ~n8773 & ~n8774 ;
  assign n8778 = ~n8776 & n8777 ;
  assign n8779 = n8772 & ~n8778 ;
  assign n8805 = ~n8771 & ~n8779 ;
  assign n8806 = n8804 & n8805 ;
  assign n8807 = ~n8790 & n8806 ;
  assign n8808 = ~n8802 & n8807 ;
  assign n8809 = \sa30_reg[0]/P0002  & ~n8808 ;
  assign n8684 = \sa30_reg[5]/P0001  & ~\sa30_reg[6]/NET0131  ;
  assign n8685 = \sa30_reg[4]/P0001  & n8684 ;
  assign n8687 = ~\sa30_reg[4]/P0001  & n8686 ;
  assign n8688 = ~n8685 & ~n8687 ;
  assign n8689 = ~\sa30_reg[3]/P0001  & ~n8688 ;
  assign n8690 = ~n8683 & ~n8689 ;
  assign n8691 = ~\sa30_reg[2]/P0001  & ~n8690 ;
  assign n8704 = \sa30_reg[3]/P0001  & n8694 ;
  assign n8706 = \sa30_reg[4]/P0001  & n8705 ;
  assign n8707 = ~n8704 & ~n8706 ;
  assign n8708 = \sa30_reg[2]/P0001  & ~n8707 ;
  assign n8692 = \sa30_reg[7]/P0001  & n8684 ;
  assign n8693 = ~\sa30_reg[4]/P0001  & n8692 ;
  assign n8696 = n8694 & n8695 ;
  assign n8703 = n8701 & n8702 ;
  assign n8712 = ~n8696 & ~n8703 ;
  assign n8713 = ~n8693 & n8712 ;
  assign n8698 = ~\sa30_reg[3]/P0001  & ~\sa30_reg[4]/P0001  ;
  assign n8699 = n8697 & n8698 ;
  assign n8700 = ~\sa30_reg[7]/P0001  & n8699 ;
  assign n8711 = ~\sa30_reg[3]/P0001  & n8710 ;
  assign n8714 = ~n8700 & ~n8711 ;
  assign n8715 = n8713 & n8714 ;
  assign n8716 = ~n8708 & n8715 ;
  assign n8717 = ~n8691 & n8716 ;
  assign n8718 = \sa30_reg[1]/P0001  & ~n8717 ;
  assign n8719 = \sa30_reg[7]/P0001  & n8698 ;
  assign n8720 = n8697 & n8719 ;
  assign n8726 = ~\sa30_reg[6]/NET0131  & n8725 ;
  assign n8722 = n8682 & n8721 ;
  assign n8724 = ~\sa30_reg[3]/P0001  & n8701 ;
  assign n8727 = ~n8722 & ~n8724 ;
  assign n8728 = ~n8726 & n8727 ;
  assign n8723 = ~\sa30_reg[2]/P0001  & ~n8722 ;
  assign n8729 = ~\sa30_reg[5]/P0001  & ~n8723 ;
  assign n8730 = ~n8728 & n8729 ;
  assign n8731 = ~n8720 & ~n8730 ;
  assign n8732 = ~\sa30_reg[1]/P0001  & ~n8731 ;
  assign n8736 = ~n8725 & ~n8735 ;
  assign n8737 = n8734 & ~n8736 ;
  assign n8733 = ~\sa30_reg[4]/P0001  & n8701 ;
  assign n8738 = ~n8696 & ~n8733 ;
  assign n8739 = ~n8737 & n8738 ;
  assign n8740 = \sa30_reg[2]/P0001  & ~n8739 ;
  assign n8743 = ~\sa30_reg[4]/P0001  & n8709 ;
  assign n8744 = ~\sa30_reg[5]/P0001  & n8743 ;
  assign n8745 = n8695 & n8734 ;
  assign n8746 = ~n8744 & ~n8745 ;
  assign n8747 = ~\sa30_reg[2]/P0001  & ~n8746 ;
  assign n8742 = n8692 & n8741 ;
  assign n8748 = ~\sa30_reg[4]/P0001  & n8734 ;
  assign n8749 = ~\sa30_reg[6]/NET0131  & n8748 ;
  assign n8750 = ~n8742 & ~n8749 ;
  assign n8751 = ~n8747 & n8750 ;
  assign n8752 = ~n8740 & n8751 ;
  assign n8753 = ~n8732 & n8752 ;
  assign n8754 = ~n8718 & n8753 ;
  assign n8755 = ~\sa30_reg[0]/P0002  & ~n8754 ;
  assign n8823 = \sa30_reg[4]/P0001  & n8710 ;
  assign n8821 = n8695 & n8697 ;
  assign n8822 = ~\sa30_reg[7]/P0001  & n8821 ;
  assign n8824 = n8694 & n8698 ;
  assign n8825 = ~n8822 & ~n8824 ;
  assign n8826 = ~n8823 & n8825 ;
  assign n8827 = ~\sa30_reg[2]/P0001  & ~n8826 ;
  assign n8810 = n8698 & n8701 ;
  assign n8813 = ~\sa30_reg[5]/P0001  & n8682 ;
  assign n8814 = ~\sa30_reg[5]/P0001  & n8686 ;
  assign n8815 = ~n8813 & ~n8814 ;
  assign n8816 = \sa30_reg[6]/NET0131  & n8694 ;
  assign n8817 = ~\sa30_reg[3]/P0001  & ~n8816 ;
  assign n8818 = n8815 & n8817 ;
  assign n8811 = \sa30_reg[2]/P0001  & \sa30_reg[4]/P0001  ;
  assign n8812 = \sa30_reg[3]/P0001  & ~n8684 ;
  assign n8819 = n8811 & ~n8812 ;
  assign n8820 = ~n8818 & n8819 ;
  assign n8828 = ~n8810 & ~n8820 ;
  assign n8829 = ~n8827 & n8828 ;
  assign n8830 = ~\sa30_reg[1]/P0001  & ~n8829 ;
  assign n8838 = ~\sa30_reg[7]/P0001  & n8725 ;
  assign n8839 = ~\sa30_reg[5]/P0001  & n8838 ;
  assign n8840 = ~\sa30_reg[6]/NET0131  & n8839 ;
  assign n8835 = ~\sa30_reg[3]/P0001  & n8686 ;
  assign n8836 = n8811 & n8835 ;
  assign n8837 = \sa30_reg[5]/P0001  & n8836 ;
  assign n8841 = ~n8742 & ~n8837 ;
  assign n8842 = ~n8840 & n8841 ;
  assign n8843 = \sa30_reg[1]/P0001  & ~n8842 ;
  assign n8844 = \sa30_reg[2]/P0001  & \sa30_reg[3]/P0001  ;
  assign n8845 = \sa30_reg[5]/P0001  & n8701 ;
  assign n8846 = n8844 & n8845 ;
  assign n8847 = \sa30_reg[4]/P0001  & n8846 ;
  assign n8831 = n8726 & n8756 ;
  assign n8832 = ~\sa30_reg[2]/P0001  & n8831 ;
  assign n8833 = ~\sa30_reg[2]/P0001  & ~\sa30_reg[3]/P0001  ;
  assign n8834 = n8710 & n8833 ;
  assign n8848 = ~n8832 & ~n8834 ;
  assign n8849 = ~n8847 & n8848 ;
  assign n8850 = ~n8843 & n8849 ;
  assign n8851 = ~n8830 & n8850 ;
  assign n8852 = ~n8755 & n8851 ;
  assign n8853 = ~n8809 & n8852 ;
  assign n8854 = \u0_w_reg[1][29]/P0002  & ~n8853 ;
  assign n8855 = ~\u0_w_reg[1][29]/P0002  & n8853 ;
  assign n8856 = ~n8854 & ~n8855 ;
  assign n8857 = n8681 & n8856 ;
  assign n8858 = ~n8681 & ~n8856 ;
  assign n8859 = ~n8857 & ~n8858 ;
  assign n8861 = n8379 & ~n8859 ;
  assign n8860 = ~n8379 & n8859 ;
  assign n8862 = ~\ld_r_reg/P0001  & ~n8860 ;
  assign n8863 = ~n8861 & n8862 ;
  assign n8865 = ~\text_in_r_reg[93]/P0001  & \u0_w_reg[1][29]/P0002  ;
  assign n8864 = \text_in_r_reg[93]/P0001  & ~\u0_w_reg[1][29]/P0002  ;
  assign n8866 = \ld_r_reg/P0001  & ~n8864 ;
  assign n8867 = ~n8865 & n8866 ;
  assign n8868 = ~n8863 & ~n8867 ;
  assign n8896 = \sa30_reg[7]/P0001  & n8695 ;
  assign n8897 = ~n8814 & ~n8896 ;
  assign n8898 = \sa30_reg[2]/P0001  & ~n8897 ;
  assign n8894 = ~\sa30_reg[3]/P0001  & n8845 ;
  assign n8895 = ~\sa30_reg[2]/P0001  & n8894 ;
  assign n8899 = \sa30_reg[7]/P0001  & n8685 ;
  assign n8900 = ~n8895 & ~n8899 ;
  assign n8901 = ~n8898 & n8900 ;
  assign n8902 = ~n8747 & n8901 ;
  assign n8903 = ~\sa30_reg[1]/P0001  & ~n8902 ;
  assign n8874 = ~\sa30_reg[5]/P0001  & \sa30_reg[7]/P0001  ;
  assign n8875 = n8698 & n8874 ;
  assign n8876 = \sa30_reg[6]/NET0131  & n8875 ;
  assign n8873 = \sa30_reg[4]/P0001  & n8686 ;
  assign n8877 = ~n8693 & ~n8873 ;
  assign n8878 = ~n8876 & n8877 ;
  assign n8879 = \sa30_reg[2]/P0001  & ~n8878 ;
  assign n8869 = n8694 & n8725 ;
  assign n8870 = ~n8781 & ~n8869 ;
  assign n8871 = ~\sa30_reg[5]/P0001  & n8833 ;
  assign n8872 = ~n8766 & n8871 ;
  assign n8880 = n8870 & ~n8872 ;
  assign n8881 = ~n8879 & n8880 ;
  assign n8882 = \sa30_reg[1]/P0001  & ~n8881 ;
  assign n8883 = n8756 & n8766 ;
  assign n8884 = ~\sa30_reg[3]/P0001  & n8684 ;
  assign n8885 = \sa30_reg[4]/P0001  & n8884 ;
  assign n8886 = ~n8883 & ~n8885 ;
  assign n8887 = ~\sa30_reg[2]/P0001  & ~n8886 ;
  assign n8888 = \sa30_reg[3]/P0001  & n8686 ;
  assign n8889 = \sa30_reg[4]/P0001  & n8888 ;
  assign n8890 = ~n8769 & ~n8889 ;
  assign n8891 = ~n8749 & ~n8796 ;
  assign n8892 = n8890 & n8891 ;
  assign n8893 = \sa30_reg[2]/P0001  & ~n8892 ;
  assign n8904 = ~n8887 & ~n8893 ;
  assign n8905 = ~n8882 & n8904 ;
  assign n8906 = ~n8903 & n8905 ;
  assign n8907 = \sa30_reg[0]/P0002  & ~n8906 ;
  assign n8911 = ~n8705 & ~n8775 ;
  assign n8912 = n8721 & ~n8911 ;
  assign n8908 = \sa30_reg[4]/P0001  & ~n8709 ;
  assign n8909 = ~n8701 & n8702 ;
  assign n8910 = ~n8908 & n8909 ;
  assign n8913 = ~\sa30_reg[2]/P0001  & ~n8910 ;
  assign n8914 = ~n8912 & n8913 ;
  assign n8915 = n8710 & n8721 ;
  assign n8916 = n8698 & n8775 ;
  assign n8917 = \sa30_reg[2]/P0001  & ~n8916 ;
  assign n8918 = ~n8915 & n8917 ;
  assign n8919 = ~n8914 & ~n8918 ;
  assign n8923 = ~\sa30_reg[1]/P0001  & ~n8883 ;
  assign n8920 = n8682 & n8698 ;
  assign n8922 = n8725 & n8874 ;
  assign n8924 = ~n8920 & ~n8922 ;
  assign n8925 = n8923 & n8924 ;
  assign n8921 = ~\sa30_reg[2]/P0001  & n8896 ;
  assign n8926 = ~n8846 & ~n8915 ;
  assign n8927 = ~n8921 & n8926 ;
  assign n8928 = n8925 & n8927 ;
  assign n8933 = ~\sa30_reg[2]/P0001  & n8749 ;
  assign n8929 = \sa30_reg[2]/P0001  & ~\sa30_reg[3]/P0001  ;
  assign n8930 = \sa30_reg[4]/P0001  & n8694 ;
  assign n8931 = ~n8748 & ~n8930 ;
  assign n8932 = n8929 & ~n8931 ;
  assign n8934 = \sa30_reg[1]/P0001  & ~n8822 ;
  assign n8935 = ~n8932 & n8934 ;
  assign n8936 = ~n8933 & n8935 ;
  assign n8937 = ~n8928 & ~n8936 ;
  assign n8938 = ~n8919 & ~n8937 ;
  assign n8939 = ~\sa30_reg[0]/P0002  & ~n8938 ;
  assign n8960 = n8692 & ~n8698 ;
  assign n8961 = ~\sa30_reg[5]/P0001  & n8873 ;
  assign n8962 = ~n8960 & ~n8961 ;
  assign n8963 = ~\sa30_reg[2]/P0001  & ~n8962 ;
  assign n8964 = n8682 & n8695 ;
  assign n8965 = ~n8699 & ~n8964 ;
  assign n8966 = ~n8963 & n8965 ;
  assign n8967 = ~\sa30_reg[1]/P0001  & ~n8966 ;
  assign n8952 = n8694 & n8766 ;
  assign n8953 = ~\sa30_reg[7]/P0001  & n8726 ;
  assign n8954 = ~n8952 & ~n8953 ;
  assign n8955 = ~\sa30_reg[1]/P0001  & ~n8954 ;
  assign n8950 = ~\sa30_reg[5]/P0001  & n8701 ;
  assign n8951 = ~\sa30_reg[3]/P0001  & n8950 ;
  assign n8956 = n8695 & n8814 ;
  assign n8957 = ~n8951 & ~n8956 ;
  assign n8958 = ~n8955 & n8957 ;
  assign n8959 = \sa30_reg[2]/P0001  & ~n8958 ;
  assign n8943 = ~\sa30_reg[7]/P0001  & n8698 ;
  assign n8944 = ~n8774 & ~n8869 ;
  assign n8945 = ~n8943 & n8944 ;
  assign n8946 = \sa30_reg[1]/P0001  & \sa30_reg[2]/P0001  ;
  assign n8947 = ~\sa30_reg[6]/NET0131  & n8946 ;
  assign n8948 = ~n8945 & n8947 ;
  assign n8942 = n8772 & n8831 ;
  assign n8940 = ~\sa30_reg[2]/P0001  & \sa30_reg[3]/P0001  ;
  assign n8941 = n8899 & n8940 ;
  assign n8949 = n8775 & n8943 ;
  assign n8968 = ~n8941 & ~n8949 ;
  assign n8969 = ~n8942 & n8968 ;
  assign n8970 = ~n8948 & n8969 ;
  assign n8971 = ~n8959 & n8970 ;
  assign n8972 = ~n8967 & n8971 ;
  assign n8973 = ~n8939 & n8972 ;
  assign n8974 = ~n8907 & n8973 ;
  assign n8975 = \u0_w_reg[1][30]/P0001  & ~n8974 ;
  assign n8976 = ~\u0_w_reg[1][30]/P0001  & n8974 ;
  assign n8977 = ~n8975 & ~n8976 ;
  assign n8997 = ~\sa12_reg[2]/P0001  & ~n8087 ;
  assign n8998 = \sa12_reg[2]/P0001  & ~n8081 ;
  assign n8999 = ~n8412 & n8998 ;
  assign n9000 = ~n8997 & ~n8999 ;
  assign n9001 = ~n8166 & ~n8424 ;
  assign n9002 = ~n9000 & n9001 ;
  assign n9003 = ~\sa12_reg[1]/P0001  & ~n9002 ;
  assign n8981 = n8084 & n8202 ;
  assign n8982 = ~n8061 & ~n8388 ;
  assign n8983 = ~n8981 & n8982 ;
  assign n8984 = \sa12_reg[2]/P0001  & ~n8983 ;
  assign n8978 = ~\sa12_reg[2]/P0001  & ~\sa12_reg[3]/P0001  ;
  assign n8979 = ~\sa12_reg[5]/P0001  & ~n8068 ;
  assign n8980 = n8978 & n8979 ;
  assign n8985 = n8078 & n8161 ;
  assign n8986 = ~n8460 & ~n8985 ;
  assign n8987 = ~n8980 & n8986 ;
  assign n8988 = ~n8984 & n8987 ;
  assign n8989 = \sa12_reg[1]/P0001  & ~n8988 ;
  assign n8990 = n8065 & n8498 ;
  assign n8991 = ~n8380 & ~n8990 ;
  assign n8992 = ~\sa12_reg[2]/P0001  & ~n8991 ;
  assign n8993 = ~n8181 & ~n8433 ;
  assign n8994 = ~n8127 & ~n8425 ;
  assign n8995 = n8993 & n8994 ;
  assign n8996 = \sa12_reg[2]/P0001  & ~n8995 ;
  assign n9004 = ~n8992 & ~n8996 ;
  assign n9005 = ~n8989 & n9004 ;
  assign n9006 = ~n9003 & n9005 ;
  assign n9007 = \sa12_reg[0]/P0001  & ~n9006 ;
  assign n9008 = ~n8165 & ~n8414 ;
  assign n9009 = n8059 & ~n9008 ;
  assign n9010 = n8142 & n8162 ;
  assign n9011 = \sa12_reg[1]/P0001  & ~n8103 ;
  assign n9012 = ~n9010 & n9011 ;
  assign n9013 = ~n9009 & n9012 ;
  assign n9016 = ~\sa12_reg[1]/P0001  & ~n8112 ;
  assign n9014 = n8080 & n8155 ;
  assign n9017 = ~n8990 & ~n9014 ;
  assign n9018 = n9016 & n9017 ;
  assign n9015 = ~\sa12_reg[6]/NET0131  & n8085 ;
  assign n9019 = ~n8058 & ~n8177 ;
  assign n9020 = ~n9015 & n9019 ;
  assign n9021 = n9018 & n9020 ;
  assign n9022 = ~n9013 & ~n9021 ;
  assign n9023 = \sa12_reg[2]/P0001  & ~n8117 ;
  assign n9024 = ~n8177 & n9023 ;
  assign n9025 = \sa12_reg[4]/P0001  & n8082 ;
  assign n9026 = ~n8116 & ~n9025 ;
  assign n9027 = ~n8180 & ~n9026 ;
  assign n9028 = n8137 & ~n8495 ;
  assign n9029 = ~n9027 & n9028 ;
  assign n9030 = ~n9024 & ~n9029 ;
  assign n9031 = ~n9022 & ~n9030 ;
  assign n9032 = ~\sa12_reg[0]/P0001  & ~n9031 ;
  assign n9048 = ~n8104 & n8185 ;
  assign n9049 = n8069 & n8390 ;
  assign n9050 = ~n9048 & ~n9049 ;
  assign n9051 = ~\sa12_reg[2]/P0001  & ~n9050 ;
  assign n9044 = n8068 & n8161 ;
  assign n9045 = ~n8195 & ~n9044 ;
  assign n9046 = \sa12_reg[2]/P0001  & ~n9045 ;
  assign n9047 = n8126 & n8180 ;
  assign n9052 = ~n8394 & ~n9047 ;
  assign n9053 = ~n9046 & n9052 ;
  assign n9054 = ~n9051 & n9053 ;
  assign n9055 = ~\sa12_reg[1]/P0001  & ~n9054 ;
  assign n9033 = \sa12_reg[1]/P0001  & \sa12_reg[2]/P0001  ;
  assign n9035 = \sa12_reg[5]/P0001  & n8381 ;
  assign n9036 = ~\sa12_reg[4]/P0001  & n9035 ;
  assign n9034 = \sa12_reg[4]/P0001  & n8142 ;
  assign n9037 = ~n8485 & ~n9034 ;
  assign n9038 = ~n9036 & n9037 ;
  assign n9039 = n9033 & ~n9038 ;
  assign n9042 = n8069 & n8075 ;
  assign n9043 = n8066 & n9042 ;
  assign n9056 = ~n8118 & ~n9043 ;
  assign n9057 = ~n8408 & n9056 ;
  assign n9040 = n8150 & n8455 ;
  assign n9041 = n8155 & n8166 ;
  assign n9058 = ~n9040 & ~n9041 ;
  assign n9059 = n9057 & n9058 ;
  assign n9060 = ~n9039 & n9059 ;
  assign n9061 = ~n9055 & n9060 ;
  assign n9062 = ~n9032 & n9061 ;
  assign n9063 = ~n9007 & n9062 ;
  assign n9074 = n8525 & n8603 ;
  assign n9073 = \sa23_reg[4]/P0001  & n8513 ;
  assign n9075 = ~n8520 & ~n9073 ;
  assign n9076 = ~n9074 & n9075 ;
  assign n9077 = \sa23_reg[2]/P0001  & ~n9076 ;
  assign n9079 = ~\sa23_reg[2]/P0001  & ~\sa23_reg[3]/P0001  ;
  assign n9080 = n8594 & n9079 ;
  assign n9078 = n8531 & n8572 ;
  assign n9081 = ~n8632 & ~n9078 ;
  assign n9082 = ~n9080 & n9081 ;
  assign n9083 = ~n9077 & n9082 ;
  assign n9084 = \sa23_reg[1]/P0001  & ~n9083 ;
  assign n9069 = ~n8567 & ~n8570 ;
  assign n9064 = ~\sa23_reg[3]/P0001  & n8631 ;
  assign n9065 = ~\sa23_reg[2]/P0001  & n9064 ;
  assign n9066 = \sa23_reg[3]/P0001  & n8569 ;
  assign n9067 = ~n8655 & ~n9066 ;
  assign n9068 = \sa23_reg[2]/P0001  & ~n9067 ;
  assign n9070 = ~n9065 & ~n9068 ;
  assign n9071 = n9069 & n9070 ;
  assign n9072 = ~\sa23_reg[1]/P0001  & ~n9071 ;
  assign n9085 = n8521 & n8577 ;
  assign n9086 = ~n8510 & ~n9085 ;
  assign n9087 = ~\sa23_reg[2]/P0001  & ~n9086 ;
  assign n9088 = ~n8604 & ~n8641 ;
  assign n9089 = ~n8568 & ~n8615 ;
  assign n9090 = n9088 & n9089 ;
  assign n9091 = \sa23_reg[2]/P0001  & ~n9090 ;
  assign n9092 = ~n9087 & ~n9091 ;
  assign n9093 = ~n9072 & n9092 ;
  assign n9094 = ~n9084 & n9093 ;
  assign n9095 = \sa23_reg[0]/P0001  & ~n9094 ;
  assign n9139 = n8519 & n8529 ;
  assign n9138 = n8511 & n8522 ;
  assign n9142 = ~n9085 & ~n9138 ;
  assign n9143 = ~n9139 & n9142 ;
  assign n9141 = n8618 & n8660 ;
  assign n9107 = ~\sa23_reg[3]/P0001  & n8602 ;
  assign n9140 = ~\sa23_reg[2]/P0001  & n9066 ;
  assign n9144 = ~n9107 & ~n9140 ;
  assign n9145 = ~n9141 & n9144 ;
  assign n9146 = n9143 & n9145 ;
  assign n9147 = ~\sa23_reg[0]/P0001  & ~n9146 ;
  assign n9148 = \sa23_reg[2]/P0001  & ~n8557 ;
  assign n9149 = n8577 & n8624 ;
  assign n9150 = n9148 & ~n9149 ;
  assign n9151 = \sa23_reg[4]/P0001  & n8525 ;
  assign n9152 = ~\sa23_reg[7]/NET0131  & n9151 ;
  assign n9153 = ~\sa23_reg[2]/P0001  & ~n9152 ;
  assign n9154 = ~\sa23_reg[6]/NET0131  & n8532 ;
  assign n9155 = ~n8570 & ~n9154 ;
  assign n9156 = n9153 & n9155 ;
  assign n9157 = ~n9150 & ~n9156 ;
  assign n9158 = n8521 & n8522 ;
  assign n9159 = n8569 & n8624 ;
  assign n9160 = ~n9158 & ~n9159 ;
  assign n9161 = ~n9157 & n9160 ;
  assign n9162 = ~n9147 & n9161 ;
  assign n9163 = ~\sa23_reg[1]/P0001  & ~n9162 ;
  assign n9096 = \sa23_reg[7]/NET0131  & n8588 ;
  assign n9097 = ~\sa23_reg[5]/P0001  & n9096 ;
  assign n9098 = ~\sa23_reg[2]/P0001  & ~n9097 ;
  assign n9101 = n8574 & n8589 ;
  assign n9099 = \sa23_reg[4]/P0001  & n8547 ;
  assign n9100 = ~n8528 & n8529 ;
  assign n9102 = ~n9099 & ~n9100 ;
  assign n9103 = ~n9101 & n9102 ;
  assign n9104 = ~n8537 & ~n9103 ;
  assign n9105 = n9098 & ~n9104 ;
  assign n9106 = n8522 & n8547 ;
  assign n9108 = \sa23_reg[2]/P0001  & ~n9106 ;
  assign n9109 = ~n9107 & n9108 ;
  assign n9110 = ~n9105 & ~n9109 ;
  assign n9112 = \sa23_reg[2]/P0001  & ~\sa23_reg[3]/P0001  ;
  assign n9113 = \sa23_reg[4]/P0001  & n8531 ;
  assign n9114 = ~\sa23_reg[4]/P0001  & n8564 ;
  assign n9115 = ~n9113 & ~n9114 ;
  assign n9116 = n9112 & ~n9115 ;
  assign n9111 = ~\sa23_reg[2]/P0001  & n8568 ;
  assign n9117 = n8537 & n8614 ;
  assign n9118 = ~n9111 & ~n9117 ;
  assign n9119 = ~n9116 & n9118 ;
  assign n9120 = \sa23_reg[1]/P0001  & ~n9119 ;
  assign n9121 = ~n9110 & ~n9120 ;
  assign n9122 = ~\sa23_reg[0]/P0001  & ~n9121 ;
  assign n9123 = ~n8523 & ~n9078 ;
  assign n9124 = ~\sa23_reg[6]/NET0131  & ~n9123 ;
  assign n9125 = ~\sa23_reg[7]/NET0131  & n9099 ;
  assign n9126 = ~n9124 & ~n9125 ;
  assign n9127 = \sa23_reg[1]/P0001  & ~n9126 ;
  assign n9128 = ~\sa23_reg[5]/P0001  & n8552 ;
  assign n9129 = n8525 & n8537 ;
  assign n9130 = ~\sa23_reg[7]/NET0131  & n9129 ;
  assign n9131 = ~n9128 & ~n9130 ;
  assign n9132 = ~n9127 & n9131 ;
  assign n9133 = \sa23_reg[2]/P0001  & ~n9132 ;
  assign n9135 = ~\sa23_reg[2]/P0001  & n8609 ;
  assign n9136 = \sa23_reg[1]/P0001  & n9135 ;
  assign n9134 = \sa23_reg[3]/P0001  & n8571 ;
  assign n9137 = n8523 & n8547 ;
  assign n9164 = ~n9134 & ~n9137 ;
  assign n9165 = ~n9136 & n9164 ;
  assign n9166 = ~n9133 & n9165 ;
  assign n9167 = ~n9122 & n9166 ;
  assign n9168 = ~n9163 & n9167 ;
  assign n9169 = ~n9095 & n9168 ;
  assign n9170 = n9063 & ~n9169 ;
  assign n9171 = ~n9063 & n9169 ;
  assign n9172 = ~n9170 & ~n9171 ;
  assign n9244 = ~\sa01_reg[2]/P0001  & ~n8277 ;
  assign n9245 = ~n8255 & n9244 ;
  assign n9246 = ~\sa01_reg[5]/P0001  & n8225 ;
  assign n9247 = \sa01_reg[2]/P0001  & ~n8305 ;
  assign n9248 = ~n9246 & n9247 ;
  assign n9249 = ~n9245 & ~n9248 ;
  assign n9243 = n8214 & n8258 ;
  assign n9250 = ~n8343 & ~n9243 ;
  assign n9251 = ~n9249 & n9250 ;
  assign n9252 = ~\sa01_reg[1]/P0001  & ~n9251 ;
  assign n9228 = ~\sa01_reg[5]/P0001  & n8226 ;
  assign n9229 = ~n8354 & ~n9228 ;
  assign n9230 = \sa01_reg[1]/P0001  & ~n9229 ;
  assign n9231 = ~\sa01_reg[4]/P0001  & n8342 ;
  assign n9232 = ~n8266 & ~n8343 ;
  assign n9233 = ~n9231 & n9232 ;
  assign n9234 = ~n9230 & n9233 ;
  assign n9235 = ~\sa01_reg[2]/P0001  & ~n9234 ;
  assign n9236 = ~\sa01_reg[6]/NET0131  & n8360 ;
  assign n9239 = ~n8217 & ~n9236 ;
  assign n9237 = n8214 & n8279 ;
  assign n9238 = \sa01_reg[7]/NET0131  & n8256 ;
  assign n9240 = ~n9237 & ~n9238 ;
  assign n9241 = n9239 & n9240 ;
  assign n9242 = \sa01_reg[1]/P0001  & ~n9241 ;
  assign n9253 = n8304 & n8368 ;
  assign n9254 = ~n9243 & ~n9253 ;
  assign n9255 = \sa01_reg[2]/P0001  & ~n9254 ;
  assign n9256 = n8276 & n8354 ;
  assign n9257 = ~n8312 & ~n9256 ;
  assign n9258 = ~n9255 & n9257 ;
  assign n9259 = ~n9242 & n9258 ;
  assign n9260 = ~n9235 & n9259 ;
  assign n9261 = ~n9252 & n9260 ;
  assign n9262 = \sa01_reg[0]/P0001  & ~n9261 ;
  assign n9184 = ~\sa01_reg[3]/P0001  & n8242 ;
  assign n9185 = \sa01_reg[4]/P0001  & n9184 ;
  assign n9182 = ~\sa01_reg[7]/NET0131  & n8304 ;
  assign n9183 = \sa01_reg[3]/P0001  & n8221 ;
  assign n9186 = ~n9182 & ~n9183 ;
  assign n9187 = ~n9185 & n9186 ;
  assign n9188 = ~\sa01_reg[2]/P0001  & ~n9187 ;
  assign n9173 = \sa01_reg[3]/P0001  & n8245 ;
  assign n9175 = \sa01_reg[4]/P0001  & n8276 ;
  assign n9176 = \sa01_reg[5]/P0001  & n9175 ;
  assign n9177 = ~n9173 & ~n9176 ;
  assign n9178 = \sa01_reg[2]/P0001  & ~n9177 ;
  assign n9180 = n8221 & n8308 ;
  assign n9179 = n8253 & n8368 ;
  assign n9189 = ~n8352 & ~n9179 ;
  assign n9190 = ~n9180 & n9189 ;
  assign n9174 = \sa01_reg[4]/P0001  & n9173 ;
  assign n9181 = n8267 & n8277 ;
  assign n9191 = ~n9174 & ~n9181 ;
  assign n9192 = n9190 & n9191 ;
  assign n9193 = ~n9178 & n9192 ;
  assign n9194 = ~n9188 & n9193 ;
  assign n9195 = \sa01_reg[1]/P0001  & ~n9194 ;
  assign n9196 = n8214 & n8221 ;
  assign n9197 = \sa01_reg[2]/P0001  & ~\sa01_reg[3]/P0001  ;
  assign n9198 = n8215 & n9197 ;
  assign n9199 = ~n9196 & ~n9198 ;
  assign n9200 = ~\sa01_reg[5]/P0001  & ~n9199 ;
  assign n9201 = ~\sa01_reg[4]/P0001  & n8227 ;
  assign n9202 = n8329 & n9201 ;
  assign n9203 = ~n8322 & ~n9202 ;
  assign n9204 = ~n9200 & n9203 ;
  assign n9205 = ~\sa01_reg[1]/P0001  & ~n9204 ;
  assign n9209 = ~\sa01_reg[2]/P0001  & \sa01_reg[4]/P0001  ;
  assign n9210 = n8279 & n9209 ;
  assign n9206 = ~\sa01_reg[5]/P0001  & n8276 ;
  assign n9207 = n8287 & n9206 ;
  assign n9208 = n8215 & n8222 ;
  assign n9219 = n8227 & n8265 ;
  assign n9220 = ~n9208 & ~n9219 ;
  assign n9221 = ~n9207 & n9220 ;
  assign n9222 = ~n9210 & n9221 ;
  assign n9211 = n8238 & n8368 ;
  assign n9212 = n8225 & n8254 ;
  assign n9213 = ~n9211 & ~n9212 ;
  assign n9214 = ~\sa01_reg[2]/P0001  & ~n9213 ;
  assign n9215 = \sa01_reg[4]/P0001  & n8245 ;
  assign n9216 = ~\sa01_reg[4]/P0001  & n8368 ;
  assign n9217 = ~n9215 & ~n9216 ;
  assign n9218 = n8329 & ~n9217 ;
  assign n9223 = ~n9214 & ~n9218 ;
  assign n9224 = n9222 & n9223 ;
  assign n9225 = ~n9205 & n9224 ;
  assign n9226 = ~n9195 & n9225 ;
  assign n9227 = ~\sa01_reg[0]/P0001  & ~n9226 ;
  assign n9268 = \sa01_reg[6]/NET0131  & n8331 ;
  assign n9269 = ~n8321 & ~n8361 ;
  assign n9270 = ~n9268 & n9269 ;
  assign n9271 = ~\sa01_reg[2]/P0001  & ~n9270 ;
  assign n9263 = ~n8344 & ~n9206 ;
  assign n9264 = ~n8258 & n9263 ;
  assign n9265 = n8287 & ~n9264 ;
  assign n9266 = \sa01_reg[5]/P0001  & n8253 ;
  assign n9267 = n8327 & n9266 ;
  assign n9272 = ~n8362 & ~n9267 ;
  assign n9273 = ~n9265 & n9272 ;
  assign n9274 = ~n9271 & n9273 ;
  assign n9275 = ~\sa01_reg[1]/P0001  & ~n9274 ;
  assign n9281 = n8253 & n9216 ;
  assign n9280 = n8277 & n8287 ;
  assign n9282 = ~n9210 & ~n9280 ;
  assign n9283 = ~n9281 & n9282 ;
  assign n9284 = \sa01_reg[1]/P0001  & ~n9283 ;
  assign n9276 = \sa01_reg[4]/P0001  & n8219 ;
  assign n9277 = n8329 & n9276 ;
  assign n9278 = ~n8220 & ~n8352 ;
  assign n9279 = ~\sa01_reg[2]/P0001  & ~n9278 ;
  assign n9285 = ~n9277 & ~n9279 ;
  assign n9286 = ~n9284 & n9285 ;
  assign n9287 = ~n9275 & n9286 ;
  assign n9288 = ~n9227 & n9287 ;
  assign n9289 = ~n9262 & n9288 ;
  assign n9290 = n8507 & ~n9289 ;
  assign n9291 = ~n8507 & n9289 ;
  assign n9292 = ~n9290 & ~n9291 ;
  assign n9293 = n9172 & n9292 ;
  assign n9294 = ~n9172 & ~n9292 ;
  assign n9295 = ~n9293 & ~n9294 ;
  assign n9297 = n8977 & ~n9295 ;
  assign n9296 = ~n8977 & n9295 ;
  assign n9298 = ~\ld_r_reg/P0001  & ~n9296 ;
  assign n9299 = ~n9297 & n9298 ;
  assign n9301 = ~\text_in_r_reg[94]/P0001  & \u0_w_reg[1][30]/P0001  ;
  assign n9300 = \text_in_r_reg[94]/P0001  & ~\u0_w_reg[1][30]/P0001  ;
  assign n9302 = \ld_r_reg/P0001  & ~n9300 ;
  assign n9303 = ~n9301 & n9302 ;
  assign n9304 = ~n9299 & ~n9303 ;
  assign n9324 = n8254 & n8304 ;
  assign n9325 = ~n9175 & ~n9180 ;
  assign n9326 = ~n9324 & n9325 ;
  assign n9327 = \sa01_reg[1]/P0001  & ~n9326 ;
  assign n9323 = ~n8286 & ~n9243 ;
  assign n9328 = ~n9219 & n9323 ;
  assign n9329 = ~n9327 & n9328 ;
  assign n9330 = \sa01_reg[2]/P0001  & ~n9329 ;
  assign n9310 = \sa01_reg[1]/P0001  & ~n8225 ;
  assign n9311 = n8351 & n9310 ;
  assign n9309 = n8276 & n8308 ;
  assign n9312 = ~n9185 & ~n9309 ;
  assign n9313 = ~n9311 & n9312 ;
  assign n9314 = ~\sa01_reg[2]/P0001  & ~n9313 ;
  assign n9305 = n8240 & n9184 ;
  assign n9306 = ~n8243 & ~n9305 ;
  assign n9307 = ~n9214 & n9306 ;
  assign n9308 = ~\sa01_reg[1]/P0001  & ~n9307 ;
  assign n9315 = n8218 & n8245 ;
  assign n9316 = ~n9236 & ~n9315 ;
  assign n9317 = \sa01_reg[1]/P0001  & ~n9316 ;
  assign n9318 = ~\sa01_reg[1]/P0001  & \sa01_reg[2]/P0001  ;
  assign n9319 = \sa01_reg[3]/P0001  & n8224 ;
  assign n9320 = ~n9206 & ~n9319 ;
  assign n9321 = n9318 & ~n9320 ;
  assign n9322 = n8329 & n8344 ;
  assign n9331 = ~n9321 & ~n9322 ;
  assign n9332 = ~n9317 & n9331 ;
  assign n9333 = ~n9308 & n9332 ;
  assign n9334 = ~n9314 & n9333 ;
  assign n9335 = ~n9330 & n9334 ;
  assign n9336 = \sa01_reg[0]/P0001  & ~n9335 ;
  assign n9339 = ~n8282 & ~n8311 ;
  assign n9340 = \sa01_reg[3]/P0001  & ~n9339 ;
  assign n9337 = n8221 & n8267 ;
  assign n9341 = ~\sa01_reg[1]/P0001  & ~n9309 ;
  assign n9342 = ~n9337 & n9341 ;
  assign n9338 = \sa01_reg[7]/NET0131  & n8356 ;
  assign n9343 = ~n8330 & ~n9338 ;
  assign n9344 = n9342 & n9343 ;
  assign n9345 = ~n9340 & n9344 ;
  assign n9346 = n9197 & ~n9217 ;
  assign n9347 = ~\sa01_reg[2]/P0001  & n9219 ;
  assign n9348 = \sa01_reg[1]/P0001  & ~n8361 ;
  assign n9349 = ~n9347 & n9348 ;
  assign n9350 = ~n9346 & n9349 ;
  assign n9351 = ~n9345 & ~n9350 ;
  assign n9352 = \sa01_reg[4]/P0001  & n8227 ;
  assign n9353 = ~\sa01_reg[3]/P0001  & n9352 ;
  assign n9358 = ~\sa01_reg[2]/P0001  & ~n9353 ;
  assign n9354 = \sa01_reg[4]/P0001  & ~n8235 ;
  assign n9355 = n8319 & ~n9354 ;
  assign n9356 = n8214 & n8342 ;
  assign n9357 = \sa01_reg[6]/NET0131  & n9356 ;
  assign n9359 = ~n9355 & ~n9357 ;
  assign n9360 = n9358 & n9359 ;
  assign n9361 = ~\sa01_reg[3]/P0001  & n9201 ;
  assign n9362 = \sa01_reg[2]/P0001  & ~n9338 ;
  assign n9363 = ~n9361 & n9362 ;
  assign n9364 = ~n9360 & ~n9363 ;
  assign n9365 = ~n9351 & ~n9364 ;
  assign n9366 = ~\sa01_reg[0]/P0001  & ~n9365 ;
  assign n9369 = ~\sa01_reg[6]/NET0131  & n9173 ;
  assign n9368 = ~\sa01_reg[5]/P0001  & n9175 ;
  assign n9370 = ~n8243 & ~n9368 ;
  assign n9371 = ~n9369 & n9370 ;
  assign n9372 = ~\sa01_reg[2]/P0001  & ~n9371 ;
  assign n9373 = n8235 & n8308 ;
  assign n9374 = \sa01_reg[2]/P0001  & n9373 ;
  assign n9367 = \sa01_reg[3]/P0001  & n9208 ;
  assign n9375 = n8224 & n8253 ;
  assign n9376 = n8257 & n8267 ;
  assign n9377 = ~n9375 & ~n9376 ;
  assign n9378 = ~n9367 & n9377 ;
  assign n9379 = ~n9374 & n9378 ;
  assign n9380 = ~n9372 & n9379 ;
  assign n9381 = ~\sa01_reg[1]/P0001  & ~n9380 ;
  assign n9388 = \sa01_reg[1]/P0001  & \sa01_reg[2]/P0001  ;
  assign n9390 = ~\sa01_reg[4]/P0001  & n9369 ;
  assign n9389 = \sa01_reg[4]/P0001  & n8216 ;
  assign n9391 = ~n8362 & ~n9389 ;
  assign n9392 = ~n9390 & n9391 ;
  assign n9393 = n9388 & ~n9392 ;
  assign n9384 = ~n8286 & ~n8339 ;
  assign n9385 = n8303 & ~n9384 ;
  assign n9382 = \sa01_reg[1]/P0001  & ~\sa01_reg[2]/P0001  ;
  assign n9383 = n8220 & n9382 ;
  assign n9386 = ~\sa01_reg[2]/P0001  & \sa01_reg[3]/P0001  ;
  assign n9387 = n8243 & n9386 ;
  assign n9394 = ~n8268 & ~n9387 ;
  assign n9395 = ~n9383 & n9394 ;
  assign n9396 = ~n9385 & n9395 ;
  assign n9397 = ~n9393 & n9396 ;
  assign n9398 = ~n9381 & n9397 ;
  assign n9399 = ~n9366 & n9398 ;
  assign n9400 = ~n9336 & n9399 ;
  assign n9401 = ~n8681 & ~n9400 ;
  assign n9402 = n8681 & n9400 ;
  assign n9403 = ~n9401 & ~n9402 ;
  assign n9404 = \u0_w_reg[1][22]/P0001  & ~n8974 ;
  assign n9405 = ~\u0_w_reg[1][22]/P0001  & n8974 ;
  assign n9406 = ~n9404 & ~n9405 ;
  assign n9407 = n9169 & n9406 ;
  assign n9408 = ~n9169 & ~n9406 ;
  assign n9409 = ~n9407 & ~n9408 ;
  assign n9411 = n9403 & n9409 ;
  assign n9410 = ~n9403 & ~n9409 ;
  assign n9412 = ~\ld_r_reg/P0001  & ~n9410 ;
  assign n9413 = ~n9411 & n9412 ;
  assign n9415 = ~\text_in_r_reg[86]/P0001  & \u0_w_reg[1][22]/P0001  ;
  assign n9414 = \text_in_r_reg[86]/P0001  & ~\u0_w_reg[1][22]/P0001  ;
  assign n9416 = \ld_r_reg/P0001  & ~n9414 ;
  assign n9417 = ~n9415 & n9416 ;
  assign n9418 = ~n9413 & ~n9417 ;
  assign n9497 = \sa23_reg[2]/P0001  & ~n8614 ;
  assign n9499 = \sa23_reg[5]/P0001  & n8511 ;
  assign n9500 = ~n8572 & n9499 ;
  assign n9498 = n8519 & n8547 ;
  assign n9501 = ~\sa23_reg[2]/P0001  & ~n9498 ;
  assign n9502 = ~n9500 & n9501 ;
  assign n9503 = ~n9497 & ~n9502 ;
  assign n9504 = n8562 & n8658 ;
  assign n9505 = ~n8604 & ~n9504 ;
  assign n9506 = ~n9503 & n9505 ;
  assign n9507 = \sa23_reg[1]/P0001  & ~n9506 ;
  assign n9492 = ~\sa23_reg[3]/P0001  & n8614 ;
  assign n9493 = ~\sa23_reg[2]/P0001  & n9492 ;
  assign n9489 = ~\sa23_reg[5]/P0001  & n8528 ;
  assign n9490 = ~n8533 & ~n9489 ;
  assign n9491 = \sa23_reg[2]/P0001  & ~n9490 ;
  assign n9494 = ~n9149 & ~n9491 ;
  assign n9495 = ~n9493 & n9494 ;
  assign n9496 = ~\sa23_reg[1]/P0001  & ~n9495 ;
  assign n9482 = n8508 & n8577 ;
  assign n9483 = ~n8646 & ~n9482 ;
  assign n9484 = ~\sa23_reg[3]/P0001  & ~n9483 ;
  assign n9485 = ~\sa23_reg[5]/P0001  & n8625 ;
  assign n9486 = ~\sa23_reg[4]/P0001  & n8642 ;
  assign n9487 = ~n9485 & ~n9486 ;
  assign n9488 = \sa23_reg[2]/P0001  & ~n9487 ;
  assign n9508 = ~n9484 & ~n9488 ;
  assign n9509 = ~n9496 & n9508 ;
  assign n9510 = ~n9507 & n9509 ;
  assign n9511 = ~\sa23_reg[0]/P0001  & ~n9510 ;
  assign n9464 = n8508 & n8523 ;
  assign n9468 = ~\sa23_reg[5]/P0001  & n8603 ;
  assign n9469 = ~\sa23_reg[6]/NET0131  & n9468 ;
  assign n9466 = n8508 & n8572 ;
  assign n9470 = ~n9064 & ~n9466 ;
  assign n9465 = \sa23_reg[2]/P0001  & ~n8590 ;
  assign n9467 = n8547 & n9066 ;
  assign n9471 = n9465 & ~n9467 ;
  assign n9472 = n9470 & n9471 ;
  assign n9473 = ~n9469 & n9472 ;
  assign n9474 = ~\sa23_reg[2]/P0001  & ~n9117 ;
  assign n9475 = ~n8577 & n8642 ;
  assign n9476 = \sa23_reg[6]/NET0131  & n9078 ;
  assign n9477 = ~n9475 & ~n9476 ;
  assign n9478 = n9474 & n9477 ;
  assign n9479 = ~n9473 & ~n9478 ;
  assign n9480 = ~n9464 & ~n9479 ;
  assign n9481 = ~\sa23_reg[1]/P0001  & ~n9480 ;
  assign n9420 = n8547 & n8569 ;
  assign n9421 = ~n8514 & ~n9420 ;
  assign n9422 = ~\sa23_reg[2]/P0001  & ~n9421 ;
  assign n9419 = n8519 & n8660 ;
  assign n9423 = \sa23_reg[1]/P0001  & ~n9419 ;
  assign n9424 = ~n8609 & n9423 ;
  assign n9425 = ~n8636 & n9424 ;
  assign n9426 = ~n9422 & n9425 ;
  assign n9431 = ~\sa23_reg[2]/P0001  & n8625 ;
  assign n9432 = ~\sa23_reg[1]/P0001  & ~n9431 ;
  assign n9433 = \sa23_reg[2]/P0001  & n8570 ;
  assign n9427 = ~\sa23_reg[2]/P0001  & ~\sa23_reg[4]/P0001  ;
  assign n9428 = ~\sa23_reg[3]/P0001  & ~n9427 ;
  assign n9429 = n8531 & ~n9428 ;
  assign n9430 = n8519 & n8588 ;
  assign n9434 = ~n9429 & ~n9430 ;
  assign n9435 = ~n9433 & n9434 ;
  assign n9436 = n9432 & n9435 ;
  assign n9437 = ~n9426 & ~n9436 ;
  assign n9439 = ~n8624 & ~n8653 ;
  assign n9440 = ~\sa23_reg[4]/P0001  & ~n9439 ;
  assign n9438 = \sa23_reg[2]/P0001  & ~n8615 ;
  assign n9441 = ~n8635 & n9438 ;
  assign n9442 = ~n9440 & n9441 ;
  assign n9443 = ~n8591 & ~n9137 ;
  assign n9444 = n9098 & n9443 ;
  assign n9445 = ~n9442 & ~n9444 ;
  assign n9446 = ~n9437 & ~n9445 ;
  assign n9447 = \sa23_reg[0]/P0001  & ~n9446 ;
  assign n9448 = ~n8558 & ~n9100 ;
  assign n9449 = ~n9137 & n9448 ;
  assign n9450 = ~\sa23_reg[2]/P0001  & ~n9449 ;
  assign n9451 = n8513 & n9112 ;
  assign n9452 = \sa23_reg[4]/P0001  & n9451 ;
  assign n9456 = ~n9141 & ~n9452 ;
  assign n9453 = ~\sa23_reg[5]/P0001  & n8519 ;
  assign n9454 = n8624 & n9453 ;
  assign n9455 = \sa23_reg[7]/NET0131  & n9129 ;
  assign n9457 = ~n9454 & ~n9455 ;
  assign n9458 = n9456 & n9457 ;
  assign n9459 = ~n9450 & n9458 ;
  assign n9460 = \sa23_reg[1]/P0001  & ~n9459 ;
  assign n9461 = n8533 & n8546 ;
  assign n9462 = n8514 & n8529 ;
  assign n9463 = ~\sa23_reg[2]/P0001  & n9462 ;
  assign n9512 = ~n9461 & ~n9463 ;
  assign n9513 = ~n9460 & n9512 ;
  assign n9514 = ~n9447 & n9513 ;
  assign n9515 = ~n9481 & n9514 ;
  assign n9516 = ~n9511 & n9515 ;
  assign n9517 = n8213 & ~n9516 ;
  assign n9518 = ~n8213 & n9516 ;
  assign n9519 = ~n9517 & ~n9518 ;
  assign n9520 = ~n9289 & ~n9519 ;
  assign n9521 = n9289 & n9519 ;
  assign n9522 = ~n9520 & ~n9521 ;
  assign n9523 = \u0_w_reg[1][21]/P0001  & ~n8853 ;
  assign n9524 = ~\u0_w_reg[1][21]/P0001  & n8853 ;
  assign n9525 = ~n9523 & ~n9524 ;
  assign n9526 = n8678 & n9525 ;
  assign n9527 = ~n8678 & ~n9525 ;
  assign n9528 = ~n9526 & ~n9527 ;
  assign n9530 = n9522 & n9528 ;
  assign n9529 = ~n9522 & ~n9528 ;
  assign n9531 = ~\ld_r_reg/P0001  & ~n9529 ;
  assign n9532 = ~n9530 & n9531 ;
  assign n9534 = ~\text_in_r_reg[85]/P0001  & \u0_w_reg[1][21]/P0001  ;
  assign n9533 = \text_in_r_reg[85]/P0001  & ~\u0_w_reg[1][21]/P0001  ;
  assign n9535 = \ld_r_reg/P0001  & ~n9533 ;
  assign n9536 = ~n9534 & n9535 ;
  assign n9537 = ~n9532 & ~n9536 ;
  assign n9538 = ~n9292 & ~n9516 ;
  assign n9539 = n9292 & n9516 ;
  assign n9540 = ~n9538 & ~n9539 ;
  assign n9572 = \sa30_reg[4]/P0001  & n8813 ;
  assign n9573 = ~n8687 & ~n9572 ;
  assign n9574 = ~\sa30_reg[2]/P0001  & ~n9573 ;
  assign n9575 = \sa30_reg[2]/P0001  & ~\sa30_reg[4]/P0001  ;
  assign n9576 = n8682 & n9575 ;
  assign n9577 = \sa30_reg[1]/P0001  & ~n9576 ;
  assign n9578 = ~n8784 & n9577 ;
  assign n9579 = ~n8831 & n9578 ;
  assign n9580 = ~n9574 & n9579 ;
  assign n9586 = \sa30_reg[3]/P0001  & n8743 ;
  assign n9587 = ~\sa30_reg[1]/P0001  & ~n9586 ;
  assign n9585 = n8692 & n8811 ;
  assign n9581 = ~\sa30_reg[2]/P0001  & n8791 ;
  assign n9582 = ~\sa30_reg[2]/P0001  & ~\sa30_reg[4]/P0001  ;
  assign n9583 = ~\sa30_reg[3]/P0001  & ~n9582 ;
  assign n9584 = n8694 & ~n9583 ;
  assign n9588 = ~n9581 & ~n9584 ;
  assign n9589 = ~n9585 & n9588 ;
  assign n9590 = n9587 & n9589 ;
  assign n9591 = ~n9580 & ~n9590 ;
  assign n9592 = \sa30_reg[2]/P0001  & ~n8796 ;
  assign n9593 = ~n8726 & ~n8783 ;
  assign n9594 = ~n8952 & n9593 ;
  assign n9595 = n9592 & n9594 ;
  assign n9596 = n8758 & n8874 ;
  assign n9597 = ~\sa30_reg[2]/P0001  & ~n8760 ;
  assign n9598 = ~n9596 & n9597 ;
  assign n9599 = ~n8949 & n9598 ;
  assign n9600 = ~n9595 & ~n9599 ;
  assign n9601 = ~n9591 & ~n9600 ;
  assign n9602 = \sa30_reg[0]/P0002  & ~n9601 ;
  assign n9542 = n8692 & ~n8725 ;
  assign n9543 = ~\sa30_reg[4]/P0001  & n8813 ;
  assign n9544 = ~n9542 & ~n9543 ;
  assign n9545 = ~\sa30_reg[2]/P0001  & ~n9544 ;
  assign n9547 = \sa30_reg[4]/P0001  & n8874 ;
  assign n9548 = n8929 & n9547 ;
  assign n9546 = \sa30_reg[2]/P0001  & n8705 ;
  assign n9549 = ~n8889 & ~n9546 ;
  assign n9550 = ~n9548 & n9549 ;
  assign n9551 = ~n9545 & n9550 ;
  assign n9552 = \sa30_reg[1]/P0001  & ~n9551 ;
  assign n9554 = ~\sa30_reg[7]/P0001  & n8833 ;
  assign n9555 = ~n8811 & ~n9554 ;
  assign n9556 = n8697 & ~n9555 ;
  assign n9553 = \sa30_reg[2]/P0001  & n8950 ;
  assign n9557 = ~n8953 & ~n9553 ;
  assign n9558 = ~n9556 & n9557 ;
  assign n9559 = ~\sa30_reg[1]/P0001  & ~n9558 ;
  assign n9560 = ~\sa30_reg[6]/NET0131  & n8695 ;
  assign n9561 = n8734 & n9560 ;
  assign n9562 = n8698 & n8792 ;
  assign n9563 = ~n9561 & ~n9562 ;
  assign n9564 = \sa30_reg[2]/P0001  & ~n9563 ;
  assign n9541 = ~\sa30_reg[3]/P0001  & n8765 ;
  assign n9565 = n8684 & n8698 ;
  assign n9566 = ~\sa30_reg[7]/P0001  & n9565 ;
  assign n9567 = ~n9541 & ~n9566 ;
  assign n9568 = ~n9564 & n9567 ;
  assign n9569 = ~n9559 & n9568 ;
  assign n9570 = ~n9552 & n9569 ;
  assign n9571 = ~\sa30_reg[0]/P0002  & ~n9570 ;
  assign n9605 = ~n8720 & ~n8909 ;
  assign n9606 = ~n8949 & n9605 ;
  assign n9607 = ~\sa30_reg[2]/P0001  & ~n9606 ;
  assign n9609 = \sa30_reg[1]/P0001  & ~n8836 ;
  assign n9608 = ~\sa30_reg[6]/NET0131  & n8922 ;
  assign n9603 = n8695 & n8709 ;
  assign n9604 = ~\sa30_reg[5]/P0001  & n9603 ;
  assign n9610 = ~n8846 & ~n9604 ;
  assign n9611 = ~n9608 & n9610 ;
  assign n9612 = n9609 & n9611 ;
  assign n9613 = ~n9607 & n9612 ;
  assign n9614 = \sa30_reg[4]/P0001  & n8792 ;
  assign n9615 = ~n8710 & ~n9614 ;
  assign n9616 = ~\sa30_reg[3]/P0001  & ~n9615 ;
  assign n9617 = n8709 & n8773 ;
  assign n9618 = ~\sa30_reg[2]/P0001  & ~n9617 ;
  assign n9619 = ~n9616 & n9618 ;
  assign n9620 = n8684 & n8725 ;
  assign n9623 = \sa30_reg[2]/P0001  & ~n8759 ;
  assign n9624 = ~n9620 & n9623 ;
  assign n9621 = ~n8721 & ~n8725 ;
  assign n9622 = n8813 & n9621 ;
  assign n9625 = ~n8894 & ~n9622 ;
  assign n9626 = n9624 & n9625 ;
  assign n9627 = ~n9619 & ~n9626 ;
  assign n9628 = ~\sa30_reg[1]/P0001  & ~n8822 ;
  assign n9629 = ~n9566 & n9628 ;
  assign n9630 = ~n9627 & n9629 ;
  assign n9631 = ~n9613 & ~n9630 ;
  assign n9634 = \sa30_reg[2]/P0001  & ~n8821 ;
  assign n9632 = n8734 & n8758 ;
  assign n9633 = ~\sa30_reg[2]/P0001  & ~n9632 ;
  assign n9635 = ~n8741 & ~n9633 ;
  assign n9636 = ~n9634 & n9635 ;
  assign n9637 = ~n9631 & ~n9636 ;
  assign n9638 = ~n9571 & n9637 ;
  assign n9639 = ~n9602 & n9638 ;
  assign n9640 = \u0_w_reg[1][13]/P0001  & ~n9639 ;
  assign n9641 = ~\u0_w_reg[1][13]/P0001  & n9639 ;
  assign n9642 = ~n9640 & ~n9641 ;
  assign n9643 = n8853 & n9642 ;
  assign n9644 = ~n8853 & ~n9642 ;
  assign n9645 = ~n9643 & ~n9644 ;
  assign n9647 = n9540 & ~n9645 ;
  assign n9646 = ~n9540 & n9645 ;
  assign n9648 = ~\ld_r_reg/P0001  & ~n9646 ;
  assign n9649 = ~n9647 & n9648 ;
  assign n9651 = \text_in_r_reg[77]/P0001  & \u0_w_reg[1][13]/P0001  ;
  assign n9650 = ~\text_in_r_reg[77]/P0001  & ~\u0_w_reg[1][13]/P0001  ;
  assign n9652 = \ld_r_reg/P0001  & ~n9650 ;
  assign n9653 = ~n9651 & n9652 ;
  assign n9654 = ~n9649 & ~n9653 ;
  assign n9655 = n9063 & ~n9400 ;
  assign n9656 = ~n9063 & n9400 ;
  assign n9657 = ~n9655 & ~n9656 ;
  assign n9658 = ~n8678 & ~n9657 ;
  assign n9659 = n8678 & n9657 ;
  assign n9660 = ~n9658 & ~n9659 ;
  assign n9661 = \u0_w_reg[1][14]/P0001  & ~n8974 ;
  assign n9662 = ~\u0_w_reg[1][14]/P0001  & n8974 ;
  assign n9663 = ~n9661 & ~n9662 ;
  assign n9664 = n8853 & n9663 ;
  assign n9665 = ~n8853 & ~n9663 ;
  assign n9666 = ~n9664 & ~n9665 ;
  assign n9668 = n9660 & n9666 ;
  assign n9667 = ~n9660 & ~n9666 ;
  assign n9669 = ~\ld_r_reg/P0001  & ~n9667 ;
  assign n9670 = ~n9668 & n9669 ;
  assign n9672 = ~\text_in_r_reg[78]/P0001  & \u0_w_reg[1][14]/P0001  ;
  assign n9671 = \text_in_r_reg[78]/P0001  & ~\u0_w_reg[1][14]/P0001  ;
  assign n9673 = \ld_r_reg/P0001  & ~n9671 ;
  assign n9674 = ~n9672 & n9673 ;
  assign n9675 = ~n9670 & ~n9674 ;
  assign n9676 = ~n9289 & ~n9657 ;
  assign n9677 = n9289 & n9657 ;
  assign n9678 = ~n9676 & ~n9677 ;
  assign n9679 = \u0_w_reg[1][6]/P0001  & ~n9169 ;
  assign n9680 = ~\u0_w_reg[1][6]/P0001  & n9169 ;
  assign n9681 = ~n9679 & ~n9680 ;
  assign n9682 = n8853 & n9681 ;
  assign n9683 = ~n8853 & ~n9681 ;
  assign n9684 = ~n9682 & ~n9683 ;
  assign n9686 = n9678 & ~n9684 ;
  assign n9685 = ~n9678 & n9684 ;
  assign n9687 = ~\ld_r_reg/P0001  & ~n9685 ;
  assign n9688 = ~n9686 & n9687 ;
  assign n9690 = \text_in_r_reg[70]/P0001  & \u0_w_reg[1][6]/P0001  ;
  assign n9689 = ~\text_in_r_reg[70]/P0001  & ~\u0_w_reg[1][6]/P0001  ;
  assign n9691 = \ld_r_reg/P0001  & ~n9689 ;
  assign n9692 = ~n9690 & n9691 ;
  assign n9693 = ~n9688 & ~n9692 ;
  assign n9728 = ~n8369 & ~n9373 ;
  assign n9729 = n8242 & ~n8281 ;
  assign n9730 = n9728 & ~n9729 ;
  assign n9731 = n9386 & ~n9730 ;
  assign n9701 = ~n8225 & ~n9352 ;
  assign n9732 = \sa01_reg[7]/NET0131  & ~n9701 ;
  assign n9733 = ~n8309 & ~n9732 ;
  assign n9734 = ~\sa01_reg[3]/P0001  & ~n9733 ;
  assign n9735 = ~n8343 & ~n9212 ;
  assign n9736 = ~n9734 & n9735 ;
  assign n9737 = \sa01_reg[2]/P0001  & ~n9736 ;
  assign n9738 = ~n9731 & ~n9737 ;
  assign n9739 = \sa01_reg[1]/P0001  & ~n9738 ;
  assign n9714 = ~n8295 & ~n9175 ;
  assign n9715 = ~n9352 & n9714 ;
  assign n9716 = ~\sa01_reg[2]/P0001  & ~n9715 ;
  assign n9710 = n8281 & n8351 ;
  assign n9711 = \sa01_reg[2]/P0001  & ~n9710 ;
  assign n9712 = ~n9244 & ~n9711 ;
  assign n9713 = ~n8222 & n8326 ;
  assign n9717 = ~n8341 & ~n9713 ;
  assign n9718 = ~n9712 & n9717 ;
  assign n9719 = ~n9716 & n9718 ;
  assign n9720 = ~\sa01_reg[1]/P0001  & ~n9719 ;
  assign n9706 = \sa01_reg[7]/NET0131  & n8304 ;
  assign n9707 = ~n9176 & ~n9185 ;
  assign n9708 = ~n9706 & n9707 ;
  assign n9709 = \sa01_reg[2]/P0001  & ~n9708 ;
  assign n9702 = ~\sa01_reg[7]/NET0131  & n8264 ;
  assign n9703 = ~n8339 & ~n9702 ;
  assign n9704 = n9701 & n9703 ;
  assign n9705 = n9388 & ~n9704 ;
  assign n9694 = ~\sa01_reg[2]/P0001  & ~\sa01_reg[3]/P0001  ;
  assign n9695 = n8344 & n9694 ;
  assign n9696 = ~n8332 & ~n9695 ;
  assign n9697 = \sa01_reg[1]/P0001  & ~n9696 ;
  assign n9700 = n8326 & n9209 ;
  assign n9698 = \sa01_reg[2]/P0001  & n8218 ;
  assign n9699 = n8310 & n9698 ;
  assign n9721 = ~n9356 & ~n9699 ;
  assign n9722 = ~n9700 & n9721 ;
  assign n9723 = ~n9697 & n9722 ;
  assign n9724 = ~n9705 & n9723 ;
  assign n9725 = ~n9709 & n9724 ;
  assign n9726 = ~n9720 & n9725 ;
  assign n9727 = \sa01_reg[0]/P0001  & ~n9726 ;
  assign n9741 = n8276 & n8318 ;
  assign n9742 = ~n8239 & ~n9741 ;
  assign n9743 = ~\sa01_reg[2]/P0001  & ~n9742 ;
  assign n9740 = ~n8240 & n8356 ;
  assign n9744 = \sa01_reg[1]/P0001  & ~n9369 ;
  assign n9745 = ~n9740 & n9744 ;
  assign n9746 = ~n9743 & n9745 ;
  assign n9747 = ~n8215 & ~n9319 ;
  assign n9748 = n8303 & ~n9747 ;
  assign n9749 = ~\sa01_reg[2]/P0001  & n8281 ;
  assign n9750 = ~\sa01_reg[1]/P0001  & ~n9315 ;
  assign n9751 = ~n9749 & n9750 ;
  assign n9752 = ~n9748 & n9751 ;
  assign n9753 = ~n9746 & ~n9752 ;
  assign n9758 = ~n8361 & ~n9389 ;
  assign n9759 = ~\sa01_reg[2]/P0001  & ~n9758 ;
  assign n9754 = n8224 & n8257 ;
  assign n9755 = ~n9276 & ~n9754 ;
  assign n9756 = n8329 & ~n9755 ;
  assign n9757 = n8329 & n9219 ;
  assign n9760 = ~n8258 & ~n9231 ;
  assign n9761 = n9694 & ~n9760 ;
  assign n9762 = ~n9757 & ~n9761 ;
  assign n9763 = ~n9756 & n9762 ;
  assign n9764 = ~n9759 & n9763 ;
  assign n9765 = ~n9753 & n9764 ;
  assign n9766 = ~\sa01_reg[0]/P0001  & ~n9765 ;
  assign n9767 = ~\sa01_reg[5]/P0001  & n8305 ;
  assign n9768 = ~n9181 & ~n9767 ;
  assign n9769 = ~\sa01_reg[2]/P0001  & ~n9768 ;
  assign n9770 = ~\sa01_reg[3]/P0001  & n8295 ;
  assign n9771 = ~n8332 & ~n9179 ;
  assign n9772 = ~n9770 & n9771 ;
  assign n9773 = \sa01_reg[2]/P0001  & ~n9772 ;
  assign n9774 = n8214 & n8245 ;
  assign n9775 = n8282 & n9386 ;
  assign n9776 = ~n9774 & ~n9775 ;
  assign n9777 = ~n9761 & n9776 ;
  assign n9778 = ~n9773 & n9777 ;
  assign n9779 = ~\sa01_reg[1]/P0001  & ~n9778 ;
  assign n9780 = ~n9769 & ~n9779 ;
  assign n9781 = ~n9766 & n9780 ;
  assign n9782 = ~n9727 & n9781 ;
  assign n9783 = ~n9739 & n9782 ;
  assign n9788 = ~n8068 & ~n9025 ;
  assign n9816 = \sa12_reg[3]/P0001  & n8060 ;
  assign n9817 = ~\sa12_reg[3]/P0001  & n8055 ;
  assign n9818 = ~n9816 & ~n9817 ;
  assign n9819 = n9788 & n9818 ;
  assign n9820 = \sa12_reg[2]/P0001  & ~n9819 ;
  assign n9821 = n8135 & n8978 ;
  assign n9822 = ~\sa12_reg[6]/NET0131  & n9821 ;
  assign n9823 = ~n8109 & ~n9822 ;
  assign n9824 = ~n9820 & n9823 ;
  assign n9825 = \sa12_reg[1]/P0001  & ~n9824 ;
  assign n9798 = ~n8135 & n8390 ;
  assign n9799 = ~n9025 & ~n9798 ;
  assign n9800 = ~\sa12_reg[2]/P0001  & ~n9799 ;
  assign n9803 = \sa12_reg[2]/P0001  & ~n8094 ;
  assign n9804 = n8060 & ~n8110 ;
  assign n9805 = ~n9803 & n9804 ;
  assign n9801 = n8104 & n8135 ;
  assign n9802 = \sa12_reg[2]/P0001  & n9801 ;
  assign n9806 = ~n8079 & ~n9802 ;
  assign n9807 = ~n9805 & n9806 ;
  assign n9808 = ~n9800 & n9807 ;
  assign n9809 = ~\sa12_reg[1]/P0001  & ~n9808 ;
  assign n9811 = ~n8084 & ~n8110 ;
  assign n9812 = n8068 & ~n9811 ;
  assign n9813 = ~n8380 & ~n8391 ;
  assign n9814 = ~n9812 & n9813 ;
  assign n9815 = \sa12_reg[2]/P0001  & ~n9814 ;
  assign n9810 = n8061 & n8978 ;
  assign n9826 = ~n8494 & ~n9810 ;
  assign n9827 = ~n9815 & n9826 ;
  assign n9828 = ~n9809 & n9827 ;
  assign n9829 = ~n9825 & n9828 ;
  assign n9830 = \sa12_reg[0]/P0001  & ~n9829 ;
  assign n9784 = ~n8070 & ~n9044 ;
  assign n9785 = n8077 & ~n8111 ;
  assign n9786 = n9784 & ~n9785 ;
  assign n9787 = n8155 & ~n9786 ;
  assign n9789 = \sa12_reg[7]/NET0131  & ~n9788 ;
  assign n9790 = n8077 & n8498 ;
  assign n9791 = ~n9789 & ~n9790 ;
  assign n9792 = ~\sa12_reg[3]/P0001  & ~n9791 ;
  assign n9793 = ~n8076 & ~n8422 ;
  assign n9794 = ~n9792 & n9793 ;
  assign n9795 = \sa12_reg[2]/P0001  & ~n9794 ;
  assign n9796 = ~n9787 & ~n9795 ;
  assign n9797 = \sa12_reg[1]/P0001  & ~n9796 ;
  assign n9833 = ~n8103 & ~n9034 ;
  assign n9834 = ~\sa12_reg[2]/P0001  & ~n9833 ;
  assign n9831 = ~n8432 & ~n8490 ;
  assign n9832 = n8057 & ~n9831 ;
  assign n9835 = ~n8130 & ~n8443 ;
  assign n9836 = n8978 & ~n9835 ;
  assign n9837 = n8055 & n8144 ;
  assign n9838 = n8110 & n9837 ;
  assign n9852 = ~n9836 & ~n9838 ;
  assign n9853 = ~n9832 & n9852 ;
  assign n9854 = ~n9834 & n9853 ;
  assign n9839 = ~n8459 & ~n9042 ;
  assign n9840 = ~\sa12_reg[2]/P0001  & ~n9839 ;
  assign n9841 = ~\sa12_reg[2]/P0001  & ~\sa12_reg[7]/NET0131  ;
  assign n9842 = n8095 & ~n9841 ;
  assign n9843 = ~n9035 & ~n9842 ;
  assign n9844 = ~n9840 & n9843 ;
  assign n9845 = \sa12_reg[1]/P0001  & ~n9844 ;
  assign n9847 = n8135 & n8479 ;
  assign n9846 = ~\sa12_reg[2]/P0001  & n8111 ;
  assign n9848 = ~n8985 & ~n9846 ;
  assign n9849 = ~n8194 & n9848 ;
  assign n9850 = ~n9847 & n9849 ;
  assign n9851 = ~\sa12_reg[1]/P0001  & ~n9850 ;
  assign n9855 = ~n9845 & ~n9851 ;
  assign n9856 = n9854 & n9855 ;
  assign n9857 = ~\sa12_reg[0]/P0001  & ~n9856 ;
  assign n9858 = ~n8201 & ~n8395 ;
  assign n9859 = ~\sa12_reg[2]/P0001  & ~n9858 ;
  assign n9860 = \sa12_reg[4]/P0001  & n8065 ;
  assign n9861 = ~\sa12_reg[3]/P0001  & n9860 ;
  assign n9862 = ~n8109 & ~n8387 ;
  assign n9863 = ~n9861 & n9862 ;
  assign n9864 = \sa12_reg[2]/P0001  & ~n9863 ;
  assign n9865 = n8094 & n8161 ;
  assign n9866 = n8110 & n9846 ;
  assign n9867 = ~n9865 & ~n9866 ;
  assign n9868 = ~n9836 & n9867 ;
  assign n9869 = ~n9864 & n9868 ;
  assign n9870 = ~\sa12_reg[1]/P0001  & ~n9869 ;
  assign n9871 = ~n9859 & ~n9870 ;
  assign n9872 = ~n9857 & n9871 ;
  assign n9873 = ~n9797 & n9872 ;
  assign n9874 = ~n9830 & n9873 ;
  assign n9875 = ~n9783 & ~n9874 ;
  assign n9876 = n9783 & n9874 ;
  assign n9877 = ~n9875 & ~n9876 ;
  assign n9878 = ~n9400 & ~n9877 ;
  assign n9879 = n9400 & n9877 ;
  assign n9880 = ~n9878 & ~n9879 ;
  assign n9905 = ~n8519 & n8521 ;
  assign n9906 = ~n9073 & ~n9099 ;
  assign n9907 = ~n9905 & n9906 ;
  assign n9908 = ~\sa23_reg[2]/P0001  & ~n9907 ;
  assign n9900 = \sa23_reg[2]/P0001  & ~\sa23_reg[4]/P0001  ;
  assign n9901 = n8513 & ~n9900 ;
  assign n9902 = \sa23_reg[2]/P0001  & n9453 ;
  assign n9903 = ~n9901 & ~n9902 ;
  assign n9904 = ~\sa23_reg[3]/P0001  & ~n9903 ;
  assign n9909 = ~n9466 & ~n9904 ;
  assign n9910 = ~n9908 & n9909 ;
  assign n9911 = ~\sa23_reg[1]/P0001  & ~n9910 ;
  assign n9882 = ~n8552 & ~n8556 ;
  assign n9881 = \sa23_reg[3]/P0001  & n8513 ;
  assign n9883 = ~n9099 & ~n9881 ;
  assign n9884 = n9882 & n9883 ;
  assign n9885 = \sa23_reg[1]/P0001  & ~n9884 ;
  assign n9886 = \sa23_reg[7]/NET0131  & n8556 ;
  assign n9887 = ~\sa23_reg[3]/P0001  & n9886 ;
  assign n9888 = ~n8510 & ~n8534 ;
  assign n9889 = ~n9887 & n9888 ;
  assign n9890 = ~n9885 & n9889 ;
  assign n9891 = \sa23_reg[2]/P0001  & ~n9890 ;
  assign n9893 = ~\sa23_reg[5]/P0001  & n8550 ;
  assign n9894 = ~\sa23_reg[2]/P0001  & n9893 ;
  assign n9895 = ~n9455 & ~n9894 ;
  assign n9896 = \sa23_reg[1]/P0001  & ~n9895 ;
  assign n9899 = \sa23_reg[5]/P0001  & n8635 ;
  assign n9892 = n9073 & n9079 ;
  assign n9897 = \sa23_reg[2]/P0001  & n8572 ;
  assign n9898 = n8525 & n9897 ;
  assign n9912 = ~n9892 & ~n9898 ;
  assign n9913 = ~n9899 & n9912 ;
  assign n9914 = ~n9896 & n9913 ;
  assign n9915 = ~n9891 & n9914 ;
  assign n9916 = ~n9911 & n9915 ;
  assign n9917 = \sa23_reg[0]/P0001  & ~n9916 ;
  assign n9920 = \sa23_reg[4]/P0001  & n8562 ;
  assign n9921 = n8546 & n9920 ;
  assign n9923 = ~\sa23_reg[1]/P0001  & ~n9078 ;
  assign n9918 = n8564 & n8660 ;
  assign n9922 = \sa23_reg[7]/NET0131  & n9427 ;
  assign n9924 = ~n9918 & ~n9922 ;
  assign n9925 = n9923 & n9924 ;
  assign n9926 = ~n9921 & n9925 ;
  assign n9927 = n8513 & n8529 ;
  assign n9928 = ~\sa23_reg[6]/NET0131  & n8537 ;
  assign n9929 = ~n9927 & ~n9928 ;
  assign n9930 = ~\sa23_reg[2]/P0001  & ~n9929 ;
  assign n9931 = \sa23_reg[2]/P0001  & \sa23_reg[4]/P0001  ;
  assign n9932 = ~n8569 & ~n9931 ;
  assign n9933 = n8642 & ~n9932 ;
  assign n9934 = \sa23_reg[1]/P0001  & ~n9154 ;
  assign n9935 = ~n9933 & n9934 ;
  assign n9936 = ~n9930 & n9935 ;
  assign n9937 = ~n9926 & ~n9936 ;
  assign n9919 = n8572 & n9918 ;
  assign n9938 = n8521 & n8569 ;
  assign n9939 = ~n8667 & ~n9938 ;
  assign n9940 = \sa23_reg[3]/P0001  & ~n9939 ;
  assign n9941 = \sa23_reg[2]/P0001  & ~n9940 ;
  assign n9942 = n8521 & n8526 ;
  assign n9943 = n8522 & n8589 ;
  assign n9944 = ~n9942 & ~n9943 ;
  assign n9945 = ~n9125 & n9944 ;
  assign n9946 = n9474 & n9945 ;
  assign n9947 = ~n9941 & ~n9946 ;
  assign n9948 = ~n9919 & ~n9947 ;
  assign n9949 = ~n9937 & n9948 ;
  assign n9950 = ~\sa23_reg[0]/P0001  & ~n9949 ;
  assign n9969 = ~n9420 & ~n9482 ;
  assign n9970 = ~n9886 & n9969 ;
  assign n9971 = ~\sa23_reg[3]/P0001  & ~n9970 ;
  assign n9972 = ~n8563 & n9465 ;
  assign n9973 = ~n9971 & n9972 ;
  assign n9963 = n8508 & ~n8519 ;
  assign n9964 = n8525 & n8577 ;
  assign n9965 = ~n8557 & ~n9964 ;
  assign n9966 = ~n9963 & n9965 ;
  assign n9967 = \sa23_reg[3]/P0001  & ~n9966 ;
  assign n9968 = ~\sa23_reg[2]/P0001  & ~n9967 ;
  assign n9974 = \sa23_reg[1]/P0001  & ~n9968 ;
  assign n9975 = ~n9973 & n9974 ;
  assign n9958 = ~\sa23_reg[1]/P0001  & \sa23_reg[2]/P0001  ;
  assign n9959 = \sa23_reg[5]/P0001  & n8574 ;
  assign n9960 = ~n8530 & ~n9455 ;
  assign n9961 = ~n9959 & n9960 ;
  assign n9962 = n9958 & ~n9961 ;
  assign n9951 = ~n8524 & ~n9485 ;
  assign n9952 = ~\sa23_reg[2]/P0001  & ~n9951 ;
  assign n9953 = \sa23_reg[2]/P0001  & ~n8619 ;
  assign n9954 = ~\sa23_reg[1]/P0001  & ~n9953 ;
  assign n9955 = ~n8619 & ~n9139 ;
  assign n9956 = n9944 & n9955 ;
  assign n9957 = n9954 & ~n9956 ;
  assign n9976 = ~n9952 & ~n9957 ;
  assign n9977 = ~n9962 & n9976 ;
  assign n9978 = ~n9975 & n9977 ;
  assign n9979 = ~n9950 & n9978 ;
  assign n9980 = ~n9917 & n9979 ;
  assign n9981 = \u0_w_reg[1][7]/P0001  & ~n9980 ;
  assign n9982 = ~\u0_w_reg[1][7]/P0001  & n9980 ;
  assign n9983 = ~n9981 & ~n9982 ;
  assign n9984 = n8974 & n9983 ;
  assign n9985 = ~n8974 & ~n9983 ;
  assign n9986 = ~n9984 & ~n9985 ;
  assign n9988 = n9880 & ~n9986 ;
  assign n9987 = ~n9880 & n9986 ;
  assign n9989 = ~\ld_r_reg/P0001  & ~n9987 ;
  assign n9990 = ~n9988 & n9989 ;
  assign n9992 = ~\text_in_r_reg[71]/P0001  & \u0_w_reg[1][7]/P0001  ;
  assign n9991 = \text_in_r_reg[71]/P0001  & ~\u0_w_reg[1][7]/P0001  ;
  assign n9993 = \ld_r_reg/P0001  & ~n9991 ;
  assign n9994 = ~n9992 & n9993 ;
  assign n9995 = ~n9990 & ~n9994 ;
  assign n10025 = ~n8136 & ~n8175 ;
  assign n10026 = \sa12_reg[2]/P0001  & ~n10025 ;
  assign n10022 = ~n8981 & ~n9049 ;
  assign n10023 = ~\sa12_reg[2]/P0001  & ~n10022 ;
  assign n10024 = \sa12_reg[4]/P0001  & n9042 ;
  assign n10027 = ~n8098 & ~n10024 ;
  assign n10028 = ~n10023 & n10027 ;
  assign n10029 = ~n10026 & n10028 ;
  assign n10030 = ~\sa12_reg[1]/P0001  & ~n10029 ;
  assign n10031 = \sa12_reg[4]/P0001  & ~n8075 ;
  assign n10032 = n8979 & ~n10031 ;
  assign n10033 = ~n8404 & ~n10032 ;
  assign n10034 = ~\sa12_reg[2]/P0001  & ~n10033 ;
  assign n10035 = ~n8114 & ~n8165 ;
  assign n10036 = \sa12_reg[2]/P0001  & ~n10035 ;
  assign n10037 = ~n8387 & n8444 ;
  assign n10038 = ~n10036 & n10037 ;
  assign n10039 = ~n10034 & n10038 ;
  assign n10040 = \sa12_reg[1]/P0001  & ~n10039 ;
  assign n10043 = ~n8098 & ~n8461 ;
  assign n10044 = ~\sa12_reg[2]/P0001  & ~n10043 ;
  assign n10041 = ~n8142 & ~n8498 ;
  assign n10042 = n8059 & ~n10041 ;
  assign n10045 = ~n8485 & ~n8491 ;
  assign n10046 = ~n10042 & n10045 ;
  assign n10047 = ~n10044 & n10046 ;
  assign n10048 = ~n10040 & n10047 ;
  assign n10049 = ~n10030 & n10048 ;
  assign n10050 = ~\sa12_reg[0]/P0001  & ~n10049 ;
  assign n9996 = n8075 & n8165 ;
  assign n9997 = ~n8422 & ~n9996 ;
  assign n9998 = ~n8111 & ~n8390 ;
  assign n9999 = ~\sa12_reg[5]/P0001  & ~n9998 ;
  assign n10000 = ~n8159 & ~n9999 ;
  assign n10001 = \sa12_reg[2]/P0001  & ~n10000 ;
  assign n10002 = n9997 & ~n10001 ;
  assign n10003 = \sa12_reg[1]/P0001  & ~n10002 ;
  assign n10013 = ~n8070 & ~n8175 ;
  assign n10014 = ~n8490 & ~n9035 ;
  assign n10015 = n10013 & n10014 ;
  assign n10016 = ~\sa12_reg[2]/P0001  & ~n10015 ;
  assign n10004 = \sa12_reg[5]/P0001  & n9015 ;
  assign n10006 = ~n8144 & n8381 ;
  assign n10005 = n8074 & n8180 ;
  assign n10007 = ~n8070 & ~n10005 ;
  assign n10008 = ~n10006 & n10007 ;
  assign n10009 = ~n10004 & n10008 ;
  assign n10010 = ~\sa12_reg[1]/P0001  & ~n10009 ;
  assign n10011 = n8096 & ~n8162 ;
  assign n10012 = \sa12_reg[4]/P0001  & n8087 ;
  assign n10017 = ~n10011 & ~n10012 ;
  assign n10018 = ~n10010 & n10017 ;
  assign n10019 = ~n10016 & n10018 ;
  assign n10020 = ~n10003 & n10019 ;
  assign n10021 = \sa12_reg[0]/P0001  & ~n10020 ;
  assign n10069 = ~n8985 & ~n9042 ;
  assign n10070 = ~n8143 & n10069 ;
  assign n10071 = ~\sa12_reg[2]/P0001  & ~n10070 ;
  assign n10072 = ~n8083 & ~n8460 ;
  assign n10073 = ~n10071 & n10072 ;
  assign n10074 = ~\sa12_reg[1]/P0001  & ~n10073 ;
  assign n10055 = ~\sa12_reg[3]/P0001  & n8077 ;
  assign n10056 = ~n8425 & ~n10055 ;
  assign n10057 = ~n8080 & ~n10056 ;
  assign n10058 = ~n8990 & ~n10057 ;
  assign n10059 = n8455 & ~n10058 ;
  assign n10051 = ~n8422 & ~n9860 ;
  assign n10052 = \sa12_reg[3]/P0001  & ~n10051 ;
  assign n10053 = ~n8177 & ~n10052 ;
  assign n10054 = n9033 & ~n10053 ;
  assign n10065 = ~n8417 & ~n8432 ;
  assign n10066 = ~n8481 & n10065 ;
  assign n10064 = ~\sa12_reg[1]/P0001  & \sa12_reg[2]/P0001  ;
  assign n10067 = ~\sa12_reg[3]/P0001  & n10064 ;
  assign n10068 = ~n10066 & n10067 ;
  assign n10060 = ~\sa12_reg[1]/P0001  & ~\sa12_reg[2]/P0001  ;
  assign n10061 = ~n8066 & ~n10060 ;
  assign n10062 = n8387 & n10061 ;
  assign n10063 = \sa12_reg[2]/P0001  & n8083 ;
  assign n10075 = ~n10062 & ~n10063 ;
  assign n10076 = ~n10068 & n10075 ;
  assign n10077 = ~n10054 & n10076 ;
  assign n10078 = ~n10059 & n10077 ;
  assign n10079 = ~n10074 & n10078 ;
  assign n10080 = ~n10021 & n10079 ;
  assign n10081 = ~n10050 & n10080 ;
  assign n10086 = \sa01_reg[4]/P0001  & n8310 ;
  assign n10109 = \sa01_reg[3]/P0001  & n10086 ;
  assign n10108 = ~\sa01_reg[3]/P0001  & n8221 ;
  assign n10110 = ~n9201 & ~n10108 ;
  assign n10111 = ~n10109 & n10110 ;
  assign n10112 = ~\sa01_reg[2]/P0001  & ~n10111 ;
  assign n10113 = \sa01_reg[1]/P0001  & ~n9179 ;
  assign n10114 = n9232 & n10113 ;
  assign n10115 = ~n10112 & n10114 ;
  assign n10117 = ~n9324 & ~n9368 ;
  assign n10118 = ~\sa01_reg[2]/P0001  & ~n10117 ;
  assign n10116 = n8238 & n9206 ;
  assign n10119 = ~\sa01_reg[1]/P0001  & ~n8355 ;
  assign n10120 = ~n10116 & n10119 ;
  assign n10121 = ~n10118 & n10120 ;
  assign n10122 = ~n10115 & ~n10121 ;
  assign n10130 = ~n8216 & ~n8265 ;
  assign n10131 = n9197 & ~n10130 ;
  assign n10132 = ~n8362 & ~n9277 ;
  assign n10133 = ~n10131 & n10132 ;
  assign n10128 = ~n8269 & ~n8293 ;
  assign n10129 = n9318 & ~n10128 ;
  assign n10123 = ~\sa01_reg[3]/P0001  & n8258 ;
  assign n10124 = ~n9215 & ~n10123 ;
  assign n10125 = n9388 & ~n10124 ;
  assign n10126 = ~n8355 & ~n9237 ;
  assign n10127 = ~\sa01_reg[2]/P0001  & ~n10126 ;
  assign n10134 = ~n10125 & ~n10127 ;
  assign n10135 = ~n10129 & n10134 ;
  assign n10136 = n10133 & n10135 ;
  assign n10137 = ~n10122 & n10136 ;
  assign n10138 = ~\sa01_reg[0]/P0001  & ~n10137 ;
  assign n10083 = n8238 & n8258 ;
  assign n10084 = ~n9212 & ~n10083 ;
  assign n10085 = \sa01_reg[3]/P0001  & n8235 ;
  assign n10087 = ~n8282 & ~n10085 ;
  assign n10088 = ~n10086 & n10087 ;
  assign n10089 = \sa01_reg[2]/P0001  & ~n10088 ;
  assign n10090 = n10084 & ~n10089 ;
  assign n10091 = \sa01_reg[1]/P0001  & ~n10090 ;
  assign n10099 = ~\sa01_reg[6]/NET0131  & n8321 ;
  assign n10098 = ~n8222 & n9183 ;
  assign n10100 = ~n8360 & ~n8369 ;
  assign n10101 = ~n10098 & n10100 ;
  assign n10102 = ~n10099 & n10101 ;
  assign n10103 = ~\sa01_reg[1]/P0001  & ~n10102 ;
  assign n10082 = ~n8246 & n8352 ;
  assign n10092 = ~\sa01_reg[3]/P0001  & n9276 ;
  assign n10093 = \sa01_reg[2]/P0001  & ~n10092 ;
  assign n10094 = ~n8293 & ~n8369 ;
  assign n10095 = ~n9276 & ~n9369 ;
  assign n10096 = n10094 & n10095 ;
  assign n10097 = ~n10093 & ~n10096 ;
  assign n10104 = ~n10082 & ~n10097 ;
  assign n10105 = ~n10103 & n10104 ;
  assign n10106 = ~n10091 & n10105 ;
  assign n10107 = \sa01_reg[0]/P0001  & ~n10106 ;
  assign n10153 = n8221 & n8351 ;
  assign n10154 = ~n8362 & ~n10153 ;
  assign n10155 = ~n9243 & n10154 ;
  assign n10156 = \sa01_reg[2]/P0001  & ~n10155 ;
  assign n10157 = n8239 & n8254 ;
  assign n10158 = ~n9236 & ~n10157 ;
  assign n10159 = ~n10156 & n10158 ;
  assign n10160 = ~\sa01_reg[1]/P0001  & ~n10159 ;
  assign n10149 = ~n8295 & ~n9212 ;
  assign n10150 = \sa01_reg[3]/P0001  & ~n10149 ;
  assign n10151 = ~n9338 & ~n10150 ;
  assign n10152 = n9388 & ~n10151 ;
  assign n10139 = ~n9184 & ~n9219 ;
  assign n10140 = ~n8224 & ~n10139 ;
  assign n10141 = ~n9179 & ~n9309 ;
  assign n10142 = ~n10140 & n10141 ;
  assign n10143 = n9382 & ~n10142 ;
  assign n10145 = ~\sa01_reg[1]/P0001  & ~\sa01_reg[2]/P0001  ;
  assign n10146 = ~n9315 & ~n9741 ;
  assign n10147 = ~n8217 & n10146 ;
  assign n10148 = n10145 & ~n10147 ;
  assign n10144 = n8303 & n9375 ;
  assign n10161 = ~n9757 & ~n10144 ;
  assign n10162 = ~n10148 & n10161 ;
  assign n10163 = ~n10143 & n10162 ;
  assign n10164 = ~n10152 & n10163 ;
  assign n10165 = ~n10160 & n10164 ;
  assign n10166 = ~n10107 & n10165 ;
  assign n10167 = ~n10138 & n10166 ;
  assign n10168 = ~n10081 & ~n10167 ;
  assign n10169 = n10081 & n10167 ;
  assign n10170 = ~n10168 & ~n10169 ;
  assign n10186 = n8215 & n8351 ;
  assign n10187 = ~n9176 & ~n10186 ;
  assign n10188 = ~n9268 & n10187 ;
  assign n10189 = \sa01_reg[2]/P0001  & ~n10188 ;
  assign n10183 = \sa01_reg[5]/P0001  & ~n8221 ;
  assign n10184 = n8218 & ~n10183 ;
  assign n10182 = n9209 & n10153 ;
  assign n10185 = n8267 & n8342 ;
  assign n10190 = ~n10182 & ~n10185 ;
  assign n10191 = ~n10184 & n10190 ;
  assign n10192 = ~n10189 & n10191 ;
  assign n10193 = ~\sa01_reg[1]/P0001  & ~n10192 ;
  assign n10179 = ~n8283 & ~n9237 ;
  assign n10180 = n9316 & n10179 ;
  assign n10181 = \sa01_reg[2]/P0001  & ~n10180 ;
  assign n10171 = ~n8216 & ~n8257 ;
  assign n10172 = ~\sa01_reg[2]/P0001  & ~n10171 ;
  assign n10173 = ~n9368 & ~n10172 ;
  assign n10174 = \sa01_reg[1]/P0001  & ~n10173 ;
  assign n10177 = ~n9356 & ~n9754 ;
  assign n10178 = ~\sa01_reg[2]/P0001  & ~n10177 ;
  assign n10175 = ~n8265 & ~n8310 ;
  assign n10176 = n9386 & ~n10175 ;
  assign n10194 = ~n8293 & ~n8333 ;
  assign n10195 = ~n10176 & n10194 ;
  assign n10196 = ~n10178 & n10195 ;
  assign n10197 = ~n10174 & n10196 ;
  assign n10198 = ~n10181 & n10197 ;
  assign n10199 = ~n10193 & n10198 ;
  assign n10200 = \sa01_reg[0]/P0001  & ~n10199 ;
  assign n10202 = \sa01_reg[6]/NET0131  & n9173 ;
  assign n10203 = ~n9237 & ~n10202 ;
  assign n10204 = ~n9361 & n10203 ;
  assign n10205 = ~\sa01_reg[2]/P0001  & ~n10204 ;
  assign n10206 = ~n8219 & ~n8310 ;
  assign n10207 = n9698 & ~n10206 ;
  assign n10208 = n8245 & ~n8264 ;
  assign n10209 = n9318 & n10208 ;
  assign n10221 = ~n10207 & ~n10209 ;
  assign n10222 = ~n10205 & n10221 ;
  assign n10210 = ~\sa01_reg[3]/P0001  & ~n9728 ;
  assign n10211 = ~n8241 & ~n10210 ;
  assign n10212 = ~\sa01_reg[1]/P0001  & ~n10211 ;
  assign n10216 = n8277 & n8329 ;
  assign n10215 = n8235 & n8238 ;
  assign n10213 = n8254 & n9694 ;
  assign n10214 = n8215 & ~n8238 ;
  assign n10217 = ~n10213 & ~n10214 ;
  assign n10218 = ~n10215 & n10217 ;
  assign n10219 = ~n10216 & n10218 ;
  assign n10220 = \sa01_reg[1]/P0001  & ~n10219 ;
  assign n10223 = ~n10212 & ~n10220 ;
  assign n10224 = n10222 & n10223 ;
  assign n10225 = ~\sa01_reg[0]/P0001  & ~n10224 ;
  assign n10226 = ~n8308 & n8326 ;
  assign n10227 = ~n8363 & ~n10226 ;
  assign n10228 = ~\sa01_reg[2]/P0001  & ~n10227 ;
  assign n10230 = \sa01_reg[2]/P0001  & n8267 ;
  assign n10231 = ~n8257 & ~n8344 ;
  assign n10232 = n10230 & ~n10231 ;
  assign n10229 = ~\sa01_reg[2]/P0001  & n9256 ;
  assign n10233 = ~n9277 & ~n10229 ;
  assign n10234 = ~n10232 & n10233 ;
  assign n10235 = ~n10228 & n10234 ;
  assign n10236 = ~\sa01_reg[1]/P0001  & ~n10235 ;
  assign n10240 = ~n8220 & ~n8268 ;
  assign n10241 = ~n9207 & ~n9322 ;
  assign n10242 = n10240 & n10241 ;
  assign n10243 = \sa01_reg[1]/P0001  & ~n10242 ;
  assign n10201 = n8222 & n8293 ;
  assign n10237 = \sa01_reg[1]/P0001  & n9774 ;
  assign n10238 = ~n10215 & ~n10237 ;
  assign n10239 = ~\sa01_reg[2]/P0001  & ~n10238 ;
  assign n10244 = ~n10201 & ~n10239 ;
  assign n10245 = ~n10243 & n10244 ;
  assign n10246 = ~n10236 & n10245 ;
  assign n10247 = ~n10225 & n10246 ;
  assign n10248 = ~n10200 & n10247 ;
  assign n10249 = ~n9783 & ~n10248 ;
  assign n10250 = n9783 & n10248 ;
  assign n10251 = ~n10249 & ~n10250 ;
  assign n10252 = n10170 & ~n10251 ;
  assign n10253 = ~n10170 & n10251 ;
  assign n10254 = ~n10252 & ~n10253 ;
  assign n10258 = ~n8706 & ~n8823 ;
  assign n10259 = ~n8951 & n10258 ;
  assign n10260 = \sa30_reg[2]/P0001  & ~n10259 ;
  assign n10255 = ~\sa30_reg[3]/P0001  & n8682 ;
  assign n10256 = ~\sa30_reg[5]/P0001  & n10255 ;
  assign n10257 = n8741 & n10256 ;
  assign n10261 = \sa30_reg[5]/P0001  & ~n8682 ;
  assign n10262 = n8725 & ~n10261 ;
  assign n10263 = n8698 & n8756 ;
  assign n10264 = ~n10262 & ~n10263 ;
  assign n10265 = ~n10257 & n10264 ;
  assign n10266 = ~n10260 & n10265 ;
  assign n10267 = ~\sa30_reg[1]/P0001  & ~n10266 ;
  assign n10280 = ~n8786 & ~n9543 ;
  assign n10281 = n8870 & n10280 ;
  assign n10282 = \sa30_reg[2]/P0001  & ~n10281 ;
  assign n10268 = ~n8697 & ~n8950 ;
  assign n10269 = ~\sa30_reg[2]/P0001  & ~n10268 ;
  assign n10270 = ~n8961 & ~n10269 ;
  assign n10271 = \sa30_reg[1]/P0001  & ~n10270 ;
  assign n10275 = \sa30_reg[6]/NET0131  & n8930 ;
  assign n10276 = n8721 & n8756 ;
  assign n10277 = ~n10275 & ~n10276 ;
  assign n10278 = ~\sa30_reg[2]/P0001  & ~n10277 ;
  assign n10272 = \sa30_reg[3]/P0001  & n8792 ;
  assign n10273 = ~n8838 & ~n10272 ;
  assign n10274 = ~\sa30_reg[2]/P0001  & ~n10273 ;
  assign n10279 = \sa30_reg[5]/P0001  & n8835 ;
  assign n10283 = ~n9608 & ~n10279 ;
  assign n10284 = ~n10274 & n10283 ;
  assign n10285 = ~n10278 & n10284 ;
  assign n10286 = ~n10271 & n10285 ;
  assign n10287 = ~n10282 & n10286 ;
  assign n10288 = ~n10267 & n10287 ;
  assign n10289 = \sa30_reg[0]/P0002  & ~n10288 ;
  assign n10290 = \sa30_reg[6]/NET0131  & n8704 ;
  assign n10291 = ~n8786 & ~n10290 ;
  assign n10292 = ~n8916 & n10291 ;
  assign n10293 = ~\sa30_reg[2]/P0001  & ~n10292 ;
  assign n10294 = ~\sa30_reg[1]/P0001  & \sa30_reg[2]/P0001  ;
  assign n10295 = n8694 & ~n8758 ;
  assign n10296 = n10294 & n10295 ;
  assign n10297 = \sa30_reg[3]/P0001  & n9575 ;
  assign n10298 = ~n8792 & ~n8845 ;
  assign n10299 = n10297 & ~n10298 ;
  assign n10311 = ~n10296 & ~n10299 ;
  assign n10312 = ~n10293 & n10311 ;
  assign n10300 = ~n8767 & ~n8952 ;
  assign n10301 = ~\sa30_reg[3]/P0001  & ~n10300 ;
  assign n10302 = ~n9581 & ~n10301 ;
  assign n10303 = ~\sa30_reg[1]/P0001  & ~n10302 ;
  assign n10304 = n8705 & n8844 ;
  assign n10306 = ~n8724 & ~n8733 ;
  assign n10305 = n8833 & n8874 ;
  assign n10307 = ~n9603 & ~n10305 ;
  assign n10308 = n10306 & n10307 ;
  assign n10309 = ~n10304 & n10308 ;
  assign n10310 = \sa30_reg[1]/P0001  & ~n10309 ;
  assign n10313 = ~n10303 & ~n10310 ;
  assign n10314 = n10312 & n10313 ;
  assign n10315 = ~\sa30_reg[0]/P0002  & ~n10314 ;
  assign n10326 = ~n8735 & ~n9565 ;
  assign n10327 = ~\sa30_reg[7]/P0001  & ~n10326 ;
  assign n10328 = ~\sa30_reg[3]/P0001  & n8814 ;
  assign n10329 = ~n10327 & ~n10328 ;
  assign n10330 = ~\sa30_reg[2]/P0001  & ~n10329 ;
  assign n10333 = \sa30_reg[7]/P0001  & n8916 ;
  assign n10334 = ~n8699 & ~n10333 ;
  assign n10335 = \sa30_reg[2]/P0001  & ~n10334 ;
  assign n10331 = ~\sa30_reg[2]/P0001  & n8705 ;
  assign n10332 = n8725 & n10331 ;
  assign n10336 = ~n8847 & ~n10332 ;
  assign n10337 = ~n10335 & n10336 ;
  assign n10338 = ~n10330 & n10337 ;
  assign n10339 = ~\sa30_reg[1]/P0001  & ~n10338 ;
  assign n10316 = ~\sa30_reg[2]/P0001  & ~n8785 ;
  assign n10317 = ~n9592 & ~n10316 ;
  assign n10318 = n8929 & n9614 ;
  assign n10319 = ~n8916 & ~n9620 ;
  assign n10320 = ~n10318 & n10319 ;
  assign n10321 = ~\sa30_reg[7]/P0001  & ~n10320 ;
  assign n10322 = ~n10317 & ~n10321 ;
  assign n10323 = \sa30_reg[1]/P0001  & ~n10322 ;
  assign n10324 = ~\sa30_reg[2]/P0001  & n9603 ;
  assign n10325 = n9575 & n10279 ;
  assign n10340 = ~n10324 & ~n10325 ;
  assign n10341 = ~n10323 & n10340 ;
  assign n10342 = ~n10339 & n10341 ;
  assign n10343 = ~n10315 & n10342 ;
  assign n10344 = ~n10289 & n10343 ;
  assign n10377 = ~n9620 & ~n10331 ;
  assign n10375 = ~\sa30_reg[4]/P0001  & n8874 ;
  assign n10376 = n8929 & n10375 ;
  assign n10372 = ~n8684 & n8741 ;
  assign n10373 = ~n8710 & n10372 ;
  assign n10374 = n8835 & ~n9575 ;
  assign n10378 = ~n10373 & ~n10374 ;
  assign n10379 = ~n10376 & n10378 ;
  assign n10380 = n10377 & n10379 ;
  assign n10381 = ~\sa30_reg[1]/P0001  & ~n10380 ;
  assign n10385 = ~n8685 & ~n8743 ;
  assign n10386 = ~\sa30_reg[3]/P0001  & ~n10385 ;
  assign n10387 = ~n8706 & ~n10386 ;
  assign n10388 = \sa30_reg[2]/P0001  & ~n10387 ;
  assign n10390 = ~n8724 & ~n8766 ;
  assign n10389 = \sa30_reg[4]/P0001  & n8775 ;
  assign n10391 = ~n8888 & ~n10389 ;
  assign n10392 = n10390 & n10391 ;
  assign n10393 = n8946 & ~n10392 ;
  assign n10382 = n8682 & n8871 ;
  assign n10383 = ~n9604 & ~n10382 ;
  assign n10384 = \sa30_reg[1]/P0001  & ~n10383 ;
  assign n10395 = n8741 & n8835 ;
  assign n10394 = n8792 & n10297 ;
  assign n10396 = ~n10276 & ~n10394 ;
  assign n10397 = ~n10395 & n10396 ;
  assign n10398 = ~n10384 & n10397 ;
  assign n10399 = ~n10393 & n10398 ;
  assign n10400 = ~n10388 & n10399 ;
  assign n10401 = ~n10381 & n10400 ;
  assign n10402 = \sa30_reg[0]/P0002  & ~n10401 ;
  assign n10361 = ~n9560 & ~n9632 ;
  assign n10362 = ~\sa30_reg[2]/P0001  & ~n10361 ;
  assign n10363 = \sa30_reg[3]/P0001  & n8692 ;
  assign n10364 = ~n8915 & ~n10318 ;
  assign n10365 = ~n10363 & n10364 ;
  assign n10366 = ~n10362 & n10365 ;
  assign n10367 = \sa30_reg[1]/P0001  & ~n10366 ;
  assign n10355 = ~\sa30_reg[3]/P0001  & n8816 ;
  assign n10356 = ~n10263 & ~n10355 ;
  assign n10357 = ~\sa30_reg[6]/NET0131  & n8774 ;
  assign n10358 = ~n8822 & ~n10357 ;
  assign n10359 = n10356 & n10358 ;
  assign n10360 = ~\sa30_reg[2]/P0001  & ~n10359 ;
  assign n10345 = ~n8773 & ~n9582 ;
  assign n10346 = \sa30_reg[7]/P0001  & ~n10345 ;
  assign n10347 = n8844 & n9547 ;
  assign n10348 = ~n9553 & ~n10347 ;
  assign n10349 = ~n10346 & n10348 ;
  assign n10350 = ~\sa30_reg[1]/P0001  & ~n10349 ;
  assign n10351 = \sa30_reg[4]/P0001  & n8845 ;
  assign n10352 = ~n8749 & ~n10275 ;
  assign n10353 = ~n10351 & n10352 ;
  assign n10354 = n8844 & ~n10353 ;
  assign n10368 = ~n10350 & ~n10354 ;
  assign n10369 = ~n10360 & n10368 ;
  assign n10370 = ~n10367 & n10369 ;
  assign n10371 = ~\sa30_reg[0]/P0002  & ~n10370 ;
  assign n10418 = ~\sa30_reg[6]/NET0131  & n8757 ;
  assign n10419 = ~n8743 & ~n9572 ;
  assign n10420 = ~n10418 & n10419 ;
  assign n10421 = ~\sa30_reg[3]/P0001  & ~n10420 ;
  assign n10422 = ~n8744 & ~n8759 ;
  assign n10423 = ~n10421 & n10422 ;
  assign n10424 = n8946 & ~n10423 ;
  assign n10414 = ~n8785 & ~n8922 ;
  assign n10415 = n10356 & n10414 ;
  assign n10413 = \sa30_reg[2]/P0001  & ~n8785 ;
  assign n10416 = ~\sa30_reg[1]/P0001  & ~n10413 ;
  assign n10417 = ~n10415 & n10416 ;
  assign n10403 = \sa30_reg[5]/P0001  & n8735 ;
  assign n10404 = ~n8703 & ~n9604 ;
  assign n10405 = ~n10403 & n10404 ;
  assign n10406 = n10294 & ~n10405 ;
  assign n10407 = ~n8685 & ~n8845 ;
  assign n10408 = n10300 & n10407 ;
  assign n10409 = \sa30_reg[1]/P0001  & n8940 ;
  assign n10410 = ~n10408 & n10409 ;
  assign n10411 = ~n8700 & ~n9561 ;
  assign n10412 = ~\sa30_reg[2]/P0001  & ~n10411 ;
  assign n10425 = ~n10410 & ~n10412 ;
  assign n10426 = ~n10406 & n10425 ;
  assign n10427 = ~n10417 & n10426 ;
  assign n10428 = ~n10424 & n10427 ;
  assign n10429 = ~n10371 & n10428 ;
  assign n10430 = ~n10402 & n10429 ;
  assign n10431 = n10344 & ~n10430 ;
  assign n10432 = ~n10344 & n10430 ;
  assign n10433 = ~n10431 & ~n10432 ;
  assign n10435 = n8509 & n8519 ;
  assign n10438 = ~\sa23_reg[1]/P0001  & ~n9964 ;
  assign n10439 = ~n10435 & n10438 ;
  assign n10436 = \sa23_reg[4]/P0001  & n8618 ;
  assign n10437 = n8512 & ~n9900 ;
  assign n10440 = ~n10436 & ~n10437 ;
  assign n10441 = n10439 & n10440 ;
  assign n10444 = ~n9096 & ~n9151 ;
  assign n10445 = ~n9453 & n10444 ;
  assign n10446 = \sa23_reg[2]/P0001  & ~n10445 ;
  assign n10442 = n8521 & n9066 ;
  assign n10443 = ~n8563 & ~n10442 ;
  assign n10447 = \sa23_reg[1]/P0001  & n10443 ;
  assign n10448 = ~n10446 & n10447 ;
  assign n10449 = ~n10441 & ~n10448 ;
  assign n10450 = ~n9154 & ~n9964 ;
  assign n10451 = ~n9492 & n10450 ;
  assign n10452 = ~\sa23_reg[2]/P0001  & ~n10451 ;
  assign n10453 = n8527 & ~n9427 ;
  assign n10434 = ~n8546 & n8667 ;
  assign n10454 = \sa23_reg[0]/P0001  & ~n10434 ;
  assign n10455 = ~n10453 & n10454 ;
  assign n10456 = ~n10452 & n10455 ;
  assign n10457 = ~n10449 & n10456 ;
  assign n10458 = ~n9074 & n9153 ;
  assign n10459 = \sa23_reg[2]/P0001  & ~n9097 ;
  assign n10460 = ~n9492 & n10459 ;
  assign n10461 = ~n10458 & ~n10460 ;
  assign n10462 = ~\sa23_reg[1]/P0001  & ~n9130 ;
  assign n10463 = ~n9476 & n10462 ;
  assign n10464 = ~n10461 & n10463 ;
  assign n10466 = ~\sa23_reg[2]/P0001  & ~n8548 ;
  assign n10467 = ~n8550 & ~n9129 ;
  assign n10468 = n10466 & n10467 ;
  assign n10469 = \sa23_reg[2]/P0001  & ~n9113 ;
  assign n10470 = ~n9942 & n10469 ;
  assign n10471 = ~n10468 & ~n10470 ;
  assign n10465 = \sa23_reg[1]/P0001  & ~n8530 ;
  assign n10472 = n8592 & n10465 ;
  assign n10473 = ~n10471 & n10472 ;
  assign n10474 = ~n10464 & ~n10473 ;
  assign n10475 = \sa23_reg[2]/P0001  & ~n8523 ;
  assign n10476 = ~n9128 & n10475 ;
  assign n10477 = ~\sa23_reg[2]/P0001  & ~n8663 ;
  assign n10478 = ~n8633 & ~n9476 ;
  assign n10479 = n10477 & n10478 ;
  assign n10480 = ~n10476 & ~n10479 ;
  assign n10481 = ~\sa23_reg[0]/P0001  & ~n8668 ;
  assign n10482 = ~n10480 & n10481 ;
  assign n10483 = ~n10474 & n10482 ;
  assign n10484 = ~n10457 & ~n10483 ;
  assign n10485 = ~\sa23_reg[1]/P0001  & ~n8632 ;
  assign n10486 = ~n8641 & ~n8663 ;
  assign n10487 = ~n9893 & n10486 ;
  assign n10488 = n10485 & n10487 ;
  assign n10489 = ~n8533 & ~n8563 ;
  assign n10490 = \sa23_reg[3]/P0001  & ~n10489 ;
  assign n10491 = \sa23_reg[1]/P0001  & ~n9107 ;
  assign n10492 = ~n10490 & n10491 ;
  assign n10493 = ~n10488 & ~n10492 ;
  assign n10494 = ~n8670 & ~n9467 ;
  assign n10495 = ~n10493 & n10494 ;
  assign n10496 = \sa23_reg[2]/P0001  & ~n10495 ;
  assign n10501 = ~n9078 & ~n9927 ;
  assign n10502 = ~n8636 & n10501 ;
  assign n10503 = ~n9467 & n10502 ;
  assign n10504 = n10485 & n10503 ;
  assign n10497 = ~n8509 & ~n8568 ;
  assign n10498 = ~n8569 & ~n10497 ;
  assign n10499 = ~n9085 & n10465 ;
  assign n10500 = ~n10498 & n10499 ;
  assign n10505 = ~\sa23_reg[2]/P0001  & ~n10500 ;
  assign n10506 = ~n10504 & n10505 ;
  assign n10507 = ~n10496 & ~n10506 ;
  assign n10508 = ~n10484 & n10507 ;
  assign n10509 = \u0_w_reg[1][1]/P0001  & ~n10508 ;
  assign n10510 = ~\u0_w_reg[1][1]/P0001  & n10508 ;
  assign n10511 = ~n10509 & ~n10510 ;
  assign n10512 = n10433 & n10511 ;
  assign n10513 = ~n10433 & ~n10511 ;
  assign n10514 = ~n10512 & ~n10513 ;
  assign n10516 = n10254 & n10514 ;
  assign n10515 = ~n10254 & ~n10514 ;
  assign n10517 = ~\ld_r_reg/P0001  & ~n10515 ;
  assign n10518 = ~n10516 & n10517 ;
  assign n10520 = \text_in_r_reg[65]/P0001  & \u0_w_reg[1][1]/P0001  ;
  assign n10519 = ~\text_in_r_reg[65]/P0001  & ~\u0_w_reg[1][1]/P0001  ;
  assign n10521 = \ld_r_reg/P0001  & ~n10519 ;
  assign n10522 = ~n10520 & n10521 ;
  assign n10523 = ~n10518 & ~n10522 ;
  assign n10524 = \u0_w_reg[1][28]/P0001  & ~n9639 ;
  assign n10525 = ~\u0_w_reg[1][28]/P0001  & n9639 ;
  assign n10526 = ~n10524 & ~n10525 ;
  assign n10527 = n9519 & n10526 ;
  assign n10528 = ~n9519 & ~n10526 ;
  assign n10529 = ~n10527 & ~n10528 ;
  assign n10569 = ~n8279 & ~n8331 ;
  assign n10570 = ~n9184 & n10569 ;
  assign n10571 = \sa01_reg[2]/P0001  & ~n10570 ;
  assign n10566 = n8240 & ~n8242 ;
  assign n10567 = ~n9215 & ~n10566 ;
  assign n10568 = ~n8264 & ~n10567 ;
  assign n10572 = ~n8269 & ~n10568 ;
  assign n10573 = ~n10571 & n10572 ;
  assign n10574 = \sa01_reg[1]/P0001  & ~n10573 ;
  assign n10553 = n8353 & ~n9741 ;
  assign n10554 = \sa01_reg[2]/P0001  & ~n8277 ;
  assign n10555 = ~n9231 & n10554 ;
  assign n10556 = ~n10553 & ~n10555 ;
  assign n10557 = ~n8362 & ~n9376 ;
  assign n10558 = ~n9322 & n10557 ;
  assign n10559 = ~n10157 & n10558 ;
  assign n10560 = ~n10556 & n10559 ;
  assign n10561 = ~\sa01_reg[1]/P0001  & ~n10560 ;
  assign n10562 = ~n9710 & n10203 ;
  assign n10563 = ~\sa01_reg[2]/P0001  & ~n10562 ;
  assign n10564 = ~n9183 & n9263 ;
  assign n10565 = n8327 & ~n10564 ;
  assign n10575 = ~n9256 & ~n10565 ;
  assign n10576 = ~n10563 & n10575 ;
  assign n10577 = ~n10561 & n10576 ;
  assign n10578 = ~n10574 & n10577 ;
  assign n10579 = \sa01_reg[0]/P0001  & ~n10578 ;
  assign n10537 = ~n9216 & ~n9357 ;
  assign n10538 = \sa01_reg[2]/P0001  & ~n10537 ;
  assign n10539 = n8246 & n8279 ;
  assign n10540 = ~n8255 & ~n10083 ;
  assign n10541 = ~n10539 & n10540 ;
  assign n10542 = ~n8322 & n10541 ;
  assign n10543 = ~n10538 & n10542 ;
  assign n10544 = \sa01_reg[1]/P0001  & ~n10543 ;
  assign n10531 = n8215 & n8327 ;
  assign n10532 = ~n9710 & ~n10531 ;
  assign n10533 = ~n9387 & n10532 ;
  assign n10530 = n8228 & n9197 ;
  assign n10534 = ~n9389 & ~n10530 ;
  assign n10535 = n10533 & n10534 ;
  assign n10536 = ~\sa01_reg[1]/P0001  & ~n10535 ;
  assign n10545 = ~\sa01_reg[2]/P0001  & ~n9323 ;
  assign n10546 = n8329 & n9216 ;
  assign n10547 = ~n9253 & ~n9374 ;
  assign n10548 = ~n10546 & n10547 ;
  assign n10549 = ~n10545 & n10548 ;
  assign n10550 = ~n10536 & n10549 ;
  assign n10551 = ~n10544 & n10550 ;
  assign n10552 = ~\sa01_reg[0]/P0001  & ~n10551 ;
  assign n10582 = \sa01_reg[6]/NET0131  & n8265 ;
  assign n10583 = ~n9180 & ~n9352 ;
  assign n10584 = ~n10582 & n10583 ;
  assign n10585 = n9694 & ~n10584 ;
  assign n10581 = ~\sa01_reg[2]/P0001  & n8333 ;
  assign n10586 = ~n8244 & ~n10581 ;
  assign n10587 = ~n10585 & n10586 ;
  assign n10588 = \sa01_reg[1]/P0001  & ~n10587 ;
  assign n10589 = ~n8217 & ~n9253 ;
  assign n10590 = n9318 & ~n10589 ;
  assign n10580 = n8236 & n10145 ;
  assign n10595 = ~n10116 & ~n10144 ;
  assign n10596 = ~n10580 & n10595 ;
  assign n10591 = n8218 & n8257 ;
  assign n10592 = ~n8269 & ~n10591 ;
  assign n10593 = n9388 & ~n10592 ;
  assign n10594 = \sa01_reg[7]/NET0131  & n9699 ;
  assign n10597 = ~n10593 & ~n10594 ;
  assign n10598 = n10596 & n10597 ;
  assign n10599 = ~n10590 & n10598 ;
  assign n10600 = ~n10588 & n10599 ;
  assign n10601 = ~n10552 & n10600 ;
  assign n10602 = ~n10579 & n10601 ;
  assign n10603 = n9783 & ~n10602 ;
  assign n10604 = ~n9783 & n10602 ;
  assign n10605 = ~n10603 & ~n10604 ;
  assign n10648 = ~n8127 & ~n8443 ;
  assign n10649 = ~n8162 & ~n10648 ;
  assign n10646 = ~n8096 & ~n9042 ;
  assign n10647 = ~\sa12_reg[2]/P0001  & ~n10646 ;
  assign n10650 = ~n8394 & ~n8485 ;
  assign n10651 = ~n8189 & n10650 ;
  assign n10652 = ~n10647 & n10651 ;
  assign n10653 = ~n10649 & n10652 ;
  assign n10654 = ~\sa12_reg[1]/P0001  & ~n10653 ;
  assign n10634 = ~n8182 & ~n8185 ;
  assign n10635 = ~n10055 & n10634 ;
  assign n10636 = \sa12_reg[2]/P0001  & ~n10635 ;
  assign n10631 = ~n8077 & n9841 ;
  assign n10632 = ~n8165 & ~n10631 ;
  assign n10633 = ~n8075 & ~n10632 ;
  assign n10637 = ~n8136 & ~n10633 ;
  assign n10638 = ~n10636 & n10637 ;
  assign n10639 = \sa12_reg[1]/P0001  & ~n10638 ;
  assign n10640 = \sa12_reg[6]/NET0131  & n8389 ;
  assign n10641 = ~n8461 & ~n10640 ;
  assign n10642 = ~n9801 & n10641 ;
  assign n10643 = ~\sa12_reg[2]/P0001  & ~n10642 ;
  assign n10644 = ~n8381 & n8482 ;
  assign n10645 = n8066 & ~n10644 ;
  assign n10655 = ~n8449 & ~n10645 ;
  assign n10656 = ~n10643 & n10655 ;
  assign n10657 = ~n10639 & n10656 ;
  assign n10658 = ~n10654 & n10657 ;
  assign n10659 = \sa12_reg[0]/P0001  & ~n10658 ;
  assign n10607 = ~n8414 & ~n8495 ;
  assign n10608 = \sa12_reg[2]/P0001  & ~n10607 ;
  assign n10610 = \sa12_reg[1]/P0001  & ~n8127 ;
  assign n10611 = ~n8115 & n10610 ;
  assign n10609 = n8077 & n9846 ;
  assign n10612 = ~n9996 & ~n10609 ;
  assign n10613 = n10611 & n10612 ;
  assign n10614 = ~n10608 & n10613 ;
  assign n10615 = ~n8082 & n8084 ;
  assign n10616 = ~n8156 & ~n10615 ;
  assign n10617 = \sa12_reg[2]/P0001  & ~n10616 ;
  assign n10618 = ~\sa12_reg[1]/P0001  & ~n9801 ;
  assign n10619 = ~n9034 & n10618 ;
  assign n10620 = ~n9041 & n10619 ;
  assign n10621 = ~n10617 & n10620 ;
  assign n10622 = ~n10614 & ~n10621 ;
  assign n10623 = ~\sa12_reg[2]/P0001  & ~n8993 ;
  assign n10606 = ~\sa12_reg[4]/P0001  & n8413 ;
  assign n10624 = n8110 & n8498 ;
  assign n10625 = ~n9044 & ~n10624 ;
  assign n10626 = \sa12_reg[2]/P0001  & ~n10625 ;
  assign n10627 = ~n10606 & ~n10626 ;
  assign n10628 = ~n10623 & n10627 ;
  assign n10629 = ~n10622 & n10628 ;
  assign n10630 = ~\sa12_reg[0]/P0001  & ~n10629 ;
  assign n10669 = ~n8146 & ~n8388 ;
  assign n10670 = ~n9025 & n10669 ;
  assign n10671 = n8978 & ~n10670 ;
  assign n10672 = ~\sa12_reg[2]/P0001  & n8113 ;
  assign n10673 = ~n8167 & ~n10672 ;
  assign n10674 = ~n10671 & n10673 ;
  assign n10675 = \sa12_reg[1]/P0001  & ~n10674 ;
  assign n10666 = n8059 & n9034 ;
  assign n10667 = ~n8448 & ~n10666 ;
  assign n10668 = ~\sa12_reg[1]/P0001  & ~n10667 ;
  assign n10660 = \sa12_reg[2]/P0001  & n8136 ;
  assign n10661 = n8159 & n10060 ;
  assign n10662 = ~n10660 & ~n10661 ;
  assign n10663 = ~\sa12_reg[4]/P0001  & ~n10662 ;
  assign n10664 = ~n8097 & ~n8136 ;
  assign n10665 = n9033 & ~n10664 ;
  assign n10676 = ~n10024 & ~n10063 ;
  assign n10677 = ~n10665 & n10676 ;
  assign n10678 = ~n10663 & n10677 ;
  assign n10679 = ~n10668 & n10678 ;
  assign n10680 = ~n10675 & n10679 ;
  assign n10681 = ~n10630 & n10680 ;
  assign n10682 = ~n10659 & n10681 ;
  assign n10683 = n9874 & ~n10682 ;
  assign n10684 = ~n9874 & n10682 ;
  assign n10685 = ~n10683 & ~n10684 ;
  assign n10686 = ~n10605 & n10685 ;
  assign n10687 = n10605 & ~n10685 ;
  assign n10688 = ~n10686 & ~n10687 ;
  assign n10690 = ~n10529 & n10688 ;
  assign n10689 = n10529 & ~n10688 ;
  assign n10691 = ~\ld_r_reg/P0001  & ~n10689 ;
  assign n10692 = ~n10690 & n10691 ;
  assign n10694 = ~\text_in_r_reg[92]/P0001  & \u0_w_reg[1][28]/P0001  ;
  assign n10693 = \text_in_r_reg[92]/P0001  & ~\u0_w_reg[1][28]/P0001  ;
  assign n10695 = \ld_r_reg/P0001  & ~n10693 ;
  assign n10696 = ~n10694 & n10695 ;
  assign n10697 = ~n10692 & ~n10696 ;
  assign n10758 = ~\sa23_reg[1]/P0001  & ~n9468 ;
  assign n10754 = \sa23_reg[2]/P0001  & n8526 ;
  assign n10755 = ~n8547 & n10754 ;
  assign n10756 = ~n8547 & ~n8660 ;
  assign n10757 = n8623 & ~n10756 ;
  assign n10759 = ~n10755 & ~n10757 ;
  assign n10760 = n10758 & n10759 ;
  assign n10761 = ~n9134 & n10760 ;
  assign n10763 = \sa23_reg[1]/P0001  & ~n8615 ;
  assign n10764 = ~n8558 & n10763 ;
  assign n10762 = n8508 & n9922 ;
  assign n10765 = ~n10442 & ~n10762 ;
  assign n10766 = n10764 & n10765 ;
  assign n10767 = ~n10761 & ~n10766 ;
  assign n10747 = ~\sa23_reg[2]/P0001  & n9088 ;
  assign n10749 = ~n9101 & ~n9114 ;
  assign n10750 = \sa23_reg[1]/P0001  & ~n10749 ;
  assign n10748 = n8529 & n8577 ;
  assign n10751 = n9148 & ~n10748 ;
  assign n10752 = ~n10750 & n10751 ;
  assign n10753 = ~n10747 & ~n10752 ;
  assign n10768 = ~n8643 & ~n10753 ;
  assign n10769 = ~n10767 & n10768 ;
  assign n10770 = ~\sa23_reg[0]/P0001  & ~n10769 ;
  assign n10709 = ~n8598 & ~n8615 ;
  assign n10710 = n9497 & n10709 ;
  assign n10711 = ~\sa23_reg[2]/P0001  & ~n8527 ;
  assign n10712 = ~n9927 & n10711 ;
  assign n10713 = ~n10710 & ~n10712 ;
  assign n10714 = ~n8663 & ~n9158 ;
  assign n10715 = ~n9467 & n10714 ;
  assign n10716 = ~n10713 & n10715 ;
  assign n10717 = ~\sa23_reg[1]/P0001  & ~n10716 ;
  assign n10699 = ~n8509 & ~n9499 ;
  assign n10700 = ~n9920 & n10699 ;
  assign n10701 = \sa23_reg[2]/P0001  & ~n10700 ;
  assign n10703 = n8513 & n9079 ;
  assign n10704 = ~n9097 & ~n10703 ;
  assign n10698 = ~n8588 & n9113 ;
  assign n10702 = ~\sa23_reg[2]/P0001  & n9489 ;
  assign n10705 = ~n10698 & ~n10702 ;
  assign n10706 = n10704 & n10705 ;
  assign n10707 = ~n10701 & n10706 ;
  assign n10708 = \sa23_reg[1]/P0001  & ~n10707 ;
  assign n10718 = \sa23_reg[6]/NET0131  & n8532 ;
  assign n10719 = ~n8633 & ~n10718 ;
  assign n10720 = ~n9468 & n10719 ;
  assign n10721 = ~\sa23_reg[2]/P0001  & ~n10720 ;
  assign n10722 = ~n8512 & n8656 ;
  assign n10723 = n9931 & ~n10722 ;
  assign n10724 = ~n8647 & ~n10723 ;
  assign n10725 = ~n10721 & n10724 ;
  assign n10726 = ~n10708 & n10725 ;
  assign n10727 = ~n10717 & n10726 ;
  assign n10728 = \sa23_reg[0]/P0001  & ~n10727 ;
  assign n10733 = ~n8514 & ~n8520 ;
  assign n10734 = ~n9099 & n10733 ;
  assign n10735 = n9079 & ~n10734 ;
  assign n10730 = n8521 & n8572 ;
  assign n10731 = ~n9097 & ~n10730 ;
  assign n10732 = \sa23_reg[2]/P0001  & ~n10731 ;
  assign n10729 = ~\sa23_reg[2]/P0001  & n9454 ;
  assign n10736 = ~n9433 & ~n10729 ;
  assign n10737 = ~n10732 & n10736 ;
  assign n10738 = ~n10735 & n10737 ;
  assign n10739 = \sa23_reg[1]/P0001  & ~n10738 ;
  assign n10740 = ~n9125 & ~n9964 ;
  assign n10741 = n9112 & ~n10740 ;
  assign n10742 = n8588 & n9922 ;
  assign n10743 = ~n10741 & ~n10742 ;
  assign n10744 = ~\sa23_reg[1]/P0001  & ~n10743 ;
  assign n10745 = ~n8563 & ~n9420 ;
  assign n10746 = n8546 & ~n10745 ;
  assign n10771 = ~n9130 & ~n10746 ;
  assign n10772 = ~n10744 & n10771 ;
  assign n10773 = ~n10739 & n10772 ;
  assign n10774 = ~n10728 & n10773 ;
  assign n10775 = ~n10770 & n10774 ;
  assign n10776 = n8376 & ~n10775 ;
  assign n10777 = ~n8376 & n10775 ;
  assign n10778 = ~n10776 & ~n10777 ;
  assign n10779 = n10685 & n10778 ;
  assign n10780 = ~n10685 & ~n10778 ;
  assign n10781 = ~n10779 & ~n10780 ;
  assign n10782 = ~n9516 & ~n9639 ;
  assign n10783 = n9516 & n9639 ;
  assign n10784 = ~n10782 & ~n10783 ;
  assign n10785 = \u0_w_reg[1][20]/P0001  & ~n9980 ;
  assign n10786 = ~\u0_w_reg[1][20]/P0001  & n9980 ;
  assign n10787 = ~n10785 & ~n10786 ;
  assign n10788 = n10784 & n10787 ;
  assign n10789 = ~n10784 & ~n10787 ;
  assign n10790 = ~n10788 & ~n10789 ;
  assign n10792 = ~n10781 & n10790 ;
  assign n10791 = n10781 & ~n10790 ;
  assign n10793 = ~\ld_r_reg/P0001  & ~n10791 ;
  assign n10794 = ~n10792 & n10793 ;
  assign n10796 = ~\text_in_r_reg[84]/P0001  & \u0_w_reg[1][20]/P0001  ;
  assign n10795 = \text_in_r_reg[84]/P0001  & ~\u0_w_reg[1][20]/P0001  ;
  assign n10797 = \ld_r_reg/P0001  & ~n10795 ;
  assign n10798 = ~n10796 & n10797 ;
  assign n10799 = ~n10794 & ~n10798 ;
  assign n10800 = ~n8376 & ~n9292 ;
  assign n10801 = n8376 & n9292 ;
  assign n10802 = ~n10800 & ~n10801 ;
  assign n10803 = \u0_w_reg[1][5]/P0001  & ~n9639 ;
  assign n10804 = ~\u0_w_reg[1][5]/P0001  & n9639 ;
  assign n10805 = ~n10803 & ~n10804 ;
  assign n10806 = n8678 & n10805 ;
  assign n10807 = ~n8678 & ~n10805 ;
  assign n10808 = ~n10806 & ~n10807 ;
  assign n10810 = n10802 & ~n10808 ;
  assign n10809 = ~n10802 & n10808 ;
  assign n10811 = ~\ld_r_reg/P0001  & ~n10809 ;
  assign n10812 = ~n10810 & n10811 ;
  assign n10814 = \text_in_r_reg[69]/P0001  & \u0_w_reg[1][5]/P0001  ;
  assign n10813 = ~\text_in_r_reg[69]/P0001  & ~\u0_w_reg[1][5]/P0001  ;
  assign n10815 = \ld_r_reg/P0001  & ~n10813 ;
  assign n10816 = ~n10814 & n10815 ;
  assign n10817 = ~n10812 & ~n10816 ;
  assign n10818 = ~n9639 & ~n10430 ;
  assign n10819 = n9639 & n10430 ;
  assign n10820 = ~n10818 & ~n10819 ;
  assign n10861 = ~n8705 & ~n8757 ;
  assign n10862 = n9592 & n10861 ;
  assign n10863 = ~n9633 & ~n10862 ;
  assign n10864 = n8775 & n8896 ;
  assign n10865 = ~n8699 & ~n8810 ;
  assign n10866 = ~n8834 & n10865 ;
  assign n10867 = ~n10864 & n10866 ;
  assign n10868 = ~n10863 & n10867 ;
  assign n10869 = ~\sa30_reg[1]/P0001  & ~n10868 ;
  assign n10850 = ~n8692 & ~n8884 ;
  assign n10851 = ~n9547 & n10850 ;
  assign n10852 = \sa30_reg[2]/P0001  & ~n10851 ;
  assign n10847 = ~n8835 & ~n8950 ;
  assign n10848 = ~\sa30_reg[2]/P0001  & ~n10847 ;
  assign n10849 = \sa30_reg[4]/P0001  & n10295 ;
  assign n10853 = ~n9596 & ~n10849 ;
  assign n10854 = ~n10848 & n10853 ;
  assign n10855 = ~n10852 & n10854 ;
  assign n10856 = \sa30_reg[1]/P0001  & ~n10855 ;
  assign n10857 = ~n8875 & n10291 ;
  assign n10858 = ~\sa30_reg[2]/P0001  & ~n10857 ;
  assign n10859 = ~n8683 & n8815 ;
  assign n10860 = n8811 & ~n10859 ;
  assign n10870 = ~n8764 & ~n10860 ;
  assign n10871 = ~n10858 & n10870 ;
  assign n10872 = ~n10856 & n10871 ;
  assign n10873 = ~n10869 & n10872 ;
  assign n10874 = \sa30_reg[0]/P0002  & ~n10873 ;
  assign n10822 = ~\sa30_reg[3]/P0001  & n8706 ;
  assign n10823 = ~n8748 & ~n10822 ;
  assign n10824 = \sa30_reg[2]/P0001  & ~n10823 ;
  assign n10826 = \sa30_reg[1]/P0001  & ~n8796 ;
  assign n10827 = ~n8720 & n10826 ;
  assign n10821 = \sa30_reg[7]/P0001  & n8821 ;
  assign n10825 = n8692 & n9582 ;
  assign n10828 = ~n10821 & ~n10825 ;
  assign n10829 = n10827 & n10828 ;
  assign n10830 = ~n10824 & n10829 ;
  assign n10831 = n8701 & n8811 ;
  assign n10834 = ~\sa30_reg[1]/P0001  & ~n8875 ;
  assign n10835 = ~n10831 & n10834 ;
  assign n10832 = \sa30_reg[7]/P0001  & ~n8775 ;
  assign n10833 = n8929 & n10832 ;
  assign n10836 = ~n10357 & ~n10833 ;
  assign n10837 = n10835 & n10836 ;
  assign n10838 = ~n8941 & n10837 ;
  assign n10839 = ~n10830 & ~n10838 ;
  assign n10841 = ~n8839 & ~n8952 ;
  assign n10842 = \sa30_reg[2]/P0001  & ~n10841 ;
  assign n10840 = ~\sa30_reg[2]/P0001  & ~n8890 ;
  assign n10843 = ~n8768 & ~n10840 ;
  assign n10844 = ~n10842 & n10843 ;
  assign n10845 = ~n10839 & n10844 ;
  assign n10846 = ~\sa30_reg[0]/P0002  & ~n10845 ;
  assign n10876 = ~n8687 & ~n10389 ;
  assign n10877 = ~n8693 & n10876 ;
  assign n10878 = n8833 & ~n10877 ;
  assign n10875 = ~\sa30_reg[2]/P0001  & n9608 ;
  assign n10880 = n8697 & n10297 ;
  assign n10879 = n8710 & n8844 ;
  assign n10881 = ~n9585 & ~n10879 ;
  assign n10882 = ~n10880 & n10881 ;
  assign n10883 = ~n10875 & n10882 ;
  assign n10884 = ~n10878 & n10883 ;
  assign n10885 = \sa30_reg[1]/P0001  & ~n10884 ;
  assign n10886 = ~n8768 & ~n8784 ;
  assign n10887 = \sa30_reg[2]/P0001  & ~n10886 ;
  assign n10888 = \sa30_reg[7]/P0001  & n8758 ;
  assign n10889 = n9582 & n10888 ;
  assign n10890 = ~n10887 & ~n10889 ;
  assign n10891 = ~\sa30_reg[1]/P0001  & ~n10890 ;
  assign n10892 = ~n8744 & ~n9572 ;
  assign n10893 = n8844 & ~n10892 ;
  assign n10894 = ~n8956 & ~n10893 ;
  assign n10895 = ~n10891 & n10894 ;
  assign n10896 = ~n10885 & n10895 ;
  assign n10897 = ~n10846 & n10896 ;
  assign n10898 = ~n10874 & n10897 ;
  assign n10899 = \u0_w_reg[1][12]/P0001  & ~n10898 ;
  assign n10900 = ~\u0_w_reg[1][12]/P0001  & n10898 ;
  assign n10901 = ~n10899 & ~n10900 ;
  assign n10902 = n10820 & n10901 ;
  assign n10903 = ~n10820 & ~n10901 ;
  assign n10904 = ~n10902 & ~n10903 ;
  assign n10905 = n9980 & ~n10775 ;
  assign n10906 = ~n9980 & n10775 ;
  assign n10907 = ~n10905 & ~n10906 ;
  assign n10908 = ~n8379 & n10907 ;
  assign n10909 = n8379 & ~n10907 ;
  assign n10910 = ~n10908 & ~n10909 ;
  assign n10912 = n10904 & n10910 ;
  assign n10911 = ~n10904 & ~n10910 ;
  assign n10913 = ~\ld_r_reg/P0001  & ~n10911 ;
  assign n10914 = ~n10912 & n10913 ;
  assign n10916 = ~\text_in_r_reg[76]/P0001  & \u0_w_reg[1][12]/P0001  ;
  assign n10915 = \text_in_r_reg[76]/P0001  & ~\u0_w_reg[1][12]/P0001  ;
  assign n10917 = \ld_r_reg/P0001  & ~n10915 ;
  assign n10918 = ~n10916 & n10917 ;
  assign n10919 = ~n10914 & ~n10918 ;
  assign n10937 = ~\sa12_reg[3]/P0001  & n8142 ;
  assign n10938 = ~n8391 & ~n8452 ;
  assign n10939 = ~n10937 & n10938 ;
  assign n10940 = \sa12_reg[2]/P0001  & ~n10939 ;
  assign n10934 = \sa12_reg[5]/P0001  & ~n8126 ;
  assign n10935 = n8078 & ~n10934 ;
  assign n10933 = n8147 & n8978 ;
  assign n10936 = n8074 & n8104 ;
  assign n10941 = ~n10933 & ~n10936 ;
  assign n10942 = ~n10935 & n10941 ;
  assign n10943 = ~n10940 & n10942 ;
  assign n10944 = ~\sa12_reg[1]/P0001  & ~n10943 ;
  assign n10930 = ~n8184 & ~n8985 ;
  assign n10931 = n8462 & n10930 ;
  assign n10932 = \sa12_reg[2]/P0001  & ~n10931 ;
  assign n10925 = ~n8093 & ~n8498 ;
  assign n10926 = \sa12_reg[3]/P0001  & ~n10925 ;
  assign n10927 = ~n8432 & ~n8494 ;
  assign n10928 = ~n10926 & n10927 ;
  assign n10929 = ~\sa12_reg[2]/P0001  & ~n10928 ;
  assign n10920 = ~\sa12_reg[2]/P0001  & ~n8077 ;
  assign n10921 = ~\sa12_reg[5]/P0001  & ~n8055 ;
  assign n10922 = n10920 & ~n10921 ;
  assign n10923 = ~n9049 & ~n10922 ;
  assign n10924 = \sa12_reg[1]/P0001  & ~n10923 ;
  assign n10945 = ~n8113 & ~n8175 ;
  assign n10946 = ~n10924 & n10945 ;
  assign n10947 = ~n10929 & n10946 ;
  assign n10948 = ~n10932 & n10947 ;
  assign n10949 = ~n10944 & n10948 ;
  assign n10950 = \sa12_reg[0]/P0001  & ~n10949 ;
  assign n10952 = n8075 & n8080 ;
  assign n10954 = ~n9817 & ~n9821 ;
  assign n10955 = ~n10952 & n10954 ;
  assign n10951 = \sa12_reg[2]/P0001  & n8076 ;
  assign n10953 = \sa12_reg[1]/P0001  & ~n8417 ;
  assign n10956 = ~n10951 & n10953 ;
  assign n10957 = n10955 & n10956 ;
  assign n10960 = ~\sa12_reg[3]/P0001  & ~n9784 ;
  assign n10958 = \sa12_reg[2]/P0001  & ~n8075 ;
  assign n10959 = n8161 & n10958 ;
  assign n10961 = n8158 & ~n10959 ;
  assign n10962 = ~n10960 & n10961 ;
  assign n10963 = ~n10957 & ~n10962 ;
  assign n10964 = ~n8056 & ~n8093 ;
  assign n10965 = n8078 & ~n10964 ;
  assign n10966 = \sa12_reg[2]/P0001  & ~n10965 ;
  assign n10967 = ~\sa12_reg[2]/P0001  & ~n8117 ;
  assign n10968 = n10641 & n10967 ;
  assign n10969 = ~n10966 & ~n10968 ;
  assign n10970 = ~n10963 & ~n10969 ;
  assign n10971 = ~\sa12_reg[0]/P0001  & ~n10970 ;
  assign n10986 = ~n8061 & ~n8412 ;
  assign n10987 = ~n9790 & n10986 ;
  assign n10988 = n8978 & ~n10987 ;
  assign n10984 = n8074 & n8155 ;
  assign n10985 = n8068 & n10984 ;
  assign n10989 = ~n8491 & ~n10985 ;
  assign n10990 = ~n10988 & n10989 ;
  assign n10991 = ~\sa12_reg[1]/P0001  & ~n10990 ;
  assign n10979 = n8066 & n8413 ;
  assign n10977 = ~\sa12_reg[2]/P0001  & ~n9865 ;
  assign n10978 = ~n8128 & ~n10977 ;
  assign n10980 = ~n8118 & ~n8150 ;
  assign n10981 = ~n10978 & n10980 ;
  assign n10982 = ~n10979 & n10981 ;
  assign n10983 = \sa12_reg[1]/P0001  & ~n10982 ;
  assign n10972 = ~n8086 & ~n8394 ;
  assign n10973 = n10064 & ~n10972 ;
  assign n10974 = n8059 & n8174 ;
  assign n10975 = ~n10952 & ~n10974 ;
  assign n10976 = ~n8066 & ~n10975 ;
  assign n10992 = ~n10973 & ~n10976 ;
  assign n10993 = ~n10983 & n10992 ;
  assign n10994 = ~n10991 & n10993 ;
  assign n10995 = ~n10971 & n10994 ;
  assign n10996 = ~n10950 & n10995 ;
  assign n10997 = n9874 & ~n10996 ;
  assign n10998 = ~n9874 & n10996 ;
  assign n10999 = ~n10997 & ~n10998 ;
  assign n11015 = ~n8534 & ~n8602 ;
  assign n11016 = ~n9128 & n11015 ;
  assign n11017 = \sa23_reg[2]/P0001  & ~n11016 ;
  assign n11012 = \sa23_reg[4]/P0001  & n9894 ;
  assign n11013 = \sa23_reg[5]/P0001  & ~n8511 ;
  assign n11014 = n8572 & ~n11013 ;
  assign n11018 = ~n9943 & ~n11014 ;
  assign n11019 = ~n11012 & n11018 ;
  assign n11020 = ~n11017 & n11019 ;
  assign n11021 = ~\sa23_reg[1]/P0001  & ~n11020 ;
  assign n11000 = ~n8521 & ~n9489 ;
  assign n11001 = \sa23_reg[1]/P0001  & ~n11000 ;
  assign n11002 = ~n8525 & ~n8577 ;
  assign n11003 = \sa23_reg[3]/P0001  & ~n11002 ;
  assign n11004 = ~n9899 & ~n9938 ;
  assign n11005 = ~n11003 & n11004 ;
  assign n11006 = ~n11001 & n11005 ;
  assign n11007 = ~\sa23_reg[2]/P0001  & ~n11006 ;
  assign n11008 = ~n9078 & ~n9498 ;
  assign n11009 = n8634 & n11008 ;
  assign n11010 = \sa23_reg[2]/P0001  & ~n11009 ;
  assign n11011 = \sa23_reg[1]/P0001  & n9152 ;
  assign n11022 = ~n9454 & ~n9492 ;
  assign n11023 = ~n11011 & n11022 ;
  assign n11024 = ~n11010 & n11023 ;
  assign n11025 = ~n11007 & n11024 ;
  assign n11026 = ~n11021 & n11025 ;
  assign n11027 = \sa23_reg[0]/P0001  & ~n11026 ;
  assign n11049 = ~n8574 & ~n8642 ;
  assign n11050 = ~n10730 & n11049 ;
  assign n11051 = ~\sa23_reg[7]/NET0131  & ~n11050 ;
  assign n11052 = ~n9464 & ~n11051 ;
  assign n11053 = ~\sa23_reg[2]/P0001  & ~n11052 ;
  assign n11054 = ~n8521 & ~n8654 ;
  assign n11055 = \sa23_reg[2]/P0001  & n8522 ;
  assign n11056 = ~n11054 & n11055 ;
  assign n11057 = ~n8668 & ~n11056 ;
  assign n11058 = ~n11053 & n11057 ;
  assign n11059 = ~\sa23_reg[1]/P0001  & ~n11058 ;
  assign n11034 = ~\sa23_reg[3]/P0001  & ~n9965 ;
  assign n11035 = n9432 & ~n11034 ;
  assign n11038 = n8546 & n8614 ;
  assign n11036 = n8562 & n9079 ;
  assign n11040 = \sa23_reg[1]/P0001  & ~n11036 ;
  assign n11037 = n8569 & n8588 ;
  assign n11039 = n8528 & ~n8537 ;
  assign n11041 = ~n11037 & ~n11039 ;
  assign n11042 = n11040 & n11041 ;
  assign n11043 = ~n11038 & n11042 ;
  assign n11044 = ~n11035 & ~n11043 ;
  assign n11028 = ~n9106 & n10719 ;
  assign n11029 = ~\sa23_reg[2]/P0001  & ~n11028 ;
  assign n11030 = ~n8525 & ~n8631 ;
  assign n11031 = n9897 & ~n11030 ;
  assign n11032 = n8531 & ~n8588 ;
  assign n11033 = n9958 & n11032 ;
  assign n11045 = ~n11031 & ~n11033 ;
  assign n11046 = ~n11029 & n11045 ;
  assign n11047 = ~n11044 & n11046 ;
  assign n11048 = ~\sa23_reg[0]/P0001  & ~n11047 ;
  assign n11061 = ~\sa23_reg[2]/P0001  & ~n8619 ;
  assign n11062 = ~n9438 & ~n11061 ;
  assign n11060 = n9112 & n9152 ;
  assign n11063 = ~n8609 & ~n9137 ;
  assign n11064 = ~n11060 & n11063 ;
  assign n11065 = ~n11062 & n11064 ;
  assign n11066 = \sa23_reg[1]/P0001  & ~n11065 ;
  assign n11067 = \sa23_reg[2]/P0001  & n8524 ;
  assign n11068 = ~\sa23_reg[2]/P0001  & n11037 ;
  assign n11069 = ~n11067 & ~n11068 ;
  assign n11070 = ~n11066 & n11069 ;
  assign n11071 = ~n11048 & n11070 ;
  assign n11072 = ~n11059 & n11071 ;
  assign n11073 = ~n11027 & n11072 ;
  assign n11074 = n10167 & ~n11073 ;
  assign n11075 = ~n10167 & n11073 ;
  assign n11076 = ~n11074 & ~n11075 ;
  assign n11077 = n10999 & n11076 ;
  assign n11078 = ~n10999 & ~n11076 ;
  assign n11079 = ~n11077 & ~n11078 ;
  assign n11126 = ~n8930 & ~n10355 ;
  assign n11127 = \sa30_reg[2]/P0001  & ~n11126 ;
  assign n11122 = \sa30_reg[4]/P0001  & n10272 ;
  assign n11123 = ~n8776 & ~n10255 ;
  assign n11124 = ~n11122 & n11123 ;
  assign n11125 = ~\sa30_reg[2]/P0001  & ~n11124 ;
  assign n11128 = \sa30_reg[1]/P0001  & ~n8703 ;
  assign n11129 = n8761 & n11128 ;
  assign n11130 = ~n11125 & n11129 ;
  assign n11131 = ~n11127 & n11130 ;
  assign n11134 = ~n8876 & ~n8961 ;
  assign n11135 = ~\sa30_reg[2]/P0001  & ~n11134 ;
  assign n11136 = ~\sa30_reg[1]/P0001  & ~n8956 ;
  assign n11132 = n8686 & n8929 ;
  assign n11133 = \sa30_reg[5]/P0001  & n11132 ;
  assign n11137 = ~n9617 & ~n10879 ;
  assign n11138 = ~n11133 & n11137 ;
  assign n11139 = n11136 & n11138 ;
  assign n11140 = ~n11135 & n11139 ;
  assign n11141 = ~n11131 & ~n11140 ;
  assign n11142 = ~n8786 & n9618 ;
  assign n11143 = \sa30_reg[2]/P0001  & ~n8943 ;
  assign n11144 = ~n8951 & n11143 ;
  assign n11145 = ~n11142 & ~n11144 ;
  assign n11146 = ~n8810 & ~n8847 ;
  assign n11147 = ~n11145 & n11146 ;
  assign n11148 = ~n11141 & n11147 ;
  assign n11149 = ~\sa30_reg[0]/P0002  & ~n11148 ;
  assign n11080 = ~n8744 & ~n10821 ;
  assign n11081 = ~n9614 & ~n10375 ;
  assign n11082 = ~n10888 & n11081 ;
  assign n11083 = \sa30_reg[2]/P0001  & ~n11082 ;
  assign n11084 = n11080 & ~n11083 ;
  assign n11085 = \sa30_reg[1]/P0001  & ~n11084 ;
  assign n11094 = n8692 & n8698 ;
  assign n11093 = n8683 & ~n9575 ;
  assign n11095 = ~n8767 & ~n8780 ;
  assign n11096 = ~n11093 & n11095 ;
  assign n11097 = ~n11094 & n11096 ;
  assign n11098 = ~\sa30_reg[1]/P0001  & ~n11097 ;
  assign n11086 = n8710 & ~n9582 ;
  assign n11087 = ~n10351 & ~n11086 ;
  assign n11088 = ~\sa30_reg[3]/P0001  & ~n11087 ;
  assign n11089 = ~n8767 & ~n10279 ;
  assign n11090 = ~n10351 & ~n10363 ;
  assign n11091 = n11089 & n11090 ;
  assign n11092 = ~\sa30_reg[2]/P0001  & ~n11091 ;
  assign n11099 = ~n11088 & ~n11092 ;
  assign n11100 = ~n11098 & n11099 ;
  assign n11101 = ~n11085 & n11100 ;
  assign n11102 = \sa30_reg[0]/P0002  & ~n11101 ;
  assign n11116 = ~n8869 & ~n9632 ;
  assign n11117 = ~n8784 & n11116 ;
  assign n11118 = ~\sa30_reg[2]/P0001  & ~n11117 ;
  assign n11119 = ~n8781 & ~n10864 ;
  assign n11120 = ~n11118 & n11119 ;
  assign n11121 = ~\sa30_reg[1]/P0001  & ~n11120 ;
  assign n11111 = ~n8703 & ~n8883 ;
  assign n11112 = ~n9565 & n11111 ;
  assign n11113 = ~n8749 & ~n8894 ;
  assign n11114 = n11112 & n11113 ;
  assign n11115 = n8772 & ~n11114 ;
  assign n11108 = ~n8769 & ~n8810 ;
  assign n11109 = ~n10256 & n11108 ;
  assign n11110 = n10294 & ~n11109 ;
  assign n11103 = n8710 & ~n9621 ;
  assign n11104 = ~n8821 & ~n11103 ;
  assign n11105 = n8946 & ~n11104 ;
  assign n11106 = ~n8749 & ~n9572 ;
  assign n11107 = n8844 & ~n11106 ;
  assign n11150 = ~n11105 & ~n11107 ;
  assign n11151 = ~n11110 & n11150 ;
  assign n11152 = ~n11115 & n11151 ;
  assign n11153 = ~n11121 & n11152 ;
  assign n11154 = ~n11102 & n11153 ;
  assign n11155 = ~n11149 & n11154 ;
  assign n11156 = ~\u0_w_reg[1][17]/P0001  & ~n11155 ;
  assign n11157 = \u0_w_reg[1][17]/P0001  & n11155 ;
  assign n11158 = ~n11156 & ~n11157 ;
  assign n11159 = n9980 & ~n10508 ;
  assign n11160 = ~n9980 & n10508 ;
  assign n11161 = ~n11159 & ~n11160 ;
  assign n11162 = n11158 & n11161 ;
  assign n11163 = ~n11158 & ~n11161 ;
  assign n11164 = ~n11162 & ~n11163 ;
  assign n11166 = n11079 & n11164 ;
  assign n11165 = ~n11079 & ~n11164 ;
  assign n11167 = ~\ld_r_reg/P0001  & ~n11165 ;
  assign n11168 = ~n11166 & n11167 ;
  assign n11170 = \text_in_r_reg[81]/P0001  & \u0_w_reg[1][17]/P0001  ;
  assign n11169 = ~\text_in_r_reg[81]/P0001  & ~\u0_w_reg[1][17]/P0001  ;
  assign n11171 = \ld_r_reg/P0001  & ~n11169 ;
  assign n11172 = ~n11170 & n11171 ;
  assign n11173 = ~n11168 & ~n11172 ;
  assign n11220 = ~n8138 & ~n9817 ;
  assign n11221 = \sa12_reg[2]/P0001  & ~n11220 ;
  assign n11222 = ~n9035 & ~n11221 ;
  assign n11223 = \sa12_reg[1]/P0001  & ~n11222 ;
  assign n11228 = ~n8075 & ~n8498 ;
  assign n11229 = \sa12_reg[1]/P0001  & ~n8074 ;
  assign n11230 = ~n11228 & n11229 ;
  assign n11231 = ~n8150 & ~n11230 ;
  assign n11232 = ~\sa12_reg[2]/P0001  & ~n11231 ;
  assign n11224 = ~n9865 & ~n10984 ;
  assign n11225 = ~\sa12_reg[1]/P0001  & ~n11224 ;
  assign n11226 = ~n8185 & ~n10660 ;
  assign n11227 = \sa12_reg[4]/P0001  & ~n11226 ;
  assign n11233 = ~n11225 & ~n11227 ;
  assign n11234 = ~n11232 & n11233 ;
  assign n11235 = ~n11223 & n11234 ;
  assign n11236 = ~\sa12_reg[0]/P0001  & ~n11235 ;
  assign n11174 = n10031 & n10920 ;
  assign n11175 = \sa12_reg[1]/P0001  & ~n9837 ;
  assign n11176 = ~n10985 & n11175 ;
  assign n11177 = ~n11174 & n11176 ;
  assign n11179 = n8162 & n9817 ;
  assign n11184 = ~n8189 & ~n8453 ;
  assign n11185 = ~n11179 & n11184 ;
  assign n11180 = ~\sa12_reg[1]/P0001  & ~n8145 ;
  assign n11178 = n8059 & n8060 ;
  assign n11181 = ~n10936 & ~n11178 ;
  assign n11182 = n11180 & n11181 ;
  assign n11183 = ~n8087 & ~n8160 ;
  assign n11186 = n11182 & n11183 ;
  assign n11187 = n11185 & n11186 ;
  assign n11188 = ~n11177 & ~n11187 ;
  assign n11189 = ~n8130 & ~n9049 ;
  assign n11190 = ~n8490 & n11189 ;
  assign n11191 = n8057 & ~n11190 ;
  assign n11192 = ~n8086 & ~n8105 ;
  assign n11193 = ~n10974 & n11192 ;
  assign n11194 = ~n11191 & n11193 ;
  assign n11195 = ~n11188 & n11194 ;
  assign n11196 = \sa12_reg[0]/P0001  & ~n11195 ;
  assign n11199 = ~n9047 & ~n9790 ;
  assign n11200 = ~n8103 & n11199 ;
  assign n11201 = n8997 & n11200 ;
  assign n11202 = \sa12_reg[2]/P0001  & ~n8497 ;
  assign n11203 = ~n9865 & n11202 ;
  assign n11204 = ~n8098 & n11203 ;
  assign n11205 = ~n11201 & ~n11204 ;
  assign n11197 = n8082 & ~n8094 ;
  assign n11198 = ~n8498 & n11197 ;
  assign n11206 = ~\sa12_reg[1]/P0001  & ~n11198 ;
  assign n11207 = ~n11205 & n11206 ;
  assign n11208 = ~n8084 & ~n9042 ;
  assign n11209 = ~\sa12_reg[4]/P0001  & ~n11208 ;
  assign n11210 = \sa12_reg[2]/P0001  & ~n8452 ;
  assign n11211 = ~n11209 & n11210 ;
  assign n11212 = ~\sa12_reg[2]/P0001  & ~n8405 ;
  assign n11213 = n9997 & n11212 ;
  assign n11214 = ~n11211 & ~n11213 ;
  assign n11215 = \sa12_reg[1]/P0001  & ~n8096 ;
  assign n11216 = ~n11214 & n11215 ;
  assign n11217 = ~n11207 & ~n11216 ;
  assign n11218 = ~n8056 & ~n8135 ;
  assign n11219 = n8447 & ~n11218 ;
  assign n11237 = ~n10672 & ~n11219 ;
  assign n11238 = ~n11217 & n11237 ;
  assign n11239 = ~n11196 & n11238 ;
  assign n11240 = ~n11236 & n11239 ;
  assign n11245 = ~n8223 & ~n10185 ;
  assign n11246 = n8237 & n11245 ;
  assign n11243 = ~\sa01_reg[5]/P0001  & ~n8246 ;
  assign n11244 = n8339 & ~n11243 ;
  assign n11241 = \sa01_reg[2]/P0001  & n8276 ;
  assign n11242 = ~n8318 & n11241 ;
  assign n11247 = ~n8312 & ~n11242 ;
  assign n11248 = ~n11244 & n11247 ;
  assign n11249 = n11246 & n11248 ;
  assign n11250 = ~n8242 & ~n8264 ;
  assign n11251 = n9209 & n11250 ;
  assign n11252 = \sa01_reg[1]/P0001  & ~n9208 ;
  assign n11253 = ~n11251 & n11252 ;
  assign n11254 = ~n10229 & n11253 ;
  assign n11255 = ~n11249 & ~n11254 ;
  assign n11256 = ~n8278 & ~n8309 ;
  assign n11257 = ~n8283 & n11256 ;
  assign n11258 = ~\sa01_reg[3]/P0001  & ~n11257 ;
  assign n11259 = ~n8258 & ~n9276 ;
  assign n11260 = ~n9368 & n11259 ;
  assign n11261 = n8329 & ~n11260 ;
  assign n11262 = ~n11258 & ~n11261 ;
  assign n11263 = ~n11255 & n11262 ;
  assign n11264 = \sa01_reg[0]/P0001  & ~n11263 ;
  assign n11265 = ~n9196 & n10084 ;
  assign n11266 = ~\sa01_reg[2]/P0001  & ~n11265 ;
  assign n11267 = ~n8352 & ~n11266 ;
  assign n11268 = \sa01_reg[1]/P0001  & ~n11267 ;
  assign n11269 = ~n8320 & ~n9268 ;
  assign n11270 = n9388 & ~n11269 ;
  assign n11273 = ~n8219 & ~n8254 ;
  assign n11274 = n10230 & ~n11273 ;
  assign n11271 = \sa01_reg[1]/P0001  & n8329 ;
  assign n11272 = n8369 & n11271 ;
  assign n11306 = ~n10581 & ~n11272 ;
  assign n11307 = ~n11274 & n11306 ;
  assign n11308 = ~n11270 & n11307 ;
  assign n11309 = ~n11268 & n11308 ;
  assign n11275 = ~n8227 & ~n9373 ;
  assign n11276 = \sa01_reg[3]/P0001  & ~n11275 ;
  assign n11277 = ~n9774 & ~n11276 ;
  assign n11278 = \sa01_reg[2]/P0001  & ~n11277 ;
  assign n11281 = ~n8309 & ~n9375 ;
  assign n11282 = ~n8361 & n11281 ;
  assign n11283 = ~\sa01_reg[2]/P0001  & ~n11282 ;
  assign n11279 = ~n8214 & n8227 ;
  assign n11280 = ~n8265 & n11279 ;
  assign n11284 = ~n9305 & ~n11280 ;
  assign n11285 = ~n11283 & n11284 ;
  assign n11286 = ~n11278 & n11285 ;
  assign n11287 = ~\sa01_reg[1]/P0001  & ~n11286 ;
  assign n11288 = ~n8266 & ~n8339 ;
  assign n11289 = \sa01_reg[2]/P0001  & ~n11288 ;
  assign n11290 = ~n8264 & ~n8265 ;
  assign n11291 = ~\sa01_reg[2]/P0001  & ~n8342 ;
  assign n11292 = ~n11290 & n11291 ;
  assign n11293 = ~n9369 & ~n11292 ;
  assign n11294 = ~n11289 & n11293 ;
  assign n11295 = \sa01_reg[1]/P0001  & ~n11294 ;
  assign n11296 = \sa01_reg[2]/P0001  & n8332 ;
  assign n11301 = ~n8243 & ~n11296 ;
  assign n11297 = n8342 & n9386 ;
  assign n11298 = ~n9774 & ~n11297 ;
  assign n11299 = ~\sa01_reg[1]/P0001  & ~n11298 ;
  assign n11300 = ~\sa01_reg[2]/P0001  & n8220 ;
  assign n11302 = ~n11299 & ~n11300 ;
  assign n11303 = n11301 & n11302 ;
  assign n11304 = ~n11295 & n11303 ;
  assign n11305 = ~\sa01_reg[0]/P0001  & ~n11304 ;
  assign n11310 = ~n11287 & ~n11305 ;
  assign n11311 = n11309 & n11310 ;
  assign n11312 = ~n11264 & n11311 ;
  assign n11313 = n11240 & ~n11312 ;
  assign n11314 = ~n11240 & n11312 ;
  assign n11315 = ~n11313 & ~n11314 ;
  assign n11316 = ~n10167 & ~n11315 ;
  assign n11317 = n10167 & n11315 ;
  assign n11318 = ~n11316 & ~n11317 ;
  assign n11327 = ~n8653 & ~n8667 ;
  assign n11328 = ~n9152 & n11327 ;
  assign n11329 = \sa23_reg[3]/P0001  & ~n11328 ;
  assign n11330 = ~n9492 & ~n11329 ;
  assign n11331 = \sa23_reg[2]/P0001  & ~n11330 ;
  assign n11319 = ~n8602 & n10477 ;
  assign n11320 = ~n9497 & ~n11319 ;
  assign n11321 = ~n9419 & ~n9430 ;
  assign n11322 = ~n9451 & ~n9943 ;
  assign n11323 = n11321 & n11322 ;
  assign n11324 = ~n9064 & n11323 ;
  assign n11325 = ~n11320 & n11324 ;
  assign n11326 = ~\sa23_reg[1]/P0001  & ~n11325 ;
  assign n11333 = ~\sa23_reg[2]/P0001  & ~n8574 ;
  assign n11334 = ~n9099 & n11333 ;
  assign n11335 = ~n8647 & n11334 ;
  assign n11332 = \sa23_reg[2]/P0001  & ~n8578 ;
  assign n11336 = \sa23_reg[1]/P0001  & ~n11332 ;
  assign n11337 = ~n11335 & n11336 ;
  assign n11338 = ~n9464 & ~n9469 ;
  assign n11339 = ~n11337 & n11338 ;
  assign n11340 = ~n11326 & n11339 ;
  assign n11341 = ~n11331 & n11340 ;
  assign n11342 = \sa23_reg[0]/P0001  & ~n11341 ;
  assign n11343 = ~n9159 & ~n9482 ;
  assign n11344 = ~n9064 & n11343 ;
  assign n11345 = n9474 & n11344 ;
  assign n11346 = \sa23_reg[3]/P0001  & n8547 ;
  assign n11347 = ~n9476 & ~n11346 ;
  assign n11348 = n9953 & n11347 ;
  assign n11349 = ~n11345 & ~n11348 ;
  assign n11350 = n8547 & ~n8573 ;
  assign n11351 = ~n8577 & n11350 ;
  assign n11352 = ~n11349 & ~n11351 ;
  assign n11353 = ~\sa23_reg[1]/P0001  & ~n11352 ;
  assign n11373 = ~n8562 & ~n8631 ;
  assign n11374 = n8522 & ~n11373 ;
  assign n11375 = ~n8602 & ~n8603 ;
  assign n11376 = ~n9462 & n11375 ;
  assign n11377 = \sa23_reg[1]/P0001  & ~n11376 ;
  assign n11378 = ~n11374 & ~n11377 ;
  assign n11379 = \sa23_reg[2]/P0001  & ~n11378 ;
  assign n11380 = ~n10729 & ~n11379 ;
  assign n11381 = ~n11353 & n11380 ;
  assign n11354 = ~n8552 & ~n8591 ;
  assign n11355 = \sa23_reg[2]/P0001  & ~n11354 ;
  assign n11356 = ~n8577 & ~n8588 ;
  assign n11357 = ~\sa23_reg[2]/P0001  & ~n8589 ;
  assign n11358 = ~n11356 & n11357 ;
  assign n11359 = ~n9154 & ~n11358 ;
  assign n11360 = ~n11355 & n11359 ;
  assign n11361 = \sa23_reg[1]/P0001  & ~n11360 ;
  assign n11362 = ~n8620 & n9954 ;
  assign n11363 = n8546 & n8602 ;
  assign n11364 = ~n8570 & ~n11363 ;
  assign n11365 = ~n9135 & n11364 ;
  assign n11366 = ~n11362 & n11365 ;
  assign n11367 = ~n11361 & n11366 ;
  assign n11368 = ~\sa23_reg[0]/P0001  & ~n11367 ;
  assign n11369 = ~n8551 & n10443 ;
  assign n11370 = ~\sa23_reg[2]/P0001  & ~n11369 ;
  assign n11371 = ~n8527 & ~n11370 ;
  assign n11372 = \sa23_reg[1]/P0001  & ~n11371 ;
  assign n11382 = ~n11368 & ~n11372 ;
  assign n11383 = n11381 & n11382 ;
  assign n11384 = ~n11342 & n11383 ;
  assign n11385 = \u0_w_reg[1][2]/P0001  & ~n11384 ;
  assign n11386 = ~\u0_w_reg[1][2]/P0001  & n11384 ;
  assign n11387 = ~n11385 & ~n11386 ;
  assign n11388 = n11155 & n11387 ;
  assign n11389 = ~n11155 & ~n11387 ;
  assign n11390 = ~n11388 & ~n11389 ;
  assign n11392 = n11318 & ~n11390 ;
  assign n11391 = ~n11318 & n11390 ;
  assign n11393 = ~\ld_r_reg/P0001  & ~n11391 ;
  assign n11394 = ~n11392 & n11393 ;
  assign n11396 = \text_in_r_reg[66]/P0001  & \u0_w_reg[1][2]/P0001  ;
  assign n11395 = ~\text_in_r_reg[66]/P0001  & ~\u0_w_reg[1][2]/P0001  ;
  assign n11397 = \ld_r_reg/P0001  & ~n11395 ;
  assign n11398 = ~n11396 & n11397 ;
  assign n11399 = ~n11394 & ~n11398 ;
  assign n11400 = n10081 & ~n10508 ;
  assign n11401 = ~n10081 & n10508 ;
  assign n11402 = ~n11400 & ~n11401 ;
  assign n11403 = \u0_w_reg[1][25]/P0001  & ~n11155 ;
  assign n11404 = ~\u0_w_reg[1][25]/P0001  & n11155 ;
  assign n11405 = ~n11403 & ~n11404 ;
  assign n11406 = n11402 & n11405 ;
  assign n11407 = ~n11402 & ~n11405 ;
  assign n11408 = ~n11406 & ~n11407 ;
  assign n11409 = n10251 & n10999 ;
  assign n11410 = ~n10251 & ~n10999 ;
  assign n11411 = ~n11409 & ~n11410 ;
  assign n11413 = n11408 & n11411 ;
  assign n11412 = ~n11408 & ~n11411 ;
  assign n11414 = ~\ld_r_reg/P0001  & ~n11412 ;
  assign n11415 = ~n11413 & n11414 ;
  assign n11417 = \text_in_r_reg[89]/P0001  & \u0_w_reg[1][25]/P0001  ;
  assign n11416 = ~\text_in_r_reg[89]/P0001  & ~\u0_w_reg[1][25]/P0001  ;
  assign n11418 = \ld_r_reg/P0001  & ~n11416 ;
  assign n11419 = ~n11417 & n11418 ;
  assign n11420 = ~n11415 & ~n11419 ;
  assign n11421 = ~n9169 & ~n9877 ;
  assign n11422 = n9169 & n9877 ;
  assign n11423 = ~n11421 & ~n11422 ;
  assign n11424 = \u0_w_reg[1][15]/P0001  & ~n10430 ;
  assign n11425 = ~\u0_w_reg[1][15]/P0001  & n10430 ;
  assign n11426 = ~n11424 & ~n11425 ;
  assign n11427 = n8974 & n11426 ;
  assign n11428 = ~n8974 & ~n11426 ;
  assign n11429 = ~n11427 & ~n11428 ;
  assign n11431 = n11423 & ~n11429 ;
  assign n11430 = ~n11423 & n11429 ;
  assign n11432 = ~\ld_r_reg/P0001  & ~n11430 ;
  assign n11433 = ~n11431 & n11432 ;
  assign n11435 = ~\text_in_r_reg[79]/P0001  & \u0_w_reg[1][15]/P0001  ;
  assign n11434 = \text_in_r_reg[79]/P0001  & ~\u0_w_reg[1][15]/P0001  ;
  assign n11436 = \ld_r_reg/P0001  & ~n11434 ;
  assign n11437 = ~n11435 & n11436 ;
  assign n11438 = ~n11433 & ~n11437 ;
  assign n11439 = ~\u0_w_reg[1][27]/P0001  & ~n10898 ;
  assign n11440 = \u0_w_reg[1][27]/P0001  & n10898 ;
  assign n11441 = ~n11439 & ~n11440 ;
  assign n11442 = n10682 & ~n10775 ;
  assign n11443 = ~n10682 & n10775 ;
  assign n11444 = ~n11442 & ~n11443 ;
  assign n11445 = n11441 & n11444 ;
  assign n11446 = ~n11441 & ~n11444 ;
  assign n11447 = ~n11445 & ~n11446 ;
  assign n11448 = n9783 & ~n11312 ;
  assign n11449 = ~n9783 & n11312 ;
  assign n11450 = ~n11448 & ~n11449 ;
  assign n11451 = n9874 & ~n11240 ;
  assign n11452 = ~n9874 & n11240 ;
  assign n11453 = ~n11451 & ~n11452 ;
  assign n11454 = n11450 & ~n11453 ;
  assign n11455 = ~n11450 & n11453 ;
  assign n11456 = ~n11454 & ~n11455 ;
  assign n11458 = n11447 & n11456 ;
  assign n11457 = ~n11447 & ~n11456 ;
  assign n11459 = ~\ld_r_reg/P0001  & ~n11457 ;
  assign n11460 = ~n11458 & n11459 ;
  assign n11462 = ~\text_in_r_reg[91]/P0001  & \u0_w_reg[1][27]/P0001  ;
  assign n11461 = \text_in_r_reg[91]/P0001  & ~\u0_w_reg[1][27]/P0001  ;
  assign n11463 = \ld_r_reg/P0001  & ~n11461 ;
  assign n11464 = ~n11462 & n11463 ;
  assign n11465 = ~n11460 & ~n11464 ;
  assign n11466 = \u0_w_reg[1][19]/P0001  & ~n10898 ;
  assign n11467 = ~\u0_w_reg[1][19]/P0001  & n10898 ;
  assign n11468 = ~n11466 & ~n11467 ;
  assign n11469 = n10907 & n11468 ;
  assign n11470 = ~n10907 & ~n11468 ;
  assign n11471 = ~n11469 & ~n11470 ;
  assign n11472 = n10602 & ~n11384 ;
  assign n11473 = ~n10602 & n11384 ;
  assign n11474 = ~n11472 & ~n11473 ;
  assign n11475 = n11453 & n11474 ;
  assign n11476 = ~n11453 & ~n11474 ;
  assign n11477 = ~n11475 & ~n11476 ;
  assign n11479 = n11471 & n11477 ;
  assign n11478 = ~n11471 & ~n11477 ;
  assign n11480 = ~\ld_r_reg/P0001  & ~n11478 ;
  assign n11481 = ~n11479 & n11480 ;
  assign n11483 = ~\text_in_r_reg[83]/P0001  & \u0_w_reg[1][19]/P0001  ;
  assign n11482 = \text_in_r_reg[83]/P0001  & ~\u0_w_reg[1][19]/P0001  ;
  assign n11484 = \ld_r_reg/P0001  & ~n11482 ;
  assign n11485 = ~n11483 & n11484 ;
  assign n11486 = ~n11481 & ~n11485 ;
  assign n11487 = n10602 & ~n10682 ;
  assign n11488 = ~n10602 & n10682 ;
  assign n11489 = ~n11487 & ~n11488 ;
  assign n11490 = n9980 & ~n11384 ;
  assign n11491 = ~n9980 & n11384 ;
  assign n11492 = ~n11490 & ~n11491 ;
  assign n11493 = n11489 & n11492 ;
  assign n11494 = ~n11489 & ~n11492 ;
  assign n11495 = ~n11493 & ~n11494 ;
  assign n11500 = ~n8758 & n10372 ;
  assign n11499 = \sa30_reg[2]/P0001  & n8733 ;
  assign n11501 = \sa30_reg[1]/P0001  & ~n11499 ;
  assign n11502 = ~n11500 & n11501 ;
  assign n11503 = ~n10332 & n11502 ;
  assign n11507 = ~n8765 & ~n8894 ;
  assign n11504 = n8724 & n9582 ;
  assign n11508 = ~n9546 & ~n11504 ;
  assign n11509 = n11507 & n11508 ;
  assign n11505 = ~n9576 & ~n10263 ;
  assign n11506 = ~n11132 & n11505 ;
  assign n11510 = n9587 & n11506 ;
  assign n11511 = n11509 & n11510 ;
  assign n11512 = ~n11503 & ~n11511 ;
  assign n11496 = ~n8816 & ~n8961 ;
  assign n11497 = ~n10351 & n11496 ;
  assign n11498 = n8844 & ~n11497 ;
  assign n11513 = \sa30_reg[0]/P0002  & ~n9566 ;
  assign n11514 = ~n10333 & ~n11133 ;
  assign n11515 = n11513 & n11514 ;
  assign n11516 = ~n11498 & n11515 ;
  assign n11517 = ~n11512 & n11516 ;
  assign n11518 = n8756 & n8940 ;
  assign n11519 = ~\sa30_reg[1]/P0001  & ~n8785 ;
  assign n11520 = ~n11518 & n11519 ;
  assign n11521 = \sa30_reg[2]/P0001  & ~n8724 ;
  assign n11522 = ~n8760 & n11521 ;
  assign n11523 = ~n8756 & n8758 ;
  assign n11524 = ~\sa30_reg[2]/P0001  & ~n8748 ;
  assign n11525 = ~n11523 & n11524 ;
  assign n11526 = ~n11522 & ~n11525 ;
  assign n11527 = \sa30_reg[1]/P0001  & ~n10363 ;
  assign n11528 = ~n11526 & n11527 ;
  assign n11529 = ~n11520 & ~n11528 ;
  assign n11530 = n8811 & n9596 ;
  assign n11531 = ~\sa30_reg[0]/P0002  & ~n8899 ;
  assign n11532 = ~n11530 & n11531 ;
  assign n11533 = ~n8832 & n11532 ;
  assign n11534 = ~n11529 & n11533 ;
  assign n11535 = ~n11517 & ~n11534 ;
  assign n11539 = ~n8775 & ~n8952 ;
  assign n11540 = \sa30_reg[3]/P0001  & ~n11539 ;
  assign n11541 = n10413 & ~n11540 ;
  assign n11542 = ~\sa30_reg[2]/P0001  & ~n8964 ;
  assign n11543 = ~n8822 & n11542 ;
  assign n11544 = ~n8894 & ~n10418 ;
  assign n11545 = n11543 & n11544 ;
  assign n11546 = ~n11541 & ~n11545 ;
  assign n11547 = n8695 & n8775 ;
  assign n11548 = ~\sa30_reg[1]/P0001  & ~n11547 ;
  assign n11549 = ~n9543 & n11548 ;
  assign n11550 = ~n11546 & n11549 ;
  assign n11551 = n8723 & n11080 ;
  assign n11552 = n8792 & n8838 ;
  assign n11553 = \sa30_reg[2]/P0001  & ~n8719 ;
  assign n11554 = ~n8823 & n11553 ;
  assign n11555 = ~n11552 & n11554 ;
  assign n11556 = ~n11551 & ~n11555 ;
  assign n11557 = \sa30_reg[1]/P0001  & ~n8711 ;
  assign n11558 = ~n11556 & n11557 ;
  assign n11559 = ~n11550 & ~n11558 ;
  assign n11536 = ~n8845 & ~n8874 ;
  assign n11537 = ~\sa30_reg[3]/P0001  & n9575 ;
  assign n11538 = ~n11536 & n11537 ;
  assign n11560 = ~n10875 & ~n11538 ;
  assign n11561 = ~n11559 & n11560 ;
  assign n11562 = ~n11535 & n11561 ;
  assign n11563 = n10430 & ~n11562 ;
  assign n11564 = ~n10430 & n11562 ;
  assign n11565 = ~n11563 & ~n11564 ;
  assign n11566 = \u0_w_reg[1][11]/P0001  & ~n10898 ;
  assign n11567 = ~\u0_w_reg[1][11]/P0001  & n10898 ;
  assign n11568 = ~n11566 & ~n11567 ;
  assign n11569 = n11565 & n11568 ;
  assign n11570 = ~n11565 & ~n11568 ;
  assign n11571 = ~n11569 & ~n11570 ;
  assign n11573 = n11495 & n11571 ;
  assign n11572 = ~n11495 & ~n11571 ;
  assign n11574 = ~\ld_r_reg/P0001  & ~n11572 ;
  assign n11575 = ~n11573 & n11574 ;
  assign n11577 = ~\text_in_r_reg[75]/P0001  & \u0_w_reg[1][11]/P0001  ;
  assign n11576 = \text_in_r_reg[75]/P0001  & ~\u0_w_reg[1][11]/P0001  ;
  assign n11578 = \ld_r_reg/P0001  & ~n11576 ;
  assign n11579 = ~n11577 & n11578 ;
  assign n11580 = ~n11575 & ~n11579 ;
  assign n11581 = ~n9516 & ~n10430 ;
  assign n11582 = n9516 & n10430 ;
  assign n11583 = ~n11581 & ~n11582 ;
  assign n11584 = \u0_w_reg[1][4]/P0001  & ~n10898 ;
  assign n11585 = ~\u0_w_reg[1][4]/P0001  & n10898 ;
  assign n11586 = ~n11584 & ~n11585 ;
  assign n11587 = n11583 & n11586 ;
  assign n11588 = ~n11583 & ~n11586 ;
  assign n11589 = ~n11587 & ~n11588 ;
  assign n11590 = ~n8379 & n10605 ;
  assign n11591 = n8379 & ~n10605 ;
  assign n11592 = ~n11590 & ~n11591 ;
  assign n11594 = n11589 & n11592 ;
  assign n11593 = ~n11589 & ~n11592 ;
  assign n11595 = ~\ld_r_reg/P0001  & ~n11593 ;
  assign n11596 = ~n11594 & n11595 ;
  assign n11598 = ~\text_in_r_reg[68]/P0001  & \u0_w_reg[1][4]/P0001  ;
  assign n11597 = \text_in_r_reg[68]/P0001  & ~\u0_w_reg[1][4]/P0001  ;
  assign n11599 = \ld_r_reg/P0001  & ~n11597 ;
  assign n11600 = ~n11598 & n11599 ;
  assign n11601 = ~n11596 & ~n11600 ;
  assign n11602 = ~\u0_w_reg[1][26]/P0001  & ~n11562 ;
  assign n11603 = \u0_w_reg[1][26]/P0001  & n11562 ;
  assign n11604 = ~n11602 & ~n11603 ;
  assign n11605 = ~n11240 & n11384 ;
  assign n11606 = n11240 & ~n11384 ;
  assign n11607 = ~n11605 & ~n11606 ;
  assign n11608 = n11604 & n11607 ;
  assign n11609 = ~n11604 & ~n11607 ;
  assign n11610 = ~n11608 & ~n11609 ;
  assign n11612 = n10170 & n11610 ;
  assign n11611 = ~n10170 & ~n11610 ;
  assign n11613 = ~\ld_r_reg/P0001  & ~n11611 ;
  assign n11614 = ~n11612 & n11613 ;
  assign n11616 = \text_in_r_reg[90]/P0001  & \u0_w_reg[1][26]/P0001  ;
  assign n11615 = ~\text_in_r_reg[90]/P0001  & ~\u0_w_reg[1][26]/P0001  ;
  assign n11617 = \ld_r_reg/P0001  & ~n11615 ;
  assign n11618 = ~n11616 & n11617 ;
  assign n11619 = ~n11614 & ~n11618 ;
  assign n11620 = \u0_w_reg[1][31]/P0001  & ~n10430 ;
  assign n11621 = ~\u0_w_reg[1][31]/P0001  & n10430 ;
  assign n11622 = ~n11620 & ~n11621 ;
  assign n11623 = ~n9874 & n9980 ;
  assign n11624 = n9874 & ~n9980 ;
  assign n11625 = ~n11623 & ~n11624 ;
  assign n11626 = n9657 & n11625 ;
  assign n11627 = ~n9657 & ~n11625 ;
  assign n11628 = ~n11626 & ~n11627 ;
  assign n11630 = n11622 & ~n11628 ;
  assign n11629 = ~n11622 & n11628 ;
  assign n11631 = ~\ld_r_reg/P0001  & ~n11629 ;
  assign n11632 = ~n11630 & n11631 ;
  assign n11634 = ~\text_in_r_reg[95]/P0001  & \u0_w_reg[1][31]/P0001  ;
  assign n11633 = \text_in_r_reg[95]/P0001  & ~\u0_w_reg[1][31]/P0001  ;
  assign n11635 = \ld_r_reg/P0001  & ~n11633 ;
  assign n11636 = ~n11634 & n11635 ;
  assign n11637 = ~n11632 & ~n11636 ;
  assign n11638 = ~\u0_w_reg[1][16]/P0001  & ~n10344 ;
  assign n11639 = \u0_w_reg[1][16]/P0001  & n10344 ;
  assign n11640 = ~n11638 & ~n11639 ;
  assign n11641 = n9980 & ~n11073 ;
  assign n11642 = ~n9980 & n11073 ;
  assign n11643 = ~n11641 & ~n11642 ;
  assign n11644 = n9874 & ~n10248 ;
  assign n11645 = ~n9874 & n10248 ;
  assign n11646 = ~n11644 & ~n11645 ;
  assign n11647 = n11643 & n11646 ;
  assign n11648 = ~n11643 & ~n11646 ;
  assign n11649 = ~n11647 & ~n11648 ;
  assign n11651 = n11640 & ~n11649 ;
  assign n11650 = ~n11640 & n11649 ;
  assign n11652 = ~\ld_r_reg/P0001  & ~n11650 ;
  assign n11653 = ~n11651 & n11652 ;
  assign n11655 = \text_in_r_reg[80]/P0001  & \u0_w_reg[1][16]/P0001  ;
  assign n11654 = ~\text_in_r_reg[80]/P0001  & ~\u0_w_reg[1][16]/P0001  ;
  assign n11656 = \ld_r_reg/P0001  & ~n11654 ;
  assign n11657 = ~n11655 & n11656 ;
  assign n11658 = ~n11653 & ~n11657 ;
  assign n11659 = ~n11312 & ~n11402 ;
  assign n11660 = n11312 & n11402 ;
  assign n11661 = ~n11659 & ~n11660 ;
  assign n11662 = \u0_w_reg[1][18]/P0001  & ~n11562 ;
  assign n11663 = ~\u0_w_reg[1][18]/P0001  & n11562 ;
  assign n11664 = ~n11662 & ~n11663 ;
  assign n11665 = n11384 & n11664 ;
  assign n11666 = ~n11384 & ~n11664 ;
  assign n11667 = ~n11665 & ~n11666 ;
  assign n11669 = n11661 & n11667 ;
  assign n11668 = ~n11661 & ~n11667 ;
  assign n11670 = ~\ld_r_reg/P0001  & ~n11668 ;
  assign n11671 = ~n11669 & n11670 ;
  assign n11673 = ~\text_in_r_reg[82]/P0001  & \u0_w_reg[1][18]/P0001  ;
  assign n11672 = \text_in_r_reg[82]/P0001  & ~\u0_w_reg[1][18]/P0001  ;
  assign n11674 = \ld_r_reg/P0001  & ~n11672 ;
  assign n11675 = ~n11673 & n11674 ;
  assign n11676 = ~n11671 & ~n11675 ;
  assign n11677 = ~n9172 & ~n9783 ;
  assign n11678 = n9172 & n9783 ;
  assign n11679 = ~n11677 & ~n11678 ;
  assign n11680 = n9980 & ~n10430 ;
  assign n11681 = ~n9980 & n10430 ;
  assign n11682 = ~n11680 & ~n11681 ;
  assign n11683 = ~\u0_w_reg[1][23]/P0001  & ~n11682 ;
  assign n11684 = \u0_w_reg[1][23]/P0001  & n11682 ;
  assign n11685 = ~n11683 & ~n11684 ;
  assign n11687 = n11679 & n11685 ;
  assign n11686 = ~n11679 & ~n11685 ;
  assign n11688 = ~\ld_r_reg/P0001  & ~n11686 ;
  assign n11689 = ~n11687 & n11688 ;
  assign n11691 = ~\text_in_r_reg[87]/P0001  & \u0_w_reg[1][23]/P0001  ;
  assign n11690 = \text_in_r_reg[87]/P0001  & ~\u0_w_reg[1][23]/P0001  ;
  assign n11692 = \ld_r_reg/P0001  & ~n11690 ;
  assign n11693 = ~n11691 & n11692 ;
  assign n11694 = ~n11689 & ~n11693 ;
  assign n11695 = ~\u0_w_reg[1][24]/P0002  & ~n10344 ;
  assign n11696 = \u0_w_reg[1][24]/P0002  & n10344 ;
  assign n11697 = ~n11695 & ~n11696 ;
  assign n11698 = n10996 & ~n11073 ;
  assign n11699 = ~n10996 & n11073 ;
  assign n11700 = ~n11698 & ~n11699 ;
  assign n11701 = n9877 & n11700 ;
  assign n11702 = ~n9877 & ~n11700 ;
  assign n11703 = ~n11701 & ~n11702 ;
  assign n11705 = n11697 & n11703 ;
  assign n11704 = ~n11697 & ~n11703 ;
  assign n11706 = ~\ld_r_reg/P0001  & ~n11704 ;
  assign n11707 = ~n11705 & n11706 ;
  assign n11709 = \text_in_r_reg[88]/P0001  & \u0_w_reg[1][24]/P0002  ;
  assign n11708 = ~\text_in_r_reg[88]/P0001  & ~\u0_w_reg[1][24]/P0002  ;
  assign n11710 = \ld_r_reg/P0001  & ~n11708 ;
  assign n11711 = ~n11709 & n11710 ;
  assign n11712 = ~n11707 & ~n11711 ;
  assign n11713 = ~\u0_w_reg[1][8]/P0001  & ~n10344 ;
  assign n11714 = \u0_w_reg[1][8]/P0001  & n10344 ;
  assign n11715 = ~n11713 & ~n11714 ;
  assign n11716 = n10248 & ~n10996 ;
  assign n11717 = ~n10248 & n10996 ;
  assign n11718 = ~n11716 & ~n11717 ;
  assign n11719 = n11682 & n11718 ;
  assign n11720 = ~n11682 & ~n11718 ;
  assign n11721 = ~n11719 & ~n11720 ;
  assign n11723 = n11715 & n11721 ;
  assign n11722 = ~n11715 & ~n11721 ;
  assign n11724 = ~\ld_r_reg/P0001  & ~n11722 ;
  assign n11725 = ~n11723 & n11724 ;
  assign n11727 = ~\text_in_r_reg[72]/P0001  & \u0_w_reg[1][8]/P0001  ;
  assign n11726 = \text_in_r_reg[72]/P0001  & ~\u0_w_reg[1][8]/P0001  ;
  assign n11728 = \ld_r_reg/P0001  & ~n11726 ;
  assign n11729 = ~n11727 & n11728 ;
  assign n11730 = ~n11725 & ~n11729 ;
  assign n11731 = ~n10508 & ~n11315 ;
  assign n11732 = n10508 & n11315 ;
  assign n11733 = ~n11731 & ~n11732 ;
  assign n11734 = \u0_w_reg[1][10]/P0001  & ~n11562 ;
  assign n11735 = ~\u0_w_reg[1][10]/P0001  & n11562 ;
  assign n11736 = ~n11734 & ~n11735 ;
  assign n11737 = n11155 & n11736 ;
  assign n11738 = ~n11155 & ~n11736 ;
  assign n11739 = ~n11737 & ~n11738 ;
  assign n11741 = n11733 & n11739 ;
  assign n11740 = ~n11733 & ~n11739 ;
  assign n11742 = ~\ld_r_reg/P0001  & ~n11740 ;
  assign n11743 = ~n11741 & n11742 ;
  assign n11745 = ~\text_in_r_reg[74]/P0001  & \u0_w_reg[1][10]/P0001  ;
  assign n11744 = \text_in_r_reg[74]/P0001  & ~\u0_w_reg[1][10]/P0001  ;
  assign n11746 = \ld_r_reg/P0001  & ~n11744 ;
  assign n11747 = ~n11745 & n11746 ;
  assign n11748 = ~n11743 & ~n11747 ;
  assign n11749 = \u0_w_reg[1][3]/P0001  & ~n10775 ;
  assign n11750 = ~\u0_w_reg[1][3]/P0001  & n10775 ;
  assign n11751 = ~n11749 & ~n11750 ;
  assign n11752 = n11565 & n11751 ;
  assign n11753 = ~n11565 & ~n11751 ;
  assign n11754 = ~n11752 & ~n11753 ;
  assign n11755 = n11450 & n11489 ;
  assign n11756 = ~n11450 & ~n11489 ;
  assign n11757 = ~n11755 & ~n11756 ;
  assign n11759 = n11754 & n11757 ;
  assign n11758 = ~n11754 & ~n11757 ;
  assign n11760 = ~\ld_r_reg/P0001  & ~n11758 ;
  assign n11761 = ~n11759 & n11760 ;
  assign n11763 = ~\text_in_r_reg[67]/P0001  & \u0_w_reg[1][3]/P0001  ;
  assign n11762 = \text_in_r_reg[67]/P0001  & ~\u0_w_reg[1][3]/P0001  ;
  assign n11764 = \ld_r_reg/P0001  & ~n11762 ;
  assign n11765 = ~n11763 & n11764 ;
  assign n11766 = ~n11761 & ~n11765 ;
  assign n11767 = ~\u0_w_reg[1][5]/P0001  & ~n8853 ;
  assign n11768 = \u0_w_reg[1][5]/P0001  & n8853 ;
  assign n11769 = ~n11767 & ~n11768 ;
  assign n11770 = ~\u0_w_reg[1][6]/P0001  & ~n8974 ;
  assign n11771 = \u0_w_reg[1][6]/P0001  & n8974 ;
  assign n11772 = ~n11770 & ~n11771 ;
  assign n11773 = ~\u0_w_reg[1][4]/P0001  & ~n9639 ;
  assign n11774 = \u0_w_reg[1][4]/P0001  & n9639 ;
  assign n11775 = ~n11773 & ~n11774 ;
  assign n11776 = ~\u0_w_reg[1][0]/P0001  & ~n10344 ;
  assign n11777 = \u0_w_reg[1][0]/P0001  & n10344 ;
  assign n11778 = ~n11776 & ~n11777 ;
  assign n11779 = ~\u0_w_reg[1][3]/P0001  & ~n10898 ;
  assign n11780 = \u0_w_reg[1][3]/P0001  & n10898 ;
  assign n11781 = ~n11779 & ~n11780 ;
  assign n11782 = ~\u0_w_reg[1][1]/P0001  & ~n11155 ;
  assign n11783 = \u0_w_reg[1][1]/P0001  & n11155 ;
  assign n11784 = ~n11782 & ~n11783 ;
  assign n11785 = ~\u0_w_reg[1][2]/P0001  & ~n11562 ;
  assign n11786 = \u0_w_reg[1][2]/P0001  & n11562 ;
  assign n11787 = ~n11785 & ~n11786 ;
  assign n11788 = ~\u0_w_reg[1][7]/P0001  & ~n10430 ;
  assign n11789 = \u0_w_reg[1][7]/P0001  & n10430 ;
  assign n11790 = ~n11788 & ~n11789 ;
  assign n11796 = \sa11_reg[3]/P0001  & ~\sa11_reg[4]/P0001  ;
  assign n11797 = \sa11_reg[5]/P0001  & ~\sa11_reg[6]/NET0131  ;
  assign n11798 = \sa11_reg[7]/NET0131  & n11797 ;
  assign n11799 = ~n11796 & n11798 ;
  assign n11800 = ~\sa11_reg[4]/P0001  & ~\sa11_reg[6]/NET0131  ;
  assign n11801 = ~\sa11_reg[5]/P0001  & \sa11_reg[7]/NET0131  ;
  assign n11802 = n11800 & n11801 ;
  assign n11803 = ~n11799 & ~n11802 ;
  assign n11804 = ~\sa11_reg[2]/P0001  & ~n11803 ;
  assign n11805 = \sa11_reg[2]/P0001  & ~\sa11_reg[3]/P0001  ;
  assign n11806 = \sa11_reg[4]/P0001  & n11801 ;
  assign n11807 = n11805 & n11806 ;
  assign n11791 = \sa11_reg[6]/NET0131  & ~\sa11_reg[7]/NET0131  ;
  assign n11792 = \sa11_reg[5]/P0001  & n11791 ;
  assign n11793 = \sa11_reg[2]/P0001  & n11792 ;
  assign n11794 = \sa11_reg[3]/P0001  & \sa11_reg[4]/P0001  ;
  assign n11795 = n11791 & n11794 ;
  assign n11808 = ~n11793 & ~n11795 ;
  assign n11809 = ~n11807 & n11808 ;
  assign n11810 = ~n11804 & n11809 ;
  assign n11811 = \sa11_reg[1]/P0001  & ~n11810 ;
  assign n11836 = ~\sa11_reg[3]/P0001  & n11792 ;
  assign n11837 = ~\sa11_reg[2]/P0001  & n11836 ;
  assign n11833 = \sa11_reg[5]/P0001  & \sa11_reg[6]/NET0131  ;
  assign n11834 = \sa11_reg[2]/P0001  & \sa11_reg[4]/P0001  ;
  assign n11835 = n11833 & n11834 ;
  assign n11829 = ~\sa11_reg[6]/NET0131  & ~\sa11_reg[7]/NET0131  ;
  assign n11830 = n11796 & n11829 ;
  assign n11812 = ~\sa11_reg[5]/P0001  & ~\sa11_reg[7]/NET0131  ;
  assign n11831 = \sa11_reg[2]/P0001  & ~\sa11_reg[6]/NET0131  ;
  assign n11832 = n11812 & n11831 ;
  assign n11838 = ~n11830 & ~n11832 ;
  assign n11839 = ~n11835 & n11838 ;
  assign n11840 = ~n11837 & n11839 ;
  assign n11841 = ~\sa11_reg[1]/P0001  & ~n11840 ;
  assign n11813 = \sa11_reg[4]/P0001  & n11812 ;
  assign n11814 = \sa11_reg[3]/P0001  & n11813 ;
  assign n11815 = ~\sa11_reg[6]/NET0131  & n11814 ;
  assign n11816 = ~\sa11_reg[5]/P0001  & \sa11_reg[6]/NET0131  ;
  assign n11817 = ~\sa11_reg[4]/P0001  & n11816 ;
  assign n11818 = ~\sa11_reg[3]/P0001  & n11817 ;
  assign n11819 = ~n11815 & ~n11818 ;
  assign n11820 = \sa11_reg[2]/P0001  & ~n11819 ;
  assign n11821 = \sa11_reg[6]/NET0131  & \sa11_reg[7]/NET0131  ;
  assign n11822 = ~\sa11_reg[5]/P0001  & n11821 ;
  assign n11823 = ~\sa11_reg[2]/P0001  & \sa11_reg[4]/P0001  ;
  assign n11824 = n11822 & n11823 ;
  assign n11825 = \sa11_reg[5]/P0001  & ~\sa11_reg[7]/NET0131  ;
  assign n11826 = n11800 & n11825 ;
  assign n11827 = ~n11824 & ~n11826 ;
  assign n11828 = ~\sa11_reg[3]/P0001  & ~n11827 ;
  assign n11842 = ~n11820 & ~n11828 ;
  assign n11843 = ~n11841 & n11842 ;
  assign n11844 = ~n11811 & n11843 ;
  assign n11845 = ~\sa11_reg[0]/P0001  & ~n11844 ;
  assign n11921 = ~\sa11_reg[3]/P0001  & n11802 ;
  assign n11858 = \sa11_reg[3]/P0001  & \sa11_reg[6]/NET0131  ;
  assign n11925 = n11825 & n11858 ;
  assign n11928 = \sa11_reg[2]/P0001  & ~n11925 ;
  assign n11929 = ~n11921 & n11928 ;
  assign n11876 = ~\sa11_reg[5]/P0001  & ~\sa11_reg[6]/NET0131  ;
  assign n11926 = \sa11_reg[7]/NET0131  & n11794 ;
  assign n11927 = n11876 & n11926 ;
  assign n11847 = \sa11_reg[5]/P0001  & n11829 ;
  assign n11922 = ~\sa11_reg[3]/P0001  & n11847 ;
  assign n11923 = \sa11_reg[5]/P0001  & n11796 ;
  assign n11924 = ~\sa11_reg[6]/NET0131  & n11923 ;
  assign n11930 = ~n11922 & ~n11924 ;
  assign n11931 = ~n11927 & n11930 ;
  assign n11932 = n11929 & n11931 ;
  assign n11935 = ~\sa11_reg[3]/P0001  & n11822 ;
  assign n11933 = \sa11_reg[7]/NET0131  & n11833 ;
  assign n11934 = n11796 & n11933 ;
  assign n11877 = ~\sa11_reg[3]/P0001  & \sa11_reg[4]/P0001  ;
  assign n11936 = n11816 & n11877 ;
  assign n11937 = ~\sa11_reg[2]/P0001  & ~n11936 ;
  assign n11938 = ~n11934 & n11937 ;
  assign n11939 = ~n11935 & n11938 ;
  assign n11940 = ~n11932 & ~n11939 ;
  assign n11941 = n11792 & n11794 ;
  assign n11860 = ~\sa11_reg[3]/P0001  & ~\sa11_reg[4]/P0001  ;
  assign n11942 = n11825 & n11860 ;
  assign n11943 = ~\sa11_reg[6]/NET0131  & n11942 ;
  assign n11944 = ~n11941 & ~n11943 ;
  assign n11945 = ~n11940 & n11944 ;
  assign n11946 = ~\sa11_reg[1]/P0001  & ~n11945 ;
  assign n11882 = ~\sa11_reg[4]/P0001  & n11791 ;
  assign n11870 = ~\sa11_reg[6]/NET0131  & \sa11_reg[7]/NET0131  ;
  assign n11871 = ~\sa11_reg[5]/P0001  & n11870 ;
  assign n11883 = \sa11_reg[4]/P0001  & n11871 ;
  assign n11884 = ~n11882 & ~n11883 ;
  assign n11885 = ~\sa11_reg[2]/P0001  & ~n11884 ;
  assign n11880 = ~\sa11_reg[6]/NET0131  & n11796 ;
  assign n11881 = n11825 & n11880 ;
  assign n11878 = ~\sa11_reg[7]/NET0131  & n11877 ;
  assign n11879 = n11876 & n11878 ;
  assign n11886 = ~\sa11_reg[4]/P0001  & \sa11_reg[7]/NET0131  ;
  assign n11887 = n11831 & n11886 ;
  assign n11888 = \sa11_reg[1]/P0001  & ~n11887 ;
  assign n11889 = ~n11879 & n11888 ;
  assign n11890 = ~n11881 & n11889 ;
  assign n11891 = ~n11885 & n11890 ;
  assign n11900 = ~\sa11_reg[6]/NET0131  & n11794 ;
  assign n11901 = ~\sa11_reg[7]/NET0131  & n11900 ;
  assign n11902 = ~\sa11_reg[2]/P0001  & n11901 ;
  assign n11898 = \sa11_reg[4]/P0001  & n11798 ;
  assign n11899 = \sa11_reg[2]/P0001  & n11898 ;
  assign n11892 = \sa11_reg[5]/P0001  & \sa11_reg[7]/NET0131  ;
  assign n11893 = ~\sa11_reg[2]/P0001  & ~\sa11_reg[4]/P0001  ;
  assign n11894 = ~\sa11_reg[3]/P0001  & ~n11893 ;
  assign n11895 = n11892 & ~n11894 ;
  assign n11896 = n11858 & n11886 ;
  assign n11897 = ~\sa11_reg[1]/P0001  & ~n11896 ;
  assign n11903 = ~n11895 & n11897 ;
  assign n11904 = ~n11899 & n11903 ;
  assign n11905 = ~n11902 & n11904 ;
  assign n11906 = ~n11891 & ~n11905 ;
  assign n11853 = ~\sa11_reg[4]/P0001  & \sa11_reg[6]/NET0131  ;
  assign n11907 = n11853 & n11892 ;
  assign n11908 = \sa11_reg[2]/P0001  & ~n11907 ;
  assign n11863 = \sa11_reg[3]/P0001  & ~\sa11_reg[5]/P0001  ;
  assign n11909 = n11863 & n11870 ;
  assign n11910 = ~n11878 & ~n11880 ;
  assign n11911 = ~n11909 & n11910 ;
  assign n11912 = n11908 & n11911 ;
  assign n11913 = n11801 & n11858 ;
  assign n11914 = ~\sa11_reg[2]/P0001  & ~n11913 ;
  assign n11865 = n11829 & n11860 ;
  assign n11866 = ~\sa11_reg[5]/P0001  & n11865 ;
  assign n11915 = n11791 & n11796 ;
  assign n11916 = ~n11866 & ~n11915 ;
  assign n11917 = n11914 & n11916 ;
  assign n11918 = ~n11912 & ~n11917 ;
  assign n11919 = ~n11906 & ~n11918 ;
  assign n11920 = \sa11_reg[0]/P0001  & ~n11919 ;
  assign n11861 = \sa11_reg[7]/NET0131  & n11860 ;
  assign n11862 = n11833 & n11861 ;
  assign n11864 = ~n11829 & n11863 ;
  assign n11867 = ~n11862 & ~n11864 ;
  assign n11868 = ~n11866 & n11867 ;
  assign n11869 = ~\sa11_reg[2]/P0001  & ~n11868 ;
  assign n11859 = n11806 & n11858 ;
  assign n11872 = n11796 & n11871 ;
  assign n11873 = ~n11859 & ~n11872 ;
  assign n11874 = ~n11869 & n11873 ;
  assign n11875 = \sa11_reg[1]/P0001  & ~n11874 ;
  assign n11846 = \sa11_reg[2]/P0001  & \sa11_reg[3]/P0001  ;
  assign n11848 = n11846 & n11847 ;
  assign n11849 = n11791 & n11805 ;
  assign n11850 = \sa11_reg[4]/P0001  & n11849 ;
  assign n11851 = ~n11848 & ~n11850 ;
  assign n11852 = \sa11_reg[1]/P0001  & ~n11851 ;
  assign n11854 = n11812 & n11853 ;
  assign n11855 = ~\sa11_reg[2]/P0001  & n11854 ;
  assign n11856 = ~n11835 & ~n11855 ;
  assign n11857 = \sa11_reg[3]/P0001  & ~n11856 ;
  assign n11947 = ~n11852 & ~n11857 ;
  assign n11948 = ~n11875 & n11947 ;
  assign n11949 = ~n11920 & n11948 ;
  assign n11950 = ~n11946 & n11949 ;
  assign n11951 = ~n11845 & n11950 ;
  assign n11966 = \sa00_reg[3]/P0001  & ~\sa00_reg[4]/P0001  ;
  assign n11952 = ~\sa00_reg[6]/NET0131  & \sa00_reg[7]/NET0131  ;
  assign n12088 = \sa00_reg[5]/P0001  & n11952 ;
  assign n12089 = ~n11966 & n12088 ;
  assign n11978 = ~\sa00_reg[4]/P0001  & \sa00_reg[7]/NET0131  ;
  assign n12090 = ~\sa00_reg[5]/P0001  & n11978 ;
  assign n12091 = ~\sa00_reg[6]/NET0131  & n12090 ;
  assign n12092 = ~n12089 & ~n12091 ;
  assign n12093 = ~\sa00_reg[2]/P0001  & ~n12092 ;
  assign n12096 = ~\sa00_reg[5]/P0001  & \sa00_reg[7]/NET0131  ;
  assign n11955 = ~\sa00_reg[3]/P0001  & \sa00_reg[4]/P0001  ;
  assign n12097 = \sa00_reg[2]/P0001  & n11955 ;
  assign n12098 = n12096 & n12097 ;
  assign n11962 = \sa00_reg[6]/NET0131  & ~\sa00_reg[7]/NET0131  ;
  assign n11982 = \sa00_reg[3]/P0001  & \sa00_reg[4]/P0001  ;
  assign n12017 = n11962 & n11982 ;
  assign n12094 = \sa00_reg[2]/P0001  & \sa00_reg[5]/P0001  ;
  assign n12095 = n11962 & n12094 ;
  assign n12099 = ~n12017 & ~n12095 ;
  assign n12100 = ~n12098 & n12099 ;
  assign n12101 = ~n12093 & n12100 ;
  assign n12102 = \sa00_reg[1]/P0001  & ~n12101 ;
  assign n11994 = ~\sa00_reg[6]/NET0131  & n11966 ;
  assign n11995 = \sa00_reg[5]/P0001  & \sa00_reg[6]/NET0131  ;
  assign n12072 = ~\sa00_reg[2]/P0001  & n11995 ;
  assign n12073 = ~\sa00_reg[3]/P0001  & n12072 ;
  assign n12074 = ~n11994 & ~n12073 ;
  assign n12075 = ~\sa00_reg[7]/NET0131  & ~n12074 ;
  assign n11956 = ~\sa00_reg[6]/NET0131  & ~\sa00_reg[7]/NET0131  ;
  assign n11957 = ~\sa00_reg[5]/P0001  & n11956 ;
  assign n12068 = \sa00_reg[4]/P0001  & n11995 ;
  assign n12076 = ~n11957 & ~n12068 ;
  assign n12077 = \sa00_reg[2]/P0001  & ~n12076 ;
  assign n12078 = ~n12075 & ~n12077 ;
  assign n12079 = ~\sa00_reg[1]/P0001  & ~n12078 ;
  assign n11992 = \sa00_reg[3]/P0001  & ~\sa00_reg[5]/P0001  ;
  assign n12080 = \sa00_reg[4]/P0001  & n11956 ;
  assign n12081 = n11992 & n12080 ;
  assign n12035 = ~\sa00_reg[5]/P0001  & \sa00_reg[6]/NET0131  ;
  assign n12082 = ~\sa00_reg[4]/P0001  & n12035 ;
  assign n12083 = ~\sa00_reg[3]/P0001  & n12082 ;
  assign n12084 = ~n12081 & ~n12083 ;
  assign n12085 = \sa00_reg[2]/P0001  & ~n12084 ;
  assign n12014 = ~\sa00_reg[4]/P0001  & \sa00_reg[5]/P0001  ;
  assign n12015 = ~\sa00_reg[3]/P0001  & n11956 ;
  assign n12016 = n12014 & n12015 ;
  assign n12002 = \sa00_reg[6]/NET0131  & \sa00_reg[7]/NET0131  ;
  assign n12020 = ~\sa00_reg[3]/P0001  & ~\sa00_reg[5]/P0001  ;
  assign n12033 = n12002 & n12020 ;
  assign n12086 = ~\sa00_reg[2]/P0001  & \sa00_reg[4]/P0001  ;
  assign n12087 = n12033 & n12086 ;
  assign n12103 = ~n12016 & ~n12087 ;
  assign n12104 = ~n12085 & n12103 ;
  assign n12105 = ~n12079 & n12104 ;
  assign n12106 = ~n12102 & n12105 ;
  assign n12107 = ~\sa00_reg[0]/P0001  & ~n12106 ;
  assign n11979 = \sa00_reg[3]/P0001  & \sa00_reg[6]/NET0131  ;
  assign n12026 = \sa00_reg[5]/P0001  & ~\sa00_reg[7]/NET0131  ;
  assign n12027 = n11979 & n12026 ;
  assign n11975 = \sa00_reg[5]/P0001  & ~\sa00_reg[6]/NET0131  ;
  assign n12019 = n11966 & n11975 ;
  assign n12028 = \sa00_reg[2]/P0001  & ~n12019 ;
  assign n12029 = ~n12027 & n12028 ;
  assign n11959 = \sa00_reg[4]/P0001  & \sa00_reg[7]/NET0131  ;
  assign n11960 = ~\sa00_reg[5]/P0001  & ~\sa00_reg[6]/NET0131  ;
  assign n12024 = \sa00_reg[3]/P0001  & n11960 ;
  assign n12025 = n11959 & n12024 ;
  assign n12021 = n11978 & n12020 ;
  assign n12022 = ~\sa00_reg[6]/NET0131  & n12021 ;
  assign n11967 = \sa00_reg[5]/P0001  & n11956 ;
  assign n12023 = ~\sa00_reg[3]/P0001  & n11967 ;
  assign n12030 = ~n12022 & ~n12023 ;
  assign n12031 = ~n12025 & n12030 ;
  assign n12032 = n12029 & n12031 ;
  assign n11996 = \sa00_reg[7]/NET0131  & n11995 ;
  assign n12034 = n11966 & n11996 ;
  assign n12036 = n11955 & n12035 ;
  assign n12037 = ~\sa00_reg[2]/P0001  & ~n12033 ;
  assign n12038 = ~n12036 & n12037 ;
  assign n12039 = ~n12034 & n12038 ;
  assign n12040 = ~n12032 & ~n12039 ;
  assign n12018 = \sa00_reg[5]/P0001  & n12017 ;
  assign n12041 = ~n12016 & ~n12018 ;
  assign n12042 = ~n12040 & n12041 ;
  assign n12043 = ~\sa00_reg[1]/P0001  & ~n12042 ;
  assign n11961 = n11959 & n11960 ;
  assign n11963 = ~\sa00_reg[4]/P0001  & n11962 ;
  assign n11964 = ~n11961 & ~n11963 ;
  assign n11965 = ~\sa00_reg[2]/P0001  & ~n11964 ;
  assign n11968 = n11966 & n11967 ;
  assign n11958 = n11955 & n11957 ;
  assign n11953 = \sa00_reg[2]/P0001  & ~\sa00_reg[4]/P0001  ;
  assign n11954 = n11952 & n11953 ;
  assign n11969 = \sa00_reg[1]/P0001  & ~n11954 ;
  assign n11970 = ~n11958 & n11969 ;
  assign n11971 = ~n11968 & n11970 ;
  assign n11972 = ~n11965 & n11971 ;
  assign n11976 = n11959 & n11975 ;
  assign n11977 = \sa00_reg[2]/P0001  & n11976 ;
  assign n11973 = \sa00_reg[5]/P0001  & \sa00_reg[7]/NET0131  ;
  assign n11974 = \sa00_reg[3]/P0001  & n11973 ;
  assign n11985 = ~\sa00_reg[2]/P0001  & \sa00_reg[5]/P0001  ;
  assign n11986 = n11978 & n11985 ;
  assign n11987 = ~n11974 & ~n11986 ;
  assign n11988 = ~n11977 & n11987 ;
  assign n11980 = n11978 & n11979 ;
  assign n11981 = ~\sa00_reg[1]/P0001  & ~n11980 ;
  assign n11983 = n11956 & n11982 ;
  assign n11984 = ~\sa00_reg[2]/P0001  & n11983 ;
  assign n11989 = n11981 & ~n11984 ;
  assign n11990 = n11988 & n11989 ;
  assign n11991 = ~n11972 & ~n11990 ;
  assign n11997 = ~n11955 & ~n11996 ;
  assign n11998 = ~n11959 & ~n11997 ;
  assign n11993 = n11952 & n11992 ;
  assign n11999 = \sa00_reg[2]/P0001  & ~n11993 ;
  assign n12000 = ~n11994 & n11999 ;
  assign n12001 = ~n11998 & n12000 ;
  assign n12005 = ~\sa00_reg[3]/P0001  & ~\sa00_reg[4]/P0001  ;
  assign n12006 = n11957 & n12005 ;
  assign n12003 = n11992 & n12002 ;
  assign n12004 = ~\sa00_reg[2]/P0001  & ~n12003 ;
  assign n12007 = ~\sa00_reg[4]/P0001  & ~\sa00_reg[7]/NET0131  ;
  assign n12008 = n11979 & n12007 ;
  assign n12009 = n12004 & ~n12008 ;
  assign n12010 = ~n12006 & n12009 ;
  assign n12011 = ~n12001 & ~n12010 ;
  assign n12012 = ~n11991 & ~n12011 ;
  assign n12013 = \sa00_reg[0]/P0001  & ~n12012 ;
  assign n12045 = n12002 & n12005 ;
  assign n12046 = \sa00_reg[5]/P0001  & n12045 ;
  assign n12044 = ~n11956 & n11992 ;
  assign n12047 = ~n12006 & ~n12044 ;
  assign n12048 = ~n12046 & n12047 ;
  assign n12049 = ~\sa00_reg[2]/P0001  & ~n12048 ;
  assign n12050 = \sa00_reg[7]/NET0131  & n11982 ;
  assign n12051 = n12035 & n12050 ;
  assign n12052 = n11978 & n11992 ;
  assign n12053 = ~\sa00_reg[6]/NET0131  & n12052 ;
  assign n12059 = ~n12051 & ~n12053 ;
  assign n12054 = \sa00_reg[2]/P0001  & \sa00_reg[3]/P0001  ;
  assign n12055 = n11967 & n12054 ;
  assign n12056 = \sa00_reg[2]/P0001  & ~\sa00_reg[3]/P0001  ;
  assign n12057 = \sa00_reg[4]/P0001  & n11962 ;
  assign n12058 = n12056 & n12057 ;
  assign n12060 = ~n12055 & ~n12058 ;
  assign n12061 = n12059 & n12060 ;
  assign n12062 = ~n12049 & n12061 ;
  assign n12063 = \sa00_reg[1]/P0001  & ~n12062 ;
  assign n12069 = \sa00_reg[2]/P0001  & ~n12068 ;
  assign n12064 = ~\sa00_reg[5]/P0001  & ~\sa00_reg[7]/NET0131  ;
  assign n12065 = ~\sa00_reg[4]/P0001  & \sa00_reg[6]/NET0131  ;
  assign n12066 = n12064 & n12065 ;
  assign n12067 = ~\sa00_reg[2]/P0001  & ~n12066 ;
  assign n12070 = \sa00_reg[3]/P0001  & ~n12067 ;
  assign n12071 = ~n12069 & n12070 ;
  assign n12108 = ~n12063 & ~n12071 ;
  assign n12109 = ~n12013 & n12108 ;
  assign n12110 = ~n12043 & n12109 ;
  assign n12111 = ~n12107 & n12110 ;
  assign n12112 = n11951 & ~n12111 ;
  assign n12113 = ~n11951 & n12111 ;
  assign n12114 = ~n12112 & ~n12113 ;
  assign n12183 = ~n11817 & ~n11901 ;
  assign n12184 = \sa11_reg[2]/P0001  & ~n12183 ;
  assign n12188 = ~\sa11_reg[2]/P0001  & \sa11_reg[3]/P0001  ;
  assign n12189 = n11871 & n12188 ;
  assign n12127 = \sa11_reg[4]/P0001  & \sa11_reg[6]/NET0131  ;
  assign n12185 = n11892 & n12127 ;
  assign n12186 = ~\sa11_reg[3]/P0001  & n12185 ;
  assign n12187 = n11792 & ~n11805 ;
  assign n12190 = ~n12186 & ~n12187 ;
  assign n12191 = ~n12189 & n12190 ;
  assign n12192 = ~n12184 & n12191 ;
  assign n12193 = ~\sa11_reg[1]/P0001  & ~n12192 ;
  assign n12169 = ~\sa11_reg[4]/P0001  & n11876 ;
  assign n12170 = ~n11813 & ~n11923 ;
  assign n12171 = ~n12169 & n12170 ;
  assign n12172 = \sa11_reg[1]/P0001  & ~n12171 ;
  assign n12167 = ~n11915 & ~n11925 ;
  assign n12168 = ~\sa11_reg[4]/P0001  & n11825 ;
  assign n12173 = n12167 & ~n12168 ;
  assign n12174 = ~n12172 & n12173 ;
  assign n12175 = ~\sa11_reg[2]/P0001  & ~n12174 ;
  assign n12176 = n11798 & n11877 ;
  assign n12177 = n11794 & n11847 ;
  assign n12178 = ~n12176 & ~n12177 ;
  assign n12179 = n11796 & n11870 ;
  assign n12180 = ~n11879 & ~n12179 ;
  assign n12181 = n12178 & n12180 ;
  assign n12182 = \sa11_reg[1]/P0001  & ~n12181 ;
  assign n12194 = ~\sa11_reg[5]/P0001  & n11791 ;
  assign n12195 = n11860 & n12194 ;
  assign n12196 = ~n12186 & ~n12195 ;
  assign n12197 = \sa11_reg[2]/P0001  & ~n12196 ;
  assign n12198 = n11792 & n11796 ;
  assign n12199 = ~n11824 & ~n12198 ;
  assign n12200 = ~n12197 & n12199 ;
  assign n12201 = ~n12182 & n12200 ;
  assign n12202 = ~n12175 & n12201 ;
  assign n12203 = ~n12193 & n12202 ;
  assign n12204 = \sa11_reg[0]/P0001  & ~n12203 ;
  assign n12119 = n11829 & n11863 ;
  assign n12132 = ~n11935 & ~n12119 ;
  assign n12124 = n11833 & n11860 ;
  assign n12125 = ~\sa11_reg[7]/NET0131  & n12124 ;
  assign n12120 = \sa11_reg[3]/P0001  & n11870 ;
  assign n12121 = ~\sa11_reg[2]/P0001  & n12120 ;
  assign n12122 = ~n11853 & ~n11877 ;
  assign n12123 = n11892 & n12122 ;
  assign n12133 = ~n12121 & ~n12123 ;
  assign n12134 = ~n12125 & n12133 ;
  assign n12135 = n12132 & n12134 ;
  assign n12115 = n11797 & n11877 ;
  assign n12116 = ~\sa11_reg[3]/P0001  & n11882 ;
  assign n12117 = ~n12115 & ~n12116 ;
  assign n12118 = ~\sa11_reg[2]/P0001  & ~n12117 ;
  assign n12126 = \sa11_reg[3]/P0001  & n11892 ;
  assign n12128 = \sa11_reg[5]/P0001  & n12127 ;
  assign n12129 = ~\sa11_reg[7]/NET0131  & n12128 ;
  assign n12130 = ~n12126 & ~n12129 ;
  assign n12131 = \sa11_reg[2]/P0001  & ~n12130 ;
  assign n12136 = ~n12118 & ~n12131 ;
  assign n12137 = n12135 & n12136 ;
  assign n12138 = \sa11_reg[1]/P0001  & ~n12137 ;
  assign n12152 = \sa11_reg[4]/P0001  & n11892 ;
  assign n12153 = ~\sa11_reg[4]/P0001  & n11812 ;
  assign n12154 = ~n12152 & ~n12153 ;
  assign n12155 = \sa11_reg[3]/P0001  & ~n12154 ;
  assign n12156 = ~n11800 & ~n11936 ;
  assign n12157 = ~\sa11_reg[7]/NET0131  & ~n12156 ;
  assign n12158 = ~n12155 & ~n12157 ;
  assign n12159 = \sa11_reg[2]/P0001  & ~n12158 ;
  assign n12142 = n11876 & n11877 ;
  assign n12143 = ~n12124 & ~n12142 ;
  assign n12144 = \sa11_reg[7]/NET0131  & ~n12143 ;
  assign n12145 = \sa11_reg[2]/P0001  & ~\sa11_reg[5]/P0001  ;
  assign n12146 = ~\sa11_reg[3]/P0001  & n11829 ;
  assign n12147 = ~n11880 & ~n12146 ;
  assign n12148 = n12145 & ~n12147 ;
  assign n12149 = ~n12144 & ~n12148 ;
  assign n12150 = ~\sa11_reg[1]/P0001  & ~n12149 ;
  assign n12139 = n11801 & n11853 ;
  assign n12140 = ~n11814 & ~n12139 ;
  assign n12141 = ~\sa11_reg[2]/P0001  & ~n12140 ;
  assign n12151 = n11800 & n11812 ;
  assign n12160 = n11798 & n11823 ;
  assign n12161 = ~n12151 & ~n12160 ;
  assign n12162 = ~n12141 & n12161 ;
  assign n12163 = ~n12150 & n12162 ;
  assign n12164 = ~n12159 & n12163 ;
  assign n12165 = ~n12138 & n12164 ;
  assign n12166 = ~\sa11_reg[0]/P0001  & ~n12165 ;
  assign n12206 = \sa11_reg[2]/P0001  & n11877 ;
  assign n12207 = ~n11871 & ~n12194 ;
  assign n12208 = ~n11933 & n12207 ;
  assign n12209 = n12206 & ~n12208 ;
  assign n12210 = \sa11_reg[5]/P0001  & n11794 ;
  assign n12211 = n11831 & n12210 ;
  assign n12212 = ~n11865 & ~n12211 ;
  assign n12213 = ~n12209 & n12212 ;
  assign n12214 = ~\sa11_reg[1]/P0001  & ~n12213 ;
  assign n12222 = ~\sa11_reg[1]/P0001  & ~\sa11_reg[2]/P0001  ;
  assign n12224 = \sa11_reg[5]/P0001  & n11861 ;
  assign n12223 = n11801 & n12127 ;
  assign n12225 = ~n11941 & ~n12223 ;
  assign n12226 = ~n12224 & n12225 ;
  assign n12227 = n12222 & ~n12226 ;
  assign n12218 = n11792 & n12206 ;
  assign n12217 = \sa11_reg[3]/P0001  & n12151 ;
  assign n12219 = ~n12160 & ~n12217 ;
  assign n12220 = ~n12218 & n12219 ;
  assign n12221 = \sa11_reg[1]/P0001  & ~n12220 ;
  assign n12205 = \sa11_reg[4]/P0001  & n11848 ;
  assign n12215 = ~n11881 & ~n11935 ;
  assign n12216 = ~\sa11_reg[2]/P0001  & ~n12215 ;
  assign n12228 = ~n12205 & ~n12216 ;
  assign n12229 = ~n12221 & n12228 ;
  assign n12230 = ~n12227 & n12229 ;
  assign n12231 = ~n12214 & n12230 ;
  assign n12232 = ~n12166 & n12231 ;
  assign n12233 = ~n12204 & n12232 ;
  assign n12303 = \sa22_reg[3]/P0001  & ~\sa22_reg[4]/P0001  ;
  assign n12355 = \sa22_reg[5]/P0001  & n12303 ;
  assign n12297 = \sa22_reg[4]/P0001  & \sa22_reg[7]/NET0131  ;
  assign n12290 = ~\sa22_reg[4]/P0001  & \sa22_reg[6]/NET0131  ;
  assign n12356 = ~\sa22_reg[5]/P0001  & ~n12290 ;
  assign n12357 = ~n12297 & n12356 ;
  assign n12358 = ~n12355 & ~n12357 ;
  assign n12359 = \sa22_reg[1]/P0001  & ~n12358 ;
  assign n12349 = \sa22_reg[5]/P0001  & ~\sa22_reg[7]/NET0131  ;
  assign n12350 = \sa22_reg[3]/P0001  & n12349 ;
  assign n12351 = \sa22_reg[6]/NET0131  & n12350 ;
  assign n12251 = \sa22_reg[6]/NET0131  & ~\sa22_reg[7]/NET0131  ;
  assign n12352 = \sa22_reg[3]/P0001  & n12251 ;
  assign n12353 = ~\sa22_reg[4]/P0001  & n12352 ;
  assign n12354 = ~n12351 & ~n12353 ;
  assign n12360 = ~\sa22_reg[4]/P0001  & n12349 ;
  assign n12361 = n12354 & ~n12360 ;
  assign n12362 = ~n12359 & n12361 ;
  assign n12363 = ~\sa22_reg[2]/P0001  & ~n12362 ;
  assign n12257 = ~\sa22_reg[5]/P0001  & \sa22_reg[6]/NET0131  ;
  assign n12314 = ~\sa22_reg[4]/P0001  & n12257 ;
  assign n12260 = \sa22_reg[3]/P0001  & \sa22_reg[4]/P0001  ;
  assign n12315 = ~\sa22_reg[6]/NET0131  & n12260 ;
  assign n12316 = ~\sa22_reg[7]/NET0131  & n12315 ;
  assign n12317 = ~n12314 & ~n12316 ;
  assign n12318 = \sa22_reg[2]/P0001  & ~n12317 ;
  assign n12263 = \sa22_reg[3]/P0001  & ~\sa22_reg[6]/NET0131  ;
  assign n12291 = ~\sa22_reg[5]/P0001  & \sa22_reg[7]/NET0131  ;
  assign n12324 = n12263 & n12291 ;
  assign n12325 = ~\sa22_reg[2]/P0001  & n12324 ;
  assign n12244 = ~\sa22_reg[3]/P0001  & \sa22_reg[4]/P0001  ;
  assign n12239 = \sa22_reg[5]/P0001  & \sa22_reg[6]/NET0131  ;
  assign n12319 = \sa22_reg[7]/NET0131  & n12239 ;
  assign n12320 = n12244 & n12319 ;
  assign n12321 = \sa22_reg[5]/P0001  & n12251 ;
  assign n12322 = \sa22_reg[2]/P0001  & ~\sa22_reg[3]/P0001  ;
  assign n12323 = n12321 & ~n12322 ;
  assign n12326 = ~n12320 & ~n12323 ;
  assign n12327 = ~n12325 & n12326 ;
  assign n12328 = ~n12318 & n12327 ;
  assign n12329 = ~\sa22_reg[1]/P0001  & ~n12328 ;
  assign n12245 = \sa22_reg[5]/P0001  & ~\sa22_reg[6]/NET0131  ;
  assign n12330 = ~\sa22_reg[3]/P0001  & n12245 ;
  assign n12331 = n12297 & n12330 ;
  assign n12300 = ~\sa22_reg[6]/NET0131  & ~\sa22_reg[7]/NET0131  ;
  assign n12332 = \sa22_reg[5]/P0001  & n12300 ;
  assign n12333 = n12260 & n12332 ;
  assign n12338 = ~n12331 & ~n12333 ;
  assign n12234 = ~\sa22_reg[5]/P0001  & ~\sa22_reg[6]/NET0131  ;
  assign n12334 = ~\sa22_reg[7]/NET0131  & n12244 ;
  assign n12335 = n12234 & n12334 ;
  assign n12336 = ~\sa22_reg[4]/P0001  & n12263 ;
  assign n12337 = \sa22_reg[7]/NET0131  & n12336 ;
  assign n12339 = ~n12335 & ~n12337 ;
  assign n12340 = n12338 & n12339 ;
  assign n12341 = \sa22_reg[1]/P0001  & ~n12340 ;
  assign n12344 = \sa22_reg[4]/P0001  & n12291 ;
  assign n12345 = \sa22_reg[6]/NET0131  & n12344 ;
  assign n12346 = ~\sa22_reg[2]/P0001  & n12345 ;
  assign n12342 = \sa22_reg[2]/P0001  & n12320 ;
  assign n12343 = n12303 & n12321 ;
  assign n12277 = ~\sa22_reg[5]/P0001  & ~\sa22_reg[7]/NET0131  ;
  assign n12347 = n12277 & n12290 ;
  assign n12348 = n12322 & n12347 ;
  assign n12364 = ~n12343 & ~n12348 ;
  assign n12365 = ~n12342 & n12364 ;
  assign n12366 = ~n12346 & n12365 ;
  assign n12367 = ~n12341 & n12366 ;
  assign n12368 = ~n12329 & n12367 ;
  assign n12369 = ~n12363 & n12368 ;
  assign n12370 = \sa22_reg[0]/P0001  & ~n12369 ;
  assign n12238 = ~\sa22_reg[3]/P0001  & ~\sa22_reg[4]/P0001  ;
  assign n12242 = ~\sa22_reg[7]/NET0131  & n12238 ;
  assign n12243 = \sa22_reg[6]/NET0131  & n12242 ;
  assign n12246 = n12244 & n12245 ;
  assign n12247 = ~\sa22_reg[2]/P0001  & ~n12246 ;
  assign n12248 = ~n12243 & n12247 ;
  assign n12252 = \sa22_reg[4]/P0001  & n12251 ;
  assign n12253 = \sa22_reg[5]/P0001  & n12252 ;
  assign n12249 = \sa22_reg[5]/P0001  & \sa22_reg[7]/NET0131  ;
  assign n12250 = \sa22_reg[3]/P0001  & n12249 ;
  assign n12254 = \sa22_reg[2]/P0001  & ~n12250 ;
  assign n12255 = ~n12253 & n12254 ;
  assign n12256 = ~n12248 & ~n12255 ;
  assign n12235 = \sa22_reg[3]/P0001  & n12234 ;
  assign n12236 = ~\sa22_reg[7]/NET0131  & n12235 ;
  assign n12237 = \sa22_reg[1]/P0001  & ~n12236 ;
  assign n12240 = n12238 & n12239 ;
  assign n12241 = ~\sa22_reg[7]/NET0131  & n12240 ;
  assign n12258 = ~\sa22_reg[3]/P0001  & \sa22_reg[7]/NET0131  ;
  assign n12259 = n12257 & n12258 ;
  assign n12266 = ~\sa22_reg[6]/NET0131  & \sa22_reg[7]/NET0131  ;
  assign n12267 = ~\sa22_reg[4]/P0001  & \sa22_reg[5]/P0001  ;
  assign n12268 = n12266 & n12267 ;
  assign n12269 = ~n12259 & ~n12268 ;
  assign n12270 = ~n12241 & n12269 ;
  assign n12261 = \sa22_reg[5]/P0001  & n12260 ;
  assign n12262 = \sa22_reg[7]/NET0131  & n12261 ;
  assign n12264 = \sa22_reg[7]/NET0131  & n12263 ;
  assign n12265 = ~\sa22_reg[2]/P0001  & n12264 ;
  assign n12271 = ~n12262 & ~n12265 ;
  assign n12272 = n12270 & n12271 ;
  assign n12273 = n12237 & n12272 ;
  assign n12274 = ~n12256 & n12273 ;
  assign n12275 = n12234 & n12258 ;
  assign n12276 = \sa22_reg[4]/P0001  & n12275 ;
  assign n12284 = ~\sa22_reg[1]/P0001  & ~n12276 ;
  assign n12282 = \sa22_reg[2]/P0001  & ~\sa22_reg[4]/P0001  ;
  assign n12283 = n12235 & n12282 ;
  assign n12278 = \sa22_reg[2]/P0001  & ~\sa22_reg[6]/NET0131  ;
  assign n12279 = n12277 & n12278 ;
  assign n12280 = ~\sa22_reg[3]/P0001  & n12279 ;
  assign n12281 = \sa22_reg[7]/NET0131  & n12240 ;
  assign n12285 = ~n12280 & ~n12281 ;
  assign n12286 = ~n12283 & n12285 ;
  assign n12287 = n12284 & n12286 ;
  assign n12288 = ~n12274 & ~n12287 ;
  assign n12302 = \sa22_reg[6]/NET0131  & n12244 ;
  assign n12304 = ~n12302 & ~n12303 ;
  assign n12305 = n12277 & ~n12304 ;
  assign n12301 = ~\sa22_reg[4]/P0001  & n12300 ;
  assign n12306 = ~n12262 & ~n12301 ;
  assign n12307 = ~n12305 & n12306 ;
  assign n12308 = \sa22_reg[2]/P0001  & ~n12307 ;
  assign n12289 = n12260 & n12277 ;
  assign n12292 = n12290 & n12291 ;
  assign n12293 = ~n12289 & ~n12292 ;
  assign n12294 = ~\sa22_reg[2]/P0001  & ~n12293 ;
  assign n12295 = ~\sa22_reg[4]/P0001  & n12234 ;
  assign n12296 = ~\sa22_reg[7]/NET0131  & n12295 ;
  assign n12298 = n12245 & n12297 ;
  assign n12299 = ~\sa22_reg[2]/P0001  & n12298 ;
  assign n12309 = ~n12296 & ~n12299 ;
  assign n12310 = ~n12294 & n12309 ;
  assign n12311 = ~n12308 & n12310 ;
  assign n12312 = ~n12288 & n12311 ;
  assign n12313 = ~\sa22_reg[0]/P0001  & ~n12312 ;
  assign n12373 = ~n12251 & ~n12266 ;
  assign n12374 = ~\sa22_reg[5]/P0001  & ~n12373 ;
  assign n12375 = ~n12319 & ~n12374 ;
  assign n12376 = \sa22_reg[2]/P0001  & n12244 ;
  assign n12377 = ~n12375 & n12376 ;
  assign n12371 = ~\sa22_reg[6]/NET0131  & n12242 ;
  assign n12372 = n12261 & n12278 ;
  assign n12378 = ~n12371 & ~n12372 ;
  assign n12379 = ~n12377 & n12378 ;
  assign n12380 = ~\sa22_reg[1]/P0001  & ~n12379 ;
  assign n12393 = n12239 & n12334 ;
  assign n12394 = \sa22_reg[2]/P0001  & n12393 ;
  assign n12395 = ~\sa22_reg[4]/P0001  & n12277 ;
  assign n12396 = n12263 & n12395 ;
  assign n12397 = ~n12299 & ~n12396 ;
  assign n12398 = ~n12394 & n12397 ;
  assign n12399 = \sa22_reg[1]/P0001  & ~n12398 ;
  assign n12383 = ~\sa22_reg[1]/P0001  & ~\sa22_reg[2]/P0001  ;
  assign n12385 = ~\sa22_reg[4]/P0001  & n12258 ;
  assign n12386 = \sa22_reg[5]/P0001  & n12385 ;
  assign n12384 = n12251 & n12261 ;
  assign n12387 = ~n12345 & ~n12384 ;
  assign n12388 = ~n12386 & n12387 ;
  assign n12389 = n12383 & ~n12388 ;
  assign n12381 = ~\sa22_reg[7]/NET0131  & n12261 ;
  assign n12382 = n12278 & n12381 ;
  assign n12390 = n12303 & n12332 ;
  assign n12391 = ~n12259 & ~n12390 ;
  assign n12392 = ~\sa22_reg[2]/P0001  & ~n12391 ;
  assign n12400 = ~n12382 & ~n12392 ;
  assign n12401 = ~n12389 & n12400 ;
  assign n12402 = ~n12399 & n12401 ;
  assign n12403 = ~n12380 & n12402 ;
  assign n12404 = ~n12313 & n12403 ;
  assign n12405 = ~n12370 & n12404 ;
  assign n12406 = n12233 & ~n12405 ;
  assign n12407 = ~n12233 & n12405 ;
  assign n12408 = ~n12406 & ~n12407 ;
  assign n12476 = \sa33_reg[3]/P0001  & ~\sa33_reg[4]/P0001  ;
  assign n12526 = \sa33_reg[5]/P0001  & n12476 ;
  assign n12460 = ~\sa33_reg[4]/P0001  & \sa33_reg[6]/P0001  ;
  assign n12467 = \sa33_reg[4]/P0001  & \sa33_reg[7]/NET0131  ;
  assign n12527 = ~n12460 & ~n12467 ;
  assign n12528 = ~\sa33_reg[5]/P0001  & n12527 ;
  assign n12529 = ~n12526 & ~n12528 ;
  assign n12530 = \sa33_reg[1]/P0001  & ~n12529 ;
  assign n12510 = \sa33_reg[5]/P0001  & ~\sa33_reg[7]/NET0131  ;
  assign n12525 = ~\sa33_reg[4]/P0001  & n12510 ;
  assign n12457 = \sa33_reg[4]/P0001  & ~\sa33_reg[5]/P0001  ;
  assign n12414 = \sa33_reg[6]/P0001  & ~\sa33_reg[7]/NET0131  ;
  assign n12531 = \sa33_reg[3]/P0001  & n12414 ;
  assign n12532 = ~n12457 & n12531 ;
  assign n12533 = ~n12525 & ~n12532 ;
  assign n12534 = ~n12530 & n12533 ;
  assign n12535 = ~\sa33_reg[2]/P0001  & ~n12534 ;
  assign n12419 = \sa33_reg[3]/P0001  & \sa33_reg[4]/P0001  ;
  assign n12465 = ~\sa33_reg[6]/P0001  & ~\sa33_reg[7]/NET0131  ;
  assign n12495 = n12419 & n12465 ;
  assign n12446 = ~\sa33_reg[4]/P0001  & ~\sa33_reg[5]/P0001  ;
  assign n12496 = \sa33_reg[6]/P0001  & n12446 ;
  assign n12497 = ~n12495 & ~n12496 ;
  assign n12498 = \sa33_reg[2]/P0001  & ~n12497 ;
  assign n12418 = \sa33_reg[5]/P0001  & \sa33_reg[7]/NET0131  ;
  assign n12448 = ~\sa33_reg[3]/P0001  & \sa33_reg[4]/P0001  ;
  assign n12449 = \sa33_reg[6]/P0001  & n12448 ;
  assign n12501 = n12418 & n12449 ;
  assign n12409 = ~\sa33_reg[6]/P0001  & \sa33_reg[7]/NET0131  ;
  assign n12426 = \sa33_reg[3]/P0001  & ~\sa33_reg[5]/P0001  ;
  assign n12493 = n12409 & n12426 ;
  assign n12494 = ~\sa33_reg[2]/P0001  & n12493 ;
  assign n12472 = \sa33_reg[2]/P0001  & ~\sa33_reg[3]/P0001  ;
  assign n12499 = \sa33_reg[5]/P0001  & n12414 ;
  assign n12500 = ~n12472 & n12499 ;
  assign n12502 = ~n12494 & ~n12500 ;
  assign n12503 = ~n12501 & n12502 ;
  assign n12504 = ~n12498 & n12503 ;
  assign n12505 = ~\sa33_reg[1]/P0001  & ~n12504 ;
  assign n12506 = n12418 & n12448 ;
  assign n12507 = ~\sa33_reg[6]/P0001  & n12506 ;
  assign n12509 = n12409 & n12476 ;
  assign n12513 = ~n12507 & ~n12509 ;
  assign n12473 = ~\sa33_reg[5]/P0001  & n12465 ;
  assign n12508 = n12448 & n12473 ;
  assign n12511 = n12419 & n12510 ;
  assign n12512 = ~\sa33_reg[6]/P0001  & n12511 ;
  assign n12514 = ~n12508 & ~n12512 ;
  assign n12515 = n12513 & n12514 ;
  assign n12516 = \sa33_reg[1]/P0001  & ~n12515 ;
  assign n12479 = ~\sa33_reg[3]/P0001  & ~\sa33_reg[4]/P0001  ;
  assign n12517 = ~\sa33_reg[5]/P0001  & n12414 ;
  assign n12518 = n12479 & n12517 ;
  assign n12519 = ~n12501 & ~n12518 ;
  assign n12520 = \sa33_reg[2]/P0001  & ~n12519 ;
  assign n12521 = ~\sa33_reg[5]/P0001  & \sa33_reg[6]/P0001  ;
  assign n12522 = n12467 & n12521 ;
  assign n12523 = ~\sa33_reg[2]/P0001  & n12522 ;
  assign n12524 = n12476 & n12499 ;
  assign n12536 = ~n12523 & ~n12524 ;
  assign n12537 = ~n12520 & n12536 ;
  assign n12538 = ~n12516 & n12537 ;
  assign n12539 = ~n12505 & n12538 ;
  assign n12540 = ~n12535 & n12539 ;
  assign n12541 = \sa33_reg[0]/P0001  & ~n12540 ;
  assign n12433 = ~\sa33_reg[3]/P0001  & n12414 ;
  assign n12434 = ~\sa33_reg[4]/P0001  & n12433 ;
  assign n12429 = \sa33_reg[5]/P0001  & ~\sa33_reg[6]/P0001  ;
  assign n12430 = ~\sa33_reg[3]/P0001  & n12429 ;
  assign n12431 = \sa33_reg[4]/P0001  & n12430 ;
  assign n12432 = \sa33_reg[3]/P0001  & n12409 ;
  assign n12435 = ~n12431 & ~n12432 ;
  assign n12436 = ~n12434 & n12435 ;
  assign n12437 = ~\sa33_reg[2]/P0001  & ~n12436 ;
  assign n12421 = \sa33_reg[3]/P0001  & n12418 ;
  assign n12422 = \sa33_reg[4]/P0001  & n12414 ;
  assign n12423 = \sa33_reg[5]/P0001  & n12422 ;
  assign n12424 = ~n12421 & ~n12423 ;
  assign n12425 = \sa33_reg[2]/P0001  & ~n12424 ;
  assign n12412 = \sa33_reg[6]/P0001  & \sa33_reg[7]/NET0131  ;
  assign n12413 = ~\sa33_reg[5]/P0001  & n12412 ;
  assign n12410 = ~\sa33_reg[4]/P0001  & \sa33_reg[5]/P0001  ;
  assign n12415 = n12410 & n12414 ;
  assign n12416 = ~n12413 & ~n12415 ;
  assign n12417 = ~\sa33_reg[3]/P0001  & ~n12416 ;
  assign n12427 = ~\sa33_reg[6]/P0001  & n12426 ;
  assign n12428 = ~\sa33_reg[7]/NET0131  & n12427 ;
  assign n12411 = n12409 & n12410 ;
  assign n12420 = n12418 & n12419 ;
  assign n12438 = ~n12411 & ~n12420 ;
  assign n12439 = ~n12428 & n12438 ;
  assign n12440 = ~n12417 & n12439 ;
  assign n12441 = ~n12425 & n12440 ;
  assign n12442 = ~n12437 & n12441 ;
  assign n12443 = \sa33_reg[1]/P0001  & ~n12442 ;
  assign n12447 = \sa33_reg[3]/P0001  & n12446 ;
  assign n12450 = ~\sa33_reg[5]/P0001  & n12449 ;
  assign n12451 = ~n12447 & ~n12450 ;
  assign n12452 = ~\sa33_reg[7]/NET0131  & ~n12451 ;
  assign n12444 = ~\sa33_reg[4]/P0001  & ~\sa33_reg[7]/NET0131  ;
  assign n12445 = ~\sa33_reg[6]/P0001  & n12444 ;
  assign n12453 = ~n12420 & ~n12445 ;
  assign n12454 = ~n12452 & n12453 ;
  assign n12455 = \sa33_reg[2]/P0001  & ~n12454 ;
  assign n12470 = ~\sa33_reg[3]/P0001  & n12409 ;
  assign n12471 = n12457 & n12470 ;
  assign n12474 = n12472 & n12473 ;
  assign n12483 = ~n12471 & ~n12474 ;
  assign n12475 = ~\sa33_reg[5]/P0001  & ~\sa33_reg[6]/P0001  ;
  assign n12477 = \sa33_reg[2]/P0001  & n12476 ;
  assign n12478 = n12475 & n12477 ;
  assign n12480 = \sa33_reg[5]/P0001  & \sa33_reg[6]/P0001  ;
  assign n12481 = \sa33_reg[7]/NET0131  & n12480 ;
  assign n12482 = n12479 & n12481 ;
  assign n12484 = ~n12478 & ~n12482 ;
  assign n12485 = n12483 & n12484 ;
  assign n12486 = ~\sa33_reg[1]/P0001  & ~n12485 ;
  assign n12456 = ~\sa33_reg[2]/P0001  & \sa33_reg[3]/P0001  ;
  assign n12458 = ~\sa33_reg[7]/NET0131  & n12457 ;
  assign n12459 = n12456 & n12458 ;
  assign n12461 = ~\sa33_reg[5]/P0001  & \sa33_reg[7]/NET0131  ;
  assign n12462 = n12460 & n12461 ;
  assign n12463 = ~\sa33_reg[2]/P0001  & n12462 ;
  assign n12464 = ~n12459 & ~n12463 ;
  assign n12466 = n12446 & n12465 ;
  assign n12468 = n12429 & n12467 ;
  assign n12469 = ~\sa33_reg[2]/P0001  & n12468 ;
  assign n12487 = ~n12466 & ~n12469 ;
  assign n12488 = n12464 & n12487 ;
  assign n12489 = ~n12486 & n12488 ;
  assign n12490 = ~n12455 & n12489 ;
  assign n12491 = ~n12443 & n12490 ;
  assign n12492 = ~\sa33_reg[0]/P0001  & ~n12491 ;
  assign n12551 = \sa33_reg[7]/NET0131  & n12479 ;
  assign n12552 = \sa33_reg[5]/P0001  & n12551 ;
  assign n12550 = \sa33_reg[6]/P0001  & n12511 ;
  assign n12553 = ~n12522 & ~n12550 ;
  assign n12554 = ~n12552 & n12553 ;
  assign n12555 = ~\sa33_reg[2]/P0001  & ~n12554 ;
  assign n12544 = ~\sa33_reg[5]/P0001  & n12409 ;
  assign n12545 = ~n12517 & ~n12544 ;
  assign n12546 = ~n12481 & n12545 ;
  assign n12547 = \sa33_reg[4]/P0001  & n12472 ;
  assign n12548 = ~n12546 & n12547 ;
  assign n12542 = \sa33_reg[2]/P0001  & n12419 ;
  assign n12543 = n12429 & n12542 ;
  assign n12549 = n12465 & n12479 ;
  assign n12556 = ~n12543 & ~n12549 ;
  assign n12557 = ~n12548 & n12556 ;
  assign n12558 = ~n12555 & n12557 ;
  assign n12559 = ~\sa33_reg[1]/P0001  & ~n12558 ;
  assign n12569 = n12448 & n12510 ;
  assign n12570 = \sa33_reg[6]/P0001  & n12569 ;
  assign n12571 = \sa33_reg[2]/P0001  & n12570 ;
  assign n12572 = n12427 & n12444 ;
  assign n12573 = ~n12469 & ~n12572 ;
  assign n12574 = ~n12571 & n12573 ;
  assign n12575 = \sa33_reg[1]/P0001  & ~n12574 ;
  assign n12560 = \sa33_reg[2]/P0001  & \sa33_reg[3]/P0001  ;
  assign n12561 = \sa33_reg[5]/P0001  & n12465 ;
  assign n12562 = n12560 & n12561 ;
  assign n12563 = \sa33_reg[4]/P0001  & n12562 ;
  assign n12564 = ~\sa33_reg[3]/P0001  & n12413 ;
  assign n12565 = n12429 & n12476 ;
  assign n12566 = ~\sa33_reg[7]/NET0131  & n12565 ;
  assign n12567 = ~n12564 & ~n12566 ;
  assign n12568 = ~\sa33_reg[2]/P0001  & ~n12567 ;
  assign n12576 = ~n12563 & ~n12568 ;
  assign n12577 = ~n12575 & n12576 ;
  assign n12578 = ~n12559 & n12577 ;
  assign n12579 = ~n12492 & n12578 ;
  assign n12580 = ~n12541 & n12579 ;
  assign n12581 = \u0_w_reg[0][29]/P0001  & ~n12580 ;
  assign n12582 = ~\u0_w_reg[0][29]/P0001  & n12580 ;
  assign n12583 = ~n12581 & ~n12582 ;
  assign n12584 = n12408 & n12583 ;
  assign n12585 = ~n12408 & ~n12583 ;
  assign n12586 = ~n12584 & ~n12585 ;
  assign n12588 = n12114 & n12586 ;
  assign n12587 = ~n12114 & ~n12586 ;
  assign n12589 = ~\ld_r_reg/P0001  & ~n12587 ;
  assign n12590 = ~n12588 & n12589 ;
  assign n12592 = \text_in_r_reg[125]/P0001  & \u0_w_reg[0][29]/P0001  ;
  assign n12591 = ~\text_in_r_reg[125]/P0001  & ~\u0_w_reg[0][29]/P0001  ;
  assign n12593 = \ld_r_reg/P0001  & ~n12591 ;
  assign n12594 = ~n12592 & n12593 ;
  assign n12595 = ~n12590 & ~n12594 ;
  assign n12614 = n11955 & n11975 ;
  assign n12608 = n11962 & n12005 ;
  assign n12613 = \sa00_reg[3]/P0001  & n11952 ;
  assign n12615 = ~n12608 & ~n12613 ;
  assign n12616 = ~n12614 & n12615 ;
  assign n12617 = ~\sa00_reg[2]/P0001  & ~n12616 ;
  assign n12605 = \sa00_reg[5]/P0001  & n12057 ;
  assign n12606 = ~n11974 & ~n12605 ;
  assign n12607 = \sa00_reg[2]/P0001  & ~n12606 ;
  assign n12609 = ~n12050 & ~n12608 ;
  assign n12610 = \sa00_reg[5]/P0001  & ~n12609 ;
  assign n12612 = n11952 & n12014 ;
  assign n12611 = n11956 & n11992 ;
  assign n12618 = ~n12033 & ~n12611 ;
  assign n12619 = ~n12612 & n12618 ;
  assign n12620 = ~n12610 & n12619 ;
  assign n12621 = ~n12607 & n12620 ;
  assign n12622 = ~n12617 & n12621 ;
  assign n12623 = \sa00_reg[1]/P0001  & ~n12622 ;
  assign n12596 = \sa00_reg[2]/P0001  & n11966 ;
  assign n12597 = ~\sa00_reg[7]/NET0131  & n12056 ;
  assign n12598 = ~n12596 & ~n12597 ;
  assign n12599 = ~\sa00_reg[6]/NET0131  & ~n12598 ;
  assign n12600 = n11952 & n11955 ;
  assign n12601 = ~n12599 & ~n12600 ;
  assign n12602 = ~\sa00_reg[5]/P0001  & ~n12601 ;
  assign n12603 = ~n12046 & ~n12602 ;
  assign n12604 = ~\sa00_reg[1]/P0001  & ~n12603 ;
  assign n12632 = \sa00_reg[4]/P0001  & n11973 ;
  assign n12633 = ~\sa00_reg[4]/P0001  & n12064 ;
  assign n12634 = ~n12632 & ~n12633 ;
  assign n12635 = \sa00_reg[3]/P0001  & ~n12634 ;
  assign n12636 = ~\sa00_reg[4]/P0001  & n11956 ;
  assign n12637 = ~\sa00_reg[7]/NET0131  & n12036 ;
  assign n12638 = ~n12636 & ~n12637 ;
  assign n12639 = ~n12635 & n12638 ;
  assign n12640 = \sa00_reg[2]/P0001  & ~n12639 ;
  assign n12624 = n11978 & n12035 ;
  assign n12625 = \sa00_reg[4]/P0001  & n12064 ;
  assign n12626 = \sa00_reg[3]/P0001  & n12625 ;
  assign n12627 = ~n12624 & ~n12626 ;
  assign n12628 = ~\sa00_reg[2]/P0001  & ~n12627 ;
  assign n12629 = ~\sa00_reg[4]/P0001  & n11960 ;
  assign n12630 = ~\sa00_reg[7]/NET0131  & n12629 ;
  assign n12631 = n12086 & n12088 ;
  assign n12641 = ~n12630 & ~n12631 ;
  assign n12642 = ~n12628 & n12641 ;
  assign n12643 = ~n12640 & n12642 ;
  assign n12644 = ~n12604 & n12643 ;
  assign n12645 = ~n12623 & n12644 ;
  assign n12646 = ~\sa00_reg[0]/P0001  & ~n12645 ;
  assign n12673 = ~n11983 & ~n12082 ;
  assign n12674 = \sa00_reg[2]/P0001  & ~n12673 ;
  assign n12672 = ~\sa00_reg[2]/P0001  & n11993 ;
  assign n12647 = n11955 & n11996 ;
  assign n12651 = \sa00_reg[5]/P0001  & n11962 ;
  assign n12671 = ~n12056 & n12651 ;
  assign n12675 = ~n12647 & ~n12671 ;
  assign n12676 = ~n12672 & n12675 ;
  assign n12677 = ~n12674 & n12676 ;
  assign n12678 = ~\sa00_reg[1]/P0001  & ~n12677 ;
  assign n12664 = ~n11994 & ~n12614 ;
  assign n12665 = \sa00_reg[7]/NET0131  & ~n12664 ;
  assign n12666 = ~\sa00_reg[6]/NET0131  & n11982 ;
  assign n12667 = n12026 & n12666 ;
  assign n12668 = ~n11958 & ~n12667 ;
  assign n12669 = ~n12665 & n12668 ;
  assign n12670 = \sa00_reg[1]/P0001  & ~n12669 ;
  assign n12648 = ~\sa00_reg[5]/P0001  & n12608 ;
  assign n12649 = ~n12647 & ~n12648 ;
  assign n12650 = \sa00_reg[2]/P0001  & ~n12649 ;
  assign n12652 = n11966 & n12651 ;
  assign n12679 = ~n12650 & ~n12652 ;
  assign n12653 = ~n12008 & ~n12027 ;
  assign n12654 = ~n12007 & ~n12035 ;
  assign n12655 = ~\sa00_reg[5]/P0001  & ~n11959 ;
  assign n12656 = ~n12654 & ~n12655 ;
  assign n12657 = n12653 & ~n12656 ;
  assign n12658 = ~\sa00_reg[2]/P0001  & ~n12657 ;
  assign n12659 = \sa00_reg[1]/P0001  & ~\sa00_reg[2]/P0001  ;
  assign n12660 = \sa00_reg[5]/P0001  & n11966 ;
  assign n12661 = ~n12625 & ~n12629 ;
  assign n12662 = ~n12660 & n12661 ;
  assign n12663 = n12659 & ~n12662 ;
  assign n12680 = ~n12658 & ~n12663 ;
  assign n12681 = n12679 & n12680 ;
  assign n12682 = ~n12670 & n12681 ;
  assign n12683 = ~n12678 & n12682 ;
  assign n12684 = \sa00_reg[0]/P0001  & ~n12683 ;
  assign n12693 = ~\sa00_reg[3]/P0001  & n12014 ;
  assign n12694 = \sa00_reg[7]/NET0131  & n12693 ;
  assign n12692 = n11959 & n12035 ;
  assign n12695 = ~n12018 & ~n12692 ;
  assign n12696 = ~n12694 & n12695 ;
  assign n12697 = ~\sa00_reg[2]/P0001  & ~n12696 ;
  assign n12685 = ~\sa00_reg[5]/P0001  & n11952 ;
  assign n12686 = ~\sa00_reg[5]/P0001  & n11962 ;
  assign n12687 = ~n12685 & ~n12686 ;
  assign n12688 = ~n11996 & n12687 ;
  assign n12689 = n12097 & ~n12688 ;
  assign n12690 = n12094 & n12666 ;
  assign n12691 = n11956 & n12005 ;
  assign n12698 = ~n12690 & ~n12691 ;
  assign n12699 = ~n12689 & n12698 ;
  assign n12700 = ~n12697 & n12699 ;
  assign n12701 = ~\sa00_reg[1]/P0001  & ~n12700 ;
  assign n12706 = n12056 & n12605 ;
  assign n12705 = n11994 & n12064 ;
  assign n12707 = ~n12631 & ~n12705 ;
  assign n12708 = ~n12706 & n12707 ;
  assign n12709 = \sa00_reg[1]/P0001  & ~n12708 ;
  assign n12702 = ~\sa00_reg[7]/NET0131  & n12690 ;
  assign n12703 = ~n11968 & ~n12033 ;
  assign n12704 = ~\sa00_reg[2]/P0001  & ~n12703 ;
  assign n12710 = ~n12702 & ~n12704 ;
  assign n12711 = ~n12709 & n12710 ;
  assign n12712 = ~n12701 & n12711 ;
  assign n12713 = ~n12684 & n12712 ;
  assign n12714 = ~n12646 & n12713 ;
  assign n12753 = \sa22_reg[5]/P0001  & n12266 ;
  assign n12754 = ~n12303 & n12753 ;
  assign n12755 = ~\sa22_reg[4]/P0001  & \sa22_reg[7]/NET0131  ;
  assign n12756 = n12234 & n12755 ;
  assign n12757 = ~n12754 & ~n12756 ;
  assign n12758 = ~\sa22_reg[2]/P0001  & ~n12757 ;
  assign n12761 = n12322 & n12344 ;
  assign n12759 = n12251 & n12260 ;
  assign n12760 = \sa22_reg[2]/P0001  & n12321 ;
  assign n12762 = ~n12759 & ~n12760 ;
  assign n12763 = ~n12761 & n12762 ;
  assign n12764 = ~n12758 & n12763 ;
  assign n12765 = \sa22_reg[1]/P0001  & ~n12764 ;
  assign n12747 = ~\sa22_reg[3]/P0001  & n12321 ;
  assign n12748 = ~\sa22_reg[2]/P0001  & n12747 ;
  assign n12736 = \sa22_reg[4]/P0001  & n12239 ;
  assign n12746 = \sa22_reg[2]/P0001  & n12736 ;
  assign n12745 = ~\sa22_reg[7]/NET0131  & n12336 ;
  assign n12749 = ~n12279 & ~n12745 ;
  assign n12750 = ~n12746 & n12749 ;
  assign n12751 = ~n12748 & n12750 ;
  assign n12752 = ~\sa22_reg[1]/P0001  & ~n12751 ;
  assign n12738 = n12267 & n12300 ;
  assign n12739 = ~n12346 & ~n12738 ;
  assign n12740 = ~\sa22_reg[3]/P0001  & ~n12739 ;
  assign n12741 = ~\sa22_reg[3]/P0001  & n12314 ;
  assign n12742 = ~\sa22_reg[6]/NET0131  & n12289 ;
  assign n12743 = ~n12741 & ~n12742 ;
  assign n12744 = \sa22_reg[2]/P0001  & ~n12743 ;
  assign n12766 = ~n12740 & ~n12744 ;
  assign n12767 = ~n12752 & n12766 ;
  assign n12768 = ~n12765 & n12767 ;
  assign n12769 = ~\sa22_reg[0]/P0001  & ~n12768 ;
  assign n12803 = ~n12244 & ~n12258 ;
  assign n12804 = n12257 & ~n12803 ;
  assign n12732 = \sa22_reg[3]/P0001  & \sa22_reg[6]/NET0131  ;
  assign n12805 = \sa22_reg[7]/NET0131  & n12732 ;
  assign n12806 = n12267 & n12805 ;
  assign n12807 = ~\sa22_reg[2]/P0001  & ~n12806 ;
  assign n12808 = ~n12804 & n12807 ;
  assign n12809 = n12234 & n12385 ;
  assign n12810 = \sa22_reg[2]/P0001  & ~n12809 ;
  assign n12814 = n12263 & n12267 ;
  assign n12815 = ~n12351 & ~n12814 ;
  assign n12811 = \sa22_reg[3]/P0001  & n12297 ;
  assign n12812 = n12234 & n12811 ;
  assign n12813 = ~\sa22_reg[3]/P0001  & n12332 ;
  assign n12816 = ~n12812 & ~n12813 ;
  assign n12817 = n12815 & n12816 ;
  assign n12818 = n12810 & n12817 ;
  assign n12819 = ~n12808 & ~n12818 ;
  assign n12802 = ~\sa22_reg[3]/P0001  & n12738 ;
  assign n12820 = ~n12384 & ~n12802 ;
  assign n12821 = ~n12819 & n12820 ;
  assign n12822 = ~\sa22_reg[1]/P0001  & ~n12821 ;
  assign n12772 = ~\sa22_reg[4]/P0001  & n12251 ;
  assign n12773 = n12234 & n12297 ;
  assign n12774 = ~n12772 & ~n12773 ;
  assign n12775 = ~\sa22_reg[2]/P0001  & ~n12774 ;
  assign n12770 = \sa22_reg[1]/P0001  & ~n12390 ;
  assign n12771 = n12278 & n12755 ;
  assign n12776 = ~n12335 & ~n12771 ;
  assign n12777 = n12770 & n12776 ;
  assign n12778 = ~n12775 & n12777 ;
  assign n12779 = ~\sa22_reg[2]/P0001  & ~\sa22_reg[7]/NET0131  ;
  assign n12780 = n12315 & n12779 ;
  assign n12781 = ~\sa22_reg[1]/P0001  & ~n12780 ;
  assign n12785 = \sa22_reg[2]/P0001  & n12298 ;
  assign n12782 = n12732 & n12755 ;
  assign n12731 = ~\sa22_reg[2]/P0001  & ~\sa22_reg[4]/P0001  ;
  assign n12783 = ~\sa22_reg[3]/P0001  & ~n12731 ;
  assign n12784 = n12249 & ~n12783 ;
  assign n12786 = ~n12782 & ~n12784 ;
  assign n12787 = ~n12785 & n12786 ;
  assign n12788 = n12781 & n12787 ;
  assign n12789 = ~n12778 & ~n12788 ;
  assign n12717 = ~\sa22_reg[3]/P0001  & n12296 ;
  assign n12790 = n12291 & n12732 ;
  assign n12791 = ~\sa22_reg[2]/P0001  & ~n12790 ;
  assign n12792 = ~n12353 & n12791 ;
  assign n12793 = ~n12717 & n12792 ;
  assign n12794 = \sa22_reg[2]/P0001  & ~n12324 ;
  assign n12795 = n12249 & n12290 ;
  assign n12796 = ~n12334 & ~n12336 ;
  assign n12797 = ~n12795 & n12796 ;
  assign n12798 = n12794 & n12797 ;
  assign n12799 = ~n12793 & ~n12798 ;
  assign n12800 = ~n12789 & ~n12799 ;
  assign n12801 = \sa22_reg[0]/P0001  & ~n12800 ;
  assign n12715 = ~\sa22_reg[5]/P0001  & ~n12300 ;
  assign n12716 = \sa22_reg[3]/P0001  & n12715 ;
  assign n12718 = ~n12281 & ~n12716 ;
  assign n12719 = ~n12717 & n12718 ;
  assign n12720 = ~\sa22_reg[2]/P0001  & ~n12719 ;
  assign n12721 = \sa22_reg[3]/P0001  & n12257 ;
  assign n12722 = n12297 & n12721 ;
  assign n12723 = n12278 & n12350 ;
  assign n12726 = ~n12722 & ~n12723 ;
  assign n12724 = ~\sa22_reg[4]/P0001  & n12324 ;
  assign n12725 = n12252 & n12322 ;
  assign n12727 = ~n12724 & ~n12725 ;
  assign n12728 = n12726 & n12727 ;
  assign n12729 = ~n12720 & n12728 ;
  assign n12730 = \sa22_reg[1]/P0001  & ~n12729 ;
  assign n12733 = n12277 & n12732 ;
  assign n12734 = n12731 & n12733 ;
  assign n12735 = \sa22_reg[2]/P0001  & \sa22_reg[3]/P0001  ;
  assign n12737 = n12735 & n12736 ;
  assign n12823 = ~n12734 & ~n12737 ;
  assign n12824 = ~n12730 & n12823 ;
  assign n12825 = ~n12801 & n12824 ;
  assign n12826 = ~n12822 & n12825 ;
  assign n12827 = ~n12769 & n12826 ;
  assign n12828 = n11951 & ~n12827 ;
  assign n12829 = ~n11951 & n12827 ;
  assign n12830 = ~n12828 & ~n12829 ;
  assign n12831 = ~n12714 & ~n12830 ;
  assign n12832 = n12714 & n12830 ;
  assign n12833 = ~n12831 & ~n12832 ;
  assign n12834 = \u0_w_reg[0][21]/P0001  & ~n12580 ;
  assign n12835 = ~\u0_w_reg[0][21]/P0001  & n12580 ;
  assign n12836 = ~n12834 & ~n12835 ;
  assign n12837 = n12405 & n12836 ;
  assign n12838 = ~n12405 & ~n12836 ;
  assign n12839 = ~n12837 & ~n12838 ;
  assign n12841 = n12833 & n12839 ;
  assign n12840 = ~n12833 & ~n12839 ;
  assign n12842 = ~\ld_r_reg/P0001  & ~n12840 ;
  assign n12843 = ~n12841 & n12842 ;
  assign n12845 = ~\text_in_r_reg[117]/P0001  & \u0_w_reg[0][21]/P0001  ;
  assign n12844 = \text_in_r_reg[117]/P0001  & ~\u0_w_reg[0][21]/P0001  ;
  assign n12846 = \ld_r_reg/P0001  & ~n12844 ;
  assign n12847 = ~n12845 & n12846 ;
  assign n12848 = ~n12843 & ~n12847 ;
  assign n12849 = n12233 & ~n12714 ;
  assign n12850 = ~n12233 & n12714 ;
  assign n12851 = ~n12849 & ~n12850 ;
  assign n12852 = ~n12827 & ~n12851 ;
  assign n12853 = n12827 & n12851 ;
  assign n12854 = ~n12852 & ~n12853 ;
  assign n12942 = ~\sa33_reg[2]/P0001  & n12409 ;
  assign n12943 = ~n12457 & ~n12526 ;
  assign n12944 = n12942 & n12943 ;
  assign n12948 = \sa33_reg[4]/P0001  & n12531 ;
  assign n12945 = \sa33_reg[2]/P0001  & \sa33_reg[6]/P0001  ;
  assign n12946 = n12510 & n12945 ;
  assign n12947 = n12461 & n12547 ;
  assign n12949 = ~n12946 & ~n12947 ;
  assign n12950 = ~n12948 & n12949 ;
  assign n12951 = ~n12944 & n12950 ;
  assign n12952 = \sa33_reg[1]/P0001  & ~n12951 ;
  assign n12932 = \sa33_reg[4]/P0001  & n12480 ;
  assign n12933 = ~n12473 & ~n12932 ;
  assign n12934 = \sa33_reg[2]/P0001  & ~n12933 ;
  assign n12935 = n12465 & n12476 ;
  assign n12936 = ~n12934 & ~n12935 ;
  assign n12937 = ~\sa33_reg[1]/P0001  & ~n12936 ;
  assign n12927 = ~\sa33_reg[3]/P0001  & n12499 ;
  assign n12928 = ~\sa33_reg[1]/P0001  & n12927 ;
  assign n12929 = \sa33_reg[4]/P0001  & n12564 ;
  assign n12930 = ~n12928 & ~n12929 ;
  assign n12931 = ~\sa33_reg[2]/P0001  & ~n12930 ;
  assign n12909 = n12479 & n12561 ;
  assign n12938 = n12479 & n12521 ;
  assign n12939 = n12419 & n12473 ;
  assign n12940 = ~n12938 & ~n12939 ;
  assign n12941 = \sa33_reg[2]/P0001  & ~n12940 ;
  assign n12953 = ~n12909 & ~n12941 ;
  assign n12954 = ~n12931 & n12953 ;
  assign n12955 = ~n12937 & n12954 ;
  assign n12956 = ~n12952 & n12955 ;
  assign n12957 = ~\sa33_reg[0]/P0001  & ~n12956 ;
  assign n12910 = n12475 & n12551 ;
  assign n12911 = \sa33_reg[2]/P0001  & ~n12910 ;
  assign n12912 = ~\sa33_reg[3]/P0001  & n12561 ;
  assign n12915 = ~n12565 & ~n12912 ;
  assign n12913 = \sa33_reg[5]/P0001  & n12531 ;
  assign n12914 = n12432 & n12457 ;
  assign n12916 = ~n12913 & ~n12914 ;
  assign n12917 = n12915 & n12916 ;
  assign n12918 = n12911 & n12917 ;
  assign n12920 = ~\sa33_reg[2]/P0001  & ~n12450 ;
  assign n12919 = n12476 & n12481 ;
  assign n12921 = ~n12564 & ~n12919 ;
  assign n12922 = n12920 & n12921 ;
  assign n12923 = ~n12918 & ~n12922 ;
  assign n12924 = ~n12550 & ~n12909 ;
  assign n12925 = ~n12923 & n12924 ;
  assign n12926 = ~\sa33_reg[1]/P0001  & ~n12925 ;
  assign n12871 = \sa33_reg[1]/P0001  & ~n12566 ;
  assign n12868 = \sa33_reg[7]/NET0131  & ~n12475 ;
  assign n12869 = ~\sa33_reg[2]/P0001  & ~n12527 ;
  assign n12870 = ~n12868 & n12869 ;
  assign n12855 = \sa33_reg[2]/P0001  & ~\sa33_reg[4]/P0001  ;
  assign n12872 = n12409 & n12855 ;
  assign n12873 = ~n12508 & ~n12872 ;
  assign n12874 = ~n12870 & n12873 ;
  assign n12875 = n12871 & n12874 ;
  assign n12876 = ~\sa33_reg[4]/P0001  & \sa33_reg[7]/NET0131  ;
  assign n12877 = \sa33_reg[3]/P0001  & \sa33_reg[6]/P0001  ;
  assign n12878 = n12876 & n12877 ;
  assign n12879 = ~\sa33_reg[1]/P0001  & ~n12878 ;
  assign n12880 = ~\sa33_reg[6]/P0001  & n12419 ;
  assign n12881 = ~\sa33_reg[2]/P0001  & ~\sa33_reg[7]/NET0131  ;
  assign n12882 = n12880 & n12881 ;
  assign n12887 = n12879 & ~n12882 ;
  assign n12883 = \sa33_reg[2]/P0001  & n12468 ;
  assign n12884 = ~\sa33_reg[2]/P0001  & ~\sa33_reg[4]/P0001  ;
  assign n12885 = ~\sa33_reg[3]/P0001  & ~n12884 ;
  assign n12886 = n12418 & ~n12885 ;
  assign n12888 = ~n12883 & ~n12886 ;
  assign n12889 = n12887 & n12888 ;
  assign n12890 = ~n12875 & ~n12889 ;
  assign n12856 = n12481 & n12855 ;
  assign n12857 = ~n12419 & ~n12479 ;
  assign n12858 = n12527 & n12857 ;
  assign n12859 = \sa33_reg[2]/P0001  & ~n12493 ;
  assign n12860 = ~n12858 & n12859 ;
  assign n12863 = ~\sa33_reg[5]/P0001  & n12549 ;
  assign n12861 = n12412 & n12426 ;
  assign n12862 = ~\sa33_reg[2]/P0001  & ~n12861 ;
  assign n12864 = n12414 & n12476 ;
  assign n12865 = n12862 & ~n12864 ;
  assign n12866 = ~n12863 & n12865 ;
  assign n12867 = ~n12860 & ~n12866 ;
  assign n12891 = ~n12856 & ~n12867 ;
  assign n12892 = ~n12890 & n12891 ;
  assign n12893 = \sa33_reg[0]/P0001  & ~n12892 ;
  assign n12894 = n12426 & ~n12465 ;
  assign n12895 = ~n12482 & ~n12894 ;
  assign n12896 = ~n12863 & n12895 ;
  assign n12897 = ~\sa33_reg[2]/P0001  & ~n12896 ;
  assign n12898 = n12422 & n12472 ;
  assign n12901 = ~n12562 & ~n12898 ;
  assign n12899 = n12476 & n12544 ;
  assign n12900 = n12413 & n12419 ;
  assign n12902 = ~n12899 & ~n12900 ;
  assign n12903 = n12901 & n12902 ;
  assign n12904 = ~n12897 & n12903 ;
  assign n12905 = \sa33_reg[1]/P0001  & ~n12904 ;
  assign n12906 = n12414 & n12446 ;
  assign n12907 = n12456 & n12906 ;
  assign n12908 = n12480 & n12542 ;
  assign n12958 = ~n12907 & ~n12908 ;
  assign n12959 = ~n12905 & n12958 ;
  assign n12960 = ~n12893 & n12959 ;
  assign n12961 = ~n12926 & n12960 ;
  assign n12962 = ~n12957 & n12961 ;
  assign n12963 = \u0_w_reg[0][13]/P0001  & ~n12962 ;
  assign n12964 = ~\u0_w_reg[0][13]/P0001  & n12962 ;
  assign n12965 = ~n12963 & ~n12964 ;
  assign n12966 = n12580 & n12965 ;
  assign n12967 = ~n12580 & ~n12965 ;
  assign n12968 = ~n12966 & ~n12967 ;
  assign n12970 = n12854 & ~n12968 ;
  assign n12969 = ~n12854 & n12968 ;
  assign n12971 = ~\ld_r_reg/P0001  & ~n12969 ;
  assign n12972 = ~n12970 & n12971 ;
  assign n12974 = \text_in_r_reg[109]/P0001  & \u0_w_reg[0][13]/P0001  ;
  assign n12973 = ~\text_in_r_reg[109]/P0001  & ~\u0_w_reg[0][13]/P0001  ;
  assign n12975 = \ld_r_reg/P0001  & ~n12973 ;
  assign n12976 = ~n12974 & n12975 ;
  assign n12977 = ~n12972 & ~n12976 ;
  assign n12978 = ~n12111 & ~n12851 ;
  assign n12979 = n12111 & n12851 ;
  assign n12980 = ~n12978 & ~n12979 ;
  assign n12981 = \u0_w_reg[0][5]/P0001  & ~n12962 ;
  assign n12982 = ~\u0_w_reg[0][5]/P0001  & n12962 ;
  assign n12983 = ~n12981 & ~n12982 ;
  assign n12984 = n12405 & n12983 ;
  assign n12985 = ~n12405 & ~n12983 ;
  assign n12986 = ~n12984 & ~n12985 ;
  assign n12988 = n12980 & ~n12986 ;
  assign n12987 = ~n12980 & n12986 ;
  assign n12989 = ~\ld_r_reg/P0001  & ~n12987 ;
  assign n12990 = ~n12988 & n12989 ;
  assign n12992 = \text_in_r_reg[101]/P0001  & \u0_w_reg[0][5]/P0001  ;
  assign n12991 = ~\text_in_r_reg[101]/P0001  & ~\u0_w_reg[0][5]/P0001  ;
  assign n12993 = \ld_r_reg/P0001  & ~n12991 ;
  assign n12994 = ~n12992 & n12993 ;
  assign n12995 = ~n12990 & ~n12994 ;
  assign n13018 = n11985 & n12015 ;
  assign n13019 = ~n11976 & ~n13018 ;
  assign n13020 = ~n12628 & n13019 ;
  assign n13021 = ~\sa00_reg[1]/P0001  & ~n13020 ;
  assign n12997 = ~\sa00_reg[4]/P0001  & n12033 ;
  assign n12998 = ~n12057 & ~n12612 ;
  assign n12999 = ~n12997 & n12998 ;
  assign n13000 = \sa00_reg[1]/P0001  & ~n12999 ;
  assign n12996 = ~n12017 & ~n12647 ;
  assign n13001 = ~n12630 & n12996 ;
  assign n13002 = ~n13000 & n13001 ;
  assign n13003 = \sa00_reg[2]/P0001  & ~n13002 ;
  assign n13012 = ~\sa00_reg[4]/P0001  & n11974 ;
  assign n13013 = ~n12667 & ~n13012 ;
  assign n13014 = \sa00_reg[1]/P0001  & ~n13013 ;
  assign n13007 = \sa00_reg[1]/P0001  & n12020 ;
  assign n13008 = ~n12065 & n13007 ;
  assign n13006 = n11962 & n12014 ;
  assign n13009 = ~n12614 & ~n13006 ;
  assign n13010 = ~n13008 & n13009 ;
  assign n13011 = ~\sa00_reg[2]/P0001  & ~n13010 ;
  assign n13004 = \sa00_reg[2]/P0001  & ~\sa00_reg[5]/P0001  ;
  assign n13005 = n12613 & n13004 ;
  assign n13015 = ~\sa00_reg[1]/P0001  & \sa00_reg[2]/P0001  ;
  assign n13016 = ~n12050 & ~n12686 ;
  assign n13017 = n13015 & ~n13016 ;
  assign n13022 = ~n13005 & ~n13017 ;
  assign n13023 = ~n13011 & n13022 ;
  assign n13024 = ~n13014 & n13023 ;
  assign n13025 = ~n13003 & n13024 ;
  assign n13026 = ~n13021 & n13025 ;
  assign n13027 = \sa00_reg[0]/P0001  & ~n13026 ;
  assign n13028 = \sa00_reg[4]/P0001  & n11960 ;
  assign n13029 = ~\sa00_reg[3]/P0001  & n13028 ;
  assign n13033 = n12004 & ~n13029 ;
  assign n13030 = ~\sa00_reg[4]/P0001  & n12044 ;
  assign n13031 = n11955 & n12026 ;
  assign n13032 = \sa00_reg[6]/NET0131  & n13031 ;
  assign n13034 = ~n13030 & ~n13032 ;
  assign n13035 = n13033 & n13034 ;
  assign n13038 = ~\sa00_reg[3]/P0001  & n12629 ;
  assign n13036 = \sa00_reg[6]/NET0131  & n11955 ;
  assign n13037 = n12096 & n13036 ;
  assign n13039 = \sa00_reg[2]/P0001  & ~n13037 ;
  assign n13040 = ~n13038 & n13039 ;
  assign n13041 = ~n13035 & ~n13040 ;
  assign n13046 = ~\sa00_reg[1]/P0001  & ~n12052 ;
  assign n13044 = ~\sa00_reg[2]/P0001  & \sa00_reg[3]/P0001  ;
  assign n13045 = n11959 & n13044 ;
  assign n13047 = ~n13006 & ~n13045 ;
  assign n13048 = n13046 & n13047 ;
  assign n13042 = ~\sa00_reg[3]/P0001  & n11952 ;
  assign n13043 = ~\sa00_reg[4]/P0001  & n13042 ;
  assign n13049 = ~n12055 & ~n13037 ;
  assign n13050 = ~n13043 & n13049 ;
  assign n13051 = n13048 & n13050 ;
  assign n13053 = ~\sa00_reg[2]/P0001  & n12630 ;
  assign n13052 = n12056 & ~n12634 ;
  assign n13054 = \sa00_reg[1]/P0001  & ~n12018 ;
  assign n13055 = ~n13052 & n13054 ;
  assign n13056 = ~n13053 & n13055 ;
  assign n13057 = ~n13051 & ~n13056 ;
  assign n13058 = ~n13041 & ~n13057 ;
  assign n13059 = ~\sa00_reg[0]/P0001  & ~n13058 ;
  assign n13069 = ~\sa00_reg[6]/NET0131  & n11974 ;
  assign n13068 = ~\sa00_reg[5]/P0001  & n12057 ;
  assign n13070 = ~n11976 & ~n13068 ;
  assign n13071 = ~n13069 & n13070 ;
  assign n13072 = ~\sa00_reg[2]/P0001  & ~n13071 ;
  assign n13073 = n11995 & n12005 ;
  assign n13074 = ~\sa00_reg[4]/P0001  & n12002 ;
  assign n13075 = n12094 & n13074 ;
  assign n13078 = ~n13073 & ~n13075 ;
  assign n13076 = n12054 & n12636 ;
  assign n13077 = ~\sa00_reg[6]/NET0131  & n12050 ;
  assign n13079 = ~n13076 & ~n13077 ;
  assign n13080 = n13078 & n13079 ;
  assign n13081 = ~n13072 & n13080 ;
  assign n13082 = ~\sa00_reg[1]/P0001  & ~n13081 ;
  assign n13060 = ~\sa00_reg[2]/P0001  & n11968 ;
  assign n13062 = ~\sa00_reg[6]/NET0131  & n12625 ;
  assign n13061 = n11973 & n11994 ;
  assign n13063 = ~n12691 & ~n13061 ;
  assign n13064 = ~n13062 & n13063 ;
  assign n13065 = \sa00_reg[2]/P0001  & ~n13064 ;
  assign n13066 = ~n13060 & ~n13065 ;
  assign n13067 = \sa00_reg[1]/P0001  & ~n13066 ;
  assign n13083 = ~n12015 & ~n12017 ;
  assign n13084 = n13004 & ~n13083 ;
  assign n13085 = n11976 & n13044 ;
  assign n13086 = ~n12006 & ~n13085 ;
  assign n13087 = ~n13084 & n13086 ;
  assign n13088 = ~n13067 & n13087 ;
  assign n13089 = ~n13082 & n13088 ;
  assign n13090 = ~n13059 & n13089 ;
  assign n13091 = ~n13027 & n13090 ;
  assign n13116 = ~\sa11_reg[2]/P0001  & n11922 ;
  assign n13114 = ~n11926 & ~n12194 ;
  assign n13115 = \sa11_reg[2]/P0001  & ~n13114 ;
  assign n13117 = ~n11898 & ~n13115 ;
  assign n13118 = ~n13116 & n13117 ;
  assign n13119 = ~n12141 & n13118 ;
  assign n13120 = ~\sa11_reg[1]/P0001  & ~n13119 ;
  assign n13101 = ~\sa11_reg[3]/P0001  & n12139 ;
  assign n13100 = ~\sa11_reg[7]/NET0131  & n12127 ;
  assign n13102 = n11800 & n11892 ;
  assign n13103 = ~n13100 & ~n13102 ;
  assign n13104 = ~n13101 & n13103 ;
  assign n13105 = \sa11_reg[2]/P0001  & ~n13104 ;
  assign n13106 = ~\sa11_reg[2]/P0001  & ~\sa11_reg[3]/P0001  ;
  assign n13107 = ~\sa11_reg[5]/P0001  & n13106 ;
  assign n13108 = ~n11853 & n13107 ;
  assign n13109 = n11796 & n11892 ;
  assign n13110 = ~n12177 & ~n13109 ;
  assign n13111 = ~n13108 & n13110 ;
  assign n13112 = ~n13105 & n13111 ;
  assign n13113 = \sa11_reg[1]/P0001  & ~n13112 ;
  assign n13092 = ~\sa11_reg[4]/P0001  & ~\sa11_reg[7]/NET0131  ;
  assign n13093 = n11833 & n13092 ;
  assign n13094 = ~n12115 & ~n13093 ;
  assign n13095 = ~\sa11_reg[2]/P0001  & ~n13094 ;
  assign n13096 = ~n11795 & ~n12186 ;
  assign n13097 = ~n11909 & ~n12151 ;
  assign n13098 = n13096 & n13097 ;
  assign n13099 = \sa11_reg[2]/P0001  & ~n13098 ;
  assign n13121 = ~n13095 & ~n13099 ;
  assign n13122 = ~n13113 & n13121 ;
  assign n13123 = ~n13120 & n13122 ;
  assign n13124 = \sa11_reg[0]/P0001  & ~n13123 ;
  assign n13128 = n11914 & ~n12142 ;
  assign n13125 = ~\sa11_reg[4]/P0001  & n11864 ;
  assign n13126 = n11825 & n11877 ;
  assign n13127 = \sa11_reg[6]/NET0131  & n13126 ;
  assign n13129 = ~n13125 & ~n13127 ;
  assign n13130 = n13128 & n13129 ;
  assign n13131 = \sa11_reg[6]/NET0131  & n11877 ;
  assign n13132 = n11801 & n13131 ;
  assign n13133 = n11860 & n11876 ;
  assign n13134 = \sa11_reg[2]/P0001  & ~n13133 ;
  assign n13135 = ~n13132 & n13134 ;
  assign n13136 = ~n13130 & ~n13135 ;
  assign n13138 = n11796 & n11801 ;
  assign n13141 = ~\sa11_reg[1]/P0001  & ~n13093 ;
  assign n13142 = ~n13138 & n13141 ;
  assign n13143 = ~n11848 & ~n13132 ;
  assign n13137 = ~\sa11_reg[2]/P0001  & n11926 ;
  assign n13139 = ~\sa11_reg[3]/P0001  & n11870 ;
  assign n13140 = ~\sa11_reg[4]/P0001  & n13139 ;
  assign n13144 = ~n13137 & ~n13140 ;
  assign n13145 = n13143 & n13144 ;
  assign n13146 = n13142 & n13145 ;
  assign n13147 = n11805 & ~n12154 ;
  assign n13148 = ~\sa11_reg[2]/P0001  & n12151 ;
  assign n13149 = \sa11_reg[1]/P0001  & ~n11941 ;
  assign n13150 = ~n13148 & n13149 ;
  assign n13151 = ~n13147 & n13150 ;
  assign n13152 = ~n13146 & ~n13151 ;
  assign n13153 = ~n13136 & ~n13152 ;
  assign n13154 = ~\sa11_reg[0]/P0001  & ~n13153 ;
  assign n13158 = n11798 & ~n11860 ;
  assign n13159 = ~\sa11_reg[5]/P0001  & n13100 ;
  assign n13160 = ~n13158 & ~n13159 ;
  assign n13161 = ~\sa11_reg[2]/P0001  & ~n13160 ;
  assign n13156 = ~n11830 & ~n11907 ;
  assign n13157 = \sa11_reg[2]/P0001  & ~n13156 ;
  assign n13155 = ~\sa11_reg[6]/NET0131  & n11926 ;
  assign n13162 = ~n12124 & ~n13155 ;
  assign n13163 = ~n13157 & n13162 ;
  assign n13164 = ~n13161 & n13163 ;
  assign n13165 = ~\sa11_reg[1]/P0001  & ~n13164 ;
  assign n13171 = \sa11_reg[1]/P0001  & \sa11_reg[2]/P0001  ;
  assign n13173 = \sa11_reg[3]/P0001  & n13102 ;
  assign n13172 = ~\sa11_reg[6]/NET0131  & n11813 ;
  assign n13174 = ~n11865 & ~n13172 ;
  assign n13175 = ~n13173 & n13174 ;
  assign n13176 = n13171 & ~n13175 ;
  assign n13166 = \sa11_reg[1]/P0001  & ~\sa11_reg[2]/P0001  ;
  assign n13167 = n11881 & n13166 ;
  assign n13177 = ~n11866 & ~n13167 ;
  assign n13168 = ~n11795 & ~n12146 ;
  assign n13169 = n12145 & ~n13168 ;
  assign n13170 = \sa11_reg[3]/P0001  & n12160 ;
  assign n13178 = ~n13169 & ~n13170 ;
  assign n13179 = n13177 & n13178 ;
  assign n13180 = ~n13176 & n13179 ;
  assign n13181 = ~n13165 & n13180 ;
  assign n13182 = ~n13154 & n13181 ;
  assign n13183 = ~n13124 & n13182 ;
  assign n13184 = n13091 & ~n13183 ;
  assign n13185 = ~n13091 & n13183 ;
  assign n13186 = ~n13184 & ~n13185 ;
  assign n13187 = ~n12714 & ~n13186 ;
  assign n13188 = n12714 & n13186 ;
  assign n13189 = ~n13187 & ~n13188 ;
  assign n13209 = n12257 & n12385 ;
  assign n13210 = ~n12252 & ~n12268 ;
  assign n13211 = ~n13209 & n13210 ;
  assign n13212 = \sa22_reg[2]/P0001  & ~n13211 ;
  assign n13206 = n12249 & n12303 ;
  assign n13207 = ~n12333 & ~n13206 ;
  assign n13200 = ~\sa22_reg[2]/P0001  & ~\sa22_reg[3]/P0001  ;
  assign n13208 = n12356 & n13200 ;
  assign n13213 = n13207 & ~n13208 ;
  assign n13214 = ~n13212 & n13213 ;
  assign n13215 = \sa22_reg[1]/P0001  & ~n13214 ;
  assign n13197 = ~\sa22_reg[7]/NET0131  & n12257 ;
  assign n13198 = ~n12811 & ~n13197 ;
  assign n13199 = \sa22_reg[2]/P0001  & ~n13198 ;
  assign n13201 = n12332 & n13200 ;
  assign n13202 = ~n12298 & ~n13201 ;
  assign n13203 = ~n12294 & n13202 ;
  assign n13204 = ~n13199 & n13203 ;
  assign n13205 = ~\sa22_reg[1]/P0001  & ~n13204 ;
  assign n13190 = n12251 & n12267 ;
  assign n13191 = ~n12246 & ~n13190 ;
  assign n13192 = ~\sa22_reg[2]/P0001  & ~n13191 ;
  assign n13193 = ~n12320 & ~n12759 ;
  assign n13194 = ~n12296 & ~n12324 ;
  assign n13195 = n13193 & n13194 ;
  assign n13196 = \sa22_reg[2]/P0001  & ~n13195 ;
  assign n13216 = ~n13192 & ~n13196 ;
  assign n13217 = ~n13205 & n13216 ;
  assign n13218 = ~n13215 & n13217 ;
  assign n13219 = \sa22_reg[0]/P0001  & ~n13218 ;
  assign n13220 = \sa22_reg[4]/P0001  & n12249 ;
  assign n13221 = ~n12395 & ~n13220 ;
  assign n13222 = n12322 & ~n13221 ;
  assign n13223 = n12295 & n12779 ;
  assign n13224 = \sa22_reg[1]/P0001  & ~n12384 ;
  assign n13225 = ~n13223 & n13224 ;
  assign n13226 = ~n13222 & n13225 ;
  assign n13231 = ~\sa22_reg[6]/NET0131  & n12258 ;
  assign n13232 = ~n12321 & ~n13231 ;
  assign n13233 = ~\sa22_reg[4]/P0001  & ~n13232 ;
  assign n13229 = n12291 & n12303 ;
  assign n13227 = ~\sa22_reg[2]/P0001  & \sa22_reg[3]/P0001  ;
  assign n13228 = n12297 & n13227 ;
  assign n13234 = ~\sa22_reg[1]/P0001  & ~n13228 ;
  assign n13235 = ~n13229 & n13234 ;
  assign n13230 = \sa22_reg[4]/P0001  & n12259 ;
  assign n13236 = ~n12723 & ~n13230 ;
  assign n13237 = n13235 & n13236 ;
  assign n13238 = ~n13233 & n13237 ;
  assign n13239 = ~n13226 & ~n13238 ;
  assign n13240 = \sa22_reg[4]/P0001  & n12234 ;
  assign n13241 = ~n12716 & ~n13240 ;
  assign n13242 = ~n12260 & ~n13241 ;
  assign n13243 = ~n12393 & n12791 ;
  assign n13244 = ~n13242 & n13243 ;
  assign n13245 = ~\sa22_reg[3]/P0001  & n12295 ;
  assign n13246 = \sa22_reg[2]/P0001  & ~n13230 ;
  assign n13247 = ~n13245 & n13246 ;
  assign n13248 = ~n13244 & ~n13247 ;
  assign n13249 = ~n13239 & ~n13248 ;
  assign n13250 = ~\sa22_reg[0]/P0001  & ~n13249 ;
  assign n13252 = ~\sa22_reg[6]/NET0131  & n12250 ;
  assign n13251 = \sa22_reg[4]/P0001  & n13197 ;
  assign n13253 = ~n12298 & ~n13251 ;
  assign n13254 = ~n13252 & n13253 ;
  assign n13255 = ~\sa22_reg[2]/P0001  & ~n13254 ;
  assign n13258 = n12282 & n12319 ;
  assign n13256 = n12301 & n12735 ;
  assign n13257 = n12263 & n12297 ;
  assign n13259 = ~n12240 & ~n13257 ;
  assign n13260 = ~n13256 & n13259 ;
  assign n13261 = ~n13258 & n13260 ;
  assign n13262 = ~n13255 & n13261 ;
  assign n13263 = ~\sa22_reg[1]/P0001  & ~n13262 ;
  assign n13264 = \sa22_reg[1]/P0001  & \sa22_reg[2]/P0001  ;
  assign n13265 = ~\sa22_reg[3]/P0001  & n12300 ;
  assign n13266 = ~n13252 & ~n13265 ;
  assign n13267 = ~\sa22_reg[4]/P0001  & ~n13266 ;
  assign n13268 = \sa22_reg[4]/P0001  & n12300 ;
  assign n13269 = ~\sa22_reg[5]/P0001  & n13268 ;
  assign n13270 = ~n13267 & ~n13269 ;
  assign n13271 = n13264 & ~n13270 ;
  assign n13272 = n12298 & n13227 ;
  assign n13277 = ~n12280 & ~n13272 ;
  assign n13278 = ~n12717 & n13277 ;
  assign n13273 = n12738 & n13227 ;
  assign n13274 = \sa22_reg[1]/P0001  & n13273 ;
  assign n13275 = n12260 & n13197 ;
  assign n13276 = \sa22_reg[2]/P0001  & n13275 ;
  assign n13279 = ~n13274 & ~n13276 ;
  assign n13280 = n13278 & n13279 ;
  assign n13281 = ~n13271 & n13280 ;
  assign n13282 = ~n13263 & n13281 ;
  assign n13283 = ~n13250 & n13282 ;
  assign n13284 = ~n13219 & n13283 ;
  assign n13285 = \u0_w_reg[0][6]/P0001  & ~n13284 ;
  assign n13286 = ~\u0_w_reg[0][6]/P0001  & n13284 ;
  assign n13287 = ~n13285 & ~n13286 ;
  assign n13288 = n12580 & n13287 ;
  assign n13289 = ~n12580 & ~n13287 ;
  assign n13290 = ~n13288 & ~n13289 ;
  assign n13292 = n13189 & ~n13290 ;
  assign n13291 = ~n13189 & n13290 ;
  assign n13293 = ~\ld_r_reg/P0001  & ~n13291 ;
  assign n13294 = ~n13292 & n13293 ;
  assign n13296 = \text_in_r_reg[102]/P0001  & \u0_w_reg[0][6]/P0001  ;
  assign n13295 = ~\text_in_r_reg[102]/P0001  & ~\u0_w_reg[0][6]/P0001  ;
  assign n13297 = \ld_r_reg/P0001  & ~n13295 ;
  assign n13298 = ~n13296 & n13297 ;
  assign n13299 = ~n13294 & ~n13298 ;
  assign n13304 = ~\sa22_reg[5]/P0001  & n13265 ;
  assign n13305 = ~n12253 & ~n12345 ;
  assign n13306 = ~n13304 & n13305 ;
  assign n13307 = \sa22_reg[2]/P0001  & ~n13306 ;
  assign n13302 = n12773 & n13200 ;
  assign n13300 = \sa22_reg[5]/P0001  & ~n12266 ;
  assign n13301 = n12303 & ~n13300 ;
  assign n13303 = n12238 & n12349 ;
  assign n13308 = ~n13301 & ~n13303 ;
  assign n13309 = ~n13302 & n13308 ;
  assign n13310 = ~n13307 & n13309 ;
  assign n13311 = ~\sa22_reg[1]/P0001  & ~n13310 ;
  assign n13317 = ~n12303 & ~n12319 ;
  assign n13318 = ~n12755 & ~n13317 ;
  assign n13316 = n12244 & n12349 ;
  assign n13319 = ~\sa22_reg[2]/P0001  & ~n12721 ;
  assign n13320 = ~n13316 & n13319 ;
  assign n13321 = ~n13318 & n13320 ;
  assign n13322 = \sa22_reg[2]/P0001  & ~n12756 ;
  assign n13323 = ~n12331 & n13322 ;
  assign n13324 = n13207 & n13323 ;
  assign n13325 = ~n13321 & ~n13324 ;
  assign n13312 = ~\sa22_reg[2]/P0001  & ~n12245 ;
  assign n13313 = ~n12715 & n13312 ;
  assign n13314 = ~n13251 & ~n13313 ;
  assign n13315 = \sa22_reg[1]/P0001  & ~n13314 ;
  assign n13326 = ~n12724 & ~n12747 ;
  assign n13327 = ~n13315 & n13326 ;
  assign n13328 = ~n13325 & n13327 ;
  assign n13329 = ~n13311 & n13328 ;
  assign n13330 = \sa22_reg[0]/P0001  & ~n13329 ;
  assign n13332 = ~n12347 & ~n12795 ;
  assign n13333 = ~\sa22_reg[3]/P0001  & ~n13332 ;
  assign n13334 = n12781 & ~n13333 ;
  assign n13335 = ~n12300 & ~n12811 ;
  assign n13336 = ~n12263 & ~n13335 ;
  assign n13337 = n12321 & n12735 ;
  assign n13338 = n12291 & n13200 ;
  assign n13339 = \sa22_reg[1]/P0001  & ~n12301 ;
  assign n13340 = ~n13338 & n13339 ;
  assign n13341 = ~n13337 & n13340 ;
  assign n13342 = ~n13336 & n13341 ;
  assign n13343 = ~n13334 & ~n13342 ;
  assign n13346 = ~n12257 & ~n12332 ;
  assign n13347 = n12303 & ~n13346 ;
  assign n13344 = ~\sa22_reg[1]/P0001  & n12249 ;
  assign n13345 = ~n12732 & n13344 ;
  assign n13348 = \sa22_reg[2]/P0001  & ~n13345 ;
  assign n13349 = ~n13347 & n13348 ;
  assign n13350 = n12249 & n12732 ;
  assign n13351 = ~n12331 & ~n13350 ;
  assign n13352 = ~\sa22_reg[2]/P0001  & ~n13245 ;
  assign n13353 = n13351 & n13352 ;
  assign n13354 = ~n13349 & ~n13353 ;
  assign n13355 = ~n13343 & ~n13354 ;
  assign n13356 = ~\sa22_reg[0]/P0001  & ~n13355 ;
  assign n13360 = n12244 & n13197 ;
  assign n13361 = ~n12324 & ~n13360 ;
  assign n13362 = \sa22_reg[2]/P0001  & ~n13361 ;
  assign n13358 = n12244 & n12249 ;
  assign n13359 = ~\sa22_reg[2]/P0001  & n13358 ;
  assign n13363 = ~n12717 & ~n13359 ;
  assign n13364 = n12770 & n13363 ;
  assign n13365 = ~n13362 & n13364 ;
  assign n13366 = ~n12240 & n12810 ;
  assign n13367 = ~\sa22_reg[2]/P0001  & ~n12343 ;
  assign n13368 = ~\sa22_reg[3]/P0001  & n12251 ;
  assign n13369 = ~n12267 & n13368 ;
  assign n13370 = ~n12802 & ~n13369 ;
  assign n13371 = n13367 & n13370 ;
  assign n13372 = ~n13366 & ~n13371 ;
  assign n13373 = ~\sa22_reg[1]/P0001  & ~n12382 ;
  assign n13374 = ~n13372 & n13373 ;
  assign n13375 = ~n13365 & ~n13374 ;
  assign n13331 = n12282 & n12747 ;
  assign n13357 = \sa22_reg[6]/NET0131  & n13228 ;
  assign n13376 = ~n13331 & ~n13357 ;
  assign n13377 = ~n13375 & n13376 ;
  assign n13378 = ~n13356 & n13377 ;
  assign n13379 = ~n13330 & n13378 ;
  assign n13413 = \sa11_reg[4]/P0001  & n11858 ;
  assign n13414 = ~n13107 & ~n13413 ;
  assign n13415 = \sa11_reg[7]/NET0131  & ~n13414 ;
  assign n13412 = \sa11_reg[3]/P0001  & n11793 ;
  assign n13416 = ~n11794 & n11829 ;
  assign n13417 = ~n13412 & ~n13416 ;
  assign n13418 = ~n13415 & n13417 ;
  assign n13419 = \sa11_reg[1]/P0001  & ~n13418 ;
  assign n13430 = ~n11854 & ~n11907 ;
  assign n13431 = ~\sa11_reg[3]/P0001  & ~n13430 ;
  assign n13432 = ~n11902 & ~n13431 ;
  assign n13433 = ~\sa11_reg[1]/P0001  & ~n13432 ;
  assign n13420 = \sa11_reg[6]/NET0131  & n12126 ;
  assign n13421 = ~n12176 & ~n13420 ;
  assign n13422 = ~n13133 & n13421 ;
  assign n13423 = ~\sa11_reg[2]/P0001  & ~n13422 ;
  assign n13424 = ~n11816 & ~n11847 ;
  assign n13425 = n11796 & ~n13424 ;
  assign n13426 = ~\sa11_reg[1]/P0001  & ~n11858 ;
  assign n13427 = n11892 & n13426 ;
  assign n13428 = ~n13425 & ~n13427 ;
  assign n13429 = \sa11_reg[2]/P0001  & ~n13428 ;
  assign n13434 = ~n13423 & ~n13429 ;
  assign n13435 = ~n13433 & n13434 ;
  assign n13436 = ~n13419 & n13435 ;
  assign n13437 = ~\sa11_reg[0]/P0001  & ~n13436 ;
  assign n13389 = ~\sa11_reg[5]/P0001  & n11829 ;
  assign n13398 = ~\sa11_reg[3]/P0001  & n13389 ;
  assign n13399 = ~n12129 & ~n12223 ;
  assign n13400 = ~n13398 & n13399 ;
  assign n13401 = \sa11_reg[2]/P0001  & ~n13400 ;
  assign n13394 = ~\sa11_reg[5]/P0001  & n13139 ;
  assign n13395 = n11823 & n13394 ;
  assign n13396 = \sa11_reg[5]/P0001  & ~n11870 ;
  assign n13397 = n11796 & ~n13396 ;
  assign n13402 = ~n11942 & ~n13397 ;
  assign n13403 = ~n13395 & n13402 ;
  assign n13404 = ~n13401 & n13403 ;
  assign n13405 = ~\sa11_reg[1]/P0001  & ~n13404 ;
  assign n13390 = ~\sa11_reg[2]/P0001  & n13389 ;
  assign n13388 = ~\sa11_reg[2]/P0001  & n11833 ;
  assign n13391 = ~n13159 & ~n13388 ;
  assign n13392 = ~n13390 & n13391 ;
  assign n13393 = \sa11_reg[1]/P0001  & ~n13392 ;
  assign n13380 = ~n11802 & ~n13109 ;
  assign n13381 = n12178 & n13380 ;
  assign n13382 = \sa11_reg[2]/P0001  & ~n13381 ;
  assign n13383 = ~n11816 & ~n13092 ;
  assign n13384 = \sa11_reg[3]/P0001  & ~n13383 ;
  assign n13385 = ~n12185 & ~n13126 ;
  assign n13386 = ~n13384 & n13385 ;
  assign n13387 = ~\sa11_reg[2]/P0001  & ~n13386 ;
  assign n13406 = ~n11836 & ~n11872 ;
  assign n13407 = ~n13387 & n13406 ;
  assign n13408 = ~n13382 & n13407 ;
  assign n13409 = ~n13393 & n13408 ;
  assign n13410 = ~n13405 & n13409 ;
  assign n13411 = \sa11_reg[0]/P0001  & ~n13410 ;
  assign n13447 = ~\sa11_reg[3]/P0001  & n12152 ;
  assign n13448 = ~\sa11_reg[2]/P0001  & n13447 ;
  assign n13451 = ~n11866 & ~n11881 ;
  assign n13449 = n12194 & n12206 ;
  assign n13450 = n11846 & n11871 ;
  assign n13452 = ~n13449 & ~n13450 ;
  assign n13453 = n13451 & n13452 ;
  assign n13454 = ~n13448 & n13453 ;
  assign n13455 = \sa11_reg[1]/P0001  & ~n13454 ;
  assign n13441 = ~n11826 & ~n12194 ;
  assign n13442 = ~n13100 & n13441 ;
  assign n13443 = n13106 & ~n13442 ;
  assign n13439 = n11825 & n12188 ;
  assign n13440 = n11853 & n13439 ;
  assign n13444 = ~n12205 & ~n13440 ;
  assign n13445 = ~n13443 & n13444 ;
  assign n13446 = ~\sa11_reg[1]/P0001  & ~n13445 ;
  assign n13438 = \sa11_reg[6]/NET0131  & n13137 ;
  assign n13456 = \sa11_reg[1]/P0001  & ~n12125 ;
  assign n13457 = \sa11_reg[2]/P0001  & n11860 ;
  assign n13458 = ~n11833 & ~n11871 ;
  assign n13459 = n13457 & ~n13458 ;
  assign n13460 = ~n13456 & n13459 ;
  assign n13461 = ~n13438 & ~n13460 ;
  assign n13462 = ~n13446 & n13461 ;
  assign n13463 = ~n13455 & n13462 ;
  assign n13464 = ~n13411 & n13463 ;
  assign n13465 = ~n13437 & n13464 ;
  assign n13466 = n13379 & ~n13465 ;
  assign n13467 = ~n13379 & n13465 ;
  assign n13468 = ~n13466 & ~n13467 ;
  assign n13490 = ~n11853 & ~n12146 ;
  assign n13488 = \sa11_reg[3]/P0001  & n11791 ;
  assign n13489 = \sa11_reg[4]/P0001  & n11876 ;
  assign n13491 = ~n13488 & ~n13489 ;
  assign n13492 = n13490 & n13491 ;
  assign n13493 = \sa11_reg[2]/P0001  & ~n13492 ;
  assign n13487 = n11870 & n13107 ;
  assign n13494 = ~n11859 & ~n13487 ;
  assign n13495 = ~n13493 & n13494 ;
  assign n13496 = \sa11_reg[1]/P0001  & ~n13495 ;
  assign n13469 = ~n13131 & ~n13388 ;
  assign n13470 = ~\sa11_reg[7]/NET0131  & ~n13469 ;
  assign n13473 = n11791 & n13106 ;
  assign n13475 = ~n11924 & ~n13473 ;
  assign n13471 = ~n11797 & n11823 ;
  assign n13472 = ~n11822 & n13471 ;
  assign n13474 = n11801 & n13457 ;
  assign n13476 = ~n13472 & ~n13474 ;
  assign n13477 = n13475 & n13476 ;
  assign n13478 = ~n13470 & n13477 ;
  assign n13479 = ~\sa11_reg[1]/P0001  & ~n13478 ;
  assign n13481 = ~\sa11_reg[5]/P0001  & n11796 ;
  assign n13482 = ~n11861 & ~n13481 ;
  assign n13483 = \sa11_reg[6]/NET0131  & ~n13482 ;
  assign n13484 = ~n12115 & ~n12129 ;
  assign n13485 = ~n13483 & n13484 ;
  assign n13486 = \sa11_reg[2]/P0001  & ~n13485 ;
  assign n13480 = n13100 & n13106 ;
  assign n13497 = ~n13126 & ~n13480 ;
  assign n13498 = ~n13486 & n13497 ;
  assign n13499 = ~n13479 & n13498 ;
  assign n13500 = ~n13496 & n13499 ;
  assign n13501 = \sa11_reg[0]/P0001  & ~n13500 ;
  assign n13530 = n11797 & ~n11886 ;
  assign n13531 = n13430 & ~n13530 ;
  assign n13532 = n12188 & ~n13531 ;
  assign n13533 = \sa11_reg[7]/NET0131  & n11853 ;
  assign n13534 = ~n11826 & ~n13533 ;
  assign n13535 = ~n11883 & n13534 ;
  assign n13536 = ~\sa11_reg[3]/P0001  & ~n13535 ;
  assign n13537 = ~n11925 & ~n12139 ;
  assign n13538 = ~n13536 & n13537 ;
  assign n13539 = \sa11_reg[2]/P0001  & ~n13538 ;
  assign n13540 = ~n13532 & ~n13539 ;
  assign n13541 = \sa11_reg[1]/P0001  & ~n13540 ;
  assign n13503 = n11806 & n11846 ;
  assign n13504 = ~\sa11_reg[1]/P0001  & ~n11832 ;
  assign n13502 = ~\sa11_reg[2]/P0001  & n11886 ;
  assign n13505 = ~n13109 & ~n13502 ;
  assign n13506 = n13504 & n13505 ;
  assign n13507 = ~n13503 & n13506 ;
  assign n13508 = \sa11_reg[2]/P0001  & ~n11936 ;
  assign n13509 = n11791 & n11863 ;
  assign n13510 = ~\sa11_reg[2]/P0001  & ~n11900 ;
  assign n13511 = ~n13509 & n13510 ;
  assign n13512 = ~n13508 & ~n13511 ;
  assign n13513 = \sa11_reg[3]/P0001  & n11798 ;
  assign n13514 = \sa11_reg[1]/P0001  & ~n13132 ;
  assign n13515 = ~n13513 & n13514 ;
  assign n13516 = ~n13512 & n13515 ;
  assign n13517 = ~n13507 & ~n13516 ;
  assign n13518 = ~n11791 & n11794 ;
  assign n13519 = n13396 & n13518 ;
  assign n13520 = \sa11_reg[2]/P0001  & ~n12217 ;
  assign n13521 = ~n13519 & n13520 ;
  assign n13524 = ~\sa11_reg[2]/P0001  & ~n11941 ;
  assign n13522 = ~\sa11_reg[3]/P0001  & n11933 ;
  assign n13523 = ~n11942 & ~n13522 ;
  assign n13525 = ~n13172 & n13523 ;
  assign n13526 = n13524 & n13525 ;
  assign n13527 = ~n13521 & ~n13526 ;
  assign n13528 = ~n13517 & ~n13527 ;
  assign n13529 = ~\sa11_reg[0]/P0001  & ~n13528 ;
  assign n13550 = ~n13138 & ~n13447 ;
  assign n13551 = n13523 & n13550 ;
  assign n13549 = \sa11_reg[2]/P0001  & ~n13447 ;
  assign n13552 = ~\sa11_reg[1]/P0001  & ~n13549 ;
  assign n13553 = ~n13551 & n13552 ;
  assign n13542 = ~n11815 & ~n12125 ;
  assign n13543 = ~\sa11_reg[2]/P0001  & ~n13542 ;
  assign n13544 = ~\sa11_reg[1]/P0001  & \sa11_reg[2]/P0001  ;
  assign n13545 = \sa11_reg[5]/P0001  & n13131 ;
  assign n13546 = ~n11859 & ~n12119 ;
  assign n13547 = ~n13545 & n13546 ;
  assign n13548 = n13544 & ~n13547 ;
  assign n13554 = ~n13543 & ~n13548 ;
  assign n13555 = ~n13553 & n13554 ;
  assign n13556 = ~n13529 & n13555 ;
  assign n13557 = ~n13541 & n13556 ;
  assign n13558 = ~n13501 & n13557 ;
  assign n13593 = n11982 & n11996 ;
  assign n13594 = ~n12624 & ~n13593 ;
  assign n13595 = \sa00_reg[7]/NET0131  & n11979 ;
  assign n13559 = \sa00_reg[4]/P0001  & n12035 ;
  assign n13596 = ~n12090 & ~n13559 ;
  assign n13597 = ~n13595 & n13596 ;
  assign n13598 = \sa00_reg[2]/P0001  & ~n13597 ;
  assign n13599 = n13594 & ~n13598 ;
  assign n13600 = \sa00_reg[1]/P0001  & ~n13599 ;
  assign n13611 = ~n12066 & ~n13069 ;
  assign n13575 = ~\sa00_reg[3]/P0001  & n12651 ;
  assign n13610 = \sa00_reg[4]/P0001  & n11967 ;
  assign n13612 = ~n13575 & ~n13610 ;
  assign n13613 = n13611 & n13612 ;
  assign n13614 = ~\sa00_reg[2]/P0001  & ~n13613 ;
  assign n13601 = ~n12693 & ~n13044 ;
  assign n13602 = n11952 & ~n13601 ;
  assign n13603 = n11982 & ~n12002 ;
  assign n13604 = ~n12064 & n13603 ;
  assign n13605 = ~n12066 & ~n13604 ;
  assign n13606 = ~n13602 & n13605 ;
  assign n13607 = ~\sa00_reg[1]/P0001  & ~n13606 ;
  assign n13609 = \sa00_reg[2]/P0001  & n12033 ;
  assign n13608 = ~\sa00_reg[6]/NET0131  & n13031 ;
  assign n13615 = ~n13037 & ~n13608 ;
  assign n13616 = ~n13609 & n13615 ;
  assign n13617 = ~n13607 & n13616 ;
  assign n13618 = ~n13614 & n13617 ;
  assign n13619 = ~n13600 & n13618 ;
  assign n13620 = \sa00_reg[0]/P0001  & ~n13619 ;
  assign n13578 = ~n12997 & ~n13068 ;
  assign n13579 = ~\sa00_reg[2]/P0001  & ~n13578 ;
  assign n13580 = n11979 & n12064 ;
  assign n13581 = \sa00_reg[4]/P0001  & n13580 ;
  assign n13582 = ~n12034 & ~n13581 ;
  assign n13583 = ~n13579 & n13582 ;
  assign n13584 = ~\sa00_reg[1]/P0001  & ~n13583 ;
  assign n13560 = \sa00_reg[3]/P0001  & n13559 ;
  assign n13561 = ~n12629 & ~n13042 ;
  assign n13562 = ~n13560 & n13561 ;
  assign n13563 = ~\sa00_reg[2]/P0001  & ~n13562 ;
  assign n13564 = ~n12611 & n12653 ;
  assign n13565 = ~n13563 & n13564 ;
  assign n13566 = \sa00_reg[1]/P0001  & ~n13565 ;
  assign n13585 = ~n12691 & ~n12702 ;
  assign n13567 = ~n11957 & ~n12007 ;
  assign n13568 = n12056 & ~n13567 ;
  assign n13569 = ~n11980 & ~n12600 ;
  assign n13570 = n11985 & ~n13569 ;
  assign n13586 = ~n13568 & ~n13570 ;
  assign n13587 = n13585 & n13586 ;
  assign n13571 = \sa00_reg[1]/P0001  & \sa00_reg[2]/P0001  ;
  assign n13572 = ~\sa00_reg[3]/P0001  & n11996 ;
  assign n13573 = ~n12632 & ~n13572 ;
  assign n13574 = n13571 & ~n13573 ;
  assign n13576 = ~n12003 & ~n13575 ;
  assign n13577 = n13015 & ~n13576 ;
  assign n13588 = ~n13574 & ~n13577 ;
  assign n13589 = n13587 & n13588 ;
  assign n13590 = ~n13566 & n13589 ;
  assign n13591 = ~n13584 & n13590 ;
  assign n13592 = ~\sa00_reg[0]/P0001  & ~n13591 ;
  assign n13635 = ~\sa00_reg[5]/P0001  & n13042 ;
  assign n13636 = \sa00_reg[2]/P0001  & ~n12691 ;
  assign n13637 = ~n12647 & n13636 ;
  assign n13638 = ~n13635 & n13637 ;
  assign n13639 = ~\sa00_reg[2]/P0001  & ~n13580 ;
  assign n13640 = ~n11958 & ~n13012 ;
  assign n13641 = n13639 & n13640 ;
  assign n13642 = ~n13638 & ~n13641 ;
  assign n13643 = ~n12025 & ~n12667 ;
  assign n13644 = ~n13642 & n13643 ;
  assign n13645 = ~\sa00_reg[1]/P0001  & ~n13644 ;
  assign n13621 = ~n12068 & ~n12624 ;
  assign n13622 = \sa00_reg[3]/P0001  & ~n13621 ;
  assign n13623 = ~n13037 & ~n13622 ;
  assign n13624 = n13571 & ~n13623 ;
  assign n13625 = \sa00_reg[2]/P0001  & n12025 ;
  assign n13626 = ~n12630 & ~n13625 ;
  assign n13627 = n12054 & ~n13626 ;
  assign n13628 = ~n12659 & ~n13627 ;
  assign n13629 = ~\sa00_reg[3]/P0001  & n11975 ;
  assign n13630 = ~n11959 & n13629 ;
  assign n13631 = ~n12611 & ~n13006 ;
  assign n13632 = ~n13630 & n13631 ;
  assign n13633 = n13626 & n13632 ;
  assign n13634 = ~n13628 & ~n13633 ;
  assign n13646 = ~n13624 & ~n13634 ;
  assign n13647 = ~n13645 & n13646 ;
  assign n13648 = ~n13592 & n13647 ;
  assign n13649 = ~n13620 & n13648 ;
  assign n13650 = n13558 & ~n13649 ;
  assign n13651 = ~n13558 & n13649 ;
  assign n13652 = ~n13650 & ~n13651 ;
  assign n13653 = n13468 & n13652 ;
  assign n13654 = ~n13468 & ~n13652 ;
  assign n13655 = ~n13653 & ~n13654 ;
  assign n13689 = ~\sa33_reg[5]/P0001  & ~n12460 ;
  assign n13690 = \sa33_reg[4]/P0001  & ~n12877 ;
  assign n13691 = n13689 & ~n13690 ;
  assign n13692 = ~n12470 & ~n13691 ;
  assign n13693 = ~\sa33_reg[2]/P0001  & ~n13692 ;
  assign n13685 = \sa33_reg[4]/P0001  & n12418 ;
  assign n13686 = ~\sa33_reg[3]/P0001  & n12481 ;
  assign n13687 = ~n13685 & ~n13686 ;
  assign n13688 = \sa33_reg[2]/P0001  & ~n13687 ;
  assign n13694 = ~n12428 & ~n12532 ;
  assign n13695 = ~n13688 & n13694 ;
  assign n13696 = ~n13693 & n13695 ;
  assign n13697 = \sa33_reg[1]/P0001  & ~n13696 ;
  assign n13698 = n12414 & n12457 ;
  assign n13699 = n12521 & n12551 ;
  assign n13700 = ~n13698 & ~n13699 ;
  assign n13701 = ~\sa33_reg[2]/P0001  & ~n13700 ;
  assign n13702 = n12472 & n12499 ;
  assign n13705 = ~n12919 & ~n13702 ;
  assign n13703 = n12413 & n12560 ;
  assign n13704 = n12458 & n12877 ;
  assign n13706 = ~n13703 & ~n13704 ;
  assign n13707 = n13705 & n13706 ;
  assign n13708 = ~n13701 & n13707 ;
  assign n13709 = ~\sa33_reg[1]/P0001  & ~n13708 ;
  assign n13712 = ~n12507 & ~n12919 ;
  assign n13713 = ~\sa33_reg[2]/P0001  & ~n13712 ;
  assign n13710 = ~n12444 & ~n12473 ;
  assign n13711 = n12472 & ~n13710 ;
  assign n13714 = ~n12549 & ~n12563 ;
  assign n13715 = ~n13711 & n13714 ;
  assign n13716 = ~n13713 & n13715 ;
  assign n13717 = ~n13709 & n13716 ;
  assign n13718 = ~n13697 & n13717 ;
  assign n13719 = ~\sa33_reg[0]/P0001  & ~n13718 ;
  assign n13657 = \sa33_reg[6]/P0001  & n12457 ;
  assign n13658 = ~n12446 & ~n12877 ;
  assign n13659 = \sa33_reg[7]/NET0131  & ~n13658 ;
  assign n13660 = ~n13657 & ~n13659 ;
  assign n13661 = \sa33_reg[2]/P0001  & ~n13660 ;
  assign n13662 = n12418 & n12877 ;
  assign n13663 = \sa33_reg[4]/P0001  & n13662 ;
  assign n13664 = ~n12462 & ~n13663 ;
  assign n13665 = ~n13661 & n13664 ;
  assign n13666 = \sa33_reg[1]/P0001  & ~n13665 ;
  assign n13675 = n12410 & n12470 ;
  assign n13674 = n12432 & ~n12855 ;
  assign n13676 = ~n12511 & ~n12906 ;
  assign n13677 = ~n13674 & n13676 ;
  assign n13678 = ~n13675 & n13677 ;
  assign n13679 = ~\sa33_reg[1]/P0001  & ~n13678 ;
  assign n13669 = ~n12906 & ~n12927 ;
  assign n13667 = \sa33_reg[4]/P0001  & n12561 ;
  assign n13668 = ~\sa33_reg[6]/P0001  & n12421 ;
  assign n13670 = ~n13667 & ~n13668 ;
  assign n13671 = n13669 & n13670 ;
  assign n13672 = ~\sa33_reg[2]/P0001  & ~n13671 ;
  assign n13656 = n12564 & ~n12884 ;
  assign n13673 = n12448 & n12561 ;
  assign n13680 = ~n13656 & ~n13673 ;
  assign n13681 = ~n13672 & n13680 ;
  assign n13682 = ~n13679 & n13681 ;
  assign n13683 = ~n13666 & n13682 ;
  assign n13684 = \sa33_reg[0]/P0001  & ~n13683 ;
  assign n13721 = ~\sa33_reg[4]/P0001  & n12421 ;
  assign n13720 = n12414 & n12426 ;
  assign n13722 = ~n12508 & ~n13720 ;
  assign n13723 = ~n13721 & n13722 ;
  assign n13724 = ~\sa33_reg[2]/P0001  & ~n13723 ;
  assign n13725 = ~n12512 & ~n12914 ;
  assign n13726 = ~n13724 & n13725 ;
  assign n13727 = ~\sa33_reg[1]/P0001  & ~n13726 ;
  assign n13733 = ~n12462 & ~n12932 ;
  assign n13734 = \sa33_reg[3]/P0001  & ~n13733 ;
  assign n13735 = \sa33_reg[2]/P0001  & ~n12929 ;
  assign n13736 = ~n13734 & n13735 ;
  assign n13729 = ~n12448 & n12473 ;
  assign n13728 = n12430 & ~n12467 ;
  assign n13730 = ~\sa33_reg[2]/P0001  & ~n12415 ;
  assign n13731 = ~n13728 & n13730 ;
  assign n13732 = ~n13729 & n13731 ;
  assign n13737 = \sa33_reg[1]/P0001  & ~n13732 ;
  assign n13738 = ~n13736 & n13737 ;
  assign n13741 = ~\sa33_reg[1]/P0001  & \sa33_reg[2]/P0001  ;
  assign n13742 = ~n12445 & ~n12544 ;
  assign n13743 = ~\sa33_reg[3]/P0001  & ~n13742 ;
  assign n13744 = ~n12501 & ~n13743 ;
  assign n13745 = n13741 & ~n13744 ;
  assign n13739 = n12544 & n12560 ;
  assign n13740 = \sa33_reg[4]/P0001  & n13739 ;
  assign n13746 = ~\sa33_reg[7]/NET0131  & n12478 ;
  assign n13747 = ~n13740 & ~n13746 ;
  assign n13748 = ~n13745 & n13747 ;
  assign n13749 = ~n13738 & n13748 ;
  assign n13750 = ~n13727 & n13749 ;
  assign n13751 = ~n13684 & n13750 ;
  assign n13752 = ~n13719 & n13751 ;
  assign n13755 = ~n13209 & ~n13251 ;
  assign n13756 = ~\sa22_reg[2]/P0001  & ~n13755 ;
  assign n13754 = ~\sa22_reg[3]/P0001  & n12760 ;
  assign n13757 = ~\sa22_reg[1]/P0001  & ~n12806 ;
  assign n13753 = \sa22_reg[2]/P0001  & n12790 ;
  assign n13758 = ~n13275 & ~n13753 ;
  assign n13759 = n13757 & n13758 ;
  assign n13760 = ~n13754 & n13759 ;
  assign n13761 = ~n13756 & n13760 ;
  assign n13766 = ~\sa22_reg[3]/P0001  & n12319 ;
  assign n13767 = ~n13220 & ~n13766 ;
  assign n13768 = \sa22_reg[2]/P0001  & ~n13767 ;
  assign n13762 = \sa22_reg[4]/P0001  & n12721 ;
  assign n13763 = ~n12295 & ~n13231 ;
  assign n13764 = ~n13762 & n13763 ;
  assign n13765 = ~\sa22_reg[2]/P0001  & ~n13764 ;
  assign n13769 = n12237 & n12354 ;
  assign n13770 = ~n13765 & n13769 ;
  assign n13771 = ~n13768 & n13770 ;
  assign n13772 = ~n13761 & ~n13771 ;
  assign n13773 = ~n12331 & ~n12371 ;
  assign n13774 = n12807 & n13773 ;
  assign n13775 = \sa22_reg[2]/P0001  & ~n12242 ;
  assign n13776 = ~n13304 & n13775 ;
  assign n13777 = ~n13774 & ~n13776 ;
  assign n13778 = ~n12382 & ~n13777 ;
  assign n13779 = ~n13772 & n13778 ;
  assign n13780 = ~\sa22_reg[0]/P0001  & ~n13779 ;
  assign n13798 = ~n12296 & ~n12330 ;
  assign n13799 = ~n12297 & ~n13798 ;
  assign n13800 = ~n12236 & ~n13190 ;
  assign n13801 = ~n13799 & n13800 ;
  assign n13802 = ~\sa22_reg[2]/P0001  & ~n13801 ;
  assign n13803 = \sa22_reg[6]/NET0131  & n12262 ;
  assign n13804 = ~n12292 & ~n13803 ;
  assign n13806 = \sa22_reg[4]/P0001  & n12257 ;
  assign n13805 = ~\sa22_reg[5]/P0001  & n12755 ;
  assign n13807 = ~n12805 & ~n13805 ;
  assign n13808 = ~n13806 & n13807 ;
  assign n13809 = \sa22_reg[2]/P0001  & ~n13808 ;
  assign n13810 = n13804 & ~n13809 ;
  assign n13811 = \sa22_reg[0]/P0001  & ~n13810 ;
  assign n13812 = ~n13802 & ~n13811 ;
  assign n13813 = \sa22_reg[1]/P0001  & ~n13812 ;
  assign n13787 = n12264 & ~n12282 ;
  assign n13786 = n12238 & n12753 ;
  assign n13788 = ~n12381 & ~n13786 ;
  assign n13789 = ~n13787 & n13788 ;
  assign n13790 = ~\sa22_reg[1]/P0001  & ~n13789 ;
  assign n13782 = \sa22_reg[5]/P0001  & n13268 ;
  assign n13783 = ~n12747 & ~n13252 ;
  assign n13784 = ~n13782 & n13783 ;
  assign n13785 = ~\sa22_reg[2]/P0001  & ~n13784 ;
  assign n13781 = \sa22_reg[4]/P0001  & n12813 ;
  assign n13791 = n12347 & ~n13264 ;
  assign n13792 = n12259 & ~n12731 ;
  assign n13793 = ~n13791 & ~n13792 ;
  assign n13794 = ~n13781 & n13793 ;
  assign n13795 = ~n13785 & n13794 ;
  assign n13796 = ~n13790 & n13795 ;
  assign n13797 = \sa22_reg[0]/P0001  & ~n13796 ;
  assign n13824 = ~n12733 & ~n13206 ;
  assign n13825 = ~n12335 & n13824 ;
  assign n13826 = ~\sa22_reg[2]/P0001  & ~n13825 ;
  assign n13827 = ~n12333 & ~n12812 ;
  assign n13828 = ~n13826 & n13827 ;
  assign n13829 = ~\sa22_reg[1]/P0001  & ~n13828 ;
  assign n13820 = ~\sa22_reg[1]/P0001  & \sa22_reg[2]/P0001  ;
  assign n13821 = ~n12275 & ~n12320 ;
  assign n13822 = ~n12371 & n13821 ;
  assign n13823 = n13820 & ~n13822 ;
  assign n13814 = ~n12292 & ~n12736 ;
  assign n13815 = \sa22_reg[3]/P0001  & ~n13814 ;
  assign n13816 = ~n13230 & ~n13815 ;
  assign n13817 = n13264 & ~n13816 ;
  assign n13818 = ~n12396 & ~n12812 ;
  assign n13819 = \sa22_reg[2]/P0001  & ~n13818 ;
  assign n13830 = ~n13817 & ~n13819 ;
  assign n13831 = ~n13823 & n13830 ;
  assign n13832 = ~n13829 & n13831 ;
  assign n13833 = ~n13797 & n13832 ;
  assign n13834 = ~n13813 & n13833 ;
  assign n13835 = ~n13780 & n13834 ;
  assign n13836 = n13752 & ~n13835 ;
  assign n13837 = ~n13752 & n13835 ;
  assign n13838 = ~n13836 & ~n13837 ;
  assign n13875 = ~n12290 & ~n12352 ;
  assign n13876 = ~n13240 & ~n13265 ;
  assign n13877 = n13875 & n13876 ;
  assign n13878 = \sa22_reg[2]/P0001  & ~n13877 ;
  assign n13879 = ~\sa22_reg[2]/P0001  & n12275 ;
  assign n13880 = ~n12722 & ~n13879 ;
  assign n13881 = ~n13878 & n13880 ;
  assign n13882 = \sa22_reg[1]/P0001  & ~n13881 ;
  assign n13866 = n12239 & ~n12755 ;
  assign n13867 = ~n12252 & ~n13240 ;
  assign n13868 = ~n13866 & n13867 ;
  assign n13869 = ~\sa22_reg[2]/P0001  & ~n13868 ;
  assign n13870 = ~n12282 & n13368 ;
  assign n13865 = n12322 & n13805 ;
  assign n13871 = ~n12814 & ~n13865 ;
  assign n13872 = ~n13870 & n13871 ;
  assign n13873 = ~n13869 & n13872 ;
  assign n13874 = ~\sa22_reg[1]/P0001  & ~n13873 ;
  assign n13883 = \sa22_reg[6]/NET0131  & n12385 ;
  assign n13884 = n12257 & n12303 ;
  assign n13885 = ~n12246 & ~n13884 ;
  assign n13886 = ~n12253 & n13885 ;
  assign n13887 = ~n13883 & n13886 ;
  assign n13888 = \sa22_reg[2]/P0001  & ~n13887 ;
  assign n13889 = n12252 & n13200 ;
  assign n13890 = ~n13316 & ~n13889 ;
  assign n13891 = ~n13888 & n13890 ;
  assign n13892 = ~n13874 & n13891 ;
  assign n13893 = ~n13882 & n13892 ;
  assign n13894 = \sa22_reg[0]/P0001  & ~n13893 ;
  assign n13846 = ~n12315 & ~n12733 ;
  assign n13847 = ~\sa22_reg[2]/P0001  & ~n13846 ;
  assign n13844 = n12244 & n12257 ;
  assign n13845 = ~n12779 & n13844 ;
  assign n13848 = \sa22_reg[1]/P0001  & ~n13252 ;
  assign n13849 = ~n13845 & n13848 ;
  assign n13850 = ~n13847 & n13849 ;
  assign n13851 = n12344 & n12735 ;
  assign n13853 = ~\sa22_reg[1]/P0001  & ~n12279 ;
  assign n13852 = ~\sa22_reg[2]/P0001  & n12755 ;
  assign n13854 = ~n13206 & ~n13852 ;
  assign n13855 = n13853 & n13854 ;
  assign n13856 = ~n13851 & n13855 ;
  assign n13857 = ~n13850 & ~n13856 ;
  assign n13839 = n12239 & n12297 ;
  assign n13840 = ~n13782 & ~n13839 ;
  assign n13841 = \sa22_reg[3]/P0001  & ~n13840 ;
  assign n13842 = ~n12396 & ~n13841 ;
  assign n13843 = \sa22_reg[2]/P0001  & ~n13842 ;
  assign n13858 = ~n13303 & ~n13766 ;
  assign n13859 = ~n12384 & ~n13269 ;
  assign n13860 = n13858 & n13859 ;
  assign n13861 = ~\sa22_reg[2]/P0001  & ~n13860 ;
  assign n13862 = ~n13843 & ~n13861 ;
  assign n13863 = ~n13857 & n13862 ;
  assign n13864 = ~\sa22_reg[0]/P0001  & ~n13863 ;
  assign n13895 = n12245 & ~n12755 ;
  assign n13896 = n13332 & ~n13895 ;
  assign n13897 = n13227 & ~n13896 ;
  assign n13898 = \sa22_reg[7]/NET0131  & n12290 ;
  assign n13899 = ~n12738 & ~n12773 ;
  assign n13900 = ~n13898 & n13899 ;
  assign n13901 = ~\sa22_reg[3]/P0001  & ~n13900 ;
  assign n13902 = ~n12292 & ~n12351 ;
  assign n13903 = ~n13901 & n13902 ;
  assign n13904 = \sa22_reg[2]/P0001  & ~n13903 ;
  assign n13905 = ~n13897 & ~n13904 ;
  assign n13906 = \sa22_reg[1]/P0001  & ~n13905 ;
  assign n13907 = ~n13229 & n13858 ;
  assign n13908 = ~\sa22_reg[2]/P0001  & ~n13907 ;
  assign n13909 = ~n13358 & ~n13908 ;
  assign n13910 = ~\sa22_reg[1]/P0001  & ~n13909 ;
  assign n13911 = n12234 & n12260 ;
  assign n13912 = ~n12240 & ~n13911 ;
  assign n13913 = n12779 & ~n13912 ;
  assign n13914 = n12239 & n12244 ;
  assign n13915 = ~n12236 & ~n13914 ;
  assign n13916 = ~n12722 & n13915 ;
  assign n13917 = n13820 & ~n13916 ;
  assign n13918 = ~n13913 & ~n13917 ;
  assign n13919 = ~n13910 & n13918 ;
  assign n13920 = ~n13906 & n13919 ;
  assign n13921 = ~n13864 & n13920 ;
  assign n13922 = ~n13894 & n13921 ;
  assign n13923 = \u0_w_reg[0][17]/P0001  & ~n13922 ;
  assign n13924 = ~\u0_w_reg[0][17]/P0001  & n13922 ;
  assign n13925 = ~n13923 & ~n13924 ;
  assign n13926 = n13838 & n13925 ;
  assign n13927 = ~n13838 & ~n13925 ;
  assign n13928 = ~n13926 & ~n13927 ;
  assign n13930 = ~n13655 & n13928 ;
  assign n13929 = n13655 & ~n13928 ;
  assign n13931 = ~\ld_r_reg/P0001  & ~n13929 ;
  assign n13932 = ~n13930 & n13931 ;
  assign n13934 = \text_in_r_reg[113]/P0001  & \u0_w_reg[0][17]/P0001  ;
  assign n13933 = ~\text_in_r_reg[113]/P0001  & ~\u0_w_reg[0][17]/P0001  ;
  assign n13935 = \ld_r_reg/P0001  & ~n13933 ;
  assign n13936 = ~n13934 & n13935 ;
  assign n13937 = ~n13932 & ~n13936 ;
  assign n13970 = \sa33_reg[4]/P0001  & n12475 ;
  assign n13985 = ~n12460 & ~n13970 ;
  assign n13986 = ~\sa33_reg[3]/P0001  & n12465 ;
  assign n13987 = ~n12531 & ~n13986 ;
  assign n13988 = n13985 & n13987 ;
  assign n13989 = \sa33_reg[1]/P0001  & ~n13988 ;
  assign n13990 = \sa33_reg[6]/P0001  & n12551 ;
  assign n13991 = ~n12423 & ~n12431 ;
  assign n13992 = ~n13990 & n13991 ;
  assign n13993 = ~n13989 & n13992 ;
  assign n13994 = \sa33_reg[2]/P0001  & ~n13993 ;
  assign n13971 = n12480 & ~n12876 ;
  assign n13972 = ~n12422 & ~n13970 ;
  assign n13973 = ~n13971 & n13972 ;
  assign n13974 = ~\sa33_reg[2]/P0001  & ~n13973 ;
  assign n13938 = \sa33_reg[2]/P0001  & ~\sa33_reg[5]/P0001  ;
  assign n13969 = n12551 & n13938 ;
  assign n13968 = n12433 & ~n12855 ;
  assign n13975 = ~n12565 & ~n13968 ;
  assign n13976 = ~n13969 & n13975 ;
  assign n13977 = ~n13974 & n13976 ;
  assign n13978 = ~\sa33_reg[1]/P0001  & ~n13977 ;
  assign n13952 = ~\sa33_reg[2]/P0001  & ~\sa33_reg[3]/P0001  ;
  assign n13980 = n12461 & n13952 ;
  assign n13981 = ~\sa33_reg[6]/P0001  & n13980 ;
  assign n13982 = ~n12900 & ~n13981 ;
  assign n13983 = \sa33_reg[1]/P0001  & ~n13982 ;
  assign n13984 = n12477 & n12521 ;
  assign n13979 = n12422 & n13952 ;
  assign n13995 = ~n12569 & ~n13979 ;
  assign n13996 = ~n13984 & n13995 ;
  assign n13997 = ~n13983 & n13996 ;
  assign n13998 = ~n13978 & n13997 ;
  assign n13999 = ~n13994 & n13998 ;
  assign n14000 = \sa33_reg[0]/P0001  & ~n13999 ;
  assign n13956 = ~n12880 & ~n13720 ;
  assign n13957 = ~\sa33_reg[2]/P0001  & ~n13956 ;
  assign n13955 = n12450 & ~n12881 ;
  assign n13958 = ~n13668 & ~n13955 ;
  assign n13959 = ~n13957 & n13958 ;
  assign n13960 = \sa33_reg[1]/P0001  & ~n13959 ;
  assign n13939 = \sa33_reg[3]/P0001  & n12467 ;
  assign n13940 = ~n12465 & ~n13939 ;
  assign n13941 = n13938 & ~n13940 ;
  assign n13942 = ~n13721 & ~n13941 ;
  assign n13943 = ~\sa33_reg[1]/P0001  & ~n13942 ;
  assign n13953 = ~n12481 & ~n12525 ;
  assign n13954 = n13952 & ~n13953 ;
  assign n13947 = ~\sa33_reg[1]/P0001  & ~\sa33_reg[2]/P0001  ;
  assign n13948 = n12876 & n13947 ;
  assign n13961 = ~n13746 & ~n13948 ;
  assign n13962 = ~n13954 & n13961 ;
  assign n13944 = \sa33_reg[7]/NET0131  & n12932 ;
  assign n13945 = ~n13667 & ~n13944 ;
  assign n13946 = n12560 & ~n13945 ;
  assign n13949 = n12457 & n12465 ;
  assign n13950 = ~n12550 & ~n13949 ;
  assign n13951 = ~\sa33_reg[2]/P0001  & ~n13950 ;
  assign n13963 = ~n13946 & ~n13951 ;
  assign n13964 = n13962 & n13963 ;
  assign n13965 = ~n13943 & n13964 ;
  assign n13966 = ~n13960 & n13965 ;
  assign n13967 = ~\sa33_reg[0]/P0001  & ~n13966 ;
  assign n14021 = \sa33_reg[1]/P0001  & \sa33_reg[2]/P0001  ;
  assign n14022 = \sa33_reg[7]/NET0131  & ~n13985 ;
  assign n14023 = n12429 & n12444 ;
  assign n14024 = ~n14022 & ~n14023 ;
  assign n14025 = ~\sa33_reg[3]/P0001  & ~n14024 ;
  assign n14026 = ~n12462 & ~n12913 ;
  assign n14027 = ~n14025 & n14026 ;
  assign n14028 = n14021 & ~n14027 ;
  assign n14001 = n12448 & n12480 ;
  assign n14002 = ~n12428 & ~n14001 ;
  assign n14003 = ~n12900 & n14002 ;
  assign n14004 = \sa33_reg[2]/P0001  & ~n14003 ;
  assign n14005 = \sa33_reg[3]/P0001  & n12461 ;
  assign n14006 = n12884 & n14005 ;
  assign n14007 = ~n12506 & ~n14006 ;
  assign n14008 = ~n13954 & n14007 ;
  assign n14009 = ~n14004 & n14008 ;
  assign n14010 = ~\sa33_reg[1]/P0001  & ~n14009 ;
  assign n14011 = n12479 & n12480 ;
  assign n14012 = n12419 & n12475 ;
  assign n14013 = ~n14011 & ~n14012 ;
  assign n14014 = n12881 & ~n14013 ;
  assign n14015 = n12429 & ~n12876 ;
  assign n14016 = n12480 & n12876 ;
  assign n14017 = ~n12906 & ~n14016 ;
  assign n14018 = ~n14015 & n14017 ;
  assign n14019 = \sa33_reg[1]/P0001  & n12456 ;
  assign n14020 = ~n14018 & n14019 ;
  assign n14029 = ~n14014 & ~n14020 ;
  assign n14030 = ~n14010 & n14029 ;
  assign n14031 = ~n14028 & n14030 ;
  assign n14032 = ~n13967 & n14031 ;
  assign n14033 = ~n14000 & n14032 ;
  assign n14053 = ~n12423 & ~n12522 ;
  assign n14054 = \sa33_reg[2]/P0001  & ~n14053 ;
  assign n14048 = n12448 & n12942 ;
  assign n14049 = \sa33_reg[2]/P0001  & n13986 ;
  assign n14050 = ~n14048 & ~n14049 ;
  assign n14051 = ~\sa33_reg[5]/P0001  & ~n14050 ;
  assign n14052 = n12479 & n12510 ;
  assign n14055 = ~n12447 & ~n12509 ;
  assign n14056 = ~n14052 & n14055 ;
  assign n14057 = ~n14051 & n14056 ;
  assign n14058 = ~n14054 & n14057 ;
  assign n14059 = ~\sa33_reg[1]/P0001  & ~n14058 ;
  assign n14043 = ~n12512 & ~n13721 ;
  assign n14044 = n12475 & n12876 ;
  assign n14045 = ~n12507 & ~n14044 ;
  assign n14046 = n14043 & n14045 ;
  assign n14047 = \sa33_reg[2]/P0001  & ~n14046 ;
  assign n14041 = ~n12569 & ~n13944 ;
  assign n14042 = ~\sa33_reg[2]/P0001  & ~n14041 ;
  assign n14034 = ~\sa33_reg[2]/P0001  & ~n12429 ;
  assign n14035 = ~\sa33_reg[5]/P0001  & ~n12465 ;
  assign n14036 = n14034 & ~n14035 ;
  assign n14037 = ~n13698 & ~n14036 ;
  assign n14038 = \sa33_reg[1]/P0001  & ~n14037 ;
  assign n14039 = ~n12444 & ~n12521 ;
  assign n14040 = n12456 & ~n14039 ;
  assign n14060 = ~n12899 & ~n12927 ;
  assign n14061 = ~n14040 & n14060 ;
  assign n14062 = ~n14038 & n14061 ;
  assign n14063 = ~n14042 & n14062 ;
  assign n14064 = ~n14047 & n14063 ;
  assign n14065 = ~n14059 & n14064 ;
  assign n14066 = \sa33_reg[0]/P0001  & ~n14065 ;
  assign n14079 = \sa33_reg[2]/P0001  & n12913 ;
  assign n14080 = \sa33_reg[1]/P0001  & ~n13980 ;
  assign n14077 = n12412 & n12419 ;
  assign n14078 = ~n12419 & n12465 ;
  assign n14081 = ~n14077 & ~n14078 ;
  assign n14082 = n14080 & n14081 ;
  assign n14083 = ~n14079 & n14082 ;
  assign n14084 = ~\sa33_reg[3]/P0001  & ~n14017 ;
  assign n14085 = ~\sa33_reg[1]/P0001  & ~n12882 ;
  assign n14086 = ~n14084 & n14085 ;
  assign n14087 = ~n14083 & ~n14086 ;
  assign n14067 = ~n12521 & ~n12561 ;
  assign n14068 = n12476 & ~n14067 ;
  assign n14069 = ~\sa33_reg[1]/P0001  & n12418 ;
  assign n14070 = ~n12877 & n14069 ;
  assign n14071 = ~n14068 & ~n14070 ;
  assign n14072 = \sa33_reg[2]/P0001  & ~n14071 ;
  assign n14073 = n12475 & n12479 ;
  assign n14074 = ~n12507 & ~n13662 ;
  assign n14075 = ~n14073 & n14074 ;
  assign n14076 = ~\sa33_reg[2]/P0001  & ~n14075 ;
  assign n14088 = ~n14072 & ~n14076 ;
  assign n14089 = ~n14087 & n14088 ;
  assign n14090 = ~\sa33_reg[0]/P0001  & ~n14089 ;
  assign n14091 = ~\sa33_reg[2]/P0001  & n13939 ;
  assign n14092 = n12472 & n12525 ;
  assign n14093 = ~n14091 & ~n14092 ;
  assign n14094 = \sa33_reg[6]/P0001  & ~n14093 ;
  assign n14095 = n13685 & n13952 ;
  assign n14097 = ~n12863 & ~n13739 ;
  assign n14098 = ~n14095 & n14097 ;
  assign n14096 = ~\sa33_reg[5]/P0001  & n12898 ;
  assign n14099 = n12871 & ~n14096 ;
  assign n14100 = n14098 & n14099 ;
  assign n14101 = n12911 & ~n14011 ;
  assign n14102 = ~n12410 & n12433 ;
  assign n14103 = ~\sa33_reg[2]/P0001  & ~n12909 ;
  assign n14104 = ~n14102 & n14103 ;
  assign n14105 = ~n14101 & ~n14104 ;
  assign n14106 = n12415 & n12456 ;
  assign n14107 = ~\sa33_reg[1]/P0001  & ~n14106 ;
  assign n14108 = ~n12563 & n14107 ;
  assign n14109 = ~n14105 & n14108 ;
  assign n14110 = ~n14100 & ~n14109 ;
  assign n14111 = ~n14094 & ~n14110 ;
  assign n14112 = ~n14090 & n14111 ;
  assign n14113 = ~n14066 & n14112 ;
  assign n14114 = n14033 & ~n14113 ;
  assign n14115 = ~n14033 & n14113 ;
  assign n14116 = ~n14114 & ~n14115 ;
  assign n14117 = \u0_w_reg[0][9]/P0001  & ~n13752 ;
  assign n14118 = ~\u0_w_reg[0][9]/P0001  & n13752 ;
  assign n14119 = ~n14117 & ~n14118 ;
  assign n14120 = n14116 & n14119 ;
  assign n14121 = ~n14116 & ~n14119 ;
  assign n14122 = ~n14120 & ~n14121 ;
  assign n14123 = n13379 & ~n13922 ;
  assign n14124 = ~n13379 & n13922 ;
  assign n14125 = ~n14123 & ~n14124 ;
  assign n14139 = ~n13101 & ~n13159 ;
  assign n14140 = ~\sa11_reg[2]/P0001  & ~n14139 ;
  assign n14136 = ~n11836 & ~n11913 ;
  assign n14137 = \sa11_reg[2]/P0001  & ~n14136 ;
  assign n14138 = n11813 & n11858 ;
  assign n14141 = ~n11934 & ~n14138 ;
  assign n14142 = ~n14137 & n14141 ;
  assign n14143 = ~n14140 & n14142 ;
  assign n14144 = ~\sa11_reg[1]/P0001  & ~n14143 ;
  assign n14128 = n11794 & n11816 ;
  assign n14129 = ~n12169 & ~n13139 ;
  assign n14130 = ~n14128 & n14129 ;
  assign n14131 = ~\sa11_reg[2]/P0001  & ~n14130 ;
  assign n14126 = ~n12152 & ~n13522 ;
  assign n14127 = \sa11_reg[2]/P0001  & ~n14126 ;
  assign n14132 = ~n12119 & n12167 ;
  assign n14133 = ~n14127 & n14132 ;
  assign n14134 = ~n14131 & n14133 ;
  assign n14135 = \sa11_reg[1]/P0001  & ~n14134 ;
  assign n14145 = ~n11934 & ~n12176 ;
  assign n14146 = ~\sa11_reg[2]/P0001  & ~n14145 ;
  assign n14147 = ~n13092 & ~n13389 ;
  assign n14148 = n11805 & ~n14147 ;
  assign n14149 = ~n11865 & ~n12205 ;
  assign n14150 = ~n14148 & n14149 ;
  assign n14151 = ~n14146 & n14150 ;
  assign n14152 = ~n14135 & n14151 ;
  assign n14153 = ~n14144 & n14152 ;
  assign n14154 = ~\sa11_reg[0]/P0001  & ~n14153 ;
  assign n14155 = n12126 & n12127 ;
  assign n14156 = ~n12139 & ~n14155 ;
  assign n14157 = ~n11886 & ~n12127 ;
  assign n14158 = ~\sa11_reg[5]/P0001  & ~n14157 ;
  assign n14159 = \sa11_reg[3]/P0001  & n11821 ;
  assign n14160 = ~n14158 & ~n14159 ;
  assign n14161 = \sa11_reg[2]/P0001  & ~n14160 ;
  assign n14162 = n14156 & ~n14161 ;
  assign n14163 = \sa11_reg[1]/P0001  & ~n14162 ;
  assign n14174 = n11794 & ~n11812 ;
  assign n14175 = ~n11821 & n14174 ;
  assign n14176 = ~n11854 & ~n12121 ;
  assign n14177 = ~n14175 & n14176 ;
  assign n14178 = ~\sa11_reg[1]/P0001  & ~n14177 ;
  assign n14165 = ~n11836 & ~n11854 ;
  assign n14164 = \sa11_reg[4]/P0001  & n11847 ;
  assign n14166 = ~n13513 & ~n14164 ;
  assign n14167 = n14165 & n14166 ;
  assign n14168 = ~\sa11_reg[2]/P0001  & ~n14167 ;
  assign n14170 = ~\sa11_reg[1]/P0001  & n13102 ;
  assign n14169 = n11822 & ~n11893 ;
  assign n14171 = ~n14164 & ~n14169 ;
  assign n14172 = ~n14170 & n14171 ;
  assign n14173 = ~\sa11_reg[3]/P0001  & ~n14172 ;
  assign n14179 = ~n14168 & ~n14173 ;
  assign n14180 = ~n14178 & n14179 ;
  assign n14181 = ~n14163 & n14180 ;
  assign n14182 = \sa11_reg[0]/P0001  & ~n14181 ;
  assign n14183 = ~n13109 & ~n13509 ;
  assign n14184 = ~n11879 & n14183 ;
  assign n14185 = ~\sa11_reg[2]/P0001  & ~n14184 ;
  assign n14186 = ~n11927 & ~n12177 ;
  assign n14187 = ~n14185 & n14186 ;
  assign n14188 = ~\sa11_reg[1]/P0001  & ~n14187 ;
  assign n14190 = ~n12128 & ~n12139 ;
  assign n14191 = \sa11_reg[3]/P0001  & ~n14190 ;
  assign n14192 = ~n13132 & ~n14191 ;
  assign n14193 = n13171 & ~n14192 ;
  assign n14189 = \sa11_reg[4]/P0001  & n13450 ;
  assign n14199 = ~n11834 & ~n12222 ;
  assign n14200 = n12119 & n14199 ;
  assign n14204 = ~n14189 & ~n14200 ;
  assign n14205 = ~n14193 & n14204 ;
  assign n14194 = n11797 & n11860 ;
  assign n14195 = ~n12151 & ~n13093 ;
  assign n14196 = ~n14194 & n14195 ;
  assign n14197 = ~n11922 & n14196 ;
  assign n14198 = n13166 & ~n14197 ;
  assign n14201 = ~n11865 & ~n12186 ;
  assign n14202 = ~n13394 & n14201 ;
  assign n14203 = n13544 & ~n14202 ;
  assign n14206 = ~n14198 & ~n14203 ;
  assign n14207 = n14205 & n14206 ;
  assign n14208 = ~n14188 & n14207 ;
  assign n14209 = ~n14182 & n14208 ;
  assign n14210 = ~n14154 & n14209 ;
  assign n14211 = n13649 & ~n14210 ;
  assign n14212 = ~n13649 & n14210 ;
  assign n14213 = ~n14211 & ~n14212 ;
  assign n14214 = ~n14125 & n14213 ;
  assign n14215 = n14125 & ~n14213 ;
  assign n14216 = ~n14214 & ~n14215 ;
  assign n14218 = n14122 & n14216 ;
  assign n14217 = ~n14122 & ~n14216 ;
  assign n14219 = ~\ld_r_reg/P0001  & ~n14217 ;
  assign n14220 = ~n14218 & n14219 ;
  assign n14222 = \text_in_r_reg[105]/P0001  & \u0_w_reg[0][9]/P0001  ;
  assign n14221 = ~\text_in_r_reg[105]/P0001  & ~\u0_w_reg[0][9]/P0001  ;
  assign n14223 = \ld_r_reg/P0001  & ~n14221 ;
  assign n14224 = ~n14222 & n14223 ;
  assign n14225 = ~n14220 & ~n14224 ;
  assign n14226 = \u0_w_reg[0][1]/P0001  & ~n13835 ;
  assign n14227 = ~\u0_w_reg[0][1]/P0001  & n13835 ;
  assign n14228 = ~n14226 & ~n14227 ;
  assign n14229 = n14116 & n14228 ;
  assign n14230 = ~n14116 & ~n14228 ;
  assign n14231 = ~n14229 & ~n14230 ;
  assign n14264 = ~\sa00_reg[4]/P0001  & n11996 ;
  assign n14265 = ~n12066 & ~n14264 ;
  assign n14266 = ~\sa00_reg[3]/P0001  & ~n14265 ;
  assign n14267 = ~n11984 & ~n14266 ;
  assign n14268 = ~\sa00_reg[1]/P0001  & ~n14267 ;
  assign n14278 = \sa00_reg[3]/P0001  & n12095 ;
  assign n14280 = ~n12015 & ~n12636 ;
  assign n14246 = ~\sa00_reg[2]/P0001  & ~\sa00_reg[3]/P0001  ;
  assign n14277 = n12096 & n14246 ;
  assign n14279 = n11982 & n12002 ;
  assign n14281 = ~n14277 & ~n14279 ;
  assign n14282 = n14280 & n14281 ;
  assign n14283 = ~n14278 & n14282 ;
  assign n14284 = \sa00_reg[1]/P0001  & ~n14283 ;
  assign n14240 = n11959 & n13629 ;
  assign n14269 = \sa00_reg[6]/NET0131  & n11974 ;
  assign n14270 = ~n14240 & ~n14269 ;
  assign n14271 = ~n13038 & n14270 ;
  assign n14272 = ~\sa00_reg[2]/P0001  & ~n14271 ;
  assign n14273 = ~n11967 & ~n12035 ;
  assign n14274 = n12596 & ~n14273 ;
  assign n14275 = n11973 & ~n11979 ;
  assign n14276 = n13015 & n14275 ;
  assign n14285 = ~n14274 & ~n14276 ;
  assign n14286 = ~n14272 & n14285 ;
  assign n14287 = ~n14284 & n14286 ;
  assign n14288 = ~n14268 & n14287 ;
  assign n14289 = ~\sa00_reg[0]/P0001  & ~n14288 ;
  assign n14249 = ~\sa00_reg[5]/P0001  & n12015 ;
  assign n14250 = ~n12605 & ~n12692 ;
  assign n14251 = ~n14249 & n14250 ;
  assign n14252 = \sa00_reg[2]/P0001  & ~n14251 ;
  assign n14247 = n11961 & n14246 ;
  assign n14244 = \sa00_reg[5]/P0001  & ~n11952 ;
  assign n14245 = n11966 & ~n14244 ;
  assign n14248 = n12005 & n12026 ;
  assign n14253 = ~n14245 & ~n14248 ;
  assign n14254 = ~n14247 & n14253 ;
  assign n14255 = ~n14252 & n14254 ;
  assign n14256 = ~\sa00_reg[1]/P0001  & ~n14255 ;
  assign n14241 = ~n12091 & ~n14240 ;
  assign n14242 = n13013 & n14241 ;
  assign n14243 = \sa00_reg[2]/P0001  & ~n14242 ;
  assign n14232 = ~\sa00_reg[2]/P0001  & n11957 ;
  assign n14233 = ~n12072 & ~n13068 ;
  assign n14234 = ~n14232 & n14233 ;
  assign n14235 = \sa00_reg[1]/P0001  & ~n14234 ;
  assign n14237 = n11959 & n11995 ;
  assign n14238 = ~n13031 & ~n14237 ;
  assign n14239 = ~\sa00_reg[2]/P0001  & ~n14238 ;
  assign n14236 = ~n12654 & n13044 ;
  assign n14257 = ~n12053 & ~n13575 ;
  assign n14258 = ~n14236 & n14257 ;
  assign n14259 = ~n14239 & n14258 ;
  assign n14260 = ~n14235 & n14259 ;
  assign n14261 = ~n14243 & n14260 ;
  assign n14262 = ~n14256 & n14261 ;
  assign n14263 = \sa00_reg[0]/P0001  & ~n14262 ;
  assign n14301 = ~\sa00_reg[3]/P0001  & n11962 ;
  assign n14302 = ~n12014 & n14301 ;
  assign n14303 = ~n12016 & ~n14302 ;
  assign n14304 = ~\sa00_reg[2]/P0001  & ~n14303 ;
  assign n14305 = \sa00_reg[2]/P0001  & n12005 ;
  assign n14306 = ~n11995 & ~n12685 ;
  assign n14307 = n14305 & ~n14306 ;
  assign n14308 = n13006 & n13044 ;
  assign n14309 = ~n12702 & ~n14308 ;
  assign n14310 = ~n14307 & n14309 ;
  assign n14311 = ~n14304 & n14310 ;
  assign n14312 = ~\sa00_reg[1]/P0001  & ~n14311 ;
  assign n14290 = ~\sa00_reg[4]/P0001  & n12026 ;
  assign n14291 = n12056 & n14290 ;
  assign n14292 = ~n13045 & ~n14291 ;
  assign n14293 = \sa00_reg[6]/NET0131  & ~n14292 ;
  assign n14294 = ~n11993 & ~n12637 ;
  assign n14295 = \sa00_reg[2]/P0001  & ~n14294 ;
  assign n14296 = n12632 & n14246 ;
  assign n14297 = ~n11968 & ~n12006 ;
  assign n14298 = ~n14296 & n14297 ;
  assign n14299 = ~n14295 & n14298 ;
  assign n14300 = \sa00_reg[1]/P0001  & ~n14299 ;
  assign n14313 = ~n14293 & ~n14300 ;
  assign n14314 = ~n14312 & n14313 ;
  assign n14315 = ~n14263 & n14314 ;
  assign n14316 = ~n14289 & n14315 ;
  assign n14354 = ~n12057 & ~n12068 ;
  assign n14355 = ~n13028 & ~n14301 ;
  assign n14356 = n14354 & n14355 ;
  assign n14357 = ~\sa00_reg[2]/P0001  & ~n14356 ;
  assign n14358 = ~n12072 & ~n13036 ;
  assign n14359 = ~\sa00_reg[7]/NET0131  & ~n14358 ;
  assign n14360 = n12056 & n12090 ;
  assign n14361 = ~n12019 & ~n14360 ;
  assign n14362 = ~n14359 & n14361 ;
  assign n14363 = ~n14357 & n14362 ;
  assign n14364 = ~\sa00_reg[1]/P0001  & ~n14363 ;
  assign n14341 = ~n12015 & ~n12065 ;
  assign n14340 = \sa00_reg[3]/P0001  & n11962 ;
  assign n14342 = ~n13028 & ~n14340 ;
  assign n14343 = n14341 & n14342 ;
  assign n14344 = \sa00_reg[1]/P0001  & ~n14343 ;
  assign n14345 = ~n12045 & ~n12614 ;
  assign n14346 = ~n12605 & n14345 ;
  assign n14347 = ~n14344 & n14346 ;
  assign n14348 = \sa00_reg[2]/P0001  & ~n14347 ;
  assign n14350 = n12685 & n14246 ;
  assign n14351 = ~n12051 & ~n14350 ;
  assign n14352 = \sa00_reg[1]/P0001  & ~n14351 ;
  assign n14353 = n12086 & n14301 ;
  assign n14349 = n12054 & n12082 ;
  assign n14365 = ~n13031 & ~n14349 ;
  assign n14366 = ~n14353 & n14365 ;
  assign n14367 = ~n14352 & n14366 ;
  assign n14368 = ~n14348 & n14367 ;
  assign n14369 = ~n14364 & n14368 ;
  assign n14370 = \sa00_reg[0]/P0001  & ~n14369 ;
  assign n14330 = \sa00_reg[2]/P0001  & ~n12036 ;
  assign n14331 = ~n12666 & n13639 ;
  assign n14332 = ~n14330 & ~n14331 ;
  assign n14333 = ~n13037 & ~n13069 ;
  assign n14334 = ~n14332 & n14333 ;
  assign n14335 = \sa00_reg[1]/P0001  & ~n14334 ;
  assign n14326 = ~n13572 & ~n14248 ;
  assign n14327 = ~n12018 & ~n13062 ;
  assign n14328 = n14326 & n14327 ;
  assign n14329 = ~\sa00_reg[2]/P0001  & ~n14328 ;
  assign n14317 = ~n12630 & ~n14237 ;
  assign n14318 = ~n13610 & n14317 ;
  assign n14319 = n12054 & ~n14318 ;
  assign n14320 = ~n11956 & ~n12050 ;
  assign n14321 = n13004 & ~n14320 ;
  assign n14322 = ~\sa00_reg[2]/P0001  & n11978 ;
  assign n14323 = ~n13012 & ~n14322 ;
  assign n14324 = ~n14321 & n14323 ;
  assign n14325 = ~\sa00_reg[1]/P0001  & ~n14324 ;
  assign n14336 = ~n14319 & ~n14325 ;
  assign n14337 = ~n14329 & n14336 ;
  assign n14338 = ~n14335 & n14337 ;
  assign n14339 = ~\sa00_reg[0]/P0001  & ~n14338 ;
  assign n14371 = n11956 & n12014 ;
  assign n14372 = ~n11961 & ~n13074 ;
  assign n14373 = ~n14371 & n14372 ;
  assign n14374 = ~\sa00_reg[3]/P0001  & ~n14373 ;
  assign n14375 = ~n12027 & ~n12624 ;
  assign n14376 = ~n14374 & n14375 ;
  assign n14377 = \sa00_reg[2]/P0001  & ~n14376 ;
  assign n14378 = n11975 & ~n11978 ;
  assign n14379 = n14265 & ~n14378 ;
  assign n14380 = n13044 & ~n14379 ;
  assign n14381 = ~n14377 & ~n14380 ;
  assign n14382 = \sa00_reg[1]/P0001  & ~n14381 ;
  assign n14390 = n11955 & n11973 ;
  assign n14392 = ~n12052 & ~n14390 ;
  assign n14393 = n14326 & n14392 ;
  assign n14391 = \sa00_reg[2]/P0001  & ~n14390 ;
  assign n14394 = ~\sa00_reg[1]/P0001  & ~n14391 ;
  assign n14395 = ~n14393 & n14394 ;
  assign n14383 = n11962 & n12693 ;
  assign n14384 = ~n12081 & ~n14383 ;
  assign n14385 = ~\sa00_reg[2]/P0001  & ~n14384 ;
  assign n14386 = \sa00_reg[5]/P0001  & n13036 ;
  assign n14387 = ~n12051 & ~n12611 ;
  assign n14388 = ~n14386 & n14387 ;
  assign n14389 = n13015 & ~n14388 ;
  assign n14396 = ~n14385 & ~n14389 ;
  assign n14397 = ~n14395 & n14396 ;
  assign n14398 = ~n14382 & n14397 ;
  assign n14399 = ~n14339 & n14398 ;
  assign n14400 = ~n14370 & n14399 ;
  assign n14401 = n14316 & ~n14400 ;
  assign n14402 = ~n14316 & n14400 ;
  assign n14403 = ~n14401 & ~n14402 ;
  assign n14404 = ~n14213 & n14403 ;
  assign n14405 = n14213 & ~n14403 ;
  assign n14406 = ~n14404 & ~n14405 ;
  assign n14408 = n14231 & n14406 ;
  assign n14407 = ~n14231 & ~n14406 ;
  assign n14409 = ~\ld_r_reg/P0001  & ~n14407 ;
  assign n14410 = ~n14408 & n14409 ;
  assign n14412 = \text_in_r_reg[97]/P0001  & \u0_w_reg[0][1]/P0001  ;
  assign n14411 = ~\text_in_r_reg[97]/P0001  & ~\u0_w_reg[0][1]/P0001  ;
  assign n14413 = \ld_r_reg/P0001  & ~n14411 ;
  assign n14414 = ~n14412 & n14413 ;
  assign n14415 = ~n14410 & ~n14414 ;
  assign n14416 = ~n11935 & ~n13509 ;
  assign n14417 = ~\sa11_reg[2]/P0001  & ~n14416 ;
  assign n14418 = ~n11792 & ~n12168 ;
  assign n14419 = \sa11_reg[2]/P0001  & ~n14418 ;
  assign n14420 = ~n11865 & ~n12124 ;
  assign n14421 = ~n11927 & n14420 ;
  assign n14422 = ~n13450 & n14421 ;
  assign n14423 = ~n14419 & n14422 ;
  assign n14424 = ~n14417 & n14423 ;
  assign n14425 = ~\sa11_reg[1]/P0001  & ~n14424 ;
  assign n14426 = \sa11_reg[3]/P0001  & ~\sa11_reg[7]/NET0131  ;
  assign n14427 = n11797 & ~n14426 ;
  assign n14428 = ~n11806 & ~n14427 ;
  assign n14429 = \sa11_reg[2]/P0001  & ~n14428 ;
  assign n14430 = ~n11913 & ~n13473 ;
  assign n14431 = ~n11898 & n14430 ;
  assign n14432 = ~n13390 & ~n13447 ;
  assign n14433 = n14431 & n14432 ;
  assign n14434 = ~n14429 & n14433 ;
  assign n14435 = \sa11_reg[1]/P0001  & ~n14434 ;
  assign n14436 = n11801 & n11860 ;
  assign n14437 = n13421 & ~n14436 ;
  assign n14438 = ~\sa11_reg[2]/P0001  & ~n14437 ;
  assign n14439 = ~n12120 & n12207 ;
  assign n14440 = n11834 & ~n14439 ;
  assign n14441 = ~n12198 & ~n14440 ;
  assign n14442 = ~n14438 & n14441 ;
  assign n14443 = ~n14435 & n14442 ;
  assign n14444 = ~n14425 & n14443 ;
  assign n14445 = \sa11_reg[0]/P0001  & ~n14444 ;
  assign n14466 = ~n12153 & ~n13127 ;
  assign n14467 = \sa11_reg[2]/P0001  & ~n14466 ;
  assign n14468 = \sa11_reg[1]/P0001  & ~n11909 ;
  assign n14469 = ~n11862 & n14468 ;
  assign n14465 = n11797 & n13502 ;
  assign n14470 = ~n14155 & ~n14465 ;
  assign n14471 = n14469 & n14470 ;
  assign n14472 = ~n14467 & n14471 ;
  assign n14475 = n11829 & n11834 ;
  assign n14476 = ~\sa11_reg[1]/P0001  & ~n14436 ;
  assign n14477 = ~n14475 & n14476 ;
  assign n14473 = \sa11_reg[7]/NET0131  & n11805 ;
  assign n14474 = ~n11876 & n14473 ;
  assign n14478 = ~n13172 & ~n14474 ;
  assign n14479 = n14477 & n14478 ;
  assign n14480 = ~n13170 & n14479 ;
  assign n14481 = ~n14472 & ~n14480 ;
  assign n14461 = ~\sa11_reg[2]/P0001  & n13096 ;
  assign n14462 = n11863 & n13092 ;
  assign n14463 = n11908 & ~n14462 ;
  assign n14464 = ~n14461 & ~n14463 ;
  assign n14482 = ~n12195 & ~n14464 ;
  assign n14483 = ~n14481 & n14482 ;
  assign n14484 = ~\sa11_reg[0]/P0001  & ~n14483 ;
  assign n14447 = ~n11882 & ~n13102 ;
  assign n14448 = ~n13489 & n14447 ;
  assign n14449 = n13106 & ~n14448 ;
  assign n14446 = n11893 & n11909 ;
  assign n14450 = ~n11899 & ~n14446 ;
  assign n14451 = ~n14449 & n14450 ;
  assign n14452 = \sa11_reg[1]/P0001  & ~n14451 ;
  assign n14453 = ~n11879 & ~n12195 ;
  assign n14454 = n13544 & ~n14453 ;
  assign n14457 = n11896 & n12222 ;
  assign n14485 = ~n14138 & ~n14457 ;
  assign n14486 = ~n14454 & n14485 ;
  assign n14455 = ~n11883 & ~n12139 ;
  assign n14456 = n11846 & ~n14455 ;
  assign n14458 = \sa11_reg[6]/NET0131  & n11923 ;
  assign n14459 = ~n11913 & ~n14458 ;
  assign n14460 = n13171 & ~n14459 ;
  assign n14487 = ~n14456 & ~n14460 ;
  assign n14488 = n14486 & n14487 ;
  assign n14489 = ~n14452 & n14488 ;
  assign n14490 = ~n14484 & n14489 ;
  assign n14491 = ~n14445 & n14490 ;
  assign n14526 = ~n12330 & ~n12344 ;
  assign n14527 = ~n12753 & n14526 ;
  assign n14528 = \sa22_reg[2]/P0001  & ~n14527 ;
  assign n14530 = ~n12298 & ~n12790 ;
  assign n14531 = n12251 & n13200 ;
  assign n14529 = n12234 & n12779 ;
  assign n14532 = ~n13358 & ~n14529 ;
  assign n14533 = ~n14531 & n14532 ;
  assign n14534 = n14530 & n14533 ;
  assign n14535 = ~n14528 & n14534 ;
  assign n14536 = \sa22_reg[1]/P0001  & ~n14535 ;
  assign n14517 = ~n12321 & ~n12360 ;
  assign n14518 = n12794 & n14517 ;
  assign n14519 = ~\sa22_reg[2]/P0001  & ~n12259 ;
  assign n14520 = ~n12733 & n14519 ;
  assign n14521 = ~n14518 & ~n14520 ;
  assign n14522 = ~n12240 & ~n12371 ;
  assign n14523 = ~n12812 & n14522 ;
  assign n14524 = ~n14521 & n14523 ;
  assign n14525 = ~\sa22_reg[1]/P0001  & ~n14524 ;
  assign n14495 = n12238 & n12291 ;
  assign n14537 = n13351 & ~n14495 ;
  assign n14538 = ~\sa22_reg[2]/P0001  & ~n14537 ;
  assign n14539 = ~n12264 & ~n12374 ;
  assign n14540 = \sa22_reg[2]/P0001  & \sa22_reg[4]/P0001  ;
  assign n14541 = ~n14539 & n14540 ;
  assign n14542 = ~n12343 & ~n14541 ;
  assign n14543 = ~n14538 & n14542 ;
  assign n14544 = ~n14525 & n14543 ;
  assign n14545 = ~n14536 & n14544 ;
  assign n14546 = \sa22_reg[0]/P0001  & ~n14545 ;
  assign n14501 = ~n12393 & ~n12395 ;
  assign n14502 = \sa22_reg[2]/P0001  & ~n14501 ;
  assign n14500 = ~\sa22_reg[2]/P0001  & n12268 ;
  assign n14503 = ~n12281 & ~n12324 ;
  assign n14504 = ~n14500 & n14503 ;
  assign n14505 = ~n13803 & n14504 ;
  assign n14506 = ~n14502 & n14505 ;
  assign n14507 = \sa22_reg[1]/P0001  & ~n14506 ;
  assign n14492 = ~n12234 & n12258 ;
  assign n14493 = ~n13268 & ~n14492 ;
  assign n14494 = \sa22_reg[2]/P0001  & ~n14493 ;
  assign n14496 = ~n13269 & ~n14495 ;
  assign n14497 = ~n13272 & n14496 ;
  assign n14498 = ~n14494 & n14497 ;
  assign n14499 = ~\sa22_reg[1]/P0001  & ~n14498 ;
  assign n14509 = ~\sa22_reg[2]/P0001  & ~n13193 ;
  assign n14510 = n12395 & n12735 ;
  assign n14508 = n12238 & n13197 ;
  assign n14511 = ~n13258 & ~n14508 ;
  assign n14512 = ~n14510 & n14511 ;
  assign n14513 = ~n14509 & n14512 ;
  assign n14514 = ~n14499 & n14513 ;
  assign n14515 = ~n14507 & n14514 ;
  assign n14516 = ~\sa22_reg[0]/P0001  & ~n14515 ;
  assign n14551 = ~n12268 & ~n12772 ;
  assign n14552 = ~n13240 & n14551 ;
  assign n14553 = n13200 & ~n14552 ;
  assign n14547 = n12756 & n13227 ;
  assign n14548 = \sa22_reg[6]/NET0131  & n12355 ;
  assign n14549 = n14530 & ~n14548 ;
  assign n14550 = \sa22_reg[2]/P0001  & ~n14549 ;
  assign n14554 = ~n14547 & ~n14550 ;
  assign n14555 = ~n14553 & n14554 ;
  assign n14556 = \sa22_reg[1]/P0001  & ~n14555 ;
  assign n14557 = ~n12335 & ~n14508 ;
  assign n14558 = n13820 & ~n14557 ;
  assign n14559 = ~n12292 & ~n12773 ;
  assign n14560 = n12735 & ~n14559 ;
  assign n14561 = n12383 & n12782 ;
  assign n14562 = ~n13275 & ~n14561 ;
  assign n14563 = ~n14560 & n14562 ;
  assign n14564 = ~n14558 & n14563 ;
  assign n14565 = ~n14556 & n14564 ;
  assign n14566 = ~n14516 & n14565 ;
  assign n14567 = ~n14546 & n14566 ;
  assign n14568 = n14491 & ~n14567 ;
  assign n14569 = ~n14491 & n14567 ;
  assign n14570 = ~n14568 & ~n14569 ;
  assign n14572 = ~n12564 & ~n13720 ;
  assign n14573 = ~\sa33_reg[2]/P0001  & ~n14572 ;
  assign n14574 = ~n12549 & ~n12946 ;
  assign n14575 = ~n14011 & n14574 ;
  assign n14571 = \sa33_reg[2]/P0001  & n12525 ;
  assign n14576 = ~n12914 & ~n13739 ;
  assign n14577 = ~n14571 & n14576 ;
  assign n14578 = n14575 & n14577 ;
  assign n14579 = ~n14573 & n14578 ;
  assign n14580 = ~\sa33_reg[1]/P0001  & ~n14579 ;
  assign n14582 = \sa33_reg[7]/NET0131  & ~n12446 ;
  assign n14583 = ~n12480 & n14582 ;
  assign n14584 = ~n12430 & ~n14583 ;
  assign n14585 = \sa33_reg[2]/P0001  & ~n14584 ;
  assign n14586 = ~n12433 & ~n12473 ;
  assign n14587 = ~\sa33_reg[2]/P0001  & ~n14586 ;
  assign n14581 = n12418 & n13690 ;
  assign n14588 = ~n12861 & ~n14581 ;
  assign n14589 = ~n14587 & n14588 ;
  assign n14590 = ~n14585 & n14589 ;
  assign n14591 = \sa33_reg[1]/P0001  & ~n14590 ;
  assign n14592 = n12461 & n12479 ;
  assign n14593 = n14074 & ~n14592 ;
  assign n14594 = ~\sa33_reg[2]/P0001  & ~n14593 ;
  assign n14595 = \sa33_reg[2]/P0001  & \sa33_reg[4]/P0001  ;
  assign n14596 = ~n12432 & n12545 ;
  assign n14597 = n14595 & ~n14596 ;
  assign n14598 = ~n12524 & ~n14597 ;
  assign n14599 = ~n14594 & n14598 ;
  assign n14600 = ~n14591 & n14599 ;
  assign n14601 = ~n14580 & n14600 ;
  assign n14602 = \sa33_reg[0]/P0001  & ~n14601 ;
  assign n14603 = ~\sa33_reg[7]/NET0131  & n12446 ;
  assign n14604 = ~n12570 & ~n14603 ;
  assign n14605 = \sa33_reg[2]/P0001  & ~n14604 ;
  assign n14607 = ~\sa33_reg[2]/P0001  & n12411 ;
  assign n14606 = n12481 & ~n12857 ;
  assign n14608 = \sa33_reg[1]/P0001  & ~n12493 ;
  assign n14609 = ~n14606 & n14608 ;
  assign n14610 = ~n14607 & n14609 ;
  assign n14611 = ~n14605 & n14610 ;
  assign n14612 = n12456 & n12468 ;
  assign n14616 = ~\sa33_reg[1]/P0001  & ~n14592 ;
  assign n14617 = ~n14612 & n14616 ;
  assign n14613 = n12472 & n12868 ;
  assign n14614 = ~n12457 & ~n14595 ;
  assign n14615 = n12465 & ~n14614 ;
  assign n14618 = ~n14613 & ~n14615 ;
  assign n14619 = n14617 & n14618 ;
  assign n14620 = ~n14611 & ~n14619 ;
  assign n14621 = ~n12501 & ~n12948 ;
  assign n14622 = ~\sa33_reg[2]/P0001  & ~n14621 ;
  assign n14623 = ~\sa33_reg[7]/NET0131  & n12476 ;
  assign n14624 = n13938 & n14623 ;
  assign n14625 = ~n12518 & ~n12856 ;
  assign n14626 = ~n14624 & n14625 ;
  assign n14627 = ~n14622 & n14626 ;
  assign n14628 = ~n14620 & n14627 ;
  assign n14629 = ~\sa33_reg[0]/P0001  & ~n14628 ;
  assign n14633 = \sa33_reg[6]/P0001  & n12444 ;
  assign n14634 = ~n12411 & ~n13970 ;
  assign n14635 = ~n14633 & n14634 ;
  assign n14636 = n13952 & ~n14635 ;
  assign n14630 = ~n12526 & ~n14005 ;
  assign n14631 = n12945 & ~n14630 ;
  assign n14632 = n12456 & n14044 ;
  assign n14637 = ~n12883 & ~n14632 ;
  assign n14638 = ~n14631 & n14637 ;
  assign n14639 = ~n14636 & n14638 ;
  assign n14640 = \sa33_reg[1]/P0001  & ~n14639 ;
  assign n14641 = ~n12508 & ~n12518 ;
  assign n14642 = n13741 & ~n14641 ;
  assign n14643 = ~n12458 & ~n13948 ;
  assign n14644 = n12877 & ~n14643 ;
  assign n14645 = n12462 & n12560 ;
  assign n14646 = ~n13740 & ~n14645 ;
  assign n14647 = ~n14644 & n14646 ;
  assign n14648 = ~n14642 & n14647 ;
  assign n14649 = ~n14640 & n14648 ;
  assign n14650 = ~n14629 & n14649 ;
  assign n14651 = ~n14602 & n14650 ;
  assign n14652 = \u0_w_reg[0][27]/P0001  & ~n14651 ;
  assign n14653 = ~\u0_w_reg[0][27]/P0001  & n14651 ;
  assign n14654 = ~n14652 & ~n14653 ;
  assign n14655 = n14570 & n14654 ;
  assign n14656 = ~n14570 & ~n14654 ;
  assign n14657 = ~n14655 & ~n14656 ;
  assign n14658 = n13558 & ~n14400 ;
  assign n14659 = ~n13558 & n14400 ;
  assign n14660 = ~n14658 & ~n14659 ;
  assign n14688 = ~n11849 & ~n11887 ;
  assign n14689 = ~n11942 & n14688 ;
  assign n14690 = ~n11793 & ~n11824 ;
  assign n14686 = ~\sa11_reg[5]/P0001  & ~n11893 ;
  assign n14687 = n12146 & ~n14686 ;
  assign n14691 = n11897 & ~n14687 ;
  assign n14692 = n14690 & n14691 ;
  assign n14693 = n14689 & n14692 ;
  assign n14695 = ~n13131 & ~n13489 ;
  assign n14696 = ~\sa11_reg[2]/P0001  & ~n14695 ;
  assign n14694 = n11831 & n13092 ;
  assign n14697 = \sa11_reg[1]/P0001  & ~n14694 ;
  assign n14698 = ~n13440 & n14697 ;
  assign n14699 = ~n14696 & n14698 ;
  assign n14700 = ~n14693 & ~n14699 ;
  assign n14683 = ~n11933 & ~n13159 ;
  assign n14684 = ~n14164 & n14683 ;
  assign n14685 = n11846 & ~n14684 ;
  assign n14701 = ~n11849 & ~n11865 ;
  assign n14702 = \sa11_reg[5]/P0001  & ~n14701 ;
  assign n14703 = \sa11_reg[0]/P0001  & ~n11921 ;
  assign n14704 = ~n14702 & n14703 ;
  assign n14705 = ~n14685 & n14704 ;
  assign n14706 = ~n14700 & n14705 ;
  assign n14708 = ~n11915 & ~n12146 ;
  assign n14709 = \sa11_reg[2]/P0001  & ~n14708 ;
  assign n14710 = ~n13513 & ~n14709 ;
  assign n14711 = \sa11_reg[1]/P0001  & ~n14710 ;
  assign n14717 = ~n13439 & ~n13447 ;
  assign n14718 = ~\sa11_reg[1]/P0001  & ~n14717 ;
  assign n14712 = ~n11858 & ~n13092 ;
  assign n14713 = \sa11_reg[1]/P0001  & ~n11825 ;
  assign n14714 = ~n14712 & n14713 ;
  assign n14715 = ~n11881 & ~n14714 ;
  assign n14716 = ~\sa11_reg[2]/P0001  & ~n14715 ;
  assign n14707 = n11846 & n12223 ;
  assign n14719 = ~\sa11_reg[0]/P0001  & ~n11898 ;
  assign n14720 = ~n14707 & n14719 ;
  assign n14721 = ~n14716 & n14720 ;
  assign n14722 = ~n14718 & n14721 ;
  assign n14723 = ~n14711 & n14722 ;
  assign n14724 = ~n14706 & ~n14723 ;
  assign n14666 = ~n11826 & ~n11922 ;
  assign n14667 = ~n13155 & n14666 ;
  assign n14668 = n13524 & n14667 ;
  assign n14669 = \sa11_reg[3]/P0001  & n11876 ;
  assign n14670 = ~n11934 & ~n14669 ;
  assign n14671 = n13549 & n14670 ;
  assign n14672 = ~n14668 & ~n14671 ;
  assign n14673 = n11876 & ~n11877 ;
  assign n14674 = ~n13092 & n14673 ;
  assign n14675 = ~n14672 & ~n14674 ;
  assign n14676 = ~\sa11_reg[1]/P0001  & ~n14675 ;
  assign n14661 = \sa11_reg[4]/P0001  & n13139 ;
  assign n14662 = n14156 & ~n14661 ;
  assign n14663 = ~\sa11_reg[2]/P0001  & ~n14662 ;
  assign n14664 = ~n11935 & ~n14663 ;
  assign n14665 = \sa11_reg[1]/P0001  & ~n14664 ;
  assign n14677 = n11796 & n12194 ;
  assign n14678 = ~n11861 & ~n12223 ;
  assign n14679 = ~n14677 & n14678 ;
  assign n14680 = n13171 & ~n14679 ;
  assign n14681 = ~n11801 & ~n11847 ;
  assign n14682 = n13457 & ~n14681 ;
  assign n14725 = ~n14446 & ~n14682 ;
  assign n14726 = ~n14680 & n14725 ;
  assign n14727 = ~n14665 & n14726 ;
  assign n14728 = ~n14676 & n14727 ;
  assign n14729 = ~n14724 & n14728 ;
  assign n14771 = ~n12691 & ~n12692 ;
  assign n14772 = ~\sa00_reg[2]/P0001  & ~n14771 ;
  assign n14774 = ~n11954 & ~n12095 ;
  assign n14773 = n11962 & n12056 ;
  assign n14775 = ~n14248 & ~n14773 ;
  assign n14776 = n14774 & n14775 ;
  assign n14777 = n11981 & ~n12023 ;
  assign n14778 = n14776 & n14777 ;
  assign n14779 = ~n14772 & n14778 ;
  assign n14781 = ~n13028 & ~n13036 ;
  assign n14782 = ~\sa00_reg[2]/P0001  & ~n14781 ;
  assign n14780 = \sa00_reg[2]/P0001  & n12636 ;
  assign n14783 = \sa00_reg[1]/P0001  & ~n14308 ;
  assign n14784 = ~n14780 & n14783 ;
  assign n14785 = ~n14782 & n14784 ;
  assign n14786 = ~n14779 & ~n14785 ;
  assign n14788 = ~n11996 & ~n13068 ;
  assign n14789 = ~n13610 & n14788 ;
  assign n14790 = n12054 & ~n14789 ;
  assign n14787 = n12056 & n12651 ;
  assign n14791 = ~n12016 & ~n12022 ;
  assign n14792 = ~n14787 & n14791 ;
  assign n14793 = ~n14790 & n14792 ;
  assign n14794 = ~n14786 & n14793 ;
  assign n14795 = \sa00_reg[0]/P0001  & ~n14794 ;
  assign n14755 = ~n12024 & ~n12034 ;
  assign n14756 = n14391 & n14755 ;
  assign n14757 = ~\sa00_reg[2]/P0001  & ~n14371 ;
  assign n14758 = ~n12018 & n14757 ;
  assign n14759 = ~n13077 & n14758 ;
  assign n14760 = ~n14756 & ~n14759 ;
  assign n14761 = ~n11955 & n11960 ;
  assign n14762 = ~n12007 & n14761 ;
  assign n14763 = ~\sa00_reg[1]/P0001  & ~n13018 ;
  assign n14764 = ~n14762 & n14763 ;
  assign n14765 = ~n14760 & n14764 ;
  assign n14766 = ~n12600 & n13594 ;
  assign n14767 = ~\sa00_reg[2]/P0001  & ~n14766 ;
  assign n14768 = \sa00_reg[1]/P0001  & ~n12033 ;
  assign n14769 = ~n14767 & n14768 ;
  assign n14770 = ~n14765 & ~n14769 ;
  assign n14730 = ~n12008 & ~n12015 ;
  assign n14731 = \sa00_reg[2]/P0001  & ~n14730 ;
  assign n14732 = ~n11979 & ~n12007 ;
  assign n14733 = ~\sa00_reg[2]/P0001  & ~n12026 ;
  assign n14734 = ~n14732 & n14733 ;
  assign n14735 = ~n13069 & ~n14734 ;
  assign n14736 = ~n14731 & n14735 ;
  assign n14737 = \sa00_reg[1]/P0001  & ~n14736 ;
  assign n14739 = n12026 & n13044 ;
  assign n14740 = ~n14390 & ~n14739 ;
  assign n14741 = ~\sa00_reg[1]/P0001  & ~n14740 ;
  assign n14738 = n13004 & n14279 ;
  assign n14742 = ~n11976 & ~n14738 ;
  assign n14743 = ~n13060 & n14742 ;
  assign n14744 = ~n14741 & n14743 ;
  assign n14745 = ~n14737 & n14744 ;
  assign n14746 = ~\sa00_reg[0]/P0001  & ~n14745 ;
  assign n14747 = \sa00_reg[1]/P0001  & n12054 ;
  assign n14748 = n12066 & n14747 ;
  assign n14749 = ~n11967 & ~n12096 ;
  assign n14750 = n14305 & ~n14749 ;
  assign n14796 = ~n14748 & ~n14750 ;
  assign n14751 = n12091 & n13044 ;
  assign n14752 = ~n12005 & ~n13559 ;
  assign n14753 = \sa00_reg[7]/NET0131  & n13571 ;
  assign n14754 = ~n14752 & n14753 ;
  assign n14797 = ~n14751 & ~n14754 ;
  assign n14798 = n14796 & n14797 ;
  assign n14799 = ~n14746 & n14798 ;
  assign n14800 = ~n14770 & n14799 ;
  assign n14801 = ~n14795 & n14800 ;
  assign n14802 = n14729 & ~n14801 ;
  assign n14803 = ~n14729 & n14801 ;
  assign n14804 = ~n14802 & ~n14803 ;
  assign n14805 = ~n14660 & n14804 ;
  assign n14806 = n14660 & ~n14804 ;
  assign n14807 = ~n14805 & ~n14806 ;
  assign n14809 = ~n14657 & n14807 ;
  assign n14808 = n14657 & ~n14807 ;
  assign n14810 = ~\ld_r_reg/P0001  & ~n14808 ;
  assign n14811 = ~n14809 & n14810 ;
  assign n14813 = ~\text_in_r_reg[123]/P0001  & \u0_w_reg[0][27]/P0001  ;
  assign n14812 = \text_in_r_reg[123]/P0001  & ~\u0_w_reg[0][27]/P0001  ;
  assign n14814 = \ld_r_reg/P0001  & ~n14812 ;
  assign n14815 = ~n14813 & n14814 ;
  assign n14816 = ~n14811 & ~n14815 ;
  assign n14817 = n13922 & ~n14567 ;
  assign n14818 = ~n13922 & n14567 ;
  assign n14819 = ~n14817 & ~n14818 ;
  assign n14820 = \u0_w_reg[0][19]/P0001  & ~n14651 ;
  assign n14821 = ~\u0_w_reg[0][19]/P0001  & n14651 ;
  assign n14822 = ~n14820 & ~n14821 ;
  assign n14823 = n14819 & n14822 ;
  assign n14824 = ~n14819 & ~n14822 ;
  assign n14825 = ~n14823 & ~n14824 ;
  assign n14866 = n12301 & n13200 ;
  assign n14870 = ~n12760 & ~n12813 ;
  assign n14871 = ~n14866 & n14870 ;
  assign n14867 = ~n12771 & ~n12782 ;
  assign n14865 = n12251 & n12322 ;
  assign n14868 = ~n13303 & ~n14865 ;
  assign n14869 = n14867 & n14868 ;
  assign n14872 = ~n12346 & n14869 ;
  assign n14873 = n14871 & n14872 ;
  assign n14874 = ~\sa22_reg[1]/P0001  & ~n14873 ;
  assign n14880 = ~n12319 & ~n13251 ;
  assign n14881 = ~n13782 & n14880 ;
  assign n14882 = n12735 & ~n14881 ;
  assign n14875 = ~n12302 & ~n13240 ;
  assign n14876 = n13367 & n14875 ;
  assign n14877 = \sa22_reg[2]/P0001  & ~n12301 ;
  assign n14878 = \sa22_reg[1]/P0001  & ~n14877 ;
  assign n14879 = ~n14876 & n14878 ;
  assign n14883 = ~n12802 & ~n12809 ;
  assign n14884 = ~n13754 & n14883 ;
  assign n14885 = ~n14879 & n14884 ;
  assign n14886 = ~n14882 & n14885 ;
  assign n14887 = ~n14874 & n14886 ;
  assign n14888 = \sa22_reg[0]/P0001  & ~n14887 ;
  assign n14849 = ~n12395 & ~n12805 ;
  assign n14850 = n13319 & n14849 ;
  assign n14851 = \sa22_reg[2]/P0001  & ~n13265 ;
  assign n14852 = ~n12353 & n14851 ;
  assign n14853 = ~n14850 & ~n14852 ;
  assign n14854 = ~n13252 & ~n14853 ;
  assign n14855 = \sa22_reg[1]/P0001  & ~n14854 ;
  assign n14857 = n12349 & n13227 ;
  assign n14858 = ~n13358 & ~n14857 ;
  assign n14859 = ~\sa22_reg[1]/P0001  & ~n14858 ;
  assign n14856 = \sa22_reg[2]/P0001  & n12722 ;
  assign n14860 = ~n12298 & ~n13273 ;
  assign n14861 = ~n14856 & n14860 ;
  assign n14862 = ~n14859 & n14861 ;
  assign n14863 = ~n14855 & n14862 ;
  assign n14864 = ~\sa22_reg[0]/P0001  & ~n14863 ;
  assign n14826 = n12244 & n12266 ;
  assign n14827 = n13804 & ~n14826 ;
  assign n14828 = ~\sa22_reg[2]/P0001  & ~n14827 ;
  assign n14829 = ~n12259 & ~n14828 ;
  assign n14830 = \sa22_reg[1]/P0001  & ~n14829 ;
  assign n14834 = ~n12738 & ~n13257 ;
  assign n14835 = ~n12384 & n14834 ;
  assign n14836 = ~\sa22_reg[2]/P0001  & ~n14835 ;
  assign n14831 = ~n12235 & ~n13358 ;
  assign n14832 = ~n12806 & n14831 ;
  assign n14833 = \sa22_reg[2]/P0001  & ~n14832 ;
  assign n14837 = ~n12756 & ~n13911 ;
  assign n14838 = ~n13201 & n14837 ;
  assign n14839 = ~n14833 & n14838 ;
  assign n14840 = ~n14836 & n14839 ;
  assign n14841 = ~\sa22_reg[1]/P0001  & ~n14840 ;
  assign n14842 = n12303 & n13197 ;
  assign n14843 = ~n12345 & ~n12385 ;
  assign n14844 = ~n14842 & n14843 ;
  assign n14845 = n13264 & ~n14844 ;
  assign n14846 = ~n12291 & ~n12332 ;
  assign n14847 = \sa22_reg[2]/P0001  & n12238 ;
  assign n14848 = ~n14846 & n14847 ;
  assign n14889 = ~n14547 & ~n14848 ;
  assign n14890 = ~n14845 & n14889 ;
  assign n14891 = ~n14841 & n14890 ;
  assign n14892 = ~n14830 & n14891 ;
  assign n14893 = ~n14864 & n14892 ;
  assign n14894 = ~n14888 & n14893 ;
  assign n14895 = n14729 & ~n14894 ;
  assign n14896 = ~n14729 & n14894 ;
  assign n14897 = ~n14895 & ~n14896 ;
  assign n14931 = ~n12655 & ~n14244 ;
  assign n14932 = ~n13629 & ~n14931 ;
  assign n14933 = \sa00_reg[2]/P0001  & ~n14932 ;
  assign n14935 = ~n11976 & ~n12003 ;
  assign n14936 = ~n14390 & n14935 ;
  assign n14934 = ~\sa00_reg[2]/P0001  & n14301 ;
  assign n14937 = ~n14232 & ~n14934 ;
  assign n14938 = n14936 & n14937 ;
  assign n14939 = ~n14933 & n14938 ;
  assign n14940 = \sa00_reg[1]/P0001  & ~n14939 ;
  assign n14923 = ~n11993 & ~n12651 ;
  assign n14924 = ~n14290 & n14923 ;
  assign n14925 = \sa00_reg[2]/P0001  & ~n14924 ;
  assign n14921 = ~n12033 & ~n13580 ;
  assign n14922 = ~\sa00_reg[2]/P0001  & ~n14921 ;
  assign n14926 = ~n12691 & ~n13073 ;
  assign n14927 = ~n12025 & n14926 ;
  assign n14928 = ~n14922 & n14927 ;
  assign n14929 = ~n14925 & n14928 ;
  assign n14930 = ~\sa00_reg[1]/P0001  & ~n14929 ;
  assign n14941 = ~n12021 & n14270 ;
  assign n14942 = ~\sa00_reg[2]/P0001  & ~n14941 ;
  assign n14943 = ~n12613 & n12687 ;
  assign n14944 = \sa00_reg[2]/P0001  & \sa00_reg[4]/P0001  ;
  assign n14945 = ~n14943 & n14944 ;
  assign n14946 = ~n12652 & ~n14945 ;
  assign n14947 = ~n14942 & n14946 ;
  assign n14948 = ~n14930 & n14947 ;
  assign n14949 = ~n14940 & n14948 ;
  assign n14950 = \sa00_reg[0]/P0001  & ~n14949 ;
  assign n14899 = ~n12633 & ~n13032 ;
  assign n14900 = \sa00_reg[2]/P0001  & ~n14899 ;
  assign n14901 = ~n11993 & ~n12046 ;
  assign n14898 = ~\sa00_reg[2]/P0001  & n12612 ;
  assign n14902 = ~n13593 & ~n14898 ;
  assign n14903 = n14901 & n14902 ;
  assign n14904 = ~n14900 & n14903 ;
  assign n14905 = \sa00_reg[1]/P0001  & ~n14904 ;
  assign n14911 = ~n12021 & ~n13085 ;
  assign n14908 = ~n11985 & n12080 ;
  assign n14909 = \sa00_reg[7]/NET0131  & ~n11960 ;
  assign n14910 = n12056 & n14909 ;
  assign n14912 = ~n14908 & ~n14910 ;
  assign n14913 = n14911 & n14912 ;
  assign n14914 = ~\sa00_reg[1]/P0001  & ~n14913 ;
  assign n14907 = ~\sa00_reg[2]/P0001  & ~n12996 ;
  assign n14906 = n12054 & n12633 ;
  assign n14915 = ~n12648 & ~n13075 ;
  assign n14916 = ~n14906 & n14915 ;
  assign n14917 = ~n14907 & n14916 ;
  assign n14918 = ~n14914 & n14917 ;
  assign n14919 = ~n14905 & n14918 ;
  assign n14920 = ~\sa00_reg[0]/P0001  & ~n14919 ;
  assign n14951 = ~n11963 & ~n12612 ;
  assign n14952 = ~n13028 & n14951 ;
  assign n14953 = n14246 & ~n14952 ;
  assign n14954 = ~n11977 & ~n14751 ;
  assign n14955 = ~n14953 & n14954 ;
  assign n14956 = \sa00_reg[1]/P0001  & ~n14955 ;
  assign n14961 = \sa00_reg[6]/NET0131  & n12660 ;
  assign n14962 = ~n12003 & ~n14961 ;
  assign n14963 = n13571 & ~n14962 ;
  assign n14957 = ~n11958 & ~n12648 ;
  assign n14958 = n13015 & ~n14957 ;
  assign n14959 = ~n12094 & ~n12659 ;
  assign n14960 = n11980 & n14959 ;
  assign n14964 = ~n13581 & ~n14960 ;
  assign n14965 = ~n13625 & n14964 ;
  assign n14966 = ~n14958 & n14965 ;
  assign n14967 = ~n14963 & n14966 ;
  assign n14968 = ~n14956 & n14967 ;
  assign n14969 = ~n14920 & n14968 ;
  assign n14970 = ~n14950 & n14969 ;
  assign n14971 = n13558 & ~n14970 ;
  assign n14972 = ~n13558 & n14970 ;
  assign n14973 = ~n14971 & ~n14972 ;
  assign n14974 = n14897 & n14973 ;
  assign n14975 = ~n14897 & ~n14973 ;
  assign n14976 = ~n14974 & ~n14975 ;
  assign n14978 = n14825 & n14976 ;
  assign n14977 = ~n14825 & ~n14976 ;
  assign n14979 = ~\ld_r_reg/P0001  & ~n14977 ;
  assign n14980 = ~n14978 & n14979 ;
  assign n14982 = ~\text_in_r_reg[115]/P0001  & \u0_w_reg[0][19]/P0001  ;
  assign n14981 = \text_in_r_reg[115]/P0001  & ~\u0_w_reg[0][19]/P0001  ;
  assign n14983 = \ld_r_reg/P0001  & ~n14981 ;
  assign n14984 = ~n14982 & n14983 ;
  assign n14985 = ~n14980 & ~n14984 ;
  assign n14986 = n14491 & ~n14970 ;
  assign n14987 = ~n14491 & n14970 ;
  assign n14988 = ~n14986 & ~n14987 ;
  assign n14989 = n13922 & ~n14894 ;
  assign n14990 = ~n13922 & n14894 ;
  assign n14991 = ~n14989 & ~n14990 ;
  assign n14992 = n14988 & n14991 ;
  assign n14993 = ~n14988 & ~n14991 ;
  assign n14994 = ~n14992 & ~n14993 ;
  assign n14995 = n14033 & ~n14651 ;
  assign n14996 = ~n14033 & n14651 ;
  assign n14997 = ~n14995 & ~n14996 ;
  assign n15000 = \sa33_reg[1]/P0001  & ~n14106 ;
  assign n14998 = \sa33_reg[2]/P0001  & n12445 ;
  assign n14999 = n13690 & n14034 ;
  assign n15001 = ~n14998 & ~n14999 ;
  assign n15002 = n15000 & n15001 ;
  assign n15006 = ~n12872 & ~n14052 ;
  assign n15007 = ~n12523 & n15006 ;
  assign n15008 = n12879 & ~n12912 ;
  assign n15003 = \sa33_reg[2]/P0001  & n12414 ;
  assign n15004 = ~n12426 & n15003 ;
  assign n15005 = n12884 & n13986 ;
  assign n15009 = ~n15004 & ~n15005 ;
  assign n15010 = n15008 & n15009 ;
  assign n15011 = n15007 & n15010 ;
  assign n15012 = ~n15002 & ~n15011 ;
  assign n15013 = ~n12481 & ~n13698 ;
  assign n15014 = ~n13667 & n15013 ;
  assign n15015 = n12560 & ~n15014 ;
  assign n15016 = \sa33_reg[0]/P0001  & ~n12909 ;
  assign n15017 = ~n12910 & ~n13702 ;
  assign n15018 = n15016 & n15017 ;
  assign n15019 = ~n15015 & n15018 ;
  assign n15020 = ~n15012 & n15019 ;
  assign n15024 = ~n12864 & ~n13986 ;
  assign n15025 = \sa33_reg[2]/P0001  & ~n15024 ;
  assign n15021 = ~n12444 & ~n12877 ;
  assign n15022 = ~\sa33_reg[2]/P0001  & ~n12510 ;
  assign n15023 = ~n15021 & n15022 ;
  assign n15026 = \sa33_reg[1]/P0001  & ~n13668 ;
  assign n15027 = ~n15023 & n15026 ;
  assign n15028 = ~n15025 & n15027 ;
  assign n15029 = n12456 & n12510 ;
  assign n15030 = ~\sa33_reg[1]/P0001  & ~n12506 ;
  assign n15031 = ~n15029 & n15030 ;
  assign n15032 = ~n15028 & ~n15031 ;
  assign n15034 = n12861 & n14595 ;
  assign n15033 = n12565 & n12881 ;
  assign n15035 = ~\sa33_reg[0]/P0001  & ~n12468 ;
  assign n15036 = ~n15033 & n15035 ;
  assign n15037 = ~n15034 & n15036 ;
  assign n15038 = ~n15032 & n15037 ;
  assign n15039 = ~n15020 & ~n15038 ;
  assign n15043 = n12409 & n12419 ;
  assign n15044 = ~\sa33_reg[2]/P0001  & ~n14023 ;
  assign n15045 = ~n15043 & n15044 ;
  assign n15046 = ~n12550 & ~n12912 ;
  assign n15047 = n15045 & n15046 ;
  assign n15048 = \sa33_reg[2]/P0001  & ~n12427 ;
  assign n15049 = ~n12506 & n15048 ;
  assign n15050 = ~n12919 & n15049 ;
  assign n15051 = ~n15047 & ~n15050 ;
  assign n15052 = ~\sa33_reg[1]/P0001  & ~n14012 ;
  assign n15053 = ~n14044 & n15052 ;
  assign n15054 = ~n15051 & n15053 ;
  assign n15055 = \sa33_reg[5]/P0001  & n14091 ;
  assign n15056 = ~n14624 & ~n15055 ;
  assign n15057 = \sa33_reg[6]/P0001  & ~n15056 ;
  assign n15058 = ~n12522 & ~n12551 ;
  assign n15059 = \sa33_reg[2]/P0001  & ~n15058 ;
  assign n15060 = \sa33_reg[1]/P0001  & ~n12463 ;
  assign n15061 = ~n12564 & ~n14048 ;
  assign n15062 = n15060 & n15061 ;
  assign n15063 = ~n15059 & n15062 ;
  assign n15064 = ~n15057 & n15063 ;
  assign n15065 = ~n15054 & ~n15064 ;
  assign n15040 = ~n12461 & ~n12561 ;
  assign n15041 = \sa33_reg[2]/P0001  & n12479 ;
  assign n15042 = ~n15040 & n15041 ;
  assign n15066 = ~n14632 & ~n15042 ;
  assign n15067 = ~n15065 & n15066 ;
  assign n15068 = ~n15039 & n15067 ;
  assign n15069 = \u0_w_reg[0][11]/P0001  & ~n15068 ;
  assign n15070 = ~\u0_w_reg[0][11]/P0001  & n15068 ;
  assign n15071 = ~n15069 & ~n15070 ;
  assign n15072 = n14997 & n15071 ;
  assign n15073 = ~n14997 & ~n15071 ;
  assign n15074 = ~n15072 & ~n15073 ;
  assign n15076 = n14994 & n15074 ;
  assign n15075 = ~n14994 & ~n15074 ;
  assign n15077 = ~\ld_r_reg/P0001  & ~n15075 ;
  assign n15078 = ~n15076 & n15077 ;
  assign n15080 = ~\text_in_r_reg[107]/P0001  & \u0_w_reg[0][11]/P0001  ;
  assign n15079 = \text_in_r_reg[107]/P0001  & ~\u0_w_reg[0][11]/P0001  ;
  assign n15081 = \ld_r_reg/P0001  & ~n15079 ;
  assign n15082 = ~n15080 & n15081 ;
  assign n15083 = ~n15078 & ~n15082 ;
  assign n15084 = \u0_w_reg[0][12]/P0001  & ~n12962 ;
  assign n15085 = ~\u0_w_reg[0][12]/P0001  & n12962 ;
  assign n15086 = ~n15084 & ~n15085 ;
  assign n15087 = n14997 & n15086 ;
  assign n15088 = ~n14997 & ~n15086 ;
  assign n15089 = ~n15087 & ~n15088 ;
  assign n15090 = n12114 & n14819 ;
  assign n15091 = ~n12114 & ~n14819 ;
  assign n15092 = ~n15090 & ~n15091 ;
  assign n15094 = n15089 & n15092 ;
  assign n15093 = ~n15089 & ~n15092 ;
  assign n15095 = ~\ld_r_reg/P0001  & ~n15093 ;
  assign n15096 = ~n15094 & n15095 ;
  assign n15098 = ~\text_in_r_reg[108]/P0001  & \u0_w_reg[0][12]/P0001  ;
  assign n15097 = \text_in_r_reg[108]/P0001  & ~\u0_w_reg[0][12]/P0001  ;
  assign n15099 = \ld_r_reg/P0001  & ~n15097 ;
  assign n15100 = ~n15098 & n15099 ;
  assign n15101 = ~n15096 & ~n15100 ;
  assign n15102 = \u0_w_reg[0][4]/P0001  & ~n12827 ;
  assign n15103 = ~\u0_w_reg[0][4]/P0001  & n12827 ;
  assign n15104 = ~n15102 & ~n15103 ;
  assign n15105 = n14997 & n15104 ;
  assign n15106 = ~n14997 & ~n15104 ;
  assign n15107 = ~n15105 & ~n15106 ;
  assign n15108 = n14400 & ~n14970 ;
  assign n15109 = ~n14400 & n14970 ;
  assign n15110 = ~n15108 & ~n15109 ;
  assign n15111 = n12114 & n15110 ;
  assign n15112 = ~n12114 & ~n15110 ;
  assign n15113 = ~n15111 & ~n15112 ;
  assign n15115 = n15107 & n15113 ;
  assign n15114 = ~n15107 & ~n15113 ;
  assign n15116 = ~\ld_r_reg/P0001  & ~n15114 ;
  assign n15117 = ~n15115 & n15116 ;
  assign n15119 = ~\text_in_r_reg[100]/P0001  & \u0_w_reg[0][4]/P0001  ;
  assign n15118 = \text_in_r_reg[100]/P0001  & ~\u0_w_reg[0][4]/P0001  ;
  assign n15120 = \ld_r_reg/P0001  & ~n15118 ;
  assign n15121 = ~n15119 & n15120 ;
  assign n15122 = ~n15117 & ~n15121 ;
  assign n15123 = \u0_w_reg[0][25]/P0001  & ~n14210 ;
  assign n15124 = ~\u0_w_reg[0][25]/P0001  & n14210 ;
  assign n15125 = ~n15123 & ~n15124 ;
  assign n15126 = n13838 & n15125 ;
  assign n15127 = ~n13838 & ~n15125 ;
  assign n15128 = ~n15126 & ~n15127 ;
  assign n15129 = n13465 & ~n14316 ;
  assign n15130 = ~n13465 & n14316 ;
  assign n15131 = ~n15129 & ~n15130 ;
  assign n15132 = n14660 & ~n15131 ;
  assign n15133 = ~n14660 & n15131 ;
  assign n15134 = ~n15132 & ~n15133 ;
  assign n15136 = n15128 & n15134 ;
  assign n15135 = ~n15128 & ~n15134 ;
  assign n15137 = ~\ld_r_reg/P0001  & ~n15135 ;
  assign n15138 = ~n15136 & n15137 ;
  assign n15140 = \text_in_r_reg[121]/P0001  & \u0_w_reg[0][25]/P0001  ;
  assign n15139 = ~\text_in_r_reg[121]/P0001  & ~\u0_w_reg[0][25]/P0001  ;
  assign n15141 = \ld_r_reg/P0001  & ~n15139 ;
  assign n15142 = ~n15140 & n15141 ;
  assign n15143 = ~n15138 & ~n15142 ;
  assign n15144 = \u0_w_reg[0][28]/P0001  & ~n12962 ;
  assign n15145 = ~\u0_w_reg[0][28]/P0001  & n12962 ;
  assign n15146 = ~n15144 & ~n15145 ;
  assign n15147 = n12830 & n15146 ;
  assign n15148 = ~n12830 & ~n15146 ;
  assign n15149 = ~n15147 & ~n15148 ;
  assign n15150 = ~n14660 & n14988 ;
  assign n15151 = n14660 & ~n14988 ;
  assign n15152 = ~n15150 & ~n15151 ;
  assign n15154 = ~n15149 & n15152 ;
  assign n15153 = n15149 & ~n15152 ;
  assign n15155 = ~\ld_r_reg/P0001  & ~n15153 ;
  assign n15156 = ~n15154 & n15155 ;
  assign n15158 = ~\text_in_r_reg[124]/P0001  & \u0_w_reg[0][28]/P0001  ;
  assign n15157 = \text_in_r_reg[124]/P0001  & ~\u0_w_reg[0][28]/P0001  ;
  assign n15159 = \ld_r_reg/P0001  & ~n15157 ;
  assign n15160 = ~n15158 & n15159 ;
  assign n15161 = ~n15156 & ~n15160 ;
  assign n15162 = ~\u0_w_reg[0][24]/P0001  & ~n14113 ;
  assign n15163 = \u0_w_reg[0][24]/P0001  & n14113 ;
  assign n15164 = ~n15162 & ~n15163 ;
  assign n15165 = ~n13468 & n14660 ;
  assign n15166 = n13468 & ~n14660 ;
  assign n15167 = ~n15165 & ~n15166 ;
  assign n15169 = n15164 & n15167 ;
  assign n15168 = ~n15164 & ~n15167 ;
  assign n15170 = ~\ld_r_reg/P0001  & ~n15168 ;
  assign n15171 = ~n15169 & n15170 ;
  assign n15173 = \text_in_r_reg[120]/P0001  & \u0_w_reg[0][24]/P0001  ;
  assign n15172 = ~\text_in_r_reg[120]/P0001  & ~\u0_w_reg[0][24]/P0001  ;
  assign n15174 = \ld_r_reg/P0001  & ~n15172 ;
  assign n15175 = ~n15173 & n15174 ;
  assign n15176 = ~n15171 & ~n15175 ;
  assign n15177 = ~\u0_w_reg[0][16]/P0001  & ~n14113 ;
  assign n15178 = \u0_w_reg[0][16]/P0001  & n14113 ;
  assign n15179 = ~n15177 & ~n15178 ;
  assign n15180 = n13558 & ~n14316 ;
  assign n15181 = ~n13558 & n14316 ;
  assign n15182 = ~n15180 & ~n15181 ;
  assign n15183 = n14125 & n15182 ;
  assign n15184 = ~n14125 & ~n15182 ;
  assign n15185 = ~n15183 & ~n15184 ;
  assign n15187 = n15179 & ~n15185 ;
  assign n15186 = ~n15179 & n15185 ;
  assign n15188 = ~\ld_r_reg/P0001  & ~n15186 ;
  assign n15189 = ~n15187 & n15188 ;
  assign n15191 = \text_in_r_reg[112]/P0001  & \u0_w_reg[0][16]/P0001  ;
  assign n15190 = ~\text_in_r_reg[112]/P0001  & ~\u0_w_reg[0][16]/P0001  ;
  assign n15192 = \ld_r_reg/P0001  & ~n15190 ;
  assign n15193 = ~n15191 & n15192 ;
  assign n15194 = ~n15189 & ~n15193 ;
  assign n15195 = n12111 & ~n13558 ;
  assign n15196 = ~n12111 & n13558 ;
  assign n15197 = ~n15195 & ~n15196 ;
  assign n15198 = n14570 & n15197 ;
  assign n15199 = ~n14570 & ~n15197 ;
  assign n15200 = ~n15198 & ~n15199 ;
  assign n15201 = ~n12827 & ~n12962 ;
  assign n15202 = n12827 & n12962 ;
  assign n15203 = ~n15201 & ~n15202 ;
  assign n15204 = \u0_w_reg[0][20]/P0001  & ~n13922 ;
  assign n15205 = ~\u0_w_reg[0][20]/P0001  & n13922 ;
  assign n15206 = ~n15204 & ~n15205 ;
  assign n15207 = n15203 & n15206 ;
  assign n15208 = ~n15203 & ~n15206 ;
  assign n15209 = ~n15207 & ~n15208 ;
  assign n15211 = ~n15200 & n15209 ;
  assign n15210 = n15200 & ~n15209 ;
  assign n15212 = ~\ld_r_reg/P0001  & ~n15210 ;
  assign n15213 = ~n15211 & n15212 ;
  assign n15215 = ~\text_in_r_reg[116]/P0001  & \u0_w_reg[0][20]/P0001  ;
  assign n15214 = \text_in_r_reg[116]/P0001  & ~\u0_w_reg[0][20]/P0001  ;
  assign n15216 = \ld_r_reg/P0001  & ~n15214 ;
  assign n15217 = ~n15215 & n15216 ;
  assign n15218 = ~n15213 & ~n15217 ;
  assign n15219 = ~n12408 & ~n13091 ;
  assign n15220 = n12408 & n13091 ;
  assign n15221 = ~n15219 & ~n15220 ;
  assign n15235 = ~n12411 & ~n12422 ;
  assign n15236 = ~n13699 & n15235 ;
  assign n15237 = \sa33_reg[2]/P0001  & ~n15236 ;
  assign n15234 = n13689 & n13952 ;
  assign n15238 = n14043 & ~n15234 ;
  assign n15239 = ~n15237 & n15238 ;
  assign n15240 = \sa33_reg[1]/P0001  & ~n15239 ;
  assign n15227 = ~n12517 & ~n13939 ;
  assign n15228 = \sa33_reg[2]/P0001  & ~n15227 ;
  assign n15229 = n12430 & n12881 ;
  assign n15230 = ~n12468 & ~n15229 ;
  assign n15231 = n12464 & n15230 ;
  assign n15232 = ~n15228 & n15231 ;
  assign n15233 = ~\sa33_reg[1]/P0001  & ~n15232 ;
  assign n15222 = ~n12415 & ~n12431 ;
  assign n15223 = ~\sa33_reg[2]/P0001  & ~n15222 ;
  assign n15224 = ~n12466 & ~n12493 ;
  assign n15225 = n14621 & n15224 ;
  assign n15226 = \sa33_reg[2]/P0001  & ~n15225 ;
  assign n15241 = ~n15223 & ~n15226 ;
  assign n15242 = ~n15233 & n15241 ;
  assign n15243 = ~n15240 & n15242 ;
  assign n15244 = \sa33_reg[0]/P0001  & ~n15243 ;
  assign n15247 = ~\sa33_reg[1]/P0001  & ~n12415 ;
  assign n15248 = ~n12562 & n15247 ;
  assign n15249 = ~n14091 & n15248 ;
  assign n15245 = ~n12470 & ~n14005 ;
  assign n15246 = ~\sa33_reg[4]/P0001  & ~n15245 ;
  assign n15250 = ~n12929 & ~n15246 ;
  assign n15251 = n15249 & n15250 ;
  assign n15253 = ~n13685 & ~n14603 ;
  assign n15254 = n12472 & ~n15253 ;
  assign n15252 = n12473 & n12884 ;
  assign n15255 = \sa33_reg[1]/P0001  & ~n12550 ;
  assign n15256 = ~n15252 & n15255 ;
  assign n15257 = ~n15254 & n15256 ;
  assign n15258 = ~n15251 & ~n15257 ;
  assign n15259 = n13735 & ~n14073 ;
  assign n15260 = ~n12894 & ~n13970 ;
  assign n15261 = ~n12419 & ~n15260 ;
  assign n15262 = ~n12570 & n12862 ;
  assign n15263 = ~n15261 & n15262 ;
  assign n15264 = ~n15259 & ~n15263 ;
  assign n15265 = ~n15258 & ~n15264 ;
  assign n15266 = ~\sa33_reg[0]/P0001  & ~n15265 ;
  assign n15267 = \sa33_reg[2]/P0001  & ~n12935 ;
  assign n15268 = ~n14016 & n15267 ;
  assign n15269 = ~\sa33_reg[2]/P0001  & ~n12468 ;
  assign n15270 = ~n13698 & n15269 ;
  assign n15271 = ~n13668 & n15270 ;
  assign n15272 = ~n15268 & ~n15271 ;
  assign n15273 = ~n14011 & ~n15043 ;
  assign n15274 = ~n15272 & n15273 ;
  assign n15275 = ~\sa33_reg[1]/P0001  & ~n15274 ;
  assign n15276 = ~n13668 & ~n13986 ;
  assign n15277 = ~\sa33_reg[4]/P0001  & ~n15276 ;
  assign n15278 = ~n13949 & ~n15277 ;
  assign n15279 = n14021 & ~n15278 ;
  assign n15280 = \sa33_reg[1]/P0001  & n15033 ;
  assign n15282 = ~n12474 & ~n12863 ;
  assign n15281 = n13720 & n14595 ;
  assign n15283 = ~n14612 & ~n15281 ;
  assign n15284 = n15282 & n15283 ;
  assign n15285 = ~n15280 & n15284 ;
  assign n15286 = ~n15279 & n15285 ;
  assign n15287 = ~n15275 & n15286 ;
  assign n15288 = ~n15266 & n15287 ;
  assign n15289 = ~n15244 & n15288 ;
  assign n15290 = \u0_w_reg[0][22]/P0001  & ~n15289 ;
  assign n15291 = ~\u0_w_reg[0][22]/P0001  & n15289 ;
  assign n15292 = ~n15290 & ~n15291 ;
  assign n15293 = n13284 & n15292 ;
  assign n15294 = ~n13284 & ~n15292 ;
  assign n15295 = ~n15293 & ~n15294 ;
  assign n15297 = n15221 & n15295 ;
  assign n15296 = ~n15221 & ~n15295 ;
  assign n15298 = ~\ld_r_reg/P0001  & ~n15296 ;
  assign n15299 = ~n15297 & n15298 ;
  assign n15301 = ~\text_in_r_reg[118]/P0001  & \u0_w_reg[0][22]/P0001  ;
  assign n15300 = \text_in_r_reg[118]/P0001  & ~\u0_w_reg[0][22]/P0001  ;
  assign n15302 = \ld_r_reg/P0001  & ~n15300 ;
  assign n15303 = ~n15301 & n15302 ;
  assign n15304 = ~n15299 & ~n15303 ;
  assign n15305 = ~\u0_w_reg[0][8]/P0001  & ~n14113 ;
  assign n15306 = \u0_w_reg[0][8]/P0001  & n14113 ;
  assign n15307 = ~n15305 & ~n15306 ;
  assign n15308 = n13922 & ~n14033 ;
  assign n15309 = ~n13922 & n14033 ;
  assign n15310 = ~n15308 & ~n15309 ;
  assign n15311 = n15131 & ~n15310 ;
  assign n15312 = ~n15131 & n15310 ;
  assign n15313 = ~n15311 & ~n15312 ;
  assign n15315 = n15307 & ~n15313 ;
  assign n15314 = ~n15307 & n15313 ;
  assign n15316 = ~\ld_r_reg/P0001  & ~n15314 ;
  assign n15317 = ~n15315 & n15316 ;
  assign n15319 = ~\text_in_r_reg[104]/P0001  & \u0_w_reg[0][8]/P0001  ;
  assign n15318 = \text_in_r_reg[104]/P0001  & ~\u0_w_reg[0][8]/P0001  ;
  assign n15320 = \ld_r_reg/P0001  & ~n15318 ;
  assign n15321 = ~n15319 & n15320 ;
  assign n15322 = ~n15317 & ~n15321 ;
  assign n15323 = n14491 & ~n14801 ;
  assign n15324 = ~n14491 & n14801 ;
  assign n15325 = ~n15323 & ~n15324 ;
  assign n15326 = n15110 & n15325 ;
  assign n15327 = ~n15110 & ~n15325 ;
  assign n15328 = ~n15326 & ~n15327 ;
  assign n15329 = ~n14033 & ~n14567 ;
  assign n15330 = n14033 & n14567 ;
  assign n15331 = ~n15329 & ~n15330 ;
  assign n15332 = \u0_w_reg[0][3]/P0001  & ~n15068 ;
  assign n15333 = ~\u0_w_reg[0][3]/P0001  & n15068 ;
  assign n15334 = ~n15332 & ~n15333 ;
  assign n15335 = n15331 & n15334 ;
  assign n15336 = ~n15331 & ~n15334 ;
  assign n15337 = ~n15335 & ~n15336 ;
  assign n15339 = ~n15328 & n15337 ;
  assign n15338 = n15328 & ~n15337 ;
  assign n15340 = ~\ld_r_reg/P0001  & ~n15338 ;
  assign n15341 = ~n15339 & n15340 ;
  assign n15343 = ~\text_in_r_reg[99]/P0001  & \u0_w_reg[0][3]/P0001  ;
  assign n15342 = \text_in_r_reg[99]/P0001  & ~\u0_w_reg[0][3]/P0001  ;
  assign n15344 = \ld_r_reg/P0001  & ~n15342 ;
  assign n15345 = ~n15343 & n15344 ;
  assign n15346 = ~n15341 & ~n15345 ;
  assign n15347 = \u0_w_reg[0][26]/P0001  & ~n15068 ;
  assign n15348 = ~\u0_w_reg[0][26]/P0001  & n15068 ;
  assign n15349 = ~n15347 & ~n15348 ;
  assign n15350 = n14897 & n15349 ;
  assign n15351 = ~n14897 & ~n15349 ;
  assign n15352 = ~n15350 & ~n15351 ;
  assign n15354 = n14213 & n15352 ;
  assign n15353 = ~n14213 & ~n15352 ;
  assign n15355 = ~\ld_r_reg/P0001  & ~n15353 ;
  assign n15356 = ~n15354 & n15355 ;
  assign n15358 = \text_in_r_reg[122]/P0001  & \u0_w_reg[0][26]/P0001  ;
  assign n15357 = ~\text_in_r_reg[122]/P0001  & ~\u0_w_reg[0][26]/P0001  ;
  assign n15359 = \ld_r_reg/P0001  & ~n15357 ;
  assign n15360 = ~n15358 & n15359 ;
  assign n15361 = ~n15356 & ~n15360 ;
  assign n15362 = ~n13649 & ~n14804 ;
  assign n15363 = n13649 & n14804 ;
  assign n15364 = ~n15362 & ~n15363 ;
  assign n15365 = \u0_w_reg[0][2]/P0001  & ~n14894 ;
  assign n15366 = ~\u0_w_reg[0][2]/P0001  & n14894 ;
  assign n15367 = ~n15365 & ~n15366 ;
  assign n15368 = n13752 & n15367 ;
  assign n15369 = ~n13752 & ~n15367 ;
  assign n15370 = ~n15368 & ~n15369 ;
  assign n15372 = n15364 & n15370 ;
  assign n15371 = ~n15364 & ~n15370 ;
  assign n15373 = ~\ld_r_reg/P0001  & ~n15371 ;
  assign n15374 = ~n15372 & n15373 ;
  assign n15376 = ~\text_in_r_reg[98]/P0001  & \u0_w_reg[0][2]/P0001  ;
  assign n15375 = \text_in_r_reg[98]/P0001  & ~\u0_w_reg[0][2]/P0001  ;
  assign n15377 = \ld_r_reg/P0001  & ~n15375 ;
  assign n15378 = ~n15376 & n15377 ;
  assign n15379 = ~n15374 & ~n15378 ;
  assign n15380 = n13183 & ~n13284 ;
  assign n15381 = ~n13183 & n13284 ;
  assign n15382 = ~n15380 & ~n15381 ;
  assign n15383 = \u0_w_reg[0][30]/P0001  & ~n15289 ;
  assign n15384 = ~\u0_w_reg[0][30]/P0001  & n15289 ;
  assign n15385 = ~n15383 & ~n15384 ;
  assign n15386 = n15382 & n15385 ;
  assign n15387 = ~n15382 & ~n15385 ;
  assign n15388 = ~n15386 & ~n15387 ;
  assign n15390 = n12851 & n15388 ;
  assign n15389 = ~n12851 & ~n15388 ;
  assign n15391 = ~\ld_r_reg/P0001  & ~n15389 ;
  assign n15392 = ~n15390 & n15391 ;
  assign n15394 = \text_in_r_reg[126]/P0001  & \u0_w_reg[0][30]/P0001  ;
  assign n15393 = ~\text_in_r_reg[126]/P0001  & ~\u0_w_reg[0][30]/P0001  ;
  assign n15395 = \ld_r_reg/P0001  & ~n15393 ;
  assign n15396 = ~n15394 & n15395 ;
  assign n15397 = ~n15392 & ~n15396 ;
  assign n15398 = \u0_w_reg[0][31]/P0001  & ~n13558 ;
  assign n15399 = ~\u0_w_reg[0][31]/P0001  & n13558 ;
  assign n15400 = ~n15398 & ~n15399 ;
  assign n15401 = n13186 & n15310 ;
  assign n15402 = ~n13186 & ~n15310 ;
  assign n15403 = ~n15401 & ~n15402 ;
  assign n15405 = n15400 & ~n15403 ;
  assign n15404 = ~n15400 & n15403 ;
  assign n15406 = ~\ld_r_reg/P0001  & ~n15404 ;
  assign n15407 = ~n15405 & n15406 ;
  assign n15409 = ~\text_in_r_reg[127]/P0001  & \u0_w_reg[0][31]/P0001  ;
  assign n15408 = \text_in_r_reg[127]/P0001  & ~\u0_w_reg[0][31]/P0001  ;
  assign n15410 = \ld_r_reg/P0001  & ~n15408 ;
  assign n15411 = ~n15409 & n15410 ;
  assign n15412 = ~n15407 & ~n15411 ;
  assign n15413 = ~n13835 & ~n14801 ;
  assign n15414 = n13835 & n14801 ;
  assign n15415 = ~n15413 & ~n15414 ;
  assign n15416 = ~n14210 & ~n15415 ;
  assign n15417 = n14210 & n15415 ;
  assign n15418 = ~n15416 & ~n15417 ;
  assign n15419 = \u0_w_reg[0][18]/P0001  & ~n15068 ;
  assign n15420 = ~\u0_w_reg[0][18]/P0001  & n15068 ;
  assign n15421 = ~n15419 & ~n15420 ;
  assign n15422 = n14894 & n15421 ;
  assign n15423 = ~n14894 & ~n15421 ;
  assign n15424 = ~n15422 & ~n15423 ;
  assign n15426 = n15418 & ~n15424 ;
  assign n15425 = ~n15418 & n15424 ;
  assign n15427 = ~\ld_r_reg/P0001  & ~n15425 ;
  assign n15428 = ~n15426 & n15427 ;
  assign n15430 = ~\text_in_r_reg[114]/P0001  & \u0_w_reg[0][18]/P0001  ;
  assign n15429 = \text_in_r_reg[114]/P0001  & ~\u0_w_reg[0][18]/P0001  ;
  assign n15431 = \ld_r_reg/P0001  & ~n15429 ;
  assign n15432 = ~n15430 & n15431 ;
  assign n15433 = ~n15428 & ~n15432 ;
  assign n15434 = ~n14400 & ~n15382 ;
  assign n15435 = n14400 & n15382 ;
  assign n15436 = ~n15434 & ~n15435 ;
  assign n15437 = ~\u0_w_reg[0][23]/P0001  & ~n15310 ;
  assign n15438 = \u0_w_reg[0][23]/P0001  & n15310 ;
  assign n15439 = ~n15437 & ~n15438 ;
  assign n15441 = n15436 & n15439 ;
  assign n15440 = ~n15436 & ~n15439 ;
  assign n15442 = ~\ld_r_reg/P0001  & ~n15440 ;
  assign n15443 = ~n15441 & n15442 ;
  assign n15445 = ~\text_in_r_reg[119]/P0001  & \u0_w_reg[0][23]/P0001  ;
  assign n15444 = \text_in_r_reg[119]/P0001  & ~\u0_w_reg[0][23]/P0001  ;
  assign n15446 = \ld_r_reg/P0001  & ~n15444 ;
  assign n15447 = ~n15445 & n15446 ;
  assign n15448 = ~n15443 & ~n15447 ;
  assign n15449 = ~n12405 & ~n13186 ;
  assign n15450 = n12405 & n13186 ;
  assign n15451 = ~n15449 & ~n15450 ;
  assign n15452 = \u0_w_reg[0][14]/P0001  & ~n15289 ;
  assign n15453 = ~\u0_w_reg[0][14]/P0001  & n15289 ;
  assign n15454 = ~n15452 & ~n15453 ;
  assign n15455 = n12580 & n15454 ;
  assign n15456 = ~n12580 & ~n15454 ;
  assign n15457 = ~n15455 & ~n15456 ;
  assign n15459 = n15451 & n15457 ;
  assign n15458 = ~n15451 & ~n15457 ;
  assign n15460 = ~\ld_r_reg/P0001  & ~n15458 ;
  assign n15461 = ~n15459 & n15460 ;
  assign n15463 = ~\text_in_r_reg[110]/P0001  & \u0_w_reg[0][14]/P0001  ;
  assign n15462 = \text_in_r_reg[110]/P0001  & ~\u0_w_reg[0][14]/P0001  ;
  assign n15464 = \ld_r_reg/P0001  & ~n15462 ;
  assign n15465 = ~n15463 & n15464 ;
  assign n15466 = ~n15461 & ~n15465 ;
  assign n15467 = ~n13284 & ~n14660 ;
  assign n15468 = n13284 & n14660 ;
  assign n15469 = ~n15467 & ~n15468 ;
  assign n15470 = \u0_w_reg[0][15]/P0001  & ~n14033 ;
  assign n15471 = ~\u0_w_reg[0][15]/P0001  & n14033 ;
  assign n15472 = ~n15470 & ~n15471 ;
  assign n15473 = n15289 & n15472 ;
  assign n15474 = ~n15289 & ~n15472 ;
  assign n15475 = ~n15473 & ~n15474 ;
  assign n15477 = n15469 & n15475 ;
  assign n15476 = ~n15469 & ~n15475 ;
  assign n15478 = ~\ld_r_reg/P0001  & ~n15476 ;
  assign n15479 = ~n15477 & n15478 ;
  assign n15481 = ~\text_in_r_reg[111]/P0001  & \u0_w_reg[0][15]/P0001  ;
  assign n15480 = \text_in_r_reg[111]/P0001  & ~\u0_w_reg[0][15]/P0001  ;
  assign n15482 = \ld_r_reg/P0001  & ~n15480 ;
  assign n15483 = ~n15481 & n15482 ;
  assign n15484 = ~n15479 & ~n15483 ;
  assign n15485 = ~n13091 & ~n14660 ;
  assign n15486 = n13091 & n14660 ;
  assign n15487 = ~n15485 & ~n15486 ;
  assign n15488 = \u0_w_reg[0][7]/P0001  & ~n15289 ;
  assign n15489 = ~\u0_w_reg[0][7]/P0001  & n15289 ;
  assign n15490 = ~n15488 & ~n15489 ;
  assign n15491 = n13922 & n15490 ;
  assign n15492 = ~n13922 & ~n15490 ;
  assign n15493 = ~n15491 & ~n15492 ;
  assign n15495 = n15487 & n15493 ;
  assign n15494 = ~n15487 & ~n15493 ;
  assign n15496 = ~\ld_r_reg/P0001  & ~n15494 ;
  assign n15497 = ~n15495 & n15496 ;
  assign n15499 = ~\text_in_r_reg[103]/P0001  & \u0_w_reg[0][7]/P0001  ;
  assign n15498 = \text_in_r_reg[103]/P0001  & ~\u0_w_reg[0][7]/P0001  ;
  assign n15500 = \ld_r_reg/P0001  & ~n15498 ;
  assign n15501 = ~n15499 & n15500 ;
  assign n15502 = ~n15497 & ~n15501 ;
  assign n15525 = ~\u0_w_reg[3][19]/P0001  & \u0_w_reg[3][20]/P0001  ;
  assign n15559 = \u0_w_reg[3][21]/P0001  & ~\u0_w_reg[3][22]/P0001  ;
  assign n15576 = n15525 & n15559 ;
  assign n15503 = \u0_w_reg[3][22]/P0001  & ~\u0_w_reg[3][23]/P0001  ;
  assign n15506 = ~\u0_w_reg[3][19]/P0001  & ~\u0_w_reg[3][20]/P0001  ;
  assign n15574 = n15503 & n15506 ;
  assign n15530 = ~\u0_w_reg[3][22]/P0001  & \u0_w_reg[3][23]/P0001  ;
  assign n15575 = \u0_w_reg[3][19]/P0001  & n15530 ;
  assign n15577 = ~n15574 & ~n15575 ;
  assign n15578 = ~n15576 & n15577 ;
  assign n15579 = ~\u0_w_reg[3][18]/P0001  & ~n15578 ;
  assign n15512 = \u0_w_reg[3][21]/P0001  & \u0_w_reg[3][22]/P0001  ;
  assign n15580 = n15506 & n15512 ;
  assign n15581 = ~\u0_w_reg[3][23]/P0001  & n15580 ;
  assign n15537 = \u0_w_reg[3][19]/P0001  & ~\u0_w_reg[3][23]/P0001  ;
  assign n15549 = ~\u0_w_reg[3][21]/P0001  & ~\u0_w_reg[3][22]/P0001  ;
  assign n15584 = n15537 & n15549 ;
  assign n15593 = ~n15581 & ~n15584 ;
  assign n15526 = \u0_w_reg[3][21]/P0001  & \u0_w_reg[3][23]/P0001  ;
  assign n15582 = ~\u0_w_reg[3][20]/P0001  & n15526 ;
  assign n15583 = ~\u0_w_reg[3][22]/P0001  & n15582 ;
  assign n15551 = \u0_w_reg[3][20]/P0001  & ~\u0_w_reg[3][23]/P0001  ;
  assign n15585 = n15512 & n15551 ;
  assign n15586 = \u0_w_reg[3][18]/P0001  & n15585 ;
  assign n15594 = ~n15583 & ~n15586 ;
  assign n15587 = \u0_w_reg[3][19]/P0001  & n15526 ;
  assign n15588 = ~\u0_w_reg[3][18]/P0001  & ~\u0_w_reg[3][20]/P0001  ;
  assign n15589 = n15587 & ~n15588 ;
  assign n15590 = \u0_w_reg[3][22]/P0001  & \u0_w_reg[3][23]/P0001  ;
  assign n15591 = ~\u0_w_reg[3][21]/P0001  & n15590 ;
  assign n15592 = ~\u0_w_reg[3][19]/P0001  & n15591 ;
  assign n15595 = ~n15589 & ~n15592 ;
  assign n15596 = n15594 & n15595 ;
  assign n15597 = n15593 & n15596 ;
  assign n15598 = ~n15579 & n15597 ;
  assign n15599 = \u0_w_reg[3][17]/P0001  & ~n15598 ;
  assign n15520 = ~\u0_w_reg[3][22]/P0001  & ~\u0_w_reg[3][23]/P0001  ;
  assign n15557 = ~\u0_w_reg[3][21]/P0001  & n15520 ;
  assign n15600 = \u0_w_reg[3][18]/P0001  & n15557 ;
  assign n15601 = ~\u0_w_reg[3][21]/P0001  & \u0_w_reg[3][23]/P0001  ;
  assign n15602 = \u0_w_reg[3][20]/P0001  & n15601 ;
  assign n15603 = ~\u0_w_reg[3][22]/P0001  & n15602 ;
  assign n15604 = ~n15600 & ~n15603 ;
  assign n15605 = ~\u0_w_reg[3][19]/P0001  & ~n15604 ;
  assign n15606 = \u0_w_reg[3][21]/P0001  & n15590 ;
  assign n15607 = n15506 & n15606 ;
  assign n15550 = ~\u0_w_reg[3][20]/P0001  & n15549 ;
  assign n15608 = \u0_w_reg[3][18]/P0001  & \u0_w_reg[3][19]/P0001  ;
  assign n15609 = n15550 & n15608 ;
  assign n15610 = ~n15607 & ~n15609 ;
  assign n15611 = ~n15605 & n15610 ;
  assign n15612 = ~\u0_w_reg[3][17]/P0001  & ~n15611 ;
  assign n15613 = ~\u0_w_reg[3][20]/P0001  & ~\u0_w_reg[3][23]/P0001  ;
  assign n15614 = ~\u0_w_reg[3][21]/P0001  & n15613 ;
  assign n15615 = \u0_w_reg[3][20]/P0001  & n15526 ;
  assign n15616 = ~n15614 & ~n15615 ;
  assign n15617 = \u0_w_reg[3][19]/P0001  & ~n15616 ;
  assign n15518 = ~\u0_w_reg[3][21]/P0001  & \u0_w_reg[3][22]/P0001  ;
  assign n15618 = n15518 & n15551 ;
  assign n15619 = ~\u0_w_reg[3][19]/P0001  & n15618 ;
  assign n15620 = ~\u0_w_reg[3][20]/P0001  & n15520 ;
  assign n15621 = ~n15619 & ~n15620 ;
  assign n15622 = ~n15617 & n15621 ;
  assign n15623 = \u0_w_reg[3][18]/P0001  & ~n15622 ;
  assign n15552 = ~\u0_w_reg[3][21]/P0001  & n15551 ;
  assign n15624 = \u0_w_reg[3][19]/P0001  & n15552 ;
  assign n15539 = ~\u0_w_reg[3][20]/P0001  & \u0_w_reg[3][22]/P0001  ;
  assign n15625 = n15539 & n15601 ;
  assign n15626 = ~n15624 & ~n15625 ;
  assign n15627 = ~\u0_w_reg[3][18]/P0001  & ~n15626 ;
  assign n15544 = \u0_w_reg[3][20]/P0001  & \u0_w_reg[3][23]/P0001  ;
  assign n15628 = n15544 & n15559 ;
  assign n15629 = ~\u0_w_reg[3][18]/P0001  & n15628 ;
  assign n15630 = n15549 & n15613 ;
  assign n15631 = ~n15629 & ~n15630 ;
  assign n15632 = ~n15627 & n15631 ;
  assign n15633 = ~n15623 & n15632 ;
  assign n15634 = ~n15612 & n15633 ;
  assign n15635 = ~n15599 & n15634 ;
  assign n15636 = ~\u0_w_reg[3][16]/P0001  & ~n15635 ;
  assign n15504 = \u0_w_reg[3][19]/P0001  & ~\u0_w_reg[3][20]/P0001  ;
  assign n15505 = \u0_w_reg[3][21]/P0001  & n15504 ;
  assign n15553 = ~n15505 & ~n15550 ;
  assign n15554 = ~n15552 & n15553 ;
  assign n15555 = ~\u0_w_reg[3][18]/P0001  & ~n15554 ;
  assign n15556 = n15504 & n15530 ;
  assign n15558 = n15525 & n15557 ;
  assign n15564 = ~n15556 & ~n15558 ;
  assign n15560 = ~\u0_w_reg[3][19]/P0001  & n15559 ;
  assign n15561 = n15544 & n15560 ;
  assign n15542 = \u0_w_reg[3][21]/P0001  & ~\u0_w_reg[3][23]/P0001  ;
  assign n15521 = \u0_w_reg[3][19]/P0001  & \u0_w_reg[3][20]/P0001  ;
  assign n15562 = ~\u0_w_reg[3][22]/P0001  & n15521 ;
  assign n15563 = n15542 & n15562 ;
  assign n15565 = ~n15561 & ~n15563 ;
  assign n15566 = n15564 & n15565 ;
  assign n15567 = ~n15555 & n15566 ;
  assign n15568 = \u0_w_reg[3][17]/P0001  & ~n15567 ;
  assign n15519 = ~\u0_w_reg[3][20]/P0001  & n15518 ;
  assign n15522 = n15520 & n15521 ;
  assign n15523 = ~n15519 & ~n15522 ;
  assign n15524 = \u0_w_reg[3][18]/P0001  & ~n15523 ;
  assign n15529 = ~\u0_w_reg[3][18]/P0001  & \u0_w_reg[3][19]/P0001  ;
  assign n15531 = ~\u0_w_reg[3][21]/P0001  & n15530 ;
  assign n15532 = n15529 & n15531 ;
  assign n15511 = \u0_w_reg[3][18]/P0001  & ~\u0_w_reg[3][19]/P0001  ;
  assign n15516 = \u0_w_reg[3][21]/P0001  & n15503 ;
  assign n15517 = ~n15511 & n15516 ;
  assign n15527 = n15525 & n15526 ;
  assign n15528 = \u0_w_reg[3][22]/P0001  & n15527 ;
  assign n15533 = ~n15517 & ~n15528 ;
  assign n15534 = ~n15532 & n15533 ;
  assign n15535 = ~n15524 & n15534 ;
  assign n15536 = ~\u0_w_reg[3][17]/P0001  & ~n15535 ;
  assign n15538 = n15512 & n15537 ;
  assign n15540 = n15537 & n15539 ;
  assign n15541 = ~n15538 & ~n15540 ;
  assign n15543 = ~\u0_w_reg[3][20]/P0001  & n15542 ;
  assign n15545 = n15518 & n15544 ;
  assign n15546 = ~n15543 & ~n15545 ;
  assign n15547 = n15541 & n15546 ;
  assign n15548 = ~\u0_w_reg[3][18]/P0001  & ~n15547 ;
  assign n15507 = \u0_w_reg[3][18]/P0001  & n15506 ;
  assign n15508 = ~\u0_w_reg[3][21]/P0001  & n15507 ;
  assign n15509 = ~n15505 & ~n15508 ;
  assign n15510 = n15503 & ~n15509 ;
  assign n15513 = \u0_w_reg[3][20]/P0001  & n15512 ;
  assign n15514 = \u0_w_reg[3][23]/P0001  & n15513 ;
  assign n15515 = n15511 & n15514 ;
  assign n15569 = ~n15510 & ~n15515 ;
  assign n15570 = ~n15548 & n15569 ;
  assign n15571 = ~n15536 & n15570 ;
  assign n15572 = ~n15568 & n15571 ;
  assign n15573 = \u0_w_reg[3][16]/P0001  & ~n15572 ;
  assign n15637 = n15506 & n15520 ;
  assign n15638 = ~\u0_w_reg[3][21]/P0001  & n15503 ;
  assign n15639 = ~n15531 & ~n15638 ;
  assign n15640 = n15525 & ~n15639 ;
  assign n15641 = n15521 & n15559 ;
  assign n15642 = ~n15528 & ~n15641 ;
  assign n15643 = ~n15640 & n15642 ;
  assign n15644 = \u0_w_reg[3][18]/P0001  & ~n15643 ;
  assign n15645 = ~n15637 & ~n15644 ;
  assign n15646 = ~\u0_w_reg[3][17]/P0001  & ~n15645 ;
  assign n15664 = n15511 & n15585 ;
  assign n15662 = ~\u0_w_reg[3][21]/P0001  & n15504 ;
  assign n15663 = n15520 & n15662 ;
  assign n15665 = ~n15629 & ~n15663 ;
  assign n15666 = ~n15664 & n15665 ;
  assign n15667 = \u0_w_reg[3][17]/P0001  & ~n15666 ;
  assign n15650 = n15513 & n15537 ;
  assign n15651 = ~\u0_w_reg[3][18]/P0001  & n15650 ;
  assign n15647 = ~\u0_w_reg[3][18]/P0001  & n15545 ;
  assign n15648 = ~\u0_w_reg[3][18]/P0001  & ~\u0_w_reg[3][19]/P0001  ;
  assign n15649 = n15582 & n15648 ;
  assign n15652 = ~n15647 & ~n15649 ;
  assign n15653 = ~n15651 & n15652 ;
  assign n15654 = ~\u0_w_reg[3][17]/P0001  & ~n15653 ;
  assign n15657 = n15504 & n15559 ;
  assign n15658 = ~\u0_w_reg[3][23]/P0001  & n15657 ;
  assign n15659 = ~\u0_w_reg[3][18]/P0001  & n15658 ;
  assign n15655 = n15551 & n15559 ;
  assign n15656 = n15608 & n15655 ;
  assign n15660 = ~\u0_w_reg[3][21]/P0001  & n15648 ;
  assign n15661 = n15590 & n15660 ;
  assign n15668 = ~n15656 & ~n15661 ;
  assign n15669 = ~n15659 & n15668 ;
  assign n15670 = ~n15654 & n15669 ;
  assign n15671 = ~n15667 & n15670 ;
  assign n15672 = ~n15646 & n15671 ;
  assign n15673 = ~n15573 & n15672 ;
  assign n15674 = ~n15636 & n15673 ;
  assign n15675 = \u0_r0_out_reg[29]/P0001  & ~n15674 ;
  assign n15676 = ~\u0_r0_out_reg[29]/P0001  & n15674 ;
  assign n15677 = ~n15675 & ~n15676 ;
  assign n15679 = \u0_w_reg[0][29]/P0001  & n15677 ;
  assign n15678 = ~\u0_w_reg[0][29]/P0001  & ~n15677 ;
  assign n15680 = ~ld_pad & ~n15678 ;
  assign n15681 = ~n15679 & n15680 ;
  assign n15682 = \key[125]_pad  & ld_pad ;
  assign n15683 = ~n15681 & ~n15682 ;
  assign n15684 = ~\key[61]_pad  & ld_pad ;
  assign n15685 = \u0_w_reg[0][29]/P0001  & ~\u0_w_reg[1][29]/P0002  ;
  assign n15686 = ~\u0_w_reg[0][29]/P0001  & \u0_w_reg[1][29]/P0002  ;
  assign n15687 = ~n15685 & ~n15686 ;
  assign n15688 = \u0_w_reg[2][29]/P0001  & n15687 ;
  assign n15689 = ~\u0_w_reg[2][29]/P0001  & ~n15687 ;
  assign n15690 = ~n15688 & ~n15689 ;
  assign n15691 = n15677 & n15690 ;
  assign n15692 = ~n15677 & ~n15690 ;
  assign n15693 = ~n15691 & ~n15692 ;
  assign n15694 = ~ld_pad & n15693 ;
  assign n15695 = ~n15684 & ~n15694 ;
  assign n15697 = \u0_w_reg[3][29]/P0001  & ~n15693 ;
  assign n15696 = ~\u0_w_reg[3][29]/P0001  & n15693 ;
  assign n15698 = ~ld_pad & ~n15696 ;
  assign n15699 = ~n15697 & n15698 ;
  assign n15700 = \key[29]_pad  & ld_pad ;
  assign n15701 = ~n15699 & ~n15700 ;
  assign n15702 = ~\key[53]_pad  & ld_pad ;
  assign n15725 = \u0_w_reg[3][14]/P0001  & ~\u0_w_reg[3][15]/P0001  ;
  assign n15741 = \u0_w_reg[3][13]/P0001  & n15725 ;
  assign n15742 = ~\u0_w_reg[3][14]/P0001  & \u0_w_reg[3][15]/P0001  ;
  assign n15743 = \u0_w_reg[3][11]/P0001  & n15742 ;
  assign n15744 = ~\u0_w_reg[3][13]/P0001  & n15743 ;
  assign n15745 = ~n15741 & ~n15744 ;
  assign n15746 = ~\u0_w_reg[3][10]/P0001  & ~n15745 ;
  assign n15735 = \u0_w_reg[3][11]/P0001  & \u0_w_reg[3][12]/P0001  ;
  assign n15736 = ~\u0_w_reg[3][14]/P0001  & ~\u0_w_reg[3][15]/P0001  ;
  assign n15737 = n15735 & n15736 ;
  assign n15708 = ~\u0_w_reg[3][13]/P0001  & \u0_w_reg[3][14]/P0001  ;
  assign n15738 = ~\u0_w_reg[3][12]/P0001  & n15708 ;
  assign n15739 = ~n15737 & ~n15738 ;
  assign n15740 = \u0_w_reg[3][10]/P0001  & ~n15739 ;
  assign n15703 = \u0_w_reg[3][12]/P0001  & \u0_w_reg[3][15]/P0001  ;
  assign n15704 = \u0_w_reg[3][14]/P0001  & n15703 ;
  assign n15705 = \u0_w_reg[3][13]/P0001  & n15704 ;
  assign n15706 = ~\u0_w_reg[3][11]/P0001  & n15705 ;
  assign n15713 = \u0_w_reg[3][13]/P0001  & \u0_w_reg[3][14]/P0001  ;
  assign n15714 = \u0_w_reg[3][11]/P0001  & ~\u0_w_reg[3][15]/P0001  ;
  assign n15715 = n15713 & n15714 ;
  assign n15747 = ~\u0_w_reg[3][9]/P0001  & ~n15715 ;
  assign n15748 = ~n15706 & n15747 ;
  assign n15749 = ~n15740 & n15748 ;
  assign n15750 = ~n15746 & n15749 ;
  assign n15756 = ~\u0_w_reg[3][13]/P0001  & ~\u0_w_reg[3][14]/P0001  ;
  assign n15757 = \u0_w_reg[3][12]/P0001  & ~\u0_w_reg[3][15]/P0001  ;
  assign n15758 = n15756 & n15757 ;
  assign n15759 = ~\u0_w_reg[3][11]/P0001  & n15758 ;
  assign n15760 = \u0_w_reg[3][9]/P0001  & ~n15759 ;
  assign n15761 = ~\u0_w_reg[3][12]/P0001  & n15743 ;
  assign n15751 = ~\u0_w_reg[3][11]/P0001  & \u0_w_reg[3][12]/P0001  ;
  assign n15752 = n15742 & n15751 ;
  assign n15753 = \u0_w_reg[3][13]/P0001  & n15752 ;
  assign n15719 = \u0_w_reg[3][13]/P0001  & ~\u0_w_reg[3][15]/P0001  ;
  assign n15754 = ~\u0_w_reg[3][14]/P0001  & n15735 ;
  assign n15755 = n15719 & n15754 ;
  assign n15762 = ~n15753 & ~n15755 ;
  assign n15763 = ~n15761 & n15762 ;
  assign n15764 = n15760 & n15763 ;
  assign n15765 = ~n15750 & ~n15764 ;
  assign n15707 = \u0_w_reg[3][10]/P0001  & ~n15706 ;
  assign n15709 = ~\u0_w_reg[3][11]/P0001  & ~\u0_w_reg[3][12]/P0001  ;
  assign n15710 = n15708 & n15709 ;
  assign n15711 = ~\u0_w_reg[3][15]/P0001  & n15710 ;
  assign n15712 = n15707 & ~n15711 ;
  assign n15716 = ~\u0_w_reg[3][12]/P0001  & \u0_w_reg[3][14]/P0001  ;
  assign n15717 = n15714 & n15716 ;
  assign n15718 = ~n15715 & ~n15717 ;
  assign n15720 = ~\u0_w_reg[3][12]/P0001  & n15719 ;
  assign n15721 = ~\u0_w_reg[3][10]/P0001  & ~n15720 ;
  assign n15722 = n15718 & n15721 ;
  assign n15723 = ~n15712 & ~n15722 ;
  assign n15726 = ~\u0_w_reg[3][10]/P0001  & \u0_w_reg[3][9]/P0001  ;
  assign n15727 = ~n15725 & ~n15726 ;
  assign n15724 = \u0_w_reg[3][11]/P0001  & ~\u0_w_reg[3][12]/P0001  ;
  assign n15728 = \u0_w_reg[3][13]/P0001  & n15724 ;
  assign n15729 = ~n15727 & n15728 ;
  assign n15766 = \u0_w_reg[3][8]/P0001  & ~n15729 ;
  assign n15730 = ~\u0_w_reg[3][10]/P0001  & n15708 ;
  assign n15731 = n15703 & n15730 ;
  assign n15732 = ~\u0_w_reg[3][13]/P0001  & ~n15716 ;
  assign n15733 = ~n15703 & n15726 ;
  assign n15734 = n15732 & n15733 ;
  assign n15767 = ~n15731 & ~n15734 ;
  assign n15768 = n15766 & n15767 ;
  assign n15769 = ~n15723 & n15768 ;
  assign n15770 = ~n15765 & n15769 ;
  assign n15771 = ~\u0_w_reg[3][12]/P0001  & n15725 ;
  assign n15772 = ~\u0_w_reg[3][11]/P0001  & n15771 ;
  assign n15773 = \u0_w_reg[3][13]/P0001  & ~\u0_w_reg[3][14]/P0001  ;
  assign n15774 = n15751 & n15773 ;
  assign n15775 = ~n15743 & ~n15774 ;
  assign n15776 = ~n15772 & n15775 ;
  assign n15777 = ~\u0_w_reg[3][10]/P0001  & ~n15776 ;
  assign n15791 = \u0_w_reg[3][10]/P0001  & n15713 ;
  assign n15792 = n15757 & n15791 ;
  assign n15786 = \u0_w_reg[3][14]/P0001  & \u0_w_reg[3][15]/P0001  ;
  assign n15787 = ~\u0_w_reg[3][13]/P0001  & n15786 ;
  assign n15788 = ~\u0_w_reg[3][11]/P0001  & n15787 ;
  assign n15789 = n15714 & n15756 ;
  assign n15790 = \u0_w_reg[3][9]/P0001  & ~n15789 ;
  assign n15794 = ~n15788 & n15790 ;
  assign n15795 = ~n15792 & n15794 ;
  assign n15784 = ~\u0_w_reg[3][11]/P0001  & n15741 ;
  assign n15785 = ~\u0_w_reg[3][12]/P0001  & n15784 ;
  assign n15778 = ~\u0_w_reg[3][12]/P0001  & \u0_w_reg[3][15]/P0001  ;
  assign n15779 = n15773 & n15778 ;
  assign n15780 = \u0_w_reg[3][13]/P0001  & \u0_w_reg[3][15]/P0001  ;
  assign n15781 = \u0_w_reg[3][11]/P0001  & n15780 ;
  assign n15782 = ~\u0_w_reg[3][10]/P0001  & ~\u0_w_reg[3][12]/P0001  ;
  assign n15783 = n15781 & ~n15782 ;
  assign n15793 = ~n15779 & ~n15783 ;
  assign n15796 = ~n15785 & n15793 ;
  assign n15797 = n15795 & n15796 ;
  assign n15798 = ~n15777 & n15797 ;
  assign n15805 = n15716 & n15780 ;
  assign n15802 = n15703 & n15756 ;
  assign n15803 = \u0_w_reg[3][10]/P0001  & ~\u0_w_reg[3][13]/P0001  ;
  assign n15804 = n15736 & n15803 ;
  assign n15806 = ~n15802 & ~n15804 ;
  assign n15807 = ~n15805 & n15806 ;
  assign n15808 = ~\u0_w_reg[3][11]/P0001  & ~n15807 ;
  assign n15799 = \u0_w_reg[3][10]/P0001  & \u0_w_reg[3][11]/P0001  ;
  assign n15800 = ~\u0_w_reg[3][12]/P0001  & n15799 ;
  assign n15801 = n15756 & n15800 ;
  assign n15809 = ~\u0_w_reg[3][9]/P0001  & ~n15801 ;
  assign n15810 = ~n15808 & n15809 ;
  assign n15811 = ~n15798 & ~n15810 ;
  assign n15812 = ~\u0_w_reg[3][13]/P0001  & n15757 ;
  assign n15813 = \u0_w_reg[3][11]/P0001  & n15812 ;
  assign n15814 = ~\u0_w_reg[3][13]/P0001  & \u0_w_reg[3][15]/P0001  ;
  assign n15815 = n15716 & n15814 ;
  assign n15816 = ~n15813 & ~n15815 ;
  assign n15817 = n15703 & n15773 ;
  assign n15818 = ~\u0_w_reg[3][10]/P0001  & ~n15817 ;
  assign n15819 = n15816 & n15818 ;
  assign n15821 = \u0_w_reg[3][12]/P0001  & n15780 ;
  assign n15822 = ~\u0_w_reg[3][12]/P0001  & ~\u0_w_reg[3][15]/P0001  ;
  assign n15823 = ~\u0_w_reg[3][13]/P0001  & n15822 ;
  assign n15824 = ~n15821 & ~n15823 ;
  assign n15825 = \u0_w_reg[3][11]/P0001  & ~n15824 ;
  assign n15826 = n15708 & n15757 ;
  assign n15827 = ~\u0_w_reg[3][11]/P0001  & n15826 ;
  assign n15820 = ~\u0_w_reg[3][12]/P0001  & n15736 ;
  assign n15828 = \u0_w_reg[3][10]/P0001  & ~n15820 ;
  assign n15829 = ~n15827 & n15828 ;
  assign n15830 = ~n15825 & n15829 ;
  assign n15831 = ~n15819 & ~n15830 ;
  assign n15832 = n15756 & n15822 ;
  assign n15833 = ~\u0_w_reg[3][8]/P0001  & ~n15832 ;
  assign n15834 = ~n15831 & n15833 ;
  assign n15835 = ~n15811 & n15834 ;
  assign n15836 = ~n15770 & ~n15835 ;
  assign n15837 = n15735 & n15773 ;
  assign n15840 = \u0_w_reg[3][13]/P0001  & n15786 ;
  assign n15838 = ~\u0_w_reg[3][13]/P0001  & n15725 ;
  assign n15839 = ~\u0_w_reg[3][13]/P0001  & n15742 ;
  assign n15841 = ~n15838 & ~n15839 ;
  assign n15842 = ~n15840 & n15841 ;
  assign n15843 = n15751 & ~n15842 ;
  assign n15844 = ~n15837 & ~n15843 ;
  assign n15845 = \u0_w_reg[3][10]/P0001  & ~n15844 ;
  assign n15849 = ~\u0_w_reg[3][10]/P0001  & \u0_w_reg[3][11]/P0001  ;
  assign n15850 = \u0_w_reg[3][12]/P0001  & n15725 ;
  assign n15851 = \u0_w_reg[3][13]/P0001  & n15850 ;
  assign n15852 = n15849 & n15851 ;
  assign n15846 = ~\u0_w_reg[3][12]/P0001  & n15780 ;
  assign n15847 = ~\u0_w_reg[3][10]/P0001  & ~\u0_w_reg[3][11]/P0001  ;
  assign n15848 = n15846 & n15847 ;
  assign n15853 = n15709 & n15736 ;
  assign n15854 = ~n15731 & ~n15853 ;
  assign n15855 = ~n15848 & n15854 ;
  assign n15856 = ~n15852 & n15855 ;
  assign n15857 = ~n15845 & n15856 ;
  assign n15858 = ~\u0_w_reg[3][9]/P0001  & ~n15857 ;
  assign n15868 = ~\u0_w_reg[3][11]/P0001  & n15792 ;
  assign n15865 = n15724 & n15736 ;
  assign n15866 = ~\u0_w_reg[3][13]/P0001  & n15865 ;
  assign n15867 = ~\u0_w_reg[3][10]/P0001  & n15817 ;
  assign n15869 = ~n15866 & ~n15867 ;
  assign n15870 = ~n15868 & n15869 ;
  assign n15871 = \u0_w_reg[3][9]/P0001  & ~n15870 ;
  assign n15872 = ~\u0_w_reg[3][10]/P0001  & n15788 ;
  assign n15859 = n15719 & n15735 ;
  assign n15860 = \u0_w_reg[3][10]/P0001  & ~\u0_w_reg[3][14]/P0001  ;
  assign n15861 = n15859 & n15860 ;
  assign n15862 = ~\u0_w_reg[3][14]/P0001  & n15724 ;
  assign n15863 = n15719 & n15862 ;
  assign n15864 = ~\u0_w_reg[3][10]/P0001  & n15863 ;
  assign n15873 = ~n15861 & ~n15864 ;
  assign n15874 = ~n15872 & n15873 ;
  assign n15875 = ~n15871 & n15874 ;
  assign n15876 = ~n15858 & n15875 ;
  assign n15877 = ~n15836 & n15876 ;
  assign n15878 = \u0_w_reg[0][21]/P0001  & ~n15877 ;
  assign n15879 = ~\u0_w_reg[0][21]/P0001  & n15877 ;
  assign n15880 = ~n15878 & ~n15879 ;
  assign n15881 = \u0_w_reg[1][21]/P0001  & ~\u0_w_reg[2][21]/P0001  ;
  assign n15882 = ~\u0_w_reg[1][21]/P0001  & \u0_w_reg[2][21]/P0001  ;
  assign n15883 = ~n15881 & ~n15882 ;
  assign n15884 = n15880 & n15883 ;
  assign n15885 = ~n15880 & ~n15883 ;
  assign n15886 = ~n15884 & ~n15885 ;
  assign n15887 = ~ld_pad & n15886 ;
  assign n15888 = ~n15702 & ~n15887 ;
  assign n15889 = ~\key[51]_pad  & ld_pad ;
  assign n15927 = ~n15720 & n15745 ;
  assign n15928 = \u0_w_reg[3][10]/P0001  & ~n15927 ;
  assign n15929 = \u0_w_reg[3][13]/P0001  & n15709 ;
  assign n15930 = \u0_w_reg[3][14]/P0001  & n15929 ;
  assign n15933 = ~n15853 & ~n15930 ;
  assign n15931 = n15838 & n15849 ;
  assign n15932 = \u0_w_reg[3][11]/P0001  & n15802 ;
  assign n15934 = ~n15931 & ~n15932 ;
  assign n15935 = n15933 & n15934 ;
  assign n15936 = ~n15872 & n15935 ;
  assign n15937 = ~n15928 & n15936 ;
  assign n15938 = ~\u0_w_reg[3][9]/P0001  & ~n15937 ;
  assign n15943 = ~\u0_w_reg[3][13]/P0001  & n15736 ;
  assign n15942 = ~\u0_w_reg[3][11]/P0001  & n15725 ;
  assign n15944 = ~\u0_w_reg[3][10]/P0001  & ~n15942 ;
  assign n15945 = ~n15943 & n15944 ;
  assign n15947 = ~n15714 & n15773 ;
  assign n15946 = \u0_w_reg[3][12]/P0001  & n15814 ;
  assign n15948 = \u0_w_reg[3][10]/P0001  & ~n15946 ;
  assign n15949 = ~n15947 & n15948 ;
  assign n15950 = ~n15945 & ~n15949 ;
  assign n15919 = \u0_w_reg[3][11]/P0001  & \u0_w_reg[3][14]/P0001  ;
  assign n15939 = n15814 & n15919 ;
  assign n15940 = ~n15817 & ~n15939 ;
  assign n15941 = n15751 & n15780 ;
  assign n15951 = n15940 & ~n15941 ;
  assign n15952 = ~n15950 & n15951 ;
  assign n15953 = \u0_w_reg[3][9]/P0001  & ~n15952 ;
  assign n15960 = n15735 & n15742 ;
  assign n15961 = ~n15802 & ~n15826 ;
  assign n15962 = ~n15960 & n15961 ;
  assign n15963 = \u0_w_reg[3][10]/P0001  & ~n15962 ;
  assign n15896 = ~\u0_w_reg[3][11]/P0001  & n15778 ;
  assign n15897 = ~\u0_w_reg[3][13]/P0001  & n15896 ;
  assign n15954 = n15780 & n15919 ;
  assign n15955 = ~n15897 & ~n15954 ;
  assign n15956 = ~\u0_w_reg[3][10]/P0001  & ~n15955 ;
  assign n15957 = n15713 & n15724 ;
  assign n15958 = ~\u0_w_reg[3][15]/P0001  & n15957 ;
  assign n15959 = ~\u0_w_reg[3][11]/P0001  & n15867 ;
  assign n15964 = ~n15958 & ~n15959 ;
  assign n15965 = ~n15956 & n15964 ;
  assign n15966 = ~n15963 & n15965 ;
  assign n15967 = ~n15953 & n15966 ;
  assign n15968 = ~n15938 & n15967 ;
  assign n15969 = \u0_w_reg[3][8]/P0001  & ~n15968 ;
  assign n15892 = \u0_w_reg[3][11]/P0001  & n15867 ;
  assign n15890 = ~n15756 & ~n15860 ;
  assign n15891 = n15757 & ~n15890 ;
  assign n15898 = ~\u0_w_reg[3][9]/P0001  & ~n15891 ;
  assign n15893 = \u0_w_reg[3][10]/P0001  & ~\u0_w_reg[3][11]/P0001  ;
  assign n15894 = \u0_w_reg[3][15]/P0001  & ~n15756 ;
  assign n15895 = n15893 & n15894 ;
  assign n15899 = ~n15895 & ~n15897 ;
  assign n15900 = n15898 & n15899 ;
  assign n15901 = ~n15892 & n15900 ;
  assign n15902 = n15713 & n15751 ;
  assign n15903 = ~\u0_w_reg[3][15]/P0001  & n15902 ;
  assign n15904 = ~n15823 & ~n15903 ;
  assign n15905 = \u0_w_reg[3][10]/P0001  & ~n15904 ;
  assign n15906 = \u0_w_reg[3][15]/P0001  & n15735 ;
  assign n15907 = ~n15896 & ~n15906 ;
  assign n15908 = n15713 & ~n15907 ;
  assign n15909 = ~\u0_w_reg[3][10]/P0001  & n15779 ;
  assign n15910 = \u0_w_reg[3][9]/P0001  & ~n15744 ;
  assign n15911 = ~n15909 & n15910 ;
  assign n15912 = ~n15908 & n15911 ;
  assign n15913 = ~n15905 & n15912 ;
  assign n15914 = ~n15901 & ~n15913 ;
  assign n15920 = n15757 & n15919 ;
  assign n15921 = ~n15706 & ~n15920 ;
  assign n15922 = ~\u0_w_reg[3][10]/P0001  & ~n15921 ;
  assign n15915 = ~\u0_w_reg[3][12]/P0001  & n15714 ;
  assign n15916 = ~\u0_w_reg[3][13]/P0001  & n15915 ;
  assign n15917 = ~n15805 & ~n15916 ;
  assign n15918 = \u0_w_reg[3][10]/P0001  & ~n15917 ;
  assign n15923 = ~n15711 & ~n15918 ;
  assign n15924 = ~n15922 & n15923 ;
  assign n15925 = ~n15914 & n15924 ;
  assign n15926 = ~\u0_w_reg[3][8]/P0001  & ~n15925 ;
  assign n15987 = n15940 & ~n15957 ;
  assign n15988 = \u0_w_reg[3][10]/P0001  & ~n15987 ;
  assign n15983 = \u0_w_reg[3][12]/P0001  & n15756 ;
  assign n15984 = ~n15771 & ~n15779 ;
  assign n15985 = ~n15983 & n15984 ;
  assign n15986 = n15847 & ~n15985 ;
  assign n15989 = n15756 & n15778 ;
  assign n15990 = n15849 & n15989 ;
  assign n15991 = ~n15986 & ~n15990 ;
  assign n15992 = ~n15988 & n15991 ;
  assign n15993 = \u0_w_reg[3][9]/P0001  & ~n15992 ;
  assign n15970 = n15724 & n15786 ;
  assign n15971 = ~\u0_w_reg[3][13]/P0001  & n15970 ;
  assign n15972 = ~n15932 & ~n15971 ;
  assign n15973 = \u0_w_reg[3][10]/P0001  & ~n15972 ;
  assign n15974 = \u0_w_reg[3][10]/P0001  & ~\u0_w_reg[3][9]/P0001  ;
  assign n15975 = ~\u0_w_reg[3][11]/P0001  & n15974 ;
  assign n15976 = n15708 & n15822 ;
  assign n15977 = ~n15758 & ~n15976 ;
  assign n15978 = n15975 & ~n15977 ;
  assign n15979 = ~\u0_w_reg[3][10]/P0001  & ~\u0_w_reg[3][9]/P0001  ;
  assign n15980 = n15778 & n15979 ;
  assign n15981 = ~n15812 & ~n15980 ;
  assign n15982 = n15919 & ~n15981 ;
  assign n15994 = ~n15978 & ~n15982 ;
  assign n15995 = ~n15973 & n15994 ;
  assign n15996 = ~n15993 & n15995 ;
  assign n15997 = ~n15926 & n15996 ;
  assign n15998 = ~n15969 & n15997 ;
  assign n15999 = \u0_w_reg[0][19]/P0001  & ~n15998 ;
  assign n16000 = ~\u0_w_reg[0][19]/P0001  & n15998 ;
  assign n16001 = ~n15999 & ~n16000 ;
  assign n16002 = \u0_w_reg[1][19]/P0001  & ~\u0_w_reg[2][19]/P0001  ;
  assign n16003 = ~\u0_w_reg[1][19]/P0001  & \u0_w_reg[2][19]/P0001  ;
  assign n16004 = ~n16002 & ~n16003 ;
  assign n16005 = n16001 & n16004 ;
  assign n16006 = ~n16001 & ~n16004 ;
  assign n16007 = ~n16005 & ~n16006 ;
  assign n16008 = ~ld_pad & n16007 ;
  assign n16009 = ~n15889 & ~n16008 ;
  assign n16010 = ~\key[37]_pad  & ld_pad ;
  assign n16043 = ~\u0_w_reg[3][30]/P0001  & \u0_w_reg[3][31]/P0001  ;
  assign n16048 = ~\u0_w_reg[3][27]/P0001  & \u0_w_reg[3][28]/P0001  ;
  assign n16124 = n16043 & n16048 ;
  assign n16051 = ~\u0_w_reg[3][30]/P0001  & ~\u0_w_reg[3][31]/P0001  ;
  assign n16125 = ~\u0_w_reg[3][27]/P0001  & n16051 ;
  assign n16126 = \u0_w_reg[3][26]/P0001  & n16125 ;
  assign n16127 = ~n16124 & ~n16126 ;
  assign n16128 = ~\u0_w_reg[3][29]/P0001  & ~n16127 ;
  assign n16011 = \u0_w_reg[3][29]/P0001  & \u0_w_reg[3][30]/P0001  ;
  assign n16037 = \u0_w_reg[3][31]/P0001  & n16011 ;
  assign n16129 = ~\u0_w_reg[3][27]/P0001  & n16037 ;
  assign n16130 = ~\u0_w_reg[3][28]/P0001  & n16129 ;
  assign n16094 = ~\u0_w_reg[3][29]/P0001  & ~\u0_w_reg[3][30]/P0001  ;
  assign n16121 = ~\u0_w_reg[3][28]/P0001  & n16094 ;
  assign n16122 = \u0_w_reg[3][26]/P0001  & \u0_w_reg[3][27]/P0001  ;
  assign n16123 = n16121 & n16122 ;
  assign n16131 = ~\u0_w_reg[3][25]/P0001  & ~n16123 ;
  assign n16132 = ~n16130 & n16131 ;
  assign n16133 = ~n16128 & n16132 ;
  assign n16079 = \u0_w_reg[3][29]/P0001  & ~\u0_w_reg[3][30]/P0001  ;
  assign n16134 = n16048 & n16079 ;
  assign n16087 = ~\u0_w_reg[3][27]/P0001  & ~\u0_w_reg[3][28]/P0001  ;
  assign n16135 = ~n16043 & ~n16087 ;
  assign n16025 = \u0_w_reg[3][30]/P0001  & ~\u0_w_reg[3][31]/P0001  ;
  assign n16136 = ~\u0_w_reg[3][27]/P0001  & ~n16025 ;
  assign n16137 = ~n16135 & ~n16136 ;
  assign n16138 = ~n16134 & ~n16137 ;
  assign n16139 = ~\u0_w_reg[3][26]/P0001  & ~n16138 ;
  assign n16098 = \u0_w_reg[3][30]/P0001  & \u0_w_reg[3][31]/P0001  ;
  assign n16099 = ~\u0_w_reg[3][29]/P0001  & n16098 ;
  assign n16100 = ~\u0_w_reg[3][27]/P0001  & n16099 ;
  assign n16149 = \u0_w_reg[3][25]/P0001  & ~n16100 ;
  assign n16026 = ~\u0_w_reg[3][28]/P0001  & \u0_w_reg[3][29]/P0001  ;
  assign n16140 = ~\u0_w_reg[3][27]/P0001  & n16025 ;
  assign n16141 = n16026 & n16140 ;
  assign n16012 = \u0_w_reg[3][27]/P0001  & ~\u0_w_reg[3][31]/P0001  ;
  assign n16144 = n16012 & n16094 ;
  assign n16150 = n16026 & n16043 ;
  assign n16151 = ~n16144 & ~n16150 ;
  assign n16152 = ~n16141 & n16151 ;
  assign n16105 = \u0_w_reg[3][28]/P0001  & ~\u0_w_reg[3][31]/P0001  ;
  assign n16142 = \u0_w_reg[3][26]/P0001  & n16011 ;
  assign n16143 = n16105 & n16142 ;
  assign n16145 = \u0_w_reg[3][29]/P0001  & \u0_w_reg[3][31]/P0001  ;
  assign n16146 = \u0_w_reg[3][27]/P0001  & n16145 ;
  assign n16147 = ~\u0_w_reg[3][26]/P0001  & ~\u0_w_reg[3][28]/P0001  ;
  assign n16148 = n16146 & ~n16147 ;
  assign n16153 = ~n16143 & ~n16148 ;
  assign n16154 = n16152 & n16153 ;
  assign n16155 = n16149 & n16154 ;
  assign n16156 = ~n16139 & n16155 ;
  assign n16157 = ~n16133 & ~n16156 ;
  assign n16039 = ~\u0_w_reg[3][28]/P0001  & ~\u0_w_reg[3][31]/P0001  ;
  assign n16120 = n16039 & n16094 ;
  assign n16019 = ~\u0_w_reg[3][29]/P0001  & \u0_w_reg[3][30]/P0001  ;
  assign n16160 = \u0_w_reg[3][28]/P0001  & n16019 ;
  assign n16161 = ~\u0_w_reg[3][31]/P0001  & n16160 ;
  assign n16162 = ~\u0_w_reg[3][27]/P0001  & n16161 ;
  assign n16093 = ~\u0_w_reg[3][28]/P0001  & n16012 ;
  assign n16165 = ~\u0_w_reg[3][29]/P0001  & n16093 ;
  assign n16045 = \u0_w_reg[3][27]/P0001  & \u0_w_reg[3][28]/P0001  ;
  assign n16158 = \u0_w_reg[3][31]/P0001  & n16045 ;
  assign n16159 = \u0_w_reg[3][29]/P0001  & n16158 ;
  assign n16163 = ~\u0_w_reg[3][28]/P0001  & n16051 ;
  assign n16164 = \u0_w_reg[3][26]/P0001  & ~n16163 ;
  assign n16166 = ~n16159 & n16164 ;
  assign n16167 = ~n16165 & n16166 ;
  assign n16168 = ~n16162 & n16167 ;
  assign n16169 = ~\u0_w_reg[3][29]/P0001  & n16105 ;
  assign n16170 = \u0_w_reg[3][27]/P0001  & n16169 ;
  assign n16014 = ~\u0_w_reg[3][28]/P0001  & \u0_w_reg[3][30]/P0001  ;
  assign n16171 = ~\u0_w_reg[3][29]/P0001  & \u0_w_reg[3][31]/P0001  ;
  assign n16172 = n16014 & n16171 ;
  assign n16173 = ~n16170 & ~n16172 ;
  assign n16020 = \u0_w_reg[3][28]/P0001  & \u0_w_reg[3][31]/P0001  ;
  assign n16091 = n16020 & n16079 ;
  assign n16174 = ~\u0_w_reg[3][26]/P0001  & ~n16091 ;
  assign n16175 = n16173 & n16174 ;
  assign n16176 = ~n16168 & ~n16175 ;
  assign n16177 = ~n16120 & ~n16176 ;
  assign n16178 = ~n16157 & n16177 ;
  assign n16179 = ~\u0_w_reg[3][24]/P0001  & ~n16178 ;
  assign n16058 = \u0_w_reg[3][29]/P0001  & n16025 ;
  assign n16059 = ~\u0_w_reg[3][29]/P0001  & n16043 ;
  assign n16060 = \u0_w_reg[3][27]/P0001  & n16059 ;
  assign n16061 = ~n16058 & ~n16060 ;
  assign n16062 = ~\u0_w_reg[3][26]/P0001  & ~n16061 ;
  assign n16065 = ~\u0_w_reg[3][29]/P0001  & n16014 ;
  assign n16066 = n16045 & n16051 ;
  assign n16067 = ~n16065 & ~n16066 ;
  assign n16068 = \u0_w_reg[3][26]/P0001  & ~n16067 ;
  assign n16013 = n16011 & n16012 ;
  assign n16063 = n16011 & n16048 ;
  assign n16064 = \u0_w_reg[3][31]/P0001  & n16063 ;
  assign n16069 = ~n16013 & ~n16064 ;
  assign n16070 = ~n16068 & n16069 ;
  assign n16071 = ~n16062 & n16070 ;
  assign n16072 = ~\u0_w_reg[3][25]/P0001  & ~n16071 ;
  assign n16032 = \u0_w_reg[3][27]/P0001  & ~\u0_w_reg[3][28]/P0001  ;
  assign n16044 = n16032 & n16043 ;
  assign n16017 = \u0_w_reg[3][29]/P0001  & ~\u0_w_reg[3][31]/P0001  ;
  assign n16046 = ~\u0_w_reg[3][30]/P0001  & n16045 ;
  assign n16047 = n16017 & n16046 ;
  assign n16054 = ~n16044 & ~n16047 ;
  assign n16049 = \u0_w_reg[3][29]/P0001  & n16043 ;
  assign n16050 = n16048 & n16049 ;
  assign n16052 = ~\u0_w_reg[3][29]/P0001  & n16051 ;
  assign n16053 = n16048 & n16052 ;
  assign n16055 = ~n16050 & ~n16053 ;
  assign n16056 = n16054 & n16055 ;
  assign n16057 = \u0_w_reg[3][25]/P0001  & ~n16056 ;
  assign n16015 = n16012 & n16014 ;
  assign n16016 = ~n16013 & ~n16015 ;
  assign n16018 = ~\u0_w_reg[3][28]/P0001  & n16017 ;
  assign n16021 = n16019 & n16020 ;
  assign n16022 = ~n16018 & ~n16021 ;
  assign n16023 = n16016 & n16022 ;
  assign n16024 = ~\u0_w_reg[3][26]/P0001  & ~n16023 ;
  assign n16027 = n16025 & n16026 ;
  assign n16028 = \u0_w_reg[3][27]/P0001  & n16027 ;
  assign n16073 = ~n16024 & ~n16028 ;
  assign n16029 = \u0_w_reg[3][25]/P0001  & ~\u0_w_reg[3][26]/P0001  ;
  assign n16030 = ~\u0_w_reg[3][29]/P0001  & ~n16014 ;
  assign n16031 = ~n16020 & n16030 ;
  assign n16033 = \u0_w_reg[3][29]/P0001  & n16032 ;
  assign n16034 = ~n16031 & ~n16033 ;
  assign n16035 = n16029 & ~n16034 ;
  assign n16036 = \u0_w_reg[3][26]/P0001  & ~\u0_w_reg[3][27]/P0001  ;
  assign n16038 = \u0_w_reg[3][28]/P0001  & n16037 ;
  assign n16040 = n16019 & n16039 ;
  assign n16041 = ~n16038 & ~n16040 ;
  assign n16042 = n16036 & ~n16041 ;
  assign n16074 = ~n16035 & ~n16042 ;
  assign n16075 = n16073 & n16074 ;
  assign n16076 = ~n16057 & n16075 ;
  assign n16077 = ~n16072 & n16076 ;
  assign n16078 = \u0_w_reg[3][24]/P0001  & ~n16077 ;
  assign n16080 = n16045 & n16079 ;
  assign n16081 = ~\u0_w_reg[3][29]/P0001  & n16025 ;
  assign n16082 = ~n16037 & ~n16059 ;
  assign n16083 = ~n16081 & n16082 ;
  assign n16084 = n16048 & ~n16083 ;
  assign n16085 = ~n16080 & ~n16084 ;
  assign n16086 = \u0_w_reg[3][26]/P0001  & ~n16085 ;
  assign n16088 = n16051 & n16087 ;
  assign n16089 = ~n16086 & ~n16088 ;
  assign n16090 = ~\u0_w_reg[3][25]/P0001  & ~n16089 ;
  assign n16109 = ~\u0_w_reg[3][25]/P0001  & ~\u0_w_reg[3][26]/P0001  ;
  assign n16112 = \u0_w_reg[3][29]/P0001  & n16087 ;
  assign n16113 = \u0_w_reg[3][31]/P0001  & n16112 ;
  assign n16110 = n16011 & n16045 ;
  assign n16111 = ~\u0_w_reg[3][31]/P0001  & n16110 ;
  assign n16114 = ~n16021 & ~n16111 ;
  assign n16115 = ~n16113 & n16114 ;
  assign n16116 = n16109 & ~n16115 ;
  assign n16092 = ~\u0_w_reg[3][26]/P0001  & n16091 ;
  assign n16095 = n16093 & n16094 ;
  assign n16096 = ~n16092 & ~n16095 ;
  assign n16097 = \u0_w_reg[3][25]/P0001  & ~n16096 ;
  assign n16101 = ~\u0_w_reg[3][26]/P0001  & n16100 ;
  assign n16117 = ~\u0_w_reg[3][26]/P0001  & \u0_w_reg[3][27]/P0001  ;
  assign n16118 = n16026 & n16051 ;
  assign n16119 = n16117 & n16118 ;
  assign n16102 = n16017 & n16045 ;
  assign n16103 = \u0_w_reg[3][26]/P0001  & ~\u0_w_reg[3][30]/P0001  ;
  assign n16104 = n16102 & n16103 ;
  assign n16106 = n16036 & n16105 ;
  assign n16107 = \u0_w_reg[3][25]/P0001  & n16011 ;
  assign n16108 = n16106 & n16107 ;
  assign n16180 = ~n16104 & ~n16108 ;
  assign n16181 = ~n16119 & n16180 ;
  assign n16182 = ~n16101 & n16181 ;
  assign n16183 = ~n16097 & n16182 ;
  assign n16184 = ~n16116 & n16183 ;
  assign n16185 = ~n16090 & n16184 ;
  assign n16186 = ~n16078 & n16185 ;
  assign n16187 = ~n16179 & n16186 ;
  assign n16188 = \u0_w_reg[0][5]/P0001  & ~n16187 ;
  assign n16189 = ~\u0_w_reg[0][5]/P0001  & n16187 ;
  assign n16190 = ~n16188 & ~n16189 ;
  assign n16191 = \u0_w_reg[1][5]/P0001  & ~\u0_w_reg[2][5]/P0001  ;
  assign n16192 = ~\u0_w_reg[1][5]/P0001  & \u0_w_reg[2][5]/P0001  ;
  assign n16193 = ~n16191 & ~n16192 ;
  assign n16194 = n16190 & n16193 ;
  assign n16195 = ~n16190 & ~n16193 ;
  assign n16196 = ~n16194 & ~n16195 ;
  assign n16197 = ~ld_pad & n16196 ;
  assign n16198 = ~n16010 & ~n16197 ;
  assign n16199 = \u0_w_reg[0][10]/P0001  & ~n15068 ;
  assign n16200 = ~\u0_w_reg[0][10]/P0001  & n15068 ;
  assign n16201 = ~n16199 & ~n16200 ;
  assign n16202 = n13752 & n16201 ;
  assign n16203 = ~n13752 & ~n16201 ;
  assign n16204 = ~n16202 & ~n16203 ;
  assign n16205 = n13835 & n14804 ;
  assign n16206 = ~n13835 & ~n14804 ;
  assign n16207 = ~n16205 & ~n16206 ;
  assign n16209 = n16204 & n16207 ;
  assign n16208 = ~n16204 & ~n16207 ;
  assign n16210 = ~\ld_r_reg/P0001  & ~n16208 ;
  assign n16211 = ~n16209 & n16210 ;
  assign n16213 = ~\text_in_r_reg[106]/P0001  & \u0_w_reg[0][10]/P0001  ;
  assign n16212 = \text_in_r_reg[106]/P0001  & ~\u0_w_reg[0][10]/P0001  ;
  assign n16214 = \ld_r_reg/P0001  & ~n16212 ;
  assign n16215 = ~n16213 & n16214 ;
  assign n16216 = ~n16211 & ~n16215 ;
  assign n16287 = n15503 & n15521 ;
  assign n16306 = ~n15528 & ~n16287 ;
  assign n16307 = ~\u0_w_reg[3][18]/P0001  & n16306 ;
  assign n16309 = \u0_w_reg[3][22]/P0001  & n15525 ;
  assign n16310 = n15542 & n16309 ;
  assign n16311 = ~n15614 & ~n16310 ;
  assign n16312 = \u0_w_reg[3][17]/P0001  & ~n16311 ;
  assign n16308 = \u0_w_reg[3][19]/P0001  & n15614 ;
  assign n16313 = n15526 & n15539 ;
  assign n16314 = \u0_w_reg[3][18]/P0001  & ~n16313 ;
  assign n16315 = ~n16308 & n16314 ;
  assign n16316 = ~n16312 & n16315 ;
  assign n16317 = ~n16307 & ~n16316 ;
  assign n16290 = ~\u0_w_reg[3][18]/P0001  & n15583 ;
  assign n16291 = \u0_w_reg[3][17]/P0001  & ~n15607 ;
  assign n16217 = \u0_w_reg[3][19]/P0001  & n15531 ;
  assign n16229 = \u0_w_reg[3][19]/P0001  & \u0_w_reg[3][22]/P0001  ;
  assign n16242 = n15526 & n16229 ;
  assign n16289 = \u0_w_reg[3][20]/P0001  & n16242 ;
  assign n16292 = ~n16217 & ~n16289 ;
  assign n16293 = n16291 & n16292 ;
  assign n16294 = ~n16290 & n16293 ;
  assign n16300 = \u0_w_reg[3][19]/P0001  & n15629 ;
  assign n16297 = \u0_w_reg[3][18]/P0001  & ~\u0_w_reg[3][22]/P0001  ;
  assign n16298 = ~n15549 & ~n16297 ;
  assign n16299 = n15551 & ~n16298 ;
  assign n16295 = \u0_w_reg[3][23]/P0001  & n15511 ;
  assign n16296 = ~n15549 & n16295 ;
  assign n16241 = n15506 & n15601 ;
  assign n16301 = ~\u0_w_reg[3][17]/P0001  & ~n16241 ;
  assign n16302 = ~n16296 & n16301 ;
  assign n16303 = ~n16299 & n16302 ;
  assign n16304 = ~n16300 & n16303 ;
  assign n16305 = ~n16294 & ~n16304 ;
  assign n16318 = ~\u0_w_reg[3][21]/P0001  & n15574 ;
  assign n16319 = ~n16305 & ~n16318 ;
  assign n16320 = ~n16317 & n16319 ;
  assign n16321 = ~\u0_w_reg[3][16]/P0001  & ~n16320 ;
  assign n16245 = ~n15537 & n15559 ;
  assign n16246 = ~n15602 & ~n16245 ;
  assign n16247 = \u0_w_reg[3][17]/P0001  & ~n16246 ;
  assign n16248 = \u0_w_reg[3][23]/P0001  & n15521 ;
  assign n16249 = ~\u0_w_reg[3][22]/P0001  & n16248 ;
  assign n16250 = ~n15603 & ~n15618 ;
  assign n16251 = ~n16249 & n16250 ;
  assign n16252 = ~n16247 & n16251 ;
  assign n16253 = \u0_w_reg[3][18]/P0001  & ~n16252 ;
  assign n16218 = ~n15516 & ~n15543 ;
  assign n16219 = ~n16217 & n16218 ;
  assign n16220 = \u0_w_reg[3][18]/P0001  & ~n16219 ;
  assign n16223 = ~n15580 & ~n15637 ;
  assign n16224 = ~n15661 & n16223 ;
  assign n16221 = n15529 & n15638 ;
  assign n16222 = n15562 & n15601 ;
  assign n16225 = ~n16221 & ~n16222 ;
  assign n16226 = n16224 & n16225 ;
  assign n16227 = ~n16220 & n16226 ;
  assign n16228 = ~\u0_w_reg[3][17]/P0001  & ~n16227 ;
  assign n16232 = ~\u0_w_reg[3][18]/P0001  & n15557 ;
  assign n16230 = n15601 & n16229 ;
  assign n16231 = ~n15628 & ~n16230 ;
  assign n16233 = n15503 & n15648 ;
  assign n16234 = ~n15527 & ~n16233 ;
  assign n16235 = n16231 & n16234 ;
  assign n16236 = ~n16232 & n16235 ;
  assign n16237 = \u0_w_reg[3][17]/P0001  & ~n16236 ;
  assign n16243 = ~n16241 & ~n16242 ;
  assign n16244 = ~\u0_w_reg[3][18]/P0001  & ~n16243 ;
  assign n16238 = n15503 & n15505 ;
  assign n16239 = ~\u0_w_reg[3][18]/P0001  & n15527 ;
  assign n16240 = ~\u0_w_reg[3][22]/P0001  & n16239 ;
  assign n16254 = ~n16238 & ~n16240 ;
  assign n16255 = ~n16244 & n16254 ;
  assign n16256 = ~n16237 & n16255 ;
  assign n16257 = ~n16228 & n16256 ;
  assign n16258 = ~n16253 & n16257 ;
  assign n16259 = \u0_w_reg[3][16]/P0001  & ~n16258 ;
  assign n16261 = \u0_w_reg[3][20]/P0001  & n15549 ;
  assign n16262 = ~\u0_w_reg[3][20]/P0001  & n15503 ;
  assign n16263 = ~n16261 & ~n16262 ;
  assign n16264 = ~n15583 & n16263 ;
  assign n16265 = n15648 & ~n16264 ;
  assign n16260 = \u0_w_reg[3][18]/P0001  & ~n16231 ;
  assign n16266 = ~\u0_w_reg[3][20]/P0001  & n15608 ;
  assign n16267 = n15512 & n16266 ;
  assign n16268 = ~\u0_w_reg[3][20]/P0001  & \u0_w_reg[3][23]/P0001  ;
  assign n16269 = n15549 & n16268 ;
  assign n16270 = n15529 & n16269 ;
  assign n16271 = ~n16267 & ~n16270 ;
  assign n16272 = ~n16260 & n16271 ;
  assign n16273 = ~n16265 & n16272 ;
  assign n16274 = \u0_w_reg[3][17]/P0001  & ~n16273 ;
  assign n16281 = ~\u0_w_reg[3][17]/P0001  & \u0_w_reg[3][18]/P0001  ;
  assign n16282 = ~\u0_w_reg[3][19]/P0001  & n16281 ;
  assign n16283 = ~\u0_w_reg[3][23]/P0001  & n15519 ;
  assign n16284 = n15549 & n15551 ;
  assign n16285 = ~n16283 & ~n16284 ;
  assign n16286 = n16282 & ~n16285 ;
  assign n16276 = \u0_w_reg[3][18]/P0001  & n16230 ;
  assign n16277 = ~\u0_w_reg[3][17]/P0001  & n15529 ;
  assign n16278 = n15590 & n16277 ;
  assign n16279 = ~n16276 & ~n16278 ;
  assign n16280 = ~\u0_w_reg[3][20]/P0001  & ~n16279 ;
  assign n16275 = n15603 & n15608 ;
  assign n16288 = ~\u0_w_reg[3][21]/P0001  & n16287 ;
  assign n16322 = ~n16275 & ~n16288 ;
  assign n16323 = ~n16280 & n16322 ;
  assign n16324 = ~n16286 & n16323 ;
  assign n16325 = ~n16274 & n16324 ;
  assign n16326 = ~n16259 & n16325 ;
  assign n16327 = ~n16321 & n16326 ;
  assign n16328 = \u0_r0_out_reg[27]/P0001  & ~\u0_w_reg[0][27]/P0001  ;
  assign n16329 = ~\u0_r0_out_reg[27]/P0001  & \u0_w_reg[0][27]/P0001  ;
  assign n16330 = ~n16328 & ~n16329 ;
  assign n16332 = n16327 & n16330 ;
  assign n16331 = ~n16327 & ~n16330 ;
  assign n16333 = ~ld_pad & ~n16331 ;
  assign n16334 = ~n16332 & n16333 ;
  assign n16335 = \key[123]_pad  & ld_pad ;
  assign n16336 = ~n16334 & ~n16335 ;
  assign n16337 = ~\key[91]_pad  & ld_pad ;
  assign n16338 = \u0_w_reg[1][27]/P0001  & ~n16330 ;
  assign n16339 = ~\u0_w_reg[1][27]/P0001  & n16330 ;
  assign n16340 = ~n16338 & ~n16339 ;
  assign n16341 = n16327 & n16340 ;
  assign n16342 = ~n16327 & ~n16340 ;
  assign n16343 = ~n16341 & ~n16342 ;
  assign n16344 = ~ld_pad & n16343 ;
  assign n16345 = ~n16337 & ~n16344 ;
  assign n16346 = ~\key[59]_pad  & ld_pad ;
  assign n16347 = \u0_w_reg[2][27]/P0001  & n16343 ;
  assign n16348 = ~\u0_w_reg[2][27]/P0001  & ~n16343 ;
  assign n16349 = ~n16347 & ~n16348 ;
  assign n16350 = ~ld_pad & n16349 ;
  assign n16351 = ~n16346 & ~n16350 ;
  assign n16353 = \u0_w_reg[3][27]/P0001  & ~n16349 ;
  assign n16352 = ~\u0_w_reg[3][27]/P0001  & n16349 ;
  assign n16354 = ~ld_pad & ~n16352 ;
  assign n16355 = ~n16353 & n16354 ;
  assign n16356 = \key[27]_pad  & ld_pad ;
  assign n16357 = ~n16355 & ~n16356 ;
  assign n16358 = ~\key[35]_pad  & ld_pad ;
  assign n16372 = ~n16018 & n16061 ;
  assign n16373 = \u0_w_reg[3][26]/P0001  & ~n16372 ;
  assign n16374 = n16081 & n16117 ;
  assign n16377 = ~\u0_w_reg[3][25]/P0001  & ~n16088 ;
  assign n16378 = ~n16374 & n16377 ;
  assign n16375 = \u0_w_reg[3][30]/P0001  & n16112 ;
  assign n16376 = n16094 & n16158 ;
  assign n16379 = ~n16375 & ~n16376 ;
  assign n16380 = n16378 & n16379 ;
  assign n16381 = ~n16101 & n16380 ;
  assign n16382 = ~n16373 & n16381 ;
  assign n16388 = \u0_w_reg[3][28]/P0001  & n16171 ;
  assign n16389 = ~n16012 & n16079 ;
  assign n16390 = ~n16388 & ~n16389 ;
  assign n16391 = \u0_w_reg[3][26]/P0001  & ~n16390 ;
  assign n16383 = ~\u0_w_reg[3][26]/P0001  & n16052 ;
  assign n16384 = \u0_w_reg[3][25]/P0001  & ~n16383 ;
  assign n16392 = \u0_w_reg[3][27]/P0001  & \u0_w_reg[3][30]/P0001  ;
  assign n16393 = n16171 & n16392 ;
  assign n16394 = ~n16091 & ~n16393 ;
  assign n16385 = n16048 & n16145 ;
  assign n16386 = ~\u0_w_reg[3][26]/P0001  & ~\u0_w_reg[3][27]/P0001  ;
  assign n16387 = n16025 & n16386 ;
  assign n16395 = ~n16385 & ~n16387 ;
  assign n16396 = n16394 & n16395 ;
  assign n16397 = n16384 & n16396 ;
  assign n16398 = ~n16391 & n16397 ;
  assign n16399 = ~n16382 & ~n16398 ;
  assign n16362 = \u0_w_reg[3][30]/P0001  & n16146 ;
  assign n16363 = ~n16050 & ~n16362 ;
  assign n16359 = ~\u0_w_reg[3][28]/P0001  & \u0_w_reg[3][31]/P0001  ;
  assign n16360 = ~\u0_w_reg[3][27]/P0001  & n16359 ;
  assign n16361 = ~\u0_w_reg[3][29]/P0001  & n16360 ;
  assign n16364 = ~\u0_w_reg[3][26]/P0001  & ~n16361 ;
  assign n16365 = n16363 & n16364 ;
  assign n16367 = ~\u0_w_reg[3][30]/P0001  & n16158 ;
  assign n16366 = n16020 & n16094 ;
  assign n16368 = \u0_w_reg[3][26]/P0001  & ~n16366 ;
  assign n16369 = ~n16161 & n16368 ;
  assign n16370 = ~n16367 & n16369 ;
  assign n16371 = ~n16365 & ~n16370 ;
  assign n16400 = ~n16028 & ~n16371 ;
  assign n16401 = ~n16399 & n16400 ;
  assign n16402 = \u0_w_reg[3][24]/P0001  & ~n16401 ;
  assign n16406 = ~\u0_w_reg[3][29]/P0001  & n16039 ;
  assign n16407 = n16017 & n16048 ;
  assign n16408 = \u0_w_reg[3][30]/P0001  & n16407 ;
  assign n16409 = ~n16406 & ~n16408 ;
  assign n16410 = \u0_w_reg[3][26]/P0001  & ~n16409 ;
  assign n16414 = \u0_w_reg[3][25]/P0001  & ~n16060 ;
  assign n16411 = ~n16045 & ~n16087 ;
  assign n16412 = n16037 & ~n16411 ;
  assign n16413 = ~\u0_w_reg[3][26]/P0001  & n16150 ;
  assign n16415 = ~n16412 & ~n16413 ;
  assign n16416 = n16414 & n16415 ;
  assign n16417 = ~n16410 & n16416 ;
  assign n16420 = \u0_w_reg[3][27]/P0001  & n16092 ;
  assign n16423 = ~\u0_w_reg[3][25]/P0001  & ~n16361 ;
  assign n16418 = ~n16094 & ~n16103 ;
  assign n16419 = n16105 & ~n16418 ;
  assign n16421 = \u0_w_reg[3][31]/P0001  & n16036 ;
  assign n16422 = ~n16094 & n16421 ;
  assign n16424 = ~n16419 & ~n16422 ;
  assign n16425 = n16423 & n16424 ;
  assign n16426 = ~n16420 & n16425 ;
  assign n16427 = ~n16417 & ~n16426 ;
  assign n16428 = n16026 & n16098 ;
  assign n16429 = ~n16165 & ~n16428 ;
  assign n16430 = \u0_w_reg[3][26]/P0001  & ~n16429 ;
  assign n16403 = n16105 & n16392 ;
  assign n16404 = ~n16064 & ~n16403 ;
  assign n16405 = ~\u0_w_reg[3][26]/P0001  & ~n16404 ;
  assign n16431 = ~\u0_w_reg[3][27]/P0001  & n16040 ;
  assign n16432 = ~n16405 & ~n16431 ;
  assign n16433 = ~n16430 & n16432 ;
  assign n16434 = ~n16427 & n16433 ;
  assign n16435 = ~\u0_w_reg[3][24]/P0001  & ~n16434 ;
  assign n16439 = ~\u0_w_reg[3][28]/P0001  & n16025 ;
  assign n16438 = \u0_w_reg[3][28]/P0001  & n16094 ;
  assign n16440 = ~n16150 & ~n16438 ;
  assign n16441 = ~n16439 & n16440 ;
  assign n16442 = n16386 & ~n16441 ;
  assign n16436 = \u0_w_reg[3][26]/P0001  & ~n16394 ;
  assign n16437 = n16032 & n16142 ;
  assign n16443 = n16094 & n16359 ;
  assign n16444 = n16117 & n16443 ;
  assign n16445 = ~n16437 & ~n16444 ;
  assign n16446 = ~n16436 & n16445 ;
  assign n16447 = ~n16442 & n16446 ;
  assign n16448 = \u0_w_reg[3][25]/P0001  & ~n16447 ;
  assign n16455 = ~n16053 & ~n16431 ;
  assign n16456 = ~\u0_w_reg[3][25]/P0001  & \u0_w_reg[3][26]/P0001  ;
  assign n16457 = ~n16455 & n16456 ;
  assign n16450 = \u0_w_reg[3][26]/P0001  & n16099 ;
  assign n16451 = n16098 & n16109 ;
  assign n16452 = ~n16450 & ~n16451 ;
  assign n16453 = n16032 & ~n16452 ;
  assign n16449 = n16169 & n16392 ;
  assign n16454 = \u0_w_reg[3][26]/P0001  & n16376 ;
  assign n16458 = ~n16449 & ~n16454 ;
  assign n16459 = ~n16453 & n16458 ;
  assign n16460 = ~n16457 & n16459 ;
  assign n16461 = ~n16448 & n16460 ;
  assign n16462 = ~n16435 & n16461 ;
  assign n16463 = ~n16402 & n16462 ;
  assign n16464 = \u0_w_reg[0][3]/P0001  & ~n16463 ;
  assign n16465 = ~\u0_w_reg[0][3]/P0001  & n16463 ;
  assign n16466 = ~n16464 & ~n16465 ;
  assign n16467 = \u0_w_reg[1][3]/P0001  & ~\u0_w_reg[2][3]/P0001  ;
  assign n16468 = ~\u0_w_reg[1][3]/P0001  & \u0_w_reg[2][3]/P0001  ;
  assign n16469 = ~n16467 & ~n16468 ;
  assign n16470 = n16466 & n16469 ;
  assign n16471 = ~n16466 & ~n16469 ;
  assign n16472 = ~n16470 & ~n16471 ;
  assign n16473 = ~ld_pad & n16472 ;
  assign n16474 = ~n16358 & ~n16473 ;
  assign n16475 = ~\key[43]_pad  & ld_pad ;
  assign n16480 = ~\u0_w_reg[3][5]/P0001  & ~\u0_w_reg[3][7]/P0001  ;
  assign n16481 = ~\u0_w_reg[3][4]/P0001  & n16480 ;
  assign n16482 = ~\u0_w_reg[3][3]/P0001  & \u0_w_reg[3][5]/P0001  ;
  assign n16483 = \u0_w_reg[3][6]/P0001  & ~\u0_w_reg[3][7]/P0001  ;
  assign n16484 = n16482 & n16483 ;
  assign n16485 = \u0_w_reg[3][4]/P0001  & n16484 ;
  assign n16486 = ~n16481 & ~n16485 ;
  assign n16487 = \u0_w_reg[3][2]/P0001  & ~n16486 ;
  assign n16476 = \u0_w_reg[3][5]/P0001  & \u0_w_reg[3][7]/P0001  ;
  assign n16477 = ~\u0_w_reg[3][4]/P0001  & \u0_w_reg[3][6]/P0001  ;
  assign n16478 = n16476 & n16477 ;
  assign n16479 = ~\u0_w_reg[3][3]/P0001  & n16478 ;
  assign n16492 = \u0_w_reg[3][3]/P0001  & \u0_w_reg[3][7]/P0001  ;
  assign n16493 = ~\u0_w_reg[3][5]/P0001  & ~\u0_w_reg[3][6]/P0001  ;
  assign n16494 = n16492 & n16493 ;
  assign n16498 = \u0_w_reg[3][1]/P0001  & ~n16494 ;
  assign n16499 = ~n16479 & n16498 ;
  assign n16488 = \u0_w_reg[3][5]/P0001  & ~\u0_w_reg[3][6]/P0001  ;
  assign n16489 = ~\u0_w_reg[3][4]/P0001  & \u0_w_reg[3][7]/P0001  ;
  assign n16490 = n16488 & n16489 ;
  assign n16491 = ~\u0_w_reg[3][2]/P0001  & n16490 ;
  assign n16495 = \u0_w_reg[3][5]/P0001  & \u0_w_reg[3][6]/P0001  ;
  assign n16496 = \u0_w_reg[3][4]/P0001  & n16492 ;
  assign n16497 = n16495 & n16496 ;
  assign n16500 = ~n16491 & ~n16497 ;
  assign n16501 = n16499 & n16500 ;
  assign n16502 = ~n16487 & n16501 ;
  assign n16503 = ~\u0_w_reg[3][5]/P0001  & n16489 ;
  assign n16504 = ~\u0_w_reg[3][3]/P0001  & n16503 ;
  assign n16515 = ~\u0_w_reg[3][1]/P0001  & ~n16504 ;
  assign n16512 = \u0_w_reg[3][2]/P0001  & ~\u0_w_reg[3][3]/P0001  ;
  assign n16513 = \u0_w_reg[3][7]/P0001  & ~n16493 ;
  assign n16514 = n16512 & n16513 ;
  assign n16505 = \u0_w_reg[3][4]/P0001  & ~\u0_w_reg[3][6]/P0001  ;
  assign n16506 = \u0_w_reg[3][2]/P0001  & ~\u0_w_reg[3][7]/P0001  ;
  assign n16507 = ~n16480 & ~n16506 ;
  assign n16508 = n16505 & ~n16507 ;
  assign n16509 = ~\u0_w_reg[3][2]/P0001  & \u0_w_reg[3][4]/P0001  ;
  assign n16510 = n16492 & n16509 ;
  assign n16511 = n16488 & n16510 ;
  assign n16516 = ~n16508 & ~n16511 ;
  assign n16517 = ~n16514 & n16516 ;
  assign n16518 = n16515 & n16517 ;
  assign n16519 = ~n16502 & ~n16518 ;
  assign n16528 = \u0_w_reg[3][4]/P0001  & \u0_w_reg[3][7]/P0001  ;
  assign n16529 = n16482 & n16528 ;
  assign n16530 = \u0_w_reg[3][6]/P0001  & n16529 ;
  assign n16531 = \u0_w_reg[3][3]/P0001  & ~\u0_w_reg[3][7]/P0001  ;
  assign n16532 = \u0_w_reg[3][4]/P0001  & n16531 ;
  assign n16533 = \u0_w_reg[3][6]/P0001  & n16532 ;
  assign n16534 = ~n16530 & ~n16533 ;
  assign n16535 = ~\u0_w_reg[3][2]/P0001  & ~n16534 ;
  assign n16520 = ~\u0_w_reg[3][3]/P0001  & ~\u0_w_reg[3][4]/P0001  ;
  assign n16521 = ~\u0_w_reg[3][5]/P0001  & \u0_w_reg[3][6]/P0001  ;
  assign n16522 = ~\u0_w_reg[3][7]/P0001  & n16521 ;
  assign n16523 = n16520 & n16522 ;
  assign n16536 = ~\u0_w_reg[3][0]/P0001  & ~n16523 ;
  assign n16524 = \u0_w_reg[3][2]/P0001  & \u0_w_reg[3][3]/P0001  ;
  assign n16525 = n16481 & n16524 ;
  assign n16526 = \u0_w_reg[3][2]/P0001  & n16476 ;
  assign n16527 = n16477 & n16526 ;
  assign n16537 = ~n16525 & ~n16527 ;
  assign n16538 = n16536 & n16537 ;
  assign n16539 = ~n16535 & n16538 ;
  assign n16540 = ~n16519 & n16539 ;
  assign n16574 = ~\u0_w_reg[3][5]/P0001  & \u0_w_reg[3][7]/P0001  ;
  assign n16582 = \u0_w_reg[3][4]/P0001  & n16574 ;
  assign n16583 = n16488 & ~n16531 ;
  assign n16584 = ~n16582 & ~n16583 ;
  assign n16585 = \u0_w_reg[3][2]/P0001  & ~n16584 ;
  assign n16544 = \u0_w_reg[3][3]/P0001  & \u0_w_reg[3][6]/P0001  ;
  assign n16580 = \u0_w_reg[3][4]/P0001  & ~n16544 ;
  assign n16581 = n16476 & n16580 ;
  assign n16590 = n16544 & n16574 ;
  assign n16586 = ~\u0_w_reg[3][2]/P0001  & ~\u0_w_reg[3][7]/P0001  ;
  assign n16587 = n16493 & n16586 ;
  assign n16588 = ~\u0_w_reg[3][2]/P0001  & ~\u0_w_reg[3][3]/P0001  ;
  assign n16589 = n16483 & n16588 ;
  assign n16591 = ~n16587 & ~n16589 ;
  assign n16592 = ~n16590 & n16591 ;
  assign n16593 = ~n16581 & n16592 ;
  assign n16594 = ~n16585 & n16593 ;
  assign n16595 = \u0_w_reg[3][1]/P0001  & ~n16594 ;
  assign n16541 = \u0_w_reg[3][6]/P0001  & \u0_w_reg[3][7]/P0001  ;
  assign n16542 = ~\u0_w_reg[3][5]/P0001  & n16541 ;
  assign n16543 = ~\u0_w_reg[3][3]/P0001  & n16542 ;
  assign n16545 = n16480 & n16544 ;
  assign n16546 = ~n16543 & ~n16545 ;
  assign n16547 = ~\u0_w_reg[3][2]/P0001  & ~n16546 ;
  assign n16554 = ~\u0_w_reg[3][2]/P0001  & ~\u0_w_reg[3][4]/P0001  ;
  assign n16555 = n16494 & ~n16554 ;
  assign n16548 = ~\u0_w_reg[3][6]/P0001  & ~\u0_w_reg[3][7]/P0001  ;
  assign n16549 = n16520 & n16548 ;
  assign n16550 = n16495 & n16506 ;
  assign n16557 = ~n16549 & ~n16550 ;
  assign n16551 = \u0_w_reg[3][5]/P0001  & ~\u0_w_reg[3][7]/P0001  ;
  assign n16552 = \u0_w_reg[3][2]/P0001  & ~\u0_w_reg[3][4]/P0001  ;
  assign n16553 = n16551 & n16552 ;
  assign n16556 = n16495 & n16520 ;
  assign n16558 = ~n16553 & ~n16556 ;
  assign n16559 = n16557 & n16558 ;
  assign n16560 = ~n16555 & n16559 ;
  assign n16561 = ~n16547 & n16560 ;
  assign n16562 = ~\u0_w_reg[3][1]/P0001  & ~n16561 ;
  assign n16563 = n16488 & n16528 ;
  assign n16564 = ~\u0_w_reg[3][3]/P0001  & n16563 ;
  assign n16565 = \u0_w_reg[3][3]/P0001  & n16476 ;
  assign n16566 = \u0_w_reg[3][6]/P0001  & n16565 ;
  assign n16567 = ~n16564 & ~n16566 ;
  assign n16568 = ~\u0_w_reg[3][2]/P0001  & ~n16504 ;
  assign n16569 = n16567 & n16568 ;
  assign n16573 = \u0_w_reg[3][4]/P0001  & n16522 ;
  assign n16575 = n16505 & n16574 ;
  assign n16570 = ~\u0_w_reg[3][6]/P0001  & \u0_w_reg[3][7]/P0001  ;
  assign n16571 = \u0_w_reg[3][3]/P0001  & \u0_w_reg[3][4]/P0001  ;
  assign n16572 = n16570 & n16571 ;
  assign n16576 = \u0_w_reg[3][2]/P0001  & ~n16572 ;
  assign n16577 = ~n16575 & n16576 ;
  assign n16578 = ~n16573 & n16577 ;
  assign n16579 = ~n16569 & ~n16578 ;
  assign n16596 = ~\u0_w_reg[3][4]/P0001  & n16551 ;
  assign n16597 = n16544 & n16596 ;
  assign n16598 = \u0_w_reg[3][0]/P0001  & ~n16597 ;
  assign n16599 = ~n16579 & n16598 ;
  assign n16600 = ~n16562 & n16599 ;
  assign n16601 = ~n16595 & n16600 ;
  assign n16602 = ~n16540 & ~n16601 ;
  assign n16608 = \u0_w_reg[3][4]/P0001  & n16493 ;
  assign n16607 = ~\u0_w_reg[3][4]/P0001  & n16483 ;
  assign n16609 = ~n16490 & ~n16607 ;
  assign n16610 = ~n16608 & n16609 ;
  assign n16611 = n16588 & ~n16610 ;
  assign n16612 = \u0_w_reg[3][3]/P0001  & ~\u0_w_reg[3][4]/P0001  ;
  assign n16613 = n16495 & n16612 ;
  assign n16614 = ~n16563 & ~n16613 ;
  assign n16615 = \u0_w_reg[3][2]/P0001  & ~n16614 ;
  assign n16606 = n16494 & n16554 ;
  assign n16616 = n16524 & n16542 ;
  assign n16617 = ~n16606 & ~n16616 ;
  assign n16618 = ~n16615 & n16617 ;
  assign n16619 = ~n16611 & n16618 ;
  assign n16620 = \u0_w_reg[3][1]/P0001  & ~n16619 ;
  assign n16621 = ~\u0_w_reg[3][1]/P0001  & \u0_w_reg[3][2]/P0001  ;
  assign n16622 = ~\u0_w_reg[3][3]/P0001  & n16548 ;
  assign n16623 = ~\u0_w_reg[3][5]/P0001  & n16622 ;
  assign n16624 = \u0_w_reg[3][4]/P0001  & n16623 ;
  assign n16625 = ~n16523 & ~n16624 ;
  assign n16626 = n16621 & ~n16625 ;
  assign n16630 = ~\u0_w_reg[3][5]/P0001  & n16532 ;
  assign n16631 = \u0_w_reg[3][6]/P0001  & n16630 ;
  assign n16603 = ~\u0_w_reg[3][1]/P0001  & ~\u0_w_reg[3][2]/P0001  ;
  assign n16604 = n16489 & n16544 ;
  assign n16605 = n16603 & n16604 ;
  assign n16627 = n16477 & n16574 ;
  assign n16628 = ~n16575 & ~n16627 ;
  assign n16629 = n16524 & ~n16628 ;
  assign n16632 = ~n16605 & ~n16629 ;
  assign n16633 = ~n16631 & n16632 ;
  assign n16634 = ~n16626 & n16633 ;
  assign n16635 = ~n16620 & n16634 ;
  assign n16636 = ~n16602 & n16635 ;
  assign n16637 = \u0_w_reg[0][11]/P0001  & ~n16636 ;
  assign n16638 = ~\u0_w_reg[0][11]/P0001  & n16636 ;
  assign n16639 = ~n16637 & ~n16638 ;
  assign n16640 = \u0_w_reg[1][11]/P0001  & ~\u0_w_reg[2][11]/P0001  ;
  assign n16641 = ~\u0_w_reg[1][11]/P0001  & \u0_w_reg[2][11]/P0001  ;
  assign n16642 = ~n16640 & ~n16641 ;
  assign n16643 = n16639 & n16642 ;
  assign n16644 = ~n16639 & ~n16642 ;
  assign n16645 = ~n16643 & ~n16644 ;
  assign n16646 = ~ld_pad & n16645 ;
  assign n16647 = ~n16475 & ~n16646 ;
  assign n16648 = ~\key[44]_pad  & ld_pad ;
  assign n16672 = ~n16575 & ~n16607 ;
  assign n16673 = ~\u0_w_reg[3][2]/P0001  & ~n16672 ;
  assign n16674 = n16552 & n16570 ;
  assign n16658 = ~\u0_w_reg[3][4]/P0001  & ~\u0_w_reg[3][7]/P0001  ;
  assign n16675 = \u0_w_reg[3][3]/P0001  & n16658 ;
  assign n16676 = n16488 & n16675 ;
  assign n16677 = ~n16674 & ~n16676 ;
  assign n16678 = ~n16624 & n16677 ;
  assign n16679 = ~n16673 & n16678 ;
  assign n16680 = \u0_w_reg[3][1]/P0001  & ~n16679 ;
  assign n16649 = ~\u0_w_reg[3][4]/P0001  & n16476 ;
  assign n16650 = n16548 & n16571 ;
  assign n16651 = ~n16649 & ~n16650 ;
  assign n16652 = ~\u0_w_reg[3][2]/P0001  & ~n16651 ;
  assign n16653 = ~\u0_w_reg[3][5]/P0001  & ~n16477 ;
  assign n16654 = n16492 & ~n16653 ;
  assign n16655 = ~n16652 & ~n16654 ;
  assign n16656 = ~\u0_w_reg[3][1]/P0001  & ~n16655 ;
  assign n16666 = ~\u0_w_reg[3][1]/P0001  & n16563 ;
  assign n16667 = ~\u0_w_reg[3][3]/P0001  & \u0_w_reg[3][4]/P0001  ;
  assign n16668 = ~\u0_w_reg[3][7]/P0001  & n16667 ;
  assign n16669 = ~n16494 & ~n16668 ;
  assign n16670 = ~n16666 & n16669 ;
  assign n16671 = \u0_w_reg[3][2]/P0001  & ~n16670 ;
  assign n16659 = n16493 & n16658 ;
  assign n16660 = ~\u0_w_reg[3][3]/P0001  & n16659 ;
  assign n16657 = n16483 & n16612 ;
  assign n16661 = ~n16590 & ~n16657 ;
  assign n16662 = ~n16660 & n16661 ;
  assign n16663 = ~\u0_w_reg[3][2]/P0001  & ~n16662 ;
  assign n16664 = ~\u0_w_reg[3][4]/P0001  & n16524 ;
  assign n16665 = ~\u0_w_reg[3][6]/P0001  & n16664 ;
  assign n16681 = \u0_w_reg[3][0]/P0001  & ~n16527 ;
  assign n16682 = ~n16665 & n16681 ;
  assign n16683 = ~n16663 & n16682 ;
  assign n16684 = ~n16671 & n16683 ;
  assign n16685 = ~n16656 & n16684 ;
  assign n16686 = ~n16680 & n16685 ;
  assign n16705 = n16489 & n16493 ;
  assign n16706 = \u0_w_reg[3][5]/P0001  & n16570 ;
  assign n16707 = ~n16612 & n16706 ;
  assign n16708 = ~n16705 & ~n16707 ;
  assign n16709 = ~\u0_w_reg[3][2]/P0001  & ~n16708 ;
  assign n16710 = n16512 & n16582 ;
  assign n16711 = ~n16533 & ~n16550 ;
  assign n16712 = ~n16710 & n16711 ;
  assign n16713 = ~n16709 & n16712 ;
  assign n16714 = \u0_w_reg[3][1]/P0001  & ~n16713 ;
  assign n16692 = \u0_w_reg[3][5]/P0001  & n16589 ;
  assign n16687 = \u0_w_reg[3][4]/P0001  & n16495 ;
  assign n16688 = \u0_w_reg[3][2]/P0001  & n16687 ;
  assign n16689 = \u0_w_reg[3][2]/P0001  & ~\u0_w_reg[3][5]/P0001  ;
  assign n16690 = ~n16612 & ~n16689 ;
  assign n16691 = n16548 & ~n16690 ;
  assign n16693 = ~n16688 & ~n16691 ;
  assign n16694 = ~n16692 & n16693 ;
  assign n16695 = ~\u0_w_reg[3][1]/P0001  & ~n16694 ;
  assign n16696 = n16509 & n16542 ;
  assign n16697 = n16488 & n16658 ;
  assign n16698 = ~n16696 & ~n16697 ;
  assign n16699 = ~\u0_w_reg[3][3]/P0001  & ~n16698 ;
  assign n16700 = ~\u0_w_reg[3][4]/P0001  & n16521 ;
  assign n16701 = n16493 & n16531 ;
  assign n16702 = ~n16700 & ~n16701 ;
  assign n16703 = \u0_w_reg[3][2]/P0001  & ~n16612 ;
  assign n16704 = ~n16702 & n16703 ;
  assign n16715 = ~\u0_w_reg[3][0]/P0001  & ~n16704 ;
  assign n16716 = ~n16699 & n16715 ;
  assign n16717 = ~n16695 & n16716 ;
  assign n16718 = ~n16714 & n16717 ;
  assign n16719 = ~n16686 & ~n16718 ;
  assign n16720 = n16522 & n16554 ;
  assign n16721 = ~n16688 & ~n16720 ;
  assign n16722 = \u0_w_reg[3][3]/P0001  & ~n16721 ;
  assign n16723 = n16544 & n16649 ;
  assign n16724 = ~\u0_w_reg[3][2]/P0001  & ~n16723 ;
  assign n16725 = ~\u0_w_reg[3][3]/P0001  & n16521 ;
  assign n16726 = ~n16658 & n16725 ;
  assign n16727 = n16724 & ~n16726 ;
  assign n16730 = ~\u0_w_reg[3][3]/P0001  & n16705 ;
  assign n16731 = \u0_w_reg[3][2]/P0001  & ~n16730 ;
  assign n16732 = n16492 & n16608 ;
  assign n16728 = n16544 & n16551 ;
  assign n16729 = n16488 & n16612 ;
  assign n16733 = ~n16728 & ~n16729 ;
  assign n16734 = ~n16732 & n16733 ;
  assign n16735 = n16731 & n16734 ;
  assign n16736 = ~n16727 & ~n16735 ;
  assign n16738 = n16482 & ~n16509 ;
  assign n16739 = n16548 & n16738 ;
  assign n16737 = n16495 & n16532 ;
  assign n16740 = ~\u0_w_reg[3][1]/P0001  & ~n16737 ;
  assign n16741 = ~n16739 & n16740 ;
  assign n16742 = ~n16736 & n16741 ;
  assign n16748 = \u0_w_reg[3][3]/P0001  & ~n16548 ;
  assign n16749 = ~n16549 & ~n16748 ;
  assign n16750 = ~\u0_w_reg[3][5]/P0001  & ~n16749 ;
  assign n16751 = ~n16479 & ~n16750 ;
  assign n16752 = ~\u0_w_reg[3][2]/P0001  & ~n16751 ;
  assign n16745 = n16483 & n16512 ;
  assign n16746 = ~n16590 & ~n16745 ;
  assign n16747 = \u0_w_reg[3][4]/P0001  & ~n16746 ;
  assign n16753 = \u0_w_reg[3][5]/P0001  & n16548 ;
  assign n16754 = n16524 & n16753 ;
  assign n16743 = ~\u0_w_reg[3][5]/P0001  & n16612 ;
  assign n16744 = n16570 & n16743 ;
  assign n16755 = \u0_w_reg[3][1]/P0001  & ~n16744 ;
  assign n16756 = ~n16754 & n16755 ;
  assign n16757 = ~n16747 & n16756 ;
  assign n16758 = ~n16752 & n16757 ;
  assign n16759 = ~n16742 & ~n16758 ;
  assign n16760 = ~n16722 & ~n16759 ;
  assign n16761 = ~n16719 & n16760 ;
  assign n16762 = \u0_w_reg[0][12]/P0001  & ~n16761 ;
  assign n16763 = ~\u0_w_reg[0][12]/P0001  & n16761 ;
  assign n16764 = ~n16762 & ~n16763 ;
  assign n16765 = \u0_w_reg[1][12]/P0001  & ~\u0_w_reg[2][12]/P0001  ;
  assign n16766 = ~\u0_w_reg[1][12]/P0001  & \u0_w_reg[2][12]/P0001  ;
  assign n16767 = ~n16765 & ~n16766 ;
  assign n16768 = n16764 & n16767 ;
  assign n16769 = ~n16764 & ~n16767 ;
  assign n16770 = ~n16768 & ~n16769 ;
  assign n16771 = ~ld_pad & n16770 ;
  assign n16772 = ~n16648 & ~n16771 ;
  assign n16773 = \key[120]_pad  & ld_pad ;
  assign n16818 = ~n15543 & ~n15600 ;
  assign n16819 = ~\u0_w_reg[3][19]/P0001  & ~n16818 ;
  assign n16820 = n15530 & n15660 ;
  assign n16821 = \u0_w_reg[3][20]/P0001  & n16820 ;
  assign n16816 = ~n15545 & ~n15585 ;
  assign n16817 = \u0_w_reg[3][18]/P0001  & ~n16816 ;
  assign n16822 = ~\u0_w_reg[3][17]/P0001  & ~n15556 ;
  assign n16823 = ~n15662 & n16822 ;
  assign n16824 = ~n16817 & n16823 ;
  assign n16825 = ~n16821 & n16824 ;
  assign n16826 = ~n16819 & n16825 ;
  assign n16827 = ~\u0_w_reg[3][18]/P0001  & n15512 ;
  assign n16828 = \u0_w_reg[3][17]/P0001  & ~n15618 ;
  assign n16829 = ~n16827 & n16828 ;
  assign n16830 = ~n16232 & n16829 ;
  assign n16831 = ~n16826 & ~n16830 ;
  assign n16802 = ~\u0_w_reg[3][20]/P0001  & n15587 ;
  assign n16803 = ~n15563 & ~n16802 ;
  assign n16804 = \u0_w_reg[3][18]/P0001  & ~n16269 ;
  assign n16805 = ~n15561 & n16804 ;
  assign n16806 = n16803 & n16805 ;
  assign n16808 = ~n15518 & ~n15613 ;
  assign n16809 = \u0_w_reg[3][19]/P0001  & ~n16808 ;
  assign n16807 = n15525 & n15542 ;
  assign n16810 = ~\u0_w_reg[3][18]/P0001  & ~n16807 ;
  assign n16811 = ~n15514 & n16810 ;
  assign n16812 = ~n16809 & n16811 ;
  assign n16813 = ~n16806 & ~n16812 ;
  assign n16814 = ~\u0_w_reg[3][19]/P0001  & n15516 ;
  assign n16815 = n15530 & n15662 ;
  assign n16832 = ~n16814 & ~n16815 ;
  assign n16833 = ~n16813 & n16832 ;
  assign n16834 = ~n16831 & n16833 ;
  assign n16835 = \u0_w_reg[3][16]/P0001  & ~n16834 ;
  assign n16779 = \u0_w_reg[3][20]/P0001  & n16229 ;
  assign n16780 = ~n15660 & ~n16779 ;
  assign n16781 = \u0_w_reg[3][23]/P0001  & ~n16780 ;
  assign n16777 = \u0_w_reg[3][18]/P0001  & n15516 ;
  assign n16778 = \u0_w_reg[3][19]/P0001  & n16777 ;
  assign n16782 = n15520 & ~n15521 ;
  assign n16783 = \u0_w_reg[3][17]/P0001  & ~n16782 ;
  assign n16784 = ~n16778 & n16783 ;
  assign n16785 = ~n16781 & n16784 ;
  assign n16786 = ~n16283 & ~n16313 ;
  assign n16787 = ~\u0_w_reg[3][19]/P0001  & ~n16786 ;
  assign n16788 = n15526 & ~n16229 ;
  assign n16789 = \u0_w_reg[3][18]/P0001  & ~n16788 ;
  assign n16790 = ~\u0_w_reg[3][18]/P0001  & ~n15522 ;
  assign n16791 = ~n16789 & ~n16790 ;
  assign n16792 = ~\u0_w_reg[3][17]/P0001  & ~n16791 ;
  assign n16793 = ~n16787 & n16792 ;
  assign n16794 = ~n16785 & ~n16793 ;
  assign n16774 = \u0_w_reg[3][21]/P0001  & n15520 ;
  assign n16775 = ~n15518 & ~n16774 ;
  assign n16776 = n16266 & ~n16775 ;
  assign n16795 = n15506 & n15549 ;
  assign n16796 = ~n16242 & ~n16795 ;
  assign n16797 = ~n15561 & n16796 ;
  assign n16798 = ~\u0_w_reg[3][18]/P0001  & ~n16797 ;
  assign n16799 = ~n16776 & ~n16798 ;
  assign n16800 = ~n16794 & n16799 ;
  assign n16801 = ~\u0_w_reg[3][16]/P0001  & ~n16800 ;
  assign n16836 = n15529 & n15544 ;
  assign n16837 = n15507 & n15542 ;
  assign n16838 = ~n16836 & ~n16837 ;
  assign n16839 = \u0_w_reg[3][22]/P0001  & ~n16838 ;
  assign n16840 = \u0_w_reg[3][20]/P0001  & n15518 ;
  assign n16841 = n15511 & n16840 ;
  assign n16842 = ~n15657 & ~n16795 ;
  assign n16843 = ~n16841 & n16842 ;
  assign n16844 = ~\u0_w_reg[3][23]/P0001  & ~n16843 ;
  assign n16845 = n15531 & n15608 ;
  assign n16846 = \u0_w_reg[3][17]/P0001  & ~n16239 ;
  assign n16847 = ~n16845 & n16846 ;
  assign n16848 = ~n16844 & n16847 ;
  assign n16854 = \u0_w_reg[3][20]/P0001  & n15503 ;
  assign n16853 = n15559 & n15613 ;
  assign n16855 = ~n15638 & ~n16853 ;
  assign n16856 = ~n16854 & n16855 ;
  assign n16857 = n15648 & ~n16856 ;
  assign n16849 = ~n15512 & ~n15531 ;
  assign n16850 = n15507 & ~n16849 ;
  assign n16851 = n15512 & n15613 ;
  assign n16852 = n15529 & n16851 ;
  assign n16858 = ~\u0_w_reg[3][17]/P0001  & ~n15656 ;
  assign n16859 = ~n16852 & n16858 ;
  assign n16860 = ~n16850 & n16859 ;
  assign n16861 = ~n16857 & n16860 ;
  assign n16862 = ~n16848 & ~n16861 ;
  assign n16863 = ~n16839 & ~n16862 ;
  assign n16864 = ~n16801 & n16863 ;
  assign n16865 = ~n16835 & n16864 ;
  assign n16866 = \u0_r0_out_reg[24]/P0001  & ~\u0_w_reg[0][24]/P0001  ;
  assign n16867 = ~\u0_r0_out_reg[24]/P0001  & \u0_w_reg[0][24]/P0001  ;
  assign n16868 = ~n16866 & ~n16867 ;
  assign n16869 = ~n16865 & ~n16868 ;
  assign n16870 = n16865 & n16868 ;
  assign n16871 = ~n16869 & ~n16870 ;
  assign n16872 = ~ld_pad & n16871 ;
  assign n16873 = ~n16773 & ~n16872 ;
  assign n16913 = ~\u0_w_reg[3][21]/P0001  & ~n15588 ;
  assign n16914 = n15520 & ~n16913 ;
  assign n16915 = ~n15543 & ~n16914 ;
  assign n16916 = ~\u0_w_reg[3][19]/P0001  & ~n16915 ;
  assign n16917 = n15503 & n15511 ;
  assign n16920 = ~\u0_w_reg[3][17]/P0001  & ~n16917 ;
  assign n16918 = n16268 & n16297 ;
  assign n16919 = n15504 & n15590 ;
  assign n16921 = ~n16918 & ~n16919 ;
  assign n16922 = n16920 & n16921 ;
  assign n16923 = ~n15647 & ~n16777 ;
  assign n16924 = n16922 & n16923 ;
  assign n16925 = ~n16916 & n16924 ;
  assign n16926 = n15613 & n16297 ;
  assign n16927 = \u0_w_reg[3][17]/P0001  & ~n16926 ;
  assign n16928 = ~n16852 & n16927 ;
  assign n16929 = ~n16925 & ~n16928 ;
  assign n16904 = ~n15606 & ~n15618 ;
  assign n16905 = ~n15655 & n16904 ;
  assign n16906 = n15608 & ~n16905 ;
  assign n16910 = \u0_w_reg[3][17]/P0001  & ~\u0_w_reg[3][18]/P0001  ;
  assign n16911 = ~n16261 & ~n16309 ;
  assign n16912 = n16910 & ~n16911 ;
  assign n16907 = ~n15531 & ~n16774 ;
  assign n16908 = n15506 & ~n16907 ;
  assign n16909 = n15511 & n15516 ;
  assign n16930 = \u0_w_reg[3][16]/P0001  & ~n16909 ;
  assign n16931 = ~n16908 & n16930 ;
  assign n16932 = ~n16912 & n16931 ;
  assign n16933 = ~n16906 & n16932 ;
  assign n16934 = ~n16929 & n16933 ;
  assign n16935 = n15529 & n15542 ;
  assign n16936 = ~\u0_w_reg[3][17]/P0001  & ~n15527 ;
  assign n16937 = ~n16935 & n16936 ;
  assign n16944 = \u0_w_reg[3][21]/P0001  & n15575 ;
  assign n16945 = \u0_w_reg[3][17]/P0001  & ~n16944 ;
  assign n16938 = ~n15613 & ~n16229 ;
  assign n16939 = ~\u0_w_reg[3][18]/P0001  & ~n15542 ;
  assign n16940 = ~n16938 & n16939 ;
  assign n16941 = ~\u0_w_reg[3][19]/P0001  & n15520 ;
  assign n16942 = ~n15540 & ~n16941 ;
  assign n16943 = \u0_w_reg[3][18]/P0001  & ~n16942 ;
  assign n16946 = ~n16940 & ~n16943 ;
  assign n16947 = n16945 & n16946 ;
  assign n16948 = ~n16937 & ~n16947 ;
  assign n16949 = n15602 & n15608 ;
  assign n16950 = \u0_w_reg[3][22]/P0001  & n16949 ;
  assign n16951 = ~\u0_w_reg[3][16]/P0001  & ~n15628 ;
  assign n16952 = ~n15659 & n16951 ;
  assign n16953 = ~n16950 & n16952 ;
  assign n16954 = ~n16948 & n16953 ;
  assign n16955 = ~n16934 & ~n16954 ;
  assign n16887 = ~n15650 & ~n16853 ;
  assign n16888 = ~n16249 & n16887 ;
  assign n16889 = ~\u0_w_reg[3][18]/P0001  & ~n16888 ;
  assign n16881 = ~n15549 & ~n16313 ;
  assign n16882 = n15608 & ~n16881 ;
  assign n16886 = \u0_w_reg[3][18]/P0001  & n15527 ;
  assign n16883 = ~n15525 & n15549 ;
  assign n16884 = ~n15613 & n16883 ;
  assign n16885 = n15648 & n16774 ;
  assign n16890 = ~n16884 & ~n16885 ;
  assign n16891 = ~n16886 & n16890 ;
  assign n16892 = ~n16882 & n16891 ;
  assign n16893 = ~n16889 & n16892 ;
  assign n16894 = ~\u0_w_reg[3][17]/P0001  & ~n16893 ;
  assign n16874 = ~n15625 & ~n16289 ;
  assign n16875 = ~\u0_w_reg[3][19]/P0001  & n15530 ;
  assign n16876 = \u0_w_reg[3][20]/P0001  & n16875 ;
  assign n16877 = n16874 & ~n16876 ;
  assign n16878 = ~\u0_w_reg[3][18]/P0001  & ~n16877 ;
  assign n16879 = ~n15592 & ~n16878 ;
  assign n16880 = \u0_w_reg[3][17]/P0001  & ~n16879 ;
  assign n16895 = n15518 & n16266 ;
  assign n16896 = \u0_w_reg[3][17]/P0001  & ~\u0_w_reg[3][23]/P0001  ;
  assign n16897 = n16895 & n16896 ;
  assign n16956 = ~n16270 & ~n16897 ;
  assign n16898 = ~n15601 & ~n16774 ;
  assign n16899 = n15507 & ~n16898 ;
  assign n16900 = ~n15506 & ~n16840 ;
  assign n16901 = \u0_w_reg[3][17]/P0001  & \u0_w_reg[3][18]/P0001  ;
  assign n16902 = \u0_w_reg[3][23]/P0001  & n16901 ;
  assign n16903 = ~n16900 & n16902 ;
  assign n16957 = ~n16899 & ~n16903 ;
  assign n16958 = n16956 & n16957 ;
  assign n16959 = ~n16880 & n16958 ;
  assign n16960 = ~n16894 & n16959 ;
  assign n16961 = ~n16955 & n16960 ;
  assign n16962 = \u0_w_reg[0][26]/P0001  & ~n16961 ;
  assign n16963 = ~\u0_w_reg[0][26]/P0001  & n16961 ;
  assign n16964 = ~n16962 & ~n16963 ;
  assign n16966 = \u0_r0_out_reg[26]/P0001  & n16964 ;
  assign n16965 = ~\u0_r0_out_reg[26]/P0001  & ~n16964 ;
  assign n16967 = ~ld_pad & ~n16965 ;
  assign n16968 = ~n16966 & n16967 ;
  assign n16969 = \key[122]_pad  & ld_pad ;
  assign n16970 = ~n16968 & ~n16969 ;
  assign n16972 = ~\u0_w_reg[3][20]/P0001  & n15592 ;
  assign n16973 = ~n15583 & ~n16854 ;
  assign n16974 = ~n16972 & n16973 ;
  assign n16975 = \u0_w_reg[3][18]/P0001  & ~n16974 ;
  assign n16971 = ~n15539 & n15660 ;
  assign n16976 = n16803 & ~n16971 ;
  assign n16977 = ~n16975 & n16976 ;
  assign n16978 = \u0_w_reg[3][17]/P0001  & ~n16977 ;
  assign n16984 = ~n15638 & ~n16248 ;
  assign n16985 = \u0_w_reg[3][18]/P0001  & ~n16984 ;
  assign n16986 = ~n15628 & ~n16885 ;
  assign n16987 = ~n16985 & n16986 ;
  assign n16988 = ~n15627 & n16987 ;
  assign n16989 = ~\u0_w_reg[3][17]/P0001  & ~n16988 ;
  assign n16979 = ~n15576 & ~n16851 ;
  assign n16980 = ~\u0_w_reg[3][18]/P0001  & ~n16979 ;
  assign n16981 = ~n15630 & ~n16217 ;
  assign n16982 = n16306 & n16981 ;
  assign n16983 = \u0_w_reg[3][18]/P0001  & ~n16982 ;
  assign n16990 = ~n16980 & ~n16983 ;
  assign n16991 = ~n16989 & n16990 ;
  assign n16992 = ~n16978 & n16991 ;
  assign n16993 = \u0_w_reg[3][16]/P0001  & ~n16992 ;
  assign n16996 = ~n16230 & ~n16310 ;
  assign n16994 = ~\u0_w_reg[3][19]/P0001  & n16261 ;
  assign n16995 = ~n15520 & n15662 ;
  assign n16997 = ~n16994 & ~n16995 ;
  assign n16998 = n16996 & n16997 ;
  assign n16999 = ~\u0_w_reg[3][18]/P0001  & ~n16998 ;
  assign n17001 = ~n15504 & ~n16309 ;
  assign n17002 = n15601 & ~n17001 ;
  assign n17004 = ~\u0_w_reg[3][17]/P0001  & ~n16836 ;
  assign n17005 = ~n16851 & n17004 ;
  assign n17000 = ~\u0_w_reg[3][20]/P0001  & n16875 ;
  assign n17003 = n15608 & n16774 ;
  assign n17006 = ~n17000 & ~n17003 ;
  assign n17007 = n17005 & n17006 ;
  assign n17008 = ~n17002 & n17007 ;
  assign n17009 = n15511 & ~n15616 ;
  assign n17010 = ~\u0_w_reg[3][18]/P0001  & n15630 ;
  assign n17011 = \u0_w_reg[3][17]/P0001  & ~n15650 ;
  assign n17012 = ~n17010 & n17011 ;
  assign n17013 = ~n17009 & n17012 ;
  assign n17014 = ~n17008 & ~n17013 ;
  assign n17015 = ~n16999 & ~n17014 ;
  assign n17016 = ~\u0_w_reg[3][16]/P0001  & ~n17015 ;
  assign n17020 = \u0_w_reg[3][21]/P0001  & n15530 ;
  assign n17035 = n15504 & n17020 ;
  assign n17036 = ~n15637 & ~n16284 ;
  assign n17037 = ~n17035 & n17036 ;
  assign n17038 = \u0_w_reg[3][17]/P0001  & ~n17037 ;
  assign n17032 = n15525 & n15591 ;
  assign n17033 = ~n16795 & ~n17032 ;
  assign n17034 = ~\u0_w_reg[3][16]/P0001  & ~n17033 ;
  assign n17039 = ~n16288 & ~n17034 ;
  assign n17040 = ~n17038 & n17039 ;
  assign n17041 = \u0_w_reg[3][18]/P0001  & ~n17040 ;
  assign n17021 = n15529 & n17020 ;
  assign n17018 = ~\u0_w_reg[3][18]/P0001  & n15618 ;
  assign n17019 = \u0_w_reg[3][18]/P0001  & n16313 ;
  assign n17024 = ~n17018 & ~n17019 ;
  assign n17025 = ~n17021 & n17024 ;
  assign n17022 = ~n15580 & ~n15629 ;
  assign n17017 = n15520 & n16266 ;
  assign n17023 = ~n16249 & ~n17017 ;
  assign n17026 = n17022 & n17023 ;
  assign n17027 = n17025 & n17026 ;
  assign n17028 = ~\u0_w_reg[3][17]/P0001  & ~n17027 ;
  assign n17030 = ~n15600 & ~n15630 ;
  assign n17031 = ~\u0_w_reg[3][19]/P0001  & ~n17030 ;
  assign n17029 = \u0_w_reg[3][17]/P0001  & n15659 ;
  assign n17042 = ~n16300 & ~n17029 ;
  assign n17043 = ~n17031 & n17042 ;
  assign n17044 = ~n17028 & n17043 ;
  assign n17045 = ~n17041 & n17044 ;
  assign n17046 = ~n17016 & n17045 ;
  assign n17047 = ~n16993 & n17046 ;
  assign n17048 = \u0_r0_out_reg[30]/P0001  & ~n17047 ;
  assign n17049 = ~\u0_r0_out_reg[30]/P0001  & n17047 ;
  assign n17050 = ~n17048 & ~n17049 ;
  assign n17052 = \u0_w_reg[0][30]/P0001  & n17050 ;
  assign n17051 = ~\u0_w_reg[0][30]/P0001  & ~n17050 ;
  assign n17053 = ~ld_pad & ~n17051 ;
  assign n17054 = ~n17052 & n17053 ;
  assign n17055 = \key[126]_pad  & ld_pad ;
  assign n17056 = ~n17054 & ~n17055 ;
  assign n17089 = \u0_w_reg[3][20]/P0001  & n15559 ;
  assign n17090 = \u0_w_reg[3][23]/P0001  & n15539 ;
  assign n17091 = ~n17089 & ~n17090 ;
  assign n17092 = n15511 & ~n17091 ;
  assign n17093 = ~n15586 & ~n16807 ;
  assign n17088 = \u0_w_reg[3][20]/P0001  & n16233 ;
  assign n17094 = ~n16895 & ~n17088 ;
  assign n17095 = n17093 & n17094 ;
  assign n17096 = ~n17092 & n17095 ;
  assign n17102 = ~n15513 & ~n16261 ;
  assign n17103 = ~n16854 & n17102 ;
  assign n17104 = ~\u0_w_reg[3][18]/P0001  & ~n17103 ;
  assign n17097 = ~n15525 & ~n15648 ;
  assign n17098 = \u0_w_reg[3][22]/P0001  & ~n17097 ;
  assign n17099 = ~n16827 & ~n17098 ;
  assign n17100 = ~\u0_w_reg[3][23]/P0001  & ~n17099 ;
  assign n17101 = \u0_w_reg[3][23]/P0001  & n15508 ;
  assign n17105 = ~n15657 & ~n17101 ;
  assign n17106 = ~n17100 & n17105 ;
  assign n17107 = ~n17104 & n17106 ;
  assign n17108 = n17096 & n17107 ;
  assign n17109 = \u0_w_reg[3][16]/P0001  & ~n17108 ;
  assign n17057 = ~n15543 & ~n15606 ;
  assign n17058 = n15648 & ~n17057 ;
  assign n17110 = ~\u0_w_reg[3][20]/P0001  & n15601 ;
  assign n17111 = n15529 & n17110 ;
  assign n17112 = n16936 & ~n17111 ;
  assign n17113 = ~n17058 & n17112 ;
  assign n17114 = ~n17109 & n17113 ;
  assign n17124 = n15559 & ~n16268 ;
  assign n17125 = n16786 & ~n17124 ;
  assign n17126 = \u0_w_reg[3][19]/P0001  & ~n17125 ;
  assign n17127 = ~\u0_w_reg[3][18]/P0001  & ~n17126 ;
  assign n17115 = ~n15539 & ~n16261 ;
  assign n17128 = \u0_w_reg[3][23]/P0001  & ~n17115 ;
  assign n17129 = ~n16853 & ~n17128 ;
  assign n17130 = ~\u0_w_reg[3][19]/P0001  & ~n17129 ;
  assign n17131 = \u0_w_reg[3][18]/P0001  & ~n15538 ;
  assign n17132 = ~n15625 & n17131 ;
  assign n17133 = ~n17130 & n17132 ;
  assign n17134 = ~n17127 & ~n17133 ;
  assign n17116 = \u0_w_reg[3][19]/P0001  & n15503 ;
  assign n17117 = ~n16941 & ~n17116 ;
  assign n17118 = n17115 & n17117 ;
  assign n17119 = \u0_w_reg[3][18]/P0001  & ~n17118 ;
  assign n17083 = n15518 & n16248 ;
  assign n17120 = ~n16820 & ~n17083 ;
  assign n17121 = ~n17119 & n17120 ;
  assign n17122 = n17096 & n17121 ;
  assign n17123 = \u0_w_reg[3][16]/P0001  & ~n17122 ;
  assign n17135 = \u0_w_reg[3][17]/P0001  & ~n17123 ;
  assign n17136 = ~n17134 & n17135 ;
  assign n17137 = ~n17114 & ~n17136 ;
  assign n17059 = n15518 & n15537 ;
  assign n17060 = ~n15562 & ~n17059 ;
  assign n17061 = ~\u0_w_reg[3][18]/P0001  & ~n17060 ;
  assign n17062 = ~n16841 & ~n17032 ;
  assign n17063 = n16945 & n17062 ;
  assign n17064 = ~n17061 & n17063 ;
  assign n17065 = ~\u0_w_reg[3][17]/P0001  & ~n15600 ;
  assign n17066 = ~n16802 & ~n16949 ;
  assign n17067 = n17065 & n17066 ;
  assign n17068 = ~n17064 & ~n17067 ;
  assign n17069 = ~n15663 & ~n16289 ;
  assign n17070 = \u0_w_reg[3][18]/P0001  & ~n17069 ;
  assign n17074 = ~n15651 & ~n15656 ;
  assign n17071 = ~\u0_w_reg[3][17]/P0001  & n16268 ;
  assign n17072 = ~n16284 & ~n17071 ;
  assign n17073 = ~\u0_w_reg[3][18]/P0001  & ~n17072 ;
  assign n17075 = ~n17058 & ~n17073 ;
  assign n17076 = n17074 & n17075 ;
  assign n17077 = ~n17070 & n17076 ;
  assign n17078 = ~n17068 & n17077 ;
  assign n17079 = ~\u0_w_reg[3][16]/P0001  & ~n17078 ;
  assign n17080 = ~\u0_w_reg[3][21]/P0001  & n15522 ;
  assign n17081 = ~n15581 & ~n17080 ;
  assign n17082 = ~\u0_w_reg[3][18]/P0001  & ~n17081 ;
  assign n17084 = \u0_w_reg[3][21]/P0001  & n16309 ;
  assign n17085 = ~n15584 & ~n17083 ;
  assign n17086 = ~n17084 & n17085 ;
  assign n17087 = n16281 & ~n17086 ;
  assign n17138 = ~n17082 & ~n17087 ;
  assign n17139 = ~n17079 & n17138 ;
  assign n17140 = ~n17137 & n17139 ;
  assign n17141 = \u0_w_reg[0][31]/P0001  & ~n17140 ;
  assign n17142 = ~\u0_w_reg[0][31]/P0001  & n17140 ;
  assign n17143 = ~n17141 & ~n17142 ;
  assign n17145 = \u0_r0_out_reg[31]/P0001  & n17143 ;
  assign n17144 = ~\u0_r0_out_reg[31]/P0001  & ~n17143 ;
  assign n17146 = ~ld_pad & ~n17144 ;
  assign n17147 = ~n17145 & n17146 ;
  assign n17148 = \key[127]_pad  & ld_pad ;
  assign n17149 = ~n17147 & ~n17148 ;
  assign n17150 = \u0_r0_out_reg[26]/P0001  & ~\u0_w_reg[1][26]/P0001  ;
  assign n17151 = ~\u0_r0_out_reg[26]/P0001  & \u0_w_reg[1][26]/P0001  ;
  assign n17152 = ~n17150 & ~n17151 ;
  assign n17154 = n16964 & ~n17152 ;
  assign n17153 = ~n16964 & n17152 ;
  assign n17155 = ~ld_pad & ~n17153 ;
  assign n17156 = ~n17154 & n17155 ;
  assign n17157 = \key[90]_pad  & ld_pad ;
  assign n17158 = ~n17156 & ~n17157 ;
  assign n17159 = \u0_w_reg[0][30]/P0001  & ~\u0_w_reg[1][30]/P0001  ;
  assign n17160 = ~\u0_w_reg[0][30]/P0001  & \u0_w_reg[1][30]/P0001  ;
  assign n17161 = ~n17159 & ~n17160 ;
  assign n17163 = n17050 & ~n17161 ;
  assign n17162 = ~n17050 & n17161 ;
  assign n17164 = ~ld_pad & ~n17162 ;
  assign n17165 = ~n17163 & n17164 ;
  assign n17166 = \key[94]_pad  & ld_pad ;
  assign n17167 = ~n17165 & ~n17166 ;
  assign n17168 = \u0_r0_out_reg[31]/P0001  & ~\u0_w_reg[1][31]/P0001  ;
  assign n17169 = ~\u0_r0_out_reg[31]/P0001  & \u0_w_reg[1][31]/P0001  ;
  assign n17170 = ~n17168 & ~n17169 ;
  assign n17172 = n17143 & ~n17170 ;
  assign n17171 = ~n17143 & n17170 ;
  assign n17173 = ~ld_pad & ~n17171 ;
  assign n17174 = ~n17172 & n17173 ;
  assign n17175 = \key[95]_pad  & ld_pad ;
  assign n17176 = ~n17174 & ~n17175 ;
  assign n17177 = \key[56]_pad  & ld_pad ;
  assign n17178 = \u0_w_reg[1][24]/P0002  & ~\u0_w_reg[2][24]/P0001  ;
  assign n17179 = ~\u0_w_reg[1][24]/P0002  & \u0_w_reg[2][24]/P0001  ;
  assign n17180 = ~n17178 & ~n17179 ;
  assign n17181 = ~n16868 & n17180 ;
  assign n17182 = n16868 & ~n17180 ;
  assign n17183 = ~n17181 & ~n17182 ;
  assign n17185 = ~n16865 & ~n17183 ;
  assign n17184 = n16865 & n17183 ;
  assign n17186 = ~ld_pad & ~n17184 ;
  assign n17187 = ~n17185 & n17186 ;
  assign n17188 = ~n17177 & ~n17187 ;
  assign n17189 = ~\key[58]_pad  & ld_pad ;
  assign n17190 = \u0_w_reg[2][26]/P0001  & n17152 ;
  assign n17191 = ~\u0_w_reg[2][26]/P0001  & ~n17152 ;
  assign n17192 = ~n17190 & ~n17191 ;
  assign n17193 = n16964 & n17192 ;
  assign n17194 = ~n16964 & ~n17192 ;
  assign n17195 = ~n17193 & ~n17194 ;
  assign n17196 = ~ld_pad & n17195 ;
  assign n17197 = ~n17189 & ~n17196 ;
  assign n17198 = ~\key[62]_pad  & ld_pad ;
  assign n17199 = \u0_w_reg[2][30]/P0001  & n17161 ;
  assign n17200 = ~\u0_w_reg[2][30]/P0001  & ~n17161 ;
  assign n17201 = ~n17199 & ~n17200 ;
  assign n17202 = n17050 & n17201 ;
  assign n17203 = ~n17050 & ~n17201 ;
  assign n17204 = ~n17202 & ~n17203 ;
  assign n17205 = ~ld_pad & n17204 ;
  assign n17206 = ~n17198 & ~n17205 ;
  assign n17207 = ~\key[63]_pad  & ld_pad ;
  assign n17208 = \u0_w_reg[2][31]/P0001  & n17170 ;
  assign n17209 = ~\u0_w_reg[2][31]/P0001  & ~n17170 ;
  assign n17210 = ~n17208 & ~n17209 ;
  assign n17211 = n17143 & n17210 ;
  assign n17212 = ~n17143 & ~n17210 ;
  assign n17213 = ~n17211 & ~n17212 ;
  assign n17214 = ~ld_pad & n17213 ;
  assign n17215 = ~n17207 & ~n17214 ;
  assign n17216 = \key[24]_pad  & ld_pad ;
  assign n17217 = ~\u0_w_reg[3][24]/P0001  & ~n16871 ;
  assign n17218 = \u0_w_reg[3][24]/P0001  & n16871 ;
  assign n17219 = ~n17217 & ~n17218 ;
  assign n17221 = ~n17180 & n17219 ;
  assign n17220 = n17180 & ~n17219 ;
  assign n17222 = ~ld_pad & ~n17220 ;
  assign n17223 = ~n17221 & n17222 ;
  assign n17224 = ~n17216 & ~n17223 ;
  assign n17226 = \u0_w_reg[3][26]/P0001  & ~n17195 ;
  assign n17225 = ~\u0_w_reg[3][26]/P0001  & n17195 ;
  assign n17227 = ~ld_pad & ~n17225 ;
  assign n17228 = ~n17226 & n17227 ;
  assign n17229 = \key[26]_pad  & ld_pad ;
  assign n17230 = ~n17228 & ~n17229 ;
  assign n17232 = \u0_w_reg[3][30]/P0001  & ~n17204 ;
  assign n17231 = ~\u0_w_reg[3][30]/P0001  & n17204 ;
  assign n17233 = ~ld_pad & ~n17231 ;
  assign n17234 = ~n17232 & n17233 ;
  assign n17235 = \key[30]_pad  & ld_pad ;
  assign n17236 = ~n17234 & ~n17235 ;
  assign n17238 = \u0_w_reg[3][31]/P0001  & ~n17213 ;
  assign n17237 = ~\u0_w_reg[3][31]/P0001  & n17213 ;
  assign n17239 = ~ld_pad & ~n17237 ;
  assign n17240 = ~n17238 & n17239 ;
  assign n17241 = \key[31]_pad  & ld_pad ;
  assign n17242 = ~n17240 & ~n17241 ;
  assign n17243 = ~ld_pad & n15880 ;
  assign n17244 = \key[117]_pad  & ld_pad ;
  assign n17245 = ~n17243 & ~n17244 ;
  assign n17247 = \u0_w_reg[1][21]/P0001  & n15880 ;
  assign n17246 = ~\u0_w_reg[1][21]/P0001  & ~n15880 ;
  assign n17248 = ~ld_pad & ~n17246 ;
  assign n17249 = ~n17247 & n17248 ;
  assign n17250 = \key[85]_pad  & ld_pad ;
  assign n17251 = ~n17249 & ~n17250 ;
  assign n17253 = \u0_w_reg[3][21]/P0001  & ~n15886 ;
  assign n17252 = ~\u0_w_reg[3][21]/P0001  & n15886 ;
  assign n17254 = ~ld_pad & ~n17252 ;
  assign n17255 = ~n17253 & n17254 ;
  assign n17256 = \key[21]_pad  & ld_pad ;
  assign n17257 = ~n17255 & ~n17256 ;
  assign n17258 = ~\key[39]_pad  & ld_pad ;
  assign n17264 = ~\u0_w_reg[3][28]/P0001  & ~n16098 ;
  assign n17263 = \u0_w_reg[3][28]/P0001  & ~n16079 ;
  assign n17265 = n16036 & ~n17263 ;
  assign n17266 = ~n17264 & n17265 ;
  assign n17267 = ~n16143 & ~n16407 ;
  assign n17259 = \u0_w_reg[3][30]/P0001  & n16105 ;
  assign n17260 = n16386 & n17259 ;
  assign n17261 = ~\u0_w_reg[3][28]/P0001  & n16122 ;
  assign n17262 = n16019 & n17261 ;
  assign n17268 = ~n17260 & ~n17262 ;
  assign n17269 = n17267 & n17268 ;
  assign n17270 = ~n17266 & n17269 ;
  assign n17272 = ~n16099 & n17263 ;
  assign n17273 = ~n16058 & ~n16140 ;
  assign n17274 = ~n17272 & n17273 ;
  assign n17275 = ~\u0_w_reg[3][26]/P0001  & ~n17274 ;
  assign n17277 = ~\u0_w_reg[3][28]/P0001  & n16171 ;
  assign n17278 = n16036 & n17277 ;
  assign n17271 = \u0_w_reg[3][28]/P0001  & n16140 ;
  assign n17276 = n16032 & n16079 ;
  assign n17279 = ~n17271 & ~n17276 ;
  assign n17280 = ~n17278 & n17279 ;
  assign n17281 = ~n17275 & n17280 ;
  assign n17282 = n17270 & n17281 ;
  assign n17283 = \u0_w_reg[3][24]/P0001  & ~n17282 ;
  assign n17285 = n16017 & n16087 ;
  assign n17286 = ~n16129 & ~n17285 ;
  assign n17287 = ~\u0_w_reg[3][29]/P0001  & n16066 ;
  assign n17288 = ~\u0_w_reg[3][26]/P0001  & ~n16141 ;
  assign n17289 = ~n17287 & n17288 ;
  assign n17290 = n17286 & n17289 ;
  assign n17291 = n16388 & n16392 ;
  assign n17292 = \u0_w_reg[3][26]/P0001  & ~n16063 ;
  assign n17293 = ~n16144 & n17292 ;
  assign n17294 = ~n17291 & n17293 ;
  assign n17295 = ~n17290 & ~n17294 ;
  assign n17284 = n16117 & n17277 ;
  assign n17296 = ~\u0_w_reg[3][25]/P0001  & ~n16385 ;
  assign n17297 = ~n17284 & n17296 ;
  assign n17298 = ~n17295 & n17297 ;
  assign n17299 = ~n17283 & n17298 ;
  assign n17300 = ~n16014 & ~n16438 ;
  assign n17311 = \u0_w_reg[3][31]/P0001  & ~n17300 ;
  assign n17312 = ~n16118 & ~n17311 ;
  assign n17313 = ~\u0_w_reg[3][27]/P0001  & ~n17312 ;
  assign n17314 = \u0_w_reg[3][26]/P0001  & ~n16013 ;
  assign n17315 = ~n16172 & n17314 ;
  assign n17316 = ~n17313 & n17315 ;
  assign n17317 = ~n16040 & ~n16428 ;
  assign n17318 = \u0_w_reg[3][29]/P0001  & n16051 ;
  assign n17319 = n17317 & ~n17318 ;
  assign n17320 = \u0_w_reg[3][27]/P0001  & ~n17319 ;
  assign n17321 = ~n16080 & n17289 ;
  assign n17322 = ~n17320 & n17321 ;
  assign n17323 = ~n17316 & ~n17322 ;
  assign n17301 = \u0_w_reg[3][27]/P0001  & n16025 ;
  assign n17302 = ~n16125 & ~n17301 ;
  assign n17303 = n17300 & n17302 ;
  assign n17304 = \u0_w_reg[3][26]/P0001  & ~n17303 ;
  assign n17305 = n16171 & n16386 ;
  assign n17306 = ~\u0_w_reg[3][30]/P0001  & n17305 ;
  assign n17307 = ~n17291 & ~n17306 ;
  assign n17308 = ~n17304 & n17307 ;
  assign n17309 = n17270 & n17308 ;
  assign n17310 = \u0_w_reg[3][24]/P0001  & ~n17309 ;
  assign n17324 = \u0_w_reg[3][25]/P0001  & ~n17310 ;
  assign n17325 = ~n17323 & n17324 ;
  assign n17326 = ~n17299 & ~n17325 ;
  assign n17346 = ~\u0_w_reg[3][26]/P0001  & ~n16111 ;
  assign n17345 = n16094 & n16105 ;
  assign n17347 = ~\u0_w_reg[3][25]/P0001  & n16359 ;
  assign n17348 = ~n17345 & ~n17347 ;
  assign n17349 = n17286 & n17348 ;
  assign n17350 = n17346 & n17349 ;
  assign n17351 = n16011 & n16158 ;
  assign n17352 = \u0_w_reg[3][26]/P0001  & ~n16047 ;
  assign n17353 = ~n17351 & n17352 ;
  assign n17354 = ~n17350 & ~n17353 ;
  assign n17332 = n16036 & n16160 ;
  assign n17331 = ~\u0_w_reg[3][30]/P0001  & n16146 ;
  assign n17333 = \u0_w_reg[3][25]/P0001  & ~n17331 ;
  assign n17334 = ~n17332 & n17333 ;
  assign n17327 = \u0_w_reg[3][28]/P0001  & n16100 ;
  assign n17328 = n16012 & n16019 ;
  assign n17329 = ~n16046 & ~n17328 ;
  assign n17330 = ~\u0_w_reg[3][26]/P0001  & ~n17329 ;
  assign n17335 = ~n17327 & ~n17330 ;
  assign n17336 = n17334 & n17335 ;
  assign n17337 = ~\u0_w_reg[3][28]/P0001  & n16146 ;
  assign n17340 = ~\u0_w_reg[3][25]/P0001  & ~n17337 ;
  assign n17338 = n16122 & n16388 ;
  assign n17339 = \u0_w_reg[3][26]/P0001  & n16052 ;
  assign n17341 = ~n17338 & ~n17339 ;
  assign n17342 = n17340 & n17341 ;
  assign n17343 = ~n17336 & ~n17342 ;
  assign n17344 = ~\u0_w_reg[3][31]/P0001  & n16123 ;
  assign n17355 = ~n17343 & ~n17344 ;
  assign n17356 = ~n17354 & n17355 ;
  assign n17357 = ~\u0_w_reg[3][24]/P0001  & ~n17356 ;
  assign n17358 = ~n17326 & ~n17357 ;
  assign n17359 = \u0_w_reg[0][7]/P0001  & ~n17358 ;
  assign n17360 = ~\u0_w_reg[0][7]/P0001  & n17358 ;
  assign n17361 = ~n17359 & ~n17360 ;
  assign n17362 = \u0_w_reg[1][7]/P0001  & ~\u0_w_reg[2][7]/P0001  ;
  assign n17363 = ~\u0_w_reg[1][7]/P0001  & \u0_w_reg[2][7]/P0001  ;
  assign n17364 = ~n17362 & ~n17363 ;
  assign n17365 = n17361 & n17364 ;
  assign n17366 = ~n17361 & ~n17364 ;
  assign n17367 = ~n17365 & ~n17366 ;
  assign n17368 = ~ld_pad & n17367 ;
  assign n17369 = ~n17258 & ~n17368 ;
  assign n17370 = ~ld_pad & n16001 ;
  assign n17371 = \key[115]_pad  & ld_pad ;
  assign n17372 = ~n17370 & ~n17371 ;
  assign n17374 = \u0_w_reg[1][19]/P0001  & n16001 ;
  assign n17373 = ~\u0_w_reg[1][19]/P0001  & ~n16001 ;
  assign n17375 = ~ld_pad & ~n17373 ;
  assign n17376 = ~n17374 & n17375 ;
  assign n17377 = \key[83]_pad  & ld_pad ;
  assign n17378 = ~n17376 & ~n17377 ;
  assign n17380 = \u0_w_reg[3][19]/P0001  & ~n16007 ;
  assign n17379 = ~\u0_w_reg[3][19]/P0001  & n16007 ;
  assign n17381 = ~ld_pad & ~n17379 ;
  assign n17382 = ~n17380 & n17381 ;
  assign n17383 = \key[19]_pad  & ld_pad ;
  assign n17384 = ~n17382 & ~n17383 ;
  assign n17385 = ~ld_pad & n16190 ;
  assign n17386 = \key[101]_pad  & ld_pad ;
  assign n17387 = ~n17385 & ~n17386 ;
  assign n17389 = \u0_w_reg[1][5]/P0001  & n16190 ;
  assign n17388 = ~\u0_w_reg[1][5]/P0001  & ~n16190 ;
  assign n17390 = ~ld_pad & ~n17388 ;
  assign n17391 = ~n17389 & n17390 ;
  assign n17392 = \key[69]_pad  & ld_pad ;
  assign n17393 = ~n17391 & ~n17392 ;
  assign n17395 = \u0_w_reg[3][5]/P0001  & ~n16196 ;
  assign n17394 = ~\u0_w_reg[3][5]/P0001  & n16196 ;
  assign n17396 = ~ld_pad & ~n17394 ;
  assign n17397 = ~n17395 & n17396 ;
  assign n17398 = \key[5]_pad  & ld_pad ;
  assign n17399 = ~n17397 & ~n17398 ;
  assign n17400 = ~\key[32]_pad  & ld_pad ;
  assign n17406 = ~n16450 & ~n17306 ;
  assign n17407 = \u0_w_reg[3][28]/P0001  & ~n17406 ;
  assign n17402 = ~\u0_w_reg[3][27]/P0001  & n16052 ;
  assign n17403 = \u0_w_reg[3][29]/P0001  & n17259 ;
  assign n17404 = ~n17402 & ~n17403 ;
  assign n17405 = \u0_w_reg[3][26]/P0001  & ~n17404 ;
  assign n17408 = ~\u0_w_reg[3][25]/P0001  & ~n17285 ;
  assign n17401 = ~\u0_w_reg[3][29]/P0001  & n16032 ;
  assign n17409 = ~n16044 & ~n17401 ;
  assign n17410 = n17408 & n17409 ;
  assign n17411 = ~n17405 & n17410 ;
  assign n17412 = ~n17407 & n17411 ;
  assign n17413 = ~\u0_w_reg[3][26]/P0001  & n16011 ;
  assign n17414 = ~n16161 & ~n17413 ;
  assign n17415 = n16384 & n17414 ;
  assign n17416 = ~n17412 & ~n17415 ;
  assign n17418 = ~n16047 & ~n17337 ;
  assign n17419 = \u0_w_reg[3][26]/P0001  & ~n16443 ;
  assign n17420 = ~n16050 & n17419 ;
  assign n17421 = n17418 & n17420 ;
  assign n17422 = \u0_w_reg[3][27]/P0001  & n16019 ;
  assign n17423 = ~\u0_w_reg[3][26]/P0001  & ~n17422 ;
  assign n17424 = ~n16093 & ~n16407 ;
  assign n17425 = ~n16038 & n17424 ;
  assign n17426 = n17423 & n17425 ;
  assign n17427 = ~n17421 & ~n17426 ;
  assign n17417 = ~\u0_w_reg[3][28]/P0001  & n16060 ;
  assign n17428 = ~\u0_w_reg[3][27]/P0001  & n16058 ;
  assign n17429 = \u0_w_reg[3][24]/P0001  & ~n17428 ;
  assign n17430 = ~n17417 & n17429 ;
  assign n17431 = ~n17427 & n17430 ;
  assign n17432 = ~n17416 & n17431 ;
  assign n17437 = ~\u0_w_reg[3][27]/P0001  & ~n17317 ;
  assign n17438 = ~\u0_w_reg[3][26]/P0001  & n16066 ;
  assign n17435 = \u0_w_reg[3][26]/P0001  & n16145 ;
  assign n17436 = ~n16392 & n17435 ;
  assign n17439 = ~\u0_w_reg[3][25]/P0001  & ~n17436 ;
  assign n17440 = ~n17438 & n17439 ;
  assign n17441 = ~n17437 & n17440 ;
  assign n17442 = n16012 & n16142 ;
  assign n17445 = \u0_w_reg[3][25]/P0001  & ~n17305 ;
  assign n17443 = n16020 & n16392 ;
  assign n17444 = ~n16045 & n16051 ;
  assign n17446 = ~n17443 & ~n17444 ;
  assign n17447 = n17445 & n17446 ;
  assign n17448 = ~n17442 & n17447 ;
  assign n17449 = ~n17441 & ~n17448 ;
  assign n17450 = n16087 & n16094 ;
  assign n17451 = n16363 & ~n17450 ;
  assign n17452 = ~\u0_w_reg[3][26]/P0001  & ~n17451 ;
  assign n17433 = ~n16019 & ~n17318 ;
  assign n17434 = n17261 & ~n17433 ;
  assign n17453 = ~\u0_w_reg[3][24]/P0001  & ~n17434 ;
  assign n17454 = ~n17452 & n17453 ;
  assign n17455 = ~n17449 & n17454 ;
  assign n17456 = ~n17432 & ~n17455 ;
  assign n17474 = n16051 & n16112 ;
  assign n17473 = ~n16026 & n16140 ;
  assign n17475 = ~n16028 & ~n17473 ;
  assign n17476 = ~n17474 & n17475 ;
  assign n17477 = ~\u0_w_reg[3][26]/P0001  & ~n17476 ;
  assign n17470 = \u0_w_reg[3][26]/P0001  & n16087 ;
  assign n17471 = ~n16011 & ~n16059 ;
  assign n17472 = n17470 & ~n17471 ;
  assign n17478 = ~n16104 & ~n17472 ;
  assign n17479 = ~n17477 & n17478 ;
  assign n17480 = ~\u0_w_reg[3][25]/P0001  & ~n17479 ;
  assign n17457 = n16020 & n16117 ;
  assign n17458 = n16018 & n16036 ;
  assign n17459 = ~n17457 & ~n17458 ;
  assign n17460 = \u0_w_reg[3][30]/P0001  & ~n17459 ;
  assign n17461 = ~n16060 & ~n16162 ;
  assign n17462 = \u0_w_reg[3][26]/P0001  & ~n17461 ;
  assign n17465 = ~\u0_w_reg[3][26]/P0001  & n16385 ;
  assign n17463 = ~\u0_w_reg[3][31]/P0001  & n17450 ;
  assign n17464 = \u0_w_reg[3][27]/P0001  & n16118 ;
  assign n17466 = ~n17463 & ~n17464 ;
  assign n17467 = ~n17465 & n17466 ;
  assign n17468 = ~n17462 & n17467 ;
  assign n17469 = \u0_w_reg[3][25]/P0001  & ~n17468 ;
  assign n17481 = ~n17460 & ~n17469 ;
  assign n17482 = ~n17480 & n17481 ;
  assign n17483 = ~n17456 & n17482 ;
  assign n17484 = \u0_w_reg[0][0]/P0001  & ~n17483 ;
  assign n17485 = ~\u0_w_reg[0][0]/P0001  & n17483 ;
  assign n17486 = ~n17484 & ~n17485 ;
  assign n17487 = \u0_w_reg[1][0]/P0001  & ~\u0_w_reg[2][0]/P0001  ;
  assign n17488 = ~\u0_w_reg[1][0]/P0001  & \u0_w_reg[2][0]/P0001  ;
  assign n17489 = ~n17487 & ~n17488 ;
  assign n17490 = n17486 & n17489 ;
  assign n17491 = ~n17486 & ~n17489 ;
  assign n17492 = ~n17490 & ~n17491 ;
  assign n17493 = ~ld_pad & n17492 ;
  assign n17494 = ~n17400 & ~n17493 ;
  assign n17495 = ~\key[42]_pad  & ld_pad ;
  assign n17552 = ~n16572 & ~n16697 ;
  assign n17553 = ~n16737 & n17552 ;
  assign n17554 = ~\u0_w_reg[3][2]/P0001  & ~n17553 ;
  assign n17555 = ~n16478 & ~n16493 ;
  assign n17556 = n16524 & ~n17555 ;
  assign n17557 = n16493 & ~n16658 ;
  assign n17558 = ~n16667 & n17557 ;
  assign n17561 = ~\u0_w_reg[3][1]/P0001  & ~n17558 ;
  assign n17559 = n16588 & n16753 ;
  assign n17560 = n16526 & n16667 ;
  assign n17562 = ~n17559 & ~n17560 ;
  assign n17563 = n17561 & n17562 ;
  assign n17564 = ~n17556 & n17563 ;
  assign n17565 = ~n17554 & n17564 ;
  assign n17572 = ~n16497 & ~n16627 ;
  assign n17573 = n16570 & n16667 ;
  assign n17574 = n17572 & ~n17573 ;
  assign n17575 = ~\u0_w_reg[3][2]/P0001  & ~n17574 ;
  assign n17566 = \u0_w_reg[3][4]/P0001  & n16521 ;
  assign n17567 = ~n16520 & ~n17566 ;
  assign n17568 = \u0_w_reg[3][7]/P0001  & ~n17567 ;
  assign n17533 = \u0_w_reg[3][3]/P0001  & n16521 ;
  assign n17569 = n16658 & n17533 ;
  assign n17570 = ~n17568 & ~n17569 ;
  assign n17571 = \u0_w_reg[3][2]/P0001  & ~n17570 ;
  assign n17576 = \u0_w_reg[3][1]/P0001  & ~n16543 ;
  assign n17577 = ~n17571 & n17576 ;
  assign n17578 = ~n17575 & n17577 ;
  assign n17579 = ~n17565 & ~n17578 ;
  assign n17510 = ~n16604 & ~n16674 ;
  assign n17505 = n16520 & n16551 ;
  assign n17511 = ~n16745 & ~n17505 ;
  assign n17512 = n17510 & n17511 ;
  assign n17507 = ~\u0_w_reg[3][5]/P0001  & ~n16554 ;
  assign n17508 = n16622 & ~n17507 ;
  assign n17509 = ~\u0_w_reg[3][1]/P0001  & ~n16550 ;
  assign n17513 = ~n16696 & n17509 ;
  assign n17514 = ~n17508 & n17513 ;
  assign n17515 = n17512 & n17514 ;
  assign n17519 = ~\u0_w_reg[3][4]/P0001  & n16548 ;
  assign n17520 = \u0_w_reg[3][2]/P0001  & n17519 ;
  assign n17516 = ~\u0_w_reg[3][2]/P0001  & \u0_w_reg[3][3]/P0001  ;
  assign n17517 = n16495 & n16658 ;
  assign n17518 = n17516 & n17517 ;
  assign n17521 = \u0_w_reg[3][1]/P0001  & ~n17518 ;
  assign n17522 = ~n17520 & n17521 ;
  assign n17523 = ~n17515 & ~n17522 ;
  assign n17500 = n16505 & n16551 ;
  assign n17501 = \u0_w_reg[3][5]/P0001  & n16541 ;
  assign n17502 = ~n17500 & ~n17501 ;
  assign n17503 = ~n16573 & n17502 ;
  assign n17504 = n16524 & ~n17503 ;
  assign n17524 = \u0_w_reg[3][0]/P0001  & ~n16730 ;
  assign n17506 = ~\u0_w_reg[3][6]/P0001  & n17505 ;
  assign n17496 = \u0_w_reg[3][5]/P0001  & n16745 ;
  assign n17497 = \u0_w_reg[3][1]/P0001  & ~\u0_w_reg[3][2]/P0001  ;
  assign n17498 = ~n16488 & n17497 ;
  assign n17499 = n16580 & n17498 ;
  assign n17525 = ~n17496 & ~n17499 ;
  assign n17526 = ~n17506 & n17525 ;
  assign n17527 = n17524 & n17526 ;
  assign n17528 = ~n17504 & n17527 ;
  assign n17529 = ~n17523 & n17528 ;
  assign n17530 = n16488 & n16492 ;
  assign n17531 = \u0_w_reg[3][1]/P0001  & ~n17530 ;
  assign n17534 = ~\u0_w_reg[3][2]/P0001  & ~n17533 ;
  assign n17532 = \u0_w_reg[3][3]/P0001  & n16541 ;
  assign n17535 = ~n16481 & ~n17532 ;
  assign n17536 = n17534 & n17535 ;
  assign n17537 = \u0_w_reg[3][2]/P0001  & ~n16622 ;
  assign n17538 = ~n16657 & n17537 ;
  assign n17539 = ~n17536 & ~n17538 ;
  assign n17540 = n17531 & ~n17539 ;
  assign n17541 = n16551 & n17516 ;
  assign n17542 = ~\u0_w_reg[3][1]/P0001  & ~n16529 ;
  assign n17543 = ~n17541 & n17542 ;
  assign n17544 = ~n17540 & ~n17543 ;
  assign n17545 = \u0_w_reg[3][4]/P0001  & n16616 ;
  assign n17546 = n16586 & n16729 ;
  assign n17547 = ~\u0_w_reg[3][0]/P0001  & ~n16563 ;
  assign n17548 = ~n17546 & n17547 ;
  assign n17549 = ~n17545 & n17548 ;
  assign n17550 = ~n17544 & n17549 ;
  assign n17551 = ~n17529 & ~n17550 ;
  assign n17580 = ~n16574 & ~n16753 ;
  assign n17581 = \u0_w_reg[3][2]/P0001  & n16520 ;
  assign n17582 = ~n17580 & n17581 ;
  assign n17583 = ~n16606 & ~n17582 ;
  assign n17584 = ~n17551 & n17583 ;
  assign n17585 = ~n17579 & n17584 ;
  assign n17586 = \u0_w_reg[0][10]/P0001  & ~n17585 ;
  assign n17587 = ~\u0_w_reg[0][10]/P0001  & n17585 ;
  assign n17588 = ~n17586 & ~n17587 ;
  assign n17589 = \u0_w_reg[1][10]/P0001  & ~\u0_w_reg[2][10]/P0001  ;
  assign n17590 = ~\u0_w_reg[1][10]/P0001  & \u0_w_reg[2][10]/P0001  ;
  assign n17591 = ~n17589 & ~n17590 ;
  assign n17592 = n17588 & n17591 ;
  assign n17593 = ~n17588 & ~n17591 ;
  assign n17594 = ~n17592 & ~n17593 ;
  assign n17595 = ~ld_pad & n17594 ;
  assign n17596 = ~n17495 & ~n17595 ;
  assign n17597 = ~\key[48]_pad  & ld_pad ;
  assign n17601 = ~n15805 & ~n15976 ;
  assign n17602 = ~\u0_w_reg[3][11]/P0001  & ~n17601 ;
  assign n17604 = \u0_w_reg[3][10]/P0001  & n15780 ;
  assign n17605 = ~n15919 & n17604 ;
  assign n17603 = ~\u0_w_reg[3][10]/P0001  & n15737 ;
  assign n17606 = ~\u0_w_reg[3][9]/P0001  & ~n17603 ;
  assign n17607 = ~n17605 & n17606 ;
  assign n17608 = ~n17602 & n17607 ;
  assign n17611 = ~\u0_w_reg[3][15]/P0001  & n15791 ;
  assign n17612 = ~n15704 & ~n17611 ;
  assign n17613 = \u0_w_reg[3][11]/P0001  & ~n17612 ;
  assign n17614 = \u0_w_reg[3][9]/P0001  & ~n15820 ;
  assign n17609 = ~\u0_w_reg[3][11]/P0001  & n15736 ;
  assign n17610 = n15814 & n15847 ;
  assign n17615 = ~n17609 & ~n17610 ;
  assign n17616 = n17614 & n17615 ;
  assign n17617 = ~n17613 & n17616 ;
  assign n17618 = ~n17608 & ~n17617 ;
  assign n17619 = n15709 & n15756 ;
  assign n17620 = ~n15954 & ~n17619 ;
  assign n17621 = ~n15753 & n17620 ;
  assign n17622 = ~\u0_w_reg[3][10]/P0001  & ~n17621 ;
  assign n17598 = \u0_w_reg[3][13]/P0001  & n15736 ;
  assign n17599 = ~n15708 & ~n17598 ;
  assign n17600 = n15800 & ~n17599 ;
  assign n17623 = ~\u0_w_reg[3][8]/P0001  & ~n17600 ;
  assign n17624 = ~n17622 & n17623 ;
  assign n17625 = ~n17618 & n17624 ;
  assign n17626 = ~n15704 & ~n17609 ;
  assign n17627 = ~\u0_w_reg[3][13]/P0001  & ~n17626 ;
  assign n17628 = ~n15851 & ~n17627 ;
  assign n17629 = \u0_w_reg[3][10]/P0001  & ~n17628 ;
  assign n17633 = n15802 & n15847 ;
  assign n17630 = n15709 & n15719 ;
  assign n17631 = \u0_w_reg[3][13]/P0001  & ~n15742 ;
  assign n17632 = n15724 & ~n17631 ;
  assign n17634 = ~n17630 & ~n17632 ;
  assign n17635 = ~n17633 & n17634 ;
  assign n17636 = ~n17629 & n17635 ;
  assign n17637 = ~\u0_w_reg[3][9]/P0001  & ~n17636 ;
  assign n17638 = n15724 & n15780 ;
  assign n17639 = ~n15755 & ~n17638 ;
  assign n17640 = \u0_w_reg[3][10]/P0001  & ~n15989 ;
  assign n17641 = ~n15753 & n17640 ;
  assign n17642 = n17639 & n17641 ;
  assign n17644 = \u0_w_reg[3][11]/P0001  & n15708 ;
  assign n17645 = ~\u0_w_reg[3][10]/P0001  & ~n17644 ;
  assign n17643 = n15719 & n15751 ;
  assign n17646 = ~n15915 & ~n17643 ;
  assign n17647 = ~n15705 & n17646 ;
  assign n17648 = n17645 & n17647 ;
  assign n17649 = ~n17642 & ~n17648 ;
  assign n17650 = ~\u0_w_reg[3][13]/P0001  & ~n15736 ;
  assign n17651 = ~\u0_w_reg[3][10]/P0001  & ~n15773 ;
  assign n17652 = ~n17650 & n17651 ;
  assign n17653 = ~n15826 & ~n17652 ;
  assign n17654 = \u0_w_reg[3][9]/P0001  & ~n17653 ;
  assign n17655 = n15724 & n15814 ;
  assign n17656 = ~\u0_w_reg[3][14]/P0001  & n17655 ;
  assign n17657 = \u0_w_reg[3][8]/P0001  & ~n15784 ;
  assign n17658 = ~n17656 & n17657 ;
  assign n17659 = ~n17654 & n17658 ;
  assign n17660 = ~n17649 & n17659 ;
  assign n17661 = ~n17637 & n17660 ;
  assign n17662 = ~n17625 & ~n17661 ;
  assign n17663 = n15720 & n15893 ;
  assign n17664 = n15703 & n15849 ;
  assign n17665 = ~n17663 & ~n17664 ;
  assign n17666 = \u0_w_reg[3][14]/P0001  & ~n17665 ;
  assign n17672 = n15773 & n15822 ;
  assign n17673 = ~n15838 & ~n15850 ;
  assign n17674 = ~n17672 & n17673 ;
  assign n17675 = n15847 & ~n17674 ;
  assign n17669 = n15756 & n15896 ;
  assign n17670 = ~n15930 & ~n17669 ;
  assign n17671 = \u0_w_reg[3][10]/P0001  & ~n17670 ;
  assign n17667 = n15713 & n15822 ;
  assign n17668 = n15849 & n17667 ;
  assign n17676 = ~\u0_w_reg[3][9]/P0001  & ~n15861 ;
  assign n17677 = ~n17668 & n17676 ;
  assign n17678 = ~n17671 & n17677 ;
  assign n17679 = ~n17675 & n17678 ;
  assign n17683 = \u0_w_reg[3][12]/P0001  & n15708 ;
  assign n17684 = n15893 & n17683 ;
  assign n17682 = n15724 & n15773 ;
  assign n17685 = ~n17619 & ~n17682 ;
  assign n17686 = ~n17684 & n17685 ;
  assign n17687 = ~\u0_w_reg[3][15]/P0001  & ~n17686 ;
  assign n17681 = n15743 & n15803 ;
  assign n17680 = ~\u0_w_reg[3][10]/P0001  & n15941 ;
  assign n17688 = \u0_w_reg[3][9]/P0001  & ~n17680 ;
  assign n17689 = ~n17681 & n17688 ;
  assign n17690 = ~n17687 & n17689 ;
  assign n17691 = ~n17679 & ~n17690 ;
  assign n17692 = ~n17666 & ~n17691 ;
  assign n17693 = ~n17662 & n17692 ;
  assign n17694 = \u0_w_reg[0][16]/P0001  & ~n17693 ;
  assign n17695 = ~\u0_w_reg[0][16]/P0001  & n17693 ;
  assign n17696 = ~n17694 & ~n17695 ;
  assign n17697 = \u0_w_reg[1][16]/P0001  & ~\u0_w_reg[2][16]/P0001  ;
  assign n17698 = ~\u0_w_reg[1][16]/P0001  & \u0_w_reg[2][16]/P0001  ;
  assign n17699 = ~n17697 & ~n17698 ;
  assign n17700 = n17696 & n17699 ;
  assign n17701 = ~n17696 & ~n17699 ;
  assign n17702 = ~n17700 & ~n17701 ;
  assign n17703 = ~ld_pad & n17702 ;
  assign n17704 = ~n17597 & ~n17703 ;
  assign n17705 = ~\key[50]_pad  & ld_pad ;
  assign n17743 = n15725 & n15893 ;
  assign n17742 = n15778 & n15860 ;
  assign n17747 = ~n17630 & ~n17742 ;
  assign n17748 = ~n17743 & n17747 ;
  assign n17749 = ~n15731 & ~n17611 ;
  assign n17744 = ~\u0_w_reg[3][13]/P0001  & ~n15782 ;
  assign n17745 = n17609 & ~n17744 ;
  assign n17746 = ~\u0_w_reg[3][9]/P0001  & ~n15970 ;
  assign n17750 = ~n17745 & n17746 ;
  assign n17751 = n17749 & n17750 ;
  assign n17752 = n17748 & n17751 ;
  assign n17753 = n15822 & n15860 ;
  assign n17754 = \u0_w_reg[3][9]/P0001  & ~n17753 ;
  assign n17755 = ~n17668 & n17754 ;
  assign n17756 = ~n17752 & ~n17755 ;
  assign n17737 = \u0_w_reg[3][12]/P0001  & n15773 ;
  assign n17738 = ~\u0_w_reg[3][15]/P0001  & n17737 ;
  assign n17739 = ~n15826 & ~n15840 ;
  assign n17740 = ~n17738 & n17739 ;
  assign n17741 = n15799 & ~n17740 ;
  assign n17757 = \u0_w_reg[3][10]/P0001  & n15784 ;
  assign n17762 = \u0_w_reg[3][8]/P0001  & ~n17669 ;
  assign n17758 = n15736 & n15929 ;
  assign n17759 = \u0_w_reg[3][12]/P0001  & ~n15919 ;
  assign n17760 = n15726 & ~n15773 ;
  assign n17761 = n17759 & n17760 ;
  assign n17763 = ~n17758 & ~n17761 ;
  assign n17764 = n17762 & n17763 ;
  assign n17765 = ~n17757 & n17764 ;
  assign n17766 = ~n17741 & n17765 ;
  assign n17767 = ~n17756 & n17766 ;
  assign n17768 = n15719 & n15849 ;
  assign n17769 = ~\u0_w_reg[3][9]/P0001  & ~n15941 ;
  assign n17770 = ~n17768 & n17769 ;
  assign n17772 = \u0_w_reg[3][11]/P0001  & n15786 ;
  assign n17773 = ~n15823 & ~n17772 ;
  assign n17774 = n17645 & n17773 ;
  assign n17775 = \u0_w_reg[3][10]/P0001  & ~n15717 ;
  assign n17776 = ~n17609 & n17775 ;
  assign n17777 = ~n17774 & ~n17776 ;
  assign n17771 = ~\u0_w_reg[3][14]/P0001  & n15781 ;
  assign n17778 = \u0_w_reg[3][9]/P0001  & ~n17771 ;
  assign n17779 = ~n17777 & n17778 ;
  assign n17780 = ~n17770 & ~n17779 ;
  assign n17781 = n15708 & n15906 ;
  assign n17782 = \u0_w_reg[3][10]/P0001  & n17781 ;
  assign n17783 = ~\u0_w_reg[3][8]/P0001  & ~n15817 ;
  assign n17784 = ~n15864 & n17783 ;
  assign n17785 = ~n17782 & n17784 ;
  assign n17786 = ~n17780 & n17785 ;
  assign n17787 = ~n17767 & ~n17786 ;
  assign n17708 = ~n15703 & ~n15915 ;
  assign n17709 = n15708 & ~n17708 ;
  assign n17706 = ~n15814 & ~n17598 ;
  assign n17707 = n15709 & ~n17706 ;
  assign n17710 = ~n15896 & ~n17707 ;
  assign n17711 = ~n17709 & n17710 ;
  assign n17712 = \u0_w_reg[3][10]/P0001  & ~n17711 ;
  assign n17713 = \u0_w_reg[3][9]/P0001  & ~n17712 ;
  assign n17714 = ~n15756 & ~n15805 ;
  assign n17715 = \u0_w_reg[3][11]/P0001  & ~n17714 ;
  assign n17716 = ~n15941 & n15974 ;
  assign n17717 = ~n17707 & n17716 ;
  assign n17718 = ~n17715 & n17717 ;
  assign n17719 = \u0_w_reg[3][13]/P0001  & n17609 ;
  assign n17720 = ~\u0_w_reg[3][10]/P0001  & ~n17719 ;
  assign n17721 = n15713 & n15735 ;
  assign n17722 = ~\u0_w_reg[3][15]/P0001  & n17721 ;
  assign n17723 = ~n15960 & ~n17672 ;
  assign n17724 = ~n17722 & n17723 ;
  assign n17725 = n17720 & n17724 ;
  assign n17726 = ~n17718 & ~n17725 ;
  assign n17727 = ~n15751 & n15756 ;
  assign n17728 = ~n15822 & n17727 ;
  assign n17729 = ~n17726 & ~n17728 ;
  assign n17730 = ~n17713 & ~n17729 ;
  assign n17731 = \u0_w_reg[3][15]/P0001  & n17721 ;
  assign n17732 = ~n15815 & ~n17731 ;
  assign n17733 = ~n15752 & n17732 ;
  assign n17734 = ~\u0_w_reg[3][10]/P0001  & ~n17733 ;
  assign n17735 = ~n15788 & ~n17734 ;
  assign n17736 = \u0_w_reg[3][9]/P0001  & ~n17735 ;
  assign n17788 = ~n15990 & ~n17736 ;
  assign n17789 = ~n17730 & n17788 ;
  assign n17790 = ~n17787 & n17789 ;
  assign n17791 = \u0_w_reg[0][18]/P0001  & ~n17790 ;
  assign n17792 = ~\u0_w_reg[0][18]/P0001  & n17790 ;
  assign n17793 = ~n17791 & ~n17792 ;
  assign n17794 = \u0_w_reg[1][18]/P0001  & ~\u0_w_reg[2][18]/P0001  ;
  assign n17795 = ~\u0_w_reg[1][18]/P0001  & \u0_w_reg[2][18]/P0001  ;
  assign n17796 = ~n17794 & ~n17795 ;
  assign n17797 = n17793 & n17796 ;
  assign n17798 = ~n17793 & ~n17796 ;
  assign n17799 = ~n17797 & ~n17798 ;
  assign n17800 = ~ld_pad & n17799 ;
  assign n17801 = ~n17705 & ~n17800 ;
  assign n17808 = n16125 & n16147 ;
  assign n17805 = ~\u0_w_reg[3][27]/P0001  & n16079 ;
  assign n17806 = ~\u0_w_reg[3][31]/P0001  & n17805 ;
  assign n17807 = ~\u0_w_reg[3][26]/P0001  & n16021 ;
  assign n17811 = ~n17806 & ~n17807 ;
  assign n17812 = ~n17808 & n17811 ;
  assign n17802 = \u0_w_reg[3][26]/P0001  & ~n17273 ;
  assign n17803 = n16103 & n16359 ;
  assign n17804 = n16359 & n16392 ;
  assign n17809 = ~n17803 & ~n17804 ;
  assign n17810 = n17408 & n17809 ;
  assign n17813 = ~n17802 & n17810 ;
  assign n17814 = n17812 & n17813 ;
  assign n17815 = ~\u0_w_reg[3][26]/P0001  & ~n16027 ;
  assign n17816 = ~n16164 & ~n16386 ;
  assign n17817 = ~n17815 & n17816 ;
  assign n17818 = \u0_w_reg[3][25]/P0001  & ~n17817 ;
  assign n17819 = ~n17814 & ~n17818 ;
  assign n17820 = \u0_w_reg[3][28]/P0001  & n17318 ;
  assign n17821 = ~n16037 & ~n16161 ;
  assign n17822 = ~n17820 & n17821 ;
  assign n17823 = n16122 & ~n17822 ;
  assign n17825 = ~\u0_w_reg[3][30]/P0001  & n16360 ;
  assign n17826 = ~\u0_w_reg[3][29]/P0001  & n17825 ;
  assign n17829 = \u0_w_reg[3][24]/P0001  & ~n17474 ;
  assign n17824 = n16036 & n16058 ;
  assign n17827 = n16029 & ~n16392 ;
  assign n17828 = n17263 & n17827 ;
  assign n17830 = ~n17824 & ~n17828 ;
  assign n17831 = n17829 & n17830 ;
  assign n17832 = ~n17826 & n17831 ;
  assign n17833 = ~n17823 & n17832 ;
  assign n17834 = ~n17819 & n17833 ;
  assign n17835 = \u0_w_reg[3][27]/P0001  & n16098 ;
  assign n17836 = ~n16406 & ~n17835 ;
  assign n17837 = n17423 & n17836 ;
  assign n17838 = \u0_w_reg[3][26]/P0001  & ~n16015 ;
  assign n17839 = ~n16125 & n17838 ;
  assign n17840 = ~n17837 & ~n17839 ;
  assign n17841 = ~n17331 & ~n17840 ;
  assign n17842 = \u0_w_reg[3][25]/P0001  & ~n17841 ;
  assign n17844 = n16017 & n16117 ;
  assign n17845 = ~n16385 & ~n17844 ;
  assign n17846 = ~\u0_w_reg[3][25]/P0001  & ~n17845 ;
  assign n17843 = n16045 & n16450 ;
  assign n17847 = ~\u0_w_reg[3][24]/P0001  & ~n16091 ;
  assign n17848 = ~n16119 & n17847 ;
  assign n17849 = ~n17843 & n17848 ;
  assign n17850 = ~n17846 & n17849 ;
  assign n17851 = ~n17842 & n17850 ;
  assign n17852 = ~n17834 & ~n17851 ;
  assign n17853 = ~n16172 & ~n17351 ;
  assign n17854 = ~n16124 & n17853 ;
  assign n17855 = ~\u0_w_reg[3][26]/P0001  & ~n17854 ;
  assign n17856 = n16149 & ~n17855 ;
  assign n17857 = ~n16118 & ~n16367 ;
  assign n17858 = n17346 & n17857 ;
  assign n17859 = ~n16094 & ~n16428 ;
  assign n17860 = \u0_w_reg[3][27]/P0001  & ~n17859 ;
  assign n17861 = \u0_w_reg[3][26]/P0001  & ~n16385 ;
  assign n17862 = ~n17860 & n17861 ;
  assign n17863 = ~n17858 & ~n17862 ;
  assign n17864 = n16386 & n17318 ;
  assign n17865 = ~\u0_w_reg[3][25]/P0001  & ~n17864 ;
  assign n17866 = ~n16048 & n16094 ;
  assign n17867 = ~n16039 & n17866 ;
  assign n17868 = n17865 & ~n17867 ;
  assign n17869 = ~n17863 & n17868 ;
  assign n17870 = ~n17856 & ~n17869 ;
  assign n17876 = ~n16171 & ~n17318 ;
  assign n17877 = n17470 & ~n17876 ;
  assign n17871 = \u0_w_reg[3][25]/P0001  & \u0_w_reg[3][26]/P0001  ;
  assign n17872 = ~n16021 & ~n16360 ;
  assign n17873 = n17871 & ~n17872 ;
  assign n17874 = \u0_w_reg[3][25]/P0001  & n16122 ;
  assign n17875 = n16040 & n17874 ;
  assign n17878 = ~n16444 & ~n17875 ;
  assign n17879 = ~n17873 & n17878 ;
  assign n17880 = ~n17877 & n17879 ;
  assign n17881 = ~n17870 & n17880 ;
  assign n17882 = ~n17852 & n17881 ;
  assign n17883 = \u0_w_reg[0][2]/P0001  & ~n17882 ;
  assign n17884 = ~\u0_w_reg[0][2]/P0001  & n17882 ;
  assign n17885 = ~n17883 & ~n17884 ;
  assign n17886 = \u0_w_reg[1][2]/P0001  & n17885 ;
  assign n17887 = ~\u0_w_reg[1][2]/P0001  & ~n17885 ;
  assign n17888 = ~n17886 & ~n17887 ;
  assign n17889 = \u0_w_reg[2][2]/P0001  & n17888 ;
  assign n17890 = ~\u0_w_reg[2][2]/P0001  & ~n17888 ;
  assign n17891 = ~n17889 & ~n17890 ;
  assign n17892 = ~ld_pad & n17891 ;
  assign n17893 = \key[34]_pad  & ld_pad ;
  assign n17894 = ~n17892 & ~n17893 ;
  assign n17895 = ~\key[46]_pad  & ld_pad ;
  assign n17960 = ~\u0_w_reg[3][3]/P0001  & n16627 ;
  assign n17961 = \u0_w_reg[3][4]/P0001  & n16483 ;
  assign n17962 = ~n16490 & ~n17961 ;
  assign n17963 = ~n17960 & n17962 ;
  assign n17964 = \u0_w_reg[3][2]/P0001  & ~n17963 ;
  assign n17959 = n16488 & n16532 ;
  assign n17957 = n16588 & n16653 ;
  assign n17958 = n16476 & n16612 ;
  assign n17965 = ~n17957 & ~n17958 ;
  assign n17966 = ~n17959 & n17965 ;
  assign n17967 = ~n17964 & n17966 ;
  assign n17968 = \u0_w_reg[3][1]/P0001  & ~n17967 ;
  assign n17944 = ~n16627 & ~n16630 ;
  assign n17945 = ~\u0_w_reg[3][2]/P0001  & ~n17944 ;
  assign n17946 = ~n16496 & ~n16522 ;
  assign n17947 = \u0_w_reg[3][2]/P0001  & ~n17946 ;
  assign n17948 = ~n16563 & ~n17559 ;
  assign n17949 = ~n17947 & n17948 ;
  assign n17950 = ~n17945 & n17949 ;
  assign n17951 = ~\u0_w_reg[3][1]/P0001  & ~n17950 ;
  assign n17954 = ~n16494 & ~n16659 ;
  assign n17955 = n16534 & n17954 ;
  assign n17956 = \u0_w_reg[3][2]/P0001  & ~n17955 ;
  assign n17952 = \u0_w_reg[3][4]/P0001  & n16488 ;
  assign n17953 = n16588 & n17952 ;
  assign n17969 = ~\u0_w_reg[3][2]/P0001  & n16495 ;
  assign n17970 = n16658 & n17969 ;
  assign n17971 = ~n17953 & ~n17970 ;
  assign n17972 = ~n17956 & n17971 ;
  assign n17973 = ~n17951 & n17972 ;
  assign n17974 = ~n17968 & n17973 ;
  assign n17975 = \u0_w_reg[3][0]/P0001  & ~n17974 ;
  assign n17896 = n16493 & n16520 ;
  assign n17897 = n16542 & n16667 ;
  assign n17898 = \u0_w_reg[3][2]/P0001  & ~n17897 ;
  assign n17899 = ~n17896 & n17898 ;
  assign n17902 = ~\u0_w_reg[3][2]/P0001  & ~n16590 ;
  assign n17903 = ~n16485 & n17902 ;
  assign n17900 = ~\u0_w_reg[3][3]/P0001  & n16608 ;
  assign n17901 = ~n16548 & n16743 ;
  assign n17904 = ~n17900 & ~n17901 ;
  assign n17905 = n17903 & n17904 ;
  assign n17906 = ~n17899 & ~n17905 ;
  assign n17909 = ~\u0_w_reg[3][1]/P0001  & ~n16510 ;
  assign n17908 = n16520 & n16570 ;
  assign n17910 = ~n17517 & ~n17908 ;
  assign n17911 = n17909 & n17910 ;
  assign n17907 = \u0_w_reg[3][7]/P0001  & n16743 ;
  assign n17912 = ~n16754 & ~n17897 ;
  assign n17913 = ~n17907 & n17912 ;
  assign n17914 = n17911 & n17913 ;
  assign n17917 = ~\u0_w_reg[3][2]/P0001  & ~n16659 ;
  assign n17915 = \u0_w_reg[3][4]/P0001  & n16476 ;
  assign n17916 = ~n16481 & ~n17915 ;
  assign n17918 = ~n16524 & ~n17916 ;
  assign n17919 = ~n17917 & n17918 ;
  assign n17920 = \u0_w_reg[3][1]/P0001  & ~n16737 ;
  assign n17921 = ~n17919 & n17920 ;
  assign n17922 = ~n17914 & ~n17921 ;
  assign n17923 = ~n17906 & ~n17922 ;
  assign n17924 = ~\u0_w_reg[3][0]/P0001  & ~n17923 ;
  assign n17925 = ~n16622 & ~n17530 ;
  assign n17926 = ~\u0_w_reg[3][4]/P0001  & ~n17925 ;
  assign n17927 = ~\u0_w_reg[3][7]/P0001  & n16608 ;
  assign n17928 = ~n17926 & ~n17927 ;
  assign n17929 = \u0_w_reg[3][2]/P0001  & ~n17928 ;
  assign n17930 = ~n17546 & ~n17929 ;
  assign n17931 = \u0_w_reg[3][1]/P0001  & ~n17930 ;
  assign n17933 = ~n16573 & ~n17530 ;
  assign n17934 = ~\u0_w_reg[3][2]/P0001  & ~n17933 ;
  assign n17936 = ~n16556 & ~n16572 ;
  assign n17937 = ~n16527 & n17936 ;
  assign n17932 = n16548 & n16664 ;
  assign n17935 = ~\u0_w_reg[3][2]/P0001  & n16563 ;
  assign n17938 = ~n17932 & ~n17935 ;
  assign n17939 = n17937 & n17938 ;
  assign n17940 = ~n17934 & n17939 ;
  assign n17941 = ~\u0_w_reg[3][1]/P0001  & ~n17940 ;
  assign n17942 = ~n16623 & ~n16631 ;
  assign n17943 = ~n16509 & ~n17942 ;
  assign n17976 = ~n16511 & ~n17943 ;
  assign n17977 = ~n17941 & n17976 ;
  assign n17978 = ~n17931 & n17977 ;
  assign n17979 = ~n17924 & n17978 ;
  assign n17980 = ~n17975 & n17979 ;
  assign n17981 = \u0_w_reg[0][14]/P0001  & ~n17980 ;
  assign n17982 = ~\u0_w_reg[0][14]/P0001  & n17980 ;
  assign n17983 = ~n17981 & ~n17982 ;
  assign n17984 = \u0_w_reg[1][14]/P0001  & ~\u0_w_reg[2][14]/P0001  ;
  assign n17985 = ~\u0_w_reg[1][14]/P0001  & \u0_w_reg[2][14]/P0001  ;
  assign n17986 = ~n17984 & ~n17985 ;
  assign n17987 = n17983 & n17986 ;
  assign n17988 = ~n17983 & ~n17986 ;
  assign n17989 = ~n17987 & ~n17988 ;
  assign n17990 = ~ld_pad & n17989 ;
  assign n17991 = ~n17895 & ~n17990 ;
  assign n17992 = ~\key[54]_pad  & ld_pad ;
  assign n17996 = ~\u0_w_reg[3][10]/P0001  & ~n15816 ;
  assign n17993 = \u0_w_reg[3][10]/P0001  & ~n15838 ;
  assign n17994 = ~n15906 & n17993 ;
  assign n17995 = ~n17720 & ~n17994 ;
  assign n17997 = ~\u0_w_reg[3][9]/P0001  & ~n15817 ;
  assign n17998 = ~n17995 & n17997 ;
  assign n17999 = ~n17996 & n17998 ;
  assign n18000 = \u0_w_reg[3][15]/P0001  & n15710 ;
  assign n18001 = ~n15779 & ~n15850 ;
  assign n18002 = ~n18000 & n18001 ;
  assign n18003 = \u0_w_reg[3][10]/P0001  & ~n18002 ;
  assign n18004 = n15732 & n15847 ;
  assign n18005 = \u0_w_reg[3][9]/P0001  & ~n18004 ;
  assign n18006 = n17639 & n18005 ;
  assign n18007 = ~n18003 & n18006 ;
  assign n18008 = ~n17999 & ~n18007 ;
  assign n18009 = ~n15832 & ~n15920 ;
  assign n18010 = ~n15744 & n18009 ;
  assign n18011 = n15707 & n18010 ;
  assign n18012 = ~\u0_w_reg[3][10]/P0001  & ~n15774 ;
  assign n18013 = ~n17667 & n18012 ;
  assign n18014 = ~n18011 & ~n18013 ;
  assign n18015 = ~n18008 & ~n18014 ;
  assign n18016 = \u0_w_reg[3][8]/P0001  & ~n18015 ;
  assign n18027 = n15709 & n15742 ;
  assign n18029 = ~n17664 & ~n17667 ;
  assign n18030 = ~n18027 & n18029 ;
  assign n18026 = n15799 & n17598 ;
  assign n18017 = n15751 & n15787 ;
  assign n18028 = ~\u0_w_reg[3][9]/P0001  & ~n17655 ;
  assign n18031 = ~n18017 & n18028 ;
  assign n18032 = ~n18026 & n18031 ;
  assign n18033 = n18030 & n18032 ;
  assign n18034 = ~n15824 & n15893 ;
  assign n18035 = ~\u0_w_reg[3][10]/P0001  & n15832 ;
  assign n18036 = \u0_w_reg[3][9]/P0001  & ~n17722 ;
  assign n18037 = ~n18035 & n18036 ;
  assign n18038 = ~n18034 & n18037 ;
  assign n18039 = ~n18033 & ~n18038 ;
  assign n18018 = ~n17619 & ~n18017 ;
  assign n18019 = \u0_w_reg[3][10]/P0001  & ~n18018 ;
  assign n18020 = ~n15741 & ~n15756 ;
  assign n18021 = n15751 & ~n18020 ;
  assign n18022 = n15724 & n17650 ;
  assign n18023 = ~n15939 & ~n18022 ;
  assign n18024 = ~n18021 & n18023 ;
  assign n18025 = ~\u0_w_reg[3][10]/P0001  & ~n18024 ;
  assign n18040 = ~n18019 & ~n18025 ;
  assign n18041 = ~n18039 & n18040 ;
  assign n18042 = ~\u0_w_reg[3][8]/P0001  & ~n18041 ;
  assign n18043 = \u0_w_reg[3][10]/P0001  & ~n15805 ;
  assign n18044 = ~n15865 & n18043 ;
  assign n18045 = n15818 & ~n15826 ;
  assign n18046 = ~n17771 & n18045 ;
  assign n18047 = ~n18044 & ~n18046 ;
  assign n18048 = ~n15930 & ~n15960 ;
  assign n18049 = ~n18047 & n18048 ;
  assign n18050 = ~\u0_w_reg[3][9]/P0001  & ~n18049 ;
  assign n18055 = \u0_w_reg[3][10]/P0001  & \u0_w_reg[3][9]/P0001  ;
  assign n18056 = ~n17609 & ~n17771 ;
  assign n18057 = ~\u0_w_reg[3][12]/P0001  & ~n18056 ;
  assign n18058 = ~n15758 & ~n18057 ;
  assign n18059 = n18055 & ~n18058 ;
  assign n18051 = ~\u0_w_reg[3][15]/P0001  & n17619 ;
  assign n18060 = ~n15892 & ~n18051 ;
  assign n18052 = ~n15920 & ~n17609 ;
  assign n18053 = n15803 & ~n18052 ;
  assign n18054 = n15726 & n15863 ;
  assign n18061 = ~n18053 & ~n18054 ;
  assign n18062 = n18060 & n18061 ;
  assign n18063 = ~n18059 & n18062 ;
  assign n18064 = ~n18050 & n18063 ;
  assign n18065 = ~n18042 & n18064 ;
  assign n18066 = ~n18016 & n18065 ;
  assign n18067 = \u0_w_reg[0][22]/P0001  & ~n18066 ;
  assign n18068 = ~\u0_w_reg[0][22]/P0001  & n18066 ;
  assign n18069 = ~n18067 & ~n18068 ;
  assign n18070 = \u0_w_reg[1][22]/P0001  & ~\u0_w_reg[2][22]/P0001  ;
  assign n18071 = ~\u0_w_reg[1][22]/P0001  & \u0_w_reg[2][22]/P0001  ;
  assign n18072 = ~n18070 & ~n18071 ;
  assign n18073 = n18069 & n18072 ;
  assign n18074 = ~n18069 & ~n18072 ;
  assign n18075 = ~n18073 & ~n18074 ;
  assign n18076 = ~ld_pad & n18075 ;
  assign n18077 = ~n17992 & ~n18076 ;
  assign n18078 = ~\key[38]_pad  & ld_pad ;
  assign n18079 = n16030 & n16386 ;
  assign n18080 = \u0_w_reg[3][25]/P0001  & ~n18079 ;
  assign n18081 = n17418 & n18080 ;
  assign n18086 = ~n16091 & n17865 ;
  assign n18094 = n16173 & n18086 ;
  assign n18095 = ~n18081 & ~n18094 ;
  assign n18096 = ~n16134 & n17815 ;
  assign n18097 = ~n18095 & n18096 ;
  assign n18082 = n16019 & n16360 ;
  assign n18083 = ~n16150 & ~n17259 ;
  assign n18084 = ~n18082 & n18083 ;
  assign n18085 = n18081 & n18084 ;
  assign n18087 = ~n16081 & ~n16158 ;
  assign n18088 = n18086 & n18087 ;
  assign n18089 = ~n18085 & ~n18088 ;
  assign n18090 = \u0_w_reg[3][26]/P0001  & ~n16060 ;
  assign n18091 = ~n16120 & n16404 ;
  assign n18092 = n18090 & n18091 ;
  assign n18093 = ~n18089 & n18092 ;
  assign n18098 = \u0_w_reg[3][24]/P0001  & ~n18093 ;
  assign n18099 = ~n18097 & n18098 ;
  assign n18100 = ~n16051 & n17401 ;
  assign n18103 = ~n16408 & ~n18100 ;
  assign n18101 = ~\u0_w_reg[3][26]/P0001  & ~n16393 ;
  assign n18102 = ~\u0_w_reg[3][27]/P0001  & n16438 ;
  assign n18104 = n18101 & ~n18102 ;
  assign n18105 = n18103 & n18104 ;
  assign n18106 = \u0_w_reg[3][26]/P0001  & ~n17450 ;
  assign n18107 = ~n17327 & n18106 ;
  assign n18108 = ~n18105 & ~n18107 ;
  assign n18110 = n16122 & n17318 ;
  assign n18109 = \u0_w_reg[3][31]/P0001  & n17401 ;
  assign n18113 = ~n17825 & ~n18109 ;
  assign n18114 = ~n18110 & n18113 ;
  assign n18111 = ~\u0_w_reg[3][25]/P0001  & ~n16027 ;
  assign n18112 = ~n17457 & n18111 ;
  assign n18115 = ~n17327 & n18112 ;
  assign n18116 = n18114 & n18115 ;
  assign n18118 = \u0_w_reg[3][28]/P0001  & n16145 ;
  assign n18119 = ~n16406 & ~n18118 ;
  assign n18120 = n16036 & ~n18119 ;
  assign n18117 = ~\u0_w_reg[3][26]/P0001  & n16120 ;
  assign n18121 = \u0_w_reg[3][25]/P0001  & ~n16111 ;
  assign n18122 = ~n18117 & n18121 ;
  assign n18123 = ~n18120 & n18122 ;
  assign n18124 = ~n18116 & ~n18123 ;
  assign n18125 = ~n18108 & ~n18124 ;
  assign n18126 = ~\u0_w_reg[3][24]/P0001  & ~n18125 ;
  assign n18127 = ~\u0_w_reg[3][26]/P0001  & ~n16161 ;
  assign n18128 = ~n16091 & ~n17331 ;
  assign n18129 = n18127 & n18128 ;
  assign n18130 = n16032 & n16051 ;
  assign n18131 = \u0_w_reg[3][26]/P0001  & ~n16428 ;
  assign n18132 = ~n18130 & n18131 ;
  assign n18133 = ~n18129 & ~n18132 ;
  assign n18134 = ~n16367 & ~n16375 ;
  assign n18135 = ~n18133 & n18134 ;
  assign n18136 = ~\u0_w_reg[3][25]/P0001  & ~n18135 ;
  assign n18140 = ~n16169 & ~n17337 ;
  assign n18141 = ~\u0_w_reg[3][30]/P0001  & ~n18140 ;
  assign n18142 = ~n16088 & ~n18141 ;
  assign n18143 = n17871 & ~n18142 ;
  assign n18137 = ~n16449 & ~n17402 ;
  assign n18138 = \u0_w_reg[3][26]/P0001  & ~n18137 ;
  assign n18139 = \u0_w_reg[3][25]/P0001  & n16119 ;
  assign n18144 = ~n16420 & ~n17463 ;
  assign n18145 = ~n18139 & n18144 ;
  assign n18146 = ~n18138 & n18145 ;
  assign n18147 = ~n18143 & n18146 ;
  assign n18148 = ~n18136 & n18147 ;
  assign n18149 = ~n18126 & n18148 ;
  assign n18150 = ~n18099 & n18149 ;
  assign n18151 = \u0_w_reg[0][6]/P0001  & ~n18150 ;
  assign n18152 = ~\u0_w_reg[0][6]/P0001  & n18150 ;
  assign n18153 = ~n18151 & ~n18152 ;
  assign n18154 = \u0_w_reg[1][6]/P0001  & ~\u0_w_reg[2][6]/P0001  ;
  assign n18155 = ~\u0_w_reg[1][6]/P0001  & \u0_w_reg[2][6]/P0001  ;
  assign n18156 = ~n18154 & ~n18155 ;
  assign n18157 = n18153 & n18156 ;
  assign n18158 = ~n18153 & ~n18156 ;
  assign n18159 = ~n18157 & ~n18158 ;
  assign n18160 = ~ld_pad & n18159 ;
  assign n18161 = ~n18078 & ~n18160 ;
  assign n18162 = ~\key[45]_pad  & ld_pad ;
  assign n18194 = \u0_w_reg[3][3]/P0001  & n16570 ;
  assign n18195 = ~n16607 & ~n17952 ;
  assign n18196 = ~\u0_w_reg[3][3]/P0001  & ~n18195 ;
  assign n18197 = ~n18194 & ~n18196 ;
  assign n18198 = ~\u0_w_reg[3][2]/P0001  & ~n18197 ;
  assign n18199 = ~n16556 & ~n16688 ;
  assign n18200 = ~\u0_w_reg[3][7]/P0001  & ~n18199 ;
  assign n18201 = ~n16554 & n16565 ;
  assign n18202 = ~n16490 & ~n16701 ;
  assign n18203 = ~n16543 & n18202 ;
  assign n18204 = ~n18201 & n18203 ;
  assign n18205 = ~n18200 & n18204 ;
  assign n18206 = ~n18198 & n18205 ;
  assign n18207 = \u0_w_reg[3][1]/P0001  & ~n18206 ;
  assign n18208 = ~n16665 & ~n17573 ;
  assign n18209 = ~\u0_w_reg[3][5]/P0001  & ~n18208 ;
  assign n18210 = \u0_w_reg[3][2]/P0001  & n16623 ;
  assign n18211 = ~n16479 & ~n18210 ;
  assign n18212 = ~n18209 & n18211 ;
  assign n18213 = ~\u0_w_reg[3][1]/P0001  & ~n18212 ;
  assign n18214 = \u0_w_reg[3][3]/P0001  & ~n17916 ;
  assign n18215 = n16521 & n16668 ;
  assign n18216 = ~n17519 & ~n18215 ;
  assign n18217 = ~n18214 & n18216 ;
  assign n18218 = \u0_w_reg[3][2]/P0001  & ~n18217 ;
  assign n18219 = ~n16659 & ~n17935 ;
  assign n18220 = ~n17945 & n18219 ;
  assign n18221 = ~n18218 & n18220 ;
  assign n18222 = ~n18213 & n18221 ;
  assign n18223 = ~n18207 & n18222 ;
  assign n18224 = ~\u0_w_reg[3][0]/P0001  & ~n18223 ;
  assign n18176 = ~n16564 & ~n17959 ;
  assign n18175 = n16570 & n16612 ;
  assign n18177 = \u0_w_reg[3][1]/P0001  & ~n18175 ;
  assign n18178 = ~n16624 & n18177 ;
  assign n18179 = n18176 & n18178 ;
  assign n18182 = ~n16650 & ~n16700 ;
  assign n18183 = \u0_w_reg[3][2]/P0001  & ~n18182 ;
  assign n18185 = ~n16530 & ~n16728 ;
  assign n18180 = n16495 & n16586 ;
  assign n18181 = ~\u0_w_reg[3][1]/P0001  & ~n18180 ;
  assign n18184 = ~\u0_w_reg[3][2]/P0001  & n16494 ;
  assign n18186 = n18181 & ~n18184 ;
  assign n18187 = n18185 & n18186 ;
  assign n18188 = ~n18183 & n18187 ;
  assign n18189 = ~n18179 & ~n18188 ;
  assign n18163 = \u0_w_reg[3][4]/P0001  & n16480 ;
  assign n18164 = ~\u0_w_reg[3][4]/P0001  & ~n16482 ;
  assign n18165 = ~n16521 & n18164 ;
  assign n18166 = ~n18163 & ~n18165 ;
  assign n18167 = \u0_w_reg[3][1]/P0001  & ~n18166 ;
  assign n18168 = ~n16657 & ~n16728 ;
  assign n18169 = ~\u0_w_reg[3][2]/P0001  & ~n16596 ;
  assign n18170 = n18168 & n18169 ;
  assign n18171 = ~n18167 & n18170 ;
  assign n18172 = \u0_w_reg[3][2]/P0001  & ~n16523 ;
  assign n18173 = ~n16530 & n18172 ;
  assign n18174 = ~n18171 & ~n18173 ;
  assign n18190 = ~n16597 & ~n16696 ;
  assign n18191 = ~n18174 & n18190 ;
  assign n18192 = ~n18189 & n18191 ;
  assign n18193 = \u0_w_reg[3][0]/P0001  & ~n18192 ;
  assign n18225 = \u0_w_reg[3][3]/P0001  & n17952 ;
  assign n18226 = ~\u0_w_reg[3][5]/P0001  & n16570 ;
  assign n18227 = ~n16522 & ~n17501 ;
  assign n18228 = ~n18226 & n18227 ;
  assign n18229 = n16667 & ~n18228 ;
  assign n18230 = ~n18225 & ~n18229 ;
  assign n18231 = \u0_w_reg[3][2]/P0001  & ~n18230 ;
  assign n18234 = ~n16549 & ~n16696 ;
  assign n18232 = n16588 & n16649 ;
  assign n18233 = n16509 & n16728 ;
  assign n18235 = ~n18232 & ~n18233 ;
  assign n18236 = n18234 & n18235 ;
  assign n18237 = ~n18231 & n18236 ;
  assign n18238 = ~\u0_w_reg[3][1]/P0001  & ~n18237 ;
  assign n18243 = \u0_w_reg[3][3]/P0001  & n16659 ;
  assign n18244 = ~n17935 & ~n18243 ;
  assign n18245 = \u0_w_reg[3][1]/P0001  & ~n18244 ;
  assign n18239 = ~n16543 & ~n16676 ;
  assign n18240 = ~\u0_w_reg[3][2]/P0001  & ~n18239 ;
  assign n18241 = \u0_w_reg[3][1]/P0001  & \u0_w_reg[3][2]/P0001  ;
  assign n18242 = n16485 & n18241 ;
  assign n18246 = n16506 & n18225 ;
  assign n18247 = ~n18242 & ~n18246 ;
  assign n18248 = ~n18240 & n18247 ;
  assign n18249 = ~n18245 & n18248 ;
  assign n18250 = ~n18238 & n18249 ;
  assign n18251 = ~n18193 & n18250 ;
  assign n18252 = ~n18224 & n18251 ;
  assign n18253 = \u0_w_reg[0][13]/P0001  & ~n18252 ;
  assign n18254 = ~\u0_w_reg[0][13]/P0001  & n18252 ;
  assign n18255 = ~n18253 & ~n18254 ;
  assign n18256 = \u0_w_reg[1][13]/P0001  & ~\u0_w_reg[2][13]/P0001  ;
  assign n18257 = ~\u0_w_reg[1][13]/P0001  & \u0_w_reg[2][13]/P0001  ;
  assign n18258 = ~n18256 & ~n18257 ;
  assign n18259 = n18255 & n18258 ;
  assign n18260 = ~n18255 & ~n18258 ;
  assign n18261 = ~n18259 & ~n18260 ;
  assign n18262 = ~ld_pad & n18261 ;
  assign n18263 = ~n18162 & ~n18262 ;
  assign n18265 = ~n16505 & ~n16522 ;
  assign n18266 = n17516 & ~n18265 ;
  assign n18264 = n16512 & n17566 ;
  assign n18267 = n17531 & ~n17897 ;
  assign n18268 = ~n18264 & n18267 ;
  assign n18269 = ~n18266 & n18268 ;
  assign n18271 = n16524 & n16582 ;
  assign n18270 = n16493 & n16506 ;
  assign n18272 = ~\u0_w_reg[3][1]/P0001  & ~n17958 ;
  assign n18273 = ~n18270 & n18272 ;
  assign n18274 = ~n18271 & n18273 ;
  assign n18275 = ~n18269 & ~n18274 ;
  assign n18282 = \u0_w_reg[3][4]/P0001  & n16587 ;
  assign n18278 = n16489 & n16603 ;
  assign n18283 = ~\u0_w_reg[3][0]/P0001  & ~n18278 ;
  assign n18284 = ~n18233 & n18283 ;
  assign n18285 = ~n18282 & n18284 ;
  assign n18279 = n16495 & n16528 ;
  assign n18280 = ~n16659 & ~n18279 ;
  assign n18281 = n16524 & ~n18280 ;
  assign n18276 = ~n16596 & ~n17501 ;
  assign n18277 = n16588 & ~n18276 ;
  assign n18286 = ~n18246 & ~n18277 ;
  assign n18287 = ~n18281 & n18286 ;
  assign n18288 = n18285 & n18287 ;
  assign n18289 = ~n18275 & n18288 ;
  assign n18290 = \u0_w_reg[3][2]/P0001  & ~n16504 ;
  assign n18291 = ~\u0_w_reg[3][2]/P0001  & ~n16608 ;
  assign n18292 = ~n16687 & ~n17961 ;
  assign n18293 = n18291 & n18292 ;
  assign n18294 = ~n18290 & ~n18293 ;
  assign n18295 = ~\u0_w_reg[3][3]/P0001  & n16483 ;
  assign n18296 = ~n16552 & n18295 ;
  assign n18297 = ~n16729 & n18181 ;
  assign n18298 = ~n18296 & n18297 ;
  assign n18299 = ~n18294 & n18298 ;
  assign n18301 = ~n16477 & ~n16608 ;
  assign n18300 = \u0_w_reg[3][3]/P0001  & n16483 ;
  assign n18302 = ~n16622 & ~n18300 ;
  assign n18303 = n18301 & n18302 ;
  assign n18304 = \u0_w_reg[3][2]/P0001  & ~n18303 ;
  assign n18306 = n16496 & n16521 ;
  assign n18305 = n16588 & n18226 ;
  assign n18307 = \u0_w_reg[3][1]/P0001  & ~n18305 ;
  assign n18308 = ~n18306 & n18307 ;
  assign n18309 = ~n18304 & n18308 ;
  assign n18310 = ~n18299 & ~n18309 ;
  assign n18317 = \u0_w_reg[3][5]/P0001  & n16668 ;
  assign n18313 = n16524 & n16700 ;
  assign n18318 = \u0_w_reg[3][0]/P0001  & ~n18313 ;
  assign n18319 = ~n18317 & n18318 ;
  assign n18311 = ~n16550 & ~n16589 ;
  assign n18312 = \u0_w_reg[3][4]/P0001  & ~n18311 ;
  assign n18314 = ~\u0_w_reg[3][4]/P0001  & n16541 ;
  assign n18315 = ~n17952 & ~n18314 ;
  assign n18316 = n16512 & ~n18315 ;
  assign n18320 = ~n18312 & ~n18316 ;
  assign n18321 = n18319 & n18320 ;
  assign n18322 = ~n18310 & n18321 ;
  assign n18323 = ~n18289 & ~n18322 ;
  assign n18330 = ~n16575 & ~n16697 ;
  assign n18331 = ~n18314 & n18330 ;
  assign n18332 = ~\u0_w_reg[3][3]/P0001  & ~n18331 ;
  assign n18333 = \u0_w_reg[3][2]/P0001  & ~n16627 ;
  assign n18334 = ~n16728 & n18333 ;
  assign n18335 = ~n18332 & n18334 ;
  assign n18324 = n16521 & n16658 ;
  assign n18325 = ~n16478 & ~n18324 ;
  assign n18326 = n16488 & ~n16489 ;
  assign n18327 = n18325 & ~n18326 ;
  assign n18328 = \u0_w_reg[3][3]/P0001  & ~n18327 ;
  assign n18329 = ~\u0_w_reg[3][2]/P0001  & ~n18328 ;
  assign n18336 = \u0_w_reg[3][1]/P0001  & ~n18329 ;
  assign n18337 = ~n18335 & n18336 ;
  assign n18338 = ~\u0_w_reg[3][2]/P0001  & n17907 ;
  assign n18339 = ~n16529 & ~n18277 ;
  assign n18340 = ~n18338 & n18339 ;
  assign n18341 = ~\u0_w_reg[3][1]/P0001  & ~n18340 ;
  assign n18346 = ~n16701 & ~n18306 ;
  assign n18347 = n16621 & ~n18346 ;
  assign n18342 = n17516 & n17927 ;
  assign n18343 = n16621 & n16687 ;
  assign n18344 = ~n17970 & ~n18343 ;
  assign n18345 = ~\u0_w_reg[3][3]/P0001  & ~n18344 ;
  assign n18348 = ~n18342 & ~n18345 ;
  assign n18349 = ~n18347 & n18348 ;
  assign n18350 = ~n18341 & n18349 ;
  assign n18351 = ~n18337 & n18350 ;
  assign n18352 = ~n18323 & n18351 ;
  assign n18353 = \u0_w_reg[0][15]/P0001  & ~n18352 ;
  assign n18354 = ~\u0_w_reg[0][15]/P0001  & n18352 ;
  assign n18355 = ~n18353 & ~n18354 ;
  assign n18356 = \u0_w_reg[1][15]/P0001  & n18355 ;
  assign n18357 = ~\u0_w_reg[1][15]/P0001  & ~n18355 ;
  assign n18358 = ~n18356 & ~n18357 ;
  assign n18359 = \u0_w_reg[2][15]/P0001  & n18358 ;
  assign n18360 = ~\u0_w_reg[2][15]/P0001  & ~n18358 ;
  assign n18361 = ~n18359 & ~n18360 ;
  assign n18362 = ~ld_pad & n18361 ;
  assign n18363 = \key[47]_pad  & ld_pad ;
  assign n18364 = ~n18362 & ~n18363 ;
  assign n18365 = ~\key[40]_pad  & ld_pad ;
  assign n18391 = ~\u0_w_reg[3][3]/P0001  & ~n18325 ;
  assign n18392 = n16526 & ~n16544 ;
  assign n18390 = ~\u0_w_reg[3][2]/P0001  & n16650 ;
  assign n18393 = ~\u0_w_reg[3][1]/P0001  & ~n18390 ;
  assign n18394 = ~n18392 & n18393 ;
  assign n18395 = ~n18391 & n18394 ;
  assign n18396 = \u0_w_reg[3][4]/P0001  & n16541 ;
  assign n18397 = ~n16550 & ~n18396 ;
  assign n18398 = \u0_w_reg[3][3]/P0001  & ~n18397 ;
  assign n18400 = \u0_w_reg[3][1]/P0001  & ~n16622 ;
  assign n18399 = n16574 & n16588 ;
  assign n18401 = ~n17519 & ~n18399 ;
  assign n18402 = n18400 & n18401 ;
  assign n18403 = ~n18398 & n18402 ;
  assign n18404 = ~n18395 & ~n18403 ;
  assign n18386 = n16567 & ~n17896 ;
  assign n18387 = ~\u0_w_reg[3][2]/P0001  & ~n18386 ;
  assign n18388 = ~n16521 & ~n16753 ;
  assign n18389 = n16664 & ~n18388 ;
  assign n18405 = ~\u0_w_reg[3][0]/P0001  & ~n18389 ;
  assign n18406 = ~n18387 & n18405 ;
  assign n18407 = ~n18404 & n18406 ;
  assign n18417 = ~n16550 & ~n18305 ;
  assign n18418 = \u0_w_reg[3][4]/P0001  & ~n18417 ;
  assign n18415 = ~n16622 & ~n18396 ;
  assign n18416 = n16689 & ~n18415 ;
  assign n18419 = ~\u0_w_reg[3][1]/P0001  & ~n16743 ;
  assign n18420 = ~n17505 & ~n18175 ;
  assign n18421 = n18419 & n18420 ;
  assign n18422 = ~n18416 & n18421 ;
  assign n18423 = ~n18418 & n18422 ;
  assign n18424 = \u0_w_reg[3][1]/P0001  & ~n16587 ;
  assign n18425 = ~n17969 & n18424 ;
  assign n18426 = ~n16573 & n18425 ;
  assign n18427 = ~n18423 & ~n18426 ;
  assign n18408 = ~n16675 & ~n18279 ;
  assign n18409 = n17534 & n18408 ;
  assign n18410 = ~n18317 & n18409 ;
  assign n18411 = \u0_w_reg[3][2]/P0001  & ~n16705 ;
  assign n18412 = ~n17958 & n18411 ;
  assign n18413 = n18176 & n18412 ;
  assign n18414 = ~n18410 & ~n18413 ;
  assign n18428 = \u0_w_reg[3][0]/P0001  & ~n16484 ;
  assign n18429 = ~n16744 & n18428 ;
  assign n18430 = ~n18414 & n18429 ;
  assign n18431 = ~n18427 & n18430 ;
  assign n18432 = ~n18407 & ~n18431 ;
  assign n18366 = ~\u0_w_reg[3][3]/P0001  & n17517 ;
  assign n18367 = ~n16494 & ~n18215 ;
  assign n18368 = ~n18366 & n18367 ;
  assign n18369 = \u0_w_reg[3][2]/P0001  & ~n18368 ;
  assign n18371 = \u0_w_reg[3][1]/P0001  & ~n16660 ;
  assign n18370 = ~\u0_w_reg[3][2]/P0001  & n16529 ;
  assign n18372 = ~n16676 & ~n18370 ;
  assign n18373 = n18371 & n18372 ;
  assign n18374 = ~n18369 & n18373 ;
  assign n18375 = ~n16556 & ~n17959 ;
  assign n18376 = n16731 & n18375 ;
  assign n18377 = ~n16522 & ~n17961 ;
  assign n18378 = ~\u0_w_reg[3][3]/P0001  & ~n18377 ;
  assign n18379 = ~\u0_w_reg[3][2]/P0001  & ~n17506 ;
  assign n18380 = ~n18378 & n18379 ;
  assign n18381 = ~n18376 & ~n18380 ;
  assign n18382 = ~\u0_w_reg[3][1]/P0001  & ~n17518 ;
  assign n18383 = ~n18381 & n18382 ;
  assign n18384 = ~n18374 & ~n18383 ;
  assign n18385 = n16509 & n17532 ;
  assign n18433 = ~n18384 & ~n18385 ;
  assign n18434 = ~n18432 & n18433 ;
  assign n18435 = \u0_w_reg[0][8]/P0001  & ~n18434 ;
  assign n18436 = ~\u0_w_reg[0][8]/P0001  & n18434 ;
  assign n18437 = ~n18435 & ~n18436 ;
  assign n18438 = \u0_w_reg[1][8]/P0001  & ~\u0_w_reg[2][8]/P0001  ;
  assign n18439 = ~\u0_w_reg[1][8]/P0001  & \u0_w_reg[2][8]/P0001  ;
  assign n18440 = ~n18438 & ~n18439 ;
  assign n18441 = n18437 & n18440 ;
  assign n18442 = ~n18437 & ~n18440 ;
  assign n18443 = ~n18441 & ~n18442 ;
  assign n18444 = ~ld_pad & n18443 ;
  assign n18445 = ~n18365 & ~n18444 ;
  assign n18474 = ~\u0_w_reg[3][19]/P0001  & n15606 ;
  assign n18475 = ~n15615 & ~n18474 ;
  assign n18476 = \u0_w_reg[3][18]/P0001  & ~n18475 ;
  assign n18470 = \u0_w_reg[3][19]/P0001  & n16840 ;
  assign n18471 = ~n15550 & ~n16875 ;
  assign n18472 = ~n18470 & n18471 ;
  assign n18473 = ~\u0_w_reg[3][18]/P0001  & ~n18472 ;
  assign n18477 = \u0_w_reg[3][17]/P0001  & ~n15584 ;
  assign n18478 = n15541 & n18477 ;
  assign n18479 = ~n18473 & n18478 ;
  assign n18480 = ~n18476 & n18479 ;
  assign n18482 = n15660 & n17090 ;
  assign n18481 = ~\u0_w_reg[3][20]/P0001  & n16242 ;
  assign n18485 = ~n17018 & ~n18481 ;
  assign n18486 = ~n18482 & n18485 ;
  assign n18483 = ~\u0_w_reg[3][17]/P0001  & ~n16276 ;
  assign n18484 = ~n16288 & ~n16909 ;
  assign n18487 = n18483 & n18484 ;
  assign n18488 = n18486 & n18487 ;
  assign n18489 = ~n18480 & ~n18488 ;
  assign n18490 = n15529 & n16313 ;
  assign n18493 = ~n15637 & ~n15656 ;
  assign n18494 = ~n18490 & n18493 ;
  assign n18491 = ~n15557 & ~n15613 ;
  assign n18492 = n15511 & ~n18491 ;
  assign n18495 = ~n16240 & ~n18492 ;
  assign n18496 = n18494 & n18495 ;
  assign n18497 = ~n18489 & n18496 ;
  assign n18498 = ~\u0_w_reg[3][16]/P0001  & ~n18497 ;
  assign n18447 = \u0_w_reg[3][19]/P0001  & n15590 ;
  assign n18448 = ~n16840 & ~n17110 ;
  assign n18449 = ~n18447 & n18448 ;
  assign n18450 = \u0_w_reg[3][18]/P0001  & ~n18449 ;
  assign n18451 = n16874 & ~n18450 ;
  assign n18452 = \u0_w_reg[3][17]/P0001  & ~n18451 ;
  assign n18455 = ~n15530 & ~n15542 ;
  assign n18456 = n15521 & ~n18455 ;
  assign n18453 = n15529 & n15530 ;
  assign n18454 = n15560 & n16268 ;
  assign n18457 = ~n18453 & ~n18454 ;
  assign n18458 = ~n18456 & n18457 ;
  assign n18459 = ~\u0_w_reg[3][17]/P0001  & ~n18458 ;
  assign n18460 = ~n16814 & ~n16944 ;
  assign n18461 = ~\u0_w_reg[3][18]/P0001  & ~n18460 ;
  assign n18462 = n16283 & ~n16901 ;
  assign n18446 = ~n15588 & n15592 ;
  assign n18463 = ~n15608 & n15655 ;
  assign n18464 = ~n18446 & ~n18463 ;
  assign n18465 = ~n18462 & n18464 ;
  assign n18466 = ~n18461 & n18465 ;
  assign n18467 = ~n18459 & n18466 ;
  assign n18468 = ~n18452 & n18467 ;
  assign n18469 = \u0_w_reg[3][16]/P0001  & ~n18468 ;
  assign n18513 = ~n15558 & ~n17059 ;
  assign n18514 = ~n16802 & n18513 ;
  assign n18515 = ~\u0_w_reg[3][18]/P0001  & ~n18514 ;
  assign n18516 = ~n15563 & ~n16222 ;
  assign n18517 = ~n18515 & n18516 ;
  assign n18518 = ~\u0_w_reg[3][17]/P0001  & ~n18517 ;
  assign n18508 = ~n15560 & ~n15630 ;
  assign n18509 = ~n15544 & ~n18508 ;
  assign n18510 = ~n15584 & ~n16851 ;
  assign n18511 = ~n18509 & n18510 ;
  assign n18512 = n16910 & ~n18511 ;
  assign n18499 = ~n15513 & ~n15625 ;
  assign n18500 = \u0_w_reg[3][19]/P0001  & ~n18499 ;
  assign n18501 = ~n17032 & ~n18500 ;
  assign n18502 = n16901 & ~n18501 ;
  assign n18503 = ~n15603 & ~n15630 ;
  assign n18504 = n15608 & ~n18503 ;
  assign n18505 = ~n15531 & ~n15620 ;
  assign n18506 = ~n15514 & n18505 ;
  assign n18507 = n16282 & ~n18506 ;
  assign n18519 = ~n18504 & ~n18507 ;
  assign n18520 = ~n18502 & n18519 ;
  assign n18521 = ~n18512 & n18520 ;
  assign n18522 = ~n18518 & n18521 ;
  assign n18523 = ~n18469 & n18522 ;
  assign n18524 = ~n18498 & n18523 ;
  assign n18525 = \u0_w_reg[0][25]/P0001  & ~n18524 ;
  assign n18526 = ~\u0_w_reg[0][25]/P0001  & n18524 ;
  assign n18527 = ~n18525 & ~n18526 ;
  assign n18529 = \u0_r0_out_reg[25]/P0001  & n18527 ;
  assign n18528 = ~\u0_r0_out_reg[25]/P0001  & ~n18527 ;
  assign n18530 = ~ld_pad & ~n18528 ;
  assign n18531 = ~n18529 & n18530 ;
  assign n18532 = \key[121]_pad  & ld_pad ;
  assign n18533 = ~n18531 & ~n18532 ;
  assign n18534 = \u0_r0_out_reg[25]/P0001  & ~\u0_w_reg[1][25]/P0001  ;
  assign n18535 = ~\u0_r0_out_reg[25]/P0001  & \u0_w_reg[1][25]/P0001  ;
  assign n18536 = ~n18534 & ~n18535 ;
  assign n18538 = n18527 & ~n18536 ;
  assign n18537 = ~n18527 & n18536 ;
  assign n18539 = ~ld_pad & ~n18537 ;
  assign n18540 = ~n18538 & n18539 ;
  assign n18541 = \key[89]_pad  & ld_pad ;
  assign n18542 = ~n18540 & ~n18541 ;
  assign n18543 = ~\key[57]_pad  & ld_pad ;
  assign n18544 = \u0_w_reg[2][25]/P0001  & n18536 ;
  assign n18545 = ~\u0_w_reg[2][25]/P0001  & ~n18536 ;
  assign n18546 = ~n18544 & ~n18545 ;
  assign n18547 = n18527 & n18546 ;
  assign n18548 = ~n18527 & ~n18546 ;
  assign n18549 = ~n18547 & ~n18548 ;
  assign n18550 = ~ld_pad & n18549 ;
  assign n18551 = ~n18543 & ~n18550 ;
  assign n18553 = \u0_w_reg[3][25]/P0001  & ~n18549 ;
  assign n18552 = ~\u0_w_reg[3][25]/P0001  & n18549 ;
  assign n18554 = ~ld_pad & ~n18552 ;
  assign n18555 = ~n18553 & n18554 ;
  assign n18556 = \key[25]_pad  & ld_pad ;
  assign n18557 = ~n18555 & ~n18556 ;
  assign n18558 = ~\u0_w_reg[3][15]/P0001  & n17644 ;
  assign n18559 = ~n15754 & ~n18558 ;
  assign n18560 = ~\u0_w_reg[3][10]/P0001  & ~n18559 ;
  assign n18561 = ~n17684 & ~n17771 ;
  assign n18562 = ~n18017 & n18561 ;
  assign n18563 = ~n18560 & n18562 ;
  assign n18564 = \u0_w_reg[3][9]/P0001  & ~n18563 ;
  assign n18571 = \u0_w_reg[3][10]/P0001  & n17731 ;
  assign n18575 = ~\u0_w_reg[3][8]/P0001  & ~n15980 ;
  assign n18576 = ~n15861 & n18575 ;
  assign n18572 = ~n15757 & n15847 ;
  assign n18573 = n17631 & n18572 ;
  assign n18574 = n15803 & n15865 ;
  assign n18577 = ~n18573 & ~n18574 ;
  assign n18578 = n18576 & n18577 ;
  assign n18579 = ~n18571 & n18578 ;
  assign n18565 = n15799 & n15946 ;
  assign n18566 = ~n15804 & ~n17638 ;
  assign n18567 = ~n18565 & n18566 ;
  assign n18568 = ~\u0_w_reg[3][9]/P0001  & ~n18567 ;
  assign n18569 = ~n15758 & ~n17722 ;
  assign n18570 = ~\u0_w_reg[3][10]/P0001  & ~n18569 ;
  assign n18580 = ~n18568 & ~n18570 ;
  assign n18581 = n18579 & n18580 ;
  assign n18582 = ~n18564 & n18581 ;
  assign n18583 = ~n15787 & n17651 ;
  assign n18584 = ~n15942 & ~n18583 ;
  assign n18585 = \u0_w_reg[3][12]/P0001  & ~n18584 ;
  assign n18588 = n15725 & n15847 ;
  assign n18589 = ~\u0_w_reg[3][9]/P0001  & ~n17682 ;
  assign n18590 = ~n18588 & n18589 ;
  assign n18586 = ~\u0_w_reg[3][10]/P0001  & n15741 ;
  assign n18587 = n15803 & n15896 ;
  assign n18591 = ~n18586 & ~n18587 ;
  assign n18592 = n18590 & n18591 ;
  assign n18593 = ~n18585 & n18592 ;
  assign n18595 = ~n15716 & ~n15983 ;
  assign n18594 = \u0_w_reg[3][11]/P0001  & n15725 ;
  assign n18596 = ~n17609 & ~n18594 ;
  assign n18597 = n18595 & n18596 ;
  assign n18598 = \u0_w_reg[3][10]/P0001  & ~n18597 ;
  assign n18599 = \u0_w_reg[3][9]/P0001  & ~n17781 ;
  assign n18600 = ~\u0_w_reg[3][14]/P0001  & n17610 ;
  assign n18601 = n18599 & ~n18600 ;
  assign n18602 = ~n18598 & n18601 ;
  assign n18603 = ~n18593 & ~n18602 ;
  assign n18605 = \u0_w_reg[3][15]/P0001  & n15716 ;
  assign n18606 = ~n17737 & ~n18605 ;
  assign n18607 = n15893 & ~n18606 ;
  assign n18609 = \u0_w_reg[3][8]/P0001  & ~n17643 ;
  assign n18610 = ~n15792 & n18609 ;
  assign n18604 = \u0_w_reg[3][12]/P0001  & n18588 ;
  assign n18608 = n15738 & n15799 ;
  assign n18611 = ~n18604 & ~n18608 ;
  assign n18612 = n18610 & n18611 ;
  assign n18613 = ~n18607 & n18612 ;
  assign n18614 = ~n18603 & n18613 ;
  assign n18615 = ~n18582 & ~n18614 ;
  assign n18620 = ~n15802 & ~n17672 ;
  assign n18621 = ~n18605 & n18620 ;
  assign n18622 = ~\u0_w_reg[3][11]/P0001  & ~n18621 ;
  assign n18623 = \u0_w_reg[3][10]/P0001  & ~n15715 ;
  assign n18624 = ~n15815 & n18623 ;
  assign n18625 = ~n18622 & n18624 ;
  assign n18616 = ~n17598 & n17601 ;
  assign n18617 = \u0_w_reg[3][11]/P0001  & ~n18616 ;
  assign n18618 = ~\u0_w_reg[3][10]/P0001  & ~n15837 ;
  assign n18619 = ~n18617 & n18618 ;
  assign n18626 = \u0_w_reg[3][9]/P0001  & ~n18619 ;
  assign n18627 = ~n18625 & n18626 ;
  assign n18634 = ~\u0_w_reg[3][12]/P0001  & n15814 ;
  assign n18635 = n15849 & n18634 ;
  assign n18636 = ~n15941 & ~n18573 ;
  assign n18637 = ~n18635 & n18636 ;
  assign n18638 = ~\u0_w_reg[3][9]/P0001  & ~n18637 ;
  assign n18628 = n15735 & n15943 ;
  assign n18629 = ~n15785 & ~n18628 ;
  assign n18630 = ~\u0_w_reg[3][10]/P0001  & ~n18629 ;
  assign n18631 = ~n15789 & ~n15902 ;
  assign n18632 = ~n17781 & n18631 ;
  assign n18633 = n15974 & ~n18632 ;
  assign n18639 = ~n18630 & ~n18633 ;
  assign n18640 = ~n18638 & n18639 ;
  assign n18641 = ~n18627 & n18640 ;
  assign n18642 = ~n18615 & n18641 ;
  assign n18643 = \u0_w_reg[0][23]/P0001  & ~n18642 ;
  assign n18644 = ~\u0_w_reg[0][23]/P0001  & n18642 ;
  assign n18645 = ~n18643 & ~n18644 ;
  assign n18646 = \u0_w_reg[1][23]/P0001  & n18645 ;
  assign n18647 = ~\u0_w_reg[1][23]/P0001  & ~n18645 ;
  assign n18648 = ~n18646 & ~n18647 ;
  assign n18649 = \u0_w_reg[2][23]/P0001  & n18648 ;
  assign n18650 = ~\u0_w_reg[2][23]/P0001  & ~n18648 ;
  assign n18651 = ~n18649 & ~n18650 ;
  assign n18652 = ~ld_pad & n18651 ;
  assign n18653 = \key[55]_pad  & ld_pad ;
  assign n18654 = ~n18652 & ~n18653 ;
  assign n18655 = ~ld_pad & n16466 ;
  assign n18656 = \key[99]_pad  & ld_pad ;
  assign n18657 = ~n18655 & ~n18656 ;
  assign n18659 = \u0_w_reg[1][3]/P0001  & n16466 ;
  assign n18658 = ~\u0_w_reg[1][3]/P0001  & ~n16466 ;
  assign n18660 = ~ld_pad & ~n18658 ;
  assign n18661 = ~n18659 & n18660 ;
  assign n18662 = \key[67]_pad  & ld_pad ;
  assign n18663 = ~n18661 & ~n18662 ;
  assign n18665 = \u0_w_reg[3][3]/P0001  & ~n16472 ;
  assign n18664 = ~\u0_w_reg[3][3]/P0001  & n16472 ;
  assign n18666 = ~ld_pad & ~n18664 ;
  assign n18667 = ~n18665 & n18666 ;
  assign n18668 = \key[3]_pad  & ld_pad ;
  assign n18669 = ~n18667 & ~n18668 ;
  assign n18670 = ~ld_pad & n16639 ;
  assign n18671 = \key[107]_pad  & ld_pad ;
  assign n18672 = ~n18670 & ~n18671 ;
  assign n18674 = \u0_w_reg[1][11]/P0001  & n16639 ;
  assign n18673 = ~\u0_w_reg[1][11]/P0001  & ~n16639 ;
  assign n18675 = ~ld_pad & ~n18673 ;
  assign n18676 = ~n18674 & n18675 ;
  assign n18677 = \key[75]_pad  & ld_pad ;
  assign n18678 = ~n18676 & ~n18677 ;
  assign n18680 = \u0_w_reg[3][11]/P0001  & ~n16645 ;
  assign n18679 = ~\u0_w_reg[3][11]/P0001  & n16645 ;
  assign n18681 = ~ld_pad & ~n18679 ;
  assign n18682 = ~n18680 & n18681 ;
  assign n18683 = \key[11]_pad  & ld_pad ;
  assign n18684 = ~n18682 & ~n18683 ;
  assign n18685 = ~\key[49]_pad  & ld_pad ;
  assign n18735 = ~n17683 & ~n17772 ;
  assign n18736 = ~n18634 & n18735 ;
  assign n18737 = \u0_w_reg[3][10]/P0001  & ~n18736 ;
  assign n18738 = n17732 & ~n18737 ;
  assign n18739 = \u0_w_reg[3][9]/P0001  & ~n18738 ;
  assign n18749 = ~n15784 & ~n15976 ;
  assign n18750 = ~n17738 & ~n17771 ;
  assign n18751 = n18749 & n18750 ;
  assign n18752 = ~\u0_w_reg[3][10]/P0001  & ~n18751 ;
  assign n18740 = ~n15742 & ~n15859 ;
  assign n18741 = ~n15735 & ~n15849 ;
  assign n18742 = ~n15929 & n18741 ;
  assign n18743 = ~n18740 & ~n18742 ;
  assign n18744 = ~n15976 & ~n18743 ;
  assign n18745 = ~\u0_w_reg[3][9]/P0001  & ~n18744 ;
  assign n18746 = ~n15782 & n15787 ;
  assign n18747 = ~n17738 & ~n18746 ;
  assign n18748 = ~\u0_w_reg[3][11]/P0001  & ~n18747 ;
  assign n18753 = ~n18745 & ~n18748 ;
  assign n18754 = ~n18752 & n18753 ;
  assign n18755 = ~n18739 & n18754 ;
  assign n18756 = \u0_w_reg[3][8]/P0001  & ~n18755 ;
  assign n18686 = n15732 & ~n17759 ;
  assign n18687 = ~\u0_w_reg[3][11]/P0001  & n15742 ;
  assign n18688 = ~\u0_w_reg[3][10]/P0001  & ~n18687 ;
  assign n18689 = ~n18686 & n18688 ;
  assign n18690 = ~\u0_w_reg[3][11]/P0001  & n15840 ;
  assign n18691 = \u0_w_reg[3][10]/P0001  & ~n15821 ;
  assign n18692 = ~n18690 & n18691 ;
  assign n18693 = ~n18689 & ~n18692 ;
  assign n18694 = n15718 & n15790 ;
  assign n18695 = ~n18693 & n18694 ;
  assign n18700 = n15787 & n15799 ;
  assign n18701 = ~\u0_w_reg[3][9]/P0001  & ~n18700 ;
  assign n18702 = ~n17757 & n18701 ;
  assign n18696 = ~n15812 & ~n15846 ;
  assign n18697 = n15919 & ~n18696 ;
  assign n18698 = ~n15757 & ~n15896 ;
  assign n18699 = n15730 & ~n18698 ;
  assign n18703 = ~n18697 & ~n18699 ;
  assign n18704 = n18702 & n18703 ;
  assign n18705 = ~n18695 & ~n18704 ;
  assign n18708 = n15805 & n15849 ;
  assign n18709 = ~n15853 & ~n15861 ;
  assign n18710 = ~n18708 & n18709 ;
  assign n18706 = ~n15822 & ~n15943 ;
  assign n18707 = n15893 & ~n18706 ;
  assign n18711 = ~n15959 & ~n18707 ;
  assign n18712 = n18710 & n18711 ;
  assign n18713 = ~n18705 & n18712 ;
  assign n18714 = ~\u0_w_reg[3][8]/P0001  & ~n18713 ;
  assign n18729 = ~n15759 & ~n17638 ;
  assign n18730 = ~n18558 & n18729 ;
  assign n18731 = ~\u0_w_reg[3][10]/P0001  & ~n18730 ;
  assign n18732 = ~n15755 & ~n15932 ;
  assign n18733 = ~n18731 & n18732 ;
  assign n18734 = ~\u0_w_reg[3][9]/P0001  & ~n18733 ;
  assign n18726 = ~n15971 & ~n17721 ;
  assign n18727 = ~n18017 & n18726 ;
  assign n18728 = n18055 & ~n18727 ;
  assign n18720 = ~n15823 & ~n15929 ;
  assign n18721 = ~\u0_w_reg[3][14]/P0001  & ~n18720 ;
  assign n18722 = ~n15789 & ~n17667 ;
  assign n18723 = ~n17719 & n18722 ;
  assign n18724 = ~n18721 & n18723 ;
  assign n18725 = n15726 & ~n18724 ;
  assign n18715 = ~n15865 & ~n15960 ;
  assign n18716 = n15803 & ~n18715 ;
  assign n18717 = ~n15820 & ~n15839 ;
  assign n18718 = ~n15705 & n18717 ;
  assign n18719 = n15975 & ~n18718 ;
  assign n18757 = ~n18716 & ~n18719 ;
  assign n18758 = ~n18725 & n18757 ;
  assign n18759 = ~n18728 & n18758 ;
  assign n18760 = ~n18734 & n18759 ;
  assign n18761 = ~n18714 & n18760 ;
  assign n18762 = ~n18756 & n18761 ;
  assign n18763 = \u0_w_reg[0][17]/P0001  & ~n18762 ;
  assign n18764 = ~\u0_w_reg[0][17]/P0001  & n18762 ;
  assign n18765 = ~n18763 & ~n18764 ;
  assign n18766 = \u0_w_reg[1][17]/P0001  & ~\u0_w_reg[2][17]/P0001  ;
  assign n18767 = ~\u0_w_reg[1][17]/P0001  & \u0_w_reg[2][17]/P0001  ;
  assign n18768 = ~n18766 & ~n18767 ;
  assign n18769 = n18765 & n18768 ;
  assign n18770 = ~n18765 & ~n18768 ;
  assign n18771 = ~n18769 & ~n18770 ;
  assign n18772 = ~ld_pad & n18771 ;
  assign n18773 = ~n18685 & ~n18772 ;
  assign n18774 = ~\key[33]_pad  & ld_pad ;
  assign n18797 = \u0_w_reg[3][26]/P0001  & ~n16393 ;
  assign n18798 = ~n18082 & n18127 ;
  assign n18799 = ~n18797 & ~n18798 ;
  assign n18801 = ~\u0_w_reg[3][25]/P0001  & ~n16449 ;
  assign n18800 = n16033 & n16098 ;
  assign n18802 = ~n17824 & ~n18800 ;
  assign n18803 = n18801 & n18802 ;
  assign n18804 = ~n18799 & n18803 ;
  assign n18808 = \u0_w_reg[3][28]/P0001  & n17422 ;
  assign n18807 = ~\u0_w_reg[3][27]/P0001  & n16043 ;
  assign n18809 = ~n16121 & ~n18807 ;
  assign n18810 = ~n18808 & n18809 ;
  assign n18811 = ~\u0_w_reg[3][26]/P0001  & ~n18810 ;
  assign n18805 = ~n16129 & ~n18118 ;
  assign n18806 = \u0_w_reg[3][26]/P0001  & ~n18805 ;
  assign n18812 = \u0_w_reg[3][25]/P0001  & ~n16144 ;
  assign n18813 = n16016 & n18812 ;
  assign n18814 = ~n18806 & n18813 ;
  assign n18815 = ~n18811 & n18814 ;
  assign n18816 = ~n18804 & ~n18815 ;
  assign n18818 = ~n16039 & ~n16052 ;
  assign n18819 = n16036 & ~n18818 ;
  assign n18821 = ~n16088 & ~n16104 ;
  assign n18817 = n16091 & n16386 ;
  assign n18820 = n16117 & n16428 ;
  assign n18822 = ~n18817 & ~n18820 ;
  assign n18823 = n18821 & n18822 ;
  assign n18824 = ~n18819 & n18823 ;
  assign n18825 = ~n18816 & n18824 ;
  assign n18826 = ~\u0_w_reg[3][24]/P0001  & ~n18825 ;
  assign n18775 = ~n16160 & ~n17277 ;
  assign n18776 = ~n17835 & n18775 ;
  assign n18777 = \u0_w_reg[3][26]/P0001  & ~n18776 ;
  assign n18778 = n17853 & ~n18777 ;
  assign n18779 = \u0_w_reg[3][25]/P0001  & ~n18778 ;
  assign n18789 = ~n16040 & ~n17331 ;
  assign n18790 = ~n17428 & ~n17820 ;
  assign n18791 = n18789 & n18790 ;
  assign n18792 = ~\u0_w_reg[3][26]/P0001  & ~n18791 ;
  assign n18780 = ~n16043 & ~n16102 ;
  assign n18781 = ~n16045 & ~n16117 ;
  assign n18782 = ~n16112 & n18781 ;
  assign n18783 = ~n18780 & ~n18782 ;
  assign n18784 = ~n16040 & ~n18783 ;
  assign n18785 = ~\u0_w_reg[3][25]/P0001  & ~n18784 ;
  assign n18786 = n16099 & ~n16147 ;
  assign n18787 = ~n17820 & ~n18786 ;
  assign n18788 = ~\u0_w_reg[3][27]/P0001  & ~n18787 ;
  assign n18793 = ~n18785 & ~n18788 ;
  assign n18794 = ~n18792 & n18793 ;
  assign n18795 = ~n18779 & n18794 ;
  assign n18796 = \u0_w_reg[3][24]/P0001  & ~n18795 ;
  assign n18839 = ~n16053 & ~n17328 ;
  assign n18840 = ~n17337 & n18839 ;
  assign n18841 = ~\u0_w_reg[3][26]/P0001  & ~n18840 ;
  assign n18842 = ~n16047 & ~n16376 ;
  assign n18843 = ~n18841 & n18842 ;
  assign n18844 = ~\u0_w_reg[3][25]/P0001  & ~n18843 ;
  assign n18828 = ~\u0_w_reg[3][31]/P0001  & n17866 ;
  assign n18827 = ~n16020 & n17805 ;
  assign n18829 = ~n16027 & ~n18827 ;
  assign n18830 = ~n18828 & n18829 ;
  assign n18831 = n16029 & ~n18830 ;
  assign n18835 = ~n16059 & ~n16163 ;
  assign n18836 = ~n16038 & n18835 ;
  assign n18837 = ~\u0_w_reg[3][25]/P0001  & n16036 ;
  assign n18838 = ~n18836 & n18837 ;
  assign n18832 = n16099 & n16411 ;
  assign n18833 = ~n16110 & ~n18832 ;
  assign n18834 = n17871 & ~n18833 ;
  assign n18845 = ~n16454 & ~n17344 ;
  assign n18846 = ~n18834 & n18845 ;
  assign n18847 = ~n18838 & n18846 ;
  assign n18848 = ~n18831 & n18847 ;
  assign n18849 = ~n18844 & n18848 ;
  assign n18850 = ~n18796 & n18849 ;
  assign n18851 = ~n18826 & n18850 ;
  assign n18852 = \u0_w_reg[0][1]/P0001  & ~n18851 ;
  assign n18853 = ~\u0_w_reg[0][1]/P0001  & n18851 ;
  assign n18854 = ~n18852 & ~n18853 ;
  assign n18855 = \u0_w_reg[1][1]/P0001  & ~\u0_w_reg[2][1]/P0001  ;
  assign n18856 = ~\u0_w_reg[1][1]/P0001  & \u0_w_reg[2][1]/P0001  ;
  assign n18857 = ~n18855 & ~n18856 ;
  assign n18858 = n18854 & n18857 ;
  assign n18859 = ~n18854 & ~n18857 ;
  assign n18860 = ~n18858 & ~n18859 ;
  assign n18861 = ~ld_pad & n18860 ;
  assign n18862 = ~n18774 & ~n18861 ;
  assign n18863 = ~\key[41]_pad  & ld_pad ;
  assign n18887 = n16588 & n16627 ;
  assign n18889 = ~n16723 & ~n17496 ;
  assign n18890 = ~n18887 & n18889 ;
  assign n18886 = ~n16512 & n16573 ;
  assign n18888 = ~\u0_w_reg[3][1]/P0001  & ~n16616 ;
  assign n18891 = ~n18886 & n18888 ;
  assign n18892 = n18890 & n18891 ;
  assign n18893 = ~\u0_w_reg[3][3]/P0001  & n16570 ;
  assign n18894 = ~n16580 & n16653 ;
  assign n18895 = ~n18893 & ~n18894 ;
  assign n18896 = ~\u0_w_reg[3][2]/P0001  & ~n18895 ;
  assign n18897 = n16482 & n16541 ;
  assign n18898 = ~n17915 & ~n18897 ;
  assign n18899 = \u0_w_reg[3][2]/P0001  & ~n18898 ;
  assign n18900 = \u0_w_reg[3][1]/P0001  & ~n16701 ;
  assign n18901 = n18168 & n18900 ;
  assign n18902 = ~n18899 & n18901 ;
  assign n18903 = ~n18896 & n18902 ;
  assign n18904 = ~n18892 & ~n18903 ;
  assign n18906 = \u0_w_reg[3][2]/P0001  & ~n17959 ;
  assign n18907 = ~n16724 & ~n18906 ;
  assign n18905 = ~\u0_w_reg[3][3]/P0001  & n17935 ;
  assign n18908 = ~n16506 & ~n16548 ;
  assign n18909 = n16520 & ~n18908 ;
  assign n18910 = ~n18210 & ~n18909 ;
  assign n18911 = ~n18905 & n18910 ;
  assign n18912 = ~n18907 & n18911 ;
  assign n18913 = ~n18904 & n18912 ;
  assign n18914 = ~\u0_w_reg[3][0]/P0001  & ~n18913 ;
  assign n18864 = ~n16503 & ~n17532 ;
  assign n18865 = ~n17566 & n18864 ;
  assign n18866 = \u0_w_reg[3][2]/P0001  & ~n18865 ;
  assign n18867 = n17572 & ~n18866 ;
  assign n18868 = \u0_w_reg[3][1]/P0001  & ~n18867 ;
  assign n18877 = ~n16532 & ~n17908 ;
  assign n18878 = \u0_w_reg[3][5]/P0001  & ~n18877 ;
  assign n18876 = ~n16552 & n18194 ;
  assign n18879 = ~n18324 & ~n18876 ;
  assign n18880 = ~n18878 & n18879 ;
  assign n18881 = ~\u0_w_reg[3][1]/P0001  & ~n18880 ;
  assign n18869 = n16542 & ~n16554 ;
  assign n18870 = ~n17500 & ~n18869 ;
  assign n18871 = ~\u0_w_reg[3][3]/P0001  & ~n18870 ;
  assign n18872 = ~n16484 & ~n17500 ;
  assign n18873 = ~n17530 & ~n18324 ;
  assign n18874 = n18872 & n18873 ;
  assign n18875 = ~\u0_w_reg[3][2]/P0001  & ~n18874 ;
  assign n18882 = ~n18871 & ~n18875 ;
  assign n18883 = ~n18881 & n18882 ;
  assign n18884 = ~n18868 & n18883 ;
  assign n18885 = \u0_w_reg[3][0]/P0001  & ~n18884 ;
  assign n18915 = ~n16545 & ~n17958 ;
  assign n18916 = ~n16624 & n18915 ;
  assign n18917 = ~\u0_w_reg[3][2]/P0001  & ~n18916 ;
  assign n18918 = ~n16732 & ~n17959 ;
  assign n18919 = ~n18917 & n18918 ;
  assign n18920 = ~\u0_w_reg[3][1]/P0001  & ~n18919 ;
  assign n18930 = ~n16481 & ~n16482 ;
  assign n18931 = ~\u0_w_reg[3][6]/P0001  & ~n16528 ;
  assign n18932 = ~n18930 & n18931 ;
  assign n18933 = ~\u0_w_reg[3][2]/P0001  & ~n16701 ;
  assign n18934 = ~n17517 & n18933 ;
  assign n18935 = ~n18932 & n18934 ;
  assign n18927 = ~n16627 & ~n16687 ;
  assign n18928 = \u0_w_reg[3][3]/P0001  & ~n18927 ;
  assign n18929 = n17898 & ~n18928 ;
  assign n18936 = \u0_w_reg[3][1]/P0001  & ~n18929 ;
  assign n18937 = ~n18935 & n18936 ;
  assign n18921 = ~n16525 & ~n18271 ;
  assign n18922 = ~\u0_w_reg[3][6]/P0001  & ~n18921 ;
  assign n18923 = ~n17519 & ~n18226 ;
  assign n18924 = ~n18279 & n18923 ;
  assign n18925 = ~\u0_w_reg[3][3]/P0001  & n16621 ;
  assign n18926 = ~n18924 & n18925 ;
  assign n18938 = ~n18922 & ~n18926 ;
  assign n18939 = ~n18937 & n18938 ;
  assign n18940 = ~n18920 & n18939 ;
  assign n18941 = ~n18885 & n18940 ;
  assign n18942 = ~n18914 & n18941 ;
  assign n18943 = \u0_w_reg[0][9]/P0001  & ~n18942 ;
  assign n18944 = ~\u0_w_reg[0][9]/P0001  & n18942 ;
  assign n18945 = ~n18943 & ~n18944 ;
  assign n18946 = \u0_w_reg[1][9]/P0001  & ~\u0_w_reg[2][9]/P0001  ;
  assign n18947 = ~\u0_w_reg[1][9]/P0001  & \u0_w_reg[2][9]/P0001  ;
  assign n18948 = ~n18946 & ~n18947 ;
  assign n18949 = n18945 & n18948 ;
  assign n18950 = ~n18945 & ~n18948 ;
  assign n18951 = ~n18949 & ~n18950 ;
  assign n18952 = ~ld_pad & n18951 ;
  assign n18953 = ~n18863 & ~n18952 ;
  assign n18954 = ~ld_pad & n16764 ;
  assign n18955 = \key[108]_pad  & ld_pad ;
  assign n18956 = ~n18954 & ~n18955 ;
  assign n18958 = \u0_w_reg[1][12]/P0001  & n16764 ;
  assign n18957 = ~\u0_w_reg[1][12]/P0001  & ~n16764 ;
  assign n18959 = ~ld_pad & ~n18957 ;
  assign n18960 = ~n18958 & n18959 ;
  assign n18961 = \key[76]_pad  & ld_pad ;
  assign n18962 = ~n18960 & ~n18961 ;
  assign n18971 = ~n15771 & ~n15802 ;
  assign n18972 = ~\u0_w_reg[3][10]/P0001  & ~n18971 ;
  assign n18973 = ~n15863 & ~n17742 ;
  assign n18974 = n15760 & n18973 ;
  assign n18975 = ~n18972 & n18974 ;
  assign n18976 = ~n15737 & ~n15846 ;
  assign n18977 = ~\u0_w_reg[3][10]/P0001  & ~n18976 ;
  assign n18978 = ~n15781 & n17746 ;
  assign n18979 = ~n18977 & n18978 ;
  assign n18980 = ~n18975 & ~n18979 ;
  assign n18967 = ~\u0_w_reg[3][15]/P0001  & n15751 ;
  assign n18968 = ~n15805 & ~n15862 ;
  assign n18969 = ~n18967 & n18968 ;
  assign n18970 = \u0_w_reg[3][10]/P0001  & ~n18969 ;
  assign n18963 = ~n15717 & ~n15939 ;
  assign n18964 = ~n18051 & n18963 ;
  assign n18965 = ~\u0_w_reg[3][10]/P0001  & ~n18964 ;
  assign n18966 = n15817 & n15974 ;
  assign n18981 = \u0_w_reg[3][8]/P0001  & ~n17681 ;
  assign n18982 = ~n18966 & n18981 ;
  assign n18983 = ~n18965 & n18982 ;
  assign n18984 = ~n18970 & n18983 ;
  assign n18985 = ~n18980 & n18984 ;
  assign n18986 = \u0_w_reg[3][13]/P0001  & ~n15724 ;
  assign n18987 = n15742 & n18986 ;
  assign n18988 = ~n15989 & ~n18987 ;
  assign n18989 = ~\u0_w_reg[3][10]/P0001  & ~n18988 ;
  assign n18990 = n15893 & n15946 ;
  assign n18991 = \u0_w_reg[3][9]/P0001  & ~n15920 ;
  assign n18992 = ~n17611 & n18991 ;
  assign n18993 = ~n18990 & n18992 ;
  assign n18994 = ~n18989 & n18993 ;
  assign n18997 = ~\u0_w_reg[3][9]/P0001  & ~n15804 ;
  assign n18998 = ~n15865 & n18997 ;
  assign n18995 = n15741 & n15847 ;
  assign n18996 = \u0_w_reg[3][12]/P0001  & n15791 ;
  assign n18999 = ~n18995 & ~n18996 ;
  assign n19000 = n18998 & n18999 ;
  assign n19001 = ~n18994 & ~n19000 ;
  assign n19004 = ~n15710 & ~n18628 ;
  assign n19005 = \u0_w_reg[3][10]/P0001  & ~n19004 ;
  assign n19002 = ~n15731 & ~n17672 ;
  assign n19003 = ~\u0_w_reg[3][11]/P0001  & ~n19002 ;
  assign n19006 = ~\u0_w_reg[3][8]/P0001  & ~n19003 ;
  assign n19007 = ~n19005 & n19006 ;
  assign n19008 = ~n19001 & n19007 ;
  assign n19009 = ~n18985 & ~n19008 ;
  assign n19010 = ~\u0_w_reg[3][10]/P0001  & n15976 ;
  assign n19011 = ~n18996 & ~n19010 ;
  assign n19012 = \u0_w_reg[3][11]/P0001  & ~n19011 ;
  assign n19013 = n15756 & ~n15907 ;
  assign n19014 = ~n15715 & ~n17682 ;
  assign n19015 = ~n17719 & n19014 ;
  assign n19016 = ~n19013 & n19015 ;
  assign n19017 = \u0_w_reg[3][10]/P0001  & ~n19016 ;
  assign n19020 = ~\u0_w_reg[3][9]/P0001  & ~n17722 ;
  assign n19018 = n15708 & ~n15822 ;
  assign n19019 = n15847 & n19018 ;
  assign n19021 = ~n17758 & ~n18708 ;
  assign n19022 = ~n19019 & n19021 ;
  assign n19023 = n19020 & n19022 ;
  assign n19024 = ~n19017 & n19023 ;
  assign n19029 = ~n17656 & ~n18026 ;
  assign n19027 = \u0_w_reg[3][12]/P0001  & n17743 ;
  assign n19028 = n15849 & n17650 ;
  assign n19030 = ~n19027 & ~n19028 ;
  assign n19031 = n19029 & n19030 ;
  assign n19025 = ~n15805 & ~n15832 ;
  assign n19026 = n15847 & ~n19025 ;
  assign n19032 = n18599 & ~n19026 ;
  assign n19033 = n19031 & n19032 ;
  assign n19034 = ~n19024 & ~n19033 ;
  assign n19035 = ~n19012 & ~n19034 ;
  assign n19036 = ~n19009 & n19035 ;
  assign n19037 = \u0_w_reg[0][20]/P0001  & ~n19036 ;
  assign n19038 = ~\u0_w_reg[0][20]/P0001  & n19036 ;
  assign n19039 = ~n19037 & ~n19038 ;
  assign n19040 = \u0_w_reg[1][20]/P0001  & n19039 ;
  assign n19041 = ~\u0_w_reg[1][20]/P0001  & ~n19039 ;
  assign n19042 = ~n19040 & ~n19041 ;
  assign n19043 = \u0_w_reg[2][20]/P0001  & n19042 ;
  assign n19044 = ~\u0_w_reg[2][20]/P0001  & ~n19042 ;
  assign n19045 = ~n19043 & ~n19044 ;
  assign n19046 = ~ld_pad & n19045 ;
  assign n19047 = \key[52]_pad  & ld_pad ;
  assign n19048 = ~n19046 & ~n19047 ;
  assign n19049 = ~\key[36]_pad  & ld_pad ;
  assign n19063 = ~n16032 & n16049 ;
  assign n19064 = ~n16443 & ~n19063 ;
  assign n19065 = ~\u0_w_reg[3][26]/P0001  & ~n19064 ;
  assign n19062 = \u0_w_reg[3][26]/P0001  & n16058 ;
  assign n19061 = n16036 & n16388 ;
  assign n19066 = ~n16403 & ~n19061 ;
  assign n19067 = ~n19062 & n19066 ;
  assign n19068 = ~n19065 & n19067 ;
  assign n19069 = \u0_w_reg[3][25]/P0001  & ~n19068 ;
  assign n19056 = ~\u0_w_reg[3][26]/P0001  & n17428 ;
  assign n19055 = \u0_w_reg[3][28]/P0001  & n16142 ;
  assign n19057 = ~n17339 & ~n18130 ;
  assign n19058 = ~n19055 & n19057 ;
  assign n19059 = ~n19056 & n19058 ;
  assign n19060 = ~\u0_w_reg[3][25]/P0001  & ~n19059 ;
  assign n19050 = ~n16118 & ~n17807 ;
  assign n19051 = ~\u0_w_reg[3][27]/P0001  & ~n19050 ;
  assign n19052 = n16019 & n16087 ;
  assign n19053 = ~n17287 & ~n19052 ;
  assign n19054 = \u0_w_reg[3][26]/P0001  & ~n19053 ;
  assign n19070 = ~n19051 & ~n19054 ;
  assign n19071 = ~n19060 & n19070 ;
  assign n19072 = ~n19069 & n19071 ;
  assign n19073 = ~\u0_w_reg[3][24]/P0001  & ~n19072 ;
  assign n19107 = \u0_w_reg[3][31]/P0001  & n16026 ;
  assign n19108 = ~n16066 & ~n19107 ;
  assign n19109 = ~\u0_w_reg[3][26]/P0001  & ~n19108 ;
  assign n19110 = ~\u0_w_reg[3][25]/P0001  & ~n16146 ;
  assign n19111 = ~n17804 & n19110 ;
  assign n19112 = ~n19109 & n19111 ;
  assign n19113 = ~n16366 & ~n16439 ;
  assign n19114 = ~\u0_w_reg[3][26]/P0001  & ~n19113 ;
  assign n19115 = \u0_w_reg[3][25]/P0001  & ~n17803 ;
  assign n19116 = ~n16053 & n19115 ;
  assign n19117 = ~n17464 & n19116 ;
  assign n19118 = ~n19114 & n19117 ;
  assign n19119 = ~n19112 & ~n19118 ;
  assign n19101 = ~\u0_w_reg[3][25]/P0001  & n16091 ;
  assign n19102 = ~n16428 & ~n19101 ;
  assign n19103 = n18090 & n19102 ;
  assign n19104 = ~n16015 & ~n17463 ;
  assign n19105 = n18101 & n19104 ;
  assign n19106 = ~n19103 & ~n19105 ;
  assign n19100 = n16032 & n16103 ;
  assign n19120 = ~n16106 & ~n19100 ;
  assign n19121 = ~n19106 & n19120 ;
  assign n19122 = ~n19119 & n19121 ;
  assign n19123 = \u0_w_reg[3][24]/P0001  & ~n19122 ;
  assign n19074 = ~n16013 & ~n17276 ;
  assign n19075 = ~n16376 & n19074 ;
  assign n19076 = ~n17806 & n19075 ;
  assign n19077 = ~n17826 & n19076 ;
  assign n19078 = \u0_w_reg[3][26]/P0001  & ~n19077 ;
  assign n19081 = ~n16111 & ~n17474 ;
  assign n19079 = n16019 & ~n16039 ;
  assign n19080 = n16386 & n19079 ;
  assign n19082 = ~n18820 & ~n19080 ;
  assign n19083 = n19081 & n19082 ;
  assign n19084 = ~n19078 & n19083 ;
  assign n19085 = ~\u0_w_reg[3][25]/P0001  & ~n19084 ;
  assign n19089 = ~n16051 & n16117 ;
  assign n19090 = ~n16044 & ~n17443 ;
  assign n19091 = ~n19089 & n19090 ;
  assign n19092 = ~\u0_w_reg[3][29]/P0001  & ~n19091 ;
  assign n19087 = ~n16120 & ~n16428 ;
  assign n19088 = n16386 & ~n19087 ;
  assign n19086 = n16036 & n17259 ;
  assign n19093 = ~n18110 & ~n19086 ;
  assign n19094 = ~n19088 & n19093 ;
  assign n19095 = ~n19092 & n19094 ;
  assign n19096 = \u0_w_reg[3][25]/P0001  & ~n19095 ;
  assign n19097 = ~\u0_w_reg[3][26]/P0001  & n16040 ;
  assign n19098 = ~n19055 & ~n19097 ;
  assign n19099 = \u0_w_reg[3][27]/P0001  & ~n19098 ;
  assign n19124 = ~n19096 & ~n19099 ;
  assign n19125 = ~n19085 & n19124 ;
  assign n19126 = ~n19123 & n19125 ;
  assign n19127 = ~n19073 & n19126 ;
  assign n19128 = \u0_w_reg[0][4]/P0001  & ~n19127 ;
  assign n19129 = ~\u0_w_reg[0][4]/P0001  & n19127 ;
  assign n19130 = ~n19128 & ~n19129 ;
  assign n19131 = \u0_w_reg[1][4]/P0001  & ~\u0_w_reg[2][4]/P0001  ;
  assign n19132 = ~\u0_w_reg[1][4]/P0001  & \u0_w_reg[2][4]/P0001  ;
  assign n19133 = ~n19131 & ~n19132 ;
  assign n19134 = n19130 & n19133 ;
  assign n19135 = ~n19130 & ~n19133 ;
  assign n19136 = ~n19134 & ~n19135 ;
  assign n19137 = ~ld_pad & n19136 ;
  assign n19138 = ~n19049 & ~n19137 ;
  assign n19140 = \u0_w_reg[3][12]/P0001  & ~n16770 ;
  assign n19139 = ~\u0_w_reg[3][12]/P0001  & n16770 ;
  assign n19141 = ~ld_pad & ~n19139 ;
  assign n19142 = ~n19140 & n19141 ;
  assign n19143 = \key[12]_pad  & ld_pad ;
  assign n19144 = ~n19142 & ~n19143 ;
  assign n19157 = ~n15603 & ~n16262 ;
  assign n19158 = ~\u0_w_reg[3][18]/P0001  & ~n19157 ;
  assign n19159 = ~n15558 & ~n16918 ;
  assign n19160 = ~n15658 & n19159 ;
  assign n19161 = ~n19158 & n19160 ;
  assign n19162 = \u0_w_reg[3][17]/P0001  & ~n19161 ;
  assign n19152 = ~n15522 & ~n15582 ;
  assign n19153 = ~\u0_w_reg[3][18]/P0001  & ~n19152 ;
  assign n19154 = ~n15587 & ~n16919 ;
  assign n19155 = ~n19153 & n19154 ;
  assign n19156 = ~\u0_w_reg[3][17]/P0001  & ~n19155 ;
  assign n19145 = ~n15637 & ~n18447 ;
  assign n19146 = ~\u0_w_reg[3][21]/P0001  & ~n19145 ;
  assign n19147 = ~n15540 & ~n19146 ;
  assign n19148 = ~\u0_w_reg[3][18]/P0001  & ~n19147 ;
  assign n19150 = n15504 & n16297 ;
  assign n19151 = n15511 & n15551 ;
  assign n19163 = ~n19150 & ~n19151 ;
  assign n19164 = ~n16845 & n19163 ;
  assign n19149 = n15628 & n16281 ;
  assign n19165 = ~n17019 & ~n19149 ;
  assign n19166 = n19164 & n19165 ;
  assign n19167 = ~n19148 & n19166 ;
  assign n19168 = ~n19156 & n19167 ;
  assign n19169 = ~n19162 & n19168 ;
  assign n19170 = \u0_w_reg[3][16]/P0001  & ~n19169 ;
  assign n19185 = ~n15504 & n17020 ;
  assign n19186 = ~n16269 & ~n19185 ;
  assign n19187 = ~\u0_w_reg[3][18]/P0001  & ~n19186 ;
  assign n19188 = n15511 & n15602 ;
  assign n19189 = \u0_w_reg[3][17]/P0001  & ~n16287 ;
  assign n19190 = ~n16777 & n19189 ;
  assign n19191 = ~n19188 & n19190 ;
  assign n19192 = ~n19187 & n19191 ;
  assign n19195 = ~\u0_w_reg[3][18]/P0001  & n16814 ;
  assign n19193 = \u0_w_reg[3][18]/P0001  & n15513 ;
  assign n19194 = n15504 & n15520 ;
  assign n19196 = ~n19193 & ~n19194 ;
  assign n19197 = n17065 & n19196 ;
  assign n19198 = ~n19195 & n19197 ;
  assign n19199 = ~n19192 & ~n19198 ;
  assign n19200 = ~\u0_w_reg[3][19]/P0001  & n15519 ;
  assign n19201 = ~n17080 & ~n19200 ;
  assign n19202 = \u0_w_reg[3][18]/P0001  & ~n19201 ;
  assign n19203 = ~n15647 & ~n16853 ;
  assign n19204 = ~\u0_w_reg[3][19]/P0001  & ~n19203 ;
  assign n19205 = ~n19202 & ~n19204 ;
  assign n19206 = ~n19199 & n19205 ;
  assign n19207 = ~\u0_w_reg[3][16]/P0001  & ~n19206 ;
  assign n19171 = ~n16269 & ~n16774 ;
  assign n19172 = ~\u0_w_reg[3][19]/P0001  & ~n19171 ;
  assign n19173 = ~n15538 & ~n15657 ;
  assign n19174 = ~n16222 & n19173 ;
  assign n19175 = ~n19172 & n19174 ;
  assign n19176 = \u0_w_reg[3][18]/P0001  & ~n19175 ;
  assign n19180 = ~n15650 & ~n18490 ;
  assign n19177 = \u0_w_reg[3][21]/P0001  & n15637 ;
  assign n19178 = \u0_w_reg[3][22]/P0001  & ~n15613 ;
  assign n19179 = n15660 & n19178 ;
  assign n19181 = ~n19177 & ~n19179 ;
  assign n19182 = n19180 & n19181 ;
  assign n19183 = ~n19176 & n19182 ;
  assign n19184 = ~\u0_w_reg[3][17]/P0001  & ~n19183 ;
  assign n19208 = ~\u0_w_reg[3][18]/P0001  & n16283 ;
  assign n19209 = ~n19193 & ~n19208 ;
  assign n19210 = \u0_w_reg[3][19]/P0001  & ~n19209 ;
  assign n19211 = \u0_w_reg[3][20]/P0001  & n16917 ;
  assign n19217 = ~n17003 & ~n17083 ;
  assign n19218 = ~n19211 & n19217 ;
  assign n19212 = ~n15520 & n15529 ;
  assign n19213 = ~n15556 & ~n19212 ;
  assign n19214 = ~\u0_w_reg[3][21]/P0001  & ~n19213 ;
  assign n19215 = ~n15630 & ~n16313 ;
  assign n19216 = n15648 & ~n19215 ;
  assign n19219 = ~n19214 & ~n19216 ;
  assign n19220 = n19218 & n19219 ;
  assign n19221 = \u0_w_reg[3][17]/P0001  & ~n19220 ;
  assign n19222 = ~n19210 & ~n19221 ;
  assign n19223 = ~n19184 & n19222 ;
  assign n19224 = ~n19207 & n19223 ;
  assign n19225 = ~n19170 & n19224 ;
  assign n19226 = ~\u0_r0_out_reg[28]/P0001  & n19225 ;
  assign n19227 = \u0_r0_out_reg[28]/P0001  & ~n19225 ;
  assign n19228 = ~n19226 & ~n19227 ;
  assign n19229 = \u0_w_reg[0][28]/P0001  & n19228 ;
  assign n19230 = ~\u0_w_reg[0][28]/P0001  & ~n19228 ;
  assign n19231 = ~n19229 & ~n19230 ;
  assign n19232 = ~ld_pad & n19231 ;
  assign n19233 = \key[124]_pad  & ld_pad ;
  assign n19234 = ~n19232 & ~n19233 ;
  assign n19236 = \u0_w_reg[1][28]/P0001  & n19231 ;
  assign n19235 = ~\u0_w_reg[1][28]/P0001  & ~n19231 ;
  assign n19237 = ~ld_pad & ~n19235 ;
  assign n19238 = ~n19236 & n19237 ;
  assign n19239 = \key[92]_pad  & ld_pad ;
  assign n19240 = ~n19238 & ~n19239 ;
  assign n19241 = \u0_w_reg[0][28]/P0001  & ~\u0_w_reg[2][28]/P0001  ;
  assign n19242 = ~\u0_w_reg[0][28]/P0001  & \u0_w_reg[2][28]/P0001  ;
  assign n19243 = ~n19241 & ~n19242 ;
  assign n19244 = n19228 & n19243 ;
  assign n19245 = ~n19228 & ~n19243 ;
  assign n19246 = ~n19244 & ~n19245 ;
  assign n19248 = \u0_w_reg[1][28]/P0001  & ~n19246 ;
  assign n19247 = ~\u0_w_reg[1][28]/P0001  & n19246 ;
  assign n19249 = ~ld_pad & ~n19247 ;
  assign n19250 = ~n19248 & n19249 ;
  assign n19251 = \key[60]_pad  & ld_pad ;
  assign n19252 = ~n19250 & ~n19251 ;
  assign n19253 = \key[28]_pad  & ld_pad ;
  assign n19254 = \u0_w_reg[1][28]/P0001  & ~\u0_w_reg[3][28]/P0001  ;
  assign n19255 = ~\u0_w_reg[1][28]/P0001  & \u0_w_reg[3][28]/P0001  ;
  assign n19256 = ~n19254 & ~n19255 ;
  assign n19258 = ~n19246 & ~n19256 ;
  assign n19257 = n19246 & n19256 ;
  assign n19259 = ~ld_pad & ~n19257 ;
  assign n19260 = ~n19258 & n19259 ;
  assign n19261 = ~n19253 & ~n19260 ;
  assign n19262 = ~ld_pad & n17361 ;
  assign n19263 = \key[103]_pad  & ld_pad ;
  assign n19264 = ~n19262 & ~n19263 ;
  assign n19266 = \u0_w_reg[1][7]/P0001  & n17361 ;
  assign n19265 = ~\u0_w_reg[1][7]/P0001  & ~n17361 ;
  assign n19267 = ~ld_pad & ~n19265 ;
  assign n19268 = ~n19266 & n19267 ;
  assign n19269 = \key[71]_pad  & ld_pad ;
  assign n19270 = ~n19268 & ~n19269 ;
  assign n19272 = \u0_w_reg[3][7]/P0001  & ~n17367 ;
  assign n19271 = ~\u0_w_reg[3][7]/P0001  & n17367 ;
  assign n19273 = ~ld_pad & ~n19271 ;
  assign n19274 = ~n19272 & n19273 ;
  assign n19275 = \key[7]_pad  & ld_pad ;
  assign n19276 = ~n19274 & ~n19275 ;
  assign n19277 = ~ld_pad & n17486 ;
  assign n19278 = \key[96]_pad  & ld_pad ;
  assign n19279 = ~n19277 & ~n19278 ;
  assign n19280 = ~ld_pad & n17588 ;
  assign n19281 = \key[106]_pad  & ld_pad ;
  assign n19282 = ~n19280 & ~n19281 ;
  assign n19283 = ~ld_pad & n17696 ;
  assign n19284 = \key[112]_pad  & ld_pad ;
  assign n19285 = ~n19283 & ~n19284 ;
  assign n19286 = ~ld_pad & n17793 ;
  assign n19287 = \key[114]_pad  & ld_pad ;
  assign n19288 = ~n19286 & ~n19287 ;
  assign n19289 = ~ld_pad & n17885 ;
  assign n19290 = \key[98]_pad  & ld_pad ;
  assign n19291 = ~n19289 & ~n19290 ;
  assign n19293 = \u0_w_reg[1][0]/P0001  & n17486 ;
  assign n19292 = ~\u0_w_reg[1][0]/P0001  & ~n17486 ;
  assign n19294 = ~ld_pad & ~n19292 ;
  assign n19295 = ~n19293 & n19294 ;
  assign n19296 = \key[64]_pad  & ld_pad ;
  assign n19297 = ~n19295 & ~n19296 ;
  assign n19299 = \u0_w_reg[1][10]/P0001  & n17588 ;
  assign n19298 = ~\u0_w_reg[1][10]/P0001  & ~n17588 ;
  assign n19300 = ~ld_pad & ~n19298 ;
  assign n19301 = ~n19299 & n19300 ;
  assign n19302 = \key[74]_pad  & ld_pad ;
  assign n19303 = ~n19301 & ~n19302 ;
  assign n19305 = \u0_w_reg[1][16]/P0001  & n17696 ;
  assign n19304 = ~\u0_w_reg[1][16]/P0001  & ~n17696 ;
  assign n19306 = ~ld_pad & ~n19304 ;
  assign n19307 = ~n19305 & n19306 ;
  assign n19308 = \key[80]_pad  & ld_pad ;
  assign n19309 = ~n19307 & ~n19308 ;
  assign n19311 = \u0_w_reg[1][18]/P0001  & n17793 ;
  assign n19310 = ~\u0_w_reg[1][18]/P0001  & ~n17793 ;
  assign n19312 = ~ld_pad & ~n19310 ;
  assign n19313 = ~n19311 & n19312 ;
  assign n19314 = \key[82]_pad  & ld_pad ;
  assign n19315 = ~n19313 & ~n19314 ;
  assign n19316 = ~ld_pad & n17888 ;
  assign n19317 = \key[66]_pad  & ld_pad ;
  assign n19318 = ~n19316 & ~n19317 ;
  assign n19320 = \u0_w_reg[3][0]/P0001  & ~n17492 ;
  assign n19319 = ~\u0_w_reg[3][0]/P0001  & n17492 ;
  assign n19321 = ~ld_pad & ~n19319 ;
  assign n19322 = ~n19320 & n19321 ;
  assign n19323 = \key[0]_pad  & ld_pad ;
  assign n19324 = ~n19322 & ~n19323 ;
  assign n19326 = \u0_w_reg[3][10]/P0001  & ~n17594 ;
  assign n19325 = ~\u0_w_reg[3][10]/P0001  & n17594 ;
  assign n19327 = ~ld_pad & ~n19325 ;
  assign n19328 = ~n19326 & n19327 ;
  assign n19329 = \key[10]_pad  & ld_pad ;
  assign n19330 = ~n19328 & ~n19329 ;
  assign n19332 = \u0_w_reg[3][16]/P0001  & ~n17702 ;
  assign n19331 = ~\u0_w_reg[3][16]/P0001  & n17702 ;
  assign n19333 = ~ld_pad & ~n19331 ;
  assign n19334 = ~n19332 & n19333 ;
  assign n19335 = \key[16]_pad  & ld_pad ;
  assign n19336 = ~n19334 & ~n19335 ;
  assign n19338 = \u0_w_reg[3][18]/P0001  & ~n17799 ;
  assign n19337 = ~\u0_w_reg[3][18]/P0001  & n17799 ;
  assign n19339 = ~ld_pad & ~n19337 ;
  assign n19340 = ~n19338 & n19339 ;
  assign n19341 = \key[18]_pad  & ld_pad ;
  assign n19342 = ~n19340 & ~n19341 ;
  assign n19344 = \u0_w_reg[3][2]/P0001  & n17891 ;
  assign n19343 = ~\u0_w_reg[3][2]/P0001  & ~n17891 ;
  assign n19345 = ~ld_pad & ~n19343 ;
  assign n19346 = ~n19344 & n19345 ;
  assign n19347 = \key[2]_pad  & ld_pad ;
  assign n19348 = ~n19346 & ~n19347 ;
  assign n19349 = ~\u0_w_reg[0][5]/P0001  & ~n12580 ;
  assign n19350 = \u0_w_reg[0][5]/P0001  & n12580 ;
  assign n19351 = ~n19349 & ~n19350 ;
  assign n19352 = ~ld_pad & n17983 ;
  assign n19353 = \key[110]_pad  & ld_pad ;
  assign n19354 = ~n19352 & ~n19353 ;
  assign n19355 = ~ld_pad & n18069 ;
  assign n19356 = \key[118]_pad  & ld_pad ;
  assign n19357 = ~n19355 & ~n19356 ;
  assign n19358 = ~ld_pad & n18153 ;
  assign n19359 = \key[102]_pad  & ld_pad ;
  assign n19360 = ~n19358 & ~n19359 ;
  assign n19362 = \u0_w_reg[1][14]/P0001  & n17983 ;
  assign n19361 = ~\u0_w_reg[1][14]/P0001  & ~n17983 ;
  assign n19363 = ~ld_pad & ~n19361 ;
  assign n19364 = ~n19362 & n19363 ;
  assign n19365 = \key[78]_pad  & ld_pad ;
  assign n19366 = ~n19364 & ~n19365 ;
  assign n19368 = \u0_w_reg[1][22]/P0001  & n18069 ;
  assign n19367 = ~\u0_w_reg[1][22]/P0001  & ~n18069 ;
  assign n19369 = ~ld_pad & ~n19367 ;
  assign n19370 = ~n19368 & n19369 ;
  assign n19371 = \key[86]_pad  & ld_pad ;
  assign n19372 = ~n19370 & ~n19371 ;
  assign n19374 = \u0_w_reg[1][6]/P0001  & n18153 ;
  assign n19373 = ~\u0_w_reg[1][6]/P0001  & ~n18153 ;
  assign n19375 = ~ld_pad & ~n19373 ;
  assign n19376 = ~n19374 & n19375 ;
  assign n19377 = \key[70]_pad  & ld_pad ;
  assign n19378 = ~n19376 & ~n19377 ;
  assign n19380 = \u0_w_reg[3][14]/P0001  & ~n17989 ;
  assign n19379 = ~\u0_w_reg[3][14]/P0001  & n17989 ;
  assign n19381 = ~ld_pad & ~n19379 ;
  assign n19382 = ~n19380 & n19381 ;
  assign n19383 = \key[14]_pad  & ld_pad ;
  assign n19384 = ~n19382 & ~n19383 ;
  assign n19386 = \u0_w_reg[3][22]/P0001  & ~n18075 ;
  assign n19385 = ~\u0_w_reg[3][22]/P0001  & n18075 ;
  assign n19387 = ~ld_pad & ~n19385 ;
  assign n19388 = ~n19386 & n19387 ;
  assign n19389 = \key[22]_pad  & ld_pad ;
  assign n19390 = ~n19388 & ~n19389 ;
  assign n19392 = \u0_w_reg[3][6]/P0001  & ~n18159 ;
  assign n19391 = ~\u0_w_reg[3][6]/P0001  & n18159 ;
  assign n19393 = ~ld_pad & ~n19391 ;
  assign n19394 = ~n19392 & n19393 ;
  assign n19395 = \key[6]_pad  & ld_pad ;
  assign n19396 = ~n19394 & ~n19395 ;
  assign n19397 = ~ld_pad & n18255 ;
  assign n19398 = \key[109]_pad  & ld_pad ;
  assign n19399 = ~n19397 & ~n19398 ;
  assign n19400 = ~ld_pad & n18355 ;
  assign n19401 = \key[111]_pad  & ld_pad ;
  assign n19402 = ~n19400 & ~n19401 ;
  assign n19403 = ~ld_pad & n18437 ;
  assign n19404 = \key[104]_pad  & ld_pad ;
  assign n19405 = ~n19403 & ~n19404 ;
  assign n19407 = \u0_w_reg[1][13]/P0001  & n18255 ;
  assign n19406 = ~\u0_w_reg[1][13]/P0001  & ~n18255 ;
  assign n19408 = ~ld_pad & ~n19406 ;
  assign n19409 = ~n19407 & n19408 ;
  assign n19410 = \key[77]_pad  & ld_pad ;
  assign n19411 = ~n19409 & ~n19410 ;
  assign n19412 = ~ld_pad & n18358 ;
  assign n19413 = \key[79]_pad  & ld_pad ;
  assign n19414 = ~n19412 & ~n19413 ;
  assign n19416 = \u0_w_reg[1][8]/P0001  & n18437 ;
  assign n19415 = ~\u0_w_reg[1][8]/P0001  & ~n18437 ;
  assign n19417 = ~ld_pad & ~n19415 ;
  assign n19418 = ~n19416 & n19417 ;
  assign n19419 = \key[72]_pad  & ld_pad ;
  assign n19420 = ~n19418 & ~n19419 ;
  assign n19422 = \u0_w_reg[3][13]/P0001  & ~n18261 ;
  assign n19421 = ~\u0_w_reg[3][13]/P0001  & n18261 ;
  assign n19423 = ~ld_pad & ~n19421 ;
  assign n19424 = ~n19422 & n19423 ;
  assign n19425 = \key[13]_pad  & ld_pad ;
  assign n19426 = ~n19424 & ~n19425 ;
  assign n19428 = \u0_w_reg[3][15]/P0001  & n18361 ;
  assign n19427 = ~\u0_w_reg[3][15]/P0001  & ~n18361 ;
  assign n19429 = ~ld_pad & ~n19427 ;
  assign n19430 = ~n19428 & n19429 ;
  assign n19431 = \key[15]_pad  & ld_pad ;
  assign n19432 = ~n19430 & ~n19431 ;
  assign n19434 = \u0_w_reg[3][8]/P0001  & ~n18443 ;
  assign n19433 = ~\u0_w_reg[3][8]/P0001  & n18443 ;
  assign n19435 = ~ld_pad & ~n19433 ;
  assign n19436 = ~n19434 & n19435 ;
  assign n19437 = \key[8]_pad  & ld_pad ;
  assign n19438 = ~n19436 & ~n19437 ;
  assign n19439 = ~\u0_w_reg[0][29]/P0001  & ~n12714 ;
  assign n19440 = \u0_w_reg[0][29]/P0001  & n12714 ;
  assign n19441 = ~n19439 & ~n19440 ;
  assign n19442 = ~\u0_w_reg[3][29]/P0001  & ~n1479 ;
  assign n19443 = \u0_w_reg[3][29]/P0001  & n1479 ;
  assign n19444 = ~n19442 & ~n19443 ;
  assign n19445 = ~\u0_w_reg[2][29]/P0001  & ~n1142 ;
  assign n19446 = \u0_w_reg[2][29]/P0001  & n1142 ;
  assign n19447 = ~n19445 & ~n19446 ;
  assign n19448 = ~\u0_w_reg[1][29]/P0002  & ~n9289 ;
  assign n19449 = \u0_w_reg[1][29]/P0002  & n9289 ;
  assign n19450 = ~n19448 & ~n19449 ;
  assign n19451 = ~ld_pad & n18645 ;
  assign n19452 = \key[119]_pad  & ld_pad ;
  assign n19453 = ~n19451 & ~n19452 ;
  assign n19454 = ~ld_pad & n18648 ;
  assign n19455 = \key[87]_pad  & ld_pad ;
  assign n19456 = ~n19454 & ~n19455 ;
  assign n19458 = \u0_w_reg[3][23]/P0001  & n18651 ;
  assign n19457 = ~\u0_w_reg[3][23]/P0001  & ~n18651 ;
  assign n19459 = ~ld_pad & ~n19457 ;
  assign n19460 = ~n19458 & n19459 ;
  assign n19461 = \key[23]_pad  & ld_pad ;
  assign n19462 = ~n19460 & ~n19461 ;
  assign n19463 = ~\u0_w_reg[3][8]/P0001  & ~n3592 ;
  assign n19464 = \u0_w_reg[3][8]/P0001  & n3592 ;
  assign n19465 = ~n19463 & ~n19464 ;
  assign n19466 = ~\u0_w_reg[0][11]/P0001  & ~n14567 ;
  assign n19467 = \u0_w_reg[0][11]/P0001  & n14567 ;
  assign n19468 = ~n19466 & ~n19467 ;
  assign n19469 = ~\u0_w_reg[3][11]/P0001  & ~n4059 ;
  assign n19470 = \u0_w_reg[3][11]/P0001  & n4059 ;
  assign n19471 = ~n19469 & ~n19470 ;
  assign n19472 = ~\u0_w_reg[2][11]/P0001  & ~n7206 ;
  assign n19473 = \u0_w_reg[2][11]/P0001  & n7206 ;
  assign n19474 = ~n19472 & ~n19473 ;
  assign n19475 = ~\u0_w_reg[1][11]/P0001  & ~n10775 ;
  assign n19476 = \u0_w_reg[1][11]/P0001  & n10775 ;
  assign n19477 = ~n19475 & ~n19476 ;
  assign n19478 = ~\u0_w_reg[0][12]/P0001  & ~n12827 ;
  assign n19479 = \u0_w_reg[0][12]/P0001  & n12827 ;
  assign n19480 = ~n19478 & ~n19479 ;
  assign n19481 = ~\u0_w_reg[2][12]/P0001  & ~n6055 ;
  assign n19482 = \u0_w_reg[2][12]/P0001  & n6055 ;
  assign n19483 = ~n19481 & ~n19482 ;
  assign n19484 = ~\u0_w_reg[1][12]/P0001  & ~n9516 ;
  assign n19485 = \u0_w_reg[1][12]/P0001  & n9516 ;
  assign n19486 = ~n19484 & ~n19485 ;
  assign n19487 = ~\u0_w_reg[0][8]/P0001  & ~n13379 ;
  assign n19488 = \u0_w_reg[0][8]/P0001  & n13379 ;
  assign n19489 = ~n19487 & ~n19488 ;
  assign n19490 = ~\u0_w_reg[0][24]/P0001  & ~n14316 ;
  assign n19491 = \u0_w_reg[0][24]/P0001  & n14316 ;
  assign n19492 = ~n19490 & ~n19491 ;
  assign n19493 = ~\u0_w_reg[0][27]/P0001  & ~n14970 ;
  assign n19494 = \u0_w_reg[0][27]/P0001  & n14970 ;
  assign n19495 = ~n19493 & ~n19494 ;
  assign n19496 = ~\u0_w_reg[3][24]/P0001  & ~n4161 ;
  assign n19497 = \u0_w_reg[3][24]/P0001  & n4161 ;
  assign n19498 = ~n19496 & ~n19497 ;
  assign n19499 = ~\u0_w_reg[3][27]/P0001  & ~n3888 ;
  assign n19500 = \u0_w_reg[3][27]/P0001  & n3888 ;
  assign n19501 = ~n19499 & ~n19500 ;
  assign n19502 = ~\u0_w_reg[2][8]/P0001  & ~n6927 ;
  assign n19503 = \u0_w_reg[2][8]/P0001  & n6927 ;
  assign n19504 = ~n19502 & ~n19503 ;
  assign n19505 = ~\u0_w_reg[2][24]/P0001  & ~n6472 ;
  assign n19506 = \u0_w_reg[2][24]/P0001  & n6472 ;
  assign n19507 = ~n19505 & ~n19506 ;
  assign n19508 = ~\u0_w_reg[2][27]/P0001  & ~n7040 ;
  assign n19509 = \u0_w_reg[2][27]/P0001  & n7040 ;
  assign n19510 = ~n19508 & ~n19509 ;
  assign n19511 = ~\u0_w_reg[1][8]/P0001  & ~n11073 ;
  assign n19512 = \u0_w_reg[1][8]/P0001  & n11073 ;
  assign n19513 = ~n19511 & ~n19512 ;
  assign n19514 = ~\u0_w_reg[1][24]/P0002  & ~n10248 ;
  assign n19515 = \u0_w_reg[1][24]/P0002  & n10248 ;
  assign n19516 = ~n19514 & ~n19515 ;
  assign n19517 = ~\u0_w_reg[1][27]/P0001  & ~n10602 ;
  assign n19518 = \u0_w_reg[1][27]/P0001  & n10602 ;
  assign n19519 = ~n19517 & ~n19518 ;
  assign n19520 = ~ld_pad & n18765 ;
  assign n19521 = \key[113]_pad  & ld_pad ;
  assign n19522 = ~n19520 & ~n19521 ;
  assign n19523 = ~ld_pad & n18854 ;
  assign n19524 = \key[97]_pad  & ld_pad ;
  assign n19525 = ~n19523 & ~n19524 ;
  assign n19526 = ~ld_pad & n18945 ;
  assign n19527 = \key[105]_pad  & ld_pad ;
  assign n19528 = ~n19526 & ~n19527 ;
  assign n19530 = \u0_w_reg[1][17]/P0001  & n18765 ;
  assign n19529 = ~\u0_w_reg[1][17]/P0001  & ~n18765 ;
  assign n19531 = ~ld_pad & ~n19529 ;
  assign n19532 = ~n19530 & n19531 ;
  assign n19533 = \key[81]_pad  & ld_pad ;
  assign n19534 = ~n19532 & ~n19533 ;
  assign n19536 = \u0_w_reg[1][1]/P0001  & n18854 ;
  assign n19535 = ~\u0_w_reg[1][1]/P0001  & ~n18854 ;
  assign n19537 = ~ld_pad & ~n19535 ;
  assign n19538 = ~n19536 & n19537 ;
  assign n19539 = \key[65]_pad  & ld_pad ;
  assign n19540 = ~n19538 & ~n19539 ;
  assign n19542 = \u0_w_reg[1][9]/P0001  & n18945 ;
  assign n19541 = ~\u0_w_reg[1][9]/P0001  & ~n18945 ;
  assign n19543 = ~ld_pad & ~n19541 ;
  assign n19544 = ~n19542 & n19543 ;
  assign n19545 = \key[73]_pad  & ld_pad ;
  assign n19546 = ~n19544 & ~n19545 ;
  assign n19548 = \u0_w_reg[3][17]/P0001  & ~n18771 ;
  assign n19547 = ~\u0_w_reg[3][17]/P0001  & n18771 ;
  assign n19549 = ~ld_pad & ~n19547 ;
  assign n19550 = ~n19548 & n19549 ;
  assign n19551 = \key[17]_pad  & ld_pad ;
  assign n19552 = ~n19550 & ~n19551 ;
  assign n19554 = \u0_w_reg[3][1]/P0001  & ~n18860 ;
  assign n19553 = ~\u0_w_reg[3][1]/P0001  & n18860 ;
  assign n19555 = ~ld_pad & ~n19553 ;
  assign n19556 = ~n19554 & n19555 ;
  assign n19557 = \key[1]_pad  & ld_pad ;
  assign n19558 = ~n19556 & ~n19557 ;
  assign n19560 = \u0_w_reg[3][9]/P0001  & ~n18951 ;
  assign n19559 = ~\u0_w_reg[3][9]/P0001  & n18951 ;
  assign n19561 = ~ld_pad & ~n19559 ;
  assign n19562 = ~n19560 & n19561 ;
  assign n19563 = \key[9]_pad  & ld_pad ;
  assign n19564 = ~n19562 & ~n19563 ;
  assign n19565 = ~\u0_w_reg[0][19]/P0001  & ~n14491 ;
  assign n19566 = \u0_w_reg[0][19]/P0001  & n14491 ;
  assign n19567 = ~n19565 & ~n19566 ;
  assign n19568 = ~\u0_w_reg[3][19]/P0001  & ~n3966 ;
  assign n19569 = \u0_w_reg[3][19]/P0001  & n3966 ;
  assign n19570 = ~n19568 & ~n19569 ;
  assign n19571 = ~\u0_w_reg[2][19]/P0001  & ~n7115 ;
  assign n19572 = \u0_w_reg[2][19]/P0001  & n7115 ;
  assign n19573 = ~n19571 & ~n19572 ;
  assign n19574 = ~\u0_w_reg[1][19]/P0001  & ~n10682 ;
  assign n19575 = \u0_w_reg[1][19]/P0001  & n10682 ;
  assign n19576 = ~n19574 & ~n19575 ;
  assign n19577 = ~\u0_w_reg[0][9]/P0001  & ~n13835 ;
  assign n19578 = \u0_w_reg[0][9]/P0001  & n13835 ;
  assign n19579 = ~n19577 & ~n19578 ;
  assign n19580 = ~\u0_w_reg[2][9]/P0001  & ~n6743 ;
  assign n19581 = \u0_w_reg[2][9]/P0001  & n6743 ;
  assign n19582 = ~n19580 & ~n19581 ;
  assign n19583 = ~\u0_w_reg[1][9]/P0001  & ~n10508 ;
  assign n19584 = \u0_w_reg[1][9]/P0001  & n10508 ;
  assign n19585 = ~n19583 & ~n19584 ;
  assign n19586 = ~\u0_w_reg[0][13]/P0001  & ~n12405 ;
  assign n19587 = \u0_w_reg[0][13]/P0001  & n12405 ;
  assign n19588 = ~n19586 & ~n19587 ;
  assign n19589 = ~\u0_w_reg[0][21]/P0001  & ~n12233 ;
  assign n19590 = \u0_w_reg[0][21]/P0001  & n12233 ;
  assign n19591 = ~n19589 & ~n19590 ;
  assign n19592 = ~\u0_w_reg[3][13]/P0001  & ~n2939 ;
  assign n19593 = \u0_w_reg[3][13]/P0001  & n2939 ;
  assign n19594 = ~n19592 & ~n19593 ;
  assign n19595 = ~\u0_w_reg[3][21]/P0001  & ~n2835 ;
  assign n19596 = \u0_w_reg[3][21]/P0001  & n2835 ;
  assign n19597 = ~n19595 & ~n19596 ;
  assign n19598 = ~\u0_w_reg[2][13]/P0001  & ~n5931 ;
  assign n19599 = \u0_w_reg[2][13]/P0001  & n5931 ;
  assign n19600 = ~n19598 & ~n19599 ;
  assign n19601 = ~\u0_w_reg[2][21]/P0001  & ~n973 ;
  assign n19602 = \u0_w_reg[2][21]/P0001  & n973 ;
  assign n19603 = ~n19601 & ~n19602 ;
  assign n19604 = ~\u0_w_reg[1][13]/P0001  & ~n8678 ;
  assign n19605 = \u0_w_reg[1][13]/P0001  & n8678 ;
  assign n19606 = ~n19604 & ~n19605 ;
  assign n19607 = ~\u0_w_reg[1][21]/P0001  & ~n8507 ;
  assign n19608 = \u0_w_reg[1][21]/P0001  & n8507 ;
  assign n19609 = ~n19607 & ~n19608 ;
  assign n19610 = ~ld_pad & n19039 ;
  assign n19611 = \key[116]_pad  & ld_pad ;
  assign n19612 = ~n19610 & ~n19611 ;
  assign n19613 = ~ld_pad & n19130 ;
  assign n19614 = \key[100]_pad  & ld_pad ;
  assign n19615 = ~n19613 & ~n19614 ;
  assign n19616 = ~ld_pad & n19042 ;
  assign n19617 = \key[84]_pad  & ld_pad ;
  assign n19618 = ~n19616 & ~n19617 ;
  assign n19620 = \u0_w_reg[1][4]/P0001  & n19130 ;
  assign n19619 = ~\u0_w_reg[1][4]/P0001  & ~n19130 ;
  assign n19621 = ~ld_pad & ~n19619 ;
  assign n19622 = ~n19620 & n19621 ;
  assign n19623 = \key[68]_pad  & ld_pad ;
  assign n19624 = ~n19622 & ~n19623 ;
  assign n19626 = \u0_w_reg[3][20]/P0001  & n19045 ;
  assign n19625 = ~\u0_w_reg[3][20]/P0001  & ~n19045 ;
  assign n19627 = ~ld_pad & ~n19625 ;
  assign n19628 = ~n19626 & n19627 ;
  assign n19629 = \key[20]_pad  & ld_pad ;
  assign n19630 = ~n19628 & ~n19629 ;
  assign n19632 = \u0_w_reg[3][4]/P0001  & ~n19136 ;
  assign n19631 = ~\u0_w_reg[3][4]/P0001  & n19136 ;
  assign n19633 = ~ld_pad & ~n19631 ;
  assign n19634 = ~n19632 & n19633 ;
  assign n19635 = \key[4]_pad  & ld_pad ;
  assign n19636 = ~n19634 & ~n19635 ;
  assign n19637 = ~\u0_w_reg[0][3]/P0001  & ~n14651 ;
  assign n19638 = \u0_w_reg[0][3]/P0001  & n14651 ;
  assign n19639 = ~n19637 & ~n19638 ;
  assign n19640 = ~\u0_w_reg[3][9]/P0001  & ~n4248 ;
  assign n19641 = \u0_w_reg[3][9]/P0001  & n4248 ;
  assign n19642 = ~n19640 & ~n19641 ;
  assign n19643 = ~\u0_w_reg[0][17]/P0001  & ~n14210 ;
  assign n19644 = \u0_w_reg[0][17]/P0001  & n14210 ;
  assign n19645 = ~n19643 & ~n19644 ;
  assign n19646 = ~\u0_w_reg[3][17]/P0001  & ~n3681 ;
  assign n19647 = \u0_w_reg[3][17]/P0001  & n3681 ;
  assign n19648 = ~n19646 & ~n19647 ;
  assign n19649 = ~\u0_w_reg[2][17]/P0001  & ~n6304 ;
  assign n19650 = \u0_w_reg[2][17]/P0001  & n6304 ;
  assign n19651 = ~n19649 & ~n19650 ;
  assign n19652 = ~\u0_w_reg[1][17]/P0001  & ~n10081 ;
  assign n19653 = \u0_w_reg[1][17]/P0001  & n10081 ;
  assign n19654 = ~n19652 & ~n19653 ;
  assign n19655 = ~\u0_w_reg[0][4]/P0001  & ~n12962 ;
  assign n19656 = \u0_w_reg[0][4]/P0001  & n12962 ;
  assign n19657 = ~n19655 & ~n19656 ;
  assign n19658 = ~\u0_w_reg[3][12]/P0001  & ~n3069 ;
  assign n19659 = \u0_w_reg[3][12]/P0001  & n3069 ;
  assign n19660 = ~n19658 & ~n19659 ;
  assign n19661 = ~\u0_w_reg[0][16]/P0001  & ~n13465 ;
  assign n19662 = \u0_w_reg[0][16]/P0001  & n13465 ;
  assign n19663 = ~n19661 & ~n19662 ;
  assign n19664 = ~\u0_w_reg[3][16]/P0001  & ~n4674 ;
  assign n19665 = \u0_w_reg[3][16]/P0001  & n4674 ;
  assign n19666 = ~n19664 & ~n19665 ;
  assign n19667 = ~\u0_w_reg[2][16]/P0001  & ~n7408 ;
  assign n19668 = \u0_w_reg[2][16]/P0001  & n7408 ;
  assign n19669 = ~n19667 & ~n19668 ;
  assign n19670 = ~\u0_w_reg[1][16]/P0001  & ~n10996 ;
  assign n19671 = \u0_w_reg[1][16]/P0001  & n10996 ;
  assign n19672 = ~n19670 & ~n19671 ;
  assign n19673 = ~\u0_w_reg[0][1]/P0001  & ~n13752 ;
  assign n19674 = \u0_w_reg[0][1]/P0001  & n13752 ;
  assign n19675 = ~n19673 & ~n19674 ;
  assign n19676 = ~\u0_w_reg[0][6]/P0001  & ~n15289 ;
  assign n19677 = \u0_w_reg[0][6]/P0001  & n15289 ;
  assign n19678 = ~n19676 & ~n19677 ;
  assign n19679 = ~\u0_w_reg[0][0]/P0001  & ~n14113 ;
  assign n19680 = \u0_w_reg[0][0]/P0001  & n14113 ;
  assign n19681 = ~n19679 & ~n19680 ;
  assign n19682 = ~\u0_w_reg[0][10]/P0001  & ~n14894 ;
  assign n19683 = \u0_w_reg[0][10]/P0001  & n14894 ;
  assign n19684 = ~n19682 & ~n19683 ;
  assign n19685 = ~\u0_w_reg[0][15]/P0001  & ~n13922 ;
  assign n19686 = \u0_w_reg[0][15]/P0001  & n13922 ;
  assign n19687 = ~n19685 & ~n19686 ;
  assign n19688 = ~\u0_w_reg[0][31]/P0001  & ~n14400 ;
  assign n19689 = \u0_w_reg[0][31]/P0001  & n14400 ;
  assign n19690 = ~n19688 & ~n19689 ;
  assign n19691 = ~\u0_w_reg[3][31]/P0001  & ~n2304 ;
  assign n19692 = \u0_w_reg[3][31]/P0001  & n2304 ;
  assign n19693 = ~n19691 & ~n19692 ;
  assign n19694 = ~\u0_w_reg[2][10]/P0001  & ~n7655 ;
  assign n19695 = \u0_w_reg[2][10]/P0001  & n7655 ;
  assign n19696 = ~n19694 & ~n19695 ;
  assign n19697 = ~\u0_w_reg[2][15]/P0001  & ~n5631 ;
  assign n19698 = \u0_w_reg[2][15]/P0001  & n5631 ;
  assign n19699 = ~n19697 & ~n19698 ;
  assign n19700 = ~\u0_w_reg[2][31]/P0001  & ~n5417 ;
  assign n19701 = \u0_w_reg[2][31]/P0001  & n5417 ;
  assign n19702 = ~n19700 & ~n19701 ;
  assign n19703 = ~\u0_w_reg[1][10]/P0001  & ~n11384 ;
  assign n19704 = \u0_w_reg[1][10]/P0001  & n11384 ;
  assign n19705 = ~n19703 & ~n19704 ;
  assign n19706 = ~\u0_w_reg[1][15]/P0001  & ~n9980 ;
  assign n19707 = \u0_w_reg[1][15]/P0001  & n9980 ;
  assign n19708 = ~n19706 & ~n19707 ;
  assign n19709 = ~\u0_w_reg[1][31]/P0001  & ~n9783 ;
  assign n19710 = \u0_w_reg[1][31]/P0001  & n9783 ;
  assign n19711 = ~n19709 & ~n19710 ;
  assign n19712 = ~\u0_w_reg[0][18]/P0001  & ~n14729 ;
  assign n19713 = \u0_w_reg[0][18]/P0001  & n14729 ;
  assign n19714 = ~n19712 & ~n19713 ;
  assign n19715 = ~\u0_w_reg[3][18]/P0001  & ~n4433 ;
  assign n19716 = \u0_w_reg[3][18]/P0001  & n4433 ;
  assign n19717 = ~n19715 & ~n19716 ;
  assign n19718 = ~\u0_w_reg[2][18]/P0001  & ~n7508 ;
  assign n19719 = \u0_w_reg[2][18]/P0001  & n7508 ;
  assign n19720 = ~n19718 & ~n19719 ;
  assign n19721 = ~\u0_w_reg[1][18]/P0001  & ~n11240 ;
  assign n19722 = \u0_w_reg[1][18]/P0001  & n11240 ;
  assign n19723 = ~n19721 & ~n19722 ;
  assign n19724 = ~\u0_w_reg[0][23]/P0001  & ~n13558 ;
  assign n19725 = \u0_w_reg[0][23]/P0001  & n13558 ;
  assign n19726 = ~n19724 & ~n19725 ;
  assign n19727 = ~\u0_w_reg[3][15]/P0001  & ~n2529 ;
  assign n19728 = \u0_w_reg[3][15]/P0001  & n2529 ;
  assign n19729 = ~n19727 & ~n19728 ;
  assign n19730 = ~\u0_w_reg[3][23]/P0001  & ~n2199 ;
  assign n19731 = \u0_w_reg[3][23]/P0001  & n2199 ;
  assign n19732 = ~n19730 & ~n19731 ;
  assign n19733 = ~\u0_w_reg[2][23]/P0001  & ~n5516 ;
  assign n19734 = \u0_w_reg[2][23]/P0001  & n5516 ;
  assign n19735 = ~n19733 & ~n19734 ;
  assign n19736 = ~\u0_w_reg[1][23]/P0001  & ~n9874 ;
  assign n19737 = \u0_w_reg[1][23]/P0001  & n9874 ;
  assign n19738 = ~n19736 & ~n19737 ;
  assign n19739 = ~\u0_w_reg[0][26]/P0001  & ~n14801 ;
  assign n19740 = \u0_w_reg[0][26]/P0001  & n14801 ;
  assign n19741 = ~n19739 & ~n19740 ;
  assign n19742 = ~\u0_w_reg[3][26]/P0001  & ~n4505 ;
  assign n19743 = \u0_w_reg[3][26]/P0001  & n4505 ;
  assign n19744 = ~n19742 & ~n19743 ;
  assign n19745 = ~\u0_w_reg[2][26]/P0001  & ~n7580 ;
  assign n19746 = \u0_w_reg[2][26]/P0001  & n7580 ;
  assign n19747 = ~n19745 & ~n19746 ;
  assign n19748 = ~\u0_w_reg[1][26]/P0001  & ~n11312 ;
  assign n19749 = \u0_w_reg[1][26]/P0001  & n11312 ;
  assign n19750 = ~n19748 & ~n19749 ;
  assign n19751 = ~\u0_w_reg[0][7]/P0001  & ~n14033 ;
  assign n19752 = \u0_w_reg[0][7]/P0001  & n14033 ;
  assign n19753 = ~n19751 & ~n19752 ;
  assign n19754 = ~\u0_w_reg[0][30]/P0001  & ~n13091 ;
  assign n19755 = \u0_w_reg[0][30]/P0001  & n13091 ;
  assign n19756 = ~n19754 & ~n19755 ;
  assign n19757 = ~\u0_w_reg[3][30]/P0001  & ~n1581 ;
  assign n19758 = \u0_w_reg[3][30]/P0001  & n1581 ;
  assign n19759 = ~n19757 & ~n19758 ;
  assign n19760 = ~\u0_w_reg[2][30]/P0001  & ~n5191 ;
  assign n19761 = \u0_w_reg[2][30]/P0001  & n5191 ;
  assign n19762 = ~n19760 & ~n19761 ;
  assign n19763 = ~\u0_w_reg[1][30]/P0001  & ~n9400 ;
  assign n19764 = \u0_w_reg[1][30]/P0001  & n9400 ;
  assign n19765 = ~n19763 & ~n19764 ;
  assign n19766 = ~\u0_w_reg[3][10]/P0001  & ~n4578 ;
  assign n19767 = \u0_w_reg[3][10]/P0001  & n4578 ;
  assign n19768 = ~n19766 & ~n19767 ;
  assign n19769 = ~\u0_w_reg[0][14]/P0001  & ~n13284 ;
  assign n19770 = \u0_w_reg[0][14]/P0001  & n13284 ;
  assign n19771 = ~n19769 & ~n19770 ;
  assign n19772 = ~\u0_w_reg[0][22]/P0001  & ~n13183 ;
  assign n19773 = \u0_w_reg[0][22]/P0001  & n13183 ;
  assign n19774 = ~n19772 & ~n19773 ;
  assign n19775 = ~\u0_w_reg[3][14]/P0001  & ~n1908 ;
  assign n19776 = \u0_w_reg[3][14]/P0001  & n1908 ;
  assign n19777 = ~n19775 & ~n19776 ;
  assign n19778 = ~\u0_w_reg[3][22]/P0001  & ~n1738 ;
  assign n19779 = \u0_w_reg[3][22]/P0001  & n1738 ;
  assign n19780 = ~n19778 & ~n19779 ;
  assign n19781 = ~\u0_w_reg[2][14]/P0001  & ~n850 ;
  assign n19782 = \u0_w_reg[2][14]/P0001  & n850 ;
  assign n19783 = ~n19781 & ~n19782 ;
  assign n19784 = ~\u0_w_reg[2][22]/P0001  & ~n689 ;
  assign n19785 = \u0_w_reg[2][22]/P0001  & n689 ;
  assign n19786 = ~n19784 & ~n19785 ;
  assign n19787 = ~\u0_w_reg[1][14]/P0001  & ~n9169 ;
  assign n19788 = \u0_w_reg[1][14]/P0001  & n9169 ;
  assign n19789 = ~n19787 & ~n19788 ;
  assign n19790 = ~\u0_w_reg[1][22]/P0001  & ~n9063 ;
  assign n19791 = \u0_w_reg[1][22]/P0001  & n9063 ;
  assign n19792 = ~n19790 & ~n19791 ;
  assign n19793 = ~\u0_w_reg[0][2]/P0001  & ~n15068 ;
  assign n19794 = \u0_w_reg[0][2]/P0001  & n15068 ;
  assign n19795 = ~n19793 & ~n19794 ;
  assign n19796 = ~\u0_w_reg[0][25]/P0001  & ~n13649 ;
  assign n19797 = \u0_w_reg[0][25]/P0001  & n13649 ;
  assign n19798 = ~n19796 & ~n19797 ;
  assign n19799 = ~\u0_w_reg[3][25]/P0001  & ~n3768 ;
  assign n19800 = \u0_w_reg[3][25]/P0001  & n3768 ;
  assign n19801 = ~n19799 & ~n19800 ;
  assign n19802 = ~\u0_w_reg[2][25]/P0001  & ~n6392 ;
  assign n19803 = \u0_w_reg[2][25]/P0001  & n6392 ;
  assign n19804 = ~n19802 & ~n19803 ;
  assign n19805 = ~\u0_w_reg[1][25]/P0001  & ~n10167 ;
  assign n19806 = \u0_w_reg[1][25]/P0001  & n10167 ;
  assign n19807 = ~n19805 & ~n19806 ;
  assign n19808 = ~\u0_w_reg[0][20]/P0001  & ~n11951 ;
  assign n19809 = \u0_w_reg[0][20]/P0001  & n11951 ;
  assign n19810 = ~n19808 & ~n19809 ;
  assign n19811 = ~\u0_w_reg[3][20]/P0001  & ~n2647 ;
  assign n19812 = \u0_w_reg[3][20]/P0001  & n2647 ;
  assign n19813 = ~n19811 & ~n19812 ;
  assign n19814 = ~\u0_w_reg[2][20]/P0001  & ~n5737 ;
  assign n19815 = \u0_w_reg[2][20]/P0001  & n5737 ;
  assign n19816 = ~n19814 & ~n19815 ;
  assign n19817 = ~\u0_w_reg[1][20]/P0001  & ~n8213 ;
  assign n19818 = \u0_w_reg[1][20]/P0001  & n8213 ;
  assign n19819 = ~n19817 & ~n19818 ;
  assign n19820 = ~\u0_w_reg[0][28]/P0001  & ~n12111 ;
  assign n19821 = \u0_w_reg[0][28]/P0001  & n12111 ;
  assign n19822 = ~n19820 & ~n19821 ;
  assign n19823 = ~\u0_w_reg[3][28]/P0001  & ~n2736 ;
  assign n19824 = \u0_w_reg[3][28]/P0001  & n2736 ;
  assign n19825 = ~n19823 & ~n19824 ;
  assign n19826 = ~\u0_w_reg[2][28]/P0001  & ~n5830 ;
  assign n19827 = \u0_w_reg[2][28]/P0001  & n5830 ;
  assign n19828 = ~n19826 & ~n19827 ;
  assign n19829 = ~\u0_w_reg[1][28]/P0001  & ~n8376 ;
  assign n19830 = \u0_w_reg[1][28]/P0001  & n8376 ;
  assign n19831 = ~n19829 & ~n19830 ;
  assign n19832 = \u0_r0_rcnt_reg[0]/P0001  & \u0_r0_rcnt_reg[1]/P0001  ;
  assign n19833 = ~\u0_r0_rcnt_reg[0]/P0001  & ~\u0_r0_rcnt_reg[1]/P0001  ;
  assign n19834 = ~n19832 & ~n19833 ;
  assign n19835 = \u0_r0_rcnt_reg[2]/P0001  & n19832 ;
  assign n19836 = ~\u0_r0_rcnt_reg[2]/P0001  & ~n19832 ;
  assign n19837 = ~n19835 & ~n19836 ;
  assign n19838 = ~\u0_r0_rcnt_reg[3]/P0001  & n19837 ;
  assign n19839 = ~n19834 & n19838 ;
  assign n19840 = \u0_r0_rcnt_reg[3]/P0001  & ~n19835 ;
  assign n19841 = ~\u0_r0_rcnt_reg[3]/P0001  & n19835 ;
  assign n19842 = ~n19840 & ~n19841 ;
  assign n19843 = ~n19834 & ~n19837 ;
  assign n19844 = ~n19842 & n19843 ;
  assign n19845 = ~n19839 & ~n19844 ;
  assign n19846 = ~\u0_r0_rcnt_reg[0]/P0001  & ~n19844 ;
  assign n19847 = ~ld_pad & ~n19846 ;
  assign n19848 = ~n19845 & n19847 ;
  assign n19849 = n19834 & ~n19837 ;
  assign n19850 = n19842 & n19849 ;
  assign n19851 = \u0_r0_rcnt_reg[0]/P0001  & ~n19850 ;
  assign n19852 = n19847 & ~n19851 ;
  assign n19854 = \u0_r0_rcnt_reg[0]/P0001  & ~n19844 ;
  assign n19853 = ~\u0_r0_rcnt_reg[0]/P0001  & ~n19850 ;
  assign n19855 = ~ld_pad & ~n19853 ;
  assign n19856 = ~n19854 & n19855 ;
  assign n19857 = ~ld_pad & ~\u0_r0_rcnt_reg[0]/P0001  ;
  assign n19858 = ~n19845 & n19857 ;
  assign n19859 = ~\u0_r0_rcnt_reg[2]/P0001  & n19833 ;
  assign n19860 = ~n19844 & ~n19859 ;
  assign n19861 = ~ld_pad & ~n19860 ;
  assign n19862 = ~ld_pad & n19834 ;
  assign n19863 = ~\u0_r0_rcnt_reg[0]/P0001  & n19862 ;
  assign n19864 = n19838 & n19863 ;
  assign n19865 = \u0_r0_rcnt_reg[0]/P0001  & n19862 ;
  assign n19866 = n19838 & n19865 ;
  assign n19867 = ~\dcnt_reg[0]/P0001  & ~\dcnt_reg[1]/P0001  ;
  assign n19868 = ~\dcnt_reg[2]/P0001  & n19867 ;
  assign n19869 = \dcnt_reg[3]/P0001  & ~n19868 ;
  assign n19870 = ~ld_pad & ~n19869 ;
  assign n19871 = rst_pad & ~n19870 ;
  assign n19872 = ~ld_pad & ~n19842 ;
  assign n19873 = ~ld_pad & ~n19835 ;
  assign n19874 = \dcnt_reg[2]/P0001  & ~n19867 ;
  assign n19875 = \dcnt_reg[3]/P0001  & n19868 ;
  assign n19876 = ~n19874 & ~n19875 ;
  assign n19877 = ~ld_pad & rst_pad ;
  assign n19878 = ~n19876 & n19877 ;
  assign n19879 = ld_pad & rst_pad ;
  assign n19880 = ~\dcnt_reg[2]/P0001  & ~\dcnt_reg[3]/P0001  ;
  assign n19881 = n19867 & n19880 ;
  assign n19882 = rst_pad & ~n19881 ;
  assign n19883 = ~\dcnt_reg[0]/P0001  & n19882 ;
  assign n19884 = ~n19879 & ~n19883 ;
  assign n19885 = \dcnt_reg[0]/P0001  & \dcnt_reg[1]/P0001  ;
  assign n19886 = ~n19867 & ~n19885 ;
  assign n19887 = n19882 & ~n19886 ;
  assign n19888 = ~n19879 & ~n19887 ;
  assign n19889 = ~ld_pad & n19837 ;
  assign n19890 = \dcnt_reg[0]/P0001  & ~\dcnt_reg[1]/P0001  ;
  assign n19891 = ~ld_pad & n19890 ;
  assign n19892 = n19880 & n19891 ;
  assign n19893 = \u0_w_reg[1][9]/P0001  & ~n11155 ;
  assign n19894 = ~\u0_w_reg[1][9]/P0001  & n11155 ;
  assign n19895 = ~n19893 & ~n19894 ;
  assign n19896 = n10433 & n19895 ;
  assign n19897 = ~n10433 & ~n19895 ;
  assign n19898 = ~n19896 & ~n19897 ;
  assign n19899 = n10170 & n11643 ;
  assign n19900 = ~n10170 & ~n11643 ;
  assign n19901 = ~n19899 & ~n19900 ;
  assign n19903 = n19898 & n19901 ;
  assign n19902 = ~n19898 & ~n19901 ;
  assign n19904 = ~\ld_r_reg/P0001  & ~n19902 ;
  assign n19905 = ~n19903 & n19904 ;
  assign n19907 = \text_in_r_reg[73]/P0001  & \u0_w_reg[1][9]/P0001  ;
  assign n19906 = ~\text_in_r_reg[73]/P0001  & ~\u0_w_reg[1][9]/P0001  ;
  assign n19908 = \ld_r_reg/P0001  & ~n19906 ;
  assign n19909 = ~n19907 & n19908 ;
  assign n19910 = ~n19905 & ~n19909 ;
  assign n19911 = \u0_w_reg[0][0]/P0001  & ~n14033 ;
  assign n19912 = ~\u0_w_reg[0][0]/P0001  & n14033 ;
  assign n19913 = ~n19911 & ~n19912 ;
  assign n19914 = ~n13468 & n14403 ;
  assign n19915 = n13468 & ~n14403 ;
  assign n19916 = ~n19914 & ~n19915 ;
  assign n19918 = n19913 & n19916 ;
  assign n19917 = ~n19913 & ~n19916 ;
  assign n19919 = ~\ld_r_reg/P0001  & ~n19917 ;
  assign n19920 = ~n19918 & n19919 ;
  assign n19922 = ~\text_in_r_reg[96]/P0001  & \u0_w_reg[0][0]/P0001  ;
  assign n19921 = \text_in_r_reg[96]/P0001  & ~\u0_w_reg[0][0]/P0001  ;
  assign n19923 = \ld_r_reg/P0001  & ~n19921 ;
  assign n19924 = ~n19922 & n19923 ;
  assign n19925 = ~n19920 & ~n19924 ;
  assign n19926 = \u0_w_reg[1][0]/P0001  & ~n10430 ;
  assign n19927 = ~\u0_w_reg[1][0]/P0001  & n10430 ;
  assign n19928 = ~n19926 & ~n19927 ;
  assign n19929 = n10251 & n11700 ;
  assign n19930 = ~n10251 & ~n11700 ;
  assign n19931 = ~n19929 & ~n19930 ;
  assign n19933 = n19928 & n19931 ;
  assign n19932 = ~n19928 & ~n19931 ;
  assign n19934 = ~\ld_r_reg/P0001  & ~n19932 ;
  assign n19935 = ~n19933 & n19934 ;
  assign n19937 = ~\text_in_r_reg[64]/P0001  & \u0_w_reg[1][0]/P0001  ;
  assign n19936 = \text_in_r_reg[64]/P0001  & ~\u0_w_reg[1][0]/P0001  ;
  assign n19938 = \ld_r_reg/P0001  & ~n19936 ;
  assign n19939 = ~n19937 & n19938 ;
  assign n19940 = ~n19935 & ~n19939 ;
  assign n19941 = \u0_w_reg[2][0]/P0001  & ~n6657 ;
  assign n19942 = ~\u0_w_reg[2][0]/P0001  & n6657 ;
  assign n19943 = ~n19941 & ~n19942 ;
  assign n19944 = n6475 & n7931 ;
  assign n19945 = ~n6475 & ~n7931 ;
  assign n19946 = ~n19944 & ~n19945 ;
  assign n19948 = n19943 & n19946 ;
  assign n19947 = ~n19943 & ~n19946 ;
  assign n19949 = ~\ld_r_reg/P0001  & ~n19947 ;
  assign n19950 = ~n19948 & n19949 ;
  assign n19952 = ~\text_in_r_reg[32]/P0001  & \u0_w_reg[2][0]/P0001  ;
  assign n19951 = \text_in_r_reg[32]/P0001  & ~\u0_w_reg[2][0]/P0001  ;
  assign n19953 = \ld_r_reg/P0001  & ~n19951 ;
  assign n19954 = ~n19952 & n19953 ;
  assign n19955 = ~n19950 & ~n19954 ;
  assign n19957 = \u0_w_reg[1][24]/P0002  & n16871 ;
  assign n19956 = ~\u0_w_reg[1][24]/P0002  & ~n16871 ;
  assign n19958 = ~ld_pad & ~n19956 ;
  assign n19959 = ~n19957 & n19958 ;
  assign n19960 = \key[88]_pad  & ld_pad ;
  assign n19961 = ~n19959 & ~n19960 ;
  assign n19963 = n15677 & ~n15687 ;
  assign n19962 = ~n15677 & n15687 ;
  assign n19964 = ~ld_pad & ~n19962 ;
  assign n19965 = ~n19963 & n19964 ;
  assign n19966 = \key[93]_pad  & ld_pad ;
  assign n19967 = ~n19965 & ~n19966 ;
  assign \_al_n0  = 1'b0 ;
  assign \_al_n1  = ~1'b0 ;
  assign \g21/_0_  = n1315 ;
  assign \g56610/_0_  = n2092 ;
  assign \g56611/_0_  = n2544 ;
  assign \g56612/_0_  = ~n2957 ;
  assign \g56613/_0_  = n2978 ;
  assign \g56614/_0_  = n3090 ;
  assign \g56615/_0_  = n3108 ;
  assign \g56616/_0_  = ~n3220 ;
  assign \g56617/_0_  = ~n3238 ;
  assign \g56630/_0_  = ~n3783 ;
  assign \g56631/_0_  = ~n3801 ;
  assign \g56632/_0_  = n3981 ;
  assign \g56633/_0_  = n4086 ;
  assign \g56634/_0_  = ~n4263 ;
  assign \g56635/_0_  = n4362 ;
  assign \g56645/_0_  = ~n4593 ;
  assign \g56646/_0_  = ~n4689 ;
  assign \g56647/_0_  = n4707 ;
  assign \g56648/_0_  = n4728 ;
  assign \g56649/_0_  = n4746 ;
  assign \g56650/_0_  = n4770 ;
  assign \g56651/_0_  = ~n4797 ;
  assign \g56652/_0_  = n4884 ;
  assign \g56666/_0_  = n4899 ;
  assign \g56667/_0_  = n4923 ;
  assign \g56668/_0_  = ~n4938 ;
  assign \g56669/_0_  = ~n4956 ;
  assign \g56670/_0_  = ~n4974 ;
  assign \g56671/_0_  = n4992 ;
  assign \g56672/_0_  = n5007 ;
  assign \g56674/_0_  = n5025 ;
  assign \g56675/_0_  = n5040 ;
  assign \g56704/_0_  = ~n5055 ;
  assign \g56739/_0_  = ~n5058 ;
  assign \g56743/_0_  = ~n5061 ;
  assign \g56763/_0_  = ~n5064 ;
  assign \g56776/_0_  = ~n5067 ;
  assign \g56812/_0_  = ~n5070 ;
  assign \g56818/_0_  = ~n5073 ;
  assign \g56861/_0_  = ~n5076 ;
  assign \g56874/_0_  = ~n5079 ;
  assign \g56919/_0_  = ~n5322 ;
  assign \g56920/_0_  = n5646 ;
  assign \g56921/_0_  = n5949 ;
  assign \g56923/_0_  = n5967 ;
  assign \g56924/_0_  = n6076 ;
  assign \g56925/_0_  = ~n6195 ;
  assign \g56926/_0_  = n6213 ;
  assign \g56956/_0_  = ~n6758 ;
  assign \g56957/_0_  = ~n6942 ;
  assign \g56958/_0_  = ~n6960 ;
  assign \g56959/_0_  = n7130 ;
  assign \g56960/_0_  = n7233 ;
  assign \g56961/_0_  = n7334 ;
  assign \g56972/_0_  = ~n7435 ;
  assign \g56973/_0_  = ~n7670 ;
  assign \g56974/_0_  = ~n7691 ;
  assign \g56976/_0_  = n7709 ;
  assign \g56977/_0_  = n7733 ;
  assign \g56978/_0_  = n7751 ;
  assign \g56979/_0_  = n7775 ;
  assign \g56980/_0_  = n7871 ;
  assign \g57008/_0_  = ~n7886 ;
  assign \g57010/_0_  = n7907 ;
  assign \g57011/_0_  = n7925 ;
  assign \g57012/_0_  = ~n7943 ;
  assign \g57013/_0_  = ~n7961 ;
  assign \g57014/_0_  = n7979 ;
  assign \g57015/_0_  = n7994 ;
  assign \g57016/_0_  = n8012 ;
  assign \g57017/_0_  = n8030 ;
  assign \g57086/_0_  = ~n8033 ;
  assign \g57091/_0_  = ~n8036 ;
  assign \g57114/_0_  = ~n8039 ;
  assign \g57129/_0_  = ~n8042 ;
  assign \g57163/_0_  = ~n8045 ;
  assign \g57171/_0_  = ~n8048 ;
  assign \g57204/_0_  = ~n8051 ;
  assign \g57218/_0_  = ~n8054 ;
  assign \g57262/_0_  = n8868 ;
  assign \g57263/_0_  = n9304 ;
  assign \g57264/_0_  = n9418 ;
  assign \g57265/_0_  = n9537 ;
  assign \g57266/_0_  = ~n9654 ;
  assign \g57267/_0_  = n9675 ;
  assign \g57268/_0_  = ~n9693 ;
  assign \g57269/_0_  = n9995 ;
  assign \g57300/_0_  = ~n10523 ;
  assign \g57301/_0_  = n10697 ;
  assign \g57302/_0_  = n10799 ;
  assign \g57303/_0_  = ~n10817 ;
  assign \g57304/_0_  = n10919 ;
  assign \g57316/_0_  = ~n11173 ;
  assign \g57317/_0_  = ~n11399 ;
  assign \g57319/_0_  = ~n11420 ;
  assign \g57320/_0_  = n11438 ;
  assign \g57321/_0_  = n11465 ;
  assign \g57322/_0_  = n11486 ;
  assign \g57323/_0_  = n11580 ;
  assign \g57324/_0_  = n11601 ;
  assign \g57350/_0_  = ~n11619 ;
  assign \g57353/_0_  = n11637 ;
  assign \g57354/_0_  = ~n11658 ;
  assign \g57355/_0_  = n11676 ;
  assign \g57356/_0_  = n11694 ;
  assign \g57357/_0_  = ~n11712 ;
  assign \g57358/_0_  = n11730 ;
  assign \g57359/_0_  = n11748 ;
  assign \g57360/_0_  = n11766 ;
  assign \g57427/_0_  = ~n11769 ;
  assign \g57432/_0_  = ~n11772 ;
  assign \g57456/_0_  = ~n11775 ;
  assign \g57471/_0_  = ~n11778 ;
  assign \g57506/_0_  = ~n11781 ;
  assign \g57512/_0_  = ~n11784 ;
  assign \g57540/_0_  = ~n11787 ;
  assign \g57547/_0_  = ~n11790 ;
  assign \g57654/_0_  = ~n12595 ;
  assign \g57655/_0_  = n12848 ;
  assign \g57656/_0_  = ~n12977 ;
  assign \g57657/_0_  = ~n12995 ;
  assign \g57658/_0_  = ~n13299 ;
  assign \g57676/_0_  = ~n13937 ;
  assign \g57677/_0_  = ~n14225 ;
  assign \g57678/_0_  = ~n14415 ;
  assign \g57679/_0_  = n14816 ;
  assign \g57680/_0_  = n14985 ;
  assign \g57681/_0_  = n15083 ;
  assign \g57682/_0_  = n15101 ;
  assign \g57683/_0_  = n15122 ;
  assign \g57684/_0_  = ~n15143 ;
  assign \g57685/_0_  = n15161 ;
  assign \g57686/_0_  = ~n15176 ;
  assign \g57687/_0_  = ~n15194 ;
  assign \g57688/_0_  = n15218 ;
  assign \g57689/_0_  = n15304 ;
  assign \g57690/_0_  = n15322 ;
  assign \g57691/_0_  = n15346 ;
  assign \g57700/_0_  = ~n15361 ;
  assign \g57701/_0_  = n15379 ;
  assign \g57702/_0_  = ~n15397 ;
  assign \g57703/_0_  = n15412 ;
  assign \g57704/_0_  = n15433 ;
  assign \g57705/_0_  = n15448 ;
  assign \g57706/_0_  = n15466 ;
  assign \g57707/_0_  = n15484 ;
  assign \g57708/_0_  = n15502 ;
  assign \g57709/_3_  = ~n15683 ;
  assign \g57710/_3_  = n15695 ;
  assign \g57711/_0_  = ~n15701 ;
  assign \g57712/_3_  = n15888 ;
  assign \g57715/_3_  = n16009 ;
  assign \g57716/_3_  = n16198 ;
  assign \g57767/_0_  = n16216 ;
  assign \g57768/_3_  = ~n16336 ;
  assign \g57769/_3_  = n16345 ;
  assign \g57770/_3_  = n16351 ;
  assign \g57771/_3_  = ~n16357 ;
  assign \g57777/_3_  = n16474 ;
  assign \g57779/_3_  = n16647 ;
  assign \g57804/_3_  = n16772 ;
  assign \g57805/_3_  = ~n16873 ;
  assign \g57806/_3_  = ~n16970 ;
  assign \g57807/_3_  = ~n17056 ;
  assign \g57808/_3_  = ~n17149 ;
  assign \g57809/_3_  = ~n17158 ;
  assign \g57810/_3_  = ~n17167 ;
  assign \g57811/_3_  = ~n17176 ;
  assign \g57812/_3_  = ~n17188 ;
  assign \g57813/_3_  = n17197 ;
  assign \g57814/_3_  = n17206 ;
  assign \g57815/_3_  = n17215 ;
  assign \g57816/_0_  = ~n17224 ;
  assign \g57817/_3_  = ~n17230 ;
  assign \g57818/_3_  = ~n17236 ;
  assign \g57819/_3_  = ~n17242 ;
  assign \g57822/_3_  = ~n17245 ;
  assign \g57823/_3_  = ~n17251 ;
  assign \g57824/_3_  = ~n17257 ;
  assign \g57830/_3_  = n17369 ;
  assign \g57835/_3_  = ~n17372 ;
  assign \g57836/_3_  = ~n17378 ;
  assign \g57837/_3_  = ~n17384 ;
  assign \g57841/_3_  = ~n17387 ;
  assign \g57842/_3_  = ~n17393 ;
  assign \g57843/_3_  = ~n17399 ;
  assign \g57854/_3_  = n17494 ;
  assign \g57855/_3_  = n17596 ;
  assign \g57856/_3_  = n17704 ;
  assign \g57857/_3_  = n17801 ;
  assign \g57858/_3_  = ~n17894 ;
  assign \g57859/_3_  = n17991 ;
  assign \g57860/_3_  = n18077 ;
  assign \g57861/_3_  = n18161 ;
  assign \g57871/_3_  = n18263 ;
  assign \g57872/_3_  = ~n18364 ;
  assign \g57874/_3_  = n18445 ;
  assign \g57968/_3_  = ~n18533 ;
  assign \g57969/_3_  = ~n18542 ;
  assign \g57970/_3_  = n18551 ;
  assign \g57971/_3_  = ~n18557 ;
  assign \g57980/_3_  = ~n18654 ;
  assign \g57983/_3_  = ~n18657 ;
  assign \g57984/_3_  = ~n18663 ;
  assign \g57985/_3_  = ~n18669 ;
  assign \g58012/_3_  = ~n18672 ;
  assign \g58013/_3_  = ~n18678 ;
  assign \g58015/_3_  = ~n18684 ;
  assign \g58057/_3_  = n18773 ;
  assign \g58058/_3_  = n18862 ;
  assign \g58059/_3_  = n18953 ;
  assign \g58189/_3_  = ~n18956 ;
  assign \g58190/_3_  = ~n18962 ;
  assign \g58191/_3_  = ~n19048 ;
  assign \g58192/_3_  = n19138 ;
  assign \g58193/_3_  = ~n19144 ;
  assign \g58194/_3_  = ~n19234 ;
  assign \g58195/_3_  = ~n19240 ;
  assign \g58196/_3_  = ~n19252 ;
  assign \g58197/_3_  = ~n19261 ;
  assign \g58224/_3_  = ~n19264 ;
  assign \g58226/_3_  = ~n19270 ;
  assign \g58229/_3_  = ~n19276 ;
  assign \g58255/_3_  = ~n19279 ;
  assign \g58256/_3_  = ~n19282 ;
  assign \g58257/_3_  = ~n19285 ;
  assign \g58258/_3_  = ~n19288 ;
  assign \g58259/_3_  = ~n19291 ;
  assign \g58260/_3_  = ~n19297 ;
  assign \g58261/_3_  = ~n19303 ;
  assign \g58262/_3_  = ~n19309 ;
  assign \g58263/_3_  = ~n19315 ;
  assign \g58264/_3_  = ~n19318 ;
  assign \g58265/_3_  = ~n19324 ;
  assign \g58266/_3_  = ~n19330 ;
  assign \g58267/_3_  = ~n19336 ;
  assign \g58268/_3_  = ~n19342 ;
  assign \g58269/_3_  = ~n19348 ;
  assign \g58270/_0_  = ~n19351 ;
  assign \g58271/_3_  = ~n19354 ;
  assign \g58272/_3_  = ~n19357 ;
  assign \g58273/_3_  = ~n19360 ;
  assign \g58274/_3_  = ~n19366 ;
  assign \g58275/_3_  = ~n19372 ;
  assign \g58276/_3_  = ~n19378 ;
  assign \g58277/_3_  = ~n19384 ;
  assign \g58278/_3_  = ~n19390 ;
  assign \g58279/_3_  = ~n19396 ;
  assign \g58285/_3_  = ~n19399 ;
  assign \g58286/_3_  = ~n19402 ;
  assign \g58288/_3_  = ~n19405 ;
  assign \g58289/_3_  = ~n19411 ;
  assign \g58290/_3_  = ~n19414 ;
  assign \g58292/_3_  = ~n19420 ;
  assign \g58294/_3_  = ~n19426 ;
  assign \g58295/_3_  = ~n19432 ;
  assign \g58297/_3_  = ~n19438 ;
  assign \g58330/_0_  = ~n19441 ;
  assign \g58331/_0_  = ~n19444 ;
  assign \g58332/_0_  = ~n19447 ;
  assign \g58333/_0_  = ~n19450 ;
  assign \g58444/_3_  = ~n19453 ;
  assign \g58445/_3_  = ~n19456 ;
  assign \g58446/_3_  = ~n19462 ;
  assign \g58462/_0_  = ~n19465 ;
  assign \g58506/_0_  = ~n19468 ;
  assign \g58507/_0_  = ~n19471 ;
  assign \g58508/_0_  = ~n19474 ;
  assign \g58509/_0_  = ~n19477 ;
  assign \g58531/_0_  = ~n19480 ;
  assign \g58532/_0_  = ~n19483 ;
  assign \g58533/_0_  = ~n19486 ;
  assign \g58550/_0_  = ~n19489 ;
  assign \g58551/_0_  = ~n19492 ;
  assign \g58552/_0_  = ~n19495 ;
  assign \g58553/_0_  = ~n19498 ;
  assign \g58554/_0_  = ~n19501 ;
  assign \g58555/_0_  = ~n19504 ;
  assign \g58556/_0_  = ~n19507 ;
  assign \g58557/_0_  = ~n19510 ;
  assign \g58558/_0_  = ~n19513 ;
  assign \g58559/_0_  = ~n19516 ;
  assign \g58560/_0_  = ~n19519 ;
  assign \g58600/_3_  = ~n19522 ;
  assign \g58601/_3_  = ~n19525 ;
  assign \g58602/_3_  = ~n19528 ;
  assign \g58603/_3_  = ~n19534 ;
  assign \g58604/_3_  = ~n19540 ;
  assign \g58605/_3_  = ~n19546 ;
  assign \g58606/_3_  = ~n19552 ;
  assign \g58607/_3_  = ~n19558 ;
  assign \g58608/_3_  = ~n19564 ;
  assign \g58611/_0_  = ~n19567 ;
  assign \g58612/_0_  = ~n19570 ;
  assign \g58613/_0_  = ~n19573 ;
  assign \g58614/_0_  = ~n19576 ;
  assign \g58617/_0_  = ~n19579 ;
  assign \g58618/_0_  = ~n19582 ;
  assign \g58619/_0_  = ~n19585 ;
  assign \g58634/_0_  = ~n19588 ;
  assign \g58635/_0_  = ~n19591 ;
  assign \g58636/_0_  = ~n19594 ;
  assign \g58637/_0_  = ~n19597 ;
  assign \g58638/_0_  = ~n19600 ;
  assign \g58639/_0_  = ~n19603 ;
  assign \g58640/_0_  = ~n19606 ;
  assign \g58641/_0_  = ~n19609 ;
  assign \g58829/_3_  = ~n19612 ;
  assign \g58830/_3_  = ~n19615 ;
  assign \g58831/_3_  = ~n19618 ;
  assign \g58832/_3_  = ~n19624 ;
  assign \g58833/_3_  = ~n19630 ;
  assign \g58834/_3_  = ~n19636 ;
  assign \g58835/_0_  = ~n19639 ;
  assign \g58844/_0_  = ~n19642 ;
  assign \g58902/_0_  = ~n19645 ;
  assign \g58903/_0_  = ~n19648 ;
  assign \g58904/_0_  = ~n19651 ;
  assign \g58905/_0_  = ~n19654 ;
  assign \g58910/_0_  = ~n19657 ;
  assign \g58913/_0_  = ~n19660 ;
  assign \g58934/_0_  = ~n19663 ;
  assign \g58935/_0_  = ~n19666 ;
  assign \g58936/_0_  = ~n19669 ;
  assign \g58937/_0_  = ~n19672 ;
  assign \g58938/_0_  = ~n19675 ;
  assign \g58970/_0_  = ~n19678 ;
  assign \g58972/_0_  = ~n19681 ;
  assign \g58994/_0_  = ~n19684 ;
  assign \g58995/_0_  = ~n19687 ;
  assign \g58996/_0_  = ~n19690 ;
  assign \g58997/_0_  = ~n19693 ;
  assign \g58998/_0_  = ~n19696 ;
  assign \g58999/_0_  = ~n19699 ;
  assign \g59000/_0_  = ~n19702 ;
  assign \g59002/_0_  = ~n19705 ;
  assign \g59003/_0_  = ~n19708 ;
  assign \g59004/_0_  = ~n19711 ;
  assign \g59254/_0_  = ~n19714 ;
  assign \g59257/_0_  = ~n19717 ;
  assign \g59258/_0_  = ~n19720 ;
  assign \g59259/_0_  = ~n19723 ;
  assign \g59276/_0_  = ~n19726 ;
  assign \g59277/_0_  = ~n19729 ;
  assign \g59278/_0_  = ~n19732 ;
  assign \g59279/_0_  = ~n19735 ;
  assign \g59280/_0_  = ~n19738 ;
  assign \g59291/_0_  = ~n19741 ;
  assign \g59292/_0_  = ~n19744 ;
  assign \g59293/_0_  = ~n19747 ;
  assign \g59294/_0_  = ~n19750 ;
  assign \g59295/_0_  = ~n19753 ;
  assign \g59308/_0_  = ~n19756 ;
  assign \g59309/_0_  = ~n19759 ;
  assign \g59310/_0_  = ~n19762 ;
  assign \g59311/_0_  = ~n19765 ;
  assign \g59330/_0_  = ~n19768 ;
  assign \g59331/_0_  = ~n19771 ;
  assign \g59332/_0_  = ~n19774 ;
  assign \g59333/_0_  = ~n19777 ;
  assign \g59334/_0_  = ~n19780 ;
  assign \g59335/_0_  = ~n19783 ;
  assign \g59336/_0_  = ~n19786 ;
  assign \g59337/_0_  = ~n19789 ;
  assign \g59338/_0_  = ~n19792 ;
  assign \g59339/_0_  = ~n19795 ;
  assign \g59596/_0_  = ~n19798 ;
  assign \g59597/_0_  = ~n19801 ;
  assign \g59598/_0_  = ~n19804 ;
  assign \g59599/_0_  = ~n19807 ;
  assign \g59625/_0_  = ~n19810 ;
  assign \g59626/_0_  = ~n19813 ;
  assign \g59627/_0_  = ~n19816 ;
  assign \g59628/_0_  = ~n19819 ;
  assign \g59837/_0_  = ~n19822 ;
  assign \g59838/_0_  = ~n19825 ;
  assign \g59839/_0_  = ~n19828 ;
  assign \g59840/_0_  = ~n19831 ;
  assign \g60090/_0_  = n19848 ;
  assign \g60320/_0_  = n19852 ;
  assign \g60321/_0_  = n19856 ;
  assign \g60409/_0_  = n19858 ;
  assign \g60539/_0_  = n19861 ;
  assign \g60860/_0_  = n19864 ;
  assign \g60977/_0_  = n19866 ;
  assign \g61012/_0_  = n19871 ;
  assign \g61185/_0_  = n19872 ;
  assign \g61524/_2_  = ~n19873 ;
  assign \g61776/_0_  = n19878 ;
  assign \g61895/_0_  = ~n19884 ;
  assign \g61897/_0_  = ~n19888 ;
  assign \g62220/_0_  = n19889 ;
  assign \g65958/_0_  = n19862 ;
  assign \g72347/_3_  = n19892 ;
  assign \g77848/_0_  = n19857 ;
  assign \g85056/_0_  = ~n19910 ;
  assign \sa30_reg[0]/_05_  = n19925 ;
  assign \sa31_reg[0]/_05_  = n19940 ;
  assign \sa32_reg[0]/_05_  = n19955 ;
  assign \u0_w_reg[1][24]/_05_  = ~n19961 ;
  assign \u0_w_reg[1][29]/_05_  = ~n19967 ;
endmodule
