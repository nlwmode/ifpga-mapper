module top (\P1_B_reg/NET0131 , \P1_IR_reg[0]/NET0131 , \P1_IR_reg[10]/NET0131 , \P1_IR_reg[11]/NET0131 , \P1_IR_reg[12]/NET0131 , \P1_IR_reg[13]/NET0131 , \P1_IR_reg[14]/NET0131 , \P1_IR_reg[15]/NET0131 , \P1_IR_reg[16]/NET0131 , \P1_IR_reg[17]/NET0131 , \P1_IR_reg[18]/NET0131 , \P1_IR_reg[19]/NET0131 , \P1_IR_reg[1]/NET0131 , \P1_IR_reg[20]/NET0131 , \P1_IR_reg[21]/NET0131 , \P1_IR_reg[22]/NET0131 , \P1_IR_reg[23]/NET0131 , \P1_IR_reg[24]/NET0131 , \P1_IR_reg[25]/NET0131 , \P1_IR_reg[26]/NET0131 , \P1_IR_reg[27]/NET0131 , \P1_IR_reg[28]/NET0131 , \P1_IR_reg[29]/NET0131 , \P1_IR_reg[2]/NET0131 , \P1_IR_reg[30]/NET0131 , \P1_IR_reg[31]/NET0131 , \P1_IR_reg[3]/NET0131 , \P1_IR_reg[4]/NET0131 , \P1_IR_reg[5]/NET0131 , \P1_IR_reg[6]/NET0131 , \P1_IR_reg[7]/NET0131 , \P1_IR_reg[8]/NET0131 , \P1_IR_reg[9]/NET0131 , \P1_addr_reg[0]/NET0131 , \P1_addr_reg[10]/NET0131 , \P1_addr_reg[11]/NET0131 , \P1_addr_reg[12]/NET0131 , \P1_addr_reg[13]/NET0131 , \P1_addr_reg[14]/NET0131 , \P1_addr_reg[15]/NET0131 , \P1_addr_reg[16]/NET0131 , \P1_addr_reg[17]/NET0131 , \P1_addr_reg[18]/NET0131 , \P1_addr_reg[19]/NET0131 , \P1_addr_reg[1]/NET0131 , \P1_addr_reg[2]/NET0131 , \P1_addr_reg[3]/NET0131 , \P1_addr_reg[4]/NET0131 , \P1_addr_reg[5]/NET0131 , \P1_addr_reg[6]/NET0131 , \P1_addr_reg[7]/NET0131 , \P1_addr_reg[8]/NET0131 , \P1_addr_reg[9]/NET0131 , \P1_d_reg[0]/NET0131 , \P1_d_reg[1]/NET0131 , \P1_datao_reg[0]/NET0131 , \P1_datao_reg[10]/NET0131 , \P1_datao_reg[11]/NET0131 , \P1_datao_reg[12]/NET0131 , \P1_datao_reg[13]/NET0131 , \P1_datao_reg[14]/NET0131 , \P1_datao_reg[15]/NET0131 , \P1_datao_reg[16]/NET0131 , \P1_datao_reg[17]/NET0131 , \P1_datao_reg[18]/NET0131 , \P1_datao_reg[19]/NET0131 , \P1_datao_reg[1]/NET0131 , \P1_datao_reg[20]/NET0131 , \P1_datao_reg[21]/NET0131 , \P1_datao_reg[22]/NET0131 , \P1_datao_reg[23]/NET0131 , \P1_datao_reg[24]/NET0131 , \P1_datao_reg[25]/NET0131 , \P1_datao_reg[26]/NET0131 , \P1_datao_reg[27]/NET0131 , \P1_datao_reg[28]/NET0131 , \P1_datao_reg[29]/NET0131 , \P1_datao_reg[2]/NET0131 , \P1_datao_reg[30]/NET0131 , \P1_datao_reg[31]/NET0131 , \P1_datao_reg[3]/NET0131 , \P1_datao_reg[4]/NET0131 , \P1_datao_reg[5]/NET0131 , \P1_datao_reg[6]/NET0131 , \P1_datao_reg[7]/NET0131 , \P1_datao_reg[8]/NET0131 , \P1_datao_reg[9]/NET0131 , \P1_rd_reg/NET0131 , \P1_reg0_reg[0]/NET0131 , \P1_reg0_reg[10]/NET0131 , \P1_reg0_reg[11]/NET0131 , \P1_reg0_reg[12]/NET0131 , \P1_reg0_reg[13]/NET0131 , \P1_reg0_reg[14]/NET0131 , \P1_reg0_reg[15]/NET0131 , \P1_reg0_reg[16]/NET0131 , \P1_reg0_reg[17]/NET0131 , \P1_reg0_reg[18]/NET0131 , \P1_reg0_reg[19]/NET0131 , \P1_reg0_reg[1]/NET0131 , \P1_reg0_reg[20]/NET0131 , \P1_reg0_reg[21]/NET0131 , \P1_reg0_reg[22]/NET0131 , \P1_reg0_reg[23]/NET0131 , \P1_reg0_reg[24]/NET0131 , \P1_reg0_reg[25]/NET0131 , \P1_reg0_reg[26]/NET0131 , \P1_reg0_reg[27]/NET0131 , \P1_reg0_reg[28]/NET0131 , \P1_reg0_reg[29]/NET0131 , \P1_reg0_reg[2]/NET0131 , \P1_reg0_reg[30]/NET0131 , \P1_reg0_reg[31]/NET0131 , \P1_reg0_reg[3]/NET0131 , \P1_reg0_reg[4]/NET0131 , \P1_reg0_reg[5]/NET0131 , \P1_reg0_reg[6]/NET0131 , \P1_reg0_reg[7]/NET0131 , \P1_reg0_reg[8]/NET0131 , \P1_reg0_reg[9]/NET0131 , \P1_reg1_reg[0]/NET0131 , \P1_reg1_reg[10]/NET0131 , \P1_reg1_reg[11]/NET0131 , \P1_reg1_reg[12]/NET0131 , \P1_reg1_reg[13]/NET0131 , \P1_reg1_reg[14]/NET0131 , \P1_reg1_reg[15]/NET0131 , \P1_reg1_reg[16]/NET0131 , \P1_reg1_reg[17]/NET0131 , \P1_reg1_reg[18]/NET0131 , \P1_reg1_reg[19]/NET0131 , \P1_reg1_reg[1]/NET0131 , \P1_reg1_reg[20]/NET0131 , \P1_reg1_reg[21]/NET0131 , \P1_reg1_reg[22]/NET0131 , \P1_reg1_reg[23]/NET0131 , \P1_reg1_reg[24]/NET0131 , \P1_reg1_reg[25]/NET0131 , \P1_reg1_reg[26]/NET0131 , \P1_reg1_reg[27]/NET0131 , \P1_reg1_reg[28]/NET0131 , \P1_reg1_reg[29]/NET0131 , \P1_reg1_reg[2]/NET0131 , \P1_reg1_reg[30]/NET0131 , \P1_reg1_reg[31]/NET0131 , \P1_reg1_reg[3]/NET0131 , \P1_reg1_reg[4]/NET0131 , \P1_reg1_reg[5]/NET0131 , \P1_reg1_reg[6]/NET0131 , \P1_reg1_reg[7]/NET0131 , \P1_reg1_reg[8]/NET0131 , \P1_reg1_reg[9]/NET0131 , \P1_reg2_reg[0]/NET0131 , \P1_reg2_reg[10]/NET0131 , \P1_reg2_reg[11]/NET0131 , \P1_reg2_reg[12]/NET0131 , \P1_reg2_reg[13]/NET0131 , \P1_reg2_reg[14]/NET0131 , \P1_reg2_reg[15]/NET0131 , \P1_reg2_reg[16]/NET0131 , \P1_reg2_reg[17]/NET0131 , \P1_reg2_reg[18]/NET0131 , \P1_reg2_reg[19]/NET0131 , \P1_reg2_reg[1]/NET0131 , \P1_reg2_reg[20]/NET0131 , \P1_reg2_reg[21]/NET0131 , \P1_reg2_reg[22]/NET0131 , \P1_reg2_reg[23]/NET0131 , \P1_reg2_reg[24]/NET0131 , \P1_reg2_reg[25]/NET0131 , \P1_reg2_reg[26]/NET0131 , \P1_reg2_reg[27]/NET0131 , \P1_reg2_reg[28]/NET0131 , \P1_reg2_reg[29]/NET0131 , \P1_reg2_reg[2]/NET0131 , \P1_reg2_reg[30]/NET0131 , \P1_reg2_reg[31]/NET0131 , \P1_reg2_reg[3]/NET0131 , \P1_reg2_reg[4]/NET0131 , \P1_reg2_reg[5]/NET0131 , \P1_reg2_reg[6]/NET0131 , \P1_reg2_reg[7]/NET0131 , \P1_reg2_reg[8]/NET0131 , \P1_reg2_reg[9]/NET0131 , \P1_reg3_reg[0]/NET0131 , \P1_reg3_reg[10]/NET0131 , \P1_reg3_reg[11]/NET0131 , \P1_reg3_reg[12]/NET0131 , \P1_reg3_reg[13]/NET0131 , \P1_reg3_reg[14]/NET0131 , \P1_reg3_reg[15]/NET0131 , \P1_reg3_reg[16]/NET0131 , \P1_reg3_reg[17]/NET0131 , \P1_reg3_reg[18]/NET0131 , \P1_reg3_reg[19]/NET0131 , \P1_reg3_reg[1]/NET0131 , \P1_reg3_reg[20]/NET0131 , \P1_reg3_reg[21]/NET0131 , \P1_reg3_reg[22]/NET0131 , \P1_reg3_reg[23]/NET0131 , \P1_reg3_reg[24]/NET0131 , \P1_reg3_reg[25]/NET0131 , \P1_reg3_reg[26]/NET0131 , \P1_reg3_reg[27]/NET0131 , \P1_reg3_reg[28]/NET0131 , \P1_reg3_reg[2]/NET0131 , \P1_reg3_reg[3]/NET0131 , \P1_reg3_reg[4]/NET0131 , \P1_reg3_reg[5]/NET0131 , \P1_reg3_reg[6]/NET0131 , \P1_reg3_reg[7]/NET0131 , \P1_reg3_reg[8]/NET0131 , \P1_reg3_reg[9]/NET0131 , \P1_state_reg[0]/NET0131 , \P1_wr_reg/NET0131 , \P2_B_reg/NET0131 , \P2_IR_reg[0]/NET0131 , \P2_IR_reg[10]/NET0131 , \P2_IR_reg[11]/NET0131 , \P2_IR_reg[12]/NET0131 , \P2_IR_reg[13]/NET0131 , \P2_IR_reg[14]/NET0131 , \P2_IR_reg[15]/NET0131 , \P2_IR_reg[16]/NET0131 , \P2_IR_reg[17]/NET0131 , \P2_IR_reg[18]/NET0131 , \P2_IR_reg[19]/NET0131 , \P2_IR_reg[1]/NET0131 , \P2_IR_reg[20]/NET0131 , \P2_IR_reg[21]/NET0131 , \P2_IR_reg[22]/NET0131 , \P2_IR_reg[23]/NET0131 , \P2_IR_reg[24]/NET0131 , \P2_IR_reg[25]/NET0131 , \P2_IR_reg[26]/NET0131 , \P2_IR_reg[27]/NET0131 , \P2_IR_reg[28]/NET0131 , \P2_IR_reg[29]/NET0131 , \P2_IR_reg[2]/NET0131 , \P2_IR_reg[30]/NET0131 , \P2_IR_reg[31]/NET0131 , \P2_IR_reg[3]/NET0131 , \P2_IR_reg[4]/NET0131 , \P2_IR_reg[5]/NET0131 , \P2_IR_reg[6]/NET0131 , \P2_IR_reg[7]/NET0131 , \P2_IR_reg[8]/NET0131 , \P2_IR_reg[9]/NET0131 , \P2_addr_reg[0]/NET0131 , \P2_addr_reg[10]/NET0131 , \P2_addr_reg[11]/NET0131 , \P2_addr_reg[12]/NET0131 , \P2_addr_reg[13]/NET0131 , \P2_addr_reg[14]/NET0131 , \P2_addr_reg[15]/NET0131 , \P2_addr_reg[16]/NET0131 , \P2_addr_reg[17]/NET0131 , \P2_addr_reg[18]/NET0131 , \P2_addr_reg[19]/NET0131 , \P2_addr_reg[1]/NET0131 , \P2_addr_reg[2]/NET0131 , \P2_addr_reg[3]/NET0131 , \P2_addr_reg[4]/NET0131 , \P2_addr_reg[5]/NET0131 , \P2_addr_reg[6]/NET0131 , \P2_addr_reg[7]/NET0131 , \P2_addr_reg[8]/NET0131 , \P2_addr_reg[9]/NET0131 , \P2_d_reg[0]/NET0131 , \P2_d_reg[1]/NET0131 , \P2_datao_reg[0]/NET0131 , \P2_datao_reg[10]/NET0131 , \P2_datao_reg[11]/NET0131 , \P2_datao_reg[12]/NET0131 , \P2_datao_reg[13]/NET0131 , \P2_datao_reg[14]/NET0131 , \P2_datao_reg[15]/NET0131 , \P2_datao_reg[16]/NET0131 , \P2_datao_reg[17]/NET0131 , \P2_datao_reg[18]/NET0131 , \P2_datao_reg[19]/NET0131 , \P2_datao_reg[1]/NET0131 , \P2_datao_reg[20]/NET0131 , \P2_datao_reg[21]/NET0131 , \P2_datao_reg[22]/NET0131 , \P2_datao_reg[23]/NET0131 , \P2_datao_reg[24]/NET0131 , \P2_datao_reg[25]/NET0131 , \P2_datao_reg[26]/NET0131 , \P2_datao_reg[27]/NET0131 , \P2_datao_reg[28]/NET0131 , \P2_datao_reg[29]/NET0131 , \P2_datao_reg[2]/NET0131 , \P2_datao_reg[30]/NET0131 , \P2_datao_reg[31]/NET0131 , \P2_datao_reg[3]/NET0131 , \P2_datao_reg[4]/NET0131 , \P2_datao_reg[5]/NET0131 , \P2_datao_reg[6]/NET0131 , \P2_datao_reg[7]/NET0131 , \P2_datao_reg[8]/NET0131 , \P2_datao_reg[9]/NET0131 , \P2_rd_reg/NET0131 , \P2_reg0_reg[0]/NET0131 , \P2_reg0_reg[10]/NET0131 , \P2_reg0_reg[11]/NET0131 , \P2_reg0_reg[12]/NET0131 , \P2_reg0_reg[13]/NET0131 , \P2_reg0_reg[14]/NET0131 , \P2_reg0_reg[15]/NET0131 , \P2_reg0_reg[16]/NET0131 , \P2_reg0_reg[17]/NET0131 , \P2_reg0_reg[18]/NET0131 , \P2_reg0_reg[19]/NET0131 , \P2_reg0_reg[1]/NET0131 , \P2_reg0_reg[20]/NET0131 , \P2_reg0_reg[21]/NET0131 , \P2_reg0_reg[22]/NET0131 , \P2_reg0_reg[23]/NET0131 , \P2_reg0_reg[24]/NET0131 , \P2_reg0_reg[25]/NET0131 , \P2_reg0_reg[26]/NET0131 , \P2_reg0_reg[27]/NET0131 , \P2_reg0_reg[28]/NET0131 , \P2_reg0_reg[29]/NET0131 , \P2_reg0_reg[2]/NET0131 , \P2_reg0_reg[30]/NET0131 , \P2_reg0_reg[31]/NET0131 , \P2_reg0_reg[3]/NET0131 , \P2_reg0_reg[4]/NET0131 , \P2_reg0_reg[5]/NET0131 , \P2_reg0_reg[6]/NET0131 , \P2_reg0_reg[7]/NET0131 , \P2_reg0_reg[8]/NET0131 , \P2_reg0_reg[9]/NET0131 , \P2_reg1_reg[0]/NET0131 , \P2_reg1_reg[10]/NET0131 , \P2_reg1_reg[11]/NET0131 , \P2_reg1_reg[12]/NET0131 , \P2_reg1_reg[13]/NET0131 , \P2_reg1_reg[14]/NET0131 , \P2_reg1_reg[15]/NET0131 , \P2_reg1_reg[16]/NET0131 , \P2_reg1_reg[17]/NET0131 , \P2_reg1_reg[18]/NET0131 , \P2_reg1_reg[19]/NET0131 , \P2_reg1_reg[1]/NET0131 , \P2_reg1_reg[20]/NET0131 , \P2_reg1_reg[21]/NET0131 , \P2_reg1_reg[22]/NET0131 , \P2_reg1_reg[23]/NET0131 , \P2_reg1_reg[24]/NET0131 , \P2_reg1_reg[25]/NET0131 , \P2_reg1_reg[26]/NET0131 , \P2_reg1_reg[27]/NET0131 , \P2_reg1_reg[28]/NET0131 , \P2_reg1_reg[29]/NET0131 , \P2_reg1_reg[2]/NET0131 , \P2_reg1_reg[30]/NET0131 , \P2_reg1_reg[31]/NET0131 , \P2_reg1_reg[3]/NET0131 , \P2_reg1_reg[4]/NET0131 , \P2_reg1_reg[5]/NET0131 , \P2_reg1_reg[6]/NET0131 , \P2_reg1_reg[7]/NET0131 , \P2_reg1_reg[8]/NET0131 , \P2_reg1_reg[9]/NET0131 , \P2_reg2_reg[0]/NET0131 , \P2_reg2_reg[10]/NET0131 , \P2_reg2_reg[11]/NET0131 , \P2_reg2_reg[12]/NET0131 , \P2_reg2_reg[13]/NET0131 , \P2_reg2_reg[14]/NET0131 , \P2_reg2_reg[15]/NET0131 , \P2_reg2_reg[16]/NET0131 , \P2_reg2_reg[17]/NET0131 , \P2_reg2_reg[18]/NET0131 , \P2_reg2_reg[19]/NET0131 , \P2_reg2_reg[1]/NET0131 , \P2_reg2_reg[20]/NET0131 , \P2_reg2_reg[21]/NET0131 , \P2_reg2_reg[22]/NET0131 , \P2_reg2_reg[23]/NET0131 , \P2_reg2_reg[24]/NET0131 , \P2_reg2_reg[25]/NET0131 , \P2_reg2_reg[26]/NET0131 , \P2_reg2_reg[27]/NET0131 , \P2_reg2_reg[28]/NET0131 , \P2_reg2_reg[29]/NET0131 , \P2_reg2_reg[2]/NET0131 , \P2_reg2_reg[30]/NET0131 , \P2_reg2_reg[31]/NET0131 , \P2_reg2_reg[3]/NET0131 , \P2_reg2_reg[4]/NET0131 , \P2_reg2_reg[5]/NET0131 , \P2_reg2_reg[6]/NET0131 , \P2_reg2_reg[7]/NET0131 , \P2_reg2_reg[8]/NET0131 , \P2_reg2_reg[9]/NET0131 , \P2_reg3_reg[0]/NET0131 , \P2_reg3_reg[10]/NET0131 , \P2_reg3_reg[11]/NET0131 , \P2_reg3_reg[12]/NET0131 , \P2_reg3_reg[13]/NET0131 , \P2_reg3_reg[14]/NET0131 , \P2_reg3_reg[15]/NET0131 , \P2_reg3_reg[16]/NET0131 , \P2_reg3_reg[17]/NET0131 , \P2_reg3_reg[18]/NET0131 , \P2_reg3_reg[19]/NET0131 , \P2_reg3_reg[1]/NET0131 , \P2_reg3_reg[20]/NET0131 , \P2_reg3_reg[21]/NET0131 , \P2_reg3_reg[22]/NET0131 , \P2_reg3_reg[23]/NET0131 , \P2_reg3_reg[24]/NET0131 , \P2_reg3_reg[25]/NET0131 , \P2_reg3_reg[26]/NET0131 , \P2_reg3_reg[27]/NET0131 , \P2_reg3_reg[28]/NET0131 , \P2_reg3_reg[2]/NET0131 , \P2_reg3_reg[3]/NET0131 , \P2_reg3_reg[4]/NET0131 , \P2_reg3_reg[5]/NET0131 , \P2_reg3_reg[6]/NET0131 , \P2_reg3_reg[7]/NET0131 , \P2_reg3_reg[8]/NET0131 , \P2_reg3_reg[9]/NET0131 , \P2_wr_reg/NET0131 , \si[0]_pad , \si[10]_pad , \si[11]_pad , \si[12]_pad , \si[13]_pad , \si[14]_pad , \si[15]_pad , \si[16]_pad , \si[17]_pad , \si[18]_pad , \si[19]_pad , \si[1]_pad , \si[20]_pad , \si[21]_pad , \si[22]_pad , \si[23]_pad , \si[24]_pad , \si[25]_pad , \si[26]_pad , \si[27]_pad , \si[28]_pad , \si[29]_pad , \si[2]_pad , \si[30]_pad , \si[31]_pad , \si[3]_pad , \si[4]_pad , \si[5]_pad , \si[6]_pad , \si[7]_pad , \si[8]_pad , \si[9]_pad , \P1_state_reg[0]/NET0131_syn_2 , \_al_n0 , \_al_n1 , \g21_dup/_0_ , \g71037/_0_ , \g71048/_0_ , \g71049/_0_ , \g71050/_0_ , \g71052/_0_ , \g71053/_0_ , \g71054/_0_ , \g71055/_0_ , \g71080/_0_ , \g71081/_0_ , \g71082/_0_ , \g71084/_0_ , \g71085/_0_ , \g71086/_0_ , \g71087/_0_ , \g71088/_0_ , \g71089/_0_ , \g71121/_0_ , \g71122/_0_ , \g71123/_0_ , \g71130/_0_ , \g71131/_0_ , \g71132/_0_ , \g71135/_0_ , \g71136/_0_ , \g71137/_0_ , \g71138/_0_ , \g71139/_0_ , \g71141/_0_ , \g71142/_0_ , \g71143/_0_ , \g71144/_0_ , \g71145/_0_ , \g71146/_0_ , \g71147/_0_ , \g71179/_0_ , \g71186/_0_ , \g71194/_0_ , \g71195/_0_ , \g71196/_0_ , \g71197/_0_ , \g71200/_0_ , \g71201/_0_ , \g71202/_0_ , \g71203/_0_ , \g71204/_0_ , \g71205/_0_ , \g71206/_0_ , \g71207/_0_ , \g71208/_0_ , \g71209/_0_ , \g71210/_0_ , \g71211/_0_ , \g71212/_0_ , \g71213/_0_ , \g71214/_0_ , \g71215/_0_ , \g71262/_0_ , \g71263/_0_ , \g71264/_0_ , \g71291/_0_ , \g71294/_0_ , \g71295/_0_ , \g71296/_0_ , \g71297/_0_ , \g71298/_0_ , \g71299/_0_ , \g71300/_0_ , \g71302/_0_ , \g71303/_0_ , \g71304/_0_ , \g71305/_0_ , \g71306/_0_ , \g71307/_0_ , \g71308/_0_ , \g71354/_0_ , \g71359/_0_ , \g71400/_0_ , \g71401/_0_ , \g71402/_0_ , \g71403/_0_ , \g71404/_0_ , \g71405/_0_ , \g71406/_0_ , \g71407/_0_ , \g71408/_0_ , \g71409/_0_ , \g71410/_0_ , \g71411/_0_ , \g71412/_0_ , \g71413/_0_ , \g71414/_0_ , \g71415/_0_ , \g71416/_0_ , \g71417/_0_ , \g71418/_0_ , \g71420/_0_ , \g71421/_0_ , \g71422/_0_ , \g71423/_0_ , \g71424/_0_ , \g71484/_0_ , \g71485/_0_ , \g71486/_0_ , \g71488/_0_ , \g71489/_0_ , \g71490/_0_ , \g71492/_0_ , \g71493/_0_ , \g71537/_0_ , \g71538/_0_ , \g71539/_0_ , \g71540/_0_ , \g71541/_0_ , \g71542/_0_ , \g71543/_0_ , \g71544/_0_ , \g71545/_0_ , \g71546/_0_ , \g71547/_0_ , \g71548/_0_ , \g71549/_0_ , \g71550/_0_ , \g71551/_0_ , \g71552/_0_ , \g71553/_0_ , \g71554/_0_ , \g71555/_0_ , \g71608/_0_ , \g71609/_0_ , \g71613/_0_ , \g71615/_0_ , \g71617/_0_ , \g71619/_0_ , \g71620/_0_ , \g71621/_0_ , \g71690/_0_ , \g71691/_0_ , \g71692/_0_ , \g71693/_0_ , \g71694/_0_ , \g71696/_0_ , \g71697/_0_ , \g71698/_0_ , \g71699/_0_ , \g71700/_0_ , \g71701/_0_ , \g71702/_0_ , \g71703/_0_ , \g71704/_0_ , \g71705/_0_ , \g71707/_0_ , \g71708/_0_ , \g71709/_0_ , \g71710/_0_ , \g71711/_0_ , \g71712/_0_ , \g71713/_0_ , \g71788/_0_ , \g71789/_0_ , \g71792/_0_ , \g71793/_0_ , \g71794/_0_ , \g71859/_0_ , \g71860/_0_ , \g71861/_0_ , \g71862/_0_ , \g71863/_0_ , \g71864/_0_ , \g71865/_0_ , \g71866/_0_ , \g71867/_0_ , \g71868/_0_ , \g71869/_0_ , \g71870/_0_ , \g71871/_0_ , \g71872/_0_ , \g71873/_0_ , \g71874/_0_ , \g71875/_0_ , \g71876/_0_ , \g71877/_0_ , \g71878/_0_ , \g71879/_0_ , \g71918/_0_ , \g71921/_0_ , \g72042/_0_ , \g72045/_0_ , \g72046/_0_ , \g72047/_0_ , \g72048/_0_ , \g72049/_0_ , \g72050/_0_ , \g72051/_0_ , \g72052/_0_ , \g72053/_0_ , \g72054/_0_ , \g72055/_0_ , \g72056/_0_ , \g72059/_0_ , \g72060/_0_ , \g72061/_0_ , \g72062/_0_ , \g72063/_0_ , \g72064/_0_ , \g72065/_0_ , \g72185/_0_ , \g72302/_0_ , \g72304/_0_ , \g72468/_0_ , \g72577/_0_ , \g72578/_0_ , \g72579/_0_ , \g72580/_0_ , \g72585/_0_ , \g72742/_0_ , \g72758/_0_ , \g72947/_0_ , \g72948/_0_ , \g72952/_0_ , \g72954/_0_ , \g72955/_0_ , \g72956/_0_ , \g72957/_0_ , \g73346/_0_ , \g73349/_0_ , \g73350/_0_ , \g73357/_0_ , \g73618/_0_ , \g74419/_0_ , \g74422/_0_ , \g74426/_0_ , \g74671/_0_ , \g75421/_0_ , \g75424/_0_ , \g75430/_0_ , \g76173/_0_ , \g76175/_0_ , \g76177/_0_ , \g76178/_0_ , \g76179/_0_ , \g76506/_0_ , \g80645/_3_ , \g80646/_3_ , \g80647/_3_ , \g80648/_3_ , \g80649/_0_ , \g80650/_0_ , \g80952/_0_ , \g80956/_0_ , \g80957/_0_ , \g80958/_0_ , \g80959/_0_ , \g80960/_0_ , \g80961/_0_ , \g80962/_0_ , \g80963/_0_ , \g80964/_0_ , \g80965/_0_ , \g80966/_3_ , \g80967/_0_ , \g80968/_0_ , \g80969/_0_ , \g80970/_0_ , \g80971/_0_ , \g80972/_0_ , \g80973/_0_ , \g80974/_3_ , \g80975/_0_ , \g80976/_0_ , \g80977/_0_ , \g80978/_3_ , \g80979/_0_ , \g80980/_0_ , \g80981/_0_ , \g80982/_3_ , \g81025/_3_ , \g81026/_3_ , \g81027/_3_ , \g81028/_3_ , \g81029/_3_ , \g81030/_3_ , \g81031/_3_ , \g81032/_3_ , \g81033/_3_ , \g81034/_3_ , \g81035/_3_ , \g81036/_3_ , \g81037/_3_ , \g81038/_3_ , \g81039/_3_ , \g81040/_3_ , \g81041/_3_ , \g81042/_3_ , \g81043/_0_ , \g81044/_3_ , \g81045/_0_ , \g81046/_3_ , \g81047/_3_ , \g81048/_0_ , \g81049/_3_ , \g81050/_3_ , \g81051/_3_ , \g81052/_3_ , \g81524/_0_ , \g81534/_0_ , \g82411/_0_ , \g82413/_0_ , \g82414/_0_ , \g82415/_0_ , \g82416/_0_ , \g82417/_0_ , \g82418/_0_ , \g82419/_0_ , \g82420/_0_ , \g82421/_0_ , \g82422/_0_ , \g82423/_0_ , \g82424/_0_ , \g82425/_0_ , \g82426/_0_ , \g82427/_0_ , \g82428/_0_ , \g82429/_0_ , \g82430/_0_ , \g82432/_0_ , \g82435/_0_ , \g82436/_0_ , \g83031/u3_syn_4 , \g83221/_0_ , \g83364/_0_ , \g83474/_0_ , \g83478/_0_ , \g83479/_0_ , \g83480/_0_ , \g83481/_0_ , \g83482/_0_ , \g83484/_0_ , \g83486/_0_ , \g83487/_0_ , \g83488/_0_ , \g83489/_0_ , \g83490/_0_ , \g83491/_0_ , \g83492/_0_ , \g83493/_0_ , \g83494/_0_ , \g83495/_0_ , \g83496/_0_ , \g83505/_0_ , \g83622/u3_syn_4 , \g83853/_0_ , \g83905/_0_ , \g84145/u3_syn_4 , \g84148/u3_syn_4 , \g85427/_2_ , \g85433/_0_ , \g85458/_0_ , \g85512/_0_ , \g85517/_0_ , \g85963/_0_ , \g85996/_0_ , \g86064/_0_ , \g86079/_0_ , \g86088/_0_ , \g86096/_0_ , \g86107/_0_ , \g86159/_0_ , \g86232_dup/_0_ , \g86249/_0_ , \g86258/_0_ , \g86268/_0_ , \g86278/_0_ , \g86281/_0_ , \g86293/_0_ , \g86305/_0_ , \g86313/_0_ , \g86329/_0_ , \g86338/_0_ , \g86355/_0_ , \g86362/_0_ , \g86375/_0_ , \g86385/_0_ , \g86394/_0_ , \g86405/_0_ , \g86413/_0_ , \g86425/_0_ , \g86433_dup/_0_ , \g86441/_0_ , \g86448/_0_ , \g86484/_0_ , \g86493/_0_ , \g86501/_0_ , \g86509/_0_ , \g86518/_0_ , \g86527/_0_ , \g86531/_0_ , \g86541/_0_ , \g86549/_0_ , \g86577/_0_ , \g86598/_0_ , \g86607/_0_ , \g87968/_0_ , \g93740/_0_ , \g93779/_0_ , \g93782/_0_ , \g93859/_0_ , \g93950/_0_ , \g93972/_0_ , \g94026/_0_ , \g94078/_0_ , \g94095/_0_ , \g94136/_0_ , \g94238/_0_ , \g94252/_0_ , \g94278/_0_ , \g94380/_0_ , \g94545/_0_ , \g94586/_0_ , \g94640/_0_ , \g94710/_0_ , \g94743/_0_ , \g94877/_0_ , \g95093/_0_ , \g95139/_0_ , \g95161/_0_ , \g95165/_0_ , \g95204/_0_ , \g95395/_0_ , \g95447/_0_ , rd_pad, \so[0]_pad , \so[10]_pad , \so[11]_pad , \so[12]_pad , \so[13]_pad , \so[14]_pad , \so[15]_pad , \so[16]_pad , \so[17]_pad , \so[18]_pad , \so[19]_pad , \so[1]_pad , \so[2]_pad , \so[3]_pad , \so[4]_pad , \so[5]_pad , \so[6]_pad , \so[7]_pad , \so[8]_pad , \so[9]_pad , wr_pad);
	input \P1_B_reg/NET0131  ;
	input \P1_IR_reg[0]/NET0131  ;
	input \P1_IR_reg[10]/NET0131  ;
	input \P1_IR_reg[11]/NET0131  ;
	input \P1_IR_reg[12]/NET0131  ;
	input \P1_IR_reg[13]/NET0131  ;
	input \P1_IR_reg[14]/NET0131  ;
	input \P1_IR_reg[15]/NET0131  ;
	input \P1_IR_reg[16]/NET0131  ;
	input \P1_IR_reg[17]/NET0131  ;
	input \P1_IR_reg[18]/NET0131  ;
	input \P1_IR_reg[19]/NET0131  ;
	input \P1_IR_reg[1]/NET0131  ;
	input \P1_IR_reg[20]/NET0131  ;
	input \P1_IR_reg[21]/NET0131  ;
	input \P1_IR_reg[22]/NET0131  ;
	input \P1_IR_reg[23]/NET0131  ;
	input \P1_IR_reg[24]/NET0131  ;
	input \P1_IR_reg[25]/NET0131  ;
	input \P1_IR_reg[26]/NET0131  ;
	input \P1_IR_reg[27]/NET0131  ;
	input \P1_IR_reg[28]/NET0131  ;
	input \P1_IR_reg[29]/NET0131  ;
	input \P1_IR_reg[2]/NET0131  ;
	input \P1_IR_reg[30]/NET0131  ;
	input \P1_IR_reg[31]/NET0131  ;
	input \P1_IR_reg[3]/NET0131  ;
	input \P1_IR_reg[4]/NET0131  ;
	input \P1_IR_reg[5]/NET0131  ;
	input \P1_IR_reg[6]/NET0131  ;
	input \P1_IR_reg[7]/NET0131  ;
	input \P1_IR_reg[8]/NET0131  ;
	input \P1_IR_reg[9]/NET0131  ;
	input \P1_addr_reg[0]/NET0131  ;
	input \P1_addr_reg[10]/NET0131  ;
	input \P1_addr_reg[11]/NET0131  ;
	input \P1_addr_reg[12]/NET0131  ;
	input \P1_addr_reg[13]/NET0131  ;
	input \P1_addr_reg[14]/NET0131  ;
	input \P1_addr_reg[15]/NET0131  ;
	input \P1_addr_reg[16]/NET0131  ;
	input \P1_addr_reg[17]/NET0131  ;
	input \P1_addr_reg[18]/NET0131  ;
	input \P1_addr_reg[19]/NET0131  ;
	input \P1_addr_reg[1]/NET0131  ;
	input \P1_addr_reg[2]/NET0131  ;
	input \P1_addr_reg[3]/NET0131  ;
	input \P1_addr_reg[4]/NET0131  ;
	input \P1_addr_reg[5]/NET0131  ;
	input \P1_addr_reg[6]/NET0131  ;
	input \P1_addr_reg[7]/NET0131  ;
	input \P1_addr_reg[8]/NET0131  ;
	input \P1_addr_reg[9]/NET0131  ;
	input \P1_d_reg[0]/NET0131  ;
	input \P1_d_reg[1]/NET0131  ;
	input \P1_datao_reg[0]/NET0131  ;
	input \P1_datao_reg[10]/NET0131  ;
	input \P1_datao_reg[11]/NET0131  ;
	input \P1_datao_reg[12]/NET0131  ;
	input \P1_datao_reg[13]/NET0131  ;
	input \P1_datao_reg[14]/NET0131  ;
	input \P1_datao_reg[15]/NET0131  ;
	input \P1_datao_reg[16]/NET0131  ;
	input \P1_datao_reg[17]/NET0131  ;
	input \P1_datao_reg[18]/NET0131  ;
	input \P1_datao_reg[19]/NET0131  ;
	input \P1_datao_reg[1]/NET0131  ;
	input \P1_datao_reg[20]/NET0131  ;
	input \P1_datao_reg[21]/NET0131  ;
	input \P1_datao_reg[22]/NET0131  ;
	input \P1_datao_reg[23]/NET0131  ;
	input \P1_datao_reg[24]/NET0131  ;
	input \P1_datao_reg[25]/NET0131  ;
	input \P1_datao_reg[26]/NET0131  ;
	input \P1_datao_reg[27]/NET0131  ;
	input \P1_datao_reg[28]/NET0131  ;
	input \P1_datao_reg[29]/NET0131  ;
	input \P1_datao_reg[2]/NET0131  ;
	input \P1_datao_reg[30]/NET0131  ;
	input \P1_datao_reg[31]/NET0131  ;
	input \P1_datao_reg[3]/NET0131  ;
	input \P1_datao_reg[4]/NET0131  ;
	input \P1_datao_reg[5]/NET0131  ;
	input \P1_datao_reg[6]/NET0131  ;
	input \P1_datao_reg[7]/NET0131  ;
	input \P1_datao_reg[8]/NET0131  ;
	input \P1_datao_reg[9]/NET0131  ;
	input \P1_rd_reg/NET0131  ;
	input \P1_reg0_reg[0]/NET0131  ;
	input \P1_reg0_reg[10]/NET0131  ;
	input \P1_reg0_reg[11]/NET0131  ;
	input \P1_reg0_reg[12]/NET0131  ;
	input \P1_reg0_reg[13]/NET0131  ;
	input \P1_reg0_reg[14]/NET0131  ;
	input \P1_reg0_reg[15]/NET0131  ;
	input \P1_reg0_reg[16]/NET0131  ;
	input \P1_reg0_reg[17]/NET0131  ;
	input \P1_reg0_reg[18]/NET0131  ;
	input \P1_reg0_reg[19]/NET0131  ;
	input \P1_reg0_reg[1]/NET0131  ;
	input \P1_reg0_reg[20]/NET0131  ;
	input \P1_reg0_reg[21]/NET0131  ;
	input \P1_reg0_reg[22]/NET0131  ;
	input \P1_reg0_reg[23]/NET0131  ;
	input \P1_reg0_reg[24]/NET0131  ;
	input \P1_reg0_reg[25]/NET0131  ;
	input \P1_reg0_reg[26]/NET0131  ;
	input \P1_reg0_reg[27]/NET0131  ;
	input \P1_reg0_reg[28]/NET0131  ;
	input \P1_reg0_reg[29]/NET0131  ;
	input \P1_reg0_reg[2]/NET0131  ;
	input \P1_reg0_reg[30]/NET0131  ;
	input \P1_reg0_reg[31]/NET0131  ;
	input \P1_reg0_reg[3]/NET0131  ;
	input \P1_reg0_reg[4]/NET0131  ;
	input \P1_reg0_reg[5]/NET0131  ;
	input \P1_reg0_reg[6]/NET0131  ;
	input \P1_reg0_reg[7]/NET0131  ;
	input \P1_reg0_reg[8]/NET0131  ;
	input \P1_reg0_reg[9]/NET0131  ;
	input \P1_reg1_reg[0]/NET0131  ;
	input \P1_reg1_reg[10]/NET0131  ;
	input \P1_reg1_reg[11]/NET0131  ;
	input \P1_reg1_reg[12]/NET0131  ;
	input \P1_reg1_reg[13]/NET0131  ;
	input \P1_reg1_reg[14]/NET0131  ;
	input \P1_reg1_reg[15]/NET0131  ;
	input \P1_reg1_reg[16]/NET0131  ;
	input \P1_reg1_reg[17]/NET0131  ;
	input \P1_reg1_reg[18]/NET0131  ;
	input \P1_reg1_reg[19]/NET0131  ;
	input \P1_reg1_reg[1]/NET0131  ;
	input \P1_reg1_reg[20]/NET0131  ;
	input \P1_reg1_reg[21]/NET0131  ;
	input \P1_reg1_reg[22]/NET0131  ;
	input \P1_reg1_reg[23]/NET0131  ;
	input \P1_reg1_reg[24]/NET0131  ;
	input \P1_reg1_reg[25]/NET0131  ;
	input \P1_reg1_reg[26]/NET0131  ;
	input \P1_reg1_reg[27]/NET0131  ;
	input \P1_reg1_reg[28]/NET0131  ;
	input \P1_reg1_reg[29]/NET0131  ;
	input \P1_reg1_reg[2]/NET0131  ;
	input \P1_reg1_reg[30]/NET0131  ;
	input \P1_reg1_reg[31]/NET0131  ;
	input \P1_reg1_reg[3]/NET0131  ;
	input \P1_reg1_reg[4]/NET0131  ;
	input \P1_reg1_reg[5]/NET0131  ;
	input \P1_reg1_reg[6]/NET0131  ;
	input \P1_reg1_reg[7]/NET0131  ;
	input \P1_reg1_reg[8]/NET0131  ;
	input \P1_reg1_reg[9]/NET0131  ;
	input \P1_reg2_reg[0]/NET0131  ;
	input \P1_reg2_reg[10]/NET0131  ;
	input \P1_reg2_reg[11]/NET0131  ;
	input \P1_reg2_reg[12]/NET0131  ;
	input \P1_reg2_reg[13]/NET0131  ;
	input \P1_reg2_reg[14]/NET0131  ;
	input \P1_reg2_reg[15]/NET0131  ;
	input \P1_reg2_reg[16]/NET0131  ;
	input \P1_reg2_reg[17]/NET0131  ;
	input \P1_reg2_reg[18]/NET0131  ;
	input \P1_reg2_reg[19]/NET0131  ;
	input \P1_reg2_reg[1]/NET0131  ;
	input \P1_reg2_reg[20]/NET0131  ;
	input \P1_reg2_reg[21]/NET0131  ;
	input \P1_reg2_reg[22]/NET0131  ;
	input \P1_reg2_reg[23]/NET0131  ;
	input \P1_reg2_reg[24]/NET0131  ;
	input \P1_reg2_reg[25]/NET0131  ;
	input \P1_reg2_reg[26]/NET0131  ;
	input \P1_reg2_reg[27]/NET0131  ;
	input \P1_reg2_reg[28]/NET0131  ;
	input \P1_reg2_reg[29]/NET0131  ;
	input \P1_reg2_reg[2]/NET0131  ;
	input \P1_reg2_reg[30]/NET0131  ;
	input \P1_reg2_reg[31]/NET0131  ;
	input \P1_reg2_reg[3]/NET0131  ;
	input \P1_reg2_reg[4]/NET0131  ;
	input \P1_reg2_reg[5]/NET0131  ;
	input \P1_reg2_reg[6]/NET0131  ;
	input \P1_reg2_reg[7]/NET0131  ;
	input \P1_reg2_reg[8]/NET0131  ;
	input \P1_reg2_reg[9]/NET0131  ;
	input \P1_reg3_reg[0]/NET0131  ;
	input \P1_reg3_reg[10]/NET0131  ;
	input \P1_reg3_reg[11]/NET0131  ;
	input \P1_reg3_reg[12]/NET0131  ;
	input \P1_reg3_reg[13]/NET0131  ;
	input \P1_reg3_reg[14]/NET0131  ;
	input \P1_reg3_reg[15]/NET0131  ;
	input \P1_reg3_reg[16]/NET0131  ;
	input \P1_reg3_reg[17]/NET0131  ;
	input \P1_reg3_reg[18]/NET0131  ;
	input \P1_reg3_reg[19]/NET0131  ;
	input \P1_reg3_reg[1]/NET0131  ;
	input \P1_reg3_reg[20]/NET0131  ;
	input \P1_reg3_reg[21]/NET0131  ;
	input \P1_reg3_reg[22]/NET0131  ;
	input \P1_reg3_reg[23]/NET0131  ;
	input \P1_reg3_reg[24]/NET0131  ;
	input \P1_reg3_reg[25]/NET0131  ;
	input \P1_reg3_reg[26]/NET0131  ;
	input \P1_reg3_reg[27]/NET0131  ;
	input \P1_reg3_reg[28]/NET0131  ;
	input \P1_reg3_reg[2]/NET0131  ;
	input \P1_reg3_reg[3]/NET0131  ;
	input \P1_reg3_reg[4]/NET0131  ;
	input \P1_reg3_reg[5]/NET0131  ;
	input \P1_reg3_reg[6]/NET0131  ;
	input \P1_reg3_reg[7]/NET0131  ;
	input \P1_reg3_reg[8]/NET0131  ;
	input \P1_reg3_reg[9]/NET0131  ;
	input \P1_state_reg[0]/NET0131  ;
	input \P1_wr_reg/NET0131  ;
	input \P2_B_reg/NET0131  ;
	input \P2_IR_reg[0]/NET0131  ;
	input \P2_IR_reg[10]/NET0131  ;
	input \P2_IR_reg[11]/NET0131  ;
	input \P2_IR_reg[12]/NET0131  ;
	input \P2_IR_reg[13]/NET0131  ;
	input \P2_IR_reg[14]/NET0131  ;
	input \P2_IR_reg[15]/NET0131  ;
	input \P2_IR_reg[16]/NET0131  ;
	input \P2_IR_reg[17]/NET0131  ;
	input \P2_IR_reg[18]/NET0131  ;
	input \P2_IR_reg[19]/NET0131  ;
	input \P2_IR_reg[1]/NET0131  ;
	input \P2_IR_reg[20]/NET0131  ;
	input \P2_IR_reg[21]/NET0131  ;
	input \P2_IR_reg[22]/NET0131  ;
	input \P2_IR_reg[23]/NET0131  ;
	input \P2_IR_reg[24]/NET0131  ;
	input \P2_IR_reg[25]/NET0131  ;
	input \P2_IR_reg[26]/NET0131  ;
	input \P2_IR_reg[27]/NET0131  ;
	input \P2_IR_reg[28]/NET0131  ;
	input \P2_IR_reg[29]/NET0131  ;
	input \P2_IR_reg[2]/NET0131  ;
	input \P2_IR_reg[30]/NET0131  ;
	input \P2_IR_reg[31]/NET0131  ;
	input \P2_IR_reg[3]/NET0131  ;
	input \P2_IR_reg[4]/NET0131  ;
	input \P2_IR_reg[5]/NET0131  ;
	input \P2_IR_reg[6]/NET0131  ;
	input \P2_IR_reg[7]/NET0131  ;
	input \P2_IR_reg[8]/NET0131  ;
	input \P2_IR_reg[9]/NET0131  ;
	input \P2_addr_reg[0]/NET0131  ;
	input \P2_addr_reg[10]/NET0131  ;
	input \P2_addr_reg[11]/NET0131  ;
	input \P2_addr_reg[12]/NET0131  ;
	input \P2_addr_reg[13]/NET0131  ;
	input \P2_addr_reg[14]/NET0131  ;
	input \P2_addr_reg[15]/NET0131  ;
	input \P2_addr_reg[16]/NET0131  ;
	input \P2_addr_reg[17]/NET0131  ;
	input \P2_addr_reg[18]/NET0131  ;
	input \P2_addr_reg[19]/NET0131  ;
	input \P2_addr_reg[1]/NET0131  ;
	input \P2_addr_reg[2]/NET0131  ;
	input \P2_addr_reg[3]/NET0131  ;
	input \P2_addr_reg[4]/NET0131  ;
	input \P2_addr_reg[5]/NET0131  ;
	input \P2_addr_reg[6]/NET0131  ;
	input \P2_addr_reg[7]/NET0131  ;
	input \P2_addr_reg[8]/NET0131  ;
	input \P2_addr_reg[9]/NET0131  ;
	input \P2_d_reg[0]/NET0131  ;
	input \P2_d_reg[1]/NET0131  ;
	input \P2_datao_reg[0]/NET0131  ;
	input \P2_datao_reg[10]/NET0131  ;
	input \P2_datao_reg[11]/NET0131  ;
	input \P2_datao_reg[12]/NET0131  ;
	input \P2_datao_reg[13]/NET0131  ;
	input \P2_datao_reg[14]/NET0131  ;
	input \P2_datao_reg[15]/NET0131  ;
	input \P2_datao_reg[16]/NET0131  ;
	input \P2_datao_reg[17]/NET0131  ;
	input \P2_datao_reg[18]/NET0131  ;
	input \P2_datao_reg[19]/NET0131  ;
	input \P2_datao_reg[1]/NET0131  ;
	input \P2_datao_reg[20]/NET0131  ;
	input \P2_datao_reg[21]/NET0131  ;
	input \P2_datao_reg[22]/NET0131  ;
	input \P2_datao_reg[23]/NET0131  ;
	input \P2_datao_reg[24]/NET0131  ;
	input \P2_datao_reg[25]/NET0131  ;
	input \P2_datao_reg[26]/NET0131  ;
	input \P2_datao_reg[27]/NET0131  ;
	input \P2_datao_reg[28]/NET0131  ;
	input \P2_datao_reg[29]/NET0131  ;
	input \P2_datao_reg[2]/NET0131  ;
	input \P2_datao_reg[30]/NET0131  ;
	input \P2_datao_reg[31]/NET0131  ;
	input \P2_datao_reg[3]/NET0131  ;
	input \P2_datao_reg[4]/NET0131  ;
	input \P2_datao_reg[5]/NET0131  ;
	input \P2_datao_reg[6]/NET0131  ;
	input \P2_datao_reg[7]/NET0131  ;
	input \P2_datao_reg[8]/NET0131  ;
	input \P2_datao_reg[9]/NET0131  ;
	input \P2_rd_reg/NET0131  ;
	input \P2_reg0_reg[0]/NET0131  ;
	input \P2_reg0_reg[10]/NET0131  ;
	input \P2_reg0_reg[11]/NET0131  ;
	input \P2_reg0_reg[12]/NET0131  ;
	input \P2_reg0_reg[13]/NET0131  ;
	input \P2_reg0_reg[14]/NET0131  ;
	input \P2_reg0_reg[15]/NET0131  ;
	input \P2_reg0_reg[16]/NET0131  ;
	input \P2_reg0_reg[17]/NET0131  ;
	input \P2_reg0_reg[18]/NET0131  ;
	input \P2_reg0_reg[19]/NET0131  ;
	input \P2_reg0_reg[1]/NET0131  ;
	input \P2_reg0_reg[20]/NET0131  ;
	input \P2_reg0_reg[21]/NET0131  ;
	input \P2_reg0_reg[22]/NET0131  ;
	input \P2_reg0_reg[23]/NET0131  ;
	input \P2_reg0_reg[24]/NET0131  ;
	input \P2_reg0_reg[25]/NET0131  ;
	input \P2_reg0_reg[26]/NET0131  ;
	input \P2_reg0_reg[27]/NET0131  ;
	input \P2_reg0_reg[28]/NET0131  ;
	input \P2_reg0_reg[29]/NET0131  ;
	input \P2_reg0_reg[2]/NET0131  ;
	input \P2_reg0_reg[30]/NET0131  ;
	input \P2_reg0_reg[31]/NET0131  ;
	input \P2_reg0_reg[3]/NET0131  ;
	input \P2_reg0_reg[4]/NET0131  ;
	input \P2_reg0_reg[5]/NET0131  ;
	input \P2_reg0_reg[6]/NET0131  ;
	input \P2_reg0_reg[7]/NET0131  ;
	input \P2_reg0_reg[8]/NET0131  ;
	input \P2_reg0_reg[9]/NET0131  ;
	input \P2_reg1_reg[0]/NET0131  ;
	input \P2_reg1_reg[10]/NET0131  ;
	input \P2_reg1_reg[11]/NET0131  ;
	input \P2_reg1_reg[12]/NET0131  ;
	input \P2_reg1_reg[13]/NET0131  ;
	input \P2_reg1_reg[14]/NET0131  ;
	input \P2_reg1_reg[15]/NET0131  ;
	input \P2_reg1_reg[16]/NET0131  ;
	input \P2_reg1_reg[17]/NET0131  ;
	input \P2_reg1_reg[18]/NET0131  ;
	input \P2_reg1_reg[19]/NET0131  ;
	input \P2_reg1_reg[1]/NET0131  ;
	input \P2_reg1_reg[20]/NET0131  ;
	input \P2_reg1_reg[21]/NET0131  ;
	input \P2_reg1_reg[22]/NET0131  ;
	input \P2_reg1_reg[23]/NET0131  ;
	input \P2_reg1_reg[24]/NET0131  ;
	input \P2_reg1_reg[25]/NET0131  ;
	input \P2_reg1_reg[26]/NET0131  ;
	input \P2_reg1_reg[27]/NET0131  ;
	input \P2_reg1_reg[28]/NET0131  ;
	input \P2_reg1_reg[29]/NET0131  ;
	input \P2_reg1_reg[2]/NET0131  ;
	input \P2_reg1_reg[30]/NET0131  ;
	input \P2_reg1_reg[31]/NET0131  ;
	input \P2_reg1_reg[3]/NET0131  ;
	input \P2_reg1_reg[4]/NET0131  ;
	input \P2_reg1_reg[5]/NET0131  ;
	input \P2_reg1_reg[6]/NET0131  ;
	input \P2_reg1_reg[7]/NET0131  ;
	input \P2_reg1_reg[8]/NET0131  ;
	input \P2_reg1_reg[9]/NET0131  ;
	input \P2_reg2_reg[0]/NET0131  ;
	input \P2_reg2_reg[10]/NET0131  ;
	input \P2_reg2_reg[11]/NET0131  ;
	input \P2_reg2_reg[12]/NET0131  ;
	input \P2_reg2_reg[13]/NET0131  ;
	input \P2_reg2_reg[14]/NET0131  ;
	input \P2_reg2_reg[15]/NET0131  ;
	input \P2_reg2_reg[16]/NET0131  ;
	input \P2_reg2_reg[17]/NET0131  ;
	input \P2_reg2_reg[18]/NET0131  ;
	input \P2_reg2_reg[19]/NET0131  ;
	input \P2_reg2_reg[1]/NET0131  ;
	input \P2_reg2_reg[20]/NET0131  ;
	input \P2_reg2_reg[21]/NET0131  ;
	input \P2_reg2_reg[22]/NET0131  ;
	input \P2_reg2_reg[23]/NET0131  ;
	input \P2_reg2_reg[24]/NET0131  ;
	input \P2_reg2_reg[25]/NET0131  ;
	input \P2_reg2_reg[26]/NET0131  ;
	input \P2_reg2_reg[27]/NET0131  ;
	input \P2_reg2_reg[28]/NET0131  ;
	input \P2_reg2_reg[29]/NET0131  ;
	input \P2_reg2_reg[2]/NET0131  ;
	input \P2_reg2_reg[30]/NET0131  ;
	input \P2_reg2_reg[31]/NET0131  ;
	input \P2_reg2_reg[3]/NET0131  ;
	input \P2_reg2_reg[4]/NET0131  ;
	input \P2_reg2_reg[5]/NET0131  ;
	input \P2_reg2_reg[6]/NET0131  ;
	input \P2_reg2_reg[7]/NET0131  ;
	input \P2_reg2_reg[8]/NET0131  ;
	input \P2_reg2_reg[9]/NET0131  ;
	input \P2_reg3_reg[0]/NET0131  ;
	input \P2_reg3_reg[10]/NET0131  ;
	input \P2_reg3_reg[11]/NET0131  ;
	input \P2_reg3_reg[12]/NET0131  ;
	input \P2_reg3_reg[13]/NET0131  ;
	input \P2_reg3_reg[14]/NET0131  ;
	input \P2_reg3_reg[15]/NET0131  ;
	input \P2_reg3_reg[16]/NET0131  ;
	input \P2_reg3_reg[17]/NET0131  ;
	input \P2_reg3_reg[18]/NET0131  ;
	input \P2_reg3_reg[19]/NET0131  ;
	input \P2_reg3_reg[1]/NET0131  ;
	input \P2_reg3_reg[20]/NET0131  ;
	input \P2_reg3_reg[21]/NET0131  ;
	input \P2_reg3_reg[22]/NET0131  ;
	input \P2_reg3_reg[23]/NET0131  ;
	input \P2_reg3_reg[24]/NET0131  ;
	input \P2_reg3_reg[25]/NET0131  ;
	input \P2_reg3_reg[26]/NET0131  ;
	input \P2_reg3_reg[27]/NET0131  ;
	input \P2_reg3_reg[28]/NET0131  ;
	input \P2_reg3_reg[2]/NET0131  ;
	input \P2_reg3_reg[3]/NET0131  ;
	input \P2_reg3_reg[4]/NET0131  ;
	input \P2_reg3_reg[5]/NET0131  ;
	input \P2_reg3_reg[6]/NET0131  ;
	input \P2_reg3_reg[7]/NET0131  ;
	input \P2_reg3_reg[8]/NET0131  ;
	input \P2_reg3_reg[9]/NET0131  ;
	input \P2_wr_reg/NET0131  ;
	input \si[0]_pad  ;
	input \si[10]_pad  ;
	input \si[11]_pad  ;
	input \si[12]_pad  ;
	input \si[13]_pad  ;
	input \si[14]_pad  ;
	input \si[15]_pad  ;
	input \si[16]_pad  ;
	input \si[17]_pad  ;
	input \si[18]_pad  ;
	input \si[19]_pad  ;
	input \si[1]_pad  ;
	input \si[20]_pad  ;
	input \si[21]_pad  ;
	input \si[22]_pad  ;
	input \si[23]_pad  ;
	input \si[24]_pad  ;
	input \si[25]_pad  ;
	input \si[26]_pad  ;
	input \si[27]_pad  ;
	input \si[28]_pad  ;
	input \si[29]_pad  ;
	input \si[2]_pad  ;
	input \si[30]_pad  ;
	input \si[31]_pad  ;
	input \si[3]_pad  ;
	input \si[4]_pad  ;
	input \si[5]_pad  ;
	input \si[6]_pad  ;
	input \si[7]_pad  ;
	input \si[8]_pad  ;
	input \si[9]_pad  ;
	output \P1_state_reg[0]/NET0131_syn_2  ;
	output \_al_n0  ;
	output \_al_n1  ;
	output \g21_dup/_0_  ;
	output \g71037/_0_  ;
	output \g71048/_0_  ;
	output \g71049/_0_  ;
	output \g71050/_0_  ;
	output \g71052/_0_  ;
	output \g71053/_0_  ;
	output \g71054/_0_  ;
	output \g71055/_0_  ;
	output \g71080/_0_  ;
	output \g71081/_0_  ;
	output \g71082/_0_  ;
	output \g71084/_0_  ;
	output \g71085/_0_  ;
	output \g71086/_0_  ;
	output \g71087/_0_  ;
	output \g71088/_0_  ;
	output \g71089/_0_  ;
	output \g71121/_0_  ;
	output \g71122/_0_  ;
	output \g71123/_0_  ;
	output \g71130/_0_  ;
	output \g71131/_0_  ;
	output \g71132/_0_  ;
	output \g71135/_0_  ;
	output \g71136/_0_  ;
	output \g71137/_0_  ;
	output \g71138/_0_  ;
	output \g71139/_0_  ;
	output \g71141/_0_  ;
	output \g71142/_0_  ;
	output \g71143/_0_  ;
	output \g71144/_0_  ;
	output \g71145/_0_  ;
	output \g71146/_0_  ;
	output \g71147/_0_  ;
	output \g71179/_0_  ;
	output \g71186/_0_  ;
	output \g71194/_0_  ;
	output \g71195/_0_  ;
	output \g71196/_0_  ;
	output \g71197/_0_  ;
	output \g71200/_0_  ;
	output \g71201/_0_  ;
	output \g71202/_0_  ;
	output \g71203/_0_  ;
	output \g71204/_0_  ;
	output \g71205/_0_  ;
	output \g71206/_0_  ;
	output \g71207/_0_  ;
	output \g71208/_0_  ;
	output \g71209/_0_  ;
	output \g71210/_0_  ;
	output \g71211/_0_  ;
	output \g71212/_0_  ;
	output \g71213/_0_  ;
	output \g71214/_0_  ;
	output \g71215/_0_  ;
	output \g71262/_0_  ;
	output \g71263/_0_  ;
	output \g71264/_0_  ;
	output \g71291/_0_  ;
	output \g71294/_0_  ;
	output \g71295/_0_  ;
	output \g71296/_0_  ;
	output \g71297/_0_  ;
	output \g71298/_0_  ;
	output \g71299/_0_  ;
	output \g71300/_0_  ;
	output \g71302/_0_  ;
	output \g71303/_0_  ;
	output \g71304/_0_  ;
	output \g71305/_0_  ;
	output \g71306/_0_  ;
	output \g71307/_0_  ;
	output \g71308/_0_  ;
	output \g71354/_0_  ;
	output \g71359/_0_  ;
	output \g71400/_0_  ;
	output \g71401/_0_  ;
	output \g71402/_0_  ;
	output \g71403/_0_  ;
	output \g71404/_0_  ;
	output \g71405/_0_  ;
	output \g71406/_0_  ;
	output \g71407/_0_  ;
	output \g71408/_0_  ;
	output \g71409/_0_  ;
	output \g71410/_0_  ;
	output \g71411/_0_  ;
	output \g71412/_0_  ;
	output \g71413/_0_  ;
	output \g71414/_0_  ;
	output \g71415/_0_  ;
	output \g71416/_0_  ;
	output \g71417/_0_  ;
	output \g71418/_0_  ;
	output \g71420/_0_  ;
	output \g71421/_0_  ;
	output \g71422/_0_  ;
	output \g71423/_0_  ;
	output \g71424/_0_  ;
	output \g71484/_0_  ;
	output \g71485/_0_  ;
	output \g71486/_0_  ;
	output \g71488/_0_  ;
	output \g71489/_0_  ;
	output \g71490/_0_  ;
	output \g71492/_0_  ;
	output \g71493/_0_  ;
	output \g71537/_0_  ;
	output \g71538/_0_  ;
	output \g71539/_0_  ;
	output \g71540/_0_  ;
	output \g71541/_0_  ;
	output \g71542/_0_  ;
	output \g71543/_0_  ;
	output \g71544/_0_  ;
	output \g71545/_0_  ;
	output \g71546/_0_  ;
	output \g71547/_0_  ;
	output \g71548/_0_  ;
	output \g71549/_0_  ;
	output \g71550/_0_  ;
	output \g71551/_0_  ;
	output \g71552/_0_  ;
	output \g71553/_0_  ;
	output \g71554/_0_  ;
	output \g71555/_0_  ;
	output \g71608/_0_  ;
	output \g71609/_0_  ;
	output \g71613/_0_  ;
	output \g71615/_0_  ;
	output \g71617/_0_  ;
	output \g71619/_0_  ;
	output \g71620/_0_  ;
	output \g71621/_0_  ;
	output \g71690/_0_  ;
	output \g71691/_0_  ;
	output \g71692/_0_  ;
	output \g71693/_0_  ;
	output \g71694/_0_  ;
	output \g71696/_0_  ;
	output \g71697/_0_  ;
	output \g71698/_0_  ;
	output \g71699/_0_  ;
	output \g71700/_0_  ;
	output \g71701/_0_  ;
	output \g71702/_0_  ;
	output \g71703/_0_  ;
	output \g71704/_0_  ;
	output \g71705/_0_  ;
	output \g71707/_0_  ;
	output \g71708/_0_  ;
	output \g71709/_0_  ;
	output \g71710/_0_  ;
	output \g71711/_0_  ;
	output \g71712/_0_  ;
	output \g71713/_0_  ;
	output \g71788/_0_  ;
	output \g71789/_0_  ;
	output \g71792/_0_  ;
	output \g71793/_0_  ;
	output \g71794/_0_  ;
	output \g71859/_0_  ;
	output \g71860/_0_  ;
	output \g71861/_0_  ;
	output \g71862/_0_  ;
	output \g71863/_0_  ;
	output \g71864/_0_  ;
	output \g71865/_0_  ;
	output \g71866/_0_  ;
	output \g71867/_0_  ;
	output \g71868/_0_  ;
	output \g71869/_0_  ;
	output \g71870/_0_  ;
	output \g71871/_0_  ;
	output \g71872/_0_  ;
	output \g71873/_0_  ;
	output \g71874/_0_  ;
	output \g71875/_0_  ;
	output \g71876/_0_  ;
	output \g71877/_0_  ;
	output \g71878/_0_  ;
	output \g71879/_0_  ;
	output \g71918/_0_  ;
	output \g71921/_0_  ;
	output \g72042/_0_  ;
	output \g72045/_0_  ;
	output \g72046/_0_  ;
	output \g72047/_0_  ;
	output \g72048/_0_  ;
	output \g72049/_0_  ;
	output \g72050/_0_  ;
	output \g72051/_0_  ;
	output \g72052/_0_  ;
	output \g72053/_0_  ;
	output \g72054/_0_  ;
	output \g72055/_0_  ;
	output \g72056/_0_  ;
	output \g72059/_0_  ;
	output \g72060/_0_  ;
	output \g72061/_0_  ;
	output \g72062/_0_  ;
	output \g72063/_0_  ;
	output \g72064/_0_  ;
	output \g72065/_0_  ;
	output \g72185/_0_  ;
	output \g72302/_0_  ;
	output \g72304/_0_  ;
	output \g72468/_0_  ;
	output \g72577/_0_  ;
	output \g72578/_0_  ;
	output \g72579/_0_  ;
	output \g72580/_0_  ;
	output \g72585/_0_  ;
	output \g72742/_0_  ;
	output \g72758/_0_  ;
	output \g72947/_0_  ;
	output \g72948/_0_  ;
	output \g72952/_0_  ;
	output \g72954/_0_  ;
	output \g72955/_0_  ;
	output \g72956/_0_  ;
	output \g72957/_0_  ;
	output \g73346/_0_  ;
	output \g73349/_0_  ;
	output \g73350/_0_  ;
	output \g73357/_0_  ;
	output \g73618/_0_  ;
	output \g74419/_0_  ;
	output \g74422/_0_  ;
	output \g74426/_0_  ;
	output \g74671/_0_  ;
	output \g75421/_0_  ;
	output \g75424/_0_  ;
	output \g75430/_0_  ;
	output \g76173/_0_  ;
	output \g76175/_0_  ;
	output \g76177/_0_  ;
	output \g76178/_0_  ;
	output \g76179/_0_  ;
	output \g76506/_0_  ;
	output \g80645/_3_  ;
	output \g80646/_3_  ;
	output \g80647/_3_  ;
	output \g80648/_3_  ;
	output \g80649/_0_  ;
	output \g80650/_0_  ;
	output \g80952/_0_  ;
	output \g80956/_0_  ;
	output \g80957/_0_  ;
	output \g80958/_0_  ;
	output \g80959/_0_  ;
	output \g80960/_0_  ;
	output \g80961/_0_  ;
	output \g80962/_0_  ;
	output \g80963/_0_  ;
	output \g80964/_0_  ;
	output \g80965/_0_  ;
	output \g80966/_3_  ;
	output \g80967/_0_  ;
	output \g80968/_0_  ;
	output \g80969/_0_  ;
	output \g80970/_0_  ;
	output \g80971/_0_  ;
	output \g80972/_0_  ;
	output \g80973/_0_  ;
	output \g80974/_3_  ;
	output \g80975/_0_  ;
	output \g80976/_0_  ;
	output \g80977/_0_  ;
	output \g80978/_3_  ;
	output \g80979/_0_  ;
	output \g80980/_0_  ;
	output \g80981/_0_  ;
	output \g80982/_3_  ;
	output \g81025/_3_  ;
	output \g81026/_3_  ;
	output \g81027/_3_  ;
	output \g81028/_3_  ;
	output \g81029/_3_  ;
	output \g81030/_3_  ;
	output \g81031/_3_  ;
	output \g81032/_3_  ;
	output \g81033/_3_  ;
	output \g81034/_3_  ;
	output \g81035/_3_  ;
	output \g81036/_3_  ;
	output \g81037/_3_  ;
	output \g81038/_3_  ;
	output \g81039/_3_  ;
	output \g81040/_3_  ;
	output \g81041/_3_  ;
	output \g81042/_3_  ;
	output \g81043/_0_  ;
	output \g81044/_3_  ;
	output \g81045/_0_  ;
	output \g81046/_3_  ;
	output \g81047/_3_  ;
	output \g81048/_0_  ;
	output \g81049/_3_  ;
	output \g81050/_3_  ;
	output \g81051/_3_  ;
	output \g81052/_3_  ;
	output \g81524/_0_  ;
	output \g81534/_0_  ;
	output \g82411/_0_  ;
	output \g82413/_0_  ;
	output \g82414/_0_  ;
	output \g82415/_0_  ;
	output \g82416/_0_  ;
	output \g82417/_0_  ;
	output \g82418/_0_  ;
	output \g82419/_0_  ;
	output \g82420/_0_  ;
	output \g82421/_0_  ;
	output \g82422/_0_  ;
	output \g82423/_0_  ;
	output \g82424/_0_  ;
	output \g82425/_0_  ;
	output \g82426/_0_  ;
	output \g82427/_0_  ;
	output \g82428/_0_  ;
	output \g82429/_0_  ;
	output \g82430/_0_  ;
	output \g82432/_0_  ;
	output \g82435/_0_  ;
	output \g82436/_0_  ;
	output \g83031/u3_syn_4  ;
	output \g83221/_0_  ;
	output \g83364/_0_  ;
	output \g83474/_0_  ;
	output \g83478/_0_  ;
	output \g83479/_0_  ;
	output \g83480/_0_  ;
	output \g83481/_0_  ;
	output \g83482/_0_  ;
	output \g83484/_0_  ;
	output \g83486/_0_  ;
	output \g83487/_0_  ;
	output \g83488/_0_  ;
	output \g83489/_0_  ;
	output \g83490/_0_  ;
	output \g83491/_0_  ;
	output \g83492/_0_  ;
	output \g83493/_0_  ;
	output \g83494/_0_  ;
	output \g83495/_0_  ;
	output \g83496/_0_  ;
	output \g83505/_0_  ;
	output \g83622/u3_syn_4  ;
	output \g83853/_0_  ;
	output \g83905/_0_  ;
	output \g84145/u3_syn_4  ;
	output \g84148/u3_syn_4  ;
	output \g85427/_2_  ;
	output \g85433/_0_  ;
	output \g85458/_0_  ;
	output \g85512/_0_  ;
	output \g85517/_0_  ;
	output \g85963/_0_  ;
	output \g85996/_0_  ;
	output \g86064/_0_  ;
	output \g86079/_0_  ;
	output \g86088/_0_  ;
	output \g86096/_0_  ;
	output \g86107/_0_  ;
	output \g86159/_0_  ;
	output \g86232_dup/_0_  ;
	output \g86249/_0_  ;
	output \g86258/_0_  ;
	output \g86268/_0_  ;
	output \g86278/_0_  ;
	output \g86281/_0_  ;
	output \g86293/_0_  ;
	output \g86305/_0_  ;
	output \g86313/_0_  ;
	output \g86329/_0_  ;
	output \g86338/_0_  ;
	output \g86355/_0_  ;
	output \g86362/_0_  ;
	output \g86375/_0_  ;
	output \g86385/_0_  ;
	output \g86394/_0_  ;
	output \g86405/_0_  ;
	output \g86413/_0_  ;
	output \g86425/_0_  ;
	output \g86433_dup/_0_  ;
	output \g86441/_0_  ;
	output \g86448/_0_  ;
	output \g86484/_0_  ;
	output \g86493/_0_  ;
	output \g86501/_0_  ;
	output \g86509/_0_  ;
	output \g86518/_0_  ;
	output \g86527/_0_  ;
	output \g86531/_0_  ;
	output \g86541/_0_  ;
	output \g86549/_0_  ;
	output \g86577/_0_  ;
	output \g86598/_0_  ;
	output \g86607/_0_  ;
	output \g87968/_0_  ;
	output \g93740/_0_  ;
	output \g93779/_0_  ;
	output \g93782/_0_  ;
	output \g93859/_0_  ;
	output \g93950/_0_  ;
	output \g93972/_0_  ;
	output \g94026/_0_  ;
	output \g94078/_0_  ;
	output \g94095/_0_  ;
	output \g94136/_0_  ;
	output \g94238/_0_  ;
	output \g94252/_0_  ;
	output \g94278/_0_  ;
	output \g94380/_0_  ;
	output \g94545/_0_  ;
	output \g94586/_0_  ;
	output \g94640/_0_  ;
	output \g94710/_0_  ;
	output \g94743/_0_  ;
	output \g94877/_0_  ;
	output \g95093/_0_  ;
	output \g95139/_0_  ;
	output \g95161/_0_  ;
	output \g95165/_0_  ;
	output \g95204/_0_  ;
	output \g95395/_0_  ;
	output \g95447/_0_  ;
	output rd_pad ;
	output \so[0]_pad  ;
	output \so[10]_pad  ;
	output \so[11]_pad  ;
	output \so[12]_pad  ;
	output \so[13]_pad  ;
	output \so[14]_pad  ;
	output \so[15]_pad  ;
	output \so[16]_pad  ;
	output \so[17]_pad  ;
	output \so[18]_pad  ;
	output \so[19]_pad  ;
	output \so[1]_pad  ;
	output \so[2]_pad  ;
	output \so[3]_pad  ;
	output \so[4]_pad  ;
	output \so[5]_pad  ;
	output \so[6]_pad  ;
	output \so[7]_pad  ;
	output \so[8]_pad  ;
	output \so[9]_pad  ;
	output wr_pad ;
	wire _w7215_ ;
	wire _w7214_ ;
	wire _w7213_ ;
	wire _w7212_ ;
	wire _w7211_ ;
	wire _w7210_ ;
	wire _w7209_ ;
	wire _w7208_ ;
	wire _w7207_ ;
	wire _w7206_ ;
	wire _w7205_ ;
	wire _w7204_ ;
	wire _w7203_ ;
	wire _w7202_ ;
	wire _w7201_ ;
	wire _w7200_ ;
	wire _w7199_ ;
	wire _w7198_ ;
	wire _w7197_ ;
	wire _w7196_ ;
	wire _w7195_ ;
	wire _w7194_ ;
	wire _w7193_ ;
	wire _w7192_ ;
	wire _w7191_ ;
	wire _w7190_ ;
	wire _w7189_ ;
	wire _w7188_ ;
	wire _w7187_ ;
	wire _w7186_ ;
	wire _w7185_ ;
	wire _w7184_ ;
	wire _w7183_ ;
	wire _w7182_ ;
	wire _w7181_ ;
	wire _w7180_ ;
	wire _w7179_ ;
	wire _w7178_ ;
	wire _w7177_ ;
	wire _w7176_ ;
	wire _w7175_ ;
	wire _w7174_ ;
	wire _w7173_ ;
	wire _w7172_ ;
	wire _w7171_ ;
	wire _w7170_ ;
	wire _w7169_ ;
	wire _w7168_ ;
	wire _w7167_ ;
	wire _w7166_ ;
	wire _w7165_ ;
	wire _w7164_ ;
	wire _w7163_ ;
	wire _w7162_ ;
	wire _w7161_ ;
	wire _w7160_ ;
	wire _w7159_ ;
	wire _w7158_ ;
	wire _w7157_ ;
	wire _w7156_ ;
	wire _w7155_ ;
	wire _w7154_ ;
	wire _w7153_ ;
	wire _w7152_ ;
	wire _w7151_ ;
	wire _w7150_ ;
	wire _w7149_ ;
	wire _w7148_ ;
	wire _w7147_ ;
	wire _w7146_ ;
	wire _w7145_ ;
	wire _w7144_ ;
	wire _w7143_ ;
	wire _w7142_ ;
	wire _w7141_ ;
	wire _w7140_ ;
	wire _w7139_ ;
	wire _w7138_ ;
	wire _w7137_ ;
	wire _w7136_ ;
	wire _w7135_ ;
	wire _w7134_ ;
	wire _w7133_ ;
	wire _w7132_ ;
	wire _w7131_ ;
	wire _w7130_ ;
	wire _w7129_ ;
	wire _w7128_ ;
	wire _w7127_ ;
	wire _w7126_ ;
	wire _w7125_ ;
	wire _w7124_ ;
	wire _w7123_ ;
	wire _w7122_ ;
	wire _w7121_ ;
	wire _w7120_ ;
	wire _w7119_ ;
	wire _w7118_ ;
	wire _w7117_ ;
	wire _w7116_ ;
	wire _w7115_ ;
	wire _w7114_ ;
	wire _w7113_ ;
	wire _w7112_ ;
	wire _w7111_ ;
	wire _w7110_ ;
	wire _w7109_ ;
	wire _w7108_ ;
	wire _w7107_ ;
	wire _w7106_ ;
	wire _w7105_ ;
	wire _w7104_ ;
	wire _w7103_ ;
	wire _w7102_ ;
	wire _w7101_ ;
	wire _w7100_ ;
	wire _w7099_ ;
	wire _w7098_ ;
	wire _w7097_ ;
	wire _w7096_ ;
	wire _w7095_ ;
	wire _w7094_ ;
	wire _w7093_ ;
	wire _w7092_ ;
	wire _w7091_ ;
	wire _w7090_ ;
	wire _w7089_ ;
	wire _w7088_ ;
	wire _w7087_ ;
	wire _w7086_ ;
	wire _w7085_ ;
	wire _w7084_ ;
	wire _w7083_ ;
	wire _w7082_ ;
	wire _w7081_ ;
	wire _w7080_ ;
	wire _w7079_ ;
	wire _w7078_ ;
	wire _w7077_ ;
	wire _w7076_ ;
	wire _w7075_ ;
	wire _w7074_ ;
	wire _w7073_ ;
	wire _w7072_ ;
	wire _w7071_ ;
	wire _w7070_ ;
	wire _w7069_ ;
	wire _w7068_ ;
	wire _w7067_ ;
	wire _w7066_ ;
	wire _w7065_ ;
	wire _w7064_ ;
	wire _w7063_ ;
	wire _w7062_ ;
	wire _w7061_ ;
	wire _w7060_ ;
	wire _w7059_ ;
	wire _w7058_ ;
	wire _w7057_ ;
	wire _w7056_ ;
	wire _w7055_ ;
	wire _w7054_ ;
	wire _w7053_ ;
	wire _w7052_ ;
	wire _w7051_ ;
	wire _w7050_ ;
	wire _w7049_ ;
	wire _w7048_ ;
	wire _w7047_ ;
	wire _w7046_ ;
	wire _w7045_ ;
	wire _w7044_ ;
	wire _w7043_ ;
	wire _w7042_ ;
	wire _w7041_ ;
	wire _w7040_ ;
	wire _w7039_ ;
	wire _w7038_ ;
	wire _w7037_ ;
	wire _w7036_ ;
	wire _w7035_ ;
	wire _w7034_ ;
	wire _w7033_ ;
	wire _w7032_ ;
	wire _w7031_ ;
	wire _w7030_ ;
	wire _w7029_ ;
	wire _w7028_ ;
	wire _w7027_ ;
	wire _w7026_ ;
	wire _w7025_ ;
	wire _w7024_ ;
	wire _w7023_ ;
	wire _w7022_ ;
	wire _w7021_ ;
	wire _w7020_ ;
	wire _w7019_ ;
	wire _w7018_ ;
	wire _w7017_ ;
	wire _w7016_ ;
	wire _w7015_ ;
	wire _w7014_ ;
	wire _w7013_ ;
	wire _w7012_ ;
	wire _w7011_ ;
	wire _w7010_ ;
	wire _w7009_ ;
	wire _w7008_ ;
	wire _w7007_ ;
	wire _w7006_ ;
	wire _w7005_ ;
	wire _w7004_ ;
	wire _w7003_ ;
	wire _w7002_ ;
	wire _w7001_ ;
	wire _w7000_ ;
	wire _w6999_ ;
	wire _w6998_ ;
	wire _w6997_ ;
	wire _w6996_ ;
	wire _w6995_ ;
	wire _w6994_ ;
	wire _w6993_ ;
	wire _w6992_ ;
	wire _w6991_ ;
	wire _w6990_ ;
	wire _w6989_ ;
	wire _w6988_ ;
	wire _w6987_ ;
	wire _w6986_ ;
	wire _w6985_ ;
	wire _w6984_ ;
	wire _w6983_ ;
	wire _w6982_ ;
	wire _w6981_ ;
	wire _w6980_ ;
	wire _w6979_ ;
	wire _w6978_ ;
	wire _w6977_ ;
	wire _w6976_ ;
	wire _w6975_ ;
	wire _w6974_ ;
	wire _w6973_ ;
	wire _w6972_ ;
	wire _w6971_ ;
	wire _w6970_ ;
	wire _w6969_ ;
	wire _w6968_ ;
	wire _w6967_ ;
	wire _w6966_ ;
	wire _w6965_ ;
	wire _w6964_ ;
	wire _w6963_ ;
	wire _w6962_ ;
	wire _w6961_ ;
	wire _w6960_ ;
	wire _w6959_ ;
	wire _w6958_ ;
	wire _w6957_ ;
	wire _w6956_ ;
	wire _w6955_ ;
	wire _w6954_ ;
	wire _w6953_ ;
	wire _w6952_ ;
	wire _w6951_ ;
	wire _w6950_ ;
	wire _w6949_ ;
	wire _w6948_ ;
	wire _w6947_ ;
	wire _w6946_ ;
	wire _w6945_ ;
	wire _w6944_ ;
	wire _w6943_ ;
	wire _w6942_ ;
	wire _w6941_ ;
	wire _w6940_ ;
	wire _w6939_ ;
	wire _w6938_ ;
	wire _w6937_ ;
	wire _w6936_ ;
	wire _w6935_ ;
	wire _w6934_ ;
	wire _w6933_ ;
	wire _w6932_ ;
	wire _w6931_ ;
	wire _w6930_ ;
	wire _w6929_ ;
	wire _w6928_ ;
	wire _w6927_ ;
	wire _w6926_ ;
	wire _w6925_ ;
	wire _w6924_ ;
	wire _w6923_ ;
	wire _w6922_ ;
	wire _w6921_ ;
	wire _w6920_ ;
	wire _w6919_ ;
	wire _w6918_ ;
	wire _w6917_ ;
	wire _w6916_ ;
	wire _w6915_ ;
	wire _w6914_ ;
	wire _w6913_ ;
	wire _w6912_ ;
	wire _w6911_ ;
	wire _w6910_ ;
	wire _w6909_ ;
	wire _w6908_ ;
	wire _w6907_ ;
	wire _w6906_ ;
	wire _w6905_ ;
	wire _w6904_ ;
	wire _w6903_ ;
	wire _w6902_ ;
	wire _w6901_ ;
	wire _w6900_ ;
	wire _w6899_ ;
	wire _w6898_ ;
	wire _w6897_ ;
	wire _w6896_ ;
	wire _w6895_ ;
	wire _w6894_ ;
	wire _w6893_ ;
	wire _w6892_ ;
	wire _w6891_ ;
	wire _w6890_ ;
	wire _w6889_ ;
	wire _w6888_ ;
	wire _w6887_ ;
	wire _w6886_ ;
	wire _w6885_ ;
	wire _w6884_ ;
	wire _w6883_ ;
	wire _w6882_ ;
	wire _w6881_ ;
	wire _w6880_ ;
	wire _w6879_ ;
	wire _w6878_ ;
	wire _w6877_ ;
	wire _w6876_ ;
	wire _w6875_ ;
	wire _w6874_ ;
	wire _w6873_ ;
	wire _w6872_ ;
	wire _w6871_ ;
	wire _w6870_ ;
	wire _w6869_ ;
	wire _w6868_ ;
	wire _w6867_ ;
	wire _w6866_ ;
	wire _w6865_ ;
	wire _w6864_ ;
	wire _w6863_ ;
	wire _w6862_ ;
	wire _w6861_ ;
	wire _w6860_ ;
	wire _w6859_ ;
	wire _w6858_ ;
	wire _w6857_ ;
	wire _w6856_ ;
	wire _w6855_ ;
	wire _w6854_ ;
	wire _w6853_ ;
	wire _w6852_ ;
	wire _w6851_ ;
	wire _w6850_ ;
	wire _w6849_ ;
	wire _w6848_ ;
	wire _w6847_ ;
	wire _w6846_ ;
	wire _w6845_ ;
	wire _w6844_ ;
	wire _w6843_ ;
	wire _w6842_ ;
	wire _w6841_ ;
	wire _w6840_ ;
	wire _w6839_ ;
	wire _w6838_ ;
	wire _w6837_ ;
	wire _w6836_ ;
	wire _w6835_ ;
	wire _w6834_ ;
	wire _w6833_ ;
	wire _w6832_ ;
	wire _w6831_ ;
	wire _w6830_ ;
	wire _w6829_ ;
	wire _w6828_ ;
	wire _w6827_ ;
	wire _w6826_ ;
	wire _w6825_ ;
	wire _w6824_ ;
	wire _w6823_ ;
	wire _w6822_ ;
	wire _w6821_ ;
	wire _w6820_ ;
	wire _w6819_ ;
	wire _w6818_ ;
	wire _w6817_ ;
	wire _w6816_ ;
	wire _w6815_ ;
	wire _w6814_ ;
	wire _w6813_ ;
	wire _w6812_ ;
	wire _w6811_ ;
	wire _w6810_ ;
	wire _w6809_ ;
	wire _w6808_ ;
	wire _w6807_ ;
	wire _w6806_ ;
	wire _w6805_ ;
	wire _w6804_ ;
	wire _w6803_ ;
	wire _w6802_ ;
	wire _w6801_ ;
	wire _w6800_ ;
	wire _w6799_ ;
	wire _w6798_ ;
	wire _w6797_ ;
	wire _w6796_ ;
	wire _w6795_ ;
	wire _w6794_ ;
	wire _w6793_ ;
	wire _w6792_ ;
	wire _w6791_ ;
	wire _w6790_ ;
	wire _w6789_ ;
	wire _w6788_ ;
	wire _w6787_ ;
	wire _w6786_ ;
	wire _w6785_ ;
	wire _w6784_ ;
	wire _w6783_ ;
	wire _w6782_ ;
	wire _w6781_ ;
	wire _w6780_ ;
	wire _w6779_ ;
	wire _w6778_ ;
	wire _w6777_ ;
	wire _w6776_ ;
	wire _w6775_ ;
	wire _w6774_ ;
	wire _w6773_ ;
	wire _w6772_ ;
	wire _w6771_ ;
	wire _w6770_ ;
	wire _w6769_ ;
	wire _w6768_ ;
	wire _w6767_ ;
	wire _w6766_ ;
	wire _w6765_ ;
	wire _w6764_ ;
	wire _w6763_ ;
	wire _w6762_ ;
	wire _w6761_ ;
	wire _w6760_ ;
	wire _w6759_ ;
	wire _w6758_ ;
	wire _w6757_ ;
	wire _w6756_ ;
	wire _w6755_ ;
	wire _w6754_ ;
	wire _w6753_ ;
	wire _w6752_ ;
	wire _w6751_ ;
	wire _w6750_ ;
	wire _w6749_ ;
	wire _w6748_ ;
	wire _w6747_ ;
	wire _w6746_ ;
	wire _w6745_ ;
	wire _w6744_ ;
	wire _w6743_ ;
	wire _w6742_ ;
	wire _w6741_ ;
	wire _w6740_ ;
	wire _w6739_ ;
	wire _w6738_ ;
	wire _w6737_ ;
	wire _w6736_ ;
	wire _w6735_ ;
	wire _w6734_ ;
	wire _w6733_ ;
	wire _w6732_ ;
	wire _w6731_ ;
	wire _w6730_ ;
	wire _w6729_ ;
	wire _w6728_ ;
	wire _w6727_ ;
	wire _w6726_ ;
	wire _w6725_ ;
	wire _w6724_ ;
	wire _w6723_ ;
	wire _w6722_ ;
	wire _w6721_ ;
	wire _w6720_ ;
	wire _w6719_ ;
	wire _w6718_ ;
	wire _w6717_ ;
	wire _w6716_ ;
	wire _w6715_ ;
	wire _w6714_ ;
	wire _w6713_ ;
	wire _w6712_ ;
	wire _w6711_ ;
	wire _w6710_ ;
	wire _w6709_ ;
	wire _w6708_ ;
	wire _w6707_ ;
	wire _w6706_ ;
	wire _w6705_ ;
	wire _w6704_ ;
	wire _w6703_ ;
	wire _w6702_ ;
	wire _w6701_ ;
	wire _w6700_ ;
	wire _w6699_ ;
	wire _w6698_ ;
	wire _w6697_ ;
	wire _w6696_ ;
	wire _w6695_ ;
	wire _w6694_ ;
	wire _w6693_ ;
	wire _w6692_ ;
	wire _w6691_ ;
	wire _w6690_ ;
	wire _w6689_ ;
	wire _w6688_ ;
	wire _w6687_ ;
	wire _w6686_ ;
	wire _w6685_ ;
	wire _w6684_ ;
	wire _w6683_ ;
	wire _w6682_ ;
	wire _w6681_ ;
	wire _w6680_ ;
	wire _w6679_ ;
	wire _w6678_ ;
	wire _w6677_ ;
	wire _w6676_ ;
	wire _w6675_ ;
	wire _w6674_ ;
	wire _w6673_ ;
	wire _w6672_ ;
	wire _w6671_ ;
	wire _w6670_ ;
	wire _w6669_ ;
	wire _w6668_ ;
	wire _w6667_ ;
	wire _w6666_ ;
	wire _w6665_ ;
	wire _w6664_ ;
	wire _w6663_ ;
	wire _w6662_ ;
	wire _w6661_ ;
	wire _w6660_ ;
	wire _w6659_ ;
	wire _w6658_ ;
	wire _w6657_ ;
	wire _w6656_ ;
	wire _w6655_ ;
	wire _w6654_ ;
	wire _w6653_ ;
	wire _w6652_ ;
	wire _w6651_ ;
	wire _w6650_ ;
	wire _w6649_ ;
	wire _w6648_ ;
	wire _w6647_ ;
	wire _w6646_ ;
	wire _w6645_ ;
	wire _w6644_ ;
	wire _w6643_ ;
	wire _w6642_ ;
	wire _w6641_ ;
	wire _w6640_ ;
	wire _w6639_ ;
	wire _w6638_ ;
	wire _w6637_ ;
	wire _w6636_ ;
	wire _w6635_ ;
	wire _w6634_ ;
	wire _w6633_ ;
	wire _w6632_ ;
	wire _w6631_ ;
	wire _w6630_ ;
	wire _w6629_ ;
	wire _w6628_ ;
	wire _w6627_ ;
	wire _w6626_ ;
	wire _w6625_ ;
	wire _w6624_ ;
	wire _w6623_ ;
	wire _w6622_ ;
	wire _w6621_ ;
	wire _w6620_ ;
	wire _w6619_ ;
	wire _w6618_ ;
	wire _w6617_ ;
	wire _w6616_ ;
	wire _w6615_ ;
	wire _w6614_ ;
	wire _w6613_ ;
	wire _w6612_ ;
	wire _w6611_ ;
	wire _w6610_ ;
	wire _w6609_ ;
	wire _w6608_ ;
	wire _w6607_ ;
	wire _w6606_ ;
	wire _w6605_ ;
	wire _w6604_ ;
	wire _w6603_ ;
	wire _w6602_ ;
	wire _w6601_ ;
	wire _w6600_ ;
	wire _w6599_ ;
	wire _w6598_ ;
	wire _w6597_ ;
	wire _w6596_ ;
	wire _w6595_ ;
	wire _w6594_ ;
	wire _w6593_ ;
	wire _w6592_ ;
	wire _w6591_ ;
	wire _w6590_ ;
	wire _w6589_ ;
	wire _w6588_ ;
	wire _w6587_ ;
	wire _w6586_ ;
	wire _w6585_ ;
	wire _w6584_ ;
	wire _w6583_ ;
	wire _w6582_ ;
	wire _w6581_ ;
	wire _w6580_ ;
	wire _w6579_ ;
	wire _w6578_ ;
	wire _w6577_ ;
	wire _w6576_ ;
	wire _w6575_ ;
	wire _w6574_ ;
	wire _w6573_ ;
	wire _w6572_ ;
	wire _w6571_ ;
	wire _w6570_ ;
	wire _w6569_ ;
	wire _w6568_ ;
	wire _w6567_ ;
	wire _w6566_ ;
	wire _w6565_ ;
	wire _w6564_ ;
	wire _w6563_ ;
	wire _w6562_ ;
	wire _w6561_ ;
	wire _w6560_ ;
	wire _w6559_ ;
	wire _w6558_ ;
	wire _w6557_ ;
	wire _w6556_ ;
	wire _w6555_ ;
	wire _w6554_ ;
	wire _w6553_ ;
	wire _w6552_ ;
	wire _w6551_ ;
	wire _w6550_ ;
	wire _w6549_ ;
	wire _w6548_ ;
	wire _w6547_ ;
	wire _w6546_ ;
	wire _w6545_ ;
	wire _w6544_ ;
	wire _w6543_ ;
	wire _w6542_ ;
	wire _w6541_ ;
	wire _w6540_ ;
	wire _w6539_ ;
	wire _w6538_ ;
	wire _w6537_ ;
	wire _w6536_ ;
	wire _w6535_ ;
	wire _w6534_ ;
	wire _w6533_ ;
	wire _w6532_ ;
	wire _w6531_ ;
	wire _w6530_ ;
	wire _w6529_ ;
	wire _w6528_ ;
	wire _w6527_ ;
	wire _w6526_ ;
	wire _w6525_ ;
	wire _w6524_ ;
	wire _w6523_ ;
	wire _w6522_ ;
	wire _w6521_ ;
	wire _w6520_ ;
	wire _w6519_ ;
	wire _w6518_ ;
	wire _w6517_ ;
	wire _w6516_ ;
	wire _w6515_ ;
	wire _w6514_ ;
	wire _w6513_ ;
	wire _w6512_ ;
	wire _w6511_ ;
	wire _w6510_ ;
	wire _w6509_ ;
	wire _w6508_ ;
	wire _w6507_ ;
	wire _w6506_ ;
	wire _w6505_ ;
	wire _w6504_ ;
	wire _w6503_ ;
	wire _w6502_ ;
	wire _w6501_ ;
	wire _w6500_ ;
	wire _w6499_ ;
	wire _w6498_ ;
	wire _w6497_ ;
	wire _w6496_ ;
	wire _w6495_ ;
	wire _w6494_ ;
	wire _w6493_ ;
	wire _w6492_ ;
	wire _w6491_ ;
	wire _w6490_ ;
	wire _w6489_ ;
	wire _w6488_ ;
	wire _w6487_ ;
	wire _w6486_ ;
	wire _w6485_ ;
	wire _w6484_ ;
	wire _w6483_ ;
	wire _w6482_ ;
	wire _w6481_ ;
	wire _w6480_ ;
	wire _w6479_ ;
	wire _w6478_ ;
	wire _w6477_ ;
	wire _w6476_ ;
	wire _w6475_ ;
	wire _w6474_ ;
	wire _w6473_ ;
	wire _w6472_ ;
	wire _w6471_ ;
	wire _w6470_ ;
	wire _w6469_ ;
	wire _w6468_ ;
	wire _w6467_ ;
	wire _w6466_ ;
	wire _w6465_ ;
	wire _w6464_ ;
	wire _w6463_ ;
	wire _w6462_ ;
	wire _w6461_ ;
	wire _w6460_ ;
	wire _w6459_ ;
	wire _w6458_ ;
	wire _w6457_ ;
	wire _w6456_ ;
	wire _w6455_ ;
	wire _w6454_ ;
	wire _w6453_ ;
	wire _w6452_ ;
	wire _w6451_ ;
	wire _w6450_ ;
	wire _w6449_ ;
	wire _w6448_ ;
	wire _w6447_ ;
	wire _w6446_ ;
	wire _w6445_ ;
	wire _w6444_ ;
	wire _w6443_ ;
	wire _w6442_ ;
	wire _w6441_ ;
	wire _w6440_ ;
	wire _w6439_ ;
	wire _w6438_ ;
	wire _w6437_ ;
	wire _w6436_ ;
	wire _w6435_ ;
	wire _w6434_ ;
	wire _w6433_ ;
	wire _w6432_ ;
	wire _w6431_ ;
	wire _w6430_ ;
	wire _w6429_ ;
	wire _w6428_ ;
	wire _w6427_ ;
	wire _w6426_ ;
	wire _w6425_ ;
	wire _w6424_ ;
	wire _w6423_ ;
	wire _w6422_ ;
	wire _w6421_ ;
	wire _w6420_ ;
	wire _w6419_ ;
	wire _w6418_ ;
	wire _w6417_ ;
	wire _w6416_ ;
	wire _w6415_ ;
	wire _w6414_ ;
	wire _w6413_ ;
	wire _w6412_ ;
	wire _w6411_ ;
	wire _w6410_ ;
	wire _w6409_ ;
	wire _w6408_ ;
	wire _w6407_ ;
	wire _w6406_ ;
	wire _w6405_ ;
	wire _w6404_ ;
	wire _w6403_ ;
	wire _w6402_ ;
	wire _w6401_ ;
	wire _w6400_ ;
	wire _w6399_ ;
	wire _w6398_ ;
	wire _w6397_ ;
	wire _w6396_ ;
	wire _w6395_ ;
	wire _w6394_ ;
	wire _w6393_ ;
	wire _w6392_ ;
	wire _w6391_ ;
	wire _w6390_ ;
	wire _w6389_ ;
	wire _w6388_ ;
	wire _w6387_ ;
	wire _w6386_ ;
	wire _w6385_ ;
	wire _w6384_ ;
	wire _w6383_ ;
	wire _w6382_ ;
	wire _w6381_ ;
	wire _w6380_ ;
	wire _w6379_ ;
	wire _w6378_ ;
	wire _w6377_ ;
	wire _w6376_ ;
	wire _w6375_ ;
	wire _w6374_ ;
	wire _w6373_ ;
	wire _w6372_ ;
	wire _w6371_ ;
	wire _w6370_ ;
	wire _w6369_ ;
	wire _w6368_ ;
	wire _w6367_ ;
	wire _w6366_ ;
	wire _w6365_ ;
	wire _w6364_ ;
	wire _w6363_ ;
	wire _w6362_ ;
	wire _w6361_ ;
	wire _w6360_ ;
	wire _w6359_ ;
	wire _w6358_ ;
	wire _w6357_ ;
	wire _w6356_ ;
	wire _w6355_ ;
	wire _w6354_ ;
	wire _w6353_ ;
	wire _w6352_ ;
	wire _w6351_ ;
	wire _w6350_ ;
	wire _w6349_ ;
	wire _w6348_ ;
	wire _w6347_ ;
	wire _w6346_ ;
	wire _w6345_ ;
	wire _w6344_ ;
	wire _w6343_ ;
	wire _w6342_ ;
	wire _w6341_ ;
	wire _w6340_ ;
	wire _w6339_ ;
	wire _w6338_ ;
	wire _w6337_ ;
	wire _w6336_ ;
	wire _w6335_ ;
	wire _w6334_ ;
	wire _w6333_ ;
	wire _w6332_ ;
	wire _w6331_ ;
	wire _w6330_ ;
	wire _w6329_ ;
	wire _w6328_ ;
	wire _w6327_ ;
	wire _w6326_ ;
	wire _w6325_ ;
	wire _w6324_ ;
	wire _w6323_ ;
	wire _w6322_ ;
	wire _w6321_ ;
	wire _w6320_ ;
	wire _w6319_ ;
	wire _w6318_ ;
	wire _w6317_ ;
	wire _w6316_ ;
	wire _w6315_ ;
	wire _w6314_ ;
	wire _w6313_ ;
	wire _w6312_ ;
	wire _w6311_ ;
	wire _w6310_ ;
	wire _w6309_ ;
	wire _w6308_ ;
	wire _w6307_ ;
	wire _w6306_ ;
	wire _w6305_ ;
	wire _w6304_ ;
	wire _w6303_ ;
	wire _w6302_ ;
	wire _w6301_ ;
	wire _w6300_ ;
	wire _w6299_ ;
	wire _w6298_ ;
	wire _w6297_ ;
	wire _w6296_ ;
	wire _w6295_ ;
	wire _w6294_ ;
	wire _w6293_ ;
	wire _w6292_ ;
	wire _w6291_ ;
	wire _w6290_ ;
	wire _w6289_ ;
	wire _w6288_ ;
	wire _w6287_ ;
	wire _w6286_ ;
	wire _w6285_ ;
	wire _w6284_ ;
	wire _w6283_ ;
	wire _w6282_ ;
	wire _w6281_ ;
	wire _w6280_ ;
	wire _w6279_ ;
	wire _w6278_ ;
	wire _w6277_ ;
	wire _w6276_ ;
	wire _w6275_ ;
	wire _w6274_ ;
	wire _w6273_ ;
	wire _w6272_ ;
	wire _w6271_ ;
	wire _w6270_ ;
	wire _w6269_ ;
	wire _w6268_ ;
	wire _w6267_ ;
	wire _w6266_ ;
	wire _w6265_ ;
	wire _w6264_ ;
	wire _w6263_ ;
	wire _w6262_ ;
	wire _w6261_ ;
	wire _w6260_ ;
	wire _w6259_ ;
	wire _w6258_ ;
	wire _w6257_ ;
	wire _w6256_ ;
	wire _w6255_ ;
	wire _w6254_ ;
	wire _w6253_ ;
	wire _w6252_ ;
	wire _w6251_ ;
	wire _w6250_ ;
	wire _w6249_ ;
	wire _w6248_ ;
	wire _w6247_ ;
	wire _w6246_ ;
	wire _w6245_ ;
	wire _w6244_ ;
	wire _w6243_ ;
	wire _w6242_ ;
	wire _w6241_ ;
	wire _w6240_ ;
	wire _w6239_ ;
	wire _w6238_ ;
	wire _w6237_ ;
	wire _w6236_ ;
	wire _w6235_ ;
	wire _w6234_ ;
	wire _w6233_ ;
	wire _w6232_ ;
	wire _w6231_ ;
	wire _w6230_ ;
	wire _w6229_ ;
	wire _w6228_ ;
	wire _w6227_ ;
	wire _w6226_ ;
	wire _w6225_ ;
	wire _w6224_ ;
	wire _w6223_ ;
	wire _w6222_ ;
	wire _w6221_ ;
	wire _w6220_ ;
	wire _w6219_ ;
	wire _w6218_ ;
	wire _w6217_ ;
	wire _w6216_ ;
	wire _w6215_ ;
	wire _w6214_ ;
	wire _w6213_ ;
	wire _w6212_ ;
	wire _w6211_ ;
	wire _w6210_ ;
	wire _w6209_ ;
	wire _w6208_ ;
	wire _w6207_ ;
	wire _w6206_ ;
	wire _w6205_ ;
	wire _w6204_ ;
	wire _w6203_ ;
	wire _w6202_ ;
	wire _w6201_ ;
	wire _w6200_ ;
	wire _w6199_ ;
	wire _w6198_ ;
	wire _w6197_ ;
	wire _w6196_ ;
	wire _w6195_ ;
	wire _w6194_ ;
	wire _w6193_ ;
	wire _w6192_ ;
	wire _w6191_ ;
	wire _w6190_ ;
	wire _w6189_ ;
	wire _w6188_ ;
	wire _w6187_ ;
	wire _w6186_ ;
	wire _w6185_ ;
	wire _w6184_ ;
	wire _w6183_ ;
	wire _w6182_ ;
	wire _w6181_ ;
	wire _w6180_ ;
	wire _w6179_ ;
	wire _w6178_ ;
	wire _w6177_ ;
	wire _w6176_ ;
	wire _w6175_ ;
	wire _w6174_ ;
	wire _w6173_ ;
	wire _w6172_ ;
	wire _w6171_ ;
	wire _w6170_ ;
	wire _w6169_ ;
	wire _w6168_ ;
	wire _w6167_ ;
	wire _w6166_ ;
	wire _w6165_ ;
	wire _w6164_ ;
	wire _w6163_ ;
	wire _w6162_ ;
	wire _w6161_ ;
	wire _w6160_ ;
	wire _w6159_ ;
	wire _w6158_ ;
	wire _w6157_ ;
	wire _w6156_ ;
	wire _w6155_ ;
	wire _w6154_ ;
	wire _w6153_ ;
	wire _w6152_ ;
	wire _w6151_ ;
	wire _w6150_ ;
	wire _w6149_ ;
	wire _w6148_ ;
	wire _w6147_ ;
	wire _w6146_ ;
	wire _w6145_ ;
	wire _w6144_ ;
	wire _w6143_ ;
	wire _w6142_ ;
	wire _w6141_ ;
	wire _w6140_ ;
	wire _w6139_ ;
	wire _w6138_ ;
	wire _w6137_ ;
	wire _w6136_ ;
	wire _w6135_ ;
	wire _w6134_ ;
	wire _w6133_ ;
	wire _w6132_ ;
	wire _w6131_ ;
	wire _w6130_ ;
	wire _w6129_ ;
	wire _w6128_ ;
	wire _w6127_ ;
	wire _w6126_ ;
	wire _w6125_ ;
	wire _w6124_ ;
	wire _w6123_ ;
	wire _w6122_ ;
	wire _w6121_ ;
	wire _w6120_ ;
	wire _w6119_ ;
	wire _w6118_ ;
	wire _w6117_ ;
	wire _w6116_ ;
	wire _w6115_ ;
	wire _w6114_ ;
	wire _w6113_ ;
	wire _w6112_ ;
	wire _w6111_ ;
	wire _w6110_ ;
	wire _w6109_ ;
	wire _w6108_ ;
	wire _w6107_ ;
	wire _w6106_ ;
	wire _w6105_ ;
	wire _w6104_ ;
	wire _w6103_ ;
	wire _w6102_ ;
	wire _w6101_ ;
	wire _w6100_ ;
	wire _w6099_ ;
	wire _w6098_ ;
	wire _w6097_ ;
	wire _w6096_ ;
	wire _w6095_ ;
	wire _w6094_ ;
	wire _w6093_ ;
	wire _w6092_ ;
	wire _w6091_ ;
	wire _w6090_ ;
	wire _w6089_ ;
	wire _w6088_ ;
	wire _w6087_ ;
	wire _w6086_ ;
	wire _w6085_ ;
	wire _w6084_ ;
	wire _w6083_ ;
	wire _w6082_ ;
	wire _w6081_ ;
	wire _w6080_ ;
	wire _w6079_ ;
	wire _w6078_ ;
	wire _w6077_ ;
	wire _w6076_ ;
	wire _w6075_ ;
	wire _w6074_ ;
	wire _w6073_ ;
	wire _w6072_ ;
	wire _w6071_ ;
	wire _w6070_ ;
	wire _w6069_ ;
	wire _w6068_ ;
	wire _w6067_ ;
	wire _w6066_ ;
	wire _w6065_ ;
	wire _w6064_ ;
	wire _w6063_ ;
	wire _w6062_ ;
	wire _w6061_ ;
	wire _w6060_ ;
	wire _w6059_ ;
	wire _w6058_ ;
	wire _w6057_ ;
	wire _w6056_ ;
	wire _w6055_ ;
	wire _w6054_ ;
	wire _w6053_ ;
	wire _w6052_ ;
	wire _w6051_ ;
	wire _w6050_ ;
	wire _w6049_ ;
	wire _w6048_ ;
	wire _w6047_ ;
	wire _w6046_ ;
	wire _w6045_ ;
	wire _w6044_ ;
	wire _w6043_ ;
	wire _w6042_ ;
	wire _w6041_ ;
	wire _w6040_ ;
	wire _w6039_ ;
	wire _w6038_ ;
	wire _w6037_ ;
	wire _w6036_ ;
	wire _w6035_ ;
	wire _w6034_ ;
	wire _w6033_ ;
	wire _w6032_ ;
	wire _w6031_ ;
	wire _w6030_ ;
	wire _w6029_ ;
	wire _w6028_ ;
	wire _w6027_ ;
	wire _w6026_ ;
	wire _w6025_ ;
	wire _w6024_ ;
	wire _w6023_ ;
	wire _w6022_ ;
	wire _w6021_ ;
	wire _w6020_ ;
	wire _w6019_ ;
	wire _w6018_ ;
	wire _w6017_ ;
	wire _w6016_ ;
	wire _w6015_ ;
	wire _w6014_ ;
	wire _w6013_ ;
	wire _w6012_ ;
	wire _w6011_ ;
	wire _w6010_ ;
	wire _w6009_ ;
	wire _w6008_ ;
	wire _w6007_ ;
	wire _w6006_ ;
	wire _w6005_ ;
	wire _w6004_ ;
	wire _w6003_ ;
	wire _w6002_ ;
	wire _w6001_ ;
	wire _w6000_ ;
	wire _w5999_ ;
	wire _w5998_ ;
	wire _w5997_ ;
	wire _w5996_ ;
	wire _w5995_ ;
	wire _w5994_ ;
	wire _w5993_ ;
	wire _w5992_ ;
	wire _w5991_ ;
	wire _w5990_ ;
	wire _w5989_ ;
	wire _w5988_ ;
	wire _w5987_ ;
	wire _w5986_ ;
	wire _w5985_ ;
	wire _w5984_ ;
	wire _w5983_ ;
	wire _w5982_ ;
	wire _w5981_ ;
	wire _w5980_ ;
	wire _w5979_ ;
	wire _w5978_ ;
	wire _w5977_ ;
	wire _w5976_ ;
	wire _w5975_ ;
	wire _w5974_ ;
	wire _w5973_ ;
	wire _w5972_ ;
	wire _w5971_ ;
	wire _w5970_ ;
	wire _w5969_ ;
	wire _w5968_ ;
	wire _w5967_ ;
	wire _w5966_ ;
	wire _w5965_ ;
	wire _w5964_ ;
	wire _w5963_ ;
	wire _w5962_ ;
	wire _w5961_ ;
	wire _w5960_ ;
	wire _w5959_ ;
	wire _w5958_ ;
	wire _w5957_ ;
	wire _w5956_ ;
	wire _w5955_ ;
	wire _w5954_ ;
	wire _w5953_ ;
	wire _w5952_ ;
	wire _w5951_ ;
	wire _w5950_ ;
	wire _w5949_ ;
	wire _w5948_ ;
	wire _w5947_ ;
	wire _w5946_ ;
	wire _w5945_ ;
	wire _w5944_ ;
	wire _w5943_ ;
	wire _w5942_ ;
	wire _w5941_ ;
	wire _w5940_ ;
	wire _w5939_ ;
	wire _w5938_ ;
	wire _w5937_ ;
	wire _w5936_ ;
	wire _w5935_ ;
	wire _w5934_ ;
	wire _w5933_ ;
	wire _w5932_ ;
	wire _w5931_ ;
	wire _w5930_ ;
	wire _w5929_ ;
	wire _w5928_ ;
	wire _w5927_ ;
	wire _w5926_ ;
	wire _w5925_ ;
	wire _w5924_ ;
	wire _w5923_ ;
	wire _w5922_ ;
	wire _w5921_ ;
	wire _w5920_ ;
	wire _w5919_ ;
	wire _w5918_ ;
	wire _w5917_ ;
	wire _w5916_ ;
	wire _w5915_ ;
	wire _w5914_ ;
	wire _w5913_ ;
	wire _w5912_ ;
	wire _w5911_ ;
	wire _w5910_ ;
	wire _w5909_ ;
	wire _w5908_ ;
	wire _w5907_ ;
	wire _w5906_ ;
	wire _w5905_ ;
	wire _w5904_ ;
	wire _w5903_ ;
	wire _w5902_ ;
	wire _w5901_ ;
	wire _w5900_ ;
	wire _w5899_ ;
	wire _w5898_ ;
	wire _w5897_ ;
	wire _w5896_ ;
	wire _w5895_ ;
	wire _w5894_ ;
	wire _w5893_ ;
	wire _w5892_ ;
	wire _w5891_ ;
	wire _w5890_ ;
	wire _w5889_ ;
	wire _w5888_ ;
	wire _w5887_ ;
	wire _w5886_ ;
	wire _w5885_ ;
	wire _w5884_ ;
	wire _w5883_ ;
	wire _w5882_ ;
	wire _w5881_ ;
	wire _w5880_ ;
	wire _w5879_ ;
	wire _w5878_ ;
	wire _w5877_ ;
	wire _w5876_ ;
	wire _w5875_ ;
	wire _w5874_ ;
	wire _w5873_ ;
	wire _w5872_ ;
	wire _w5871_ ;
	wire _w5870_ ;
	wire _w5869_ ;
	wire _w5868_ ;
	wire _w5867_ ;
	wire _w5866_ ;
	wire _w5865_ ;
	wire _w5864_ ;
	wire _w5863_ ;
	wire _w5862_ ;
	wire _w5861_ ;
	wire _w5860_ ;
	wire _w5859_ ;
	wire _w5858_ ;
	wire _w5857_ ;
	wire _w5856_ ;
	wire _w5855_ ;
	wire _w5854_ ;
	wire _w5853_ ;
	wire _w5852_ ;
	wire _w5851_ ;
	wire _w5850_ ;
	wire _w5849_ ;
	wire _w5848_ ;
	wire _w5847_ ;
	wire _w5846_ ;
	wire _w5845_ ;
	wire _w5844_ ;
	wire _w5843_ ;
	wire _w5842_ ;
	wire _w5841_ ;
	wire _w5840_ ;
	wire _w5839_ ;
	wire _w5838_ ;
	wire _w5837_ ;
	wire _w5836_ ;
	wire _w5835_ ;
	wire _w5834_ ;
	wire _w5833_ ;
	wire _w5832_ ;
	wire _w5831_ ;
	wire _w5830_ ;
	wire _w5829_ ;
	wire _w5828_ ;
	wire _w5827_ ;
	wire _w5826_ ;
	wire _w5825_ ;
	wire _w5824_ ;
	wire _w5823_ ;
	wire _w5822_ ;
	wire _w5821_ ;
	wire _w5820_ ;
	wire _w5819_ ;
	wire _w5818_ ;
	wire _w5817_ ;
	wire _w5816_ ;
	wire _w5815_ ;
	wire _w5814_ ;
	wire _w5813_ ;
	wire _w5812_ ;
	wire _w5811_ ;
	wire _w5810_ ;
	wire _w5809_ ;
	wire _w5808_ ;
	wire _w5807_ ;
	wire _w5806_ ;
	wire _w5805_ ;
	wire _w5804_ ;
	wire _w5803_ ;
	wire _w5802_ ;
	wire _w5801_ ;
	wire _w5800_ ;
	wire _w5799_ ;
	wire _w5798_ ;
	wire _w5797_ ;
	wire _w5796_ ;
	wire _w5795_ ;
	wire _w5794_ ;
	wire _w5793_ ;
	wire _w5792_ ;
	wire _w5791_ ;
	wire _w5790_ ;
	wire _w5789_ ;
	wire _w5788_ ;
	wire _w5787_ ;
	wire _w5786_ ;
	wire _w5785_ ;
	wire _w5784_ ;
	wire _w5783_ ;
	wire _w5782_ ;
	wire _w5781_ ;
	wire _w5780_ ;
	wire _w5779_ ;
	wire _w5778_ ;
	wire _w5777_ ;
	wire _w5776_ ;
	wire _w5775_ ;
	wire _w5774_ ;
	wire _w5773_ ;
	wire _w5772_ ;
	wire _w5771_ ;
	wire _w5770_ ;
	wire _w5769_ ;
	wire _w5768_ ;
	wire _w5767_ ;
	wire _w5766_ ;
	wire _w5765_ ;
	wire _w5764_ ;
	wire _w5763_ ;
	wire _w5762_ ;
	wire _w5761_ ;
	wire _w5760_ ;
	wire _w5759_ ;
	wire _w5758_ ;
	wire _w5757_ ;
	wire _w5756_ ;
	wire _w5755_ ;
	wire _w5754_ ;
	wire _w5753_ ;
	wire _w5752_ ;
	wire _w5751_ ;
	wire _w5750_ ;
	wire _w5749_ ;
	wire _w5748_ ;
	wire _w5747_ ;
	wire _w5746_ ;
	wire _w5745_ ;
	wire _w5744_ ;
	wire _w5743_ ;
	wire _w5742_ ;
	wire _w5741_ ;
	wire _w5740_ ;
	wire _w5739_ ;
	wire _w5738_ ;
	wire _w5737_ ;
	wire _w5736_ ;
	wire _w5735_ ;
	wire _w5734_ ;
	wire _w5733_ ;
	wire _w5732_ ;
	wire _w5731_ ;
	wire _w5730_ ;
	wire _w5729_ ;
	wire _w5728_ ;
	wire _w5727_ ;
	wire _w5726_ ;
	wire _w5725_ ;
	wire _w5724_ ;
	wire _w5723_ ;
	wire _w5722_ ;
	wire _w5721_ ;
	wire _w5720_ ;
	wire _w5719_ ;
	wire _w5718_ ;
	wire _w5717_ ;
	wire _w5716_ ;
	wire _w5715_ ;
	wire _w5714_ ;
	wire _w5713_ ;
	wire _w5712_ ;
	wire _w5711_ ;
	wire _w5710_ ;
	wire _w5709_ ;
	wire _w5708_ ;
	wire _w5707_ ;
	wire _w5706_ ;
	wire _w5705_ ;
	wire _w5704_ ;
	wire _w5703_ ;
	wire _w5702_ ;
	wire _w5701_ ;
	wire _w5700_ ;
	wire _w5699_ ;
	wire _w5698_ ;
	wire _w5697_ ;
	wire _w5696_ ;
	wire _w5695_ ;
	wire _w5694_ ;
	wire _w5693_ ;
	wire _w5692_ ;
	wire _w5691_ ;
	wire _w5690_ ;
	wire _w5689_ ;
	wire _w5688_ ;
	wire _w5687_ ;
	wire _w5686_ ;
	wire _w5685_ ;
	wire _w5684_ ;
	wire _w5683_ ;
	wire _w5682_ ;
	wire _w5681_ ;
	wire _w5680_ ;
	wire _w5679_ ;
	wire _w5678_ ;
	wire _w5677_ ;
	wire _w5676_ ;
	wire _w5675_ ;
	wire _w5674_ ;
	wire _w5673_ ;
	wire _w5672_ ;
	wire _w5671_ ;
	wire _w5670_ ;
	wire _w5669_ ;
	wire _w5668_ ;
	wire _w5667_ ;
	wire _w5666_ ;
	wire _w5665_ ;
	wire _w5664_ ;
	wire _w5663_ ;
	wire _w5662_ ;
	wire _w5661_ ;
	wire _w5660_ ;
	wire _w5659_ ;
	wire _w5658_ ;
	wire _w5657_ ;
	wire _w5656_ ;
	wire _w5655_ ;
	wire _w5654_ ;
	wire _w5653_ ;
	wire _w5652_ ;
	wire _w5651_ ;
	wire _w5650_ ;
	wire _w5649_ ;
	wire _w5648_ ;
	wire _w5647_ ;
	wire _w5646_ ;
	wire _w5645_ ;
	wire _w5644_ ;
	wire _w5643_ ;
	wire _w5642_ ;
	wire _w5641_ ;
	wire _w5640_ ;
	wire _w5639_ ;
	wire _w5638_ ;
	wire _w5637_ ;
	wire _w5636_ ;
	wire _w5635_ ;
	wire _w5634_ ;
	wire _w5633_ ;
	wire _w5632_ ;
	wire _w5631_ ;
	wire _w5630_ ;
	wire _w5629_ ;
	wire _w5628_ ;
	wire _w5627_ ;
	wire _w5626_ ;
	wire _w5625_ ;
	wire _w5624_ ;
	wire _w5623_ ;
	wire _w5622_ ;
	wire _w5621_ ;
	wire _w5620_ ;
	wire _w5619_ ;
	wire _w5618_ ;
	wire _w5617_ ;
	wire _w5616_ ;
	wire _w5615_ ;
	wire _w5614_ ;
	wire _w5613_ ;
	wire _w5612_ ;
	wire _w5611_ ;
	wire _w5610_ ;
	wire _w5609_ ;
	wire _w5608_ ;
	wire _w5607_ ;
	wire _w5606_ ;
	wire _w5605_ ;
	wire _w5604_ ;
	wire _w5603_ ;
	wire _w5602_ ;
	wire _w5601_ ;
	wire _w5600_ ;
	wire _w5599_ ;
	wire _w5598_ ;
	wire _w5597_ ;
	wire _w5596_ ;
	wire _w5595_ ;
	wire _w5594_ ;
	wire _w5593_ ;
	wire _w5592_ ;
	wire _w5591_ ;
	wire _w5590_ ;
	wire _w5589_ ;
	wire _w5588_ ;
	wire _w5587_ ;
	wire _w5586_ ;
	wire _w5585_ ;
	wire _w5584_ ;
	wire _w5583_ ;
	wire _w5582_ ;
	wire _w5581_ ;
	wire _w5580_ ;
	wire _w5579_ ;
	wire _w5578_ ;
	wire _w5577_ ;
	wire _w5576_ ;
	wire _w5575_ ;
	wire _w5574_ ;
	wire _w5573_ ;
	wire _w5572_ ;
	wire _w5571_ ;
	wire _w5570_ ;
	wire _w5569_ ;
	wire _w5568_ ;
	wire _w5567_ ;
	wire _w5566_ ;
	wire _w5565_ ;
	wire _w5564_ ;
	wire _w5563_ ;
	wire _w5562_ ;
	wire _w5561_ ;
	wire _w5560_ ;
	wire _w5559_ ;
	wire _w5558_ ;
	wire _w5557_ ;
	wire _w5556_ ;
	wire _w5555_ ;
	wire _w5554_ ;
	wire _w5553_ ;
	wire _w5552_ ;
	wire _w5551_ ;
	wire _w5550_ ;
	wire _w2819_ ;
	wire _w2818_ ;
	wire _w2817_ ;
	wire _w2816_ ;
	wire _w2815_ ;
	wire _w2814_ ;
	wire _w2813_ ;
	wire _w2812_ ;
	wire _w2811_ ;
	wire _w2810_ ;
	wire _w2809_ ;
	wire _w2808_ ;
	wire _w2807_ ;
	wire _w2806_ ;
	wire _w2805_ ;
	wire _w2804_ ;
	wire _w2803_ ;
	wire _w2802_ ;
	wire _w2801_ ;
	wire _w2800_ ;
	wire _w2799_ ;
	wire _w2798_ ;
	wire _w2797_ ;
	wire _w2796_ ;
	wire _w2795_ ;
	wire _w2794_ ;
	wire _w2793_ ;
	wire _w2792_ ;
	wire _w2791_ ;
	wire _w2790_ ;
	wire _w2789_ ;
	wire _w2788_ ;
	wire _w2787_ ;
	wire _w2786_ ;
	wire _w2785_ ;
	wire _w2784_ ;
	wire _w2783_ ;
	wire _w2782_ ;
	wire _w2781_ ;
	wire _w2780_ ;
	wire _w2779_ ;
	wire _w2778_ ;
	wire _w2777_ ;
	wire _w2776_ ;
	wire _w2775_ ;
	wire _w2774_ ;
	wire _w2773_ ;
	wire _w2772_ ;
	wire _w2771_ ;
	wire _w2770_ ;
	wire _w2769_ ;
	wire _w2768_ ;
	wire _w2767_ ;
	wire _w2766_ ;
	wire _w2765_ ;
	wire _w2764_ ;
	wire _w2763_ ;
	wire _w2762_ ;
	wire _w2761_ ;
	wire _w2760_ ;
	wire _w2759_ ;
	wire _w2758_ ;
	wire _w2757_ ;
	wire _w2756_ ;
	wire _w2755_ ;
	wire _w2754_ ;
	wire _w2753_ ;
	wire _w2752_ ;
	wire _w2751_ ;
	wire _w2750_ ;
	wire _w2749_ ;
	wire _w2748_ ;
	wire _w2747_ ;
	wire _w2746_ ;
	wire _w2745_ ;
	wire _w2744_ ;
	wire _w2743_ ;
	wire _w2742_ ;
	wire _w2741_ ;
	wire _w2740_ ;
	wire _w2739_ ;
	wire _w2738_ ;
	wire _w2737_ ;
	wire _w2736_ ;
	wire _w2735_ ;
	wire _w2734_ ;
	wire _w2733_ ;
	wire _w2732_ ;
	wire _w2731_ ;
	wire _w2730_ ;
	wire _w2729_ ;
	wire _w2728_ ;
	wire _w2727_ ;
	wire _w2726_ ;
	wire _w2725_ ;
	wire _w2724_ ;
	wire _w2723_ ;
	wire _w2722_ ;
	wire _w2721_ ;
	wire _w2720_ ;
	wire _w2719_ ;
	wire _w2718_ ;
	wire _w2717_ ;
	wire _w2716_ ;
	wire _w2715_ ;
	wire _w2714_ ;
	wire _w2713_ ;
	wire _w2712_ ;
	wire _w2711_ ;
	wire _w2710_ ;
	wire _w2709_ ;
	wire _w2708_ ;
	wire _w2707_ ;
	wire _w2706_ ;
	wire _w2705_ ;
	wire _w2704_ ;
	wire _w2703_ ;
	wire _w2702_ ;
	wire _w2701_ ;
	wire _w2700_ ;
	wire _w2699_ ;
	wire _w2698_ ;
	wire _w2697_ ;
	wire _w2696_ ;
	wire _w2695_ ;
	wire _w2694_ ;
	wire _w2693_ ;
	wire _w2692_ ;
	wire _w2691_ ;
	wire _w2690_ ;
	wire _w2689_ ;
	wire _w2688_ ;
	wire _w2687_ ;
	wire _w2686_ ;
	wire _w2685_ ;
	wire _w2684_ ;
	wire _w2683_ ;
	wire _w2682_ ;
	wire _w2681_ ;
	wire _w2680_ ;
	wire _w2679_ ;
	wire _w2678_ ;
	wire _w2677_ ;
	wire _w2676_ ;
	wire _w2675_ ;
	wire _w2674_ ;
	wire _w2673_ ;
	wire _w2672_ ;
	wire _w2671_ ;
	wire _w2670_ ;
	wire _w2669_ ;
	wire _w2668_ ;
	wire _w2667_ ;
	wire _w2666_ ;
	wire _w2665_ ;
	wire _w2664_ ;
	wire _w2663_ ;
	wire _w2662_ ;
	wire _w2661_ ;
	wire _w2660_ ;
	wire _w2659_ ;
	wire _w2658_ ;
	wire _w2657_ ;
	wire _w2656_ ;
	wire _w2655_ ;
	wire _w2654_ ;
	wire _w2653_ ;
	wire _w2652_ ;
	wire _w2651_ ;
	wire _w2650_ ;
	wire _w2649_ ;
	wire _w2648_ ;
	wire _w2647_ ;
	wire _w2646_ ;
	wire _w2645_ ;
	wire _w2644_ ;
	wire _w2643_ ;
	wire _w2642_ ;
	wire _w2641_ ;
	wire _w2640_ ;
	wire _w2639_ ;
	wire _w2638_ ;
	wire _w2637_ ;
	wire _w2636_ ;
	wire _w2635_ ;
	wire _w2634_ ;
	wire _w2633_ ;
	wire _w2632_ ;
	wire _w2631_ ;
	wire _w2630_ ;
	wire _w2629_ ;
	wire _w2628_ ;
	wire _w2627_ ;
	wire _w2626_ ;
	wire _w2625_ ;
	wire _w2624_ ;
	wire _w2623_ ;
	wire _w2622_ ;
	wire _w2621_ ;
	wire _w2620_ ;
	wire _w2619_ ;
	wire _w2618_ ;
	wire _w2617_ ;
	wire _w2616_ ;
	wire _w2615_ ;
	wire _w2614_ ;
	wire _w2613_ ;
	wire _w2612_ ;
	wire _w2611_ ;
	wire _w2610_ ;
	wire _w2609_ ;
	wire _w2608_ ;
	wire _w2607_ ;
	wire _w2606_ ;
	wire _w2605_ ;
	wire _w2604_ ;
	wire _w2603_ ;
	wire _w2602_ ;
	wire _w2601_ ;
	wire _w2600_ ;
	wire _w2599_ ;
	wire _w2598_ ;
	wire _w2597_ ;
	wire _w2596_ ;
	wire _w2595_ ;
	wire _w2594_ ;
	wire _w2593_ ;
	wire _w2592_ ;
	wire _w2591_ ;
	wire _w2590_ ;
	wire _w2589_ ;
	wire _w2588_ ;
	wire _w2587_ ;
	wire _w2586_ ;
	wire _w2585_ ;
	wire _w2584_ ;
	wire _w2583_ ;
	wire _w2582_ ;
	wire _w2581_ ;
	wire _w2580_ ;
	wire _w2579_ ;
	wire _w2578_ ;
	wire _w2577_ ;
	wire _w2576_ ;
	wire _w2575_ ;
	wire _w2574_ ;
	wire _w2572_ ;
	wire _w2571_ ;
	wire _w2570_ ;
	wire _w2569_ ;
	wire _w2568_ ;
	wire _w2567_ ;
	wire _w2566_ ;
	wire _w2565_ ;
	wire _w2564_ ;
	wire _w2563_ ;
	wire _w2562_ ;
	wire _w2561_ ;
	wire _w2560_ ;
	wire _w2559_ ;
	wire _w2558_ ;
	wire _w2557_ ;
	wire _w2556_ ;
	wire _w2555_ ;
	wire _w2554_ ;
	wire _w2553_ ;
	wire _w2552_ ;
	wire _w2551_ ;
	wire _w2550_ ;
	wire _w2549_ ;
	wire _w2548_ ;
	wire _w2547_ ;
	wire _w2546_ ;
	wire _w2545_ ;
	wire _w2544_ ;
	wire _w2543_ ;
	wire _w2542_ ;
	wire _w2541_ ;
	wire _w2540_ ;
	wire _w2539_ ;
	wire _w2538_ ;
	wire _w2537_ ;
	wire _w2536_ ;
	wire _w2535_ ;
	wire _w2534_ ;
	wire _w2533_ ;
	wire _w2532_ ;
	wire _w2531_ ;
	wire _w2530_ ;
	wire _w2529_ ;
	wire _w2528_ ;
	wire _w2527_ ;
	wire _w2526_ ;
	wire _w2525_ ;
	wire _w2524_ ;
	wire _w2523_ ;
	wire _w2522_ ;
	wire _w2521_ ;
	wire _w2520_ ;
	wire _w2519_ ;
	wire _w2518_ ;
	wire _w2517_ ;
	wire _w2516_ ;
	wire _w2515_ ;
	wire _w2514_ ;
	wire _w2513_ ;
	wire _w2512_ ;
	wire _w2511_ ;
	wire _w2510_ ;
	wire _w2509_ ;
	wire _w2508_ ;
	wire _w2507_ ;
	wire _w2506_ ;
	wire _w2505_ ;
	wire _w2504_ ;
	wire _w2503_ ;
	wire _w2502_ ;
	wire _w2501_ ;
	wire _w2500_ ;
	wire _w2499_ ;
	wire _w2498_ ;
	wire _w2497_ ;
	wire _w2496_ ;
	wire _w2495_ ;
	wire _w2494_ ;
	wire _w2493_ ;
	wire _w2492_ ;
	wire _w2491_ ;
	wire _w2490_ ;
	wire _w2489_ ;
	wire _w2488_ ;
	wire _w2487_ ;
	wire _w2486_ ;
	wire _w2485_ ;
	wire _w2484_ ;
	wire _w2483_ ;
	wire _w2482_ ;
	wire _w2481_ ;
	wire _w2480_ ;
	wire _w2479_ ;
	wire _w2478_ ;
	wire _w2477_ ;
	wire _w2476_ ;
	wire _w2475_ ;
	wire _w2474_ ;
	wire _w2473_ ;
	wire _w2472_ ;
	wire _w2471_ ;
	wire _w2470_ ;
	wire _w2469_ ;
	wire _w2468_ ;
	wire _w2467_ ;
	wire _w2466_ ;
	wire _w2465_ ;
	wire _w2464_ ;
	wire _w2463_ ;
	wire _w2462_ ;
	wire _w2461_ ;
	wire _w2460_ ;
	wire _w2459_ ;
	wire _w2458_ ;
	wire _w2457_ ;
	wire _w2456_ ;
	wire _w2455_ ;
	wire _w2454_ ;
	wire _w2453_ ;
	wire _w2452_ ;
	wire _w2451_ ;
	wire _w2450_ ;
	wire _w2449_ ;
	wire _w2448_ ;
	wire _w2447_ ;
	wire _w2446_ ;
	wire _w2445_ ;
	wire _w2444_ ;
	wire _w2443_ ;
	wire _w2442_ ;
	wire _w2441_ ;
	wire _w2440_ ;
	wire _w2439_ ;
	wire _w2438_ ;
	wire _w2437_ ;
	wire _w2436_ ;
	wire _w2435_ ;
	wire _w2434_ ;
	wire _w2433_ ;
	wire _w2432_ ;
	wire _w2431_ ;
	wire _w2430_ ;
	wire _w2429_ ;
	wire _w2428_ ;
	wire _w2427_ ;
	wire _w2426_ ;
	wire _w2425_ ;
	wire _w2424_ ;
	wire _w2423_ ;
	wire _w2422_ ;
	wire _w2421_ ;
	wire _w2420_ ;
	wire _w2419_ ;
	wire _w2418_ ;
	wire _w2417_ ;
	wire _w2416_ ;
	wire _w2415_ ;
	wire _w2414_ ;
	wire _w2413_ ;
	wire _w2412_ ;
	wire _w2411_ ;
	wire _w2410_ ;
	wire _w2409_ ;
	wire _w2408_ ;
	wire _w2407_ ;
	wire _w2406_ ;
	wire _w2405_ ;
	wire _w2404_ ;
	wire _w2403_ ;
	wire _w2402_ ;
	wire _w2401_ ;
	wire _w2400_ ;
	wire _w2399_ ;
	wire _w2398_ ;
	wire _w2397_ ;
	wire _w2396_ ;
	wire _w2395_ ;
	wire _w2394_ ;
	wire _w2393_ ;
	wire _w2392_ ;
	wire _w2391_ ;
	wire _w2390_ ;
	wire _w2389_ ;
	wire _w2388_ ;
	wire _w2387_ ;
	wire _w2386_ ;
	wire _w2385_ ;
	wire _w2384_ ;
	wire _w2383_ ;
	wire _w2382_ ;
	wire _w2381_ ;
	wire _w2380_ ;
	wire _w2379_ ;
	wire _w2378_ ;
	wire _w2377_ ;
	wire _w2376_ ;
	wire _w2375_ ;
	wire _w2374_ ;
	wire _w2373_ ;
	wire _w2372_ ;
	wire _w2371_ ;
	wire _w2370_ ;
	wire _w2369_ ;
	wire _w2368_ ;
	wire _w2367_ ;
	wire _w2366_ ;
	wire _w2365_ ;
	wire _w2364_ ;
	wire _w2363_ ;
	wire _w2362_ ;
	wire _w2361_ ;
	wire _w2360_ ;
	wire _w2359_ ;
	wire _w2358_ ;
	wire _w2357_ ;
	wire _w2356_ ;
	wire _w2355_ ;
	wire _w2354_ ;
	wire _w2353_ ;
	wire _w2352_ ;
	wire _w2351_ ;
	wire _w2350_ ;
	wire _w2349_ ;
	wire _w2348_ ;
	wire _w2347_ ;
	wire _w2346_ ;
	wire _w2345_ ;
	wire _w2344_ ;
	wire _w2343_ ;
	wire _w2342_ ;
	wire _w2341_ ;
	wire _w2340_ ;
	wire _w2339_ ;
	wire _w2338_ ;
	wire _w2337_ ;
	wire _w2336_ ;
	wire _w2335_ ;
	wire _w2334_ ;
	wire _w2333_ ;
	wire _w2332_ ;
	wire _w2331_ ;
	wire _w2330_ ;
	wire _w2329_ ;
	wire _w2328_ ;
	wire _w2327_ ;
	wire _w2326_ ;
	wire _w2325_ ;
	wire _w2324_ ;
	wire _w2323_ ;
	wire _w2322_ ;
	wire _w2321_ ;
	wire _w2320_ ;
	wire _w2319_ ;
	wire _w2318_ ;
	wire _w2317_ ;
	wire _w2316_ ;
	wire _w2315_ ;
	wire _w2314_ ;
	wire _w2313_ ;
	wire _w2312_ ;
	wire _w2311_ ;
	wire _w2310_ ;
	wire _w2309_ ;
	wire _w2308_ ;
	wire _w2307_ ;
	wire _w2306_ ;
	wire _w2305_ ;
	wire _w2304_ ;
	wire _w2303_ ;
	wire _w2302_ ;
	wire _w2301_ ;
	wire _w2300_ ;
	wire _w2299_ ;
	wire _w2298_ ;
	wire _w2297_ ;
	wire _w2296_ ;
	wire _w2295_ ;
	wire _w2294_ ;
	wire _w2293_ ;
	wire _w2292_ ;
	wire _w2291_ ;
	wire _w2290_ ;
	wire _w2289_ ;
	wire _w2288_ ;
	wire _w2287_ ;
	wire _w2286_ ;
	wire _w2285_ ;
	wire _w2284_ ;
	wire _w2283_ ;
	wire _w2282_ ;
	wire _w2281_ ;
	wire _w2280_ ;
	wire _w2279_ ;
	wire _w2278_ ;
	wire _w2277_ ;
	wire _w2276_ ;
	wire _w2275_ ;
	wire _w2274_ ;
	wire _w2273_ ;
	wire _w2272_ ;
	wire _w2271_ ;
	wire _w2270_ ;
	wire _w2269_ ;
	wire _w2268_ ;
	wire _w2267_ ;
	wire _w2266_ ;
	wire _w2265_ ;
	wire _w2264_ ;
	wire _w2263_ ;
	wire _w2262_ ;
	wire _w2261_ ;
	wire _w2260_ ;
	wire _w2259_ ;
	wire _w2258_ ;
	wire _w2257_ ;
	wire _w2256_ ;
	wire _w2255_ ;
	wire _w2254_ ;
	wire _w2253_ ;
	wire _w2252_ ;
	wire _w2251_ ;
	wire _w2250_ ;
	wire _w2249_ ;
	wire _w2248_ ;
	wire _w2247_ ;
	wire _w2246_ ;
	wire _w2245_ ;
	wire _w2244_ ;
	wire _w2243_ ;
	wire _w2242_ ;
	wire _w2241_ ;
	wire _w2240_ ;
	wire _w2239_ ;
	wire _w2238_ ;
	wire _w2237_ ;
	wire _w2236_ ;
	wire _w2235_ ;
	wire _w2234_ ;
	wire _w2233_ ;
	wire _w2232_ ;
	wire _w2231_ ;
	wire _w2230_ ;
	wire _w2229_ ;
	wire _w2228_ ;
	wire _w2227_ ;
	wire _w2226_ ;
	wire _w2225_ ;
	wire _w2224_ ;
	wire _w2223_ ;
	wire _w2222_ ;
	wire _w2221_ ;
	wire _w2220_ ;
	wire _w2219_ ;
	wire _w2218_ ;
	wire _w2217_ ;
	wire _w2216_ ;
	wire _w2215_ ;
	wire _w2214_ ;
	wire _w2213_ ;
	wire _w2212_ ;
	wire _w2211_ ;
	wire _w2210_ ;
	wire _w2209_ ;
	wire _w2208_ ;
	wire _w2207_ ;
	wire _w2206_ ;
	wire _w2205_ ;
	wire _w2204_ ;
	wire _w2203_ ;
	wire _w2202_ ;
	wire _w2201_ ;
	wire _w2200_ ;
	wire _w2199_ ;
	wire _w2198_ ;
	wire _w2197_ ;
	wire _w2196_ ;
	wire _w2195_ ;
	wire _w2194_ ;
	wire _w2193_ ;
	wire _w2192_ ;
	wire _w2191_ ;
	wire _w2190_ ;
	wire _w2189_ ;
	wire _w2188_ ;
	wire _w2187_ ;
	wire _w2186_ ;
	wire _w2185_ ;
	wire _w2184_ ;
	wire _w2183_ ;
	wire _w2182_ ;
	wire _w2181_ ;
	wire _w2180_ ;
	wire _w2179_ ;
	wire _w2178_ ;
	wire _w2177_ ;
	wire _w2176_ ;
	wire _w2175_ ;
	wire _w2174_ ;
	wire _w2173_ ;
	wire _w2172_ ;
	wire _w2171_ ;
	wire _w2170_ ;
	wire _w2169_ ;
	wire _w2168_ ;
	wire _w2167_ ;
	wire _w2166_ ;
	wire _w2165_ ;
	wire _w2164_ ;
	wire _w2163_ ;
	wire _w2162_ ;
	wire _w2161_ ;
	wire _w2160_ ;
	wire _w2159_ ;
	wire _w2158_ ;
	wire _w2157_ ;
	wire _w2156_ ;
	wire _w2155_ ;
	wire _w2154_ ;
	wire _w2153_ ;
	wire _w2152_ ;
	wire _w2151_ ;
	wire _w2150_ ;
	wire _w2149_ ;
	wire _w2148_ ;
	wire _w2147_ ;
	wire _w2146_ ;
	wire _w2145_ ;
	wire _w2144_ ;
	wire _w2143_ ;
	wire _w2142_ ;
	wire _w2141_ ;
	wire _w2140_ ;
	wire _w2139_ ;
	wire _w2138_ ;
	wire _w2137_ ;
	wire _w2136_ ;
	wire _w2135_ ;
	wire _w2134_ ;
	wire _w2133_ ;
	wire _w2132_ ;
	wire _w2131_ ;
	wire _w2130_ ;
	wire _w2129_ ;
	wire _w2128_ ;
	wire _w2127_ ;
	wire _w2126_ ;
	wire _w2125_ ;
	wire _w2124_ ;
	wire _w2123_ ;
	wire _w2122_ ;
	wire _w2121_ ;
	wire _w2120_ ;
	wire _w2119_ ;
	wire _w2118_ ;
	wire _w2117_ ;
	wire _w2116_ ;
	wire _w2115_ ;
	wire _w2114_ ;
	wire _w2113_ ;
	wire _w2112_ ;
	wire _w2111_ ;
	wire _w2110_ ;
	wire _w2109_ ;
	wire _w2108_ ;
	wire _w2107_ ;
	wire _w2106_ ;
	wire _w2105_ ;
	wire _w2104_ ;
	wire _w2103_ ;
	wire _w2102_ ;
	wire _w2101_ ;
	wire _w2100_ ;
	wire _w2099_ ;
	wire _w2098_ ;
	wire _w2097_ ;
	wire _w2096_ ;
	wire _w2095_ ;
	wire _w2094_ ;
	wire _w2093_ ;
	wire _w2092_ ;
	wire _w2091_ ;
	wire _w2090_ ;
	wire _w2089_ ;
	wire _w2088_ ;
	wire _w2087_ ;
	wire _w2086_ ;
	wire _w2085_ ;
	wire _w2084_ ;
	wire _w2083_ ;
	wire _w2082_ ;
	wire _w2081_ ;
	wire _w2080_ ;
	wire _w2079_ ;
	wire _w2078_ ;
	wire _w2077_ ;
	wire _w2076_ ;
	wire _w2075_ ;
	wire _w2074_ ;
	wire _w2073_ ;
	wire _w2072_ ;
	wire _w2071_ ;
	wire _w2070_ ;
	wire _w2069_ ;
	wire _w2068_ ;
	wire _w2067_ ;
	wire _w2066_ ;
	wire _w2065_ ;
	wire _w2064_ ;
	wire _w2063_ ;
	wire _w2062_ ;
	wire _w2061_ ;
	wire _w2060_ ;
	wire _w2059_ ;
	wire _w2058_ ;
	wire _w2057_ ;
	wire _w2056_ ;
	wire _w2055_ ;
	wire _w2054_ ;
	wire _w2053_ ;
	wire _w2052_ ;
	wire _w2051_ ;
	wire _w2050_ ;
	wire _w2049_ ;
	wire _w2048_ ;
	wire _w2047_ ;
	wire _w2046_ ;
	wire _w2045_ ;
	wire _w2044_ ;
	wire _w2043_ ;
	wire _w2042_ ;
	wire _w2041_ ;
	wire _w2040_ ;
	wire _w2039_ ;
	wire _w2038_ ;
	wire _w2037_ ;
	wire _w2036_ ;
	wire _w2035_ ;
	wire _w2034_ ;
	wire _w2033_ ;
	wire _w2032_ ;
	wire _w2031_ ;
	wire _w2030_ ;
	wire _w2029_ ;
	wire _w2028_ ;
	wire _w2027_ ;
	wire _w2026_ ;
	wire _w2025_ ;
	wire _w2024_ ;
	wire _w2023_ ;
	wire _w2022_ ;
	wire _w2021_ ;
	wire _w2020_ ;
	wire _w2019_ ;
	wire _w2018_ ;
	wire _w2017_ ;
	wire _w2016_ ;
	wire _w2015_ ;
	wire _w2014_ ;
	wire _w2013_ ;
	wire _w2012_ ;
	wire _w2011_ ;
	wire _w2010_ ;
	wire _w2009_ ;
	wire _w2008_ ;
	wire _w2007_ ;
	wire _w2006_ ;
	wire _w2005_ ;
	wire _w2004_ ;
	wire _w2003_ ;
	wire _w2002_ ;
	wire _w2001_ ;
	wire _w2000_ ;
	wire _w1999_ ;
	wire _w1998_ ;
	wire _w1997_ ;
	wire _w1996_ ;
	wire _w1995_ ;
	wire _w1994_ ;
	wire _w1993_ ;
	wire _w1992_ ;
	wire _w1991_ ;
	wire _w1990_ ;
	wire _w1989_ ;
	wire _w1988_ ;
	wire _w1987_ ;
	wire _w1986_ ;
	wire _w1985_ ;
	wire _w1984_ ;
	wire _w1983_ ;
	wire _w1982_ ;
	wire _w1981_ ;
	wire _w1980_ ;
	wire _w1979_ ;
	wire _w1978_ ;
	wire _w1977_ ;
	wire _w1976_ ;
	wire _w1975_ ;
	wire _w1974_ ;
	wire _w1973_ ;
	wire _w1972_ ;
	wire _w1971_ ;
	wire _w1970_ ;
	wire _w1969_ ;
	wire _w1968_ ;
	wire _w1967_ ;
	wire _w1966_ ;
	wire _w1965_ ;
	wire _w1964_ ;
	wire _w1963_ ;
	wire _w1962_ ;
	wire _w1961_ ;
	wire _w1960_ ;
	wire _w1959_ ;
	wire _w1958_ ;
	wire _w1957_ ;
	wire _w1956_ ;
	wire _w1955_ ;
	wire _w1954_ ;
	wire _w1953_ ;
	wire _w1952_ ;
	wire _w1951_ ;
	wire _w1950_ ;
	wire _w1949_ ;
	wire _w1948_ ;
	wire _w1947_ ;
	wire _w1946_ ;
	wire _w1945_ ;
	wire _w1944_ ;
	wire _w1943_ ;
	wire _w1942_ ;
	wire _w1941_ ;
	wire _w1940_ ;
	wire _w1939_ ;
	wire _w1938_ ;
	wire _w1937_ ;
	wire _w1936_ ;
	wire _w1935_ ;
	wire _w1934_ ;
	wire _w1933_ ;
	wire _w1932_ ;
	wire _w1931_ ;
	wire _w1930_ ;
	wire _w1929_ ;
	wire _w1928_ ;
	wire _w1927_ ;
	wire _w1926_ ;
	wire _w1925_ ;
	wire _w1924_ ;
	wire _w1923_ ;
	wire _w1922_ ;
	wire _w1921_ ;
	wire _w1920_ ;
	wire _w1919_ ;
	wire _w1918_ ;
	wire _w1917_ ;
	wire _w1916_ ;
	wire _w1915_ ;
	wire _w1914_ ;
	wire _w1913_ ;
	wire _w1912_ ;
	wire _w1911_ ;
	wire _w1910_ ;
	wire _w1909_ ;
	wire _w1908_ ;
	wire _w1907_ ;
	wire _w1906_ ;
	wire _w1905_ ;
	wire _w1904_ ;
	wire _w1903_ ;
	wire _w1902_ ;
	wire _w1901_ ;
	wire _w1900_ ;
	wire _w1899_ ;
	wire _w1898_ ;
	wire _w1897_ ;
	wire _w1896_ ;
	wire _w1895_ ;
	wire _w1894_ ;
	wire _w1893_ ;
	wire _w1892_ ;
	wire _w1891_ ;
	wire _w1890_ ;
	wire _w1889_ ;
	wire _w1888_ ;
	wire _w1887_ ;
	wire _w1886_ ;
	wire _w1885_ ;
	wire _w1884_ ;
	wire _w1883_ ;
	wire _w1882_ ;
	wire _w1881_ ;
	wire _w1880_ ;
	wire _w1879_ ;
	wire _w1878_ ;
	wire _w1877_ ;
	wire _w1876_ ;
	wire _w1875_ ;
	wire _w1874_ ;
	wire _w1873_ ;
	wire _w1872_ ;
	wire _w1871_ ;
	wire _w1870_ ;
	wire _w1869_ ;
	wire _w1868_ ;
	wire _w1867_ ;
	wire _w1866_ ;
	wire _w1865_ ;
	wire _w1864_ ;
	wire _w1863_ ;
	wire _w1862_ ;
	wire _w1861_ ;
	wire _w1860_ ;
	wire _w1859_ ;
	wire _w1858_ ;
	wire _w1857_ ;
	wire _w1856_ ;
	wire _w1855_ ;
	wire _w1854_ ;
	wire _w1853_ ;
	wire _w1852_ ;
	wire _w1851_ ;
	wire _w1850_ ;
	wire _w1849_ ;
	wire _w1848_ ;
	wire _w1847_ ;
	wire _w1846_ ;
	wire _w1845_ ;
	wire _w1844_ ;
	wire _w1843_ ;
	wire _w1842_ ;
	wire _w1841_ ;
	wire _w1840_ ;
	wire _w1839_ ;
	wire _w1838_ ;
	wire _w1837_ ;
	wire _w1836_ ;
	wire _w1835_ ;
	wire _w1834_ ;
	wire _w1833_ ;
	wire _w1832_ ;
	wire _w1831_ ;
	wire _w1830_ ;
	wire _w1829_ ;
	wire _w1828_ ;
	wire _w1827_ ;
	wire _w1826_ ;
	wire _w1825_ ;
	wire _w1824_ ;
	wire _w1823_ ;
	wire _w1822_ ;
	wire _w1821_ ;
	wire _w1820_ ;
	wire _w1819_ ;
	wire _w1818_ ;
	wire _w1817_ ;
	wire _w1816_ ;
	wire _w1815_ ;
	wire _w1814_ ;
	wire _w1813_ ;
	wire _w1812_ ;
	wire _w1811_ ;
	wire _w1810_ ;
	wire _w1809_ ;
	wire _w1808_ ;
	wire _w1807_ ;
	wire _w1806_ ;
	wire _w1805_ ;
	wire _w1804_ ;
	wire _w1803_ ;
	wire _w1802_ ;
	wire _w1801_ ;
	wire _w1800_ ;
	wire _w1799_ ;
	wire _w1798_ ;
	wire _w1797_ ;
	wire _w1796_ ;
	wire _w1795_ ;
	wire _w1794_ ;
	wire _w1793_ ;
	wire _w1792_ ;
	wire _w1791_ ;
	wire _w1790_ ;
	wire _w1789_ ;
	wire _w1788_ ;
	wire _w1787_ ;
	wire _w1786_ ;
	wire _w1785_ ;
	wire _w1784_ ;
	wire _w1783_ ;
	wire _w1782_ ;
	wire _w1781_ ;
	wire _w1780_ ;
	wire _w1779_ ;
	wire _w1778_ ;
	wire _w1777_ ;
	wire _w1776_ ;
	wire _w1775_ ;
	wire _w1774_ ;
	wire _w1773_ ;
	wire _w1772_ ;
	wire _w1771_ ;
	wire _w1770_ ;
	wire _w1769_ ;
	wire _w1768_ ;
	wire _w1767_ ;
	wire _w1766_ ;
	wire _w1765_ ;
	wire _w1764_ ;
	wire _w1763_ ;
	wire _w1762_ ;
	wire _w1761_ ;
	wire _w1760_ ;
	wire _w1759_ ;
	wire _w1758_ ;
	wire _w1757_ ;
	wire _w1756_ ;
	wire _w1755_ ;
	wire _w1754_ ;
	wire _w1753_ ;
	wire _w1752_ ;
	wire _w1751_ ;
	wire _w1750_ ;
	wire _w1749_ ;
	wire _w1748_ ;
	wire _w1747_ ;
	wire _w1746_ ;
	wire _w1745_ ;
	wire _w1744_ ;
	wire _w1743_ ;
	wire _w1742_ ;
	wire _w1741_ ;
	wire _w1740_ ;
	wire _w1739_ ;
	wire _w1738_ ;
	wire _w1737_ ;
	wire _w1736_ ;
	wire _w1735_ ;
	wire _w1734_ ;
	wire _w1733_ ;
	wire _w1732_ ;
	wire _w1731_ ;
	wire _w1730_ ;
	wire _w1729_ ;
	wire _w1728_ ;
	wire _w1727_ ;
	wire _w1726_ ;
	wire _w1725_ ;
	wire _w1724_ ;
	wire _w1723_ ;
	wire _w1722_ ;
	wire _w1721_ ;
	wire _w1720_ ;
	wire _w1719_ ;
	wire _w1718_ ;
	wire _w1717_ ;
	wire _w1716_ ;
	wire _w1715_ ;
	wire _w1714_ ;
	wire _w1713_ ;
	wire _w1712_ ;
	wire _w1711_ ;
	wire _w1710_ ;
	wire _w1709_ ;
	wire _w1708_ ;
	wire _w1707_ ;
	wire _w1706_ ;
	wire _w1705_ ;
	wire _w1704_ ;
	wire _w1703_ ;
	wire _w1702_ ;
	wire _w1701_ ;
	wire _w1700_ ;
	wire _w1699_ ;
	wire _w1698_ ;
	wire _w1697_ ;
	wire _w1696_ ;
	wire _w1695_ ;
	wire _w1694_ ;
	wire _w1693_ ;
	wire _w1692_ ;
	wire _w1691_ ;
	wire _w1690_ ;
	wire _w1689_ ;
	wire _w1688_ ;
	wire _w1687_ ;
	wire _w1686_ ;
	wire _w1685_ ;
	wire _w1684_ ;
	wire _w1683_ ;
	wire _w1682_ ;
	wire _w1681_ ;
	wire _w1680_ ;
	wire _w1679_ ;
	wire _w1678_ ;
	wire _w1677_ ;
	wire _w1676_ ;
	wire _w1675_ ;
	wire _w1674_ ;
	wire _w1673_ ;
	wire _w1672_ ;
	wire _w1671_ ;
	wire _w1670_ ;
	wire _w1669_ ;
	wire _w1668_ ;
	wire _w1667_ ;
	wire _w1666_ ;
	wire _w1665_ ;
	wire _w1664_ ;
	wire _w1663_ ;
	wire _w1662_ ;
	wire _w1661_ ;
	wire _w1660_ ;
	wire _w1659_ ;
	wire _w1658_ ;
	wire _w1657_ ;
	wire _w1656_ ;
	wire _w1655_ ;
	wire _w1654_ ;
	wire _w1653_ ;
	wire _w1652_ ;
	wire _w1651_ ;
	wire _w1650_ ;
	wire _w1649_ ;
	wire _w1648_ ;
	wire _w1647_ ;
	wire _w1646_ ;
	wire _w1645_ ;
	wire _w1644_ ;
	wire _w1643_ ;
	wire _w1642_ ;
	wire _w1641_ ;
	wire _w1640_ ;
	wire _w1639_ ;
	wire _w1638_ ;
	wire _w1637_ ;
	wire _w1636_ ;
	wire _w1635_ ;
	wire _w1634_ ;
	wire _w1633_ ;
	wire _w1632_ ;
	wire _w1631_ ;
	wire _w1630_ ;
	wire _w1629_ ;
	wire _w1628_ ;
	wire _w1627_ ;
	wire _w1626_ ;
	wire _w1625_ ;
	wire _w1624_ ;
	wire _w1623_ ;
	wire _w1622_ ;
	wire _w1621_ ;
	wire _w1620_ ;
	wire _w1619_ ;
	wire _w1618_ ;
	wire _w1617_ ;
	wire _w1616_ ;
	wire _w1615_ ;
	wire _w1614_ ;
	wire _w1613_ ;
	wire _w1612_ ;
	wire _w1611_ ;
	wire _w1610_ ;
	wire _w1609_ ;
	wire _w1608_ ;
	wire _w1607_ ;
	wire _w1606_ ;
	wire _w1605_ ;
	wire _w1604_ ;
	wire _w1603_ ;
	wire _w1602_ ;
	wire _w1601_ ;
	wire _w1600_ ;
	wire _w1599_ ;
	wire _w1598_ ;
	wire _w1597_ ;
	wire _w1596_ ;
	wire _w1595_ ;
	wire _w1594_ ;
	wire _w1593_ ;
	wire _w1592_ ;
	wire _w1591_ ;
	wire _w1590_ ;
	wire _w1589_ ;
	wire _w1588_ ;
	wire _w1587_ ;
	wire _w1586_ ;
	wire _w1585_ ;
	wire _w1584_ ;
	wire _w1583_ ;
	wire _w1582_ ;
	wire _w1581_ ;
	wire _w1580_ ;
	wire _w1579_ ;
	wire _w1578_ ;
	wire _w1577_ ;
	wire _w1576_ ;
	wire _w1575_ ;
	wire _w1574_ ;
	wire _w1573_ ;
	wire _w1572_ ;
	wire _w1003_ ;
	wire _w1002_ ;
	wire _w1001_ ;
	wire _w1000_ ;
	wire _w999_ ;
	wire _w998_ ;
	wire _w997_ ;
	wire _w996_ ;
	wire _w995_ ;
	wire _w994_ ;
	wire _w993_ ;
	wire _w992_ ;
	wire _w991_ ;
	wire _w990_ ;
	wire _w989_ ;
	wire _w988_ ;
	wire _w987_ ;
	wire _w986_ ;
	wire _w985_ ;
	wire _w984_ ;
	wire _w983_ ;
	wire _w982_ ;
	wire _w981_ ;
	wire _w980_ ;
	wire _w979_ ;
	wire _w978_ ;
	wire _w977_ ;
	wire _w976_ ;
	wire _w975_ ;
	wire _w974_ ;
	wire _w973_ ;
	wire _w972_ ;
	wire _w971_ ;
	wire _w970_ ;
	wire _w969_ ;
	wire _w968_ ;
	wire _w967_ ;
	wire _w966_ ;
	wire _w965_ ;
	wire _w964_ ;
	wire _w963_ ;
	wire _w962_ ;
	wire _w961_ ;
	wire _w960_ ;
	wire _w959_ ;
	wire _w958_ ;
	wire _w957_ ;
	wire _w956_ ;
	wire _w955_ ;
	wire _w954_ ;
	wire _w953_ ;
	wire _w952_ ;
	wire _w951_ ;
	wire _w950_ ;
	wire _w949_ ;
	wire _w948_ ;
	wire _w947_ ;
	wire _w946_ ;
	wire _w945_ ;
	wire _w944_ ;
	wire _w943_ ;
	wire _w942_ ;
	wire _w941_ ;
	wire _w940_ ;
	wire _w939_ ;
	wire _w938_ ;
	wire _w937_ ;
	wire _w936_ ;
	wire _w935_ ;
	wire _w934_ ;
	wire _w933_ ;
	wire _w932_ ;
	wire _w931_ ;
	wire _w930_ ;
	wire _w929_ ;
	wire _w928_ ;
	wire _w927_ ;
	wire _w926_ ;
	wire _w925_ ;
	wire _w924_ ;
	wire _w923_ ;
	wire _w922_ ;
	wire _w921_ ;
	wire _w920_ ;
	wire _w919_ ;
	wire _w918_ ;
	wire _w917_ ;
	wire _w916_ ;
	wire _w915_ ;
	wire _w914_ ;
	wire _w913_ ;
	wire _w912_ ;
	wire _w911_ ;
	wire _w910_ ;
	wire _w909_ ;
	wire _w908_ ;
	wire _w907_ ;
	wire _w906_ ;
	wire _w905_ ;
	wire _w904_ ;
	wire _w903_ ;
	wire _w902_ ;
	wire _w901_ ;
	wire _w900_ ;
	wire _w899_ ;
	wire _w898_ ;
	wire _w897_ ;
	wire _w896_ ;
	wire _w895_ ;
	wire _w894_ ;
	wire _w893_ ;
	wire _w892_ ;
	wire _w891_ ;
	wire _w890_ ;
	wire _w889_ ;
	wire _w888_ ;
	wire _w887_ ;
	wire _w886_ ;
	wire _w885_ ;
	wire _w884_ ;
	wire _w883_ ;
	wire _w882_ ;
	wire _w881_ ;
	wire _w880_ ;
	wire _w879_ ;
	wire _w878_ ;
	wire _w877_ ;
	wire _w876_ ;
	wire _w875_ ;
	wire _w874_ ;
	wire _w873_ ;
	wire _w872_ ;
	wire _w871_ ;
	wire _w870_ ;
	wire _w869_ ;
	wire _w868_ ;
	wire _w867_ ;
	wire _w866_ ;
	wire _w865_ ;
	wire _w864_ ;
	wire _w863_ ;
	wire _w862_ ;
	wire _w861_ ;
	wire _w860_ ;
	wire _w859_ ;
	wire _w858_ ;
	wire _w857_ ;
	wire _w856_ ;
	wire _w855_ ;
	wire _w854_ ;
	wire _w853_ ;
	wire _w852_ ;
	wire _w851_ ;
	wire _w850_ ;
	wire _w849_ ;
	wire _w848_ ;
	wire _w847_ ;
	wire _w846_ ;
	wire _w845_ ;
	wire _w844_ ;
	wire _w843_ ;
	wire _w842_ ;
	wire _w841_ ;
	wire _w840_ ;
	wire _w839_ ;
	wire _w838_ ;
	wire _w837_ ;
	wire _w836_ ;
	wire _w835_ ;
	wire _w834_ ;
	wire _w833_ ;
	wire _w832_ ;
	wire _w831_ ;
	wire _w830_ ;
	wire _w829_ ;
	wire _w828_ ;
	wire _w827_ ;
	wire _w826_ ;
	wire _w825_ ;
	wire _w824_ ;
	wire _w823_ ;
	wire _w822_ ;
	wire _w821_ ;
	wire _w820_ ;
	wire _w819_ ;
	wire _w818_ ;
	wire _w817_ ;
	wire _w816_ ;
	wire _w815_ ;
	wire _w814_ ;
	wire _w813_ ;
	wire _w812_ ;
	wire _w811_ ;
	wire _w810_ ;
	wire _w809_ ;
	wire _w808_ ;
	wire _w807_ ;
	wire _w806_ ;
	wire _w805_ ;
	wire _w804_ ;
	wire _w803_ ;
	wire _w802_ ;
	wire _w801_ ;
	wire _w800_ ;
	wire _w799_ ;
	wire _w798_ ;
	wire _w797_ ;
	wire _w796_ ;
	wire _w795_ ;
	wire _w794_ ;
	wire _w793_ ;
	wire _w792_ ;
	wire _w791_ ;
	wire _w790_ ;
	wire _w789_ ;
	wire _w788_ ;
	wire _w787_ ;
	wire _w786_ ;
	wire _w785_ ;
	wire _w784_ ;
	wire _w783_ ;
	wire _w782_ ;
	wire _w781_ ;
	wire _w780_ ;
	wire _w779_ ;
	wire _w778_ ;
	wire _w777_ ;
	wire _w776_ ;
	wire _w775_ ;
	wire _w774_ ;
	wire _w773_ ;
	wire _w772_ ;
	wire _w771_ ;
	wire _w770_ ;
	wire _w769_ ;
	wire _w768_ ;
	wire _w767_ ;
	wire _w766_ ;
	wire _w765_ ;
	wire _w764_ ;
	wire _w763_ ;
	wire _w762_ ;
	wire _w761_ ;
	wire _w760_ ;
	wire _w759_ ;
	wire _w758_ ;
	wire _w756_ ;
	wire _w755_ ;
	wire _w754_ ;
	wire _w753_ ;
	wire _w752_ ;
	wire _w751_ ;
	wire _w750_ ;
	wire _w749_ ;
	wire _w748_ ;
	wire _w747_ ;
	wire _w746_ ;
	wire _w745_ ;
	wire _w744_ ;
	wire _w743_ ;
	wire _w742_ ;
	wire _w741_ ;
	wire _w740_ ;
	wire _w739_ ;
	wire _w738_ ;
	wire _w737_ ;
	wire _w736_ ;
	wire _w735_ ;
	wire _w734_ ;
	wire _w733_ ;
	wire _w732_ ;
	wire _w731_ ;
	wire _w730_ ;
	wire _w729_ ;
	wire _w728_ ;
	wire _w727_ ;
	wire _w726_ ;
	wire _w725_ ;
	wire _w724_ ;
	wire _w723_ ;
	wire _w722_ ;
	wire _w721_ ;
	wire _w720_ ;
	wire _w589_ ;
	wire _w588_ ;
	wire _w587_ ;
	wire _w586_ ;
	wire _w585_ ;
	wire _w584_ ;
	wire _w583_ ;
	wire _w582_ ;
	wire _w581_ ;
	wire _w580_ ;
	wire _w579_ ;
	wire _w578_ ;
	wire _w577_ ;
	wire _w576_ ;
	wire _w575_ ;
	wire _w574_ ;
	wire _w573_ ;
	wire _w572_ ;
	wire _w571_ ;
	wire _w570_ ;
	wire _w569_ ;
	wire _w568_ ;
	wire _w567_ ;
	wire _w566_ ;
	wire _w565_ ;
	wire _w564_ ;
	wire _w563_ ;
	wire _w562_ ;
	wire _w561_ ;
	wire _w560_ ;
	wire _w559_ ;
	wire _w558_ ;
	wire _w557_ ;
	wire _w556_ ;
	wire _w555_ ;
	wire _w554_ ;
	wire _w553_ ;
	wire _w552_ ;
	wire _w551_ ;
	wire _w550_ ;
	wire _w549_ ;
	wire _w548_ ;
	wire _w547_ ;
	wire _w546_ ;
	wire _w545_ ;
	wire _w544_ ;
	wire _w543_ ;
	wire _w542_ ;
	wire _w541_ ;
	wire _w540_ ;
	wire _w539_ ;
	wire _w538_ ;
	wire _w537_ ;
	wire _w536_ ;
	wire _w535_ ;
	wire _w534_ ;
	wire _w533_ ;
	wire _w532_ ;
	wire _w531_ ;
	wire _w530_ ;
	wire _w529_ ;
	wire _w528_ ;
	wire _w527_ ;
	wire _w526_ ;
	wire _w525_ ;
	wire _w524_ ;
	wire _w523_ ;
	wire _w522_ ;
	wire _w491_ ;
	wire _w490_ ;
	wire _w489_ ;
	wire _w488_ ;
	wire _w487_ ;
	wire _w486_ ;
	wire _w485_ ;
	wire _w484_ ;
	wire _w483_ ;
	wire _w482_ ;
	wire _w481_ ;
	wire _w480_ ;
	wire _w479_ ;
	wire _w478_ ;
	wire _w476_ ;
	wire _w477_ ;
	wire _w511_ ;
	wire _w464_ ;
	wire _w465_ ;
	wire _w466_ ;
	wire _w467_ ;
	wire _w468_ ;
	wire _w469_ ;
	wire _w757_ ;
	wire _w2573_ ;
	wire _w216_ ;
	wire _w5303_ ;
	wire _w1325_ ;
	wire _w473_ ;
	wire _w470_ ;
	wire _w471_ ;
	wire _w472_ ;
	wire _w474_ ;
	wire _w475_ ;
	wire _w492_ ;
	wire _w493_ ;
	wire _w494_ ;
	wire _w495_ ;
	wire _w496_ ;
	wire _w497_ ;
	wire _w498_ ;
	wire _w499_ ;
	wire _w500_ ;
	wire _w501_ ;
	wire _w502_ ;
	wire _w503_ ;
	wire _w504_ ;
	wire _w505_ ;
	wire _w506_ ;
	wire _w507_ ;
	wire _w508_ ;
	wire _w509_ ;
	wire _w510_ ;
	wire _w512_ ;
	wire _w513_ ;
	wire _w514_ ;
	wire _w515_ ;
	wire _w516_ ;
	wire _w517_ ;
	wire _w518_ ;
	wire _w519_ ;
	wire _w520_ ;
	wire _w521_ ;
	wire _w590_ ;
	wire _w591_ ;
	wire _w592_ ;
	wire _w593_ ;
	wire _w594_ ;
	wire _w595_ ;
	wire _w596_ ;
	wire _w597_ ;
	wire _w598_ ;
	wire _w599_ ;
	wire _w600_ ;
	wire _w601_ ;
	wire _w602_ ;
	wire _w603_ ;
	wire _w604_ ;
	wire _w605_ ;
	wire _w606_ ;
	wire _w607_ ;
	wire _w608_ ;
	wire _w609_ ;
	wire _w610_ ;
	wire _w611_ ;
	wire _w612_ ;
	wire _w613_ ;
	wire _w614_ ;
	wire _w615_ ;
	wire _w616_ ;
	wire _w617_ ;
	wire _w618_ ;
	wire _w619_ ;
	wire _w620_ ;
	wire _w621_ ;
	wire _w622_ ;
	wire _w623_ ;
	wire _w624_ ;
	wire _w625_ ;
	wire _w626_ ;
	wire _w627_ ;
	wire _w628_ ;
	wire _w629_ ;
	wire _w630_ ;
	wire _w631_ ;
	wire _w632_ ;
	wire _w633_ ;
	wire _w634_ ;
	wire _w635_ ;
	wire _w636_ ;
	wire _w637_ ;
	wire _w638_ ;
	wire _w639_ ;
	wire _w640_ ;
	wire _w641_ ;
	wire _w642_ ;
	wire _w643_ ;
	wire _w644_ ;
	wire _w645_ ;
	wire _w646_ ;
	wire _w647_ ;
	wire _w648_ ;
	wire _w649_ ;
	wire _w650_ ;
	wire _w651_ ;
	wire _w652_ ;
	wire _w653_ ;
	wire _w654_ ;
	wire _w655_ ;
	wire _w656_ ;
	wire _w657_ ;
	wire _w658_ ;
	wire _w659_ ;
	wire _w660_ ;
	wire _w661_ ;
	wire _w662_ ;
	wire _w663_ ;
	wire _w664_ ;
	wire _w665_ ;
	wire _w666_ ;
	wire _w667_ ;
	wire _w668_ ;
	wire _w669_ ;
	wire _w670_ ;
	wire _w671_ ;
	wire _w672_ ;
	wire _w673_ ;
	wire _w674_ ;
	wire _w675_ ;
	wire _w676_ ;
	wire _w677_ ;
	wire _w678_ ;
	wire _w679_ ;
	wire _w680_ ;
	wire _w681_ ;
	wire _w682_ ;
	wire _w683_ ;
	wire _w684_ ;
	wire _w685_ ;
	wire _w686_ ;
	wire _w687_ ;
	wire _w688_ ;
	wire _w689_ ;
	wire _w690_ ;
	wire _w691_ ;
	wire _w692_ ;
	wire _w693_ ;
	wire _w694_ ;
	wire _w695_ ;
	wire _w696_ ;
	wire _w697_ ;
	wire _w698_ ;
	wire _w699_ ;
	wire _w700_ ;
	wire _w701_ ;
	wire _w702_ ;
	wire _w703_ ;
	wire _w704_ ;
	wire _w705_ ;
	wire _w706_ ;
	wire _w707_ ;
	wire _w708_ ;
	wire _w709_ ;
	wire _w710_ ;
	wire _w711_ ;
	wire _w712_ ;
	wire _w713_ ;
	wire _w714_ ;
	wire _w715_ ;
	wire _w716_ ;
	wire _w717_ ;
	wire _w718_ ;
	wire _w719_ ;
	wire _w1004_ ;
	wire _w1005_ ;
	wire _w1006_ ;
	wire _w1007_ ;
	wire _w1008_ ;
	wire _w1009_ ;
	wire _w1010_ ;
	wire _w1011_ ;
	wire _w1012_ ;
	wire _w1013_ ;
	wire _w1014_ ;
	wire _w1015_ ;
	wire _w1016_ ;
	wire _w1017_ ;
	wire _w1018_ ;
	wire _w1019_ ;
	wire _w1020_ ;
	wire _w1021_ ;
	wire _w1022_ ;
	wire _w1023_ ;
	wire _w1024_ ;
	wire _w1025_ ;
	wire _w1026_ ;
	wire _w1027_ ;
	wire _w1028_ ;
	wire _w1029_ ;
	wire _w1030_ ;
	wire _w1031_ ;
	wire _w1032_ ;
	wire _w1033_ ;
	wire _w1034_ ;
	wire _w1035_ ;
	wire _w1036_ ;
	wire _w1037_ ;
	wire _w1038_ ;
	wire _w1039_ ;
	wire _w1040_ ;
	wire _w1041_ ;
	wire _w1042_ ;
	wire _w1043_ ;
	wire _w1044_ ;
	wire _w1045_ ;
	wire _w1046_ ;
	wire _w1047_ ;
	wire _w1048_ ;
	wire _w1049_ ;
	wire _w1050_ ;
	wire _w1051_ ;
	wire _w1052_ ;
	wire _w1053_ ;
	wire _w1054_ ;
	wire _w1055_ ;
	wire _w1056_ ;
	wire _w1057_ ;
	wire _w1058_ ;
	wire _w1059_ ;
	wire _w1060_ ;
	wire _w1061_ ;
	wire _w1062_ ;
	wire _w1063_ ;
	wire _w1064_ ;
	wire _w1065_ ;
	wire _w1066_ ;
	wire _w1067_ ;
	wire _w1068_ ;
	wire _w1069_ ;
	wire _w1070_ ;
	wire _w1071_ ;
	wire _w1072_ ;
	wire _w1073_ ;
	wire _w1074_ ;
	wire _w1075_ ;
	wire _w1076_ ;
	wire _w1077_ ;
	wire _w1078_ ;
	wire _w1079_ ;
	wire _w1080_ ;
	wire _w1081_ ;
	wire _w1082_ ;
	wire _w1083_ ;
	wire _w1084_ ;
	wire _w1085_ ;
	wire _w1086_ ;
	wire _w1087_ ;
	wire _w1088_ ;
	wire _w1089_ ;
	wire _w1090_ ;
	wire _w1091_ ;
	wire _w1092_ ;
	wire _w1093_ ;
	wire _w1094_ ;
	wire _w1095_ ;
	wire _w1096_ ;
	wire _w1097_ ;
	wire _w1098_ ;
	wire _w1099_ ;
	wire _w1100_ ;
	wire _w1101_ ;
	wire _w1102_ ;
	wire _w1103_ ;
	wire _w1104_ ;
	wire _w1105_ ;
	wire _w1106_ ;
	wire _w1107_ ;
	wire _w1108_ ;
	wire _w1109_ ;
	wire _w1110_ ;
	wire _w1111_ ;
	wire _w1112_ ;
	wire _w1113_ ;
	wire _w1114_ ;
	wire _w1115_ ;
	wire _w1116_ ;
	wire _w1117_ ;
	wire _w1118_ ;
	wire _w1119_ ;
	wire _w1120_ ;
	wire _w1121_ ;
	wire _w1122_ ;
	wire _w1123_ ;
	wire _w1124_ ;
	wire _w1125_ ;
	wire _w1126_ ;
	wire _w1127_ ;
	wire _w1128_ ;
	wire _w1129_ ;
	wire _w1130_ ;
	wire _w1131_ ;
	wire _w1132_ ;
	wire _w1133_ ;
	wire _w1134_ ;
	wire _w1135_ ;
	wire _w1136_ ;
	wire _w1137_ ;
	wire _w1138_ ;
	wire _w1139_ ;
	wire _w1140_ ;
	wire _w1141_ ;
	wire _w1142_ ;
	wire _w1143_ ;
	wire _w1144_ ;
	wire _w1145_ ;
	wire _w1146_ ;
	wire _w1147_ ;
	wire _w1148_ ;
	wire _w1149_ ;
	wire _w1150_ ;
	wire _w1151_ ;
	wire _w1152_ ;
	wire _w1153_ ;
	wire _w1154_ ;
	wire _w1155_ ;
	wire _w1156_ ;
	wire _w1157_ ;
	wire _w1158_ ;
	wire _w1159_ ;
	wire _w1160_ ;
	wire _w1161_ ;
	wire _w1162_ ;
	wire _w1163_ ;
	wire _w1164_ ;
	wire _w1165_ ;
	wire _w1166_ ;
	wire _w1167_ ;
	wire _w1168_ ;
	wire _w1169_ ;
	wire _w1170_ ;
	wire _w1171_ ;
	wire _w1172_ ;
	wire _w1173_ ;
	wire _w1174_ ;
	wire _w1175_ ;
	wire _w1176_ ;
	wire _w1177_ ;
	wire _w1178_ ;
	wire _w1179_ ;
	wire _w1180_ ;
	wire _w1181_ ;
	wire _w1182_ ;
	wire _w1183_ ;
	wire _w1184_ ;
	wire _w1185_ ;
	wire _w1186_ ;
	wire _w1187_ ;
	wire _w1188_ ;
	wire _w1189_ ;
	wire _w1190_ ;
	wire _w1191_ ;
	wire _w1192_ ;
	wire _w1193_ ;
	wire _w1194_ ;
	wire _w1195_ ;
	wire _w1196_ ;
	wire _w1197_ ;
	wire _w1198_ ;
	wire _w1199_ ;
	wire _w1200_ ;
	wire _w1201_ ;
	wire _w1202_ ;
	wire _w1203_ ;
	wire _w1204_ ;
	wire _w1205_ ;
	wire _w1206_ ;
	wire _w1207_ ;
	wire _w1208_ ;
	wire _w1209_ ;
	wire _w1210_ ;
	wire _w1211_ ;
	wire _w1212_ ;
	wire _w1213_ ;
	wire _w1214_ ;
	wire _w1215_ ;
	wire _w1216_ ;
	wire _w1217_ ;
	wire _w1218_ ;
	wire _w1219_ ;
	wire _w1220_ ;
	wire _w1221_ ;
	wire _w1222_ ;
	wire _w1223_ ;
	wire _w1224_ ;
	wire _w1225_ ;
	wire _w1226_ ;
	wire _w1227_ ;
	wire _w1228_ ;
	wire _w1229_ ;
	wire _w1230_ ;
	wire _w1231_ ;
	wire _w1232_ ;
	wire _w1233_ ;
	wire _w1234_ ;
	wire _w1235_ ;
	wire _w1236_ ;
	wire _w1237_ ;
	wire _w1238_ ;
	wire _w1239_ ;
	wire _w1240_ ;
	wire _w1241_ ;
	wire _w1242_ ;
	wire _w1243_ ;
	wire _w1244_ ;
	wire _w1245_ ;
	wire _w1246_ ;
	wire _w1247_ ;
	wire _w1248_ ;
	wire _w1249_ ;
	wire _w1250_ ;
	wire _w1251_ ;
	wire _w1252_ ;
	wire _w1253_ ;
	wire _w1254_ ;
	wire _w1255_ ;
	wire _w1256_ ;
	wire _w1257_ ;
	wire _w1258_ ;
	wire _w1259_ ;
	wire _w1260_ ;
	wire _w1261_ ;
	wire _w1262_ ;
	wire _w1263_ ;
	wire _w1264_ ;
	wire _w1265_ ;
	wire _w1266_ ;
	wire _w1267_ ;
	wire _w1268_ ;
	wire _w1269_ ;
	wire _w1270_ ;
	wire _w1271_ ;
	wire _w1272_ ;
	wire _w1273_ ;
	wire _w1274_ ;
	wire _w1275_ ;
	wire _w1276_ ;
	wire _w1277_ ;
	wire _w1278_ ;
	wire _w1279_ ;
	wire _w1280_ ;
	wire _w1281_ ;
	wire _w1282_ ;
	wire _w1283_ ;
	wire _w1284_ ;
	wire _w1285_ ;
	wire _w1286_ ;
	wire _w1287_ ;
	wire _w1288_ ;
	wire _w1289_ ;
	wire _w1290_ ;
	wire _w1291_ ;
	wire _w1292_ ;
	wire _w1293_ ;
	wire _w1294_ ;
	wire _w1295_ ;
	wire _w1296_ ;
	wire _w1297_ ;
	wire _w1298_ ;
	wire _w1299_ ;
	wire _w1300_ ;
	wire _w1301_ ;
	wire _w1302_ ;
	wire _w1303_ ;
	wire _w1304_ ;
	wire _w1305_ ;
	wire _w1306_ ;
	wire _w1307_ ;
	wire _w1308_ ;
	wire _w1309_ ;
	wire _w1310_ ;
	wire _w1311_ ;
	wire _w1312_ ;
	wire _w1313_ ;
	wire _w1314_ ;
	wire _w1315_ ;
	wire _w1316_ ;
	wire _w1317_ ;
	wire _w1318_ ;
	wire _w1319_ ;
	wire _w1320_ ;
	wire _w1321_ ;
	wire _w1322_ ;
	wire _w1323_ ;
	wire _w1324_ ;
	wire _w1326_ ;
	wire _w1327_ ;
	wire _w1328_ ;
	wire _w1329_ ;
	wire _w1330_ ;
	wire _w1331_ ;
	wire _w1332_ ;
	wire _w1333_ ;
	wire _w1334_ ;
	wire _w1335_ ;
	wire _w1336_ ;
	wire _w1337_ ;
	wire _w1338_ ;
	wire _w1339_ ;
	wire _w1340_ ;
	wire _w1341_ ;
	wire _w1342_ ;
	wire _w1343_ ;
	wire _w1344_ ;
	wire _w1345_ ;
	wire _w1346_ ;
	wire _w1347_ ;
	wire _w1348_ ;
	wire _w1349_ ;
	wire _w1350_ ;
	wire _w1351_ ;
	wire _w1352_ ;
	wire _w1353_ ;
	wire _w1354_ ;
	wire _w1355_ ;
	wire _w1356_ ;
	wire _w1357_ ;
	wire _w1358_ ;
	wire _w1359_ ;
	wire _w1360_ ;
	wire _w1361_ ;
	wire _w1362_ ;
	wire _w1363_ ;
	wire _w1364_ ;
	wire _w1365_ ;
	wire _w1366_ ;
	wire _w1367_ ;
	wire _w1368_ ;
	wire _w1369_ ;
	wire _w1370_ ;
	wire _w1371_ ;
	wire _w1372_ ;
	wire _w1373_ ;
	wire _w1374_ ;
	wire _w1375_ ;
	wire _w1376_ ;
	wire _w1377_ ;
	wire _w1378_ ;
	wire _w1379_ ;
	wire _w1380_ ;
	wire _w1381_ ;
	wire _w1382_ ;
	wire _w1383_ ;
	wire _w1384_ ;
	wire _w1385_ ;
	wire _w1386_ ;
	wire _w1387_ ;
	wire _w1388_ ;
	wire _w1389_ ;
	wire _w1390_ ;
	wire _w1391_ ;
	wire _w1392_ ;
	wire _w1393_ ;
	wire _w1394_ ;
	wire _w1395_ ;
	wire _w1396_ ;
	wire _w1397_ ;
	wire _w1398_ ;
	wire _w1399_ ;
	wire _w1400_ ;
	wire _w1401_ ;
	wire _w1402_ ;
	wire _w1403_ ;
	wire _w1404_ ;
	wire _w1405_ ;
	wire _w1406_ ;
	wire _w1407_ ;
	wire _w1408_ ;
	wire _w1409_ ;
	wire _w1410_ ;
	wire _w1411_ ;
	wire _w1412_ ;
	wire _w1413_ ;
	wire _w1414_ ;
	wire _w1415_ ;
	wire _w1416_ ;
	wire _w1417_ ;
	wire _w1418_ ;
	wire _w1419_ ;
	wire _w1420_ ;
	wire _w1421_ ;
	wire _w1422_ ;
	wire _w1423_ ;
	wire _w1424_ ;
	wire _w1425_ ;
	wire _w1426_ ;
	wire _w1427_ ;
	wire _w1428_ ;
	wire _w1429_ ;
	wire _w1430_ ;
	wire _w1431_ ;
	wire _w1432_ ;
	wire _w1433_ ;
	wire _w1434_ ;
	wire _w1435_ ;
	wire _w1436_ ;
	wire _w1437_ ;
	wire _w1438_ ;
	wire _w1439_ ;
	wire _w1440_ ;
	wire _w1441_ ;
	wire _w1442_ ;
	wire _w1443_ ;
	wire _w1444_ ;
	wire _w1445_ ;
	wire _w1446_ ;
	wire _w1447_ ;
	wire _w1448_ ;
	wire _w1449_ ;
	wire _w1450_ ;
	wire _w1451_ ;
	wire _w1452_ ;
	wire _w1453_ ;
	wire _w1454_ ;
	wire _w1455_ ;
	wire _w1456_ ;
	wire _w1457_ ;
	wire _w1458_ ;
	wire _w1459_ ;
	wire _w1460_ ;
	wire _w1461_ ;
	wire _w1462_ ;
	wire _w1463_ ;
	wire _w1464_ ;
	wire _w1465_ ;
	wire _w1466_ ;
	wire _w1467_ ;
	wire _w1468_ ;
	wire _w1469_ ;
	wire _w1470_ ;
	wire _w1471_ ;
	wire _w1472_ ;
	wire _w1473_ ;
	wire _w1474_ ;
	wire _w1475_ ;
	wire _w1476_ ;
	wire _w1477_ ;
	wire _w1478_ ;
	wire _w1479_ ;
	wire _w1480_ ;
	wire _w1481_ ;
	wire _w1482_ ;
	wire _w1483_ ;
	wire _w1484_ ;
	wire _w1485_ ;
	wire _w1486_ ;
	wire _w1487_ ;
	wire _w1488_ ;
	wire _w1489_ ;
	wire _w1490_ ;
	wire _w1491_ ;
	wire _w1492_ ;
	wire _w1493_ ;
	wire _w1494_ ;
	wire _w1495_ ;
	wire _w1496_ ;
	wire _w1497_ ;
	wire _w1498_ ;
	wire _w1499_ ;
	wire _w1500_ ;
	wire _w1501_ ;
	wire _w1502_ ;
	wire _w1503_ ;
	wire _w1504_ ;
	wire _w1505_ ;
	wire _w1506_ ;
	wire _w1507_ ;
	wire _w1508_ ;
	wire _w1509_ ;
	wire _w1510_ ;
	wire _w1511_ ;
	wire _w1512_ ;
	wire _w1513_ ;
	wire _w1514_ ;
	wire _w1515_ ;
	wire _w1516_ ;
	wire _w1517_ ;
	wire _w1518_ ;
	wire _w1519_ ;
	wire _w1520_ ;
	wire _w1521_ ;
	wire _w1522_ ;
	wire _w1523_ ;
	wire _w1524_ ;
	wire _w1525_ ;
	wire _w1526_ ;
	wire _w1527_ ;
	wire _w1528_ ;
	wire _w1529_ ;
	wire _w1530_ ;
	wire _w1531_ ;
	wire _w1532_ ;
	wire _w1533_ ;
	wire _w1534_ ;
	wire _w1535_ ;
	wire _w1536_ ;
	wire _w1537_ ;
	wire _w1538_ ;
	wire _w1539_ ;
	wire _w1540_ ;
	wire _w1541_ ;
	wire _w1542_ ;
	wire _w1543_ ;
	wire _w1544_ ;
	wire _w1545_ ;
	wire _w1546_ ;
	wire _w1547_ ;
	wire _w1548_ ;
	wire _w1549_ ;
	wire _w1550_ ;
	wire _w1551_ ;
	wire _w1552_ ;
	wire _w1553_ ;
	wire _w1554_ ;
	wire _w1555_ ;
	wire _w1556_ ;
	wire _w1557_ ;
	wire _w1558_ ;
	wire _w1559_ ;
	wire _w1560_ ;
	wire _w1561_ ;
	wire _w1562_ ;
	wire _w1563_ ;
	wire _w1564_ ;
	wire _w1565_ ;
	wire _w1566_ ;
	wire _w1567_ ;
	wire _w1568_ ;
	wire _w1569_ ;
	wire _w1570_ ;
	wire _w1571_ ;
	wire _w2820_ ;
	wire _w2821_ ;
	wire _w2822_ ;
	wire _w2823_ ;
	wire _w2824_ ;
	wire _w2825_ ;
	wire _w2826_ ;
	wire _w2827_ ;
	wire _w2828_ ;
	wire _w2829_ ;
	wire _w2830_ ;
	wire _w2831_ ;
	wire _w2832_ ;
	wire _w2833_ ;
	wire _w2834_ ;
	wire _w2835_ ;
	wire _w2836_ ;
	wire _w2837_ ;
	wire _w2838_ ;
	wire _w2839_ ;
	wire _w2840_ ;
	wire _w2841_ ;
	wire _w2842_ ;
	wire _w2843_ ;
	wire _w2844_ ;
	wire _w2845_ ;
	wire _w2846_ ;
	wire _w2847_ ;
	wire _w2848_ ;
	wire _w2849_ ;
	wire _w2850_ ;
	wire _w2851_ ;
	wire _w2852_ ;
	wire _w2853_ ;
	wire _w2854_ ;
	wire _w2855_ ;
	wire _w2856_ ;
	wire _w2857_ ;
	wire _w2858_ ;
	wire _w2859_ ;
	wire _w2860_ ;
	wire _w2861_ ;
	wire _w2862_ ;
	wire _w2863_ ;
	wire _w2864_ ;
	wire _w2865_ ;
	wire _w2866_ ;
	wire _w2867_ ;
	wire _w2868_ ;
	wire _w2869_ ;
	wire _w2870_ ;
	wire _w2871_ ;
	wire _w2872_ ;
	wire _w2873_ ;
	wire _w2874_ ;
	wire _w2875_ ;
	wire _w2876_ ;
	wire _w2877_ ;
	wire _w2878_ ;
	wire _w2879_ ;
	wire _w2880_ ;
	wire _w2881_ ;
	wire _w2882_ ;
	wire _w2883_ ;
	wire _w2884_ ;
	wire _w2885_ ;
	wire _w2886_ ;
	wire _w2887_ ;
	wire _w2888_ ;
	wire _w2889_ ;
	wire _w2890_ ;
	wire _w2891_ ;
	wire _w2892_ ;
	wire _w2893_ ;
	wire _w2894_ ;
	wire _w2895_ ;
	wire _w2896_ ;
	wire _w2897_ ;
	wire _w2898_ ;
	wire _w2899_ ;
	wire _w2900_ ;
	wire _w2901_ ;
	wire _w2902_ ;
	wire _w2903_ ;
	wire _w2904_ ;
	wire _w2905_ ;
	wire _w2906_ ;
	wire _w2907_ ;
	wire _w2908_ ;
	wire _w2909_ ;
	wire _w2910_ ;
	wire _w2911_ ;
	wire _w2912_ ;
	wire _w2913_ ;
	wire _w2914_ ;
	wire _w2915_ ;
	wire _w2916_ ;
	wire _w2917_ ;
	wire _w2918_ ;
	wire _w2919_ ;
	wire _w2920_ ;
	wire _w2921_ ;
	wire _w2922_ ;
	wire _w2923_ ;
	wire _w2924_ ;
	wire _w2925_ ;
	wire _w2926_ ;
	wire _w2927_ ;
	wire _w2928_ ;
	wire _w2929_ ;
	wire _w2930_ ;
	wire _w2931_ ;
	wire _w2932_ ;
	wire _w2933_ ;
	wire _w2934_ ;
	wire _w2935_ ;
	wire _w2936_ ;
	wire _w2937_ ;
	wire _w2938_ ;
	wire _w2939_ ;
	wire _w2940_ ;
	wire _w2941_ ;
	wire _w2942_ ;
	wire _w2943_ ;
	wire _w2944_ ;
	wire _w2945_ ;
	wire _w2946_ ;
	wire _w2947_ ;
	wire _w2948_ ;
	wire _w2949_ ;
	wire _w2950_ ;
	wire _w2951_ ;
	wire _w2952_ ;
	wire _w2953_ ;
	wire _w2954_ ;
	wire _w2955_ ;
	wire _w2956_ ;
	wire _w2957_ ;
	wire _w2958_ ;
	wire _w2959_ ;
	wire _w2960_ ;
	wire _w2961_ ;
	wire _w2962_ ;
	wire _w2963_ ;
	wire _w2964_ ;
	wire _w2965_ ;
	wire _w2966_ ;
	wire _w2967_ ;
	wire _w2968_ ;
	wire _w2969_ ;
	wire _w2970_ ;
	wire _w2971_ ;
	wire _w2972_ ;
	wire _w2973_ ;
	wire _w2974_ ;
	wire _w2975_ ;
	wire _w2976_ ;
	wire _w2977_ ;
	wire _w2978_ ;
	wire _w2979_ ;
	wire _w2980_ ;
	wire _w2981_ ;
	wire _w2982_ ;
	wire _w2983_ ;
	wire _w2984_ ;
	wire _w2985_ ;
	wire _w2986_ ;
	wire _w2987_ ;
	wire _w2988_ ;
	wire _w2989_ ;
	wire _w2990_ ;
	wire _w2991_ ;
	wire _w2992_ ;
	wire _w2993_ ;
	wire _w2994_ ;
	wire _w2995_ ;
	wire _w2996_ ;
	wire _w2997_ ;
	wire _w2998_ ;
	wire _w2999_ ;
	wire _w3000_ ;
	wire _w3001_ ;
	wire _w3002_ ;
	wire _w3003_ ;
	wire _w3004_ ;
	wire _w3005_ ;
	wire _w3006_ ;
	wire _w3007_ ;
	wire _w3008_ ;
	wire _w3009_ ;
	wire _w3010_ ;
	wire _w3011_ ;
	wire _w3012_ ;
	wire _w3013_ ;
	wire _w3014_ ;
	wire _w3015_ ;
	wire _w3016_ ;
	wire _w3017_ ;
	wire _w3018_ ;
	wire _w3019_ ;
	wire _w3020_ ;
	wire _w3021_ ;
	wire _w3022_ ;
	wire _w3023_ ;
	wire _w3024_ ;
	wire _w3025_ ;
	wire _w3026_ ;
	wire _w3027_ ;
	wire _w3028_ ;
	wire _w3029_ ;
	wire _w3030_ ;
	wire _w3031_ ;
	wire _w3032_ ;
	wire _w3033_ ;
	wire _w3034_ ;
	wire _w3035_ ;
	wire _w3036_ ;
	wire _w3037_ ;
	wire _w3038_ ;
	wire _w3039_ ;
	wire _w3040_ ;
	wire _w3041_ ;
	wire _w3042_ ;
	wire _w3043_ ;
	wire _w3044_ ;
	wire _w3045_ ;
	wire _w3046_ ;
	wire _w3047_ ;
	wire _w3048_ ;
	wire _w3049_ ;
	wire _w3050_ ;
	wire _w3051_ ;
	wire _w3052_ ;
	wire _w3053_ ;
	wire _w3054_ ;
	wire _w3055_ ;
	wire _w3056_ ;
	wire _w3057_ ;
	wire _w3058_ ;
	wire _w3059_ ;
	wire _w3060_ ;
	wire _w3061_ ;
	wire _w3062_ ;
	wire _w3063_ ;
	wire _w3064_ ;
	wire _w3065_ ;
	wire _w3066_ ;
	wire _w3067_ ;
	wire _w3068_ ;
	wire _w3069_ ;
	wire _w3070_ ;
	wire _w3071_ ;
	wire _w3072_ ;
	wire _w3073_ ;
	wire _w3074_ ;
	wire _w3075_ ;
	wire _w3076_ ;
	wire _w3077_ ;
	wire _w3078_ ;
	wire _w3079_ ;
	wire _w3080_ ;
	wire _w3081_ ;
	wire _w3082_ ;
	wire _w3083_ ;
	wire _w3084_ ;
	wire _w3085_ ;
	wire _w3086_ ;
	wire _w3087_ ;
	wire _w3088_ ;
	wire _w3089_ ;
	wire _w3090_ ;
	wire _w3091_ ;
	wire _w3092_ ;
	wire _w3093_ ;
	wire _w3094_ ;
	wire _w3095_ ;
	wire _w3096_ ;
	wire _w3097_ ;
	wire _w3098_ ;
	wire _w3099_ ;
	wire _w3100_ ;
	wire _w3101_ ;
	wire _w3102_ ;
	wire _w3103_ ;
	wire _w3104_ ;
	wire _w3105_ ;
	wire _w3106_ ;
	wire _w3107_ ;
	wire _w3108_ ;
	wire _w3109_ ;
	wire _w3110_ ;
	wire _w3111_ ;
	wire _w3112_ ;
	wire _w3113_ ;
	wire _w3114_ ;
	wire _w3115_ ;
	wire _w3116_ ;
	wire _w3117_ ;
	wire _w3118_ ;
	wire _w3119_ ;
	wire _w3120_ ;
	wire _w3121_ ;
	wire _w3122_ ;
	wire _w3123_ ;
	wire _w3124_ ;
	wire _w3125_ ;
	wire _w3126_ ;
	wire _w3127_ ;
	wire _w3128_ ;
	wire _w3129_ ;
	wire _w3130_ ;
	wire _w3131_ ;
	wire _w3132_ ;
	wire _w3133_ ;
	wire _w3134_ ;
	wire _w3135_ ;
	wire _w3136_ ;
	wire _w3137_ ;
	wire _w3138_ ;
	wire _w3139_ ;
	wire _w3140_ ;
	wire _w3141_ ;
	wire _w3142_ ;
	wire _w3143_ ;
	wire _w3144_ ;
	wire _w3145_ ;
	wire _w3146_ ;
	wire _w3147_ ;
	wire _w3148_ ;
	wire _w3149_ ;
	wire _w3150_ ;
	wire _w3151_ ;
	wire _w3152_ ;
	wire _w3153_ ;
	wire _w3154_ ;
	wire _w3155_ ;
	wire _w3156_ ;
	wire _w3157_ ;
	wire _w3158_ ;
	wire _w3159_ ;
	wire _w3160_ ;
	wire _w3161_ ;
	wire _w3162_ ;
	wire _w3163_ ;
	wire _w3164_ ;
	wire _w3165_ ;
	wire _w3166_ ;
	wire _w3167_ ;
	wire _w3168_ ;
	wire _w3169_ ;
	wire _w3170_ ;
	wire _w3171_ ;
	wire _w3172_ ;
	wire _w3173_ ;
	wire _w3174_ ;
	wire _w3175_ ;
	wire _w3176_ ;
	wire _w3177_ ;
	wire _w3178_ ;
	wire _w3179_ ;
	wire _w3180_ ;
	wire _w3181_ ;
	wire _w3182_ ;
	wire _w3183_ ;
	wire _w3184_ ;
	wire _w3185_ ;
	wire _w3186_ ;
	wire _w3187_ ;
	wire _w3188_ ;
	wire _w3189_ ;
	wire _w3190_ ;
	wire _w3191_ ;
	wire _w3192_ ;
	wire _w3193_ ;
	wire _w3194_ ;
	wire _w3195_ ;
	wire _w3196_ ;
	wire _w3197_ ;
	wire _w3198_ ;
	wire _w3199_ ;
	wire _w3200_ ;
	wire _w3201_ ;
	wire _w3202_ ;
	wire _w3203_ ;
	wire _w3204_ ;
	wire _w3205_ ;
	wire _w3206_ ;
	wire _w3207_ ;
	wire _w3208_ ;
	wire _w3209_ ;
	wire _w3210_ ;
	wire _w3211_ ;
	wire _w3212_ ;
	wire _w3213_ ;
	wire _w3214_ ;
	wire _w3215_ ;
	wire _w3216_ ;
	wire _w3217_ ;
	wire _w3218_ ;
	wire _w3219_ ;
	wire _w3220_ ;
	wire _w3221_ ;
	wire _w3222_ ;
	wire _w3223_ ;
	wire _w3224_ ;
	wire _w3225_ ;
	wire _w3226_ ;
	wire _w3227_ ;
	wire _w3228_ ;
	wire _w3229_ ;
	wire _w3230_ ;
	wire _w3231_ ;
	wire _w3232_ ;
	wire _w3233_ ;
	wire _w3234_ ;
	wire _w3235_ ;
	wire _w3236_ ;
	wire _w3237_ ;
	wire _w3238_ ;
	wire _w3239_ ;
	wire _w3240_ ;
	wire _w3241_ ;
	wire _w3242_ ;
	wire _w3243_ ;
	wire _w3244_ ;
	wire _w3245_ ;
	wire _w3246_ ;
	wire _w3247_ ;
	wire _w3248_ ;
	wire _w3249_ ;
	wire _w3250_ ;
	wire _w3251_ ;
	wire _w3252_ ;
	wire _w3253_ ;
	wire _w3254_ ;
	wire _w3255_ ;
	wire _w3256_ ;
	wire _w3257_ ;
	wire _w3258_ ;
	wire _w3259_ ;
	wire _w3260_ ;
	wire _w3261_ ;
	wire _w3262_ ;
	wire _w3263_ ;
	wire _w3264_ ;
	wire _w3265_ ;
	wire _w3266_ ;
	wire _w3267_ ;
	wire _w3268_ ;
	wire _w3269_ ;
	wire _w3270_ ;
	wire _w3271_ ;
	wire _w3272_ ;
	wire _w3273_ ;
	wire _w3274_ ;
	wire _w3275_ ;
	wire _w3276_ ;
	wire _w3277_ ;
	wire _w3278_ ;
	wire _w3279_ ;
	wire _w3280_ ;
	wire _w3281_ ;
	wire _w3282_ ;
	wire _w3283_ ;
	wire _w3284_ ;
	wire _w3285_ ;
	wire _w3286_ ;
	wire _w3287_ ;
	wire _w3288_ ;
	wire _w3289_ ;
	wire _w3290_ ;
	wire _w3291_ ;
	wire _w3292_ ;
	wire _w3293_ ;
	wire _w3294_ ;
	wire _w3295_ ;
	wire _w3296_ ;
	wire _w3297_ ;
	wire _w3298_ ;
	wire _w3299_ ;
	wire _w3300_ ;
	wire _w3301_ ;
	wire _w3302_ ;
	wire _w3303_ ;
	wire _w3304_ ;
	wire _w3305_ ;
	wire _w3306_ ;
	wire _w3307_ ;
	wire _w3308_ ;
	wire _w3309_ ;
	wire _w3310_ ;
	wire _w3311_ ;
	wire _w3312_ ;
	wire _w3313_ ;
	wire _w3314_ ;
	wire _w3315_ ;
	wire _w3316_ ;
	wire _w3317_ ;
	wire _w3318_ ;
	wire _w3319_ ;
	wire _w3320_ ;
	wire _w3321_ ;
	wire _w3322_ ;
	wire _w3323_ ;
	wire _w3324_ ;
	wire _w3325_ ;
	wire _w3326_ ;
	wire _w3327_ ;
	wire _w3328_ ;
	wire _w3329_ ;
	wire _w3330_ ;
	wire _w3331_ ;
	wire _w3332_ ;
	wire _w3333_ ;
	wire _w3334_ ;
	wire _w3335_ ;
	wire _w3336_ ;
	wire _w3337_ ;
	wire _w3338_ ;
	wire _w3339_ ;
	wire _w3340_ ;
	wire _w3341_ ;
	wire _w3342_ ;
	wire _w3343_ ;
	wire _w3344_ ;
	wire _w3345_ ;
	wire _w3346_ ;
	wire _w3347_ ;
	wire _w3348_ ;
	wire _w3349_ ;
	wire _w3350_ ;
	wire _w3351_ ;
	wire _w3352_ ;
	wire _w3353_ ;
	wire _w3354_ ;
	wire _w3355_ ;
	wire _w3356_ ;
	wire _w3357_ ;
	wire _w3358_ ;
	wire _w3359_ ;
	wire _w3360_ ;
	wire _w3361_ ;
	wire _w3362_ ;
	wire _w3363_ ;
	wire _w3364_ ;
	wire _w3365_ ;
	wire _w3366_ ;
	wire _w3367_ ;
	wire _w3368_ ;
	wire _w3369_ ;
	wire _w3370_ ;
	wire _w3371_ ;
	wire _w3372_ ;
	wire _w3373_ ;
	wire _w3374_ ;
	wire _w3375_ ;
	wire _w3376_ ;
	wire _w3377_ ;
	wire _w3378_ ;
	wire _w3379_ ;
	wire _w3380_ ;
	wire _w3381_ ;
	wire _w3382_ ;
	wire _w3383_ ;
	wire _w3384_ ;
	wire _w3385_ ;
	wire _w3386_ ;
	wire _w3387_ ;
	wire _w3388_ ;
	wire _w3389_ ;
	wire _w3390_ ;
	wire _w3391_ ;
	wire _w3392_ ;
	wire _w3393_ ;
	wire _w3394_ ;
	wire _w3395_ ;
	wire _w3396_ ;
	wire _w3397_ ;
	wire _w3398_ ;
	wire _w3399_ ;
	wire _w3400_ ;
	wire _w3401_ ;
	wire _w3402_ ;
	wire _w3403_ ;
	wire _w3404_ ;
	wire _w3405_ ;
	wire _w3406_ ;
	wire _w3407_ ;
	wire _w3408_ ;
	wire _w3409_ ;
	wire _w3410_ ;
	wire _w3411_ ;
	wire _w3412_ ;
	wire _w3413_ ;
	wire _w3414_ ;
	wire _w3415_ ;
	wire _w3416_ ;
	wire _w3417_ ;
	wire _w3418_ ;
	wire _w3419_ ;
	wire _w3420_ ;
	wire _w3421_ ;
	wire _w3422_ ;
	wire _w3423_ ;
	wire _w3424_ ;
	wire _w3425_ ;
	wire _w3426_ ;
	wire _w3427_ ;
	wire _w3428_ ;
	wire _w3429_ ;
	wire _w3430_ ;
	wire _w3431_ ;
	wire _w3432_ ;
	wire _w3433_ ;
	wire _w3434_ ;
	wire _w3435_ ;
	wire _w3436_ ;
	wire _w3437_ ;
	wire _w3438_ ;
	wire _w3439_ ;
	wire _w3440_ ;
	wire _w3441_ ;
	wire _w3442_ ;
	wire _w3443_ ;
	wire _w3444_ ;
	wire _w3445_ ;
	wire _w3446_ ;
	wire _w3447_ ;
	wire _w3448_ ;
	wire _w3449_ ;
	wire _w3450_ ;
	wire _w3451_ ;
	wire _w3452_ ;
	wire _w3453_ ;
	wire _w3454_ ;
	wire _w3455_ ;
	wire _w3456_ ;
	wire _w3457_ ;
	wire _w3458_ ;
	wire _w3459_ ;
	wire _w3460_ ;
	wire _w3461_ ;
	wire _w3462_ ;
	wire _w3463_ ;
	wire _w3464_ ;
	wire _w3465_ ;
	wire _w3466_ ;
	wire _w3467_ ;
	wire _w3468_ ;
	wire _w3469_ ;
	wire _w3470_ ;
	wire _w3471_ ;
	wire _w3472_ ;
	wire _w3473_ ;
	wire _w3474_ ;
	wire _w3475_ ;
	wire _w3476_ ;
	wire _w3477_ ;
	wire _w3478_ ;
	wire _w3479_ ;
	wire _w3480_ ;
	wire _w3481_ ;
	wire _w3482_ ;
	wire _w3483_ ;
	wire _w3484_ ;
	wire _w3485_ ;
	wire _w3486_ ;
	wire _w3487_ ;
	wire _w3488_ ;
	wire _w3489_ ;
	wire _w3490_ ;
	wire _w3491_ ;
	wire _w3492_ ;
	wire _w3493_ ;
	wire _w3494_ ;
	wire _w3495_ ;
	wire _w3496_ ;
	wire _w3497_ ;
	wire _w3498_ ;
	wire _w3499_ ;
	wire _w3500_ ;
	wire _w3501_ ;
	wire _w3502_ ;
	wire _w3503_ ;
	wire _w3504_ ;
	wire _w3505_ ;
	wire _w3506_ ;
	wire _w3507_ ;
	wire _w3508_ ;
	wire _w3509_ ;
	wire _w3510_ ;
	wire _w3511_ ;
	wire _w3512_ ;
	wire _w3513_ ;
	wire _w3514_ ;
	wire _w3515_ ;
	wire _w3516_ ;
	wire _w3517_ ;
	wire _w3518_ ;
	wire _w3519_ ;
	wire _w3520_ ;
	wire _w3521_ ;
	wire _w3522_ ;
	wire _w3523_ ;
	wire _w3524_ ;
	wire _w3525_ ;
	wire _w3526_ ;
	wire _w3527_ ;
	wire _w3528_ ;
	wire _w3529_ ;
	wire _w3530_ ;
	wire _w3531_ ;
	wire _w3532_ ;
	wire _w3533_ ;
	wire _w3534_ ;
	wire _w3535_ ;
	wire _w3536_ ;
	wire _w3537_ ;
	wire _w3538_ ;
	wire _w3539_ ;
	wire _w3540_ ;
	wire _w3541_ ;
	wire _w3542_ ;
	wire _w3543_ ;
	wire _w3544_ ;
	wire _w3545_ ;
	wire _w3546_ ;
	wire _w3547_ ;
	wire _w3548_ ;
	wire _w3549_ ;
	wire _w3550_ ;
	wire _w3551_ ;
	wire _w3552_ ;
	wire _w3553_ ;
	wire _w3554_ ;
	wire _w3555_ ;
	wire _w3556_ ;
	wire _w3557_ ;
	wire _w3558_ ;
	wire _w3559_ ;
	wire _w3560_ ;
	wire _w3561_ ;
	wire _w3562_ ;
	wire _w3563_ ;
	wire _w3564_ ;
	wire _w3565_ ;
	wire _w3566_ ;
	wire _w3567_ ;
	wire _w3568_ ;
	wire _w3569_ ;
	wire _w3570_ ;
	wire _w3571_ ;
	wire _w3572_ ;
	wire _w3573_ ;
	wire _w3574_ ;
	wire _w3575_ ;
	wire _w3576_ ;
	wire _w3577_ ;
	wire _w3578_ ;
	wire _w3579_ ;
	wire _w3580_ ;
	wire _w3581_ ;
	wire _w3582_ ;
	wire _w3583_ ;
	wire _w3584_ ;
	wire _w3585_ ;
	wire _w3586_ ;
	wire _w3587_ ;
	wire _w3588_ ;
	wire _w3589_ ;
	wire _w3590_ ;
	wire _w3591_ ;
	wire _w3592_ ;
	wire _w3593_ ;
	wire _w3594_ ;
	wire _w3595_ ;
	wire _w3596_ ;
	wire _w3597_ ;
	wire _w3598_ ;
	wire _w3599_ ;
	wire _w3600_ ;
	wire _w3601_ ;
	wire _w3602_ ;
	wire _w3603_ ;
	wire _w3604_ ;
	wire _w3605_ ;
	wire _w3606_ ;
	wire _w3607_ ;
	wire _w3608_ ;
	wire _w3609_ ;
	wire _w3610_ ;
	wire _w3611_ ;
	wire _w3612_ ;
	wire _w3613_ ;
	wire _w3614_ ;
	wire _w3615_ ;
	wire _w3616_ ;
	wire _w3617_ ;
	wire _w3618_ ;
	wire _w3619_ ;
	wire _w3620_ ;
	wire _w3621_ ;
	wire _w3622_ ;
	wire _w3623_ ;
	wire _w3624_ ;
	wire _w3625_ ;
	wire _w3626_ ;
	wire _w3627_ ;
	wire _w3628_ ;
	wire _w3629_ ;
	wire _w3630_ ;
	wire _w3631_ ;
	wire _w3632_ ;
	wire _w3633_ ;
	wire _w3634_ ;
	wire _w3635_ ;
	wire _w3636_ ;
	wire _w3637_ ;
	wire _w3638_ ;
	wire _w3639_ ;
	wire _w3640_ ;
	wire _w3641_ ;
	wire _w3642_ ;
	wire _w3643_ ;
	wire _w3644_ ;
	wire _w3645_ ;
	wire _w3646_ ;
	wire _w3647_ ;
	wire _w3648_ ;
	wire _w3649_ ;
	wire _w3650_ ;
	wire _w3651_ ;
	wire _w3652_ ;
	wire _w3653_ ;
	wire _w3654_ ;
	wire _w3655_ ;
	wire _w3656_ ;
	wire _w3657_ ;
	wire _w3658_ ;
	wire _w3659_ ;
	wire _w3660_ ;
	wire _w3661_ ;
	wire _w3662_ ;
	wire _w3663_ ;
	wire _w3664_ ;
	wire _w3665_ ;
	wire _w3666_ ;
	wire _w3667_ ;
	wire _w3668_ ;
	wire _w3669_ ;
	wire _w3670_ ;
	wire _w3671_ ;
	wire _w3672_ ;
	wire _w3673_ ;
	wire _w3674_ ;
	wire _w3675_ ;
	wire _w3676_ ;
	wire _w3677_ ;
	wire _w3678_ ;
	wire _w3679_ ;
	wire _w3680_ ;
	wire _w3681_ ;
	wire _w3682_ ;
	wire _w3683_ ;
	wire _w3684_ ;
	wire _w3685_ ;
	wire _w3686_ ;
	wire _w3687_ ;
	wire _w3688_ ;
	wire _w3689_ ;
	wire _w3690_ ;
	wire _w3691_ ;
	wire _w3692_ ;
	wire _w3693_ ;
	wire _w3694_ ;
	wire _w3695_ ;
	wire _w3696_ ;
	wire _w3697_ ;
	wire _w3698_ ;
	wire _w3699_ ;
	wire _w3700_ ;
	wire _w3701_ ;
	wire _w3702_ ;
	wire _w3703_ ;
	wire _w3704_ ;
	wire _w3705_ ;
	wire _w3706_ ;
	wire _w3707_ ;
	wire _w3708_ ;
	wire _w3709_ ;
	wire _w3710_ ;
	wire _w3711_ ;
	wire _w3712_ ;
	wire _w3713_ ;
	wire _w3714_ ;
	wire _w3715_ ;
	wire _w3716_ ;
	wire _w3717_ ;
	wire _w3718_ ;
	wire _w3719_ ;
	wire _w3720_ ;
	wire _w3721_ ;
	wire _w3722_ ;
	wire _w3723_ ;
	wire _w3724_ ;
	wire _w3725_ ;
	wire _w3726_ ;
	wire _w3727_ ;
	wire _w3728_ ;
	wire _w3729_ ;
	wire _w3730_ ;
	wire _w3731_ ;
	wire _w3732_ ;
	wire _w3733_ ;
	wire _w3734_ ;
	wire _w3735_ ;
	wire _w3736_ ;
	wire _w3737_ ;
	wire _w3738_ ;
	wire _w3739_ ;
	wire _w3740_ ;
	wire _w3741_ ;
	wire _w3742_ ;
	wire _w3743_ ;
	wire _w3744_ ;
	wire _w3745_ ;
	wire _w3746_ ;
	wire _w3747_ ;
	wire _w3748_ ;
	wire _w3749_ ;
	wire _w3750_ ;
	wire _w3751_ ;
	wire _w3752_ ;
	wire _w3753_ ;
	wire _w3754_ ;
	wire _w3755_ ;
	wire _w3756_ ;
	wire _w3757_ ;
	wire _w3758_ ;
	wire _w3759_ ;
	wire _w3760_ ;
	wire _w3761_ ;
	wire _w3762_ ;
	wire _w3763_ ;
	wire _w3764_ ;
	wire _w3765_ ;
	wire _w3766_ ;
	wire _w3767_ ;
	wire _w3768_ ;
	wire _w3769_ ;
	wire _w3770_ ;
	wire _w3771_ ;
	wire _w3772_ ;
	wire _w3773_ ;
	wire _w3774_ ;
	wire _w3775_ ;
	wire _w3776_ ;
	wire _w3777_ ;
	wire _w3778_ ;
	wire _w3779_ ;
	wire _w3780_ ;
	wire _w3781_ ;
	wire _w3782_ ;
	wire _w3783_ ;
	wire _w3784_ ;
	wire _w3785_ ;
	wire _w3786_ ;
	wire _w3787_ ;
	wire _w3788_ ;
	wire _w3789_ ;
	wire _w3790_ ;
	wire _w3791_ ;
	wire _w3792_ ;
	wire _w3793_ ;
	wire _w3794_ ;
	wire _w3795_ ;
	wire _w3796_ ;
	wire _w3797_ ;
	wire _w3798_ ;
	wire _w3799_ ;
	wire _w3800_ ;
	wire _w3801_ ;
	wire _w3802_ ;
	wire _w3803_ ;
	wire _w3804_ ;
	wire _w3805_ ;
	wire _w3806_ ;
	wire _w3807_ ;
	wire _w3808_ ;
	wire _w3809_ ;
	wire _w3810_ ;
	wire _w3811_ ;
	wire _w3812_ ;
	wire _w3813_ ;
	wire _w3814_ ;
	wire _w3815_ ;
	wire _w3816_ ;
	wire _w3817_ ;
	wire _w3818_ ;
	wire _w3819_ ;
	wire _w3820_ ;
	wire _w3821_ ;
	wire _w3822_ ;
	wire _w3823_ ;
	wire _w3824_ ;
	wire _w3825_ ;
	wire _w3826_ ;
	wire _w3827_ ;
	wire _w3828_ ;
	wire _w3829_ ;
	wire _w3830_ ;
	wire _w3831_ ;
	wire _w3832_ ;
	wire _w3833_ ;
	wire _w3834_ ;
	wire _w3835_ ;
	wire _w3836_ ;
	wire _w3837_ ;
	wire _w3838_ ;
	wire _w3839_ ;
	wire _w3840_ ;
	wire _w3841_ ;
	wire _w3842_ ;
	wire _w3843_ ;
	wire _w3844_ ;
	wire _w3845_ ;
	wire _w3846_ ;
	wire _w3847_ ;
	wire _w3848_ ;
	wire _w3849_ ;
	wire _w3850_ ;
	wire _w3851_ ;
	wire _w3852_ ;
	wire _w3853_ ;
	wire _w3854_ ;
	wire _w3855_ ;
	wire _w3856_ ;
	wire _w3857_ ;
	wire _w3858_ ;
	wire _w3859_ ;
	wire _w3860_ ;
	wire _w3861_ ;
	wire _w3862_ ;
	wire _w3863_ ;
	wire _w3864_ ;
	wire _w3865_ ;
	wire _w3866_ ;
	wire _w3867_ ;
	wire _w3868_ ;
	wire _w3869_ ;
	wire _w3870_ ;
	wire _w3871_ ;
	wire _w3872_ ;
	wire _w3873_ ;
	wire _w3874_ ;
	wire _w3875_ ;
	wire _w3876_ ;
	wire _w3877_ ;
	wire _w3878_ ;
	wire _w3879_ ;
	wire _w3880_ ;
	wire _w3881_ ;
	wire _w3882_ ;
	wire _w3883_ ;
	wire _w3884_ ;
	wire _w3885_ ;
	wire _w3886_ ;
	wire _w3887_ ;
	wire _w3888_ ;
	wire _w3889_ ;
	wire _w3890_ ;
	wire _w3891_ ;
	wire _w3892_ ;
	wire _w3893_ ;
	wire _w3894_ ;
	wire _w3895_ ;
	wire _w3896_ ;
	wire _w3897_ ;
	wire _w3898_ ;
	wire _w3899_ ;
	wire _w3900_ ;
	wire _w3901_ ;
	wire _w3902_ ;
	wire _w3903_ ;
	wire _w3904_ ;
	wire _w3905_ ;
	wire _w3906_ ;
	wire _w3907_ ;
	wire _w3908_ ;
	wire _w3909_ ;
	wire _w3910_ ;
	wire _w3911_ ;
	wire _w3912_ ;
	wire _w3913_ ;
	wire _w3914_ ;
	wire _w3915_ ;
	wire _w3916_ ;
	wire _w3917_ ;
	wire _w3918_ ;
	wire _w3919_ ;
	wire _w3920_ ;
	wire _w3921_ ;
	wire _w3922_ ;
	wire _w3923_ ;
	wire _w3924_ ;
	wire _w3925_ ;
	wire _w3926_ ;
	wire _w3927_ ;
	wire _w3928_ ;
	wire _w3929_ ;
	wire _w3930_ ;
	wire _w3931_ ;
	wire _w3932_ ;
	wire _w3933_ ;
	wire _w3934_ ;
	wire _w3935_ ;
	wire _w3936_ ;
	wire _w3937_ ;
	wire _w3938_ ;
	wire _w3939_ ;
	wire _w3940_ ;
	wire _w3941_ ;
	wire _w3942_ ;
	wire _w3943_ ;
	wire _w3944_ ;
	wire _w3945_ ;
	wire _w3946_ ;
	wire _w3947_ ;
	wire _w3948_ ;
	wire _w3949_ ;
	wire _w3950_ ;
	wire _w3951_ ;
	wire _w3952_ ;
	wire _w3953_ ;
	wire _w3954_ ;
	wire _w3955_ ;
	wire _w3956_ ;
	wire _w3957_ ;
	wire _w3958_ ;
	wire _w3959_ ;
	wire _w3960_ ;
	wire _w3961_ ;
	wire _w3962_ ;
	wire _w3963_ ;
	wire _w3964_ ;
	wire _w3965_ ;
	wire _w3966_ ;
	wire _w3967_ ;
	wire _w3968_ ;
	wire _w3969_ ;
	wire _w3970_ ;
	wire _w3971_ ;
	wire _w3972_ ;
	wire _w3973_ ;
	wire _w3974_ ;
	wire _w3975_ ;
	wire _w3976_ ;
	wire _w3977_ ;
	wire _w3978_ ;
	wire _w3979_ ;
	wire _w3980_ ;
	wire _w3981_ ;
	wire _w3982_ ;
	wire _w3983_ ;
	wire _w3984_ ;
	wire _w3985_ ;
	wire _w3986_ ;
	wire _w3987_ ;
	wire _w3988_ ;
	wire _w3989_ ;
	wire _w3990_ ;
	wire _w3991_ ;
	wire _w3992_ ;
	wire _w3993_ ;
	wire _w3994_ ;
	wire _w3995_ ;
	wire _w3996_ ;
	wire _w3997_ ;
	wire _w3998_ ;
	wire _w3999_ ;
	wire _w4000_ ;
	wire _w4001_ ;
	wire _w4002_ ;
	wire _w4003_ ;
	wire _w4004_ ;
	wire _w4005_ ;
	wire _w4006_ ;
	wire _w4007_ ;
	wire _w4008_ ;
	wire _w4009_ ;
	wire _w4010_ ;
	wire _w4011_ ;
	wire _w4012_ ;
	wire _w4013_ ;
	wire _w4014_ ;
	wire _w4015_ ;
	wire _w4016_ ;
	wire _w4017_ ;
	wire _w4018_ ;
	wire _w4019_ ;
	wire _w4020_ ;
	wire _w4021_ ;
	wire _w4022_ ;
	wire _w4023_ ;
	wire _w4024_ ;
	wire _w4025_ ;
	wire _w4026_ ;
	wire _w4027_ ;
	wire _w4028_ ;
	wire _w4029_ ;
	wire _w4030_ ;
	wire _w4031_ ;
	wire _w4032_ ;
	wire _w4033_ ;
	wire _w4034_ ;
	wire _w4035_ ;
	wire _w4036_ ;
	wire _w4037_ ;
	wire _w4038_ ;
	wire _w4039_ ;
	wire _w4040_ ;
	wire _w4041_ ;
	wire _w4042_ ;
	wire _w4043_ ;
	wire _w4044_ ;
	wire _w4045_ ;
	wire _w4046_ ;
	wire _w4047_ ;
	wire _w4048_ ;
	wire _w4049_ ;
	wire _w4050_ ;
	wire _w4051_ ;
	wire _w4052_ ;
	wire _w4053_ ;
	wire _w4054_ ;
	wire _w4055_ ;
	wire _w4056_ ;
	wire _w4057_ ;
	wire _w4058_ ;
	wire _w4059_ ;
	wire _w4060_ ;
	wire _w4061_ ;
	wire _w4062_ ;
	wire _w4063_ ;
	wire _w4064_ ;
	wire _w4065_ ;
	wire _w4066_ ;
	wire _w4067_ ;
	wire _w4068_ ;
	wire _w4069_ ;
	wire _w4070_ ;
	wire _w4071_ ;
	wire _w4072_ ;
	wire _w4073_ ;
	wire _w4074_ ;
	wire _w4075_ ;
	wire _w4076_ ;
	wire _w4077_ ;
	wire _w4078_ ;
	wire _w4079_ ;
	wire _w4080_ ;
	wire _w4081_ ;
	wire _w4082_ ;
	wire _w4083_ ;
	wire _w4084_ ;
	wire _w4085_ ;
	wire _w4086_ ;
	wire _w4087_ ;
	wire _w4088_ ;
	wire _w4089_ ;
	wire _w4090_ ;
	wire _w4091_ ;
	wire _w4092_ ;
	wire _w4093_ ;
	wire _w4094_ ;
	wire _w4095_ ;
	wire _w4096_ ;
	wire _w4097_ ;
	wire _w4098_ ;
	wire _w4099_ ;
	wire _w4100_ ;
	wire _w4101_ ;
	wire _w4102_ ;
	wire _w4103_ ;
	wire _w4104_ ;
	wire _w4105_ ;
	wire _w4106_ ;
	wire _w4107_ ;
	wire _w4108_ ;
	wire _w4109_ ;
	wire _w4110_ ;
	wire _w4111_ ;
	wire _w4112_ ;
	wire _w4113_ ;
	wire _w4114_ ;
	wire _w4115_ ;
	wire _w4116_ ;
	wire _w4117_ ;
	wire _w4118_ ;
	wire _w4119_ ;
	wire _w4120_ ;
	wire _w4121_ ;
	wire _w4122_ ;
	wire _w4123_ ;
	wire _w4124_ ;
	wire _w4125_ ;
	wire _w4126_ ;
	wire _w4127_ ;
	wire _w4128_ ;
	wire _w4129_ ;
	wire _w4130_ ;
	wire _w4131_ ;
	wire _w4132_ ;
	wire _w4133_ ;
	wire _w4134_ ;
	wire _w4135_ ;
	wire _w4136_ ;
	wire _w4137_ ;
	wire _w4138_ ;
	wire _w4139_ ;
	wire _w4140_ ;
	wire _w4141_ ;
	wire _w4142_ ;
	wire _w4143_ ;
	wire _w4144_ ;
	wire _w4145_ ;
	wire _w4146_ ;
	wire _w4147_ ;
	wire _w4148_ ;
	wire _w4149_ ;
	wire _w4150_ ;
	wire _w4151_ ;
	wire _w4152_ ;
	wire _w4153_ ;
	wire _w4154_ ;
	wire _w4155_ ;
	wire _w4156_ ;
	wire _w4157_ ;
	wire _w4158_ ;
	wire _w4159_ ;
	wire _w4160_ ;
	wire _w4161_ ;
	wire _w4162_ ;
	wire _w4163_ ;
	wire _w4164_ ;
	wire _w4165_ ;
	wire _w4166_ ;
	wire _w4167_ ;
	wire _w4168_ ;
	wire _w4169_ ;
	wire _w4170_ ;
	wire _w4171_ ;
	wire _w4172_ ;
	wire _w4173_ ;
	wire _w4174_ ;
	wire _w4175_ ;
	wire _w4176_ ;
	wire _w4177_ ;
	wire _w4178_ ;
	wire _w4179_ ;
	wire _w4180_ ;
	wire _w4181_ ;
	wire _w4182_ ;
	wire _w4183_ ;
	wire _w4184_ ;
	wire _w4185_ ;
	wire _w4186_ ;
	wire _w4187_ ;
	wire _w4188_ ;
	wire _w4189_ ;
	wire _w4190_ ;
	wire _w4191_ ;
	wire _w4192_ ;
	wire _w4193_ ;
	wire _w4194_ ;
	wire _w4195_ ;
	wire _w4196_ ;
	wire _w4197_ ;
	wire _w4198_ ;
	wire _w4199_ ;
	wire _w4200_ ;
	wire _w4201_ ;
	wire _w4202_ ;
	wire _w4203_ ;
	wire _w4204_ ;
	wire _w4205_ ;
	wire _w4206_ ;
	wire _w4207_ ;
	wire _w4208_ ;
	wire _w4209_ ;
	wire _w4210_ ;
	wire _w4211_ ;
	wire _w4212_ ;
	wire _w4213_ ;
	wire _w4214_ ;
	wire _w4215_ ;
	wire _w4216_ ;
	wire _w4217_ ;
	wire _w4218_ ;
	wire _w4219_ ;
	wire _w4220_ ;
	wire _w4221_ ;
	wire _w4222_ ;
	wire _w4223_ ;
	wire _w4224_ ;
	wire _w4225_ ;
	wire _w4226_ ;
	wire _w4227_ ;
	wire _w4228_ ;
	wire _w4229_ ;
	wire _w4230_ ;
	wire _w4231_ ;
	wire _w4232_ ;
	wire _w4233_ ;
	wire _w4234_ ;
	wire _w4235_ ;
	wire _w4236_ ;
	wire _w4237_ ;
	wire _w4238_ ;
	wire _w4239_ ;
	wire _w4240_ ;
	wire _w4241_ ;
	wire _w4242_ ;
	wire _w4243_ ;
	wire _w4244_ ;
	wire _w4245_ ;
	wire _w4246_ ;
	wire _w4247_ ;
	wire _w4248_ ;
	wire _w4249_ ;
	wire _w4250_ ;
	wire _w4251_ ;
	wire _w4252_ ;
	wire _w4253_ ;
	wire _w4254_ ;
	wire _w4255_ ;
	wire _w4256_ ;
	wire _w4257_ ;
	wire _w4258_ ;
	wire _w4259_ ;
	wire _w4260_ ;
	wire _w4261_ ;
	wire _w4262_ ;
	wire _w4263_ ;
	wire _w4264_ ;
	wire _w4265_ ;
	wire _w4266_ ;
	wire _w4267_ ;
	wire _w4268_ ;
	wire _w4269_ ;
	wire _w4270_ ;
	wire _w4271_ ;
	wire _w4272_ ;
	wire _w4273_ ;
	wire _w4274_ ;
	wire _w4275_ ;
	wire _w4276_ ;
	wire _w4277_ ;
	wire _w4278_ ;
	wire _w4279_ ;
	wire _w4280_ ;
	wire _w4281_ ;
	wire _w4282_ ;
	wire _w4283_ ;
	wire _w4284_ ;
	wire _w4285_ ;
	wire _w4286_ ;
	wire _w4287_ ;
	wire _w4288_ ;
	wire _w4289_ ;
	wire _w4290_ ;
	wire _w4291_ ;
	wire _w4292_ ;
	wire _w4293_ ;
	wire _w4294_ ;
	wire _w4295_ ;
	wire _w4296_ ;
	wire _w4297_ ;
	wire _w4298_ ;
	wire _w4299_ ;
	wire _w4300_ ;
	wire _w4301_ ;
	wire _w4302_ ;
	wire _w4303_ ;
	wire _w4304_ ;
	wire _w4305_ ;
	wire _w4306_ ;
	wire _w4307_ ;
	wire _w4308_ ;
	wire _w4309_ ;
	wire _w4310_ ;
	wire _w4311_ ;
	wire _w4312_ ;
	wire _w4313_ ;
	wire _w4314_ ;
	wire _w4315_ ;
	wire _w4316_ ;
	wire _w4317_ ;
	wire _w4318_ ;
	wire _w4319_ ;
	wire _w4320_ ;
	wire _w4321_ ;
	wire _w4322_ ;
	wire _w4323_ ;
	wire _w4324_ ;
	wire _w4325_ ;
	wire _w4326_ ;
	wire _w4327_ ;
	wire _w4328_ ;
	wire _w4329_ ;
	wire _w4330_ ;
	wire _w4331_ ;
	wire _w4332_ ;
	wire _w4333_ ;
	wire _w4334_ ;
	wire _w4335_ ;
	wire _w4336_ ;
	wire _w4337_ ;
	wire _w4338_ ;
	wire _w4339_ ;
	wire _w4340_ ;
	wire _w4341_ ;
	wire _w4342_ ;
	wire _w4343_ ;
	wire _w4344_ ;
	wire _w4345_ ;
	wire _w4346_ ;
	wire _w4347_ ;
	wire _w4348_ ;
	wire _w4349_ ;
	wire _w4350_ ;
	wire _w4351_ ;
	wire _w4352_ ;
	wire _w4353_ ;
	wire _w4354_ ;
	wire _w4355_ ;
	wire _w4356_ ;
	wire _w4357_ ;
	wire _w4358_ ;
	wire _w4359_ ;
	wire _w4360_ ;
	wire _w4361_ ;
	wire _w4362_ ;
	wire _w4363_ ;
	wire _w4364_ ;
	wire _w4365_ ;
	wire _w4366_ ;
	wire _w4367_ ;
	wire _w4368_ ;
	wire _w4369_ ;
	wire _w4370_ ;
	wire _w4371_ ;
	wire _w4372_ ;
	wire _w4373_ ;
	wire _w4374_ ;
	wire _w4375_ ;
	wire _w4376_ ;
	wire _w4377_ ;
	wire _w4378_ ;
	wire _w4379_ ;
	wire _w4380_ ;
	wire _w4381_ ;
	wire _w4382_ ;
	wire _w4383_ ;
	wire _w4384_ ;
	wire _w4385_ ;
	wire _w4386_ ;
	wire _w4387_ ;
	wire _w4388_ ;
	wire _w4389_ ;
	wire _w4390_ ;
	wire _w4391_ ;
	wire _w4392_ ;
	wire _w4393_ ;
	wire _w4394_ ;
	wire _w4395_ ;
	wire _w4396_ ;
	wire _w4397_ ;
	wire _w4398_ ;
	wire _w4399_ ;
	wire _w4400_ ;
	wire _w4401_ ;
	wire _w4402_ ;
	wire _w4403_ ;
	wire _w4404_ ;
	wire _w4405_ ;
	wire _w4406_ ;
	wire _w4407_ ;
	wire _w4408_ ;
	wire _w4409_ ;
	wire _w4410_ ;
	wire _w4411_ ;
	wire _w4412_ ;
	wire _w4413_ ;
	wire _w4414_ ;
	wire _w4415_ ;
	wire _w4416_ ;
	wire _w4417_ ;
	wire _w4418_ ;
	wire _w4419_ ;
	wire _w4420_ ;
	wire _w4421_ ;
	wire _w4422_ ;
	wire _w4423_ ;
	wire _w4424_ ;
	wire _w4425_ ;
	wire _w4426_ ;
	wire _w4427_ ;
	wire _w4428_ ;
	wire _w4429_ ;
	wire _w4430_ ;
	wire _w4431_ ;
	wire _w4432_ ;
	wire _w4433_ ;
	wire _w4434_ ;
	wire _w4435_ ;
	wire _w4436_ ;
	wire _w4437_ ;
	wire _w4438_ ;
	wire _w4439_ ;
	wire _w4440_ ;
	wire _w4441_ ;
	wire _w4442_ ;
	wire _w4443_ ;
	wire _w4444_ ;
	wire _w4445_ ;
	wire _w4446_ ;
	wire _w4447_ ;
	wire _w4448_ ;
	wire _w4449_ ;
	wire _w4450_ ;
	wire _w4451_ ;
	wire _w4452_ ;
	wire _w4453_ ;
	wire _w4454_ ;
	wire _w4455_ ;
	wire _w4456_ ;
	wire _w4457_ ;
	wire _w4458_ ;
	wire _w4459_ ;
	wire _w4460_ ;
	wire _w4461_ ;
	wire _w4462_ ;
	wire _w4463_ ;
	wire _w4464_ ;
	wire _w4465_ ;
	wire _w4466_ ;
	wire _w4467_ ;
	wire _w4468_ ;
	wire _w4469_ ;
	wire _w4470_ ;
	wire _w4471_ ;
	wire _w4472_ ;
	wire _w4473_ ;
	wire _w4474_ ;
	wire _w4475_ ;
	wire _w4476_ ;
	wire _w4477_ ;
	wire _w4478_ ;
	wire _w4479_ ;
	wire _w4480_ ;
	wire _w4481_ ;
	wire _w4482_ ;
	wire _w4483_ ;
	wire _w4484_ ;
	wire _w4485_ ;
	wire _w4486_ ;
	wire _w4487_ ;
	wire _w4488_ ;
	wire _w4489_ ;
	wire _w4490_ ;
	wire _w4491_ ;
	wire _w4492_ ;
	wire _w4493_ ;
	wire _w4494_ ;
	wire _w4495_ ;
	wire _w4496_ ;
	wire _w4497_ ;
	wire _w4498_ ;
	wire _w4499_ ;
	wire _w4500_ ;
	wire _w4501_ ;
	wire _w4502_ ;
	wire _w4503_ ;
	wire _w4504_ ;
	wire _w4505_ ;
	wire _w4506_ ;
	wire _w4507_ ;
	wire _w4508_ ;
	wire _w4509_ ;
	wire _w4510_ ;
	wire _w4511_ ;
	wire _w4512_ ;
	wire _w4513_ ;
	wire _w4514_ ;
	wire _w4515_ ;
	wire _w4516_ ;
	wire _w4517_ ;
	wire _w4518_ ;
	wire _w4519_ ;
	wire _w4520_ ;
	wire _w4521_ ;
	wire _w4522_ ;
	wire _w4523_ ;
	wire _w4524_ ;
	wire _w4525_ ;
	wire _w4526_ ;
	wire _w4527_ ;
	wire _w4528_ ;
	wire _w4529_ ;
	wire _w4530_ ;
	wire _w4531_ ;
	wire _w4532_ ;
	wire _w4533_ ;
	wire _w4534_ ;
	wire _w4535_ ;
	wire _w4536_ ;
	wire _w4537_ ;
	wire _w4538_ ;
	wire _w4539_ ;
	wire _w4540_ ;
	wire _w4541_ ;
	wire _w4542_ ;
	wire _w4543_ ;
	wire _w4544_ ;
	wire _w4545_ ;
	wire _w4546_ ;
	wire _w4547_ ;
	wire _w4548_ ;
	wire _w4549_ ;
	wire _w4550_ ;
	wire _w4551_ ;
	wire _w4552_ ;
	wire _w4553_ ;
	wire _w4554_ ;
	wire _w4555_ ;
	wire _w4556_ ;
	wire _w4557_ ;
	wire _w4558_ ;
	wire _w4559_ ;
	wire _w4560_ ;
	wire _w4561_ ;
	wire _w4562_ ;
	wire _w4563_ ;
	wire _w4564_ ;
	wire _w4565_ ;
	wire _w4566_ ;
	wire _w4567_ ;
	wire _w4568_ ;
	wire _w4569_ ;
	wire _w4570_ ;
	wire _w4571_ ;
	wire _w4572_ ;
	wire _w4573_ ;
	wire _w4574_ ;
	wire _w4575_ ;
	wire _w4576_ ;
	wire _w4577_ ;
	wire _w4578_ ;
	wire _w4579_ ;
	wire _w4580_ ;
	wire _w4581_ ;
	wire _w4582_ ;
	wire _w4583_ ;
	wire _w4584_ ;
	wire _w4585_ ;
	wire _w4586_ ;
	wire _w4587_ ;
	wire _w4588_ ;
	wire _w4589_ ;
	wire _w4590_ ;
	wire _w4591_ ;
	wire _w4592_ ;
	wire _w4593_ ;
	wire _w4594_ ;
	wire _w4595_ ;
	wire _w4596_ ;
	wire _w4597_ ;
	wire _w4598_ ;
	wire _w4599_ ;
	wire _w4600_ ;
	wire _w4601_ ;
	wire _w4602_ ;
	wire _w4603_ ;
	wire _w4604_ ;
	wire _w4605_ ;
	wire _w4606_ ;
	wire _w4607_ ;
	wire _w4608_ ;
	wire _w4609_ ;
	wire _w4610_ ;
	wire _w4611_ ;
	wire _w4612_ ;
	wire _w4613_ ;
	wire _w4614_ ;
	wire _w4615_ ;
	wire _w4616_ ;
	wire _w4617_ ;
	wire _w4618_ ;
	wire _w4619_ ;
	wire _w4620_ ;
	wire _w4621_ ;
	wire _w4622_ ;
	wire _w4623_ ;
	wire _w4624_ ;
	wire _w4625_ ;
	wire _w4626_ ;
	wire _w4627_ ;
	wire _w4628_ ;
	wire _w4629_ ;
	wire _w4630_ ;
	wire _w4631_ ;
	wire _w4632_ ;
	wire _w4633_ ;
	wire _w4634_ ;
	wire _w4635_ ;
	wire _w4636_ ;
	wire _w4637_ ;
	wire _w4638_ ;
	wire _w4639_ ;
	wire _w4640_ ;
	wire _w4641_ ;
	wire _w4642_ ;
	wire _w4643_ ;
	wire _w4644_ ;
	wire _w4645_ ;
	wire _w4646_ ;
	wire _w4647_ ;
	wire _w4648_ ;
	wire _w4649_ ;
	wire _w4650_ ;
	wire _w4651_ ;
	wire _w4652_ ;
	wire _w4653_ ;
	wire _w4654_ ;
	wire _w4655_ ;
	wire _w4656_ ;
	wire _w4657_ ;
	wire _w4658_ ;
	wire _w4659_ ;
	wire _w4660_ ;
	wire _w4661_ ;
	wire _w4662_ ;
	wire _w4663_ ;
	wire _w4664_ ;
	wire _w4665_ ;
	wire _w4666_ ;
	wire _w4667_ ;
	wire _w4668_ ;
	wire _w4669_ ;
	wire _w4670_ ;
	wire _w4671_ ;
	wire _w4672_ ;
	wire _w4673_ ;
	wire _w4674_ ;
	wire _w4675_ ;
	wire _w4676_ ;
	wire _w4677_ ;
	wire _w4678_ ;
	wire _w4679_ ;
	wire _w4680_ ;
	wire _w4681_ ;
	wire _w4682_ ;
	wire _w4683_ ;
	wire _w4684_ ;
	wire _w4685_ ;
	wire _w4686_ ;
	wire _w4687_ ;
	wire _w4688_ ;
	wire _w4689_ ;
	wire _w4690_ ;
	wire _w4691_ ;
	wire _w4692_ ;
	wire _w4693_ ;
	wire _w4694_ ;
	wire _w4695_ ;
	wire _w4696_ ;
	wire _w4697_ ;
	wire _w4698_ ;
	wire _w4699_ ;
	wire _w4700_ ;
	wire _w4701_ ;
	wire _w4702_ ;
	wire _w4703_ ;
	wire _w4704_ ;
	wire _w4705_ ;
	wire _w4706_ ;
	wire _w4707_ ;
	wire _w4708_ ;
	wire _w4709_ ;
	wire _w4710_ ;
	wire _w4711_ ;
	wire _w4712_ ;
	wire _w4713_ ;
	wire _w4714_ ;
	wire _w4715_ ;
	wire _w4716_ ;
	wire _w4717_ ;
	wire _w4718_ ;
	wire _w4719_ ;
	wire _w4720_ ;
	wire _w4721_ ;
	wire _w4722_ ;
	wire _w4723_ ;
	wire _w4724_ ;
	wire _w4725_ ;
	wire _w4726_ ;
	wire _w4727_ ;
	wire _w4728_ ;
	wire _w4729_ ;
	wire _w4730_ ;
	wire _w4731_ ;
	wire _w4732_ ;
	wire _w4733_ ;
	wire _w4734_ ;
	wire _w4735_ ;
	wire _w4736_ ;
	wire _w4737_ ;
	wire _w4738_ ;
	wire _w4739_ ;
	wire _w4740_ ;
	wire _w4741_ ;
	wire _w4742_ ;
	wire _w4743_ ;
	wire _w4744_ ;
	wire _w4745_ ;
	wire _w4746_ ;
	wire _w4747_ ;
	wire _w4748_ ;
	wire _w4749_ ;
	wire _w4750_ ;
	wire _w4751_ ;
	wire _w4752_ ;
	wire _w4753_ ;
	wire _w4754_ ;
	wire _w4755_ ;
	wire _w4756_ ;
	wire _w4757_ ;
	wire _w4758_ ;
	wire _w4759_ ;
	wire _w4760_ ;
	wire _w4761_ ;
	wire _w4762_ ;
	wire _w4763_ ;
	wire _w4764_ ;
	wire _w4765_ ;
	wire _w4766_ ;
	wire _w4767_ ;
	wire _w4768_ ;
	wire _w4769_ ;
	wire _w4770_ ;
	wire _w4771_ ;
	wire _w4772_ ;
	wire _w4773_ ;
	wire _w4774_ ;
	wire _w4775_ ;
	wire _w4776_ ;
	wire _w4777_ ;
	wire _w4778_ ;
	wire _w4779_ ;
	wire _w4780_ ;
	wire _w4781_ ;
	wire _w4782_ ;
	wire _w4783_ ;
	wire _w4784_ ;
	wire _w4785_ ;
	wire _w4786_ ;
	wire _w4787_ ;
	wire _w4788_ ;
	wire _w4789_ ;
	wire _w4790_ ;
	wire _w4791_ ;
	wire _w4792_ ;
	wire _w4793_ ;
	wire _w4794_ ;
	wire _w4795_ ;
	wire _w4796_ ;
	wire _w4797_ ;
	wire _w4798_ ;
	wire _w4799_ ;
	wire _w4800_ ;
	wire _w4801_ ;
	wire _w4802_ ;
	wire _w4803_ ;
	wire _w4804_ ;
	wire _w4805_ ;
	wire _w4806_ ;
	wire _w4807_ ;
	wire _w4808_ ;
	wire _w4809_ ;
	wire _w4810_ ;
	wire _w4811_ ;
	wire _w4812_ ;
	wire _w4813_ ;
	wire _w4814_ ;
	wire _w4815_ ;
	wire _w4816_ ;
	wire _w4817_ ;
	wire _w4818_ ;
	wire _w4819_ ;
	wire _w4820_ ;
	wire _w4821_ ;
	wire _w4822_ ;
	wire _w4823_ ;
	wire _w4824_ ;
	wire _w4825_ ;
	wire _w4826_ ;
	wire _w4827_ ;
	wire _w4828_ ;
	wire _w4829_ ;
	wire _w4830_ ;
	wire _w4831_ ;
	wire _w4832_ ;
	wire _w4833_ ;
	wire _w4834_ ;
	wire _w4835_ ;
	wire _w4836_ ;
	wire _w4837_ ;
	wire _w4838_ ;
	wire _w4839_ ;
	wire _w4840_ ;
	wire _w4841_ ;
	wire _w4842_ ;
	wire _w4843_ ;
	wire _w4844_ ;
	wire _w4845_ ;
	wire _w4846_ ;
	wire _w4847_ ;
	wire _w4848_ ;
	wire _w4849_ ;
	wire _w4850_ ;
	wire _w4851_ ;
	wire _w4852_ ;
	wire _w4853_ ;
	wire _w4854_ ;
	wire _w4855_ ;
	wire _w4856_ ;
	wire _w4857_ ;
	wire _w4858_ ;
	wire _w4859_ ;
	wire _w4860_ ;
	wire _w4861_ ;
	wire _w4862_ ;
	wire _w4863_ ;
	wire _w4864_ ;
	wire _w4865_ ;
	wire _w4866_ ;
	wire _w4867_ ;
	wire _w4868_ ;
	wire _w4869_ ;
	wire _w4870_ ;
	wire _w4871_ ;
	wire _w4872_ ;
	wire _w4873_ ;
	wire _w4874_ ;
	wire _w4875_ ;
	wire _w4876_ ;
	wire _w4877_ ;
	wire _w4878_ ;
	wire _w4879_ ;
	wire _w4880_ ;
	wire _w4881_ ;
	wire _w4882_ ;
	wire _w4883_ ;
	wire _w4884_ ;
	wire _w4885_ ;
	wire _w4886_ ;
	wire _w4887_ ;
	wire _w4888_ ;
	wire _w4889_ ;
	wire _w4890_ ;
	wire _w4891_ ;
	wire _w4892_ ;
	wire _w4893_ ;
	wire _w4894_ ;
	wire _w4895_ ;
	wire _w4896_ ;
	wire _w4897_ ;
	wire _w4898_ ;
	wire _w4899_ ;
	wire _w4900_ ;
	wire _w4901_ ;
	wire _w4902_ ;
	wire _w4903_ ;
	wire _w4904_ ;
	wire _w4905_ ;
	wire _w4906_ ;
	wire _w4907_ ;
	wire _w4908_ ;
	wire _w4909_ ;
	wire _w4910_ ;
	wire _w4911_ ;
	wire _w4912_ ;
	wire _w4913_ ;
	wire _w4914_ ;
	wire _w4915_ ;
	wire _w4916_ ;
	wire _w4917_ ;
	wire _w4918_ ;
	wire _w4919_ ;
	wire _w4920_ ;
	wire _w4921_ ;
	wire _w4922_ ;
	wire _w4923_ ;
	wire _w4924_ ;
	wire _w4925_ ;
	wire _w4926_ ;
	wire _w4927_ ;
	wire _w4928_ ;
	wire _w4929_ ;
	wire _w4930_ ;
	wire _w4931_ ;
	wire _w4932_ ;
	wire _w4933_ ;
	wire _w4934_ ;
	wire _w4935_ ;
	wire _w4936_ ;
	wire _w4937_ ;
	wire _w4938_ ;
	wire _w4939_ ;
	wire _w4940_ ;
	wire _w4941_ ;
	wire _w4942_ ;
	wire _w4943_ ;
	wire _w4944_ ;
	wire _w4945_ ;
	wire _w4946_ ;
	wire _w4947_ ;
	wire _w4948_ ;
	wire _w4949_ ;
	wire _w4950_ ;
	wire _w4951_ ;
	wire _w4952_ ;
	wire _w4953_ ;
	wire _w4954_ ;
	wire _w4955_ ;
	wire _w4956_ ;
	wire _w4957_ ;
	wire _w4958_ ;
	wire _w4959_ ;
	wire _w4960_ ;
	wire _w4961_ ;
	wire _w4962_ ;
	wire _w4963_ ;
	wire _w4964_ ;
	wire _w4965_ ;
	wire _w4966_ ;
	wire _w4967_ ;
	wire _w4968_ ;
	wire _w4969_ ;
	wire _w4970_ ;
	wire _w4971_ ;
	wire _w4972_ ;
	wire _w4973_ ;
	wire _w4974_ ;
	wire _w4975_ ;
	wire _w4976_ ;
	wire _w4977_ ;
	wire _w4978_ ;
	wire _w4979_ ;
	wire _w4980_ ;
	wire _w4981_ ;
	wire _w4982_ ;
	wire _w4983_ ;
	wire _w4984_ ;
	wire _w4985_ ;
	wire _w4986_ ;
	wire _w4987_ ;
	wire _w4988_ ;
	wire _w4989_ ;
	wire _w4990_ ;
	wire _w4991_ ;
	wire _w4992_ ;
	wire _w4993_ ;
	wire _w4994_ ;
	wire _w4995_ ;
	wire _w4996_ ;
	wire _w4997_ ;
	wire _w4998_ ;
	wire _w4999_ ;
	wire _w5000_ ;
	wire _w5001_ ;
	wire _w5002_ ;
	wire _w5003_ ;
	wire _w5004_ ;
	wire _w5005_ ;
	wire _w5006_ ;
	wire _w5007_ ;
	wire _w5008_ ;
	wire _w5009_ ;
	wire _w5010_ ;
	wire _w5011_ ;
	wire _w5012_ ;
	wire _w5013_ ;
	wire _w5014_ ;
	wire _w5015_ ;
	wire _w5016_ ;
	wire _w5017_ ;
	wire _w5018_ ;
	wire _w5019_ ;
	wire _w5020_ ;
	wire _w5021_ ;
	wire _w5022_ ;
	wire _w5023_ ;
	wire _w5024_ ;
	wire _w5025_ ;
	wire _w5026_ ;
	wire _w5027_ ;
	wire _w5028_ ;
	wire _w5029_ ;
	wire _w5030_ ;
	wire _w5031_ ;
	wire _w5032_ ;
	wire _w5033_ ;
	wire _w5034_ ;
	wire _w5035_ ;
	wire _w5036_ ;
	wire _w5037_ ;
	wire _w5038_ ;
	wire _w5039_ ;
	wire _w5040_ ;
	wire _w5041_ ;
	wire _w5042_ ;
	wire _w5043_ ;
	wire _w5044_ ;
	wire _w5045_ ;
	wire _w5046_ ;
	wire _w5047_ ;
	wire _w5048_ ;
	wire _w5049_ ;
	wire _w5050_ ;
	wire _w5051_ ;
	wire _w5052_ ;
	wire _w5053_ ;
	wire _w5054_ ;
	wire _w5055_ ;
	wire _w5056_ ;
	wire _w5057_ ;
	wire _w5058_ ;
	wire _w5059_ ;
	wire _w5060_ ;
	wire _w5061_ ;
	wire _w5062_ ;
	wire _w5063_ ;
	wire _w5064_ ;
	wire _w5065_ ;
	wire _w5066_ ;
	wire _w5067_ ;
	wire _w5068_ ;
	wire _w5069_ ;
	wire _w5070_ ;
	wire _w5071_ ;
	wire _w5072_ ;
	wire _w5073_ ;
	wire _w5074_ ;
	wire _w5075_ ;
	wire _w5076_ ;
	wire _w5077_ ;
	wire _w5078_ ;
	wire _w5079_ ;
	wire _w5080_ ;
	wire _w5081_ ;
	wire _w5082_ ;
	wire _w5083_ ;
	wire _w5084_ ;
	wire _w5085_ ;
	wire _w5086_ ;
	wire _w5087_ ;
	wire _w5088_ ;
	wire _w5089_ ;
	wire _w5090_ ;
	wire _w5091_ ;
	wire _w5092_ ;
	wire _w5093_ ;
	wire _w5094_ ;
	wire _w5095_ ;
	wire _w5096_ ;
	wire _w5097_ ;
	wire _w5098_ ;
	wire _w5099_ ;
	wire _w5100_ ;
	wire _w5101_ ;
	wire _w5102_ ;
	wire _w5103_ ;
	wire _w5104_ ;
	wire _w5105_ ;
	wire _w5106_ ;
	wire _w5107_ ;
	wire _w5108_ ;
	wire _w5109_ ;
	wire _w5110_ ;
	wire _w5111_ ;
	wire _w5112_ ;
	wire _w5113_ ;
	wire _w5114_ ;
	wire _w5115_ ;
	wire _w5116_ ;
	wire _w5117_ ;
	wire _w5118_ ;
	wire _w5119_ ;
	wire _w5120_ ;
	wire _w5121_ ;
	wire _w5122_ ;
	wire _w5123_ ;
	wire _w5124_ ;
	wire _w5125_ ;
	wire _w5126_ ;
	wire _w5127_ ;
	wire _w5128_ ;
	wire _w5129_ ;
	wire _w5130_ ;
	wire _w5131_ ;
	wire _w5132_ ;
	wire _w5133_ ;
	wire _w5134_ ;
	wire _w5135_ ;
	wire _w5136_ ;
	wire _w5137_ ;
	wire _w5138_ ;
	wire _w5139_ ;
	wire _w5140_ ;
	wire _w5141_ ;
	wire _w5142_ ;
	wire _w5143_ ;
	wire _w5144_ ;
	wire _w5145_ ;
	wire _w5146_ ;
	wire _w5147_ ;
	wire _w5148_ ;
	wire _w5149_ ;
	wire _w5150_ ;
	wire _w5151_ ;
	wire _w5152_ ;
	wire _w5153_ ;
	wire _w5154_ ;
	wire _w5155_ ;
	wire _w5156_ ;
	wire _w5157_ ;
	wire _w5158_ ;
	wire _w5159_ ;
	wire _w5160_ ;
	wire _w5161_ ;
	wire _w5162_ ;
	wire _w5163_ ;
	wire _w5164_ ;
	wire _w5165_ ;
	wire _w5166_ ;
	wire _w5167_ ;
	wire _w5168_ ;
	wire _w5169_ ;
	wire _w5170_ ;
	wire _w5171_ ;
	wire _w5172_ ;
	wire _w5173_ ;
	wire _w5174_ ;
	wire _w5175_ ;
	wire _w5176_ ;
	wire _w5177_ ;
	wire _w5178_ ;
	wire _w5179_ ;
	wire _w5180_ ;
	wire _w5181_ ;
	wire _w5182_ ;
	wire _w5183_ ;
	wire _w5184_ ;
	wire _w5185_ ;
	wire _w5186_ ;
	wire _w5187_ ;
	wire _w5188_ ;
	wire _w5189_ ;
	wire _w5190_ ;
	wire _w5191_ ;
	wire _w5192_ ;
	wire _w5193_ ;
	wire _w5194_ ;
	wire _w5195_ ;
	wire _w5196_ ;
	wire _w5197_ ;
	wire _w5198_ ;
	wire _w5199_ ;
	wire _w5200_ ;
	wire _w5201_ ;
	wire _w5202_ ;
	wire _w5203_ ;
	wire _w5204_ ;
	wire _w5205_ ;
	wire _w5206_ ;
	wire _w5207_ ;
	wire _w5208_ ;
	wire _w5209_ ;
	wire _w5210_ ;
	wire _w5211_ ;
	wire _w5212_ ;
	wire _w5213_ ;
	wire _w5214_ ;
	wire _w5215_ ;
	wire _w5216_ ;
	wire _w5217_ ;
	wire _w5218_ ;
	wire _w5219_ ;
	wire _w5220_ ;
	wire _w5221_ ;
	wire _w5222_ ;
	wire _w5223_ ;
	wire _w5224_ ;
	wire _w5225_ ;
	wire _w5226_ ;
	wire _w5227_ ;
	wire _w5228_ ;
	wire _w5229_ ;
	wire _w5230_ ;
	wire _w5231_ ;
	wire _w5232_ ;
	wire _w5233_ ;
	wire _w5234_ ;
	wire _w5235_ ;
	wire _w5236_ ;
	wire _w5237_ ;
	wire _w5238_ ;
	wire _w5239_ ;
	wire _w5240_ ;
	wire _w5241_ ;
	wire _w5242_ ;
	wire _w5243_ ;
	wire _w5244_ ;
	wire _w5245_ ;
	wire _w5246_ ;
	wire _w5247_ ;
	wire _w5248_ ;
	wire _w5249_ ;
	wire _w5250_ ;
	wire _w5251_ ;
	wire _w5252_ ;
	wire _w5253_ ;
	wire _w5254_ ;
	wire _w5255_ ;
	wire _w5256_ ;
	wire _w5257_ ;
	wire _w5258_ ;
	wire _w5259_ ;
	wire _w5260_ ;
	wire _w5261_ ;
	wire _w5262_ ;
	wire _w5263_ ;
	wire _w5264_ ;
	wire _w5265_ ;
	wire _w5266_ ;
	wire _w5267_ ;
	wire _w5268_ ;
	wire _w5269_ ;
	wire _w5270_ ;
	wire _w5271_ ;
	wire _w5272_ ;
	wire _w5273_ ;
	wire _w5274_ ;
	wire _w5275_ ;
	wire _w5276_ ;
	wire _w5277_ ;
	wire _w5278_ ;
	wire _w5279_ ;
	wire _w5280_ ;
	wire _w5281_ ;
	wire _w5282_ ;
	wire _w5283_ ;
	wire _w5284_ ;
	wire _w5285_ ;
	wire _w5286_ ;
	wire _w5287_ ;
	wire _w5288_ ;
	wire _w5289_ ;
	wire _w5290_ ;
	wire _w5291_ ;
	wire _w5292_ ;
	wire _w5293_ ;
	wire _w5294_ ;
	wire _w5295_ ;
	wire _w5296_ ;
	wire _w5297_ ;
	wire _w5298_ ;
	wire _w5299_ ;
	wire _w5300_ ;
	wire _w5301_ ;
	wire _w5302_ ;
	wire _w5304_ ;
	wire _w5305_ ;
	wire _w5306_ ;
	wire _w5307_ ;
	wire _w5308_ ;
	wire _w5309_ ;
	wire _w5310_ ;
	wire _w5311_ ;
	wire _w5312_ ;
	wire _w5313_ ;
	wire _w5314_ ;
	wire _w5315_ ;
	wire _w5316_ ;
	wire _w5317_ ;
	wire _w5318_ ;
	wire _w5319_ ;
	wire _w5320_ ;
	wire _w5321_ ;
	wire _w5322_ ;
	wire _w5323_ ;
	wire _w5324_ ;
	wire _w5325_ ;
	wire _w5326_ ;
	wire _w5327_ ;
	wire _w5328_ ;
	wire _w5329_ ;
	wire _w5330_ ;
	wire _w5331_ ;
	wire _w5332_ ;
	wire _w5333_ ;
	wire _w5334_ ;
	wire _w5335_ ;
	wire _w5336_ ;
	wire _w5337_ ;
	wire _w5338_ ;
	wire _w5339_ ;
	wire _w5340_ ;
	wire _w5341_ ;
	wire _w5342_ ;
	wire _w5343_ ;
	wire _w5344_ ;
	wire _w5345_ ;
	wire _w5346_ ;
	wire _w5347_ ;
	wire _w5348_ ;
	wire _w5349_ ;
	wire _w5350_ ;
	wire _w5351_ ;
	wire _w5352_ ;
	wire _w5353_ ;
	wire _w5354_ ;
	wire _w5355_ ;
	wire _w5356_ ;
	wire _w5357_ ;
	wire _w5358_ ;
	wire _w5359_ ;
	wire _w5360_ ;
	wire _w5361_ ;
	wire _w5362_ ;
	wire _w5363_ ;
	wire _w5364_ ;
	wire _w5365_ ;
	wire _w5366_ ;
	wire _w5367_ ;
	wire _w5368_ ;
	wire _w5369_ ;
	wire _w5370_ ;
	wire _w5371_ ;
	wire _w5372_ ;
	wire _w5373_ ;
	wire _w5374_ ;
	wire _w5375_ ;
	wire _w5376_ ;
	wire _w5377_ ;
	wire _w5378_ ;
	wire _w5379_ ;
	wire _w5380_ ;
	wire _w5381_ ;
	wire _w5382_ ;
	wire _w5383_ ;
	wire _w5384_ ;
	wire _w5385_ ;
	wire _w5386_ ;
	wire _w5387_ ;
	wire _w5388_ ;
	wire _w5389_ ;
	wire _w5390_ ;
	wire _w5391_ ;
	wire _w5392_ ;
	wire _w5393_ ;
	wire _w5394_ ;
	wire _w5395_ ;
	wire _w5396_ ;
	wire _w5397_ ;
	wire _w5398_ ;
	wire _w5399_ ;
	wire _w5400_ ;
	wire _w5401_ ;
	wire _w5402_ ;
	wire _w5403_ ;
	wire _w5404_ ;
	wire _w5405_ ;
	wire _w5406_ ;
	wire _w5407_ ;
	wire _w5408_ ;
	wire _w5409_ ;
	wire _w5410_ ;
	wire _w5411_ ;
	wire _w5412_ ;
	wire _w5413_ ;
	wire _w5414_ ;
	wire _w5415_ ;
	wire _w5416_ ;
	wire _w5417_ ;
	wire _w5418_ ;
	wire _w5419_ ;
	wire _w5420_ ;
	wire _w5421_ ;
	wire _w5422_ ;
	wire _w5423_ ;
	wire _w5424_ ;
	wire _w5425_ ;
	wire _w5426_ ;
	wire _w5427_ ;
	wire _w5428_ ;
	wire _w5429_ ;
	wire _w5430_ ;
	wire _w5431_ ;
	wire _w5432_ ;
	wire _w5433_ ;
	wire _w5434_ ;
	wire _w5435_ ;
	wire _w5436_ ;
	wire _w5437_ ;
	wire _w5438_ ;
	wire _w5439_ ;
	wire _w5440_ ;
	wire _w5441_ ;
	wire _w5442_ ;
	wire _w5443_ ;
	wire _w5444_ ;
	wire _w5445_ ;
	wire _w5446_ ;
	wire _w5447_ ;
	wire _w5448_ ;
	wire _w5449_ ;
	wire _w5450_ ;
	wire _w5451_ ;
	wire _w5452_ ;
	wire _w5453_ ;
	wire _w5454_ ;
	wire _w5455_ ;
	wire _w5456_ ;
	wire _w5457_ ;
	wire _w5458_ ;
	wire _w5459_ ;
	wire _w5460_ ;
	wire _w5461_ ;
	wire _w5462_ ;
	wire _w5463_ ;
	wire _w5464_ ;
	wire _w5465_ ;
	wire _w5466_ ;
	wire _w5467_ ;
	wire _w5468_ ;
	wire _w5469_ ;
	wire _w5470_ ;
	wire _w5471_ ;
	wire _w5472_ ;
	wire _w5473_ ;
	wire _w5474_ ;
	wire _w5475_ ;
	wire _w5476_ ;
	wire _w5477_ ;
	wire _w5478_ ;
	wire _w5479_ ;
	wire _w5480_ ;
	wire _w5481_ ;
	wire _w5482_ ;
	wire _w5483_ ;
	wire _w5484_ ;
	wire _w5485_ ;
	wire _w5486_ ;
	wire _w5487_ ;
	wire _w5488_ ;
	wire _w5489_ ;
	wire _w5490_ ;
	wire _w5491_ ;
	wire _w5492_ ;
	wire _w5493_ ;
	wire _w5494_ ;
	wire _w5495_ ;
	wire _w5496_ ;
	wire _w5497_ ;
	wire _w5498_ ;
	wire _w5499_ ;
	wire _w5500_ ;
	wire _w5501_ ;
	wire _w5502_ ;
	wire _w5503_ ;
	wire _w5504_ ;
	wire _w5505_ ;
	wire _w5506_ ;
	wire _w5507_ ;
	wire _w5508_ ;
	wire _w5509_ ;
	wire _w5510_ ;
	wire _w5511_ ;
	wire _w5512_ ;
	wire _w5513_ ;
	wire _w5514_ ;
	wire _w5515_ ;
	wire _w5516_ ;
	wire _w5517_ ;
	wire _w5518_ ;
	wire _w5519_ ;
	wire _w5520_ ;
	wire _w5521_ ;
	wire _w5522_ ;
	wire _w5523_ ;
	wire _w5524_ ;
	wire _w5525_ ;
	wire _w5526_ ;
	wire _w5527_ ;
	wire _w5528_ ;
	wire _w5529_ ;
	wire _w5530_ ;
	wire _w5531_ ;
	wire _w5532_ ;
	wire _w5533_ ;
	wire _w5534_ ;
	wire _w5535_ ;
	wire _w5536_ ;
	wire _w5537_ ;
	wire _w5538_ ;
	wire _w5539_ ;
	wire _w5540_ ;
	wire _w5541_ ;
	wire _w5542_ ;
	wire _w5543_ ;
	wire _w5544_ ;
	wire _w5545_ ;
	wire _w5546_ ;
	wire _w5547_ ;
	wire _w5548_ ;
	wire _w5549_ ;
	LUT1 #(
		.INIT('h1)
	) name0 (
		\P1_state_reg[0]/NET0131 ,
		_w216_
	);
	LUT4 #(
		.INIT('h0001)
	) name1 (
		\P2_reg3_reg[3]/NET0131 ,
		\P2_reg3_reg[4]/NET0131 ,
		\P2_reg3_reg[5]/NET0131 ,
		\P2_reg3_reg[6]/NET0131 ,
		_w464_
	);
	LUT4 #(
		.INIT('h0100)
	) name2 (
		\P2_reg3_reg[7]/NET0131 ,
		\P2_reg3_reg[8]/NET0131 ,
		\P2_reg3_reg[9]/NET0131 ,
		_w464_,
		_w465_
	);
	LUT3 #(
		.INIT('h10)
	) name3 (
		\P2_reg3_reg[10]/NET0131 ,
		\P2_reg3_reg[11]/NET0131 ,
		_w465_,
		_w466_
	);
	LUT4 #(
		.INIT('h0100)
	) name4 (
		\P2_reg3_reg[10]/NET0131 ,
		\P2_reg3_reg[11]/NET0131 ,
		\P2_reg3_reg[12]/NET0131 ,
		_w465_,
		_w467_
	);
	LUT4 #(
		.INIT('h0100)
	) name5 (
		\P2_reg3_reg[13]/NET0131 ,
		\P2_reg3_reg[14]/NET0131 ,
		\P2_reg3_reg[15]/NET0131 ,
		_w467_,
		_w468_
	);
	LUT4 #(
		.INIT('h0001)
	) name6 (
		\P2_reg3_reg[13]/NET0131 ,
		\P2_reg3_reg[14]/NET0131 ,
		\P2_reg3_reg[15]/NET0131 ,
		\P2_reg3_reg[16]/NET0131 ,
		_w469_
	);
	LUT2 #(
		.INIT('h8)
	) name7 (
		_w467_,
		_w469_,
		_w470_
	);
	LUT3 #(
		.INIT('h0d)
	) name8 (
		\P2_reg3_reg[16]/NET0131 ,
		_w468_,
		_w470_,
		_w471_
	);
	LUT4 #(
		.INIT('h0001)
	) name9 (
		\P2_IR_reg[0]/NET0131 ,
		\P2_IR_reg[1]/NET0131 ,
		\P2_IR_reg[2]/NET0131 ,
		\P2_IR_reg[3]/NET0131 ,
		_w472_
	);
	LUT3 #(
		.INIT('h01)
	) name10 (
		\P2_IR_reg[5]/NET0131 ,
		\P2_IR_reg[6]/NET0131 ,
		\P2_IR_reg[7]/NET0131 ,
		_w473_
	);
	LUT3 #(
		.INIT('h40)
	) name11 (
		\P2_IR_reg[4]/NET0131 ,
		_w472_,
		_w473_,
		_w474_
	);
	LUT3 #(
		.INIT('h01)
	) name12 (
		\P2_IR_reg[10]/NET0131 ,
		\P2_IR_reg[8]/NET0131 ,
		\P2_IR_reg[9]/NET0131 ,
		_w475_
	);
	LUT4 #(
		.INIT('h4000)
	) name13 (
		\P2_IR_reg[4]/NET0131 ,
		_w472_,
		_w473_,
		_w475_,
		_w476_
	);
	LUT2 #(
		.INIT('h1)
	) name14 (
		\P2_IR_reg[11]/NET0131 ,
		\P2_IR_reg[12]/NET0131 ,
		_w477_
	);
	LUT3 #(
		.INIT('h01)
	) name15 (
		\P2_IR_reg[11]/NET0131 ,
		\P2_IR_reg[12]/NET0131 ,
		\P2_IR_reg[13]/NET0131 ,
		_w478_
	);
	LUT3 #(
		.INIT('h2a)
	) name16 (
		\P2_IR_reg[31]/NET0131 ,
		_w476_,
		_w478_,
		_w479_
	);
	LUT4 #(
		.INIT('h0001)
	) name17 (
		\P2_IR_reg[14]/NET0131 ,
		\P2_IR_reg[15]/NET0131 ,
		\P2_IR_reg[16]/NET0131 ,
		\P2_IR_reg[17]/NET0131 ,
		_w480_
	);
	LUT4 #(
		.INIT('h0001)
	) name18 (
		\P2_IR_reg[19]/NET0131 ,
		\P2_IR_reg[20]/NET0131 ,
		\P2_IR_reg[21]/NET0131 ,
		\P2_IR_reg[22]/NET0131 ,
		_w481_
	);
	LUT4 #(
		.INIT('h1000)
	) name19 (
		\P2_IR_reg[18]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		_w480_,
		_w481_,
		_w482_
	);
	LUT2 #(
		.INIT('h1)
	) name20 (
		\P2_IR_reg[24]/NET0131 ,
		\P2_IR_reg[25]/NET0131 ,
		_w483_
	);
	LUT2 #(
		.INIT('h1)
	) name21 (
		\P2_IR_reg[27]/NET0131 ,
		\P2_IR_reg[28]/NET0131 ,
		_w484_
	);
	LUT3 #(
		.INIT('h01)
	) name22 (
		\P2_IR_reg[27]/NET0131 ,
		\P2_IR_reg[28]/NET0131 ,
		\P2_IR_reg[29]/NET0131 ,
		_w485_
	);
	LUT4 #(
		.INIT('h0001)
	) name23 (
		\P2_IR_reg[26]/NET0131 ,
		\P2_IR_reg[27]/NET0131 ,
		\P2_IR_reg[28]/NET0131 ,
		\P2_IR_reg[29]/NET0131 ,
		_w486_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name24 (
		\P2_IR_reg[31]/NET0131 ,
		_w482_,
		_w483_,
		_w486_,
		_w487_
	);
	LUT3 #(
		.INIT('h56)
	) name25 (
		\P2_IR_reg[30]/NET0131 ,
		_w479_,
		_w487_,
		_w488_
	);
	LUT3 #(
		.INIT('h2a)
	) name26 (
		\P2_IR_reg[31]/NET0131 ,
		_w476_,
		_w477_,
		_w489_
	);
	LUT4 #(
		.INIT('h1000)
	) name27 (
		\P2_IR_reg[13]/NET0131 ,
		\P2_IR_reg[18]/NET0131 ,
		_w480_,
		_w481_,
		_w490_
	);
	LUT4 #(
		.INIT('h0001)
	) name28 (
		\P2_IR_reg[23]/NET0131 ,
		\P2_IR_reg[24]/NET0131 ,
		\P2_IR_reg[25]/NET0131 ,
		\P2_IR_reg[26]/NET0131 ,
		_w491_
	);
	LUT2 #(
		.INIT('h8)
	) name29 (
		_w484_,
		_w491_,
		_w492_
	);
	LUT3 #(
		.INIT('h2a)
	) name30 (
		\P2_IR_reg[31]/NET0131 ,
		_w490_,
		_w492_,
		_w493_
	);
	LUT3 #(
		.INIT('h56)
	) name31 (
		\P2_IR_reg[29]/NET0131 ,
		_w489_,
		_w493_,
		_w494_
	);
	LUT2 #(
		.INIT('h8)
	) name32 (
		_w488_,
		_w494_,
		_w495_
	);
	LUT3 #(
		.INIT('h20)
	) name33 (
		\P2_reg1_reg[16]/NET0131 ,
		_w488_,
		_w494_,
		_w496_
	);
	LUT4 #(
		.INIT('hff35)
	) name34 (
		\P2_reg0_reg[16]/NET0131 ,
		\P2_reg2_reg[16]/NET0131 ,
		_w488_,
		_w494_,
		_w497_
	);
	LUT4 #(
		.INIT('h4500)
	) name35 (
		_w496_,
		_w471_,
		_w495_,
		_w497_,
		_w498_
	);
	LUT4 #(
		.INIT('hbaff)
	) name36 (
		_w496_,
		_w471_,
		_w495_,
		_w497_,
		_w499_
	);
	LUT4 #(
		.INIT('h0001)
	) name37 (
		\P1_IR_reg[0]/NET0131 ,
		\P1_IR_reg[1]/NET0131 ,
		\P1_IR_reg[2]/NET0131 ,
		\P1_IR_reg[3]/NET0131 ,
		_w500_
	);
	LUT2 #(
		.INIT('h1)
	) name38 (
		\P1_IR_reg[6]/NET0131 ,
		\P1_IR_reg[7]/NET0131 ,
		_w501_
	);
	LUT4 #(
		.INIT('h0001)
	) name39 (
		\P1_IR_reg[6]/NET0131 ,
		\P1_IR_reg[7]/NET0131 ,
		\P1_IR_reg[8]/NET0131 ,
		\P1_IR_reg[9]/NET0131 ,
		_w502_
	);
	LUT4 #(
		.INIT('h1000)
	) name40 (
		\P1_IR_reg[4]/NET0131 ,
		\P1_IR_reg[5]/NET0131 ,
		_w500_,
		_w502_,
		_w503_
	);
	LUT4 #(
		.INIT('h0001)
	) name41 (
		\P1_IR_reg[10]/NET0131 ,
		\P1_IR_reg[11]/NET0131 ,
		\P1_IR_reg[12]/NET0131 ,
		\P1_IR_reg[13]/NET0131 ,
		_w504_
	);
	LUT4 #(
		.INIT('h0001)
	) name42 (
		\P1_IR_reg[16]/NET0131 ,
		\P1_IR_reg[17]/NET0131 ,
		\P1_IR_reg[20]/NET0131 ,
		\P1_IR_reg[21]/NET0131 ,
		_w505_
	);
	LUT2 #(
		.INIT('h1)
	) name43 (
		\P1_IR_reg[18]/NET0131 ,
		\P1_IR_reg[19]/NET0131 ,
		_w506_
	);
	LUT4 #(
		.INIT('h0001)
	) name44 (
		\P1_IR_reg[14]/NET0131 ,
		\P1_IR_reg[15]/NET0131 ,
		\P1_IR_reg[18]/NET0131 ,
		\P1_IR_reg[19]/NET0131 ,
		_w507_
	);
	LUT2 #(
		.INIT('h8)
	) name45 (
		_w505_,
		_w507_,
		_w508_
	);
	LUT4 #(
		.INIT('h4000)
	) name46 (
		\P1_IR_reg[22]/NET0131 ,
		_w503_,
		_w504_,
		_w508_,
		_w509_
	);
	LUT3 #(
		.INIT('ha6)
	) name47 (
		\P1_IR_reg[23]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		_w509_,
		_w510_
	);
	LUT4 #(
		.INIT('h5090)
	) name48 (
		\P1_IR_reg[23]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w509_,
		_w511_
	);
	LUT2 #(
		.INIT('h2)
	) name49 (
		\P1_reg2_reg[29]/NET0131 ,
		_w511_,
		_w512_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name50 (
		\P1_IR_reg[31]/NET0131 ,
		_w503_,
		_w504_,
		_w508_,
		_w513_
	);
	LUT3 #(
		.INIT('h01)
	) name51 (
		\P1_IR_reg[22]/NET0131 ,
		\P1_IR_reg[23]/NET0131 ,
		\P1_IR_reg[24]/NET0131 ,
		_w514_
	);
	LUT4 #(
		.INIT('h0001)
	) name52 (
		\P1_IR_reg[22]/NET0131 ,
		\P1_IR_reg[23]/NET0131 ,
		\P1_IR_reg[24]/NET0131 ,
		\P1_IR_reg[25]/NET0131 ,
		_w515_
	);
	LUT2 #(
		.INIT('h2)
	) name53 (
		\P1_IR_reg[31]/NET0131 ,
		_w515_,
		_w516_
	);
	LUT3 #(
		.INIT('h56)
	) name54 (
		\P1_IR_reg[26]/NET0131 ,
		_w513_,
		_w516_,
		_w517_
	);
	LUT3 #(
		.INIT('he0)
	) name55 (
		\P1_IR_reg[22]/NET0131 ,
		\P1_IR_reg[23]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		_w518_
	);
	LUT3 #(
		.INIT('h56)
	) name56 (
		\P1_IR_reg[24]/NET0131 ,
		_w513_,
		_w518_,
		_w519_
	);
	LUT3 #(
		.INIT('h80)
	) name57 (
		_w505_,
		_w507_,
		_w514_,
		_w520_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name58 (
		\P1_IR_reg[31]/NET0131 ,
		_w503_,
		_w504_,
		_w520_,
		_w521_
	);
	LUT2 #(
		.INIT('h6)
	) name59 (
		\P1_IR_reg[25]/NET0131 ,
		_w521_,
		_w522_
	);
	LUT3 #(
		.INIT('h80)
	) name60 (
		_w519_,
		_w522_,
		_w517_,
		_w523_
	);
	LUT4 #(
		.INIT('h4000)
	) name61 (
		_w510_,
		_w519_,
		_w522_,
		_w517_,
		_w524_
	);
	LUT2 #(
		.INIT('h8)
	) name62 (
		\P1_reg2_reg[29]/NET0131 ,
		_w524_,
		_w525_
	);
	LUT4 #(
		.INIT('h1555)
	) name63 (
		_w510_,
		_w519_,
		_w522_,
		_w517_,
		_w526_
	);
	LUT4 #(
		.INIT('h8882)
	) name64 (
		\P1_B_reg/NET0131 ,
		\P1_IR_reg[24]/NET0131 ,
		_w513_,
		_w518_,
		_w527_
	);
	LUT4 #(
		.INIT('hb0a0)
	) name65 (
		\P1_d_reg[0]/NET0131 ,
		_w522_,
		_w517_,
		_w527_,
		_w528_
	);
	LUT3 #(
		.INIT('h41)
	) name66 (
		\P1_B_reg/NET0131 ,
		\P1_IR_reg[25]/NET0131 ,
		_w521_,
		_w529_
	);
	LUT3 #(
		.INIT('ha2)
	) name67 (
		_w519_,
		_w517_,
		_w529_,
		_w530_
	);
	LUT2 #(
		.INIT('he)
	) name68 (
		_w528_,
		_w530_,
		_w531_
	);
	LUT4 #(
		.INIT('h6669)
	) name69 (
		\P1_B_reg/NET0131 ,
		\P1_IR_reg[24]/NET0131 ,
		_w513_,
		_w518_,
		_w532_
	);
	LUT4 #(
		.INIT('hacbc)
	) name70 (
		\P1_d_reg[1]/NET0131 ,
		_w522_,
		_w517_,
		_w532_,
		_w533_
	);
	LUT3 #(
		.INIT('h10)
	) name71 (
		_w528_,
		_w530_,
		_w533_,
		_w534_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name72 (
		\P1_reg2_reg[29]/NET0131 ,
		_w528_,
		_w530_,
		_w533_,
		_w535_
	);
	LUT4 #(
		.INIT('he0f0)
	) name73 (
		\P1_IR_reg[26]/NET0131 ,
		\P1_IR_reg[27]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		_w515_,
		_w536_
	);
	LUT3 #(
		.INIT('h56)
	) name74 (
		\P1_IR_reg[28]/NET0131 ,
		_w513_,
		_w536_,
		_w537_
	);
	LUT4 #(
		.INIT('h0001)
	) name75 (
		\P1_IR_reg[23]/NET0131 ,
		\P1_IR_reg[24]/NET0131 ,
		\P1_IR_reg[25]/NET0131 ,
		\P1_IR_reg[26]/NET0131 ,
		_w538_
	);
	LUT2 #(
		.INIT('h2)
	) name76 (
		\P1_IR_reg[31]/NET0131 ,
		_w538_,
		_w539_
	);
	LUT4 #(
		.INIT('h55a6)
	) name77 (
		\P1_IR_reg[27]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		_w509_,
		_w539_,
		_w540_
	);
	LUT2 #(
		.INIT('h1)
	) name78 (
		_w537_,
		_w540_,
		_w541_
	);
	LUT4 #(
		.INIT('hfe5e)
	) name79 (
		\P1_addr_reg[19]/NET0131 ,
		\P1_rd_reg/NET0131 ,
		\P2_addr_reg[19]/NET0131 ,
		\P2_rd_reg/NET0131 ,
		_w542_
	);
	LUT2 #(
		.INIT('h8)
	) name80 (
		\P2_datao_reg[29]/NET0131 ,
		_w542_,
		_w543_
	);
	LUT2 #(
		.INIT('h8)
	) name81 (
		\P2_datao_reg[29]/NET0131 ,
		\si[29]_pad ,
		_w544_
	);
	LUT2 #(
		.INIT('h6)
	) name82 (
		\P2_datao_reg[29]/NET0131 ,
		\si[29]_pad ,
		_w545_
	);
	LUT2 #(
		.INIT('h1)
	) name83 (
		\P2_datao_reg[28]/NET0131 ,
		\si[28]_pad ,
		_w546_
	);
	LUT4 #(
		.INIT('h135f)
	) name84 (
		\P2_datao_reg[27]/NET0131 ,
		\P2_datao_reg[28]/NET0131 ,
		\si[27]_pad ,
		\si[28]_pad ,
		_w547_
	);
	LUT2 #(
		.INIT('h1)
	) name85 (
		\P2_datao_reg[27]/NET0131 ,
		\si[27]_pad ,
		_w548_
	);
	LUT2 #(
		.INIT('h1)
	) name86 (
		\P2_datao_reg[26]/NET0131 ,
		\si[26]_pad ,
		_w549_
	);
	LUT4 #(
		.INIT('hec80)
	) name87 (
		\P2_datao_reg[25]/NET0131 ,
		\P2_datao_reg[26]/NET0131 ,
		\si[25]_pad ,
		\si[26]_pad ,
		_w550_
	);
	LUT4 #(
		.INIT('hfac8)
	) name88 (
		\P2_datao_reg[25]/NET0131 ,
		\P2_datao_reg[26]/NET0131 ,
		\si[25]_pad ,
		\si[26]_pad ,
		_w551_
	);
	LUT2 #(
		.INIT('h1)
	) name89 (
		\P2_datao_reg[24]/NET0131 ,
		\si[24]_pad ,
		_w552_
	);
	LUT4 #(
		.INIT('hfac8)
	) name90 (
		\P2_datao_reg[23]/NET0131 ,
		\P2_datao_reg[24]/NET0131 ,
		\si[23]_pad ,
		\si[24]_pad ,
		_w553_
	);
	LUT4 #(
		.INIT('hec80)
	) name91 (
		\P2_datao_reg[21]/NET0131 ,
		\P2_datao_reg[22]/NET0131 ,
		\si[21]_pad ,
		\si[22]_pad ,
		_w554_
	);
	LUT4 #(
		.INIT('hec80)
	) name92 (
		\P2_datao_reg[23]/NET0131 ,
		\P2_datao_reg[24]/NET0131 ,
		\si[23]_pad ,
		\si[24]_pad ,
		_w555_
	);
	LUT3 #(
		.INIT('h07)
	) name93 (
		_w553_,
		_w554_,
		_w555_,
		_w556_
	);
	LUT4 #(
		.INIT('haa80)
	) name94 (
		_w551_,
		_w553_,
		_w554_,
		_w555_,
		_w557_
	);
	LUT4 #(
		.INIT('h888a)
	) name95 (
		_w547_,
		_w548_,
		_w550_,
		_w557_,
		_w558_
	);
	LUT2 #(
		.INIT('h1)
	) name96 (
		_w546_,
		_w558_,
		_w559_
	);
	LUT2 #(
		.INIT('h8)
	) name97 (
		\P2_datao_reg[4]/NET0131 ,
		\si[4]_pad ,
		_w560_
	);
	LUT2 #(
		.INIT('h8)
	) name98 (
		\P2_datao_reg[3]/NET0131 ,
		\si[3]_pad ,
		_w561_
	);
	LUT2 #(
		.INIT('h8)
	) name99 (
		\P2_datao_reg[0]/NET0131 ,
		\si[0]_pad ,
		_w562_
	);
	LUT4 #(
		.INIT('hec80)
	) name100 (
		\P2_datao_reg[0]/NET0131 ,
		\P2_datao_reg[1]/NET0131 ,
		\si[0]_pad ,
		\si[1]_pad ,
		_w563_
	);
	LUT3 #(
		.INIT('he8)
	) name101 (
		\P2_datao_reg[2]/NET0131 ,
		\si[2]_pad ,
		_w563_,
		_w564_
	);
	LUT4 #(
		.INIT('h0107)
	) name102 (
		\P2_datao_reg[2]/NET0131 ,
		\si[2]_pad ,
		_w561_,
		_w563_,
		_w565_
	);
	LUT2 #(
		.INIT('h1)
	) name103 (
		\P2_datao_reg[4]/NET0131 ,
		\si[4]_pad ,
		_w566_
	);
	LUT2 #(
		.INIT('h1)
	) name104 (
		\P2_datao_reg[3]/NET0131 ,
		\si[3]_pad ,
		_w567_
	);
	LUT4 #(
		.INIT('hfac8)
	) name105 (
		\P2_datao_reg[3]/NET0131 ,
		\P2_datao_reg[4]/NET0131 ,
		\si[3]_pad ,
		\si[4]_pad ,
		_w568_
	);
	LUT3 #(
		.INIT('h45)
	) name106 (
		_w560_,
		_w565_,
		_w568_,
		_w569_
	);
	LUT2 #(
		.INIT('h1)
	) name107 (
		\P2_datao_reg[5]/NET0131 ,
		\si[5]_pad ,
		_w570_
	);
	LUT4 #(
		.INIT('hfac8)
	) name108 (
		\P2_datao_reg[5]/NET0131 ,
		\P2_datao_reg[6]/NET0131 ,
		\si[5]_pad ,
		\si[6]_pad ,
		_w571_
	);
	LUT2 #(
		.INIT('h1)
	) name109 (
		\P2_datao_reg[7]/NET0131 ,
		\si[7]_pad ,
		_w572_
	);
	LUT4 #(
		.INIT('hfac8)
	) name110 (
		\P2_datao_reg[7]/NET0131 ,
		\P2_datao_reg[8]/NET0131 ,
		\si[7]_pad ,
		\si[8]_pad ,
		_w573_
	);
	LUT2 #(
		.INIT('h8)
	) name111 (
		_w571_,
		_w573_,
		_w574_
	);
	LUT4 #(
		.INIT('hba00)
	) name112 (
		_w560_,
		_w565_,
		_w568_,
		_w574_,
		_w575_
	);
	LUT2 #(
		.INIT('h8)
	) name113 (
		\P2_datao_reg[8]/NET0131 ,
		\si[8]_pad ,
		_w576_
	);
	LUT4 #(
		.INIT('hec80)
	) name114 (
		\P2_datao_reg[5]/NET0131 ,
		\P2_datao_reg[6]/NET0131 ,
		\si[5]_pad ,
		\si[6]_pad ,
		_w577_
	);
	LUT2 #(
		.INIT('h8)
	) name115 (
		\P2_datao_reg[7]/NET0131 ,
		\si[7]_pad ,
		_w578_
	);
	LUT4 #(
		.INIT('h1113)
	) name116 (
		_w573_,
		_w576_,
		_w577_,
		_w578_,
		_w579_
	);
	LUT2 #(
		.INIT('h1)
	) name117 (
		\P2_datao_reg[10]/NET0131 ,
		\si[10]_pad ,
		_w580_
	);
	LUT4 #(
		.INIT('hfac8)
	) name118 (
		\P2_datao_reg[10]/NET0131 ,
		\P2_datao_reg[11]/NET0131 ,
		\si[10]_pad ,
		\si[11]_pad ,
		_w581_
	);
	LUT2 #(
		.INIT('h1)
	) name119 (
		\P2_datao_reg[12]/NET0131 ,
		\si[12]_pad ,
		_w582_
	);
	LUT2 #(
		.INIT('h1)
	) name120 (
		\P2_datao_reg[9]/NET0131 ,
		\si[9]_pad ,
		_w583_
	);
	LUT4 #(
		.INIT('hfac8)
	) name121 (
		\P2_datao_reg[12]/NET0131 ,
		\P2_datao_reg[9]/NET0131 ,
		\si[12]_pad ,
		\si[9]_pad ,
		_w584_
	);
	LUT2 #(
		.INIT('h8)
	) name122 (
		_w581_,
		_w584_,
		_w585_
	);
	LUT2 #(
		.INIT('h8)
	) name123 (
		\P2_datao_reg[12]/NET0131 ,
		\si[12]_pad ,
		_w586_
	);
	LUT2 #(
		.INIT('h8)
	) name124 (
		\P2_datao_reg[10]/NET0131 ,
		\si[10]_pad ,
		_w587_
	);
	LUT4 #(
		.INIT('he8a0)
	) name125 (
		\P2_datao_reg[10]/NET0131 ,
		\P2_datao_reg[9]/NET0131 ,
		\si[10]_pad ,
		\si[9]_pad ,
		_w588_
	);
	LUT2 #(
		.INIT('h8)
	) name126 (
		\P2_datao_reg[11]/NET0131 ,
		\si[11]_pad ,
		_w589_
	);
	LUT4 #(
		.INIT('hfac8)
	) name127 (
		\P2_datao_reg[11]/NET0131 ,
		\P2_datao_reg[12]/NET0131 ,
		\si[11]_pad ,
		\si[12]_pad ,
		_w590_
	);
	LUT4 #(
		.INIT('h0155)
	) name128 (
		_w586_,
		_w588_,
		_w589_,
		_w590_,
		_w591_
	);
	LUT4 #(
		.INIT('h4f00)
	) name129 (
		_w575_,
		_w579_,
		_w585_,
		_w591_,
		_w592_
	);
	LUT2 #(
		.INIT('h1)
	) name130 (
		\P2_datao_reg[17]/NET0131 ,
		\si[17]_pad ,
		_w593_
	);
	LUT2 #(
		.INIT('h1)
	) name131 (
		\P2_datao_reg[20]/NET0131 ,
		\si[20]_pad ,
		_w594_
	);
	LUT2 #(
		.INIT('h1)
	) name132 (
		\P2_datao_reg[19]/NET0131 ,
		\si[19]_pad ,
		_w595_
	);
	LUT2 #(
		.INIT('h1)
	) name133 (
		\P2_datao_reg[18]/NET0131 ,
		\si[18]_pad ,
		_w596_
	);
	LUT4 #(
		.INIT('hfac8)
	) name134 (
		\P2_datao_reg[18]/NET0131 ,
		\P2_datao_reg[19]/NET0131 ,
		\si[18]_pad ,
		\si[19]_pad ,
		_w597_
	);
	LUT3 #(
		.INIT('h10)
	) name135 (
		_w593_,
		_w594_,
		_w597_,
		_w598_
	);
	LUT2 #(
		.INIT('h1)
	) name136 (
		\P2_datao_reg[16]/NET0131 ,
		\si[16]_pad ,
		_w599_
	);
	LUT2 #(
		.INIT('h1)
	) name137 (
		\P2_datao_reg[15]/NET0131 ,
		\si[15]_pad ,
		_w600_
	);
	LUT2 #(
		.INIT('h1)
	) name138 (
		\P2_datao_reg[14]/NET0131 ,
		\si[14]_pad ,
		_w601_
	);
	LUT4 #(
		.INIT('hfac8)
	) name139 (
		\P2_datao_reg[14]/NET0131 ,
		\P2_datao_reg[15]/NET0131 ,
		\si[14]_pad ,
		\si[15]_pad ,
		_w602_
	);
	LUT2 #(
		.INIT('h1)
	) name140 (
		\P2_datao_reg[13]/NET0131 ,
		\si[13]_pad ,
		_w603_
	);
	LUT3 #(
		.INIT('h04)
	) name141 (
		_w599_,
		_w602_,
		_w603_,
		_w604_
	);
	LUT2 #(
		.INIT('h8)
	) name142 (
		_w598_,
		_w604_,
		_w605_
	);
	LUT4 #(
		.INIT('h135f)
	) name143 (
		\P2_datao_reg[15]/NET0131 ,
		\P2_datao_reg[16]/NET0131 ,
		\si[15]_pad ,
		\si[16]_pad ,
		_w606_
	);
	LUT4 #(
		.INIT('h135f)
	) name144 (
		\P2_datao_reg[13]/NET0131 ,
		\P2_datao_reg[14]/NET0131 ,
		\si[13]_pad ,
		\si[14]_pad ,
		_w607_
	);
	LUT4 #(
		.INIT('h0545)
	) name145 (
		_w599_,
		_w602_,
		_w606_,
		_w607_,
		_w608_
	);
	LUT4 #(
		.INIT('hec80)
	) name146 (
		\P2_datao_reg[19]/NET0131 ,
		\P2_datao_reg[20]/NET0131 ,
		\si[19]_pad ,
		\si[20]_pad ,
		_w609_
	);
	LUT4 #(
		.INIT('h135f)
	) name147 (
		\P2_datao_reg[17]/NET0131 ,
		\P2_datao_reg[18]/NET0131 ,
		\si[17]_pad ,
		\si[18]_pad ,
		_w610_
	);
	LUT4 #(
		.INIT('h0f0b)
	) name148 (
		_w594_,
		_w597_,
		_w609_,
		_w610_,
		_w611_
	);
	LUT3 #(
		.INIT('h70)
	) name149 (
		_w598_,
		_w608_,
		_w611_,
		_w612_
	);
	LUT3 #(
		.INIT('hb0)
	) name150 (
		_w592_,
		_w605_,
		_w612_,
		_w613_
	);
	LUT2 #(
		.INIT('h4)
	) name151 (
		_w548_,
		_w551_,
		_w614_
	);
	LUT4 #(
		.INIT('hfac8)
	) name152 (
		\P2_datao_reg[21]/NET0131 ,
		\P2_datao_reg[22]/NET0131 ,
		\si[21]_pad ,
		\si[22]_pad ,
		_w615_
	);
	LUT2 #(
		.INIT('h8)
	) name153 (
		_w553_,
		_w615_,
		_w616_
	);
	LUT3 #(
		.INIT('h40)
	) name154 (
		_w546_,
		_w553_,
		_w615_,
		_w617_
	);
	LUT2 #(
		.INIT('h8)
	) name155 (
		_w614_,
		_w617_,
		_w618_
	);
	LUT4 #(
		.INIT('h4f00)
	) name156 (
		_w592_,
		_w605_,
		_w612_,
		_w618_,
		_w619_
	);
	LUT4 #(
		.INIT('h1114)
	) name157 (
		_w542_,
		_w545_,
		_w559_,
		_w619_,
		_w620_
	);
	LUT3 #(
		.INIT('h54)
	) name158 (
		_w541_,
		_w543_,
		_w620_,
		_w621_
	);
	LUT3 #(
		.INIT('h01)
	) name159 (
		\P1_IR_reg[27]/NET0131 ,
		\P1_IR_reg[28]/NET0131 ,
		\P1_IR_reg[29]/NET0131 ,
		_w622_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name160 (
		\P1_IR_reg[26]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		_w515_,
		_w622_,
		_w623_
	);
	LUT3 #(
		.INIT('h56)
	) name161 (
		\P1_IR_reg[30]/NET0131 ,
		_w513_,
		_w623_,
		_w624_
	);
	LUT4 #(
		.INIT('h0001)
	) name162 (
		\P1_IR_reg[25]/NET0131 ,
		\P1_IR_reg[26]/NET0131 ,
		\P1_IR_reg[27]/NET0131 ,
		\P1_IR_reg[28]/NET0131 ,
		_w625_
	);
	LUT2 #(
		.INIT('h2)
	) name163 (
		\P1_IR_reg[31]/NET0131 ,
		_w625_,
		_w626_
	);
	LUT3 #(
		.INIT('h56)
	) name164 (
		\P1_IR_reg[29]/NET0131 ,
		_w521_,
		_w626_,
		_w627_
	);
	LUT3 #(
		.INIT('h20)
	) name165 (
		\P1_reg1_reg[29]/NET0131 ,
		_w624_,
		_w627_,
		_w628_
	);
	LUT2 #(
		.INIT('h8)
	) name166 (
		_w624_,
		_w627_,
		_w629_
	);
	LUT4 #(
		.INIT('h8000)
	) name167 (
		\P1_reg3_reg[3]/NET0131 ,
		\P1_reg3_reg[4]/NET0131 ,
		\P1_reg3_reg[5]/NET0131 ,
		\P1_reg3_reg[6]/NET0131 ,
		_w630_
	);
	LUT4 #(
		.INIT('h8000)
	) name168 (
		\P1_reg3_reg[7]/NET0131 ,
		\P1_reg3_reg[8]/NET0131 ,
		\P1_reg3_reg[9]/NET0131 ,
		_w630_,
		_w631_
	);
	LUT4 #(
		.INIT('h8000)
	) name169 (
		\P1_reg3_reg[10]/NET0131 ,
		\P1_reg3_reg[11]/NET0131 ,
		\P1_reg3_reg[12]/NET0131 ,
		_w631_,
		_w632_
	);
	LUT4 #(
		.INIT('h8000)
	) name170 (
		\P1_reg3_reg[15]/NET0131 ,
		\P1_reg3_reg[16]/NET0131 ,
		\P1_reg3_reg[17]/NET0131 ,
		\P1_reg3_reg[18]/NET0131 ,
		_w633_
	);
	LUT4 #(
		.INIT('h8000)
	) name171 (
		\P1_reg3_reg[13]/NET0131 ,
		\P1_reg3_reg[14]/NET0131 ,
		_w632_,
		_w633_,
		_w634_
	);
	LUT2 #(
		.INIT('h8)
	) name172 (
		\P1_reg3_reg[19]/NET0131 ,
		\P1_reg3_reg[20]/NET0131 ,
		_w635_
	);
	LUT4 #(
		.INIT('h8000)
	) name173 (
		\P1_reg3_reg[19]/NET0131 ,
		\P1_reg3_reg[20]/NET0131 ,
		\P1_reg3_reg[21]/NET0131 ,
		\P1_reg3_reg[22]/NET0131 ,
		_w636_
	);
	LUT2 #(
		.INIT('h8)
	) name174 (
		\P1_reg3_reg[24]/NET0131 ,
		\P1_reg3_reg[25]/NET0131 ,
		_w637_
	);
	LUT4 #(
		.INIT('h8000)
	) name175 (
		\P1_reg3_reg[23]/NET0131 ,
		\P1_reg3_reg[26]/NET0131 ,
		\P1_reg3_reg[27]/NET0131 ,
		\P1_reg3_reg[28]/NET0131 ,
		_w638_
	);
	LUT3 #(
		.INIT('h80)
	) name176 (
		_w637_,
		_w636_,
		_w638_,
		_w639_
	);
	LUT2 #(
		.INIT('h8)
	) name177 (
		_w634_,
		_w639_,
		_w640_
	);
	LUT4 #(
		.INIT('h8000)
	) name178 (
		_w624_,
		_w627_,
		_w634_,
		_w639_,
		_w641_
	);
	LUT4 #(
		.INIT('hff35)
	) name179 (
		\P1_reg0_reg[29]/NET0131 ,
		\P1_reg2_reg[29]/NET0131 ,
		_w624_,
		_w627_,
		_w642_
	);
	LUT3 #(
		.INIT('h10)
	) name180 (
		_w628_,
		_w641_,
		_w642_,
		_w643_
	);
	LUT3 #(
		.INIT('hef)
	) name181 (
		_w628_,
		_w641_,
		_w642_,
		_w644_
	);
	LUT4 #(
		.INIT('h5400)
	) name182 (
		_w541_,
		_w543_,
		_w620_,
		_w643_,
		_w645_
	);
	LUT4 #(
		.INIT('h00ab)
	) name183 (
		_w541_,
		_w543_,
		_w620_,
		_w643_,
		_w646_
	);
	LUT4 #(
		.INIT('hab54)
	) name184 (
		_w541_,
		_w543_,
		_w620_,
		_w643_,
		_w647_
	);
	LUT4 #(
		.INIT('h1000)
	) name185 (
		\P1_IR_reg[14]/NET0131 ,
		\P1_IR_reg[15]/NET0131 ,
		_w503_,
		_w504_,
		_w648_
	);
	LUT3 #(
		.INIT('h10)
	) name186 (
		\P1_IR_reg[16]/NET0131 ,
		\P1_IR_reg[17]/NET0131 ,
		_w648_,
		_w649_
	);
	LUT4 #(
		.INIT('he0f0)
	) name187 (
		\P1_IR_reg[16]/NET0131 ,
		\P1_IR_reg[17]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		_w648_,
		_w650_
	);
	LUT2 #(
		.INIT('h8)
	) name188 (
		\P1_IR_reg[18]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		_w651_
	);
	LUT3 #(
		.INIT('h56)
	) name189 (
		\P1_IR_reg[19]/NET0131 ,
		_w650_,
		_w651_,
		_w652_
	);
	LUT2 #(
		.INIT('h2)
	) name190 (
		_w541_,
		_w652_,
		_w653_
	);
	LUT4 #(
		.INIT('hfac8)
	) name191 (
		\P2_datao_reg[16]/NET0131 ,
		\P2_datao_reg[17]/NET0131 ,
		\si[16]_pad ,
		\si[17]_pad ,
		_w654_
	);
	LUT3 #(
		.INIT('h10)
	) name192 (
		_w596_,
		_w600_,
		_w654_,
		_w655_
	);
	LUT2 #(
		.INIT('h4)
	) name193 (
		_w566_,
		_w571_,
		_w656_
	);
	LUT4 #(
		.INIT('h00e8)
	) name194 (
		\P2_datao_reg[2]/NET0131 ,
		\si[2]_pad ,
		_w563_,
		_w567_,
		_w657_
	);
	LUT4 #(
		.INIT('h135f)
	) name195 (
		\P2_datao_reg[3]/NET0131 ,
		\P2_datao_reg[4]/NET0131 ,
		\si[3]_pad ,
		\si[4]_pad ,
		_w658_
	);
	LUT4 #(
		.INIT('h1511)
	) name196 (
		_w577_,
		_w656_,
		_w657_,
		_w658_,
		_w659_
	);
	LUT3 #(
		.INIT('h02)
	) name197 (
		_w573_,
		_w580_,
		_w583_,
		_w660_
	);
	LUT4 #(
		.INIT('h135f)
	) name198 (
		\P2_datao_reg[7]/NET0131 ,
		\P2_datao_reg[8]/NET0131 ,
		\si[7]_pad ,
		\si[8]_pad ,
		_w661_
	);
	LUT4 #(
		.INIT('hfac8)
	) name199 (
		\P2_datao_reg[8]/NET0131 ,
		\P2_datao_reg[9]/NET0131 ,
		\si[8]_pad ,
		\si[9]_pad ,
		_w662_
	);
	LUT4 #(
		.INIT('h3323)
	) name200 (
		_w580_,
		_w588_,
		_w662_,
		_w661_,
		_w663_
	);
	LUT3 #(
		.INIT('hb0)
	) name201 (
		_w659_,
		_w660_,
		_w663_,
		_w664_
	);
	LUT3 #(
		.INIT('h02)
	) name202 (
		_w590_,
		_w601_,
		_w603_,
		_w665_
	);
	LUT4 #(
		.INIT('h4f00)
	) name203 (
		_w659_,
		_w660_,
		_w663_,
		_w665_,
		_w666_
	);
	LUT4 #(
		.INIT('h135f)
	) name204 (
		\P2_datao_reg[11]/NET0131 ,
		\P2_datao_reg[12]/NET0131 ,
		\si[11]_pad ,
		\si[12]_pad ,
		_w667_
	);
	LUT4 #(
		.INIT('hfac8)
	) name205 (
		\P2_datao_reg[12]/NET0131 ,
		\P2_datao_reg[13]/NET0131 ,
		\si[12]_pad ,
		\si[13]_pad ,
		_w668_
	);
	LUT4 #(
		.INIT('h1511)
	) name206 (
		_w601_,
		_w607_,
		_w667_,
		_w668_,
		_w669_
	);
	LUT4 #(
		.INIT('h1505)
	) name207 (
		_w596_,
		_w606_,
		_w610_,
		_w654_,
		_w670_
	);
	LUT3 #(
		.INIT('h07)
	) name208 (
		_w655_,
		_w669_,
		_w670_,
		_w671_
	);
	LUT3 #(
		.INIT('h70)
	) name209 (
		_w655_,
		_w666_,
		_w671_,
		_w672_
	);
	LUT4 #(
		.INIT('h5956)
	) name210 (
		\P2_datao_reg[19]/NET0131 ,
		\si[19]_pad ,
		_w542_,
		_w672_,
		_w673_
	);
	LUT3 #(
		.INIT('h23)
	) name211 (
		_w541_,
		_w653_,
		_w673_,
		_w674_
	);
	LUT2 #(
		.INIT('h6)
	) name212 (
		\P1_reg3_reg[19]/NET0131 ,
		_w634_,
		_w675_
	);
	LUT4 #(
		.INIT('h4080)
	) name213 (
		\P1_reg3_reg[19]/NET0131 ,
		_w624_,
		_w627_,
		_w634_,
		_w676_
	);
	LUT3 #(
		.INIT('h20)
	) name214 (
		\P1_reg1_reg[19]/NET0131 ,
		_w624_,
		_w627_,
		_w677_
	);
	LUT4 #(
		.INIT('hff35)
	) name215 (
		\P1_reg0_reg[19]/NET0131 ,
		\P1_reg2_reg[19]/NET0131 ,
		_w624_,
		_w627_,
		_w678_
	);
	LUT3 #(
		.INIT('h10)
	) name216 (
		_w677_,
		_w676_,
		_w678_,
		_w679_
	);
	LUT3 #(
		.INIT('hef)
	) name217 (
		_w677_,
		_w676_,
		_w678_,
		_w680_
	);
	LUT4 #(
		.INIT('h7200)
	) name218 (
		_w541_,
		_w652_,
		_w673_,
		_w679_,
		_w681_
	);
	LUT3 #(
		.INIT('h04)
	) name219 (
		_w566_,
		_w571_,
		_w572_,
		_w682_
	);
	LUT4 #(
		.INIT('h135f)
	) name220 (
		\P2_datao_reg[6]/NET0131 ,
		\P2_datao_reg[7]/NET0131 ,
		\si[6]_pad ,
		\si[7]_pad ,
		_w683_
	);
	LUT4 #(
		.INIT('h135f)
	) name221 (
		\P2_datao_reg[4]/NET0131 ,
		\P2_datao_reg[5]/NET0131 ,
		\si[4]_pad ,
		\si[5]_pad ,
		_w684_
	);
	LUT4 #(
		.INIT('h0323)
	) name222 (
		_w571_,
		_w572_,
		_w683_,
		_w684_,
		_w685_
	);
	LUT4 #(
		.INIT('h00ef)
	) name223 (
		_w565_,
		_w567_,
		_w682_,
		_w685_,
		_w686_
	);
	LUT2 #(
		.INIT('h8)
	) name224 (
		_w581_,
		_w662_,
		_w687_
	);
	LUT4 #(
		.INIT('hec80)
	) name225 (
		\P2_datao_reg[8]/NET0131 ,
		\P2_datao_reg[9]/NET0131 ,
		\si[8]_pad ,
		\si[9]_pad ,
		_w688_
	);
	LUT4 #(
		.INIT('h0507)
	) name226 (
		_w581_,
		_w587_,
		_w589_,
		_w688_,
		_w689_
	);
	LUT3 #(
		.INIT('hb0)
	) name227 (
		_w686_,
		_w687_,
		_w689_,
		_w690_
	);
	LUT3 #(
		.INIT('h04)
	) name228 (
		_w582_,
		_w602_,
		_w603_,
		_w691_
	);
	LUT4 #(
		.INIT('h4f00)
	) name229 (
		_w686_,
		_w687_,
		_w689_,
		_w691_,
		_w692_
	);
	LUT4 #(
		.INIT('hec80)
	) name230 (
		\P2_datao_reg[14]/NET0131 ,
		\P2_datao_reg[15]/NET0131 ,
		\si[14]_pad ,
		\si[15]_pad ,
		_w693_
	);
	LUT4 #(
		.INIT('hec80)
	) name231 (
		\P2_datao_reg[12]/NET0131 ,
		\P2_datao_reg[13]/NET0131 ,
		\si[12]_pad ,
		\si[13]_pad ,
		_w694_
	);
	LUT3 #(
		.INIT('h13)
	) name232 (
		_w602_,
		_w693_,
		_w694_,
		_w695_
	);
	LUT3 #(
		.INIT('h10)
	) name233 (
		_w595_,
		_w596_,
		_w654_,
		_w696_
	);
	LUT4 #(
		.INIT('hec80)
	) name234 (
		\P2_datao_reg[18]/NET0131 ,
		\P2_datao_reg[19]/NET0131 ,
		\si[18]_pad ,
		\si[19]_pad ,
		_w697_
	);
	LUT4 #(
		.INIT('hec80)
	) name235 (
		\P2_datao_reg[16]/NET0131 ,
		\P2_datao_reg[17]/NET0131 ,
		\si[16]_pad ,
		\si[17]_pad ,
		_w698_
	);
	LUT3 #(
		.INIT('h13)
	) name236 (
		_w597_,
		_w697_,
		_w698_,
		_w699_
	);
	LUT4 #(
		.INIT('h4f00)
	) name237 (
		_w692_,
		_w695_,
		_w696_,
		_w699_,
		_w700_
	);
	LUT4 #(
		.INIT('h5956)
	) name238 (
		\P2_datao_reg[20]/NET0131 ,
		\si[20]_pad ,
		_w542_,
		_w700_,
		_w701_
	);
	LUT2 #(
		.INIT('h1)
	) name239 (
		_w541_,
		_w701_,
		_w702_
	);
	LUT3 #(
		.INIT('h6c)
	) name240 (
		\P1_reg3_reg[19]/NET0131 ,
		\P1_reg3_reg[20]/NET0131 ,
		_w634_,
		_w703_
	);
	LUT3 #(
		.INIT('h08)
	) name241 (
		\P1_reg2_reg[20]/NET0131 ,
		_w624_,
		_w627_,
		_w704_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name242 (
		\P1_reg0_reg[20]/NET0131 ,
		\P1_reg1_reg[20]/NET0131 ,
		_w624_,
		_w627_,
		_w705_
	);
	LUT4 #(
		.INIT('h1300)
	) name243 (
		_w629_,
		_w704_,
		_w703_,
		_w705_,
		_w706_
	);
	LUT4 #(
		.INIT('hecff)
	) name244 (
		_w629_,
		_w704_,
		_w703_,
		_w705_,
		_w707_
	);
	LUT3 #(
		.INIT('he0)
	) name245 (
		_w541_,
		_w701_,
		_w706_,
		_w708_
	);
	LUT2 #(
		.INIT('h1)
	) name246 (
		_w681_,
		_w708_,
		_w709_
	);
	LUT2 #(
		.INIT('h8)
	) name247 (
		\P2_datao_reg[17]/NET0131 ,
		_w542_,
		_w710_
	);
	LUT4 #(
		.INIT('hb000)
	) name248 (
		_w575_,
		_w579_,
		_w585_,
		_w604_,
		_w711_
	);
	LUT3 #(
		.INIT('h0b)
	) name249 (
		_w591_,
		_w604_,
		_w608_,
		_w712_
	);
	LUT2 #(
		.INIT('h6)
	) name250 (
		\P2_datao_reg[17]/NET0131 ,
		\si[17]_pad ,
		_w713_
	);
	LUT4 #(
		.INIT('h1045)
	) name251 (
		_w542_,
		_w711_,
		_w712_,
		_w713_,
		_w714_
	);
	LUT4 #(
		.INIT('h6c3c)
	) name252 (
		\P1_IR_reg[16]/NET0131 ,
		\P1_IR_reg[17]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		_w648_,
		_w715_
	);
	LUT3 #(
		.INIT('h10)
	) name253 (
		_w537_,
		_w540_,
		_w715_,
		_w716_
	);
	LUT4 #(
		.INIT('h00ab)
	) name254 (
		_w541_,
		_w710_,
		_w714_,
		_w716_,
		_w717_
	);
	LUT4 #(
		.INIT('h8000)
	) name255 (
		\P1_reg3_reg[13]/NET0131 ,
		\P1_reg3_reg[14]/NET0131 ,
		\P1_reg3_reg[15]/NET0131 ,
		_w632_,
		_w718_
	);
	LUT3 #(
		.INIT('h6c)
	) name256 (
		\P1_reg3_reg[16]/NET0131 ,
		\P1_reg3_reg[17]/NET0131 ,
		_w718_,
		_w719_
	);
	LUT3 #(
		.INIT('h20)
	) name257 (
		\P1_reg1_reg[17]/NET0131 ,
		_w624_,
		_w627_,
		_w720_
	);
	LUT4 #(
		.INIT('hff35)
	) name258 (
		\P1_reg0_reg[17]/NET0131 ,
		\P1_reg2_reg[17]/NET0131 ,
		_w624_,
		_w627_,
		_w721_
	);
	LUT4 #(
		.INIT('h1300)
	) name259 (
		_w629_,
		_w720_,
		_w719_,
		_w721_,
		_w722_
	);
	LUT4 #(
		.INIT('hecff)
	) name260 (
		_w629_,
		_w720_,
		_w719_,
		_w721_,
		_w723_
	);
	LUT2 #(
		.INIT('h8)
	) name261 (
		_w717_,
		_w722_,
		_w724_
	);
	LUT4 #(
		.INIT('h135f)
	) name262 (
		\P2_datao_reg[10]/NET0131 ,
		\P2_datao_reg[11]/NET0131 ,
		\si[10]_pad ,
		\si[11]_pad ,
		_w725_
	);
	LUT4 #(
		.INIT('h0f0d)
	) name263 (
		_w590_,
		_w603_,
		_w694_,
		_w725_,
		_w726_
	);
	LUT3 #(
		.INIT('h08)
	) name264 (
		_w571_,
		_w573_,
		_w583_,
		_w727_
	);
	LUT4 #(
		.INIT('h4f00)
	) name265 (
		_w565_,
		_w568_,
		_w684_,
		_w727_,
		_w728_
	);
	LUT4 #(
		.INIT('h0f0d)
	) name266 (
		_w573_,
		_w583_,
		_w688_,
		_w683_,
		_w729_
	);
	LUT2 #(
		.INIT('h8)
	) name267 (
		_w581_,
		_w668_,
		_w730_
	);
	LUT4 #(
		.INIT('h20aa)
	) name268 (
		_w726_,
		_w728_,
		_w729_,
		_w730_,
		_w731_
	);
	LUT2 #(
		.INIT('h8)
	) name269 (
		_w602_,
		_w654_,
		_w732_
	);
	LUT3 #(
		.INIT('h13)
	) name270 (
		_w654_,
		_w698_,
		_w693_,
		_w733_
	);
	LUT3 #(
		.INIT('hb0)
	) name271 (
		_w731_,
		_w732_,
		_w733_,
		_w734_
	);
	LUT4 #(
		.INIT('h5956)
	) name272 (
		\P2_datao_reg[18]/NET0131 ,
		\si[18]_pad ,
		_w542_,
		_w734_,
		_w735_
	);
	LUT3 #(
		.INIT('ha6)
	) name273 (
		\P1_IR_reg[18]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		_w649_,
		_w736_
	);
	LUT2 #(
		.INIT('h8)
	) name274 (
		_w541_,
		_w736_,
		_w737_
	);
	LUT3 #(
		.INIT('h0e)
	) name275 (
		_w541_,
		_w735_,
		_w737_,
		_w738_
	);
	LUT4 #(
		.INIT('h070f)
	) name276 (
		\P1_reg3_reg[16]/NET0131 ,
		\P1_reg3_reg[17]/NET0131 ,
		\P1_reg3_reg[18]/NET0131 ,
		_w718_,
		_w739_
	);
	LUT2 #(
		.INIT('h1)
	) name277 (
		_w634_,
		_w739_,
		_w740_
	);
	LUT3 #(
		.INIT('h02)
	) name278 (
		_w629_,
		_w634_,
		_w739_,
		_w741_
	);
	LUT3 #(
		.INIT('h08)
	) name279 (
		\P1_reg2_reg[18]/NET0131 ,
		_w624_,
		_w627_,
		_w742_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name280 (
		\P1_reg0_reg[18]/NET0131 ,
		\P1_reg1_reg[18]/NET0131 ,
		_w624_,
		_w627_,
		_w743_
	);
	LUT2 #(
		.INIT('h4)
	) name281 (
		_w742_,
		_w743_,
		_w744_
	);
	LUT2 #(
		.INIT('h4)
	) name282 (
		_w741_,
		_w744_,
		_w745_
	);
	LUT2 #(
		.INIT('hb)
	) name283 (
		_w741_,
		_w744_,
		_w746_
	);
	LUT3 #(
		.INIT('h15)
	) name284 (
		_w724_,
		_w738_,
		_w745_,
		_w747_
	);
	LUT2 #(
		.INIT('h8)
	) name285 (
		_w709_,
		_w747_,
		_w748_
	);
	LUT2 #(
		.INIT('h6)
	) name286 (
		\P1_reg3_reg[13]/NET0131 ,
		_w632_,
		_w749_
	);
	LUT4 #(
		.INIT('h1fdf)
	) name287 (
		\P1_reg1_reg[13]/NET0131 ,
		_w624_,
		_w627_,
		_w749_,
		_w750_
	);
	LUT4 #(
		.INIT('hff35)
	) name288 (
		\P1_reg0_reg[13]/NET0131 ,
		\P1_reg2_reg[13]/NET0131 ,
		_w624_,
		_w627_,
		_w751_
	);
	LUT2 #(
		.INIT('h8)
	) name289 (
		_w750_,
		_w751_,
		_w752_
	);
	LUT2 #(
		.INIT('h7)
	) name290 (
		_w750_,
		_w751_,
		_w753_
	);
	LUT4 #(
		.INIT('h5956)
	) name291 (
		\P2_datao_reg[13]/NET0131 ,
		\si[13]_pad ,
		_w542_,
		_w592_,
		_w754_
	);
	LUT4 #(
		.INIT('hfe00)
	) name292 (
		\P1_IR_reg[10]/NET0131 ,
		\P1_IR_reg[11]/NET0131 ,
		\P1_IR_reg[12]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		_w755_
	);
	LUT4 #(
		.INIT('h55a6)
	) name293 (
		\P1_IR_reg[13]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		_w503_,
		_w755_,
		_w756_
	);
	LUT3 #(
		.INIT('h10)
	) name294 (
		_w537_,
		_w540_,
		_w756_,
		_w757_
	);
	LUT3 #(
		.INIT('h0e)
	) name295 (
		_w541_,
		_w754_,
		_w757_,
		_w758_
	);
	LUT4 #(
		.INIT('hff35)
	) name296 (
		\P1_reg0_reg[14]/NET0131 ,
		\P1_reg2_reg[14]/NET0131 ,
		_w624_,
		_w627_,
		_w759_
	);
	LUT3 #(
		.INIT('h6c)
	) name297 (
		\P1_reg3_reg[13]/NET0131 ,
		\P1_reg3_reg[14]/NET0131 ,
		_w632_,
		_w760_
	);
	LUT4 #(
		.INIT('h1fdf)
	) name298 (
		\P1_reg1_reg[14]/NET0131 ,
		_w624_,
		_w627_,
		_w760_,
		_w761_
	);
	LUT2 #(
		.INIT('h8)
	) name299 (
		_w759_,
		_w761_,
		_w762_
	);
	LUT2 #(
		.INIT('h7)
	) name300 (
		_w759_,
		_w761_,
		_w763_
	);
	LUT4 #(
		.INIT('h5956)
	) name301 (
		\P2_datao_reg[14]/NET0131 ,
		\si[14]_pad ,
		_w542_,
		_w731_,
		_w764_
	);
	LUT4 #(
		.INIT('h5999)
	) name302 (
		\P1_IR_reg[14]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		_w503_,
		_w504_,
		_w765_
	);
	LUT3 #(
		.INIT('h01)
	) name303 (
		_w537_,
		_w540_,
		_w765_,
		_w766_
	);
	LUT3 #(
		.INIT('h0e)
	) name304 (
		_w541_,
		_w764_,
		_w766_,
		_w767_
	);
	LUT4 #(
		.INIT('h0777)
	) name305 (
		_w752_,
		_w758_,
		_w762_,
		_w767_,
		_w768_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name306 (
		\P1_reg0_reg[15]/NET0131 ,
		\P1_reg1_reg[15]/NET0131 ,
		_w624_,
		_w627_,
		_w769_
	);
	LUT4 #(
		.INIT('h78f0)
	) name307 (
		\P1_reg3_reg[13]/NET0131 ,
		\P1_reg3_reg[14]/NET0131 ,
		\P1_reg3_reg[15]/NET0131 ,
		_w632_,
		_w770_
	);
	LUT4 #(
		.INIT('h37f7)
	) name308 (
		\P1_reg2_reg[15]/NET0131 ,
		_w624_,
		_w627_,
		_w770_,
		_w771_
	);
	LUT2 #(
		.INIT('h8)
	) name309 (
		_w769_,
		_w771_,
		_w772_
	);
	LUT2 #(
		.INIT('h7)
	) name310 (
		_w769_,
		_w771_,
		_w773_
	);
	LUT2 #(
		.INIT('h8)
	) name311 (
		\P2_datao_reg[15]/NET0131 ,
		_w542_,
		_w774_
	);
	LUT2 #(
		.INIT('h6)
	) name312 (
		\P2_datao_reg[15]/NET0131 ,
		\si[15]_pad ,
		_w775_
	);
	LUT4 #(
		.INIT('h0154)
	) name313 (
		_w542_,
		_w666_,
		_w669_,
		_w775_,
		_w776_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name314 (
		\P1_IR_reg[14]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		_w503_,
		_w504_,
		_w777_
	);
	LUT2 #(
		.INIT('h9)
	) name315 (
		\P1_IR_reg[15]/NET0131 ,
		_w777_,
		_w778_
	);
	LUT3 #(
		.INIT('h01)
	) name316 (
		_w537_,
		_w540_,
		_w778_,
		_w779_
	);
	LUT4 #(
		.INIT('h00ab)
	) name317 (
		_w541_,
		_w774_,
		_w776_,
		_w779_,
		_w780_
	);
	LUT2 #(
		.INIT('h8)
	) name318 (
		\P2_datao_reg[16]/NET0131 ,
		_w542_,
		_w781_
	);
	LUT2 #(
		.INIT('h6)
	) name319 (
		\P2_datao_reg[16]/NET0131 ,
		\si[16]_pad ,
		_w782_
	);
	LUT4 #(
		.INIT('h1045)
	) name320 (
		_w542_,
		_w692_,
		_w695_,
		_w782_,
		_w783_
	);
	LUT3 #(
		.INIT('ha6)
	) name321 (
		\P1_IR_reg[16]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		_w648_,
		_w784_
	);
	LUT3 #(
		.INIT('h10)
	) name322 (
		_w537_,
		_w540_,
		_w784_,
		_w785_
	);
	LUT4 #(
		.INIT('h00ab)
	) name323 (
		_w541_,
		_w781_,
		_w783_,
		_w785_,
		_w786_
	);
	LUT2 #(
		.INIT('h6)
	) name324 (
		\P1_reg3_reg[16]/NET0131 ,
		_w718_,
		_w787_
	);
	LUT4 #(
		.INIT('h4080)
	) name325 (
		\P1_reg3_reg[16]/NET0131 ,
		_w624_,
		_w627_,
		_w718_,
		_w788_
	);
	LUT3 #(
		.INIT('h08)
	) name326 (
		\P1_reg2_reg[16]/NET0131 ,
		_w624_,
		_w627_,
		_w789_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name327 (
		\P1_reg0_reg[16]/NET0131 ,
		\P1_reg1_reg[16]/NET0131 ,
		_w624_,
		_w627_,
		_w790_
	);
	LUT3 #(
		.INIT('h10)
	) name328 (
		_w789_,
		_w788_,
		_w790_,
		_w791_
	);
	LUT3 #(
		.INIT('hef)
	) name329 (
		_w789_,
		_w788_,
		_w790_,
		_w792_
	);
	LUT4 #(
		.INIT('h0777)
	) name330 (
		_w772_,
		_w780_,
		_w786_,
		_w791_,
		_w793_
	);
	LUT2 #(
		.INIT('h8)
	) name331 (
		_w768_,
		_w793_,
		_w794_
	);
	LUT3 #(
		.INIT('h80)
	) name332 (
		_w709_,
		_w747_,
		_w794_,
		_w795_
	);
	LUT3 #(
		.INIT('h6c)
	) name333 (
		\P1_reg3_reg[10]/NET0131 ,
		\P1_reg3_reg[11]/NET0131 ,
		_w631_,
		_w796_
	);
	LUT4 #(
		.INIT('h3dfd)
	) name334 (
		\P1_reg0_reg[11]/NET0131 ,
		_w624_,
		_w627_,
		_w796_,
		_w797_
	);
	LUT4 #(
		.INIT('hf53f)
	) name335 (
		\P1_reg1_reg[11]/NET0131 ,
		\P1_reg2_reg[11]/NET0131 ,
		_w624_,
		_w627_,
		_w798_
	);
	LUT2 #(
		.INIT('h8)
	) name336 (
		_w797_,
		_w798_,
		_w799_
	);
	LUT2 #(
		.INIT('h7)
	) name337 (
		_w797_,
		_w798_,
		_w800_
	);
	LUT4 #(
		.INIT('h5956)
	) name338 (
		\P2_datao_reg[11]/NET0131 ,
		\si[11]_pad ,
		_w542_,
		_w664_,
		_w801_
	);
	LUT4 #(
		.INIT('h6c3c)
	) name339 (
		\P1_IR_reg[10]/NET0131 ,
		\P1_IR_reg[11]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		_w503_,
		_w802_
	);
	LUT3 #(
		.INIT('h10)
	) name340 (
		_w537_,
		_w540_,
		_w802_,
		_w803_
	);
	LUT3 #(
		.INIT('h0e)
	) name341 (
		_w541_,
		_w801_,
		_w803_,
		_w804_
	);
	LUT4 #(
		.INIT('hf53f)
	) name342 (
		\P1_reg1_reg[12]/NET0131 ,
		\P1_reg2_reg[12]/NET0131 ,
		_w624_,
		_w627_,
		_w805_
	);
	LUT4 #(
		.INIT('h78f0)
	) name343 (
		\P1_reg3_reg[10]/NET0131 ,
		\P1_reg3_reg[11]/NET0131 ,
		\P1_reg3_reg[12]/NET0131 ,
		_w631_,
		_w806_
	);
	LUT4 #(
		.INIT('h3dfd)
	) name344 (
		\P1_reg0_reg[12]/NET0131 ,
		_w624_,
		_w627_,
		_w806_,
		_w807_
	);
	LUT2 #(
		.INIT('h8)
	) name345 (
		_w805_,
		_w807_,
		_w808_
	);
	LUT2 #(
		.INIT('h7)
	) name346 (
		_w805_,
		_w807_,
		_w809_
	);
	LUT4 #(
		.INIT('h5956)
	) name347 (
		\P2_datao_reg[12]/NET0131 ,
		\si[12]_pad ,
		_w542_,
		_w690_,
		_w810_
	);
	LUT3 #(
		.INIT('he0)
	) name348 (
		\P1_IR_reg[10]/NET0131 ,
		\P1_IR_reg[11]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		_w811_
	);
	LUT4 #(
		.INIT('h55a6)
	) name349 (
		\P1_IR_reg[12]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		_w503_,
		_w811_,
		_w812_
	);
	LUT3 #(
		.INIT('h10)
	) name350 (
		_w537_,
		_w540_,
		_w812_,
		_w813_
	);
	LUT3 #(
		.INIT('h0e)
	) name351 (
		_w541_,
		_w810_,
		_w813_,
		_w814_
	);
	LUT4 #(
		.INIT('h0777)
	) name352 (
		_w799_,
		_w804_,
		_w808_,
		_w814_,
		_w815_
	);
	LUT2 #(
		.INIT('h6)
	) name353 (
		\P1_reg3_reg[10]/NET0131 ,
		_w631_,
		_w816_
	);
	LUT4 #(
		.INIT('h3dfd)
	) name354 (
		\P1_reg0_reg[10]/NET0131 ,
		_w624_,
		_w627_,
		_w816_,
		_w817_
	);
	LUT4 #(
		.INIT('hf53f)
	) name355 (
		\P1_reg1_reg[10]/NET0131 ,
		\P1_reg2_reg[10]/NET0131 ,
		_w624_,
		_w627_,
		_w818_
	);
	LUT2 #(
		.INIT('h8)
	) name356 (
		_w817_,
		_w818_,
		_w819_
	);
	LUT2 #(
		.INIT('h7)
	) name357 (
		_w817_,
		_w818_,
		_w820_
	);
	LUT2 #(
		.INIT('h8)
	) name358 (
		\P2_datao_reg[10]/NET0131 ,
		_w542_,
		_w821_
	);
	LUT2 #(
		.INIT('h6)
	) name359 (
		\P2_datao_reg[10]/NET0131 ,
		\si[10]_pad ,
		_w822_
	);
	LUT4 #(
		.INIT('h1045)
	) name360 (
		_w542_,
		_w728_,
		_w729_,
		_w822_,
		_w823_
	);
	LUT4 #(
		.INIT('heee0)
	) name361 (
		_w537_,
		_w540_,
		_w821_,
		_w823_,
		_w824_
	);
	LUT3 #(
		.INIT('ha6)
	) name362 (
		\P1_IR_reg[10]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		_w503_,
		_w825_
	);
	LUT3 #(
		.INIT('h10)
	) name363 (
		_w537_,
		_w540_,
		_w825_,
		_w826_
	);
	LUT2 #(
		.INIT('h1)
	) name364 (
		_w824_,
		_w826_,
		_w827_
	);
	LUT4 #(
		.INIT('h0008)
	) name365 (
		_w817_,
		_w818_,
		_w824_,
		_w826_,
		_w828_
	);
	LUT4 #(
		.INIT('h7770)
	) name366 (
		_w817_,
		_w818_,
		_w824_,
		_w826_,
		_w829_
	);
	LUT4 #(
		.INIT('hff35)
	) name367 (
		\P1_reg0_reg[9]/NET0131 ,
		\P1_reg2_reg[9]/NET0131 ,
		_w624_,
		_w627_,
		_w830_
	);
	LUT4 #(
		.INIT('h78f0)
	) name368 (
		\P1_reg3_reg[7]/NET0131 ,
		\P1_reg3_reg[8]/NET0131 ,
		\P1_reg3_reg[9]/NET0131 ,
		_w630_,
		_w831_
	);
	LUT4 #(
		.INIT('h1fdf)
	) name369 (
		\P1_reg1_reg[9]/NET0131 ,
		_w624_,
		_w627_,
		_w831_,
		_w832_
	);
	LUT2 #(
		.INIT('h8)
	) name370 (
		_w830_,
		_w832_,
		_w833_
	);
	LUT2 #(
		.INIT('h7)
	) name371 (
		_w830_,
		_w832_,
		_w834_
	);
	LUT2 #(
		.INIT('h8)
	) name372 (
		\P2_datao_reg[9]/NET0131 ,
		_w542_,
		_w835_
	);
	LUT2 #(
		.INIT('h6)
	) name373 (
		\P2_datao_reg[9]/NET0131 ,
		\si[9]_pad ,
		_w836_
	);
	LUT4 #(
		.INIT('h1045)
	) name374 (
		_w542_,
		_w575_,
		_w579_,
		_w836_,
		_w837_
	);
	LUT4 #(
		.INIT('heee0)
	) name375 (
		_w537_,
		_w540_,
		_w835_,
		_w837_,
		_w838_
	);
	LUT4 #(
		.INIT('h1000)
	) name376 (
		\P1_IR_reg[4]/NET0131 ,
		\P1_IR_reg[5]/NET0131 ,
		_w500_,
		_w501_,
		_w839_
	);
	LUT4 #(
		.INIT('h785a)
	) name377 (
		\P1_IR_reg[31]/NET0131 ,
		\P1_IR_reg[8]/NET0131 ,
		\P1_IR_reg[9]/NET0131 ,
		_w839_,
		_w840_
	);
	LUT3 #(
		.INIT('h10)
	) name378 (
		_w537_,
		_w540_,
		_w840_,
		_w841_
	);
	LUT2 #(
		.INIT('h1)
	) name379 (
		_w838_,
		_w841_,
		_w842_
	);
	LUT4 #(
		.INIT('h7770)
	) name380 (
		_w830_,
		_w832_,
		_w838_,
		_w841_,
		_w843_
	);
	LUT3 #(
		.INIT('h54)
	) name381 (
		_w828_,
		_w829_,
		_w843_,
		_w844_
	);
	LUT4 #(
		.INIT('hfee0)
	) name382 (
		_w799_,
		_w804_,
		_w808_,
		_w814_,
		_w845_
	);
	LUT3 #(
		.INIT('h70)
	) name383 (
		_w815_,
		_w844_,
		_w845_,
		_w846_
	);
	LUT4 #(
		.INIT('h3ff5)
	) name384 (
		\P1_reg0_reg[2]/NET0131 ,
		\P1_reg3_reg[2]/NET0131 ,
		_w624_,
		_w627_,
		_w847_
	);
	LUT4 #(
		.INIT('hf53f)
	) name385 (
		\P1_reg1_reg[2]/NET0131 ,
		\P1_reg2_reg[2]/NET0131 ,
		_w624_,
		_w627_,
		_w848_
	);
	LUT2 #(
		.INIT('h8)
	) name386 (
		_w847_,
		_w848_,
		_w849_
	);
	LUT2 #(
		.INIT('h7)
	) name387 (
		_w847_,
		_w848_,
		_w850_
	);
	LUT4 #(
		.INIT('h5659)
	) name388 (
		\P2_datao_reg[2]/NET0131 ,
		\si[2]_pad ,
		_w542_,
		_w563_,
		_w851_
	);
	LUT4 #(
		.INIT('h1ef0)
	) name389 (
		\P1_IR_reg[0]/NET0131 ,
		\P1_IR_reg[1]/NET0131 ,
		\P1_IR_reg[2]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		_w852_
	);
	LUT4 #(
		.INIT('he0f1)
	) name390 (
		_w537_,
		_w540_,
		_w851_,
		_w852_,
		_w853_
	);
	LUT3 #(
		.INIT('h07)
	) name391 (
		_w847_,
		_w848_,
		_w853_,
		_w854_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name392 (
		\P1_reg2_reg[1]/NET0131 ,
		\P1_reg3_reg[1]/NET0131 ,
		_w624_,
		_w627_,
		_w855_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name393 (
		\P1_reg0_reg[1]/NET0131 ,
		\P1_reg1_reg[1]/NET0131 ,
		_w624_,
		_w627_,
		_w856_
	);
	LUT2 #(
		.INIT('h8)
	) name394 (
		_w855_,
		_w856_,
		_w857_
	);
	LUT2 #(
		.INIT('h7)
	) name395 (
		_w855_,
		_w856_,
		_w858_
	);
	LUT3 #(
		.INIT('h93)
	) name396 (
		\P1_IR_reg[0]/NET0131 ,
		\P1_IR_reg[1]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		_w859_
	);
	LUT4 #(
		.INIT('ha9a6)
	) name397 (
		\P2_datao_reg[1]/NET0131 ,
		\si[1]_pad ,
		_w542_,
		_w562_,
		_w860_
	);
	LUT4 #(
		.INIT('h10fe)
	) name398 (
		_w537_,
		_w540_,
		_w859_,
		_w860_,
		_w861_
	);
	LUT3 #(
		.INIT('h80)
	) name399 (
		_w855_,
		_w856_,
		_w861_,
		_w862_
	);
	LUT3 #(
		.INIT('h07)
	) name400 (
		_w855_,
		_w856_,
		_w861_,
		_w863_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name401 (
		\P1_reg2_reg[0]/NET0131 ,
		\P1_reg3_reg[0]/NET0131 ,
		_w624_,
		_w627_,
		_w864_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name402 (
		\P1_reg0_reg[0]/NET0131 ,
		\P1_reg1_reg[0]/NET0131 ,
		_w624_,
		_w627_,
		_w865_
	);
	LUT2 #(
		.INIT('h8)
	) name403 (
		_w864_,
		_w865_,
		_w866_
	);
	LUT2 #(
		.INIT('h7)
	) name404 (
		_w864_,
		_w865_,
		_w867_
	);
	LUT3 #(
		.INIT('ha6)
	) name405 (
		\P2_datao_reg[0]/NET0131 ,
		\si[0]_pad ,
		_w542_,
		_w868_
	);
	LUT4 #(
		.INIT('h01fd)
	) name406 (
		\P1_IR_reg[0]/NET0131 ,
		_w537_,
		_w540_,
		_w868_,
		_w869_
	);
	LUT3 #(
		.INIT('h07)
	) name407 (
		_w864_,
		_w865_,
		_w869_,
		_w870_
	);
	LUT3 #(
		.INIT('h54)
	) name408 (
		_w862_,
		_w863_,
		_w870_,
		_w871_
	);
	LUT4 #(
		.INIT('h4054)
	) name409 (
		_w854_,
		_w857_,
		_w861_,
		_w870_,
		_w872_
	);
	LUT3 #(
		.INIT('h80)
	) name410 (
		_w847_,
		_w848_,
		_w853_,
		_w873_
	);
	LUT4 #(
		.INIT('hcff5)
	) name411 (
		\P1_reg0_reg[3]/NET0131 ,
		\P1_reg3_reg[3]/NET0131 ,
		_w624_,
		_w627_,
		_w874_
	);
	LUT4 #(
		.INIT('hf53f)
	) name412 (
		\P1_reg1_reg[3]/NET0131 ,
		\P1_reg2_reg[3]/NET0131 ,
		_w624_,
		_w627_,
		_w875_
	);
	LUT2 #(
		.INIT('h8)
	) name413 (
		_w874_,
		_w875_,
		_w876_
	);
	LUT2 #(
		.INIT('h7)
	) name414 (
		_w874_,
		_w875_,
		_w877_
	);
	LUT4 #(
		.INIT('hfe00)
	) name415 (
		\P1_IR_reg[0]/NET0131 ,
		\P1_IR_reg[1]/NET0131 ,
		\P1_IR_reg[2]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		_w878_
	);
	LUT2 #(
		.INIT('h9)
	) name416 (
		\P1_IR_reg[3]/NET0131 ,
		_w878_,
		_w879_
	);
	LUT4 #(
		.INIT('ha9a6)
	) name417 (
		\P2_datao_reg[3]/NET0131 ,
		\si[3]_pad ,
		_w542_,
		_w564_,
		_w880_
	);
	LUT4 #(
		.INIT('h10fe)
	) name418 (
		_w537_,
		_w540_,
		_w879_,
		_w880_,
		_w881_
	);
	LUT3 #(
		.INIT('h80)
	) name419 (
		_w874_,
		_w875_,
		_w881_,
		_w882_
	);
	LUT2 #(
		.INIT('h1)
	) name420 (
		_w873_,
		_w882_,
		_w883_
	);
	LUT4 #(
		.INIT('hf53f)
	) name421 (
		\P1_reg1_reg[4]/NET0131 ,
		\P1_reg2_reg[4]/NET0131 ,
		_w624_,
		_w627_,
		_w884_
	);
	LUT2 #(
		.INIT('h6)
	) name422 (
		\P1_reg3_reg[3]/NET0131 ,
		\P1_reg3_reg[4]/NET0131 ,
		_w885_
	);
	LUT4 #(
		.INIT('h3dfd)
	) name423 (
		\P1_reg0_reg[4]/NET0131 ,
		_w624_,
		_w627_,
		_w885_,
		_w886_
	);
	LUT2 #(
		.INIT('h8)
	) name424 (
		_w884_,
		_w886_,
		_w887_
	);
	LUT2 #(
		.INIT('h7)
	) name425 (
		_w884_,
		_w886_,
		_w888_
	);
	LUT3 #(
		.INIT('h39)
	) name426 (
		\P1_IR_reg[31]/NET0131 ,
		\P1_IR_reg[4]/NET0131 ,
		_w500_,
		_w889_
	);
	LUT2 #(
		.INIT('h4)
	) name427 (
		\P2_datao_reg[4]/NET0131 ,
		_w542_,
		_w890_
	);
	LUT2 #(
		.INIT('h6)
	) name428 (
		\P2_datao_reg[4]/NET0131 ,
		\si[4]_pad ,
		_w891_
	);
	LUT4 #(
		.INIT('h0154)
	) name429 (
		_w542_,
		_w565_,
		_w567_,
		_w891_,
		_w892_
	);
	LUT2 #(
		.INIT('h1)
	) name430 (
		_w890_,
		_w892_,
		_w893_
	);
	LUT4 #(
		.INIT('h10fe)
	) name431 (
		_w537_,
		_w540_,
		_w889_,
		_w893_,
		_w894_
	);
	LUT3 #(
		.INIT('h80)
	) name432 (
		_w884_,
		_w886_,
		_w894_,
		_w895_
	);
	LUT3 #(
		.INIT('h01)
	) name433 (
		_w873_,
		_w882_,
		_w895_,
		_w896_
	);
	LUT3 #(
		.INIT('h07)
	) name434 (
		_w884_,
		_w886_,
		_w894_,
		_w897_
	);
	LUT3 #(
		.INIT('h07)
	) name435 (
		_w874_,
		_w875_,
		_w881_,
		_w898_
	);
	LUT3 #(
		.INIT('h23)
	) name436 (
		_w895_,
		_w897_,
		_w898_,
		_w899_
	);
	LUT4 #(
		.INIT('hf53f)
	) name437 (
		\P1_reg1_reg[8]/NET0131 ,
		\P1_reg2_reg[8]/NET0131 ,
		_w624_,
		_w627_,
		_w900_
	);
	LUT3 #(
		.INIT('h6c)
	) name438 (
		\P1_reg3_reg[7]/NET0131 ,
		\P1_reg3_reg[8]/NET0131 ,
		_w630_,
		_w901_
	);
	LUT4 #(
		.INIT('h3dfd)
	) name439 (
		\P1_reg0_reg[8]/NET0131 ,
		_w624_,
		_w627_,
		_w901_,
		_w902_
	);
	LUT2 #(
		.INIT('h8)
	) name440 (
		_w900_,
		_w902_,
		_w903_
	);
	LUT2 #(
		.INIT('h7)
	) name441 (
		_w900_,
		_w902_,
		_w904_
	);
	LUT4 #(
		.INIT('h5956)
	) name442 (
		\P2_datao_reg[8]/NET0131 ,
		\si[8]_pad ,
		_w542_,
		_w686_,
		_w905_
	);
	LUT3 #(
		.INIT('hc6)
	) name443 (
		\P1_IR_reg[31]/NET0131 ,
		\P1_IR_reg[8]/NET0131 ,
		_w839_,
		_w906_
	);
	LUT4 #(
		.INIT('he0f1)
	) name444 (
		_w537_,
		_w540_,
		_w905_,
		_w906_,
		_w907_
	);
	LUT3 #(
		.INIT('h80)
	) name445 (
		_w900_,
		_w902_,
		_w907_,
		_w908_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name446 (
		\P1_reg0_reg[7]/NET0131 ,
		\P1_reg1_reg[7]/NET0131 ,
		_w624_,
		_w627_,
		_w909_
	);
	LUT2 #(
		.INIT('h6)
	) name447 (
		\P1_reg3_reg[7]/NET0131 ,
		_w630_,
		_w910_
	);
	LUT4 #(
		.INIT('h37f7)
	) name448 (
		\P1_reg2_reg[7]/NET0131 ,
		_w624_,
		_w627_,
		_w910_,
		_w911_
	);
	LUT2 #(
		.INIT('h8)
	) name449 (
		_w909_,
		_w911_,
		_w912_
	);
	LUT2 #(
		.INIT('h7)
	) name450 (
		_w909_,
		_w911_,
		_w913_
	);
	LUT4 #(
		.INIT('h5956)
	) name451 (
		\P2_datao_reg[7]/NET0131 ,
		\si[7]_pad ,
		_w542_,
		_w659_,
		_w914_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name452 (
		\P1_IR_reg[31]/NET0131 ,
		\P1_IR_reg[4]/NET0131 ,
		\P1_IR_reg[5]/NET0131 ,
		_w500_,
		_w915_
	);
	LUT2 #(
		.INIT('h8)
	) name453 (
		\P1_IR_reg[31]/NET0131 ,
		\P1_IR_reg[6]/NET0131 ,
		_w916_
	);
	LUT3 #(
		.INIT('h56)
	) name454 (
		\P1_IR_reg[7]/NET0131 ,
		_w915_,
		_w916_,
		_w917_
	);
	LUT4 #(
		.INIT('he0f1)
	) name455 (
		_w537_,
		_w540_,
		_w914_,
		_w917_,
		_w918_
	);
	LUT3 #(
		.INIT('h80)
	) name456 (
		_w909_,
		_w911_,
		_w918_,
		_w919_
	);
	LUT2 #(
		.INIT('h1)
	) name457 (
		_w908_,
		_w919_,
		_w920_
	);
	LUT4 #(
		.INIT('hf53f)
	) name458 (
		\P1_reg1_reg[6]/NET0131 ,
		\P1_reg2_reg[6]/NET0131 ,
		_w624_,
		_w627_,
		_w921_
	);
	LUT4 #(
		.INIT('h7f80)
	) name459 (
		\P1_reg3_reg[3]/NET0131 ,
		\P1_reg3_reg[4]/NET0131 ,
		\P1_reg3_reg[5]/NET0131 ,
		\P1_reg3_reg[6]/NET0131 ,
		_w922_
	);
	LUT4 #(
		.INIT('h3dfd)
	) name460 (
		\P1_reg0_reg[6]/NET0131 ,
		_w624_,
		_w627_,
		_w922_,
		_w923_
	);
	LUT2 #(
		.INIT('h8)
	) name461 (
		_w921_,
		_w923_,
		_w924_
	);
	LUT2 #(
		.INIT('h7)
	) name462 (
		_w921_,
		_w923_,
		_w925_
	);
	LUT2 #(
		.INIT('h9)
	) name463 (
		\P1_IR_reg[6]/NET0131 ,
		_w915_,
		_w926_
	);
	LUT4 #(
		.INIT('h040f)
	) name464 (
		_w565_,
		_w568_,
		_w570_,
		_w684_,
		_w927_
	);
	LUT4 #(
		.INIT('ha9a6)
	) name465 (
		\P2_datao_reg[6]/NET0131 ,
		\si[6]_pad ,
		_w542_,
		_w927_,
		_w928_
	);
	LUT4 #(
		.INIT('h10fe)
	) name466 (
		_w537_,
		_w540_,
		_w926_,
		_w928_,
		_w929_
	);
	LUT3 #(
		.INIT('h80)
	) name467 (
		_w921_,
		_w923_,
		_w929_,
		_w930_
	);
	LUT3 #(
		.INIT('h78)
	) name468 (
		\P1_reg3_reg[3]/NET0131 ,
		\P1_reg3_reg[4]/NET0131 ,
		\P1_reg3_reg[5]/NET0131 ,
		_w931_
	);
	LUT4 #(
		.INIT('h37f7)
	) name469 (
		\P1_reg2_reg[5]/NET0131 ,
		_w624_,
		_w627_,
		_w931_,
		_w932_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name470 (
		\P1_reg0_reg[5]/NET0131 ,
		\P1_reg1_reg[5]/NET0131 ,
		_w624_,
		_w627_,
		_w933_
	);
	LUT2 #(
		.INIT('h8)
	) name471 (
		_w932_,
		_w933_,
		_w934_
	);
	LUT2 #(
		.INIT('h7)
	) name472 (
		_w932_,
		_w933_,
		_w935_
	);
	LUT4 #(
		.INIT('h5956)
	) name473 (
		\P2_datao_reg[5]/NET0131 ,
		\si[5]_pad ,
		_w542_,
		_w569_,
		_w936_
	);
	LUT4 #(
		.INIT('h785a)
	) name474 (
		\P1_IR_reg[31]/NET0131 ,
		\P1_IR_reg[4]/NET0131 ,
		\P1_IR_reg[5]/NET0131 ,
		_w500_,
		_w937_
	);
	LUT4 #(
		.INIT('he0f1)
	) name475 (
		_w537_,
		_w540_,
		_w936_,
		_w937_,
		_w938_
	);
	LUT3 #(
		.INIT('h80)
	) name476 (
		_w932_,
		_w933_,
		_w938_,
		_w939_
	);
	LUT2 #(
		.INIT('h1)
	) name477 (
		_w930_,
		_w939_,
		_w940_
	);
	LUT4 #(
		.INIT('h0001)
	) name478 (
		_w908_,
		_w919_,
		_w930_,
		_w939_,
		_w941_
	);
	LUT4 #(
		.INIT('h4f00)
	) name479 (
		_w872_,
		_w896_,
		_w899_,
		_w941_,
		_w942_
	);
	LUT3 #(
		.INIT('h07)
	) name480 (
		_w921_,
		_w923_,
		_w929_,
		_w943_
	);
	LUT3 #(
		.INIT('h07)
	) name481 (
		_w932_,
		_w933_,
		_w938_,
		_w944_
	);
	LUT3 #(
		.INIT('h23)
	) name482 (
		_w930_,
		_w943_,
		_w944_,
		_w945_
	);
	LUT3 #(
		.INIT('h07)
	) name483 (
		_w900_,
		_w902_,
		_w907_,
		_w946_
	);
	LUT3 #(
		.INIT('h07)
	) name484 (
		_w909_,
		_w911_,
		_w918_,
		_w947_
	);
	LUT3 #(
		.INIT('h23)
	) name485 (
		_w908_,
		_w946_,
		_w947_,
		_w948_
	);
	LUT3 #(
		.INIT('hd0)
	) name486 (
		_w920_,
		_w945_,
		_w948_,
		_w949_
	);
	LUT4 #(
		.INIT('h0008)
	) name487 (
		_w830_,
		_w832_,
		_w838_,
		_w841_,
		_w950_
	);
	LUT2 #(
		.INIT('h1)
	) name488 (
		_w828_,
		_w950_,
		_w951_
	);
	LUT2 #(
		.INIT('h8)
	) name489 (
		_w815_,
		_w951_,
		_w952_
	);
	LUT3 #(
		.INIT('hb0)
	) name490 (
		_w942_,
		_w949_,
		_w952_,
		_w953_
	);
	LUT4 #(
		.INIT('h20aa)
	) name491 (
		_w846_,
		_w942_,
		_w949_,
		_w952_,
		_w954_
	);
	LUT4 #(
		.INIT('hfee0)
	) name492 (
		_w752_,
		_w758_,
		_w762_,
		_w767_,
		_w955_
	);
	LUT4 #(
		.INIT('hfee0)
	) name493 (
		_w772_,
		_w780_,
		_w786_,
		_w791_,
		_w956_
	);
	LUT3 #(
		.INIT('hd0)
	) name494 (
		_w793_,
		_w955_,
		_w956_,
		_w957_
	);
	LUT3 #(
		.INIT('h08)
	) name495 (
		_w709_,
		_w747_,
		_w957_,
		_w958_
	);
	LUT2 #(
		.INIT('h1)
	) name496 (
		_w717_,
		_w722_,
		_w959_
	);
	LUT3 #(
		.INIT('h8e)
	) name497 (
		_w738_,
		_w745_,
		_w959_,
		_w960_
	);
	LUT3 #(
		.INIT('h01)
	) name498 (
		_w541_,
		_w701_,
		_w706_,
		_w961_
	);
	LUT4 #(
		.INIT('h008d)
	) name499 (
		_w541_,
		_w652_,
		_w673_,
		_w679_,
		_w962_
	);
	LUT3 #(
		.INIT('h23)
	) name500 (
		_w708_,
		_w961_,
		_w962_,
		_w963_
	);
	LUT3 #(
		.INIT('hd0)
	) name501 (
		_w709_,
		_w960_,
		_w963_,
		_w964_
	);
	LUT4 #(
		.INIT('h0d00)
	) name502 (
		_w795_,
		_w954_,
		_w958_,
		_w964_,
		_w965_
	);
	LUT4 #(
		.INIT('h4c44)
	) name503 (
		_w598_,
		_w611_,
		_w711_,
		_w712_,
		_w966_
	);
	LUT3 #(
		.INIT('ha2)
	) name504 (
		_w556_,
		_w616_,
		_w966_,
		_w967_
	);
	LUT4 #(
		.INIT('h5956)
	) name505 (
		\P2_datao_reg[25]/NET0131 ,
		\si[25]_pad ,
		_w542_,
		_w967_,
		_w968_
	);
	LUT2 #(
		.INIT('h1)
	) name506 (
		_w541_,
		_w968_,
		_w969_
	);
	LUT3 #(
		.INIT('h80)
	) name507 (
		\P1_reg3_reg[23]/NET0131 ,
		_w634_,
		_w636_,
		_w970_
	);
	LUT4 #(
		.INIT('h8000)
	) name508 (
		\P1_reg3_reg[23]/NET0131 ,
		_w634_,
		_w637_,
		_w636_,
		_w971_
	);
	LUT3 #(
		.INIT('h6c)
	) name509 (
		\P1_reg3_reg[24]/NET0131 ,
		\P1_reg3_reg[25]/NET0131 ,
		_w970_,
		_w972_
	);
	LUT4 #(
		.INIT('h60c0)
	) name510 (
		\P1_reg3_reg[24]/NET0131 ,
		\P1_reg3_reg[25]/NET0131 ,
		_w629_,
		_w970_,
		_w973_
	);
	LUT3 #(
		.INIT('h08)
	) name511 (
		\P1_reg2_reg[25]/NET0131 ,
		_w624_,
		_w627_,
		_w974_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name512 (
		\P1_reg0_reg[25]/NET0131 ,
		\P1_reg1_reg[25]/NET0131 ,
		_w624_,
		_w627_,
		_w975_
	);
	LUT2 #(
		.INIT('h4)
	) name513 (
		_w974_,
		_w975_,
		_w976_
	);
	LUT2 #(
		.INIT('h4)
	) name514 (
		_w973_,
		_w976_,
		_w977_
	);
	LUT2 #(
		.INIT('hb)
	) name515 (
		_w973_,
		_w976_,
		_w978_
	);
	LUT3 #(
		.INIT('he0)
	) name516 (
		_w541_,
		_w968_,
		_w977_,
		_w979_
	);
	LUT2 #(
		.INIT('h8)
	) name517 (
		\P2_datao_reg[26]/NET0131 ,
		_w542_,
		_w980_
	);
	LUT2 #(
		.INIT('h6)
	) name518 (
		\P2_datao_reg[26]/NET0131 ,
		\si[26]_pad ,
		_w981_
	);
	LUT4 #(
		.INIT('hfac8)
	) name519 (
		\P2_datao_reg[20]/NET0131 ,
		\P2_datao_reg[21]/NET0131 ,
		\si[20]_pad ,
		\si[21]_pad ,
		_w982_
	);
	LUT2 #(
		.INIT('h8)
	) name520 (
		_w597_,
		_w982_,
		_w983_
	);
	LUT4 #(
		.INIT('hfac8)
	) name521 (
		\P2_datao_reg[22]/NET0131 ,
		\P2_datao_reg[23]/NET0131 ,
		\si[22]_pad ,
		\si[23]_pad ,
		_w984_
	);
	LUT4 #(
		.INIT('hfac8)
	) name522 (
		\P2_datao_reg[24]/NET0131 ,
		\P2_datao_reg[25]/NET0131 ,
		\si[24]_pad ,
		\si[25]_pad ,
		_w985_
	);
	LUT2 #(
		.INIT('h8)
	) name523 (
		_w984_,
		_w985_,
		_w986_
	);
	LUT4 #(
		.INIT('h8000)
	) name524 (
		_w602_,
		_w654_,
		_w984_,
		_w985_,
		_w987_
	);
	LUT2 #(
		.INIT('h8)
	) name525 (
		_w983_,
		_w987_,
		_w988_
	);
	LUT4 #(
		.INIT('hb000)
	) name526 (
		_w728_,
		_w729_,
		_w730_,
		_w988_,
		_w989_
	);
	LUT4 #(
		.INIT('hec80)
	) name527 (
		\P2_datao_reg[20]/NET0131 ,
		\P2_datao_reg[21]/NET0131 ,
		\si[20]_pad ,
		\si[21]_pad ,
		_w990_
	);
	LUT3 #(
		.INIT('h07)
	) name528 (
		_w697_,
		_w982_,
		_w990_,
		_w991_
	);
	LUT4 #(
		.INIT('h4f00)
	) name529 (
		_w726_,
		_w732_,
		_w733_,
		_w983_,
		_w992_
	);
	LUT4 #(
		.INIT('hec80)
	) name530 (
		\P2_datao_reg[22]/NET0131 ,
		\P2_datao_reg[23]/NET0131 ,
		\si[22]_pad ,
		\si[23]_pad ,
		_w993_
	);
	LUT4 #(
		.INIT('hec80)
	) name531 (
		\P2_datao_reg[24]/NET0131 ,
		\P2_datao_reg[25]/NET0131 ,
		\si[24]_pad ,
		\si[25]_pad ,
		_w994_
	);
	LUT3 #(
		.INIT('h07)
	) name532 (
		_w985_,
		_w993_,
		_w994_,
		_w995_
	);
	LUT4 #(
		.INIT('h5d00)
	) name533 (
		_w986_,
		_w991_,
		_w992_,
		_w995_,
		_w996_
	);
	LUT4 #(
		.INIT('h1411)
	) name534 (
		_w542_,
		_w981_,
		_w989_,
		_w996_,
		_w997_
	);
	LUT3 #(
		.INIT('h54)
	) name535 (
		_w541_,
		_w980_,
		_w997_,
		_w998_
	);
	LUT2 #(
		.INIT('h6)
	) name536 (
		\P1_reg3_reg[26]/NET0131 ,
		_w971_,
		_w999_
	);
	LUT3 #(
		.INIT('h48)
	) name537 (
		\P1_reg3_reg[26]/NET0131 ,
		_w629_,
		_w971_,
		_w1000_
	);
	LUT3 #(
		.INIT('h20)
	) name538 (
		\P1_reg1_reg[26]/NET0131 ,
		_w624_,
		_w627_,
		_w1001_
	);
	LUT4 #(
		.INIT('hff35)
	) name539 (
		\P1_reg0_reg[26]/NET0131 ,
		\P1_reg2_reg[26]/NET0131 ,
		_w624_,
		_w627_,
		_w1002_
	);
	LUT2 #(
		.INIT('h4)
	) name540 (
		_w1001_,
		_w1002_,
		_w1003_
	);
	LUT2 #(
		.INIT('h4)
	) name541 (
		_w1000_,
		_w1003_,
		_w1004_
	);
	LUT2 #(
		.INIT('hb)
	) name542 (
		_w1000_,
		_w1003_,
		_w1005_
	);
	LUT3 #(
		.INIT('h10)
	) name543 (
		_w998_,
		_w1000_,
		_w1003_,
		_w1006_
	);
	LUT4 #(
		.INIT('h001f)
	) name544 (
		_w541_,
		_w968_,
		_w977_,
		_w1006_,
		_w1007_
	);
	LUT2 #(
		.INIT('h8)
	) name545 (
		\P2_datao_reg[28]/NET0131 ,
		_w542_,
		_w1008_
	);
	LUT2 #(
		.INIT('h6)
	) name546 (
		\P2_datao_reg[28]/NET0131 ,
		\si[28]_pad ,
		_w1009_
	);
	LUT2 #(
		.INIT('h8)
	) name547 (
		_w984_,
		_w982_,
		_w1010_
	);
	LUT3 #(
		.INIT('h07)
	) name548 (
		_w984_,
		_w990_,
		_w993_,
		_w1011_
	);
	LUT3 #(
		.INIT('hb0)
	) name549 (
		_w700_,
		_w1010_,
		_w1011_,
		_w1012_
	);
	LUT3 #(
		.INIT('h04)
	) name550 (
		_w548_,
		_w551_,
		_w552_,
		_w1013_
	);
	LUT4 #(
		.INIT('h4f00)
	) name551 (
		_w700_,
		_w1010_,
		_w1011_,
		_w1013_,
		_w1014_
	);
	LUT4 #(
		.INIT('h135f)
	) name552 (
		\P2_datao_reg[26]/NET0131 ,
		\P2_datao_reg[27]/NET0131 ,
		\si[26]_pad ,
		\si[27]_pad ,
		_w1015_
	);
	LUT4 #(
		.INIT('h1055)
	) name553 (
		_w548_,
		_w549_,
		_w994_,
		_w1015_,
		_w1016_
	);
	LUT4 #(
		.INIT('h1114)
	) name554 (
		_w542_,
		_w1009_,
		_w1014_,
		_w1016_,
		_w1017_
	);
	LUT3 #(
		.INIT('h54)
	) name555 (
		_w541_,
		_w1008_,
		_w1017_,
		_w1018_
	);
	LUT4 #(
		.INIT('h870f)
	) name556 (
		\P1_reg3_reg[26]/NET0131 ,
		\P1_reg3_reg[27]/NET0131 ,
		\P1_reg3_reg[28]/NET0131 ,
		_w971_,
		_w1019_
	);
	LUT3 #(
		.INIT('h08)
	) name557 (
		\P1_reg2_reg[28]/NET0131 ,
		_w624_,
		_w627_,
		_w1020_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name558 (
		\P1_reg0_reg[28]/NET0131 ,
		\P1_reg1_reg[28]/NET0131 ,
		_w624_,
		_w627_,
		_w1021_
	);
	LUT2 #(
		.INIT('h4)
	) name559 (
		_w1020_,
		_w1021_,
		_w1022_
	);
	LUT3 #(
		.INIT('hd0)
	) name560 (
		_w629_,
		_w1019_,
		_w1022_,
		_w1023_
	);
	LUT3 #(
		.INIT('h2f)
	) name561 (
		_w629_,
		_w1019_,
		_w1022_,
		_w1024_
	);
	LUT4 #(
		.INIT('hab00)
	) name562 (
		_w541_,
		_w1008_,
		_w1017_,
		_w1023_,
		_w1025_
	);
	LUT3 #(
		.INIT('h15)
	) name563 (
		_w550_,
		_w551_,
		_w555_,
		_w1026_
	);
	LUT2 #(
		.INIT('h8)
	) name564 (
		_w551_,
		_w553_,
		_w1027_
	);
	LUT3 #(
		.INIT('h15)
	) name565 (
		_w554_,
		_w609_,
		_w615_,
		_w1028_
	);
	LUT4 #(
		.INIT('hfac8)
	) name566 (
		\P2_datao_reg[19]/NET0131 ,
		\P2_datao_reg[22]/NET0131 ,
		\si[19]_pad ,
		\si[22]_pad ,
		_w1029_
	);
	LUT2 #(
		.INIT('h8)
	) name567 (
		_w982_,
		_w1029_,
		_w1030_
	);
	LUT4 #(
		.INIT('h8f00)
	) name568 (
		_w655_,
		_w666_,
		_w671_,
		_w1030_,
		_w1031_
	);
	LUT4 #(
		.INIT('h22a2)
	) name569 (
		_w1026_,
		_w1027_,
		_w1028_,
		_w1031_,
		_w1032_
	);
	LUT4 #(
		.INIT('h5956)
	) name570 (
		\P2_datao_reg[27]/NET0131 ,
		\si[27]_pad ,
		_w542_,
		_w1032_,
		_w1033_
	);
	LUT2 #(
		.INIT('h1)
	) name571 (
		_w541_,
		_w1033_,
		_w1034_
	);
	LUT3 #(
		.INIT('h6c)
	) name572 (
		\P1_reg3_reg[26]/NET0131 ,
		\P1_reg3_reg[27]/NET0131 ,
		_w971_,
		_w1035_
	);
	LUT4 #(
		.INIT('h60c0)
	) name573 (
		\P1_reg3_reg[26]/NET0131 ,
		\P1_reg3_reg[27]/NET0131 ,
		_w629_,
		_w971_,
		_w1036_
	);
	LUT3 #(
		.INIT('h20)
	) name574 (
		\P1_reg1_reg[27]/NET0131 ,
		_w624_,
		_w627_,
		_w1037_
	);
	LUT4 #(
		.INIT('hff35)
	) name575 (
		\P1_reg0_reg[27]/NET0131 ,
		\P1_reg2_reg[27]/NET0131 ,
		_w624_,
		_w627_,
		_w1038_
	);
	LUT2 #(
		.INIT('h4)
	) name576 (
		_w1037_,
		_w1038_,
		_w1039_
	);
	LUT2 #(
		.INIT('h4)
	) name577 (
		_w1036_,
		_w1039_,
		_w1040_
	);
	LUT2 #(
		.INIT('hb)
	) name578 (
		_w1036_,
		_w1039_,
		_w1041_
	);
	LUT3 #(
		.INIT('he0)
	) name579 (
		_w541_,
		_w1033_,
		_w1040_,
		_w1042_
	);
	LUT3 #(
		.INIT('h02)
	) name580 (
		_w1007_,
		_w1025_,
		_w1042_,
		_w1043_
	);
	LUT4 #(
		.INIT('h0057)
	) name581 (
		_w655_,
		_w666_,
		_w669_,
		_w670_,
		_w1044_
	);
	LUT3 #(
		.INIT('ha2)
	) name582 (
		_w1028_,
		_w1030_,
		_w1044_,
		_w1045_
	);
	LUT4 #(
		.INIT('h5956)
	) name583 (
		\P2_datao_reg[23]/NET0131 ,
		\si[23]_pad ,
		_w542_,
		_w1045_,
		_w1046_
	);
	LUT2 #(
		.INIT('h1)
	) name584 (
		_w541_,
		_w1046_,
		_w1047_
	);
	LUT3 #(
		.INIT('h6a)
	) name585 (
		\P1_reg3_reg[23]/NET0131 ,
		_w634_,
		_w636_,
		_w1048_
	);
	LUT3 #(
		.INIT('h20)
	) name586 (
		\P1_reg1_reg[23]/NET0131 ,
		_w624_,
		_w627_,
		_w1049_
	);
	LUT4 #(
		.INIT('hff35)
	) name587 (
		\P1_reg0_reg[23]/NET0131 ,
		\P1_reg2_reg[23]/NET0131 ,
		_w624_,
		_w627_,
		_w1050_
	);
	LUT4 #(
		.INIT('h1300)
	) name588 (
		_w629_,
		_w1049_,
		_w1048_,
		_w1050_,
		_w1051_
	);
	LUT4 #(
		.INIT('hecff)
	) name589 (
		_w629_,
		_w1049_,
		_w1048_,
		_w1050_,
		_w1052_
	);
	LUT3 #(
		.INIT('he0)
	) name590 (
		_w541_,
		_w1046_,
		_w1051_,
		_w1053_
	);
	LUT4 #(
		.INIT('h5956)
	) name591 (
		\P2_datao_reg[24]/NET0131 ,
		\si[24]_pad ,
		_w542_,
		_w1012_,
		_w1054_
	);
	LUT2 #(
		.INIT('h1)
	) name592 (
		_w541_,
		_w1054_,
		_w1055_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name593 (
		\P1_reg3_reg[23]/NET0131 ,
		\P1_reg3_reg[24]/NET0131 ,
		_w634_,
		_w636_,
		_w1056_
	);
	LUT3 #(
		.INIT('h02)
	) name594 (
		\P1_reg0_reg[24]/NET0131 ,
		_w624_,
		_w627_,
		_w1057_
	);
	LUT4 #(
		.INIT('hf53f)
	) name595 (
		\P1_reg1_reg[24]/NET0131 ,
		\P1_reg2_reg[24]/NET0131 ,
		_w624_,
		_w627_,
		_w1058_
	);
	LUT4 #(
		.INIT('h1300)
	) name596 (
		_w629_,
		_w1057_,
		_w1056_,
		_w1058_,
		_w1059_
	);
	LUT4 #(
		.INIT('hecff)
	) name597 (
		_w629_,
		_w1057_,
		_w1056_,
		_w1058_,
		_w1060_
	);
	LUT3 #(
		.INIT('he0)
	) name598 (
		_w541_,
		_w1054_,
		_w1059_,
		_w1061_
	);
	LUT2 #(
		.INIT('h8)
	) name599 (
		\P2_datao_reg[22]/NET0131 ,
		_w542_,
		_w1062_
	);
	LUT2 #(
		.INIT('h6)
	) name600 (
		\P2_datao_reg[22]/NET0131 ,
		\si[22]_pad ,
		_w1063_
	);
	LUT4 #(
		.INIT('h4f00)
	) name601 (
		_w731_,
		_w732_,
		_w733_,
		_w983_,
		_w1064_
	);
	LUT4 #(
		.INIT('h0541)
	) name602 (
		_w542_,
		_w991_,
		_w1063_,
		_w1064_,
		_w1065_
	);
	LUT3 #(
		.INIT('h54)
	) name603 (
		_w541_,
		_w1062_,
		_w1065_,
		_w1066_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name604 (
		\P1_reg3_reg[21]/NET0131 ,
		\P1_reg3_reg[22]/NET0131 ,
		_w634_,
		_w635_,
		_w1067_
	);
	LUT3 #(
		.INIT('h20)
	) name605 (
		\P1_reg1_reg[22]/NET0131 ,
		_w624_,
		_w627_,
		_w1068_
	);
	LUT4 #(
		.INIT('hff35)
	) name606 (
		\P1_reg0_reg[22]/NET0131 ,
		\P1_reg2_reg[22]/NET0131 ,
		_w624_,
		_w627_,
		_w1069_
	);
	LUT4 #(
		.INIT('h1300)
	) name607 (
		_w629_,
		_w1068_,
		_w1067_,
		_w1069_,
		_w1070_
	);
	LUT4 #(
		.INIT('hecff)
	) name608 (
		_w629_,
		_w1068_,
		_w1067_,
		_w1069_,
		_w1071_
	);
	LUT4 #(
		.INIT('hab00)
	) name609 (
		_w541_,
		_w1062_,
		_w1065_,
		_w1070_,
		_w1072_
	);
	LUT4 #(
		.INIT('h5956)
	) name610 (
		\P2_datao_reg[21]/NET0131 ,
		\si[21]_pad ,
		_w542_,
		_w613_,
		_w1073_
	);
	LUT2 #(
		.INIT('h1)
	) name611 (
		_w541_,
		_w1073_,
		_w1074_
	);
	LUT3 #(
		.INIT('h6a)
	) name612 (
		\P1_reg3_reg[21]/NET0131 ,
		_w634_,
		_w635_,
		_w1075_
	);
	LUT3 #(
		.INIT('h08)
	) name613 (
		\P1_reg2_reg[21]/NET0131 ,
		_w624_,
		_w627_,
		_w1076_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name614 (
		\P1_reg0_reg[21]/NET0131 ,
		\P1_reg1_reg[21]/NET0131 ,
		_w624_,
		_w627_,
		_w1077_
	);
	LUT4 #(
		.INIT('h1300)
	) name615 (
		_w629_,
		_w1076_,
		_w1075_,
		_w1077_,
		_w1078_
	);
	LUT4 #(
		.INIT('hecff)
	) name616 (
		_w629_,
		_w1076_,
		_w1075_,
		_w1077_,
		_w1079_
	);
	LUT3 #(
		.INIT('he0)
	) name617 (
		_w541_,
		_w1073_,
		_w1078_,
		_w1080_
	);
	LUT2 #(
		.INIT('h1)
	) name618 (
		_w1072_,
		_w1080_,
		_w1081_
	);
	LUT3 #(
		.INIT('h10)
	) name619 (
		_w1053_,
		_w1061_,
		_w1081_,
		_w1082_
	);
	LUT2 #(
		.INIT('h8)
	) name620 (
		_w1043_,
		_w1082_,
		_w1083_
	);
	LUT4 #(
		.INIT('h0054)
	) name621 (
		_w541_,
		_w1062_,
		_w1065_,
		_w1070_,
		_w1084_
	);
	LUT3 #(
		.INIT('h01)
	) name622 (
		_w541_,
		_w1073_,
		_w1078_,
		_w1085_
	);
	LUT3 #(
		.INIT('h23)
	) name623 (
		_w1072_,
		_w1084_,
		_w1085_,
		_w1086_
	);
	LUT3 #(
		.INIT('h01)
	) name624 (
		_w1053_,
		_w1061_,
		_w1086_,
		_w1087_
	);
	LUT3 #(
		.INIT('h01)
	) name625 (
		_w541_,
		_w1054_,
		_w1059_,
		_w1088_
	);
	LUT3 #(
		.INIT('h01)
	) name626 (
		_w541_,
		_w1046_,
		_w1051_,
		_w1089_
	);
	LUT3 #(
		.INIT('h23)
	) name627 (
		_w1061_,
		_w1088_,
		_w1089_,
		_w1090_
	);
	LUT2 #(
		.INIT('h4)
	) name628 (
		_w1087_,
		_w1090_,
		_w1091_
	);
	LUT3 #(
		.INIT('h8a)
	) name629 (
		_w1043_,
		_w1087_,
		_w1090_,
		_w1092_
	);
	LUT3 #(
		.INIT('h8a)
	) name630 (
		_w998_,
		_w1000_,
		_w1003_,
		_w1093_
	);
	LUT3 #(
		.INIT('h01)
	) name631 (
		_w541_,
		_w968_,
		_w977_,
		_w1094_
	);
	LUT4 #(
		.INIT('h0001)
	) name632 (
		_w541_,
		_w968_,
		_w977_,
		_w1006_,
		_w1095_
	);
	LUT2 #(
		.INIT('h1)
	) name633 (
		_w1093_,
		_w1095_,
		_w1096_
	);
	LUT4 #(
		.INIT('h1110)
	) name634 (
		_w1025_,
		_w1042_,
		_w1093_,
		_w1095_,
		_w1097_
	);
	LUT4 #(
		.INIT('h0054)
	) name635 (
		_w541_,
		_w1008_,
		_w1017_,
		_w1023_,
		_w1098_
	);
	LUT3 #(
		.INIT('h01)
	) name636 (
		_w541_,
		_w1033_,
		_w1040_,
		_w1099_
	);
	LUT3 #(
		.INIT('h23)
	) name637 (
		_w1025_,
		_w1098_,
		_w1099_,
		_w1100_
	);
	LUT2 #(
		.INIT('h4)
	) name638 (
		_w1097_,
		_w1100_,
		_w1101_
	);
	LUT4 #(
		.INIT('h0b00)
	) name639 (
		_w965_,
		_w1083_,
		_w1092_,
		_w1101_,
		_w1102_
	);
	LUT4 #(
		.INIT('hd11d)
	) name640 (
		\P1_reg2_reg[29]/NET0131 ,
		_w534_,
		_w647_,
		_w1102_,
		_w1103_
	);
	LUT2 #(
		.INIT('h6)
	) name641 (
		\P1_IR_reg[22]/NET0131 ,
		_w513_,
		_w1104_
	);
	LUT4 #(
		.INIT('h1000)
	) name642 (
		\P1_IR_reg[16]/NET0131 ,
		\P1_IR_reg[17]/NET0131 ,
		_w506_,
		_w648_,
		_w1105_
	);
	LUT4 #(
		.INIT('h6c3c)
	) name643 (
		\P1_IR_reg[20]/NET0131 ,
		\P1_IR_reg[21]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		_w1105_,
		_w1106_
	);
	LUT2 #(
		.INIT('h1)
	) name644 (
		_w1104_,
		_w1106_,
		_w1107_
	);
	LUT2 #(
		.INIT('h8)
	) name645 (
		_w1104_,
		_w1106_,
		_w1108_
	);
	LUT2 #(
		.INIT('h6)
	) name646 (
		_w1104_,
		_w1106_,
		_w1109_
	);
	LUT4 #(
		.INIT('h5600)
	) name647 (
		\P1_IR_reg[19]/NET0131 ,
		_w650_,
		_w651_,
		_w1104_,
		_w1110_
	);
	LUT3 #(
		.INIT('h59)
	) name648 (
		\P1_IR_reg[20]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		_w1105_,
		_w1111_
	);
	LUT4 #(
		.INIT('h2818)
	) name649 (
		\P1_IR_reg[20]/NET0131 ,
		\P1_IR_reg[21]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		_w1105_,
		_w1112_
	);
	LUT2 #(
		.INIT('h1)
	) name650 (
		_w1110_,
		_w1112_,
		_w1113_
	);
	LUT4 #(
		.INIT('h0034)
	) name651 (
		_w652_,
		_w1104_,
		_w1106_,
		_w1112_,
		_w1114_
	);
	LUT4 #(
		.INIT('h8000)
	) name652 (
		_w853_,
		_w861_,
		_w869_,
		_w881_,
		_w1115_
	);
	LUT3 #(
		.INIT('h80)
	) name653 (
		_w918_,
		_w929_,
		_w938_,
		_w1116_
	);
	LUT3 #(
		.INIT('h80)
	) name654 (
		_w894_,
		_w1115_,
		_w1116_,
		_w1117_
	);
	LUT4 #(
		.INIT('h0001)
	) name655 (
		_w824_,
		_w826_,
		_w838_,
		_w841_,
		_w1118_
	);
	LUT2 #(
		.INIT('h8)
	) name656 (
		_w907_,
		_w1118_,
		_w1119_
	);
	LUT4 #(
		.INIT('h8000)
	) name657 (
		_w804_,
		_w814_,
		_w1117_,
		_w1119_,
		_w1120_
	);
	LUT2 #(
		.INIT('h8)
	) name658 (
		_w758_,
		_w767_,
		_w1121_
	);
	LUT3 #(
		.INIT('h80)
	) name659 (
		_w758_,
		_w767_,
		_w780_,
		_w1122_
	);
	LUT4 #(
		.INIT('h40c8)
	) name660 (
		_w541_,
		_w717_,
		_w735_,
		_w736_,
		_w1123_
	);
	LUT4 #(
		.INIT('h7200)
	) name661 (
		_w541_,
		_w652_,
		_w673_,
		_w786_,
		_w1124_
	);
	LUT3 #(
		.INIT('h40)
	) name662 (
		_w702_,
		_w1123_,
		_w1124_,
		_w1125_
	);
	LUT4 #(
		.INIT('habaa)
	) name663 (
		_w541_,
		_w1062_,
		_w1065_,
		_w1073_,
		_w1126_
	);
	LUT3 #(
		.INIT('he0)
	) name664 (
		_w541_,
		_w1046_,
		_w1126_,
		_w1127_
	);
	LUT4 #(
		.INIT('h8000)
	) name665 (
		_w1120_,
		_w1122_,
		_w1125_,
		_w1127_,
		_w1128_
	);
	LUT3 #(
		.INIT('hea)
	) name666 (
		_w541_,
		_w968_,
		_w1054_,
		_w1129_
	);
	LUT3 #(
		.INIT('h32)
	) name667 (
		_w541_,
		_w998_,
		_w1033_,
		_w1130_
	);
	LUT2 #(
		.INIT('h8)
	) name668 (
		_w1129_,
		_w1130_,
		_w1131_
	);
	LUT2 #(
		.INIT('h8)
	) name669 (
		_w1128_,
		_w1131_,
		_w1132_
	);
	LUT4 #(
		.INIT('h1000)
	) name670 (
		_w621_,
		_w1018_,
		_w1128_,
		_w1131_,
		_w1133_
	);
	LUT4 #(
		.INIT('h6555)
	) name671 (
		_w621_,
		_w1018_,
		_w1128_,
		_w1131_,
		_w1134_
	);
	LUT3 #(
		.INIT('h10)
	) name672 (
		_w1104_,
		_w1106_,
		_w1111_,
		_w1135_
	);
	LUT4 #(
		.INIT('h0100)
	) name673 (
		_w652_,
		_w1104_,
		_w1106_,
		_w1111_,
		_w1136_
	);
	LUT4 #(
		.INIT('he200)
	) name674 (
		\P1_reg2_reg[29]/NET0131 ,
		_w534_,
		_w1134_,
		_w1136_,
		_w1137_
	);
	LUT3 #(
		.INIT('h01)
	) name675 (
		_w1104_,
		_w1106_,
		_w1111_,
		_w1138_
	);
	LUT4 #(
		.INIT('h5400)
	) name676 (
		_w541_,
		_w543_,
		_w620_,
		_w1138_,
		_w1139_
	);
	LUT2 #(
		.INIT('h4)
	) name677 (
		_w652_,
		_w1111_,
		_w1140_
	);
	LUT4 #(
		.INIT('h80c0)
	) name678 (
		_w652_,
		_w1104_,
		_w1106_,
		_w1111_,
		_w1141_
	);
	LUT4 #(
		.INIT('haa20)
	) name679 (
		\P1_reg2_reg[29]/NET0131 ,
		_w534_,
		_w1138_,
		_w1141_,
		_w1142_
	);
	LUT4 #(
		.INIT('h0200)
	) name680 (
		_w652_,
		_w1104_,
		_w1106_,
		_w1111_,
		_w1143_
	);
	LUT2 #(
		.INIT('h8)
	) name681 (
		_w640_,
		_w1143_,
		_w1144_
	);
	LUT4 #(
		.INIT('h0007)
	) name682 (
		_w534_,
		_w1139_,
		_w1142_,
		_w1144_,
		_w1145_
	);
	LUT2 #(
		.INIT('h4)
	) name683 (
		_w1137_,
		_w1145_,
		_w1146_
	);
	LUT3 #(
		.INIT('hb0)
	) name684 (
		_w1103_,
		_w1114_,
		_w1146_,
		_w1147_
	);
	LUT4 #(
		.INIT('h08aa)
	) name685 (
		_w537_,
		_w629_,
		_w1019_,
		_w1022_,
		_w1148_
	);
	LUT3 #(
		.INIT('h08)
	) name686 (
		\P1_reg2_reg[31]/NET0131 ,
		_w624_,
		_w627_,
		_w1149_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name687 (
		\P1_reg0_reg[31]/NET0131 ,
		\P1_reg1_reg[31]/NET0131 ,
		_w624_,
		_w627_,
		_w1150_
	);
	LUT3 #(
		.INIT('h10)
	) name688 (
		_w641_,
		_w1149_,
		_w1150_,
		_w1151_
	);
	LUT3 #(
		.INIT('hef)
	) name689 (
		_w641_,
		_w1149_,
		_w1150_,
		_w1152_
	);
	LUT4 #(
		.INIT('h0001)
	) name690 (
		_w849_,
		_w857_,
		_w866_,
		_w1151_,
		_w1153_
	);
	LUT4 #(
		.INIT('h0100)
	) name691 (
		_w876_,
		_w887_,
		_w934_,
		_w1153_,
		_w1154_
	);
	LUT4 #(
		.INIT('h0777)
	) name692 (
		_w817_,
		_w818_,
		_w830_,
		_w832_,
		_w1155_
	);
	LUT4 #(
		.INIT('h0777)
	) name693 (
		_w900_,
		_w902_,
		_w909_,
		_w911_,
		_w1156_
	);
	LUT2 #(
		.INIT('h8)
	) name694 (
		_w1155_,
		_w1156_,
		_w1157_
	);
	LUT3 #(
		.INIT('h40)
	) name695 (
		_w924_,
		_w1154_,
		_w1157_,
		_w1158_
	);
	LUT4 #(
		.INIT('h0777)
	) name696 (
		_w750_,
		_w751_,
		_w797_,
		_w798_,
		_w1159_
	);
	LUT2 #(
		.INIT('h4)
	) name697 (
		_w808_,
		_w1159_,
		_w1160_
	);
	LUT4 #(
		.INIT('h4000)
	) name698 (
		_w924_,
		_w1154_,
		_w1157_,
		_w1160_,
		_w1161_
	);
	LUT4 #(
		.INIT('h0777)
	) name699 (
		_w759_,
		_w761_,
		_w769_,
		_w771_,
		_w1162_
	);
	LUT3 #(
		.INIT('h10)
	) name700 (
		_w722_,
		_w791_,
		_w1162_,
		_w1163_
	);
	LUT2 #(
		.INIT('h8)
	) name701 (
		_w1161_,
		_w1163_,
		_w1164_
	);
	LUT3 #(
		.INIT('h45)
	) name702 (
		_w679_,
		_w741_,
		_w744_,
		_w1165_
	);
	LUT2 #(
		.INIT('h1)
	) name703 (
		_w706_,
		_w1078_,
		_w1166_
	);
	LUT3 #(
		.INIT('h01)
	) name704 (
		_w706_,
		_w1070_,
		_w1078_,
		_w1167_
	);
	LUT4 #(
		.INIT('h0001)
	) name705 (
		_w706_,
		_w1051_,
		_w1070_,
		_w1078_,
		_w1168_
	);
	LUT2 #(
		.INIT('h8)
	) name706 (
		_w1165_,
		_w1168_,
		_w1169_
	);
	LUT3 #(
		.INIT('h40)
	) name707 (
		_w1059_,
		_w1165_,
		_w1168_,
		_w1170_
	);
	LUT4 #(
		.INIT('h1000)
	) name708 (
		_w977_,
		_w1059_,
		_w1165_,
		_w1168_,
		_w1171_
	);
	LUT3 #(
		.INIT('h80)
	) name709 (
		_w1161_,
		_w1163_,
		_w1171_,
		_w1172_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name710 (
		_w1000_,
		_w1003_,
		_w1036_,
		_w1039_,
		_w1173_
	);
	LUT2 #(
		.INIT('h4)
	) name711 (
		_w1023_,
		_w1173_,
		_w1174_
	);
	LUT3 #(
		.INIT('h10)
	) name712 (
		_w643_,
		_w1023_,
		_w1173_,
		_w1175_
	);
	LUT4 #(
		.INIT('h8000)
	) name713 (
		_w1161_,
		_w1163_,
		_w1171_,
		_w1175_,
		_w1176_
	);
	LUT3 #(
		.INIT('h02)
	) name714 (
		\P1_reg0_reg[30]/NET0131 ,
		_w624_,
		_w627_,
		_w1177_
	);
	LUT4 #(
		.INIT('hf53f)
	) name715 (
		\P1_reg1_reg[30]/NET0131 ,
		\P1_reg2_reg[30]/NET0131 ,
		_w624_,
		_w627_,
		_w1178_
	);
	LUT3 #(
		.INIT('h10)
	) name716 (
		_w641_,
		_w1177_,
		_w1178_,
		_w1179_
	);
	LUT3 #(
		.INIT('hef)
	) name717 (
		_w641_,
		_w1177_,
		_w1178_,
		_w1180_
	);
	LUT3 #(
		.INIT('h13)
	) name718 (
		\P1_B_reg/NET0131 ,
		_w537_,
		_w540_,
		_w1181_
	);
	LUT4 #(
		.INIT('h1455)
	) name719 (
		_w1148_,
		_w1176_,
		_w1179_,
		_w1181_,
		_w1182_
	);
	LUT4 #(
		.INIT('h4000)
	) name720 (
		_w652_,
		_w1104_,
		_w1106_,
		_w1111_,
		_w1183_
	);
	LUT4 #(
		.INIT('h2e00)
	) name721 (
		\P1_reg2_reg[29]/NET0131 ,
		_w534_,
		_w1182_,
		_w1183_,
		_w1184_
	);
	LUT3 #(
		.INIT('h10)
	) name722 (
		_w541_,
		_w701_,
		_w706_,
		_w1185_
	);
	LUT4 #(
		.INIT('h8d00)
	) name723 (
		_w541_,
		_w652_,
		_w673_,
		_w679_,
		_w1186_
	);
	LUT2 #(
		.INIT('h1)
	) name724 (
		_w1185_,
		_w1186_,
		_w1187_
	);
	LUT2 #(
		.INIT('h4)
	) name725 (
		_w717_,
		_w722_,
		_w1188_
	);
	LUT3 #(
		.INIT('h0b)
	) name726 (
		_w738_,
		_w745_,
		_w1188_,
		_w1189_
	);
	LUT2 #(
		.INIT('h8)
	) name727 (
		_w1187_,
		_w1189_,
		_w1190_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name728 (
		_w772_,
		_w780_,
		_w786_,
		_w791_,
		_w1191_
	);
	LUT4 #(
		.INIT('hdd0d)
	) name729 (
		_w752_,
		_w758_,
		_w762_,
		_w767_,
		_w1192_
	);
	LUT2 #(
		.INIT('h8)
	) name730 (
		_w1191_,
		_w1192_,
		_w1193_
	);
	LUT3 #(
		.INIT('h80)
	) name731 (
		_w1187_,
		_w1189_,
		_w1193_,
		_w1194_
	);
	LUT4 #(
		.INIT('hdd0d)
	) name732 (
		_w799_,
		_w804_,
		_w808_,
		_w814_,
		_w1195_
	);
	LUT4 #(
		.INIT('h8880)
	) name733 (
		_w817_,
		_w818_,
		_w824_,
		_w826_,
		_w1196_
	);
	LUT4 #(
		.INIT('h0007)
	) name734 (
		_w817_,
		_w818_,
		_w824_,
		_w826_,
		_w1197_
	);
	LUT4 #(
		.INIT('h0007)
	) name735 (
		_w830_,
		_w832_,
		_w838_,
		_w841_,
		_w1198_
	);
	LUT3 #(
		.INIT('h54)
	) name736 (
		_w1196_,
		_w1197_,
		_w1198_,
		_w1199_
	);
	LUT2 #(
		.INIT('h4)
	) name737 (
		_w799_,
		_w804_,
		_w1200_
	);
	LUT4 #(
		.INIT('h4f04)
	) name738 (
		_w799_,
		_w804_,
		_w808_,
		_w814_,
		_w1201_
	);
	LUT3 #(
		.INIT('h07)
	) name739 (
		_w1195_,
		_w1199_,
		_w1201_,
		_w1202_
	);
	LUT3 #(
		.INIT('h08)
	) name740 (
		_w909_,
		_w911_,
		_w918_,
		_w1203_
	);
	LUT3 #(
		.INIT('h08)
	) name741 (
		_w900_,
		_w902_,
		_w907_,
		_w1204_
	);
	LUT2 #(
		.INIT('h1)
	) name742 (
		_w1203_,
		_w1204_,
		_w1205_
	);
	LUT3 #(
		.INIT('h08)
	) name743 (
		_w864_,
		_w865_,
		_w869_,
		_w1206_
	);
	LUT3 #(
		.INIT('h08)
	) name744 (
		_w855_,
		_w856_,
		_w861_,
		_w1207_
	);
	LUT3 #(
		.INIT('h70)
	) name745 (
		_w855_,
		_w856_,
		_w861_,
		_w1208_
	);
	LUT3 #(
		.INIT('h70)
	) name746 (
		_w847_,
		_w848_,
		_w853_,
		_w1209_
	);
	LUT4 #(
		.INIT('h00b2)
	) name747 (
		_w857_,
		_w861_,
		_w1206_,
		_w1209_,
		_w1210_
	);
	LUT3 #(
		.INIT('h08)
	) name748 (
		_w884_,
		_w886_,
		_w894_,
		_w1211_
	);
	LUT3 #(
		.INIT('h08)
	) name749 (
		_w874_,
		_w875_,
		_w881_,
		_w1212_
	);
	LUT3 #(
		.INIT('h08)
	) name750 (
		_w847_,
		_w848_,
		_w853_,
		_w1213_
	);
	LUT2 #(
		.INIT('h1)
	) name751 (
		_w1212_,
		_w1213_,
		_w1214_
	);
	LUT3 #(
		.INIT('h01)
	) name752 (
		_w1211_,
		_w1212_,
		_w1213_,
		_w1215_
	);
	LUT3 #(
		.INIT('h70)
	) name753 (
		_w884_,
		_w886_,
		_w894_,
		_w1216_
	);
	LUT3 #(
		.INIT('h70)
	) name754 (
		_w874_,
		_w875_,
		_w881_,
		_w1217_
	);
	LUT2 #(
		.INIT('h1)
	) name755 (
		_w1216_,
		_w1217_,
		_w1218_
	);
	LUT3 #(
		.INIT('h54)
	) name756 (
		_w1211_,
		_w1216_,
		_w1217_,
		_w1219_
	);
	LUT3 #(
		.INIT('h0b)
	) name757 (
		_w1210_,
		_w1215_,
		_w1219_,
		_w1220_
	);
	LUT3 #(
		.INIT('h08)
	) name758 (
		_w921_,
		_w923_,
		_w929_,
		_w1221_
	);
	LUT3 #(
		.INIT('h08)
	) name759 (
		_w932_,
		_w933_,
		_w938_,
		_w1222_
	);
	LUT2 #(
		.INIT('h1)
	) name760 (
		_w1221_,
		_w1222_,
		_w1223_
	);
	LUT4 #(
		.INIT('hf400)
	) name761 (
		_w1210_,
		_w1215_,
		_w1219_,
		_w1223_,
		_w1224_
	);
	LUT3 #(
		.INIT('h70)
	) name762 (
		_w921_,
		_w923_,
		_w929_,
		_w1225_
	);
	LUT3 #(
		.INIT('h70)
	) name763 (
		_w932_,
		_w933_,
		_w938_,
		_w1226_
	);
	LUT2 #(
		.INIT('h1)
	) name764 (
		_w1225_,
		_w1226_,
		_w1227_
	);
	LUT3 #(
		.INIT('h54)
	) name765 (
		_w1221_,
		_w1225_,
		_w1226_,
		_w1228_
	);
	LUT3 #(
		.INIT('h70)
	) name766 (
		_w900_,
		_w902_,
		_w907_,
		_w1229_
	);
	LUT3 #(
		.INIT('h70)
	) name767 (
		_w909_,
		_w911_,
		_w918_,
		_w1230_
	);
	LUT3 #(
		.INIT('h23)
	) name768 (
		_w1204_,
		_w1229_,
		_w1230_,
		_w1231_
	);
	LUT3 #(
		.INIT('h70)
	) name769 (
		_w1205_,
		_w1228_,
		_w1231_,
		_w1232_
	);
	LUT3 #(
		.INIT('h70)
	) name770 (
		_w1205_,
		_w1224_,
		_w1232_,
		_w1233_
	);
	LUT4 #(
		.INIT('h8880)
	) name771 (
		_w830_,
		_w832_,
		_w838_,
		_w841_,
		_w1234_
	);
	LUT2 #(
		.INIT('h1)
	) name772 (
		_w1196_,
		_w1234_,
		_w1235_
	);
	LUT2 #(
		.INIT('h8)
	) name773 (
		_w1195_,
		_w1235_,
		_w1236_
	);
	LUT4 #(
		.INIT('h8f00)
	) name774 (
		_w1205_,
		_w1224_,
		_w1232_,
		_w1236_,
		_w1237_
	);
	LUT3 #(
		.INIT('ha2)
	) name775 (
		_w1194_,
		_w1202_,
		_w1237_,
		_w1238_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name776 (
		_w752_,
		_w758_,
		_w762_,
		_w767_,
		_w1239_
	);
	LUT4 #(
		.INIT('h4f04)
	) name777 (
		_w752_,
		_w758_,
		_w762_,
		_w767_,
		_w1240_
	);
	LUT2 #(
		.INIT('h4)
	) name778 (
		_w772_,
		_w780_,
		_w1241_
	);
	LUT4 #(
		.INIT('hbf0b)
	) name779 (
		_w772_,
		_w780_,
		_w786_,
		_w791_,
		_w1242_
	);
	LUT3 #(
		.INIT('h70)
	) name780 (
		_w1191_,
		_w1240_,
		_w1242_,
		_w1243_
	);
	LUT3 #(
		.INIT('h08)
	) name781 (
		_w1187_,
		_w1189_,
		_w1243_,
		_w1244_
	);
	LUT2 #(
		.INIT('h2)
	) name782 (
		_w717_,
		_w722_,
		_w1245_
	);
	LUT3 #(
		.INIT('hb2)
	) name783 (
		_w738_,
		_w745_,
		_w1245_,
		_w1246_
	);
	LUT3 #(
		.INIT('h0e)
	) name784 (
		_w541_,
		_w701_,
		_w706_,
		_w1247_
	);
	LUT4 #(
		.INIT('h0072)
	) name785 (
		_w541_,
		_w652_,
		_w673_,
		_w679_,
		_w1248_
	);
	LUT3 #(
		.INIT('h54)
	) name786 (
		_w1185_,
		_w1247_,
		_w1248_,
		_w1249_
	);
	LUT3 #(
		.INIT('h07)
	) name787 (
		_w1187_,
		_w1246_,
		_w1249_,
		_w1250_
	);
	LUT2 #(
		.INIT('h4)
	) name788 (
		_w1244_,
		_w1250_,
		_w1251_
	);
	LUT3 #(
		.INIT('h10)
	) name789 (
		_w541_,
		_w1073_,
		_w1078_,
		_w1252_
	);
	LUT4 #(
		.INIT('h5400)
	) name790 (
		_w541_,
		_w1062_,
		_w1065_,
		_w1070_,
		_w1253_
	);
	LUT2 #(
		.INIT('h1)
	) name791 (
		_w1252_,
		_w1253_,
		_w1254_
	);
	LUT3 #(
		.INIT('h10)
	) name792 (
		_w541_,
		_w1046_,
		_w1051_,
		_w1255_
	);
	LUT3 #(
		.INIT('h10)
	) name793 (
		_w541_,
		_w1054_,
		_w1059_,
		_w1256_
	);
	LUT3 #(
		.INIT('h02)
	) name794 (
		_w1254_,
		_w1255_,
		_w1256_,
		_w1257_
	);
	LUT4 #(
		.INIT('h5400)
	) name795 (
		_w541_,
		_w1008_,
		_w1017_,
		_w1023_,
		_w1258_
	);
	LUT3 #(
		.INIT('h20)
	) name796 (
		_w998_,
		_w1000_,
		_w1003_,
		_w1259_
	);
	LUT3 #(
		.INIT('h10)
	) name797 (
		_w541_,
		_w1033_,
		_w1040_,
		_w1260_
	);
	LUT4 #(
		.INIT('h00ef)
	) name798 (
		_w541_,
		_w1033_,
		_w1040_,
		_w1259_,
		_w1261_
	);
	LUT3 #(
		.INIT('h10)
	) name799 (
		_w541_,
		_w968_,
		_w977_,
		_w1262_
	);
	LUT3 #(
		.INIT('h02)
	) name800 (
		_w1261_,
		_w1258_,
		_w1262_,
		_w1263_
	);
	LUT2 #(
		.INIT('h8)
	) name801 (
		_w1257_,
		_w1263_,
		_w1264_
	);
	LUT3 #(
		.INIT('hb0)
	) name802 (
		_w1238_,
		_w1251_,
		_w1264_,
		_w1265_
	);
	LUT4 #(
		.INIT('h00ab)
	) name803 (
		_w541_,
		_w1062_,
		_w1065_,
		_w1070_,
		_w1266_
	);
	LUT3 #(
		.INIT('h0e)
	) name804 (
		_w541_,
		_w1073_,
		_w1078_,
		_w1267_
	);
	LUT3 #(
		.INIT('h54)
	) name805 (
		_w1253_,
		_w1266_,
		_w1267_,
		_w1268_
	);
	LUT3 #(
		.INIT('h10)
	) name806 (
		_w1255_,
		_w1256_,
		_w1268_,
		_w1269_
	);
	LUT3 #(
		.INIT('h0e)
	) name807 (
		_w541_,
		_w1054_,
		_w1059_,
		_w1270_
	);
	LUT3 #(
		.INIT('h0e)
	) name808 (
		_w541_,
		_w1046_,
		_w1051_,
		_w1271_
	);
	LUT3 #(
		.INIT('h54)
	) name809 (
		_w1256_,
		_w1270_,
		_w1271_,
		_w1272_
	);
	LUT2 #(
		.INIT('h1)
	) name810 (
		_w1269_,
		_w1272_,
		_w1273_
	);
	LUT3 #(
		.INIT('ha8)
	) name811 (
		_w1263_,
		_w1269_,
		_w1272_,
		_w1274_
	);
	LUT4 #(
		.INIT('h00ab)
	) name812 (
		_w541_,
		_w1008_,
		_w1017_,
		_w1023_,
		_w1275_
	);
	LUT3 #(
		.INIT('h0e)
	) name813 (
		_w541_,
		_w1033_,
		_w1040_,
		_w1276_
	);
	LUT2 #(
		.INIT('h1)
	) name814 (
		_w1275_,
		_w1276_,
		_w1277_
	);
	LUT3 #(
		.INIT('h45)
	) name815 (
		_w998_,
		_w1000_,
		_w1003_,
		_w1278_
	);
	LUT3 #(
		.INIT('h0e)
	) name816 (
		_w541_,
		_w968_,
		_w977_,
		_w1279_
	);
	LUT4 #(
		.INIT('h00f1)
	) name817 (
		_w541_,
		_w968_,
		_w977_,
		_w1278_,
		_w1280_
	);
	LUT2 #(
		.INIT('h1)
	) name818 (
		_w1259_,
		_w1280_,
		_w1281_
	);
	LUT3 #(
		.INIT('h01)
	) name819 (
		_w1259_,
		_w1260_,
		_w1280_,
		_w1282_
	);
	LUT3 #(
		.INIT('h51)
	) name820 (
		_w1258_,
		_w1277_,
		_w1282_,
		_w1283_
	);
	LUT2 #(
		.INIT('h1)
	) name821 (
		_w1274_,
		_w1283_,
		_w1284_
	);
	LUT4 #(
		.INIT('h2822)
	) name822 (
		_w534_,
		_w647_,
		_w1265_,
		_w1284_,
		_w1285_
	);
	LUT4 #(
		.INIT('h3f08)
	) name823 (
		_w652_,
		_w1104_,
		_w1106_,
		_w1112_,
		_w1286_
	);
	LUT4 #(
		.INIT('h0133)
	) name824 (
		_w535_,
		_w1184_,
		_w1285_,
		_w1286_,
		_w1287_
	);
	LUT4 #(
		.INIT('h5111)
	) name825 (
		_w525_,
		_w526_,
		_w1147_,
		_w1287_,
		_w1288_
	);
	LUT3 #(
		.INIT('hce)
	) name826 (
		\P1_state_reg[0]/NET0131 ,
		_w512_,
		_w1288_,
		_w1289_
	);
	LUT2 #(
		.INIT('h8)
	) name827 (
		_w537_,
		_w540_,
		_w1290_
	);
	LUT2 #(
		.INIT('h4)
	) name828 (
		_w523_,
		_w1290_,
		_w1291_
	);
	LUT4 #(
		.INIT('ha888)
	) name829 (
		\P1_state_reg[0]/NET0131 ,
		_w510_,
		_w1183_,
		_w1291_,
		_w1292_
	);
	LUT2 #(
		.INIT('h2)
	) name830 (
		\P1_B_reg/NET0131 ,
		_w1292_,
		_w1293_
	);
	LUT4 #(
		.INIT('ha060)
	) name831 (
		\P1_IR_reg[23]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w509_,
		_w1294_
	);
	LUT2 #(
		.INIT('h1)
	) name832 (
		\P2_datao_reg[30]/NET0131 ,
		\si[30]_pad ,
		_w1295_
	);
	LUT4 #(
		.INIT('hfac8)
	) name833 (
		\P2_datao_reg[28]/NET0131 ,
		\P2_datao_reg[29]/NET0131 ,
		\si[28]_pad ,
		\si[29]_pad ,
		_w1296_
	);
	LUT3 #(
		.INIT('h10)
	) name834 (
		_w548_,
		_w1295_,
		_w1296_,
		_w1297_
	);
	LUT2 #(
		.INIT('h8)
	) name835 (
		_w1027_,
		_w1297_,
		_w1298_
	);
	LUT4 #(
		.INIT('h5d00)
	) name836 (
		_w1028_,
		_w1030_,
		_w1044_,
		_w1298_,
		_w1299_
	);
	LUT4 #(
		.INIT('h0b0a)
	) name837 (
		_w544_,
		_w547_,
		_w1295_,
		_w1296_,
		_w1300_
	);
	LUT2 #(
		.INIT('h8)
	) name838 (
		\P2_datao_reg[30]/NET0131 ,
		\si[30]_pad ,
		_w1301_
	);
	LUT4 #(
		.INIT('h000b)
	) name839 (
		_w1026_,
		_w1297_,
		_w1300_,
		_w1301_,
		_w1302_
	);
	LUT4 #(
		.INIT('h1211)
	) name840 (
		\si[31]_pad ,
		_w542_,
		_w1299_,
		_w1302_,
		_w1303_
	);
	LUT3 #(
		.INIT('h12)
	) name841 (
		\P2_datao_reg[31]/NET0131 ,
		_w541_,
		_w1303_,
		_w1304_
	);
	LUT3 #(
		.INIT('h10)
	) name842 (
		_w548_,
		_w549_,
		_w1296_,
		_w1305_
	);
	LUT2 #(
		.INIT('h8)
	) name843 (
		_w986_,
		_w1305_,
		_w1306_
	);
	LUT4 #(
		.INIT('h137f)
	) name844 (
		\P2_datao_reg[28]/NET0131 ,
		\P2_datao_reg[29]/NET0131 ,
		\si[28]_pad ,
		\si[29]_pad ,
		_w1307_
	);
	LUT4 #(
		.INIT('hef00)
	) name845 (
		_w548_,
		_w1015_,
		_w1296_,
		_w1307_,
		_w1308_
	);
	LUT3 #(
		.INIT('hb0)
	) name846 (
		_w995_,
		_w1305_,
		_w1308_,
		_w1309_
	);
	LUT4 #(
		.INIT('h2f00)
	) name847 (
		_w991_,
		_w1064_,
		_w1306_,
		_w1309_,
		_w1310_
	);
	LUT4 #(
		.INIT('h5956)
	) name848 (
		\P2_datao_reg[30]/NET0131 ,
		\si[30]_pad ,
		_w542_,
		_w1310_,
		_w1311_
	);
	LUT2 #(
		.INIT('h1)
	) name849 (
		_w541_,
		_w1311_,
		_w1312_
	);
	LUT3 #(
		.INIT('h32)
	) name850 (
		_w541_,
		_w1179_,
		_w1311_,
		_w1313_
	);
	LUT4 #(
		.INIT('h3031)
	) name851 (
		_w541_,
		_w1151_,
		_w1179_,
		_w1311_,
		_w1314_
	);
	LUT2 #(
		.INIT('h2)
	) name852 (
		_w1304_,
		_w1314_,
		_w1315_
	);
	LUT3 #(
		.INIT('h54)
	) name853 (
		_w645_,
		_w646_,
		_w1275_,
		_w1316_
	);
	LUT2 #(
		.INIT('h1)
	) name854 (
		_w645_,
		_w1258_,
		_w1317_
	);
	LUT3 #(
		.INIT('h54)
	) name855 (
		_w1262_,
		_w1270_,
		_w1279_,
		_w1318_
	);
	LUT4 #(
		.INIT('h0701)
	) name856 (
		_w969_,
		_w977_,
		_w1259_,
		_w1270_,
		_w1319_
	);
	LUT4 #(
		.INIT('h00f1)
	) name857 (
		_w541_,
		_w1033_,
		_w1040_,
		_w1278_,
		_w1320_
	);
	LUT3 #(
		.INIT('h45)
	) name858 (
		_w1260_,
		_w1319_,
		_w1320_,
		_w1321_
	);
	LUT3 #(
		.INIT('h04)
	) name859 (
		_w1256_,
		_w1261_,
		_w1262_,
		_w1322_
	);
	LUT4 #(
		.INIT('h00ef)
	) name860 (
		_w541_,
		_w1046_,
		_w1051_,
		_w1253_,
		_w1323_
	);
	LUT3 #(
		.INIT('h32)
	) name861 (
		_w1247_,
		_w1252_,
		_w1267_,
		_w1324_
	);
	LUT4 #(
		.INIT('h00f1)
	) name862 (
		_w541_,
		_w1046_,
		_w1051_,
		_w1266_,
		_w1325_
	);
	LUT4 #(
		.INIT('hef0e)
	) name863 (
		_w541_,
		_w1046_,
		_w1051_,
		_w1266_,
		_w1326_
	);
	LUT3 #(
		.INIT('h07)
	) name864 (
		_w1323_,
		_w1324_,
		_w1326_,
		_w1327_
	);
	LUT3 #(
		.INIT('h0b)
	) name865 (
		_w738_,
		_w745_,
		_w1186_,
		_w1328_
	);
	LUT4 #(
		.INIT('hdd0d)
	) name866 (
		_w717_,
		_w722_,
		_w786_,
		_w791_,
		_w1329_
	);
	LUT4 #(
		.INIT('h22b2)
	) name867 (
		_w717_,
		_w722_,
		_w786_,
		_w791_,
		_w1330_
	);
	LUT4 #(
		.INIT('h0b00)
	) name868 (
		_w738_,
		_w745_,
		_w1186_,
		_w1330_,
		_w1331_
	);
	LUT4 #(
		.INIT('h0f02)
	) name869 (
		_w738_,
		_w745_,
		_w1186_,
		_w1248_,
		_w1332_
	);
	LUT2 #(
		.INIT('h1)
	) name870 (
		_w1331_,
		_w1332_,
		_w1333_
	);
	LUT2 #(
		.INIT('h1)
	) name871 (
		_w1185_,
		_w1252_,
		_w1334_
	);
	LUT4 #(
		.INIT('h00e8)
	) name872 (
		_w1074_,
		_w1078_,
		_w1185_,
		_w1266_,
		_w1335_
	);
	LUT3 #(
		.INIT('h51)
	) name873 (
		_w1271_,
		_w1323_,
		_w1335_,
		_w1336_
	);
	LUT3 #(
		.INIT('h07)
	) name874 (
		_w1327_,
		_w1333_,
		_w1336_,
		_w1337_
	);
	LUT2 #(
		.INIT('h8)
	) name875 (
		_w1323_,
		_w1334_,
		_w1338_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name876 (
		_w717_,
		_w722_,
		_w786_,
		_w791_,
		_w1339_
	);
	LUT4 #(
		.INIT('h0b00)
	) name877 (
		_w738_,
		_w745_,
		_w1186_,
		_w1339_,
		_w1340_
	);
	LUT3 #(
		.INIT('h80)
	) name878 (
		_w1323_,
		_w1334_,
		_w1340_,
		_w1341_
	);
	LUT4 #(
		.INIT('hdd0d)
	) name879 (
		_w762_,
		_w767_,
		_w772_,
		_w780_,
		_w1342_
	);
	LUT4 #(
		.INIT('h4d44)
	) name880 (
		_w752_,
		_w758_,
		_w808_,
		_w814_,
		_w1343_
	);
	LUT4 #(
		.INIT('h4f04)
	) name881 (
		_w762_,
		_w767_,
		_w772_,
		_w780_,
		_w1344_
	);
	LUT3 #(
		.INIT('h07)
	) name882 (
		_w1342_,
		_w1343_,
		_w1344_,
		_w1345_
	);
	LUT3 #(
		.INIT('h0d)
	) name883 (
		_w799_,
		_w804_,
		_w1196_,
		_w1346_
	);
	LUT2 #(
		.INIT('h1)
	) name884 (
		_w1204_,
		_w1234_,
		_w1347_
	);
	LUT4 #(
		.INIT('h0b02)
	) name885 (
		_w833_,
		_w842_,
		_w1197_,
		_w1204_,
		_w1348_
	);
	LUT3 #(
		.INIT('h51)
	) name886 (
		_w1200_,
		_w1346_,
		_w1348_,
		_w1349_
	);
	LUT4 #(
		.INIT('hdd0d)
	) name887 (
		_w752_,
		_w758_,
		_w808_,
		_w814_,
		_w1350_
	);
	LUT4 #(
		.INIT('h0323)
	) name888 (
		_w1239_,
		_w1241_,
		_w1342_,
		_w1350_,
		_w1351_
	);
	LUT3 #(
		.INIT('ha8)
	) name889 (
		_w1345_,
		_w1349_,
		_w1351_,
		_w1352_
	);
	LUT2 #(
		.INIT('h8)
	) name890 (
		_w1342_,
		_w1350_,
		_w1353_
	);
	LUT2 #(
		.INIT('h1)
	) name891 (
		_w1198_,
		_w1229_,
		_w1354_
	);
	LUT3 #(
		.INIT('h0e)
	) name892 (
		_w1198_,
		_w1229_,
		_w1234_,
		_w1355_
	);
	LUT3 #(
		.INIT('h0b)
	) name893 (
		_w799_,
		_w804_,
		_w1197_,
		_w1356_
	);
	LUT3 #(
		.INIT('hd4)
	) name894 (
		_w799_,
		_w804_,
		_w1197_,
		_w1357_
	);
	LUT3 #(
		.INIT('h07)
	) name895 (
		_w1346_,
		_w1355_,
		_w1357_,
		_w1358_
	);
	LUT2 #(
		.INIT('h2)
	) name896 (
		_w1353_,
		_w1358_,
		_w1359_
	);
	LUT3 #(
		.INIT('hb2)
	) name897 (
		_w857_,
		_w861_,
		_w1206_,
		_w1360_
	);
	LUT3 #(
		.INIT('h32)
	) name898 (
		_w1209_,
		_w1212_,
		_w1217_,
		_w1361_
	);
	LUT2 #(
		.INIT('h1)
	) name899 (
		_w1203_,
		_w1221_,
		_w1362_
	);
	LUT2 #(
		.INIT('h1)
	) name900 (
		_w1211_,
		_w1222_,
		_w1363_
	);
	LUT4 #(
		.INIT('h0001)
	) name901 (
		_w1203_,
		_w1211_,
		_w1221_,
		_w1222_,
		_w1364_
	);
	LUT4 #(
		.INIT('hf200)
	) name902 (
		_w1214_,
		_w1360_,
		_w1361_,
		_w1364_,
		_w1365_
	);
	LUT3 #(
		.INIT('h0d)
	) name903 (
		_w1216_,
		_w1222_,
		_w1226_,
		_w1366_
	);
	LUT3 #(
		.INIT('h54)
	) name904 (
		_w1203_,
		_w1225_,
		_w1230_,
		_w1367_
	);
	LUT3 #(
		.INIT('h0d)
	) name905 (
		_w1362_,
		_w1366_,
		_w1367_,
		_w1368_
	);
	LUT3 #(
		.INIT('h20)
	) name906 (
		_w1345_,
		_w1365_,
		_w1368_,
		_w1369_
	);
	LUT4 #(
		.INIT('h2022)
	) name907 (
		_w1341_,
		_w1352_,
		_w1359_,
		_w1369_,
		_w1370_
	);
	LUT4 #(
		.INIT('h0507)
	) name908 (
		_w1322_,
		_w1337_,
		_w1321_,
		_w1370_,
		_w1371_
	);
	LUT4 #(
		.INIT('h0e0d)
	) name909 (
		\P2_datao_reg[31]/NET0131 ,
		_w541_,
		_w1151_,
		_w1303_,
		_w1372_
	);
	LUT2 #(
		.INIT('h1)
	) name910 (
		_w1151_,
		_w1179_,
		_w1373_
	);
	LUT3 #(
		.INIT('h01)
	) name911 (
		_w541_,
		_w1311_,
		_w1373_,
		_w1374_
	);
	LUT2 #(
		.INIT('h1)
	) name912 (
		_w1372_,
		_w1374_,
		_w1375_
	);
	LUT4 #(
		.INIT('hae00)
	) name913 (
		_w1316_,
		_w1317_,
		_w1371_,
		_w1375_,
		_w1376_
	);
	LUT4 #(
		.INIT('h8884)
	) name914 (
		_w652_,
		_w1112_,
		_w1315_,
		_w1376_,
		_w1377_
	);
	LUT2 #(
		.INIT('h8)
	) name915 (
		_w652_,
		_w1111_,
		_w1378_
	);
	LUT3 #(
		.INIT('h20)
	) name916 (
		_w652_,
		_w1106_,
		_w1111_,
		_w1379_
	);
	LUT4 #(
		.INIT('h08a0)
	) name917 (
		\P1_B_reg/NET0131 ,
		_w652_,
		_w1106_,
		_w1111_,
		_w1380_
	);
	LUT4 #(
		.INIT('h1020)
	) name918 (
		\P2_datao_reg[31]/NET0131 ,
		_w541_,
		_w1151_,
		_w1303_,
		_w1381_
	);
	LUT2 #(
		.INIT('h1)
	) name919 (
		_w1313_,
		_w1381_,
		_w1382_
	);
	LUT3 #(
		.INIT('h04)
	) name920 (
		_w541_,
		_w1179_,
		_w1311_,
		_w1383_
	);
	LUT4 #(
		.INIT('h0071)
	) name921 (
		_w621_,
		_w643_,
		_w1275_,
		_w1383_,
		_w1384_
	);
	LUT3 #(
		.INIT('h51)
	) name922 (
		_w1372_,
		_w1382_,
		_w1384_,
		_w1385_
	);
	LUT2 #(
		.INIT('h8)
	) name923 (
		_w1346_,
		_w1347_,
		_w1386_
	);
	LUT4 #(
		.INIT('h20aa)
	) name924 (
		_w1358_,
		_w1365_,
		_w1368_,
		_w1386_,
		_w1387_
	);
	LUT4 #(
		.INIT('h22a2)
	) name925 (
		_w1341_,
		_w1345_,
		_w1353_,
		_w1387_,
		_w1388_
	);
	LUT4 #(
		.INIT('h0057)
	) name926 (
		_w1322_,
		_w1337_,
		_w1388_,
		_w1321_,
		_w1389_
	);
	LUT4 #(
		.INIT('h0001)
	) name927 (
		_w645_,
		_w1258_,
		_w1372_,
		_w1383_,
		_w1390_
	);
	LUT4 #(
		.INIT('h8a88)
	) name928 (
		_w1379_,
		_w1385_,
		_w1389_,
		_w1390_,
		_w1391_
	);
	LUT3 #(
		.INIT('ha8)
	) name929 (
		_w1104_,
		_w1380_,
		_w1391_,
		_w1392_
	);
	LUT3 #(
		.INIT('h01)
	) name930 (
		_w646_,
		_w1313_,
		_w1381_,
		_w1393_
	);
	LUT3 #(
		.INIT('h01)
	) name931 (
		_w1270_,
		_w1278_,
		_w1279_,
		_w1394_
	);
	LUT3 #(
		.INIT('h80)
	) name932 (
		_w1277_,
		_w1393_,
		_w1394_,
		_w1395_
	);
	LUT3 #(
		.INIT('h70)
	) name933 (
		_w864_,
		_w865_,
		_w869_,
		_w1396_
	);
	LUT4 #(
		.INIT('h020b)
	) name934 (
		_w857_,
		_w861_,
		_w1209_,
		_w1396_,
		_w1397_
	);
	LUT4 #(
		.INIT('h30b0)
	) name935 (
		_w1214_,
		_w1218_,
		_w1363_,
		_w1397_,
		_w1398_
	);
	LUT3 #(
		.INIT('hc4)
	) name936 (
		_w1227_,
		_w1362_,
		_w1398_,
		_w1399_
	);
	LUT3 #(
		.INIT('h0b)
	) name937 (
		_w808_,
		_w814_,
		_w1230_,
		_w1400_
	);
	LUT3 #(
		.INIT('h80)
	) name938 (
		_w1354_,
		_w1356_,
		_w1400_,
		_w1401_
	);
	LUT2 #(
		.INIT('h2)
	) name939 (
		_w1239_,
		_w1241_,
		_w1402_
	);
	LUT2 #(
		.INIT('h8)
	) name940 (
		_w1401_,
		_w1402_,
		_w1403_
	);
	LUT3 #(
		.INIT('h01)
	) name941 (
		_w1247_,
		_w1248_,
		_w1267_,
		_w1404_
	);
	LUT3 #(
		.INIT('hd0)
	) name942 (
		_w738_,
		_w745_,
		_w1329_,
		_w1405_
	);
	LUT3 #(
		.INIT('h80)
	) name943 (
		_w1325_,
		_w1404_,
		_w1405_,
		_w1406_
	);
	LUT4 #(
		.INIT('hba00)
	) name944 (
		_w1352_,
		_w1399_,
		_w1403_,
		_w1406_,
		_w1407_
	);
	LUT2 #(
		.INIT('h8)
	) name945 (
		_w1395_,
		_w1407_,
		_w1408_
	);
	LUT4 #(
		.INIT('h000d)
	) name946 (
		_w738_,
		_w745_,
		_w1245_,
		_w1339_,
		_w1409_
	);
	LUT4 #(
		.INIT('ha200)
	) name947 (
		_w1325_,
		_w1328_,
		_w1409_,
		_w1404_,
		_w1410_
	);
	LUT2 #(
		.INIT('h1)
	) name948 (
		_w1336_,
		_w1410_,
		_w1411_
	);
	LUT3 #(
		.INIT('h32)
	) name949 (
		_w1372_,
		_w1381_,
		_w1383_,
		_w1412_
	);
	LUT4 #(
		.INIT('h04cc)
	) name950 (
		_w1256_,
		_w1261_,
		_w1262_,
		_w1280_,
		_w1413_
	);
	LUT4 #(
		.INIT('h30b0)
	) name951 (
		_w1277_,
		_w1317_,
		_w1393_,
		_w1413_,
		_w1414_
	);
	LUT4 #(
		.INIT('h000b)
	) name952 (
		_w1411_,
		_w1395_,
		_w1412_,
		_w1414_,
		_w1415_
	);
	LUT4 #(
		.INIT('h8000)
	) name953 (
		_w652_,
		_w1104_,
		_w1106_,
		_w1111_,
		_w1416_
	);
	LUT4 #(
		.INIT('hba00)
	) name954 (
		\P1_B_reg/NET0131 ,
		_w1408_,
		_w1415_,
		_w1416_,
		_w1417_
	);
	LUT4 #(
		.INIT('hc8cc)
	) name955 (
		\P1_B_reg/NET0131 ,
		_w1183_,
		_w1408_,
		_w1415_,
		_w1418_
	);
	LUT4 #(
		.INIT('h54ab)
	) name956 (
		_w541_,
		_w1008_,
		_w1017_,
		_w1023_,
		_w1419_
	);
	LUT3 #(
		.INIT('h1e)
	) name957 (
		_w541_,
		_w968_,
		_w977_,
		_w1420_
	);
	LUT3 #(
		.INIT('h1e)
	) name958 (
		_w541_,
		_w701_,
		_w706_,
		_w1421_
	);
	LUT4 #(
		.INIT('h23dc)
	) name959 (
		_w541_,
		_w653_,
		_w673_,
		_w679_,
		_w1422_
	);
	LUT2 #(
		.INIT('h9)
	) name960 (
		_w738_,
		_w745_,
		_w1423_
	);
	LUT4 #(
		.INIT('h0009)
	) name961 (
		_w738_,
		_w745_,
		_w1422_,
		_w1421_,
		_w1424_
	);
	LUT3 #(
		.INIT('h1e)
	) name962 (
		_w541_,
		_w1054_,
		_w1059_,
		_w1425_
	);
	LUT3 #(
		.INIT('h1e)
	) name963 (
		_w541_,
		_w1046_,
		_w1051_,
		_w1426_
	);
	LUT4 #(
		.INIT('h0100)
	) name964 (
		_w1420_,
		_w1425_,
		_w1426_,
		_w1424_,
		_w1427_
	);
	LUT3 #(
		.INIT('h1e)
	) name965 (
		_w541_,
		_w1033_,
		_w1040_,
		_w1428_
	);
	LUT2 #(
		.INIT('h6)
	) name966 (
		_w786_,
		_w791_,
		_w1429_
	);
	LUT3 #(
		.INIT('h1e)
	) name967 (
		_w541_,
		_w1073_,
		_w1078_,
		_w1430_
	);
	LUT2 #(
		.INIT('h6)
	) name968 (
		_w717_,
		_w722_,
		_w1431_
	);
	LUT3 #(
		.INIT('h65)
	) name969 (
		_w998_,
		_w1000_,
		_w1003_,
		_w1432_
	);
	LUT4 #(
		.INIT('h0001)
	) name970 (
		_w1429_,
		_w1430_,
		_w1431_,
		_w1432_,
		_w1433_
	);
	LUT3 #(
		.INIT('h87)
	) name971 (
		_w874_,
		_w875_,
		_w881_,
		_w1434_
	);
	LUT3 #(
		.INIT('h87)
	) name972 (
		_w864_,
		_w865_,
		_w869_,
		_w1435_
	);
	LUT3 #(
		.INIT('h87)
	) name973 (
		_w855_,
		_w856_,
		_w861_,
		_w1436_
	);
	LUT3 #(
		.INIT('h80)
	) name974 (
		_w1435_,
		_w1436_,
		_w1434_,
		_w1437_
	);
	LUT4 #(
		.INIT('h7778)
	) name975 (
		_w817_,
		_w818_,
		_w824_,
		_w826_,
		_w1438_
	);
	LUT3 #(
		.INIT('h87)
	) name976 (
		_w847_,
		_w848_,
		_w853_,
		_w1439_
	);
	LUT3 #(
		.INIT('h87)
	) name977 (
		_w884_,
		_w886_,
		_w894_,
		_w1440_
	);
	LUT3 #(
		.INIT('h78)
	) name978 (
		_w909_,
		_w911_,
		_w918_,
		_w1441_
	);
	LUT4 #(
		.INIT('h0080)
	) name979 (
		_w1438_,
		_w1439_,
		_w1440_,
		_w1441_,
		_w1442_
	);
	LUT2 #(
		.INIT('h6)
	) name980 (
		_w752_,
		_w758_,
		_w1443_
	);
	LUT2 #(
		.INIT('h9)
	) name981 (
		_w762_,
		_w767_,
		_w1444_
	);
	LUT4 #(
		.INIT('h9009)
	) name982 (
		_w752_,
		_w758_,
		_w762_,
		_w767_,
		_w1445_
	);
	LUT3 #(
		.INIT('h80)
	) name983 (
		_w1437_,
		_w1442_,
		_w1445_,
		_w1446_
	);
	LUT2 #(
		.INIT('h9)
	) name984 (
		_w772_,
		_w780_,
		_w1447_
	);
	LUT3 #(
		.INIT('h87)
	) name985 (
		_w921_,
		_w923_,
		_w929_,
		_w1448_
	);
	LUT3 #(
		.INIT('h78)
	) name986 (
		_w932_,
		_w933_,
		_w938_,
		_w1449_
	);
	LUT4 #(
		.INIT('h8887)
	) name987 (
		_w830_,
		_w832_,
		_w838_,
		_w841_,
		_w1450_
	);
	LUT3 #(
		.INIT('h87)
	) name988 (
		_w900_,
		_w902_,
		_w907_,
		_w1451_
	);
	LUT4 #(
		.INIT('h0200)
	) name989 (
		_w1448_,
		_w1449_,
		_w1450_,
		_w1451_,
		_w1452_
	);
	LUT2 #(
		.INIT('h6)
	) name990 (
		_w799_,
		_w804_,
		_w1453_
	);
	LUT2 #(
		.INIT('h6)
	) name991 (
		_w808_,
		_w814_,
		_w1454_
	);
	LUT4 #(
		.INIT('h9009)
	) name992 (
		_w799_,
		_w804_,
		_w808_,
		_w814_,
		_w1455_
	);
	LUT3 #(
		.INIT('h80)
	) name993 (
		_w1447_,
		_w1452_,
		_w1455_,
		_w1456_
	);
	LUT4 #(
		.INIT('h54ab)
	) name994 (
		_w541_,
		_w1062_,
		_w1065_,
		_w1070_,
		_w1457_
	);
	LUT2 #(
		.INIT('h2)
	) name995 (
		_w647_,
		_w1457_,
		_w1458_
	);
	LUT4 #(
		.INIT('h8000)
	) name996 (
		_w1446_,
		_w1456_,
		_w1433_,
		_w1458_,
		_w1459_
	);
	LUT4 #(
		.INIT('h1000)
	) name997 (
		_w1428_,
		_w1419_,
		_w1459_,
		_w1427_,
		_w1460_
	);
	LUT4 #(
		.INIT('h0012)
	) name998 (
		_w1179_,
		_w1372_,
		_w1312_,
		_w1381_,
		_w1461_
	);
	LUT4 #(
		.INIT('h1222)
	) name999 (
		_w652_,
		_w1111_,
		_w1460_,
		_w1461_,
		_w1462_
	);
	LUT3 #(
		.INIT('h28)
	) name1000 (
		\P1_B_reg/NET0131 ,
		\P1_IR_reg[22]/NET0131 ,
		_w513_,
		_w1463_
	);
	LUT3 #(
		.INIT('h70)
	) name1001 (
		_w652_,
		_w1111_,
		_w1463_,
		_w1464_
	);
	LUT3 #(
		.INIT('h54)
	) name1002 (
		_w1106_,
		_w1462_,
		_w1464_,
		_w1465_
	);
	LUT3 #(
		.INIT('h01)
	) name1003 (
		_w1418_,
		_w1465_,
		_w1417_,
		_w1466_
	);
	LUT3 #(
		.INIT('h45)
	) name1004 (
		_w1140_,
		_w1408_,
		_w1415_,
		_w1467_
	);
	LUT2 #(
		.INIT('h4)
	) name1005 (
		_w1104_,
		_w1106_,
		_w1468_
	);
	LUT4 #(
		.INIT('hef00)
	) name1006 (
		_w1378_,
		_w1408_,
		_w1415_,
		_w1468_,
		_w1469_
	);
	LUT3 #(
		.INIT('h10)
	) name1007 (
		_w652_,
		_w1106_,
		_w1111_,
		_w1470_
	);
	LUT4 #(
		.INIT('h0045)
	) name1008 (
		_w1385_,
		_w1389_,
		_w1390_,
		_w1470_,
		_w1471_
	);
	LUT4 #(
		.INIT('h4544)
	) name1009 (
		_w1143_,
		_w1385_,
		_w1389_,
		_w1390_,
		_w1472_
	);
	LUT4 #(
		.INIT('hbbb0)
	) name1010 (
		_w1467_,
		_w1469_,
		_w1471_,
		_w1472_,
		_w1473_
	);
	LUT4 #(
		.INIT('h1000)
	) name1011 (
		_w1392_,
		_w1377_,
		_w1466_,
		_w1473_,
		_w1474_
	);
	LUT3 #(
		.INIT('hae)
	) name1012 (
		_w1293_,
		_w1294_,
		_w1474_,
		_w1475_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name1013 (
		\P2_IR_reg[31]/NET0131 ,
		_w476_,
		_w477_,
		_w490_,
		_w1476_
	);
	LUT2 #(
		.INIT('h9)
	) name1014 (
		\P2_IR_reg[23]/NET0131 ,
		_w1476_,
		_w1477_
	);
	LUT3 #(
		.INIT('h82)
	) name1015 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		_w1476_,
		_w1478_
	);
	LUT4 #(
		.INIT('h70d0)
	) name1016 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg2_reg[28]/NET0131 ,
		_w1476_,
		_w1479_
	);
	LUT3 #(
		.INIT('he0)
	) name1017 (
		\P2_IR_reg[23]/NET0131 ,
		\P2_IR_reg[24]/NET0131 ,
		\P2_IR_reg[31]/NET0131 ,
		_w1480_
	);
	LUT3 #(
		.INIT('h56)
	) name1018 (
		\P2_IR_reg[25]/NET0131 ,
		_w1476_,
		_w1480_,
		_w1481_
	);
	LUT4 #(
		.INIT('hd555)
	) name1019 (
		\P2_IR_reg[31]/NET0131 ,
		_w476_,
		_w478_,
		_w482_,
		_w1482_
	);
	LUT2 #(
		.INIT('h9)
	) name1020 (
		\P2_IR_reg[24]/NET0131 ,
		_w1482_,
		_w1483_
	);
	LUT3 #(
		.INIT('h2a)
	) name1021 (
		\P2_IR_reg[31]/NET0131 ,
		_w482_,
		_w483_,
		_w1484_
	);
	LUT3 #(
		.INIT('h56)
	) name1022 (
		\P2_IR_reg[26]/NET0131 ,
		_w479_,
		_w1484_,
		_w1485_
	);
	LUT3 #(
		.INIT('h80)
	) name1023 (
		_w1483_,
		_w1485_,
		_w1481_,
		_w1486_
	);
	LUT4 #(
		.INIT('h8000)
	) name1024 (
		_w1477_,
		_w1483_,
		_w1485_,
		_w1481_,
		_w1487_
	);
	LUT2 #(
		.INIT('h8)
	) name1025 (
		\P2_reg2_reg[28]/NET0131 ,
		_w1487_,
		_w1488_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name1026 (
		_w1477_,
		_w1483_,
		_w1485_,
		_w1481_,
		_w1489_
	);
	LUT3 #(
		.INIT('h28)
	) name1027 (
		\P2_B_reg/NET0131 ,
		\P2_IR_reg[24]/NET0131 ,
		_w1482_,
		_w1490_
	);
	LUT4 #(
		.INIT('h8c88)
	) name1028 (
		\P2_d_reg[0]/NET0131 ,
		_w1485_,
		_w1481_,
		_w1490_,
		_w1491_
	);
	LUT4 #(
		.INIT('h4441)
	) name1029 (
		\P2_B_reg/NET0131 ,
		\P2_IR_reg[25]/NET0131 ,
		_w1476_,
		_w1480_,
		_w1492_
	);
	LUT3 #(
		.INIT('ha2)
	) name1030 (
		_w1483_,
		_w1485_,
		_w1492_,
		_w1493_
	);
	LUT2 #(
		.INIT('he)
	) name1031 (
		_w1491_,
		_w1493_,
		_w1494_
	);
	LUT3 #(
		.INIT('h96)
	) name1032 (
		\P2_B_reg/NET0131 ,
		\P2_IR_reg[24]/NET0131 ,
		_w1482_,
		_w1495_
	);
	LUT4 #(
		.INIT('hb8bc)
	) name1033 (
		\P2_d_reg[1]/NET0131 ,
		_w1485_,
		_w1481_,
		_w1495_,
		_w1496_
	);
	LUT3 #(
		.INIT('h10)
	) name1034 (
		_w1491_,
		_w1493_,
		_w1496_,
		_w1497_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name1035 (
		\P2_reg2_reg[28]/NET0131 ,
		_w1491_,
		_w1493_,
		_w1496_,
		_w1498_
	);
	LUT4 #(
		.INIT('hff35)
	) name1036 (
		\P2_reg0_reg[6]/NET0131 ,
		\P2_reg2_reg[6]/NET0131 ,
		_w488_,
		_w494_,
		_w1499_
	);
	LUT4 #(
		.INIT('h01fe)
	) name1037 (
		\P2_reg3_reg[3]/NET0131 ,
		\P2_reg3_reg[4]/NET0131 ,
		\P2_reg3_reg[5]/NET0131 ,
		\P2_reg3_reg[6]/NET0131 ,
		_w1500_
	);
	LUT4 #(
		.INIT('hdf1f)
	) name1038 (
		\P2_reg1_reg[6]/NET0131 ,
		_w488_,
		_w494_,
		_w1500_,
		_w1501_
	);
	LUT2 #(
		.INIT('h8)
	) name1039 (
		_w1499_,
		_w1501_,
		_w1502_
	);
	LUT2 #(
		.INIT('h7)
	) name1040 (
		_w1499_,
		_w1501_,
		_w1503_
	);
	LUT4 #(
		.INIT('h8000)
	) name1041 (
		_w476_,
		_w477_,
		_w490_,
		_w491_,
		_w1504_
	);
	LUT3 #(
		.INIT('h59)
	) name1042 (
		\P2_IR_reg[27]/NET0131 ,
		\P2_IR_reg[31]/NET0131 ,
		_w1504_,
		_w1505_
	);
	LUT2 #(
		.INIT('h1)
	) name1043 (
		\P2_IR_reg[26]/NET0131 ,
		\P2_IR_reg[27]/NET0131 ,
		_w1506_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name1044 (
		\P2_IR_reg[31]/NET0131 ,
		_w476_,
		_w478_,
		_w1506_,
		_w1507_
	);
	LUT3 #(
		.INIT('h56)
	) name1045 (
		\P2_IR_reg[28]/NET0131 ,
		_w1484_,
		_w1507_,
		_w1508_
	);
	LUT2 #(
		.INIT('h2)
	) name1046 (
		_w1505_,
		_w1508_,
		_w1509_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name1047 (
		\P2_IR_reg[31]/NET0131 ,
		\P2_IR_reg[4]/NET0131 ,
		\P2_IR_reg[5]/NET0131 ,
		_w472_,
		_w1510_
	);
	LUT2 #(
		.INIT('h6)
	) name1048 (
		\P2_IR_reg[6]/NET0131 ,
		_w1510_,
		_w1511_
	);
	LUT2 #(
		.INIT('h1)
	) name1049 (
		\P1_datao_reg[5]/NET0131 ,
		\si[5]_pad ,
		_w1512_
	);
	LUT2 #(
		.INIT('h8)
	) name1050 (
		\P1_datao_reg[0]/NET0131 ,
		\si[0]_pad ,
		_w1513_
	);
	LUT4 #(
		.INIT('h135f)
	) name1051 (
		\P1_datao_reg[0]/NET0131 ,
		\P1_datao_reg[1]/NET0131 ,
		\si[0]_pad ,
		\si[1]_pad ,
		_w1514_
	);
	LUT4 #(
		.INIT('hfac8)
	) name1052 (
		\P1_datao_reg[1]/NET0131 ,
		\P1_datao_reg[2]/NET0131 ,
		\si[1]_pad ,
		\si[2]_pad ,
		_w1515_
	);
	LUT2 #(
		.INIT('h8)
	) name1053 (
		\P1_datao_reg[2]/NET0131 ,
		\si[2]_pad ,
		_w1516_
	);
	LUT4 #(
		.INIT('h135f)
	) name1054 (
		\P1_datao_reg[2]/NET0131 ,
		\P1_datao_reg[3]/NET0131 ,
		\si[2]_pad ,
		\si[3]_pad ,
		_w1517_
	);
	LUT2 #(
		.INIT('h1)
	) name1055 (
		\P1_datao_reg[3]/NET0131 ,
		\si[3]_pad ,
		_w1518_
	);
	LUT2 #(
		.INIT('h1)
	) name1056 (
		\P1_datao_reg[4]/NET0131 ,
		\si[4]_pad ,
		_w1519_
	);
	LUT4 #(
		.INIT('hfac8)
	) name1057 (
		\P1_datao_reg[3]/NET0131 ,
		\P1_datao_reg[4]/NET0131 ,
		\si[3]_pad ,
		\si[4]_pad ,
		_w1520_
	);
	LUT4 #(
		.INIT('h4f00)
	) name1058 (
		_w1514_,
		_w1515_,
		_w1517_,
		_w1520_,
		_w1521_
	);
	LUT2 #(
		.INIT('h8)
	) name1059 (
		\P1_datao_reg[4]/NET0131 ,
		\si[4]_pad ,
		_w1522_
	);
	LUT4 #(
		.INIT('h135f)
	) name1060 (
		\P1_datao_reg[4]/NET0131 ,
		\P1_datao_reg[5]/NET0131 ,
		\si[4]_pad ,
		\si[5]_pad ,
		_w1523_
	);
	LUT3 #(
		.INIT('h45)
	) name1061 (
		_w1512_,
		_w1521_,
		_w1523_,
		_w1524_
	);
	LUT2 #(
		.INIT('h8)
	) name1062 (
		\P1_datao_reg[6]/NET0131 ,
		\si[6]_pad ,
		_w1525_
	);
	LUT4 #(
		.INIT('h9a6a)
	) name1063 (
		\P1_datao_reg[6]/NET0131 ,
		\si[6]_pad ,
		_w542_,
		_w1524_,
		_w1526_
	);
	LUT4 #(
		.INIT('h02df)
	) name1064 (
		_w1505_,
		_w1508_,
		_w1511_,
		_w1526_,
		_w1527_
	);
	LUT3 #(
		.INIT('h80)
	) name1065 (
		_w1499_,
		_w1501_,
		_w1527_,
		_w1528_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name1066 (
		\P2_reg0_reg[7]/NET0131 ,
		\P2_reg1_reg[7]/NET0131 ,
		_w488_,
		_w494_,
		_w1529_
	);
	LUT2 #(
		.INIT('h9)
	) name1067 (
		\P2_reg3_reg[7]/NET0131 ,
		_w464_,
		_w1530_
	);
	LUT4 #(
		.INIT('hf737)
	) name1068 (
		\P2_reg2_reg[7]/NET0131 ,
		_w488_,
		_w494_,
		_w1530_,
		_w1531_
	);
	LUT2 #(
		.INIT('h8)
	) name1069 (
		_w1529_,
		_w1531_,
		_w1532_
	);
	LUT2 #(
		.INIT('h7)
	) name1070 (
		_w1529_,
		_w1531_,
		_w1533_
	);
	LUT2 #(
		.INIT('h8)
	) name1071 (
		\P1_datao_reg[7]/NET0131 ,
		\si[7]_pad ,
		_w1534_
	);
	LUT3 #(
		.INIT('h0b)
	) name1072 (
		_w1514_,
		_w1515_,
		_w1516_,
		_w1535_
	);
	LUT4 #(
		.INIT('hfac8)
	) name1073 (
		\P1_datao_reg[5]/NET0131 ,
		\P1_datao_reg[6]/NET0131 ,
		\si[5]_pad ,
		\si[6]_pad ,
		_w1536_
	);
	LUT2 #(
		.INIT('h8)
	) name1074 (
		_w1520_,
		_w1536_,
		_w1537_
	);
	LUT4 #(
		.INIT('hec80)
	) name1075 (
		\P1_datao_reg[5]/NET0131 ,
		\P1_datao_reg[6]/NET0131 ,
		\si[5]_pad ,
		\si[6]_pad ,
		_w1538_
	);
	LUT4 #(
		.INIT('h135f)
	) name1076 (
		\P1_datao_reg[3]/NET0131 ,
		\P1_datao_reg[4]/NET0131 ,
		\si[3]_pad ,
		\si[4]_pad ,
		_w1539_
	);
	LUT4 #(
		.INIT('h3323)
	) name1077 (
		_w1519_,
		_w1538_,
		_w1536_,
		_w1539_,
		_w1540_
	);
	LUT3 #(
		.INIT('hb0)
	) name1078 (
		_w1535_,
		_w1537_,
		_w1540_,
		_w1541_
	);
	LUT4 #(
		.INIT('h9565)
	) name1079 (
		\P1_datao_reg[7]/NET0131 ,
		\si[7]_pad ,
		_w542_,
		_w1541_,
		_w1542_
	);
	LUT2 #(
		.INIT('h8)
	) name1080 (
		\P2_IR_reg[31]/NET0131 ,
		\P2_IR_reg[6]/NET0131 ,
		_w1543_
	);
	LUT3 #(
		.INIT('h56)
	) name1081 (
		\P2_IR_reg[7]/NET0131 ,
		_w1510_,
		_w1543_,
		_w1544_
	);
	LUT4 #(
		.INIT('hd0f2)
	) name1082 (
		_w1505_,
		_w1508_,
		_w1542_,
		_w1544_,
		_w1545_
	);
	LUT3 #(
		.INIT('h80)
	) name1083 (
		_w1529_,
		_w1531_,
		_w1545_,
		_w1546_
	);
	LUT2 #(
		.INIT('h1)
	) name1084 (
		_w1528_,
		_w1546_,
		_w1547_
	);
	LUT4 #(
		.INIT('hc5ff)
	) name1085 (
		\P2_reg1_reg[3]/NET0131 ,
		\P2_reg3_reg[3]/NET0131 ,
		_w488_,
		_w494_,
		_w1548_
	);
	LUT4 #(
		.INIT('hff35)
	) name1086 (
		\P2_reg0_reg[3]/NET0131 ,
		\P2_reg2_reg[3]/NET0131 ,
		_w488_,
		_w494_,
		_w1549_
	);
	LUT2 #(
		.INIT('h8)
	) name1087 (
		_w1548_,
		_w1549_,
		_w1550_
	);
	LUT2 #(
		.INIT('h7)
	) name1088 (
		_w1548_,
		_w1549_,
		_w1551_
	);
	LUT4 #(
		.INIT('h9565)
	) name1089 (
		\P1_datao_reg[3]/NET0131 ,
		\si[3]_pad ,
		_w542_,
		_w1535_,
		_w1552_
	);
	LUT4 #(
		.INIT('hfe00)
	) name1090 (
		\P2_IR_reg[0]/NET0131 ,
		\P2_IR_reg[1]/NET0131 ,
		\P2_IR_reg[2]/NET0131 ,
		\P2_IR_reg[31]/NET0131 ,
		_w1553_
	);
	LUT2 #(
		.INIT('h6)
	) name1091 (
		\P2_IR_reg[3]/NET0131 ,
		_w1553_,
		_w1554_
	);
	LUT4 #(
		.INIT('hd0f2)
	) name1092 (
		_w1505_,
		_w1508_,
		_w1552_,
		_w1554_,
		_w1555_
	);
	LUT3 #(
		.INIT('h07)
	) name1093 (
		_w1548_,
		_w1549_,
		_w1555_,
		_w1556_
	);
	LUT4 #(
		.INIT('hf53f)
	) name1094 (
		\P2_reg1_reg[2]/NET0131 ,
		\P2_reg2_reg[2]/NET0131 ,
		_w488_,
		_w494_,
		_w1557_
	);
	LUT4 #(
		.INIT('h3ff5)
	) name1095 (
		\P2_reg0_reg[2]/NET0131 ,
		\P2_reg3_reg[2]/NET0131 ,
		_w488_,
		_w494_,
		_w1558_
	);
	LUT2 #(
		.INIT('h8)
	) name1096 (
		_w1557_,
		_w1558_,
		_w1559_
	);
	LUT2 #(
		.INIT('h7)
	) name1097 (
		_w1557_,
		_w1558_,
		_w1560_
	);
	LUT4 #(
		.INIT('he10f)
	) name1098 (
		\P2_IR_reg[0]/NET0131 ,
		\P2_IR_reg[1]/NET0131 ,
		\P2_IR_reg[2]/NET0131 ,
		\P2_IR_reg[31]/NET0131 ,
		_w1561_
	);
	LUT4 #(
		.INIT('hec80)
	) name1099 (
		\P1_datao_reg[0]/NET0131 ,
		\P1_datao_reg[1]/NET0131 ,
		\si[0]_pad ,
		\si[1]_pad ,
		_w1562_
	);
	LUT4 #(
		.INIT('h9a6a)
	) name1100 (
		\P1_datao_reg[2]/NET0131 ,
		\si[2]_pad ,
		_w542_,
		_w1562_,
		_w1563_
	);
	LUT4 #(
		.INIT('h20fd)
	) name1101 (
		_w1505_,
		_w1508_,
		_w1561_,
		_w1563_,
		_w1564_
	);
	LUT3 #(
		.INIT('h80)
	) name1102 (
		_w1557_,
		_w1558_,
		_w1564_,
		_w1565_
	);
	LUT3 #(
		.INIT('h07)
	) name1103 (
		_w1557_,
		_w1558_,
		_w1564_,
		_w1566_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name1104 (
		\P2_reg2_reg[1]/NET0131 ,
		\P2_reg3_reg[1]/NET0131 ,
		_w488_,
		_w494_,
		_w1567_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name1105 (
		\P2_reg0_reg[1]/NET0131 ,
		\P2_reg1_reg[1]/NET0131 ,
		_w488_,
		_w494_,
		_w1568_
	);
	LUT2 #(
		.INIT('h8)
	) name1106 (
		_w1567_,
		_w1568_,
		_w1569_
	);
	LUT2 #(
		.INIT('h7)
	) name1107 (
		_w1567_,
		_w1568_,
		_w1570_
	);
	LUT3 #(
		.INIT('h93)
	) name1108 (
		\P2_IR_reg[0]/NET0131 ,
		\P2_IR_reg[1]/NET0131 ,
		\P2_IR_reg[31]/NET0131 ,
		_w1571_
	);
	LUT4 #(
		.INIT('h9a6a)
	) name1109 (
		\P1_datao_reg[1]/NET0131 ,
		\si[1]_pad ,
		_w542_,
		_w1513_,
		_w1572_
	);
	LUT4 #(
		.INIT('h20fd)
	) name1110 (
		_w1505_,
		_w1508_,
		_w1571_,
		_w1572_,
		_w1573_
	);
	LUT3 #(
		.INIT('h80)
	) name1111 (
		_w1567_,
		_w1568_,
		_w1573_,
		_w1574_
	);
	LUT3 #(
		.INIT('h07)
	) name1112 (
		_w1567_,
		_w1568_,
		_w1573_,
		_w1575_
	);
	LUT4 #(
		.INIT('h3ff5)
	) name1113 (
		\P2_reg0_reg[0]/NET0131 ,
		\P2_reg3_reg[0]/NET0131 ,
		_w488_,
		_w494_,
		_w1576_
	);
	LUT4 #(
		.INIT('hf53f)
	) name1114 (
		\P2_reg1_reg[0]/NET0131 ,
		\P2_reg2_reg[0]/NET0131 ,
		_w488_,
		_w494_,
		_w1577_
	);
	LUT2 #(
		.INIT('h7)
	) name1115 (
		_w1576_,
		_w1577_,
		_w1578_
	);
	LUT3 #(
		.INIT('h6a)
	) name1116 (
		\P1_datao_reg[0]/NET0131 ,
		\si[0]_pad ,
		_w542_,
		_w1579_
	);
	LUT4 #(
		.INIT('h04f7)
	) name1117 (
		\P2_IR_reg[0]/NET0131 ,
		_w1505_,
		_w1508_,
		_w1579_,
		_w1580_
	);
	LUT3 #(
		.INIT('h07)
	) name1118 (
		_w1576_,
		_w1577_,
		_w1580_,
		_w1581_
	);
	LUT4 #(
		.INIT('h4054)
	) name1119 (
		_w1566_,
		_w1569_,
		_w1573_,
		_w1581_,
		_w1582_
	);
	LUT4 #(
		.INIT('hff35)
	) name1120 (
		\P2_reg0_reg[5]/NET0131 ,
		\P2_reg2_reg[5]/NET0131 ,
		_w488_,
		_w494_,
		_w1583_
	);
	LUT3 #(
		.INIT('h1e)
	) name1121 (
		\P2_reg3_reg[3]/NET0131 ,
		\P2_reg3_reg[4]/NET0131 ,
		\P2_reg3_reg[5]/NET0131 ,
		_w1584_
	);
	LUT4 #(
		.INIT('hdf1f)
	) name1122 (
		\P2_reg1_reg[5]/NET0131 ,
		_w488_,
		_w494_,
		_w1584_,
		_w1585_
	);
	LUT2 #(
		.INIT('h8)
	) name1123 (
		_w1583_,
		_w1585_,
		_w1586_
	);
	LUT2 #(
		.INIT('h7)
	) name1124 (
		_w1583_,
		_w1585_,
		_w1587_
	);
	LUT2 #(
		.INIT('h2)
	) name1125 (
		\P1_datao_reg[5]/NET0131 ,
		_w542_,
		_w1588_
	);
	LUT2 #(
		.INIT('h6)
	) name1126 (
		\P1_datao_reg[5]/NET0131 ,
		\si[5]_pad ,
		_w1589_
	);
	LUT4 #(
		.INIT('h02a8)
	) name1127 (
		_w542_,
		_w1521_,
		_w1522_,
		_w1589_,
		_w1590_
	);
	LUT2 #(
		.INIT('h1)
	) name1128 (
		_w1588_,
		_w1590_,
		_w1591_
	);
	LUT4 #(
		.INIT('h87a5)
	) name1129 (
		\P2_IR_reg[31]/NET0131 ,
		\P2_IR_reg[4]/NET0131 ,
		\P2_IR_reg[5]/NET0131 ,
		_w472_,
		_w1592_
	);
	LUT4 #(
		.INIT('hf2d0)
	) name1130 (
		_w1505_,
		_w1508_,
		_w1591_,
		_w1592_,
		_w1593_
	);
	LUT3 #(
		.INIT('h80)
	) name1131 (
		_w1583_,
		_w1585_,
		_w1593_,
		_w1594_
	);
	LUT3 #(
		.INIT('h80)
	) name1132 (
		_w1548_,
		_w1549_,
		_w1555_,
		_w1595_
	);
	LUT2 #(
		.INIT('h6)
	) name1133 (
		\P2_reg3_reg[3]/NET0131 ,
		\P2_reg3_reg[4]/NET0131 ,
		_w1596_
	);
	LUT4 #(
		.INIT('hf737)
	) name1134 (
		\P2_reg2_reg[4]/NET0131 ,
		_w488_,
		_w494_,
		_w1596_,
		_w1597_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name1135 (
		\P2_reg0_reg[4]/NET0131 ,
		\P2_reg1_reg[4]/NET0131 ,
		_w488_,
		_w494_,
		_w1598_
	);
	LUT2 #(
		.INIT('h8)
	) name1136 (
		_w1597_,
		_w1598_,
		_w1599_
	);
	LUT2 #(
		.INIT('h7)
	) name1137 (
		_w1597_,
		_w1598_,
		_w1600_
	);
	LUT3 #(
		.INIT('hc6)
	) name1138 (
		\P2_IR_reg[31]/NET0131 ,
		\P2_IR_reg[4]/NET0131 ,
		_w472_,
		_w1601_
	);
	LUT4 #(
		.INIT('h004f)
	) name1139 (
		_w1514_,
		_w1515_,
		_w1517_,
		_w1518_,
		_w1602_
	);
	LUT4 #(
		.INIT('h9a6a)
	) name1140 (
		\P1_datao_reg[4]/NET0131 ,
		\si[4]_pad ,
		_w542_,
		_w1602_,
		_w1603_
	);
	LUT4 #(
		.INIT('h02df)
	) name1141 (
		_w1505_,
		_w1508_,
		_w1601_,
		_w1603_,
		_w1604_
	);
	LUT3 #(
		.INIT('h80)
	) name1142 (
		_w1597_,
		_w1598_,
		_w1604_,
		_w1605_
	);
	LUT2 #(
		.INIT('h1)
	) name1143 (
		_w1595_,
		_w1605_,
		_w1606_
	);
	LUT3 #(
		.INIT('h01)
	) name1144 (
		_w1594_,
		_w1595_,
		_w1605_,
		_w1607_
	);
	LUT4 #(
		.INIT('hab00)
	) name1145 (
		_w1556_,
		_w1565_,
		_w1582_,
		_w1607_,
		_w1608_
	);
	LUT3 #(
		.INIT('h07)
	) name1146 (
		_w1583_,
		_w1585_,
		_w1593_,
		_w1609_
	);
	LUT3 #(
		.INIT('h07)
	) name1147 (
		_w1597_,
		_w1598_,
		_w1604_,
		_w1610_
	);
	LUT3 #(
		.INIT('h54)
	) name1148 (
		_w1594_,
		_w1609_,
		_w1610_,
		_w1611_
	);
	LUT3 #(
		.INIT('h07)
	) name1149 (
		_w1529_,
		_w1531_,
		_w1545_,
		_w1612_
	);
	LUT3 #(
		.INIT('h07)
	) name1150 (
		_w1499_,
		_w1501_,
		_w1527_,
		_w1613_
	);
	LUT3 #(
		.INIT('h23)
	) name1151 (
		_w1546_,
		_w1612_,
		_w1613_,
		_w1614_
	);
	LUT3 #(
		.INIT('h70)
	) name1152 (
		_w1547_,
		_w1611_,
		_w1614_,
		_w1615_
	);
	LUT4 #(
		.INIT('hff35)
	) name1153 (
		\P2_reg0_reg[11]/NET0131 ,
		\P2_reg2_reg[11]/NET0131 ,
		_w488_,
		_w494_,
		_w1616_
	);
	LUT3 #(
		.INIT('h63)
	) name1154 (
		\P2_reg3_reg[10]/NET0131 ,
		\P2_reg3_reg[11]/NET0131 ,
		_w465_,
		_w1617_
	);
	LUT4 #(
		.INIT('hdf1f)
	) name1155 (
		\P2_reg1_reg[11]/NET0131 ,
		_w488_,
		_w494_,
		_w1617_,
		_w1618_
	);
	LUT2 #(
		.INIT('h8)
	) name1156 (
		_w1616_,
		_w1618_,
		_w1619_
	);
	LUT2 #(
		.INIT('h7)
	) name1157 (
		_w1616_,
		_w1618_,
		_w1620_
	);
	LUT2 #(
		.INIT('h2)
	) name1158 (
		\P1_datao_reg[11]/NET0131 ,
		_w542_,
		_w1621_
	);
	LUT2 #(
		.INIT('h1)
	) name1159 (
		\P1_datao_reg[11]/NET0131 ,
		\si[11]_pad ,
		_w1622_
	);
	LUT2 #(
		.INIT('h8)
	) name1160 (
		\P1_datao_reg[11]/NET0131 ,
		\si[11]_pad ,
		_w1623_
	);
	LUT2 #(
		.INIT('h6)
	) name1161 (
		\P1_datao_reg[11]/NET0131 ,
		\si[11]_pad ,
		_w1624_
	);
	LUT2 #(
		.INIT('h1)
	) name1162 (
		\P1_datao_reg[10]/NET0131 ,
		\si[10]_pad ,
		_w1625_
	);
	LUT2 #(
		.INIT('h1)
	) name1163 (
		\P1_datao_reg[9]/NET0131 ,
		\si[9]_pad ,
		_w1626_
	);
	LUT4 #(
		.INIT('hfac8)
	) name1164 (
		\P1_datao_reg[10]/NET0131 ,
		\P1_datao_reg[9]/NET0131 ,
		\si[10]_pad ,
		\si[9]_pad ,
		_w1627_
	);
	LUT2 #(
		.INIT('h1)
	) name1165 (
		\P1_datao_reg[8]/NET0131 ,
		\si[8]_pad ,
		_w1628_
	);
	LUT4 #(
		.INIT('hfac8)
	) name1166 (
		\P1_datao_reg[7]/NET0131 ,
		\P1_datao_reg[8]/NET0131 ,
		\si[7]_pad ,
		\si[8]_pad ,
		_w1629_
	);
	LUT2 #(
		.INIT('h8)
	) name1167 (
		_w1627_,
		_w1629_,
		_w1630_
	);
	LUT4 #(
		.INIT('h4f00)
	) name1168 (
		_w1535_,
		_w1537_,
		_w1540_,
		_w1630_,
		_w1631_
	);
	LUT2 #(
		.INIT('h8)
	) name1169 (
		\P1_datao_reg[8]/NET0131 ,
		\si[8]_pad ,
		_w1632_
	);
	LUT4 #(
		.INIT('h135f)
	) name1170 (
		\P1_datao_reg[7]/NET0131 ,
		\P1_datao_reg[8]/NET0131 ,
		\si[7]_pad ,
		\si[8]_pad ,
		_w1633_
	);
	LUT2 #(
		.INIT('h8)
	) name1171 (
		\P1_datao_reg[10]/NET0131 ,
		\si[10]_pad ,
		_w1634_
	);
	LUT4 #(
		.INIT('he8a0)
	) name1172 (
		\P1_datao_reg[10]/NET0131 ,
		\P1_datao_reg[9]/NET0131 ,
		\si[10]_pad ,
		\si[9]_pad ,
		_w1635_
	);
	LUT4 #(
		.INIT('h00fd)
	) name1173 (
		_w1627_,
		_w1628_,
		_w1633_,
		_w1635_,
		_w1636_
	);
	LUT4 #(
		.INIT('h2822)
	) name1174 (
		_w542_,
		_w1624_,
		_w1631_,
		_w1636_,
		_w1637_
	);
	LUT4 #(
		.INIT('hddd0)
	) name1175 (
		_w1505_,
		_w1508_,
		_w1621_,
		_w1637_,
		_w1638_
	);
	LUT3 #(
		.INIT('ha6)
	) name1176 (
		\P2_IR_reg[11]/NET0131 ,
		\P2_IR_reg[31]/NET0131 ,
		_w476_,
		_w1639_
	);
	LUT3 #(
		.INIT('h20)
	) name1177 (
		_w1505_,
		_w1508_,
		_w1639_,
		_w1640_
	);
	LUT2 #(
		.INIT('h1)
	) name1178 (
		_w1638_,
		_w1640_,
		_w1641_
	);
	LUT4 #(
		.INIT('h0008)
	) name1179 (
		_w1616_,
		_w1618_,
		_w1638_,
		_w1640_,
		_w1642_
	);
	LUT2 #(
		.INIT('h9)
	) name1180 (
		\P2_reg3_reg[10]/NET0131 ,
		_w465_,
		_w1643_
	);
	LUT4 #(
		.INIT('hf737)
	) name1181 (
		\P2_reg2_reg[10]/NET0131 ,
		_w488_,
		_w494_,
		_w1643_,
		_w1644_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name1182 (
		\P2_reg0_reg[10]/NET0131 ,
		\P2_reg1_reg[10]/NET0131 ,
		_w488_,
		_w494_,
		_w1645_
	);
	LUT2 #(
		.INIT('h8)
	) name1183 (
		_w1644_,
		_w1645_,
		_w1646_
	);
	LUT2 #(
		.INIT('h7)
	) name1184 (
		_w1644_,
		_w1645_,
		_w1647_
	);
	LUT3 #(
		.INIT('h20)
	) name1185 (
		_w1536_,
		_w1626_,
		_w1629_,
		_w1648_
	);
	LUT4 #(
		.INIT('hec80)
	) name1186 (
		\P1_datao_reg[8]/NET0131 ,
		\P1_datao_reg[9]/NET0131 ,
		\si[8]_pad ,
		\si[9]_pad ,
		_w1649_
	);
	LUT4 #(
		.INIT('h135f)
	) name1187 (
		\P1_datao_reg[6]/NET0131 ,
		\P1_datao_reg[7]/NET0131 ,
		\si[6]_pad ,
		\si[7]_pad ,
		_w1650_
	);
	LUT4 #(
		.INIT('h0f0b)
	) name1188 (
		_w1626_,
		_w1629_,
		_w1649_,
		_w1650_,
		_w1651_
	);
	LUT4 #(
		.INIT('h4f00)
	) name1189 (
		_w1521_,
		_w1523_,
		_w1648_,
		_w1651_,
		_w1652_
	);
	LUT4 #(
		.INIT('h9565)
	) name1190 (
		\P1_datao_reg[10]/NET0131 ,
		\si[10]_pad ,
		_w542_,
		_w1652_,
		_w1653_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name1191 (
		\P2_IR_reg[31]/NET0131 ,
		\P2_IR_reg[4]/NET0131 ,
		_w472_,
		_w473_,
		_w1654_
	);
	LUT3 #(
		.INIT('ha8)
	) name1192 (
		\P2_IR_reg[31]/NET0131 ,
		\P2_IR_reg[8]/NET0131 ,
		\P2_IR_reg[9]/NET0131 ,
		_w1655_
	);
	LUT3 #(
		.INIT('h56)
	) name1193 (
		\P2_IR_reg[10]/NET0131 ,
		_w1654_,
		_w1655_,
		_w1656_
	);
	LUT4 #(
		.INIT('hd0f2)
	) name1194 (
		_w1505_,
		_w1508_,
		_w1653_,
		_w1656_,
		_w1657_
	);
	LUT3 #(
		.INIT('h80)
	) name1195 (
		_w1644_,
		_w1645_,
		_w1657_,
		_w1658_
	);
	LUT2 #(
		.INIT('h1)
	) name1196 (
		_w1642_,
		_w1658_,
		_w1659_
	);
	LUT4 #(
		.INIT('h1e0f)
	) name1197 (
		\P2_reg3_reg[7]/NET0131 ,
		\P2_reg3_reg[8]/NET0131 ,
		\P2_reg3_reg[9]/NET0131 ,
		_w464_,
		_w1660_
	);
	LUT4 #(
		.INIT('hfd3d)
	) name1198 (
		\P2_reg0_reg[9]/NET0131 ,
		_w488_,
		_w494_,
		_w1660_,
		_w1661_
	);
	LUT4 #(
		.INIT('hf53f)
	) name1199 (
		\P2_reg1_reg[9]/NET0131 ,
		\P2_reg2_reg[9]/NET0131 ,
		_w488_,
		_w494_,
		_w1662_
	);
	LUT2 #(
		.INIT('h8)
	) name1200 (
		_w1661_,
		_w1662_,
		_w1663_
	);
	LUT2 #(
		.INIT('h7)
	) name1201 (
		_w1661_,
		_w1662_,
		_w1664_
	);
	LUT2 #(
		.INIT('h1)
	) name1202 (
		_w1534_,
		_w1538_,
		_w1665_
	);
	LUT4 #(
		.INIT('h1f00)
	) name1203 (
		_w1521_,
		_w1522_,
		_w1536_,
		_w1665_,
		_w1666_
	);
	LUT3 #(
		.INIT('h51)
	) name1204 (
		_w1632_,
		_w1629_,
		_w1666_,
		_w1667_
	);
	LUT4 #(
		.INIT('h9565)
	) name1205 (
		\P1_datao_reg[9]/NET0131 ,
		\si[9]_pad ,
		_w542_,
		_w1667_,
		_w1668_
	);
	LUT2 #(
		.INIT('h8)
	) name1206 (
		\P2_IR_reg[31]/NET0131 ,
		\P2_IR_reg[8]/NET0131 ,
		_w1669_
	);
	LUT3 #(
		.INIT('h56)
	) name1207 (
		\P2_IR_reg[9]/NET0131 ,
		_w1654_,
		_w1669_,
		_w1670_
	);
	LUT3 #(
		.INIT('h20)
	) name1208 (
		_w1505_,
		_w1508_,
		_w1670_,
		_w1671_
	);
	LUT3 #(
		.INIT('h0e)
	) name1209 (
		_w1509_,
		_w1668_,
		_w1671_,
		_w1672_
	);
	LUT4 #(
		.INIT('hff35)
	) name1210 (
		\P2_reg0_reg[8]/NET0131 ,
		\P2_reg2_reg[8]/NET0131 ,
		_w488_,
		_w494_,
		_w1673_
	);
	LUT3 #(
		.INIT('h63)
	) name1211 (
		\P2_reg3_reg[7]/NET0131 ,
		\P2_reg3_reg[8]/NET0131 ,
		_w464_,
		_w1674_
	);
	LUT4 #(
		.INIT('hdf1f)
	) name1212 (
		\P2_reg1_reg[8]/NET0131 ,
		_w488_,
		_w494_,
		_w1674_,
		_w1675_
	);
	LUT2 #(
		.INIT('h8)
	) name1213 (
		_w1673_,
		_w1675_,
		_w1676_
	);
	LUT2 #(
		.INIT('h7)
	) name1214 (
		_w1673_,
		_w1675_,
		_w1677_
	);
	LUT4 #(
		.INIT('h00ba)
	) name1215 (
		_w1512_,
		_w1521_,
		_w1523_,
		_w1525_,
		_w1678_
	);
	LUT4 #(
		.INIT('hfac8)
	) name1216 (
		\P1_datao_reg[6]/NET0131 ,
		\P1_datao_reg[7]/NET0131 ,
		\si[6]_pad ,
		\si[7]_pad ,
		_w1679_
	);
	LUT3 #(
		.INIT('h45)
	) name1217 (
		_w1534_,
		_w1678_,
		_w1679_,
		_w1680_
	);
	LUT4 #(
		.INIT('h9565)
	) name1218 (
		\P1_datao_reg[8]/NET0131 ,
		\si[8]_pad ,
		_w542_,
		_w1680_,
		_w1681_
	);
	LUT3 #(
		.INIT('hc6)
	) name1219 (
		\P2_IR_reg[31]/NET0131 ,
		\P2_IR_reg[8]/NET0131 ,
		_w474_,
		_w1682_
	);
	LUT3 #(
		.INIT('h20)
	) name1220 (
		_w1505_,
		_w1508_,
		_w1682_,
		_w1683_
	);
	LUT3 #(
		.INIT('h0e)
	) name1221 (
		_w1509_,
		_w1681_,
		_w1683_,
		_w1684_
	);
	LUT4 #(
		.INIT('h0777)
	) name1222 (
		_w1663_,
		_w1672_,
		_w1676_,
		_w1684_,
		_w1685_
	);
	LUT2 #(
		.INIT('h8)
	) name1223 (
		_w1659_,
		_w1685_,
		_w1686_
	);
	LUT4 #(
		.INIT('h8f00)
	) name1224 (
		_w1547_,
		_w1608_,
		_w1615_,
		_w1686_,
		_w1687_
	);
	LUT4 #(
		.INIT('heee8)
	) name1225 (
		_w1663_,
		_w1672_,
		_w1676_,
		_w1684_,
		_w1688_
	);
	LUT4 #(
		.INIT('h7770)
	) name1226 (
		_w1616_,
		_w1618_,
		_w1638_,
		_w1640_,
		_w1689_
	);
	LUT3 #(
		.INIT('h07)
	) name1227 (
		_w1644_,
		_w1645_,
		_w1657_,
		_w1690_
	);
	LUT3 #(
		.INIT('h54)
	) name1228 (
		_w1642_,
		_w1689_,
		_w1690_,
		_w1691_
	);
	LUT3 #(
		.INIT('h0d)
	) name1229 (
		_w1659_,
		_w1688_,
		_w1691_,
		_w1692_
	);
	LUT4 #(
		.INIT('h1e0f)
	) name1230 (
		\P2_reg3_reg[13]/NET0131 ,
		\P2_reg3_reg[14]/NET0131 ,
		\P2_reg3_reg[15]/NET0131 ,
		_w467_,
		_w1693_
	);
	LUT3 #(
		.INIT('h08)
	) name1231 (
		_w488_,
		_w494_,
		_w1693_,
		_w1694_
	);
	LUT3 #(
		.INIT('h02)
	) name1232 (
		\P2_reg0_reg[15]/NET0131 ,
		_w488_,
		_w494_,
		_w1695_
	);
	LUT4 #(
		.INIT('hf53f)
	) name1233 (
		\P2_reg1_reg[15]/NET0131 ,
		\P2_reg2_reg[15]/NET0131 ,
		_w488_,
		_w494_,
		_w1696_
	);
	LUT3 #(
		.INIT('h10)
	) name1234 (
		_w1694_,
		_w1695_,
		_w1696_,
		_w1697_
	);
	LUT3 #(
		.INIT('hef)
	) name1235 (
		_w1694_,
		_w1695_,
		_w1696_,
		_w1698_
	);
	LUT2 #(
		.INIT('h1)
	) name1236 (
		\P1_datao_reg[15]/NET0131 ,
		\si[15]_pad ,
		_w1699_
	);
	LUT2 #(
		.INIT('h8)
	) name1237 (
		\P1_datao_reg[15]/NET0131 ,
		\si[15]_pad ,
		_w1700_
	);
	LUT2 #(
		.INIT('h1)
	) name1238 (
		\P1_datao_reg[12]/NET0131 ,
		\si[12]_pad ,
		_w1701_
	);
	LUT2 #(
		.INIT('h1)
	) name1239 (
		\P1_datao_reg[13]/NET0131 ,
		\si[13]_pad ,
		_w1702_
	);
	LUT4 #(
		.INIT('hfac8)
	) name1240 (
		\P1_datao_reg[13]/NET0131 ,
		\P1_datao_reg[14]/NET0131 ,
		\si[13]_pad ,
		\si[14]_pad ,
		_w1703_
	);
	LUT2 #(
		.INIT('h8)
	) name1241 (
		\P1_datao_reg[12]/NET0131 ,
		\si[12]_pad ,
		_w1704_
	);
	LUT4 #(
		.INIT('h135f)
	) name1242 (
		\P1_datao_reg[11]/NET0131 ,
		\P1_datao_reg[12]/NET0131 ,
		\si[11]_pad ,
		\si[12]_pad ,
		_w1705_
	);
	LUT4 #(
		.INIT('hec80)
	) name1243 (
		\P1_datao_reg[13]/NET0131 ,
		\P1_datao_reg[14]/NET0131 ,
		\si[13]_pad ,
		\si[14]_pad ,
		_w1706_
	);
	LUT4 #(
		.INIT('h00fb)
	) name1244 (
		_w1701_,
		_w1703_,
		_w1705_,
		_w1706_,
		_w1707_
	);
	LUT4 #(
		.INIT('hfac8)
	) name1245 (
		\P1_datao_reg[11]/NET0131 ,
		\P1_datao_reg[12]/NET0131 ,
		\si[11]_pad ,
		\si[12]_pad ,
		_w1708_
	);
	LUT2 #(
		.INIT('h8)
	) name1246 (
		_w1703_,
		_w1708_,
		_w1709_
	);
	LUT4 #(
		.INIT('h40f0)
	) name1247 (
		_w1631_,
		_w1636_,
		_w1707_,
		_w1709_,
		_w1710_
	);
	LUT4 #(
		.INIT('h9565)
	) name1248 (
		\P1_datao_reg[15]/NET0131 ,
		\si[15]_pad ,
		_w542_,
		_w1710_,
		_w1711_
	);
	LUT4 #(
		.INIT('h7333)
	) name1249 (
		\P2_IR_reg[14]/NET0131 ,
		\P2_IR_reg[31]/NET0131 ,
		_w476_,
		_w478_,
		_w1712_
	);
	LUT2 #(
		.INIT('h9)
	) name1250 (
		\P2_IR_reg[15]/NET0131 ,
		_w1712_,
		_w1713_
	);
	LUT3 #(
		.INIT('h20)
	) name1251 (
		_w1505_,
		_w1508_,
		_w1713_,
		_w1714_
	);
	LUT3 #(
		.INIT('h0e)
	) name1252 (
		_w1509_,
		_w1711_,
		_w1714_,
		_w1715_
	);
	LUT2 #(
		.INIT('h8)
	) name1253 (
		_w1697_,
		_w1715_,
		_w1716_
	);
	LUT4 #(
		.INIT('hff35)
	) name1254 (
		\P2_reg0_reg[14]/NET0131 ,
		\P2_reg2_reg[14]/NET0131 ,
		_w488_,
		_w494_,
		_w1717_
	);
	LUT3 #(
		.INIT('h63)
	) name1255 (
		\P2_reg3_reg[13]/NET0131 ,
		\P2_reg3_reg[14]/NET0131 ,
		_w467_,
		_w1718_
	);
	LUT4 #(
		.INIT('hdf1f)
	) name1256 (
		\P2_reg1_reg[14]/NET0131 ,
		_w488_,
		_w494_,
		_w1718_,
		_w1719_
	);
	LUT2 #(
		.INIT('h8)
	) name1257 (
		_w1717_,
		_w1719_,
		_w1720_
	);
	LUT2 #(
		.INIT('h7)
	) name1258 (
		_w1717_,
		_w1719_,
		_w1721_
	);
	LUT3 #(
		.INIT('h10)
	) name1259 (
		_w1625_,
		_w1702_,
		_w1708_,
		_w1722_
	);
	LUT4 #(
		.INIT('hec80)
	) name1260 (
		\P1_datao_reg[12]/NET0131 ,
		\P1_datao_reg[13]/NET0131 ,
		\si[12]_pad ,
		\si[13]_pad ,
		_w1723_
	);
	LUT4 #(
		.INIT('h135f)
	) name1261 (
		\P1_datao_reg[10]/NET0131 ,
		\P1_datao_reg[11]/NET0131 ,
		\si[10]_pad ,
		\si[11]_pad ,
		_w1724_
	);
	LUT4 #(
		.INIT('h0f0b)
	) name1262 (
		_w1702_,
		_w1708_,
		_w1723_,
		_w1724_,
		_w1725_
	);
	LUT3 #(
		.INIT('hb0)
	) name1263 (
		_w1652_,
		_w1722_,
		_w1725_,
		_w1726_
	);
	LUT4 #(
		.INIT('h9565)
	) name1264 (
		\P1_datao_reg[14]/NET0131 ,
		\si[14]_pad ,
		_w542_,
		_w1726_,
		_w1727_
	);
	LUT4 #(
		.INIT('h5999)
	) name1265 (
		\P2_IR_reg[14]/NET0131 ,
		\P2_IR_reg[31]/NET0131 ,
		_w476_,
		_w478_,
		_w1728_
	);
	LUT3 #(
		.INIT('h02)
	) name1266 (
		_w1505_,
		_w1508_,
		_w1728_,
		_w1729_
	);
	LUT3 #(
		.INIT('h0e)
	) name1267 (
		_w1509_,
		_w1727_,
		_w1729_,
		_w1730_
	);
	LUT4 #(
		.INIT('h0777)
	) name1268 (
		_w1697_,
		_w1715_,
		_w1720_,
		_w1730_,
		_w1731_
	);
	LUT4 #(
		.INIT('h1e0f)
	) name1269 (
		\P2_reg3_reg[10]/NET0131 ,
		\P2_reg3_reg[11]/NET0131 ,
		\P2_reg3_reg[12]/NET0131 ,
		_w465_,
		_w1732_
	);
	LUT4 #(
		.INIT('hdf1f)
	) name1270 (
		\P2_reg1_reg[12]/NET0131 ,
		_w488_,
		_w494_,
		_w1732_,
		_w1733_
	);
	LUT4 #(
		.INIT('hff35)
	) name1271 (
		\P2_reg0_reg[12]/NET0131 ,
		\P2_reg2_reg[12]/NET0131 ,
		_w488_,
		_w494_,
		_w1734_
	);
	LUT2 #(
		.INIT('h8)
	) name1272 (
		_w1733_,
		_w1734_,
		_w1735_
	);
	LUT2 #(
		.INIT('h7)
	) name1273 (
		_w1733_,
		_w1734_,
		_w1736_
	);
	LUT2 #(
		.INIT('h2)
	) name1274 (
		\P1_datao_reg[12]/NET0131 ,
		_w542_,
		_w1737_
	);
	LUT2 #(
		.INIT('h6)
	) name1275 (
		\P1_datao_reg[12]/NET0131 ,
		\si[12]_pad ,
		_w1738_
	);
	LUT3 #(
		.INIT('h04)
	) name1276 (
		_w1622_,
		_w1627_,
		_w1628_,
		_w1739_
	);
	LUT4 #(
		.INIT('hba00)
	) name1277 (
		_w1534_,
		_w1678_,
		_w1679_,
		_w1739_,
		_w1740_
	);
	LUT4 #(
		.INIT('hfac8)
	) name1278 (
		\P1_datao_reg[10]/NET0131 ,
		\P1_datao_reg[11]/NET0131 ,
		\si[10]_pad ,
		\si[11]_pad ,
		_w1741_
	);
	LUT4 #(
		.INIT('h0155)
	) name1279 (
		_w1623_,
		_w1634_,
		_w1649_,
		_w1741_,
		_w1742_
	);
	LUT4 #(
		.INIT('h2822)
	) name1280 (
		_w542_,
		_w1738_,
		_w1740_,
		_w1742_,
		_w1743_
	);
	LUT4 #(
		.INIT('h6c3c)
	) name1281 (
		\P2_IR_reg[11]/NET0131 ,
		\P2_IR_reg[12]/NET0131 ,
		\P2_IR_reg[31]/NET0131 ,
		_w476_,
		_w1744_
	);
	LUT3 #(
		.INIT('h20)
	) name1282 (
		_w1505_,
		_w1508_,
		_w1744_,
		_w1745_
	);
	LUT4 #(
		.INIT('h00ab)
	) name1283 (
		_w1509_,
		_w1737_,
		_w1743_,
		_w1745_,
		_w1746_
	);
	LUT4 #(
		.INIT('hff35)
	) name1284 (
		\P2_reg0_reg[13]/NET0131 ,
		\P2_reg2_reg[13]/NET0131 ,
		_w488_,
		_w494_,
		_w1747_
	);
	LUT3 #(
		.INIT('he0)
	) name1285 (
		\P2_reg3_reg[1]/NET0131 ,
		\P2_reg3_reg[2]/NET0131 ,
		\P2_reg3_reg[3]/NET0131 ,
		_w1748_
	);
	LUT3 #(
		.INIT('h19)
	) name1286 (
		\P2_reg3_reg[13]/NET0131 ,
		_w467_,
		_w1748_,
		_w1749_
	);
	LUT4 #(
		.INIT('hdf1f)
	) name1287 (
		\P2_reg1_reg[13]/NET0131 ,
		_w488_,
		_w494_,
		_w1749_,
		_w1750_
	);
	LUT2 #(
		.INIT('h8)
	) name1288 (
		_w1747_,
		_w1750_,
		_w1751_
	);
	LUT2 #(
		.INIT('h7)
	) name1289 (
		_w1747_,
		_w1750_,
		_w1752_
	);
	LUT2 #(
		.INIT('h2)
	) name1290 (
		\P1_datao_reg[13]/NET0131 ,
		_w542_,
		_w1753_
	);
	LUT2 #(
		.INIT('h6)
	) name1291 (
		\P1_datao_reg[13]/NET0131 ,
		\si[13]_pad ,
		_w1754_
	);
	LUT4 #(
		.INIT('h010f)
	) name1292 (
		_w1623_,
		_w1635_,
		_w1704_,
		_w1708_,
		_w1755_
	);
	LUT2 #(
		.INIT('h8)
	) name1293 (
		_w1627_,
		_w1708_,
		_w1756_
	);
	LUT4 #(
		.INIT('hae00)
	) name1294 (
		_w1632_,
		_w1629_,
		_w1666_,
		_w1756_,
		_w1757_
	);
	LUT4 #(
		.INIT('h2282)
	) name1295 (
		_w542_,
		_w1754_,
		_w1755_,
		_w1757_,
		_w1758_
	);
	LUT4 #(
		.INIT('ha666)
	) name1296 (
		\P2_IR_reg[13]/NET0131 ,
		\P2_IR_reg[31]/NET0131 ,
		_w476_,
		_w477_,
		_w1759_
	);
	LUT3 #(
		.INIT('h20)
	) name1297 (
		_w1505_,
		_w1508_,
		_w1759_,
		_w1760_
	);
	LUT4 #(
		.INIT('h00ab)
	) name1298 (
		_w1509_,
		_w1753_,
		_w1758_,
		_w1760_,
		_w1761_
	);
	LUT4 #(
		.INIT('h0777)
	) name1299 (
		_w1735_,
		_w1746_,
		_w1751_,
		_w1761_,
		_w1762_
	);
	LUT2 #(
		.INIT('h8)
	) name1300 (
		_w1731_,
		_w1762_,
		_w1763_
	);
	LUT2 #(
		.INIT('h8)
	) name1301 (
		\P1_datao_reg[17]/NET0131 ,
		\si[17]_pad ,
		_w1764_
	);
	LUT2 #(
		.INIT('h8)
	) name1302 (
		\P1_datao_reg[16]/NET0131 ,
		\si[16]_pad ,
		_w1765_
	);
	LUT2 #(
		.INIT('h1)
	) name1303 (
		\P1_datao_reg[16]/NET0131 ,
		\si[16]_pad ,
		_w1766_
	);
	LUT4 #(
		.INIT('hfac8)
	) name1304 (
		\P1_datao_reg[15]/NET0131 ,
		\P1_datao_reg[16]/NET0131 ,
		\si[15]_pad ,
		\si[16]_pad ,
		_w1767_
	);
	LUT4 #(
		.INIT('h010f)
	) name1305 (
		_w1700_,
		_w1706_,
		_w1765_,
		_w1767_,
		_w1768_
	);
	LUT2 #(
		.INIT('h8)
	) name1306 (
		_w1703_,
		_w1767_,
		_w1769_
	);
	LUT4 #(
		.INIT('h20f0)
	) name1307 (
		_w1755_,
		_w1757_,
		_w1768_,
		_w1769_,
		_w1770_
	);
	LUT4 #(
		.INIT('h9565)
	) name1308 (
		\P1_datao_reg[17]/NET0131 ,
		\si[17]_pad ,
		_w542_,
		_w1770_,
		_w1771_
	);
	LUT4 #(
		.INIT('hfe00)
	) name1309 (
		\P2_IR_reg[14]/NET0131 ,
		\P2_IR_reg[15]/NET0131 ,
		\P2_IR_reg[16]/NET0131 ,
		\P2_IR_reg[31]/NET0131 ,
		_w1772_
	);
	LUT4 #(
		.INIT('h00d5)
	) name1310 (
		\P2_IR_reg[31]/NET0131 ,
		_w476_,
		_w478_,
		_w1772_,
		_w1773_
	);
	LUT2 #(
		.INIT('h9)
	) name1311 (
		\P2_IR_reg[17]/NET0131 ,
		_w1773_,
		_w1774_
	);
	LUT3 #(
		.INIT('h20)
	) name1312 (
		_w1505_,
		_w1508_,
		_w1774_,
		_w1775_
	);
	LUT3 #(
		.INIT('h0e)
	) name1313 (
		_w1509_,
		_w1771_,
		_w1775_,
		_w1776_
	);
	LUT4 #(
		.INIT('h5595)
	) name1314 (
		\P2_reg3_reg[17]/NET0131 ,
		_w467_,
		_w469_,
		_w1748_,
		_w1777_
	);
	LUT3 #(
		.INIT('h08)
	) name1315 (
		_w488_,
		_w494_,
		_w1777_,
		_w1778_
	);
	LUT3 #(
		.INIT('h20)
	) name1316 (
		\P2_reg1_reg[17]/NET0131 ,
		_w488_,
		_w494_,
		_w1779_
	);
	LUT4 #(
		.INIT('hff35)
	) name1317 (
		\P2_reg0_reg[17]/NET0131 ,
		\P2_reg2_reg[17]/NET0131 ,
		_w488_,
		_w494_,
		_w1780_
	);
	LUT3 #(
		.INIT('h10)
	) name1318 (
		_w1779_,
		_w1778_,
		_w1780_,
		_w1781_
	);
	LUT3 #(
		.INIT('hef)
	) name1319 (
		_w1779_,
		_w1778_,
		_w1780_,
		_w1782_
	);
	LUT4 #(
		.INIT('h0e00)
	) name1320 (
		_w1509_,
		_w1771_,
		_w1775_,
		_w1781_,
		_w1783_
	);
	LUT3 #(
		.INIT('h10)
	) name1321 (
		_w1699_,
		_w1701_,
		_w1703_,
		_w1784_
	);
	LUT4 #(
		.INIT('hfac8)
	) name1322 (
		\P1_datao_reg[14]/NET0131 ,
		\P1_datao_reg[15]/NET0131 ,
		\si[14]_pad ,
		\si[15]_pad ,
		_w1785_
	);
	LUT4 #(
		.INIT('hec80)
	) name1323 (
		\P1_datao_reg[14]/NET0131 ,
		\P1_datao_reg[15]/NET0131 ,
		\si[14]_pad ,
		\si[15]_pad ,
		_w1786_
	);
	LUT3 #(
		.INIT('h07)
	) name1324 (
		_w1723_,
		_w1785_,
		_w1786_,
		_w1787_
	);
	LUT3 #(
		.INIT('hb0)
	) name1325 (
		_w1742_,
		_w1784_,
		_w1787_,
		_w1788_
	);
	LUT3 #(
		.INIT('h70)
	) name1326 (
		_w1740_,
		_w1784_,
		_w1788_,
		_w1789_
	);
	LUT4 #(
		.INIT('h9565)
	) name1327 (
		\P1_datao_reg[16]/NET0131 ,
		\si[16]_pad ,
		_w542_,
		_w1789_,
		_w1790_
	);
	LUT3 #(
		.INIT('he0)
	) name1328 (
		\P2_IR_reg[14]/NET0131 ,
		\P2_IR_reg[15]/NET0131 ,
		\P2_IR_reg[31]/NET0131 ,
		_w1791_
	);
	LUT4 #(
		.INIT('h00d5)
	) name1329 (
		\P2_IR_reg[31]/NET0131 ,
		_w476_,
		_w478_,
		_w1791_,
		_w1792_
	);
	LUT2 #(
		.INIT('h9)
	) name1330 (
		\P2_IR_reg[16]/NET0131 ,
		_w1792_,
		_w1793_
	);
	LUT3 #(
		.INIT('h20)
	) name1331 (
		_w1505_,
		_w1508_,
		_w1793_,
		_w1794_
	);
	LUT3 #(
		.INIT('h0e)
	) name1332 (
		_w1509_,
		_w1790_,
		_w1794_,
		_w1795_
	);
	LUT4 #(
		.INIT('h00a8)
	) name1333 (
		_w498_,
		_w1509_,
		_w1790_,
		_w1794_,
		_w1796_
	);
	LUT2 #(
		.INIT('h2)
	) name1334 (
		\P1_datao_reg[19]/NET0131 ,
		_w542_,
		_w1797_
	);
	LUT2 #(
		.INIT('h1)
	) name1335 (
		\P1_datao_reg[19]/NET0131 ,
		\si[19]_pad ,
		_w1798_
	);
	LUT2 #(
		.INIT('h6)
	) name1336 (
		\P1_datao_reg[19]/NET0131 ,
		\si[19]_pad ,
		_w1799_
	);
	LUT4 #(
		.INIT('hfac8)
	) name1337 (
		\P1_datao_reg[17]/NET0131 ,
		\P1_datao_reg[18]/NET0131 ,
		\si[17]_pad ,
		\si[18]_pad ,
		_w1800_
	);
	LUT2 #(
		.INIT('h8)
	) name1338 (
		_w1767_,
		_w1800_,
		_w1801_
	);
	LUT4 #(
		.INIT('hec80)
	) name1339 (
		\P1_datao_reg[17]/NET0131 ,
		\P1_datao_reg[18]/NET0131 ,
		\si[17]_pad ,
		\si[18]_pad ,
		_w1802_
	);
	LUT4 #(
		.INIT('h137f)
	) name1340 (
		\P1_datao_reg[15]/NET0131 ,
		\P1_datao_reg[16]/NET0131 ,
		\si[15]_pad ,
		\si[16]_pad ,
		_w1803_
	);
	LUT2 #(
		.INIT('h4)
	) name1341 (
		_w1802_,
		_w1803_,
		_w1804_
	);
	LUT4 #(
		.INIT('h0137)
	) name1342 (
		\P1_datao_reg[17]/NET0131 ,
		\P1_datao_reg[18]/NET0131 ,
		\si[17]_pad ,
		\si[18]_pad ,
		_w1805_
	);
	LUT4 #(
		.INIT('h004f)
	) name1343 (
		_w1707_,
		_w1801_,
		_w1804_,
		_w1805_,
		_w1806_
	);
	LUT4 #(
		.INIT('hb000)
	) name1344 (
		_w1631_,
		_w1636_,
		_w1709_,
		_w1801_,
		_w1807_
	);
	LUT4 #(
		.INIT('h2228)
	) name1345 (
		_w542_,
		_w1799_,
		_w1806_,
		_w1807_,
		_w1808_
	);
	LUT4 #(
		.INIT('he0f0)
	) name1346 (
		\P2_IR_reg[13]/NET0131 ,
		\P2_IR_reg[18]/NET0131 ,
		\P2_IR_reg[31]/NET0131 ,
		_w480_,
		_w1809_
	);
	LUT4 #(
		.INIT('h00d5)
	) name1347 (
		\P2_IR_reg[31]/NET0131 ,
		_w476_,
		_w477_,
		_w1809_,
		_w1810_
	);
	LUT2 #(
		.INIT('h9)
	) name1348 (
		\P2_IR_reg[19]/NET0131 ,
		_w1810_,
		_w1811_
	);
	LUT3 #(
		.INIT('h20)
	) name1349 (
		_w1505_,
		_w1508_,
		_w1811_,
		_w1812_
	);
	LUT4 #(
		.INIT('h00ab)
	) name1350 (
		_w1509_,
		_w1797_,
		_w1808_,
		_w1812_,
		_w1813_
	);
	LUT4 #(
		.INIT('h1000)
	) name1351 (
		\P2_reg3_reg[17]/NET0131 ,
		\P2_reg3_reg[18]/NET0131 ,
		_w467_,
		_w469_,
		_w1814_
	);
	LUT2 #(
		.INIT('h9)
	) name1352 (
		\P2_reg3_reg[19]/NET0131 ,
		_w1814_,
		_w1815_
	);
	LUT4 #(
		.INIT('h4080)
	) name1353 (
		\P2_reg3_reg[19]/NET0131 ,
		_w488_,
		_w494_,
		_w1814_,
		_w1816_
	);
	LUT3 #(
		.INIT('h20)
	) name1354 (
		\P2_reg1_reg[19]/NET0131 ,
		_w488_,
		_w494_,
		_w1817_
	);
	LUT4 #(
		.INIT('hff35)
	) name1355 (
		\P2_reg0_reg[19]/NET0131 ,
		\P2_reg2_reg[19]/NET0131 ,
		_w488_,
		_w494_,
		_w1818_
	);
	LUT3 #(
		.INIT('h10)
	) name1356 (
		_w1817_,
		_w1816_,
		_w1818_,
		_w1819_
	);
	LUT3 #(
		.INIT('hef)
	) name1357 (
		_w1817_,
		_w1816_,
		_w1818_,
		_w1820_
	);
	LUT2 #(
		.INIT('h8)
	) name1358 (
		_w1813_,
		_w1819_,
		_w1821_
	);
	LUT2 #(
		.INIT('h2)
	) name1359 (
		\P1_datao_reg[18]/NET0131 ,
		_w542_,
		_w1822_
	);
	LUT2 #(
		.INIT('h6)
	) name1360 (
		\P1_datao_reg[18]/NET0131 ,
		\si[18]_pad ,
		_w1823_
	);
	LUT4 #(
		.INIT('hfac8)
	) name1361 (
		\P1_datao_reg[16]/NET0131 ,
		\P1_datao_reg[17]/NET0131 ,
		\si[16]_pad ,
		\si[17]_pad ,
		_w1824_
	);
	LUT4 #(
		.INIT('h0155)
	) name1362 (
		_w1764_,
		_w1765_,
		_w1786_,
		_w1824_,
		_w1825_
	);
	LUT2 #(
		.INIT('h8)
	) name1363 (
		_w1785_,
		_w1824_,
		_w1826_
	);
	LUT4 #(
		.INIT('h4f00)
	) name1364 (
		_w1652_,
		_w1722_,
		_w1725_,
		_w1826_,
		_w1827_
	);
	LUT4 #(
		.INIT('h2282)
	) name1365 (
		_w542_,
		_w1823_,
		_w1825_,
		_w1827_,
		_w1828_
	);
	LUT2 #(
		.INIT('h2)
	) name1366 (
		\P2_IR_reg[31]/NET0131 ,
		_w480_,
		_w1829_
	);
	LUT4 #(
		.INIT('h00d5)
	) name1367 (
		\P2_IR_reg[31]/NET0131 ,
		_w476_,
		_w478_,
		_w1829_,
		_w1830_
	);
	LUT2 #(
		.INIT('h9)
	) name1368 (
		\P2_IR_reg[18]/NET0131 ,
		_w1830_,
		_w1831_
	);
	LUT3 #(
		.INIT('h20)
	) name1369 (
		_w1505_,
		_w1508_,
		_w1831_,
		_w1832_
	);
	LUT4 #(
		.INIT('h00ab)
	) name1370 (
		_w1509_,
		_w1822_,
		_w1828_,
		_w1832_,
		_w1833_
	);
	LUT4 #(
		.INIT('h6333)
	) name1371 (
		\P2_reg3_reg[17]/NET0131 ,
		\P2_reg3_reg[18]/NET0131 ,
		_w467_,
		_w469_,
		_w1834_
	);
	LUT3 #(
		.INIT('h08)
	) name1372 (
		_w488_,
		_w494_,
		_w1834_,
		_w1835_
	);
	LUT3 #(
		.INIT('h20)
	) name1373 (
		\P2_reg1_reg[18]/NET0131 ,
		_w488_,
		_w494_,
		_w1836_
	);
	LUT4 #(
		.INIT('hff35)
	) name1374 (
		\P2_reg0_reg[18]/NET0131 ,
		\P2_reg2_reg[18]/NET0131 ,
		_w488_,
		_w494_,
		_w1837_
	);
	LUT3 #(
		.INIT('h10)
	) name1375 (
		_w1836_,
		_w1835_,
		_w1837_,
		_w1838_
	);
	LUT3 #(
		.INIT('hef)
	) name1376 (
		_w1836_,
		_w1835_,
		_w1837_,
		_w1839_
	);
	LUT2 #(
		.INIT('h8)
	) name1377 (
		_w1833_,
		_w1838_,
		_w1840_
	);
	LUT4 #(
		.INIT('h0777)
	) name1378 (
		_w1813_,
		_w1819_,
		_w1833_,
		_w1838_,
		_w1841_
	);
	LUT3 #(
		.INIT('h10)
	) name1379 (
		_w1783_,
		_w1796_,
		_w1841_,
		_w1842_
	);
	LUT2 #(
		.INIT('h8)
	) name1380 (
		_w1763_,
		_w1842_,
		_w1843_
	);
	LUT4 #(
		.INIT('hfee0)
	) name1381 (
		_w1735_,
		_w1746_,
		_w1751_,
		_w1761_,
		_w1844_
	);
	LUT2 #(
		.INIT('h1)
	) name1382 (
		_w1697_,
		_w1715_,
		_w1845_
	);
	LUT4 #(
		.INIT('heee8)
	) name1383 (
		_w1697_,
		_w1715_,
		_w1720_,
		_w1730_,
		_w1846_
	);
	LUT3 #(
		.INIT('hd0)
	) name1384 (
		_w1731_,
		_w1844_,
		_w1846_,
		_w1847_
	);
	LUT4 #(
		.INIT('h00f1)
	) name1385 (
		_w1509_,
		_w1771_,
		_w1775_,
		_w1781_,
		_w1848_
	);
	LUT4 #(
		.INIT('h5501)
	) name1386 (
		_w498_,
		_w1509_,
		_w1790_,
		_w1794_,
		_w1849_
	);
	LUT3 #(
		.INIT('h23)
	) name1387 (
		_w1783_,
		_w1848_,
		_w1849_,
		_w1850_
	);
	LUT4 #(
		.INIT('h7010)
	) name1388 (
		_w1776_,
		_w1781_,
		_w1841_,
		_w1849_,
		_w1851_
	);
	LUT2 #(
		.INIT('h1)
	) name1389 (
		_w1813_,
		_w1819_,
		_w1852_
	);
	LUT2 #(
		.INIT('h1)
	) name1390 (
		_w1833_,
		_w1838_,
		_w1853_
	);
	LUT4 #(
		.INIT('heee8)
	) name1391 (
		_w1813_,
		_w1819_,
		_w1833_,
		_w1838_,
		_w1854_
	);
	LUT2 #(
		.INIT('h4)
	) name1392 (
		_w1851_,
		_w1854_,
		_w1855_
	);
	LUT4 #(
		.INIT('h0d00)
	) name1393 (
		_w1842_,
		_w1847_,
		_w1851_,
		_w1854_,
		_w1856_
	);
	LUT4 #(
		.INIT('h4f00)
	) name1394 (
		_w1687_,
		_w1692_,
		_w1843_,
		_w1856_,
		_w1857_
	);
	LUT2 #(
		.INIT('h2)
	) name1395 (
		\P1_datao_reg[20]/NET0131 ,
		_w542_,
		_w1858_
	);
	LUT3 #(
		.INIT('h10)
	) name1396 (
		_w1766_,
		_w1798_,
		_w1800_,
		_w1859_
	);
	LUT4 #(
		.INIT('h8f00)
	) name1397 (
		_w1740_,
		_w1784_,
		_w1788_,
		_w1859_,
		_w1860_
	);
	LUT4 #(
		.INIT('hec80)
	) name1398 (
		\P1_datao_reg[18]/NET0131 ,
		\P1_datao_reg[19]/NET0131 ,
		\si[18]_pad ,
		\si[19]_pad ,
		_w1861_
	);
	LUT4 #(
		.INIT('h135f)
	) name1399 (
		\P1_datao_reg[16]/NET0131 ,
		\P1_datao_reg[17]/NET0131 ,
		\si[16]_pad ,
		\si[17]_pad ,
		_w1862_
	);
	LUT4 #(
		.INIT('h0f0b)
	) name1400 (
		_w1798_,
		_w1800_,
		_w1861_,
		_w1862_,
		_w1863_
	);
	LUT2 #(
		.INIT('h6)
	) name1401 (
		\P1_datao_reg[20]/NET0131 ,
		\si[20]_pad ,
		_w1864_
	);
	LUT4 #(
		.INIT('h208a)
	) name1402 (
		_w542_,
		_w1860_,
		_w1863_,
		_w1864_,
		_w1865_
	);
	LUT3 #(
		.INIT('h54)
	) name1403 (
		_w1509_,
		_w1858_,
		_w1865_,
		_w1866_
	);
	LUT4 #(
		.INIT('h0001)
	) name1404 (
		\P2_reg3_reg[17]/NET0131 ,
		\P2_reg3_reg[18]/NET0131 ,
		\P2_reg3_reg[19]/NET0131 ,
		\P2_reg3_reg[20]/NET0131 ,
		_w1867_
	);
	LUT3 #(
		.INIT('h80)
	) name1405 (
		_w467_,
		_w469_,
		_w1867_,
		_w1868_
	);
	LUT4 #(
		.INIT('h0073)
	) name1406 (
		\P2_reg3_reg[19]/NET0131 ,
		\P2_reg3_reg[20]/NET0131 ,
		_w1814_,
		_w1868_,
		_w1869_
	);
	LUT3 #(
		.INIT('h08)
	) name1407 (
		\P2_reg2_reg[20]/NET0131 ,
		_w488_,
		_w494_,
		_w1870_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name1408 (
		\P2_reg0_reg[20]/NET0131 ,
		\P2_reg1_reg[20]/NET0131 ,
		_w488_,
		_w494_,
		_w1871_
	);
	LUT4 #(
		.INIT('h3100)
	) name1409 (
		_w495_,
		_w1870_,
		_w1869_,
		_w1871_,
		_w1872_
	);
	LUT4 #(
		.INIT('hceff)
	) name1410 (
		_w495_,
		_w1870_,
		_w1869_,
		_w1871_,
		_w1873_
	);
	LUT4 #(
		.INIT('hab00)
	) name1411 (
		_w1509_,
		_w1858_,
		_w1865_,
		_w1872_,
		_w1874_
	);
	LUT4 #(
		.INIT('hfac8)
	) name1412 (
		\P1_datao_reg[19]/NET0131 ,
		\P1_datao_reg[20]/NET0131 ,
		\si[19]_pad ,
		\si[20]_pad ,
		_w1875_
	);
	LUT2 #(
		.INIT('h8)
	) name1413 (
		_w1800_,
		_w1875_,
		_w1876_
	);
	LUT4 #(
		.INIT('h8000)
	) name1414 (
		_w1703_,
		_w1767_,
		_w1800_,
		_w1875_,
		_w1877_
	);
	LUT4 #(
		.INIT('hec80)
	) name1415 (
		\P1_datao_reg[19]/NET0131 ,
		\P1_datao_reg[20]/NET0131 ,
		\si[19]_pad ,
		\si[20]_pad ,
		_w1878_
	);
	LUT3 #(
		.INIT('h07)
	) name1416 (
		_w1802_,
		_w1875_,
		_w1878_,
		_w1879_
	);
	LUT3 #(
		.INIT('hb0)
	) name1417 (
		_w1768_,
		_w1876_,
		_w1879_,
		_w1880_
	);
	LUT4 #(
		.INIT('h2f00)
	) name1418 (
		_w1755_,
		_w1757_,
		_w1877_,
		_w1880_,
		_w1881_
	);
	LUT4 #(
		.INIT('h9565)
	) name1419 (
		\P1_datao_reg[21]/NET0131 ,
		\si[21]_pad ,
		_w542_,
		_w1881_,
		_w1882_
	);
	LUT2 #(
		.INIT('h1)
	) name1420 (
		_w1509_,
		_w1882_,
		_w1883_
	);
	LUT4 #(
		.INIT('h4000)
	) name1421 (
		\P2_reg3_reg[21]/NET0131 ,
		_w467_,
		_w469_,
		_w1867_,
		_w1884_
	);
	LUT4 #(
		.INIT('h9555)
	) name1422 (
		\P2_reg3_reg[21]/NET0131 ,
		_w467_,
		_w469_,
		_w1867_,
		_w1885_
	);
	LUT3 #(
		.INIT('h08)
	) name1423 (
		_w488_,
		_w494_,
		_w1885_,
		_w1886_
	);
	LUT3 #(
		.INIT('h20)
	) name1424 (
		\P2_reg1_reg[21]/NET0131 ,
		_w488_,
		_w494_,
		_w1887_
	);
	LUT4 #(
		.INIT('hff35)
	) name1425 (
		\P2_reg0_reg[21]/NET0131 ,
		\P2_reg2_reg[21]/NET0131 ,
		_w488_,
		_w494_,
		_w1888_
	);
	LUT3 #(
		.INIT('h10)
	) name1426 (
		_w1887_,
		_w1886_,
		_w1888_,
		_w1889_
	);
	LUT3 #(
		.INIT('hef)
	) name1427 (
		_w1887_,
		_w1886_,
		_w1888_,
		_w1890_
	);
	LUT3 #(
		.INIT('he0)
	) name1428 (
		_w1509_,
		_w1882_,
		_w1889_,
		_w1891_
	);
	LUT2 #(
		.INIT('h8)
	) name1429 (
		\P1_datao_reg[23]/NET0131 ,
		\si[23]_pad ,
		_w1892_
	);
	LUT2 #(
		.INIT('h1)
	) name1430 (
		\P1_datao_reg[23]/NET0131 ,
		\si[23]_pad ,
		_w1893_
	);
	LUT4 #(
		.INIT('hfac8)
	) name1431 (
		\P1_datao_reg[21]/NET0131 ,
		\P1_datao_reg[22]/NET0131 ,
		\si[21]_pad ,
		\si[22]_pad ,
		_w1894_
	);
	LUT2 #(
		.INIT('h8)
	) name1432 (
		_w1875_,
		_w1894_,
		_w1895_
	);
	LUT4 #(
		.INIT('h8000)
	) name1433 (
		_w1767_,
		_w1800_,
		_w1875_,
		_w1894_,
		_w1896_
	);
	LUT2 #(
		.INIT('h8)
	) name1434 (
		\P1_datao_reg[22]/NET0131 ,
		\si[22]_pad ,
		_w1897_
	);
	LUT4 #(
		.INIT('hec80)
	) name1435 (
		\P1_datao_reg[21]/NET0131 ,
		\P1_datao_reg[22]/NET0131 ,
		\si[21]_pad ,
		\si[22]_pad ,
		_w1898_
	);
	LUT3 #(
		.INIT('h07)
	) name1436 (
		_w1878_,
		_w1894_,
		_w1898_,
		_w1899_
	);
	LUT3 #(
		.INIT('h40)
	) name1437 (
		_w1805_,
		_w1875_,
		_w1894_,
		_w1900_
	);
	LUT3 #(
		.INIT('h8c)
	) name1438 (
		_w1804_,
		_w1899_,
		_w1900_,
		_w1901_
	);
	LUT3 #(
		.INIT('hb0)
	) name1439 (
		_w1710_,
		_w1896_,
		_w1901_,
		_w1902_
	);
	LUT4 #(
		.INIT('h9565)
	) name1440 (
		\P1_datao_reg[23]/NET0131 ,
		\si[23]_pad ,
		_w542_,
		_w1902_,
		_w1903_
	);
	LUT3 #(
		.INIT('h63)
	) name1441 (
		\P2_reg3_reg[22]/NET0131 ,
		\P2_reg3_reg[23]/NET0131 ,
		_w1884_,
		_w1904_
	);
	LUT3 #(
		.INIT('h08)
	) name1442 (
		\P2_reg2_reg[23]/NET0131 ,
		_w488_,
		_w494_,
		_w1905_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name1443 (
		\P2_reg0_reg[23]/NET0131 ,
		\P2_reg1_reg[23]/NET0131 ,
		_w488_,
		_w494_,
		_w1906_
	);
	LUT4 #(
		.INIT('h3100)
	) name1444 (
		_w495_,
		_w1905_,
		_w1904_,
		_w1906_,
		_w1907_
	);
	LUT4 #(
		.INIT('hceff)
	) name1445 (
		_w495_,
		_w1905_,
		_w1904_,
		_w1906_,
		_w1908_
	);
	LUT3 #(
		.INIT('he0)
	) name1446 (
		_w1509_,
		_w1903_,
		_w1907_,
		_w1909_
	);
	LUT4 #(
		.INIT('hec80)
	) name1447 (
		\P1_datao_reg[20]/NET0131 ,
		\P1_datao_reg[21]/NET0131 ,
		\si[20]_pad ,
		\si[21]_pad ,
		_w1910_
	);
	LUT4 #(
		.INIT('hfac8)
	) name1448 (
		\P1_datao_reg[20]/NET0131 ,
		\P1_datao_reg[21]/NET0131 ,
		\si[20]_pad ,
		\si[21]_pad ,
		_w1911_
	);
	LUT3 #(
		.INIT('h13)
	) name1449 (
		_w1861_,
		_w1910_,
		_w1911_,
		_w1912_
	);
	LUT4 #(
		.INIT('hfac8)
	) name1450 (
		\P1_datao_reg[18]/NET0131 ,
		\P1_datao_reg[21]/NET0131 ,
		\si[18]_pad ,
		\si[21]_pad ,
		_w1913_
	);
	LUT2 #(
		.INIT('h8)
	) name1451 (
		_w1875_,
		_w1913_,
		_w1914_
	);
	LUT4 #(
		.INIT('h20f0)
	) name1452 (
		_w1825_,
		_w1827_,
		_w1912_,
		_w1914_,
		_w1915_
	);
	LUT4 #(
		.INIT('h9565)
	) name1453 (
		\P1_datao_reg[22]/NET0131 ,
		\si[22]_pad ,
		_w542_,
		_w1915_,
		_w1916_
	);
	LUT2 #(
		.INIT('h9)
	) name1454 (
		\P2_reg3_reg[22]/NET0131 ,
		_w1884_,
		_w1917_
	);
	LUT4 #(
		.INIT('h4080)
	) name1455 (
		\P2_reg3_reg[22]/NET0131 ,
		_w488_,
		_w494_,
		_w1884_,
		_w1918_
	);
	LUT3 #(
		.INIT('h20)
	) name1456 (
		\P2_reg1_reg[22]/NET0131 ,
		_w488_,
		_w494_,
		_w1919_
	);
	LUT4 #(
		.INIT('hff35)
	) name1457 (
		\P2_reg0_reg[22]/NET0131 ,
		\P2_reg2_reg[22]/NET0131 ,
		_w488_,
		_w494_,
		_w1920_
	);
	LUT3 #(
		.INIT('h10)
	) name1458 (
		_w1919_,
		_w1918_,
		_w1920_,
		_w1921_
	);
	LUT3 #(
		.INIT('hef)
	) name1459 (
		_w1919_,
		_w1918_,
		_w1920_,
		_w1922_
	);
	LUT3 #(
		.INIT('he0)
	) name1460 (
		_w1509_,
		_w1916_,
		_w1921_,
		_w1923_
	);
	LUT2 #(
		.INIT('h1)
	) name1461 (
		_w1909_,
		_w1923_,
		_w1924_
	);
	LUT4 #(
		.INIT('h0001)
	) name1462 (
		_w1874_,
		_w1891_,
		_w1909_,
		_w1923_,
		_w1925_
	);
	LUT2 #(
		.INIT('h2)
	) name1463 (
		\P1_datao_reg[25]/NET0131 ,
		_w542_,
		_w1926_
	);
	LUT2 #(
		.INIT('h6)
	) name1464 (
		\P1_datao_reg[25]/NET0131 ,
		\si[25]_pad ,
		_w1927_
	);
	LUT4 #(
		.INIT('hec80)
	) name1465 (
		\P1_datao_reg[23]/NET0131 ,
		\P1_datao_reg[24]/NET0131 ,
		\si[23]_pad ,
		\si[24]_pad ,
		_w1928_
	);
	LUT4 #(
		.INIT('hfac8)
	) name1466 (
		\P1_datao_reg[23]/NET0131 ,
		\P1_datao_reg[24]/NET0131 ,
		\si[23]_pad ,
		\si[24]_pad ,
		_w1929_
	);
	LUT3 #(
		.INIT('h13)
	) name1467 (
		_w1898_,
		_w1928_,
		_w1929_,
		_w1930_
	);
	LUT2 #(
		.INIT('h8)
	) name1468 (
		_w1894_,
		_w1929_,
		_w1931_
	);
	LUT4 #(
		.INIT('h7300)
	) name1469 (
		_w1755_,
		_w1768_,
		_w1769_,
		_w1876_,
		_w1932_
	);
	LUT2 #(
		.INIT('h2)
	) name1470 (
		_w1879_,
		_w1932_,
		_w1933_
	);
	LUT4 #(
		.INIT('h80f0)
	) name1471 (
		_w1757_,
		_w1877_,
		_w1931_,
		_w1933_,
		_w1934_
	);
	LUT4 #(
		.INIT('h2282)
	) name1472 (
		_w542_,
		_w1927_,
		_w1930_,
		_w1934_,
		_w1935_
	);
	LUT3 #(
		.INIT('h54)
	) name1473 (
		_w1509_,
		_w1926_,
		_w1935_,
		_w1936_
	);
	LUT4 #(
		.INIT('h0001)
	) name1474 (
		\P2_reg3_reg[21]/NET0131 ,
		\P2_reg3_reg[22]/NET0131 ,
		\P2_reg3_reg[23]/NET0131 ,
		\P2_reg3_reg[24]/NET0131 ,
		_w1937_
	);
	LUT4 #(
		.INIT('h8000)
	) name1475 (
		_w467_,
		_w469_,
		_w1867_,
		_w1937_,
		_w1938_
	);
	LUT2 #(
		.INIT('h9)
	) name1476 (
		\P2_reg3_reg[25]/NET0131 ,
		_w1938_,
		_w1939_
	);
	LUT4 #(
		.INIT('h4080)
	) name1477 (
		\P2_reg3_reg[25]/NET0131 ,
		_w488_,
		_w494_,
		_w1938_,
		_w1940_
	);
	LUT3 #(
		.INIT('h08)
	) name1478 (
		\P2_reg2_reg[25]/NET0131 ,
		_w488_,
		_w494_,
		_w1941_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name1479 (
		\P2_reg0_reg[25]/NET0131 ,
		\P2_reg1_reg[25]/NET0131 ,
		_w488_,
		_w494_,
		_w1942_
	);
	LUT3 #(
		.INIT('h10)
	) name1480 (
		_w1941_,
		_w1940_,
		_w1942_,
		_w1943_
	);
	LUT3 #(
		.INIT('hef)
	) name1481 (
		_w1941_,
		_w1940_,
		_w1942_,
		_w1944_
	);
	LUT4 #(
		.INIT('hab00)
	) name1482 (
		_w1509_,
		_w1926_,
		_w1935_,
		_w1943_,
		_w1945_
	);
	LUT4 #(
		.INIT('hfac8)
	) name1483 (
		\P1_datao_reg[22]/NET0131 ,
		\P1_datao_reg[23]/NET0131 ,
		\si[22]_pad ,
		\si[23]_pad ,
		_w1946_
	);
	LUT4 #(
		.INIT('h0155)
	) name1484 (
		_w1892_,
		_w1897_,
		_w1910_,
		_w1946_,
		_w1947_
	);
	LUT2 #(
		.INIT('h8)
	) name1485 (
		_w1911_,
		_w1946_,
		_w1948_
	);
	LUT4 #(
		.INIT('h4f00)
	) name1486 (
		_w1742_,
		_w1784_,
		_w1787_,
		_w1859_,
		_w1949_
	);
	LUT2 #(
		.INIT('h2)
	) name1487 (
		_w1863_,
		_w1949_,
		_w1950_
	);
	LUT4 #(
		.INIT('h7f00)
	) name1488 (
		_w1740_,
		_w1784_,
		_w1859_,
		_w1950_,
		_w1951_
	);
	LUT3 #(
		.INIT('ha2)
	) name1489 (
		_w1947_,
		_w1948_,
		_w1951_,
		_w1952_
	);
	LUT4 #(
		.INIT('h9565)
	) name1490 (
		\P1_datao_reg[24]/NET0131 ,
		\si[24]_pad ,
		_w542_,
		_w1952_,
		_w1953_
	);
	LUT4 #(
		.INIT('he0f0)
	) name1491 (
		\P2_reg3_reg[22]/NET0131 ,
		\P2_reg3_reg[23]/NET0131 ,
		\P2_reg3_reg[24]/NET0131 ,
		_w1884_,
		_w1954_
	);
	LUT2 #(
		.INIT('h1)
	) name1492 (
		_w1938_,
		_w1954_,
		_w1955_
	);
	LUT3 #(
		.INIT('ha8)
	) name1493 (
		_w495_,
		_w1938_,
		_w1954_,
		_w1956_
	);
	LUT3 #(
		.INIT('h08)
	) name1494 (
		\P2_reg2_reg[24]/NET0131 ,
		_w488_,
		_w494_,
		_w1957_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name1495 (
		\P2_reg0_reg[24]/NET0131 ,
		\P2_reg1_reg[24]/NET0131 ,
		_w488_,
		_w494_,
		_w1958_
	);
	LUT2 #(
		.INIT('h4)
	) name1496 (
		_w1957_,
		_w1958_,
		_w1959_
	);
	LUT2 #(
		.INIT('h4)
	) name1497 (
		_w1956_,
		_w1959_,
		_w1960_
	);
	LUT2 #(
		.INIT('hb)
	) name1498 (
		_w1956_,
		_w1959_,
		_w1961_
	);
	LUT4 #(
		.INIT('h0133)
	) name1499 (
		_w1509_,
		_w1945_,
		_w1953_,
		_w1960_,
		_w1962_
	);
	LUT2 #(
		.INIT('h1)
	) name1500 (
		\P1_datao_reg[27]/NET0131 ,
		\si[27]_pad ,
		_w1963_
	);
	LUT4 #(
		.INIT('hfac8)
	) name1501 (
		\P1_datao_reg[25]/NET0131 ,
		\P1_datao_reg[26]/NET0131 ,
		\si[25]_pad ,
		\si[26]_pad ,
		_w1964_
	);
	LUT4 #(
		.INIT('hec80)
	) name1502 (
		\P1_datao_reg[25]/NET0131 ,
		\P1_datao_reg[26]/NET0131 ,
		\si[25]_pad ,
		\si[26]_pad ,
		_w1965_
	);
	LUT3 #(
		.INIT('h07)
	) name1503 (
		_w1928_,
		_w1964_,
		_w1965_,
		_w1966_
	);
	LUT4 #(
		.INIT('h1f00)
	) name1504 (
		_w1806_,
		_w1807_,
		_w1895_,
		_w1899_,
		_w1967_
	);
	LUT2 #(
		.INIT('h8)
	) name1505 (
		_w1929_,
		_w1964_,
		_w1968_
	);
	LUT3 #(
		.INIT('h8a)
	) name1506 (
		_w1966_,
		_w1967_,
		_w1968_,
		_w1969_
	);
	LUT4 #(
		.INIT('h9565)
	) name1507 (
		\P1_datao_reg[27]/NET0131 ,
		\si[27]_pad ,
		_w542_,
		_w1969_,
		_w1970_
	);
	LUT3 #(
		.INIT('h10)
	) name1508 (
		\P2_reg3_reg[25]/NET0131 ,
		\P2_reg3_reg[26]/NET0131 ,
		_w1938_,
		_w1971_
	);
	LUT4 #(
		.INIT('h1e0f)
	) name1509 (
		\P2_reg3_reg[25]/NET0131 ,
		\P2_reg3_reg[26]/NET0131 ,
		\P2_reg3_reg[27]/NET0131 ,
		_w1938_,
		_w1972_
	);
	LUT3 #(
		.INIT('h20)
	) name1510 (
		\P2_reg1_reg[27]/NET0131 ,
		_w488_,
		_w494_,
		_w1973_
	);
	LUT4 #(
		.INIT('hff35)
	) name1511 (
		\P2_reg0_reg[27]/NET0131 ,
		\P2_reg2_reg[27]/NET0131 ,
		_w488_,
		_w494_,
		_w1974_
	);
	LUT4 #(
		.INIT('h3100)
	) name1512 (
		_w495_,
		_w1973_,
		_w1972_,
		_w1974_,
		_w1975_
	);
	LUT4 #(
		.INIT('hceff)
	) name1513 (
		_w495_,
		_w1973_,
		_w1972_,
		_w1974_,
		_w1976_
	);
	LUT3 #(
		.INIT('he0)
	) name1514 (
		_w1509_,
		_w1970_,
		_w1975_,
		_w1977_
	);
	LUT4 #(
		.INIT('hfac8)
	) name1515 (
		\P1_datao_reg[24]/NET0131 ,
		\P1_datao_reg[25]/NET0131 ,
		\si[24]_pad ,
		\si[25]_pad ,
		_w1978_
	);
	LUT2 #(
		.INIT('h8)
	) name1516 (
		_w1946_,
		_w1978_,
		_w1979_
	);
	LUT4 #(
		.INIT('hec80)
	) name1517 (
		\P1_datao_reg[24]/NET0131 ,
		\P1_datao_reg[25]/NET0131 ,
		\si[24]_pad ,
		\si[25]_pad ,
		_w1980_
	);
	LUT4 #(
		.INIT('h135f)
	) name1518 (
		\P1_datao_reg[22]/NET0131 ,
		\P1_datao_reg[23]/NET0131 ,
		\si[22]_pad ,
		\si[23]_pad ,
		_w1981_
	);
	LUT4 #(
		.INIT('h0f0b)
	) name1519 (
		_w1893_,
		_w1978_,
		_w1980_,
		_w1981_,
		_w1982_
	);
	LUT3 #(
		.INIT('hb0)
	) name1520 (
		_w1915_,
		_w1979_,
		_w1982_,
		_w1983_
	);
	LUT4 #(
		.INIT('h9565)
	) name1521 (
		\P1_datao_reg[26]/NET0131 ,
		\si[26]_pad ,
		_w542_,
		_w1983_,
		_w1984_
	);
	LUT3 #(
		.INIT('h63)
	) name1522 (
		\P2_reg3_reg[25]/NET0131 ,
		\P2_reg3_reg[26]/NET0131 ,
		_w1938_,
		_w1985_
	);
	LUT3 #(
		.INIT('h08)
	) name1523 (
		\P2_reg2_reg[26]/NET0131 ,
		_w488_,
		_w494_,
		_w1986_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name1524 (
		\P2_reg0_reg[26]/NET0131 ,
		\P2_reg1_reg[26]/NET0131 ,
		_w488_,
		_w494_,
		_w1987_
	);
	LUT4 #(
		.INIT('h3100)
	) name1525 (
		_w495_,
		_w1986_,
		_w1985_,
		_w1987_,
		_w1988_
	);
	LUT4 #(
		.INIT('hceff)
	) name1526 (
		_w495_,
		_w1986_,
		_w1985_,
		_w1987_,
		_w1989_
	);
	LUT3 #(
		.INIT('he0)
	) name1527 (
		_w1509_,
		_w1984_,
		_w1988_,
		_w1990_
	);
	LUT2 #(
		.INIT('h1)
	) name1528 (
		_w1977_,
		_w1990_,
		_w1991_
	);
	LUT3 #(
		.INIT('h02)
	) name1529 (
		_w1962_,
		_w1977_,
		_w1990_,
		_w1992_
	);
	LUT4 #(
		.INIT('h0008)
	) name1530 (
		_w1925_,
		_w1962_,
		_w1977_,
		_w1990_,
		_w1993_
	);
	LUT3 #(
		.INIT('h01)
	) name1531 (
		_w1509_,
		_w1984_,
		_w1988_,
		_w1994_
	);
	LUT4 #(
		.INIT('h0054)
	) name1532 (
		_w1509_,
		_w1926_,
		_w1935_,
		_w1943_,
		_w1995_
	);
	LUT4 #(
		.INIT('h0001)
	) name1533 (
		_w1509_,
		_w1945_,
		_w1953_,
		_w1960_,
		_w1996_
	);
	LUT3 #(
		.INIT('h01)
	) name1534 (
		_w1994_,
		_w1995_,
		_w1996_,
		_w1997_
	);
	LUT2 #(
		.INIT('h2)
	) name1535 (
		_w1991_,
		_w1997_,
		_w1998_
	);
	LUT3 #(
		.INIT('h01)
	) name1536 (
		_w1509_,
		_w1882_,
		_w1889_,
		_w1999_
	);
	LUT4 #(
		.INIT('h0054)
	) name1537 (
		_w1509_,
		_w1858_,
		_w1865_,
		_w1872_,
		_w2000_
	);
	LUT3 #(
		.INIT('h23)
	) name1538 (
		_w1891_,
		_w1999_,
		_w2000_,
		_w2001_
	);
	LUT3 #(
		.INIT('h01)
	) name1539 (
		_w1509_,
		_w1903_,
		_w1907_,
		_w2002_
	);
	LUT3 #(
		.INIT('h01)
	) name1540 (
		_w1509_,
		_w1916_,
		_w1921_,
		_w2003_
	);
	LUT3 #(
		.INIT('h23)
	) name1541 (
		_w1909_,
		_w2002_,
		_w2003_,
		_w2004_
	);
	LUT3 #(
		.INIT('hd0)
	) name1542 (
		_w1924_,
		_w2001_,
		_w2004_,
		_w2005_
	);
	LUT3 #(
		.INIT('h01)
	) name1543 (
		_w1509_,
		_w1970_,
		_w1975_,
		_w2006_
	);
	LUT3 #(
		.INIT('h0d)
	) name1544 (
		_w1992_,
		_w2005_,
		_w2006_,
		_w2007_
	);
	LUT4 #(
		.INIT('h0b00)
	) name1545 (
		_w1857_,
		_w1993_,
		_w1998_,
		_w2007_,
		_w2008_
	);
	LUT2 #(
		.INIT('h1)
	) name1546 (
		\P1_datao_reg[28]/NET0131 ,
		\si[28]_pad ,
		_w2009_
	);
	LUT2 #(
		.INIT('h8)
	) name1547 (
		\P1_datao_reg[28]/NET0131 ,
		\si[28]_pad ,
		_w2010_
	);
	LUT4 #(
		.INIT('hfac8)
	) name1548 (
		\P1_datao_reg[26]/NET0131 ,
		\P1_datao_reg[27]/NET0131 ,
		\si[26]_pad ,
		\si[27]_pad ,
		_w2011_
	);
	LUT4 #(
		.INIT('h8000)
	) name1549 (
		_w1911_,
		_w1946_,
		_w1978_,
		_w2011_,
		_w2012_
	);
	LUT4 #(
		.INIT('hf400)
	) name1550 (
		_w1947_,
		_w1978_,
		_w1980_,
		_w2011_,
		_w2013_
	);
	LUT4 #(
		.INIT('hec80)
	) name1551 (
		\P1_datao_reg[26]/NET0131 ,
		\P1_datao_reg[27]/NET0131 ,
		\si[26]_pad ,
		\si[27]_pad ,
		_w2014_
	);
	LUT2 #(
		.INIT('h1)
	) name1552 (
		_w2013_,
		_w2014_,
		_w2015_
	);
	LUT4 #(
		.INIT('h4f00)
	) name1553 (
		_w1860_,
		_w1863_,
		_w2012_,
		_w2015_,
		_w2016_
	);
	LUT4 #(
		.INIT('h9565)
	) name1554 (
		\P1_datao_reg[28]/NET0131 ,
		\si[28]_pad ,
		_w542_,
		_w2016_,
		_w2017_
	);
	LUT3 #(
		.INIT('h63)
	) name1555 (
		\P2_reg3_reg[27]/NET0131 ,
		\P2_reg3_reg[28]/NET0131 ,
		_w1971_,
		_w2018_
	);
	LUT4 #(
		.INIT('h90c0)
	) name1556 (
		\P2_reg3_reg[27]/NET0131 ,
		\P2_reg3_reg[28]/NET0131 ,
		_w495_,
		_w1971_,
		_w2019_
	);
	LUT3 #(
		.INIT('h02)
	) name1557 (
		\P2_reg0_reg[28]/NET0131 ,
		_w488_,
		_w494_,
		_w2020_
	);
	LUT4 #(
		.INIT('hf53f)
	) name1558 (
		\P2_reg1_reg[28]/NET0131 ,
		\P2_reg2_reg[28]/NET0131 ,
		_w488_,
		_w494_,
		_w2021_
	);
	LUT2 #(
		.INIT('h4)
	) name1559 (
		_w2020_,
		_w2021_,
		_w2022_
	);
	LUT2 #(
		.INIT('h4)
	) name1560 (
		_w2019_,
		_w2022_,
		_w2023_
	);
	LUT2 #(
		.INIT('hb)
	) name1561 (
		_w2019_,
		_w2022_,
		_w2024_
	);
	LUT3 #(
		.INIT('he0)
	) name1562 (
		_w1509_,
		_w2017_,
		_w2023_,
		_w2025_
	);
	LUT3 #(
		.INIT('h01)
	) name1563 (
		_w1509_,
		_w2017_,
		_w2023_,
		_w2026_
	);
	LUT3 #(
		.INIT('h1e)
	) name1564 (
		_w1509_,
		_w2017_,
		_w2023_,
		_w2027_
	);
	LUT4 #(
		.INIT('h1dd1)
	) name1565 (
		\P2_reg2_reg[28]/NET0131 ,
		_w1497_,
		_w2008_,
		_w2027_,
		_w2028_
	);
	LUT3 #(
		.INIT('h10)
	) name1566 (
		\P2_IR_reg[18]/NET0131 ,
		\P2_IR_reg[19]/NET0131 ,
		_w480_,
		_w2029_
	);
	LUT3 #(
		.INIT('h80)
	) name1567 (
		_w476_,
		_w478_,
		_w2029_,
		_w2030_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name1568 (
		\P2_IR_reg[31]/NET0131 ,
		_w476_,
		_w478_,
		_w2029_,
		_w2031_
	);
	LUT3 #(
		.INIT('he0)
	) name1569 (
		\P2_IR_reg[20]/NET0131 ,
		\P2_IR_reg[21]/NET0131 ,
		\P2_IR_reg[31]/NET0131 ,
		_w2032_
	);
	LUT3 #(
		.INIT('h56)
	) name1570 (
		\P2_IR_reg[22]/NET0131 ,
		_w2031_,
		_w2032_,
		_w2033_
	);
	LUT2 #(
		.INIT('h8)
	) name1571 (
		\P2_IR_reg[20]/NET0131 ,
		\P2_IR_reg[31]/NET0131 ,
		_w2034_
	);
	LUT3 #(
		.INIT('h56)
	) name1572 (
		\P2_IR_reg[21]/NET0131 ,
		_w2031_,
		_w2034_,
		_w2035_
	);
	LUT3 #(
		.INIT('ha6)
	) name1573 (
		\P2_IR_reg[20]/NET0131 ,
		\P2_IR_reg[31]/NET0131 ,
		_w2030_,
		_w2036_
	);
	LUT3 #(
		.INIT('h40)
	) name1574 (
		_w2033_,
		_w2035_,
		_w2036_,
		_w2037_
	);
	LUT4 #(
		.INIT('h3808)
	) name1575 (
		_w1811_,
		_w2033_,
		_w2035_,
		_w2036_,
		_w2038_
	);
	LUT3 #(
		.INIT('h0e)
	) name1576 (
		_w1491_,
		_w1493_,
		_w1496_,
		_w2039_
	);
	LUT4 #(
		.INIT('haa02)
	) name1577 (
		\P2_reg2_reg[28]/NET0131 ,
		_w1491_,
		_w1493_,
		_w1496_,
		_w2040_
	);
	LUT2 #(
		.INIT('h4)
	) name1578 (
		_w1505_,
		_w1508_,
		_w2041_
	);
	LUT2 #(
		.INIT('h9)
	) name1579 (
		_w1505_,
		_w1508_,
		_w2042_
	);
	LUT2 #(
		.INIT('h4)
	) name1580 (
		_w1975_,
		_w2042_,
		_w2043_
	);
	LUT4 #(
		.INIT('h0001)
	) name1581 (
		\P2_reg3_reg[25]/NET0131 ,
		\P2_reg3_reg[26]/NET0131 ,
		\P2_reg3_reg[27]/NET0131 ,
		\P2_reg3_reg[28]/NET0131 ,
		_w2044_
	);
	LUT3 #(
		.INIT('h80)
	) name1582 (
		_w1867_,
		_w1937_,
		_w2044_,
		_w2045_
	);
	LUT4 #(
		.INIT('h0800)
	) name1583 (
		_w467_,
		_w469_,
		_w1748_,
		_w2045_,
		_w2046_
	);
	LUT4 #(
		.INIT('h3dfd)
	) name1584 (
		\P2_reg0_reg[29]/NET0131 ,
		_w488_,
		_w494_,
		_w2046_,
		_w2047_
	);
	LUT4 #(
		.INIT('hf53f)
	) name1585 (
		\P2_reg1_reg[29]/NET0131 ,
		\P2_reg2_reg[29]/NET0131 ,
		_w488_,
		_w494_,
		_w2048_
	);
	LUT2 #(
		.INIT('h8)
	) name1586 (
		_w2047_,
		_w2048_,
		_w2049_
	);
	LUT2 #(
		.INIT('h7)
	) name1587 (
		_w2047_,
		_w2048_,
		_w2050_
	);
	LUT4 #(
		.INIT('h37f7)
	) name1588 (
		\P2_reg2_reg[31]/NET0131 ,
		_w488_,
		_w494_,
		_w2046_,
		_w2051_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name1589 (
		\P2_reg0_reg[31]/NET0131 ,
		\P2_reg1_reg[31]/NET0131 ,
		_w488_,
		_w494_,
		_w2052_
	);
	LUT2 #(
		.INIT('h8)
	) name1590 (
		_w2051_,
		_w2052_,
		_w2053_
	);
	LUT2 #(
		.INIT('h7)
	) name1591 (
		_w2051_,
		_w2052_,
		_w2054_
	);
	LUT4 #(
		.INIT('h0777)
	) name1592 (
		_w1576_,
		_w1577_,
		_w2051_,
		_w2052_,
		_w2055_
	);
	LUT3 #(
		.INIT('h10)
	) name1593 (
		_w1559_,
		_w1569_,
		_w2055_,
		_w2056_
	);
	LUT4 #(
		.INIT('h0100)
	) name1594 (
		_w1550_,
		_w1559_,
		_w1569_,
		_w2055_,
		_w2057_
	);
	LUT4 #(
		.INIT('h0777)
	) name1595 (
		_w1499_,
		_w1501_,
		_w1529_,
		_w1531_,
		_w2058_
	);
	LUT4 #(
		.INIT('h0777)
	) name1596 (
		_w1583_,
		_w1585_,
		_w1597_,
		_w1598_,
		_w2059_
	);
	LUT2 #(
		.INIT('h8)
	) name1597 (
		_w2058_,
		_w2059_,
		_w2060_
	);
	LUT4 #(
		.INIT('h0777)
	) name1598 (
		_w1616_,
		_w1618_,
		_w1644_,
		_w1645_,
		_w2061_
	);
	LUT4 #(
		.INIT('h0777)
	) name1599 (
		_w1661_,
		_w1662_,
		_w1673_,
		_w1675_,
		_w2062_
	);
	LUT4 #(
		.INIT('h0777)
	) name1600 (
		_w1733_,
		_w1734_,
		_w1747_,
		_w1750_,
		_w2063_
	);
	LUT3 #(
		.INIT('h80)
	) name1601 (
		_w2061_,
		_w2062_,
		_w2063_,
		_w2064_
	);
	LUT3 #(
		.INIT('h80)
	) name1602 (
		_w2057_,
		_w2060_,
		_w2064_,
		_w2065_
	);
	LUT4 #(
		.INIT('h4000)
	) name1603 (
		_w1720_,
		_w2057_,
		_w2060_,
		_w2064_,
		_w2066_
	);
	LUT2 #(
		.INIT('h1)
	) name1604 (
		_w498_,
		_w1781_,
		_w2067_
	);
	LUT3 #(
		.INIT('h01)
	) name1605 (
		_w498_,
		_w1781_,
		_w1838_,
		_w2068_
	);
	LUT3 #(
		.INIT('h40)
	) name1606 (
		_w1697_,
		_w2066_,
		_w2068_,
		_w2069_
	);
	LUT2 #(
		.INIT('h1)
	) name1607 (
		_w1872_,
		_w1889_,
		_w2070_
	);
	LUT3 #(
		.INIT('h01)
	) name1608 (
		_w1819_,
		_w1907_,
		_w1921_,
		_w2071_
	);
	LUT3 #(
		.INIT('h40)
	) name1609 (
		_w1960_,
		_w2070_,
		_w2071_,
		_w2072_
	);
	LUT4 #(
		.INIT('h4000)
	) name1610 (
		_w1697_,
		_w2066_,
		_w2068_,
		_w2072_,
		_w2073_
	);
	LUT3 #(
		.INIT('h01)
	) name1611 (
		_w1943_,
		_w1975_,
		_w1988_,
		_w2074_
	);
	LUT4 #(
		.INIT('hbf00)
	) name1612 (
		_w2023_,
		_w2073_,
		_w2074_,
		_w2049_,
		_w2075_
	);
	LUT3 #(
		.INIT('h0b)
	) name1613 (
		_w2019_,
		_w2022_,
		_w2049_,
		_w2076_
	);
	LUT3 #(
		.INIT('h80)
	) name1614 (
		_w2073_,
		_w2074_,
		_w2076_,
		_w2077_
	);
	LUT4 #(
		.INIT('h1555)
	) name1615 (
		_w2042_,
		_w2073_,
		_w2074_,
		_w2076_,
		_w2078_
	);
	LUT4 #(
		.INIT('h8a88)
	) name1616 (
		_w2039_,
		_w2043_,
		_w2075_,
		_w2078_,
		_w2079_
	);
	LUT2 #(
		.INIT('h8)
	) name1617 (
		_w2033_,
		_w2035_,
		_w2080_
	);
	LUT4 #(
		.INIT('h0040)
	) name1618 (
		_w1811_,
		_w2033_,
		_w2035_,
		_w2036_,
		_w2081_
	);
	LUT2 #(
		.INIT('h2)
	) name1619 (
		_w1811_,
		_w2036_,
		_w2082_
	);
	LUT2 #(
		.INIT('h1)
	) name1620 (
		_w2033_,
		_w2035_,
		_w2083_
	);
	LUT4 #(
		.INIT('h0301)
	) name1621 (
		_w1811_,
		_w2033_,
		_w2035_,
		_w2036_,
		_w2084_
	);
	LUT4 #(
		.INIT('h1000)
	) name1622 (
		_w1491_,
		_w1493_,
		_w1496_,
		_w2084_,
		_w2085_
	);
	LUT4 #(
		.INIT('hc080)
	) name1623 (
		_w1811_,
		_w2033_,
		_w2035_,
		_w2036_,
		_w2086_
	);
	LUT4 #(
		.INIT('hef00)
	) name1624 (
		_w1491_,
		_w1493_,
		_w1496_,
		_w2084_,
		_w2087_
	);
	LUT4 #(
		.INIT('h0002)
	) name1625 (
		_w1811_,
		_w2033_,
		_w2035_,
		_w2036_,
		_w2088_
	);
	LUT4 #(
		.INIT('h9c00)
	) name1626 (
		\P2_reg3_reg[27]/NET0131 ,
		\P2_reg3_reg[28]/NET0131 ,
		_w1971_,
		_w2088_,
		_w2089_
	);
	LUT4 #(
		.INIT('h0057)
	) name1627 (
		\P2_reg2_reg[28]/NET0131 ,
		_w2086_,
		_w2087_,
		_w2089_,
		_w2090_
	);
	LUT4 #(
		.INIT('hef00)
	) name1628 (
		_w1509_,
		_w2017_,
		_w2085_,
		_w2090_,
		_w2091_
	);
	LUT4 #(
		.INIT('h1f00)
	) name1629 (
		_w2040_,
		_w2079_,
		_w2081_,
		_w2091_,
		_w2092_
	);
	LUT3 #(
		.INIT('hb0)
	) name1630 (
		_w2028_,
		_w2038_,
		_w2092_,
		_w2093_
	);
	LUT3 #(
		.INIT('h08)
	) name1631 (
		_w1644_,
		_w1645_,
		_w1657_,
		_w2094_
	);
	LUT4 #(
		.INIT('h8880)
	) name1632 (
		_w1616_,
		_w1618_,
		_w1638_,
		_w1640_,
		_w2095_
	);
	LUT2 #(
		.INIT('h1)
	) name1633 (
		_w2094_,
		_w2095_,
		_w2096_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name1634 (
		_w1663_,
		_w1672_,
		_w1676_,
		_w1684_,
		_w2097_
	);
	LUT4 #(
		.INIT('h4d44)
	) name1635 (
		_w1663_,
		_w1672_,
		_w1676_,
		_w1684_,
		_w2098_
	);
	LUT4 #(
		.INIT('h0007)
	) name1636 (
		_w1616_,
		_w1618_,
		_w1638_,
		_w1640_,
		_w2099_
	);
	LUT3 #(
		.INIT('h70)
	) name1637 (
		_w1644_,
		_w1645_,
		_w1657_,
		_w2100_
	);
	LUT3 #(
		.INIT('h54)
	) name1638 (
		_w2095_,
		_w2099_,
		_w2100_,
		_w2101_
	);
	LUT3 #(
		.INIT('h07)
	) name1639 (
		_w2096_,
		_w2098_,
		_w2101_,
		_w2102_
	);
	LUT3 #(
		.INIT('h08)
	) name1640 (
		_w1529_,
		_w1531_,
		_w1545_,
		_w2103_
	);
	LUT3 #(
		.INIT('h08)
	) name1641 (
		_w1499_,
		_w1501_,
		_w1527_,
		_w2104_
	);
	LUT2 #(
		.INIT('h1)
	) name1642 (
		_w2103_,
		_w2104_,
		_w2105_
	);
	LUT3 #(
		.INIT('h08)
	) name1643 (
		_w1583_,
		_w1585_,
		_w1593_,
		_w2106_
	);
	LUT3 #(
		.INIT('h08)
	) name1644 (
		_w1597_,
		_w1598_,
		_w1604_,
		_w2107_
	);
	LUT2 #(
		.INIT('h1)
	) name1645 (
		_w2106_,
		_w2107_,
		_w2108_
	);
	LUT3 #(
		.INIT('h08)
	) name1646 (
		_w1548_,
		_w1549_,
		_w1555_,
		_w2109_
	);
	LUT3 #(
		.INIT('h08)
	) name1647 (
		_w1557_,
		_w1558_,
		_w1564_,
		_w2110_
	);
	LUT2 #(
		.INIT('h1)
	) name1648 (
		_w2109_,
		_w2110_,
		_w2111_
	);
	LUT3 #(
		.INIT('h08)
	) name1649 (
		_w1576_,
		_w1577_,
		_w1580_,
		_w2112_
	);
	LUT3 #(
		.INIT('hb2)
	) name1650 (
		_w1569_,
		_w1573_,
		_w2112_,
		_w2113_
	);
	LUT3 #(
		.INIT('h70)
	) name1651 (
		_w1548_,
		_w1549_,
		_w1555_,
		_w2114_
	);
	LUT3 #(
		.INIT('h70)
	) name1652 (
		_w1557_,
		_w1558_,
		_w1564_,
		_w2115_
	);
	LUT3 #(
		.INIT('h54)
	) name1653 (
		_w2109_,
		_w2114_,
		_w2115_,
		_w2116_
	);
	LUT4 #(
		.INIT('haa08)
	) name1654 (
		_w2108_,
		_w2111_,
		_w2113_,
		_w2116_,
		_w2117_
	);
	LUT3 #(
		.INIT('h70)
	) name1655 (
		_w1583_,
		_w1585_,
		_w1593_,
		_w2118_
	);
	LUT3 #(
		.INIT('h70)
	) name1656 (
		_w1597_,
		_w1598_,
		_w1604_,
		_w2119_
	);
	LUT3 #(
		.INIT('h23)
	) name1657 (
		_w2106_,
		_w2118_,
		_w2119_,
		_w2120_
	);
	LUT3 #(
		.INIT('h70)
	) name1658 (
		_w1529_,
		_w1531_,
		_w1545_,
		_w2121_
	);
	LUT3 #(
		.INIT('h70)
	) name1659 (
		_w1499_,
		_w1501_,
		_w1527_,
		_w2122_
	);
	LUT3 #(
		.INIT('h54)
	) name1660 (
		_w2103_,
		_w2121_,
		_w2122_,
		_w2123_
	);
	LUT4 #(
		.INIT('h0075)
	) name1661 (
		_w2105_,
		_w2117_,
		_w2120_,
		_w2123_,
		_w2124_
	);
	LUT4 #(
		.INIT('hdd0d)
	) name1662 (
		_w1663_,
		_w1672_,
		_w1676_,
		_w1684_,
		_w2125_
	);
	LUT2 #(
		.INIT('h8)
	) name1663 (
		_w2096_,
		_w2125_,
		_w2126_
	);
	LUT2 #(
		.INIT('h2)
	) name1664 (
		_w1697_,
		_w1715_,
		_w2127_
	);
	LUT4 #(
		.INIT('hdd0d)
	) name1665 (
		_w1697_,
		_w1715_,
		_w1720_,
		_w1730_,
		_w2128_
	);
	LUT4 #(
		.INIT('hdd0d)
	) name1666 (
		_w1735_,
		_w1746_,
		_w1751_,
		_w1761_,
		_w2129_
	);
	LUT2 #(
		.INIT('h8)
	) name1667 (
		_w2128_,
		_w2129_,
		_w2130_
	);
	LUT4 #(
		.INIT('hf100)
	) name1668 (
		_w1509_,
		_w1771_,
		_w1775_,
		_w1781_,
		_w2131_
	);
	LUT4 #(
		.INIT('haa02)
	) name1669 (
		_w498_,
		_w1509_,
		_w1790_,
		_w1794_,
		_w2132_
	);
	LUT2 #(
		.INIT('h4)
	) name1670 (
		_w1833_,
		_w1838_,
		_w2133_
	);
	LUT2 #(
		.INIT('h4)
	) name1671 (
		_w1813_,
		_w1819_,
		_w2134_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name1672 (
		_w1813_,
		_w1819_,
		_w1833_,
		_w1838_,
		_w2135_
	);
	LUT3 #(
		.INIT('h10)
	) name1673 (
		_w2131_,
		_w2132_,
		_w2135_,
		_w2136_
	);
	LUT2 #(
		.INIT('h8)
	) name1674 (
		_w2130_,
		_w2136_,
		_w2137_
	);
	LUT4 #(
		.INIT('h7500)
	) name1675 (
		_w2102_,
		_w2124_,
		_w2126_,
		_w2137_,
		_w2138_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name1676 (
		_w1735_,
		_w1746_,
		_w1751_,
		_w1761_,
		_w2139_
	);
	LUT4 #(
		.INIT('h4f04)
	) name1677 (
		_w1735_,
		_w1746_,
		_w1751_,
		_w1761_,
		_w2140_
	);
	LUT2 #(
		.INIT('h4)
	) name1678 (
		_w1697_,
		_w1715_,
		_w2141_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name1679 (
		_w1697_,
		_w1715_,
		_w1720_,
		_w1730_,
		_w2142_
	);
	LUT4 #(
		.INIT('h4d44)
	) name1680 (
		_w1697_,
		_w1715_,
		_w1720_,
		_w1730_,
		_w2143_
	);
	LUT3 #(
		.INIT('h07)
	) name1681 (
		_w2128_,
		_w2140_,
		_w2143_,
		_w2144_
	);
	LUT4 #(
		.INIT('h0054)
	) name1682 (
		_w498_,
		_w1509_,
		_w1790_,
		_w1794_,
		_w2145_
	);
	LUT4 #(
		.INIT('h000e)
	) name1683 (
		_w1509_,
		_w1771_,
		_w1775_,
		_w1781_,
		_w2146_
	);
	LUT2 #(
		.INIT('h1)
	) name1684 (
		_w2145_,
		_w2146_,
		_w2147_
	);
	LUT3 #(
		.INIT('h54)
	) name1685 (
		_w2131_,
		_w2145_,
		_w2146_,
		_w2148_
	);
	LUT4 #(
		.INIT('hb020)
	) name1686 (
		_w1776_,
		_w1781_,
		_w2135_,
		_w2145_,
		_w2149_
	);
	LUT2 #(
		.INIT('h2)
	) name1687 (
		_w1813_,
		_w1819_,
		_w2150_
	);
	LUT2 #(
		.INIT('h2)
	) name1688 (
		_w1833_,
		_w1838_,
		_w2151_
	);
	LUT4 #(
		.INIT('hdd0d)
	) name1689 (
		_w1813_,
		_w1819_,
		_w1833_,
		_w1838_,
		_w2152_
	);
	LUT4 #(
		.INIT('h22b2)
	) name1690 (
		_w1813_,
		_w1819_,
		_w1833_,
		_w1838_,
		_w2153_
	);
	LUT2 #(
		.INIT('h1)
	) name1691 (
		_w2149_,
		_w2153_,
		_w2154_
	);
	LUT4 #(
		.INIT('h000d)
	) name1692 (
		_w2136_,
		_w2144_,
		_w2149_,
		_w2153_,
		_w2155_
	);
	LUT4 #(
		.INIT('h5400)
	) name1693 (
		_w1509_,
		_w1858_,
		_w1865_,
		_w1872_,
		_w2156_
	);
	LUT3 #(
		.INIT('h10)
	) name1694 (
		_w1509_,
		_w1882_,
		_w1889_,
		_w2157_
	);
	LUT3 #(
		.INIT('h10)
	) name1695 (
		_w1509_,
		_w1916_,
		_w1921_,
		_w2158_
	);
	LUT3 #(
		.INIT('h10)
	) name1696 (
		_w1509_,
		_w1903_,
		_w1907_,
		_w2159_
	);
	LUT2 #(
		.INIT('h1)
	) name1697 (
		_w2158_,
		_w2159_,
		_w2160_
	);
	LUT4 #(
		.INIT('h0001)
	) name1698 (
		_w2156_,
		_w2157_,
		_w2158_,
		_w2159_,
		_w2161_
	);
	LUT3 #(
		.INIT('h10)
	) name1699 (
		_w1509_,
		_w1953_,
		_w1960_,
		_w2162_
	);
	LUT4 #(
		.INIT('h5400)
	) name1700 (
		_w1509_,
		_w1926_,
		_w1935_,
		_w1943_,
		_w2163_
	);
	LUT4 #(
		.INIT('h00ef)
	) name1701 (
		_w1509_,
		_w1953_,
		_w1960_,
		_w2163_,
		_w2164_
	);
	LUT3 #(
		.INIT('h10)
	) name1702 (
		_w1509_,
		_w1984_,
		_w1988_,
		_w2165_
	);
	LUT3 #(
		.INIT('h10)
	) name1703 (
		_w1509_,
		_w1970_,
		_w1975_,
		_w2166_
	);
	LUT3 #(
		.INIT('h02)
	) name1704 (
		_w2164_,
		_w2165_,
		_w2166_,
		_w2167_
	);
	LUT4 #(
		.INIT('h0008)
	) name1705 (
		_w2161_,
		_w2164_,
		_w2165_,
		_w2166_,
		_w2168_
	);
	LUT3 #(
		.INIT('hb0)
	) name1706 (
		_w2138_,
		_w2155_,
		_w2168_,
		_w2169_
	);
	LUT4 #(
		.INIT('h00ab)
	) name1707 (
		_w1509_,
		_w1858_,
		_w1865_,
		_w1872_,
		_w2170_
	);
	LUT3 #(
		.INIT('h0e)
	) name1708 (
		_w1509_,
		_w1882_,
		_w1889_,
		_w2171_
	);
	LUT2 #(
		.INIT('h1)
	) name1709 (
		_w2170_,
		_w2171_,
		_w2172_
	);
	LUT3 #(
		.INIT('h54)
	) name1710 (
		_w2157_,
		_w2170_,
		_w2171_,
		_w2173_
	);
	LUT3 #(
		.INIT('h0e)
	) name1711 (
		_w1509_,
		_w1916_,
		_w1921_,
		_w2174_
	);
	LUT3 #(
		.INIT('h0e)
	) name1712 (
		_w1509_,
		_w1903_,
		_w1907_,
		_w2175_
	);
	LUT3 #(
		.INIT('h54)
	) name1713 (
		_w2159_,
		_w2174_,
		_w2175_,
		_w2176_
	);
	LUT3 #(
		.INIT('h07)
	) name1714 (
		_w2160_,
		_w2173_,
		_w2176_,
		_w2177_
	);
	LUT2 #(
		.INIT('h2)
	) name1715 (
		_w2167_,
		_w2177_,
		_w2178_
	);
	LUT3 #(
		.INIT('h0e)
	) name1716 (
		_w1509_,
		_w1984_,
		_w1988_,
		_w2179_
	);
	LUT3 #(
		.INIT('h0e)
	) name1717 (
		_w1509_,
		_w1970_,
		_w1975_,
		_w2180_
	);
	LUT2 #(
		.INIT('h1)
	) name1718 (
		_w2179_,
		_w2180_,
		_w2181_
	);
	LUT4 #(
		.INIT('h00ab)
	) name1719 (
		_w1509_,
		_w1926_,
		_w1935_,
		_w1943_,
		_w2182_
	);
	LUT4 #(
		.INIT('h00f1)
	) name1720 (
		_w1509_,
		_w1953_,
		_w1960_,
		_w2182_,
		_w2183_
	);
	LUT3 #(
		.INIT('h01)
	) name1721 (
		_w2163_,
		_w2165_,
		_w2183_,
		_w2184_
	);
	LUT3 #(
		.INIT('h51)
	) name1722 (
		_w2166_,
		_w2181_,
		_w2184_,
		_w2185_
	);
	LUT2 #(
		.INIT('h1)
	) name1723 (
		_w2178_,
		_w2185_,
		_w2186_
	);
	LUT4 #(
		.INIT('h8488)
	) name1724 (
		_w2027_,
		_w2039_,
		_w2169_,
		_w2186_,
		_w2187_
	);
	LUT4 #(
		.INIT('h0400)
	) name1725 (
		_w1811_,
		_w2033_,
		_w2035_,
		_w2036_,
		_w2188_
	);
	LUT3 #(
		.INIT('he0)
	) name1726 (
		_w2040_,
		_w2187_,
		_w2188_,
		_w2189_
	);
	LUT4 #(
		.INIT('h8288)
	) name1727 (
		_w1497_,
		_w2027_,
		_w2169_,
		_w2186_,
		_w2190_
	);
	LUT3 #(
		.INIT('h04)
	) name1728 (
		_w2033_,
		_w2035_,
		_w2036_,
		_w2191_
	);
	LUT4 #(
		.INIT('hfbcb)
	) name1729 (
		_w1811_,
		_w2033_,
		_w2035_,
		_w2036_,
		_w2192_
	);
	LUT4 #(
		.INIT('h0034)
	) name1730 (
		_w1811_,
		_w2033_,
		_w2035_,
		_w2036_,
		_w2193_
	);
	LUT3 #(
		.INIT('he0)
	) name1731 (
		_w1498_,
		_w2190_,
		_w2193_,
		_w2194_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name1732 (
		_w1489_,
		_w2189_,
		_w2194_,
		_w2093_,
		_w2195_
	);
	LUT4 #(
		.INIT('heeec)
	) name1733 (
		\P1_state_reg[0]/NET0131 ,
		_w1479_,
		_w1488_,
		_w2195_,
		_w2196_
	);
	LUT3 #(
		.INIT('he0)
	) name1734 (
		_w528_,
		_w530_,
		_w533_,
		_w2197_
	);
	LUT2 #(
		.INIT('h1)
	) name1735 (
		_w1019_,
		_w2197_,
		_w2198_
	);
	LUT4 #(
		.INIT('h22a2)
	) name1736 (
		_w1340_,
		_w1345_,
		_w1353_,
		_w1387_,
		_w2199_
	);
	LUT2 #(
		.INIT('h8)
	) name1737 (
		_w1322_,
		_w1338_,
		_w2200_
	);
	LUT3 #(
		.INIT('hd0)
	) name1738 (
		_w1333_,
		_w2199_,
		_w2200_,
		_w2201_
	);
	LUT2 #(
		.INIT('h2)
	) name1739 (
		_w1322_,
		_w1327_,
		_w2202_
	);
	LUT2 #(
		.INIT('h1)
	) name1740 (
		_w1321_,
		_w2202_,
		_w2203_
	);
	LUT4 #(
		.INIT('h8488)
	) name1741 (
		_w1419_,
		_w2197_,
		_w2201_,
		_w2203_,
		_w2204_
	);
	LUT3 #(
		.INIT('ha8)
	) name1742 (
		_w1286_,
		_w2198_,
		_w2204_,
		_w2205_
	);
	LUT4 #(
		.INIT('h1444)
	) name1743 (
		_w537_,
		_w643_,
		_w1172_,
		_w1174_,
		_w2206_
	);
	LUT3 #(
		.INIT('h20)
	) name1744 (
		_w537_,
		_w1036_,
		_w1039_,
		_w2207_
	);
	LUT4 #(
		.INIT('h3331)
	) name1745 (
		_w2197_,
		_w2198_,
		_w2206_,
		_w2207_,
		_w2208_
	);
	LUT3 #(
		.INIT('h15)
	) name1746 (
		_w681_,
		_w738_,
		_w745_,
		_w2209_
	);
	LUT4 #(
		.INIT('h0777)
	) name1747 (
		_w717_,
		_w722_,
		_w786_,
		_w791_,
		_w2210_
	);
	LUT4 #(
		.INIT('h1500)
	) name1748 (
		_w681_,
		_w738_,
		_w745_,
		_w2210_,
		_w2211_
	);
	LUT4 #(
		.INIT('h0777)
	) name1749 (
		_w762_,
		_w767_,
		_w772_,
		_w780_,
		_w2212_
	);
	LUT4 #(
		.INIT('h0777)
	) name1750 (
		_w752_,
		_w758_,
		_w808_,
		_w814_,
		_w2213_
	);
	LUT2 #(
		.INIT('h8)
	) name1751 (
		_w2212_,
		_w2213_,
		_w2214_
	);
	LUT2 #(
		.INIT('h8)
	) name1752 (
		_w2211_,
		_w2214_,
		_w2215_
	);
	LUT3 #(
		.INIT('h07)
	) name1753 (
		_w799_,
		_w804_,
		_w828_,
		_w2216_
	);
	LUT3 #(
		.INIT('h51)
	) name1754 (
		_w843_,
		_w946_,
		_w950_,
		_w2217_
	);
	LUT3 #(
		.INIT('h8e)
	) name1755 (
		_w799_,
		_w804_,
		_w829_,
		_w2218_
	);
	LUT3 #(
		.INIT('hd0)
	) name1756 (
		_w2216_,
		_w2217_,
		_w2218_,
		_w2219_
	);
	LUT3 #(
		.INIT('h0d)
	) name1757 (
		_w854_,
		_w882_,
		_w898_,
		_w2220_
	);
	LUT2 #(
		.INIT('h1)
	) name1758 (
		_w919_,
		_w930_,
		_w2221_
	);
	LUT2 #(
		.INIT('h1)
	) name1759 (
		_w895_,
		_w939_,
		_w2222_
	);
	LUT4 #(
		.INIT('h0001)
	) name1760 (
		_w895_,
		_w919_,
		_w930_,
		_w939_,
		_w2223_
	);
	LUT4 #(
		.INIT('h8f00)
	) name1761 (
		_w871_,
		_w883_,
		_w2220_,
		_w2223_,
		_w2224_
	);
	LUT3 #(
		.INIT('h0d)
	) name1762 (
		_w897_,
		_w939_,
		_w944_,
		_w2225_
	);
	LUT3 #(
		.INIT('h0b)
	) name1763 (
		_w919_,
		_w943_,
		_w947_,
		_w2226_
	);
	LUT3 #(
		.INIT('hd0)
	) name1764 (
		_w2221_,
		_w2225_,
		_w2226_,
		_w2227_
	);
	LUT2 #(
		.INIT('h1)
	) name1765 (
		_w908_,
		_w950_,
		_w2228_
	);
	LUT2 #(
		.INIT('h8)
	) name1766 (
		_w2216_,
		_w2228_,
		_w2229_
	);
	LUT3 #(
		.INIT('hb0)
	) name1767 (
		_w2224_,
		_w2227_,
		_w2229_,
		_w2230_
	);
	LUT4 #(
		.INIT('h20aa)
	) name1768 (
		_w2219_,
		_w2224_,
		_w2227_,
		_w2229_,
		_w2231_
	);
	LUT4 #(
		.INIT('heee8)
	) name1769 (
		_w752_,
		_w758_,
		_w808_,
		_w814_,
		_w2232_
	);
	LUT4 #(
		.INIT('hfee0)
	) name1770 (
		_w762_,
		_w767_,
		_w772_,
		_w780_,
		_w2233_
	);
	LUT3 #(
		.INIT('hd0)
	) name1771 (
		_w2212_,
		_w2232_,
		_w2233_,
		_w2234_
	);
	LUT4 #(
		.INIT('h1117)
	) name1772 (
		_w717_,
		_w722_,
		_w786_,
		_w791_,
		_w2235_
	);
	LUT4 #(
		.INIT('h1500)
	) name1773 (
		_w681_,
		_w738_,
		_w745_,
		_w2235_,
		_w2236_
	);
	LUT4 #(
		.INIT('h00fe)
	) name1774 (
		_w681_,
		_w738_,
		_w745_,
		_w962_,
		_w2237_
	);
	LUT2 #(
		.INIT('h4)
	) name1775 (
		_w2236_,
		_w2237_,
		_w2238_
	);
	LUT4 #(
		.INIT('h0d00)
	) name1776 (
		_w2211_,
		_w2234_,
		_w2236_,
		_w2237_,
		_w2239_
	);
	LUT3 #(
		.INIT('hd0)
	) name1777 (
		_w2215_,
		_w2231_,
		_w2239_,
		_w2240_
	);
	LUT4 #(
		.INIT('h0133)
	) name1778 (
		_w541_,
		_w1006_,
		_w1033_,
		_w1040_,
		_w2241_
	);
	LUT3 #(
		.INIT('h10)
	) name1779 (
		_w979_,
		_w1061_,
		_w2241_,
		_w2242_
	);
	LUT4 #(
		.INIT('h001f)
	) name1780 (
		_w541_,
		_w1046_,
		_w1051_,
		_w1072_,
		_w2243_
	);
	LUT2 #(
		.INIT('h1)
	) name1781 (
		_w708_,
		_w1080_,
		_w2244_
	);
	LUT2 #(
		.INIT('h8)
	) name1782 (
		_w2243_,
		_w2244_,
		_w2245_
	);
	LUT2 #(
		.INIT('h8)
	) name1783 (
		_w2242_,
		_w2245_,
		_w2246_
	);
	LUT3 #(
		.INIT('h0d)
	) name1784 (
		_w961_,
		_w1080_,
		_w1085_,
		_w2247_
	);
	LUT4 #(
		.INIT('he0fe)
	) name1785 (
		_w541_,
		_w1046_,
		_w1051_,
		_w1084_,
		_w2248_
	);
	LUT3 #(
		.INIT('hd0)
	) name1786 (
		_w2243_,
		_w2247_,
		_w2248_,
		_w2249_
	);
	LUT3 #(
		.INIT('h0b)
	) name1787 (
		_w979_,
		_w1088_,
		_w1094_,
		_w2250_
	);
	LUT4 #(
		.INIT('hb200)
	) name1788 (
		_w969_,
		_w977_,
		_w1088_,
		_w2241_,
		_w2251_
	);
	LUT4 #(
		.INIT('he0fe)
	) name1789 (
		_w541_,
		_w1033_,
		_w1040_,
		_w1093_,
		_w2252_
	);
	LUT4 #(
		.INIT('h0d00)
	) name1790 (
		_w2242_,
		_w2249_,
		_w2251_,
		_w2252_,
		_w2253_
	);
	LUT4 #(
		.INIT('h65aa)
	) name1791 (
		_w1419_,
		_w2240_,
		_w2246_,
		_w2253_,
		_w2254_
	);
	LUT4 #(
		.INIT('h04c4)
	) name1792 (
		_w1019_,
		_w1114_,
		_w2197_,
		_w2254_,
		_w2255_
	);
	LUT4 #(
		.INIT('h9500)
	) name1793 (
		_w1018_,
		_w1128_,
		_w1131_,
		_w2197_,
		_w2256_
	);
	LUT3 #(
		.INIT('h31)
	) name1794 (
		_w1138_,
		_w1141_,
		_w2197_,
		_w2257_
	);
	LUT4 #(
		.INIT('h5054)
	) name1795 (
		_w1019_,
		_w1138_,
		_w1141_,
		_w2197_,
		_w2258_
	);
	LUT4 #(
		.INIT('h0203)
	) name1796 (
		_w652_,
		_w1104_,
		_w1106_,
		_w1111_,
		_w2259_
	);
	LUT4 #(
		.INIT('h001f)
	) name1797 (
		_w528_,
		_w530_,
		_w533_,
		_w1111_,
		_w2260_
	);
	LUT2 #(
		.INIT('h2)
	) name1798 (
		_w2259_,
		_w2260_,
		_w2261_
	);
	LUT4 #(
		.INIT('h5400)
	) name1799 (
		_w541_,
		_w1008_,
		_w1017_,
		_w2261_,
		_w2262_
	);
	LUT2 #(
		.INIT('h1)
	) name1800 (
		_w2258_,
		_w2262_,
		_w2263_
	);
	LUT4 #(
		.INIT('h5700)
	) name1801 (
		_w1136_,
		_w2198_,
		_w2256_,
		_w2263_,
		_w2264_
	);
	LUT4 #(
		.INIT('h0d00)
	) name1802 (
		_w1183_,
		_w2208_,
		_w2255_,
		_w2264_,
		_w2265_
	);
	LUT2 #(
		.INIT('h2)
	) name1803 (
		_w524_,
		_w1019_,
		_w2266_
	);
	LUT4 #(
		.INIT('h0075)
	) name1804 (
		_w526_,
		_w2205_,
		_w2265_,
		_w2266_,
		_w2267_
	);
	LUT2 #(
		.INIT('h2)
	) name1805 (
		\P1_reg3_reg[28]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w2268_
	);
	LUT3 #(
		.INIT('h0b)
	) name1806 (
		_w1019_,
		_w1294_,
		_w2268_,
		_w2269_
	);
	LUT3 #(
		.INIT('h2f)
	) name1807 (
		\P1_state_reg[0]/NET0131 ,
		_w2267_,
		_w2269_,
		_w2270_
	);
	LUT4 #(
		.INIT('h90c0)
	) name1808 (
		\P2_reg3_reg[27]/NET0131 ,
		\P2_reg3_reg[28]/NET0131 ,
		_w1487_,
		_w1971_,
		_w2271_
	);
	LUT3 #(
		.INIT('he0)
	) name1809 (
		_w1491_,
		_w1493_,
		_w1496_,
		_w2272_
	);
	LUT2 #(
		.INIT('h1)
	) name1810 (
		_w2018_,
		_w2272_,
		_w2273_
	);
	LUT4 #(
		.INIT('h006f)
	) name1811 (
		_w2008_,
		_w2027_,
		_w2272_,
		_w2273_,
		_w2274_
	);
	LUT3 #(
		.INIT('h02)
	) name1812 (
		_w1811_,
		_w2035_,
		_w2036_,
		_w2275_
	);
	LUT4 #(
		.INIT('hcff7)
	) name1813 (
		_w1811_,
		_w2033_,
		_w2035_,
		_w2036_,
		_w2276_
	);
	LUT3 #(
		.INIT('h01)
	) name1814 (
		_w1491_,
		_w1493_,
		_w1496_,
		_w2277_
	);
	LUT2 #(
		.INIT('h1)
	) name1815 (
		_w2018_,
		_w2277_,
		_w2278_
	);
	LUT4 #(
		.INIT('hba00)
	) name1816 (
		_w2043_,
		_w2075_,
		_w2078_,
		_w2277_,
		_w2279_
	);
	LUT4 #(
		.INIT('h1f00)
	) name1817 (
		_w1491_,
		_w1493_,
		_w1496_,
		_w2084_,
		_w2280_
	);
	LUT3 #(
		.INIT('h54)
	) name1818 (
		_w2018_,
		_w2086_,
		_w2280_,
		_w2281_
	);
	LUT4 #(
		.INIT('h001f)
	) name1819 (
		_w1491_,
		_w1493_,
		_w1496_,
		_w2082_,
		_w2282_
	);
	LUT2 #(
		.INIT('h2)
	) name1820 (
		_w2083_,
		_w2282_,
		_w2283_
	);
	LUT4 #(
		.INIT('h0e0f)
	) name1821 (
		_w1509_,
		_w2017_,
		_w2281_,
		_w2283_,
		_w2284_
	);
	LUT4 #(
		.INIT('h5700)
	) name1822 (
		_w2081_,
		_w2278_,
		_w2279_,
		_w2284_,
		_w2285_
	);
	LUT3 #(
		.INIT('he0)
	) name1823 (
		_w2274_,
		_w2276_,
		_w2285_,
		_w2286_
	);
	LUT4 #(
		.INIT('h9a00)
	) name1824 (
		_w2027_,
		_w2169_,
		_w2186_,
		_w2272_,
		_w2287_
	);
	LUT3 #(
		.INIT('h54)
	) name1825 (
		_w2192_,
		_w2273_,
		_w2287_,
		_w2288_
	);
	LUT4 #(
		.INIT('h006f)
	) name1826 (
		_w2008_,
		_w2027_,
		_w2277_,
		_w2278_,
		_w2289_
	);
	LUT4 #(
		.INIT('h0800)
	) name1827 (
		_w1811_,
		_w2033_,
		_w2035_,
		_w2036_,
		_w2290_
	);
	LUT2 #(
		.INIT('h4)
	) name1828 (
		_w2289_,
		_w2290_,
		_w2291_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name1829 (
		_w1489_,
		_w2288_,
		_w2291_,
		_w2286_,
		_w2292_
	);
	LUT3 #(
		.INIT('h28)
	) name1830 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		_w1476_,
		_w2293_
	);
	LUT4 #(
		.INIT('h9c00)
	) name1831 (
		\P2_reg3_reg[27]/NET0131 ,
		\P2_reg3_reg[28]/NET0131 ,
		_w1971_,
		_w2293_,
		_w2294_
	);
	LUT2 #(
		.INIT('h4)
	) name1832 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[28]/NET0131 ,
		_w2295_
	);
	LUT2 #(
		.INIT('h1)
	) name1833 (
		_w2294_,
		_w2295_,
		_w2296_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name1834 (
		\P1_state_reg[0]/NET0131 ,
		_w2271_,
		_w2292_,
		_w2296_,
		_w2297_
	);
	LUT4 #(
		.INIT('h70d0)
	) name1835 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg2_reg[27]/NET0131 ,
		_w1476_,
		_w2298_
	);
	LUT2 #(
		.INIT('h8)
	) name1836 (
		\P2_reg2_reg[27]/NET0131 ,
		_w1487_,
		_w2299_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name1837 (
		\P2_reg2_reg[27]/NET0131 ,
		_w1491_,
		_w1493_,
		_w1496_,
		_w2300_
	);
	LUT3 #(
		.INIT('h1e)
	) name1838 (
		_w1509_,
		_w1970_,
		_w1975_,
		_w2301_
	);
	LUT2 #(
		.INIT('h1)
	) name1839 (
		_w1528_,
		_w1594_,
		_w2302_
	);
	LUT3 #(
		.INIT('h32)
	) name1840 (
		_w1556_,
		_w1605_,
		_w1610_,
		_w2303_
	);
	LUT4 #(
		.INIT('h00ef)
	) name1841 (
		_w1565_,
		_w1582_,
		_w1606_,
		_w2303_,
		_w2304_
	);
	LUT3 #(
		.INIT('h54)
	) name1842 (
		_w1528_,
		_w1609_,
		_w1613_,
		_w2305_
	);
	LUT3 #(
		.INIT('h15)
	) name1843 (
		_w1658_,
		_w1663_,
		_w1672_,
		_w2306_
	);
	LUT3 #(
		.INIT('h15)
	) name1844 (
		_w1546_,
		_w1676_,
		_w1684_,
		_w2307_
	);
	LUT2 #(
		.INIT('h8)
	) name1845 (
		_w2306_,
		_w2307_,
		_w2308_
	);
	LUT4 #(
		.INIT('hf200)
	) name1846 (
		_w2302_,
		_w2304_,
		_w2305_,
		_w2308_,
		_w2309_
	);
	LUT3 #(
		.INIT('hd4)
	) name1847 (
		_w1612_,
		_w1676_,
		_w1684_,
		_w2310_
	);
	LUT4 #(
		.INIT('h00fe)
	) name1848 (
		_w1658_,
		_w1663_,
		_w1672_,
		_w1690_,
		_w2311_
	);
	LUT3 #(
		.INIT('hd0)
	) name1849 (
		_w2306_,
		_w2310_,
		_w2311_,
		_w2312_
	);
	LUT3 #(
		.INIT('h15)
	) name1850 (
		_w1642_,
		_w1735_,
		_w1746_,
		_w2313_
	);
	LUT4 #(
		.INIT('h0777)
	) name1851 (
		_w1720_,
		_w1730_,
		_w1751_,
		_w1761_,
		_w2314_
	);
	LUT2 #(
		.INIT('h8)
	) name1852 (
		_w2313_,
		_w2314_,
		_w2315_
	);
	LUT2 #(
		.INIT('h1)
	) name1853 (
		_w1783_,
		_w1840_,
		_w2316_
	);
	LUT4 #(
		.INIT('h0001)
	) name1854 (
		_w1716_,
		_w1783_,
		_w1796_,
		_w1840_,
		_w2317_
	);
	LUT2 #(
		.INIT('h8)
	) name1855 (
		_w2315_,
		_w2317_,
		_w2318_
	);
	LUT3 #(
		.INIT('hb0)
	) name1856 (
		_w2309_,
		_w2312_,
		_w2318_,
		_w2319_
	);
	LUT3 #(
		.INIT('hd4)
	) name1857 (
		_w1689_,
		_w1735_,
		_w1746_,
		_w2320_
	);
	LUT4 #(
		.INIT('h1117)
	) name1858 (
		_w1720_,
		_w1730_,
		_w1751_,
		_w1761_,
		_w2321_
	);
	LUT3 #(
		.INIT('h0d)
	) name1859 (
		_w2314_,
		_w2320_,
		_w2321_,
		_w2322_
	);
	LUT2 #(
		.INIT('h2)
	) name1860 (
		_w2317_,
		_w2322_,
		_w2323_
	);
	LUT3 #(
		.INIT('h0b)
	) name1861 (
		_w1796_,
		_w1845_,
		_w1849_,
		_w2324_
	);
	LUT3 #(
		.INIT('h0b)
	) name1862 (
		_w1840_,
		_w1848_,
		_w1853_,
		_w2325_
	);
	LUT3 #(
		.INIT('hd0)
	) name1863 (
		_w2316_,
		_w2324_,
		_w2325_,
		_w2326_
	);
	LUT2 #(
		.INIT('h4)
	) name1864 (
		_w2323_,
		_w2326_,
		_w2327_
	);
	LUT4 #(
		.INIT('h0133)
	) name1865 (
		_w1509_,
		_w1945_,
		_w1984_,
		_w1988_,
		_w2328_
	);
	LUT4 #(
		.INIT('h0133)
	) name1866 (
		_w1509_,
		_w1909_,
		_w1953_,
		_w1960_,
		_w2329_
	);
	LUT2 #(
		.INIT('h8)
	) name1867 (
		_w2328_,
		_w2329_,
		_w2330_
	);
	LUT2 #(
		.INIT('h1)
	) name1868 (
		_w1821_,
		_w1874_,
		_w2331_
	);
	LUT2 #(
		.INIT('h1)
	) name1869 (
		_w1891_,
		_w1923_,
		_w2332_
	);
	LUT4 #(
		.INIT('h0001)
	) name1870 (
		_w1821_,
		_w1874_,
		_w1891_,
		_w1923_,
		_w2333_
	);
	LUT3 #(
		.INIT('h80)
	) name1871 (
		_w2328_,
		_w2329_,
		_w2333_,
		_w2334_
	);
	LUT3 #(
		.INIT('h0d)
	) name1872 (
		_w1852_,
		_w1874_,
		_w2000_,
		_w2335_
	);
	LUT3 #(
		.INIT('h0b)
	) name1873 (
		_w1923_,
		_w1999_,
		_w2003_,
		_w2336_
	);
	LUT3 #(
		.INIT('hd0)
	) name1874 (
		_w2332_,
		_w2335_,
		_w2336_,
		_w2337_
	);
	LUT4 #(
		.INIT('he0fe)
	) name1875 (
		_w1509_,
		_w1953_,
		_w1960_,
		_w2002_,
		_w2338_
	);
	LUT4 #(
		.INIT('he0fe)
	) name1876 (
		_w1509_,
		_w1984_,
		_w1988_,
		_w1995_,
		_w2339_
	);
	LUT3 #(
		.INIT('hd0)
	) name1877 (
		_w2328_,
		_w2338_,
		_w2339_,
		_w2340_
	);
	LUT3 #(
		.INIT('hd0)
	) name1878 (
		_w2330_,
		_w2337_,
		_w2340_,
		_w2341_
	);
	LUT4 #(
		.INIT('h4f00)
	) name1879 (
		_w2319_,
		_w2327_,
		_w2334_,
		_w2341_,
		_w2342_
	);
	LUT4 #(
		.INIT('h1dd1)
	) name1880 (
		\P2_reg2_reg[27]/NET0131 ,
		_w1497_,
		_w2301_,
		_w2342_,
		_w2343_
	);
	LUT2 #(
		.INIT('h2)
	) name1881 (
		_w2038_,
		_w2343_,
		_w2344_
	);
	LUT4 #(
		.INIT('haa02)
	) name1882 (
		\P2_reg2_reg[27]/NET0131 ,
		_w1491_,
		_w1493_,
		_w1496_,
		_w2345_
	);
	LUT2 #(
		.INIT('h1)
	) name1883 (
		_w2157_,
		_w2158_,
		_w2346_
	);
	LUT3 #(
		.INIT('h0d)
	) name1884 (
		_w2150_,
		_w2156_,
		_w2170_,
		_w2347_
	);
	LUT3 #(
		.INIT('h54)
	) name1885 (
		_w2158_,
		_w2171_,
		_w2174_,
		_w2348_
	);
	LUT3 #(
		.INIT('h0d)
	) name1886 (
		_w2346_,
		_w2347_,
		_w2348_,
		_w2349_
	);
	LUT2 #(
		.INIT('h1)
	) name1887 (
		_w2118_,
		_w2122_,
		_w2350_
	);
	LUT3 #(
		.INIT('h54)
	) name1888 (
		_w2104_,
		_w2118_,
		_w2122_,
		_w2351_
	);
	LUT2 #(
		.INIT('h1)
	) name1889 (
		_w2114_,
		_w2119_,
		_w2352_
	);
	LUT4 #(
		.INIT('h00b2)
	) name1890 (
		_w1569_,
		_w1573_,
		_w2112_,
		_w2115_,
		_w2353_
	);
	LUT3 #(
		.INIT('h01)
	) name1891 (
		_w2104_,
		_w2106_,
		_w2107_,
		_w2354_
	);
	LUT4 #(
		.INIT('h3b00)
	) name1892 (
		_w2111_,
		_w2352_,
		_w2353_,
		_w2354_,
		_w2355_
	);
	LUT3 #(
		.INIT('h0d)
	) name1893 (
		_w1663_,
		_w1672_,
		_w2094_,
		_w2356_
	);
	LUT3 #(
		.INIT('h0d)
	) name1894 (
		_w1676_,
		_w1684_,
		_w2103_,
		_w2357_
	);
	LUT2 #(
		.INIT('h8)
	) name1895 (
		_w2356_,
		_w2357_,
		_w2358_
	);
	LUT3 #(
		.INIT('hd4)
	) name1896 (
		_w1676_,
		_w1684_,
		_w2121_,
		_w2359_
	);
	LUT3 #(
		.INIT('h0b)
	) name1897 (
		_w1663_,
		_w1672_,
		_w2100_,
		_w2360_
	);
	LUT4 #(
		.INIT('h0f04)
	) name1898 (
		_w1663_,
		_w1672_,
		_w2094_,
		_w2100_,
		_w2361_
	);
	LUT3 #(
		.INIT('h07)
	) name1899 (
		_w2356_,
		_w2359_,
		_w2361_,
		_w2362_
	);
	LUT4 #(
		.INIT('h1f00)
	) name1900 (
		_w2351_,
		_w2355_,
		_w2358_,
		_w2362_,
		_w2363_
	);
	LUT2 #(
		.INIT('h1)
	) name1901 (
		_w2131_,
		_w2133_,
		_w2364_
	);
	LUT4 #(
		.INIT('h0001)
	) name1902 (
		_w2127_,
		_w2131_,
		_w2132_,
		_w2133_,
		_w2365_
	);
	LUT4 #(
		.INIT('hdd0d)
	) name1903 (
		_w1720_,
		_w1730_,
		_w1751_,
		_w1761_,
		_w2366_
	);
	LUT3 #(
		.INIT('h0d)
	) name1904 (
		_w1735_,
		_w1746_,
		_w2095_,
		_w2367_
	);
	LUT2 #(
		.INIT('h8)
	) name1905 (
		_w2366_,
		_w2367_,
		_w2368_
	);
	LUT2 #(
		.INIT('h8)
	) name1906 (
		_w2365_,
		_w2368_,
		_w2369_
	);
	LUT3 #(
		.INIT('h2b)
	) name1907 (
		_w1735_,
		_w1746_,
		_w2099_,
		_w2370_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name1908 (
		_w1720_,
		_w1730_,
		_w1751_,
		_w1761_,
		_w2371_
	);
	LUT4 #(
		.INIT('h4d44)
	) name1909 (
		_w1720_,
		_w1730_,
		_w1751_,
		_w1761_,
		_w2372_
	);
	LUT3 #(
		.INIT('h0d)
	) name1910 (
		_w2366_,
		_w2370_,
		_w2372_,
		_w2373_
	);
	LUT2 #(
		.INIT('h2)
	) name1911 (
		_w2365_,
		_w2373_,
		_w2374_
	);
	LUT3 #(
		.INIT('h0b)
	) name1912 (
		_w2132_,
		_w2141_,
		_w2145_,
		_w2375_
	);
	LUT3 #(
		.INIT('h54)
	) name1913 (
		_w2133_,
		_w2146_,
		_w2151_,
		_w2376_
	);
	LUT3 #(
		.INIT('h0d)
	) name1914 (
		_w2364_,
		_w2375_,
		_w2376_,
		_w2377_
	);
	LUT4 #(
		.INIT('h0b00)
	) name1915 (
		_w2363_,
		_w2369_,
		_w2374_,
		_w2377_,
		_w2378_
	);
	LUT2 #(
		.INIT('h1)
	) name1916 (
		_w2134_,
		_w2156_,
		_w2379_
	);
	LUT4 #(
		.INIT('h0001)
	) name1917 (
		_w2134_,
		_w2156_,
		_w2157_,
		_w2158_,
		_w2380_
	);
	LUT4 #(
		.INIT('h00ef)
	) name1918 (
		_w1509_,
		_w1984_,
		_w1988_,
		_w2163_,
		_w2381_
	);
	LUT4 #(
		.INIT('h10f1)
	) name1919 (
		_w1509_,
		_w1953_,
		_w1960_,
		_w2175_,
		_w2382_
	);
	LUT4 #(
		.INIT('h00f1)
	) name1920 (
		_w1509_,
		_w1984_,
		_w1988_,
		_w2182_,
		_w2383_
	);
	LUT4 #(
		.INIT('hef0e)
	) name1921 (
		_w1509_,
		_w1984_,
		_w1988_,
		_w2182_,
		_w2384_
	);
	LUT4 #(
		.INIT('h00ef)
	) name1922 (
		_w1509_,
		_w1953_,
		_w1960_,
		_w2159_,
		_w2385_
	);
	LUT4 #(
		.INIT('h0800)
	) name1923 (
		_w2381_,
		_w2382_,
		_w2384_,
		_w2385_,
		_w2386_
	);
	LUT4 #(
		.INIT('h7500)
	) name1924 (
		_w2349_,
		_w2378_,
		_w2380_,
		_w2386_,
		_w2387_
	);
	LUT4 #(
		.INIT('h0df2)
	) name1925 (
		_w2381_,
		_w2382_,
		_w2384_,
		_w2301_,
		_w2388_
	);
	LUT4 #(
		.INIT('h80a2)
	) name1926 (
		_w2039_,
		_w2387_,
		_w2301_,
		_w2388_,
		_w2389_
	);
	LUT3 #(
		.INIT('ha8)
	) name1927 (
		_w2188_,
		_w2345_,
		_w2389_,
		_w2390_
	);
	LUT4 #(
		.INIT('h80a2)
	) name1928 (
		_w1497_,
		_w2387_,
		_w2301_,
		_w2388_,
		_w2391_
	);
	LUT4 #(
		.INIT('h2111)
	) name1929 (
		_w2023_,
		_w2042_,
		_w2073_,
		_w2074_,
		_w2392_
	);
	LUT2 #(
		.INIT('h4)
	) name1930 (
		_w1988_,
		_w2042_,
		_w2393_
	);
	LUT4 #(
		.INIT('h111d)
	) name1931 (
		\P2_reg2_reg[27]/NET0131 ,
		_w2039_,
		_w2392_,
		_w2393_,
		_w2394_
	);
	LUT2 #(
		.INIT('h4)
	) name1932 (
		_w1972_,
		_w2088_,
		_w2395_
	);
	LUT4 #(
		.INIT('h0057)
	) name1933 (
		\P2_reg2_reg[27]/NET0131 ,
		_w2086_,
		_w2087_,
		_w2395_,
		_w2396_
	);
	LUT4 #(
		.INIT('hef00)
	) name1934 (
		_w1509_,
		_w1970_,
		_w2085_,
		_w2396_,
		_w2397_
	);
	LUT3 #(
		.INIT('hd0)
	) name1935 (
		_w2081_,
		_w2394_,
		_w2397_,
		_w2398_
	);
	LUT4 #(
		.INIT('h5700)
	) name1936 (
		_w2193_,
		_w2300_,
		_w2391_,
		_w2398_,
		_w2399_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name1937 (
		_w1489_,
		_w2344_,
		_w2390_,
		_w2399_,
		_w2400_
	);
	LUT4 #(
		.INIT('heeec)
	) name1938 (
		\P1_state_reg[0]/NET0131 ,
		_w2298_,
		_w2299_,
		_w2400_,
		_w2401_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name1939 (
		\P1_reg2_reg[28]/NET0131 ,
		_w528_,
		_w530_,
		_w533_,
		_w2402_
	);
	LUT4 #(
		.INIT('h8288)
	) name1940 (
		_w534_,
		_w1419_,
		_w2201_,
		_w2203_,
		_w2403_
	);
	LUT3 #(
		.INIT('ha8)
	) name1941 (
		_w1286_,
		_w2402_,
		_w2403_,
		_w2404_
	);
	LUT4 #(
		.INIT('hddd1)
	) name1942 (
		\P1_reg2_reg[28]/NET0131 ,
		_w534_,
		_w2206_,
		_w2207_,
		_w2405_
	);
	LUT4 #(
		.INIT('h5400)
	) name1943 (
		_w541_,
		_w1008_,
		_w1017_,
		_w1138_,
		_w2406_
	);
	LUT4 #(
		.INIT('h9500)
	) name1944 (
		_w1018_,
		_w1128_,
		_w1131_,
		_w1136_,
		_w2407_
	);
	LUT2 #(
		.INIT('h1)
	) name1945 (
		_w2406_,
		_w2407_,
		_w2408_
	);
	LUT4 #(
		.INIT('h08aa)
	) name1946 (
		_w534_,
		_w1114_,
		_w2254_,
		_w2408_,
		_w2409_
	);
	LUT2 #(
		.INIT('h4)
	) name1947 (
		_w1019_,
		_w1143_,
		_w2410_
	);
	LUT4 #(
		.INIT('h00ab)
	) name1948 (
		_w534_,
		_w1136_,
		_w1138_,
		_w1141_,
		_w2411_
	);
	LUT2 #(
		.INIT('h4)
	) name1949 (
		_w534_,
		_w1114_,
		_w2412_
	);
	LUT4 #(
		.INIT('h1131)
	) name1950 (
		\P1_reg2_reg[28]/NET0131 ,
		_w2410_,
		_w2411_,
		_w2412_,
		_w2413_
	);
	LUT4 #(
		.INIT('h0d00)
	) name1951 (
		_w1183_,
		_w2405_,
		_w2409_,
		_w2413_,
		_w2414_
	);
	LUT2 #(
		.INIT('h8)
	) name1952 (
		\P1_reg2_reg[28]/NET0131 ,
		_w524_,
		_w2415_
	);
	LUT4 #(
		.INIT('h0075)
	) name1953 (
		_w526_,
		_w2404_,
		_w2414_,
		_w2415_,
		_w2416_
	);
	LUT2 #(
		.INIT('h2)
	) name1954 (
		\P1_reg2_reg[28]/NET0131 ,
		_w511_,
		_w2417_
	);
	LUT3 #(
		.INIT('hf2)
	) name1955 (
		\P1_state_reg[0]/NET0131 ,
		_w2416_,
		_w2417_,
		_w2418_
	);
	LUT2 #(
		.INIT('h2)
	) name1956 (
		\P1_reg1_reg[29]/NET0131 ,
		_w511_,
		_w2419_
	);
	LUT2 #(
		.INIT('h8)
	) name1957 (
		\P1_reg1_reg[29]/NET0131 ,
		_w524_,
		_w2420_
	);
	LUT3 #(
		.INIT('h0e)
	) name1958 (
		_w528_,
		_w530_,
		_w533_,
		_w2421_
	);
	LUT4 #(
		.INIT('haa02)
	) name1959 (
		\P1_reg1_reg[29]/NET0131 ,
		_w528_,
		_w530_,
		_w533_,
		_w2422_
	);
	LUT4 #(
		.INIT('hc355)
	) name1960 (
		\P1_reg1_reg[29]/NET0131 ,
		_w647_,
		_w1102_,
		_w2421_,
		_w2423_
	);
	LUT4 #(
		.INIT('hc0a0)
	) name1961 (
		\P1_reg1_reg[29]/NET0131 ,
		_w1134_,
		_w1136_,
		_w2421_,
		_w2424_
	);
	LUT4 #(
		.INIT('h7d3f)
	) name1962 (
		_w652_,
		_w1104_,
		_w1106_,
		_w1111_,
		_w2425_
	);
	LUT3 #(
		.INIT('hd0)
	) name1963 (
		_w1138_,
		_w2421_,
		_w2425_,
		_w2426_
	);
	LUT4 #(
		.INIT('h08aa)
	) name1964 (
		\P1_reg1_reg[29]/NET0131 ,
		_w1138_,
		_w2421_,
		_w2425_,
		_w2427_
	);
	LUT3 #(
		.INIT('h07)
	) name1965 (
		_w1139_,
		_w2421_,
		_w2427_,
		_w2428_
	);
	LUT2 #(
		.INIT('h4)
	) name1966 (
		_w2424_,
		_w2428_,
		_w2429_
	);
	LUT3 #(
		.INIT('hd0)
	) name1967 (
		_w1114_,
		_w2423_,
		_w2429_,
		_w2430_
	);
	LUT4 #(
		.INIT('h6500)
	) name1968 (
		_w647_,
		_w1265_,
		_w1284_,
		_w2421_,
		_w2431_
	);
	LUT4 #(
		.INIT('h30a0)
	) name1969 (
		\P1_reg1_reg[29]/NET0131 ,
		_w1182_,
		_w1183_,
		_w2421_,
		_w2432_
	);
	LUT4 #(
		.INIT('h0057)
	) name1970 (
		_w1286_,
		_w2422_,
		_w2431_,
		_w2432_,
		_w2433_
	);
	LUT4 #(
		.INIT('h3111)
	) name1971 (
		_w526_,
		_w2420_,
		_w2430_,
		_w2433_,
		_w2434_
	);
	LUT3 #(
		.INIT('hce)
	) name1972 (
		\P1_state_reg[0]/NET0131 ,
		_w2419_,
		_w2434_,
		_w2435_
	);
	LUT3 #(
		.INIT('ha8)
	) name1973 (
		_w1487_,
		_w1938_,
		_w1954_,
		_w2436_
	);
	LUT3 #(
		.INIT('h1e)
	) name1974 (
		_w1509_,
		_w1953_,
		_w1960_,
		_w2437_
	);
	LUT4 #(
		.INIT('h40f0)
	) name1975 (
		_w1692_,
		_w1763_,
		_w1842_,
		_w1847_,
		_w2438_
	);
	LUT4 #(
		.INIT('h0070)
	) name1976 (
		_w1687_,
		_w1843_,
		_w1855_,
		_w2438_,
		_w2439_
	);
	LUT4 #(
		.INIT('h3cb4)
	) name1977 (
		_w1925_,
		_w2005_,
		_w2437_,
		_w2439_,
		_w2440_
	);
	LUT4 #(
		.INIT('h010d)
	) name1978 (
		_w1955_,
		_w2272_,
		_w2276_,
		_w2440_,
		_w2441_
	);
	LUT2 #(
		.INIT('h4)
	) name1979 (
		_w1907_,
		_w2042_,
		_w2442_
	);
	LUT4 #(
		.INIT('h00de)
	) name1980 (
		_w1943_,
		_w2042_,
		_w2073_,
		_w2442_,
		_w2443_
	);
	LUT4 #(
		.INIT('h04c4)
	) name1981 (
		_w1955_,
		_w2081_,
		_w2277_,
		_w2443_,
		_w2444_
	);
	LUT3 #(
		.INIT('h54)
	) name1982 (
		_w1955_,
		_w2086_,
		_w2280_,
		_w2445_
	);
	LUT4 #(
		.INIT('h00ef)
	) name1983 (
		_w1509_,
		_w1953_,
		_w2283_,
		_w2445_,
		_w2446_
	);
	LUT2 #(
		.INIT('h4)
	) name1984 (
		_w2444_,
		_w2446_,
		_w2447_
	);
	LUT3 #(
		.INIT('hb0)
	) name1985 (
		_w2102_,
		_w2130_,
		_w2144_,
		_w2448_
	);
	LUT4 #(
		.INIT('h40f0)
	) name1986 (
		_w2102_,
		_w2130_,
		_w2136_,
		_w2144_,
		_w2449_
	);
	LUT3 #(
		.INIT('hc4)
	) name1987 (
		_w2154_,
		_w2161_,
		_w2449_,
		_w2450_
	);
	LUT2 #(
		.INIT('h8)
	) name1988 (
		_w2136_,
		_w2161_,
		_w2451_
	);
	LUT4 #(
		.INIT('h4000)
	) name1989 (
		_w2124_,
		_w2126_,
		_w2130_,
		_w2451_,
		_w2452_
	);
	LUT4 #(
		.INIT('h3339)
	) name1990 (
		_w2177_,
		_w2437_,
		_w2452_,
		_w2450_,
		_w2453_
	);
	LUT4 #(
		.INIT('h0131)
	) name1991 (
		_w1955_,
		_w2192_,
		_w2272_,
		_w2453_,
		_w2454_
	);
	LUT4 #(
		.INIT('h10d0)
	) name1992 (
		_w1955_,
		_w2277_,
		_w2290_,
		_w2440_,
		_w2455_
	);
	LUT4 #(
		.INIT('h0100)
	) name1993 (
		_w2441_,
		_w2454_,
		_w2455_,
		_w2447_,
		_w2456_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name1994 (
		\P1_state_reg[0]/NET0131 ,
		_w1489_,
		_w2436_,
		_w2456_,
		_w2457_
	);
	LUT2 #(
		.INIT('h4)
	) name1995 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[24]/NET0131 ,
		_w2458_
	);
	LUT4 #(
		.INIT('h001f)
	) name1996 (
		_w1938_,
		_w1954_,
		_w2293_,
		_w2458_,
		_w2459_
	);
	LUT2 #(
		.INIT('hb)
	) name1997 (
		_w2457_,
		_w2459_,
		_w2460_
	);
	LUT2 #(
		.INIT('h2)
	) name1998 (
		_w1487_,
		_w1985_,
		_w2461_
	);
	LUT4 #(
		.INIT('h001f)
	) name1999 (
		_w1491_,
		_w1493_,
		_w1496_,
		_w1985_,
		_w2462_
	);
	LUT3 #(
		.INIT('h1e)
	) name2000 (
		_w1509_,
		_w1984_,
		_w1988_,
		_w2463_
	);
	LUT3 #(
		.INIT('h02)
	) name2001 (
		_w1731_,
		_w1783_,
		_w1796_,
		_w2464_
	);
	LUT2 #(
		.INIT('h8)
	) name2002 (
		_w1547_,
		_w1685_,
		_w2465_
	);
	LUT3 #(
		.INIT('hb0)
	) name2003 (
		_w1614_,
		_w1685_,
		_w1688_,
		_w2466_
	);
	LUT4 #(
		.INIT('h1f00)
	) name2004 (
		_w1608_,
		_w1611_,
		_w2465_,
		_w2466_,
		_w2467_
	);
	LUT2 #(
		.INIT('h8)
	) name2005 (
		_w1659_,
		_w1762_,
		_w2468_
	);
	LUT3 #(
		.INIT('h70)
	) name2006 (
		_w1691_,
		_w1762_,
		_w1844_,
		_w2469_
	);
	LUT3 #(
		.INIT('h01)
	) name2007 (
		_w1783_,
		_w1796_,
		_w1846_,
		_w2470_
	);
	LUT4 #(
		.INIT('h00a2)
	) name2008 (
		_w1850_,
		_w2464_,
		_w2469_,
		_w2470_,
		_w2471_
	);
	LUT4 #(
		.INIT('hdf00)
	) name2009 (
		_w2464_,
		_w2467_,
		_w2468_,
		_w2471_,
		_w2472_
	);
	LUT3 #(
		.INIT('h02)
	) name2010 (
		_w1841_,
		_w1874_,
		_w1891_,
		_w2473_
	);
	LUT3 #(
		.INIT('h80)
	) name2011 (
		_w1924_,
		_w1962_,
		_w2473_,
		_w2474_
	);
	LUT3 #(
		.INIT('h01)
	) name2012 (
		_w1854_,
		_w1874_,
		_w1891_,
		_w2475_
	);
	LUT2 #(
		.INIT('h2)
	) name2013 (
		_w2001_,
		_w2475_,
		_w2476_
	);
	LUT4 #(
		.INIT('h8808)
	) name2014 (
		_w1924_,
		_w1962_,
		_w2001_,
		_w2475_,
		_w2477_
	);
	LUT4 #(
		.INIT('h000d)
	) name2015 (
		_w1962_,
		_w2004_,
		_w1995_,
		_w1996_,
		_w2478_
	);
	LUT2 #(
		.INIT('h4)
	) name2016 (
		_w2477_,
		_w2478_,
		_w2479_
	);
	LUT4 #(
		.INIT('h65aa)
	) name2017 (
		_w2463_,
		_w2472_,
		_w2474_,
		_w2479_,
		_w2480_
	);
	LUT4 #(
		.INIT('h010d)
	) name2018 (
		_w1985_,
		_w2272_,
		_w2276_,
		_w2480_,
		_w2481_
	);
	LUT4 #(
		.INIT('h00fe)
	) name2019 (
		_w1491_,
		_w1493_,
		_w1496_,
		_w1985_,
		_w2482_
	);
	LUT4 #(
		.INIT('hef00)
	) name2020 (
		_w1941_,
		_w1940_,
		_w1942_,
		_w2042_,
		_w2483_
	);
	LUT4 #(
		.INIT('hc8cc)
	) name2021 (
		_w1943_,
		_w1975_,
		_w1988_,
		_w2073_,
		_w2484_
	);
	LUT3 #(
		.INIT('h15)
	) name2022 (
		_w2042_,
		_w2073_,
		_w2074_,
		_w2485_
	);
	LUT4 #(
		.INIT('h8a88)
	) name2023 (
		_w2277_,
		_w2483_,
		_w2484_,
		_w2485_,
		_w2486_
	);
	LUT3 #(
		.INIT('h54)
	) name2024 (
		_w1985_,
		_w2086_,
		_w2280_,
		_w2487_
	);
	LUT4 #(
		.INIT('h00ef)
	) name2025 (
		_w1509_,
		_w1984_,
		_w2283_,
		_w2487_,
		_w2488_
	);
	LUT4 #(
		.INIT('h5700)
	) name2026 (
		_w2081_,
		_w2482_,
		_w2486_,
		_w2488_,
		_w2489_
	);
	LUT2 #(
		.INIT('h4)
	) name2027 (
		_w2481_,
		_w2489_,
		_w2490_
	);
	LUT3 #(
		.INIT('h02)
	) name2028 (
		_w2128_,
		_w2131_,
		_w2132_,
		_w2491_
	);
	LUT4 #(
		.INIT('h8a00)
	) name2029 (
		_w2105_,
		_w2117_,
		_w2120_,
		_w2125_,
		_w2492_
	);
	LUT3 #(
		.INIT('h15)
	) name2030 (
		_w2098_,
		_w2123_,
		_w2125_,
		_w2493_
	);
	LUT2 #(
		.INIT('h8)
	) name2031 (
		_w2096_,
		_w2129_,
		_w2494_
	);
	LUT4 #(
		.INIT('h8a00)
	) name2032 (
		_w2491_,
		_w2492_,
		_w2493_,
		_w2494_,
		_w2495_
	);
	LUT3 #(
		.INIT('h07)
	) name2033 (
		_w2101_,
		_w2129_,
		_w2140_,
		_w2496_
	);
	LUT3 #(
		.INIT('h10)
	) name2034 (
		_w2131_,
		_w2132_,
		_w2143_,
		_w2497_
	);
	LUT4 #(
		.INIT('h0051)
	) name2035 (
		_w2148_,
		_w2491_,
		_w2496_,
		_w2497_,
		_w2498_
	);
	LUT3 #(
		.INIT('h02)
	) name2036 (
		_w2135_,
		_w2156_,
		_w2157_,
		_w2499_
	);
	LUT3 #(
		.INIT('h80)
	) name2037 (
		_w2160_,
		_w2164_,
		_w2499_,
		_w2500_
	);
	LUT3 #(
		.INIT('h02)
	) name2038 (
		_w2153_,
		_w2156_,
		_w2157_,
		_w2501_
	);
	LUT2 #(
		.INIT('h1)
	) name2039 (
		_w2173_,
		_w2501_,
		_w2502_
	);
	LUT4 #(
		.INIT('h8880)
	) name2040 (
		_w2160_,
		_w2164_,
		_w2173_,
		_w2501_,
		_w2503_
	);
	LUT4 #(
		.INIT('hefcc)
	) name2041 (
		_w2162_,
		_w2163_,
		_w2176_,
		_w2183_,
		_w2504_
	);
	LUT2 #(
		.INIT('h4)
	) name2042 (
		_w2503_,
		_w2504_,
		_w2505_
	);
	LUT4 #(
		.INIT('h4f00)
	) name2043 (
		_w2495_,
		_w2498_,
		_w2500_,
		_w2505_,
		_w2506_
	);
	LUT4 #(
		.INIT('h3113)
	) name2044 (
		_w2272_,
		_w2462_,
		_w2463_,
		_w2506_,
		_w2507_
	);
	LUT4 #(
		.INIT('h10d0)
	) name2045 (
		_w1985_,
		_w2277_,
		_w2290_,
		_w2480_,
		_w2508_
	);
	LUT3 #(
		.INIT('h0e)
	) name2046 (
		_w2192_,
		_w2507_,
		_w2508_,
		_w2509_
	);
	LUT4 #(
		.INIT('h3111)
	) name2047 (
		_w1489_,
		_w2461_,
		_w2490_,
		_w2509_,
		_w2510_
	);
	LUT2 #(
		.INIT('h4)
	) name2048 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[26]/NET0131 ,
		_w2511_
	);
	LUT4 #(
		.INIT('h9c00)
	) name2049 (
		\P2_reg3_reg[25]/NET0131 ,
		\P2_reg3_reg[26]/NET0131 ,
		_w1938_,
		_w2293_,
		_w2512_
	);
	LUT2 #(
		.INIT('h1)
	) name2050 (
		_w2511_,
		_w2512_,
		_w2513_
	);
	LUT3 #(
		.INIT('h2f)
	) name2051 (
		\P1_state_reg[0]/NET0131 ,
		_w2510_,
		_w2513_,
		_w2514_
	);
	LUT4 #(
		.INIT('h70d0)
	) name2052 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg2_reg[24]/NET0131 ,
		_w1476_,
		_w2515_
	);
	LUT2 #(
		.INIT('h8)
	) name2053 (
		\P2_reg2_reg[24]/NET0131 ,
		_w1487_,
		_w2516_
	);
	LUT4 #(
		.INIT('h20e0)
	) name2054 (
		\P2_reg2_reg[24]/NET0131 ,
		_w1497_,
		_w2038_,
		_w2440_,
		_w2517_
	);
	LUT4 #(
		.INIT('h20e0)
	) name2055 (
		\P2_reg2_reg[24]/NET0131 ,
		_w2039_,
		_w2081_,
		_w2443_,
		_w2518_
	);
	LUT3 #(
		.INIT('he0)
	) name2056 (
		_w1938_,
		_w1954_,
		_w2088_,
		_w2519_
	);
	LUT4 #(
		.INIT('h0057)
	) name2057 (
		\P2_reg2_reg[24]/NET0131 ,
		_w2086_,
		_w2087_,
		_w2519_,
		_w2520_
	);
	LUT4 #(
		.INIT('hef00)
	) name2058 (
		_w1509_,
		_w1953_,
		_w2085_,
		_w2520_,
		_w2521_
	);
	LUT2 #(
		.INIT('h4)
	) name2059 (
		_w2518_,
		_w2521_,
		_w2522_
	);
	LUT4 #(
		.INIT('h20e0)
	) name2060 (
		\P2_reg2_reg[24]/NET0131 ,
		_w2039_,
		_w2188_,
		_w2453_,
		_w2523_
	);
	LUT4 #(
		.INIT('h20e0)
	) name2061 (
		\P2_reg2_reg[24]/NET0131 ,
		_w1497_,
		_w2193_,
		_w2453_,
		_w2524_
	);
	LUT4 #(
		.INIT('h0100)
	) name2062 (
		_w2517_,
		_w2523_,
		_w2524_,
		_w2522_,
		_w2525_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name2063 (
		\P1_state_reg[0]/NET0131 ,
		_w1489_,
		_w2516_,
		_w2525_,
		_w2526_
	);
	LUT2 #(
		.INIT('he)
	) name2064 (
		_w2515_,
		_w2526_,
		_w2527_
	);
	LUT4 #(
		.INIT('h70d0)
	) name2065 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg2_reg[25]/NET0131 ,
		_w1476_,
		_w2528_
	);
	LUT2 #(
		.INIT('h8)
	) name2066 (
		\P2_reg2_reg[25]/NET0131 ,
		_w1487_,
		_w2529_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name2067 (
		\P2_reg2_reg[25]/NET0131 ,
		_w1491_,
		_w1493_,
		_w1496_,
		_w2530_
	);
	LUT4 #(
		.INIT('h54ab)
	) name2068 (
		_w1509_,
		_w1926_,
		_w1935_,
		_w1943_,
		_w2531_
	);
	LUT3 #(
		.INIT('hc4)
	) name2069 (
		_w2329_,
		_w2338_,
		_w2336_,
		_w2532_
	);
	LUT2 #(
		.INIT('h8)
	) name2070 (
		_w2302_,
		_w2307_,
		_w2533_
	);
	LUT3 #(
		.INIT('h70)
	) name2071 (
		_w2305_,
		_w2307_,
		_w2310_,
		_w2534_
	);
	LUT2 #(
		.INIT('h8)
	) name2072 (
		_w2306_,
		_w2313_,
		_w2535_
	);
	LUT4 #(
		.INIT('h4f00)
	) name2073 (
		_w2304_,
		_w2533_,
		_w2534_,
		_w2535_,
		_w2536_
	);
	LUT4 #(
		.INIT('h0001)
	) name2074 (
		_w1783_,
		_w1821_,
		_w1840_,
		_w1874_,
		_w2537_
	);
	LUT3 #(
		.INIT('h10)
	) name2075 (
		_w1716_,
		_w1796_,
		_w2314_,
		_w2538_
	);
	LUT2 #(
		.INIT('h8)
	) name2076 (
		_w2537_,
		_w2538_,
		_w2539_
	);
	LUT2 #(
		.INIT('h8)
	) name2077 (
		_w2536_,
		_w2539_,
		_w2540_
	);
	LUT3 #(
		.INIT('hb0)
	) name2078 (
		_w2311_,
		_w2313_,
		_w2320_,
		_w2541_
	);
	LUT3 #(
		.INIT('h10)
	) name2079 (
		_w1716_,
		_w1796_,
		_w2321_,
		_w2542_
	);
	LUT2 #(
		.INIT('h2)
	) name2080 (
		_w2324_,
		_w2542_,
		_w2543_
	);
	LUT4 #(
		.INIT('h00a2)
	) name2081 (
		_w2324_,
		_w2538_,
		_w2541_,
		_w2542_,
		_w2544_
	);
	LUT3 #(
		.INIT('hb0)
	) name2082 (
		_w2325_,
		_w2331_,
		_w2335_,
		_w2545_
	);
	LUT3 #(
		.INIT('hd0)
	) name2083 (
		_w2537_,
		_w2544_,
		_w2545_,
		_w2546_
	);
	LUT2 #(
		.INIT('h8)
	) name2084 (
		_w2329_,
		_w2332_,
		_w2547_
	);
	LUT4 #(
		.INIT('h20aa)
	) name2085 (
		_w2532_,
		_w2540_,
		_w2546_,
		_w2547_,
		_w2548_
	);
	LUT4 #(
		.INIT('h1dd1)
	) name2086 (
		\P2_reg2_reg[25]/NET0131 ,
		_w1497_,
		_w2531_,
		_w2548_,
		_w2549_
	);
	LUT2 #(
		.INIT('h2)
	) name2087 (
		_w2038_,
		_w2549_,
		_w2550_
	);
	LUT2 #(
		.INIT('h8)
	) name2088 (
		_w2346_,
		_w2385_,
		_w2551_
	);
	LUT4 #(
		.INIT('h0001)
	) name2089 (
		_w2131_,
		_w2133_,
		_w2134_,
		_w2156_,
		_w2552_
	);
	LUT3 #(
		.INIT('h10)
	) name2090 (
		_w2127_,
		_w2132_,
		_w2366_,
		_w2553_
	);
	LUT3 #(
		.INIT('h70)
	) name2091 (
		_w2367_,
		_w2361_,
		_w2370_,
		_w2554_
	);
	LUT3 #(
		.INIT('h10)
	) name2092 (
		_w2127_,
		_w2132_,
		_w2372_,
		_w2555_
	);
	LUT2 #(
		.INIT('h2)
	) name2093 (
		_w2375_,
		_w2555_,
		_w2556_
	);
	LUT4 #(
		.INIT('h00a2)
	) name2094 (
		_w2375_,
		_w2553_,
		_w2554_,
		_w2555_,
		_w2557_
	);
	LUT3 #(
		.INIT('h2a)
	) name2095 (
		_w2347_,
		_w2376_,
		_w2379_,
		_w2558_
	);
	LUT4 #(
		.INIT('h08aa)
	) name2096 (
		_w2551_,
		_w2552_,
		_w2557_,
		_w2558_,
		_w2559_
	);
	LUT2 #(
		.INIT('h8)
	) name2097 (
		_w2552_,
		_w2553_,
		_w2560_
	);
	LUT3 #(
		.INIT('h15)
	) name2098 (
		_w2359_,
		_w2351_,
		_w2357_,
		_w2561_
	);
	LUT2 #(
		.INIT('h8)
	) name2099 (
		_w2367_,
		_w2356_,
		_w2562_
	);
	LUT4 #(
		.INIT('h8f00)
	) name2100 (
		_w2355_,
		_w2357_,
		_w2561_,
		_w2562_,
		_w2563_
	);
	LUT3 #(
		.INIT('h4c)
	) name2101 (
		_w2348_,
		_w2382_,
		_w2385_,
		_w2564_
	);
	LUT4 #(
		.INIT('h7f00)
	) name2102 (
		_w2563_,
		_w2551_,
		_w2560_,
		_w2564_,
		_w2565_
	);
	LUT4 #(
		.INIT('h8288)
	) name2103 (
		_w1497_,
		_w2531_,
		_w2559_,
		_w2565_,
		_w2566_
	);
	LUT4 #(
		.INIT('h5400)
	) name2104 (
		_w1509_,
		_w1926_,
		_w1935_,
		_w2084_,
		_w2567_
	);
	LUT2 #(
		.INIT('h4)
	) name2105 (
		_w1939_,
		_w2088_,
		_w2568_
	);
	LUT4 #(
		.INIT('h0057)
	) name2106 (
		\P2_reg2_reg[25]/NET0131 ,
		_w2086_,
		_w2087_,
		_w2568_,
		_w2569_
	);
	LUT3 #(
		.INIT('h70)
	) name2107 (
		_w1497_,
		_w2567_,
		_w2569_,
		_w2570_
	);
	LUT4 #(
		.INIT('h5700)
	) name2108 (
		_w2193_,
		_w2530_,
		_w2566_,
		_w2570_,
		_w2571_
	);
	LUT4 #(
		.INIT('haa02)
	) name2109 (
		\P2_reg2_reg[25]/NET0131 ,
		_w1491_,
		_w1493_,
		_w1496_,
		_w2572_
	);
	LUT3 #(
		.INIT('hb0)
	) name2110 (
		_w1956_,
		_w1959_,
		_w2042_,
		_w2573_
	);
	LUT4 #(
		.INIT('h0603)
	) name2111 (
		_w1943_,
		_w1988_,
		_w2042_,
		_w2073_,
		_w2574_
	);
	LUT4 #(
		.INIT('h111d)
	) name2112 (
		\P2_reg2_reg[25]/NET0131 ,
		_w2039_,
		_w2573_,
		_w2574_,
		_w2575_
	);
	LUT2 #(
		.INIT('h2)
	) name2113 (
		_w2081_,
		_w2575_,
		_w2576_
	);
	LUT4 #(
		.INIT('h8288)
	) name2114 (
		_w2039_,
		_w2531_,
		_w2559_,
		_w2565_,
		_w2577_
	);
	LUT3 #(
		.INIT('ha8)
	) name2115 (
		_w2188_,
		_w2572_,
		_w2577_,
		_w2578_
	);
	LUT3 #(
		.INIT('h10)
	) name2116 (
		_w2576_,
		_w2578_,
		_w2571_,
		_w2579_
	);
	LUT4 #(
		.INIT('h1311)
	) name2117 (
		_w1489_,
		_w2529_,
		_w2550_,
		_w2579_,
		_w2580_
	);
	LUT3 #(
		.INIT('hce)
	) name2118 (
		\P1_state_reg[0]/NET0131 ,
		_w2528_,
		_w2580_,
		_w2581_
	);
	LUT4 #(
		.INIT('h70d0)
	) name2119 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg2_reg[26]/NET0131 ,
		_w1476_,
		_w2582_
	);
	LUT2 #(
		.INIT('h8)
	) name2120 (
		\P2_reg2_reg[26]/NET0131 ,
		_w1487_,
		_w2583_
	);
	LUT4 #(
		.INIT('h20e0)
	) name2121 (
		\P2_reg2_reg[26]/NET0131 ,
		_w1497_,
		_w2038_,
		_w2480_,
		_w2584_
	);
	LUT4 #(
		.INIT('haa02)
	) name2122 (
		\P2_reg2_reg[26]/NET0131 ,
		_w1491_,
		_w1493_,
		_w1496_,
		_w2585_
	);
	LUT4 #(
		.INIT('h8a88)
	) name2123 (
		_w2039_,
		_w2483_,
		_w2484_,
		_w2485_,
		_w2586_
	);
	LUT2 #(
		.INIT('h4)
	) name2124 (
		_w1985_,
		_w2088_,
		_w2587_
	);
	LUT4 #(
		.INIT('h0057)
	) name2125 (
		\P2_reg2_reg[26]/NET0131 ,
		_w2086_,
		_w2087_,
		_w2587_,
		_w2588_
	);
	LUT4 #(
		.INIT('hef00)
	) name2126 (
		_w1509_,
		_w1984_,
		_w2085_,
		_w2588_,
		_w2589_
	);
	LUT4 #(
		.INIT('h5700)
	) name2127 (
		_w2081_,
		_w2585_,
		_w2586_,
		_w2589_,
		_w2590_
	);
	LUT2 #(
		.INIT('h4)
	) name2128 (
		_w2584_,
		_w2590_,
		_w2591_
	);
	LUT4 #(
		.INIT('hd11d)
	) name2129 (
		\P2_reg2_reg[26]/NET0131 ,
		_w1497_,
		_w2463_,
		_w2506_,
		_w2592_
	);
	LUT4 #(
		.INIT('hd11d)
	) name2130 (
		\P2_reg2_reg[26]/NET0131 ,
		_w2039_,
		_w2463_,
		_w2506_,
		_w2593_
	);
	LUT4 #(
		.INIT('hf351)
	) name2131 (
		_w2188_,
		_w2193_,
		_w2592_,
		_w2593_,
		_w2594_
	);
	LUT4 #(
		.INIT('h3111)
	) name2132 (
		_w1489_,
		_w2583_,
		_w2591_,
		_w2594_,
		_w2595_
	);
	LUT3 #(
		.INIT('hce)
	) name2133 (
		\P1_state_reg[0]/NET0131 ,
		_w2582_,
		_w2595_,
		_w2596_
	);
	LUT4 #(
		.INIT('h70d0)
	) name2134 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg0_reg[29]/NET0131 ,
		_w1476_,
		_w2597_
	);
	LUT2 #(
		.INIT('h8)
	) name2135 (
		\P2_reg0_reg[29]/NET0131 ,
		_w1487_,
		_w2598_
	);
	LUT3 #(
		.INIT('hb0)
	) name2136 (
		_w2019_,
		_w2022_,
		_w2042_,
		_w2599_
	);
	LUT4 #(
		.INIT('h3dfd)
	) name2137 (
		\P2_reg0_reg[30]/NET0131 ,
		_w488_,
		_w494_,
		_w2046_,
		_w2600_
	);
	LUT4 #(
		.INIT('hf53f)
	) name2138 (
		\P2_reg1_reg[30]/NET0131 ,
		\P2_reg2_reg[30]/NET0131 ,
		_w488_,
		_w494_,
		_w2601_
	);
	LUT2 #(
		.INIT('h8)
	) name2139 (
		_w2600_,
		_w2601_,
		_w2602_
	);
	LUT2 #(
		.INIT('h7)
	) name2140 (
		_w2600_,
		_w2601_,
		_w2603_
	);
	LUT4 #(
		.INIT('h0080)
	) name2141 (
		_w2073_,
		_w2074_,
		_w2076_,
		_w2602_,
		_w2604_
	);
	LUT3 #(
		.INIT('he3)
	) name2142 (
		\P2_B_reg/NET0131 ,
		_w1505_,
		_w1508_,
		_w2605_
	);
	LUT4 #(
		.INIT('h3312)
	) name2143 (
		_w2077_,
		_w2599_,
		_w2602_,
		_w2605_,
		_w2606_
	);
	LUT4 #(
		.INIT('h08c8)
	) name2144 (
		\P2_reg0_reg[29]/NET0131 ,
		_w2081_,
		_w2272_,
		_w2606_,
		_w2607_
	);
	LUT2 #(
		.INIT('h8)
	) name2145 (
		\P1_datao_reg[29]/NET0131 ,
		\si[29]_pad ,
		_w2608_
	);
	LUT4 #(
		.INIT('h135f)
	) name2146 (
		\P1_datao_reg[27]/NET0131 ,
		\P1_datao_reg[28]/NET0131 ,
		\si[27]_pad ,
		\si[28]_pad ,
		_w2609_
	);
	LUT4 #(
		.INIT('hec00)
	) name2147 (
		_w1898_,
		_w1928_,
		_w1929_,
		_w1964_,
		_w2610_
	);
	LUT4 #(
		.INIT('ha0b0)
	) name2148 (
		_w1963_,
		_w1965_,
		_w2609_,
		_w2610_,
		_w2611_
	);
	LUT2 #(
		.INIT('h1)
	) name2149 (
		_w2009_,
		_w2611_,
		_w2612_
	);
	LUT4 #(
		.INIT('hfac8)
	) name2150 (
		\P1_datao_reg[27]/NET0131 ,
		\P1_datao_reg[28]/NET0131 ,
		\si[27]_pad ,
		\si[28]_pad ,
		_w2613_
	);
	LUT4 #(
		.INIT('h8000)
	) name2151 (
		_w1894_,
		_w1929_,
		_w1964_,
		_w2613_,
		_w2614_
	);
	LUT3 #(
		.INIT('h23)
	) name2152 (
		_w1881_,
		_w2612_,
		_w2614_,
		_w2615_
	);
	LUT4 #(
		.INIT('h9565)
	) name2153 (
		\P1_datao_reg[29]/NET0131 ,
		\si[29]_pad ,
		_w542_,
		_w2615_,
		_w2616_
	);
	LUT2 #(
		.INIT('h1)
	) name2154 (
		_w1509_,
		_w2616_,
		_w2617_
	);
	LUT3 #(
		.INIT('h32)
	) name2155 (
		_w1509_,
		_w2049_,
		_w2616_,
		_w2618_
	);
	LUT3 #(
		.INIT('h04)
	) name2156 (
		_w1509_,
		_w2049_,
		_w2616_,
		_w2619_
	);
	LUT3 #(
		.INIT('hc9)
	) name2157 (
		_w1509_,
		_w2049_,
		_w2616_,
		_w2620_
	);
	LUT3 #(
		.INIT('h8c)
	) name2158 (
		_w2563_,
		_w2560_,
		_w2554_,
		_w2621_
	);
	LUT3 #(
		.INIT('hc4)
	) name2159 (
		_w2375_,
		_w2552_,
		_w2555_,
		_w2622_
	);
	LUT2 #(
		.INIT('h2)
	) name2160 (
		_w2558_,
		_w2622_,
		_w2623_
	);
	LUT3 #(
		.INIT('h10)
	) name2161 (
		_w1509_,
		_w2017_,
		_w2023_,
		_w2624_
	);
	LUT3 #(
		.INIT('h04)
	) name2162 (
		_w2166_,
		_w2381_,
		_w2624_,
		_w2625_
	);
	LUT2 #(
		.INIT('h8)
	) name2163 (
		_w2551_,
		_w2625_,
		_w2626_
	);
	LUT3 #(
		.INIT('h04)
	) name2164 (
		_w2166_,
		_w2384_,
		_w2624_,
		_w2627_
	);
	LUT3 #(
		.INIT('h0e)
	) name2165 (
		_w1509_,
		_w2017_,
		_w2023_,
		_w2628_
	);
	LUT3 #(
		.INIT('h0d)
	) name2166 (
		_w2180_,
		_w2624_,
		_w2628_,
		_w2629_
	);
	LUT4 #(
		.INIT('h0b00)
	) name2167 (
		_w2564_,
		_w2625_,
		_w2627_,
		_w2629_,
		_w2630_
	);
	LUT4 #(
		.INIT('h4f00)
	) name2168 (
		_w2621_,
		_w2623_,
		_w2626_,
		_w2630_,
		_w2631_
	);
	LUT4 #(
		.INIT('h1dd1)
	) name2169 (
		\P2_reg0_reg[29]/NET0131 ,
		_w2277_,
		_w2620_,
		_w2631_,
		_w2632_
	);
	LUT4 #(
		.INIT('h3f7d)
	) name2170 (
		_w1811_,
		_w2033_,
		_w2035_,
		_w2036_,
		_w2633_
	);
	LUT4 #(
		.INIT('hfe00)
	) name2171 (
		_w1491_,
		_w1493_,
		_w1496_,
		_w2084_,
		_w2634_
	);
	LUT2 #(
		.INIT('h2)
	) name2172 (
		_w2633_,
		_w2634_,
		_w2635_
	);
	LUT3 #(
		.INIT('ha2)
	) name2173 (
		\P2_reg0_reg[29]/NET0131 ,
		_w2633_,
		_w2634_,
		_w2636_
	);
	LUT4 #(
		.INIT('h0040)
	) name2174 (
		_w1509_,
		_w2084_,
		_w2277_,
		_w2616_,
		_w2637_
	);
	LUT2 #(
		.INIT('h1)
	) name2175 (
		_w2636_,
		_w2637_,
		_w2638_
	);
	LUT4 #(
		.INIT('h0e00)
	) name2176 (
		_w2192_,
		_w2632_,
		_w2607_,
		_w2638_,
		_w2639_
	);
	LUT3 #(
		.INIT('h8c)
	) name2177 (
		_w2536_,
		_w2539_,
		_w2541_,
		_w2640_
	);
	LUT3 #(
		.INIT('hc4)
	) name2178 (
		_w2324_,
		_w2537_,
		_w2542_,
		_w2641_
	);
	LUT2 #(
		.INIT('h2)
	) name2179 (
		_w2545_,
		_w2641_,
		_w2642_
	);
	LUT2 #(
		.INIT('h1)
	) name2180 (
		_w1977_,
		_w2025_,
		_w2643_
	);
	LUT3 #(
		.INIT('h80)
	) name2181 (
		_w2328_,
		_w2329_,
		_w2332_,
		_w2644_
	);
	LUT2 #(
		.INIT('h8)
	) name2182 (
		_w2643_,
		_w2644_,
		_w2645_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name2183 (
		_w2328_,
		_w2329_,
		_w2338_,
		_w2336_,
		_w2646_
	);
	LUT3 #(
		.INIT('h32)
	) name2184 (
		_w2006_,
		_w2025_,
		_w2026_,
		_w2647_
	);
	LUT4 #(
		.INIT('h003b)
	) name2185 (
		_w2339_,
		_w2643_,
		_w2646_,
		_w2647_,
		_w2648_
	);
	LUT4 #(
		.INIT('h4f00)
	) name2186 (
		_w2640_,
		_w2642_,
		_w2645_,
		_w2648_,
		_w2649_
	);
	LUT4 #(
		.INIT('hd11d)
	) name2187 (
		\P2_reg0_reg[29]/NET0131 ,
		_w2277_,
		_w2620_,
		_w2649_,
		_w2650_
	);
	LUT4 #(
		.INIT('hd11d)
	) name2188 (
		\P2_reg0_reg[29]/NET0131 ,
		_w2272_,
		_w2620_,
		_w2649_,
		_w2651_
	);
	LUT4 #(
		.INIT('hfa32)
	) name2189 (
		_w2276_,
		_w2290_,
		_w2650_,
		_w2651_,
		_w2652_
	);
	LUT4 #(
		.INIT('h3111)
	) name2190 (
		_w1489_,
		_w2598_,
		_w2639_,
		_w2652_,
		_w2653_
	);
	LUT3 #(
		.INIT('hce)
	) name2191 (
		\P1_state_reg[0]/NET0131 ,
		_w2597_,
		_w2653_,
		_w2654_
	);
	LUT4 #(
		.INIT('h70d0)
	) name2192 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg1_reg[29]/NET0131 ,
		_w1476_,
		_w2655_
	);
	LUT2 #(
		.INIT('h8)
	) name2193 (
		\P2_reg1_reg[29]/NET0131 ,
		_w1487_,
		_w2656_
	);
	LUT4 #(
		.INIT('hd11d)
	) name2194 (
		\P2_reg1_reg[29]/NET0131 ,
		_w2039_,
		_w2620_,
		_w2649_,
		_w2657_
	);
	LUT2 #(
		.INIT('h2)
	) name2195 (
		_w2038_,
		_w2657_,
		_w2658_
	);
	LUT4 #(
		.INIT('h1dd1)
	) name2196 (
		\P2_reg1_reg[29]/NET0131 ,
		_w2039_,
		_w2620_,
		_w2631_,
		_w2659_
	);
	LUT4 #(
		.INIT('hf100)
	) name2197 (
		_w1491_,
		_w1493_,
		_w1496_,
		_w2084_,
		_w2660_
	);
	LUT2 #(
		.INIT('h2)
	) name2198 (
		_w2633_,
		_w2660_,
		_w2661_
	);
	LUT3 #(
		.INIT('ha2)
	) name2199 (
		\P2_reg1_reg[29]/NET0131 ,
		_w2633_,
		_w2660_,
		_w2662_
	);
	LUT4 #(
		.INIT('h0040)
	) name2200 (
		_w1509_,
		_w2039_,
		_w2084_,
		_w2616_,
		_w2663_
	);
	LUT2 #(
		.INIT('h1)
	) name2201 (
		_w2662_,
		_w2663_,
		_w2664_
	);
	LUT3 #(
		.INIT('hd0)
	) name2202 (
		_w2193_,
		_w2659_,
		_w2664_,
		_w2665_
	);
	LUT4 #(
		.INIT('h20e0)
	) name2203 (
		\P2_reg1_reg[29]/NET0131 ,
		_w1497_,
		_w2081_,
		_w2606_,
		_w2666_
	);
	LUT4 #(
		.INIT('h1dd1)
	) name2204 (
		\P2_reg1_reg[29]/NET0131 ,
		_w1497_,
		_w2620_,
		_w2631_,
		_w2667_
	);
	LUT3 #(
		.INIT('h31)
	) name2205 (
		_w2188_,
		_w2666_,
		_w2667_,
		_w2668_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name2206 (
		_w1489_,
		_w2658_,
		_w2665_,
		_w2668_,
		_w2669_
	);
	LUT4 #(
		.INIT('heeec)
	) name2207 (
		\P1_state_reg[0]/NET0131 ,
		_w2655_,
		_w2656_,
		_w2669_,
		_w2670_
	);
	LUT4 #(
		.INIT('h70d0)
	) name2208 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg2_reg[29]/NET0131 ,
		_w1476_,
		_w2671_
	);
	LUT2 #(
		.INIT('h8)
	) name2209 (
		\P2_reg2_reg[29]/NET0131 ,
		_w1487_,
		_w2672_
	);
	LUT4 #(
		.INIT('hd11d)
	) name2210 (
		\P2_reg2_reg[29]/NET0131 ,
		_w1497_,
		_w2620_,
		_w2649_,
		_w2673_
	);
	LUT2 #(
		.INIT('h2)
	) name2211 (
		_w2038_,
		_w2673_,
		_w2674_
	);
	LUT4 #(
		.INIT('h1dd1)
	) name2212 (
		\P2_reg2_reg[29]/NET0131 ,
		_w1497_,
		_w2620_,
		_w2631_,
		_w2675_
	);
	LUT4 #(
		.INIT('h0020)
	) name2213 (
		_w1497_,
		_w1509_,
		_w2084_,
		_w2616_,
		_w2676_
	);
	LUT2 #(
		.INIT('h8)
	) name2214 (
		_w2046_,
		_w2088_,
		_w2677_
	);
	LUT4 #(
		.INIT('h0057)
	) name2215 (
		\P2_reg2_reg[29]/NET0131 ,
		_w2086_,
		_w2087_,
		_w2677_,
		_w2678_
	);
	LUT2 #(
		.INIT('h4)
	) name2216 (
		_w2676_,
		_w2678_,
		_w2679_
	);
	LUT3 #(
		.INIT('hd0)
	) name2217 (
		_w2193_,
		_w2675_,
		_w2679_,
		_w2680_
	);
	LUT4 #(
		.INIT('h20e0)
	) name2218 (
		\P2_reg2_reg[29]/NET0131 ,
		_w2039_,
		_w2081_,
		_w2606_,
		_w2681_
	);
	LUT4 #(
		.INIT('h1dd1)
	) name2219 (
		\P2_reg2_reg[29]/NET0131 ,
		_w2039_,
		_w2620_,
		_w2631_,
		_w2682_
	);
	LUT3 #(
		.INIT('h31)
	) name2220 (
		_w2188_,
		_w2681_,
		_w2682_,
		_w2683_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name2221 (
		_w1489_,
		_w2674_,
		_w2680_,
		_w2683_,
		_w2684_
	);
	LUT4 #(
		.INIT('heeec)
	) name2222 (
		\P1_state_reg[0]/NET0131 ,
		_w2671_,
		_w2672_,
		_w2684_,
		_w2685_
	);
	LUT2 #(
		.INIT('h2)
	) name2223 (
		\P1_reg0_reg[29]/NET0131 ,
		_w511_,
		_w2686_
	);
	LUT2 #(
		.INIT('h8)
	) name2224 (
		\P1_reg0_reg[29]/NET0131 ,
		_w524_,
		_w2687_
	);
	LUT3 #(
		.INIT('h01)
	) name2225 (
		_w528_,
		_w530_,
		_w533_,
		_w2688_
	);
	LUT4 #(
		.INIT('haaa8)
	) name2226 (
		\P1_reg0_reg[29]/NET0131 ,
		_w528_,
		_w530_,
		_w533_,
		_w2689_
	);
	LUT4 #(
		.INIT('h30a0)
	) name2227 (
		\P1_reg0_reg[29]/NET0131 ,
		_w1182_,
		_w1183_,
		_w2688_,
		_w2690_
	);
	LUT4 #(
		.INIT('hc0a0)
	) name2228 (
		\P1_reg0_reg[29]/NET0131 ,
		_w1134_,
		_w1136_,
		_w2688_,
		_w2691_
	);
	LUT3 #(
		.INIT('hc4)
	) name2229 (
		_w1138_,
		_w2425_,
		_w2688_,
		_w2692_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name2230 (
		\P1_reg0_reg[29]/NET0131 ,
		_w1138_,
		_w2425_,
		_w2688_,
		_w2693_
	);
	LUT3 #(
		.INIT('h07)
	) name2231 (
		_w1139_,
		_w2688_,
		_w2693_,
		_w2694_
	);
	LUT2 #(
		.INIT('h4)
	) name2232 (
		_w2691_,
		_w2694_,
		_w2695_
	);
	LUT2 #(
		.INIT('h4)
	) name2233 (
		_w2690_,
		_w2695_,
		_w2696_
	);
	LUT4 #(
		.INIT('h6500)
	) name2234 (
		_w647_,
		_w1265_,
		_w1284_,
		_w2688_,
		_w2697_
	);
	LUT3 #(
		.INIT('ha8)
	) name2235 (
		_w1286_,
		_w2689_,
		_w2697_,
		_w2698_
	);
	LUT4 #(
		.INIT('hc355)
	) name2236 (
		\P1_reg0_reg[29]/NET0131 ,
		_w647_,
		_w1102_,
		_w2688_,
		_w2699_
	);
	LUT2 #(
		.INIT('h2)
	) name2237 (
		_w1114_,
		_w2699_,
		_w2700_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name2238 (
		_w526_,
		_w2698_,
		_w2700_,
		_w2696_,
		_w2701_
	);
	LUT4 #(
		.INIT('heeec)
	) name2239 (
		\P1_state_reg[0]/NET0131 ,
		_w2686_,
		_w2687_,
		_w2701_,
		_w2702_
	);
	LUT2 #(
		.INIT('h2)
	) name2240 (
		_w1487_,
		_w1777_,
		_w2703_
	);
	LUT4 #(
		.INIT('h001f)
	) name2241 (
		_w1491_,
		_w1493_,
		_w1496_,
		_w1777_,
		_w2704_
	);
	LUT4 #(
		.INIT('hf10e)
	) name2242 (
		_w1509_,
		_w1771_,
		_w1775_,
		_w1781_,
		_w2705_
	);
	LUT4 #(
		.INIT('h7300)
	) name2243 (
		_w2536_,
		_w2538_,
		_w2541_,
		_w2543_,
		_w2706_
	);
	LUT4 #(
		.INIT('h007d)
	) name2244 (
		_w2272_,
		_w2705_,
		_w2706_,
		_w2704_,
		_w2707_
	);
	LUT2 #(
		.INIT('h1)
	) name2245 (
		_w2276_,
		_w2707_,
		_w2708_
	);
	LUT4 #(
		.INIT('h00fe)
	) name2246 (
		_w1491_,
		_w1493_,
		_w1496_,
		_w1777_,
		_w2709_
	);
	LUT4 #(
		.INIT('h1331)
	) name2247 (
		_w2277_,
		_w2709_,
		_w2705_,
		_w2706_,
		_w2710_
	);
	LUT2 #(
		.INIT('h2)
	) name2248 (
		_w2290_,
		_w2710_,
		_w2711_
	);
	LUT4 #(
		.INIT('h7300)
	) name2249 (
		_w2563_,
		_w2553_,
		_w2554_,
		_w2556_,
		_w2712_
	);
	LUT4 #(
		.INIT('h0d07)
	) name2250 (
		_w2272_,
		_w2705_,
		_w2704_,
		_w2712_,
		_w2713_
	);
	LUT2 #(
		.INIT('h4)
	) name2251 (
		_w498_,
		_w2042_,
		_w2714_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name2252 (
		_w1697_,
		_w1838_,
		_w2066_,
		_w2067_,
		_w2715_
	);
	LUT4 #(
		.INIT('h2333)
	) name2253 (
		_w1697_,
		_w2042_,
		_w2066_,
		_w2068_,
		_w2716_
	);
	LUT4 #(
		.INIT('h8a88)
	) name2254 (
		_w2277_,
		_w2714_,
		_w2715_,
		_w2716_,
		_w2717_
	);
	LUT3 #(
		.INIT('h54)
	) name2255 (
		_w1777_,
		_w2086_,
		_w2280_,
		_w2718_
	);
	LUT3 #(
		.INIT('h0b)
	) name2256 (
		_w1776_,
		_w2283_,
		_w2718_,
		_w2719_
	);
	LUT4 #(
		.INIT('h5700)
	) name2257 (
		_w2081_,
		_w2709_,
		_w2717_,
		_w2719_,
		_w2720_
	);
	LUT3 #(
		.INIT('he0)
	) name2258 (
		_w2192_,
		_w2713_,
		_w2720_,
		_w2721_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name2259 (
		_w1489_,
		_w2711_,
		_w2708_,
		_w2721_,
		_w2722_
	);
	LUT2 #(
		.INIT('h4)
	) name2260 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[17]/NET0131 ,
		_w2723_
	);
	LUT3 #(
		.INIT('h0b)
	) name2261 (
		_w1777_,
		_w2293_,
		_w2723_,
		_w2724_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name2262 (
		\P1_state_reg[0]/NET0131 ,
		_w2703_,
		_w2722_,
		_w2724_,
		_w2725_
	);
	LUT2 #(
		.INIT('h2)
	) name2263 (
		_w1487_,
		_w1834_,
		_w2726_
	);
	LUT4 #(
		.INIT('h00fe)
	) name2264 (
		_w1491_,
		_w1493_,
		_w1496_,
		_w1834_,
		_w2727_
	);
	LUT2 #(
		.INIT('h6)
	) name2265 (
		_w1833_,
		_w1838_,
		_w2728_
	);
	LUT4 #(
		.INIT('h070d)
	) name2266 (
		_w2277_,
		_w2472_,
		_w2727_,
		_w2728_,
		_w2729_
	);
	LUT4 #(
		.INIT('h1000)
	) name2267 (
		_w1697_,
		_w1819_,
		_w2066_,
		_w2068_,
		_w2730_
	);
	LUT4 #(
		.INIT('hef00)
	) name2268 (
		_w1779_,
		_w1778_,
		_w1780_,
		_w2042_,
		_w2731_
	);
	LUT4 #(
		.INIT('h00de)
	) name2269 (
		_w1819_,
		_w2042_,
		_w2069_,
		_w2731_,
		_w2732_
	);
	LUT4 #(
		.INIT('h04c4)
	) name2270 (
		_w1834_,
		_w2081_,
		_w2277_,
		_w2732_,
		_w2733_
	);
	LUT3 #(
		.INIT('h04)
	) name2271 (
		_w1833_,
		_w2083_,
		_w2282_,
		_w2734_
	);
	LUT3 #(
		.INIT('h54)
	) name2272 (
		_w1834_,
		_w2086_,
		_w2280_,
		_w2735_
	);
	LUT2 #(
		.INIT('h1)
	) name2273 (
		_w2734_,
		_w2735_,
		_w2736_
	);
	LUT4 #(
		.INIT('h0d00)
	) name2274 (
		_w2290_,
		_w2729_,
		_w2733_,
		_w2736_,
		_w2737_
	);
	LUT4 #(
		.INIT('h001f)
	) name2275 (
		_w1491_,
		_w1493_,
		_w1496_,
		_w1834_,
		_w2738_
	);
	LUT4 #(
		.INIT('h8a20)
	) name2276 (
		_w2272_,
		_w2495_,
		_w2498_,
		_w2728_,
		_w2739_
	);
	LUT3 #(
		.INIT('h54)
	) name2277 (
		_w2192_,
		_w2738_,
		_w2739_,
		_w2740_
	);
	LUT4 #(
		.INIT('h007d)
	) name2278 (
		_w2272_,
		_w2472_,
		_w2728_,
		_w2738_,
		_w2741_
	);
	LUT2 #(
		.INIT('h1)
	) name2279 (
		_w2276_,
		_w2741_,
		_w2742_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name2280 (
		_w1489_,
		_w2740_,
		_w2742_,
		_w2737_,
		_w2743_
	);
	LUT2 #(
		.INIT('h4)
	) name2281 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[18]/NET0131 ,
		_w2744_
	);
	LUT3 #(
		.INIT('h0b)
	) name2282 (
		_w1834_,
		_w2293_,
		_w2744_,
		_w2745_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name2283 (
		\P1_state_reg[0]/NET0131 ,
		_w2726_,
		_w2743_,
		_w2745_,
		_w2746_
	);
	LUT2 #(
		.INIT('h2)
	) name2284 (
		_w1487_,
		_w1815_,
		_w2747_
	);
	LUT4 #(
		.INIT('h001f)
	) name2285 (
		_w1491_,
		_w1493_,
		_w1496_,
		_w1815_,
		_w2748_
	);
	LUT2 #(
		.INIT('h6)
	) name2286 (
		_w1813_,
		_w1819_,
		_w2749_
	);
	LUT4 #(
		.INIT('h208a)
	) name2287 (
		_w2272_,
		_w2319_,
		_w2327_,
		_w2749_,
		_w2750_
	);
	LUT3 #(
		.INIT('h54)
	) name2288 (
		_w2276_,
		_w2748_,
		_w2750_,
		_w2751_
	);
	LUT4 #(
		.INIT('h00fe)
	) name2289 (
		_w1491_,
		_w1493_,
		_w1496_,
		_w1815_,
		_w2752_
	);
	LUT4 #(
		.INIT('h208a)
	) name2290 (
		_w2277_,
		_w2319_,
		_w2327_,
		_w2749_,
		_w2753_
	);
	LUT3 #(
		.INIT('ha8)
	) name2291 (
		_w2290_,
		_w2752_,
		_w2753_,
		_w2754_
	);
	LUT4 #(
		.INIT('hef00)
	) name2292 (
		_w1836_,
		_w1835_,
		_w1837_,
		_w2042_,
		_w2755_
	);
	LUT4 #(
		.INIT('h00de)
	) name2293 (
		_w1872_,
		_w2042_,
		_w2730_,
		_w2755_,
		_w2756_
	);
	LUT4 #(
		.INIT('h04c4)
	) name2294 (
		_w1815_,
		_w2081_,
		_w2277_,
		_w2756_,
		_w2757_
	);
	LUT4 #(
		.INIT('h00d7)
	) name2295 (
		_w2272_,
		_w2378_,
		_w2749_,
		_w2748_,
		_w2758_
	);
	LUT3 #(
		.INIT('h54)
	) name2296 (
		_w1815_,
		_w2086_,
		_w2280_,
		_w2759_
	);
	LUT3 #(
		.INIT('h04)
	) name2297 (
		_w1813_,
		_w2083_,
		_w2282_,
		_w2760_
	);
	LUT2 #(
		.INIT('h1)
	) name2298 (
		_w2759_,
		_w2760_,
		_w2761_
	);
	LUT4 #(
		.INIT('h3200)
	) name2299 (
		_w2192_,
		_w2757_,
		_w2758_,
		_w2761_,
		_w2762_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name2300 (
		_w1489_,
		_w2754_,
		_w2751_,
		_w2762_,
		_w2763_
	);
	LUT4 #(
		.INIT('hb9b3)
	) name2301 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[19]/NET0131 ,
		_w1477_,
		_w1814_,
		_w2764_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name2302 (
		\P1_state_reg[0]/NET0131 ,
		_w2747_,
		_w2763_,
		_w2764_,
		_w2765_
	);
	LUT2 #(
		.INIT('h8)
	) name2303 (
		_w524_,
		_w1056_,
		_w2766_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name2304 (
		_w1327_,
		_w1333_,
		_w1338_,
		_w2199_,
		_w2767_
	);
	LUT4 #(
		.INIT('h001f)
	) name2305 (
		_w528_,
		_w530_,
		_w533_,
		_w1056_,
		_w2768_
	);
	LUT2 #(
		.INIT('h2)
	) name2306 (
		_w1286_,
		_w2768_,
		_w2769_
	);
	LUT4 #(
		.INIT('h7b00)
	) name2307 (
		_w1425_,
		_w2197_,
		_w2767_,
		_w2769_,
		_w2770_
	);
	LUT4 #(
		.INIT('h08aa)
	) name2308 (
		_w2211_,
		_w2214_,
		_w2219_,
		_w2234_,
		_w2771_
	);
	LUT4 #(
		.INIT('h0070)
	) name2309 (
		_w2215_,
		_w2230_,
		_w2238_,
		_w2771_,
		_w2772_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name2310 (
		_w1425_,
		_w2245_,
		_w2249_,
		_w2772_,
		_w2773_
	);
	LUT4 #(
		.INIT('h5010)
	) name2311 (
		_w1425_,
		_w2245_,
		_w2249_,
		_w2772_,
		_w2774_
	);
	LUT3 #(
		.INIT('h02)
	) name2312 (
		_w1114_,
		_w2774_,
		_w2773_,
		_w2775_
	);
	LUT2 #(
		.INIT('h2)
	) name2313 (
		_w537_,
		_w1051_,
		_w2776_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name2314 (
		_w977_,
		_w1170_,
		_w1161_,
		_w1163_,
		_w2777_
	);
	LUT4 #(
		.INIT('h1555)
	) name2315 (
		_w537_,
		_w1161_,
		_w1163_,
		_w1171_,
		_w2778_
	);
	LUT4 #(
		.INIT('h8a88)
	) name2316 (
		_w1183_,
		_w2776_,
		_w2777_,
		_w2778_,
		_w2779_
	);
	LUT3 #(
		.INIT('h90)
	) name2317 (
		_w1055_,
		_w1128_,
		_w1136_,
		_w2780_
	);
	LUT2 #(
		.INIT('h1)
	) name2318 (
		_w2779_,
		_w2780_,
		_w2781_
	);
	LUT3 #(
		.INIT('h10)
	) name2319 (
		_w541_,
		_w1054_,
		_w2261_,
		_w2782_
	);
	LUT3 #(
		.INIT('h01)
	) name2320 (
		_w1286_,
		_w2197_,
		_w2259_,
		_w2783_
	);
	LUT3 #(
		.INIT('ha2)
	) name2321 (
		_w1056_,
		_w2257_,
		_w2783_,
		_w2784_
	);
	LUT2 #(
		.INIT('h1)
	) name2322 (
		_w2782_,
		_w2784_,
		_w2785_
	);
	LUT4 #(
		.INIT('h7500)
	) name2323 (
		_w2197_,
		_w2775_,
		_w2781_,
		_w2785_,
		_w2786_
	);
	LUT4 #(
		.INIT('h1311)
	) name2324 (
		_w526_,
		_w2766_,
		_w2770_,
		_w2786_,
		_w2787_
	);
	LUT2 #(
		.INIT('h2)
	) name2325 (
		\P1_reg3_reg[24]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w2788_
	);
	LUT3 #(
		.INIT('h07)
	) name2326 (
		_w1056_,
		_w1294_,
		_w2788_,
		_w2789_
	);
	LUT3 #(
		.INIT('h2f)
	) name2327 (
		\P1_state_reg[0]/NET0131 ,
		_w2787_,
		_w2789_,
		_w2790_
	);
	LUT2 #(
		.INIT('h2)
	) name2328 (
		_w1487_,
		_w1917_,
		_w2791_
	);
	LUT4 #(
		.INIT('h001f)
	) name2329 (
		_w1491_,
		_w1493_,
		_w1496_,
		_w1917_,
		_w2792_
	);
	LUT3 #(
		.INIT('h1e)
	) name2330 (
		_w1509_,
		_w1916_,
		_w1921_,
		_w2793_
	);
	LUT4 #(
		.INIT('h4f00)
	) name2331 (
		_w2492_,
		_w2493_,
		_w2494_,
		_w2496_,
		_w2794_
	);
	LUT2 #(
		.INIT('h8)
	) name2332 (
		_w2491_,
		_w2499_,
		_w2795_
	);
	LUT3 #(
		.INIT('he0)
	) name2333 (
		_w2148_,
		_w2497_,
		_w2499_,
		_w2796_
	);
	LUT2 #(
		.INIT('h2)
	) name2334 (
		_w2502_,
		_w2796_,
		_w2797_
	);
	LUT4 #(
		.INIT('h9a55)
	) name2335 (
		_w2793_,
		_w2794_,
		_w2795_,
		_w2797_,
		_w2798_
	);
	LUT4 #(
		.INIT('h0131)
	) name2336 (
		_w1917_,
		_w2192_,
		_w2272_,
		_w2798_,
		_w2799_
	);
	LUT3 #(
		.INIT('h54)
	) name2337 (
		_w1917_,
		_w2086_,
		_w2280_,
		_w2800_
	);
	LUT4 #(
		.INIT('h0010)
	) name2338 (
		_w1509_,
		_w1916_,
		_w2083_,
		_w2282_,
		_w2801_
	);
	LUT2 #(
		.INIT('h1)
	) name2339 (
		_w2800_,
		_w2801_,
		_w2802_
	);
	LUT2 #(
		.INIT('h4)
	) name2340 (
		_w2799_,
		_w2802_,
		_w2803_
	);
	LUT2 #(
		.INIT('h8)
	) name2341 (
		_w2464_,
		_w2473_,
		_w2804_
	);
	LUT4 #(
		.INIT('h4f00)
	) name2342 (
		_w2467_,
		_w2468_,
		_w2469_,
		_w2804_,
		_w2805_
	);
	LUT3 #(
		.INIT('hd0)
	) name2343 (
		_w1850_,
		_w2470_,
		_w2473_,
		_w2806_
	);
	LUT2 #(
		.INIT('h2)
	) name2344 (
		_w2476_,
		_w2806_,
		_w2807_
	);
	LUT4 #(
		.INIT('h2822)
	) name2345 (
		_w2272_,
		_w2793_,
		_w2805_,
		_w2807_,
		_w2808_
	);
	LUT3 #(
		.INIT('h54)
	) name2346 (
		_w2276_,
		_w2792_,
		_w2808_,
		_w2809_
	);
	LUT4 #(
		.INIT('h00fe)
	) name2347 (
		_w1491_,
		_w1493_,
		_w1496_,
		_w1917_,
		_w2810_
	);
	LUT4 #(
		.INIT('h2822)
	) name2348 (
		_w2277_,
		_w2793_,
		_w2805_,
		_w2807_,
		_w2811_
	);
	LUT3 #(
		.INIT('ha8)
	) name2349 (
		_w2290_,
		_w2810_,
		_w2811_,
		_w2812_
	);
	LUT3 #(
		.INIT('h40)
	) name2350 (
		_w1921_,
		_w2070_,
		_w2730_,
		_w2813_
	);
	LUT4 #(
		.INIT('h1000)
	) name2351 (
		_w1907_,
		_w1921_,
		_w2070_,
		_w2730_,
		_w2814_
	);
	LUT4 #(
		.INIT('hef00)
	) name2352 (
		_w1887_,
		_w1886_,
		_w1888_,
		_w2042_,
		_w2815_
	);
	LUT4 #(
		.INIT('h00de)
	) name2353 (
		_w1907_,
		_w2042_,
		_w2813_,
		_w2815_,
		_w2816_
	);
	LUT4 #(
		.INIT('h04c4)
	) name2354 (
		_w1917_,
		_w2081_,
		_w2277_,
		_w2816_,
		_w2817_
	);
	LUT3 #(
		.INIT('h01)
	) name2355 (
		_w2812_,
		_w2817_,
		_w2809_,
		_w2818_
	);
	LUT4 #(
		.INIT('h3111)
	) name2356 (
		_w1489_,
		_w2791_,
		_w2803_,
		_w2818_,
		_w2819_
	);
	LUT4 #(
		.INIT('hb9b3)
	) name2357 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[22]/NET0131 ,
		_w1477_,
		_w1884_,
		_w2820_
	);
	LUT3 #(
		.INIT('h2f)
	) name2358 (
		\P1_state_reg[0]/NET0131 ,
		_w2819_,
		_w2820_,
		_w2821_
	);
	LUT4 #(
		.INIT('h70d0)
	) name2359 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg2_reg[22]/NET0131 ,
		_w1476_,
		_w2822_
	);
	LUT2 #(
		.INIT('h8)
	) name2360 (
		\P2_reg2_reg[22]/NET0131 ,
		_w1487_,
		_w2823_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name2361 (
		\P2_reg2_reg[22]/NET0131 ,
		_w1491_,
		_w1493_,
		_w1496_,
		_w2824_
	);
	LUT4 #(
		.INIT('h20e0)
	) name2362 (
		\P2_reg2_reg[22]/NET0131 ,
		_w1497_,
		_w2193_,
		_w2798_,
		_w2825_
	);
	LUT3 #(
		.INIT('ha8)
	) name2363 (
		\P2_reg2_reg[22]/NET0131 ,
		_w2086_,
		_w2087_,
		_w2826_
	);
	LUT2 #(
		.INIT('h4)
	) name2364 (
		_w1917_,
		_w2088_,
		_w2827_
	);
	LUT4 #(
		.INIT('h00ef)
	) name2365 (
		_w1509_,
		_w1916_,
		_w2085_,
		_w2827_,
		_w2828_
	);
	LUT2 #(
		.INIT('h4)
	) name2366 (
		_w2826_,
		_w2828_,
		_w2829_
	);
	LUT2 #(
		.INIT('h4)
	) name2367 (
		_w2825_,
		_w2829_,
		_w2830_
	);
	LUT4 #(
		.INIT('h20e0)
	) name2368 (
		\P2_reg2_reg[22]/NET0131 ,
		_w2039_,
		_w2188_,
		_w2798_,
		_w2831_
	);
	LUT4 #(
		.INIT('h2822)
	) name2369 (
		_w1497_,
		_w2793_,
		_w2805_,
		_w2807_,
		_w2832_
	);
	LUT3 #(
		.INIT('ha8)
	) name2370 (
		_w2038_,
		_w2824_,
		_w2832_,
		_w2833_
	);
	LUT4 #(
		.INIT('h20e0)
	) name2371 (
		\P2_reg2_reg[22]/NET0131 ,
		_w2039_,
		_w2081_,
		_w2816_,
		_w2834_
	);
	LUT3 #(
		.INIT('h01)
	) name2372 (
		_w2833_,
		_w2834_,
		_w2831_,
		_w2835_
	);
	LUT4 #(
		.INIT('h3111)
	) name2373 (
		_w1489_,
		_w2823_,
		_w2830_,
		_w2835_,
		_w2836_
	);
	LUT3 #(
		.INIT('hce)
	) name2374 (
		\P1_state_reg[0]/NET0131 ,
		_w2822_,
		_w2836_,
		_w2837_
	);
	LUT4 #(
		.INIT('h60c0)
	) name2375 (
		\P1_reg3_reg[26]/NET0131 ,
		\P1_reg3_reg[27]/NET0131 ,
		_w524_,
		_w971_,
		_w2838_
	);
	LUT2 #(
		.INIT('h2)
	) name2376 (
		_w1035_,
		_w2197_,
		_w2839_
	);
	LUT4 #(
		.INIT('h0b00)
	) name2377 (
		_w738_,
		_w745_,
		_w1188_,
		_w1191_,
		_w2840_
	);
	LUT4 #(
		.INIT('h0001)
	) name2378 (
		_w1196_,
		_w1203_,
		_w1204_,
		_w1234_,
		_w2841_
	);
	LUT3 #(
		.INIT('h45)
	) name2379 (
		_w1199_,
		_w1231_,
		_w1235_,
		_w2842_
	);
	LUT4 #(
		.INIT('h1f00)
	) name2380 (
		_w1224_,
		_w1228_,
		_w2841_,
		_w2842_,
		_w2843_
	);
	LUT2 #(
		.INIT('h8)
	) name2381 (
		_w1192_,
		_w1195_,
		_w2844_
	);
	LUT3 #(
		.INIT('h07)
	) name2382 (
		_w1192_,
		_w1201_,
		_w1240_,
		_w2845_
	);
	LUT4 #(
		.INIT('h000b)
	) name2383 (
		_w738_,
		_w745_,
		_w1188_,
		_w1242_,
		_w2846_
	);
	LUT4 #(
		.INIT('h0051)
	) name2384 (
		_w1246_,
		_w2840_,
		_w2845_,
		_w2846_,
		_w2847_
	);
	LUT4 #(
		.INIT('hdf00)
	) name2385 (
		_w2840_,
		_w2843_,
		_w2844_,
		_w2847_,
		_w2848_
	);
	LUT4 #(
		.INIT('h0001)
	) name2386 (
		_w1185_,
		_w1186_,
		_w1252_,
		_w1253_,
		_w2849_
	);
	LUT4 #(
		.INIT('h00ef)
	) name2387 (
		_w541_,
		_w968_,
		_w977_,
		_w1259_,
		_w2850_
	);
	LUT3 #(
		.INIT('h10)
	) name2388 (
		_w1255_,
		_w1256_,
		_w2850_,
		_w2851_
	);
	LUT4 #(
		.INIT('h1000)
	) name2389 (
		_w1255_,
		_w1256_,
		_w2849_,
		_w2850_,
		_w2852_
	);
	LUT3 #(
		.INIT('h07)
	) name2390 (
		_w1249_,
		_w1254_,
		_w1268_,
		_w2853_
	);
	LUT4 #(
		.INIT('h7100)
	) name2391 (
		_w1055_,
		_w1059_,
		_w1271_,
		_w2850_,
		_w2854_
	);
	LUT4 #(
		.INIT('h0501)
	) name2392 (
		_w1281_,
		_w2851_,
		_w2854_,
		_w2853_,
		_w2855_
	);
	LUT4 #(
		.INIT('h9a55)
	) name2393 (
		_w1428_,
		_w2848_,
		_w2852_,
		_w2855_,
		_w2856_
	);
	LUT4 #(
		.INIT('h08c8)
	) name2394 (
		_w1035_,
		_w1286_,
		_w2197_,
		_w2856_,
		_w2857_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name2395 (
		_w998_,
		_w1034_,
		_w1128_,
		_w1129_,
		_w2858_
	);
	LUT4 #(
		.INIT('h0040)
	) name2396 (
		_w1132_,
		_w1136_,
		_w2197_,
		_w2858_,
		_w2859_
	);
	LUT4 #(
		.INIT('h0f01)
	) name2397 (
		_w1136_,
		_w1138_,
		_w1141_,
		_w2197_,
		_w2860_
	);
	LUT2 #(
		.INIT('h2)
	) name2398 (
		_w1035_,
		_w2860_,
		_w2861_
	);
	LUT3 #(
		.INIT('h10)
	) name2399 (
		_w541_,
		_w1033_,
		_w2261_,
		_w2862_
	);
	LUT2 #(
		.INIT('h1)
	) name2400 (
		_w2861_,
		_w2862_,
		_w2863_
	);
	LUT2 #(
		.INIT('h4)
	) name2401 (
		_w2859_,
		_w2863_,
		_w2864_
	);
	LUT2 #(
		.INIT('h4)
	) name2402 (
		_w2857_,
		_w2864_,
		_w2865_
	);
	LUT4 #(
		.INIT('h1500)
	) name2403 (
		_w724_,
		_w738_,
		_w745_,
		_w793_,
		_w2866_
	);
	LUT3 #(
		.INIT('h40)
	) name2404 (
		_w872_,
		_w896_,
		_w940_,
		_w2867_
	);
	LUT3 #(
		.INIT('hb0)
	) name2405 (
		_w899_,
		_w940_,
		_w945_,
		_w2868_
	);
	LUT4 #(
		.INIT('h0001)
	) name2406 (
		_w828_,
		_w908_,
		_w919_,
		_w950_,
		_w2869_
	);
	LUT3 #(
		.INIT('h45)
	) name2407 (
		_w844_,
		_w948_,
		_w951_,
		_w2870_
	);
	LUT4 #(
		.INIT('h4f00)
	) name2408 (
		_w2867_,
		_w2868_,
		_w2869_,
		_w2870_,
		_w2871_
	);
	LUT2 #(
		.INIT('h8)
	) name2409 (
		_w768_,
		_w815_,
		_w2872_
	);
	LUT3 #(
		.INIT('hd0)
	) name2410 (
		_w768_,
		_w845_,
		_w955_,
		_w2873_
	);
	LUT4 #(
		.INIT('h0015)
	) name2411 (
		_w724_,
		_w738_,
		_w745_,
		_w956_,
		_w2874_
	);
	LUT4 #(
		.INIT('h00a2)
	) name2412 (
		_w960_,
		_w2866_,
		_w2873_,
		_w2874_,
		_w2875_
	);
	LUT4 #(
		.INIT('hdf00)
	) name2413 (
		_w2866_,
		_w2871_,
		_w2872_,
		_w2875_,
		_w2876_
	);
	LUT3 #(
		.INIT('h02)
	) name2414 (
		_w1007_,
		_w1053_,
		_w1061_,
		_w2877_
	);
	LUT4 #(
		.INIT('h0001)
	) name2415 (
		_w681_,
		_w708_,
		_w1072_,
		_w1080_,
		_w2878_
	);
	LUT4 #(
		.INIT('h0200)
	) name2416 (
		_w1007_,
		_w1053_,
		_w1061_,
		_w2878_,
		_w2879_
	);
	LUT3 #(
		.INIT('hb0)
	) name2417 (
		_w963_,
		_w1081_,
		_w1086_,
		_w2880_
	);
	LUT4 #(
		.INIT('h8a08)
	) name2418 (
		_w1007_,
		_w1055_,
		_w1059_,
		_w1089_,
		_w2881_
	);
	LUT4 #(
		.INIT('h0a02)
	) name2419 (
		_w1096_,
		_w2877_,
		_w2881_,
		_w2880_,
		_w2882_
	);
	LUT4 #(
		.INIT('h65aa)
	) name2420 (
		_w1428_,
		_w2876_,
		_w2879_,
		_w2882_,
		_w2883_
	);
	LUT4 #(
		.INIT('h08c8)
	) name2421 (
		_w1035_,
		_w1114_,
		_w2197_,
		_w2883_,
		_w2884_
	);
	LUT4 #(
		.INIT('h1444)
	) name2422 (
		_w537_,
		_w1023_,
		_w1172_,
		_w1173_,
		_w2885_
	);
	LUT3 #(
		.INIT('h20)
	) name2423 (
		_w537_,
		_w1000_,
		_w1003_,
		_w2886_
	);
	LUT4 #(
		.INIT('h3331)
	) name2424 (
		_w2197_,
		_w2839_,
		_w2885_,
		_w2886_,
		_w2887_
	);
	LUT3 #(
		.INIT('h31)
	) name2425 (
		_w1183_,
		_w2884_,
		_w2887_,
		_w2888_
	);
	LUT4 #(
		.INIT('h3111)
	) name2426 (
		_w526_,
		_w2838_,
		_w2865_,
		_w2888_,
		_w2889_
	);
	LUT2 #(
		.INIT('h2)
	) name2427 (
		\P1_reg3_reg[27]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w2890_
	);
	LUT4 #(
		.INIT('h6c00)
	) name2428 (
		\P1_reg3_reg[26]/NET0131 ,
		\P1_reg3_reg[27]/NET0131 ,
		_w971_,
		_w1294_,
		_w2891_
	);
	LUT2 #(
		.INIT('h1)
	) name2429 (
		_w2890_,
		_w2891_,
		_w2892_
	);
	LUT3 #(
		.INIT('h2f)
	) name2430 (
		\P1_state_reg[0]/NET0131 ,
		_w2889_,
		_w2892_,
		_w2893_
	);
	LUT2 #(
		.INIT('h2)
	) name2431 (
		_w1487_,
		_w1972_,
		_w2894_
	);
	LUT4 #(
		.INIT('h00fe)
	) name2432 (
		_w1491_,
		_w1493_,
		_w1496_,
		_w1972_,
		_w2895_
	);
	LUT4 #(
		.INIT('h007d)
	) name2433 (
		_w2277_,
		_w2301_,
		_w2342_,
		_w2895_,
		_w2896_
	);
	LUT2 #(
		.INIT('h2)
	) name2434 (
		_w2290_,
		_w2896_,
		_w2897_
	);
	LUT4 #(
		.INIT('h001f)
	) name2435 (
		_w1491_,
		_w1493_,
		_w1496_,
		_w1972_,
		_w2898_
	);
	LUT4 #(
		.INIT('h007d)
	) name2436 (
		_w2272_,
		_w2301_,
		_w2342_,
		_w2898_,
		_w2899_
	);
	LUT2 #(
		.INIT('h1)
	) name2437 (
		_w2276_,
		_w2899_,
		_w2900_
	);
	LUT4 #(
		.INIT('h80a2)
	) name2438 (
		_w2272_,
		_w2387_,
		_w2301_,
		_w2388_,
		_w2901_
	);
	LUT4 #(
		.INIT('h0057)
	) name2439 (
		_w2277_,
		_w2392_,
		_w2393_,
		_w2895_,
		_w2902_
	);
	LUT3 #(
		.INIT('h54)
	) name2440 (
		_w1972_,
		_w2086_,
		_w2280_,
		_w2903_
	);
	LUT4 #(
		.INIT('h00ef)
	) name2441 (
		_w1509_,
		_w1970_,
		_w2283_,
		_w2903_,
		_w2904_
	);
	LUT3 #(
		.INIT('hd0)
	) name2442 (
		_w2081_,
		_w2902_,
		_w2904_,
		_w2905_
	);
	LUT4 #(
		.INIT('hab00)
	) name2443 (
		_w2192_,
		_w2898_,
		_w2901_,
		_w2905_,
		_w2906_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name2444 (
		_w1489_,
		_w2900_,
		_w2897_,
		_w2906_,
		_w2907_
	);
	LUT2 #(
		.INIT('h4)
	) name2445 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[27]/NET0131 ,
		_w2908_
	);
	LUT3 #(
		.INIT('h0b)
	) name2446 (
		_w1972_,
		_w2293_,
		_w2908_,
		_w2909_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name2447 (
		\P1_state_reg[0]/NET0131 ,
		_w2894_,
		_w2907_,
		_w2909_,
		_w2910_
	);
	LUT4 #(
		.INIT('h70d0)
	) name2448 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg0_reg[27]/NET0131 ,
		_w1476_,
		_w2911_
	);
	LUT2 #(
		.INIT('h8)
	) name2449 (
		\P2_reg0_reg[27]/NET0131 ,
		_w1487_,
		_w2912_
	);
	LUT4 #(
		.INIT('h1dd1)
	) name2450 (
		\P2_reg0_reg[27]/NET0131 ,
		_w2272_,
		_w2301_,
		_w2342_,
		_w2913_
	);
	LUT2 #(
		.INIT('h2)
	) name2451 (
		_w2290_,
		_w2913_,
		_w2914_
	);
	LUT4 #(
		.INIT('haaa8)
	) name2452 (
		\P2_reg0_reg[27]/NET0131 ,
		_w1491_,
		_w1493_,
		_w1496_,
		_w2915_
	);
	LUT4 #(
		.INIT('h1dd1)
	) name2453 (
		\P2_reg0_reg[27]/NET0131 ,
		_w2277_,
		_w2301_,
		_w2342_,
		_w2916_
	);
	LUT2 #(
		.INIT('h1)
	) name2454 (
		_w2276_,
		_w2916_,
		_w2917_
	);
	LUT4 #(
		.INIT('h80a2)
	) name2455 (
		_w2277_,
		_w2387_,
		_w2301_,
		_w2388_,
		_w2918_
	);
	LUT4 #(
		.INIT('h111d)
	) name2456 (
		\P2_reg0_reg[27]/NET0131 ,
		_w2272_,
		_w2392_,
		_w2393_,
		_w2919_
	);
	LUT4 #(
		.INIT('h0100)
	) name2457 (
		_w1491_,
		_w1493_,
		_w1496_,
		_w2084_,
		_w2920_
	);
	LUT3 #(
		.INIT('ha2)
	) name2458 (
		\P2_reg0_reg[27]/NET0131 ,
		_w2633_,
		_w2634_,
		_w2921_
	);
	LUT4 #(
		.INIT('h00ef)
	) name2459 (
		_w1509_,
		_w1970_,
		_w2920_,
		_w2921_,
		_w2922_
	);
	LUT3 #(
		.INIT('hd0)
	) name2460 (
		_w2081_,
		_w2919_,
		_w2922_,
		_w2923_
	);
	LUT4 #(
		.INIT('hab00)
	) name2461 (
		_w2192_,
		_w2915_,
		_w2918_,
		_w2923_,
		_w2924_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name2462 (
		_w1489_,
		_w2917_,
		_w2914_,
		_w2924_,
		_w2925_
	);
	LUT4 #(
		.INIT('heeec)
	) name2463 (
		\P1_state_reg[0]/NET0131 ,
		_w2911_,
		_w2912_,
		_w2925_,
		_w2926_
	);
	LUT4 #(
		.INIT('h70d0)
	) name2464 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg0_reg[28]/NET0131 ,
		_w1476_,
		_w2927_
	);
	LUT2 #(
		.INIT('h8)
	) name2465 (
		\P2_reg0_reg[28]/NET0131 ,
		_w1487_,
		_w2928_
	);
	LUT4 #(
		.INIT('haaa8)
	) name2466 (
		\P2_reg0_reg[28]/NET0131 ,
		_w1491_,
		_w1493_,
		_w1496_,
		_w2929_
	);
	LUT4 #(
		.INIT('h3c55)
	) name2467 (
		\P2_reg0_reg[28]/NET0131 ,
		_w2008_,
		_w2027_,
		_w2277_,
		_w2930_
	);
	LUT4 #(
		.INIT('h02aa)
	) name2468 (
		\P2_reg0_reg[28]/NET0131 ,
		_w1491_,
		_w1493_,
		_w1496_,
		_w2931_
	);
	LUT4 #(
		.INIT('hba00)
	) name2469 (
		_w2043_,
		_w2075_,
		_w2078_,
		_w2272_,
		_w2932_
	);
	LUT3 #(
		.INIT('ha2)
	) name2470 (
		\P2_reg0_reg[28]/NET0131 ,
		_w2633_,
		_w2634_,
		_w2933_
	);
	LUT4 #(
		.INIT('h00ef)
	) name2471 (
		_w1509_,
		_w2017_,
		_w2920_,
		_w2933_,
		_w2934_
	);
	LUT4 #(
		.INIT('h5700)
	) name2472 (
		_w2081_,
		_w2931_,
		_w2932_,
		_w2934_,
		_w2935_
	);
	LUT3 #(
		.INIT('he0)
	) name2473 (
		_w2276_,
		_w2930_,
		_w2935_,
		_w2936_
	);
	LUT4 #(
		.INIT('h9a00)
	) name2474 (
		_w2027_,
		_w2169_,
		_w2186_,
		_w2277_,
		_w2937_
	);
	LUT3 #(
		.INIT('h54)
	) name2475 (
		_w2192_,
		_w2929_,
		_w2937_,
		_w2938_
	);
	LUT4 #(
		.INIT('h3c55)
	) name2476 (
		\P2_reg0_reg[28]/NET0131 ,
		_w2008_,
		_w2027_,
		_w2272_,
		_w2939_
	);
	LUT2 #(
		.INIT('h2)
	) name2477 (
		_w2290_,
		_w2939_,
		_w2940_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name2478 (
		_w1489_,
		_w2938_,
		_w2940_,
		_w2936_,
		_w2941_
	);
	LUT4 #(
		.INIT('heeec)
	) name2479 (
		\P1_state_reg[0]/NET0131 ,
		_w2927_,
		_w2928_,
		_w2941_,
		_w2942_
	);
	LUT2 #(
		.INIT('h2)
	) name2480 (
		\P1_reg2_reg[24]/NET0131 ,
		_w511_,
		_w2943_
	);
	LUT2 #(
		.INIT('h8)
	) name2481 (
		\P1_reg2_reg[24]/NET0131 ,
		_w524_,
		_w2944_
	);
	LUT4 #(
		.INIT('h5455)
	) name2482 (
		\P1_reg2_reg[24]/NET0131 ,
		_w528_,
		_w530_,
		_w533_,
		_w2945_
	);
	LUT2 #(
		.INIT('h2)
	) name2483 (
		_w1286_,
		_w2945_,
		_w2946_
	);
	LUT4 #(
		.INIT('h7d00)
	) name2484 (
		_w534_,
		_w1425_,
		_w2767_,
		_w2946_,
		_w2947_
	);
	LUT3 #(
		.INIT('h10)
	) name2485 (
		_w541_,
		_w1054_,
		_w1138_,
		_w2948_
	);
	LUT4 #(
		.INIT('haa8a)
	) name2486 (
		_w534_,
		_w2775_,
		_w2781_,
		_w2948_,
		_w2949_
	);
	LUT2 #(
		.INIT('h8)
	) name2487 (
		_w1056_,
		_w1143_,
		_w2950_
	);
	LUT2 #(
		.INIT('h4)
	) name2488 (
		_w534_,
		_w1183_,
		_w2951_
	);
	LUT4 #(
		.INIT('haaa2)
	) name2489 (
		\P1_reg2_reg[24]/NET0131 ,
		_w2411_,
		_w2412_,
		_w2951_,
		_w2952_
	);
	LUT2 #(
		.INIT('h1)
	) name2490 (
		_w2950_,
		_w2952_,
		_w2953_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name2491 (
		_w526_,
		_w2949_,
		_w2947_,
		_w2953_,
		_w2954_
	);
	LUT4 #(
		.INIT('heeec)
	) name2492 (
		\P1_state_reg[0]/NET0131 ,
		_w2943_,
		_w2944_,
		_w2954_,
		_w2955_
	);
	LUT4 #(
		.INIT('h70d0)
	) name2493 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg1_reg[28]/NET0131 ,
		_w1476_,
		_w2956_
	);
	LUT2 #(
		.INIT('h8)
	) name2494 (
		\P2_reg1_reg[28]/NET0131 ,
		_w1487_,
		_w2957_
	);
	LUT4 #(
		.INIT('haa02)
	) name2495 (
		\P2_reg1_reg[28]/NET0131 ,
		_w1491_,
		_w1493_,
		_w1496_,
		_w2958_
	);
	LUT4 #(
		.INIT('h3c55)
	) name2496 (
		\P2_reg1_reg[28]/NET0131 ,
		_w2008_,
		_w2027_,
		_w2039_,
		_w2959_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name2497 (
		\P2_reg1_reg[28]/NET0131 ,
		_w1491_,
		_w1493_,
		_w1496_,
		_w2960_
	);
	LUT4 #(
		.INIT('h8a88)
	) name2498 (
		_w1497_,
		_w2043_,
		_w2075_,
		_w2078_,
		_w2961_
	);
	LUT3 #(
		.INIT('ha2)
	) name2499 (
		\P2_reg1_reg[28]/NET0131 ,
		_w2633_,
		_w2660_,
		_w2962_
	);
	LUT4 #(
		.INIT('h0e00)
	) name2500 (
		_w1491_,
		_w1493_,
		_w1496_,
		_w2084_,
		_w2963_
	);
	LUT4 #(
		.INIT('h0e0f)
	) name2501 (
		_w1509_,
		_w2017_,
		_w2962_,
		_w2963_,
		_w2964_
	);
	LUT4 #(
		.INIT('h5700)
	) name2502 (
		_w2081_,
		_w2960_,
		_w2961_,
		_w2964_,
		_w2965_
	);
	LUT3 #(
		.INIT('hd0)
	) name2503 (
		_w2038_,
		_w2959_,
		_w2965_,
		_w2966_
	);
	LUT3 #(
		.INIT('hc8)
	) name2504 (
		_w2187_,
		_w2193_,
		_w2958_,
		_w2967_
	);
	LUT3 #(
		.INIT('ha8)
	) name2505 (
		_w2188_,
		_w2190_,
		_w2960_,
		_w2968_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name2506 (
		_w1489_,
		_w2967_,
		_w2968_,
		_w2966_,
		_w2969_
	);
	LUT4 #(
		.INIT('heeec)
	) name2507 (
		\P1_state_reg[0]/NET0131 ,
		_w2956_,
		_w2957_,
		_w2969_,
		_w2970_
	);
	LUT4 #(
		.INIT('h70d0)
	) name2508 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg1_reg[27]/NET0131 ,
		_w1476_,
		_w2971_
	);
	LUT2 #(
		.INIT('h8)
	) name2509 (
		\P2_reg1_reg[27]/NET0131 ,
		_w1487_,
		_w2972_
	);
	LUT4 #(
		.INIT('haa02)
	) name2510 (
		\P2_reg1_reg[27]/NET0131 ,
		_w1491_,
		_w1493_,
		_w1496_,
		_w2973_
	);
	LUT4 #(
		.INIT('h1dd1)
	) name2511 (
		\P2_reg1_reg[27]/NET0131 ,
		_w2039_,
		_w2301_,
		_w2342_,
		_w2974_
	);
	LUT2 #(
		.INIT('h2)
	) name2512 (
		_w2038_,
		_w2974_,
		_w2975_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name2513 (
		\P2_reg1_reg[27]/NET0131 ,
		_w1491_,
		_w1493_,
		_w1496_,
		_w2976_
	);
	LUT3 #(
		.INIT('ha8)
	) name2514 (
		_w2188_,
		_w2391_,
		_w2976_,
		_w2977_
	);
	LUT4 #(
		.INIT('h111d)
	) name2515 (
		\P2_reg1_reg[27]/NET0131 ,
		_w1497_,
		_w2392_,
		_w2393_,
		_w2978_
	);
	LUT3 #(
		.INIT('ha2)
	) name2516 (
		\P2_reg1_reg[27]/NET0131 ,
		_w2633_,
		_w2660_,
		_w2979_
	);
	LUT4 #(
		.INIT('h00ef)
	) name2517 (
		_w1509_,
		_w1970_,
		_w2963_,
		_w2979_,
		_w2980_
	);
	LUT3 #(
		.INIT('hd0)
	) name2518 (
		_w2081_,
		_w2978_,
		_w2980_,
		_w2981_
	);
	LUT4 #(
		.INIT('h5700)
	) name2519 (
		_w2193_,
		_w2389_,
		_w2973_,
		_w2981_,
		_w2982_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name2520 (
		_w1489_,
		_w2975_,
		_w2977_,
		_w2982_,
		_w2983_
	);
	LUT4 #(
		.INIT('heeec)
	) name2521 (
		\P1_state_reg[0]/NET0131 ,
		_w2971_,
		_w2972_,
		_w2983_,
		_w2984_
	);
	LUT2 #(
		.INIT('h2)
	) name2522 (
		\P1_reg0_reg[28]/NET0131 ,
		_w511_,
		_w2985_
	);
	LUT4 #(
		.INIT('haaa8)
	) name2523 (
		\P1_reg0_reg[28]/NET0131 ,
		_w528_,
		_w530_,
		_w533_,
		_w2986_
	);
	LUT4 #(
		.INIT('h9a00)
	) name2524 (
		_w1419_,
		_w2201_,
		_w2203_,
		_w2688_,
		_w2987_
	);
	LUT3 #(
		.INIT('ha8)
	) name2525 (
		_w1286_,
		_w2986_,
		_w2987_,
		_w2988_
	);
	LUT4 #(
		.INIT('hfc55)
	) name2526 (
		\P1_reg0_reg[28]/NET0131 ,
		_w2206_,
		_w2207_,
		_w2688_,
		_w2989_
	);
	LUT4 #(
		.INIT('h2f00)
	) name2527 (
		_w1114_,
		_w2254_,
		_w2408_,
		_w2688_,
		_w2990_
	);
	LUT3 #(
		.INIT('h0e)
	) name2528 (
		_w1114_,
		_w1136_,
		_w2688_,
		_w2991_
	);
	LUT3 #(
		.INIT('ha2)
	) name2529 (
		\P1_reg0_reg[28]/NET0131 ,
		_w2692_,
		_w2991_,
		_w2992_
	);
	LUT4 #(
		.INIT('h000d)
	) name2530 (
		_w1183_,
		_w2989_,
		_w2990_,
		_w2992_,
		_w2993_
	);
	LUT2 #(
		.INIT('h8)
	) name2531 (
		\P1_reg0_reg[28]/NET0131 ,
		_w524_,
		_w2994_
	);
	LUT4 #(
		.INIT('h0075)
	) name2532 (
		_w526_,
		_w2988_,
		_w2993_,
		_w2994_,
		_w2995_
	);
	LUT3 #(
		.INIT('hce)
	) name2533 (
		\P1_state_reg[0]/NET0131 ,
		_w2985_,
		_w2995_,
		_w2996_
	);
	LUT2 #(
		.INIT('h2)
	) name2534 (
		\P1_reg0_reg[25]/NET0131 ,
		_w511_,
		_w2997_
	);
	LUT2 #(
		.INIT('h8)
	) name2535 (
		\P1_reg0_reg[25]/NET0131 ,
		_w524_,
		_w2998_
	);
	LUT4 #(
		.INIT('haaa8)
	) name2536 (
		\P1_reg0_reg[25]/NET0131 ,
		_w528_,
		_w530_,
		_w533_,
		_w2999_
	);
	LUT2 #(
		.INIT('h8)
	) name2537 (
		_w795_,
		_w953_,
		_w3000_
	);
	LUT3 #(
		.INIT('hd0)
	) name2538 (
		_w794_,
		_w846_,
		_w957_,
		_w3001_
	);
	LUT3 #(
		.INIT('hc4)
	) name2539 (
		_w748_,
		_w964_,
		_w3001_,
		_w3002_
	);
	LUT4 #(
		.INIT('h4c44)
	) name2540 (
		_w1082_,
		_w1091_,
		_w3000_,
		_w3002_,
		_w3003_
	);
	LUT4 #(
		.INIT('h35c5)
	) name2541 (
		\P1_reg0_reg[25]/NET0131 ,
		_w1420_,
		_w2688_,
		_w3003_,
		_w3004_
	);
	LUT3 #(
		.INIT('h08)
	) name2542 (
		_w1107_,
		_w1140_,
		_w2688_,
		_w3005_
	);
	LUT3 #(
		.INIT('ha2)
	) name2543 (
		\P1_reg0_reg[25]/NET0131 ,
		_w2692_,
		_w3005_,
		_w3006_
	);
	LUT3 #(
		.INIT('h10)
	) name2544 (
		_w541_,
		_w968_,
		_w1138_,
		_w3007_
	);
	LUT4 #(
		.INIT('h6500)
	) name2545 (
		_w969_,
		_w1055_,
		_w1128_,
		_w1136_,
		_w3008_
	);
	LUT4 #(
		.INIT('h1113)
	) name2546 (
		_w2688_,
		_w3006_,
		_w3007_,
		_w3008_,
		_w3009_
	);
	LUT3 #(
		.INIT('hd0)
	) name2547 (
		_w1114_,
		_w3004_,
		_w3009_,
		_w3010_
	);
	LUT4 #(
		.INIT('h9555)
	) name2548 (
		_w1004_,
		_w1161_,
		_w1163_,
		_w1171_,
		_w3011_
	);
	LUT4 #(
		.INIT('h7020)
	) name2549 (
		_w537_,
		_w1059_,
		_w2688_,
		_w3011_,
		_w3012_
	);
	LUT3 #(
		.INIT('ha8)
	) name2550 (
		_w1183_,
		_w2999_,
		_w3012_,
		_w3013_
	);
	LUT2 #(
		.INIT('h8)
	) name2551 (
		_w1194_,
		_w1237_,
		_w3014_
	);
	LUT3 #(
		.INIT('hd0)
	) name2552 (
		_w1193_,
		_w1202_,
		_w1243_,
		_w3015_
	);
	LUT3 #(
		.INIT('hc4)
	) name2553 (
		_w1190_,
		_w1250_,
		_w3015_,
		_w3016_
	);
	LUT4 #(
		.INIT('h4c44)
	) name2554 (
		_w1257_,
		_w1273_,
		_w3014_,
		_w3016_,
		_w3017_
	);
	LUT4 #(
		.INIT('hc535)
	) name2555 (
		\P1_reg0_reg[25]/NET0131 ,
		_w1420_,
		_w2688_,
		_w3017_,
		_w3018_
	);
	LUT3 #(
		.INIT('h31)
	) name2556 (
		_w1286_,
		_w3013_,
		_w3018_,
		_w3019_
	);
	LUT4 #(
		.INIT('h3111)
	) name2557 (
		_w526_,
		_w2998_,
		_w3010_,
		_w3019_,
		_w3020_
	);
	LUT3 #(
		.INIT('hce)
	) name2558 (
		\P1_state_reg[0]/NET0131 ,
		_w2997_,
		_w3020_,
		_w3021_
	);
	LUT2 #(
		.INIT('h2)
	) name2559 (
		\P1_reg1_reg[25]/NET0131 ,
		_w511_,
		_w3022_
	);
	LUT2 #(
		.INIT('h8)
	) name2560 (
		\P1_reg1_reg[25]/NET0131 ,
		_w524_,
		_w3023_
	);
	LUT4 #(
		.INIT('haa02)
	) name2561 (
		\P1_reg1_reg[25]/NET0131 ,
		_w528_,
		_w530_,
		_w533_,
		_w3024_
	);
	LUT4 #(
		.INIT('h35c5)
	) name2562 (
		\P1_reg1_reg[25]/NET0131 ,
		_w1420_,
		_w2421_,
		_w3003_,
		_w3025_
	);
	LUT4 #(
		.INIT('hf100)
	) name2563 (
		_w1136_,
		_w1138_,
		_w2421_,
		_w2425_,
		_w3026_
	);
	LUT2 #(
		.INIT('h2)
	) name2564 (
		\P1_reg1_reg[25]/NET0131 ,
		_w3026_,
		_w3027_
	);
	LUT4 #(
		.INIT('h0057)
	) name2565 (
		_w2421_,
		_w3007_,
		_w3008_,
		_w3027_,
		_w3028_
	);
	LUT3 #(
		.INIT('hd0)
	) name2566 (
		_w1114_,
		_w3025_,
		_w3028_,
		_w3029_
	);
	LUT4 #(
		.INIT('h7020)
	) name2567 (
		_w537_,
		_w1059_,
		_w2421_,
		_w3011_,
		_w3030_
	);
	LUT3 #(
		.INIT('ha8)
	) name2568 (
		_w1183_,
		_w3024_,
		_w3030_,
		_w3031_
	);
	LUT4 #(
		.INIT('hc535)
	) name2569 (
		\P1_reg1_reg[25]/NET0131 ,
		_w1420_,
		_w2421_,
		_w3017_,
		_w3032_
	);
	LUT3 #(
		.INIT('h31)
	) name2570 (
		_w1286_,
		_w3031_,
		_w3032_,
		_w3033_
	);
	LUT4 #(
		.INIT('h3111)
	) name2571 (
		_w526_,
		_w3023_,
		_w3029_,
		_w3033_,
		_w3034_
	);
	LUT3 #(
		.INIT('hce)
	) name2572 (
		\P1_state_reg[0]/NET0131 ,
		_w3022_,
		_w3034_,
		_w3035_
	);
	LUT2 #(
		.INIT('h2)
	) name2573 (
		\P1_reg1_reg[26]/NET0131 ,
		_w511_,
		_w3036_
	);
	LUT2 #(
		.INIT('h8)
	) name2574 (
		\P1_reg1_reg[26]/NET0131 ,
		_w524_,
		_w3037_
	);
	LUT4 #(
		.INIT('h4150)
	) name2575 (
		_w537_,
		_w1004_,
		_w1040_,
		_w1172_,
		_w3038_
	);
	LUT4 #(
		.INIT('hdf00)
	) name2576 (
		_w537_,
		_w973_,
		_w976_,
		_w1183_,
		_w3039_
	);
	LUT2 #(
		.INIT('h4)
	) name2577 (
		_w3038_,
		_w3039_,
		_w3040_
	);
	LUT3 #(
		.INIT('h10)
	) name2578 (
		_w979_,
		_w1061_,
		_w2243_,
		_w3041_
	);
	LUT3 #(
		.INIT('hb0)
	) name2579 (
		_w2237_,
		_w2244_,
		_w2247_,
		_w3042_
	);
	LUT2 #(
		.INIT('h8)
	) name2580 (
		_w2209_,
		_w2244_,
		_w3043_
	);
	LUT2 #(
		.INIT('h8)
	) name2581 (
		_w2210_,
		_w2212_,
		_w3044_
	);
	LUT3 #(
		.INIT('hd0)
	) name2582 (
		_w2213_,
		_w2218_,
		_w2232_,
		_w3045_
	);
	LUT3 #(
		.INIT('h0d)
	) name2583 (
		_w2210_,
		_w2233_,
		_w2235_,
		_w3046_
	);
	LUT3 #(
		.INIT('hd0)
	) name2584 (
		_w3044_,
		_w3045_,
		_w3046_,
		_w3047_
	);
	LUT4 #(
		.INIT('h22a2)
	) name2585 (
		_w3041_,
		_w3042_,
		_w3043_,
		_w3047_,
		_w3048_
	);
	LUT4 #(
		.INIT('h80f0)
	) name2586 (
		_w871_,
		_w883_,
		_w2222_,
		_w2220_,
		_w3049_
	);
	LUT4 #(
		.INIT('h0001)
	) name2587 (
		_w908_,
		_w919_,
		_w930_,
		_w950_,
		_w3050_
	);
	LUT3 #(
		.INIT('h8a)
	) name2588 (
		_w2217_,
		_w2226_,
		_w2228_,
		_w3051_
	);
	LUT4 #(
		.INIT('h2f00)
	) name2589 (
		_w2225_,
		_w3049_,
		_w3050_,
		_w3051_,
		_w3052_
	);
	LUT2 #(
		.INIT('h8)
	) name2590 (
		_w2213_,
		_w2216_,
		_w3053_
	);
	LUT3 #(
		.INIT('h80)
	) name2591 (
		_w2209_,
		_w2244_,
		_w3044_,
		_w3054_
	);
	LUT4 #(
		.INIT('h2000)
	) name2592 (
		_w3041_,
		_w3052_,
		_w3053_,
		_w3054_,
		_w3055_
	);
	LUT3 #(
		.INIT('h01)
	) name2593 (
		_w979_,
		_w1061_,
		_w2248_,
		_w3056_
	);
	LUT2 #(
		.INIT('h2)
	) name2594 (
		_w2250_,
		_w3056_,
		_w3057_
	);
	LUT4 #(
		.INIT('ha9aa)
	) name2595 (
		_w1432_,
		_w3048_,
		_w3055_,
		_w3057_,
		_w3058_
	);
	LUT4 #(
		.INIT('h9500)
	) name2596 (
		_w998_,
		_w1128_,
		_w1129_,
		_w1136_,
		_w3059_
	);
	LUT2 #(
		.INIT('h8)
	) name2597 (
		_w998_,
		_w1138_,
		_w3060_
	);
	LUT2 #(
		.INIT('h1)
	) name2598 (
		_w3059_,
		_w3060_,
		_w3061_
	);
	LUT3 #(
		.INIT('hd0)
	) name2599 (
		_w1114_,
		_w3058_,
		_w3061_,
		_w3062_
	);
	LUT3 #(
		.INIT('h8a)
	) name2600 (
		_w2421_,
		_w3040_,
		_w3062_,
		_w3063_
	);
	LUT4 #(
		.INIT('h82c3)
	) name2601 (
		_w652_,
		_w1104_,
		_w1106_,
		_w1111_,
		_w3064_
	);
	LUT2 #(
		.INIT('h1)
	) name2602 (
		_w2421_,
		_w3064_,
		_w3065_
	);
	LUT3 #(
		.INIT('h02)
	) name2603 (
		_w1113_,
		_w2421_,
		_w3064_,
		_w3066_
	);
	LUT3 #(
		.INIT('ha2)
	) name2604 (
		\P1_reg1_reg[26]/NET0131 ,
		_w2426_,
		_w3066_,
		_w3067_
	);
	LUT3 #(
		.INIT('h10)
	) name2605 (
		_w1256_,
		_w1262_,
		_w1323_,
		_w3068_
	);
	LUT3 #(
		.INIT('h15)
	) name2606 (
		_w1324_,
		_w1332_,
		_w1334_,
		_w3069_
	);
	LUT2 #(
		.INIT('h8)
	) name2607 (
		_w1328_,
		_w1334_,
		_w3070_
	);
	LUT2 #(
		.INIT('h8)
	) name2608 (
		_w1339_,
		_w1342_,
		_w3071_
	);
	LUT3 #(
		.INIT('h80)
	) name2609 (
		_w1328_,
		_w1334_,
		_w3071_,
		_w3072_
	);
	LUT4 #(
		.INIT('hf200)
	) name2610 (
		_w1214_,
		_w1360_,
		_w1361_,
		_w1363_,
		_w3073_
	);
	LUT4 #(
		.INIT('h0001)
	) name2611 (
		_w1203_,
		_w1204_,
		_w1221_,
		_w1234_,
		_w3074_
	);
	LUT3 #(
		.INIT('h15)
	) name2612 (
		_w1355_,
		_w1367_,
		_w1347_,
		_w3075_
	);
	LUT4 #(
		.INIT('h2f00)
	) name2613 (
		_w1366_,
		_w3073_,
		_w3074_,
		_w3075_,
		_w3076_
	);
	LUT2 #(
		.INIT('h8)
	) name2614 (
		_w1350_,
		_w1346_,
		_w3077_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name2615 (
		_w3069_,
		_w3072_,
		_w3076_,
		_w3077_,
		_w3078_
	);
	LUT3 #(
		.INIT('h15)
	) name2616 (
		_w1343_,
		_w1350_,
		_w1357_,
		_w3079_
	);
	LUT3 #(
		.INIT('h15)
	) name2617 (
		_w1330_,
		_w1339_,
		_w1344_,
		_w3080_
	);
	LUT3 #(
		.INIT('hd0)
	) name2618 (
		_w3071_,
		_w3079_,
		_w3080_,
		_w3081_
	);
	LUT3 #(
		.INIT('h08)
	) name2619 (
		_w3068_,
		_w3070_,
		_w3081_,
		_w3082_
	);
	LUT3 #(
		.INIT('h10)
	) name2620 (
		_w1256_,
		_w1262_,
		_w1326_,
		_w3083_
	);
	LUT2 #(
		.INIT('h1)
	) name2621 (
		_w1318_,
		_w3083_,
		_w3084_
	);
	LUT4 #(
		.INIT('h0d00)
	) name2622 (
		_w3068_,
		_w3078_,
		_w3082_,
		_w3084_,
		_w3085_
	);
	LUT4 #(
		.INIT('h5501)
	) name2623 (
		\P1_reg1_reg[26]/NET0131 ,
		_w528_,
		_w530_,
		_w533_,
		_w3086_
	);
	LUT2 #(
		.INIT('h2)
	) name2624 (
		_w1286_,
		_w3086_,
		_w3087_
	);
	LUT4 #(
		.INIT('h7b00)
	) name2625 (
		_w1432_,
		_w2421_,
		_w3085_,
		_w3087_,
		_w3088_
	);
	LUT2 #(
		.INIT('h1)
	) name2626 (
		_w3067_,
		_w3088_,
		_w3089_
	);
	LUT4 #(
		.INIT('h1311)
	) name2627 (
		_w526_,
		_w3037_,
		_w3063_,
		_w3089_,
		_w3090_
	);
	LUT3 #(
		.INIT('hce)
	) name2628 (
		\P1_state_reg[0]/NET0131 ,
		_w3036_,
		_w3090_,
		_w3091_
	);
	LUT2 #(
		.INIT('h2)
	) name2629 (
		\P1_reg1_reg[28]/NET0131 ,
		_w511_,
		_w3092_
	);
	LUT4 #(
		.INIT('haa02)
	) name2630 (
		\P1_reg1_reg[28]/NET0131 ,
		_w528_,
		_w530_,
		_w533_,
		_w3093_
	);
	LUT4 #(
		.INIT('h9a00)
	) name2631 (
		_w1419_,
		_w2201_,
		_w2203_,
		_w2421_,
		_w3094_
	);
	LUT3 #(
		.INIT('ha8)
	) name2632 (
		_w1286_,
		_w3093_,
		_w3094_,
		_w3095_
	);
	LUT4 #(
		.INIT('hfc55)
	) name2633 (
		\P1_reg1_reg[28]/NET0131 ,
		_w2206_,
		_w2207_,
		_w2421_,
		_w3096_
	);
	LUT4 #(
		.INIT('h2f00)
	) name2634 (
		_w1114_,
		_w2254_,
		_w2408_,
		_w2421_,
		_w3097_
	);
	LUT3 #(
		.INIT('h0e)
	) name2635 (
		_w1114_,
		_w1136_,
		_w2421_,
		_w3098_
	);
	LUT3 #(
		.INIT('ha2)
	) name2636 (
		\P1_reg1_reg[28]/NET0131 ,
		_w2426_,
		_w3098_,
		_w3099_
	);
	LUT4 #(
		.INIT('h000d)
	) name2637 (
		_w1183_,
		_w3096_,
		_w3097_,
		_w3099_,
		_w3100_
	);
	LUT2 #(
		.INIT('h8)
	) name2638 (
		\P1_reg1_reg[28]/NET0131 ,
		_w524_,
		_w3101_
	);
	LUT4 #(
		.INIT('h0075)
	) name2639 (
		_w526_,
		_w3095_,
		_w3100_,
		_w3101_,
		_w3102_
	);
	LUT3 #(
		.INIT('hce)
	) name2640 (
		\P1_state_reg[0]/NET0131 ,
		_w3092_,
		_w3102_,
		_w3103_
	);
	LUT2 #(
		.INIT('h8)
	) name2641 (
		_w524_,
		_w787_,
		_w3104_
	);
	LUT4 #(
		.INIT('h1f00)
	) name2642 (
		_w528_,
		_w530_,
		_w533_,
		_w787_,
		_w3105_
	);
	LUT4 #(
		.INIT('h0100)
	) name2643 (
		_w762_,
		_w772_,
		_w791_,
		_w1161_,
		_w3106_
	);
	LUT4 #(
		.INIT('h5054)
	) name2644 (
		_w537_,
		_w722_,
		_w1164_,
		_w3106_,
		_w3107_
	);
	LUT3 #(
		.INIT('h80)
	) name2645 (
		_w537_,
		_w769_,
		_w771_,
		_w3108_
	);
	LUT4 #(
		.INIT('h3331)
	) name2646 (
		_w2197_,
		_w3105_,
		_w3107_,
		_w3108_,
		_w3109_
	);
	LUT4 #(
		.INIT('h5100)
	) name2647 (
		_w1429_,
		_w2214_,
		_w2231_,
		_w2234_,
		_w3110_
	);
	LUT4 #(
		.INIT('h08aa)
	) name2648 (
		_w1429_,
		_w2214_,
		_w2231_,
		_w2234_,
		_w3111_
	);
	LUT3 #(
		.INIT('h02)
	) name2649 (
		_w1114_,
		_w3111_,
		_w3110_,
		_w3112_
	);
	LUT4 #(
		.INIT('ha200)
	) name2650 (
		_w1345_,
		_w1353_,
		_w1387_,
		_w1429_,
		_w3113_
	);
	LUT4 #(
		.INIT('h005d)
	) name2651 (
		_w1345_,
		_w1353_,
		_w1387_,
		_w1429_,
		_w3114_
	);
	LUT3 #(
		.INIT('h02)
	) name2652 (
		_w1286_,
		_w3114_,
		_w3113_,
		_w3115_
	);
	LUT3 #(
		.INIT('h80)
	) name2653 (
		_w786_,
		_w1120_,
		_w1122_,
		_w3116_
	);
	LUT4 #(
		.INIT('h6a00)
	) name2654 (
		_w786_,
		_w1120_,
		_w1122_,
		_w2197_,
		_w3117_
	);
	LUT3 #(
		.INIT('h98)
	) name2655 (
		_w1104_,
		_w1106_,
		_w1111_,
		_w3118_
	);
	LUT4 #(
		.INIT('h888a)
	) name2656 (
		_w787_,
		_w1141_,
		_w2197_,
		_w3118_,
		_w3119_
	);
	LUT3 #(
		.INIT('h04)
	) name2657 (
		_w786_,
		_w2259_,
		_w2260_,
		_w3120_
	);
	LUT2 #(
		.INIT('h1)
	) name2658 (
		_w3119_,
		_w3120_,
		_w3121_
	);
	LUT4 #(
		.INIT('h5700)
	) name2659 (
		_w1136_,
		_w3105_,
		_w3117_,
		_w3121_,
		_w3122_
	);
	LUT4 #(
		.INIT('h5700)
	) name2660 (
		_w2197_,
		_w3112_,
		_w3115_,
		_w3122_,
		_w3123_
	);
	LUT4 #(
		.INIT('h08aa)
	) name2661 (
		_w526_,
		_w1183_,
		_w3109_,
		_w3123_,
		_w3124_
	);
	LUT2 #(
		.INIT('h2)
	) name2662 (
		\P1_reg3_reg[16]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w3125_
	);
	LUT4 #(
		.INIT('h9d5d)
	) name2663 (
		\P1_reg3_reg[16]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w510_,
		_w718_,
		_w3126_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name2664 (
		\P1_state_reg[0]/NET0131 ,
		_w3104_,
		_w3124_,
		_w3126_,
		_w3127_
	);
	LUT2 #(
		.INIT('h8)
	) name2665 (
		_w524_,
		_w703_,
		_w3128_
	);
	LUT4 #(
		.INIT('ha028)
	) name2666 (
		_w1286_,
		_w1333_,
		_w1421_,
		_w2199_,
		_w3129_
	);
	LUT4 #(
		.INIT('h8000)
	) name2667 (
		_w786_,
		_w1120_,
		_w1122_,
		_w1123_,
		_w3130_
	);
	LUT4 #(
		.INIT('h7f00)
	) name2668 (
		_w1120_,
		_w1122_,
		_w1125_,
		_w1136_,
		_w3131_
	);
	LUT4 #(
		.INIT('h7300)
	) name2669 (
		_w674_,
		_w702_,
		_w3130_,
		_w3131_,
		_w3132_
	);
	LUT4 #(
		.INIT('h007d)
	) name2670 (
		_w1114_,
		_w1421_,
		_w2240_,
		_w3132_,
		_w3133_
	);
	LUT3 #(
		.INIT('h8a)
	) name2671 (
		_w2197_,
		_w3129_,
		_w3133_,
		_w3134_
	);
	LUT4 #(
		.INIT('h4000)
	) name2672 (
		_w706_,
		_w1165_,
		_w1161_,
		_w1163_,
		_w3135_
	);
	LUT4 #(
		.INIT('h8000)
	) name2673 (
		_w1166_,
		_w1165_,
		_w1161_,
		_w1163_,
		_w3136_
	);
	LUT4 #(
		.INIT('h5504)
	) name2674 (
		_w537_,
		_w1078_,
		_w3135_,
		_w3136_,
		_w3137_
	);
	LUT4 #(
		.INIT('h0200)
	) name2675 (
		_w537_,
		_w677_,
		_w676_,
		_w678_,
		_w3138_
	);
	LUT4 #(
		.INIT('h001f)
	) name2676 (
		_w528_,
		_w530_,
		_w533_,
		_w703_,
		_w3139_
	);
	LUT2 #(
		.INIT('h2)
	) name2677 (
		_w1183_,
		_w3139_,
		_w3140_
	);
	LUT4 #(
		.INIT('h5700)
	) name2678 (
		_w2197_,
		_w3137_,
		_w3138_,
		_w3140_,
		_w3141_
	);
	LUT4 #(
		.INIT('hc2c3)
	) name2679 (
		_w652_,
		_w1104_,
		_w1106_,
		_w1111_,
		_w3142_
	);
	LUT4 #(
		.INIT('h3130)
	) name2680 (
		_w1138_,
		_w1141_,
		_w2197_,
		_w3142_,
		_w3143_
	);
	LUT4 #(
		.INIT('h0010)
	) name2681 (
		_w541_,
		_w701_,
		_w2259_,
		_w2260_,
		_w3144_
	);
	LUT3 #(
		.INIT('h0d)
	) name2682 (
		_w703_,
		_w3143_,
		_w3144_,
		_w3145_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name2683 (
		_w526_,
		_w3141_,
		_w3134_,
		_w3145_,
		_w3146_
	);
	LUT2 #(
		.INIT('h2)
	) name2684 (
		\P1_reg3_reg[20]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w3147_
	);
	LUT4 #(
		.INIT('h6c00)
	) name2685 (
		\P1_reg3_reg[19]/NET0131 ,
		\P1_reg3_reg[20]/NET0131 ,
		_w634_,
		_w1294_,
		_w3148_
	);
	LUT2 #(
		.INIT('h1)
	) name2686 (
		_w3147_,
		_w3148_,
		_w3149_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name2687 (
		\P1_state_reg[0]/NET0131 ,
		_w3128_,
		_w3146_,
		_w3149_,
		_w3150_
	);
	LUT4 #(
		.INIT('h70d0)
	) name2688 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg2_reg[18]/NET0131 ,
		_w1476_,
		_w3151_
	);
	LUT2 #(
		.INIT('h8)
	) name2689 (
		\P2_reg2_reg[18]/NET0131 ,
		_w1487_,
		_w3152_
	);
	LUT4 #(
		.INIT('haa02)
	) name2690 (
		\P2_reg2_reg[18]/NET0131 ,
		_w1491_,
		_w1493_,
		_w1496_,
		_w3153_
	);
	LUT4 #(
		.INIT('h8a20)
	) name2691 (
		_w2039_,
		_w2495_,
		_w2498_,
		_w2728_,
		_w3154_
	);
	LUT3 #(
		.INIT('ha8)
	) name2692 (
		_w2188_,
		_w3153_,
		_w3154_,
		_w3155_
	);
	LUT4 #(
		.INIT('h20e0)
	) name2693 (
		\P2_reg2_reg[18]/NET0131 ,
		_w2039_,
		_w2081_,
		_w2732_,
		_w3156_
	);
	LUT3 #(
		.INIT('ha8)
	) name2694 (
		\P2_reg2_reg[18]/NET0131 ,
		_w2086_,
		_w2087_,
		_w3157_
	);
	LUT2 #(
		.INIT('h4)
	) name2695 (
		_w1834_,
		_w2088_,
		_w3158_
	);
	LUT3 #(
		.INIT('h0b)
	) name2696 (
		_w1833_,
		_w2085_,
		_w3158_,
		_w3159_
	);
	LUT2 #(
		.INIT('h4)
	) name2697 (
		_w3157_,
		_w3159_,
		_w3160_
	);
	LUT2 #(
		.INIT('h4)
	) name2698 (
		_w3156_,
		_w3160_,
		_w3161_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name2699 (
		\P2_reg2_reg[18]/NET0131 ,
		_w1491_,
		_w1493_,
		_w1496_,
		_w3162_
	);
	LUT4 #(
		.INIT('h8a20)
	) name2700 (
		_w1497_,
		_w2495_,
		_w2498_,
		_w2728_,
		_w3163_
	);
	LUT3 #(
		.INIT('ha8)
	) name2701 (
		_w2193_,
		_w3162_,
		_w3163_,
		_w3164_
	);
	LUT4 #(
		.INIT('h1dd1)
	) name2702 (
		\P2_reg2_reg[18]/NET0131 ,
		_w1497_,
		_w2472_,
		_w2728_,
		_w3165_
	);
	LUT2 #(
		.INIT('h2)
	) name2703 (
		_w2038_,
		_w3165_,
		_w3166_
	);
	LUT4 #(
		.INIT('h0100)
	) name2704 (
		_w3155_,
		_w3164_,
		_w3166_,
		_w3161_,
		_w3167_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name2705 (
		\P1_state_reg[0]/NET0131 ,
		_w1489_,
		_w3152_,
		_w3167_,
		_w3168_
	);
	LUT2 #(
		.INIT('he)
	) name2706 (
		_w3151_,
		_w3168_,
		_w3169_
	);
	LUT4 #(
		.INIT('h70d0)
	) name2707 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg2_reg[19]/NET0131 ,
		_w1476_,
		_w3170_
	);
	LUT2 #(
		.INIT('h8)
	) name2708 (
		\P2_reg2_reg[19]/NET0131 ,
		_w1487_,
		_w3171_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name2709 (
		\P2_reg2_reg[19]/NET0131 ,
		_w1491_,
		_w1493_,
		_w1496_,
		_w3172_
	);
	LUT4 #(
		.INIT('h208a)
	) name2710 (
		_w1497_,
		_w2319_,
		_w2327_,
		_w2749_,
		_w3173_
	);
	LUT3 #(
		.INIT('ha8)
	) name2711 (
		_w2038_,
		_w3172_,
		_w3173_,
		_w3174_
	);
	LUT4 #(
		.INIT('h20e0)
	) name2712 (
		\P2_reg2_reg[19]/NET0131 ,
		_w2039_,
		_w2081_,
		_w2756_,
		_w3175_
	);
	LUT4 #(
		.INIT('hd11d)
	) name2713 (
		\P2_reg2_reg[19]/NET0131 ,
		_w1497_,
		_w2378_,
		_w2749_,
		_w3176_
	);
	LUT2 #(
		.INIT('h2)
	) name2714 (
		_w2193_,
		_w3176_,
		_w3177_
	);
	LUT4 #(
		.INIT('hd11d)
	) name2715 (
		\P2_reg2_reg[19]/NET0131 ,
		_w2039_,
		_w2378_,
		_w2749_,
		_w3178_
	);
	LUT3 #(
		.INIT('ha8)
	) name2716 (
		\P2_reg2_reg[19]/NET0131 ,
		_w2086_,
		_w2087_,
		_w3179_
	);
	LUT2 #(
		.INIT('h4)
	) name2717 (
		_w1815_,
		_w2088_,
		_w3180_
	);
	LUT3 #(
		.INIT('h0b)
	) name2718 (
		_w1813_,
		_w2085_,
		_w3180_,
		_w3181_
	);
	LUT2 #(
		.INIT('h4)
	) name2719 (
		_w3179_,
		_w3181_,
		_w3182_
	);
	LUT3 #(
		.INIT('hd0)
	) name2720 (
		_w2188_,
		_w3178_,
		_w3182_,
		_w3183_
	);
	LUT4 #(
		.INIT('h0100)
	) name2721 (
		_w3174_,
		_w3175_,
		_w3177_,
		_w3183_,
		_w3184_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name2722 (
		\P1_state_reg[0]/NET0131 ,
		_w1489_,
		_w3171_,
		_w3184_,
		_w3185_
	);
	LUT2 #(
		.INIT('he)
	) name2723 (
		_w3170_,
		_w3185_,
		_w3186_
	);
	LUT4 #(
		.INIT('h70d0)
	) name2724 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg2_reg[20]/NET0131 ,
		_w1476_,
		_w3187_
	);
	LUT2 #(
		.INIT('h8)
	) name2725 (
		\P2_reg2_reg[20]/NET0131 ,
		_w1487_,
		_w3188_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name2726 (
		\P2_reg2_reg[20]/NET0131 ,
		_w1491_,
		_w1493_,
		_w1496_,
		_w3189_
	);
	LUT4 #(
		.INIT('h54ab)
	) name2727 (
		_w1509_,
		_w1858_,
		_w1865_,
		_w1872_,
		_w3190_
	);
	LUT4 #(
		.INIT('h1dd1)
	) name2728 (
		\P2_reg2_reg[20]/NET0131 ,
		_w1497_,
		_w1857_,
		_w3190_,
		_w3191_
	);
	LUT2 #(
		.INIT('h2)
	) name2729 (
		_w2038_,
		_w3191_,
		_w3192_
	);
	LUT4 #(
		.INIT('haa02)
	) name2730 (
		\P2_reg2_reg[20]/NET0131 ,
		_w1491_,
		_w1493_,
		_w1496_,
		_w3193_
	);
	LUT4 #(
		.INIT('hef00)
	) name2731 (
		_w1817_,
		_w1816_,
		_w1818_,
		_w2042_,
		_w3194_
	);
	LUT4 #(
		.INIT('h0603)
	) name2732 (
		_w1872_,
		_w1889_,
		_w2042_,
		_w2730_,
		_w3195_
	);
	LUT4 #(
		.INIT('h111d)
	) name2733 (
		\P2_reg2_reg[20]/NET0131 ,
		_w2039_,
		_w3194_,
		_w3195_,
		_w3196_
	);
	LUT4 #(
		.INIT('h5400)
	) name2734 (
		_w1509_,
		_w1858_,
		_w1865_,
		_w2085_,
		_w3197_
	);
	LUT2 #(
		.INIT('h4)
	) name2735 (
		_w1869_,
		_w2088_,
		_w3198_
	);
	LUT4 #(
		.INIT('h0057)
	) name2736 (
		\P2_reg2_reg[20]/NET0131 ,
		_w2086_,
		_w2087_,
		_w3198_,
		_w3199_
	);
	LUT2 #(
		.INIT('h4)
	) name2737 (
		_w3197_,
		_w3199_,
		_w3200_
	);
	LUT3 #(
		.INIT('hd0)
	) name2738 (
		_w2081_,
		_w3196_,
		_w3200_,
		_w3201_
	);
	LUT4 #(
		.INIT('h8a20)
	) name2739 (
		_w2039_,
		_w2138_,
		_w2155_,
		_w3190_,
		_w3202_
	);
	LUT3 #(
		.INIT('ha8)
	) name2740 (
		_w2188_,
		_w3193_,
		_w3202_,
		_w3203_
	);
	LUT4 #(
		.INIT('h8a20)
	) name2741 (
		_w1497_,
		_w2138_,
		_w2155_,
		_w3190_,
		_w3204_
	);
	LUT3 #(
		.INIT('ha8)
	) name2742 (
		_w2193_,
		_w3189_,
		_w3204_,
		_w3205_
	);
	LUT4 #(
		.INIT('h0100)
	) name2743 (
		_w3192_,
		_w3203_,
		_w3205_,
		_w3201_,
		_w3206_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name2744 (
		\P1_state_reg[0]/NET0131 ,
		_w1489_,
		_w3188_,
		_w3206_,
		_w3207_
	);
	LUT2 #(
		.INIT('he)
	) name2745 (
		_w3187_,
		_w3207_,
		_w3208_
	);
	LUT4 #(
		.INIT('h70d0)
	) name2746 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg2_reg[21]/NET0131 ,
		_w1476_,
		_w3209_
	);
	LUT2 #(
		.INIT('h8)
	) name2747 (
		\P2_reg2_reg[21]/NET0131 ,
		_w1487_,
		_w3210_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name2748 (
		\P2_reg2_reg[21]/NET0131 ,
		_w1491_,
		_w1493_,
		_w1496_,
		_w3211_
	);
	LUT3 #(
		.INIT('h1e)
	) name2749 (
		_w1509_,
		_w1882_,
		_w1889_,
		_w3212_
	);
	LUT4 #(
		.INIT('h8a20)
	) name2750 (
		_w1497_,
		_w2621_,
		_w2623_,
		_w3212_,
		_w3213_
	);
	LUT3 #(
		.INIT('ha8)
	) name2751 (
		_w2193_,
		_w3211_,
		_w3213_,
		_w3214_
	);
	LUT4 #(
		.INIT('haa02)
	) name2752 (
		\P2_reg2_reg[21]/NET0131 ,
		_w1491_,
		_w1493_,
		_w1496_,
		_w3215_
	);
	LUT4 #(
		.INIT('h8a20)
	) name2753 (
		_w2039_,
		_w2621_,
		_w2623_,
		_w3212_,
		_w3216_
	);
	LUT4 #(
		.INIT('h0200)
	) name2754 (
		_w1497_,
		_w1509_,
		_w1882_,
		_w2084_,
		_w3217_
	);
	LUT2 #(
		.INIT('h4)
	) name2755 (
		_w1885_,
		_w2088_,
		_w3218_
	);
	LUT4 #(
		.INIT('h0057)
	) name2756 (
		\P2_reg2_reg[21]/NET0131 ,
		_w2086_,
		_w2087_,
		_w3218_,
		_w3219_
	);
	LUT2 #(
		.INIT('h4)
	) name2757 (
		_w3217_,
		_w3219_,
		_w3220_
	);
	LUT4 #(
		.INIT('h5700)
	) name2758 (
		_w2188_,
		_w3215_,
		_w3216_,
		_w3220_,
		_w3221_
	);
	LUT2 #(
		.INIT('h4)
	) name2759 (
		_w1872_,
		_w2042_,
		_w3222_
	);
	LUT4 #(
		.INIT('h2111)
	) name2760 (
		_w1921_,
		_w2042_,
		_w2070_,
		_w2730_,
		_w3223_
	);
	LUT4 #(
		.INIT('h111d)
	) name2761 (
		\P2_reg2_reg[21]/NET0131 ,
		_w2039_,
		_w3222_,
		_w3223_,
		_w3224_
	);
	LUT2 #(
		.INIT('h2)
	) name2762 (
		_w2081_,
		_w3224_,
		_w3225_
	);
	LUT4 #(
		.INIT('h208a)
	) name2763 (
		_w1497_,
		_w2640_,
		_w2642_,
		_w3212_,
		_w3226_
	);
	LUT3 #(
		.INIT('ha8)
	) name2764 (
		_w2038_,
		_w3211_,
		_w3226_,
		_w3227_
	);
	LUT4 #(
		.INIT('h0100)
	) name2765 (
		_w3225_,
		_w3214_,
		_w3227_,
		_w3221_,
		_w3228_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name2766 (
		\P1_state_reg[0]/NET0131 ,
		_w1489_,
		_w3210_,
		_w3228_,
		_w3229_
	);
	LUT2 #(
		.INIT('he)
	) name2767 (
		_w3209_,
		_w3229_,
		_w3230_
	);
	LUT3 #(
		.INIT('h48)
	) name2768 (
		\P1_reg3_reg[26]/NET0131 ,
		_w524_,
		_w971_,
		_w3231_
	);
	LUT2 #(
		.INIT('h2)
	) name2769 (
		_w999_,
		_w2197_,
		_w3232_
	);
	LUT4 #(
		.INIT('h00b7)
	) name2770 (
		_w1432_,
		_w2197_,
		_w3085_,
		_w3232_,
		_w3233_
	);
	LUT4 #(
		.INIT('h08c8)
	) name2771 (
		_w999_,
		_w1114_,
		_w2197_,
		_w3058_,
		_w3234_
	);
	LUT4 #(
		.INIT('h9500)
	) name2772 (
		_w998_,
		_w1128_,
		_w1129_,
		_w2197_,
		_w3235_
	);
	LUT3 #(
		.INIT('h08)
	) name2773 (
		_w998_,
		_w2259_,
		_w2260_,
		_w3236_
	);
	LUT2 #(
		.INIT('h2)
	) name2774 (
		_w1183_,
		_w2197_,
		_w3237_
	);
	LUT4 #(
		.INIT('hdd05)
	) name2775 (
		_w1108_,
		_w1140_,
		_w1138_,
		_w2197_,
		_w3238_
	);
	LUT3 #(
		.INIT('h31)
	) name2776 (
		_w999_,
		_w3236_,
		_w3238_,
		_w3239_
	);
	LUT4 #(
		.INIT('h5700)
	) name2777 (
		_w1136_,
		_w3232_,
		_w3235_,
		_w3239_,
		_w3240_
	);
	LUT4 #(
		.INIT('hdf00)
	) name2778 (
		_w2197_,
		_w3038_,
		_w3039_,
		_w3240_,
		_w3241_
	);
	LUT4 #(
		.INIT('h0d00)
	) name2779 (
		_w1286_,
		_w3233_,
		_w3234_,
		_w3241_,
		_w3242_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name2780 (
		\P1_state_reg[0]/NET0131 ,
		_w526_,
		_w3231_,
		_w3242_,
		_w3243_
	);
	LUT4 #(
		.INIT('h9d5d)
	) name2781 (
		\P1_reg3_reg[26]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w510_,
		_w971_,
		_w3244_
	);
	LUT2 #(
		.INIT('hb)
	) name2782 (
		_w3243_,
		_w3244_,
		_w3245_
	);
	LUT2 #(
		.INIT('h2)
	) name2783 (
		_w1487_,
		_w1869_,
		_w3246_
	);
	LUT4 #(
		.INIT('h001f)
	) name2784 (
		_w1491_,
		_w1493_,
		_w1496_,
		_w1869_,
		_w3247_
	);
	LUT4 #(
		.INIT('h007b)
	) name2785 (
		_w1857_,
		_w2272_,
		_w3190_,
		_w3247_,
		_w3248_
	);
	LUT2 #(
		.INIT('h1)
	) name2786 (
		_w2276_,
		_w3248_,
		_w3249_
	);
	LUT4 #(
		.INIT('h00fe)
	) name2787 (
		_w1491_,
		_w1493_,
		_w1496_,
		_w1869_,
		_w3250_
	);
	LUT4 #(
		.INIT('h0057)
	) name2788 (
		_w2277_,
		_w3194_,
		_w3195_,
		_w3250_,
		_w3251_
	);
	LUT3 #(
		.INIT('h54)
	) name2789 (
		_w1869_,
		_w2086_,
		_w2280_,
		_w3252_
	);
	LUT3 #(
		.INIT('h07)
	) name2790 (
		_w1866_,
		_w2283_,
		_w3252_,
		_w3253_
	);
	LUT3 #(
		.INIT('hd0)
	) name2791 (
		_w2081_,
		_w3251_,
		_w3253_,
		_w3254_
	);
	LUT4 #(
		.INIT('hb040)
	) name2792 (
		_w2138_,
		_w2155_,
		_w2272_,
		_w3190_,
		_w3255_
	);
	LUT3 #(
		.INIT('h54)
	) name2793 (
		_w2192_,
		_w3247_,
		_w3255_,
		_w3256_
	);
	LUT4 #(
		.INIT('h007b)
	) name2794 (
		_w1857_,
		_w2277_,
		_w3190_,
		_w3250_,
		_w3257_
	);
	LUT2 #(
		.INIT('h2)
	) name2795 (
		_w2290_,
		_w3257_,
		_w3258_
	);
	LUT4 #(
		.INIT('h0100)
	) name2796 (
		_w3249_,
		_w3256_,
		_w3258_,
		_w3254_,
		_w3259_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name2797 (
		\P1_state_reg[0]/NET0131 ,
		_w1489_,
		_w3246_,
		_w3259_,
		_w3260_
	);
	LUT2 #(
		.INIT('h4)
	) name2798 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[20]/NET0131 ,
		_w3261_
	);
	LUT3 #(
		.INIT('h0b)
	) name2799 (
		_w1869_,
		_w2293_,
		_w3261_,
		_w3262_
	);
	LUT2 #(
		.INIT('hb)
	) name2800 (
		_w3260_,
		_w3262_,
		_w3263_
	);
	LUT2 #(
		.INIT('h2)
	) name2801 (
		_w1487_,
		_w1939_,
		_w3264_
	);
	LUT4 #(
		.INIT('h00fe)
	) name2802 (
		_w1491_,
		_w1493_,
		_w1496_,
		_w1939_,
		_w3265_
	);
	LUT4 #(
		.INIT('h0057)
	) name2803 (
		_w2277_,
		_w2573_,
		_w2574_,
		_w3265_,
		_w3266_
	);
	LUT2 #(
		.INIT('h2)
	) name2804 (
		_w2081_,
		_w3266_,
		_w3267_
	);
	LUT4 #(
		.INIT('h001f)
	) name2805 (
		_w1491_,
		_w1493_,
		_w1496_,
		_w1939_,
		_w3268_
	);
	LUT4 #(
		.INIT('h8288)
	) name2806 (
		_w2272_,
		_w2531_,
		_w2559_,
		_w2565_,
		_w3269_
	);
	LUT3 #(
		.INIT('h54)
	) name2807 (
		_w1939_,
		_w2086_,
		_w2280_,
		_w3270_
	);
	LUT3 #(
		.INIT('h07)
	) name2808 (
		_w1936_,
		_w2283_,
		_w3270_,
		_w3271_
	);
	LUT4 #(
		.INIT('hab00)
	) name2809 (
		_w2192_,
		_w3268_,
		_w3269_,
		_w3271_,
		_w3272_
	);
	LUT2 #(
		.INIT('h4)
	) name2810 (
		_w3267_,
		_w3272_,
		_w3273_
	);
	LUT4 #(
		.INIT('h007d)
	) name2811 (
		_w2277_,
		_w2531_,
		_w2548_,
		_w3265_,
		_w3274_
	);
	LUT4 #(
		.INIT('h007d)
	) name2812 (
		_w2272_,
		_w2531_,
		_w2548_,
		_w3268_,
		_w3275_
	);
	LUT4 #(
		.INIT('hf3a2)
	) name2813 (
		_w2276_,
		_w2290_,
		_w3274_,
		_w3275_,
		_w3276_
	);
	LUT4 #(
		.INIT('h3111)
	) name2814 (
		_w1489_,
		_w3264_,
		_w3273_,
		_w3276_,
		_w3277_
	);
	LUT4 #(
		.INIT('hb9b3)
	) name2815 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[25]/NET0131 ,
		_w1477_,
		_w1938_,
		_w3278_
	);
	LUT3 #(
		.INIT('h2f)
	) name2816 (
		\P1_state_reg[0]/NET0131 ,
		_w3277_,
		_w3278_,
		_w3279_
	);
	LUT2 #(
		.INIT('h2)
	) name2817 (
		\P1_reg2_reg[31]/NET0131 ,
		_w511_,
		_w3280_
	);
	LUT2 #(
		.INIT('h8)
	) name2818 (
		\P1_reg2_reg[31]/NET0131 ,
		_w524_,
		_w3281_
	);
	LUT4 #(
		.INIT('ha028)
	) name2819 (
		_w534_,
		_w1133_,
		_w1304_,
		_w1312_,
		_w3282_
	);
	LUT4 #(
		.INIT('h5455)
	) name2820 (
		\P1_reg2_reg[31]/NET0131 ,
		_w528_,
		_w530_,
		_w533_,
		_w3283_
	);
	LUT2 #(
		.INIT('h2)
	) name2821 (
		_w1136_,
		_w3283_,
		_w3284_
	);
	LUT2 #(
		.INIT('h4)
	) name2822 (
		_w3282_,
		_w3284_,
		_w3285_
	);
	LUT4 #(
		.INIT('h5100)
	) name2823 (
		_w1151_,
		_w1176_,
		_w1179_,
		_w1181_,
		_w3286_
	);
	LUT2 #(
		.INIT('h8)
	) name2824 (
		_w534_,
		_w1183_,
		_w3287_
	);
	LUT2 #(
		.INIT('h8)
	) name2825 (
		_w534_,
		_w1138_,
		_w3288_
	);
	LUT4 #(
		.INIT('h1200)
	) name2826 (
		\P2_datao_reg[31]/NET0131 ,
		_w541_,
		_w1303_,
		_w3288_,
		_w3289_
	);
	LUT4 #(
		.INIT('h0a02)
	) name2827 (
		\P1_reg2_reg[31]/NET0131 ,
		_w534_,
		_w1135_,
		_w1141_,
		_w3290_
	);
	LUT2 #(
		.INIT('h1)
	) name2828 (
		_w1144_,
		_w3290_,
		_w3291_
	);
	LUT2 #(
		.INIT('h4)
	) name2829 (
		_w3289_,
		_w3291_,
		_w3292_
	);
	LUT3 #(
		.INIT('h70)
	) name2830 (
		_w3286_,
		_w3287_,
		_w3292_,
		_w3293_
	);
	LUT4 #(
		.INIT('h1311)
	) name2831 (
		_w526_,
		_w3281_,
		_w3285_,
		_w3293_,
		_w3294_
	);
	LUT3 #(
		.INIT('hce)
	) name2832 (
		\P1_state_reg[0]/NET0131 ,
		_w3280_,
		_w3294_,
		_w3295_
	);
	LUT4 #(
		.INIT('h70d0)
	) name2833 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg0_reg[25]/NET0131 ,
		_w1476_,
		_w3296_
	);
	LUT2 #(
		.INIT('h8)
	) name2834 (
		\P2_reg0_reg[25]/NET0131 ,
		_w1487_,
		_w3297_
	);
	LUT4 #(
		.INIT('h111d)
	) name2835 (
		\P2_reg0_reg[25]/NET0131 ,
		_w2272_,
		_w2573_,
		_w2574_,
		_w3298_
	);
	LUT2 #(
		.INIT('h2)
	) name2836 (
		_w2081_,
		_w3298_,
		_w3299_
	);
	LUT4 #(
		.INIT('haaa8)
	) name2837 (
		\P2_reg0_reg[25]/NET0131 ,
		_w1491_,
		_w1493_,
		_w1496_,
		_w3300_
	);
	LUT4 #(
		.INIT('h8288)
	) name2838 (
		_w2277_,
		_w2531_,
		_w2559_,
		_w2565_,
		_w3301_
	);
	LUT3 #(
		.INIT('ha2)
	) name2839 (
		\P2_reg0_reg[25]/NET0131 ,
		_w2633_,
		_w2634_,
		_w3302_
	);
	LUT3 #(
		.INIT('h07)
	) name2840 (
		_w2277_,
		_w2567_,
		_w3302_,
		_w3303_
	);
	LUT4 #(
		.INIT('hab00)
	) name2841 (
		_w2192_,
		_w3300_,
		_w3301_,
		_w3303_,
		_w3304_
	);
	LUT2 #(
		.INIT('h4)
	) name2842 (
		_w3299_,
		_w3304_,
		_w3305_
	);
	LUT4 #(
		.INIT('h1dd1)
	) name2843 (
		\P2_reg0_reg[25]/NET0131 ,
		_w2277_,
		_w2531_,
		_w2548_,
		_w3306_
	);
	LUT4 #(
		.INIT('h1dd1)
	) name2844 (
		\P2_reg0_reg[25]/NET0131 ,
		_w2272_,
		_w2531_,
		_w2548_,
		_w3307_
	);
	LUT4 #(
		.INIT('hfa32)
	) name2845 (
		_w2276_,
		_w2290_,
		_w3306_,
		_w3307_,
		_w3308_
	);
	LUT4 #(
		.INIT('h3111)
	) name2846 (
		_w1489_,
		_w3297_,
		_w3305_,
		_w3308_,
		_w3309_
	);
	LUT3 #(
		.INIT('hce)
	) name2847 (
		\P1_state_reg[0]/NET0131 ,
		_w3296_,
		_w3309_,
		_w3310_
	);
	LUT4 #(
		.INIT('h70d0)
	) name2848 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg0_reg[24]/NET0131 ,
		_w1476_,
		_w3311_
	);
	LUT2 #(
		.INIT('h8)
	) name2849 (
		\P2_reg0_reg[24]/NET0131 ,
		_w1487_,
		_w3312_
	);
	LUT4 #(
		.INIT('h20e0)
	) name2850 (
		\P2_reg0_reg[24]/NET0131 ,
		_w2272_,
		_w2290_,
		_w2440_,
		_w3313_
	);
	LUT4 #(
		.INIT('h08c8)
	) name2851 (
		\P2_reg0_reg[24]/NET0131 ,
		_w2081_,
		_w2272_,
		_w2443_,
		_w3314_
	);
	LUT3 #(
		.INIT('ha2)
	) name2852 (
		\P2_reg0_reg[24]/NET0131 ,
		_w2633_,
		_w2634_,
		_w3315_
	);
	LUT4 #(
		.INIT('h00ef)
	) name2853 (
		_w1509_,
		_w1953_,
		_w2920_,
		_w3315_,
		_w3316_
	);
	LUT2 #(
		.INIT('h4)
	) name2854 (
		_w3314_,
		_w3316_,
		_w3317_
	);
	LUT4 #(
		.INIT('h0232)
	) name2855 (
		\P2_reg0_reg[24]/NET0131 ,
		_w2192_,
		_w2277_,
		_w2453_,
		_w3318_
	);
	LUT4 #(
		.INIT('h0232)
	) name2856 (
		\P2_reg0_reg[24]/NET0131 ,
		_w2276_,
		_w2277_,
		_w2440_,
		_w3319_
	);
	LUT4 #(
		.INIT('h0100)
	) name2857 (
		_w3313_,
		_w3318_,
		_w3319_,
		_w3317_,
		_w3320_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name2858 (
		\P1_state_reg[0]/NET0131 ,
		_w1489_,
		_w3312_,
		_w3320_,
		_w3321_
	);
	LUT2 #(
		.INIT('he)
	) name2859 (
		_w3311_,
		_w3321_,
		_w3322_
	);
	LUT4 #(
		.INIT('h70d0)
	) name2860 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg0_reg[26]/NET0131 ,
		_w1476_,
		_w3323_
	);
	LUT2 #(
		.INIT('h8)
	) name2861 (
		\P2_reg0_reg[26]/NET0131 ,
		_w1487_,
		_w3324_
	);
	LUT4 #(
		.INIT('h0232)
	) name2862 (
		\P2_reg0_reg[26]/NET0131 ,
		_w2276_,
		_w2277_,
		_w2480_,
		_w3325_
	);
	LUT4 #(
		.INIT('h02aa)
	) name2863 (
		\P2_reg0_reg[26]/NET0131 ,
		_w1491_,
		_w1493_,
		_w1496_,
		_w3326_
	);
	LUT4 #(
		.INIT('h8a88)
	) name2864 (
		_w2272_,
		_w2483_,
		_w2484_,
		_w2485_,
		_w3327_
	);
	LUT3 #(
		.INIT('ha2)
	) name2865 (
		\P2_reg0_reg[26]/NET0131 ,
		_w2633_,
		_w2634_,
		_w3328_
	);
	LUT4 #(
		.INIT('h00ef)
	) name2866 (
		_w1509_,
		_w1984_,
		_w2920_,
		_w3328_,
		_w3329_
	);
	LUT4 #(
		.INIT('h5700)
	) name2867 (
		_w2081_,
		_w3326_,
		_w3327_,
		_w3329_,
		_w3330_
	);
	LUT2 #(
		.INIT('h4)
	) name2868 (
		_w3325_,
		_w3330_,
		_w3331_
	);
	LUT4 #(
		.INIT('hd11d)
	) name2869 (
		\P2_reg0_reg[26]/NET0131 ,
		_w2277_,
		_w2463_,
		_w2506_,
		_w3332_
	);
	LUT4 #(
		.INIT('h20e0)
	) name2870 (
		\P2_reg0_reg[26]/NET0131 ,
		_w2272_,
		_w2290_,
		_w2480_,
		_w3333_
	);
	LUT3 #(
		.INIT('h0e)
	) name2871 (
		_w2192_,
		_w3332_,
		_w3333_,
		_w3334_
	);
	LUT4 #(
		.INIT('h3111)
	) name2872 (
		_w1489_,
		_w3324_,
		_w3331_,
		_w3334_,
		_w3335_
	);
	LUT3 #(
		.INIT('hce)
	) name2873 (
		\P1_state_reg[0]/NET0131 ,
		_w3323_,
		_w3335_,
		_w3336_
	);
	LUT2 #(
		.INIT('h2)
	) name2874 (
		\P1_reg2_reg[12]/NET0131 ,
		_w511_,
		_w3337_
	);
	LUT2 #(
		.INIT('h8)
	) name2875 (
		\P1_reg2_reg[12]/NET0131 ,
		_w524_,
		_w3338_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name2876 (
		\P1_reg2_reg[12]/NET0131 ,
		_w528_,
		_w530_,
		_w533_,
		_w3339_
	);
	LUT4 #(
		.INIT('h1000)
	) name2877 (
		_w799_,
		_w924_,
		_w1154_,
		_w1157_,
		_w3340_
	);
	LUT4 #(
		.INIT('h0705)
	) name2878 (
		_w752_,
		_w808_,
		_w1161_,
		_w3340_,
		_w3341_
	);
	LUT4 #(
		.INIT('h2a08)
	) name2879 (
		_w534_,
		_w537_,
		_w799_,
		_w3341_,
		_w3342_
	);
	LUT3 #(
		.INIT('ha8)
	) name2880 (
		_w1183_,
		_w3339_,
		_w3342_,
		_w3343_
	);
	LUT2 #(
		.INIT('h4)
	) name2881 (
		_w814_,
		_w1138_,
		_w3344_
	);
	LUT3 #(
		.INIT('h28)
	) name2882 (
		_w1286_,
		_w1387_,
		_w1454_,
		_w3345_
	);
	LUT3 #(
		.INIT('h82)
	) name2883 (
		_w1114_,
		_w1454_,
		_w2231_,
		_w3346_
	);
	LUT4 #(
		.INIT('haaa8)
	) name2884 (
		_w534_,
		_w3344_,
		_w3345_,
		_w3346_,
		_w3347_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name2885 (
		_w804_,
		_w814_,
		_w1117_,
		_w1119_,
		_w3348_
	);
	LUT4 #(
		.INIT('he020)
	) name2886 (
		\P1_reg2_reg[12]/NET0131 ,
		_w534_,
		_w1136_,
		_w3348_,
		_w3349_
	);
	LUT4 #(
		.INIT('h00ab)
	) name2887 (
		_w534_,
		_w1109_,
		_w1138_,
		_w1141_,
		_w3350_
	);
	LUT2 #(
		.INIT('h8)
	) name2888 (
		_w806_,
		_w1143_,
		_w3351_
	);
	LUT3 #(
		.INIT('h0d)
	) name2889 (
		\P1_reg2_reg[12]/NET0131 ,
		_w3350_,
		_w3351_,
		_w3352_
	);
	LUT2 #(
		.INIT('h4)
	) name2890 (
		_w3349_,
		_w3352_,
		_w3353_
	);
	LUT2 #(
		.INIT('h4)
	) name2891 (
		_w3347_,
		_w3353_,
		_w3354_
	);
	LUT4 #(
		.INIT('h1311)
	) name2892 (
		_w526_,
		_w3338_,
		_w3343_,
		_w3354_,
		_w3355_
	);
	LUT3 #(
		.INIT('hce)
	) name2893 (
		\P1_state_reg[0]/NET0131 ,
		_w3337_,
		_w3355_,
		_w3356_
	);
	LUT2 #(
		.INIT('h2)
	) name2894 (
		\P1_reg2_reg[26]/NET0131 ,
		_w511_,
		_w3357_
	);
	LUT2 #(
		.INIT('h8)
	) name2895 (
		\P1_reg2_reg[26]/NET0131 ,
		_w524_,
		_w3358_
	);
	LUT3 #(
		.INIT('h28)
	) name2896 (
		_w1286_,
		_w1432_,
		_w3085_,
		_w3359_
	);
	LUT4 #(
		.INIT('haa8a)
	) name2897 (
		_w534_,
		_w3040_,
		_w3062_,
		_w3359_,
		_w3360_
	);
	LUT2 #(
		.INIT('h8)
	) name2898 (
		_w999_,
		_w1143_,
		_w3361_
	);
	LUT4 #(
		.INIT('h00a2)
	) name2899 (
		\P1_reg2_reg[26]/NET0131 ,
		_w534_,
		_w1141_,
		_w1143_,
		_w3362_
	);
	LUT2 #(
		.INIT('h1)
	) name2900 (
		_w3361_,
		_w3362_,
		_w3363_
	);
	LUT4 #(
		.INIT('h1311)
	) name2901 (
		_w526_,
		_w3358_,
		_w3360_,
		_w3363_,
		_w3364_
	);
	LUT3 #(
		.INIT('hce)
	) name2902 (
		\P1_state_reg[0]/NET0131 ,
		_w3357_,
		_w3364_,
		_w3365_
	);
	LUT2 #(
		.INIT('h2)
	) name2903 (
		\P1_reg2_reg[27]/NET0131 ,
		_w511_,
		_w3366_
	);
	LUT2 #(
		.INIT('h8)
	) name2904 (
		\P1_reg2_reg[27]/NET0131 ,
		_w524_,
		_w3367_
	);
	LUT4 #(
		.INIT('h20e0)
	) name2905 (
		\P1_reg2_reg[27]/NET0131 ,
		_w534_,
		_w1286_,
		_w2856_,
		_w3368_
	);
	LUT4 #(
		.INIT('hddd1)
	) name2906 (
		\P1_reg2_reg[27]/NET0131 ,
		_w534_,
		_w1132_,
		_w2858_,
		_w3369_
	);
	LUT3 #(
		.INIT('h10)
	) name2907 (
		_w541_,
		_w1033_,
		_w1138_,
		_w3370_
	);
	LUT4 #(
		.INIT('h0200)
	) name2908 (
		_w534_,
		_w541_,
		_w1033_,
		_w1138_,
		_w3371_
	);
	LUT2 #(
		.INIT('h8)
	) name2909 (
		_w1035_,
		_w1143_,
		_w3372_
	);
	LUT4 #(
		.INIT('haa20)
	) name2910 (
		\P1_reg2_reg[27]/NET0131 ,
		_w534_,
		_w1138_,
		_w1141_,
		_w3373_
	);
	LUT2 #(
		.INIT('h1)
	) name2911 (
		_w3372_,
		_w3373_,
		_w3374_
	);
	LUT2 #(
		.INIT('h4)
	) name2912 (
		_w3371_,
		_w3374_,
		_w3375_
	);
	LUT3 #(
		.INIT('hd0)
	) name2913 (
		_w1136_,
		_w3369_,
		_w3375_,
		_w3376_
	);
	LUT2 #(
		.INIT('h4)
	) name2914 (
		_w3368_,
		_w3376_,
		_w3377_
	);
	LUT4 #(
		.INIT('h20e0)
	) name2915 (
		\P1_reg2_reg[27]/NET0131 ,
		_w534_,
		_w1114_,
		_w2883_,
		_w3378_
	);
	LUT4 #(
		.INIT('hddd1)
	) name2916 (
		\P1_reg2_reg[27]/NET0131 ,
		_w534_,
		_w2885_,
		_w2886_,
		_w3379_
	);
	LUT3 #(
		.INIT('h31)
	) name2917 (
		_w1183_,
		_w3378_,
		_w3379_,
		_w3380_
	);
	LUT4 #(
		.INIT('h3111)
	) name2918 (
		_w526_,
		_w3367_,
		_w3377_,
		_w3380_,
		_w3381_
	);
	LUT3 #(
		.INIT('hce)
	) name2919 (
		\P1_state_reg[0]/NET0131 ,
		_w3366_,
		_w3381_,
		_w3382_
	);
	LUT4 #(
		.INIT('h70d0)
	) name2920 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg1_reg[24]/NET0131 ,
		_w1476_,
		_w3383_
	);
	LUT2 #(
		.INIT('h8)
	) name2921 (
		\P2_reg1_reg[24]/NET0131 ,
		_w1487_,
		_w3384_
	);
	LUT4 #(
		.INIT('h08c8)
	) name2922 (
		\P2_reg1_reg[24]/NET0131 ,
		_w2038_,
		_w2039_,
		_w2440_,
		_w3385_
	);
	LUT4 #(
		.INIT('h20e0)
	) name2923 (
		\P2_reg1_reg[24]/NET0131 ,
		_w1497_,
		_w2081_,
		_w2443_,
		_w3386_
	);
	LUT3 #(
		.INIT('ha2)
	) name2924 (
		\P2_reg1_reg[24]/NET0131 ,
		_w2633_,
		_w2660_,
		_w3387_
	);
	LUT4 #(
		.INIT('h00ef)
	) name2925 (
		_w1509_,
		_w1953_,
		_w2963_,
		_w3387_,
		_w3388_
	);
	LUT2 #(
		.INIT('h4)
	) name2926 (
		_w3386_,
		_w3388_,
		_w3389_
	);
	LUT4 #(
		.INIT('h20e0)
	) name2927 (
		\P2_reg1_reg[24]/NET0131 ,
		_w1497_,
		_w2188_,
		_w2453_,
		_w3390_
	);
	LUT4 #(
		.INIT('h20e0)
	) name2928 (
		\P2_reg1_reg[24]/NET0131 ,
		_w2039_,
		_w2193_,
		_w2453_,
		_w3391_
	);
	LUT4 #(
		.INIT('h0100)
	) name2929 (
		_w3385_,
		_w3390_,
		_w3391_,
		_w3389_,
		_w3392_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name2930 (
		\P1_state_reg[0]/NET0131 ,
		_w1489_,
		_w3384_,
		_w3392_,
		_w3393_
	);
	LUT2 #(
		.INIT('he)
	) name2931 (
		_w3383_,
		_w3393_,
		_w3394_
	);
	LUT4 #(
		.INIT('h70d0)
	) name2932 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg1_reg[25]/NET0131 ,
		_w1476_,
		_w3395_
	);
	LUT2 #(
		.INIT('h8)
	) name2933 (
		\P2_reg1_reg[25]/NET0131 ,
		_w1487_,
		_w3396_
	);
	LUT4 #(
		.INIT('haa02)
	) name2934 (
		\P2_reg1_reg[25]/NET0131 ,
		_w1491_,
		_w1493_,
		_w1496_,
		_w3397_
	);
	LUT4 #(
		.INIT('h1dd1)
	) name2935 (
		\P2_reg1_reg[25]/NET0131 ,
		_w2039_,
		_w2531_,
		_w2548_,
		_w3398_
	);
	LUT2 #(
		.INIT('h2)
	) name2936 (
		_w2038_,
		_w3398_,
		_w3399_
	);
	LUT3 #(
		.INIT('ha2)
	) name2937 (
		\P2_reg1_reg[25]/NET0131 ,
		_w2633_,
		_w2660_,
		_w3400_
	);
	LUT3 #(
		.INIT('h07)
	) name2938 (
		_w2039_,
		_w2567_,
		_w3400_,
		_w3401_
	);
	LUT4 #(
		.INIT('h5700)
	) name2939 (
		_w2193_,
		_w2577_,
		_w3397_,
		_w3401_,
		_w3402_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name2940 (
		\P2_reg1_reg[25]/NET0131 ,
		_w1491_,
		_w1493_,
		_w1496_,
		_w3403_
	);
	LUT4 #(
		.INIT('h111d)
	) name2941 (
		\P2_reg1_reg[25]/NET0131 ,
		_w1497_,
		_w2573_,
		_w2574_,
		_w3404_
	);
	LUT2 #(
		.INIT('h2)
	) name2942 (
		_w2081_,
		_w3404_,
		_w3405_
	);
	LUT3 #(
		.INIT('ha8)
	) name2943 (
		_w2188_,
		_w2566_,
		_w3403_,
		_w3406_
	);
	LUT3 #(
		.INIT('h10)
	) name2944 (
		_w3405_,
		_w3406_,
		_w3402_,
		_w3407_
	);
	LUT4 #(
		.INIT('h1311)
	) name2945 (
		_w1489_,
		_w3396_,
		_w3399_,
		_w3407_,
		_w3408_
	);
	LUT3 #(
		.INIT('hce)
	) name2946 (
		\P1_state_reg[0]/NET0131 ,
		_w3395_,
		_w3408_,
		_w3409_
	);
	LUT4 #(
		.INIT('h70d0)
	) name2947 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg1_reg[26]/NET0131 ,
		_w1476_,
		_w3410_
	);
	LUT2 #(
		.INIT('h8)
	) name2948 (
		\P2_reg1_reg[26]/NET0131 ,
		_w1487_,
		_w3411_
	);
	LUT4 #(
		.INIT('h08c8)
	) name2949 (
		\P2_reg1_reg[26]/NET0131 ,
		_w2038_,
		_w2039_,
		_w2480_,
		_w3412_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name2950 (
		\P2_reg1_reg[26]/NET0131 ,
		_w1491_,
		_w1493_,
		_w1496_,
		_w3413_
	);
	LUT4 #(
		.INIT('h8a88)
	) name2951 (
		_w1497_,
		_w2483_,
		_w2484_,
		_w2485_,
		_w3414_
	);
	LUT3 #(
		.INIT('ha2)
	) name2952 (
		\P2_reg1_reg[26]/NET0131 ,
		_w2633_,
		_w2660_,
		_w3415_
	);
	LUT4 #(
		.INIT('h00ef)
	) name2953 (
		_w1509_,
		_w1984_,
		_w2963_,
		_w3415_,
		_w3416_
	);
	LUT4 #(
		.INIT('h5700)
	) name2954 (
		_w2081_,
		_w3413_,
		_w3414_,
		_w3416_,
		_w3417_
	);
	LUT2 #(
		.INIT('h4)
	) name2955 (
		_w3412_,
		_w3417_,
		_w3418_
	);
	LUT4 #(
		.INIT('hd11d)
	) name2956 (
		\P2_reg1_reg[26]/NET0131 ,
		_w2039_,
		_w2463_,
		_w2506_,
		_w3419_
	);
	LUT4 #(
		.INIT('hd11d)
	) name2957 (
		\P2_reg1_reg[26]/NET0131 ,
		_w1497_,
		_w2463_,
		_w2506_,
		_w3420_
	);
	LUT4 #(
		.INIT('hf351)
	) name2958 (
		_w2188_,
		_w2193_,
		_w3419_,
		_w3420_,
		_w3421_
	);
	LUT4 #(
		.INIT('h3111)
	) name2959 (
		_w1489_,
		_w3411_,
		_w3418_,
		_w3421_,
		_w3422_
	);
	LUT3 #(
		.INIT('hce)
	) name2960 (
		\P1_state_reg[0]/NET0131 ,
		_w3410_,
		_w3422_,
		_w3423_
	);
	LUT2 #(
		.INIT('h2)
	) name2961 (
		\P1_reg0_reg[26]/NET0131 ,
		_w511_,
		_w3424_
	);
	LUT2 #(
		.INIT('h8)
	) name2962 (
		\P1_reg0_reg[26]/NET0131 ,
		_w524_,
		_w3425_
	);
	LUT4 #(
		.INIT('h82c0)
	) name2963 (
		_w652_,
		_w1104_,
		_w1106_,
		_w1111_,
		_w3426_
	);
	LUT4 #(
		.INIT('h222a)
	) name2964 (
		\P1_reg0_reg[26]/NET0131 ,
		_w2425_,
		_w2688_,
		_w3426_,
		_w3427_
	);
	LUT4 #(
		.INIT('haa8a)
	) name2965 (
		_w2688_,
		_w3040_,
		_w3062_,
		_w3359_,
		_w3428_
	);
	LUT4 #(
		.INIT('h1113)
	) name2966 (
		_w526_,
		_w3425_,
		_w3427_,
		_w3428_,
		_w3429_
	);
	LUT3 #(
		.INIT('hce)
	) name2967 (
		\P1_state_reg[0]/NET0131 ,
		_w3424_,
		_w3429_,
		_w3430_
	);
	LUT2 #(
		.INIT('h2)
	) name2968 (
		\P1_reg0_reg[27]/NET0131 ,
		_w511_,
		_w3431_
	);
	LUT2 #(
		.INIT('h8)
	) name2969 (
		\P1_reg0_reg[27]/NET0131 ,
		_w524_,
		_w3432_
	);
	LUT4 #(
		.INIT('h08c8)
	) name2970 (
		\P1_reg0_reg[27]/NET0131 ,
		_w1286_,
		_w2688_,
		_w2856_,
		_w3433_
	);
	LUT4 #(
		.INIT('h00fb)
	) name2971 (
		_w1132_,
		_w1136_,
		_w2858_,
		_w3370_,
		_w3434_
	);
	LUT3 #(
		.INIT('ha2)
	) name2972 (
		\P1_reg0_reg[27]/NET0131 ,
		_w2692_,
		_w3005_,
		_w3435_
	);
	LUT3 #(
		.INIT('h0d)
	) name2973 (
		_w2688_,
		_w3434_,
		_w3435_,
		_w3436_
	);
	LUT2 #(
		.INIT('h4)
	) name2974 (
		_w3433_,
		_w3436_,
		_w3437_
	);
	LUT4 #(
		.INIT('hddd1)
	) name2975 (
		\P1_reg0_reg[27]/NET0131 ,
		_w2688_,
		_w2885_,
		_w2886_,
		_w3438_
	);
	LUT4 #(
		.INIT('h08c8)
	) name2976 (
		\P1_reg0_reg[27]/NET0131 ,
		_w1114_,
		_w2688_,
		_w2883_,
		_w3439_
	);
	LUT3 #(
		.INIT('h0d)
	) name2977 (
		_w1183_,
		_w3438_,
		_w3439_,
		_w3440_
	);
	LUT4 #(
		.INIT('h3111)
	) name2978 (
		_w526_,
		_w3432_,
		_w3437_,
		_w3440_,
		_w3441_
	);
	LUT3 #(
		.INIT('hce)
	) name2979 (
		\P1_state_reg[0]/NET0131 ,
		_w3431_,
		_w3441_,
		_w3442_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name2980 (
		_w511_,
		_w519_,
		_w522_,
		_w517_,
		_w3443_
	);
	LUT2 #(
		.INIT('h1)
	) name2981 (
		\P1_reg1_reg[27]/NET0131 ,
		_w3443_,
		_w3444_
	);
	LUT4 #(
		.INIT('hddd1)
	) name2982 (
		\P1_reg1_reg[27]/NET0131 ,
		_w2421_,
		_w2885_,
		_w2886_,
		_w3445_
	);
	LUT4 #(
		.INIT('h4c44)
	) name2983 (
		\P1_reg1_reg[27]/NET0131 ,
		_w511_,
		_w523_,
		_w3026_,
		_w3446_
	);
	LUT3 #(
		.INIT('hd0)
	) name2984 (
		_w2421_,
		_w3434_,
		_w3446_,
		_w3447_
	);
	LUT3 #(
		.INIT('hd0)
	) name2985 (
		_w1183_,
		_w3445_,
		_w3447_,
		_w3448_
	);
	LUT4 #(
		.INIT('h08c8)
	) name2986 (
		\P1_reg1_reg[27]/NET0131 ,
		_w1114_,
		_w2421_,
		_w2883_,
		_w3449_
	);
	LUT4 #(
		.INIT('h08c8)
	) name2987 (
		\P1_reg1_reg[27]/NET0131 ,
		_w1286_,
		_w2421_,
		_w2856_,
		_w3450_
	);
	LUT2 #(
		.INIT('h1)
	) name2988 (
		_w3449_,
		_w3450_,
		_w3451_
	);
	LUT3 #(
		.INIT('h15)
	) name2989 (
		_w3444_,
		_w3448_,
		_w3451_,
		_w3452_
	);
	LUT2 #(
		.INIT('h8)
	) name2990 (
		_w524_,
		_w806_,
		_w3453_
	);
	LUT4 #(
		.INIT('h1f00)
	) name2991 (
		_w528_,
		_w530_,
		_w533_,
		_w806_,
		_w3454_
	);
	LUT4 #(
		.INIT('h7020)
	) name2992 (
		_w537_,
		_w799_,
		_w2197_,
		_w3341_,
		_w3455_
	);
	LUT4 #(
		.INIT('hc808)
	) name2993 (
		_w806_,
		_w1136_,
		_w2197_,
		_w3348_,
		_w3456_
	);
	LUT4 #(
		.INIT('h888a)
	) name2994 (
		_w806_,
		_w1141_,
		_w2197_,
		_w3118_,
		_w3457_
	);
	LUT3 #(
		.INIT('h04)
	) name2995 (
		_w814_,
		_w2259_,
		_w2260_,
		_w3458_
	);
	LUT2 #(
		.INIT('h1)
	) name2996 (
		_w3457_,
		_w3458_,
		_w3459_
	);
	LUT2 #(
		.INIT('h4)
	) name2997 (
		_w3456_,
		_w3459_,
		_w3460_
	);
	LUT4 #(
		.INIT('h5700)
	) name2998 (
		_w2197_,
		_w3345_,
		_w3346_,
		_w3460_,
		_w3461_
	);
	LUT4 #(
		.INIT('h5700)
	) name2999 (
		_w1183_,
		_w3454_,
		_w3455_,
		_w3461_,
		_w3462_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name3000 (
		\P1_state_reg[0]/NET0131 ,
		_w526_,
		_w3453_,
		_w3462_,
		_w3463_
	);
	LUT2 #(
		.INIT('h2)
	) name3001 (
		\P1_reg3_reg[12]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w3464_
	);
	LUT3 #(
		.INIT('h07)
	) name3002 (
		_w806_,
		_w1294_,
		_w3464_,
		_w3465_
	);
	LUT2 #(
		.INIT('hb)
	) name3003 (
		_w3463_,
		_w3465_,
		_w3466_
	);
	LUT3 #(
		.INIT('h02)
	) name3004 (
		_w524_,
		_w634_,
		_w739_,
		_w3467_
	);
	LUT2 #(
		.INIT('h2)
	) name3005 (
		_w740_,
		_w2197_,
		_w3468_
	);
	LUT4 #(
		.INIT('h20aa)
	) name3006 (
		_w3071_,
		_w3076_,
		_w3077_,
		_w3079_,
		_w3469_
	);
	LUT4 #(
		.INIT('h4484)
	) name3007 (
		_w1423_,
		_w2197_,
		_w3080_,
		_w3469_,
		_w3470_
	);
	LUT4 #(
		.INIT('h60c0)
	) name3008 (
		_w717_,
		_w738_,
		_w2197_,
		_w3116_,
		_w3471_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name3009 (
		_w740_,
		_w1138_,
		_w1141_,
		_w2197_,
		_w3472_
	);
	LUT3 #(
		.INIT('h0b)
	) name3010 (
		_w738_,
		_w2261_,
		_w3472_,
		_w3473_
	);
	LUT4 #(
		.INIT('h5700)
	) name3011 (
		_w1136_,
		_w3468_,
		_w3471_,
		_w3473_,
		_w3474_
	);
	LUT4 #(
		.INIT('h5700)
	) name3012 (
		_w1286_,
		_w3468_,
		_w3470_,
		_w3474_,
		_w3475_
	);
	LUT4 #(
		.INIT('h2a22)
	) name3013 (
		_w3044_,
		_w3045_,
		_w3052_,
		_w3053_,
		_w3476_
	);
	LUT4 #(
		.INIT('h8848)
	) name3014 (
		_w1423_,
		_w2197_,
		_w3046_,
		_w3476_,
		_w3477_
	);
	LUT3 #(
		.INIT('ha8)
	) name3015 (
		_w1114_,
		_w3468_,
		_w3477_,
		_w3478_
	);
	LUT4 #(
		.INIT('h6555)
	) name3016 (
		_w679_,
		_w745_,
		_w1161_,
		_w1163_,
		_w3479_
	);
	LUT4 #(
		.INIT('h7020)
	) name3017 (
		_w537_,
		_w722_,
		_w2197_,
		_w3479_,
		_w3480_
	);
	LUT3 #(
		.INIT('ha8)
	) name3018 (
		_w1183_,
		_w3468_,
		_w3480_,
		_w3481_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name3019 (
		_w526_,
		_w3478_,
		_w3481_,
		_w3475_,
		_w3482_
	);
	LUT2 #(
		.INIT('h2)
	) name3020 (
		\P1_reg3_reg[18]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w3483_
	);
	LUT4 #(
		.INIT('h00ef)
	) name3021 (
		_w634_,
		_w739_,
		_w1294_,
		_w3483_,
		_w3484_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name3022 (
		\P1_state_reg[0]/NET0131 ,
		_w3467_,
		_w3482_,
		_w3484_,
		_w3485_
	);
	LUT2 #(
		.INIT('h8)
	) name3023 (
		_w524_,
		_w719_,
		_w3486_
	);
	LUT4 #(
		.INIT('h1f00)
	) name3024 (
		_w528_,
		_w530_,
		_w533_,
		_w719_,
		_w3487_
	);
	LUT4 #(
		.INIT('h1444)
	) name3025 (
		_w537_,
		_w745_,
		_w1161_,
		_w1163_,
		_w3488_
	);
	LUT4 #(
		.INIT('h0200)
	) name3026 (
		_w537_,
		_w789_,
		_w788_,
		_w790_,
		_w3489_
	);
	LUT4 #(
		.INIT('h3331)
	) name3027 (
		_w2197_,
		_w3487_,
		_w3488_,
		_w3489_,
		_w3490_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name3028 (
		_w717_,
		_w786_,
		_w1120_,
		_w1122_,
		_w3491_
	);
	LUT4 #(
		.INIT('hc808)
	) name3029 (
		_w719_,
		_w1136_,
		_w2197_,
		_w3491_,
		_w3492_
	);
	LUT3 #(
		.INIT('h04)
	) name3030 (
		_w717_,
		_w2259_,
		_w2260_,
		_w3493_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name3031 (
		_w719_,
		_w1138_,
		_w1141_,
		_w2197_,
		_w3494_
	);
	LUT2 #(
		.INIT('h1)
	) name3032 (
		_w3493_,
		_w3494_,
		_w3495_
	);
	LUT2 #(
		.INIT('h4)
	) name3033 (
		_w3492_,
		_w3495_,
		_w3496_
	);
	LUT3 #(
		.INIT('hd0)
	) name3034 (
		_w1183_,
		_w3490_,
		_w3496_,
		_w3497_
	);
	LUT4 #(
		.INIT('h5d00)
	) name3035 (
		_w1193_,
		_w1202_,
		_w1237_,
		_w1243_,
		_w3498_
	);
	LUT4 #(
		.INIT('h0b07)
	) name3036 (
		_w1431_,
		_w2197_,
		_w3487_,
		_w3498_,
		_w3499_
	);
	LUT4 #(
		.INIT('hd02f)
	) name3037 (
		_w794_,
		_w954_,
		_w957_,
		_w1431_,
		_w3500_
	);
	LUT4 #(
		.INIT('hc808)
	) name3038 (
		_w719_,
		_w1114_,
		_w2197_,
		_w3500_,
		_w3501_
	);
	LUT3 #(
		.INIT('h0d)
	) name3039 (
		_w1286_,
		_w3499_,
		_w3501_,
		_w3502_
	);
	LUT4 #(
		.INIT('h3111)
	) name3040 (
		_w526_,
		_w3486_,
		_w3497_,
		_w3502_,
		_w3503_
	);
	LUT2 #(
		.INIT('h2)
	) name3041 (
		\P1_reg3_reg[17]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w3504_
	);
	LUT4 #(
		.INIT('h6c00)
	) name3042 (
		\P1_reg3_reg[16]/NET0131 ,
		\P1_reg3_reg[17]/NET0131 ,
		_w718_,
		_w1294_,
		_w3505_
	);
	LUT2 #(
		.INIT('h1)
	) name3043 (
		_w3504_,
		_w3505_,
		_w3506_
	);
	LUT3 #(
		.INIT('h2f)
	) name3044 (
		\P1_state_reg[0]/NET0131 ,
		_w3503_,
		_w3506_,
		_w3507_
	);
	LUT4 #(
		.INIT('h70d0)
	) name3045 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg2_reg[23]/NET0131 ,
		_w1476_,
		_w3508_
	);
	LUT2 #(
		.INIT('h8)
	) name3046 (
		\P2_reg2_reg[23]/NET0131 ,
		_w1487_,
		_w3509_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name3047 (
		\P2_reg2_reg[23]/NET0131 ,
		_w1491_,
		_w1493_,
		_w1496_,
		_w3510_
	);
	LUT3 #(
		.INIT('h1e)
	) name3048 (
		_w1509_,
		_w1903_,
		_w1907_,
		_w3511_
	);
	LUT4 #(
		.INIT('h4f00)
	) name3049 (
		_w2309_,
		_w2312_,
		_w2315_,
		_w2322_,
		_w3512_
	);
	LUT2 #(
		.INIT('h8)
	) name3050 (
		_w2317_,
		_w2333_,
		_w3513_
	);
	LUT4 #(
		.INIT('h2f00)
	) name3051 (
		_w2316_,
		_w2324_,
		_w2325_,
		_w2333_,
		_w3514_
	);
	LUT2 #(
		.INIT('h2)
	) name3052 (
		_w2337_,
		_w3514_,
		_w3515_
	);
	LUT4 #(
		.INIT('h65aa)
	) name3053 (
		_w3511_,
		_w3512_,
		_w3513_,
		_w3515_,
		_w3516_
	);
	LUT4 #(
		.INIT('h20e0)
	) name3054 (
		\P2_reg2_reg[23]/NET0131 ,
		_w1497_,
		_w2038_,
		_w3516_,
		_w3517_
	);
	LUT4 #(
		.INIT('haa02)
	) name3055 (
		\P2_reg2_reg[23]/NET0131 ,
		_w1491_,
		_w1493_,
		_w1496_,
		_w3518_
	);
	LUT4 #(
		.INIT('hef00)
	) name3056 (
		_w1919_,
		_w1918_,
		_w1920_,
		_w2042_,
		_w3519_
	);
	LUT2 #(
		.INIT('h1)
	) name3057 (
		_w2042_,
		_w2073_,
		_w3520_
	);
	LUT4 #(
		.INIT('h020f)
	) name3058 (
		_w1960_,
		_w2814_,
		_w3519_,
		_w3520_,
		_w3521_
	);
	LUT4 #(
		.INIT('h20e0)
	) name3059 (
		\P2_reg2_reg[23]/NET0131 ,
		_w2039_,
		_w2081_,
		_w3521_,
		_w3522_
	);
	LUT2 #(
		.INIT('h8)
	) name3060 (
		_w2365_,
		_w2380_,
		_w3523_
	);
	LUT4 #(
		.INIT('h2f00)
	) name3061 (
		_w2368_,
		_w2363_,
		_w2373_,
		_w3523_,
		_w3524_
	);
	LUT4 #(
		.INIT('hf200)
	) name3062 (
		_w2364_,
		_w2375_,
		_w2376_,
		_w2380_,
		_w3525_
	);
	LUT2 #(
		.INIT('h2)
	) name3063 (
		_w2349_,
		_w3525_,
		_w3526_
	);
	LUT4 #(
		.INIT('h8288)
	) name3064 (
		_w2039_,
		_w3511_,
		_w3524_,
		_w3526_,
		_w3527_
	);
	LUT3 #(
		.INIT('ha8)
	) name3065 (
		_w2188_,
		_w3518_,
		_w3527_,
		_w3528_
	);
	LUT4 #(
		.INIT('h8288)
	) name3066 (
		_w1497_,
		_w3511_,
		_w3524_,
		_w3526_,
		_w3529_
	);
	LUT3 #(
		.INIT('ha8)
	) name3067 (
		\P2_reg2_reg[23]/NET0131 ,
		_w2086_,
		_w2087_,
		_w3530_
	);
	LUT2 #(
		.INIT('h4)
	) name3068 (
		_w1904_,
		_w2088_,
		_w3531_
	);
	LUT4 #(
		.INIT('h00ef)
	) name3069 (
		_w1509_,
		_w1903_,
		_w2085_,
		_w3531_,
		_w3532_
	);
	LUT2 #(
		.INIT('h4)
	) name3070 (
		_w3530_,
		_w3532_,
		_w3533_
	);
	LUT4 #(
		.INIT('h5700)
	) name3071 (
		_w2193_,
		_w3510_,
		_w3529_,
		_w3533_,
		_w3534_
	);
	LUT4 #(
		.INIT('h0100)
	) name3072 (
		_w3517_,
		_w3522_,
		_w3528_,
		_w3534_,
		_w3535_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name3073 (
		\P1_state_reg[0]/NET0131 ,
		_w1489_,
		_w3509_,
		_w3535_,
		_w3536_
	);
	LUT2 #(
		.INIT('he)
	) name3074 (
		_w3508_,
		_w3536_,
		_w3537_
	);
	LUT2 #(
		.INIT('h8)
	) name3075 (
		_w524_,
		_w1075_,
		_w3538_
	);
	LUT4 #(
		.INIT('h1f00)
	) name3076 (
		_w528_,
		_w530_,
		_w533_,
		_w1075_,
		_w3539_
	);
	LUT4 #(
		.INIT('h8000)
	) name3077 (
		_w1167_,
		_w1165_,
		_w1161_,
		_w1163_,
		_w3540_
	);
	LUT4 #(
		.INIT('h5504)
	) name3078 (
		_w537_,
		_w1070_,
		_w3136_,
		_w3540_,
		_w3541_
	);
	LUT2 #(
		.INIT('h8)
	) name3079 (
		_w537_,
		_w706_,
		_w3542_
	);
	LUT4 #(
		.INIT('h3331)
	) name3080 (
		_w2197_,
		_w3539_,
		_w3541_,
		_w3542_,
		_w3543_
	);
	LUT4 #(
		.INIT('hb040)
	) name3081 (
		_w1238_,
		_w1251_,
		_w1286_,
		_w1430_,
		_w3544_
	);
	LUT3 #(
		.INIT('h84)
	) name3082 (
		_w965_,
		_w1114_,
		_w1430_,
		_w3545_
	);
	LUT4 #(
		.INIT('h4000)
	) name3083 (
		_w1074_,
		_w1120_,
		_w1122_,
		_w1125_,
		_w3546_
	);
	LUT4 #(
		.INIT('h9555)
	) name3084 (
		_w1074_,
		_w1120_,
		_w1122_,
		_w1125_,
		_w3547_
	);
	LUT4 #(
		.INIT('hc808)
	) name3085 (
		_w1075_,
		_w1136_,
		_w2197_,
		_w3547_,
		_w3548_
	);
	LUT4 #(
		.INIT('h0010)
	) name3086 (
		_w541_,
		_w1073_,
		_w2259_,
		_w2260_,
		_w3549_
	);
	LUT4 #(
		.INIT('h888a)
	) name3087 (
		_w1075_,
		_w1141_,
		_w2197_,
		_w3118_,
		_w3550_
	);
	LUT2 #(
		.INIT('h1)
	) name3088 (
		_w3549_,
		_w3550_,
		_w3551_
	);
	LUT2 #(
		.INIT('h4)
	) name3089 (
		_w3548_,
		_w3551_,
		_w3552_
	);
	LUT4 #(
		.INIT('h5700)
	) name3090 (
		_w2197_,
		_w3544_,
		_w3545_,
		_w3552_,
		_w3553_
	);
	LUT4 #(
		.INIT('h08aa)
	) name3091 (
		_w526_,
		_w1183_,
		_w3543_,
		_w3553_,
		_w3554_
	);
	LUT4 #(
		.INIT('h6a00)
	) name3092 (
		\P1_reg3_reg[21]/NET0131 ,
		_w634_,
		_w635_,
		_w1294_,
		_w3555_
	);
	LUT2 #(
		.INIT('h2)
	) name3093 (
		\P1_reg3_reg[21]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w3556_
	);
	LUT2 #(
		.INIT('h1)
	) name3094 (
		_w3555_,
		_w3556_,
		_w3557_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name3095 (
		\P1_state_reg[0]/NET0131 ,
		_w3538_,
		_w3554_,
		_w3557_,
		_w3558_
	);
	LUT2 #(
		.INIT('h2)
	) name3096 (
		_w1487_,
		_w1904_,
		_w3559_
	);
	LUT4 #(
		.INIT('h10d0)
	) name3097 (
		_w1904_,
		_w2277_,
		_w2290_,
		_w3516_,
		_w3560_
	);
	LUT4 #(
		.INIT('h001f)
	) name3098 (
		_w1491_,
		_w1493_,
		_w1496_,
		_w1904_,
		_w3561_
	);
	LUT4 #(
		.INIT('h010d)
	) name3099 (
		_w1904_,
		_w2272_,
		_w2276_,
		_w3516_,
		_w3562_
	);
	LUT4 #(
		.INIT('h04c4)
	) name3100 (
		_w1904_,
		_w2081_,
		_w2277_,
		_w3521_,
		_w3563_
	);
	LUT4 #(
		.INIT('h8288)
	) name3101 (
		_w2272_,
		_w3511_,
		_w3524_,
		_w3526_,
		_w3564_
	);
	LUT3 #(
		.INIT('h54)
	) name3102 (
		_w1904_,
		_w2086_,
		_w2280_,
		_w3565_
	);
	LUT4 #(
		.INIT('h0010)
	) name3103 (
		_w1509_,
		_w1903_,
		_w2083_,
		_w2282_,
		_w3566_
	);
	LUT2 #(
		.INIT('h1)
	) name3104 (
		_w3565_,
		_w3566_,
		_w3567_
	);
	LUT4 #(
		.INIT('hab00)
	) name3105 (
		_w2192_,
		_w3561_,
		_w3564_,
		_w3567_,
		_w3568_
	);
	LUT4 #(
		.INIT('h0100)
	) name3106 (
		_w3563_,
		_w3562_,
		_w3560_,
		_w3568_,
		_w3569_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name3107 (
		\P1_state_reg[0]/NET0131 ,
		_w1489_,
		_w3559_,
		_w3569_,
		_w3570_
	);
	LUT2 #(
		.INIT('h4)
	) name3108 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[23]/NET0131 ,
		_w3571_
	);
	LUT4 #(
		.INIT('h9c00)
	) name3109 (
		\P2_reg3_reg[22]/NET0131 ,
		\P2_reg3_reg[23]/NET0131 ,
		_w1884_,
		_w2293_,
		_w3572_
	);
	LUT2 #(
		.INIT('h1)
	) name3110 (
		_w3571_,
		_w3572_,
		_w3573_
	);
	LUT2 #(
		.INIT('hb)
	) name3111 (
		_w3570_,
		_w3573_,
		_w3574_
	);
	LUT4 #(
		.INIT('h70d0)
	) name3112 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg0_reg[22]/NET0131 ,
		_w1476_,
		_w3575_
	);
	LUT2 #(
		.INIT('h8)
	) name3113 (
		\P2_reg0_reg[22]/NET0131 ,
		_w1487_,
		_w3576_
	);
	LUT4 #(
		.INIT('haaa8)
	) name3114 (
		\P2_reg0_reg[22]/NET0131 ,
		_w1491_,
		_w1493_,
		_w1496_,
		_w3577_
	);
	LUT3 #(
		.INIT('h10)
	) name3115 (
		_w1509_,
		_w1916_,
		_w2920_,
		_w3578_
	);
	LUT3 #(
		.INIT('ha2)
	) name3116 (
		\P2_reg0_reg[22]/NET0131 ,
		_w2633_,
		_w2634_,
		_w3579_
	);
	LUT2 #(
		.INIT('h1)
	) name3117 (
		_w3578_,
		_w3579_,
		_w3580_
	);
	LUT4 #(
		.INIT('hab00)
	) name3118 (
		_w2276_,
		_w2811_,
		_w3577_,
		_w3580_,
		_w3581_
	);
	LUT4 #(
		.INIT('h0232)
	) name3119 (
		\P2_reg0_reg[22]/NET0131 ,
		_w2192_,
		_w2277_,
		_w2798_,
		_w3582_
	);
	LUT4 #(
		.INIT('h02aa)
	) name3120 (
		\P2_reg0_reg[22]/NET0131 ,
		_w1491_,
		_w1493_,
		_w1496_,
		_w3583_
	);
	LUT3 #(
		.INIT('ha8)
	) name3121 (
		_w2290_,
		_w2808_,
		_w3583_,
		_w3584_
	);
	LUT4 #(
		.INIT('h08c8)
	) name3122 (
		\P2_reg0_reg[22]/NET0131 ,
		_w2081_,
		_w2272_,
		_w2816_,
		_w3585_
	);
	LUT4 #(
		.INIT('h0100)
	) name3123 (
		_w3584_,
		_w3585_,
		_w3582_,
		_w3581_,
		_w3586_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name3124 (
		\P1_state_reg[0]/NET0131 ,
		_w1489_,
		_w3576_,
		_w3586_,
		_w3587_
	);
	LUT2 #(
		.INIT('he)
	) name3125 (
		_w3575_,
		_w3587_,
		_w3588_
	);
	LUT2 #(
		.INIT('h2)
	) name3126 (
		\P1_reg2_reg[16]/NET0131 ,
		_w511_,
		_w3589_
	);
	LUT2 #(
		.INIT('h8)
	) name3127 (
		\P1_reg2_reg[16]/NET0131 ,
		_w524_,
		_w3590_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name3128 (
		\P1_reg2_reg[16]/NET0131 ,
		_w528_,
		_w530_,
		_w533_,
		_w3591_
	);
	LUT4 #(
		.INIT('hddd1)
	) name3129 (
		\P1_reg2_reg[16]/NET0131 ,
		_w534_,
		_w3107_,
		_w3108_,
		_w3592_
	);
	LUT2 #(
		.INIT('h4)
	) name3130 (
		_w786_,
		_w1138_,
		_w3593_
	);
	LUT4 #(
		.INIT('haaa8)
	) name3131 (
		_w534_,
		_w3112_,
		_w3115_,
		_w3593_,
		_w3594_
	);
	LUT4 #(
		.INIT('h2888)
	) name3132 (
		_w534_,
		_w786_,
		_w1120_,
		_w1122_,
		_w3595_
	);
	LUT2 #(
		.INIT('h8)
	) name3133 (
		_w787_,
		_w1143_,
		_w3596_
	);
	LUT3 #(
		.INIT('h0d)
	) name3134 (
		\P1_reg2_reg[16]/NET0131 ,
		_w3350_,
		_w3596_,
		_w3597_
	);
	LUT4 #(
		.INIT('h5700)
	) name3135 (
		_w1136_,
		_w3591_,
		_w3595_,
		_w3597_,
		_w3598_
	);
	LUT4 #(
		.INIT('h0d00)
	) name3136 (
		_w1183_,
		_w3592_,
		_w3594_,
		_w3598_,
		_w3599_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name3137 (
		\P1_state_reg[0]/NET0131 ,
		_w526_,
		_w3590_,
		_w3599_,
		_w3600_
	);
	LUT2 #(
		.INIT('he)
	) name3138 (
		_w3589_,
		_w3600_,
		_w3601_
	);
	LUT2 #(
		.INIT('h4)
	) name3139 (
		_w534_,
		_w1286_,
		_w3602_
	);
	LUT4 #(
		.INIT('h0002)
	) name3140 (
		_w2411_,
		_w2412_,
		_w2951_,
		_w3602_,
		_w3603_
	);
	LUT3 #(
		.INIT('h2a)
	) name3141 (
		\P1_reg2_reg[20]/NET0131 ,
		_w3443_,
		_w3603_,
		_w3604_
	);
	LUT2 #(
		.INIT('h8)
	) name3142 (
		_w703_,
		_w1143_,
		_w3605_
	);
	LUT3 #(
		.INIT('h02)
	) name3143 (
		_w1183_,
		_w3137_,
		_w3138_,
		_w3606_
	);
	LUT3 #(
		.INIT('h10)
	) name3144 (
		_w541_,
		_w701_,
		_w1138_,
		_w3607_
	);
	LUT3 #(
		.INIT('h04)
	) name3145 (
		_w3129_,
		_w3133_,
		_w3607_,
		_w3608_
	);
	LUT4 #(
		.INIT('h1311)
	) name3146 (
		_w534_,
		_w3605_,
		_w3606_,
		_w3608_,
		_w3609_
	);
	LUT3 #(
		.INIT('hce)
	) name3147 (
		_w3443_,
		_w3604_,
		_w3609_,
		_w3610_
	);
	LUT4 #(
		.INIT('h70d0)
	) name3148 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg1_reg[22]/NET0131 ,
		_w1476_,
		_w3611_
	);
	LUT2 #(
		.INIT('h8)
	) name3149 (
		\P2_reg1_reg[22]/NET0131 ,
		_w1487_,
		_w3612_
	);
	LUT4 #(
		.INIT('haa02)
	) name3150 (
		\P2_reg1_reg[22]/NET0131 ,
		_w1491_,
		_w1493_,
		_w1496_,
		_w3613_
	);
	LUT4 #(
		.INIT('h20e0)
	) name3151 (
		\P2_reg1_reg[22]/NET0131 ,
		_w2039_,
		_w2193_,
		_w2798_,
		_w3614_
	);
	LUT3 #(
		.INIT('ha2)
	) name3152 (
		\P2_reg1_reg[22]/NET0131 ,
		_w2633_,
		_w2660_,
		_w3615_
	);
	LUT3 #(
		.INIT('h10)
	) name3153 (
		_w1509_,
		_w1916_,
		_w2963_,
		_w3616_
	);
	LUT2 #(
		.INIT('h1)
	) name3154 (
		_w3615_,
		_w3616_,
		_w3617_
	);
	LUT2 #(
		.INIT('h4)
	) name3155 (
		_w3614_,
		_w3617_,
		_w3618_
	);
	LUT4 #(
		.INIT('h2822)
	) name3156 (
		_w2039_,
		_w2793_,
		_w2805_,
		_w2807_,
		_w3619_
	);
	LUT3 #(
		.INIT('ha8)
	) name3157 (
		_w2038_,
		_w3613_,
		_w3619_,
		_w3620_
	);
	LUT4 #(
		.INIT('h20e0)
	) name3158 (
		\P2_reg1_reg[22]/NET0131 ,
		_w1497_,
		_w2188_,
		_w2798_,
		_w3621_
	);
	LUT4 #(
		.INIT('h20e0)
	) name3159 (
		\P2_reg1_reg[22]/NET0131 ,
		_w1497_,
		_w2081_,
		_w2816_,
		_w3622_
	);
	LUT3 #(
		.INIT('h01)
	) name3160 (
		_w3621_,
		_w3622_,
		_w3620_,
		_w3623_
	);
	LUT4 #(
		.INIT('h3111)
	) name3161 (
		_w1489_,
		_w3612_,
		_w3618_,
		_w3623_,
		_w3624_
	);
	LUT3 #(
		.INIT('hce)
	) name3162 (
		\P1_state_reg[0]/NET0131 ,
		_w3611_,
		_w3624_,
		_w3625_
	);
	LUT2 #(
		.INIT('h2)
	) name3163 (
		\P1_reg0_reg[16]/NET0131 ,
		_w511_,
		_w3626_
	);
	LUT2 #(
		.INIT('h8)
	) name3164 (
		\P1_reg0_reg[16]/NET0131 ,
		_w524_,
		_w3627_
	);
	LUT4 #(
		.INIT('h5554)
	) name3165 (
		\P1_reg0_reg[16]/NET0131 ,
		_w528_,
		_w530_,
		_w533_,
		_w3628_
	);
	LUT2 #(
		.INIT('h2)
	) name3166 (
		_w1183_,
		_w3628_,
		_w3629_
	);
	LUT4 #(
		.INIT('h5700)
	) name3167 (
		_w2688_,
		_w3107_,
		_w3108_,
		_w3629_,
		_w3630_
	);
	LUT4 #(
		.INIT('h6a00)
	) name3168 (
		_w786_,
		_w1120_,
		_w1122_,
		_w1136_,
		_w3631_
	);
	LUT4 #(
		.INIT('h0001)
	) name3169 (
		_w3112_,
		_w3115_,
		_w3593_,
		_w3631_,
		_w3632_
	);
	LUT4 #(
		.INIT('hc4c0)
	) name3170 (
		_w1138_,
		_w2425_,
		_w2688_,
		_w3142_,
		_w3633_
	);
	LUT2 #(
		.INIT('h2)
	) name3171 (
		\P1_reg0_reg[16]/NET0131 ,
		_w3633_,
		_w3634_
	);
	LUT4 #(
		.INIT('h000d)
	) name3172 (
		_w2688_,
		_w3632_,
		_w3634_,
		_w3630_,
		_w3635_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name3173 (
		\P1_state_reg[0]/NET0131 ,
		_w526_,
		_w3627_,
		_w3635_,
		_w3636_
	);
	LUT2 #(
		.INIT('he)
	) name3174 (
		_w3626_,
		_w3636_,
		_w3637_
	);
	LUT2 #(
		.INIT('h2)
	) name3175 (
		\P1_reg0_reg[17]/NET0131 ,
		_w511_,
		_w3638_
	);
	LUT2 #(
		.INIT('h8)
	) name3176 (
		\P1_reg0_reg[17]/NET0131 ,
		_w524_,
		_w3639_
	);
	LUT4 #(
		.INIT('hddd1)
	) name3177 (
		\P1_reg0_reg[17]/NET0131 ,
		_w2688_,
		_w3488_,
		_w3489_,
		_w3640_
	);
	LUT2 #(
		.INIT('h4)
	) name3178 (
		_w717_,
		_w1138_,
		_w3641_
	);
	LUT4 #(
		.INIT('hcc80)
	) name3179 (
		_w1136_,
		_w2688_,
		_w3491_,
		_w3641_,
		_w3642_
	);
	LUT3 #(
		.INIT('ha2)
	) name3180 (
		\P1_reg0_reg[17]/NET0131 ,
		_w2692_,
		_w3005_,
		_w3643_
	);
	LUT2 #(
		.INIT('h1)
	) name3181 (
		_w3642_,
		_w3643_,
		_w3644_
	);
	LUT3 #(
		.INIT('hd0)
	) name3182 (
		_w1183_,
		_w3640_,
		_w3644_,
		_w3645_
	);
	LUT4 #(
		.INIT('hc535)
	) name3183 (
		\P1_reg0_reg[17]/NET0131 ,
		_w1431_,
		_w2688_,
		_w3498_,
		_w3646_
	);
	LUT4 #(
		.INIT('hc808)
	) name3184 (
		\P1_reg0_reg[17]/NET0131 ,
		_w1114_,
		_w2688_,
		_w3500_,
		_w3647_
	);
	LUT3 #(
		.INIT('h0d)
	) name3185 (
		_w1286_,
		_w3646_,
		_w3647_,
		_w3648_
	);
	LUT4 #(
		.INIT('h3111)
	) name3186 (
		_w526_,
		_w3639_,
		_w3645_,
		_w3648_,
		_w3649_
	);
	LUT3 #(
		.INIT('hce)
	) name3187 (
		\P1_state_reg[0]/NET0131 ,
		_w3638_,
		_w3649_,
		_w3650_
	);
	LUT4 #(
		.INIT('h0100)
	) name3188 (
		_w528_,
		_w530_,
		_w533_,
		_w3443_,
		_w3651_
	);
	LUT3 #(
		.INIT('h02)
	) name3189 (
		_w1183_,
		_w3541_,
		_w3542_,
		_w3652_
	);
	LUT3 #(
		.INIT('h10)
	) name3190 (
		_w541_,
		_w1073_,
		_w1138_,
		_w3653_
	);
	LUT3 #(
		.INIT('h07)
	) name3191 (
		_w1136_,
		_w3547_,
		_w3653_,
		_w3654_
	);
	LUT3 #(
		.INIT('h10)
	) name3192 (
		_w3544_,
		_w3545_,
		_w3654_,
		_w3655_
	);
	LUT4 #(
		.INIT('h0103)
	) name3193 (
		_w652_,
		_w1104_,
		_w1106_,
		_w1111_,
		_w3656_
	);
	LUT4 #(
		.INIT('hc2c0)
	) name3194 (
		_w652_,
		_w1104_,
		_w1106_,
		_w1111_,
		_w3657_
	);
	LUT4 #(
		.INIT('ha080)
	) name3195 (
		_w2425_,
		_w2688_,
		_w3443_,
		_w3657_,
		_w3658_
	);
	LUT3 #(
		.INIT('h08)
	) name3196 (
		_w1108_,
		_w1140_,
		_w2688_,
		_w3659_
	);
	LUT3 #(
		.INIT('ha2)
	) name3197 (
		\P1_reg0_reg[21]/NET0131 ,
		_w3658_,
		_w3659_,
		_w3660_
	);
	LUT4 #(
		.INIT('hff8a)
	) name3198 (
		_w3651_,
		_w3652_,
		_w3655_,
		_w3660_,
		_w3661_
	);
	LUT2 #(
		.INIT('h2)
	) name3199 (
		\P1_reg0_reg[24]/NET0131 ,
		_w511_,
		_w3662_
	);
	LUT2 #(
		.INIT('h8)
	) name3200 (
		\P1_reg0_reg[24]/NET0131 ,
		_w524_,
		_w3663_
	);
	LUT3 #(
		.INIT('h01)
	) name3201 (
		_w1107_,
		_w1141_,
		_w2688_,
		_w3664_
	);
	LUT4 #(
		.INIT('haaa2)
	) name3202 (
		\P1_reg0_reg[24]/NET0131 ,
		_w2692_,
		_w3005_,
		_w3664_,
		_w3665_
	);
	LUT3 #(
		.INIT('h28)
	) name3203 (
		_w1286_,
		_w1425_,
		_w2767_,
		_w3666_
	);
	LUT4 #(
		.INIT('h0004)
	) name3204 (
		_w2775_,
		_w2781_,
		_w2948_,
		_w3666_,
		_w3667_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name3205 (
		_w526_,
		_w2688_,
		_w3665_,
		_w3667_,
		_w3668_
	);
	LUT4 #(
		.INIT('heeec)
	) name3206 (
		\P1_state_reg[0]/NET0131 ,
		_w3662_,
		_w3663_,
		_w3668_,
		_w3669_
	);
	LUT2 #(
		.INIT('h2)
	) name3207 (
		\P1_reg0_reg[31]/NET0131 ,
		_w511_,
		_w3670_
	);
	LUT2 #(
		.INIT('h8)
	) name3208 (
		\P1_reg0_reg[31]/NET0131 ,
		_w524_,
		_w3671_
	);
	LUT4 #(
		.INIT('haaa8)
	) name3209 (
		\P1_reg0_reg[31]/NET0131 ,
		_w528_,
		_w530_,
		_w533_,
		_w3672_
	);
	LUT4 #(
		.INIT('h3900)
	) name3210 (
		_w1133_,
		_w1304_,
		_w1312_,
		_w2688_,
		_w3673_
	);
	LUT3 #(
		.INIT('ha8)
	) name3211 (
		_w1136_,
		_w3672_,
		_w3673_,
		_w3674_
	);
	LUT2 #(
		.INIT('h8)
	) name3212 (
		_w1183_,
		_w2688_,
		_w3675_
	);
	LUT4 #(
		.INIT('h1200)
	) name3213 (
		\P2_datao_reg[31]/NET0131 ,
		_w541_,
		_w1303_,
		_w2688_,
		_w3676_
	);
	LUT4 #(
		.INIT('h0a2a)
	) name3214 (
		\P1_reg0_reg[31]/NET0131 ,
		_w1107_,
		_w2425_,
		_w2688_,
		_w3677_
	);
	LUT4 #(
		.INIT('h0057)
	) name3215 (
		_w1138_,
		_w3672_,
		_w3676_,
		_w3677_,
		_w3678_
	);
	LUT3 #(
		.INIT('h70)
	) name3216 (
		_w3286_,
		_w3675_,
		_w3678_,
		_w3679_
	);
	LUT4 #(
		.INIT('h1311)
	) name3217 (
		_w526_,
		_w3671_,
		_w3674_,
		_w3679_,
		_w3680_
	);
	LUT3 #(
		.INIT('hce)
	) name3218 (
		\P1_state_reg[0]/NET0131 ,
		_w3670_,
		_w3680_,
		_w3681_
	);
	LUT2 #(
		.INIT('h2)
	) name3219 (
		\P1_reg1_reg[16]/NET0131 ,
		_w511_,
		_w3682_
	);
	LUT2 #(
		.INIT('h8)
	) name3220 (
		\P1_reg1_reg[16]/NET0131 ,
		_w524_,
		_w3683_
	);
	LUT2 #(
		.INIT('h1)
	) name3221 (
		_w2421_,
		_w3142_,
		_w3684_
	);
	LUT2 #(
		.INIT('h2)
	) name3222 (
		_w1183_,
		_w2421_,
		_w3685_
	);
	LUT3 #(
		.INIT('hdc)
	) name3223 (
		_w1183_,
		_w2421_,
		_w3142_,
		_w3686_
	);
	LUT3 #(
		.INIT('h2a)
	) name3224 (
		\P1_reg1_reg[16]/NET0131 ,
		_w2426_,
		_w3686_,
		_w3687_
	);
	LUT2 #(
		.INIT('h8)
	) name3225 (
		_w1183_,
		_w2421_,
		_w3688_
	);
	LUT4 #(
		.INIT('h0e0f)
	) name3226 (
		_w3107_,
		_w3108_,
		_w3687_,
		_w3688_,
		_w3689_
	);
	LUT4 #(
		.INIT('h08aa)
	) name3227 (
		_w526_,
		_w2421_,
		_w3632_,
		_w3689_,
		_w3690_
	);
	LUT4 #(
		.INIT('heeec)
	) name3228 (
		\P1_state_reg[0]/NET0131 ,
		_w3682_,
		_w3683_,
		_w3690_,
		_w3691_
	);
	LUT2 #(
		.INIT('h2)
	) name3229 (
		\P1_reg1_reg[24]/NET0131 ,
		_w511_,
		_w3692_
	);
	LUT2 #(
		.INIT('h8)
	) name3230 (
		\P1_reg1_reg[24]/NET0131 ,
		_w524_,
		_w3693_
	);
	LUT3 #(
		.INIT('h2a)
	) name3231 (
		\P1_reg1_reg[24]/NET0131 ,
		_w2426_,
		_w3686_,
		_w3694_
	);
	LUT4 #(
		.INIT('haa08)
	) name3232 (
		_w526_,
		_w2421_,
		_w3667_,
		_w3694_,
		_w3695_
	);
	LUT4 #(
		.INIT('heeec)
	) name3233 (
		\P1_state_reg[0]/NET0131 ,
		_w3692_,
		_w3693_,
		_w3695_,
		_w3696_
	);
	LUT2 #(
		.INIT('h2)
	) name3234 (
		\P1_reg1_reg[31]/NET0131 ,
		_w511_,
		_w3697_
	);
	LUT2 #(
		.INIT('h8)
	) name3235 (
		\P1_reg1_reg[31]/NET0131 ,
		_w524_,
		_w3698_
	);
	LUT4 #(
		.INIT('haa02)
	) name3236 (
		\P1_reg1_reg[31]/NET0131 ,
		_w528_,
		_w530_,
		_w533_,
		_w3699_
	);
	LUT4 #(
		.INIT('h3900)
	) name3237 (
		_w1133_,
		_w1304_,
		_w1312_,
		_w2421_,
		_w3700_
	);
	LUT3 #(
		.INIT('ha8)
	) name3238 (
		_w1136_,
		_w3699_,
		_w3700_,
		_w3701_
	);
	LUT4 #(
		.INIT('h1200)
	) name3239 (
		\P2_datao_reg[31]/NET0131 ,
		_w541_,
		_w1303_,
		_w2421_,
		_w3702_
	);
	LUT4 #(
		.INIT('h02aa)
	) name3240 (
		\P1_reg1_reg[31]/NET0131 ,
		_w1107_,
		_w2421_,
		_w2425_,
		_w3703_
	);
	LUT4 #(
		.INIT('h0057)
	) name3241 (
		_w1138_,
		_w3699_,
		_w3702_,
		_w3703_,
		_w3704_
	);
	LUT3 #(
		.INIT('h70)
	) name3242 (
		_w3286_,
		_w3688_,
		_w3704_,
		_w3705_
	);
	LUT4 #(
		.INIT('h1311)
	) name3243 (
		_w526_,
		_w3698_,
		_w3701_,
		_w3705_,
		_w3706_
	);
	LUT3 #(
		.INIT('hce)
	) name3244 (
		\P1_state_reg[0]/NET0131 ,
		_w3697_,
		_w3706_,
		_w3707_
	);
	LUT2 #(
		.INIT('h8)
	) name3245 (
		_w524_,
		_w675_,
		_w3708_
	);
	LUT4 #(
		.INIT('h1f00)
	) name3246 (
		_w528_,
		_w530_,
		_w533_,
		_w675_,
		_w3709_
	);
	LUT4 #(
		.INIT('h9555)
	) name3247 (
		_w706_,
		_w1165_,
		_w1161_,
		_w1163_,
		_w3710_
	);
	LUT4 #(
		.INIT('h7020)
	) name3248 (
		_w537_,
		_w745_,
		_w2197_,
		_w3710_,
		_w3711_
	);
	LUT3 #(
		.INIT('ha8)
	) name3249 (
		_w1183_,
		_w3709_,
		_w3711_,
		_w3712_
	);
	LUT4 #(
		.INIT('h00b7)
	) name3250 (
		_w1422_,
		_w2197_,
		_w2848_,
		_w3709_,
		_w3713_
	);
	LUT2 #(
		.INIT('h2)
	) name3251 (
		_w1286_,
		_w3713_,
		_w3714_
	);
	LUT4 #(
		.INIT('h007b)
	) name3252 (
		_w1422_,
		_w2197_,
		_w2876_,
		_w3709_,
		_w3715_
	);
	LUT4 #(
		.INIT('h007b)
	) name3253 (
		_w674_,
		_w2197_,
		_w3130_,
		_w3709_,
		_w3716_
	);
	LUT4 #(
		.INIT('h8d00)
	) name3254 (
		_w541_,
		_w652_,
		_w673_,
		_w1138_,
		_w3717_
	);
	LUT3 #(
		.INIT('hb0)
	) name3255 (
		_w541_,
		_w673_,
		_w1143_,
		_w3718_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name3256 (
		_w675_,
		_w1138_,
		_w1141_,
		_w2197_,
		_w3719_
	);
	LUT4 #(
		.INIT('h0013)
	) name3257 (
		_w2197_,
		_w3718_,
		_w3717_,
		_w3719_,
		_w3720_
	);
	LUT3 #(
		.INIT('hd0)
	) name3258 (
		_w1136_,
		_w3716_,
		_w3720_,
		_w3721_
	);
	LUT3 #(
		.INIT('hd0)
	) name3259 (
		_w1114_,
		_w3715_,
		_w3721_,
		_w3722_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name3260 (
		_w526_,
		_w3712_,
		_w3714_,
		_w3722_,
		_w3723_
	);
	LUT2 #(
		.INIT('h2)
	) name3261 (
		\P1_reg3_reg[19]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w3724_
	);
	LUT4 #(
		.INIT('h9d5d)
	) name3262 (
		\P1_reg3_reg[19]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w510_,
		_w634_,
		_w3725_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name3263 (
		\P1_state_reg[0]/NET0131 ,
		_w3708_,
		_w3723_,
		_w3725_,
		_w3726_
	);
	LUT2 #(
		.INIT('h8)
	) name3264 (
		_w524_,
		_w901_,
		_w3727_
	);
	LUT4 #(
		.INIT('h0100)
	) name3265 (
		_w903_,
		_w912_,
		_w924_,
		_w1154_,
		_w3728_
	);
	LUT3 #(
		.INIT('h80)
	) name3266 (
		_w537_,
		_w909_,
		_w911_,
		_w3729_
	);
	LUT4 #(
		.INIT('h00eb)
	) name3267 (
		_w537_,
		_w833_,
		_w3728_,
		_w3729_,
		_w3730_
	);
	LUT4 #(
		.INIT('hc808)
	) name3268 (
		_w901_,
		_w1183_,
		_w2197_,
		_w3730_,
		_w3731_
	);
	LUT4 #(
		.INIT('h208a)
	) name3269 (
		_w1286_,
		_w1365_,
		_w1368_,
		_w1451_,
		_w3732_
	);
	LUT4 #(
		.INIT('h8288)
	) name3270 (
		_w1114_,
		_w1451_,
		_w2224_,
		_w2227_,
		_w3733_
	);
	LUT4 #(
		.INIT('h8000)
	) name3271 (
		_w894_,
		_w907_,
		_w1115_,
		_w1116_,
		_w3734_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name3272 (
		_w894_,
		_w907_,
		_w1115_,
		_w1116_,
		_w3735_
	);
	LUT4 #(
		.INIT('hc808)
	) name3273 (
		_w901_,
		_w1136_,
		_w2197_,
		_w3735_,
		_w3736_
	);
	LUT4 #(
		.INIT('h888a)
	) name3274 (
		_w901_,
		_w1141_,
		_w2197_,
		_w3118_,
		_w3737_
	);
	LUT3 #(
		.INIT('h04)
	) name3275 (
		_w907_,
		_w2259_,
		_w2260_,
		_w3738_
	);
	LUT2 #(
		.INIT('h1)
	) name3276 (
		_w3737_,
		_w3738_,
		_w3739_
	);
	LUT2 #(
		.INIT('h4)
	) name3277 (
		_w3736_,
		_w3739_,
		_w3740_
	);
	LUT4 #(
		.INIT('h5700)
	) name3278 (
		_w2197_,
		_w3732_,
		_w3733_,
		_w3740_,
		_w3741_
	);
	LUT4 #(
		.INIT('h1311)
	) name3279 (
		_w526_,
		_w3727_,
		_w3731_,
		_w3741_,
		_w3742_
	);
	LUT2 #(
		.INIT('h2)
	) name3280 (
		\P1_reg3_reg[8]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w3743_
	);
	LUT3 #(
		.INIT('h07)
	) name3281 (
		_w901_,
		_w1294_,
		_w3743_,
		_w3744_
	);
	LUT3 #(
		.INIT('h2f)
	) name3282 (
		\P1_state_reg[0]/NET0131 ,
		_w3742_,
		_w3744_,
		_w3745_
	);
	LUT2 #(
		.INIT('h8)
	) name3283 (
		_w524_,
		_w1048_,
		_w3746_
	);
	LUT2 #(
		.INIT('h8)
	) name3284 (
		_w2866_,
		_w2878_,
		_w3747_
	);
	LUT4 #(
		.INIT('h4f00)
	) name3285 (
		_w2871_,
		_w2872_,
		_w2873_,
		_w3747_,
		_w3748_
	);
	LUT3 #(
		.INIT('hd0)
	) name3286 (
		_w960_,
		_w2874_,
		_w2878_,
		_w3749_
	);
	LUT2 #(
		.INIT('h2)
	) name3287 (
		_w2880_,
		_w3749_,
		_w3750_
	);
	LUT4 #(
		.INIT('h2822)
	) name3288 (
		_w1114_,
		_w1426_,
		_w3748_,
		_w3750_,
		_w3751_
	);
	LUT3 #(
		.INIT('h8a)
	) name3289 (
		_w1047_,
		_w1066_,
		_w3546_,
		_w3752_
	);
	LUT2 #(
		.INIT('h4)
	) name3290 (
		_w1128_,
		_w1136_,
		_w3753_
	);
	LUT2 #(
		.INIT('h4)
	) name3291 (
		_w3752_,
		_w3753_,
		_w3754_
	);
	LUT3 #(
		.INIT('h80)
	) name3292 (
		_w1169_,
		_w1161_,
		_w1163_,
		_w3755_
	);
	LUT4 #(
		.INIT('h9555)
	) name3293 (
		_w1059_,
		_w1169_,
		_w1161_,
		_w1163_,
		_w3756_
	);
	LUT4 #(
		.INIT('h7020)
	) name3294 (
		_w537_,
		_w1070_,
		_w1183_,
		_w3756_,
		_w3757_
	);
	LUT2 #(
		.INIT('h8)
	) name3295 (
		_w2840_,
		_w2849_,
		_w3758_
	);
	LUT4 #(
		.INIT('h4f00)
	) name3296 (
		_w2843_,
		_w2844_,
		_w2845_,
		_w3758_,
		_w3759_
	);
	LUT3 #(
		.INIT('he0)
	) name3297 (
		_w1246_,
		_w2846_,
		_w2849_,
		_w3760_
	);
	LUT2 #(
		.INIT('h2)
	) name3298 (
		_w2853_,
		_w3760_,
		_w3761_
	);
	LUT4 #(
		.INIT('h8288)
	) name3299 (
		_w1286_,
		_w1426_,
		_w3759_,
		_w3761_,
		_w3762_
	);
	LUT4 #(
		.INIT('h0001)
	) name3300 (
		_w3751_,
		_w3754_,
		_w3757_,
		_w3762_,
		_w3763_
	);
	LUT3 #(
		.INIT('h10)
	) name3301 (
		_w541_,
		_w1046_,
		_w2261_,
		_w3764_
	);
	LUT4 #(
		.INIT('h3130)
	) name3302 (
		_w1138_,
		_w1141_,
		_w2197_,
		_w2259_,
		_w3765_
	);
	LUT2 #(
		.INIT('h2)
	) name3303 (
		_w1048_,
		_w3765_,
		_w3766_
	);
	LUT2 #(
		.INIT('h1)
	) name3304 (
		_w3764_,
		_w3766_,
		_w3767_
	);
	LUT4 #(
		.INIT('h08aa)
	) name3305 (
		_w526_,
		_w2197_,
		_w3763_,
		_w3767_,
		_w3768_
	);
	LUT2 #(
		.INIT('h2)
	) name3306 (
		\P1_reg3_reg[23]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w3769_
	);
	LUT4 #(
		.INIT('h6a00)
	) name3307 (
		\P1_reg3_reg[23]/NET0131 ,
		_w634_,
		_w636_,
		_w1294_,
		_w3770_
	);
	LUT2 #(
		.INIT('h1)
	) name3308 (
		_w3769_,
		_w3770_,
		_w3771_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name3309 (
		\P1_state_reg[0]/NET0131 ,
		_w3746_,
		_w3768_,
		_w3771_,
		_w3772_
	);
	LUT2 #(
		.INIT('h8)
	) name3310 (
		_w524_,
		_w1067_,
		_w3773_
	);
	LUT4 #(
		.INIT('h1f00)
	) name3311 (
		_w528_,
		_w530_,
		_w533_,
		_w1067_,
		_w3774_
	);
	LUT4 #(
		.INIT('h5504)
	) name3312 (
		_w537_,
		_w1051_,
		_w3540_,
		_w3755_,
		_w3775_
	);
	LUT2 #(
		.INIT('h8)
	) name3313 (
		_w537_,
		_w1078_,
		_w3776_
	);
	LUT4 #(
		.INIT('h3331)
	) name3314 (
		_w2197_,
		_w3774_,
		_w3775_,
		_w3776_,
		_w3777_
	);
	LUT4 #(
		.INIT('h7500)
	) name3315 (
		_w3045_,
		_w3052_,
		_w3053_,
		_w3054_,
		_w3778_
	);
	LUT3 #(
		.INIT('h08)
	) name3316 (
		_w2209_,
		_w2244_,
		_w3046_,
		_w3779_
	);
	LUT2 #(
		.INIT('h2)
	) name3317 (
		_w3042_,
		_w3779_,
		_w3780_
	);
	LUT4 #(
		.INIT('h4844)
	) name3318 (
		_w1457_,
		_w2197_,
		_w3778_,
		_w3780_,
		_w3781_
	);
	LUT3 #(
		.INIT('ha8)
	) name3319 (
		_w1114_,
		_w3774_,
		_w3781_,
		_w3782_
	);
	LUT4 #(
		.INIT('h20aa)
	) name3320 (
		_w3072_,
		_w3076_,
		_w3077_,
		_w3079_,
		_w3783_
	);
	LUT3 #(
		.INIT('h08)
	) name3321 (
		_w1328_,
		_w1334_,
		_w3080_,
		_w3784_
	);
	LUT2 #(
		.INIT('h2)
	) name3322 (
		_w3069_,
		_w3784_,
		_w3785_
	);
	LUT4 #(
		.INIT('h8488)
	) name3323 (
		_w1457_,
		_w2197_,
		_w3783_,
		_w3785_,
		_w3786_
	);
	LUT4 #(
		.INIT('h8040)
	) name3324 (
		_w1066_,
		_w1136_,
		_w2197_,
		_w3546_,
		_w3787_
	);
	LUT4 #(
		.INIT('h5f13)
	) name3325 (
		_w1066_,
		_w1067_,
		_w2261_,
		_w2860_,
		_w3788_
	);
	LUT2 #(
		.INIT('h4)
	) name3326 (
		_w3787_,
		_w3788_,
		_w3789_
	);
	LUT4 #(
		.INIT('h5700)
	) name3327 (
		_w1286_,
		_w3774_,
		_w3786_,
		_w3789_,
		_w3790_
	);
	LUT4 #(
		.INIT('h0d00)
	) name3328 (
		_w1183_,
		_w3777_,
		_w3782_,
		_w3790_,
		_w3791_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name3329 (
		\P1_state_reg[0]/NET0131 ,
		_w526_,
		_w3773_,
		_w3791_,
		_w3792_
	);
	LUT2 #(
		.INIT('h2)
	) name3330 (
		\P1_reg3_reg[22]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w3793_
	);
	LUT3 #(
		.INIT('h07)
	) name3331 (
		_w1067_,
		_w1294_,
		_w3793_,
		_w3794_
	);
	LUT2 #(
		.INIT('hb)
	) name3332 (
		_w3792_,
		_w3794_,
		_w3795_
	);
	LUT2 #(
		.INIT('h2)
	) name3333 (
		_w1487_,
		_w1885_,
		_w3796_
	);
	LUT4 #(
		.INIT('h00fe)
	) name3334 (
		_w1491_,
		_w1493_,
		_w1496_,
		_w1885_,
		_w3797_
	);
	LUT4 #(
		.INIT('h208a)
	) name3335 (
		_w2277_,
		_w2640_,
		_w2642_,
		_w3212_,
		_w3798_
	);
	LUT3 #(
		.INIT('ha8)
	) name3336 (
		_w2290_,
		_w3797_,
		_w3798_,
		_w3799_
	);
	LUT4 #(
		.INIT('h001f)
	) name3337 (
		_w1491_,
		_w1493_,
		_w1496_,
		_w1885_,
		_w3800_
	);
	LUT4 #(
		.INIT('h8a20)
	) name3338 (
		_w2272_,
		_w2621_,
		_w2623_,
		_w3212_,
		_w3801_
	);
	LUT4 #(
		.INIT('h0010)
	) name3339 (
		_w1509_,
		_w1882_,
		_w2083_,
		_w2282_,
		_w3802_
	);
	LUT3 #(
		.INIT('h54)
	) name3340 (
		_w1885_,
		_w2086_,
		_w2280_,
		_w3803_
	);
	LUT2 #(
		.INIT('h1)
	) name3341 (
		_w3802_,
		_w3803_,
		_w3804_
	);
	LUT4 #(
		.INIT('hab00)
	) name3342 (
		_w2192_,
		_w3800_,
		_w3801_,
		_w3804_,
		_w3805_
	);
	LUT4 #(
		.INIT('h0057)
	) name3343 (
		_w2277_,
		_w3222_,
		_w3223_,
		_w3797_,
		_w3806_
	);
	LUT2 #(
		.INIT('h2)
	) name3344 (
		_w2081_,
		_w3806_,
		_w3807_
	);
	LUT4 #(
		.INIT('h208a)
	) name3345 (
		_w2272_,
		_w2640_,
		_w2642_,
		_w3212_,
		_w3808_
	);
	LUT3 #(
		.INIT('h54)
	) name3346 (
		_w2276_,
		_w3800_,
		_w3808_,
		_w3809_
	);
	LUT4 #(
		.INIT('h0100)
	) name3347 (
		_w3799_,
		_w3807_,
		_w3809_,
		_w3805_,
		_w3810_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name3348 (
		\P1_state_reg[0]/NET0131 ,
		_w1489_,
		_w3796_,
		_w3810_,
		_w3811_
	);
	LUT2 #(
		.INIT('h4)
	) name3349 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[21]/NET0131 ,
		_w3812_
	);
	LUT3 #(
		.INIT('h0b)
	) name3350 (
		_w1885_,
		_w2293_,
		_w3812_,
		_w3813_
	);
	LUT2 #(
		.INIT('hb)
	) name3351 (
		_w3811_,
		_w3813_,
		_w3814_
	);
	LUT4 #(
		.INIT('h70d0)
	) name3352 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg0_reg[17]/NET0131 ,
		_w1476_,
		_w3815_
	);
	LUT2 #(
		.INIT('h8)
	) name3353 (
		\P2_reg0_reg[17]/NET0131 ,
		_w1487_,
		_w3816_
	);
	LUT4 #(
		.INIT('h1dd1)
	) name3354 (
		\P2_reg0_reg[17]/NET0131 ,
		_w2277_,
		_w2705_,
		_w2706_,
		_w3817_
	);
	LUT2 #(
		.INIT('h1)
	) name3355 (
		_w2276_,
		_w3817_,
		_w3818_
	);
	LUT4 #(
		.INIT('h02aa)
	) name3356 (
		\P2_reg0_reg[17]/NET0131 ,
		_w1491_,
		_w1493_,
		_w1496_,
		_w3819_
	);
	LUT4 #(
		.INIT('h1dd1)
	) name3357 (
		\P2_reg0_reg[17]/NET0131 ,
		_w2272_,
		_w2705_,
		_w2706_,
		_w3820_
	);
	LUT2 #(
		.INIT('h2)
	) name3358 (
		_w2290_,
		_w3820_,
		_w3821_
	);
	LUT4 #(
		.INIT('hd11d)
	) name3359 (
		\P2_reg0_reg[17]/NET0131 ,
		_w2277_,
		_w2705_,
		_w2712_,
		_w3822_
	);
	LUT4 #(
		.INIT('h8a88)
	) name3360 (
		_w2272_,
		_w2714_,
		_w2715_,
		_w2716_,
		_w3823_
	);
	LUT3 #(
		.INIT('ha2)
	) name3361 (
		\P2_reg0_reg[17]/NET0131 ,
		_w2633_,
		_w2634_,
		_w3824_
	);
	LUT4 #(
		.INIT('hf100)
	) name3362 (
		_w1509_,
		_w1771_,
		_w1775_,
		_w2920_,
		_w3825_
	);
	LUT2 #(
		.INIT('h1)
	) name3363 (
		_w3824_,
		_w3825_,
		_w3826_
	);
	LUT4 #(
		.INIT('h5700)
	) name3364 (
		_w2081_,
		_w3819_,
		_w3823_,
		_w3826_,
		_w3827_
	);
	LUT3 #(
		.INIT('he0)
	) name3365 (
		_w2192_,
		_w3822_,
		_w3827_,
		_w3828_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name3366 (
		_w1489_,
		_w3821_,
		_w3818_,
		_w3828_,
		_w3829_
	);
	LUT4 #(
		.INIT('heeec)
	) name3367 (
		\P1_state_reg[0]/NET0131 ,
		_w3815_,
		_w3816_,
		_w3829_,
		_w3830_
	);
	LUT4 #(
		.INIT('h70d0)
	) name3368 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg0_reg[18]/NET0131 ,
		_w1476_,
		_w3831_
	);
	LUT2 #(
		.INIT('h8)
	) name3369 (
		\P2_reg0_reg[18]/NET0131 ,
		_w1487_,
		_w3832_
	);
	LUT4 #(
		.INIT('haaa8)
	) name3370 (
		\P2_reg0_reg[18]/NET0131 ,
		_w1491_,
		_w1493_,
		_w1496_,
		_w3833_
	);
	LUT4 #(
		.INIT('h1dd1)
	) name3371 (
		\P2_reg0_reg[18]/NET0131 ,
		_w2277_,
		_w2472_,
		_w2728_,
		_w3834_
	);
	LUT4 #(
		.INIT('h08c8)
	) name3372 (
		\P2_reg0_reg[18]/NET0131 ,
		_w2081_,
		_w2272_,
		_w2732_,
		_w3835_
	);
	LUT2 #(
		.INIT('h4)
	) name3373 (
		_w1833_,
		_w2920_,
		_w3836_
	);
	LUT3 #(
		.INIT('ha2)
	) name3374 (
		\P2_reg0_reg[18]/NET0131 ,
		_w2633_,
		_w2634_,
		_w3837_
	);
	LUT2 #(
		.INIT('h1)
	) name3375 (
		_w3836_,
		_w3837_,
		_w3838_
	);
	LUT4 #(
		.INIT('h0e00)
	) name3376 (
		_w2276_,
		_w3834_,
		_w3835_,
		_w3838_,
		_w3839_
	);
	LUT4 #(
		.INIT('h8a20)
	) name3377 (
		_w2277_,
		_w2495_,
		_w2498_,
		_w2728_,
		_w3840_
	);
	LUT3 #(
		.INIT('h54)
	) name3378 (
		_w2192_,
		_w3833_,
		_w3840_,
		_w3841_
	);
	LUT4 #(
		.INIT('h1dd1)
	) name3379 (
		\P2_reg0_reg[18]/NET0131 ,
		_w2272_,
		_w2472_,
		_w2728_,
		_w3842_
	);
	LUT2 #(
		.INIT('h2)
	) name3380 (
		_w2290_,
		_w3842_,
		_w3843_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name3381 (
		_w1489_,
		_w3841_,
		_w3843_,
		_w3839_,
		_w3844_
	);
	LUT4 #(
		.INIT('heeec)
	) name3382 (
		\P1_state_reg[0]/NET0131 ,
		_w3831_,
		_w3832_,
		_w3844_,
		_w3845_
	);
	LUT4 #(
		.INIT('h70d0)
	) name3383 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg0_reg[19]/NET0131 ,
		_w1476_,
		_w3846_
	);
	LUT2 #(
		.INIT('h8)
	) name3384 (
		\P2_reg0_reg[19]/NET0131 ,
		_w1487_,
		_w3847_
	);
	LUT4 #(
		.INIT('haaa8)
	) name3385 (
		\P2_reg0_reg[19]/NET0131 ,
		_w1491_,
		_w1493_,
		_w1496_,
		_w3848_
	);
	LUT3 #(
		.INIT('h54)
	) name3386 (
		_w2276_,
		_w2753_,
		_w3848_,
		_w3849_
	);
	LUT4 #(
		.INIT('h02aa)
	) name3387 (
		\P2_reg0_reg[19]/NET0131 ,
		_w1491_,
		_w1493_,
		_w1496_,
		_w3850_
	);
	LUT3 #(
		.INIT('ha8)
	) name3388 (
		_w2290_,
		_w2750_,
		_w3850_,
		_w3851_
	);
	LUT4 #(
		.INIT('h08c8)
	) name3389 (
		\P2_reg0_reg[19]/NET0131 ,
		_w2081_,
		_w2272_,
		_w2756_,
		_w3852_
	);
	LUT4 #(
		.INIT('hd11d)
	) name3390 (
		\P2_reg0_reg[19]/NET0131 ,
		_w2277_,
		_w2378_,
		_w2749_,
		_w3853_
	);
	LUT3 #(
		.INIT('ha2)
	) name3391 (
		\P2_reg0_reg[19]/NET0131 ,
		_w2633_,
		_w2634_,
		_w3854_
	);
	LUT2 #(
		.INIT('h4)
	) name3392 (
		_w1813_,
		_w2920_,
		_w3855_
	);
	LUT2 #(
		.INIT('h1)
	) name3393 (
		_w3854_,
		_w3855_,
		_w3856_
	);
	LUT4 #(
		.INIT('h3200)
	) name3394 (
		_w2192_,
		_w3852_,
		_w3853_,
		_w3856_,
		_w3857_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name3395 (
		_w1489_,
		_w3851_,
		_w3849_,
		_w3857_,
		_w3858_
	);
	LUT4 #(
		.INIT('heeec)
	) name3396 (
		\P1_state_reg[0]/NET0131 ,
		_w3846_,
		_w3847_,
		_w3858_,
		_w3859_
	);
	LUT4 #(
		.INIT('h70d0)
	) name3397 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg0_reg[20]/NET0131 ,
		_w1476_,
		_w3860_
	);
	LUT2 #(
		.INIT('h8)
	) name3398 (
		\P2_reg0_reg[20]/NET0131 ,
		_w1487_,
		_w3861_
	);
	LUT4 #(
		.INIT('haaa8)
	) name3399 (
		\P2_reg0_reg[20]/NET0131 ,
		_w1491_,
		_w1493_,
		_w1496_,
		_w3862_
	);
	LUT4 #(
		.INIT('h35c5)
	) name3400 (
		\P2_reg0_reg[20]/NET0131 ,
		_w1857_,
		_w2277_,
		_w3190_,
		_w3863_
	);
	LUT2 #(
		.INIT('h1)
	) name3401 (
		_w2276_,
		_w3863_,
		_w3864_
	);
	LUT4 #(
		.INIT('h111d)
	) name3402 (
		\P2_reg0_reg[20]/NET0131 ,
		_w2272_,
		_w3194_,
		_w3195_,
		_w3865_
	);
	LUT3 #(
		.INIT('ha2)
	) name3403 (
		\P2_reg0_reg[20]/NET0131 ,
		_w2633_,
		_w2634_,
		_w3866_
	);
	LUT4 #(
		.INIT('h5400)
	) name3404 (
		_w1509_,
		_w1858_,
		_w1865_,
		_w2920_,
		_w3867_
	);
	LUT2 #(
		.INIT('h1)
	) name3405 (
		_w3866_,
		_w3867_,
		_w3868_
	);
	LUT3 #(
		.INIT('hd0)
	) name3406 (
		_w2081_,
		_w3865_,
		_w3868_,
		_w3869_
	);
	LUT4 #(
		.INIT('hb040)
	) name3407 (
		_w2138_,
		_w2155_,
		_w2277_,
		_w3190_,
		_w3870_
	);
	LUT3 #(
		.INIT('h54)
	) name3408 (
		_w2192_,
		_w3862_,
		_w3870_,
		_w3871_
	);
	LUT4 #(
		.INIT('h35c5)
	) name3409 (
		\P2_reg0_reg[20]/NET0131 ,
		_w1857_,
		_w2272_,
		_w3190_,
		_w3872_
	);
	LUT2 #(
		.INIT('h2)
	) name3410 (
		_w2290_,
		_w3872_,
		_w3873_
	);
	LUT4 #(
		.INIT('h0100)
	) name3411 (
		_w3864_,
		_w3871_,
		_w3873_,
		_w3869_,
		_w3874_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name3412 (
		\P1_state_reg[0]/NET0131 ,
		_w1489_,
		_w3861_,
		_w3874_,
		_w3875_
	);
	LUT2 #(
		.INIT('he)
	) name3413 (
		_w3860_,
		_w3875_,
		_w3876_
	);
	LUT4 #(
		.INIT('h70d0)
	) name3414 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg0_reg[21]/NET0131 ,
		_w1476_,
		_w3877_
	);
	LUT2 #(
		.INIT('h8)
	) name3415 (
		\P2_reg0_reg[21]/NET0131 ,
		_w1487_,
		_w3878_
	);
	LUT4 #(
		.INIT('h02aa)
	) name3416 (
		\P2_reg0_reg[21]/NET0131 ,
		_w1491_,
		_w1493_,
		_w1496_,
		_w3879_
	);
	LUT3 #(
		.INIT('ha8)
	) name3417 (
		_w2290_,
		_w3808_,
		_w3879_,
		_w3880_
	);
	LUT4 #(
		.INIT('haaa8)
	) name3418 (
		\P2_reg0_reg[21]/NET0131 ,
		_w1491_,
		_w1493_,
		_w1496_,
		_w3881_
	);
	LUT4 #(
		.INIT('h8a20)
	) name3419 (
		_w2277_,
		_w2621_,
		_w2623_,
		_w3212_,
		_w3882_
	);
	LUT3 #(
		.INIT('ha2)
	) name3420 (
		\P2_reg0_reg[21]/NET0131 ,
		_w2633_,
		_w2634_,
		_w3883_
	);
	LUT4 #(
		.INIT('h1000)
	) name3421 (
		_w1509_,
		_w1882_,
		_w2084_,
		_w2277_,
		_w3884_
	);
	LUT2 #(
		.INIT('h1)
	) name3422 (
		_w3883_,
		_w3884_,
		_w3885_
	);
	LUT4 #(
		.INIT('hab00)
	) name3423 (
		_w2192_,
		_w3881_,
		_w3882_,
		_w3885_,
		_w3886_
	);
	LUT4 #(
		.INIT('h111d)
	) name3424 (
		\P2_reg0_reg[21]/NET0131 ,
		_w2272_,
		_w3222_,
		_w3223_,
		_w3887_
	);
	LUT2 #(
		.INIT('h2)
	) name3425 (
		_w2081_,
		_w3887_,
		_w3888_
	);
	LUT3 #(
		.INIT('h54)
	) name3426 (
		_w2276_,
		_w3798_,
		_w3881_,
		_w3889_
	);
	LUT4 #(
		.INIT('h0100)
	) name3427 (
		_w3880_,
		_w3888_,
		_w3889_,
		_w3886_,
		_w3890_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name3428 (
		\P1_state_reg[0]/NET0131 ,
		_w1489_,
		_w3878_,
		_w3890_,
		_w3891_
	);
	LUT2 #(
		.INIT('he)
	) name3429 (
		_w3877_,
		_w3891_,
		_w3892_
	);
	LUT2 #(
		.INIT('h2)
	) name3430 (
		\P1_reg2_reg[18]/NET0131 ,
		_w511_,
		_w3893_
	);
	LUT2 #(
		.INIT('h8)
	) name3431 (
		\P1_reg2_reg[18]/NET0131 ,
		_w524_,
		_w3894_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name3432 (
		\P1_reg2_reg[18]/NET0131 ,
		_w528_,
		_w530_,
		_w533_,
		_w3895_
	);
	LUT4 #(
		.INIT('h2282)
	) name3433 (
		_w534_,
		_w1423_,
		_w3080_,
		_w3469_,
		_w3896_
	);
	LUT4 #(
		.INIT('h60c0)
	) name3434 (
		_w717_,
		_w738_,
		_w1136_,
		_w3116_,
		_w3897_
	);
	LUT4 #(
		.INIT('hb100)
	) name3435 (
		_w541_,
		_w735_,
		_w736_,
		_w1138_,
		_w3898_
	);
	LUT2 #(
		.INIT('h8)
	) name3436 (
		_w740_,
		_w1143_,
		_w3899_
	);
	LUT3 #(
		.INIT('h0d)
	) name3437 (
		\P1_reg2_reg[18]/NET0131 ,
		_w2411_,
		_w3899_,
		_w3900_
	);
	LUT4 #(
		.INIT('h5700)
	) name3438 (
		_w534_,
		_w3897_,
		_w3898_,
		_w3900_,
		_w3901_
	);
	LUT4 #(
		.INIT('h5700)
	) name3439 (
		_w1286_,
		_w3895_,
		_w3896_,
		_w3901_,
		_w3902_
	);
	LUT4 #(
		.INIT('h8828)
	) name3440 (
		_w534_,
		_w1423_,
		_w3046_,
		_w3476_,
		_w3903_
	);
	LUT3 #(
		.INIT('ha8)
	) name3441 (
		_w1114_,
		_w3895_,
		_w3903_,
		_w3904_
	);
	LUT4 #(
		.INIT('h2a08)
	) name3442 (
		_w534_,
		_w537_,
		_w722_,
		_w3479_,
		_w3905_
	);
	LUT3 #(
		.INIT('ha8)
	) name3443 (
		_w1183_,
		_w3895_,
		_w3905_,
		_w3906_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name3444 (
		_w526_,
		_w3904_,
		_w3906_,
		_w3902_,
		_w3907_
	);
	LUT4 #(
		.INIT('heeec)
	) name3445 (
		\P1_state_reg[0]/NET0131 ,
		_w3893_,
		_w3894_,
		_w3907_,
		_w3908_
	);
	LUT2 #(
		.INIT('h2)
	) name3446 (
		\P1_reg2_reg[19]/NET0131 ,
		_w511_,
		_w3909_
	);
	LUT2 #(
		.INIT('h8)
	) name3447 (
		\P1_reg2_reg[19]/NET0131 ,
		_w524_,
		_w3910_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name3448 (
		\P1_reg2_reg[19]/NET0131 ,
		_w528_,
		_w530_,
		_w533_,
		_w3911_
	);
	LUT4 #(
		.INIT('h2a08)
	) name3449 (
		_w534_,
		_w537_,
		_w745_,
		_w3710_,
		_w3912_
	);
	LUT3 #(
		.INIT('ha8)
	) name3450 (
		_w1183_,
		_w3911_,
		_w3912_,
		_w3913_
	);
	LUT4 #(
		.INIT('hd11d)
	) name3451 (
		\P1_reg2_reg[19]/NET0131 ,
		_w534_,
		_w1422_,
		_w2848_,
		_w3914_
	);
	LUT2 #(
		.INIT('h2)
	) name3452 (
		_w1286_,
		_w3914_,
		_w3915_
	);
	LUT4 #(
		.INIT('h1dd1)
	) name3453 (
		\P1_reg2_reg[19]/NET0131 ,
		_w534_,
		_w1422_,
		_w2876_,
		_w3916_
	);
	LUT4 #(
		.INIT('h1dd1)
	) name3454 (
		\P1_reg2_reg[19]/NET0131 ,
		_w534_,
		_w674_,
		_w3130_,
		_w3917_
	);
	LUT2 #(
		.INIT('h8)
	) name3455 (
		_w675_,
		_w1143_,
		_w3918_
	);
	LUT4 #(
		.INIT('haa20)
	) name3456 (
		\P1_reg2_reg[19]/NET0131 ,
		_w534_,
		_w1138_,
		_w1141_,
		_w3919_
	);
	LUT4 #(
		.INIT('h0007)
	) name3457 (
		_w534_,
		_w3717_,
		_w3918_,
		_w3919_,
		_w3920_
	);
	LUT3 #(
		.INIT('hd0)
	) name3458 (
		_w1136_,
		_w3917_,
		_w3920_,
		_w3921_
	);
	LUT3 #(
		.INIT('hd0)
	) name3459 (
		_w1114_,
		_w3916_,
		_w3921_,
		_w3922_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name3460 (
		_w526_,
		_w3913_,
		_w3915_,
		_w3922_,
		_w3923_
	);
	LUT4 #(
		.INIT('heeec)
	) name3461 (
		\P1_state_reg[0]/NET0131 ,
		_w3909_,
		_w3910_,
		_w3923_,
		_w3924_
	);
	LUT2 #(
		.INIT('h2)
	) name3462 (
		\P1_reg2_reg[17]/NET0131 ,
		_w511_,
		_w3925_
	);
	LUT2 #(
		.INIT('h8)
	) name3463 (
		\P1_reg2_reg[17]/NET0131 ,
		_w524_,
		_w3926_
	);
	LUT4 #(
		.INIT('hddd1)
	) name3464 (
		\P1_reg2_reg[17]/NET0131 ,
		_w534_,
		_w3488_,
		_w3489_,
		_w3927_
	);
	LUT4 #(
		.INIT('haa80)
	) name3465 (
		_w534_,
		_w1136_,
		_w3491_,
		_w3641_,
		_w3928_
	);
	LUT2 #(
		.INIT('h8)
	) name3466 (
		_w719_,
		_w1143_,
		_w3929_
	);
	LUT3 #(
		.INIT('h0d)
	) name3467 (
		\P1_reg2_reg[17]/NET0131 ,
		_w2411_,
		_w3929_,
		_w3930_
	);
	LUT2 #(
		.INIT('h4)
	) name3468 (
		_w3928_,
		_w3930_,
		_w3931_
	);
	LUT3 #(
		.INIT('hd0)
	) name3469 (
		_w1183_,
		_w3927_,
		_w3931_,
		_w3932_
	);
	LUT4 #(
		.INIT('hd11d)
	) name3470 (
		\P1_reg2_reg[17]/NET0131 ,
		_w534_,
		_w1431_,
		_w3498_,
		_w3933_
	);
	LUT4 #(
		.INIT('he020)
	) name3471 (
		\P1_reg2_reg[17]/NET0131 ,
		_w534_,
		_w1114_,
		_w3500_,
		_w3934_
	);
	LUT3 #(
		.INIT('h0d)
	) name3472 (
		_w1286_,
		_w3933_,
		_w3934_,
		_w3935_
	);
	LUT4 #(
		.INIT('h3111)
	) name3473 (
		_w526_,
		_w3926_,
		_w3932_,
		_w3935_,
		_w3936_
	);
	LUT3 #(
		.INIT('hce)
	) name3474 (
		\P1_state_reg[0]/NET0131 ,
		_w3925_,
		_w3936_,
		_w3937_
	);
	LUT4 #(
		.INIT('h3020)
	) name3475 (
		_w534_,
		_w1141_,
		_w3443_,
		_w3657_,
		_w3938_
	);
	LUT3 #(
		.INIT('h8a)
	) name3476 (
		\P1_reg2_reg[21]/NET0131 ,
		_w2951_,
		_w3938_,
		_w3939_
	);
	LUT2 #(
		.INIT('h8)
	) name3477 (
		_w1075_,
		_w1143_,
		_w3940_
	);
	LUT4 #(
		.INIT('h0075)
	) name3478 (
		_w534_,
		_w3652_,
		_w3655_,
		_w3940_,
		_w3941_
	);
	LUT3 #(
		.INIT('hce)
	) name3479 (
		_w3443_,
		_w3939_,
		_w3941_,
		_w3942_
	);
	LUT2 #(
		.INIT('h2)
	) name3480 (
		\P1_reg2_reg[22]/NET0131 ,
		_w511_,
		_w3943_
	);
	LUT2 #(
		.INIT('h8)
	) name3481 (
		\P1_reg2_reg[22]/NET0131 ,
		_w524_,
		_w3944_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name3482 (
		\P1_reg2_reg[22]/NET0131 ,
		_w528_,
		_w530_,
		_w533_,
		_w3945_
	);
	LUT4 #(
		.INIT('hddd1)
	) name3483 (
		\P1_reg2_reg[22]/NET0131 ,
		_w534_,
		_w3775_,
		_w3776_,
		_w3946_
	);
	LUT4 #(
		.INIT('h2822)
	) name3484 (
		_w534_,
		_w1457_,
		_w3778_,
		_w3780_,
		_w3947_
	);
	LUT3 #(
		.INIT('ha8)
	) name3485 (
		_w1114_,
		_w3945_,
		_w3947_,
		_w3948_
	);
	LUT4 #(
		.INIT('h8288)
	) name3486 (
		_w534_,
		_w1457_,
		_w3783_,
		_w3785_,
		_w3949_
	);
	LUT4 #(
		.INIT('h1dd1)
	) name3487 (
		\P1_reg2_reg[22]/NET0131 ,
		_w534_,
		_w1066_,
		_w3546_,
		_w3950_
	);
	LUT4 #(
		.INIT('h5400)
	) name3488 (
		_w541_,
		_w1062_,
		_w1065_,
		_w1138_,
		_w3951_
	);
	LUT2 #(
		.INIT('h8)
	) name3489 (
		_w1067_,
		_w1143_,
		_w3952_
	);
	LUT4 #(
		.INIT('haa20)
	) name3490 (
		\P1_reg2_reg[22]/NET0131 ,
		_w534_,
		_w1138_,
		_w1141_,
		_w3953_
	);
	LUT4 #(
		.INIT('h0007)
	) name3491 (
		_w534_,
		_w3951_,
		_w3952_,
		_w3953_,
		_w3954_
	);
	LUT3 #(
		.INIT('hd0)
	) name3492 (
		_w1136_,
		_w3950_,
		_w3954_,
		_w3955_
	);
	LUT4 #(
		.INIT('h5700)
	) name3493 (
		_w1286_,
		_w3945_,
		_w3949_,
		_w3955_,
		_w3956_
	);
	LUT4 #(
		.INIT('h0d00)
	) name3494 (
		_w1183_,
		_w3946_,
		_w3948_,
		_w3956_,
		_w3957_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name3495 (
		\P1_state_reg[0]/NET0131 ,
		_w526_,
		_w3944_,
		_w3957_,
		_w3958_
	);
	LUT2 #(
		.INIT('he)
	) name3496 (
		_w3943_,
		_w3958_,
		_w3959_
	);
	LUT2 #(
		.INIT('h2)
	) name3497 (
		\P1_reg0_reg[12]/NET0131 ,
		_w511_,
		_w3960_
	);
	LUT2 #(
		.INIT('h8)
	) name3498 (
		\P1_reg0_reg[12]/NET0131 ,
		_w524_,
		_w3961_
	);
	LUT2 #(
		.INIT('h8)
	) name3499 (
		_w1136_,
		_w3348_,
		_w3962_
	);
	LUT4 #(
		.INIT('h0001)
	) name3500 (
		_w3344_,
		_w3345_,
		_w3346_,
		_w3962_,
		_w3963_
	);
	LUT4 #(
		.INIT('h7200)
	) name3501 (
		_w537_,
		_w799_,
		_w3341_,
		_w3675_,
		_w3964_
	);
	LUT3 #(
		.INIT('h02)
	) name3502 (
		_w1140_,
		_w1468_,
		_w2688_,
		_w3965_
	);
	LUT3 #(
		.INIT('h01)
	) name3503 (
		_w1107_,
		_w1108_,
		_w2688_,
		_w3966_
	);
	LUT4 #(
		.INIT('haaa2)
	) name3504 (
		\P1_reg0_reg[12]/NET0131 ,
		_w2692_,
		_w3965_,
		_w3966_,
		_w3967_
	);
	LUT4 #(
		.INIT('h0031)
	) name3505 (
		_w2688_,
		_w3964_,
		_w3963_,
		_w3967_,
		_w3968_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name3506 (
		\P1_state_reg[0]/NET0131 ,
		_w526_,
		_w3961_,
		_w3968_,
		_w3969_
	);
	LUT2 #(
		.INIT('he)
	) name3507 (
		_w3960_,
		_w3969_,
		_w3970_
	);
	LUT4 #(
		.INIT('h70d0)
	) name3508 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg1_reg[17]/NET0131 ,
		_w1476_,
		_w3971_
	);
	LUT2 #(
		.INIT('h8)
	) name3509 (
		\P2_reg1_reg[17]/NET0131 ,
		_w1487_,
		_w3972_
	);
	LUT4 #(
		.INIT('h1dd1)
	) name3510 (
		\P2_reg1_reg[17]/NET0131 ,
		_w2039_,
		_w2705_,
		_w2706_,
		_w3973_
	);
	LUT2 #(
		.INIT('h2)
	) name3511 (
		_w2038_,
		_w3973_,
		_w3974_
	);
	LUT4 #(
		.INIT('hd11d)
	) name3512 (
		\P2_reg1_reg[17]/NET0131 ,
		_w2039_,
		_w2705_,
		_w2712_,
		_w3975_
	);
	LUT2 #(
		.INIT('h2)
	) name3513 (
		_w2193_,
		_w3975_,
		_w3976_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name3514 (
		\P2_reg1_reg[17]/NET0131 ,
		_w1491_,
		_w1493_,
		_w1496_,
		_w3977_
	);
	LUT4 #(
		.INIT('hd11d)
	) name3515 (
		\P2_reg1_reg[17]/NET0131 ,
		_w1497_,
		_w2705_,
		_w2712_,
		_w3978_
	);
	LUT4 #(
		.INIT('h8a88)
	) name3516 (
		_w1497_,
		_w2714_,
		_w2715_,
		_w2716_,
		_w3979_
	);
	LUT4 #(
		.INIT('hf100)
	) name3517 (
		_w1509_,
		_w1771_,
		_w1775_,
		_w2963_,
		_w3980_
	);
	LUT3 #(
		.INIT('ha2)
	) name3518 (
		\P2_reg1_reg[17]/NET0131 ,
		_w2633_,
		_w2660_,
		_w3981_
	);
	LUT2 #(
		.INIT('h1)
	) name3519 (
		_w3980_,
		_w3981_,
		_w3982_
	);
	LUT4 #(
		.INIT('h5700)
	) name3520 (
		_w2081_,
		_w3977_,
		_w3979_,
		_w3982_,
		_w3983_
	);
	LUT3 #(
		.INIT('hd0)
	) name3521 (
		_w2188_,
		_w3978_,
		_w3983_,
		_w3984_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name3522 (
		_w1489_,
		_w3976_,
		_w3974_,
		_w3984_,
		_w3985_
	);
	LUT4 #(
		.INIT('heeec)
	) name3523 (
		\P1_state_reg[0]/NET0131 ,
		_w3971_,
		_w3972_,
		_w3985_,
		_w3986_
	);
	LUT4 #(
		.INIT('h70d0)
	) name3524 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg1_reg[18]/NET0131 ,
		_w1476_,
		_w3987_
	);
	LUT2 #(
		.INIT('h8)
	) name3525 (
		\P2_reg1_reg[18]/NET0131 ,
		_w1487_,
		_w3988_
	);
	LUT4 #(
		.INIT('haa02)
	) name3526 (
		\P2_reg1_reg[18]/NET0131 ,
		_w1491_,
		_w1493_,
		_w1496_,
		_w3989_
	);
	LUT3 #(
		.INIT('ha8)
	) name3527 (
		_w2193_,
		_w3154_,
		_w3989_,
		_w3990_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name3528 (
		\P2_reg1_reg[18]/NET0131 ,
		_w1491_,
		_w1493_,
		_w1496_,
		_w3991_
	);
	LUT4 #(
		.INIT('h20e0)
	) name3529 (
		\P2_reg1_reg[18]/NET0131 ,
		_w1497_,
		_w2081_,
		_w2732_,
		_w3992_
	);
	LUT2 #(
		.INIT('h4)
	) name3530 (
		_w1833_,
		_w2963_,
		_w3993_
	);
	LUT3 #(
		.INIT('ha2)
	) name3531 (
		\P2_reg1_reg[18]/NET0131 ,
		_w2633_,
		_w2660_,
		_w3994_
	);
	LUT2 #(
		.INIT('h1)
	) name3532 (
		_w3993_,
		_w3994_,
		_w3995_
	);
	LUT2 #(
		.INIT('h4)
	) name3533 (
		_w3992_,
		_w3995_,
		_w3996_
	);
	LUT3 #(
		.INIT('ha8)
	) name3534 (
		_w2188_,
		_w3163_,
		_w3991_,
		_w3997_
	);
	LUT4 #(
		.INIT('h1dd1)
	) name3535 (
		\P2_reg1_reg[18]/NET0131 ,
		_w2039_,
		_w2472_,
		_w2728_,
		_w3998_
	);
	LUT2 #(
		.INIT('h2)
	) name3536 (
		_w2038_,
		_w3998_,
		_w3999_
	);
	LUT4 #(
		.INIT('h0100)
	) name3537 (
		_w3990_,
		_w3997_,
		_w3999_,
		_w3996_,
		_w4000_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name3538 (
		\P1_state_reg[0]/NET0131 ,
		_w1489_,
		_w3988_,
		_w4000_,
		_w4001_
	);
	LUT2 #(
		.INIT('he)
	) name3539 (
		_w3987_,
		_w4001_,
		_w4002_
	);
	LUT4 #(
		.INIT('h70d0)
	) name3540 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg1_reg[19]/NET0131 ,
		_w1476_,
		_w4003_
	);
	LUT2 #(
		.INIT('h8)
	) name3541 (
		\P2_reg1_reg[19]/NET0131 ,
		_w1487_,
		_w4004_
	);
	LUT4 #(
		.INIT('haa02)
	) name3542 (
		\P2_reg1_reg[19]/NET0131 ,
		_w1491_,
		_w1493_,
		_w1496_,
		_w4005_
	);
	LUT4 #(
		.INIT('h208a)
	) name3543 (
		_w2039_,
		_w2319_,
		_w2327_,
		_w2749_,
		_w4006_
	);
	LUT3 #(
		.INIT('ha8)
	) name3544 (
		_w2038_,
		_w4005_,
		_w4006_,
		_w4007_
	);
	LUT4 #(
		.INIT('h20e0)
	) name3545 (
		\P2_reg1_reg[19]/NET0131 ,
		_w1497_,
		_w2081_,
		_w2756_,
		_w4008_
	);
	LUT4 #(
		.INIT('hd11d)
	) name3546 (
		\P2_reg1_reg[19]/NET0131 ,
		_w2039_,
		_w2378_,
		_w2749_,
		_w4009_
	);
	LUT2 #(
		.INIT('h2)
	) name3547 (
		_w2193_,
		_w4009_,
		_w4010_
	);
	LUT4 #(
		.INIT('hd11d)
	) name3548 (
		\P2_reg1_reg[19]/NET0131 ,
		_w1497_,
		_w2378_,
		_w2749_,
		_w4011_
	);
	LUT3 #(
		.INIT('ha2)
	) name3549 (
		\P2_reg1_reg[19]/NET0131 ,
		_w2633_,
		_w2660_,
		_w4012_
	);
	LUT2 #(
		.INIT('h4)
	) name3550 (
		_w1813_,
		_w2963_,
		_w4013_
	);
	LUT2 #(
		.INIT('h1)
	) name3551 (
		_w4012_,
		_w4013_,
		_w4014_
	);
	LUT3 #(
		.INIT('hd0)
	) name3552 (
		_w2188_,
		_w4011_,
		_w4014_,
		_w4015_
	);
	LUT4 #(
		.INIT('h0100)
	) name3553 (
		_w4007_,
		_w4008_,
		_w4010_,
		_w4015_,
		_w4016_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name3554 (
		\P1_state_reg[0]/NET0131 ,
		_w1489_,
		_w4004_,
		_w4016_,
		_w4017_
	);
	LUT2 #(
		.INIT('he)
	) name3555 (
		_w4003_,
		_w4017_,
		_w4018_
	);
	LUT4 #(
		.INIT('h70d0)
	) name3556 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg1_reg[20]/NET0131 ,
		_w1476_,
		_w4019_
	);
	LUT2 #(
		.INIT('h8)
	) name3557 (
		\P2_reg1_reg[20]/NET0131 ,
		_w1487_,
		_w4020_
	);
	LUT4 #(
		.INIT('haa02)
	) name3558 (
		\P2_reg1_reg[20]/NET0131 ,
		_w1491_,
		_w1493_,
		_w1496_,
		_w4021_
	);
	LUT4 #(
		.INIT('h35c5)
	) name3559 (
		\P2_reg1_reg[20]/NET0131 ,
		_w1857_,
		_w2039_,
		_w3190_,
		_w4022_
	);
	LUT2 #(
		.INIT('h2)
	) name3560 (
		_w2038_,
		_w4022_,
		_w4023_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name3561 (
		\P2_reg1_reg[20]/NET0131 ,
		_w1491_,
		_w1493_,
		_w1496_,
		_w4024_
	);
	LUT4 #(
		.INIT('h111d)
	) name3562 (
		\P2_reg1_reg[20]/NET0131 ,
		_w1497_,
		_w3194_,
		_w3195_,
		_w4025_
	);
	LUT4 #(
		.INIT('h5400)
	) name3563 (
		_w1509_,
		_w1858_,
		_w1865_,
		_w2963_,
		_w4026_
	);
	LUT3 #(
		.INIT('ha2)
	) name3564 (
		\P2_reg1_reg[20]/NET0131 ,
		_w2633_,
		_w2660_,
		_w4027_
	);
	LUT2 #(
		.INIT('h1)
	) name3565 (
		_w4026_,
		_w4027_,
		_w4028_
	);
	LUT3 #(
		.INIT('hd0)
	) name3566 (
		_w2081_,
		_w4025_,
		_w4028_,
		_w4029_
	);
	LUT3 #(
		.INIT('ha8)
	) name3567 (
		_w2193_,
		_w3202_,
		_w4021_,
		_w4030_
	);
	LUT3 #(
		.INIT('ha8)
	) name3568 (
		_w2188_,
		_w3204_,
		_w4024_,
		_w4031_
	);
	LUT4 #(
		.INIT('h0100)
	) name3569 (
		_w4023_,
		_w4030_,
		_w4031_,
		_w4029_,
		_w4032_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name3570 (
		\P1_state_reg[0]/NET0131 ,
		_w1489_,
		_w4020_,
		_w4032_,
		_w4033_
	);
	LUT2 #(
		.INIT('he)
	) name3571 (
		_w4019_,
		_w4033_,
		_w4034_
	);
	LUT4 #(
		.INIT('h70d0)
	) name3572 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg1_reg[21]/NET0131 ,
		_w1476_,
		_w4035_
	);
	LUT2 #(
		.INIT('h8)
	) name3573 (
		\P2_reg1_reg[21]/NET0131 ,
		_w1487_,
		_w4036_
	);
	LUT4 #(
		.INIT('haa02)
	) name3574 (
		\P2_reg1_reg[21]/NET0131 ,
		_w1491_,
		_w1493_,
		_w1496_,
		_w4037_
	);
	LUT3 #(
		.INIT('ha8)
	) name3575 (
		_w2193_,
		_w3216_,
		_w4037_,
		_w4038_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name3576 (
		\P2_reg1_reg[21]/NET0131 ,
		_w1491_,
		_w1493_,
		_w1496_,
		_w4039_
	);
	LUT3 #(
		.INIT('ha2)
	) name3577 (
		\P2_reg1_reg[21]/NET0131 ,
		_w2633_,
		_w2660_,
		_w4040_
	);
	LUT4 #(
		.INIT('h1000)
	) name3578 (
		_w1509_,
		_w1882_,
		_w2039_,
		_w2084_,
		_w4041_
	);
	LUT2 #(
		.INIT('h1)
	) name3579 (
		_w4040_,
		_w4041_,
		_w4042_
	);
	LUT4 #(
		.INIT('h5700)
	) name3580 (
		_w2188_,
		_w3213_,
		_w4039_,
		_w4042_,
		_w4043_
	);
	LUT4 #(
		.INIT('h111d)
	) name3581 (
		\P2_reg1_reg[21]/NET0131 ,
		_w1497_,
		_w3222_,
		_w3223_,
		_w4044_
	);
	LUT2 #(
		.INIT('h2)
	) name3582 (
		_w2081_,
		_w4044_,
		_w4045_
	);
	LUT4 #(
		.INIT('h208a)
	) name3583 (
		_w2039_,
		_w2640_,
		_w2642_,
		_w3212_,
		_w4046_
	);
	LUT3 #(
		.INIT('ha8)
	) name3584 (
		_w2038_,
		_w4037_,
		_w4046_,
		_w4047_
	);
	LUT4 #(
		.INIT('h0100)
	) name3585 (
		_w4045_,
		_w4038_,
		_w4047_,
		_w4043_,
		_w4048_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name3586 (
		\P1_state_reg[0]/NET0131 ,
		_w1489_,
		_w4036_,
		_w4048_,
		_w4049_
	);
	LUT2 #(
		.INIT('he)
	) name3587 (
		_w4035_,
		_w4049_,
		_w4050_
	);
	LUT4 #(
		.INIT('ha800)
	) name3588 (
		_w2425_,
		_w2688_,
		_w3426_,
		_w3443_,
		_w4051_
	);
	LUT2 #(
		.INIT('h2)
	) name3589 (
		\P1_reg0_reg[20]/NET0131 ,
		_w4051_,
		_w4052_
	);
	LUT4 #(
		.INIT('hffb0)
	) name3590 (
		_w3606_,
		_w3608_,
		_w3651_,
		_w4052_,
		_w4053_
	);
	LUT2 #(
		.INIT('h2)
	) name3591 (
		\P1_reg1_reg[12]/NET0131 ,
		_w511_,
		_w4054_
	);
	LUT2 #(
		.INIT('h8)
	) name3592 (
		\P1_reg1_reg[12]/NET0131 ,
		_w524_,
		_w4055_
	);
	LUT3 #(
		.INIT('h2a)
	) name3593 (
		\P1_reg1_reg[12]/NET0131 ,
		_w2426_,
		_w3686_,
		_w4056_
	);
	LUT4 #(
		.INIT('h7200)
	) name3594 (
		_w537_,
		_w799_,
		_w3341_,
		_w3688_,
		_w4057_
	);
	LUT4 #(
		.INIT('h000d)
	) name3595 (
		_w2421_,
		_w3963_,
		_w4056_,
		_w4057_,
		_w4058_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name3596 (
		\P1_state_reg[0]/NET0131 ,
		_w526_,
		_w4055_,
		_w4058_,
		_w4059_
	);
	LUT2 #(
		.INIT('he)
	) name3597 (
		_w4054_,
		_w4059_,
		_w4060_
	);
	LUT2 #(
		.INIT('h2)
	) name3598 (
		\P1_reg1_reg[17]/NET0131 ,
		_w511_,
		_w4061_
	);
	LUT2 #(
		.INIT('h8)
	) name3599 (
		\P1_reg1_reg[17]/NET0131 ,
		_w524_,
		_w4062_
	);
	LUT4 #(
		.INIT('hddd1)
	) name3600 (
		\P1_reg1_reg[17]/NET0131 ,
		_w2421_,
		_w3488_,
		_w3489_,
		_w4063_
	);
	LUT2 #(
		.INIT('h2)
	) name3601 (
		\P1_reg1_reg[17]/NET0131 ,
		_w3026_,
		_w4064_
	);
	LUT4 #(
		.INIT('hcc80)
	) name3602 (
		_w1136_,
		_w2421_,
		_w3491_,
		_w3641_,
		_w4065_
	);
	LUT2 #(
		.INIT('h1)
	) name3603 (
		_w4064_,
		_w4065_,
		_w4066_
	);
	LUT3 #(
		.INIT('hd0)
	) name3604 (
		_w1183_,
		_w4063_,
		_w4066_,
		_w4067_
	);
	LUT4 #(
		.INIT('hc535)
	) name3605 (
		\P1_reg1_reg[17]/NET0131 ,
		_w1431_,
		_w2421_,
		_w3498_,
		_w4068_
	);
	LUT4 #(
		.INIT('hc808)
	) name3606 (
		\P1_reg1_reg[17]/NET0131 ,
		_w1114_,
		_w2421_,
		_w3500_,
		_w4069_
	);
	LUT3 #(
		.INIT('h0d)
	) name3607 (
		_w1286_,
		_w4068_,
		_w4069_,
		_w4070_
	);
	LUT4 #(
		.INIT('h3111)
	) name3608 (
		_w526_,
		_w4062_,
		_w4067_,
		_w4070_,
		_w4071_
	);
	LUT3 #(
		.INIT('hce)
	) name3609 (
		\P1_state_reg[0]/NET0131 ,
		_w4061_,
		_w4071_,
		_w4072_
	);
	LUT4 #(
		.INIT('h00a8)
	) name3610 (
		_w526_,
		_w528_,
		_w530_,
		_w533_,
		_w4073_
	);
	LUT2 #(
		.INIT('h8)
	) name3611 (
		\P1_state_reg[0]/NET0131 ,
		_w4073_,
		_w4074_
	);
	LUT4 #(
		.INIT('hd000)
	) name3612 (
		_w1138_,
		_w2421_,
		_w2425_,
		_w3443_,
		_w4075_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name3613 (
		\P1_reg1_reg[20]/NET0131 ,
		_w3684_,
		_w3685_,
		_w4075_,
		_w4076_
	);
	LUT4 #(
		.INIT('hffb0)
	) name3614 (
		_w3606_,
		_w3608_,
		_w4074_,
		_w4076_,
		_w4077_
	);
	LUT2 #(
		.INIT('h1)
	) name3615 (
		_w2421_,
		_w3657_,
		_w4078_
	);
	LUT4 #(
		.INIT('hc080)
	) name3616 (
		_w2421_,
		_w2425_,
		_w3443_,
		_w3657_,
		_w4079_
	);
	LUT3 #(
		.INIT('h8a)
	) name3617 (
		\P1_reg1_reg[21]/NET0131 ,
		_w3685_,
		_w4079_,
		_w4080_
	);
	LUT4 #(
		.INIT('hffb0)
	) name3618 (
		_w3652_,
		_w3655_,
		_w4074_,
		_w4080_,
		_w4081_
	);
	LUT2 #(
		.INIT('h8)
	) name3619 (
		_w524_,
		_w816_,
		_w4082_
	);
	LUT4 #(
		.INIT('h1f00)
	) name3620 (
		_w528_,
		_w530_,
		_w533_,
		_w816_,
		_w4083_
	);
	LUT4 #(
		.INIT('h6555)
	) name3621 (
		_w799_,
		_w924_,
		_w1154_,
		_w1157_,
		_w4084_
	);
	LUT4 #(
		.INIT('h7020)
	) name3622 (
		_w537_,
		_w833_,
		_w2197_,
		_w4084_,
		_w4085_
	);
	LUT3 #(
		.INIT('ha8)
	) name3623 (
		_w1183_,
		_w4083_,
		_w4085_,
		_w4086_
	);
	LUT4 #(
		.INIT('h007b)
	) name3624 (
		_w1438_,
		_w2197_,
		_w3076_,
		_w4083_,
		_w4087_
	);
	LUT2 #(
		.INIT('h2)
	) name3625 (
		_w1286_,
		_w4087_,
		_w4088_
	);
	LUT4 #(
		.INIT('h00b7)
	) name3626 (
		_w1438_,
		_w2197_,
		_w3052_,
		_w4083_,
		_w4089_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name3627 (
		_w827_,
		_w842_,
		_w907_,
		_w1117_,
		_w4090_
	);
	LUT4 #(
		.INIT('hc808)
	) name3628 (
		_w816_,
		_w1136_,
		_w2197_,
		_w4090_,
		_w4091_
	);
	LUT3 #(
		.INIT('h04)
	) name3629 (
		_w827_,
		_w2259_,
		_w2260_,
		_w4092_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name3630 (
		_w816_,
		_w1138_,
		_w1141_,
		_w2197_,
		_w4093_
	);
	LUT2 #(
		.INIT('h1)
	) name3631 (
		_w4092_,
		_w4093_,
		_w4094_
	);
	LUT2 #(
		.INIT('h4)
	) name3632 (
		_w4091_,
		_w4094_,
		_w4095_
	);
	LUT3 #(
		.INIT('hd0)
	) name3633 (
		_w1114_,
		_w4089_,
		_w4095_,
		_w4096_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name3634 (
		_w526_,
		_w4086_,
		_w4088_,
		_w4096_,
		_w4097_
	);
	LUT2 #(
		.INIT('h2)
	) name3635 (
		\P1_reg3_reg[10]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w4098_
	);
	LUT3 #(
		.INIT('h07)
	) name3636 (
		_w816_,
		_w1294_,
		_w4098_,
		_w4099_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name3637 (
		\P1_state_reg[0]/NET0131 ,
		_w4082_,
		_w4097_,
		_w4099_,
		_w4100_
	);
	LUT2 #(
		.INIT('h8)
	) name3638 (
		_w524_,
		_w760_,
		_w4101_
	);
	LUT4 #(
		.INIT('h1f00)
	) name3639 (
		_w528_,
		_w530_,
		_w533_,
		_w760_,
		_w4102_
	);
	LUT4 #(
		.INIT('h4150)
	) name3640 (
		_w537_,
		_w762_,
		_w772_,
		_w1161_,
		_w4103_
	);
	LUT3 #(
		.INIT('h80)
	) name3641 (
		_w537_,
		_w750_,
		_w751_,
		_w4104_
	);
	LUT4 #(
		.INIT('h3331)
	) name3642 (
		_w2197_,
		_w4102_,
		_w4103_,
		_w4104_,
		_w4105_
	);
	LUT2 #(
		.INIT('h2)
	) name3643 (
		_w1183_,
		_w4105_,
		_w4106_
	);
	LUT4 #(
		.INIT('h9a55)
	) name3644 (
		_w1444_,
		_w3076_,
		_w3077_,
		_w3079_,
		_w4107_
	);
	LUT4 #(
		.INIT('hc808)
	) name3645 (
		_w760_,
		_w1286_,
		_w2197_,
		_w4107_,
		_w4108_
	);
	LUT4 #(
		.INIT('h9599)
	) name3646 (
		_w1444_,
		_w3045_,
		_w3052_,
		_w3053_,
		_w4109_
	);
	LUT4 #(
		.INIT('h08c8)
	) name3647 (
		_w760_,
		_w1114_,
		_w2197_,
		_w4109_,
		_w4110_
	);
	LUT4 #(
		.INIT('h6c00)
	) name3648 (
		_w758_,
		_w767_,
		_w1120_,
		_w2197_,
		_w4111_
	);
	LUT3 #(
		.INIT('h04)
	) name3649 (
		_w767_,
		_w2259_,
		_w2260_,
		_w4112_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name3650 (
		_w760_,
		_w1138_,
		_w1141_,
		_w2197_,
		_w4113_
	);
	LUT2 #(
		.INIT('h1)
	) name3651 (
		_w4112_,
		_w4113_,
		_w4114_
	);
	LUT4 #(
		.INIT('h5700)
	) name3652 (
		_w1136_,
		_w4102_,
		_w4111_,
		_w4114_,
		_w4115_
	);
	LUT3 #(
		.INIT('h10)
	) name3653 (
		_w4110_,
		_w4108_,
		_w4115_,
		_w4116_
	);
	LUT4 #(
		.INIT('h1311)
	) name3654 (
		_w526_,
		_w4101_,
		_w4106_,
		_w4116_,
		_w4117_
	);
	LUT2 #(
		.INIT('h2)
	) name3655 (
		\P1_reg3_reg[14]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w4118_
	);
	LUT3 #(
		.INIT('h07)
	) name3656 (
		_w760_,
		_w1294_,
		_w4118_,
		_w4119_
	);
	LUT3 #(
		.INIT('h2f)
	) name3657 (
		\P1_state_reg[0]/NET0131 ,
		_w4117_,
		_w4119_,
		_w4120_
	);
	LUT2 #(
		.INIT('h8)
	) name3658 (
		_w524_,
		_w770_,
		_w4121_
	);
	LUT4 #(
		.INIT('h1f00)
	) name3659 (
		_w528_,
		_w530_,
		_w533_,
		_w770_,
		_w4122_
	);
	LUT4 #(
		.INIT('h1e0f)
	) name3660 (
		_w762_,
		_w772_,
		_w791_,
		_w1161_,
		_w4123_
	);
	LUT4 #(
		.INIT('h7020)
	) name3661 (
		_w537_,
		_w762_,
		_w2197_,
		_w4123_,
		_w4124_
	);
	LUT3 #(
		.INIT('ha8)
	) name3662 (
		_w1183_,
		_w4122_,
		_w4124_,
		_w4125_
	);
	LUT4 #(
		.INIT('h9a55)
	) name3663 (
		_w1447_,
		_w2843_,
		_w2844_,
		_w2845_,
		_w4126_
	);
	LUT4 #(
		.INIT('hc808)
	) name3664 (
		_w770_,
		_w1286_,
		_w2197_,
		_w4126_,
		_w4127_
	);
	LUT4 #(
		.INIT('h9a55)
	) name3665 (
		_w1447_,
		_w2871_,
		_w2872_,
		_w2873_,
		_w4128_
	);
	LUT4 #(
		.INIT('h08c8)
	) name3666 (
		_w770_,
		_w1114_,
		_w2197_,
		_w4128_,
		_w4129_
	);
	LUT4 #(
		.INIT('h6a00)
	) name3667 (
		_w780_,
		_w1120_,
		_w1121_,
		_w2197_,
		_w4130_
	);
	LUT3 #(
		.INIT('h04)
	) name3668 (
		_w780_,
		_w2259_,
		_w2260_,
		_w4131_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name3669 (
		_w770_,
		_w1138_,
		_w1141_,
		_w2197_,
		_w4132_
	);
	LUT2 #(
		.INIT('h1)
	) name3670 (
		_w4131_,
		_w4132_,
		_w4133_
	);
	LUT4 #(
		.INIT('h5700)
	) name3671 (
		_w1136_,
		_w4122_,
		_w4130_,
		_w4133_,
		_w4134_
	);
	LUT3 #(
		.INIT('h10)
	) name3672 (
		_w4129_,
		_w4127_,
		_w4134_,
		_w4135_
	);
	LUT4 #(
		.INIT('h1311)
	) name3673 (
		_w526_,
		_w4121_,
		_w4125_,
		_w4135_,
		_w4136_
	);
	LUT2 #(
		.INIT('h2)
	) name3674 (
		\P1_reg3_reg[15]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w4137_
	);
	LUT3 #(
		.INIT('h07)
	) name3675 (
		_w770_,
		_w1294_,
		_w4137_,
		_w4138_
	);
	LUT3 #(
		.INIT('h2f)
	) name3676 (
		\P1_state_reg[0]/NET0131 ,
		_w4136_,
		_w4138_,
		_w4139_
	);
	LUT2 #(
		.INIT('h2)
	) name3677 (
		_w1487_,
		_w1643_,
		_w4140_
	);
	LUT4 #(
		.INIT('h001f)
	) name3678 (
		_w1491_,
		_w1493_,
		_w1496_,
		_w1643_,
		_w4141_
	);
	LUT3 #(
		.INIT('h78)
	) name3679 (
		_w1644_,
		_w1645_,
		_w1657_,
		_w4142_
	);
	LUT4 #(
		.INIT('h070d)
	) name3680 (
		_w2272_,
		_w2467_,
		_w4141_,
		_w4142_,
		_w4143_
	);
	LUT3 #(
		.INIT('h04)
	) name3681 (
		_w1657_,
		_w2083_,
		_w2282_,
		_w4144_
	);
	LUT3 #(
		.INIT('h54)
	) name3682 (
		_w1643_,
		_w2086_,
		_w2280_,
		_w4145_
	);
	LUT2 #(
		.INIT('h1)
	) name3683 (
		_w4144_,
		_w4145_,
		_w4146_
	);
	LUT3 #(
		.INIT('he0)
	) name3684 (
		_w2276_,
		_w4143_,
		_w4146_,
		_w4147_
	);
	LUT4 #(
		.INIT('h00fe)
	) name3685 (
		_w1491_,
		_w1493_,
		_w1496_,
		_w1643_,
		_w4148_
	);
	LUT3 #(
		.INIT('h40)
	) name3686 (
		_w1676_,
		_w2057_,
		_w2060_,
		_w4149_
	);
	LUT4 #(
		.INIT('h1000)
	) name3687 (
		_w1663_,
		_w1676_,
		_w2057_,
		_w2060_,
		_w4150_
	);
	LUT3 #(
		.INIT('h10)
	) name3688 (
		_w1619_,
		_w1646_,
		_w4150_,
		_w4151_
	);
	LUT4 #(
		.INIT('h0605)
	) name3689 (
		_w1619_,
		_w1646_,
		_w2042_,
		_w4150_,
		_w4152_
	);
	LUT3 #(
		.INIT('h70)
	) name3690 (
		_w1661_,
		_w1662_,
		_w2042_,
		_w4153_
	);
	LUT4 #(
		.INIT('h1113)
	) name3691 (
		_w2277_,
		_w4148_,
		_w4152_,
		_w4153_,
		_w4154_
	);
	LUT2 #(
		.INIT('h2)
	) name3692 (
		_w2081_,
		_w4154_,
		_w4155_
	);
	LUT4 #(
		.INIT('h8a20)
	) name3693 (
		_w2272_,
		_w2492_,
		_w2493_,
		_w4142_,
		_w4156_
	);
	LUT3 #(
		.INIT('h54)
	) name3694 (
		_w2192_,
		_w4141_,
		_w4156_,
		_w4157_
	);
	LUT4 #(
		.INIT('h007d)
	) name3695 (
		_w2277_,
		_w2467_,
		_w4142_,
		_w4148_,
		_w4158_
	);
	LUT2 #(
		.INIT('h2)
	) name3696 (
		_w2290_,
		_w4158_,
		_w4159_
	);
	LUT4 #(
		.INIT('h0100)
	) name3697 (
		_w4157_,
		_w4159_,
		_w4155_,
		_w4147_,
		_w4160_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name3698 (
		\P1_state_reg[0]/NET0131 ,
		_w1489_,
		_w4140_,
		_w4160_,
		_w4161_
	);
	LUT2 #(
		.INIT('h4)
	) name3699 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[10]/NET0131 ,
		_w4162_
	);
	LUT4 #(
		.INIT('h0028)
	) name3700 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		_w1476_,
		_w1643_,
		_w4163_
	);
	LUT2 #(
		.INIT('h1)
	) name3701 (
		_w4162_,
		_w4163_,
		_w4164_
	);
	LUT2 #(
		.INIT('hb)
	) name3702 (
		_w4161_,
		_w4164_,
		_w4165_
	);
	LUT2 #(
		.INIT('h8)
	) name3703 (
		\P1_state_reg[0]/NET0131 ,
		_w1489_,
		_w4166_
	);
	LUT4 #(
		.INIT('h00fe)
	) name3704 (
		_w1491_,
		_w1493_,
		_w1496_,
		_w1732_,
		_w4167_
	);
	LUT2 #(
		.INIT('h6)
	) name3705 (
		_w1735_,
		_w1746_,
		_w4168_
	);
	LUT4 #(
		.INIT('h40b0)
	) name3706 (
		_w1687_,
		_w1692_,
		_w2277_,
		_w4168_,
		_w4169_
	);
	LUT3 #(
		.INIT('h04)
	) name3707 (
		_w1746_,
		_w2083_,
		_w2282_,
		_w4170_
	);
	LUT3 #(
		.INIT('h54)
	) name3708 (
		_w1732_,
		_w2086_,
		_w2280_,
		_w4171_
	);
	LUT2 #(
		.INIT('h1)
	) name3709 (
		_w4170_,
		_w4171_,
		_w4172_
	);
	LUT4 #(
		.INIT('h5700)
	) name3710 (
		_w2290_,
		_w4167_,
		_w4169_,
		_w4172_,
		_w4173_
	);
	LUT4 #(
		.INIT('h001f)
	) name3711 (
		_w1491_,
		_w1493_,
		_w1496_,
		_w1732_,
		_w4174_
	);
	LUT4 #(
		.INIT('h40b0)
	) name3712 (
		_w1687_,
		_w1692_,
		_w2272_,
		_w4168_,
		_w4175_
	);
	LUT3 #(
		.INIT('h54)
	) name3713 (
		_w2276_,
		_w4174_,
		_w4175_,
		_w4176_
	);
	LUT3 #(
		.INIT('h70)
	) name3714 (
		_w1616_,
		_w1618_,
		_w2042_,
		_w4177_
	);
	LUT4 #(
		.INIT('h0100)
	) name3715 (
		_w1619_,
		_w1646_,
		_w1735_,
		_w4150_,
		_w4178_
	);
	LUT4 #(
		.INIT('h1555)
	) name3716 (
		_w2042_,
		_w2057_,
		_w2060_,
		_w2064_,
		_w4179_
	);
	LUT4 #(
		.INIT('h0233)
	) name3717 (
		_w1751_,
		_w4177_,
		_w4178_,
		_w4179_,
		_w4180_
	);
	LUT4 #(
		.INIT('h04c4)
	) name3718 (
		_w1732_,
		_w2081_,
		_w2277_,
		_w4180_,
		_w4181_
	);
	LUT4 #(
		.INIT('h8a75)
	) name3719 (
		_w2102_,
		_w2124_,
		_w2126_,
		_w4168_,
		_w4182_
	);
	LUT4 #(
		.INIT('h0131)
	) name3720 (
		_w1732_,
		_w2192_,
		_w2272_,
		_w4182_,
		_w4183_
	);
	LUT4 #(
		.INIT('h0100)
	) name3721 (
		_w4181_,
		_w4183_,
		_w4176_,
		_w4173_,
		_w4184_
	);
	LUT2 #(
		.INIT('h4)
	) name3722 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[12]/NET0131 ,
		_w4185_
	);
	LUT4 #(
		.INIT('hbb93)
	) name3723 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[12]/NET0131 ,
		_w466_,
		_w1489_,
		_w4186_
	);
	LUT3 #(
		.INIT('h2f)
	) name3724 (
		_w4166_,
		_w4184_,
		_w4186_,
		_w4187_
	);
	LUT2 #(
		.INIT('h2)
	) name3725 (
		_w1487_,
		_w1749_,
		_w4188_
	);
	LUT4 #(
		.INIT('h00fe)
	) name3726 (
		_w1491_,
		_w1493_,
		_w1496_,
		_w1749_,
		_w4189_
	);
	LUT2 #(
		.INIT('h9)
	) name3727 (
		_w1751_,
		_w1761_,
		_w4190_
	);
	LUT4 #(
		.INIT('h8a20)
	) name3728 (
		_w2277_,
		_w2536_,
		_w2541_,
		_w4190_,
		_w4191_
	);
	LUT3 #(
		.INIT('ha8)
	) name3729 (
		_w2290_,
		_w4189_,
		_w4191_,
		_w4192_
	);
	LUT4 #(
		.INIT('h001f)
	) name3730 (
		_w1491_,
		_w1493_,
		_w1496_,
		_w1749_,
		_w4193_
	);
	LUT4 #(
		.INIT('h8a20)
	) name3731 (
		_w2272_,
		_w2536_,
		_w2541_,
		_w4190_,
		_w4194_
	);
	LUT3 #(
		.INIT('h54)
	) name3732 (
		_w2276_,
		_w4193_,
		_w4194_,
		_w4195_
	);
	LUT4 #(
		.INIT('h208a)
	) name3733 (
		_w2272_,
		_w2563_,
		_w2554_,
		_w4190_,
		_w4196_
	);
	LUT3 #(
		.INIT('h54)
	) name3734 (
		_w2192_,
		_w4193_,
		_w4196_,
		_w4197_
	);
	LUT3 #(
		.INIT('h70)
	) name3735 (
		_w1733_,
		_w1734_,
		_w2042_,
		_w4198_
	);
	LUT4 #(
		.INIT('h00de)
	) name3736 (
		_w1720_,
		_w2042_,
		_w2065_,
		_w4198_,
		_w4199_
	);
	LUT4 #(
		.INIT('h04c4)
	) name3737 (
		_w1749_,
		_w2081_,
		_w2277_,
		_w4199_,
		_w4200_
	);
	LUT3 #(
		.INIT('h04)
	) name3738 (
		_w1761_,
		_w2083_,
		_w2282_,
		_w4201_
	);
	LUT3 #(
		.INIT('h54)
	) name3739 (
		_w1749_,
		_w2086_,
		_w2280_,
		_w4202_
	);
	LUT2 #(
		.INIT('h1)
	) name3740 (
		_w4201_,
		_w4202_,
		_w4203_
	);
	LUT2 #(
		.INIT('h4)
	) name3741 (
		_w4200_,
		_w4203_,
		_w4204_
	);
	LUT4 #(
		.INIT('h0100)
	) name3742 (
		_w4195_,
		_w4192_,
		_w4197_,
		_w4204_,
		_w4205_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name3743 (
		\P1_state_reg[0]/NET0131 ,
		_w1489_,
		_w4188_,
		_w4205_,
		_w4206_
	);
	LUT2 #(
		.INIT('h4)
	) name3744 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[13]/NET0131 ,
		_w4207_
	);
	LUT3 #(
		.INIT('h0b)
	) name3745 (
		_w1749_,
		_w2293_,
		_w4207_,
		_w4208_
	);
	LUT2 #(
		.INIT('hb)
	) name3746 (
		_w4206_,
		_w4208_,
		_w4209_
	);
	LUT2 #(
		.INIT('h8)
	) name3747 (
		_w524_,
		_w831_,
		_w4210_
	);
	LUT4 #(
		.INIT('h1f00)
	) name3748 (
		_w528_,
		_w530_,
		_w533_,
		_w831_,
		_w4211_
	);
	LUT4 #(
		.INIT('h0705)
	) name3749 (
		_w819_,
		_w833_,
		_w1158_,
		_w3728_,
		_w4212_
	);
	LUT4 #(
		.INIT('h7020)
	) name3750 (
		_w537_,
		_w903_,
		_w2197_,
		_w4212_,
		_w4213_
	);
	LUT4 #(
		.INIT('h40b0)
	) name3751 (
		_w942_,
		_w949_,
		_w1114_,
		_w1450_,
		_w4214_
	);
	LUT4 #(
		.INIT('h00b7)
	) name3752 (
		_w1233_,
		_w1286_,
		_w1450_,
		_w4214_,
		_w4215_
	);
	LUT4 #(
		.INIT('h00b7)
	) name3753 (
		_w842_,
		_w2197_,
		_w3734_,
		_w4211_,
		_w4216_
	);
	LUT3 #(
		.INIT('h04)
	) name3754 (
		_w842_,
		_w2259_,
		_w2260_,
		_w4217_
	);
	LUT4 #(
		.INIT('h888a)
	) name3755 (
		_w831_,
		_w1141_,
		_w2197_,
		_w3118_,
		_w4218_
	);
	LUT2 #(
		.INIT('h1)
	) name3756 (
		_w4217_,
		_w4218_,
		_w4219_
	);
	LUT3 #(
		.INIT('hd0)
	) name3757 (
		_w1136_,
		_w4216_,
		_w4219_,
		_w4220_
	);
	LUT3 #(
		.INIT('hd0)
	) name3758 (
		_w2197_,
		_w4215_,
		_w4220_,
		_w4221_
	);
	LUT4 #(
		.INIT('h5700)
	) name3759 (
		_w1183_,
		_w4211_,
		_w4213_,
		_w4221_,
		_w4222_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name3760 (
		\P1_state_reg[0]/NET0131 ,
		_w526_,
		_w4210_,
		_w4222_,
		_w4223_
	);
	LUT2 #(
		.INIT('h2)
	) name3761 (
		\P1_reg3_reg[9]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w4224_
	);
	LUT3 #(
		.INIT('h07)
	) name3762 (
		_w831_,
		_w1294_,
		_w4224_,
		_w4225_
	);
	LUT2 #(
		.INIT('hb)
	) name3763 (
		_w4223_,
		_w4225_,
		_w4226_
	);
	LUT2 #(
		.INIT('h2)
	) name3764 (
		_w1487_,
		_w1660_,
		_w4227_
	);
	LUT2 #(
		.INIT('h6)
	) name3765 (
		_w1663_,
		_w1672_,
		_w4228_
	);
	LUT4 #(
		.INIT('hb04f)
	) name3766 (
		_w2304_,
		_w2533_,
		_w2534_,
		_w4228_,
		_w4229_
	);
	LUT4 #(
		.INIT('h0d01)
	) name3767 (
		_w1660_,
		_w2272_,
		_w2276_,
		_w4229_,
		_w4230_
	);
	LUT4 #(
		.INIT('h708f)
	) name3768 (
		_w2355_,
		_w2357_,
		_w2561_,
		_w4228_,
		_w4231_
	);
	LUT4 #(
		.INIT('h0131)
	) name3769 (
		_w1660_,
		_w2192_,
		_w2272_,
		_w4231_,
		_w4232_
	);
	LUT3 #(
		.INIT('h04)
	) name3770 (
		_w1672_,
		_w2083_,
		_w2282_,
		_w4233_
	);
	LUT3 #(
		.INIT('h54)
	) name3771 (
		_w1660_,
		_w2086_,
		_w2280_,
		_w4234_
	);
	LUT2 #(
		.INIT('h1)
	) name3772 (
		_w4233_,
		_w4234_,
		_w4235_
	);
	LUT3 #(
		.INIT('h10)
	) name3773 (
		_w4230_,
		_w4232_,
		_w4235_,
		_w4236_
	);
	LUT3 #(
		.INIT('h70)
	) name3774 (
		_w1673_,
		_w1675_,
		_w2042_,
		_w4237_
	);
	LUT4 #(
		.INIT('h00de)
	) name3775 (
		_w1646_,
		_w2042_,
		_w4150_,
		_w4237_,
		_w4238_
	);
	LUT4 #(
		.INIT('h04c4)
	) name3776 (
		_w1660_,
		_w2081_,
		_w2277_,
		_w4238_,
		_w4239_
	);
	LUT4 #(
		.INIT('hd010)
	) name3777 (
		_w1660_,
		_w2277_,
		_w2290_,
		_w4229_,
		_w4240_
	);
	LUT2 #(
		.INIT('h1)
	) name3778 (
		_w4239_,
		_w4240_,
		_w4241_
	);
	LUT4 #(
		.INIT('h3111)
	) name3779 (
		_w1489_,
		_w4227_,
		_w4236_,
		_w4241_,
		_w4242_
	);
	LUT2 #(
		.INIT('h4)
	) name3780 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[9]/NET0131 ,
		_w4243_
	);
	LUT4 #(
		.INIT('h0028)
	) name3781 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		_w1476_,
		_w1660_,
		_w4244_
	);
	LUT2 #(
		.INIT('h1)
	) name3782 (
		_w4243_,
		_w4244_,
		_w4245_
	);
	LUT3 #(
		.INIT('h2f)
	) name3783 (
		\P1_state_reg[0]/NET0131 ,
		_w4242_,
		_w4245_,
		_w4246_
	);
	LUT3 #(
		.INIT('h8a)
	) name3784 (
		\P1_reg1_reg[8]/NET0131 ,
		_w3685_,
		_w4079_,
		_w4247_
	);
	LUT4 #(
		.INIT('h0001)
	) name3785 (
		_w907_,
		_w1104_,
		_w1106_,
		_w1111_,
		_w4248_
	);
	LUT3 #(
		.INIT('h07)
	) name3786 (
		_w1136_,
		_w3735_,
		_w4248_,
		_w4249_
	);
	LUT3 #(
		.INIT('h10)
	) name3787 (
		_w3732_,
		_w3733_,
		_w4249_,
		_w4250_
	);
	LUT4 #(
		.INIT('h80f0)
	) name3788 (
		_w1183_,
		_w3730_,
		_w4074_,
		_w4250_,
		_w4251_
	);
	LUT2 #(
		.INIT('he)
	) name3789 (
		_w4247_,
		_w4251_,
		_w4252_
	);
	LUT3 #(
		.INIT('h8a)
	) name3790 (
		\P1_reg1_reg[9]/NET0131 ,
		_w3685_,
		_w4079_,
		_w4253_
	);
	LUT4 #(
		.INIT('h7020)
	) name3791 (
		_w537_,
		_w903_,
		_w1183_,
		_w4212_,
		_w4254_
	);
	LUT2 #(
		.INIT('h4)
	) name3792 (
		_w842_,
		_w1138_,
		_w4255_
	);
	LUT4 #(
		.INIT('h00b7)
	) name3793 (
		_w842_,
		_w1136_,
		_w3734_,
		_w4255_,
		_w4256_
	);
	LUT2 #(
		.INIT('h8)
	) name3794 (
		_w4215_,
		_w4256_,
		_w4257_
	);
	LUT4 #(
		.INIT('hecee)
	) name3795 (
		_w4074_,
		_w4253_,
		_w4254_,
		_w4257_,
		_w4258_
	);
	LUT4 #(
		.INIT('h70d0)
	) name3796 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg0_reg[23]/NET0131 ,
		_w1476_,
		_w4259_
	);
	LUT2 #(
		.INIT('h8)
	) name3797 (
		\P2_reg0_reg[23]/NET0131 ,
		_w1487_,
		_w4260_
	);
	LUT4 #(
		.INIT('h20e0)
	) name3798 (
		\P2_reg0_reg[23]/NET0131 ,
		_w2272_,
		_w2290_,
		_w3516_,
		_w4261_
	);
	LUT4 #(
		.INIT('haaa8)
	) name3799 (
		\P2_reg0_reg[23]/NET0131 ,
		_w1491_,
		_w1493_,
		_w1496_,
		_w4262_
	);
	LUT4 #(
		.INIT('h0232)
	) name3800 (
		\P2_reg0_reg[23]/NET0131 ,
		_w2276_,
		_w2277_,
		_w3516_,
		_w4263_
	);
	LUT4 #(
		.INIT('h08c8)
	) name3801 (
		\P2_reg0_reg[23]/NET0131 ,
		_w2081_,
		_w2272_,
		_w3521_,
		_w4264_
	);
	LUT4 #(
		.INIT('h8288)
	) name3802 (
		_w2277_,
		_w3511_,
		_w3524_,
		_w3526_,
		_w4265_
	);
	LUT3 #(
		.INIT('ha2)
	) name3803 (
		\P2_reg0_reg[23]/NET0131 ,
		_w2633_,
		_w2634_,
		_w4266_
	);
	LUT3 #(
		.INIT('h10)
	) name3804 (
		_w1509_,
		_w1903_,
		_w2920_,
		_w4267_
	);
	LUT2 #(
		.INIT('h1)
	) name3805 (
		_w4266_,
		_w4267_,
		_w4268_
	);
	LUT4 #(
		.INIT('hab00)
	) name3806 (
		_w2192_,
		_w4262_,
		_w4265_,
		_w4268_,
		_w4269_
	);
	LUT4 #(
		.INIT('h0100)
	) name3807 (
		_w4264_,
		_w4263_,
		_w4261_,
		_w4269_,
		_w4270_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name3808 (
		\P1_state_reg[0]/NET0131 ,
		_w1489_,
		_w4260_,
		_w4270_,
		_w4271_
	);
	LUT2 #(
		.INIT('he)
	) name3809 (
		_w4259_,
		_w4271_,
		_w4272_
	);
	LUT2 #(
		.INIT('h2)
	) name3810 (
		\P1_reg2_reg[23]/NET0131 ,
		_w511_,
		_w4273_
	);
	LUT2 #(
		.INIT('h8)
	) name3811 (
		\P1_reg2_reg[23]/NET0131 ,
		_w524_,
		_w4274_
	);
	LUT3 #(
		.INIT('h10)
	) name3812 (
		_w541_,
		_w1046_,
		_w1138_,
		_w4275_
	);
	LUT2 #(
		.INIT('h8)
	) name3813 (
		_w1048_,
		_w1143_,
		_w4276_
	);
	LUT3 #(
		.INIT('h0d)
	) name3814 (
		\P1_reg2_reg[23]/NET0131 ,
		_w3603_,
		_w4276_,
		_w4277_
	);
	LUT4 #(
		.INIT('h5d00)
	) name3815 (
		_w534_,
		_w3763_,
		_w4275_,
		_w4277_,
		_w4278_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name3816 (
		\P1_state_reg[0]/NET0131 ,
		_w526_,
		_w4274_,
		_w4278_,
		_w4279_
	);
	LUT2 #(
		.INIT('he)
	) name3817 (
		_w4273_,
		_w4279_,
		_w4280_
	);
	LUT2 #(
		.INIT('h2)
	) name3818 (
		\P1_reg2_reg[30]/NET0131 ,
		_w511_,
		_w4281_
	);
	LUT2 #(
		.INIT('h8)
	) name3819 (
		\P1_reg2_reg[30]/NET0131 ,
		_w524_,
		_w4282_
	);
	LUT4 #(
		.INIT('h5455)
	) name3820 (
		\P1_reg2_reg[30]/NET0131 ,
		_w528_,
		_w530_,
		_w533_,
		_w4283_
	);
	LUT2 #(
		.INIT('h2)
	) name3821 (
		_w1136_,
		_w4283_,
		_w4284_
	);
	LUT4 #(
		.INIT('hd700)
	) name3822 (
		_w534_,
		_w1133_,
		_w1312_,
		_w4284_,
		_w4285_
	);
	LUT3 #(
		.INIT('h10)
	) name3823 (
		_w541_,
		_w1311_,
		_w3288_,
		_w4286_
	);
	LUT4 #(
		.INIT('h0a02)
	) name3824 (
		\P1_reg2_reg[30]/NET0131 ,
		_w534_,
		_w1135_,
		_w1141_,
		_w4287_
	);
	LUT2 #(
		.INIT('h1)
	) name3825 (
		_w1144_,
		_w4287_,
		_w4288_
	);
	LUT2 #(
		.INIT('h4)
	) name3826 (
		_w4286_,
		_w4288_,
		_w4289_
	);
	LUT4 #(
		.INIT('h0700)
	) name3827 (
		_w3286_,
		_w3287_,
		_w4285_,
		_w4289_,
		_w4290_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name3828 (
		\P1_state_reg[0]/NET0131 ,
		_w526_,
		_w4282_,
		_w4290_,
		_w4291_
	);
	LUT2 #(
		.INIT('he)
	) name3829 (
		_w4281_,
		_w4291_,
		_w4292_
	);
	LUT4 #(
		.INIT('h70d0)
	) name3830 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg1_reg[23]/NET0131 ,
		_w1476_,
		_w4293_
	);
	LUT2 #(
		.INIT('h8)
	) name3831 (
		\P2_reg1_reg[23]/NET0131 ,
		_w1487_,
		_w4294_
	);
	LUT4 #(
		.INIT('haa02)
	) name3832 (
		\P2_reg1_reg[23]/NET0131 ,
		_w1491_,
		_w1493_,
		_w1496_,
		_w4295_
	);
	LUT4 #(
		.INIT('h08c8)
	) name3833 (
		\P2_reg1_reg[23]/NET0131 ,
		_w2038_,
		_w2039_,
		_w3516_,
		_w4296_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name3834 (
		\P2_reg1_reg[23]/NET0131 ,
		_w1491_,
		_w1493_,
		_w1496_,
		_w4297_
	);
	LUT4 #(
		.INIT('h20e0)
	) name3835 (
		\P2_reg1_reg[23]/NET0131 ,
		_w1497_,
		_w2081_,
		_w3521_,
		_w4298_
	);
	LUT3 #(
		.INIT('ha8)
	) name3836 (
		_w2188_,
		_w3529_,
		_w4297_,
		_w4299_
	);
	LUT3 #(
		.INIT('ha2)
	) name3837 (
		\P2_reg1_reg[23]/NET0131 ,
		_w2633_,
		_w2660_,
		_w4300_
	);
	LUT3 #(
		.INIT('h10)
	) name3838 (
		_w1509_,
		_w1903_,
		_w2963_,
		_w4301_
	);
	LUT2 #(
		.INIT('h1)
	) name3839 (
		_w4300_,
		_w4301_,
		_w4302_
	);
	LUT4 #(
		.INIT('h5700)
	) name3840 (
		_w2193_,
		_w3527_,
		_w4295_,
		_w4302_,
		_w4303_
	);
	LUT4 #(
		.INIT('h0100)
	) name3841 (
		_w4296_,
		_w4298_,
		_w4299_,
		_w4303_,
		_w4304_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name3842 (
		\P1_state_reg[0]/NET0131 ,
		_w1489_,
		_w4294_,
		_w4304_,
		_w4305_
	);
	LUT2 #(
		.INIT('he)
	) name3843 (
		_w4293_,
		_w4305_,
		_w4306_
	);
	LUT4 #(
		.INIT('h80aa)
	) name3844 (
		_w534_,
		_w1183_,
		_w3730_,
		_w4250_,
		_w4307_
	);
	LUT2 #(
		.INIT('h8)
	) name3845 (
		_w901_,
		_w1143_,
		_w4308_
	);
	LUT3 #(
		.INIT('ha8)
	) name3846 (
		_w3443_,
		_w4307_,
		_w4308_,
		_w4309_
	);
	LUT4 #(
		.INIT('h3b00)
	) name3847 (
		_w534_,
		_w1183_,
		_w3730_,
		_w3938_,
		_w4310_
	);
	LUT2 #(
		.INIT('h2)
	) name3848 (
		\P1_reg2_reg[8]/NET0131 ,
		_w4310_,
		_w4311_
	);
	LUT2 #(
		.INIT('he)
	) name3849 (
		_w4309_,
		_w4311_,
		_w4312_
	);
	LUT2 #(
		.INIT('h2)
	) name3850 (
		\P1_reg0_reg[18]/NET0131 ,
		_w511_,
		_w4313_
	);
	LUT2 #(
		.INIT('h8)
	) name3851 (
		\P1_reg0_reg[18]/NET0131 ,
		_w524_,
		_w4314_
	);
	LUT4 #(
		.INIT('haaa8)
	) name3852 (
		\P1_reg0_reg[18]/NET0131 ,
		_w528_,
		_w530_,
		_w533_,
		_w4315_
	);
	LUT4 #(
		.INIT('h4484)
	) name3853 (
		_w1423_,
		_w2688_,
		_w3080_,
		_w3469_,
		_w4316_
	);
	LUT3 #(
		.INIT('ha2)
	) name3854 (
		\P1_reg0_reg[18]/NET0131 ,
		_w2692_,
		_w3005_,
		_w4317_
	);
	LUT4 #(
		.INIT('h0057)
	) name3855 (
		_w2688_,
		_w3897_,
		_w3898_,
		_w4317_,
		_w4318_
	);
	LUT4 #(
		.INIT('h5700)
	) name3856 (
		_w1286_,
		_w4315_,
		_w4316_,
		_w4318_,
		_w4319_
	);
	LUT4 #(
		.INIT('h8848)
	) name3857 (
		_w1423_,
		_w2688_,
		_w3046_,
		_w3476_,
		_w4320_
	);
	LUT3 #(
		.INIT('ha8)
	) name3858 (
		_w1114_,
		_w4315_,
		_w4320_,
		_w4321_
	);
	LUT4 #(
		.INIT('h7020)
	) name3859 (
		_w537_,
		_w722_,
		_w2688_,
		_w3479_,
		_w4322_
	);
	LUT3 #(
		.INIT('ha8)
	) name3860 (
		_w1183_,
		_w4315_,
		_w4322_,
		_w4323_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name3861 (
		_w526_,
		_w4321_,
		_w4323_,
		_w4319_,
		_w4324_
	);
	LUT4 #(
		.INIT('heeec)
	) name3862 (
		\P1_state_reg[0]/NET0131 ,
		_w4313_,
		_w4314_,
		_w4324_,
		_w4325_
	);
	LUT2 #(
		.INIT('h2)
	) name3863 (
		\P1_reg0_reg[19]/NET0131 ,
		_w511_,
		_w4326_
	);
	LUT2 #(
		.INIT('h8)
	) name3864 (
		\P1_reg0_reg[19]/NET0131 ,
		_w524_,
		_w4327_
	);
	LUT4 #(
		.INIT('haaa8)
	) name3865 (
		\P1_reg0_reg[19]/NET0131 ,
		_w528_,
		_w530_,
		_w533_,
		_w4328_
	);
	LUT4 #(
		.INIT('h7020)
	) name3866 (
		_w537_,
		_w745_,
		_w2688_,
		_w3710_,
		_w4329_
	);
	LUT3 #(
		.INIT('ha8)
	) name3867 (
		_w1183_,
		_w4328_,
		_w4329_,
		_w4330_
	);
	LUT4 #(
		.INIT('hc535)
	) name3868 (
		\P1_reg0_reg[19]/NET0131 ,
		_w1422_,
		_w2688_,
		_w2848_,
		_w4331_
	);
	LUT2 #(
		.INIT('h2)
	) name3869 (
		_w1286_,
		_w4331_,
		_w4332_
	);
	LUT4 #(
		.INIT('h35c5)
	) name3870 (
		\P1_reg0_reg[19]/NET0131 ,
		_w1422_,
		_w2688_,
		_w2876_,
		_w4333_
	);
	LUT4 #(
		.INIT('h35c5)
	) name3871 (
		\P1_reg0_reg[19]/NET0131 ,
		_w674_,
		_w2688_,
		_w3130_,
		_w4334_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name3872 (
		\P1_reg0_reg[19]/NET0131 ,
		_w1138_,
		_w2425_,
		_w2688_,
		_w4335_
	);
	LUT3 #(
		.INIT('h07)
	) name3873 (
		_w2688_,
		_w3717_,
		_w4335_,
		_w4336_
	);
	LUT3 #(
		.INIT('hd0)
	) name3874 (
		_w1136_,
		_w4334_,
		_w4336_,
		_w4337_
	);
	LUT3 #(
		.INIT('hd0)
	) name3875 (
		_w1114_,
		_w4333_,
		_w4337_,
		_w4338_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name3876 (
		_w526_,
		_w4330_,
		_w4332_,
		_w4338_,
		_w4339_
	);
	LUT4 #(
		.INIT('heeec)
	) name3877 (
		\P1_state_reg[0]/NET0131 ,
		_w4326_,
		_w4327_,
		_w4339_,
		_w4340_
	);
	LUT2 #(
		.INIT('h2)
	) name3878 (
		\P1_reg0_reg[22]/NET0131 ,
		_w511_,
		_w4341_
	);
	LUT2 #(
		.INIT('h8)
	) name3879 (
		\P1_reg0_reg[22]/NET0131 ,
		_w524_,
		_w4342_
	);
	LUT4 #(
		.INIT('haaa8)
	) name3880 (
		\P1_reg0_reg[22]/NET0131 ,
		_w528_,
		_w530_,
		_w533_,
		_w4343_
	);
	LUT4 #(
		.INIT('hddd1)
	) name3881 (
		\P1_reg0_reg[22]/NET0131 ,
		_w2688_,
		_w3775_,
		_w3776_,
		_w4344_
	);
	LUT4 #(
		.INIT('h4844)
	) name3882 (
		_w1457_,
		_w2688_,
		_w3778_,
		_w3780_,
		_w4345_
	);
	LUT3 #(
		.INIT('ha8)
	) name3883 (
		_w1114_,
		_w4343_,
		_w4345_,
		_w4346_
	);
	LUT4 #(
		.INIT('h8488)
	) name3884 (
		_w1457_,
		_w2688_,
		_w3783_,
		_w3785_,
		_w4347_
	);
	LUT3 #(
		.INIT('ha2)
	) name3885 (
		\P1_reg0_reg[22]/NET0131 ,
		_w2692_,
		_w3005_,
		_w4348_
	);
	LUT4 #(
		.INIT('h007b)
	) name3886 (
		_w1066_,
		_w1136_,
		_w3546_,
		_w3951_,
		_w4349_
	);
	LUT3 #(
		.INIT('h31)
	) name3887 (
		_w2688_,
		_w4348_,
		_w4349_,
		_w4350_
	);
	LUT4 #(
		.INIT('h5700)
	) name3888 (
		_w1286_,
		_w4343_,
		_w4347_,
		_w4350_,
		_w4351_
	);
	LUT4 #(
		.INIT('h0d00)
	) name3889 (
		_w1183_,
		_w4344_,
		_w4346_,
		_w4351_,
		_w4352_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name3890 (
		\P1_state_reg[0]/NET0131 ,
		_w526_,
		_w4342_,
		_w4352_,
		_w4353_
	);
	LUT2 #(
		.INIT('he)
	) name3891 (
		_w4341_,
		_w4353_,
		_w4354_
	);
	LUT2 #(
		.INIT('h2)
	) name3892 (
		\P1_reg0_reg[23]/NET0131 ,
		_w511_,
		_w4355_
	);
	LUT2 #(
		.INIT('h8)
	) name3893 (
		\P1_reg0_reg[23]/NET0131 ,
		_w524_,
		_w4356_
	);
	LUT4 #(
		.INIT('haaa2)
	) name3894 (
		\P1_reg0_reg[23]/NET0131 ,
		_w2692_,
		_w3005_,
		_w3664_,
		_w4357_
	);
	LUT4 #(
		.INIT('h005d)
	) name3895 (
		_w2688_,
		_w3763_,
		_w4275_,
		_w4357_,
		_w4358_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name3896 (
		\P1_state_reg[0]/NET0131 ,
		_w526_,
		_w4356_,
		_w4358_,
		_w4359_
	);
	LUT2 #(
		.INIT('he)
	) name3897 (
		_w4355_,
		_w4359_,
		_w4360_
	);
	LUT2 #(
		.INIT('h2)
	) name3898 (
		\P1_reg0_reg[30]/NET0131 ,
		_w511_,
		_w4361_
	);
	LUT4 #(
		.INIT('h3c55)
	) name3899 (
		\P1_reg0_reg[30]/NET0131 ,
		_w1133_,
		_w1312_,
		_w2688_,
		_w4362_
	);
	LUT2 #(
		.INIT('h2)
	) name3900 (
		_w1136_,
		_w4362_,
		_w4363_
	);
	LUT4 #(
		.INIT('h0a2a)
	) name3901 (
		\P1_reg0_reg[30]/NET0131 ,
		_w1107_,
		_w2425_,
		_w2688_,
		_w4364_
	);
	LUT4 #(
		.INIT('hfc55)
	) name3902 (
		\P1_reg0_reg[30]/NET0131 ,
		_w541_,
		_w1311_,
		_w2688_,
		_w4365_
	);
	LUT3 #(
		.INIT('h31)
	) name3903 (
		_w1138_,
		_w4364_,
		_w4365_,
		_w4366_
	);
	LUT3 #(
		.INIT('h70)
	) name3904 (
		_w3286_,
		_w3675_,
		_w4366_,
		_w4367_
	);
	LUT2 #(
		.INIT('h8)
	) name3905 (
		\P1_reg0_reg[30]/NET0131 ,
		_w524_,
		_w4368_
	);
	LUT4 #(
		.INIT('h0075)
	) name3906 (
		_w526_,
		_w4363_,
		_w4367_,
		_w4368_,
		_w4369_
	);
	LUT3 #(
		.INIT('hce)
	) name3907 (
		\P1_state_reg[0]/NET0131 ,
		_w4361_,
		_w4369_,
		_w4370_
	);
	LUT4 #(
		.INIT('h80cc)
	) name3908 (
		_w1183_,
		_w3651_,
		_w3730_,
		_w4250_,
		_w4371_
	);
	LUT4 #(
		.INIT('h0020)
	) name3909 (
		_w2692_,
		_w3005_,
		_w3443_,
		_w3664_,
		_w4372_
	);
	LUT2 #(
		.INIT('h2)
	) name3910 (
		\P1_reg0_reg[8]/NET0131 ,
		_w4372_,
		_w4373_
	);
	LUT2 #(
		.INIT('he)
	) name3911 (
		_w4371_,
		_w4373_,
		_w4374_
	);
	LUT4 #(
		.INIT('haaa8)
	) name3912 (
		\P1_reg0_reg[9]/NET0131 ,
		_w528_,
		_w530_,
		_w533_,
		_w4375_
	);
	LUT4 #(
		.INIT('h7020)
	) name3913 (
		_w537_,
		_w903_,
		_w3651_,
		_w4212_,
		_w4376_
	);
	LUT2 #(
		.INIT('h2)
	) name3914 (
		\P1_reg0_reg[9]/NET0131 ,
		_w3658_,
		_w4377_
	);
	LUT4 #(
		.INIT('h00d5)
	) name3915 (
		_w3651_,
		_w4215_,
		_w4256_,
		_w4377_,
		_w4378_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name3916 (
		_w1183_,
		_w4375_,
		_w4376_,
		_w4378_,
		_w4379_
	);
	LUT2 #(
		.INIT('h2)
	) name3917 (
		\P1_reg1_reg[18]/NET0131 ,
		_w511_,
		_w4380_
	);
	LUT2 #(
		.INIT('h8)
	) name3918 (
		\P1_reg1_reg[18]/NET0131 ,
		_w524_,
		_w4381_
	);
	LUT4 #(
		.INIT('haa02)
	) name3919 (
		\P1_reg1_reg[18]/NET0131 ,
		_w528_,
		_w530_,
		_w533_,
		_w4382_
	);
	LUT4 #(
		.INIT('h4484)
	) name3920 (
		_w1423_,
		_w2421_,
		_w3080_,
		_w3469_,
		_w4383_
	);
	LUT2 #(
		.INIT('h2)
	) name3921 (
		\P1_reg1_reg[18]/NET0131 ,
		_w3026_,
		_w4384_
	);
	LUT4 #(
		.INIT('h0057)
	) name3922 (
		_w2421_,
		_w3897_,
		_w3898_,
		_w4384_,
		_w4385_
	);
	LUT4 #(
		.INIT('h5700)
	) name3923 (
		_w1286_,
		_w4382_,
		_w4383_,
		_w4385_,
		_w4386_
	);
	LUT4 #(
		.INIT('h8848)
	) name3924 (
		_w1423_,
		_w2421_,
		_w3046_,
		_w3476_,
		_w4387_
	);
	LUT3 #(
		.INIT('ha8)
	) name3925 (
		_w1114_,
		_w4382_,
		_w4387_,
		_w4388_
	);
	LUT4 #(
		.INIT('h7020)
	) name3926 (
		_w537_,
		_w722_,
		_w2421_,
		_w3479_,
		_w4389_
	);
	LUT3 #(
		.INIT('ha8)
	) name3927 (
		_w1183_,
		_w4382_,
		_w4389_,
		_w4390_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name3928 (
		_w526_,
		_w4388_,
		_w4390_,
		_w4386_,
		_w4391_
	);
	LUT4 #(
		.INIT('heeec)
	) name3929 (
		\P1_state_reg[0]/NET0131 ,
		_w4380_,
		_w4381_,
		_w4391_,
		_w4392_
	);
	LUT2 #(
		.INIT('h2)
	) name3930 (
		\P1_reg1_reg[19]/NET0131 ,
		_w511_,
		_w4393_
	);
	LUT2 #(
		.INIT('h8)
	) name3931 (
		\P1_reg1_reg[19]/NET0131 ,
		_w524_,
		_w4394_
	);
	LUT4 #(
		.INIT('haa02)
	) name3932 (
		\P1_reg1_reg[19]/NET0131 ,
		_w528_,
		_w530_,
		_w533_,
		_w4395_
	);
	LUT4 #(
		.INIT('h7020)
	) name3933 (
		_w537_,
		_w745_,
		_w2421_,
		_w3710_,
		_w4396_
	);
	LUT3 #(
		.INIT('ha8)
	) name3934 (
		_w1183_,
		_w4395_,
		_w4396_,
		_w4397_
	);
	LUT4 #(
		.INIT('hc535)
	) name3935 (
		\P1_reg1_reg[19]/NET0131 ,
		_w1422_,
		_w2421_,
		_w2848_,
		_w4398_
	);
	LUT2 #(
		.INIT('h2)
	) name3936 (
		_w1286_,
		_w4398_,
		_w4399_
	);
	LUT4 #(
		.INIT('h35c5)
	) name3937 (
		\P1_reg1_reg[19]/NET0131 ,
		_w1422_,
		_w2421_,
		_w2876_,
		_w4400_
	);
	LUT4 #(
		.INIT('h35c5)
	) name3938 (
		\P1_reg1_reg[19]/NET0131 ,
		_w674_,
		_w2421_,
		_w3130_,
		_w4401_
	);
	LUT4 #(
		.INIT('h08aa)
	) name3939 (
		\P1_reg1_reg[19]/NET0131 ,
		_w1138_,
		_w2421_,
		_w2425_,
		_w4402_
	);
	LUT3 #(
		.INIT('h07)
	) name3940 (
		_w2421_,
		_w3717_,
		_w4402_,
		_w4403_
	);
	LUT3 #(
		.INIT('hd0)
	) name3941 (
		_w1136_,
		_w4401_,
		_w4403_,
		_w4404_
	);
	LUT3 #(
		.INIT('hd0)
	) name3942 (
		_w1114_,
		_w4400_,
		_w4404_,
		_w4405_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name3943 (
		_w526_,
		_w4397_,
		_w4399_,
		_w4405_,
		_w4406_
	);
	LUT4 #(
		.INIT('heeec)
	) name3944 (
		\P1_state_reg[0]/NET0131 ,
		_w4393_,
		_w4394_,
		_w4406_,
		_w4407_
	);
	LUT4 #(
		.INIT('h0001)
	) name3945 (
		_w3751_,
		_w3754_,
		_w3762_,
		_w4275_,
		_w4408_
	);
	LUT3 #(
		.INIT('h8a)
	) name3946 (
		\P1_reg1_reg[23]/NET0131 ,
		_w3684_,
		_w4075_,
		_w4409_
	);
	LUT4 #(
		.INIT('haa02)
	) name3947 (
		\P1_reg1_reg[23]/NET0131 ,
		_w528_,
		_w530_,
		_w533_,
		_w4410_
	);
	LUT4 #(
		.INIT('h7200)
	) name3948 (
		_w537_,
		_w1070_,
		_w3756_,
		_w4074_,
		_w4411_
	);
	LUT4 #(
		.INIT('h1113)
	) name3949 (
		_w1183_,
		_w4409_,
		_w4410_,
		_w4411_,
		_w4412_
	);
	LUT3 #(
		.INIT('h2f)
	) name3950 (
		_w4074_,
		_w4408_,
		_w4412_,
		_w4413_
	);
	LUT2 #(
		.INIT('h2)
	) name3951 (
		\P1_reg1_reg[22]/NET0131 ,
		_w511_,
		_w4414_
	);
	LUT2 #(
		.INIT('h8)
	) name3952 (
		\P1_reg1_reg[22]/NET0131 ,
		_w524_,
		_w4415_
	);
	LUT4 #(
		.INIT('haa02)
	) name3953 (
		\P1_reg1_reg[22]/NET0131 ,
		_w528_,
		_w530_,
		_w533_,
		_w4416_
	);
	LUT4 #(
		.INIT('hddd1)
	) name3954 (
		\P1_reg1_reg[22]/NET0131 ,
		_w2421_,
		_w3775_,
		_w3776_,
		_w4417_
	);
	LUT4 #(
		.INIT('h4844)
	) name3955 (
		_w1457_,
		_w2421_,
		_w3778_,
		_w3780_,
		_w4418_
	);
	LUT3 #(
		.INIT('ha8)
	) name3956 (
		_w1114_,
		_w4416_,
		_w4418_,
		_w4419_
	);
	LUT4 #(
		.INIT('h8488)
	) name3957 (
		_w1457_,
		_w2421_,
		_w3783_,
		_w3785_,
		_w4420_
	);
	LUT2 #(
		.INIT('h2)
	) name3958 (
		\P1_reg1_reg[22]/NET0131 ,
		_w3026_,
		_w4421_
	);
	LUT3 #(
		.INIT('h0d)
	) name3959 (
		_w2421_,
		_w4349_,
		_w4421_,
		_w4422_
	);
	LUT4 #(
		.INIT('h5700)
	) name3960 (
		_w1286_,
		_w4416_,
		_w4420_,
		_w4422_,
		_w4423_
	);
	LUT4 #(
		.INIT('h0d00)
	) name3961 (
		_w1183_,
		_w4417_,
		_w4419_,
		_w4423_,
		_w4424_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name3962 (
		\P1_state_reg[0]/NET0131 ,
		_w526_,
		_w4415_,
		_w4424_,
		_w4425_
	);
	LUT2 #(
		.INIT('he)
	) name3963 (
		_w4414_,
		_w4425_,
		_w4426_
	);
	LUT2 #(
		.INIT('h2)
	) name3964 (
		\P1_reg1_reg[30]/NET0131 ,
		_w511_,
		_w4427_
	);
	LUT4 #(
		.INIT('h3c55)
	) name3965 (
		\P1_reg1_reg[30]/NET0131 ,
		_w1133_,
		_w1312_,
		_w2421_,
		_w4428_
	);
	LUT2 #(
		.INIT('h2)
	) name3966 (
		_w1136_,
		_w4428_,
		_w4429_
	);
	LUT4 #(
		.INIT('h02aa)
	) name3967 (
		\P1_reg1_reg[30]/NET0131 ,
		_w1107_,
		_w2421_,
		_w2425_,
		_w4430_
	);
	LUT4 #(
		.INIT('hfc55)
	) name3968 (
		\P1_reg1_reg[30]/NET0131 ,
		_w541_,
		_w1311_,
		_w2421_,
		_w4431_
	);
	LUT3 #(
		.INIT('h31)
	) name3969 (
		_w1138_,
		_w4430_,
		_w4431_,
		_w4432_
	);
	LUT3 #(
		.INIT('h70)
	) name3970 (
		_w3286_,
		_w3688_,
		_w4432_,
		_w4433_
	);
	LUT2 #(
		.INIT('h8)
	) name3971 (
		\P1_reg1_reg[30]/NET0131 ,
		_w524_,
		_w4434_
	);
	LUT4 #(
		.INIT('h0075)
	) name3972 (
		_w526_,
		_w4429_,
		_w4433_,
		_w4434_,
		_w4435_
	);
	LUT3 #(
		.INIT('hce)
	) name3973 (
		\P1_state_reg[0]/NET0131 ,
		_w4427_,
		_w4435_,
		_w4436_
	);
	LUT2 #(
		.INIT('h8)
	) name3974 (
		_w524_,
		_w796_,
		_w4437_
	);
	LUT4 #(
		.INIT('h1f00)
	) name3975 (
		_w528_,
		_w530_,
		_w533_,
		_w796_,
		_w4438_
	);
	LUT3 #(
		.INIT('h80)
	) name3976 (
		_w537_,
		_w817_,
		_w818_,
		_w4439_
	);
	LUT4 #(
		.INIT('h00eb)
	) name3977 (
		_w537_,
		_w808_,
		_w3340_,
		_w4439_,
		_w4440_
	);
	LUT4 #(
		.INIT('hc808)
	) name3978 (
		_w796_,
		_w1183_,
		_w2197_,
		_w4440_,
		_w4441_
	);
	LUT4 #(
		.INIT('h00b7)
	) name3979 (
		_w1453_,
		_w2197_,
		_w2843_,
		_w4438_,
		_w4442_
	);
	LUT2 #(
		.INIT('h2)
	) name3980 (
		_w1286_,
		_w4442_,
		_w4443_
	);
	LUT4 #(
		.INIT('h007b)
	) name3981 (
		_w1453_,
		_w2197_,
		_w2871_,
		_w4438_,
		_w4444_
	);
	LUT4 #(
		.INIT('h6a00)
	) name3982 (
		_w804_,
		_w1117_,
		_w1119_,
		_w1136_,
		_w4445_
	);
	LUT3 #(
		.INIT('h04)
	) name3983 (
		_w804_,
		_w2259_,
		_w2260_,
		_w4446_
	);
	LUT3 #(
		.INIT('h0d)
	) name3984 (
		_w796_,
		_w2860_,
		_w4446_,
		_w4447_
	);
	LUT3 #(
		.INIT('h70)
	) name3985 (
		_w2197_,
		_w4445_,
		_w4447_,
		_w4448_
	);
	LUT3 #(
		.INIT('hd0)
	) name3986 (
		_w1114_,
		_w4444_,
		_w4448_,
		_w4449_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name3987 (
		_w526_,
		_w4443_,
		_w4441_,
		_w4449_,
		_w4450_
	);
	LUT2 #(
		.INIT('h2)
	) name3988 (
		\P1_reg3_reg[11]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w4451_
	);
	LUT3 #(
		.INIT('h07)
	) name3989 (
		_w796_,
		_w1294_,
		_w4451_,
		_w4452_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name3990 (
		\P1_state_reg[0]/NET0131 ,
		_w4437_,
		_w4450_,
		_w4452_,
		_w4453_
	);
	LUT2 #(
		.INIT('h8)
	) name3991 (
		_w524_,
		_w749_,
		_w4454_
	);
	LUT4 #(
		.INIT('h1f00)
	) name3992 (
		_w528_,
		_w530_,
		_w533_,
		_w749_,
		_w4455_
	);
	LUT3 #(
		.INIT('h80)
	) name3993 (
		_w537_,
		_w805_,
		_w807_,
		_w4456_
	);
	LUT4 #(
		.INIT('h00eb)
	) name3994 (
		_w537_,
		_w762_,
		_w1161_,
		_w4456_,
		_w4457_
	);
	LUT4 #(
		.INIT('hc808)
	) name3995 (
		_w749_,
		_w1183_,
		_w2197_,
		_w4457_,
		_w4458_
	);
	LUT4 #(
		.INIT('h006f)
	) name3996 (
		_w954_,
		_w1443_,
		_w2197_,
		_w4455_,
		_w4459_
	);
	LUT2 #(
		.INIT('h2)
	) name3997 (
		_w1114_,
		_w4459_,
		_w4460_
	);
	LUT4 #(
		.INIT('hd200)
	) name3998 (
		_w1202_,
		_w1237_,
		_w1443_,
		_w2197_,
		_w4461_
	);
	LUT4 #(
		.INIT('h009f)
	) name3999 (
		_w758_,
		_w1120_,
		_w2197_,
		_w4455_,
		_w4462_
	);
	LUT3 #(
		.INIT('h04)
	) name4000 (
		_w758_,
		_w2259_,
		_w2260_,
		_w4463_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name4001 (
		_w749_,
		_w1138_,
		_w1141_,
		_w2197_,
		_w4464_
	);
	LUT2 #(
		.INIT('h1)
	) name4002 (
		_w4463_,
		_w4464_,
		_w4465_
	);
	LUT3 #(
		.INIT('hd0)
	) name4003 (
		_w1136_,
		_w4462_,
		_w4465_,
		_w4466_
	);
	LUT4 #(
		.INIT('h5700)
	) name4004 (
		_w1286_,
		_w4455_,
		_w4461_,
		_w4466_,
		_w4467_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name4005 (
		_w526_,
		_w4458_,
		_w4460_,
		_w4467_,
		_w4468_
	);
	LUT2 #(
		.INIT('h2)
	) name4006 (
		\P1_reg3_reg[13]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w4469_
	);
	LUT3 #(
		.INIT('h07)
	) name4007 (
		_w749_,
		_w1294_,
		_w4469_,
		_w4470_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name4008 (
		\P1_state_reg[0]/NET0131 ,
		_w4454_,
		_w4468_,
		_w4470_,
		_w4471_
	);
	LUT2 #(
		.INIT('h2)
	) name4009 (
		_w1487_,
		_w1617_,
		_w4472_
	);
	LUT4 #(
		.INIT('h001f)
	) name4010 (
		_w1491_,
		_w1493_,
		_w1496_,
		_w1617_,
		_w4473_
	);
	LUT4 #(
		.INIT('h7778)
	) name4011 (
		_w1616_,
		_w1618_,
		_w1638_,
		_w1640_,
		_w4474_
	);
	LUT4 #(
		.INIT('h8a20)
	) name4012 (
		_w2272_,
		_w2309_,
		_w2312_,
		_w4474_,
		_w4475_
	);
	LUT3 #(
		.INIT('h54)
	) name4013 (
		_w2276_,
		_w4473_,
		_w4475_,
		_w4476_
	);
	LUT4 #(
		.INIT('h070d)
	) name4014 (
		_w2272_,
		_w2363_,
		_w4473_,
		_w4474_,
		_w4477_
	);
	LUT3 #(
		.INIT('h04)
	) name4015 (
		_w1641_,
		_w2083_,
		_w2282_,
		_w4478_
	);
	LUT3 #(
		.INIT('h54)
	) name4016 (
		_w1617_,
		_w2086_,
		_w2280_,
		_w4479_
	);
	LUT2 #(
		.INIT('h1)
	) name4017 (
		_w4478_,
		_w4479_,
		_w4480_
	);
	LUT3 #(
		.INIT('he0)
	) name4018 (
		_w2192_,
		_w4477_,
		_w4480_,
		_w4481_
	);
	LUT4 #(
		.INIT('h00fe)
	) name4019 (
		_w1491_,
		_w1493_,
		_w1496_,
		_w1617_,
		_w4482_
	);
	LUT4 #(
		.INIT('h8a20)
	) name4020 (
		_w2277_,
		_w2309_,
		_w2312_,
		_w4474_,
		_w4483_
	);
	LUT3 #(
		.INIT('ha8)
	) name4021 (
		_w2290_,
		_w4482_,
		_w4483_,
		_w4484_
	);
	LUT3 #(
		.INIT('h70)
	) name4022 (
		_w1644_,
		_w1645_,
		_w2042_,
		_w4485_
	);
	LUT4 #(
		.INIT('h00de)
	) name4023 (
		_w1735_,
		_w2042_,
		_w4151_,
		_w4485_,
		_w4486_
	);
	LUT4 #(
		.INIT('h04c4)
	) name4024 (
		_w1617_,
		_w2081_,
		_w2277_,
		_w4486_,
		_w4487_
	);
	LUT4 #(
		.INIT('h0100)
	) name4025 (
		_w4476_,
		_w4484_,
		_w4487_,
		_w4481_,
		_w4488_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name4026 (
		\P1_state_reg[0]/NET0131 ,
		_w1489_,
		_w4472_,
		_w4488_,
		_w4489_
	);
	LUT2 #(
		.INIT('h4)
	) name4027 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[11]/NET0131 ,
		_w4490_
	);
	LUT4 #(
		.INIT('h0028)
	) name4028 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		_w1476_,
		_w1617_,
		_w4491_
	);
	LUT2 #(
		.INIT('h1)
	) name4029 (
		_w4490_,
		_w4491_,
		_w4492_
	);
	LUT2 #(
		.INIT('hb)
	) name4030 (
		_w4489_,
		_w4492_,
		_w4493_
	);
	LUT2 #(
		.INIT('h2)
	) name4031 (
		_w1487_,
		_w1718_,
		_w4494_
	);
	LUT4 #(
		.INIT('h001f)
	) name4032 (
		_w1491_,
		_w1493_,
		_w1496_,
		_w1718_,
		_w4495_
	);
	LUT2 #(
		.INIT('h9)
	) name4033 (
		_w1720_,
		_w1730_,
		_w4496_
	);
	LUT4 #(
		.INIT('h070d)
	) name4034 (
		_w2272_,
		_w2794_,
		_w4495_,
		_w4496_,
		_w4497_
	);
	LUT3 #(
		.INIT('h70)
	) name4035 (
		_w1747_,
		_w1750_,
		_w2042_,
		_w4498_
	);
	LUT4 #(
		.INIT('h00de)
	) name4036 (
		_w1697_,
		_w2042_,
		_w2066_,
		_w4498_,
		_w4499_
	);
	LUT4 #(
		.INIT('h04c4)
	) name4037 (
		_w1718_,
		_w2081_,
		_w2277_,
		_w4499_,
		_w4500_
	);
	LUT3 #(
		.INIT('h04)
	) name4038 (
		_w1730_,
		_w2083_,
		_w2282_,
		_w4501_
	);
	LUT3 #(
		.INIT('h54)
	) name4039 (
		_w1718_,
		_w2086_,
		_w2280_,
		_w4502_
	);
	LUT2 #(
		.INIT('h1)
	) name4040 (
		_w4501_,
		_w4502_,
		_w4503_
	);
	LUT2 #(
		.INIT('h4)
	) name4041 (
		_w4500_,
		_w4503_,
		_w4504_
	);
	LUT3 #(
		.INIT('he0)
	) name4042 (
		_w2192_,
		_w4497_,
		_w4504_,
		_w4505_
	);
	LUT4 #(
		.INIT('hb04f)
	) name4043 (
		_w2467_,
		_w2468_,
		_w2469_,
		_w4496_,
		_w4506_
	);
	LUT4 #(
		.INIT('h10d0)
	) name4044 (
		_w1718_,
		_w2277_,
		_w2290_,
		_w4506_,
		_w4507_
	);
	LUT4 #(
		.INIT('h010d)
	) name4045 (
		_w1718_,
		_w2272_,
		_w2276_,
		_w4506_,
		_w4508_
	);
	LUT2 #(
		.INIT('h1)
	) name4046 (
		_w4507_,
		_w4508_,
		_w4509_
	);
	LUT4 #(
		.INIT('h3111)
	) name4047 (
		_w1489_,
		_w4494_,
		_w4505_,
		_w4509_,
		_w4510_
	);
	LUT2 #(
		.INIT('h4)
	) name4048 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[14]/NET0131 ,
		_w4511_
	);
	LUT3 #(
		.INIT('h0b)
	) name4049 (
		_w1718_,
		_w2293_,
		_w4511_,
		_w4512_
	);
	LUT3 #(
		.INIT('h2f)
	) name4050 (
		\P1_state_reg[0]/NET0131 ,
		_w4510_,
		_w4512_,
		_w4513_
	);
	LUT2 #(
		.INIT('h2)
	) name4051 (
		_w1487_,
		_w1693_,
		_w4514_
	);
	LUT4 #(
		.INIT('h00fe)
	) name4052 (
		_w1491_,
		_w1493_,
		_w1496_,
		_w1693_,
		_w4515_
	);
	LUT2 #(
		.INIT('h6)
	) name4053 (
		_w1697_,
		_w1715_,
		_w4516_
	);
	LUT4 #(
		.INIT('h007d)
	) name4054 (
		_w2277_,
		_w3512_,
		_w4516_,
		_w4515_,
		_w4517_
	);
	LUT2 #(
		.INIT('h2)
	) name4055 (
		_w2290_,
		_w4517_,
		_w4518_
	);
	LUT4 #(
		.INIT('h001f)
	) name4056 (
		_w1491_,
		_w1493_,
		_w1496_,
		_w1693_,
		_w4519_
	);
	LUT4 #(
		.INIT('h070d)
	) name4057 (
		_w2272_,
		_w3512_,
		_w4519_,
		_w4516_,
		_w4520_
	);
	LUT4 #(
		.INIT('hd02f)
	) name4058 (
		_w2368_,
		_w2363_,
		_w2373_,
		_w4516_,
		_w4521_
	);
	LUT4 #(
		.INIT('h0131)
	) name4059 (
		_w1693_,
		_w2192_,
		_w2272_,
		_w4521_,
		_w4522_
	);
	LUT3 #(
		.INIT('h70)
	) name4060 (
		_w1717_,
		_w1719_,
		_w2042_,
		_w4523_
	);
	LUT4 #(
		.INIT('h0e0f)
	) name4061 (
		_w498_,
		_w1697_,
		_w2042_,
		_w2066_,
		_w4524_
	);
	LUT4 #(
		.INIT('h0605)
	) name4062 (
		_w498_,
		_w1697_,
		_w2042_,
		_w2066_,
		_w4525_
	);
	LUT4 #(
		.INIT('h1113)
	) name4063 (
		_w2277_,
		_w4515_,
		_w4523_,
		_w4525_,
		_w4526_
	);
	LUT3 #(
		.INIT('h04)
	) name4064 (
		_w1715_,
		_w2083_,
		_w2282_,
		_w4527_
	);
	LUT3 #(
		.INIT('h54)
	) name4065 (
		_w1693_,
		_w2086_,
		_w2280_,
		_w4528_
	);
	LUT2 #(
		.INIT('h1)
	) name4066 (
		_w4527_,
		_w4528_,
		_w4529_
	);
	LUT3 #(
		.INIT('hd0)
	) name4067 (
		_w2081_,
		_w4526_,
		_w4529_,
		_w4530_
	);
	LUT4 #(
		.INIT('h0e00)
	) name4068 (
		_w2276_,
		_w4520_,
		_w4522_,
		_w4530_,
		_w4531_
	);
	LUT4 #(
		.INIT('h1311)
	) name4069 (
		_w1489_,
		_w4514_,
		_w4518_,
		_w4531_,
		_w4532_
	);
	LUT2 #(
		.INIT('h4)
	) name4070 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[15]/NET0131 ,
		_w4533_
	);
	LUT3 #(
		.INIT('h0b)
	) name4071 (
		_w1693_,
		_w2293_,
		_w4533_,
		_w4534_
	);
	LUT3 #(
		.INIT('h2f)
	) name4072 (
		\P1_state_reg[0]/NET0131 ,
		_w4532_,
		_w4534_,
		_w4535_
	);
	LUT3 #(
		.INIT('h04)
	) name4073 (
		_w894_,
		_w2259_,
		_w2260_,
		_w4536_
	);
	LUT4 #(
		.INIT('h1e0f)
	) name4074 (
		_w876_,
		_w887_,
		_w934_,
		_w1153_,
		_w4537_
	);
	LUT4 #(
		.INIT('h7020)
	) name4075 (
		_w537_,
		_w876_,
		_w1183_,
		_w4537_,
		_w4538_
	);
	LUT4 #(
		.INIT('h780f)
	) name4076 (
		_w871_,
		_w883_,
		_w1440_,
		_w2220_,
		_w4539_
	);
	LUT2 #(
		.INIT('h2)
	) name4077 (
		_w1114_,
		_w4539_,
		_w4540_
	);
	LUT4 #(
		.INIT('h0df2)
	) name4078 (
		_w1214_,
		_w1360_,
		_w1361_,
		_w1440_,
		_w4541_
	);
	LUT3 #(
		.INIT('h60)
	) name4079 (
		_w894_,
		_w1115_,
		_w1136_,
		_w4542_
	);
	LUT3 #(
		.INIT('h07)
	) name4080 (
		_w1286_,
		_w4541_,
		_w4542_,
		_w4543_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name4081 (
		_w2197_,
		_w4540_,
		_w4538_,
		_w4543_,
		_w4544_
	);
	LUT4 #(
		.INIT('h3130)
	) name4082 (
		_w1136_,
		_w1141_,
		_w2197_,
		_w3118_,
		_w4545_
	);
	LUT3 #(
		.INIT('h51)
	) name4083 (
		_w523_,
		_w1183_,
		_w2197_,
		_w4546_
	);
	LUT4 #(
		.INIT('h5900)
	) name4084 (
		\P1_IR_reg[23]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		_w509_,
		_w885_,
		_w4547_
	);
	LUT3 #(
		.INIT('h70)
	) name4085 (
		_w4545_,
		_w4546_,
		_w4547_,
		_w4548_
	);
	LUT4 #(
		.INIT('h0057)
	) name4086 (
		_w526_,
		_w4536_,
		_w4544_,
		_w4548_,
		_w4549_
	);
	LUT3 #(
		.INIT('h6c)
	) name4087 (
		\P1_reg3_reg[3]/NET0131 ,
		\P1_reg3_reg[4]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w4550_
	);
	LUT2 #(
		.INIT('h4)
	) name4088 (
		_w511_,
		_w4550_,
		_w4551_
	);
	LUT3 #(
		.INIT('hf2)
	) name4089 (
		\P1_state_reg[0]/NET0131 ,
		_w4549_,
		_w4551_,
		_w4552_
	);
	LUT2 #(
		.INIT('h8)
	) name4090 (
		_w524_,
		_w931_,
		_w4553_
	);
	LUT3 #(
		.INIT('h80)
	) name4091 (
		_w537_,
		_w884_,
		_w886_,
		_w4554_
	);
	LUT4 #(
		.INIT('h00eb)
	) name4092 (
		_w537_,
		_w924_,
		_w1154_,
		_w4554_,
		_w4555_
	);
	LUT4 #(
		.INIT('h001f)
	) name4093 (
		_w528_,
		_w530_,
		_w533_,
		_w931_,
		_w4556_
	);
	LUT2 #(
		.INIT('h2)
	) name4094 (
		_w1183_,
		_w4556_,
		_w4557_
	);
	LUT3 #(
		.INIT('hd0)
	) name4095 (
		_w2197_,
		_w4555_,
		_w4557_,
		_w4558_
	);
	LUT4 #(
		.INIT('h00b0)
	) name4096 (
		_w872_,
		_w896_,
		_w899_,
		_w1449_,
		_w4559_
	);
	LUT4 #(
		.INIT('h4f00)
	) name4097 (
		_w872_,
		_w896_,
		_w899_,
		_w1449_,
		_w4560_
	);
	LUT3 #(
		.INIT('h02)
	) name4098 (
		_w1114_,
		_w4560_,
		_w4559_,
		_w4561_
	);
	LUT4 #(
		.INIT('h6c00)
	) name4099 (
		_w894_,
		_w938_,
		_w1115_,
		_w1136_,
		_w4562_
	);
	LUT4 #(
		.INIT('h00b7)
	) name4100 (
		_w1220_,
		_w1286_,
		_w1449_,
		_w4562_,
		_w4563_
	);
	LUT3 #(
		.INIT('h04)
	) name4101 (
		_w938_,
		_w2259_,
		_w2260_,
		_w4564_
	);
	LUT3 #(
		.INIT('h0d)
	) name4102 (
		_w931_,
		_w4545_,
		_w4564_,
		_w4565_
	);
	LUT4 #(
		.INIT('h7500)
	) name4103 (
		_w2197_,
		_w4561_,
		_w4563_,
		_w4565_,
		_w4566_
	);
	LUT4 #(
		.INIT('h1311)
	) name4104 (
		_w526_,
		_w4553_,
		_w4558_,
		_w4566_,
		_w4567_
	);
	LUT2 #(
		.INIT('h2)
	) name4105 (
		\P1_reg3_reg[5]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w4568_
	);
	LUT3 #(
		.INIT('h07)
	) name4106 (
		_w931_,
		_w1294_,
		_w4568_,
		_w4569_
	);
	LUT3 #(
		.INIT('h2f)
	) name4107 (
		\P1_state_reg[0]/NET0131 ,
		_w4567_,
		_w4569_,
		_w4570_
	);
	LUT2 #(
		.INIT('h4)
	) name4108 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[8]/NET0131 ,
		_w4571_
	);
	LUT4 #(
		.INIT('h001f)
	) name4109 (
		_w1491_,
		_w1493_,
		_w1496_,
		_w1674_,
		_w4572_
	);
	LUT2 #(
		.INIT('h9)
	) name4110 (
		_w1676_,
		_w1684_,
		_w4573_
	);
	LUT4 #(
		.INIT('h708f)
	) name4111 (
		_w1547_,
		_w1608_,
		_w1615_,
		_w4573_,
		_w4574_
	);
	LUT4 #(
		.INIT('h010d)
	) name4112 (
		_w1674_,
		_w2272_,
		_w2276_,
		_w4574_,
		_w4575_
	);
	LUT3 #(
		.INIT('h70)
	) name4113 (
		_w1529_,
		_w1531_,
		_w2042_,
		_w4576_
	);
	LUT4 #(
		.INIT('h00de)
	) name4114 (
		_w1663_,
		_w2042_,
		_w4149_,
		_w4576_,
		_w4577_
	);
	LUT4 #(
		.INIT('h04c4)
	) name4115 (
		_w1674_,
		_w2081_,
		_w2277_,
		_w4577_,
		_w4578_
	);
	LUT4 #(
		.INIT('h3050)
	) name4116 (
		_w1674_,
		_w1684_,
		_w2084_,
		_w2272_,
		_w4579_
	);
	LUT4 #(
		.INIT('h3332)
	) name4117 (
		_w1487_,
		_w1674_,
		_w2086_,
		_w2293_,
		_w4580_
	);
	LUT4 #(
		.INIT('hf100)
	) name4118 (
		_w1509_,
		_w1681_,
		_w1683_,
		_w2088_,
		_w4581_
	);
	LUT2 #(
		.INIT('h1)
	) name4119 (
		_w4580_,
		_w4581_,
		_w4582_
	);
	LUT2 #(
		.INIT('h4)
	) name4120 (
		_w4579_,
		_w4582_,
		_w4583_
	);
	LUT3 #(
		.INIT('h10)
	) name4121 (
		_w4575_,
		_w4578_,
		_w4583_,
		_w4584_
	);
	LUT4 #(
		.INIT('h10d0)
	) name4122 (
		_w1674_,
		_w2277_,
		_w2290_,
		_w4574_,
		_w4585_
	);
	LUT4 #(
		.INIT('h070b)
	) name4123 (
		_w2124_,
		_w2272_,
		_w4572_,
		_w4573_,
		_w4586_
	);
	LUT3 #(
		.INIT('h32)
	) name4124 (
		_w2192_,
		_w4585_,
		_w4586_,
		_w4587_
	);
	LUT3 #(
		.INIT('h8a)
	) name4125 (
		\P1_state_reg[0]/NET0131 ,
		_w1489_,
		_w1674_,
		_w4588_
	);
	LUT4 #(
		.INIT('hbfaa)
	) name4126 (
		_w4571_,
		_w4584_,
		_w4587_,
		_w4588_,
		_w4589_
	);
	LUT4 #(
		.INIT('h70d0)
	) name4127 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg0_reg[16]/NET0131 ,
		_w1476_,
		_w4590_
	);
	LUT2 #(
		.INIT('h8)
	) name4128 (
		\P2_reg0_reg[16]/NET0131 ,
		_w1487_,
		_w4591_
	);
	LUT4 #(
		.INIT('h02aa)
	) name4129 (
		\P2_reg0_reg[16]/NET0131 ,
		_w1491_,
		_w1493_,
		_w1496_,
		_w4592_
	);
	LUT4 #(
		.INIT('haa56)
	) name4130 (
		_w498_,
		_w1509_,
		_w1790_,
		_w1794_,
		_w4593_
	);
	LUT4 #(
		.INIT('h4f00)
	) name4131 (
		_w1687_,
		_w1692_,
		_w1763_,
		_w1847_,
		_w4594_
	);
	LUT4 #(
		.INIT('h1dd1)
	) name4132 (
		\P2_reg0_reg[16]/NET0131 ,
		_w2272_,
		_w4593_,
		_w4594_,
		_w4595_
	);
	LUT2 #(
		.INIT('h2)
	) name4133 (
		_w2290_,
		_w4595_,
		_w4596_
	);
	LUT4 #(
		.INIT('h1dd1)
	) name4134 (
		\P2_reg0_reg[16]/NET0131 ,
		_w2277_,
		_w4593_,
		_w4594_,
		_w4597_
	);
	LUT2 #(
		.INIT('h1)
	) name4135 (
		_w2276_,
		_w4597_,
		_w4598_
	);
	LUT4 #(
		.INIT('hbf00)
	) name4136 (
		_w2124_,
		_w2126_,
		_w2130_,
		_w2448_,
		_w4599_
	);
	LUT4 #(
		.INIT('hd11d)
	) name4137 (
		\P2_reg0_reg[16]/NET0131 ,
		_w2277_,
		_w4593_,
		_w4599_,
		_w4600_
	);
	LUT2 #(
		.INIT('h4)
	) name4138 (
		_w498_,
		_w1781_,
		_w4601_
	);
	LUT4 #(
		.INIT('h5444)
	) name4139 (
		_w1697_,
		_w2042_,
		_w2066_,
		_w4601_,
		_w4602_
	);
	LUT4 #(
		.INIT('hcc40)
	) name4140 (
		_w1781_,
		_w2272_,
		_w4524_,
		_w4602_,
		_w4603_
	);
	LUT3 #(
		.INIT('ha2)
	) name4141 (
		\P2_reg0_reg[16]/NET0131 ,
		_w2633_,
		_w2634_,
		_w4604_
	);
	LUT4 #(
		.INIT('hf100)
	) name4142 (
		_w1509_,
		_w1790_,
		_w1794_,
		_w2920_,
		_w4605_
	);
	LUT2 #(
		.INIT('h1)
	) name4143 (
		_w4604_,
		_w4605_,
		_w4606_
	);
	LUT4 #(
		.INIT('h5700)
	) name4144 (
		_w2081_,
		_w4592_,
		_w4603_,
		_w4606_,
		_w4607_
	);
	LUT3 #(
		.INIT('he0)
	) name4145 (
		_w2192_,
		_w4600_,
		_w4607_,
		_w4608_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name4146 (
		_w1489_,
		_w4598_,
		_w4596_,
		_w4608_,
		_w4609_
	);
	LUT4 #(
		.INIT('heeec)
	) name4147 (
		\P1_state_reg[0]/NET0131 ,
		_w4590_,
		_w4591_,
		_w4609_,
		_w4610_
	);
	LUT2 #(
		.INIT('h2)
	) name4148 (
		\P1_reg2_reg[10]/NET0131 ,
		_w511_,
		_w4611_
	);
	LUT2 #(
		.INIT('h8)
	) name4149 (
		\P1_reg2_reg[10]/NET0131 ,
		_w524_,
		_w4612_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name4150 (
		\P1_reg2_reg[10]/NET0131 ,
		_w528_,
		_w530_,
		_w533_,
		_w4613_
	);
	LUT4 #(
		.INIT('h2a08)
	) name4151 (
		_w534_,
		_w537_,
		_w833_,
		_w4084_,
		_w4614_
	);
	LUT3 #(
		.INIT('ha8)
	) name4152 (
		_w1183_,
		_w4613_,
		_w4614_,
		_w4615_
	);
	LUT4 #(
		.INIT('h1dd1)
	) name4153 (
		\P1_reg2_reg[10]/NET0131 ,
		_w534_,
		_w1438_,
		_w3076_,
		_w4616_
	);
	LUT2 #(
		.INIT('h2)
	) name4154 (
		_w1286_,
		_w4616_,
		_w4617_
	);
	LUT4 #(
		.INIT('hd11d)
	) name4155 (
		\P1_reg2_reg[10]/NET0131 ,
		_w534_,
		_w1438_,
		_w3052_,
		_w4618_
	);
	LUT4 #(
		.INIT('he020)
	) name4156 (
		\P1_reg2_reg[10]/NET0131 ,
		_w534_,
		_w1136_,
		_w4090_,
		_w4619_
	);
	LUT4 #(
		.INIT('haa20)
	) name4157 (
		\P1_reg2_reg[10]/NET0131 ,
		_w534_,
		_w1138_,
		_w1141_,
		_w4620_
	);
	LUT3 #(
		.INIT('h20)
	) name4158 (
		_w534_,
		_w827_,
		_w1138_,
		_w4621_
	);
	LUT2 #(
		.INIT('h8)
	) name4159 (
		_w816_,
		_w1143_,
		_w4622_
	);
	LUT3 #(
		.INIT('h01)
	) name4160 (
		_w4621_,
		_w4622_,
		_w4620_,
		_w4623_
	);
	LUT2 #(
		.INIT('h4)
	) name4161 (
		_w4619_,
		_w4623_,
		_w4624_
	);
	LUT3 #(
		.INIT('hd0)
	) name4162 (
		_w1114_,
		_w4618_,
		_w4624_,
		_w4625_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name4163 (
		_w526_,
		_w4615_,
		_w4617_,
		_w4625_,
		_w4626_
	);
	LUT4 #(
		.INIT('heeec)
	) name4164 (
		\P1_state_reg[0]/NET0131 ,
		_w4611_,
		_w4612_,
		_w4626_,
		_w4627_
	);
	LUT2 #(
		.INIT('h8)
	) name4165 (
		_w749_,
		_w1143_,
		_w4628_
	);
	LUT2 #(
		.INIT('h8)
	) name4166 (
		_w1183_,
		_w4457_,
		_w4629_
	);
	LUT3 #(
		.INIT('h84)
	) name4167 (
		_w954_,
		_w1114_,
		_w1443_,
		_w4630_
	);
	LUT4 #(
		.INIT('hd020)
	) name4168 (
		_w1202_,
		_w1237_,
		_w1286_,
		_w1443_,
		_w4631_
	);
	LUT2 #(
		.INIT('h4)
	) name4169 (
		_w758_,
		_w1138_,
		_w4632_
	);
	LUT4 #(
		.INIT('h009f)
	) name4170 (
		_w758_,
		_w1120_,
		_w1136_,
		_w4632_,
		_w4633_
	);
	LUT3 #(
		.INIT('h10)
	) name4171 (
		_w4631_,
		_w4630_,
		_w4633_,
		_w4634_
	);
	LUT4 #(
		.INIT('h1311)
	) name4172 (
		_w534_,
		_w4628_,
		_w4629_,
		_w4634_,
		_w4635_
	);
	LUT3 #(
		.INIT('h2a)
	) name4173 (
		\P1_reg2_reg[13]/NET0131 ,
		_w3443_,
		_w3603_,
		_w4636_
	);
	LUT3 #(
		.INIT('hf2)
	) name4174 (
		_w3443_,
		_w4635_,
		_w4636_,
		_w4637_
	);
	LUT2 #(
		.INIT('h2)
	) name4175 (
		\P1_reg2_reg[14]/NET0131 ,
		_w511_,
		_w4638_
	);
	LUT2 #(
		.INIT('h8)
	) name4176 (
		\P1_reg2_reg[14]/NET0131 ,
		_w524_,
		_w4639_
	);
	LUT4 #(
		.INIT('hddd1)
	) name4177 (
		\P1_reg2_reg[14]/NET0131 ,
		_w534_,
		_w4103_,
		_w4104_,
		_w4640_
	);
	LUT2 #(
		.INIT('h2)
	) name4178 (
		_w1183_,
		_w4640_,
		_w4641_
	);
	LUT4 #(
		.INIT('he020)
	) name4179 (
		\P1_reg2_reg[14]/NET0131 ,
		_w534_,
		_w1286_,
		_w4107_,
		_w4642_
	);
	LUT4 #(
		.INIT('h20e0)
	) name4180 (
		\P1_reg2_reg[14]/NET0131 ,
		_w534_,
		_w1114_,
		_w4109_,
		_w4643_
	);
	LUT2 #(
		.INIT('h4)
	) name4181 (
		_w767_,
		_w1138_,
		_w4644_
	);
	LUT4 #(
		.INIT('h6c00)
	) name4182 (
		_w758_,
		_w767_,
		_w1120_,
		_w1136_,
		_w4645_
	);
	LUT2 #(
		.INIT('h1)
	) name4183 (
		_w4644_,
		_w4645_,
		_w4646_
	);
	LUT2 #(
		.INIT('h8)
	) name4184 (
		_w760_,
		_w1143_,
		_w4647_
	);
	LUT3 #(
		.INIT('h0d)
	) name4185 (
		\P1_reg2_reg[14]/NET0131 ,
		_w2411_,
		_w4647_,
		_w4648_
	);
	LUT4 #(
		.INIT('h5700)
	) name4186 (
		_w534_,
		_w4644_,
		_w4645_,
		_w4648_,
		_w4649_
	);
	LUT3 #(
		.INIT('h10)
	) name4187 (
		_w4643_,
		_w4642_,
		_w4649_,
		_w4650_
	);
	LUT4 #(
		.INIT('h1311)
	) name4188 (
		_w526_,
		_w4639_,
		_w4641_,
		_w4650_,
		_w4651_
	);
	LUT3 #(
		.INIT('hce)
	) name4189 (
		\P1_state_reg[0]/NET0131 ,
		_w4638_,
		_w4651_,
		_w4652_
	);
	LUT2 #(
		.INIT('h2)
	) name4190 (
		\P1_reg2_reg[15]/NET0131 ,
		_w511_,
		_w4653_
	);
	LUT2 #(
		.INIT('h8)
	) name4191 (
		\P1_reg2_reg[15]/NET0131 ,
		_w524_,
		_w4654_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name4192 (
		\P1_reg2_reg[15]/NET0131 ,
		_w528_,
		_w530_,
		_w533_,
		_w4655_
	);
	LUT4 #(
		.INIT('h2a08)
	) name4193 (
		_w534_,
		_w537_,
		_w762_,
		_w4123_,
		_w4656_
	);
	LUT3 #(
		.INIT('ha8)
	) name4194 (
		_w1183_,
		_w4655_,
		_w4656_,
		_w4657_
	);
	LUT4 #(
		.INIT('he020)
	) name4195 (
		\P1_reg2_reg[15]/NET0131 ,
		_w534_,
		_w1286_,
		_w4126_,
		_w4658_
	);
	LUT4 #(
		.INIT('h20e0)
	) name4196 (
		\P1_reg2_reg[15]/NET0131 ,
		_w534_,
		_w1114_,
		_w4128_,
		_w4659_
	);
	LUT4 #(
		.INIT('h6a00)
	) name4197 (
		_w780_,
		_w1120_,
		_w1121_,
		_w1136_,
		_w4660_
	);
	LUT2 #(
		.INIT('h4)
	) name4198 (
		_w780_,
		_w1138_,
		_w4661_
	);
	LUT2 #(
		.INIT('h1)
	) name4199 (
		_w4660_,
		_w4661_,
		_w4662_
	);
	LUT2 #(
		.INIT('h8)
	) name4200 (
		_w770_,
		_w1143_,
		_w4663_
	);
	LUT3 #(
		.INIT('h0d)
	) name4201 (
		\P1_reg2_reg[15]/NET0131 ,
		_w2411_,
		_w4663_,
		_w4664_
	);
	LUT4 #(
		.INIT('h5700)
	) name4202 (
		_w534_,
		_w4660_,
		_w4661_,
		_w4664_,
		_w4665_
	);
	LUT3 #(
		.INIT('h10)
	) name4203 (
		_w4659_,
		_w4658_,
		_w4665_,
		_w4666_
	);
	LUT4 #(
		.INIT('h1311)
	) name4204 (
		_w526_,
		_w4654_,
		_w4657_,
		_w4666_,
		_w4667_
	);
	LUT3 #(
		.INIT('hce)
	) name4205 (
		\P1_state_reg[0]/NET0131 ,
		_w4653_,
		_w4667_,
		_w4668_
	);
	LUT4 #(
		.INIT('h70d0)
	) name4206 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg1_reg[10]/NET0131 ,
		_w1476_,
		_w4669_
	);
	LUT2 #(
		.INIT('h8)
	) name4207 (
		\P2_reg1_reg[10]/NET0131 ,
		_w1487_,
		_w4670_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name4208 (
		\P2_reg1_reg[10]/NET0131 ,
		_w1491_,
		_w1493_,
		_w1496_,
		_w4671_
	);
	LUT4 #(
		.INIT('h8a20)
	) name4209 (
		_w1497_,
		_w2492_,
		_w2493_,
		_w4142_,
		_w4672_
	);
	LUT2 #(
		.INIT('h4)
	) name4210 (
		_w1657_,
		_w2084_,
		_w4673_
	);
	LUT2 #(
		.INIT('h8)
	) name4211 (
		_w2039_,
		_w4673_,
		_w4674_
	);
	LUT3 #(
		.INIT('ha2)
	) name4212 (
		\P2_reg1_reg[10]/NET0131 ,
		_w2633_,
		_w2660_,
		_w4675_
	);
	LUT2 #(
		.INIT('h1)
	) name4213 (
		_w4674_,
		_w4675_,
		_w4676_
	);
	LUT4 #(
		.INIT('h5700)
	) name4214 (
		_w2188_,
		_w4671_,
		_w4672_,
		_w4676_,
		_w4677_
	);
	LUT4 #(
		.INIT('h111d)
	) name4215 (
		\P2_reg1_reg[10]/NET0131 ,
		_w1497_,
		_w4152_,
		_w4153_,
		_w4678_
	);
	LUT2 #(
		.INIT('h2)
	) name4216 (
		_w2081_,
		_w4678_,
		_w4679_
	);
	LUT4 #(
		.INIT('haa02)
	) name4217 (
		\P2_reg1_reg[10]/NET0131 ,
		_w1491_,
		_w1493_,
		_w1496_,
		_w4680_
	);
	LUT4 #(
		.INIT('h1dd1)
	) name4218 (
		\P2_reg1_reg[10]/NET0131 ,
		_w2039_,
		_w2467_,
		_w4142_,
		_w4681_
	);
	LUT2 #(
		.INIT('h2)
	) name4219 (
		_w2038_,
		_w4681_,
		_w4682_
	);
	LUT4 #(
		.INIT('h8a20)
	) name4220 (
		_w2039_,
		_w2492_,
		_w2493_,
		_w4142_,
		_w4683_
	);
	LUT3 #(
		.INIT('ha8)
	) name4221 (
		_w2193_,
		_w4680_,
		_w4683_,
		_w4684_
	);
	LUT4 #(
		.INIT('h0100)
	) name4222 (
		_w4682_,
		_w4684_,
		_w4679_,
		_w4677_,
		_w4685_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name4223 (
		\P1_state_reg[0]/NET0131 ,
		_w1489_,
		_w4670_,
		_w4685_,
		_w4686_
	);
	LUT2 #(
		.INIT('he)
	) name4224 (
		_w4669_,
		_w4686_,
		_w4687_
	);
	LUT4 #(
		.INIT('h70d0)
	) name4225 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg1_reg[12]/NET0131 ,
		_w1476_,
		_w4688_
	);
	LUT2 #(
		.INIT('h8)
	) name4226 (
		\P2_reg1_reg[12]/NET0131 ,
		_w1487_,
		_w4689_
	);
	LUT4 #(
		.INIT('h20e0)
	) name4227 (
		\P2_reg1_reg[12]/NET0131 ,
		_w1497_,
		_w2081_,
		_w4180_,
		_w4690_
	);
	LUT3 #(
		.INIT('h40)
	) name4228 (
		_w1746_,
		_w2039_,
		_w2084_,
		_w4691_
	);
	LUT3 #(
		.INIT('ha2)
	) name4229 (
		\P2_reg1_reg[12]/NET0131 ,
		_w2633_,
		_w2660_,
		_w4692_
	);
	LUT2 #(
		.INIT('h1)
	) name4230 (
		_w4691_,
		_w4692_,
		_w4693_
	);
	LUT2 #(
		.INIT('h4)
	) name4231 (
		_w4690_,
		_w4693_,
		_w4694_
	);
	LUT4 #(
		.INIT('haa02)
	) name4232 (
		\P2_reg1_reg[12]/NET0131 ,
		_w1491_,
		_w1493_,
		_w1496_,
		_w4695_
	);
	LUT4 #(
		.INIT('h20e0)
	) name4233 (
		\P2_reg1_reg[12]/NET0131 ,
		_w2039_,
		_w2193_,
		_w4182_,
		_w4696_
	);
	LUT4 #(
		.INIT('h20e0)
	) name4234 (
		\P2_reg1_reg[12]/NET0131 ,
		_w1497_,
		_w2188_,
		_w4182_,
		_w4697_
	);
	LUT4 #(
		.INIT('h40b0)
	) name4235 (
		_w1687_,
		_w1692_,
		_w2039_,
		_w4168_,
		_w4698_
	);
	LUT3 #(
		.INIT('ha8)
	) name4236 (
		_w2038_,
		_w4695_,
		_w4698_,
		_w4699_
	);
	LUT3 #(
		.INIT('h01)
	) name4237 (
		_w4697_,
		_w4699_,
		_w4696_,
		_w4700_
	);
	LUT4 #(
		.INIT('h3111)
	) name4238 (
		_w1489_,
		_w4689_,
		_w4694_,
		_w4700_,
		_w4701_
	);
	LUT3 #(
		.INIT('hce)
	) name4239 (
		\P1_state_reg[0]/NET0131 ,
		_w4688_,
		_w4701_,
		_w4702_
	);
	LUT4 #(
		.INIT('h70d0)
	) name4240 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg1_reg[13]/NET0131 ,
		_w1476_,
		_w4703_
	);
	LUT2 #(
		.INIT('h8)
	) name4241 (
		\P2_reg1_reg[13]/NET0131 ,
		_w1487_,
		_w4704_
	);
	LUT4 #(
		.INIT('haa02)
	) name4242 (
		\P2_reg1_reg[13]/NET0131 ,
		_w1491_,
		_w1493_,
		_w1496_,
		_w4705_
	);
	LUT4 #(
		.INIT('h8a20)
	) name4243 (
		_w2039_,
		_w2536_,
		_w2541_,
		_w4190_,
		_w4706_
	);
	LUT3 #(
		.INIT('ha8)
	) name4244 (
		_w2038_,
		_w4705_,
		_w4706_,
		_w4707_
	);
	LUT4 #(
		.INIT('h208a)
	) name4245 (
		_w2039_,
		_w2563_,
		_w2554_,
		_w4190_,
		_w4708_
	);
	LUT3 #(
		.INIT('ha8)
	) name4246 (
		_w2193_,
		_w4705_,
		_w4708_,
		_w4709_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name4247 (
		\P2_reg1_reg[13]/NET0131 ,
		_w1491_,
		_w1493_,
		_w1496_,
		_w4710_
	);
	LUT4 #(
		.INIT('h208a)
	) name4248 (
		_w1497_,
		_w2563_,
		_w2554_,
		_w4190_,
		_w4711_
	);
	LUT3 #(
		.INIT('ha8)
	) name4249 (
		_w2188_,
		_w4710_,
		_w4711_,
		_w4712_
	);
	LUT4 #(
		.INIT('h20e0)
	) name4250 (
		\P2_reg1_reg[13]/NET0131 ,
		_w1497_,
		_w2081_,
		_w4199_,
		_w4713_
	);
	LUT3 #(
		.INIT('h40)
	) name4251 (
		_w1761_,
		_w2039_,
		_w2084_,
		_w4714_
	);
	LUT3 #(
		.INIT('ha2)
	) name4252 (
		\P2_reg1_reg[13]/NET0131 ,
		_w2633_,
		_w2660_,
		_w4715_
	);
	LUT2 #(
		.INIT('h1)
	) name4253 (
		_w4714_,
		_w4715_,
		_w4716_
	);
	LUT2 #(
		.INIT('h4)
	) name4254 (
		_w4713_,
		_w4716_,
		_w4717_
	);
	LUT4 #(
		.INIT('h0100)
	) name4255 (
		_w4712_,
		_w4709_,
		_w4707_,
		_w4717_,
		_w4718_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name4256 (
		\P1_state_reg[0]/NET0131 ,
		_w1489_,
		_w4704_,
		_w4718_,
		_w4719_
	);
	LUT2 #(
		.INIT('he)
	) name4257 (
		_w4703_,
		_w4719_,
		_w4720_
	);
	LUT4 #(
		.INIT('h70d0)
	) name4258 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg1_reg[16]/NET0131 ,
		_w1476_,
		_w4721_
	);
	LUT2 #(
		.INIT('h8)
	) name4259 (
		\P2_reg1_reg[16]/NET0131 ,
		_w1487_,
		_w4722_
	);
	LUT4 #(
		.INIT('h1dd1)
	) name4260 (
		\P2_reg1_reg[16]/NET0131 ,
		_w2039_,
		_w4593_,
		_w4594_,
		_w4723_
	);
	LUT2 #(
		.INIT('h2)
	) name4261 (
		_w2038_,
		_w4723_,
		_w4724_
	);
	LUT4 #(
		.INIT('hd11d)
	) name4262 (
		\P2_reg1_reg[16]/NET0131 ,
		_w2039_,
		_w4593_,
		_w4599_,
		_w4725_
	);
	LUT2 #(
		.INIT('h2)
	) name4263 (
		_w2193_,
		_w4725_,
		_w4726_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name4264 (
		\P2_reg1_reg[16]/NET0131 ,
		_w1491_,
		_w1493_,
		_w1496_,
		_w4727_
	);
	LUT4 #(
		.INIT('hd11d)
	) name4265 (
		\P2_reg1_reg[16]/NET0131 ,
		_w1497_,
		_w4593_,
		_w4599_,
		_w4728_
	);
	LUT4 #(
		.INIT('haa20)
	) name4266 (
		_w1497_,
		_w1781_,
		_w4524_,
		_w4602_,
		_w4729_
	);
	LUT4 #(
		.INIT('hf100)
	) name4267 (
		_w1509_,
		_w1790_,
		_w1794_,
		_w2963_,
		_w4730_
	);
	LUT3 #(
		.INIT('ha2)
	) name4268 (
		\P2_reg1_reg[16]/NET0131 ,
		_w2633_,
		_w2660_,
		_w4731_
	);
	LUT2 #(
		.INIT('h1)
	) name4269 (
		_w4730_,
		_w4731_,
		_w4732_
	);
	LUT4 #(
		.INIT('h5700)
	) name4270 (
		_w2081_,
		_w4727_,
		_w4729_,
		_w4732_,
		_w4733_
	);
	LUT3 #(
		.INIT('hd0)
	) name4271 (
		_w2188_,
		_w4728_,
		_w4733_,
		_w4734_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name4272 (
		_w1489_,
		_w4726_,
		_w4724_,
		_w4734_,
		_w4735_
	);
	LUT4 #(
		.INIT('heeec)
	) name4273 (
		\P1_state_reg[0]/NET0131 ,
		_w4721_,
		_w4722_,
		_w4735_,
		_w4736_
	);
	LUT2 #(
		.INIT('h2)
	) name4274 (
		\P1_reg2_reg[9]/NET0131 ,
		_w511_,
		_w4737_
	);
	LUT2 #(
		.INIT('h8)
	) name4275 (
		\P1_reg2_reg[9]/NET0131 ,
		_w524_,
		_w4738_
	);
	LUT2 #(
		.INIT('h8)
	) name4276 (
		_w831_,
		_w1143_,
		_w4739_
	);
	LUT4 #(
		.INIT('h00a2)
	) name4277 (
		\P1_reg2_reg[9]/NET0131 ,
		_w534_,
		_w1141_,
		_w1143_,
		_w4740_
	);
	LUT2 #(
		.INIT('h1)
	) name4278 (
		_w4739_,
		_w4740_,
		_w4741_
	);
	LUT4 #(
		.INIT('h7500)
	) name4279 (
		_w534_,
		_w4254_,
		_w4257_,
		_w4741_,
		_w4742_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name4280 (
		\P1_state_reg[0]/NET0131 ,
		_w526_,
		_w4738_,
		_w4742_,
		_w4743_
	);
	LUT2 #(
		.INIT('he)
	) name4281 (
		_w4737_,
		_w4743_,
		_w4744_
	);
	LUT4 #(
		.INIT('h70d0)
	) name4282 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg1_reg[9]/NET0131 ,
		_w1476_,
		_w4745_
	);
	LUT2 #(
		.INIT('h8)
	) name4283 (
		\P2_reg1_reg[9]/NET0131 ,
		_w1487_,
		_w4746_
	);
	LUT4 #(
		.INIT('h20e0)
	) name4284 (
		\P2_reg1_reg[9]/NET0131 ,
		_w1497_,
		_w2188_,
		_w4231_,
		_w4747_
	);
	LUT4 #(
		.INIT('h20e0)
	) name4285 (
		\P2_reg1_reg[9]/NET0131 ,
		_w2039_,
		_w2193_,
		_w4231_,
		_w4748_
	);
	LUT4 #(
		.INIT('hf100)
	) name4286 (
		_w1509_,
		_w1668_,
		_w1671_,
		_w2084_,
		_w4749_
	);
	LUT2 #(
		.INIT('h8)
	) name4287 (
		_w2039_,
		_w4749_,
		_w4750_
	);
	LUT3 #(
		.INIT('ha2)
	) name4288 (
		\P2_reg1_reg[9]/NET0131 ,
		_w2633_,
		_w2660_,
		_w4751_
	);
	LUT2 #(
		.INIT('h1)
	) name4289 (
		_w4750_,
		_w4751_,
		_w4752_
	);
	LUT3 #(
		.INIT('h10)
	) name4290 (
		_w4748_,
		_w4747_,
		_w4752_,
		_w4753_
	);
	LUT4 #(
		.INIT('hc808)
	) name4291 (
		\P2_reg1_reg[9]/NET0131 ,
		_w2038_,
		_w2039_,
		_w4229_,
		_w4754_
	);
	LUT4 #(
		.INIT('h20e0)
	) name4292 (
		\P2_reg1_reg[9]/NET0131 ,
		_w1497_,
		_w2081_,
		_w4238_,
		_w4755_
	);
	LUT2 #(
		.INIT('h1)
	) name4293 (
		_w4754_,
		_w4755_,
		_w4756_
	);
	LUT4 #(
		.INIT('h3111)
	) name4294 (
		_w1489_,
		_w4746_,
		_w4753_,
		_w4756_,
		_w4757_
	);
	LUT3 #(
		.INIT('hce)
	) name4295 (
		\P1_state_reg[0]/NET0131 ,
		_w4745_,
		_w4757_,
		_w4758_
	);
	LUT4 #(
		.INIT('h70d0)
	) name4296 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg2_reg[10]/NET0131 ,
		_w1476_,
		_w4759_
	);
	LUT2 #(
		.INIT('h8)
	) name4297 (
		\P2_reg2_reg[10]/NET0131 ,
		_w1487_,
		_w4760_
	);
	LUT4 #(
		.INIT('haa02)
	) name4298 (
		\P2_reg2_reg[10]/NET0131 ,
		_w1491_,
		_w1493_,
		_w1496_,
		_w4761_
	);
	LUT3 #(
		.INIT('ha8)
	) name4299 (
		\P2_reg2_reg[10]/NET0131 ,
		_w2086_,
		_w2087_,
		_w4762_
	);
	LUT2 #(
		.INIT('h4)
	) name4300 (
		_w1643_,
		_w2088_,
		_w4763_
	);
	LUT3 #(
		.INIT('h07)
	) name4301 (
		_w1497_,
		_w4673_,
		_w4763_,
		_w4764_
	);
	LUT2 #(
		.INIT('h4)
	) name4302 (
		_w4762_,
		_w4764_,
		_w4765_
	);
	LUT4 #(
		.INIT('h5700)
	) name4303 (
		_w2188_,
		_w4683_,
		_w4761_,
		_w4765_,
		_w4766_
	);
	LUT4 #(
		.INIT('h111d)
	) name4304 (
		\P2_reg2_reg[10]/NET0131 ,
		_w2039_,
		_w4152_,
		_w4153_,
		_w4767_
	);
	LUT2 #(
		.INIT('h2)
	) name4305 (
		_w2081_,
		_w4767_,
		_w4768_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name4306 (
		\P2_reg2_reg[10]/NET0131 ,
		_w1491_,
		_w1493_,
		_w1496_,
		_w4769_
	);
	LUT3 #(
		.INIT('ha8)
	) name4307 (
		_w2193_,
		_w4672_,
		_w4769_,
		_w4770_
	);
	LUT4 #(
		.INIT('h1dd1)
	) name4308 (
		\P2_reg2_reg[10]/NET0131 ,
		_w1497_,
		_w2467_,
		_w4142_,
		_w4771_
	);
	LUT2 #(
		.INIT('h2)
	) name4309 (
		_w2038_,
		_w4771_,
		_w4772_
	);
	LUT4 #(
		.INIT('h0100)
	) name4310 (
		_w4770_,
		_w4772_,
		_w4768_,
		_w4766_,
		_w4773_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name4311 (
		\P1_state_reg[0]/NET0131 ,
		_w1489_,
		_w4760_,
		_w4773_,
		_w4774_
	);
	LUT2 #(
		.INIT('he)
	) name4312 (
		_w4759_,
		_w4774_,
		_w4775_
	);
	LUT4 #(
		.INIT('h70d0)
	) name4313 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg2_reg[12]/NET0131 ,
		_w1476_,
		_w4776_
	);
	LUT2 #(
		.INIT('h8)
	) name4314 (
		\P2_reg2_reg[12]/NET0131 ,
		_w1487_,
		_w4777_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name4315 (
		\P2_reg2_reg[12]/NET0131 ,
		_w1491_,
		_w1493_,
		_w1496_,
		_w4778_
	);
	LUT4 #(
		.INIT('h20e0)
	) name4316 (
		\P2_reg2_reg[12]/NET0131 ,
		_w1497_,
		_w2193_,
		_w4182_,
		_w4779_
	);
	LUT3 #(
		.INIT('ha8)
	) name4317 (
		\P2_reg2_reg[12]/NET0131 ,
		_w2086_,
		_w2087_,
		_w4780_
	);
	LUT2 #(
		.INIT('h4)
	) name4318 (
		_w1732_,
		_w2088_,
		_w4781_
	);
	LUT4 #(
		.INIT('h00df)
	) name4319 (
		_w1497_,
		_w1746_,
		_w2084_,
		_w4781_,
		_w4782_
	);
	LUT2 #(
		.INIT('h4)
	) name4320 (
		_w4780_,
		_w4782_,
		_w4783_
	);
	LUT2 #(
		.INIT('h4)
	) name4321 (
		_w4779_,
		_w4783_,
		_w4784_
	);
	LUT4 #(
		.INIT('h20e0)
	) name4322 (
		\P2_reg2_reg[12]/NET0131 ,
		_w2039_,
		_w2081_,
		_w4180_,
		_w4785_
	);
	LUT4 #(
		.INIT('h208a)
	) name4323 (
		_w1497_,
		_w1687_,
		_w1692_,
		_w4168_,
		_w4786_
	);
	LUT3 #(
		.INIT('ha8)
	) name4324 (
		_w2038_,
		_w4778_,
		_w4786_,
		_w4787_
	);
	LUT4 #(
		.INIT('h20e0)
	) name4325 (
		\P2_reg2_reg[12]/NET0131 ,
		_w2039_,
		_w2188_,
		_w4182_,
		_w4788_
	);
	LUT3 #(
		.INIT('h01)
	) name4326 (
		_w4787_,
		_w4788_,
		_w4785_,
		_w4789_
	);
	LUT4 #(
		.INIT('h3111)
	) name4327 (
		_w1489_,
		_w4777_,
		_w4784_,
		_w4789_,
		_w4790_
	);
	LUT3 #(
		.INIT('hce)
	) name4328 (
		\P1_state_reg[0]/NET0131 ,
		_w4776_,
		_w4790_,
		_w4791_
	);
	LUT4 #(
		.INIT('h70d0)
	) name4329 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg2_reg[13]/NET0131 ,
		_w1476_,
		_w4792_
	);
	LUT2 #(
		.INIT('h8)
	) name4330 (
		\P2_reg2_reg[13]/NET0131 ,
		_w1487_,
		_w4793_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name4331 (
		\P2_reg2_reg[13]/NET0131 ,
		_w1491_,
		_w1493_,
		_w1496_,
		_w4794_
	);
	LUT4 #(
		.INIT('h8a20)
	) name4332 (
		_w1497_,
		_w2536_,
		_w2541_,
		_w4190_,
		_w4795_
	);
	LUT3 #(
		.INIT('ha8)
	) name4333 (
		_w2038_,
		_w4794_,
		_w4795_,
		_w4796_
	);
	LUT3 #(
		.INIT('ha8)
	) name4334 (
		_w2193_,
		_w4711_,
		_w4794_,
		_w4797_
	);
	LUT4 #(
		.INIT('haa02)
	) name4335 (
		\P2_reg2_reg[13]/NET0131 ,
		_w1491_,
		_w1493_,
		_w1496_,
		_w4798_
	);
	LUT3 #(
		.INIT('ha8)
	) name4336 (
		_w2188_,
		_w4708_,
		_w4798_,
		_w4799_
	);
	LUT4 #(
		.INIT('h20e0)
	) name4337 (
		\P2_reg2_reg[13]/NET0131 ,
		_w2039_,
		_w2081_,
		_w4199_,
		_w4800_
	);
	LUT3 #(
		.INIT('ha8)
	) name4338 (
		\P2_reg2_reg[13]/NET0131 ,
		_w2086_,
		_w2087_,
		_w4801_
	);
	LUT2 #(
		.INIT('h4)
	) name4339 (
		_w1749_,
		_w2088_,
		_w4802_
	);
	LUT4 #(
		.INIT('h00df)
	) name4340 (
		_w1497_,
		_w1761_,
		_w2084_,
		_w4802_,
		_w4803_
	);
	LUT2 #(
		.INIT('h4)
	) name4341 (
		_w4801_,
		_w4803_,
		_w4804_
	);
	LUT2 #(
		.INIT('h4)
	) name4342 (
		_w4800_,
		_w4804_,
		_w4805_
	);
	LUT4 #(
		.INIT('h0100)
	) name4343 (
		_w4799_,
		_w4797_,
		_w4796_,
		_w4805_,
		_w4806_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name4344 (
		\P1_state_reg[0]/NET0131 ,
		_w1489_,
		_w4793_,
		_w4806_,
		_w4807_
	);
	LUT2 #(
		.INIT('he)
	) name4345 (
		_w4792_,
		_w4807_,
		_w4808_
	);
	LUT4 #(
		.INIT('h70d0)
	) name4346 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg2_reg[16]/NET0131 ,
		_w1476_,
		_w4809_
	);
	LUT2 #(
		.INIT('h8)
	) name4347 (
		\P2_reg2_reg[16]/NET0131 ,
		_w1487_,
		_w4810_
	);
	LUT4 #(
		.INIT('h1dd1)
	) name4348 (
		\P2_reg2_reg[16]/NET0131 ,
		_w1497_,
		_w4593_,
		_w4594_,
		_w4811_
	);
	LUT2 #(
		.INIT('h2)
	) name4349 (
		_w2038_,
		_w4811_,
		_w4812_
	);
	LUT4 #(
		.INIT('hd11d)
	) name4350 (
		\P2_reg2_reg[16]/NET0131 ,
		_w1497_,
		_w4593_,
		_w4599_,
		_w4813_
	);
	LUT2 #(
		.INIT('h2)
	) name4351 (
		_w2193_,
		_w4813_,
		_w4814_
	);
	LUT4 #(
		.INIT('haa02)
	) name4352 (
		\P2_reg2_reg[16]/NET0131 ,
		_w1491_,
		_w1493_,
		_w1496_,
		_w4815_
	);
	LUT4 #(
		.INIT('hd11d)
	) name4353 (
		\P2_reg2_reg[16]/NET0131 ,
		_w2039_,
		_w4593_,
		_w4599_,
		_w4816_
	);
	LUT4 #(
		.INIT('hcc40)
	) name4354 (
		_w1781_,
		_w2039_,
		_w4524_,
		_w4602_,
		_w4817_
	);
	LUT3 #(
		.INIT('ha8)
	) name4355 (
		\P2_reg2_reg[16]/NET0131 ,
		_w2086_,
		_w2087_,
		_w4818_
	);
	LUT4 #(
		.INIT('hf100)
	) name4356 (
		_w1509_,
		_w1790_,
		_w1794_,
		_w2085_,
		_w4819_
	);
	LUT2 #(
		.INIT('h4)
	) name4357 (
		_w471_,
		_w2088_,
		_w4820_
	);
	LUT3 #(
		.INIT('h01)
	) name4358 (
		_w4819_,
		_w4820_,
		_w4818_,
		_w4821_
	);
	LUT4 #(
		.INIT('h5700)
	) name4359 (
		_w2081_,
		_w4815_,
		_w4817_,
		_w4821_,
		_w4822_
	);
	LUT3 #(
		.INIT('hd0)
	) name4360 (
		_w2188_,
		_w4816_,
		_w4822_,
		_w4823_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name4361 (
		_w1489_,
		_w4814_,
		_w4812_,
		_w4823_,
		_w4824_
	);
	LUT4 #(
		.INIT('heeec)
	) name4362 (
		\P1_state_reg[0]/NET0131 ,
		_w4809_,
		_w4810_,
		_w4824_,
		_w4825_
	);
	LUT2 #(
		.INIT('h2)
	) name4363 (
		\P1_reg0_reg[15]/NET0131 ,
		_w511_,
		_w4826_
	);
	LUT2 #(
		.INIT('h8)
	) name4364 (
		\P1_reg0_reg[15]/NET0131 ,
		_w524_,
		_w4827_
	);
	LUT4 #(
		.INIT('haaa2)
	) name4365 (
		\P1_reg0_reg[15]/NET0131 ,
		_w2692_,
		_w3005_,
		_w3664_,
		_w4828_
	);
	LUT4 #(
		.INIT('h7020)
	) name4366 (
		_w537_,
		_w762_,
		_w1183_,
		_w4123_,
		_w4829_
	);
	LUT2 #(
		.INIT('h8)
	) name4367 (
		_w1286_,
		_w4126_,
		_w4830_
	);
	LUT3 #(
		.INIT('hd0)
	) name4368 (
		_w1114_,
		_w4128_,
		_w4662_,
		_w4831_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name4369 (
		_w2688_,
		_w4829_,
		_w4830_,
		_w4831_,
		_w4832_
	);
	LUT4 #(
		.INIT('h1113)
	) name4370 (
		_w526_,
		_w4827_,
		_w4828_,
		_w4832_,
		_w4833_
	);
	LUT3 #(
		.INIT('hce)
	) name4371 (
		\P1_state_reg[0]/NET0131 ,
		_w4826_,
		_w4833_,
		_w4834_
	);
	LUT2 #(
		.INIT('h2)
	) name4372 (
		\P1_reg0_reg[4]/NET0131 ,
		_w511_,
		_w4835_
	);
	LUT2 #(
		.INIT('h8)
	) name4373 (
		\P1_reg0_reg[4]/NET0131 ,
		_w524_,
		_w4836_
	);
	LUT4 #(
		.INIT('haaa8)
	) name4374 (
		\P1_reg0_reg[4]/NET0131 ,
		_w528_,
		_w530_,
		_w533_,
		_w4837_
	);
	LUT4 #(
		.INIT('h7020)
	) name4375 (
		_w537_,
		_w876_,
		_w2688_,
		_w4537_,
		_w4838_
	);
	LUT3 #(
		.INIT('ha8)
	) name4376 (
		_w1183_,
		_w4837_,
		_w4838_,
		_w4839_
	);
	LUT4 #(
		.INIT('h08c8)
	) name4377 (
		\P1_reg0_reg[4]/NET0131 ,
		_w1114_,
		_w2688_,
		_w4539_,
		_w4840_
	);
	LUT4 #(
		.INIT('hc808)
	) name4378 (
		\P1_reg0_reg[4]/NET0131 ,
		_w1286_,
		_w2688_,
		_w4541_,
		_w4841_
	);
	LUT4 #(
		.INIT('hc355)
	) name4379 (
		\P1_reg0_reg[4]/NET0131 ,
		_w894_,
		_w1115_,
		_w2688_,
		_w4842_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name4380 (
		\P1_reg0_reg[4]/NET0131 ,
		_w1138_,
		_w2425_,
		_w2688_,
		_w4843_
	);
	LUT4 #(
		.INIT('h0001)
	) name4381 (
		_w894_,
		_w1104_,
		_w1106_,
		_w1111_,
		_w4844_
	);
	LUT2 #(
		.INIT('h8)
	) name4382 (
		_w2688_,
		_w4844_,
		_w4845_
	);
	LUT4 #(
		.INIT('h0031)
	) name4383 (
		_w1136_,
		_w4843_,
		_w4842_,
		_w4845_,
		_w4846_
	);
	LUT3 #(
		.INIT('h10)
	) name4384 (
		_w4841_,
		_w4840_,
		_w4846_,
		_w4847_
	);
	LUT4 #(
		.INIT('h1311)
	) name4385 (
		_w526_,
		_w4836_,
		_w4839_,
		_w4847_,
		_w4848_
	);
	LUT3 #(
		.INIT('hce)
	) name4386 (
		\P1_state_reg[0]/NET0131 ,
		_w4835_,
		_w4848_,
		_w4849_
	);
	LUT2 #(
		.INIT('h8)
	) name4387 (
		\P1_reg1_reg[15]/NET0131 ,
		_w524_,
		_w4850_
	);
	LUT3 #(
		.INIT('h2a)
	) name4388 (
		\P1_reg1_reg[15]/NET0131 ,
		_w2426_,
		_w3686_,
		_w4851_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name4389 (
		_w2421_,
		_w4829_,
		_w4830_,
		_w4831_,
		_w4852_
	);
	LUT4 #(
		.INIT('h1113)
	) name4390 (
		_w526_,
		_w4850_,
		_w4851_,
		_w4852_,
		_w4853_
	);
	LUT2 #(
		.INIT('h2)
	) name4391 (
		\P1_reg1_reg[15]/NET0131 ,
		_w511_,
		_w4854_
	);
	LUT3 #(
		.INIT('hf2)
	) name4392 (
		\P1_state_reg[0]/NET0131 ,
		_w4853_,
		_w4854_,
		_w4855_
	);
	LUT4 #(
		.INIT('h70d0)
	) name4393 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg0_reg[10]/NET0131 ,
		_w1476_,
		_w4856_
	);
	LUT2 #(
		.INIT('h8)
	) name4394 (
		\P2_reg0_reg[10]/NET0131 ,
		_w1487_,
		_w4857_
	);
	LUT4 #(
		.INIT('haaa8)
	) name4395 (
		\P2_reg0_reg[10]/NET0131 ,
		_w1491_,
		_w1493_,
		_w1496_,
		_w4858_
	);
	LUT4 #(
		.INIT('h1dd1)
	) name4396 (
		\P2_reg0_reg[10]/NET0131 ,
		_w2277_,
		_w2467_,
		_w4142_,
		_w4859_
	);
	LUT2 #(
		.INIT('h8)
	) name4397 (
		_w2277_,
		_w4673_,
		_w4860_
	);
	LUT3 #(
		.INIT('ha2)
	) name4398 (
		\P2_reg0_reg[10]/NET0131 ,
		_w2633_,
		_w2634_,
		_w4861_
	);
	LUT2 #(
		.INIT('h1)
	) name4399 (
		_w4860_,
		_w4861_,
		_w4862_
	);
	LUT3 #(
		.INIT('he0)
	) name4400 (
		_w2276_,
		_w4859_,
		_w4862_,
		_w4863_
	);
	LUT4 #(
		.INIT('h111d)
	) name4401 (
		\P2_reg0_reg[10]/NET0131 ,
		_w2272_,
		_w4152_,
		_w4153_,
		_w4864_
	);
	LUT2 #(
		.INIT('h2)
	) name4402 (
		_w2081_,
		_w4864_,
		_w4865_
	);
	LUT4 #(
		.INIT('h8a20)
	) name4403 (
		_w2277_,
		_w2492_,
		_w2493_,
		_w4142_,
		_w4866_
	);
	LUT3 #(
		.INIT('h54)
	) name4404 (
		_w2192_,
		_w4858_,
		_w4866_,
		_w4867_
	);
	LUT4 #(
		.INIT('h1dd1)
	) name4405 (
		\P2_reg0_reg[10]/NET0131 ,
		_w2272_,
		_w2467_,
		_w4142_,
		_w4868_
	);
	LUT2 #(
		.INIT('h2)
	) name4406 (
		_w2290_,
		_w4868_,
		_w4869_
	);
	LUT4 #(
		.INIT('h0100)
	) name4407 (
		_w4867_,
		_w4869_,
		_w4865_,
		_w4863_,
		_w4870_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name4408 (
		\P1_state_reg[0]/NET0131 ,
		_w1489_,
		_w4857_,
		_w4870_,
		_w4871_
	);
	LUT2 #(
		.INIT('he)
	) name4409 (
		_w4856_,
		_w4871_,
		_w4872_
	);
	LUT4 #(
		.INIT('h70d0)
	) name4410 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg0_reg[12]/NET0131 ,
		_w1476_,
		_w4873_
	);
	LUT2 #(
		.INIT('h8)
	) name4411 (
		\P2_reg0_reg[12]/NET0131 ,
		_w1487_,
		_w4874_
	);
	LUT4 #(
		.INIT('h02aa)
	) name4412 (
		\P2_reg0_reg[12]/NET0131 ,
		_w1491_,
		_w1493_,
		_w1496_,
		_w4875_
	);
	LUT4 #(
		.INIT('h08c8)
	) name4413 (
		\P2_reg0_reg[12]/NET0131 ,
		_w2081_,
		_w2272_,
		_w4180_,
		_w4876_
	);
	LUT3 #(
		.INIT('h40)
	) name4414 (
		_w1746_,
		_w2084_,
		_w2277_,
		_w4877_
	);
	LUT3 #(
		.INIT('ha2)
	) name4415 (
		\P2_reg0_reg[12]/NET0131 ,
		_w2633_,
		_w2634_,
		_w4878_
	);
	LUT2 #(
		.INIT('h1)
	) name4416 (
		_w4877_,
		_w4878_,
		_w4879_
	);
	LUT2 #(
		.INIT('h4)
	) name4417 (
		_w4876_,
		_w4879_,
		_w4880_
	);
	LUT4 #(
		.INIT('haaa8)
	) name4418 (
		\P2_reg0_reg[12]/NET0131 ,
		_w1491_,
		_w1493_,
		_w1496_,
		_w4881_
	);
	LUT4 #(
		.INIT('h0232)
	) name4419 (
		\P2_reg0_reg[12]/NET0131 ,
		_w2192_,
		_w2277_,
		_w4182_,
		_w4882_
	);
	LUT3 #(
		.INIT('ha8)
	) name4420 (
		_w2290_,
		_w4175_,
		_w4875_,
		_w4883_
	);
	LUT3 #(
		.INIT('h54)
	) name4421 (
		_w2276_,
		_w4169_,
		_w4881_,
		_w4884_
	);
	LUT3 #(
		.INIT('h01)
	) name4422 (
		_w4883_,
		_w4884_,
		_w4882_,
		_w4885_
	);
	LUT4 #(
		.INIT('h3111)
	) name4423 (
		_w1489_,
		_w4874_,
		_w4880_,
		_w4885_,
		_w4886_
	);
	LUT3 #(
		.INIT('hce)
	) name4424 (
		\P1_state_reg[0]/NET0131 ,
		_w4873_,
		_w4886_,
		_w4887_
	);
	LUT4 #(
		.INIT('h70d0)
	) name4425 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg0_reg[13]/NET0131 ,
		_w1476_,
		_w4888_
	);
	LUT2 #(
		.INIT('h8)
	) name4426 (
		\P2_reg0_reg[13]/NET0131 ,
		_w1487_,
		_w4889_
	);
	LUT4 #(
		.INIT('h02aa)
	) name4427 (
		\P2_reg0_reg[13]/NET0131 ,
		_w1491_,
		_w1493_,
		_w1496_,
		_w4890_
	);
	LUT3 #(
		.INIT('ha8)
	) name4428 (
		_w2290_,
		_w4194_,
		_w4890_,
		_w4891_
	);
	LUT4 #(
		.INIT('haaa8)
	) name4429 (
		\P2_reg0_reg[13]/NET0131 ,
		_w1491_,
		_w1493_,
		_w1496_,
		_w4892_
	);
	LUT3 #(
		.INIT('h54)
	) name4430 (
		_w2276_,
		_w4191_,
		_w4892_,
		_w4893_
	);
	LUT4 #(
		.INIT('h208a)
	) name4431 (
		_w2277_,
		_w2563_,
		_w2554_,
		_w4190_,
		_w4894_
	);
	LUT3 #(
		.INIT('h54)
	) name4432 (
		_w2192_,
		_w4892_,
		_w4894_,
		_w4895_
	);
	LUT4 #(
		.INIT('h08c8)
	) name4433 (
		\P2_reg0_reg[13]/NET0131 ,
		_w2081_,
		_w2272_,
		_w4199_,
		_w4896_
	);
	LUT3 #(
		.INIT('h40)
	) name4434 (
		_w1761_,
		_w2084_,
		_w2277_,
		_w4897_
	);
	LUT3 #(
		.INIT('ha2)
	) name4435 (
		\P2_reg0_reg[13]/NET0131 ,
		_w2633_,
		_w2634_,
		_w4898_
	);
	LUT2 #(
		.INIT('h1)
	) name4436 (
		_w4897_,
		_w4898_,
		_w4899_
	);
	LUT2 #(
		.INIT('h4)
	) name4437 (
		_w4896_,
		_w4899_,
		_w4900_
	);
	LUT4 #(
		.INIT('h0100)
	) name4438 (
		_w4893_,
		_w4891_,
		_w4895_,
		_w4900_,
		_w4901_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name4439 (
		\P1_state_reg[0]/NET0131 ,
		_w1489_,
		_w4889_,
		_w4901_,
		_w4902_
	);
	LUT2 #(
		.INIT('he)
	) name4440 (
		_w4888_,
		_w4902_,
		_w4903_
	);
	LUT2 #(
		.INIT('h2)
	) name4441 (
		\P1_reg1_reg[4]/NET0131 ,
		_w511_,
		_w4904_
	);
	LUT2 #(
		.INIT('h8)
	) name4442 (
		\P1_reg1_reg[4]/NET0131 ,
		_w524_,
		_w4905_
	);
	LUT4 #(
		.INIT('haa02)
	) name4443 (
		\P1_reg1_reg[4]/NET0131 ,
		_w528_,
		_w530_,
		_w533_,
		_w4906_
	);
	LUT4 #(
		.INIT('h7020)
	) name4444 (
		_w537_,
		_w876_,
		_w2421_,
		_w4537_,
		_w4907_
	);
	LUT3 #(
		.INIT('ha8)
	) name4445 (
		_w1183_,
		_w4906_,
		_w4907_,
		_w4908_
	);
	LUT4 #(
		.INIT('h08c8)
	) name4446 (
		\P1_reg1_reg[4]/NET0131 ,
		_w1114_,
		_w2421_,
		_w4539_,
		_w4909_
	);
	LUT4 #(
		.INIT('hc808)
	) name4447 (
		\P1_reg1_reg[4]/NET0131 ,
		_w1286_,
		_w2421_,
		_w4541_,
		_w4910_
	);
	LUT4 #(
		.INIT('hc355)
	) name4448 (
		\P1_reg1_reg[4]/NET0131 ,
		_w894_,
		_w1115_,
		_w2421_,
		_w4911_
	);
	LUT4 #(
		.INIT('h08aa)
	) name4449 (
		\P1_reg1_reg[4]/NET0131 ,
		_w1138_,
		_w2421_,
		_w2425_,
		_w4912_
	);
	LUT2 #(
		.INIT('h8)
	) name4450 (
		_w2421_,
		_w4844_,
		_w4913_
	);
	LUT4 #(
		.INIT('h0031)
	) name4451 (
		_w1136_,
		_w4912_,
		_w4911_,
		_w4913_,
		_w4914_
	);
	LUT3 #(
		.INIT('h10)
	) name4452 (
		_w4910_,
		_w4909_,
		_w4914_,
		_w4915_
	);
	LUT4 #(
		.INIT('h1311)
	) name4453 (
		_w526_,
		_w4905_,
		_w4908_,
		_w4915_,
		_w4916_
	);
	LUT3 #(
		.INIT('hce)
	) name4454 (
		\P1_state_reg[0]/NET0131 ,
		_w4904_,
		_w4916_,
		_w4917_
	);
	LUT2 #(
		.INIT('h4)
	) name4455 (
		\P1_reg3_reg[3]/NET0131 ,
		_w524_,
		_w4918_
	);
	LUT4 #(
		.INIT('h4150)
	) name4456 (
		_w537_,
		_w876_,
		_w887_,
		_w1153_,
		_w4919_
	);
	LUT3 #(
		.INIT('h80)
	) name4457 (
		_w537_,
		_w847_,
		_w848_,
		_w4920_
	);
	LUT3 #(
		.INIT('h02)
	) name4458 (
		_w1183_,
		_w4919_,
		_w4920_,
		_w4921_
	);
	LUT4 #(
		.INIT('h10e0)
	) name4459 (
		_w872_,
		_w873_,
		_w1114_,
		_w1434_,
		_w4922_
	);
	LUT4 #(
		.INIT('h7f80)
	) name4460 (
		_w853_,
		_w861_,
		_w869_,
		_w881_,
		_w4923_
	);
	LUT2 #(
		.INIT('h8)
	) name4461 (
		_w1136_,
		_w4923_,
		_w4924_
	);
	LUT4 #(
		.INIT('he010)
	) name4462 (
		_w1210_,
		_w1213_,
		_w1286_,
		_w1434_,
		_w4925_
	);
	LUT3 #(
		.INIT('h01)
	) name4463 (
		_w4924_,
		_w4922_,
		_w4925_,
		_w4926_
	);
	LUT3 #(
		.INIT('h04)
	) name4464 (
		_w881_,
		_w2259_,
		_w2260_,
		_w4927_
	);
	LUT4 #(
		.INIT('h00ae)
	) name4465 (
		\P1_reg3_reg[3]/NET0131 ,
		_w3143_,
		_w3237_,
		_w4927_,
		_w4928_
	);
	LUT4 #(
		.INIT('h7500)
	) name4466 (
		_w2197_,
		_w4921_,
		_w4926_,
		_w4928_,
		_w4929_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name4467 (
		\P1_state_reg[0]/NET0131 ,
		_w526_,
		_w4918_,
		_w4929_,
		_w4930_
	);
	LUT2 #(
		.INIT('h2)
	) name4468 (
		\P1_reg3_reg[3]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w4931_
	);
	LUT3 #(
		.INIT('h9d)
	) name4469 (
		\P1_reg3_reg[3]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w510_,
		_w4932_
	);
	LUT2 #(
		.INIT('hb)
	) name4470 (
		_w4930_,
		_w4932_,
		_w4933_
	);
	LUT2 #(
		.INIT('h8)
	) name4471 (
		_w524_,
		_w910_,
		_w4934_
	);
	LUT4 #(
		.INIT('h5655)
	) name4472 (
		_w903_,
		_w912_,
		_w924_,
		_w1154_,
		_w4935_
	);
	LUT4 #(
		.INIT('h80d0)
	) name4473 (
		_w537_,
		_w924_,
		_w2197_,
		_w4935_,
		_w4936_
	);
	LUT4 #(
		.INIT('h001f)
	) name4474 (
		_w528_,
		_w530_,
		_w533_,
		_w910_,
		_w4937_
	);
	LUT2 #(
		.INIT('h2)
	) name4475 (
		_w1183_,
		_w4937_,
		_w4938_
	);
	LUT4 #(
		.INIT('he010)
	) name4476 (
		_w1224_,
		_w1228_,
		_w1286_,
		_w1441_,
		_w4939_
	);
	LUT4 #(
		.INIT('h2822)
	) name4477 (
		_w1114_,
		_w1441_,
		_w2867_,
		_w2868_,
		_w4940_
	);
	LUT4 #(
		.INIT('h8000)
	) name4478 (
		_w894_,
		_w929_,
		_w938_,
		_w1115_,
		_w4941_
	);
	LUT4 #(
		.INIT('h7f00)
	) name4479 (
		_w894_,
		_w1115_,
		_w1116_,
		_w1136_,
		_w4942_
	);
	LUT3 #(
		.INIT('he0)
	) name4480 (
		_w918_,
		_w4941_,
		_w4942_,
		_w4943_
	);
	LUT4 #(
		.INIT('haaa8)
	) name4481 (
		_w2197_,
		_w4940_,
		_w4943_,
		_w4939_,
		_w4944_
	);
	LUT3 #(
		.INIT('h04)
	) name4482 (
		_w918_,
		_w2259_,
		_w2260_,
		_w4945_
	);
	LUT3 #(
		.INIT('h0d)
	) name4483 (
		_w910_,
		_w4545_,
		_w4945_,
		_w4946_
	);
	LUT4 #(
		.INIT('h0b00)
	) name4484 (
		_w4936_,
		_w4938_,
		_w4944_,
		_w4946_,
		_w4947_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name4485 (
		\P1_state_reg[0]/NET0131 ,
		_w526_,
		_w4934_,
		_w4947_,
		_w4948_
	);
	LUT2 #(
		.INIT('h2)
	) name4486 (
		\P1_reg3_reg[7]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w4949_
	);
	LUT3 #(
		.INIT('h07)
	) name4487 (
		_w910_,
		_w1294_,
		_w4949_,
		_w4950_
	);
	LUT2 #(
		.INIT('hb)
	) name4488 (
		_w4948_,
		_w4950_,
		_w4951_
	);
	LUT2 #(
		.INIT('h2)
	) name4489 (
		_w1487_,
		_w1584_,
		_w4952_
	);
	LUT4 #(
		.INIT('h00fe)
	) name4490 (
		_w1491_,
		_w1493_,
		_w1496_,
		_w1584_,
		_w4953_
	);
	LUT3 #(
		.INIT('h10)
	) name4491 (
		_w1586_,
		_w1599_,
		_w2057_,
		_w4954_
	);
	LUT4 #(
		.INIT('h0100)
	) name4492 (
		_w1502_,
		_w1586_,
		_w1599_,
		_w2057_,
		_w4955_
	);
	LUT3 #(
		.INIT('h70)
	) name4493 (
		_w1597_,
		_w1598_,
		_w2042_,
		_w4956_
	);
	LUT4 #(
		.INIT('h00de)
	) name4494 (
		_w1502_,
		_w2042_,
		_w4954_,
		_w4956_,
		_w4957_
	);
	LUT4 #(
		.INIT('h04c4)
	) name4495 (
		_w1584_,
		_w2081_,
		_w2277_,
		_w4957_,
		_w4958_
	);
	LUT3 #(
		.INIT('h87)
	) name4496 (
		_w1583_,
		_w1585_,
		_w1593_,
		_w4959_
	);
	LUT4 #(
		.INIT('h00d7)
	) name4497 (
		_w2277_,
		_w2304_,
		_w4959_,
		_w4953_,
		_w4960_
	);
	LUT2 #(
		.INIT('h2)
	) name4498 (
		_w2290_,
		_w4960_,
		_w4961_
	);
	LUT4 #(
		.INIT('h001f)
	) name4499 (
		_w1491_,
		_w1493_,
		_w1496_,
		_w1584_,
		_w4962_
	);
	LUT4 #(
		.INIT('h0d07)
	) name4500 (
		_w2272_,
		_w2304_,
		_w4962_,
		_w4959_,
		_w4963_
	);
	LUT2 #(
		.INIT('h1)
	) name4501 (
		_w2276_,
		_w4963_,
		_w4964_
	);
	LUT4 #(
		.INIT('h0545)
	) name4502 (
		_w2107_,
		_w2111_,
		_w2352_,
		_w2353_,
		_w4965_
	);
	LUT4 #(
		.INIT('h3113)
	) name4503 (
		_w2272_,
		_w4962_,
		_w4959_,
		_w4965_,
		_w4966_
	);
	LUT3 #(
		.INIT('h04)
	) name4504 (
		_w1593_,
		_w2083_,
		_w2282_,
		_w4967_
	);
	LUT3 #(
		.INIT('h54)
	) name4505 (
		_w1584_,
		_w2086_,
		_w2280_,
		_w4968_
	);
	LUT2 #(
		.INIT('h1)
	) name4506 (
		_w4967_,
		_w4968_,
		_w4969_
	);
	LUT3 #(
		.INIT('he0)
	) name4507 (
		_w2192_,
		_w4966_,
		_w4969_,
		_w4970_
	);
	LUT4 #(
		.INIT('h0100)
	) name4508 (
		_w4964_,
		_w4961_,
		_w4958_,
		_w4970_,
		_w4971_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name4509 (
		\P1_state_reg[0]/NET0131 ,
		_w1489_,
		_w4952_,
		_w4971_,
		_w4972_
	);
	LUT2 #(
		.INIT('h4)
	) name4510 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[5]/NET0131 ,
		_w4973_
	);
	LUT4 #(
		.INIT('h0028)
	) name4511 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		_w1476_,
		_w1584_,
		_w4974_
	);
	LUT2 #(
		.INIT('h1)
	) name4512 (
		_w4973_,
		_w4974_,
		_w4975_
	);
	LUT2 #(
		.INIT('hb)
	) name4513 (
		_w4972_,
		_w4975_,
		_w4976_
	);
	LUT2 #(
		.INIT('h4)
	) name4514 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[6]/NET0131 ,
		_w4977_
	);
	LUT4 #(
		.INIT('h00fe)
	) name4515 (
		_w1491_,
		_w1493_,
		_w1496_,
		_w1500_,
		_w4978_
	);
	LUT3 #(
		.INIT('h70)
	) name4516 (
		_w1583_,
		_w1585_,
		_w2042_,
		_w4979_
	);
	LUT3 #(
		.INIT('h15)
	) name4517 (
		_w2042_,
		_w2057_,
		_w2060_,
		_w4980_
	);
	LUT4 #(
		.INIT('h020f)
	) name4518 (
		_w1532_,
		_w4955_,
		_w4979_,
		_w4980_,
		_w4981_
	);
	LUT4 #(
		.INIT('h04c4)
	) name4519 (
		_w1500_,
		_w2081_,
		_w2277_,
		_w4981_,
		_w4982_
	);
	LUT4 #(
		.INIT('h001f)
	) name4520 (
		_w1491_,
		_w1493_,
		_w1496_,
		_w1500_,
		_w4983_
	);
	LUT3 #(
		.INIT('h87)
	) name4521 (
		_w1499_,
		_w1501_,
		_w1527_,
		_w4984_
	);
	LUT4 #(
		.INIT('h40b0)
	) name4522 (
		_w2117_,
		_w2120_,
		_w2272_,
		_w4984_,
		_w4985_
	);
	LUT4 #(
		.INIT('h00e0)
	) name4523 (
		_w1491_,
		_w1493_,
		_w1496_,
		_w1527_,
		_w4986_
	);
	LUT3 #(
		.INIT('ha8)
	) name4524 (
		_w2084_,
		_w4983_,
		_w4986_,
		_w4987_
	);
	LUT2 #(
		.INIT('h4)
	) name4525 (
		_w1527_,
		_w2088_,
		_w4988_
	);
	LUT4 #(
		.INIT('h3332)
	) name4526 (
		_w1487_,
		_w1500_,
		_w2086_,
		_w2293_,
		_w4989_
	);
	LUT2 #(
		.INIT('h1)
	) name4527 (
		_w4988_,
		_w4989_,
		_w4990_
	);
	LUT2 #(
		.INIT('h4)
	) name4528 (
		_w4987_,
		_w4990_,
		_w4991_
	);
	LUT4 #(
		.INIT('hab00)
	) name4529 (
		_w2192_,
		_w4983_,
		_w4985_,
		_w4991_,
		_w4992_
	);
	LUT4 #(
		.INIT('he010)
	) name4530 (
		_w1608_,
		_w1611_,
		_w2277_,
		_w4984_,
		_w4993_
	);
	LUT3 #(
		.INIT('ha8)
	) name4531 (
		_w2290_,
		_w4978_,
		_w4993_,
		_w4994_
	);
	LUT4 #(
		.INIT('he010)
	) name4532 (
		_w1608_,
		_w1611_,
		_w2272_,
		_w4984_,
		_w4995_
	);
	LUT3 #(
		.INIT('h54)
	) name4533 (
		_w2276_,
		_w4983_,
		_w4995_,
		_w4996_
	);
	LUT4 #(
		.INIT('h0100)
	) name4534 (
		_w4982_,
		_w4994_,
		_w4996_,
		_w4992_,
		_w4997_
	);
	LUT3 #(
		.INIT('h8a)
	) name4535 (
		\P1_state_reg[0]/NET0131 ,
		_w1489_,
		_w1500_,
		_w4998_
	);
	LUT3 #(
		.INIT('hba)
	) name4536 (
		_w4977_,
		_w4997_,
		_w4998_,
		_w4999_
	);
	LUT2 #(
		.INIT('h2)
	) name4537 (
		_w1487_,
		_w1530_,
		_w5000_
	);
	LUT4 #(
		.INIT('h00fe)
	) name4538 (
		_w1491_,
		_w1493_,
		_w1496_,
		_w1530_,
		_w5001_
	);
	LUT3 #(
		.INIT('h78)
	) name4539 (
		_w1529_,
		_w1531_,
		_w1545_,
		_w5002_
	);
	LUT4 #(
		.INIT('h0df2)
	) name4540 (
		_w2302_,
		_w2304_,
		_w2305_,
		_w5002_,
		_w5003_
	);
	LUT4 #(
		.INIT('hd010)
	) name4541 (
		_w1530_,
		_w2277_,
		_w2290_,
		_w5003_,
		_w5004_
	);
	LUT4 #(
		.INIT('h001f)
	) name4542 (
		_w1491_,
		_w1493_,
		_w1496_,
		_w1530_,
		_w5005_
	);
	LUT4 #(
		.INIT('h0d01)
	) name4543 (
		_w1530_,
		_w2272_,
		_w2276_,
		_w5003_,
		_w5006_
	);
	LUT4 #(
		.INIT('h2111)
	) name4544 (
		_w1676_,
		_w2042_,
		_w2057_,
		_w2060_,
		_w5007_
	);
	LUT3 #(
		.INIT('h70)
	) name4545 (
		_w1499_,
		_w1501_,
		_w2042_,
		_w5008_
	);
	LUT4 #(
		.INIT('h1113)
	) name4546 (
		_w2277_,
		_w5001_,
		_w5007_,
		_w5008_,
		_w5009_
	);
	LUT2 #(
		.INIT('h2)
	) name4547 (
		_w2081_,
		_w5009_,
		_w5010_
	);
	LUT4 #(
		.INIT('ha802)
	) name4548 (
		_w2272_,
		_w2351_,
		_w2355_,
		_w5002_,
		_w5011_
	);
	LUT3 #(
		.INIT('h04)
	) name4549 (
		_w1545_,
		_w2083_,
		_w2282_,
		_w5012_
	);
	LUT3 #(
		.INIT('h54)
	) name4550 (
		_w1530_,
		_w2086_,
		_w2280_,
		_w5013_
	);
	LUT2 #(
		.INIT('h1)
	) name4551 (
		_w5012_,
		_w5013_,
		_w5014_
	);
	LUT4 #(
		.INIT('hab00)
	) name4552 (
		_w2192_,
		_w5005_,
		_w5011_,
		_w5014_,
		_w5015_
	);
	LUT4 #(
		.INIT('h0100)
	) name4553 (
		_w5006_,
		_w5004_,
		_w5010_,
		_w5015_,
		_w5016_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name4554 (
		\P1_state_reg[0]/NET0131 ,
		_w1489_,
		_w5000_,
		_w5016_,
		_w5017_
	);
	LUT2 #(
		.INIT('h4)
	) name4555 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[7]/NET0131 ,
		_w5018_
	);
	LUT4 #(
		.INIT('h0028)
	) name4556 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		_w1476_,
		_w1530_,
		_w5019_
	);
	LUT2 #(
		.INIT('h1)
	) name4557 (
		_w5018_,
		_w5019_,
		_w5020_
	);
	LUT2 #(
		.INIT('hb)
	) name4558 (
		_w5017_,
		_w5020_,
		_w5021_
	);
	LUT2 #(
		.INIT('h2)
	) name4559 (
		\P1_reg2_reg[4]/NET0131 ,
		_w511_,
		_w5022_
	);
	LUT2 #(
		.INIT('h8)
	) name4560 (
		\P1_reg2_reg[4]/NET0131 ,
		_w524_,
		_w5023_
	);
	LUT4 #(
		.INIT('h0010)
	) name4561 (
		_w4540_,
		_w4538_,
		_w4543_,
		_w4844_,
		_w5024_
	);
	LUT3 #(
		.INIT('hab)
	) name4562 (
		_w534_,
		_w1109_,
		_w1183_,
		_w5025_
	);
	LUT2 #(
		.INIT('h8)
	) name4563 (
		_w885_,
		_w1143_,
		_w5026_
	);
	LUT4 #(
		.INIT('h00d5)
	) name4564 (
		\P1_reg2_reg[4]/NET0131 ,
		_w2411_,
		_w5025_,
		_w5026_,
		_w5027_
	);
	LUT4 #(
		.INIT('h08aa)
	) name4565 (
		_w526_,
		_w534_,
		_w5024_,
		_w5027_,
		_w5028_
	);
	LUT4 #(
		.INIT('heeec)
	) name4566 (
		\P1_state_reg[0]/NET0131 ,
		_w5022_,
		_w5023_,
		_w5028_,
		_w5029_
	);
	LUT3 #(
		.INIT('h2a)
	) name4567 (
		\P1_reg2_reg[11]/NET0131 ,
		_w3443_,
		_w3603_,
		_w5030_
	);
	LUT2 #(
		.INIT('h8)
	) name4568 (
		_w796_,
		_w1143_,
		_w5031_
	);
	LUT3 #(
		.INIT('h28)
	) name4569 (
		_w1286_,
		_w1453_,
		_w2843_,
		_w5032_
	);
	LUT2 #(
		.INIT('h4)
	) name4570 (
		_w804_,
		_w1138_,
		_w5033_
	);
	LUT2 #(
		.INIT('h1)
	) name4571 (
		_w4445_,
		_w5033_,
		_w5034_
	);
	LUT4 #(
		.INIT('h7d00)
	) name4572 (
		_w1114_,
		_w1453_,
		_w2871_,
		_w5034_,
		_w5035_
	);
	LUT4 #(
		.INIT('h0700)
	) name4573 (
		_w1183_,
		_w4440_,
		_w5032_,
		_w5035_,
		_w5036_
	);
	LUT4 #(
		.INIT('hc0c8)
	) name4574 (
		_w534_,
		_w3443_,
		_w5031_,
		_w5036_,
		_w5037_
	);
	LUT2 #(
		.INIT('he)
	) name4575 (
		_w5030_,
		_w5037_,
		_w5038_
	);
	LUT4 #(
		.INIT('h70d0)
	) name4576 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg1_reg[11]/NET0131 ,
		_w1476_,
		_w5039_
	);
	LUT2 #(
		.INIT('h8)
	) name4577 (
		\P2_reg1_reg[11]/NET0131 ,
		_w1487_,
		_w5040_
	);
	LUT4 #(
		.INIT('h20e0)
	) name4578 (
		\P2_reg1_reg[11]/NET0131 ,
		_w1497_,
		_w2081_,
		_w4486_,
		_w5041_
	);
	LUT4 #(
		.INIT('haa02)
	) name4579 (
		\P2_reg1_reg[11]/NET0131 ,
		_w1491_,
		_w1493_,
		_w1496_,
		_w5042_
	);
	LUT4 #(
		.INIT('h8a20)
	) name4580 (
		_w2039_,
		_w2309_,
		_w2312_,
		_w4474_,
		_w5043_
	);
	LUT3 #(
		.INIT('ha8)
	) name4581 (
		_w2038_,
		_w5042_,
		_w5043_,
		_w5044_
	);
	LUT4 #(
		.INIT('h1dd1)
	) name4582 (
		\P2_reg1_reg[11]/NET0131 ,
		_w2039_,
		_w2363_,
		_w4474_,
		_w5045_
	);
	LUT2 #(
		.INIT('h2)
	) name4583 (
		_w2193_,
		_w5045_,
		_w5046_
	);
	LUT4 #(
		.INIT('h1dd1)
	) name4584 (
		\P2_reg1_reg[11]/NET0131 ,
		_w1497_,
		_w2363_,
		_w4474_,
		_w5047_
	);
	LUT3 #(
		.INIT('he0)
	) name4585 (
		_w1638_,
		_w1640_,
		_w2084_,
		_w5048_
	);
	LUT2 #(
		.INIT('h8)
	) name4586 (
		_w2039_,
		_w5048_,
		_w5049_
	);
	LUT3 #(
		.INIT('ha2)
	) name4587 (
		\P2_reg1_reg[11]/NET0131 ,
		_w2633_,
		_w2660_,
		_w5050_
	);
	LUT2 #(
		.INIT('h1)
	) name4588 (
		_w5049_,
		_w5050_,
		_w5051_
	);
	LUT3 #(
		.INIT('hd0)
	) name4589 (
		_w2188_,
		_w5047_,
		_w5051_,
		_w5052_
	);
	LUT4 #(
		.INIT('h0100)
	) name4590 (
		_w5044_,
		_w5041_,
		_w5046_,
		_w5052_,
		_w5053_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name4591 (
		\P1_state_reg[0]/NET0131 ,
		_w1489_,
		_w5040_,
		_w5053_,
		_w5054_
	);
	LUT2 #(
		.INIT('he)
	) name4592 (
		_w5039_,
		_w5054_,
		_w5055_
	);
	LUT4 #(
		.INIT('h70d0)
	) name4593 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg1_reg[14]/NET0131 ,
		_w1476_,
		_w5056_
	);
	LUT2 #(
		.INIT('h8)
	) name4594 (
		\P2_reg1_reg[14]/NET0131 ,
		_w1487_,
		_w5057_
	);
	LUT4 #(
		.INIT('h08c8)
	) name4595 (
		\P2_reg1_reg[14]/NET0131 ,
		_w2038_,
		_w2039_,
		_w4506_,
		_w5058_
	);
	LUT4 #(
		.INIT('h20e0)
	) name4596 (
		\P2_reg1_reg[14]/NET0131 ,
		_w1497_,
		_w2081_,
		_w4499_,
		_w5059_
	);
	LUT4 #(
		.INIT('hf100)
	) name4597 (
		_w1509_,
		_w1727_,
		_w1729_,
		_w2084_,
		_w5060_
	);
	LUT2 #(
		.INIT('h8)
	) name4598 (
		_w2039_,
		_w5060_,
		_w5061_
	);
	LUT3 #(
		.INIT('ha2)
	) name4599 (
		\P2_reg1_reg[14]/NET0131 ,
		_w2633_,
		_w2660_,
		_w5062_
	);
	LUT2 #(
		.INIT('h1)
	) name4600 (
		_w5061_,
		_w5062_,
		_w5063_
	);
	LUT2 #(
		.INIT('h4)
	) name4601 (
		_w5059_,
		_w5063_,
		_w5064_
	);
	LUT2 #(
		.INIT('h4)
	) name4602 (
		_w5058_,
		_w5064_,
		_w5065_
	);
	LUT4 #(
		.INIT('h1dd1)
	) name4603 (
		\P2_reg1_reg[14]/NET0131 ,
		_w2039_,
		_w2794_,
		_w4496_,
		_w5066_
	);
	LUT4 #(
		.INIT('h1dd1)
	) name4604 (
		\P2_reg1_reg[14]/NET0131 ,
		_w1497_,
		_w2794_,
		_w4496_,
		_w5067_
	);
	LUT4 #(
		.INIT('hf351)
	) name4605 (
		_w2188_,
		_w2193_,
		_w5066_,
		_w5067_,
		_w5068_
	);
	LUT4 #(
		.INIT('h3111)
	) name4606 (
		_w1489_,
		_w5057_,
		_w5065_,
		_w5068_,
		_w5069_
	);
	LUT3 #(
		.INIT('hce)
	) name4607 (
		\P1_state_reg[0]/NET0131 ,
		_w5056_,
		_w5069_,
		_w5070_
	);
	LUT4 #(
		.INIT('h70d0)
	) name4608 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg1_reg[15]/NET0131 ,
		_w1476_,
		_w5071_
	);
	LUT2 #(
		.INIT('h8)
	) name4609 (
		\P2_reg1_reg[15]/NET0131 ,
		_w1487_,
		_w5072_
	);
	LUT4 #(
		.INIT('h1dd1)
	) name4610 (
		\P2_reg1_reg[15]/NET0131 ,
		_w2039_,
		_w3512_,
		_w4516_,
		_w5073_
	);
	LUT2 #(
		.INIT('h2)
	) name4611 (
		_w2038_,
		_w5073_,
		_w5074_
	);
	LUT4 #(
		.INIT('h20e0)
	) name4612 (
		\P2_reg1_reg[15]/NET0131 ,
		_w2039_,
		_w2193_,
		_w4521_,
		_w5075_
	);
	LUT4 #(
		.INIT('h20e0)
	) name4613 (
		\P2_reg1_reg[15]/NET0131 ,
		_w1497_,
		_w2188_,
		_w4521_,
		_w5076_
	);
	LUT4 #(
		.INIT('h111d)
	) name4614 (
		\P2_reg1_reg[15]/NET0131 ,
		_w1497_,
		_w4523_,
		_w4525_,
		_w5077_
	);
	LUT4 #(
		.INIT('hf100)
	) name4615 (
		_w1509_,
		_w1711_,
		_w1714_,
		_w2084_,
		_w5078_
	);
	LUT2 #(
		.INIT('h8)
	) name4616 (
		_w2039_,
		_w5078_,
		_w5079_
	);
	LUT3 #(
		.INIT('ha2)
	) name4617 (
		\P2_reg1_reg[15]/NET0131 ,
		_w2633_,
		_w2660_,
		_w5080_
	);
	LUT2 #(
		.INIT('h1)
	) name4618 (
		_w5079_,
		_w5080_,
		_w5081_
	);
	LUT3 #(
		.INIT('hd0)
	) name4619 (
		_w2081_,
		_w5077_,
		_w5081_,
		_w5082_
	);
	LUT3 #(
		.INIT('h10)
	) name4620 (
		_w5076_,
		_w5075_,
		_w5082_,
		_w5083_
	);
	LUT4 #(
		.INIT('h1311)
	) name4621 (
		_w1489_,
		_w5072_,
		_w5074_,
		_w5083_,
		_w5084_
	);
	LUT3 #(
		.INIT('hce)
	) name4622 (
		\P1_state_reg[0]/NET0131 ,
		_w5071_,
		_w5084_,
		_w5085_
	);
	LUT2 #(
		.INIT('h2)
	) name4623 (
		\P1_reg0_reg[10]/NET0131 ,
		_w511_,
		_w5086_
	);
	LUT2 #(
		.INIT('h8)
	) name4624 (
		\P1_reg0_reg[10]/NET0131 ,
		_w524_,
		_w5087_
	);
	LUT4 #(
		.INIT('haaa8)
	) name4625 (
		\P1_reg0_reg[10]/NET0131 ,
		_w528_,
		_w530_,
		_w533_,
		_w5088_
	);
	LUT4 #(
		.INIT('h7020)
	) name4626 (
		_w537_,
		_w833_,
		_w2688_,
		_w4084_,
		_w5089_
	);
	LUT3 #(
		.INIT('ha8)
	) name4627 (
		_w1183_,
		_w5088_,
		_w5089_,
		_w5090_
	);
	LUT4 #(
		.INIT('hc535)
	) name4628 (
		\P1_reg0_reg[10]/NET0131 ,
		_w1438_,
		_w2688_,
		_w3052_,
		_w5091_
	);
	LUT2 #(
		.INIT('h2)
	) name4629 (
		_w1114_,
		_w5091_,
		_w5092_
	);
	LUT4 #(
		.INIT('h35c5)
	) name4630 (
		\P1_reg0_reg[10]/NET0131 ,
		_w1438_,
		_w2688_,
		_w3076_,
		_w5093_
	);
	LUT4 #(
		.INIT('hc808)
	) name4631 (
		\P1_reg0_reg[10]/NET0131 ,
		_w1136_,
		_w2688_,
		_w4090_,
		_w5094_
	);
	LUT3 #(
		.INIT('h40)
	) name4632 (
		_w827_,
		_w1138_,
		_w2688_,
		_w5095_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name4633 (
		\P1_reg0_reg[10]/NET0131 ,
		_w1138_,
		_w2425_,
		_w2688_,
		_w5096_
	);
	LUT2 #(
		.INIT('h1)
	) name4634 (
		_w5095_,
		_w5096_,
		_w5097_
	);
	LUT2 #(
		.INIT('h4)
	) name4635 (
		_w5094_,
		_w5097_,
		_w5098_
	);
	LUT3 #(
		.INIT('hd0)
	) name4636 (
		_w1286_,
		_w5093_,
		_w5098_,
		_w5099_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name4637 (
		_w526_,
		_w5090_,
		_w5092_,
		_w5099_,
		_w5100_
	);
	LUT4 #(
		.INIT('heeec)
	) name4638 (
		\P1_state_reg[0]/NET0131 ,
		_w5086_,
		_w5087_,
		_w5100_,
		_w5101_
	);
	LUT2 #(
		.INIT('h2)
	) name4639 (
		_w1286_,
		_w2688_,
		_w5102_
	);
	LUT4 #(
		.INIT('hf700)
	) name4640 (
		_w1108_,
		_w1140_,
		_w2688_,
		_w3443_,
		_w5103_
	);
	LUT4 #(
		.INIT('h0200)
	) name4641 (
		_w2692_,
		_w2991_,
		_w5102_,
		_w5103_,
		_w5104_
	);
	LUT2 #(
		.INIT('h2)
	) name4642 (
		\P1_reg0_reg[11]/NET0131 ,
		_w5104_,
		_w5105_
	);
	LUT3 #(
		.INIT('hf2)
	) name4643 (
		_w3651_,
		_w5036_,
		_w5105_,
		_w5106_
	);
	LUT4 #(
		.INIT('h70d0)
	) name4644 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg2_reg[11]/NET0131 ,
		_w1476_,
		_w5107_
	);
	LUT2 #(
		.INIT('h8)
	) name4645 (
		\P2_reg2_reg[11]/NET0131 ,
		_w1487_,
		_w5108_
	);
	LUT4 #(
		.INIT('h20e0)
	) name4646 (
		\P2_reg2_reg[11]/NET0131 ,
		_w2039_,
		_w2081_,
		_w4486_,
		_w5109_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name4647 (
		\P2_reg2_reg[11]/NET0131 ,
		_w1491_,
		_w1493_,
		_w1496_,
		_w5110_
	);
	LUT4 #(
		.INIT('h8a20)
	) name4648 (
		_w1497_,
		_w2309_,
		_w2312_,
		_w4474_,
		_w5111_
	);
	LUT3 #(
		.INIT('ha8)
	) name4649 (
		_w2038_,
		_w5110_,
		_w5111_,
		_w5112_
	);
	LUT4 #(
		.INIT('h1dd1)
	) name4650 (
		\P2_reg2_reg[11]/NET0131 ,
		_w1497_,
		_w2363_,
		_w4474_,
		_w5113_
	);
	LUT2 #(
		.INIT('h2)
	) name4651 (
		_w2193_,
		_w5113_,
		_w5114_
	);
	LUT4 #(
		.INIT('h1dd1)
	) name4652 (
		\P2_reg2_reg[11]/NET0131 ,
		_w2039_,
		_w2363_,
		_w4474_,
		_w5115_
	);
	LUT3 #(
		.INIT('ha8)
	) name4653 (
		\P2_reg2_reg[11]/NET0131 ,
		_w2086_,
		_w2087_,
		_w5116_
	);
	LUT2 #(
		.INIT('h4)
	) name4654 (
		_w1617_,
		_w2088_,
		_w5117_
	);
	LUT3 #(
		.INIT('h07)
	) name4655 (
		_w1497_,
		_w5048_,
		_w5117_,
		_w5118_
	);
	LUT2 #(
		.INIT('h4)
	) name4656 (
		_w5116_,
		_w5118_,
		_w5119_
	);
	LUT3 #(
		.INIT('hd0)
	) name4657 (
		_w2188_,
		_w5115_,
		_w5119_,
		_w5120_
	);
	LUT4 #(
		.INIT('h0100)
	) name4658 (
		_w5112_,
		_w5109_,
		_w5114_,
		_w5120_,
		_w5121_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name4659 (
		\P1_state_reg[0]/NET0131 ,
		_w1489_,
		_w5108_,
		_w5121_,
		_w5122_
	);
	LUT2 #(
		.INIT('he)
	) name4660 (
		_w5107_,
		_w5122_,
		_w5123_
	);
	LUT4 #(
		.INIT('h70d0)
	) name4661 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg2_reg[14]/NET0131 ,
		_w1476_,
		_w5124_
	);
	LUT2 #(
		.INIT('h8)
	) name4662 (
		\P2_reg2_reg[14]/NET0131 ,
		_w1487_,
		_w5125_
	);
	LUT4 #(
		.INIT('h20e0)
	) name4663 (
		\P2_reg2_reg[14]/NET0131 ,
		_w1497_,
		_w2038_,
		_w4506_,
		_w5126_
	);
	LUT4 #(
		.INIT('h20e0)
	) name4664 (
		\P2_reg2_reg[14]/NET0131 ,
		_w2039_,
		_w2081_,
		_w4499_,
		_w5127_
	);
	LUT3 #(
		.INIT('ha8)
	) name4665 (
		\P2_reg2_reg[14]/NET0131 ,
		_w2086_,
		_w2087_,
		_w5128_
	);
	LUT2 #(
		.INIT('h4)
	) name4666 (
		_w1718_,
		_w2088_,
		_w5129_
	);
	LUT3 #(
		.INIT('h07)
	) name4667 (
		_w1497_,
		_w5060_,
		_w5129_,
		_w5130_
	);
	LUT2 #(
		.INIT('h4)
	) name4668 (
		_w5128_,
		_w5130_,
		_w5131_
	);
	LUT2 #(
		.INIT('h4)
	) name4669 (
		_w5127_,
		_w5131_,
		_w5132_
	);
	LUT2 #(
		.INIT('h4)
	) name4670 (
		_w5126_,
		_w5132_,
		_w5133_
	);
	LUT4 #(
		.INIT('h1dd1)
	) name4671 (
		\P2_reg2_reg[14]/NET0131 ,
		_w1497_,
		_w2794_,
		_w4496_,
		_w5134_
	);
	LUT4 #(
		.INIT('h1dd1)
	) name4672 (
		\P2_reg2_reg[14]/NET0131 ,
		_w2039_,
		_w2794_,
		_w4496_,
		_w5135_
	);
	LUT4 #(
		.INIT('hf351)
	) name4673 (
		_w2188_,
		_w2193_,
		_w5134_,
		_w5135_,
		_w5136_
	);
	LUT4 #(
		.INIT('h3111)
	) name4674 (
		_w1489_,
		_w5125_,
		_w5133_,
		_w5136_,
		_w5137_
	);
	LUT3 #(
		.INIT('hce)
	) name4675 (
		\P1_state_reg[0]/NET0131 ,
		_w5124_,
		_w5137_,
		_w5138_
	);
	LUT4 #(
		.INIT('h70d0)
	) name4676 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg2_reg[15]/NET0131 ,
		_w1476_,
		_w5139_
	);
	LUT2 #(
		.INIT('h8)
	) name4677 (
		\P2_reg2_reg[15]/NET0131 ,
		_w1487_,
		_w5140_
	);
	LUT4 #(
		.INIT('h1dd1)
	) name4678 (
		\P2_reg2_reg[15]/NET0131 ,
		_w1497_,
		_w3512_,
		_w4516_,
		_w5141_
	);
	LUT2 #(
		.INIT('h2)
	) name4679 (
		_w2038_,
		_w5141_,
		_w5142_
	);
	LUT4 #(
		.INIT('h20e0)
	) name4680 (
		\P2_reg2_reg[15]/NET0131 ,
		_w2039_,
		_w2188_,
		_w4521_,
		_w5143_
	);
	LUT4 #(
		.INIT('h20e0)
	) name4681 (
		\P2_reg2_reg[15]/NET0131 ,
		_w1497_,
		_w2193_,
		_w4521_,
		_w5144_
	);
	LUT4 #(
		.INIT('h111d)
	) name4682 (
		\P2_reg2_reg[15]/NET0131 ,
		_w2039_,
		_w4523_,
		_w4525_,
		_w5145_
	);
	LUT3 #(
		.INIT('ha8)
	) name4683 (
		\P2_reg2_reg[15]/NET0131 ,
		_w2086_,
		_w2087_,
		_w5146_
	);
	LUT2 #(
		.INIT('h4)
	) name4684 (
		_w1693_,
		_w2088_,
		_w5147_
	);
	LUT3 #(
		.INIT('h07)
	) name4685 (
		_w1497_,
		_w5078_,
		_w5147_,
		_w5148_
	);
	LUT2 #(
		.INIT('h4)
	) name4686 (
		_w5146_,
		_w5148_,
		_w5149_
	);
	LUT3 #(
		.INIT('hd0)
	) name4687 (
		_w2081_,
		_w5145_,
		_w5149_,
		_w5150_
	);
	LUT3 #(
		.INIT('h10)
	) name4688 (
		_w5144_,
		_w5143_,
		_w5150_,
		_w5151_
	);
	LUT4 #(
		.INIT('h1311)
	) name4689 (
		_w1489_,
		_w5140_,
		_w5142_,
		_w5151_,
		_w5152_
	);
	LUT3 #(
		.INIT('hce)
	) name4690 (
		\P1_state_reg[0]/NET0131 ,
		_w5139_,
		_w5152_,
		_w5153_
	);
	LUT2 #(
		.INIT('h2)
	) name4691 (
		\P1_reg0_reg[13]/NET0131 ,
		_w4051_,
		_w5154_
	);
	LUT4 #(
		.INIT('hff8a)
	) name4692 (
		_w3651_,
		_w4629_,
		_w4634_,
		_w5154_,
		_w5155_
	);
	LUT2 #(
		.INIT('h2)
	) name4693 (
		\P1_reg0_reg[14]/NET0131 ,
		_w511_,
		_w5156_
	);
	LUT2 #(
		.INIT('h8)
	) name4694 (
		\P1_reg0_reg[14]/NET0131 ,
		_w524_,
		_w5157_
	);
	LUT4 #(
		.INIT('haaa2)
	) name4695 (
		\P1_reg0_reg[14]/NET0131 ,
		_w2692_,
		_w3005_,
		_w3664_,
		_w5158_
	);
	LUT3 #(
		.INIT('h02)
	) name4696 (
		_w1183_,
		_w4103_,
		_w4104_,
		_w5159_
	);
	LUT2 #(
		.INIT('h2)
	) name4697 (
		_w1114_,
		_w4109_,
		_w5160_
	);
	LUT3 #(
		.INIT('h70)
	) name4698 (
		_w1286_,
		_w4107_,
		_w4646_,
		_w5161_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name4699 (
		_w2688_,
		_w5160_,
		_w5159_,
		_w5161_,
		_w5162_
	);
	LUT4 #(
		.INIT('h1113)
	) name4700 (
		_w526_,
		_w5157_,
		_w5158_,
		_w5162_,
		_w5163_
	);
	LUT3 #(
		.INIT('hce)
	) name4701 (
		\P1_state_reg[0]/NET0131 ,
		_w5156_,
		_w5163_,
		_w5164_
	);
	LUT3 #(
		.INIT('ha2)
	) name4702 (
		\P1_reg0_reg[5]/NET0131 ,
		_w3658_,
		_w3659_,
		_w5165_
	);
	LUT2 #(
		.INIT('h8)
	) name4703 (
		_w1183_,
		_w4555_,
		_w5166_
	);
	LUT4 #(
		.INIT('h0001)
	) name4704 (
		_w938_,
		_w1104_,
		_w1106_,
		_w1111_,
		_w5167_
	);
	LUT3 #(
		.INIT('h04)
	) name4705 (
		_w4561_,
		_w4563_,
		_w5167_,
		_w5168_
	);
	LUT4 #(
		.INIT('hecee)
	) name4706 (
		_w3651_,
		_w5165_,
		_w5166_,
		_w5168_,
		_w5169_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name4707 (
		\P1_reg1_reg[11]/NET0131 ,
		_w3684_,
		_w3685_,
		_w4075_,
		_w5170_
	);
	LUT3 #(
		.INIT('hf2)
	) name4708 (
		_w4074_,
		_w5036_,
		_w5170_,
		_w5171_
	);
	LUT2 #(
		.INIT('h2)
	) name4709 (
		\P1_reg1_reg[10]/NET0131 ,
		_w511_,
		_w5172_
	);
	LUT2 #(
		.INIT('h8)
	) name4710 (
		\P1_reg1_reg[10]/NET0131 ,
		_w524_,
		_w5173_
	);
	LUT4 #(
		.INIT('haa02)
	) name4711 (
		\P1_reg1_reg[10]/NET0131 ,
		_w528_,
		_w530_,
		_w533_,
		_w5174_
	);
	LUT4 #(
		.INIT('h7020)
	) name4712 (
		_w537_,
		_w833_,
		_w2421_,
		_w4084_,
		_w5175_
	);
	LUT3 #(
		.INIT('ha8)
	) name4713 (
		_w1183_,
		_w5174_,
		_w5175_,
		_w5176_
	);
	LUT4 #(
		.INIT('hc535)
	) name4714 (
		\P1_reg1_reg[10]/NET0131 ,
		_w1438_,
		_w2421_,
		_w3052_,
		_w5177_
	);
	LUT2 #(
		.INIT('h2)
	) name4715 (
		_w1114_,
		_w5177_,
		_w5178_
	);
	LUT4 #(
		.INIT('h35c5)
	) name4716 (
		\P1_reg1_reg[10]/NET0131 ,
		_w1438_,
		_w2421_,
		_w3076_,
		_w5179_
	);
	LUT4 #(
		.INIT('hc808)
	) name4717 (
		\P1_reg1_reg[10]/NET0131 ,
		_w1136_,
		_w2421_,
		_w4090_,
		_w5180_
	);
	LUT3 #(
		.INIT('h40)
	) name4718 (
		_w827_,
		_w1138_,
		_w2421_,
		_w5181_
	);
	LUT4 #(
		.INIT('h08aa)
	) name4719 (
		\P1_reg1_reg[10]/NET0131 ,
		_w1138_,
		_w2421_,
		_w2425_,
		_w5182_
	);
	LUT2 #(
		.INIT('h1)
	) name4720 (
		_w5181_,
		_w5182_,
		_w5183_
	);
	LUT2 #(
		.INIT('h4)
	) name4721 (
		_w5180_,
		_w5183_,
		_w5184_
	);
	LUT3 #(
		.INIT('hd0)
	) name4722 (
		_w1286_,
		_w5179_,
		_w5184_,
		_w5185_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name4723 (
		_w526_,
		_w5176_,
		_w5178_,
		_w5185_,
		_w5186_
	);
	LUT4 #(
		.INIT('heeec)
	) name4724 (
		\P1_state_reg[0]/NET0131 ,
		_w5172_,
		_w5173_,
		_w5186_,
		_w5187_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name4725 (
		\P1_reg1_reg[13]/NET0131 ,
		_w3684_,
		_w3685_,
		_w4075_,
		_w5188_
	);
	LUT4 #(
		.INIT('hff8a)
	) name4726 (
		_w4074_,
		_w4629_,
		_w4634_,
		_w5188_,
		_w5189_
	);
	LUT2 #(
		.INIT('h2)
	) name4727 (
		\P1_reg1_reg[14]/NET0131 ,
		_w511_,
		_w5190_
	);
	LUT2 #(
		.INIT('h8)
	) name4728 (
		\P1_reg1_reg[14]/NET0131 ,
		_w524_,
		_w5191_
	);
	LUT3 #(
		.INIT('h2a)
	) name4729 (
		\P1_reg1_reg[14]/NET0131 ,
		_w2426_,
		_w3686_,
		_w5192_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name4730 (
		_w2421_,
		_w5160_,
		_w5159_,
		_w5161_,
		_w5193_
	);
	LUT4 #(
		.INIT('h1113)
	) name4731 (
		_w526_,
		_w5191_,
		_w5192_,
		_w5193_,
		_w5194_
	);
	LUT3 #(
		.INIT('hce)
	) name4732 (
		\P1_state_reg[0]/NET0131 ,
		_w5190_,
		_w5194_,
		_w5195_
	);
	LUT4 #(
		.INIT('h70d0)
	) name4733 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg0_reg[11]/NET0131 ,
		_w1476_,
		_w5196_
	);
	LUT2 #(
		.INIT('h8)
	) name4734 (
		\P2_reg0_reg[11]/NET0131 ,
		_w1487_,
		_w5197_
	);
	LUT4 #(
		.INIT('haaa8)
	) name4735 (
		\P2_reg0_reg[11]/NET0131 ,
		_w1491_,
		_w1493_,
		_w1496_,
		_w5198_
	);
	LUT3 #(
		.INIT('h54)
	) name4736 (
		_w2276_,
		_w4483_,
		_w5198_,
		_w5199_
	);
	LUT4 #(
		.INIT('h1dd1)
	) name4737 (
		\P2_reg0_reg[11]/NET0131 ,
		_w2277_,
		_w2363_,
		_w4474_,
		_w5200_
	);
	LUT2 #(
		.INIT('h8)
	) name4738 (
		_w2277_,
		_w5048_,
		_w5201_
	);
	LUT3 #(
		.INIT('ha2)
	) name4739 (
		\P2_reg0_reg[11]/NET0131 ,
		_w2633_,
		_w2634_,
		_w5202_
	);
	LUT2 #(
		.INIT('h1)
	) name4740 (
		_w5201_,
		_w5202_,
		_w5203_
	);
	LUT3 #(
		.INIT('he0)
	) name4741 (
		_w2192_,
		_w5200_,
		_w5203_,
		_w5204_
	);
	LUT4 #(
		.INIT('h02aa)
	) name4742 (
		\P2_reg0_reg[11]/NET0131 ,
		_w1491_,
		_w1493_,
		_w1496_,
		_w5205_
	);
	LUT3 #(
		.INIT('ha8)
	) name4743 (
		_w2290_,
		_w4475_,
		_w5205_,
		_w5206_
	);
	LUT4 #(
		.INIT('h08c8)
	) name4744 (
		\P2_reg0_reg[11]/NET0131 ,
		_w2081_,
		_w2272_,
		_w4486_,
		_w5207_
	);
	LUT4 #(
		.INIT('h0100)
	) name4745 (
		_w5199_,
		_w5206_,
		_w5207_,
		_w5204_,
		_w5208_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name4746 (
		\P1_state_reg[0]/NET0131 ,
		_w1489_,
		_w5197_,
		_w5208_,
		_w5209_
	);
	LUT2 #(
		.INIT('he)
	) name4747 (
		_w5196_,
		_w5209_,
		_w5210_
	);
	LUT4 #(
		.INIT('h70d0)
	) name4748 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg0_reg[14]/NET0131 ,
		_w1476_,
		_w5211_
	);
	LUT2 #(
		.INIT('h8)
	) name4749 (
		\P2_reg0_reg[14]/NET0131 ,
		_w1487_,
		_w5212_
	);
	LUT4 #(
		.INIT('h1dd1)
	) name4750 (
		\P2_reg0_reg[14]/NET0131 ,
		_w2277_,
		_w2794_,
		_w4496_,
		_w5213_
	);
	LUT4 #(
		.INIT('h08c8)
	) name4751 (
		\P2_reg0_reg[14]/NET0131 ,
		_w2081_,
		_w2272_,
		_w4499_,
		_w5214_
	);
	LUT2 #(
		.INIT('h8)
	) name4752 (
		_w2277_,
		_w5060_,
		_w5215_
	);
	LUT3 #(
		.INIT('ha2)
	) name4753 (
		\P2_reg0_reg[14]/NET0131 ,
		_w2633_,
		_w2634_,
		_w5216_
	);
	LUT2 #(
		.INIT('h1)
	) name4754 (
		_w5215_,
		_w5216_,
		_w5217_
	);
	LUT2 #(
		.INIT('h4)
	) name4755 (
		_w5214_,
		_w5217_,
		_w5218_
	);
	LUT3 #(
		.INIT('he0)
	) name4756 (
		_w2192_,
		_w5213_,
		_w5218_,
		_w5219_
	);
	LUT4 #(
		.INIT('h20e0)
	) name4757 (
		\P2_reg0_reg[14]/NET0131 ,
		_w2272_,
		_w2290_,
		_w4506_,
		_w5220_
	);
	LUT4 #(
		.INIT('h0232)
	) name4758 (
		\P2_reg0_reg[14]/NET0131 ,
		_w2276_,
		_w2277_,
		_w4506_,
		_w5221_
	);
	LUT2 #(
		.INIT('h1)
	) name4759 (
		_w5220_,
		_w5221_,
		_w5222_
	);
	LUT4 #(
		.INIT('h3111)
	) name4760 (
		_w1489_,
		_w5212_,
		_w5219_,
		_w5222_,
		_w5223_
	);
	LUT3 #(
		.INIT('hce)
	) name4761 (
		\P1_state_reg[0]/NET0131 ,
		_w5211_,
		_w5223_,
		_w5224_
	);
	LUT4 #(
		.INIT('h70d0)
	) name4762 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg0_reg[15]/NET0131 ,
		_w1476_,
		_w5225_
	);
	LUT2 #(
		.INIT('h8)
	) name4763 (
		\P2_reg0_reg[15]/NET0131 ,
		_w1487_,
		_w5226_
	);
	LUT4 #(
		.INIT('h1dd1)
	) name4764 (
		\P2_reg0_reg[15]/NET0131 ,
		_w2272_,
		_w3512_,
		_w4516_,
		_w5227_
	);
	LUT2 #(
		.INIT('h2)
	) name4765 (
		_w2290_,
		_w5227_,
		_w5228_
	);
	LUT4 #(
		.INIT('h1dd1)
	) name4766 (
		\P2_reg0_reg[15]/NET0131 ,
		_w2277_,
		_w3512_,
		_w4516_,
		_w5229_
	);
	LUT4 #(
		.INIT('h0232)
	) name4767 (
		\P2_reg0_reg[15]/NET0131 ,
		_w2192_,
		_w2277_,
		_w4521_,
		_w5230_
	);
	LUT4 #(
		.INIT('h111d)
	) name4768 (
		\P2_reg0_reg[15]/NET0131 ,
		_w2272_,
		_w4523_,
		_w4525_,
		_w5231_
	);
	LUT2 #(
		.INIT('h8)
	) name4769 (
		_w2277_,
		_w5078_,
		_w5232_
	);
	LUT3 #(
		.INIT('ha2)
	) name4770 (
		\P2_reg0_reg[15]/NET0131 ,
		_w2633_,
		_w2634_,
		_w5233_
	);
	LUT2 #(
		.INIT('h1)
	) name4771 (
		_w5232_,
		_w5233_,
		_w5234_
	);
	LUT3 #(
		.INIT('hd0)
	) name4772 (
		_w2081_,
		_w5231_,
		_w5234_,
		_w5235_
	);
	LUT4 #(
		.INIT('h0e00)
	) name4773 (
		_w2276_,
		_w5229_,
		_w5230_,
		_w5235_,
		_w5236_
	);
	LUT4 #(
		.INIT('h1311)
	) name4774 (
		_w1489_,
		_w5226_,
		_w5228_,
		_w5236_,
		_w5237_
	);
	LUT3 #(
		.INIT('hce)
	) name4775 (
		\P1_state_reg[0]/NET0131 ,
		_w5225_,
		_w5237_,
		_w5238_
	);
	LUT3 #(
		.INIT('h8a)
	) name4776 (
		\P1_reg1_reg[5]/NET0131 ,
		_w3065_,
		_w4075_,
		_w5239_
	);
	LUT4 #(
		.INIT('hff8a)
	) name4777 (
		_w4074_,
		_w5166_,
		_w5168_,
		_w5239_,
		_w5240_
	);
	LUT2 #(
		.INIT('h8)
	) name4778 (
		_w524_,
		_w922_,
		_w5241_
	);
	LUT4 #(
		.INIT('h1f00)
	) name4779 (
		_w528_,
		_w530_,
		_w533_,
		_w922_,
		_w5242_
	);
	LUT4 #(
		.INIT('h4144)
	) name4780 (
		_w537_,
		_w912_,
		_w924_,
		_w1154_,
		_w5243_
	);
	LUT3 #(
		.INIT('h80)
	) name4781 (
		_w537_,
		_w932_,
		_w933_,
		_w5244_
	);
	LUT4 #(
		.INIT('h3331)
	) name4782 (
		_w2197_,
		_w5242_,
		_w5243_,
		_w5244_,
		_w5245_
	);
	LUT4 #(
		.INIT('h3090)
	) name4783 (
		_w1366_,
		_w1448_,
		_w2197_,
		_w3073_,
		_w5246_
	);
	LUT3 #(
		.INIT('ha8)
	) name4784 (
		_w1286_,
		_w5242_,
		_w5246_,
		_w5247_
	);
	LUT4 #(
		.INIT('h8848)
	) name4785 (
		_w1448_,
		_w2197_,
		_w2225_,
		_w3049_,
		_w5248_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name4786 (
		_w894_,
		_w929_,
		_w938_,
		_w1115_,
		_w5249_
	);
	LUT4 #(
		.INIT('hc808)
	) name4787 (
		_w922_,
		_w1136_,
		_w2197_,
		_w5249_,
		_w5250_
	);
	LUT3 #(
		.INIT('h04)
	) name4788 (
		_w929_,
		_w2259_,
		_w2260_,
		_w5251_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name4789 (
		_w922_,
		_w1138_,
		_w1141_,
		_w2197_,
		_w5252_
	);
	LUT2 #(
		.INIT('h1)
	) name4790 (
		_w5251_,
		_w5252_,
		_w5253_
	);
	LUT2 #(
		.INIT('h4)
	) name4791 (
		_w5250_,
		_w5253_,
		_w5254_
	);
	LUT4 #(
		.INIT('h5700)
	) name4792 (
		_w1114_,
		_w5242_,
		_w5248_,
		_w5254_,
		_w5255_
	);
	LUT4 #(
		.INIT('h3100)
	) name4793 (
		_w1183_,
		_w5247_,
		_w5245_,
		_w5255_,
		_w5256_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name4794 (
		\P1_state_reg[0]/NET0131 ,
		_w526_,
		_w5241_,
		_w5256_,
		_w5257_
	);
	LUT2 #(
		.INIT('h2)
	) name4795 (
		\P1_reg3_reg[6]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w5258_
	);
	LUT3 #(
		.INIT('h07)
	) name4796 (
		_w922_,
		_w1294_,
		_w5258_,
		_w5259_
	);
	LUT2 #(
		.INIT('hb)
	) name4797 (
		_w5257_,
		_w5259_,
		_w5260_
	);
	LUT2 #(
		.INIT('h2)
	) name4798 (
		_w1487_,
		_w1596_,
		_w5261_
	);
	LUT4 #(
		.INIT('h001f)
	) name4799 (
		_w1491_,
		_w1493_,
		_w1496_,
		_w1596_,
		_w5262_
	);
	LUT3 #(
		.INIT('h78)
	) name4800 (
		_w1597_,
		_w1598_,
		_w1604_,
		_w5263_
	);
	LUT4 #(
		.INIT('h1117)
	) name4801 (
		_w1550_,
		_w1555_,
		_w1565_,
		_w1582_,
		_w5264_
	);
	LUT4 #(
		.INIT('h3113)
	) name4802 (
		_w2272_,
		_w5262_,
		_w5263_,
		_w5264_,
		_w5265_
	);
	LUT4 #(
		.INIT('h0df2)
	) name4803 (
		_w2111_,
		_w2113_,
		_w2116_,
		_w5263_,
		_w5266_
	);
	LUT4 #(
		.INIT('h0131)
	) name4804 (
		_w1596_,
		_w2192_,
		_w2272_,
		_w5266_,
		_w5267_
	);
	LUT3 #(
		.INIT('h04)
	) name4805 (
		_w1604_,
		_w2083_,
		_w2282_,
		_w5268_
	);
	LUT3 #(
		.INIT('h54)
	) name4806 (
		_w1596_,
		_w2086_,
		_w2280_,
		_w5269_
	);
	LUT2 #(
		.INIT('h1)
	) name4807 (
		_w5268_,
		_w5269_,
		_w5270_
	);
	LUT4 #(
		.INIT('h0e00)
	) name4808 (
		_w2276_,
		_w5265_,
		_w5267_,
		_w5270_,
		_w5271_
	);
	LUT4 #(
		.INIT('h00fe)
	) name4809 (
		_w1491_,
		_w1493_,
		_w1496_,
		_w1596_,
		_w5272_
	);
	LUT4 #(
		.INIT('h00d7)
	) name4810 (
		_w2277_,
		_w5263_,
		_w5264_,
		_w5272_,
		_w5273_
	);
	LUT4 #(
		.INIT('h0605)
	) name4811 (
		_w1586_,
		_w1599_,
		_w2042_,
		_w2057_,
		_w5274_
	);
	LUT3 #(
		.INIT('h70)
	) name4812 (
		_w1548_,
		_w1549_,
		_w2042_,
		_w5275_
	);
	LUT4 #(
		.INIT('h1113)
	) name4813 (
		_w2277_,
		_w5272_,
		_w5274_,
		_w5275_,
		_w5276_
	);
	LUT4 #(
		.INIT('hf351)
	) name4814 (
		_w2081_,
		_w2290_,
		_w5273_,
		_w5276_,
		_w5277_
	);
	LUT4 #(
		.INIT('h3111)
	) name4815 (
		_w1489_,
		_w5261_,
		_w5271_,
		_w5277_,
		_w5278_
	);
	LUT2 #(
		.INIT('h4)
	) name4816 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[4]/NET0131 ,
		_w5279_
	);
	LUT4 #(
		.INIT('h0028)
	) name4817 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		_w1476_,
		_w1596_,
		_w5280_
	);
	LUT2 #(
		.INIT('h1)
	) name4818 (
		_w5279_,
		_w5280_,
		_w5281_
	);
	LUT3 #(
		.INIT('h2f)
	) name4819 (
		\P1_state_reg[0]/NET0131 ,
		_w5278_,
		_w5281_,
		_w5282_
	);
	LUT3 #(
		.INIT('h8a)
	) name4820 (
		\P1_reg1_reg[7]/NET0131 ,
		_w3685_,
		_w4079_,
		_w5283_
	);
	LUT4 #(
		.INIT('h7020)
	) name4821 (
		_w537_,
		_w924_,
		_w1183_,
		_w4935_,
		_w5284_
	);
	LUT4 #(
		.INIT('h0001)
	) name4822 (
		_w918_,
		_w1104_,
		_w1106_,
		_w1111_,
		_w5285_
	);
	LUT4 #(
		.INIT('h0001)
	) name4823 (
		_w4940_,
		_w4943_,
		_w4939_,
		_w5285_,
		_w5286_
	);
	LUT4 #(
		.INIT('hecee)
	) name4824 (
		_w4074_,
		_w5283_,
		_w5284_,
		_w5286_,
		_w5287_
	);
	LUT4 #(
		.INIT('h70d0)
	) name4825 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg0_reg[5]/NET0131 ,
		_w1476_,
		_w5288_
	);
	LUT2 #(
		.INIT('h8)
	) name4826 (
		\P2_reg0_reg[5]/NET0131 ,
		_w1487_,
		_w5289_
	);
	LUT4 #(
		.INIT('h08c8)
	) name4827 (
		\P2_reg0_reg[5]/NET0131 ,
		_w2081_,
		_w2272_,
		_w4957_,
		_w5290_
	);
	LUT4 #(
		.INIT('hd11d)
	) name4828 (
		\P2_reg0_reg[5]/NET0131 ,
		_w2272_,
		_w2304_,
		_w4959_,
		_w5291_
	);
	LUT2 #(
		.INIT('h2)
	) name4829 (
		_w2290_,
		_w5291_,
		_w5292_
	);
	LUT4 #(
		.INIT('hd11d)
	) name4830 (
		\P2_reg0_reg[5]/NET0131 ,
		_w2277_,
		_w2304_,
		_w4959_,
		_w5293_
	);
	LUT2 #(
		.INIT('h1)
	) name4831 (
		_w2276_,
		_w5293_,
		_w5294_
	);
	LUT4 #(
		.INIT('hd11d)
	) name4832 (
		\P2_reg0_reg[5]/NET0131 ,
		_w2277_,
		_w4959_,
		_w4965_,
		_w5295_
	);
	LUT2 #(
		.INIT('h4)
	) name4833 (
		_w1593_,
		_w2084_,
		_w5296_
	);
	LUT2 #(
		.INIT('h8)
	) name4834 (
		_w2277_,
		_w5296_,
		_w5297_
	);
	LUT3 #(
		.INIT('ha2)
	) name4835 (
		\P2_reg0_reg[5]/NET0131 ,
		_w2633_,
		_w2634_,
		_w5298_
	);
	LUT2 #(
		.INIT('h1)
	) name4836 (
		_w5297_,
		_w5298_,
		_w5299_
	);
	LUT3 #(
		.INIT('he0)
	) name4837 (
		_w2192_,
		_w5295_,
		_w5299_,
		_w5300_
	);
	LUT4 #(
		.INIT('h0100)
	) name4838 (
		_w5294_,
		_w5292_,
		_w5290_,
		_w5300_,
		_w5301_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name4839 (
		\P1_state_reg[0]/NET0131 ,
		_w1489_,
		_w5289_,
		_w5301_,
		_w5302_
	);
	LUT2 #(
		.INIT('he)
	) name4840 (
		_w5288_,
		_w5302_,
		_w5303_
	);
	LUT4 #(
		.INIT('h70d0)
	) name4841 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg0_reg[6]/NET0131 ,
		_w1476_,
		_w5304_
	);
	LUT2 #(
		.INIT('h8)
	) name4842 (
		\P2_reg0_reg[6]/NET0131 ,
		_w1487_,
		_w5305_
	);
	LUT4 #(
		.INIT('haaa8)
	) name4843 (
		\P2_reg0_reg[6]/NET0131 ,
		_w1491_,
		_w1493_,
		_w1496_,
		_w5306_
	);
	LUT3 #(
		.INIT('h54)
	) name4844 (
		_w2276_,
		_w4993_,
		_w5306_,
		_w5307_
	);
	LUT4 #(
		.INIT('h40b0)
	) name4845 (
		_w2117_,
		_w2120_,
		_w2277_,
		_w4984_,
		_w5308_
	);
	LUT2 #(
		.INIT('h4)
	) name4846 (
		_w1527_,
		_w2084_,
		_w5309_
	);
	LUT2 #(
		.INIT('h8)
	) name4847 (
		_w2277_,
		_w5309_,
		_w5310_
	);
	LUT3 #(
		.INIT('ha2)
	) name4848 (
		\P2_reg0_reg[6]/NET0131 ,
		_w2633_,
		_w2634_,
		_w5311_
	);
	LUT2 #(
		.INIT('h1)
	) name4849 (
		_w5310_,
		_w5311_,
		_w5312_
	);
	LUT4 #(
		.INIT('hab00)
	) name4850 (
		_w2192_,
		_w5306_,
		_w5308_,
		_w5312_,
		_w5313_
	);
	LUT4 #(
		.INIT('h02aa)
	) name4851 (
		\P2_reg0_reg[6]/NET0131 ,
		_w1491_,
		_w1493_,
		_w1496_,
		_w5314_
	);
	LUT3 #(
		.INIT('ha8)
	) name4852 (
		_w2290_,
		_w4995_,
		_w5314_,
		_w5315_
	);
	LUT4 #(
		.INIT('h08c8)
	) name4853 (
		\P2_reg0_reg[6]/NET0131 ,
		_w2081_,
		_w2272_,
		_w4981_,
		_w5316_
	);
	LUT4 #(
		.INIT('h0100)
	) name4854 (
		_w5307_,
		_w5315_,
		_w5316_,
		_w5313_,
		_w5317_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name4855 (
		\P1_state_reg[0]/NET0131 ,
		_w1489_,
		_w5305_,
		_w5317_,
		_w5318_
	);
	LUT2 #(
		.INIT('he)
	) name4856 (
		_w5304_,
		_w5318_,
		_w5319_
	);
	LUT4 #(
		.INIT('h70d0)
	) name4857 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg0_reg[7]/NET0131 ,
		_w1476_,
		_w5320_
	);
	LUT2 #(
		.INIT('h8)
	) name4858 (
		\P2_reg0_reg[7]/NET0131 ,
		_w1487_,
		_w5321_
	);
	LUT4 #(
		.INIT('he020)
	) name4859 (
		\P2_reg0_reg[7]/NET0131 ,
		_w2272_,
		_w2290_,
		_w5003_,
		_w5322_
	);
	LUT4 #(
		.INIT('haaa8)
	) name4860 (
		\P2_reg0_reg[7]/NET0131 ,
		_w1491_,
		_w1493_,
		_w1496_,
		_w5323_
	);
	LUT4 #(
		.INIT('h3202)
	) name4861 (
		\P2_reg0_reg[7]/NET0131 ,
		_w2276_,
		_w2277_,
		_w5003_,
		_w5324_
	);
	LUT4 #(
		.INIT('h111d)
	) name4862 (
		\P2_reg0_reg[7]/NET0131 ,
		_w2272_,
		_w5007_,
		_w5008_,
		_w5325_
	);
	LUT2 #(
		.INIT('h2)
	) name4863 (
		_w2081_,
		_w5325_,
		_w5326_
	);
	LUT4 #(
		.INIT('ha802)
	) name4864 (
		_w2277_,
		_w2351_,
		_w2355_,
		_w5002_,
		_w5327_
	);
	LUT2 #(
		.INIT('h4)
	) name4865 (
		_w1545_,
		_w2084_,
		_w5328_
	);
	LUT2 #(
		.INIT('h8)
	) name4866 (
		_w2277_,
		_w5328_,
		_w5329_
	);
	LUT3 #(
		.INIT('ha2)
	) name4867 (
		\P2_reg0_reg[7]/NET0131 ,
		_w2633_,
		_w2634_,
		_w5330_
	);
	LUT2 #(
		.INIT('h1)
	) name4868 (
		_w5329_,
		_w5330_,
		_w5331_
	);
	LUT4 #(
		.INIT('hab00)
	) name4869 (
		_w2192_,
		_w5323_,
		_w5327_,
		_w5331_,
		_w5332_
	);
	LUT4 #(
		.INIT('h0100)
	) name4870 (
		_w5324_,
		_w5322_,
		_w5326_,
		_w5332_,
		_w5333_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name4871 (
		\P1_state_reg[0]/NET0131 ,
		_w1489_,
		_w5321_,
		_w5333_,
		_w5334_
	);
	LUT2 #(
		.INIT('he)
	) name4872 (
		_w5320_,
		_w5334_,
		_w5335_
	);
	LUT4 #(
		.INIT('h70d0)
	) name4873 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg0_reg[8]/NET0131 ,
		_w1476_,
		_w5336_
	);
	LUT2 #(
		.INIT('h8)
	) name4874 (
		\P2_reg0_reg[8]/NET0131 ,
		_w1487_,
		_w5337_
	);
	LUT4 #(
		.INIT('h35c5)
	) name4875 (
		\P2_reg0_reg[8]/NET0131 ,
		_w2124_,
		_w2277_,
		_w4573_,
		_w5338_
	);
	LUT4 #(
		.INIT('h08c8)
	) name4876 (
		\P2_reg0_reg[8]/NET0131 ,
		_w2081_,
		_w2272_,
		_w4577_,
		_w5339_
	);
	LUT4 #(
		.INIT('hf100)
	) name4877 (
		_w1509_,
		_w1681_,
		_w1683_,
		_w2084_,
		_w5340_
	);
	LUT2 #(
		.INIT('h8)
	) name4878 (
		_w2277_,
		_w5340_,
		_w5341_
	);
	LUT3 #(
		.INIT('ha2)
	) name4879 (
		\P2_reg0_reg[8]/NET0131 ,
		_w2633_,
		_w2634_,
		_w5342_
	);
	LUT2 #(
		.INIT('h1)
	) name4880 (
		_w5341_,
		_w5342_,
		_w5343_
	);
	LUT4 #(
		.INIT('h0e00)
	) name4881 (
		_w2192_,
		_w5338_,
		_w5339_,
		_w5343_,
		_w5344_
	);
	LUT4 #(
		.INIT('h20e0)
	) name4882 (
		\P2_reg0_reg[8]/NET0131 ,
		_w2272_,
		_w2290_,
		_w4574_,
		_w5345_
	);
	LUT4 #(
		.INIT('h0232)
	) name4883 (
		\P2_reg0_reg[8]/NET0131 ,
		_w2276_,
		_w2277_,
		_w4574_,
		_w5346_
	);
	LUT2 #(
		.INIT('h1)
	) name4884 (
		_w5345_,
		_w5346_,
		_w5347_
	);
	LUT4 #(
		.INIT('h3111)
	) name4885 (
		_w1489_,
		_w5337_,
		_w5344_,
		_w5347_,
		_w5348_
	);
	LUT3 #(
		.INIT('hce)
	) name4886 (
		\P1_state_reg[0]/NET0131 ,
		_w5336_,
		_w5348_,
		_w5349_
	);
	LUT4 #(
		.INIT('h0001)
	) name4887 (
		_w881_,
		_w1104_,
		_w1106_,
		_w1111_,
		_w5350_
	);
	LUT4 #(
		.INIT('h0001)
	) name4888 (
		_w4924_,
		_w4922_,
		_w4925_,
		_w5350_,
		_w5351_
	);
	LUT2 #(
		.INIT('h4)
	) name4889 (
		\P1_reg3_reg[3]/NET0131 ,
		_w1143_,
		_w5352_
	);
	LUT4 #(
		.INIT('h5455)
	) name4890 (
		\P1_reg2_reg[3]/NET0131 ,
		_w528_,
		_w530_,
		_w533_,
		_w5353_
	);
	LUT2 #(
		.INIT('h2)
	) name4891 (
		_w1183_,
		_w5353_,
		_w5354_
	);
	LUT4 #(
		.INIT('h5700)
	) name4892 (
		_w534_,
		_w4919_,
		_w4920_,
		_w5354_,
		_w5355_
	);
	LUT4 #(
		.INIT('h0031)
	) name4893 (
		_w534_,
		_w5352_,
		_w5351_,
		_w5355_,
		_w5356_
	);
	LUT3 #(
		.INIT('hb0)
	) name4894 (
		_w534_,
		_w1286_,
		_w3443_,
		_w5357_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name4895 (
		\P1_reg2_reg[3]/NET0131 ,
		_w2411_,
		_w2412_,
		_w5357_,
		_w5358_
	);
	LUT3 #(
		.INIT('hf2)
	) name4896 (
		_w3443_,
		_w5356_,
		_w5358_,
		_w5359_
	);
	LUT3 #(
		.INIT('h8a)
	) name4897 (
		\P1_reg2_reg[5]/NET0131 ,
		_w2951_,
		_w3938_,
		_w5360_
	);
	LUT2 #(
		.INIT('h8)
	) name4898 (
		_w931_,
		_w1143_,
		_w5361_
	);
	LUT4 #(
		.INIT('h0075)
	) name4899 (
		_w534_,
		_w5166_,
		_w5168_,
		_w5361_,
		_w5362_
	);
	LUT3 #(
		.INIT('hce)
	) name4900 (
		_w3443_,
		_w5360_,
		_w5362_,
		_w5363_
	);
	LUT2 #(
		.INIT('h2)
	) name4901 (
		\P1_reg2_reg[6]/NET0131 ,
		_w511_,
		_w5364_
	);
	LUT2 #(
		.INIT('h8)
	) name4902 (
		\P1_reg2_reg[6]/NET0131 ,
		_w524_,
		_w5365_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name4903 (
		\P1_reg2_reg[6]/NET0131 ,
		_w528_,
		_w530_,
		_w533_,
		_w5366_
	);
	LUT4 #(
		.INIT('hddd1)
	) name4904 (
		\P1_reg2_reg[6]/NET0131 ,
		_w534_,
		_w5243_,
		_w5244_,
		_w5367_
	);
	LUT4 #(
		.INIT('h8828)
	) name4905 (
		_w534_,
		_w1448_,
		_w2225_,
		_w3049_,
		_w5368_
	);
	LUT3 #(
		.INIT('ha8)
	) name4906 (
		_w1114_,
		_w5366_,
		_w5368_,
		_w5369_
	);
	LUT4 #(
		.INIT('h0a82)
	) name4907 (
		_w534_,
		_w1366_,
		_w1448_,
		_w3073_,
		_w5370_
	);
	LUT4 #(
		.INIT('he020)
	) name4908 (
		\P1_reg2_reg[6]/NET0131 ,
		_w534_,
		_w1136_,
		_w5249_,
		_w5371_
	);
	LUT4 #(
		.INIT('haa20)
	) name4909 (
		\P1_reg2_reg[6]/NET0131 ,
		_w534_,
		_w1138_,
		_w1141_,
		_w5372_
	);
	LUT4 #(
		.INIT('h0001)
	) name4910 (
		_w929_,
		_w1104_,
		_w1106_,
		_w1111_,
		_w5373_
	);
	LUT4 #(
		.INIT('h153f)
	) name4911 (
		_w534_,
		_w922_,
		_w1143_,
		_w5373_,
		_w5374_
	);
	LUT2 #(
		.INIT('h4)
	) name4912 (
		_w5372_,
		_w5374_,
		_w5375_
	);
	LUT2 #(
		.INIT('h4)
	) name4913 (
		_w5371_,
		_w5375_,
		_w5376_
	);
	LUT4 #(
		.INIT('h5700)
	) name4914 (
		_w1286_,
		_w5366_,
		_w5370_,
		_w5376_,
		_w5377_
	);
	LUT4 #(
		.INIT('h3100)
	) name4915 (
		_w1183_,
		_w5369_,
		_w5367_,
		_w5377_,
		_w5378_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name4916 (
		\P1_state_reg[0]/NET0131 ,
		_w526_,
		_w5365_,
		_w5378_,
		_w5379_
	);
	LUT2 #(
		.INIT('he)
	) name4917 (
		_w5364_,
		_w5379_,
		_w5380_
	);
	LUT4 #(
		.INIT('hf200)
	) name4918 (
		_w534_,
		_w1141_,
		_w1143_,
		_w3443_,
		_w5381_
	);
	LUT2 #(
		.INIT('h2)
	) name4919 (
		\P1_reg2_reg[7]/NET0131 ,
		_w5381_,
		_w5382_
	);
	LUT2 #(
		.INIT('h8)
	) name4920 (
		_w910_,
		_w1143_,
		_w5383_
	);
	LUT4 #(
		.INIT('h0075)
	) name4921 (
		_w534_,
		_w5284_,
		_w5286_,
		_w5383_,
		_w5384_
	);
	LUT3 #(
		.INIT('hce)
	) name4922 (
		_w3443_,
		_w5382_,
		_w5384_,
		_w5385_
	);
	LUT4 #(
		.INIT('h70d0)
	) name4923 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg1_reg[5]/NET0131 ,
		_w1476_,
		_w5386_
	);
	LUT2 #(
		.INIT('h8)
	) name4924 (
		\P2_reg1_reg[5]/NET0131 ,
		_w1487_,
		_w5387_
	);
	LUT4 #(
		.INIT('h20e0)
	) name4925 (
		\P2_reg1_reg[5]/NET0131 ,
		_w1497_,
		_w2081_,
		_w4957_,
		_w5388_
	);
	LUT4 #(
		.INIT('hd11d)
	) name4926 (
		\P2_reg1_reg[5]/NET0131 ,
		_w2039_,
		_w2304_,
		_w4959_,
		_w5389_
	);
	LUT2 #(
		.INIT('h2)
	) name4927 (
		_w2038_,
		_w5389_,
		_w5390_
	);
	LUT4 #(
		.INIT('hd11d)
	) name4928 (
		\P2_reg1_reg[5]/NET0131 ,
		_w2039_,
		_w4959_,
		_w4965_,
		_w5391_
	);
	LUT2 #(
		.INIT('h2)
	) name4929 (
		_w2193_,
		_w5391_,
		_w5392_
	);
	LUT4 #(
		.INIT('hd11d)
	) name4930 (
		\P2_reg1_reg[5]/NET0131 ,
		_w1497_,
		_w4959_,
		_w4965_,
		_w5393_
	);
	LUT2 #(
		.INIT('h8)
	) name4931 (
		_w2039_,
		_w5296_,
		_w5394_
	);
	LUT3 #(
		.INIT('ha2)
	) name4932 (
		\P2_reg1_reg[5]/NET0131 ,
		_w2633_,
		_w2660_,
		_w5395_
	);
	LUT2 #(
		.INIT('h1)
	) name4933 (
		_w5394_,
		_w5395_,
		_w5396_
	);
	LUT3 #(
		.INIT('hd0)
	) name4934 (
		_w2188_,
		_w5393_,
		_w5396_,
		_w5397_
	);
	LUT4 #(
		.INIT('h0100)
	) name4935 (
		_w5388_,
		_w5390_,
		_w5392_,
		_w5397_,
		_w5398_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name4936 (
		\P1_state_reg[0]/NET0131 ,
		_w1489_,
		_w5387_,
		_w5398_,
		_w5399_
	);
	LUT2 #(
		.INIT('he)
	) name4937 (
		_w5386_,
		_w5399_,
		_w5400_
	);
	LUT4 #(
		.INIT('h70d0)
	) name4938 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg1_reg[6]/NET0131 ,
		_w1476_,
		_w5401_
	);
	LUT2 #(
		.INIT('h8)
	) name4939 (
		\P2_reg1_reg[6]/NET0131 ,
		_w1487_,
		_w5402_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name4940 (
		\P2_reg1_reg[6]/NET0131 ,
		_w1491_,
		_w1493_,
		_w1496_,
		_w5403_
	);
	LUT4 #(
		.INIT('h208a)
	) name4941 (
		_w1497_,
		_w2117_,
		_w2120_,
		_w4984_,
		_w5404_
	);
	LUT3 #(
		.INIT('ha8)
	) name4942 (
		_w2188_,
		_w5403_,
		_w5404_,
		_w5405_
	);
	LUT4 #(
		.INIT('haa02)
	) name4943 (
		\P2_reg1_reg[6]/NET0131 ,
		_w1491_,
		_w1493_,
		_w1496_,
		_w5406_
	);
	LUT4 #(
		.INIT('h208a)
	) name4944 (
		_w2039_,
		_w2117_,
		_w2120_,
		_w4984_,
		_w5407_
	);
	LUT2 #(
		.INIT('h8)
	) name4945 (
		_w2039_,
		_w5309_,
		_w5408_
	);
	LUT3 #(
		.INIT('ha2)
	) name4946 (
		\P2_reg1_reg[6]/NET0131 ,
		_w2633_,
		_w2660_,
		_w5409_
	);
	LUT2 #(
		.INIT('h1)
	) name4947 (
		_w5408_,
		_w5409_,
		_w5410_
	);
	LUT4 #(
		.INIT('h5700)
	) name4948 (
		_w2193_,
		_w5406_,
		_w5407_,
		_w5410_,
		_w5411_
	);
	LUT4 #(
		.INIT('he010)
	) name4949 (
		_w1608_,
		_w1611_,
		_w2039_,
		_w4984_,
		_w5412_
	);
	LUT3 #(
		.INIT('ha8)
	) name4950 (
		_w2038_,
		_w5406_,
		_w5412_,
		_w5413_
	);
	LUT4 #(
		.INIT('h20e0)
	) name4951 (
		\P2_reg1_reg[6]/NET0131 ,
		_w1497_,
		_w2081_,
		_w4981_,
		_w5414_
	);
	LUT4 #(
		.INIT('h0100)
	) name4952 (
		_w5413_,
		_w5414_,
		_w5405_,
		_w5411_,
		_w5415_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name4953 (
		\P1_state_reg[0]/NET0131 ,
		_w1489_,
		_w5402_,
		_w5415_,
		_w5416_
	);
	LUT2 #(
		.INIT('he)
	) name4954 (
		_w5401_,
		_w5416_,
		_w5417_
	);
	LUT4 #(
		.INIT('h70d0)
	) name4955 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg1_reg[7]/NET0131 ,
		_w1476_,
		_w5418_
	);
	LUT2 #(
		.INIT('h8)
	) name4956 (
		\P2_reg1_reg[7]/NET0131 ,
		_w1487_,
		_w5419_
	);
	LUT4 #(
		.INIT('haa02)
	) name4957 (
		\P2_reg1_reg[7]/NET0131 ,
		_w1491_,
		_w1493_,
		_w1496_,
		_w5420_
	);
	LUT4 #(
		.INIT('hc808)
	) name4958 (
		\P2_reg1_reg[7]/NET0131 ,
		_w2038_,
		_w2039_,
		_w5003_,
		_w5421_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name4959 (
		\P2_reg1_reg[7]/NET0131 ,
		_w1491_,
		_w1493_,
		_w1496_,
		_w5422_
	);
	LUT4 #(
		.INIT('h111d)
	) name4960 (
		\P2_reg1_reg[7]/NET0131 ,
		_w1497_,
		_w5007_,
		_w5008_,
		_w5423_
	);
	LUT2 #(
		.INIT('h4)
	) name4961 (
		_w1545_,
		_w2963_,
		_w5424_
	);
	LUT3 #(
		.INIT('ha2)
	) name4962 (
		\P2_reg1_reg[7]/NET0131 ,
		_w2633_,
		_w2660_,
		_w5425_
	);
	LUT2 #(
		.INIT('h1)
	) name4963 (
		_w5424_,
		_w5425_,
		_w5426_
	);
	LUT3 #(
		.INIT('hd0)
	) name4964 (
		_w2081_,
		_w5423_,
		_w5426_,
		_w5427_
	);
	LUT4 #(
		.INIT('ha802)
	) name4965 (
		_w1497_,
		_w2351_,
		_w2355_,
		_w5002_,
		_w5428_
	);
	LUT3 #(
		.INIT('ha8)
	) name4966 (
		_w2188_,
		_w5422_,
		_w5428_,
		_w5429_
	);
	LUT4 #(
		.INIT('ha802)
	) name4967 (
		_w2039_,
		_w2351_,
		_w2355_,
		_w5002_,
		_w5430_
	);
	LUT3 #(
		.INIT('ha8)
	) name4968 (
		_w2193_,
		_w5420_,
		_w5430_,
		_w5431_
	);
	LUT4 #(
		.INIT('h0100)
	) name4969 (
		_w5429_,
		_w5421_,
		_w5431_,
		_w5427_,
		_w5432_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name4970 (
		\P1_state_reg[0]/NET0131 ,
		_w1489_,
		_w5419_,
		_w5432_,
		_w5433_
	);
	LUT2 #(
		.INIT('he)
	) name4971 (
		_w5418_,
		_w5433_,
		_w5434_
	);
	LUT4 #(
		.INIT('h70d0)
	) name4972 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg1_reg[8]/NET0131 ,
		_w1476_,
		_w5435_
	);
	LUT2 #(
		.INIT('h8)
	) name4973 (
		\P2_reg1_reg[8]/NET0131 ,
		_w1487_,
		_w5436_
	);
	LUT4 #(
		.INIT('h1dd1)
	) name4974 (
		\P2_reg1_reg[8]/NET0131 ,
		_w1497_,
		_w2124_,
		_w4573_,
		_w5437_
	);
	LUT4 #(
		.INIT('h20e0)
	) name4975 (
		\P2_reg1_reg[8]/NET0131 ,
		_w1497_,
		_w2081_,
		_w4577_,
		_w5438_
	);
	LUT2 #(
		.INIT('h8)
	) name4976 (
		_w2039_,
		_w5340_,
		_w5439_
	);
	LUT3 #(
		.INIT('ha2)
	) name4977 (
		\P2_reg1_reg[8]/NET0131 ,
		_w2633_,
		_w2660_,
		_w5440_
	);
	LUT2 #(
		.INIT('h1)
	) name4978 (
		_w5439_,
		_w5440_,
		_w5441_
	);
	LUT4 #(
		.INIT('h0d00)
	) name4979 (
		_w2188_,
		_w5437_,
		_w5438_,
		_w5441_,
		_w5442_
	);
	LUT4 #(
		.INIT('h1dd1)
	) name4980 (
		\P2_reg1_reg[8]/NET0131 ,
		_w2039_,
		_w2124_,
		_w4573_,
		_w5443_
	);
	LUT4 #(
		.INIT('h08c8)
	) name4981 (
		\P2_reg1_reg[8]/NET0131 ,
		_w2038_,
		_w2039_,
		_w4574_,
		_w5444_
	);
	LUT3 #(
		.INIT('h0d)
	) name4982 (
		_w2193_,
		_w5443_,
		_w5444_,
		_w5445_
	);
	LUT4 #(
		.INIT('h3111)
	) name4983 (
		_w1489_,
		_w5436_,
		_w5442_,
		_w5445_,
		_w5446_
	);
	LUT3 #(
		.INIT('hce)
	) name4984 (
		\P1_state_reg[0]/NET0131 ,
		_w5435_,
		_w5446_,
		_w5447_
	);
	LUT4 #(
		.INIT('h70d0)
	) name4985 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg2_reg[5]/NET0131 ,
		_w1476_,
		_w5448_
	);
	LUT2 #(
		.INIT('h8)
	) name4986 (
		\P2_reg2_reg[5]/NET0131 ,
		_w1487_,
		_w5449_
	);
	LUT4 #(
		.INIT('h20e0)
	) name4987 (
		\P2_reg2_reg[5]/NET0131 ,
		_w2039_,
		_w2081_,
		_w4957_,
		_w5450_
	);
	LUT4 #(
		.INIT('hd11d)
	) name4988 (
		\P2_reg2_reg[5]/NET0131 ,
		_w1497_,
		_w2304_,
		_w4959_,
		_w5451_
	);
	LUT2 #(
		.INIT('h2)
	) name4989 (
		_w2038_,
		_w5451_,
		_w5452_
	);
	LUT4 #(
		.INIT('hd11d)
	) name4990 (
		\P2_reg2_reg[5]/NET0131 ,
		_w2039_,
		_w4959_,
		_w4965_,
		_w5453_
	);
	LUT2 #(
		.INIT('h2)
	) name4991 (
		_w2188_,
		_w5453_,
		_w5454_
	);
	LUT4 #(
		.INIT('hd11d)
	) name4992 (
		\P2_reg2_reg[5]/NET0131 ,
		_w1497_,
		_w4959_,
		_w4965_,
		_w5455_
	);
	LUT3 #(
		.INIT('ha8)
	) name4993 (
		\P2_reg2_reg[5]/NET0131 ,
		_w2086_,
		_w2087_,
		_w5456_
	);
	LUT2 #(
		.INIT('h4)
	) name4994 (
		_w1584_,
		_w2088_,
		_w5457_
	);
	LUT3 #(
		.INIT('h07)
	) name4995 (
		_w1497_,
		_w5296_,
		_w5457_,
		_w5458_
	);
	LUT2 #(
		.INIT('h4)
	) name4996 (
		_w5456_,
		_w5458_,
		_w5459_
	);
	LUT3 #(
		.INIT('hd0)
	) name4997 (
		_w2193_,
		_w5455_,
		_w5459_,
		_w5460_
	);
	LUT4 #(
		.INIT('h0100)
	) name4998 (
		_w5450_,
		_w5452_,
		_w5454_,
		_w5460_,
		_w5461_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name4999 (
		\P1_state_reg[0]/NET0131 ,
		_w1489_,
		_w5449_,
		_w5461_,
		_w5462_
	);
	LUT2 #(
		.INIT('he)
	) name5000 (
		_w5448_,
		_w5462_,
		_w5463_
	);
	LUT4 #(
		.INIT('h70d0)
	) name5001 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg2_reg[6]/NET0131 ,
		_w1476_,
		_w5464_
	);
	LUT2 #(
		.INIT('h8)
	) name5002 (
		\P2_reg2_reg[6]/NET0131 ,
		_w1487_,
		_w5465_
	);
	LUT4 #(
		.INIT('haa02)
	) name5003 (
		\P2_reg2_reg[6]/NET0131 ,
		_w1491_,
		_w1493_,
		_w1496_,
		_w5466_
	);
	LUT3 #(
		.INIT('ha8)
	) name5004 (
		_w2188_,
		_w5407_,
		_w5466_,
		_w5467_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name5005 (
		\P2_reg2_reg[6]/NET0131 ,
		_w1491_,
		_w1493_,
		_w1496_,
		_w5468_
	);
	LUT3 #(
		.INIT('ha8)
	) name5006 (
		\P2_reg2_reg[6]/NET0131 ,
		_w2086_,
		_w2087_,
		_w5469_
	);
	LUT2 #(
		.INIT('h4)
	) name5007 (
		_w1500_,
		_w2088_,
		_w5470_
	);
	LUT3 #(
		.INIT('h07)
	) name5008 (
		_w1497_,
		_w5309_,
		_w5470_,
		_w5471_
	);
	LUT2 #(
		.INIT('h4)
	) name5009 (
		_w5469_,
		_w5471_,
		_w5472_
	);
	LUT4 #(
		.INIT('h5700)
	) name5010 (
		_w2193_,
		_w5404_,
		_w5468_,
		_w5472_,
		_w5473_
	);
	LUT4 #(
		.INIT('ha802)
	) name5011 (
		_w1497_,
		_w1608_,
		_w1611_,
		_w4984_,
		_w5474_
	);
	LUT3 #(
		.INIT('ha8)
	) name5012 (
		_w2038_,
		_w5468_,
		_w5474_,
		_w5475_
	);
	LUT4 #(
		.INIT('h20e0)
	) name5013 (
		\P2_reg2_reg[6]/NET0131 ,
		_w2039_,
		_w2081_,
		_w4981_,
		_w5476_
	);
	LUT4 #(
		.INIT('h0100)
	) name5014 (
		_w5475_,
		_w5476_,
		_w5467_,
		_w5473_,
		_w5477_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name5015 (
		\P1_state_reg[0]/NET0131 ,
		_w1489_,
		_w5465_,
		_w5477_,
		_w5478_
	);
	LUT2 #(
		.INIT('he)
	) name5016 (
		_w5464_,
		_w5478_,
		_w5479_
	);
	LUT4 #(
		.INIT('h70d0)
	) name5017 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg2_reg[7]/NET0131 ,
		_w1476_,
		_w5480_
	);
	LUT2 #(
		.INIT('h8)
	) name5018 (
		\P2_reg2_reg[7]/NET0131 ,
		_w1487_,
		_w5481_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name5019 (
		\P2_reg2_reg[7]/NET0131 ,
		_w1491_,
		_w1493_,
		_w1496_,
		_w5482_
	);
	LUT4 #(
		.INIT('he020)
	) name5020 (
		\P2_reg2_reg[7]/NET0131 ,
		_w1497_,
		_w2038_,
		_w5003_,
		_w5483_
	);
	LUT4 #(
		.INIT('haa02)
	) name5021 (
		\P2_reg2_reg[7]/NET0131 ,
		_w1491_,
		_w1493_,
		_w1496_,
		_w5484_
	);
	LUT4 #(
		.INIT('h111d)
	) name5022 (
		\P2_reg2_reg[7]/NET0131 ,
		_w2039_,
		_w5007_,
		_w5008_,
		_w5485_
	);
	LUT3 #(
		.INIT('ha8)
	) name5023 (
		\P2_reg2_reg[7]/NET0131 ,
		_w2086_,
		_w2087_,
		_w5486_
	);
	LUT2 #(
		.INIT('h4)
	) name5024 (
		_w1530_,
		_w2088_,
		_w5487_
	);
	LUT3 #(
		.INIT('h07)
	) name5025 (
		_w1497_,
		_w5328_,
		_w5487_,
		_w5488_
	);
	LUT2 #(
		.INIT('h4)
	) name5026 (
		_w5486_,
		_w5488_,
		_w5489_
	);
	LUT3 #(
		.INIT('hd0)
	) name5027 (
		_w2081_,
		_w5485_,
		_w5489_,
		_w5490_
	);
	LUT3 #(
		.INIT('ha8)
	) name5028 (
		_w2188_,
		_w5430_,
		_w5484_,
		_w5491_
	);
	LUT3 #(
		.INIT('ha8)
	) name5029 (
		_w2193_,
		_w5428_,
		_w5482_,
		_w5492_
	);
	LUT4 #(
		.INIT('h0100)
	) name5030 (
		_w5491_,
		_w5483_,
		_w5492_,
		_w5490_,
		_w5493_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name5031 (
		\P1_state_reg[0]/NET0131 ,
		_w1489_,
		_w5481_,
		_w5493_,
		_w5494_
	);
	LUT2 #(
		.INIT('he)
	) name5032 (
		_w5480_,
		_w5494_,
		_w5495_
	);
	LUT4 #(
		.INIT('h70d0)
	) name5033 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg2_reg[8]/NET0131 ,
		_w1476_,
		_w5496_
	);
	LUT2 #(
		.INIT('h8)
	) name5034 (
		\P2_reg2_reg[8]/NET0131 ,
		_w1487_,
		_w5497_
	);
	LUT4 #(
		.INIT('h1dd1)
	) name5035 (
		\P2_reg2_reg[8]/NET0131 ,
		_w1497_,
		_w2124_,
		_w4573_,
		_w5498_
	);
	LUT4 #(
		.INIT('h20e0)
	) name5036 (
		\P2_reg2_reg[8]/NET0131 ,
		_w2039_,
		_w2081_,
		_w4577_,
		_w5499_
	);
	LUT3 #(
		.INIT('ha8)
	) name5037 (
		\P2_reg2_reg[8]/NET0131 ,
		_w2086_,
		_w2087_,
		_w5500_
	);
	LUT2 #(
		.INIT('h4)
	) name5038 (
		_w1674_,
		_w2088_,
		_w5501_
	);
	LUT3 #(
		.INIT('h07)
	) name5039 (
		_w1497_,
		_w5340_,
		_w5501_,
		_w5502_
	);
	LUT2 #(
		.INIT('h4)
	) name5040 (
		_w5500_,
		_w5502_,
		_w5503_
	);
	LUT4 #(
		.INIT('h3100)
	) name5041 (
		_w2193_,
		_w5499_,
		_w5498_,
		_w5503_,
		_w5504_
	);
	LUT4 #(
		.INIT('h1dd1)
	) name5042 (
		\P2_reg2_reg[8]/NET0131 ,
		_w2039_,
		_w2124_,
		_w4573_,
		_w5505_
	);
	LUT4 #(
		.INIT('h20e0)
	) name5043 (
		\P2_reg2_reg[8]/NET0131 ,
		_w1497_,
		_w2038_,
		_w4574_,
		_w5506_
	);
	LUT3 #(
		.INIT('h0d)
	) name5044 (
		_w2188_,
		_w5505_,
		_w5506_,
		_w5507_
	);
	LUT4 #(
		.INIT('h3111)
	) name5045 (
		_w1489_,
		_w5497_,
		_w5504_,
		_w5507_,
		_w5508_
	);
	LUT3 #(
		.INIT('hce)
	) name5046 (
		\P1_state_reg[0]/NET0131 ,
		_w5496_,
		_w5508_,
		_w5509_
	);
	LUT2 #(
		.INIT('h2)
	) name5047 (
		\P1_reg0_reg[3]/NET0131 ,
		_w511_,
		_w5510_
	);
	LUT2 #(
		.INIT('h8)
	) name5048 (
		\P1_reg0_reg[3]/NET0131 ,
		_w524_,
		_w5511_
	);
	LUT4 #(
		.INIT('hddd1)
	) name5049 (
		\P1_reg0_reg[3]/NET0131 ,
		_w2688_,
		_w4919_,
		_w4920_,
		_w5512_
	);
	LUT4 #(
		.INIT('haaa8)
	) name5050 (
		_w2688_,
		_w4922_,
		_w4925_,
		_w5350_,
		_w5513_
	);
	LUT4 #(
		.INIT('hc808)
	) name5051 (
		\P1_reg0_reg[3]/NET0131 ,
		_w1136_,
		_w2688_,
		_w4923_,
		_w5514_
	);
	LUT4 #(
		.INIT('h005d)
	) name5052 (
		\P1_reg0_reg[3]/NET0131 ,
		_w2692_,
		_w3966_,
		_w5514_,
		_w5515_
	);
	LUT4 #(
		.INIT('h0d00)
	) name5053 (
		_w1183_,
		_w5512_,
		_w5513_,
		_w5515_,
		_w5516_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name5054 (
		\P1_state_reg[0]/NET0131 ,
		_w526_,
		_w5511_,
		_w5516_,
		_w5517_
	);
	LUT2 #(
		.INIT('he)
	) name5055 (
		_w5510_,
		_w5517_,
		_w5518_
	);
	LUT3 #(
		.INIT('hd0)
	) name5056 (
		_w1140_,
		_w2688_,
		_w3443_,
		_w5519_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name5057 (
		\P1_reg0_reg[7]/NET0131 ,
		_w2692_,
		_w3966_,
		_w5519_,
		_w5520_
	);
	LUT4 #(
		.INIT('hff8a)
	) name5058 (
		_w3651_,
		_w5284_,
		_w5286_,
		_w5520_,
		_w5521_
	);
	LUT2 #(
		.INIT('h2)
	) name5059 (
		\P1_reg1_reg[3]/NET0131 ,
		_w511_,
		_w5522_
	);
	LUT4 #(
		.INIT('h5100)
	) name5060 (
		_w523_,
		_w1183_,
		_w2421_,
		_w2425_,
		_w5523_
	);
	LUT4 #(
		.INIT('h5090)
	) name5061 (
		\P1_IR_reg[23]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		\P1_reg1_reg[3]/NET0131 ,
		_w509_,
		_w5524_
	);
	LUT3 #(
		.INIT('hb0)
	) name5062 (
		_w4078_,
		_w5523_,
		_w5524_,
		_w5525_
	);
	LUT4 #(
		.INIT('h0075)
	) name5063 (
		_w4073_,
		_w4921_,
		_w5351_,
		_w5525_,
		_w5526_
	);
	LUT3 #(
		.INIT('hce)
	) name5064 (
		\P1_state_reg[0]/NET0131 ,
		_w5522_,
		_w5526_,
		_w5527_
	);
	LUT4 #(
		.INIT('h5554)
	) name5065 (
		\P2_reg3_reg[3]/NET0131 ,
		_w1491_,
		_w1493_,
		_w1496_,
		_w5528_
	);
	LUT3 #(
		.INIT('h70)
	) name5066 (
		_w1557_,
		_w1558_,
		_w2042_,
		_w5529_
	);
	LUT4 #(
		.INIT('h00de)
	) name5067 (
		_w1599_,
		_w2042_,
		_w2057_,
		_w5529_,
		_w5530_
	);
	LUT4 #(
		.INIT('h04c4)
	) name5068 (
		\P2_reg3_reg[3]/NET0131 ,
		_w2081_,
		_w2277_,
		_w5530_,
		_w5531_
	);
	LUT4 #(
		.INIT('h0155)
	) name5069 (
		\P2_reg3_reg[3]/NET0131 ,
		_w1491_,
		_w1493_,
		_w1496_,
		_w5532_
	);
	LUT3 #(
		.INIT('h78)
	) name5070 (
		_w1548_,
		_w1549_,
		_w1555_,
		_w5533_
	);
	LUT4 #(
		.INIT('he010)
	) name5071 (
		_w1565_,
		_w1582_,
		_w2272_,
		_w5533_,
		_w5534_
	);
	LUT3 #(
		.INIT('h54)
	) name5072 (
		_w2276_,
		_w5532_,
		_w5534_,
		_w5535_
	);
	LUT4 #(
		.INIT('he010)
	) name5073 (
		_w1565_,
		_w1582_,
		_w2277_,
		_w5533_,
		_w5536_
	);
	LUT3 #(
		.INIT('ha8)
	) name5074 (
		_w2290_,
		_w5528_,
		_w5536_,
		_w5537_
	);
	LUT4 #(
		.INIT('h04c8)
	) name5075 (
		_w2110_,
		_w2272_,
		_w2353_,
		_w5533_,
		_w5538_
	);
	LUT3 #(
		.INIT('h04)
	) name5076 (
		_w1555_,
		_w2083_,
		_w2282_,
		_w5539_
	);
	LUT3 #(
		.INIT('h54)
	) name5077 (
		\P2_reg3_reg[3]/NET0131 ,
		_w2086_,
		_w2280_,
		_w5540_
	);
	LUT2 #(
		.INIT('h1)
	) name5078 (
		_w5539_,
		_w5540_,
		_w5541_
	);
	LUT4 #(
		.INIT('hab00)
	) name5079 (
		_w2192_,
		_w5532_,
		_w5538_,
		_w5541_,
		_w5542_
	);
	LUT4 #(
		.INIT('h0100)
	) name5080 (
		_w5531_,
		_w5537_,
		_w5535_,
		_w5542_,
		_w5543_
	);
	LUT2 #(
		.INIT('h4)
	) name5081 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[3]/NET0131 ,
		_w5544_
	);
	LUT3 #(
		.INIT('hb9)
	) name5082 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[3]/NET0131 ,
		_w1489_,
		_w5545_
	);
	LUT3 #(
		.INIT('h2f)
	) name5083 (
		_w4166_,
		_w5543_,
		_w5545_,
		_w5546_
	);
	LUT2 #(
		.INIT('h2)
	) name5084 (
		\P1_reg1_reg[6]/NET0131 ,
		_w511_,
		_w5547_
	);
	LUT2 #(
		.INIT('h8)
	) name5085 (
		\P1_reg1_reg[6]/NET0131 ,
		_w524_,
		_w5548_
	);
	LUT4 #(
		.INIT('haa02)
	) name5086 (
		\P1_reg1_reg[6]/NET0131 ,
		_w528_,
		_w530_,
		_w533_,
		_w5549_
	);
	LUT4 #(
		.INIT('hddd1)
	) name5087 (
		\P1_reg1_reg[6]/NET0131 ,
		_w2421_,
		_w5243_,
		_w5244_,
		_w5550_
	);
	LUT4 #(
		.INIT('h3090)
	) name5088 (
		_w1366_,
		_w1448_,
		_w2421_,
		_w3073_,
		_w5551_
	);
	LUT3 #(
		.INIT('ha8)
	) name5089 (
		_w1286_,
		_w5549_,
		_w5551_,
		_w5552_
	);
	LUT4 #(
		.INIT('ha060)
	) name5090 (
		_w1448_,
		_w2225_,
		_w2421_,
		_w3049_,
		_w5553_
	);
	LUT4 #(
		.INIT('hc808)
	) name5091 (
		\P1_reg1_reg[6]/NET0131 ,
		_w1136_,
		_w2421_,
		_w5249_,
		_w5554_
	);
	LUT2 #(
		.INIT('h8)
	) name5092 (
		_w2421_,
		_w5373_,
		_w5555_
	);
	LUT4 #(
		.INIT('h08aa)
	) name5093 (
		\P1_reg1_reg[6]/NET0131 ,
		_w1138_,
		_w2421_,
		_w2425_,
		_w5556_
	);
	LUT2 #(
		.INIT('h1)
	) name5094 (
		_w5555_,
		_w5556_,
		_w5557_
	);
	LUT2 #(
		.INIT('h4)
	) name5095 (
		_w5554_,
		_w5557_,
		_w5558_
	);
	LUT4 #(
		.INIT('h5700)
	) name5096 (
		_w1114_,
		_w5549_,
		_w5553_,
		_w5558_,
		_w5559_
	);
	LUT4 #(
		.INIT('h3100)
	) name5097 (
		_w1183_,
		_w5552_,
		_w5550_,
		_w5559_,
		_w5560_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name5098 (
		\P1_state_reg[0]/NET0131 ,
		_w526_,
		_w5548_,
		_w5560_,
		_w5561_
	);
	LUT2 #(
		.INIT('he)
	) name5099 (
		_w5547_,
		_w5561_,
		_w5562_
	);
	LUT2 #(
		.INIT('h2)
	) name5100 (
		\P1_reg0_reg[6]/NET0131 ,
		_w511_,
		_w5563_
	);
	LUT2 #(
		.INIT('h8)
	) name5101 (
		\P1_reg0_reg[6]/NET0131 ,
		_w524_,
		_w5564_
	);
	LUT4 #(
		.INIT('haaa8)
	) name5102 (
		\P1_reg0_reg[6]/NET0131 ,
		_w528_,
		_w530_,
		_w533_,
		_w5565_
	);
	LUT4 #(
		.INIT('hddd1)
	) name5103 (
		\P1_reg0_reg[6]/NET0131 ,
		_w2688_,
		_w5243_,
		_w5244_,
		_w5566_
	);
	LUT4 #(
		.INIT('h3090)
	) name5104 (
		_w1366_,
		_w1448_,
		_w2688_,
		_w3073_,
		_w5567_
	);
	LUT3 #(
		.INIT('ha8)
	) name5105 (
		_w1286_,
		_w5565_,
		_w5567_,
		_w5568_
	);
	LUT4 #(
		.INIT('ha060)
	) name5106 (
		_w1448_,
		_w2225_,
		_w2688_,
		_w3049_,
		_w5569_
	);
	LUT4 #(
		.INIT('hc808)
	) name5107 (
		\P1_reg0_reg[6]/NET0131 ,
		_w1136_,
		_w2688_,
		_w5249_,
		_w5570_
	);
	LUT2 #(
		.INIT('h8)
	) name5108 (
		_w2688_,
		_w5373_,
		_w5571_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name5109 (
		\P1_reg0_reg[6]/NET0131 ,
		_w1138_,
		_w2425_,
		_w2688_,
		_w5572_
	);
	LUT2 #(
		.INIT('h1)
	) name5110 (
		_w5571_,
		_w5572_,
		_w5573_
	);
	LUT2 #(
		.INIT('h4)
	) name5111 (
		_w5570_,
		_w5573_,
		_w5574_
	);
	LUT4 #(
		.INIT('h5700)
	) name5112 (
		_w1114_,
		_w5565_,
		_w5569_,
		_w5574_,
		_w5575_
	);
	LUT4 #(
		.INIT('h3100)
	) name5113 (
		_w1183_,
		_w5568_,
		_w5566_,
		_w5575_,
		_w5576_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name5114 (
		\P1_state_reg[0]/NET0131 ,
		_w526_,
		_w5564_,
		_w5576_,
		_w5577_
	);
	LUT2 #(
		.INIT('he)
	) name5115 (
		_w5563_,
		_w5577_,
		_w5578_
	);
	LUT2 #(
		.INIT('h4)
	) name5116 (
		_w853_,
		_w1143_,
		_w5579_
	);
	LUT3 #(
		.INIT('h80)
	) name5117 (
		_w537_,
		_w855_,
		_w856_,
		_w5580_
	);
	LUT4 #(
		.INIT('h00eb)
	) name5118 (
		_w537_,
		_w876_,
		_w1153_,
		_w5580_,
		_w5581_
	);
	LUT4 #(
		.INIT('hf100)
	) name5119 (
		_w1206_,
		_w1207_,
		_w1208_,
		_w1439_,
		_w5582_
	);
	LUT4 #(
		.INIT('h000e)
	) name5120 (
		_w1206_,
		_w1207_,
		_w1208_,
		_w1439_,
		_w5583_
	);
	LUT3 #(
		.INIT('h02)
	) name5121 (
		_w1286_,
		_w5583_,
		_w5582_,
		_w5584_
	);
	LUT4 #(
		.INIT('h0001)
	) name5122 (
		_w853_,
		_w1104_,
		_w1106_,
		_w1111_,
		_w5585_
	);
	LUT3 #(
		.INIT('h6a)
	) name5123 (
		_w853_,
		_w861_,
		_w869_,
		_w5586_
	);
	LUT3 #(
		.INIT('h13)
	) name5124 (
		_w1136_,
		_w5585_,
		_w5586_,
		_w5587_
	);
	LUT4 #(
		.INIT('h7b00)
	) name5125 (
		_w871_,
		_w1114_,
		_w1439_,
		_w5587_,
		_w5588_
	);
	LUT4 #(
		.INIT('h0700)
	) name5126 (
		_w1183_,
		_w5581_,
		_w5584_,
		_w5588_,
		_w5589_
	);
	LUT4 #(
		.INIT('hc0c8)
	) name5127 (
		_w2197_,
		_w3443_,
		_w5579_,
		_w5589_,
		_w5590_
	);
	LUT4 #(
		.INIT('h5400)
	) name5128 (
		_w1141_,
		_w2197_,
		_w3426_,
		_w3443_,
		_w5591_
	);
	LUT2 #(
		.INIT('h2)
	) name5129 (
		\P1_reg3_reg[2]/NET0131 ,
		_w5591_,
		_w5592_
	);
	LUT2 #(
		.INIT('he)
	) name5130 (
		_w5590_,
		_w5592_,
		_w5593_
	);
	LUT4 #(
		.INIT('h70d0)
	) name5131 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg0_reg[3]/NET0131 ,
		_w1476_,
		_w5594_
	);
	LUT2 #(
		.INIT('h8)
	) name5132 (
		\P2_reg0_reg[3]/NET0131 ,
		_w1487_,
		_w5595_
	);
	LUT4 #(
		.INIT('h02aa)
	) name5133 (
		\P2_reg0_reg[3]/NET0131 ,
		_w1491_,
		_w1493_,
		_w1496_,
		_w5596_
	);
	LUT4 #(
		.INIT('h08c8)
	) name5134 (
		\P2_reg0_reg[3]/NET0131 ,
		_w2081_,
		_w2272_,
		_w5530_,
		_w5597_
	);
	LUT3 #(
		.INIT('ha8)
	) name5135 (
		_w2290_,
		_w5534_,
		_w5596_,
		_w5598_
	);
	LUT4 #(
		.INIT('haaa8)
	) name5136 (
		\P2_reg0_reg[3]/NET0131 ,
		_w1491_,
		_w1493_,
		_w1496_,
		_w5599_
	);
	LUT3 #(
		.INIT('h54)
	) name5137 (
		_w2276_,
		_w5536_,
		_w5599_,
		_w5600_
	);
	LUT4 #(
		.INIT('h04c8)
	) name5138 (
		_w2110_,
		_w2277_,
		_w2353_,
		_w5533_,
		_w5601_
	);
	LUT2 #(
		.INIT('h4)
	) name5139 (
		_w1555_,
		_w2084_,
		_w5602_
	);
	LUT2 #(
		.INIT('h8)
	) name5140 (
		_w2277_,
		_w5602_,
		_w5603_
	);
	LUT3 #(
		.INIT('ha2)
	) name5141 (
		\P2_reg0_reg[3]/NET0131 ,
		_w2633_,
		_w2634_,
		_w5604_
	);
	LUT2 #(
		.INIT('h1)
	) name5142 (
		_w5603_,
		_w5604_,
		_w5605_
	);
	LUT4 #(
		.INIT('hab00)
	) name5143 (
		_w2192_,
		_w5599_,
		_w5601_,
		_w5605_,
		_w5606_
	);
	LUT4 #(
		.INIT('h0100)
	) name5144 (
		_w5600_,
		_w5598_,
		_w5597_,
		_w5606_,
		_w5607_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name5145 (
		\P1_state_reg[0]/NET0131 ,
		_w1489_,
		_w5595_,
		_w5607_,
		_w5608_
	);
	LUT2 #(
		.INIT('he)
	) name5146 (
		_w5594_,
		_w5608_,
		_w5609_
	);
	LUT4 #(
		.INIT('h70d0)
	) name5147 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg0_reg[4]/NET0131 ,
		_w1476_,
		_w5610_
	);
	LUT2 #(
		.INIT('h8)
	) name5148 (
		\P2_reg0_reg[4]/NET0131 ,
		_w1487_,
		_w5611_
	);
	LUT4 #(
		.INIT('hd11d)
	) name5149 (
		\P2_reg0_reg[4]/NET0131 ,
		_w2277_,
		_w5263_,
		_w5264_,
		_w5612_
	);
	LUT4 #(
		.INIT('h0232)
	) name5150 (
		\P2_reg0_reg[4]/NET0131 ,
		_w2192_,
		_w2277_,
		_w5266_,
		_w5613_
	);
	LUT2 #(
		.INIT('h4)
	) name5151 (
		_w1604_,
		_w2084_,
		_w5614_
	);
	LUT2 #(
		.INIT('h8)
	) name5152 (
		_w2277_,
		_w5614_,
		_w5615_
	);
	LUT3 #(
		.INIT('ha2)
	) name5153 (
		\P2_reg0_reg[4]/NET0131 ,
		_w2633_,
		_w2634_,
		_w5616_
	);
	LUT2 #(
		.INIT('h1)
	) name5154 (
		_w5615_,
		_w5616_,
		_w5617_
	);
	LUT4 #(
		.INIT('h0e00)
	) name5155 (
		_w2276_,
		_w5612_,
		_w5613_,
		_w5617_,
		_w5618_
	);
	LUT4 #(
		.INIT('hd11d)
	) name5156 (
		\P2_reg0_reg[4]/NET0131 ,
		_w2272_,
		_w5263_,
		_w5264_,
		_w5619_
	);
	LUT4 #(
		.INIT('h111d)
	) name5157 (
		\P2_reg0_reg[4]/NET0131 ,
		_w2272_,
		_w5274_,
		_w5275_,
		_w5620_
	);
	LUT4 #(
		.INIT('hf351)
	) name5158 (
		_w2081_,
		_w2290_,
		_w5619_,
		_w5620_,
		_w5621_
	);
	LUT4 #(
		.INIT('h3111)
	) name5159 (
		_w1489_,
		_w5611_,
		_w5618_,
		_w5621_,
		_w5622_
	);
	LUT3 #(
		.INIT('hce)
	) name5160 (
		\P1_state_reg[0]/NET0131 ,
		_w5610_,
		_w5622_,
		_w5623_
	);
	LUT4 #(
		.INIT('h70d0)
	) name5161 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg1_reg[3]/NET0131 ,
		_w1476_,
		_w5624_
	);
	LUT2 #(
		.INIT('h8)
	) name5162 (
		\P2_reg1_reg[3]/NET0131 ,
		_w1487_,
		_w5625_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name5163 (
		\P2_reg1_reg[3]/NET0131 ,
		_w1491_,
		_w1493_,
		_w1496_,
		_w5626_
	);
	LUT4 #(
		.INIT('h20e0)
	) name5164 (
		\P2_reg1_reg[3]/NET0131 ,
		_w1497_,
		_w2081_,
		_w5530_,
		_w5627_
	);
	LUT4 #(
		.INIT('haa02)
	) name5165 (
		\P2_reg1_reg[3]/NET0131 ,
		_w1491_,
		_w1493_,
		_w1496_,
		_w5628_
	);
	LUT4 #(
		.INIT('he010)
	) name5166 (
		_w1565_,
		_w1582_,
		_w2039_,
		_w5533_,
		_w5629_
	);
	LUT3 #(
		.INIT('ha8)
	) name5167 (
		_w2038_,
		_w5628_,
		_w5629_,
		_w5630_
	);
	LUT4 #(
		.INIT('h02a8)
	) name5168 (
		_w2039_,
		_w2110_,
		_w2353_,
		_w5533_,
		_w5631_
	);
	LUT3 #(
		.INIT('ha8)
	) name5169 (
		_w2193_,
		_w5628_,
		_w5631_,
		_w5632_
	);
	LUT4 #(
		.INIT('h02a8)
	) name5170 (
		_w1497_,
		_w2110_,
		_w2353_,
		_w5533_,
		_w5633_
	);
	LUT2 #(
		.INIT('h8)
	) name5171 (
		_w2039_,
		_w5602_,
		_w5634_
	);
	LUT3 #(
		.INIT('ha2)
	) name5172 (
		\P2_reg1_reg[3]/NET0131 ,
		_w2633_,
		_w2660_,
		_w5635_
	);
	LUT2 #(
		.INIT('h1)
	) name5173 (
		_w5634_,
		_w5635_,
		_w5636_
	);
	LUT4 #(
		.INIT('h5700)
	) name5174 (
		_w2188_,
		_w5626_,
		_w5633_,
		_w5636_,
		_w5637_
	);
	LUT4 #(
		.INIT('h0100)
	) name5175 (
		_w5627_,
		_w5630_,
		_w5632_,
		_w5637_,
		_w5638_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name5176 (
		\P1_state_reg[0]/NET0131 ,
		_w1489_,
		_w5625_,
		_w5638_,
		_w5639_
	);
	LUT2 #(
		.INIT('he)
	) name5177 (
		_w5624_,
		_w5639_,
		_w5640_
	);
	LUT4 #(
		.INIT('h70d0)
	) name5178 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg1_reg[4]/NET0131 ,
		_w1476_,
		_w5641_
	);
	LUT2 #(
		.INIT('h8)
	) name5179 (
		\P2_reg1_reg[4]/NET0131 ,
		_w1487_,
		_w5642_
	);
	LUT4 #(
		.INIT('hd11d)
	) name5180 (
		\P2_reg1_reg[4]/NET0131 ,
		_w2039_,
		_w5263_,
		_w5264_,
		_w5643_
	);
	LUT2 #(
		.INIT('h2)
	) name5181 (
		_w2038_,
		_w5643_,
		_w5644_
	);
	LUT4 #(
		.INIT('h111d)
	) name5182 (
		\P2_reg1_reg[4]/NET0131 ,
		_w1497_,
		_w5274_,
		_w5275_,
		_w5645_
	);
	LUT2 #(
		.INIT('h2)
	) name5183 (
		_w2081_,
		_w5645_,
		_w5646_
	);
	LUT4 #(
		.INIT('h20e0)
	) name5184 (
		\P2_reg1_reg[4]/NET0131 ,
		_w1497_,
		_w2188_,
		_w5266_,
		_w5647_
	);
	LUT4 #(
		.INIT('h20e0)
	) name5185 (
		\P2_reg1_reg[4]/NET0131 ,
		_w2039_,
		_w2193_,
		_w5266_,
		_w5648_
	);
	LUT2 #(
		.INIT('h8)
	) name5186 (
		_w2039_,
		_w5614_,
		_w5649_
	);
	LUT3 #(
		.INIT('ha2)
	) name5187 (
		\P2_reg1_reg[4]/NET0131 ,
		_w2633_,
		_w2660_,
		_w5650_
	);
	LUT2 #(
		.INIT('h1)
	) name5188 (
		_w5649_,
		_w5650_,
		_w5651_
	);
	LUT3 #(
		.INIT('h10)
	) name5189 (
		_w5648_,
		_w5647_,
		_w5651_,
		_w5652_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name5190 (
		_w1489_,
		_w5646_,
		_w5644_,
		_w5652_,
		_w5653_
	);
	LUT4 #(
		.INIT('heeec)
	) name5191 (
		\P1_state_reg[0]/NET0131 ,
		_w5641_,
		_w5642_,
		_w5653_,
		_w5654_
	);
	LUT4 #(
		.INIT('h70d0)
	) name5192 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg2_reg[4]/NET0131 ,
		_w1476_,
		_w5655_
	);
	LUT2 #(
		.INIT('h8)
	) name5193 (
		\P2_reg2_reg[4]/NET0131 ,
		_w1487_,
		_w5656_
	);
	LUT4 #(
		.INIT('hd11d)
	) name5194 (
		\P2_reg2_reg[4]/NET0131 ,
		_w1497_,
		_w5263_,
		_w5264_,
		_w5657_
	);
	LUT2 #(
		.INIT('h2)
	) name5195 (
		_w2038_,
		_w5657_,
		_w5658_
	);
	LUT4 #(
		.INIT('h111d)
	) name5196 (
		\P2_reg2_reg[4]/NET0131 ,
		_w2039_,
		_w5274_,
		_w5275_,
		_w5659_
	);
	LUT2 #(
		.INIT('h2)
	) name5197 (
		_w2081_,
		_w5659_,
		_w5660_
	);
	LUT4 #(
		.INIT('h20e0)
	) name5198 (
		\P2_reg2_reg[4]/NET0131 ,
		_w1497_,
		_w2193_,
		_w5266_,
		_w5661_
	);
	LUT4 #(
		.INIT('h20e0)
	) name5199 (
		\P2_reg2_reg[4]/NET0131 ,
		_w2039_,
		_w2188_,
		_w5266_,
		_w5662_
	);
	LUT3 #(
		.INIT('ha8)
	) name5200 (
		\P2_reg2_reg[4]/NET0131 ,
		_w2086_,
		_w2087_,
		_w5663_
	);
	LUT2 #(
		.INIT('h4)
	) name5201 (
		_w1596_,
		_w2088_,
		_w5664_
	);
	LUT3 #(
		.INIT('h07)
	) name5202 (
		_w1497_,
		_w5614_,
		_w5664_,
		_w5665_
	);
	LUT2 #(
		.INIT('h4)
	) name5203 (
		_w5663_,
		_w5665_,
		_w5666_
	);
	LUT3 #(
		.INIT('h10)
	) name5204 (
		_w5662_,
		_w5661_,
		_w5666_,
		_w5667_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name5205 (
		_w1489_,
		_w5660_,
		_w5658_,
		_w5667_,
		_w5668_
	);
	LUT4 #(
		.INIT('heeec)
	) name5206 (
		\P1_state_reg[0]/NET0131 ,
		_w5655_,
		_w5656_,
		_w5668_,
		_w5669_
	);
	LUT4 #(
		.INIT('h0001)
	) name5207 (
		_w861_,
		_w1104_,
		_w1106_,
		_w1111_,
		_w5670_
	);
	LUT4 #(
		.INIT('h5556)
	) name5208 (
		_w849_,
		_w857_,
		_w866_,
		_w1151_,
		_w5671_
	);
	LUT4 #(
		.INIT('h7020)
	) name5209 (
		_w537_,
		_w866_,
		_w1183_,
		_w5671_,
		_w5672_
	);
	LUT3 #(
		.INIT('h84)
	) name5210 (
		_w1206_,
		_w1286_,
		_w1436_,
		_w5673_
	);
	LUT3 #(
		.INIT('h84)
	) name5211 (
		_w870_,
		_w1114_,
		_w1436_,
		_w5674_
	);
	LUT2 #(
		.INIT('h6)
	) name5212 (
		_w861_,
		_w869_,
		_w5675_
	);
	LUT2 #(
		.INIT('h8)
	) name5213 (
		_w1136_,
		_w5675_,
		_w5676_
	);
	LUT3 #(
		.INIT('h01)
	) name5214 (
		_w5674_,
		_w5676_,
		_w5673_,
		_w5677_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name5215 (
		_w2197_,
		_w5670_,
		_w5672_,
		_w5677_,
		_w5678_
	);
	LUT2 #(
		.INIT('h4)
	) name5216 (
		_w861_,
		_w1143_,
		_w5679_
	);
	LUT4 #(
		.INIT('h80d0)
	) name5217 (
		_w537_,
		_w866_,
		_w2197_,
		_w5671_,
		_w5680_
	);
	LUT2 #(
		.INIT('h8)
	) name5218 (
		_w3143_,
		_w3443_,
		_w5681_
	);
	LUT4 #(
		.INIT('h08aa)
	) name5219 (
		\P1_reg3_reg[1]/NET0131 ,
		_w1183_,
		_w5680_,
		_w5681_,
		_w5682_
	);
	LUT4 #(
		.INIT('hffa8)
	) name5220 (
		_w3443_,
		_w5678_,
		_w5679_,
		_w5682_,
		_w5683_
	);
	LUT4 #(
		.INIT('h70d0)
	) name5221 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg3_reg[1]/NET0131 ,
		_w1476_,
		_w5684_
	);
	LUT2 #(
		.INIT('h8)
	) name5222 (
		\P2_reg3_reg[1]/NET0131 ,
		_w1487_,
		_w5685_
	);
	LUT4 #(
		.INIT('h0605)
	) name5223 (
		_w1559_,
		_w1569_,
		_w2042_,
		_w2055_,
		_w5686_
	);
	LUT3 #(
		.INIT('h70)
	) name5224 (
		_w1576_,
		_w1577_,
		_w2042_,
		_w5687_
	);
	LUT4 #(
		.INIT('h111d)
	) name5225 (
		\P2_reg3_reg[1]/NET0131 ,
		_w2277_,
		_w5686_,
		_w5687_,
		_w5688_
	);
	LUT4 #(
		.INIT('h02aa)
	) name5226 (
		\P2_reg3_reg[1]/NET0131 ,
		_w1491_,
		_w1493_,
		_w1496_,
		_w5689_
	);
	LUT3 #(
		.INIT('h87)
	) name5227 (
		_w1567_,
		_w1568_,
		_w1573_,
		_w5690_
	);
	LUT4 #(
		.INIT('h35c5)
	) name5228 (
		\P2_reg3_reg[1]/NET0131 ,
		_w2112_,
		_w2272_,
		_w5690_,
		_w5691_
	);
	LUT4 #(
		.INIT('h00e0)
	) name5229 (
		_w1491_,
		_w1493_,
		_w1496_,
		_w1573_,
		_w5692_
	);
	LUT4 #(
		.INIT('h4c5f)
	) name5230 (
		\P2_reg3_reg[1]/NET0131 ,
		_w1573_,
		_w2086_,
		_w2088_,
		_w5693_
	);
	LUT4 #(
		.INIT('h5700)
	) name5231 (
		_w2084_,
		_w5689_,
		_w5692_,
		_w5693_,
		_w5694_
	);
	LUT3 #(
		.INIT('he0)
	) name5232 (
		_w2192_,
		_w5691_,
		_w5694_,
		_w5695_
	);
	LUT4 #(
		.INIT('h35c5)
	) name5233 (
		\P2_reg3_reg[1]/NET0131 ,
		_w1581_,
		_w2277_,
		_w5690_,
		_w5696_
	);
	LUT4 #(
		.INIT('h35c5)
	) name5234 (
		\P2_reg3_reg[1]/NET0131 ,
		_w1581_,
		_w2272_,
		_w5690_,
		_w5697_
	);
	LUT4 #(
		.INIT('hf3a2)
	) name5235 (
		_w2276_,
		_w2290_,
		_w5696_,
		_w5697_,
		_w5698_
	);
	LUT4 #(
		.INIT('hd000)
	) name5236 (
		_w2081_,
		_w5688_,
		_w5695_,
		_w5698_,
		_w5699_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name5237 (
		\P1_state_reg[0]/NET0131 ,
		_w1489_,
		_w5685_,
		_w5699_,
		_w5700_
	);
	LUT2 #(
		.INIT('he)
	) name5238 (
		_w5684_,
		_w5700_,
		_w5701_
	);
	LUT2 #(
		.INIT('h2)
	) name5239 (
		\P1_reg2_reg[2]/NET0131 ,
		_w5381_,
		_w5702_
	);
	LUT2 #(
		.INIT('h8)
	) name5240 (
		\P1_reg3_reg[2]/NET0131 ,
		_w1143_,
		_w5703_
	);
	LUT4 #(
		.INIT('hcc08)
	) name5241 (
		_w534_,
		_w3443_,
		_w5589_,
		_w5703_,
		_w5704_
	);
	LUT2 #(
		.INIT('he)
	) name5242 (
		_w5702_,
		_w5704_,
		_w5705_
	);
	LUT4 #(
		.INIT('h70d0)
	) name5243 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg1_reg[2]/NET0131 ,
		_w1476_,
		_w5706_
	);
	LUT2 #(
		.INIT('h8)
	) name5244 (
		\P2_reg1_reg[2]/NET0131 ,
		_w1487_,
		_w5707_
	);
	LUT3 #(
		.INIT('h70)
	) name5245 (
		_w1567_,
		_w1568_,
		_w2042_,
		_w5708_
	);
	LUT4 #(
		.INIT('h00de)
	) name5246 (
		_w1550_,
		_w2042_,
		_w2056_,
		_w5708_,
		_w5709_
	);
	LUT4 #(
		.INIT('h20e0)
	) name5247 (
		\P2_reg1_reg[2]/NET0131 ,
		_w1497_,
		_w2081_,
		_w5709_,
		_w5710_
	);
	LUT3 #(
		.INIT('h87)
	) name5248 (
		_w1557_,
		_w1558_,
		_w1564_,
		_w5711_
	);
	LUT4 #(
		.INIT('hb24d)
	) name5249 (
		_w1569_,
		_w1573_,
		_w2112_,
		_w5711_,
		_w5712_
	);
	LUT4 #(
		.INIT('he020)
	) name5250 (
		\P2_reg1_reg[2]/NET0131 ,
		_w1497_,
		_w2188_,
		_w5712_,
		_w5713_
	);
	LUT2 #(
		.INIT('h4)
	) name5251 (
		_w1564_,
		_w2084_,
		_w5714_
	);
	LUT2 #(
		.INIT('h8)
	) name5252 (
		_w2039_,
		_w5714_,
		_w5715_
	);
	LUT3 #(
		.INIT('ha2)
	) name5253 (
		\P2_reg1_reg[2]/NET0131 ,
		_w2633_,
		_w2660_,
		_w5716_
	);
	LUT2 #(
		.INIT('h1)
	) name5254 (
		_w5715_,
		_w5716_,
		_w5717_
	);
	LUT4 #(
		.INIT('hab54)
	) name5255 (
		_w1574_,
		_w1575_,
		_w1581_,
		_w5711_,
		_w5718_
	);
	LUT4 #(
		.INIT('h08c8)
	) name5256 (
		\P2_reg1_reg[2]/NET0131 ,
		_w2038_,
		_w2039_,
		_w5718_,
		_w5719_
	);
	LUT4 #(
		.INIT('he020)
	) name5257 (
		\P2_reg1_reg[2]/NET0131 ,
		_w2039_,
		_w2193_,
		_w5712_,
		_w5720_
	);
	LUT4 #(
		.INIT('h0100)
	) name5258 (
		_w5713_,
		_w5719_,
		_w5720_,
		_w5717_,
		_w5721_
	);
	LUT4 #(
		.INIT('h1311)
	) name5259 (
		_w1489_,
		_w5707_,
		_w5710_,
		_w5721_,
		_w5722_
	);
	LUT3 #(
		.INIT('hce)
	) name5260 (
		\P1_state_reg[0]/NET0131 ,
		_w5706_,
		_w5722_,
		_w5723_
	);
	LUT4 #(
		.INIT('h70d0)
	) name5261 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg2_reg[2]/NET0131 ,
		_w1476_,
		_w5724_
	);
	LUT2 #(
		.INIT('h8)
	) name5262 (
		\P2_reg2_reg[2]/NET0131 ,
		_w1487_,
		_w5725_
	);
	LUT4 #(
		.INIT('h20e0)
	) name5263 (
		\P2_reg2_reg[2]/NET0131 ,
		_w2039_,
		_w2081_,
		_w5709_,
		_w5726_
	);
	LUT4 #(
		.INIT('he020)
	) name5264 (
		\P2_reg2_reg[2]/NET0131 ,
		_w1497_,
		_w2193_,
		_w5712_,
		_w5727_
	);
	LUT3 #(
		.INIT('ha8)
	) name5265 (
		\P2_reg2_reg[2]/NET0131 ,
		_w2086_,
		_w2087_,
		_w5728_
	);
	LUT2 #(
		.INIT('h8)
	) name5266 (
		\P2_reg3_reg[2]/NET0131 ,
		_w2088_,
		_w5729_
	);
	LUT3 #(
		.INIT('h07)
	) name5267 (
		_w1497_,
		_w5714_,
		_w5729_,
		_w5730_
	);
	LUT2 #(
		.INIT('h4)
	) name5268 (
		_w5728_,
		_w5730_,
		_w5731_
	);
	LUT4 #(
		.INIT('he020)
	) name5269 (
		\P2_reg2_reg[2]/NET0131 ,
		_w2039_,
		_w2188_,
		_w5712_,
		_w5732_
	);
	LUT4 #(
		.INIT('h20e0)
	) name5270 (
		\P2_reg2_reg[2]/NET0131 ,
		_w1497_,
		_w2038_,
		_w5718_,
		_w5733_
	);
	LUT4 #(
		.INIT('h0100)
	) name5271 (
		_w5727_,
		_w5732_,
		_w5733_,
		_w5731_,
		_w5734_
	);
	LUT4 #(
		.INIT('h1311)
	) name5272 (
		_w1489_,
		_w5725_,
		_w5726_,
		_w5734_,
		_w5735_
	);
	LUT3 #(
		.INIT('hce)
	) name5273 (
		\P1_state_reg[0]/NET0131 ,
		_w5724_,
		_w5735_,
		_w5736_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name5274 (
		_w3651_,
		_w5670_,
		_w5672_,
		_w5677_,
		_w5737_
	);
	LUT3 #(
		.INIT('h2a)
	) name5275 (
		\P1_reg0_reg[1]/NET0131 ,
		_w3633_,
		_w5103_,
		_w5738_
	);
	LUT2 #(
		.INIT('he)
	) name5276 (
		_w5737_,
		_w5738_,
		_w5739_
	);
	LUT3 #(
		.INIT('ha2)
	) name5277 (
		\P1_reg0_reg[2]/NET0131 ,
		_w3658_,
		_w3659_,
		_w5740_
	);
	LUT3 #(
		.INIT('hf2)
	) name5278 (
		_w3651_,
		_w5589_,
		_w5740_,
		_w5741_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name5279 (
		_w4074_,
		_w5670_,
		_w5672_,
		_w5677_,
		_w5742_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name5280 (
		\P1_reg1_reg[1]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w2425_,
		_w4073_,
		_w5743_
	);
	LUT2 #(
		.INIT('he)
	) name5281 (
		_w5742_,
		_w5743_,
		_w5744_
	);
	LUT2 #(
		.INIT('h8)
	) name5282 (
		\P1_reg1_reg[2]/NET0131 ,
		_w1183_,
		_w5745_
	);
	LUT3 #(
		.INIT('hd0)
	) name5283 (
		_w2421_,
		_w5581_,
		_w5745_,
		_w5746_
	);
	LUT4 #(
		.INIT('hcc08)
	) name5284 (
		_w2421_,
		_w3443_,
		_w5589_,
		_w5746_,
		_w5747_
	);
	LUT2 #(
		.INIT('h2)
	) name5285 (
		\P1_reg1_reg[2]/NET0131 ,
		_w4079_,
		_w5748_
	);
	LUT2 #(
		.INIT('he)
	) name5286 (
		_w5747_,
		_w5748_,
		_w5749_
	);
	LUT4 #(
		.INIT('h70d0)
	) name5287 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg0_reg[1]/NET0131 ,
		_w1476_,
		_w5750_
	);
	LUT2 #(
		.INIT('h8)
	) name5288 (
		\P2_reg0_reg[1]/NET0131 ,
		_w1487_,
		_w5751_
	);
	LUT4 #(
		.INIT('h111d)
	) name5289 (
		\P2_reg0_reg[1]/NET0131 ,
		_w2272_,
		_w5686_,
		_w5687_,
		_w5752_
	);
	LUT4 #(
		.INIT('haaa8)
	) name5290 (
		\P2_reg0_reg[1]/NET0131 ,
		_w1491_,
		_w1493_,
		_w1496_,
		_w5753_
	);
	LUT4 #(
		.INIT('h35c5)
	) name5291 (
		\P2_reg0_reg[1]/NET0131 ,
		_w1581_,
		_w2277_,
		_w5690_,
		_w5754_
	);
	LUT2 #(
		.INIT('h2)
	) name5292 (
		\P2_reg0_reg[1]/NET0131 ,
		_w2633_,
		_w5755_
	);
	LUT4 #(
		.INIT('h0001)
	) name5293 (
		_w1491_,
		_w1493_,
		_w1496_,
		_w1573_,
		_w5756_
	);
	LUT4 #(
		.INIT('h1113)
	) name5294 (
		_w2084_,
		_w5755_,
		_w5753_,
		_w5756_,
		_w5757_
	);
	LUT3 #(
		.INIT('he0)
	) name5295 (
		_w2276_,
		_w5754_,
		_w5757_,
		_w5758_
	);
	LUT4 #(
		.INIT('h35c5)
	) name5296 (
		\P2_reg0_reg[1]/NET0131 ,
		_w1581_,
		_w2272_,
		_w5690_,
		_w5759_
	);
	LUT4 #(
		.INIT('h35c5)
	) name5297 (
		\P2_reg0_reg[1]/NET0131 ,
		_w2112_,
		_w2277_,
		_w5690_,
		_w5760_
	);
	LUT4 #(
		.INIT('hf3a2)
	) name5298 (
		_w2192_,
		_w2290_,
		_w5759_,
		_w5760_,
		_w5761_
	);
	LUT4 #(
		.INIT('hd000)
	) name5299 (
		_w2081_,
		_w5752_,
		_w5758_,
		_w5761_,
		_w5762_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name5300 (
		\P1_state_reg[0]/NET0131 ,
		_w1489_,
		_w5751_,
		_w5762_,
		_w5763_
	);
	LUT2 #(
		.INIT('he)
	) name5301 (
		_w5750_,
		_w5763_,
		_w5764_
	);
	LUT2 #(
		.INIT('h2)
	) name5302 (
		\P1_reg2_reg[1]/NET0131 ,
		_w511_,
		_w5765_
	);
	LUT2 #(
		.INIT('h8)
	) name5303 (
		\P1_reg2_reg[1]/NET0131 ,
		_w524_,
		_w5766_
	);
	LUT3 #(
		.INIT('ha2)
	) name5304 (
		\P1_reg2_reg[1]/NET0131 ,
		_w534_,
		_w1141_,
		_w5767_
	);
	LUT3 #(
		.INIT('h31)
	) name5305 (
		\P1_reg2_reg[1]/NET0131 ,
		_w534_,
		_w2259_,
		_w5768_
	);
	LUT4 #(
		.INIT('h00fb)
	) name5306 (
		_w5672_,
		_w5677_,
		_w5767_,
		_w5768_,
		_w5769_
	);
	LUT4 #(
		.INIT('h1000)
	) name5307 (
		_w528_,
		_w530_,
		_w533_,
		_w861_,
		_w5770_
	);
	LUT4 #(
		.INIT('h5455)
	) name5308 (
		\P1_reg2_reg[1]/NET0131 ,
		_w528_,
		_w530_,
		_w533_,
		_w5771_
	);
	LUT3 #(
		.INIT('h02)
	) name5309 (
		_w1138_,
		_w5771_,
		_w5770_,
		_w5772_
	);
	LUT2 #(
		.INIT('h8)
	) name5310 (
		\P1_reg3_reg[1]/NET0131 ,
		_w1143_,
		_w5773_
	);
	LUT2 #(
		.INIT('h1)
	) name5311 (
		_w5772_,
		_w5773_,
		_w5774_
	);
	LUT4 #(
		.INIT('h1311)
	) name5312 (
		_w526_,
		_w5766_,
		_w5769_,
		_w5774_,
		_w5775_
	);
	LUT3 #(
		.INIT('hce)
	) name5313 (
		\P1_state_reg[0]/NET0131 ,
		_w5765_,
		_w5775_,
		_w5776_
	);
	LUT4 #(
		.INIT('h70d0)
	) name5314 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg1_reg[1]/NET0131 ,
		_w1476_,
		_w5777_
	);
	LUT2 #(
		.INIT('h8)
	) name5315 (
		\P2_reg1_reg[1]/NET0131 ,
		_w1487_,
		_w5778_
	);
	LUT4 #(
		.INIT('h111d)
	) name5316 (
		\P2_reg1_reg[1]/NET0131 ,
		_w1497_,
		_w5686_,
		_w5687_,
		_w5779_
	);
	LUT4 #(
		.INIT('haa02)
	) name5317 (
		\P2_reg1_reg[1]/NET0131 ,
		_w1491_,
		_w1493_,
		_w1496_,
		_w5780_
	);
	LUT4 #(
		.INIT('h1dd1)
	) name5318 (
		\P2_reg1_reg[1]/NET0131 ,
		_w2039_,
		_w2112_,
		_w5690_,
		_w5781_
	);
	LUT2 #(
		.INIT('h2)
	) name5319 (
		\P2_reg1_reg[1]/NET0131 ,
		_w2633_,
		_w5782_
	);
	LUT4 #(
		.INIT('h000e)
	) name5320 (
		_w1491_,
		_w1493_,
		_w1496_,
		_w1573_,
		_w5783_
	);
	LUT4 #(
		.INIT('h1113)
	) name5321 (
		_w2084_,
		_w5782_,
		_w5780_,
		_w5783_,
		_w5784_
	);
	LUT3 #(
		.INIT('hd0)
	) name5322 (
		_w2193_,
		_w5781_,
		_w5784_,
		_w5785_
	);
	LUT4 #(
		.INIT('h1dd1)
	) name5323 (
		\P2_reg1_reg[1]/NET0131 ,
		_w1497_,
		_w2112_,
		_w5690_,
		_w5786_
	);
	LUT4 #(
		.INIT('h35c5)
	) name5324 (
		\P2_reg1_reg[1]/NET0131 ,
		_w1581_,
		_w2039_,
		_w5690_,
		_w5787_
	);
	LUT4 #(
		.INIT('hf351)
	) name5325 (
		_w2038_,
		_w2188_,
		_w5786_,
		_w5787_,
		_w5788_
	);
	LUT4 #(
		.INIT('hd000)
	) name5326 (
		_w2081_,
		_w5779_,
		_w5785_,
		_w5788_,
		_w5789_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name5327 (
		\P1_state_reg[0]/NET0131 ,
		_w1489_,
		_w5778_,
		_w5789_,
		_w5790_
	);
	LUT2 #(
		.INIT('he)
	) name5328 (
		_w5777_,
		_w5790_,
		_w5791_
	);
	LUT4 #(
		.INIT('h70d0)
	) name5329 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg2_reg[1]/NET0131 ,
		_w1476_,
		_w5792_
	);
	LUT2 #(
		.INIT('h8)
	) name5330 (
		\P2_reg2_reg[1]/NET0131 ,
		_w1487_,
		_w5793_
	);
	LUT4 #(
		.INIT('h111d)
	) name5331 (
		\P2_reg2_reg[1]/NET0131 ,
		_w2039_,
		_w5686_,
		_w5687_,
		_w5794_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name5332 (
		\P2_reg2_reg[1]/NET0131 ,
		_w1491_,
		_w1493_,
		_w1496_,
		_w5795_
	);
	LUT4 #(
		.INIT('h1dd1)
	) name5333 (
		\P2_reg2_reg[1]/NET0131 ,
		_w1497_,
		_w2112_,
		_w5690_,
		_w5796_
	);
	LUT4 #(
		.INIT('h0010)
	) name5334 (
		_w1491_,
		_w1493_,
		_w1496_,
		_w1573_,
		_w5797_
	);
	LUT4 #(
		.INIT('h135f)
	) name5335 (
		\P2_reg2_reg[1]/NET0131 ,
		\P2_reg3_reg[1]/NET0131 ,
		_w2086_,
		_w2088_,
		_w5798_
	);
	LUT4 #(
		.INIT('h5700)
	) name5336 (
		_w2084_,
		_w5795_,
		_w5797_,
		_w5798_,
		_w5799_
	);
	LUT3 #(
		.INIT('hd0)
	) name5337 (
		_w2193_,
		_w5796_,
		_w5799_,
		_w5800_
	);
	LUT4 #(
		.INIT('h1dd1)
	) name5338 (
		\P2_reg2_reg[1]/NET0131 ,
		_w2039_,
		_w2112_,
		_w5690_,
		_w5801_
	);
	LUT4 #(
		.INIT('h1dd1)
	) name5339 (
		\P2_reg2_reg[1]/NET0131 ,
		_w1497_,
		_w1581_,
		_w5690_,
		_w5802_
	);
	LUT4 #(
		.INIT('hf351)
	) name5340 (
		_w2038_,
		_w2188_,
		_w5801_,
		_w5802_,
		_w5803_
	);
	LUT4 #(
		.INIT('hd000)
	) name5341 (
		_w2081_,
		_w5794_,
		_w5800_,
		_w5803_,
		_w5804_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name5342 (
		\P1_state_reg[0]/NET0131 ,
		_w1489_,
		_w5793_,
		_w5804_,
		_w5805_
	);
	LUT2 #(
		.INIT('he)
	) name5343 (
		_w5792_,
		_w5805_,
		_w5806_
	);
	LUT4 #(
		.INIT('h70d0)
	) name5344 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg3_reg[0]/NET0131 ,
		_w1476_,
		_w5807_
	);
	LUT2 #(
		.INIT('h8)
	) name5345 (
		\P2_reg3_reg[0]/NET0131 ,
		_w1487_,
		_w5808_
	);
	LUT4 #(
		.INIT('haaa8)
	) name5346 (
		\P2_reg3_reg[0]/NET0131 ,
		_w1491_,
		_w1493_,
		_w1496_,
		_w5809_
	);
	LUT4 #(
		.INIT('h2100)
	) name5347 (
		_w1569_,
		_w2042_,
		_w2055_,
		_w2277_,
		_w5810_
	);
	LUT3 #(
		.INIT('ha8)
	) name5348 (
		_w2081_,
		_w5809_,
		_w5810_,
		_w5811_
	);
	LUT4 #(
		.INIT('h02aa)
	) name5349 (
		\P2_reg3_reg[0]/NET0131 ,
		_w1491_,
		_w1493_,
		_w1496_,
		_w5812_
	);
	LUT3 #(
		.INIT('h70)
	) name5350 (
		_w1576_,
		_w1577_,
		_w1580_,
		_w5813_
	);
	LUT3 #(
		.INIT('h87)
	) name5351 (
		_w1576_,
		_w1577_,
		_w1580_,
		_w5814_
	);
	LUT4 #(
		.INIT('hcbc3)
	) name5352 (
		_w1811_,
		_w2033_,
		_w2035_,
		_w2036_,
		_w5815_
	);
	LUT4 #(
		.INIT('h002e)
	) name5353 (
		\P2_reg3_reg[0]/NET0131 ,
		_w2272_,
		_w5814_,
		_w5815_,
		_w5816_
	);
	LUT4 #(
		.INIT('h4c5f)
	) name5354 (
		\P2_reg3_reg[0]/NET0131 ,
		_w1580_,
		_w2086_,
		_w2088_,
		_w5817_
	);
	LUT4 #(
		.INIT('h00e0)
	) name5355 (
		_w1491_,
		_w1493_,
		_w1496_,
		_w1580_,
		_w5818_
	);
	LUT3 #(
		.INIT('ha8)
	) name5356 (
		_w2084_,
		_w5812_,
		_w5818_,
		_w5819_
	);
	LUT4 #(
		.INIT('h20e0)
	) name5357 (
		\P2_reg3_reg[0]/NET0131 ,
		_w2277_,
		_w2290_,
		_w5814_,
		_w5820_
	);
	LUT4 #(
		.INIT('h0100)
	) name5358 (
		_w5816_,
		_w5819_,
		_w5820_,
		_w5817_,
		_w5821_
	);
	LUT4 #(
		.INIT('h1311)
	) name5359 (
		_w1489_,
		_w5808_,
		_w5811_,
		_w5821_,
		_w5822_
	);
	LUT3 #(
		.INIT('hce)
	) name5360 (
		\P1_state_reg[0]/NET0131 ,
		_w5807_,
		_w5822_,
		_w5823_
	);
	LUT4 #(
		.INIT('h70d0)
	) name5361 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg1_reg[0]/NET0131 ,
		_w1476_,
		_w5824_
	);
	LUT2 #(
		.INIT('h8)
	) name5362 (
		\P2_reg1_reg[0]/NET0131 ,
		_w1487_,
		_w5825_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name5363 (
		\P2_reg1_reg[0]/NET0131 ,
		_w1491_,
		_w1493_,
		_w1496_,
		_w5826_
	);
	LUT4 #(
		.INIT('h0802)
	) name5364 (
		_w1497_,
		_w1569_,
		_w2042_,
		_w2055_,
		_w5827_
	);
	LUT3 #(
		.INIT('ha8)
	) name5365 (
		_w2081_,
		_w5826_,
		_w5827_,
		_w5828_
	);
	LUT4 #(
		.INIT('haa02)
	) name5366 (
		\P2_reg1_reg[0]/NET0131 ,
		_w1491_,
		_w1493_,
		_w1496_,
		_w5829_
	);
	LUT4 #(
		.INIT('h383c)
	) name5367 (
		_w1811_,
		_w2033_,
		_w2035_,
		_w2036_,
		_w5830_
	);
	LUT4 #(
		.INIT('h2e00)
	) name5368 (
		\P2_reg1_reg[0]/NET0131 ,
		_w2039_,
		_w5814_,
		_w5830_,
		_w5831_
	);
	LUT2 #(
		.INIT('h2)
	) name5369 (
		\P2_reg1_reg[0]/NET0131 ,
		_w2633_,
		_w5832_
	);
	LUT4 #(
		.INIT('h20e0)
	) name5370 (
		\P2_reg1_reg[0]/NET0131 ,
		_w1497_,
		_w2188_,
		_w5814_,
		_w5833_
	);
	LUT4 #(
		.INIT('h000e)
	) name5371 (
		_w1491_,
		_w1493_,
		_w1496_,
		_w1580_,
		_w5834_
	);
	LUT3 #(
		.INIT('ha8)
	) name5372 (
		_w2084_,
		_w5829_,
		_w5834_,
		_w5835_
	);
	LUT4 #(
		.INIT('h0001)
	) name5373 (
		_w5831_,
		_w5833_,
		_w5835_,
		_w5832_,
		_w5836_
	);
	LUT4 #(
		.INIT('h1311)
	) name5374 (
		_w1489_,
		_w5825_,
		_w5828_,
		_w5836_,
		_w5837_
	);
	LUT3 #(
		.INIT('hce)
	) name5375 (
		\P1_state_reg[0]/NET0131 ,
		_w5824_,
		_w5837_,
		_w5838_
	);
	LUT4 #(
		.INIT('h70d0)
	) name5376 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg2_reg[0]/NET0131 ,
		_w1476_,
		_w5839_
	);
	LUT2 #(
		.INIT('h8)
	) name5377 (
		\P2_reg2_reg[0]/NET0131 ,
		_w1487_,
		_w5840_
	);
	LUT4 #(
		.INIT('haa02)
	) name5378 (
		\P2_reg2_reg[0]/NET0131 ,
		_w1491_,
		_w1493_,
		_w1496_,
		_w5841_
	);
	LUT4 #(
		.INIT('h0804)
	) name5379 (
		_w1569_,
		_w2039_,
		_w2042_,
		_w2055_,
		_w5842_
	);
	LUT3 #(
		.INIT('ha8)
	) name5380 (
		_w2081_,
		_w5841_,
		_w5842_,
		_w5843_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name5381 (
		\P2_reg2_reg[0]/NET0131 ,
		_w1491_,
		_w1493_,
		_w1496_,
		_w5844_
	);
	LUT4 #(
		.INIT('h2e00)
	) name5382 (
		\P2_reg2_reg[0]/NET0131 ,
		_w1497_,
		_w5814_,
		_w5830_,
		_w5845_
	);
	LUT4 #(
		.INIT('h135f)
	) name5383 (
		\P2_reg2_reg[0]/NET0131 ,
		\P2_reg3_reg[0]/NET0131 ,
		_w2086_,
		_w2088_,
		_w5846_
	);
	LUT4 #(
		.INIT('h20e0)
	) name5384 (
		\P2_reg2_reg[0]/NET0131 ,
		_w2039_,
		_w2188_,
		_w5814_,
		_w5847_
	);
	LUT4 #(
		.INIT('h0010)
	) name5385 (
		_w1491_,
		_w1493_,
		_w1496_,
		_w1580_,
		_w5848_
	);
	LUT3 #(
		.INIT('ha8)
	) name5386 (
		_w2084_,
		_w5844_,
		_w5848_,
		_w5849_
	);
	LUT4 #(
		.INIT('h0100)
	) name5387 (
		_w5845_,
		_w5847_,
		_w5849_,
		_w5846_,
		_w5850_
	);
	LUT4 #(
		.INIT('h1311)
	) name5388 (
		_w1489_,
		_w5840_,
		_w5843_,
		_w5850_,
		_w5851_
	);
	LUT3 #(
		.INIT('hce)
	) name5389 (
		\P1_state_reg[0]/NET0131 ,
		_w5839_,
		_w5851_,
		_w5852_
	);
	LUT4 #(
		.INIT('h70d0)
	) name5390 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg0_reg[0]/NET0131 ,
		_w1476_,
		_w5853_
	);
	LUT2 #(
		.INIT('h8)
	) name5391 (
		\P2_reg0_reg[0]/NET0131 ,
		_w1487_,
		_w5854_
	);
	LUT4 #(
		.INIT('h02aa)
	) name5392 (
		\P2_reg0_reg[0]/NET0131 ,
		_w1491_,
		_w1493_,
		_w1496_,
		_w5855_
	);
	LUT4 #(
		.INIT('h2100)
	) name5393 (
		_w1569_,
		_w2042_,
		_w2055_,
		_w2272_,
		_w5856_
	);
	LUT3 #(
		.INIT('ha8)
	) name5394 (
		_w2081_,
		_w5855_,
		_w5856_,
		_w5857_
	);
	LUT4 #(
		.INIT('haaa8)
	) name5395 (
		\P2_reg0_reg[0]/NET0131 ,
		_w1491_,
		_w1493_,
		_w1496_,
		_w5858_
	);
	LUT4 #(
		.INIT('h0001)
	) name5396 (
		_w1491_,
		_w1493_,
		_w1496_,
		_w1580_,
		_w5859_
	);
	LUT2 #(
		.INIT('h2)
	) name5397 (
		\P2_reg0_reg[0]/NET0131 ,
		_w2633_,
		_w5860_
	);
	LUT4 #(
		.INIT('h0057)
	) name5398 (
		_w2084_,
		_w5858_,
		_w5859_,
		_w5860_,
		_w5861_
	);
	LUT4 #(
		.INIT('h20e0)
	) name5399 (
		\P2_reg0_reg[0]/NET0131 ,
		_w2272_,
		_w2290_,
		_w5814_,
		_w5862_
	);
	LUT4 #(
		.INIT('h002e)
	) name5400 (
		\P2_reg0_reg[0]/NET0131 ,
		_w2277_,
		_w5814_,
		_w5815_,
		_w5863_
	);
	LUT3 #(
		.INIT('h10)
	) name5401 (
		_w5862_,
		_w5863_,
		_w5861_,
		_w5864_
	);
	LUT4 #(
		.INIT('h1311)
	) name5402 (
		_w1489_,
		_w5854_,
		_w5857_,
		_w5864_,
		_w5865_
	);
	LUT3 #(
		.INIT('hce)
	) name5403 (
		\P1_state_reg[0]/NET0131 ,
		_w5853_,
		_w5865_,
		_w5866_
	);
	LUT2 #(
		.INIT('h2)
	) name5404 (
		\P1_reg3_reg[0]/NET0131 ,
		_w511_,
		_w5867_
	);
	LUT2 #(
		.INIT('h8)
	) name5405 (
		\P1_reg3_reg[0]/NET0131 ,
		_w524_,
		_w5868_
	);
	LUT4 #(
		.INIT('h02aa)
	) name5406 (
		\P1_reg3_reg[0]/NET0131 ,
		_w528_,
		_w530_,
		_w533_,
		_w5869_
	);
	LUT4 #(
		.INIT('h1114)
	) name5407 (
		_w537_,
		_w857_,
		_w866_,
		_w1151_,
		_w5870_
	);
	LUT4 #(
		.INIT('hc808)
	) name5408 (
		\P1_reg3_reg[0]/NET0131 ,
		_w1183_,
		_w2197_,
		_w5870_,
		_w5871_
	);
	LUT4 #(
		.INIT('h0c88)
	) name5409 (
		\P1_reg3_reg[0]/NET0131 ,
		_w1109_,
		_w1435_,
		_w2197_,
		_w5872_
	);
	LUT4 #(
		.INIT('h00e0)
	) name5410 (
		_w528_,
		_w530_,
		_w533_,
		_w869_,
		_w5873_
	);
	LUT3 #(
		.INIT('ha8)
	) name5411 (
		_w3656_,
		_w5869_,
		_w5873_,
		_w5874_
	);
	LUT4 #(
		.INIT('h4c5f)
	) name5412 (
		\P1_reg3_reg[0]/NET0131 ,
		_w869_,
		_w1141_,
		_w1143_,
		_w5875_
	);
	LUT3 #(
		.INIT('h10)
	) name5413 (
		_w5874_,
		_w5872_,
		_w5875_,
		_w5876_
	);
	LUT4 #(
		.INIT('h1311)
	) name5414 (
		_w526_,
		_w5868_,
		_w5871_,
		_w5876_,
		_w5877_
	);
	LUT3 #(
		.INIT('hce)
	) name5415 (
		\P1_state_reg[0]/NET0131 ,
		_w5867_,
		_w5877_,
		_w5878_
	);
	LUT2 #(
		.INIT('h2)
	) name5416 (
		\P1_reg2_reg[0]/NET0131 ,
		_w511_,
		_w5879_
	);
	LUT2 #(
		.INIT('h8)
	) name5417 (
		\P1_reg2_reg[0]/NET0131 ,
		_w524_,
		_w5880_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name5418 (
		\P1_reg2_reg[0]/NET0131 ,
		_w528_,
		_w530_,
		_w533_,
		_w5881_
	);
	LUT4 #(
		.INIT('he020)
	) name5419 (
		\P1_reg2_reg[0]/NET0131 ,
		_w534_,
		_w1183_,
		_w5870_,
		_w5882_
	);
	LUT4 #(
		.INIT('h20e0)
	) name5420 (
		\P1_reg2_reg[0]/NET0131 ,
		_w534_,
		_w1109_,
		_w1435_,
		_w5883_
	);
	LUT4 #(
		.INIT('h0010)
	) name5421 (
		_w528_,
		_w530_,
		_w533_,
		_w869_,
		_w5884_
	);
	LUT3 #(
		.INIT('ha8)
	) name5422 (
		_w3656_,
		_w5881_,
		_w5884_,
		_w5885_
	);
	LUT4 #(
		.INIT('h135f)
	) name5423 (
		\P1_reg2_reg[0]/NET0131 ,
		\P1_reg3_reg[0]/NET0131 ,
		_w1141_,
		_w1143_,
		_w5886_
	);
	LUT3 #(
		.INIT('h10)
	) name5424 (
		_w5885_,
		_w5883_,
		_w5886_,
		_w5887_
	);
	LUT4 #(
		.INIT('h1311)
	) name5425 (
		_w526_,
		_w5880_,
		_w5882_,
		_w5887_,
		_w5888_
	);
	LUT3 #(
		.INIT('hce)
	) name5426 (
		\P1_state_reg[0]/NET0131 ,
		_w5879_,
		_w5888_,
		_w5889_
	);
	LUT2 #(
		.INIT('h2)
	) name5427 (
		\P1_reg0_reg[0]/NET0131 ,
		_w511_,
		_w5890_
	);
	LUT2 #(
		.INIT('h8)
	) name5428 (
		\P1_reg0_reg[0]/NET0131 ,
		_w524_,
		_w5891_
	);
	LUT4 #(
		.INIT('haaa8)
	) name5429 (
		\P1_reg0_reg[0]/NET0131 ,
		_w528_,
		_w530_,
		_w533_,
		_w5892_
	);
	LUT4 #(
		.INIT('hc808)
	) name5430 (
		\P1_reg0_reg[0]/NET0131 ,
		_w1183_,
		_w2688_,
		_w5870_,
		_w5893_
	);
	LUT4 #(
		.INIT('h0001)
	) name5431 (
		_w528_,
		_w530_,
		_w533_,
		_w869_,
		_w5894_
	);
	LUT3 #(
		.INIT('ha8)
	) name5432 (
		_w3656_,
		_w5892_,
		_w5894_,
		_w5895_
	);
	LUT2 #(
		.INIT('h2)
	) name5433 (
		\P1_reg0_reg[0]/NET0131 ,
		_w2425_,
		_w5896_
	);
	LUT4 #(
		.INIT('h0c88)
	) name5434 (
		\P1_reg0_reg[0]/NET0131 ,
		_w1109_,
		_w1435_,
		_w2688_,
		_w5897_
	);
	LUT3 #(
		.INIT('h01)
	) name5435 (
		_w5896_,
		_w5897_,
		_w5895_,
		_w5898_
	);
	LUT4 #(
		.INIT('h1311)
	) name5436 (
		_w526_,
		_w5891_,
		_w5893_,
		_w5898_,
		_w5899_
	);
	LUT3 #(
		.INIT('hce)
	) name5437 (
		\P1_state_reg[0]/NET0131 ,
		_w5890_,
		_w5899_,
		_w5900_
	);
	LUT2 #(
		.INIT('h2)
	) name5438 (
		\P1_reg1_reg[0]/NET0131 ,
		_w511_,
		_w5901_
	);
	LUT2 #(
		.INIT('h8)
	) name5439 (
		\P1_reg1_reg[0]/NET0131 ,
		_w524_,
		_w5902_
	);
	LUT4 #(
		.INIT('haa02)
	) name5440 (
		\P1_reg1_reg[0]/NET0131 ,
		_w528_,
		_w530_,
		_w533_,
		_w5903_
	);
	LUT4 #(
		.INIT('hc808)
	) name5441 (
		\P1_reg1_reg[0]/NET0131 ,
		_w1183_,
		_w2421_,
		_w5870_,
		_w5904_
	);
	LUT4 #(
		.INIT('h000e)
	) name5442 (
		_w528_,
		_w530_,
		_w533_,
		_w869_,
		_w5905_
	);
	LUT3 #(
		.INIT('ha8)
	) name5443 (
		_w3656_,
		_w5903_,
		_w5905_,
		_w5906_
	);
	LUT2 #(
		.INIT('h2)
	) name5444 (
		\P1_reg1_reg[0]/NET0131 ,
		_w2425_,
		_w5907_
	);
	LUT4 #(
		.INIT('h0c88)
	) name5445 (
		\P1_reg1_reg[0]/NET0131 ,
		_w1109_,
		_w1435_,
		_w2421_,
		_w5908_
	);
	LUT3 #(
		.INIT('h01)
	) name5446 (
		_w5907_,
		_w5908_,
		_w5906_,
		_w5909_
	);
	LUT4 #(
		.INIT('h1311)
	) name5447 (
		_w526_,
		_w5902_,
		_w5904_,
		_w5909_,
		_w5910_
	);
	LUT3 #(
		.INIT('hce)
	) name5448 (
		\P1_state_reg[0]/NET0131 ,
		_w5901_,
		_w5910_,
		_w5911_
	);
	LUT2 #(
		.INIT('h8)
	) name5449 (
		\P1_datao_reg[30]/NET0131 ,
		\si[30]_pad ,
		_w5912_
	);
	LUT2 #(
		.INIT('h1)
	) name5450 (
		\P1_datao_reg[30]/NET0131 ,
		\si[30]_pad ,
		_w5913_
	);
	LUT4 #(
		.INIT('hfac8)
	) name5451 (
		\P1_datao_reg[28]/NET0131 ,
		\P1_datao_reg[29]/NET0131 ,
		\si[28]_pad ,
		\si[29]_pad ,
		_w5914_
	);
	LUT2 #(
		.INIT('h8)
	) name5452 (
		_w2011_,
		_w5914_,
		_w5915_
	);
	LUT4 #(
		.INIT('h8000)
	) name5453 (
		_w1875_,
		_w1913_,
		_w1946_,
		_w1978_,
		_w5916_
	);
	LUT2 #(
		.INIT('h8)
	) name5454 (
		_w5915_,
		_w5916_,
		_w5917_
	);
	LUT4 #(
		.INIT('h7300)
	) name5455 (
		_w1825_,
		_w1912_,
		_w1914_,
		_w1979_,
		_w5918_
	);
	LUT4 #(
		.INIT('h010f)
	) name5456 (
		_w2010_,
		_w2014_,
		_w2608_,
		_w5914_,
		_w5919_
	);
	LUT4 #(
		.INIT('h3b00)
	) name5457 (
		_w1982_,
		_w5915_,
		_w5918_,
		_w5919_,
		_w5920_
	);
	LUT3 #(
		.INIT('h70)
	) name5458 (
		_w1827_,
		_w5917_,
		_w5920_,
		_w5921_
	);
	LUT4 #(
		.INIT('h9565)
	) name5459 (
		\P1_datao_reg[30]/NET0131 ,
		\si[30]_pad ,
		_w542_,
		_w5921_,
		_w5922_
	);
	LUT3 #(
		.INIT('h04)
	) name5460 (
		_w1509_,
		_w2920_,
		_w5922_,
		_w5923_
	);
	LUT3 #(
		.INIT('h70)
	) name5461 (
		_w2051_,
		_w2052_,
		_w2081_,
		_w5924_
	);
	LUT4 #(
		.INIT('h0200)
	) name5462 (
		_w2272_,
		_w2604_,
		_w2605_,
		_w5924_,
		_w5925_
	);
	LUT4 #(
		.INIT('h00fe)
	) name5463 (
		_w1491_,
		_w1493_,
		_w1496_,
		_w5815_,
		_w5926_
	);
	LUT4 #(
		.INIT('hf7bf)
	) name5464 (
		_w1811_,
		_w2033_,
		_w2035_,
		_w2036_,
		_w5927_
	);
	LUT4 #(
		.INIT('h001f)
	) name5465 (
		_w1491_,
		_w1493_,
		_w1496_,
		_w5927_,
		_w5928_
	);
	LUT3 #(
		.INIT('h02)
	) name5466 (
		_w4166_,
		_w5928_,
		_w5926_,
		_w5929_
	);
	LUT3 #(
		.INIT('h2a)
	) name5467 (
		\P2_reg0_reg[30]/NET0131 ,
		_w2635_,
		_w5929_,
		_w5930_
	);
	LUT4 #(
		.INIT('hffa8)
	) name5468 (
		_w4166_,
		_w5923_,
		_w5925_,
		_w5930_,
		_w5931_
	);
	LUT4 #(
		.INIT('hfac8)
	) name5469 (
		\P1_datao_reg[29]/NET0131 ,
		\P1_datao_reg[30]/NET0131 ,
		\si[29]_pad ,
		\si[30]_pad ,
		_w5932_
	);
	LUT2 #(
		.INIT('h8)
	) name5470 (
		_w2613_,
		_w5932_,
		_w5933_
	);
	LUT4 #(
		.INIT('h8000)
	) name5471 (
		_w1929_,
		_w1964_,
		_w2613_,
		_w5932_,
		_w5934_
	);
	LUT4 #(
		.INIT('h7300)
	) name5472 (
		_w1804_,
		_w1899_,
		_w1900_,
		_w1968_,
		_w5935_
	);
	LUT4 #(
		.INIT('h0b0a)
	) name5473 (
		_w2608_,
		_w2609_,
		_w5913_,
		_w5914_,
		_w5936_
	);
	LUT2 #(
		.INIT('h1)
	) name5474 (
		_w5912_,
		_w5936_,
		_w5937_
	);
	LUT4 #(
		.INIT('h3b00)
	) name5475 (
		_w1966_,
		_w5933_,
		_w5935_,
		_w5937_,
		_w5938_
	);
	LUT4 #(
		.INIT('hbf00)
	) name5476 (
		_w1710_,
		_w1896_,
		_w5934_,
		_w5938_,
		_w5939_
	);
	LUT4 #(
		.INIT('h6a9a)
	) name5477 (
		\P1_datao_reg[31]/NET0131 ,
		\si[31]_pad ,
		_w542_,
		_w5939_,
		_w5940_
	);
	LUT2 #(
		.INIT('h4)
	) name5478 (
		_w1509_,
		_w5940_,
		_w5941_
	);
	LUT4 #(
		.INIT('h4000)
	) name5479 (
		_w1509_,
		_w2084_,
		_w2277_,
		_w5940_,
		_w5942_
	);
	LUT3 #(
		.INIT('h2a)
	) name5480 (
		\P2_reg0_reg[31]/NET0131 ,
		_w2635_,
		_w5929_,
		_w5943_
	);
	LUT4 #(
		.INIT('hffa8)
	) name5481 (
		_w4166_,
		_w5925_,
		_w5942_,
		_w5943_,
		_w5944_
	);
	LUT3 #(
		.INIT('h04)
	) name5482 (
		_w1509_,
		_w2963_,
		_w5922_,
		_w5945_
	);
	LUT4 #(
		.INIT('h0200)
	) name5483 (
		_w1497_,
		_w2604_,
		_w2605_,
		_w5924_,
		_w5946_
	);
	LUT4 #(
		.INIT('hf100)
	) name5484 (
		_w1491_,
		_w1493_,
		_w1496_,
		_w5830_,
		_w5947_
	);
	LUT4 #(
		.INIT('hfbbf)
	) name5485 (
		_w1811_,
		_w2033_,
		_w2035_,
		_w2036_,
		_w5948_
	);
	LUT4 #(
		.INIT('h00ef)
	) name5486 (
		_w1491_,
		_w1493_,
		_w1496_,
		_w5948_,
		_w5949_
	);
	LUT3 #(
		.INIT('h02)
	) name5487 (
		_w4166_,
		_w5949_,
		_w5947_,
		_w5950_
	);
	LUT3 #(
		.INIT('h2a)
	) name5488 (
		\P2_reg1_reg[30]/NET0131 ,
		_w2661_,
		_w5950_,
		_w5951_
	);
	LUT4 #(
		.INIT('hffa8)
	) name5489 (
		_w4166_,
		_w5945_,
		_w5946_,
		_w5951_,
		_w5952_
	);
	LUT3 #(
		.INIT('h40)
	) name5490 (
		_w1509_,
		_w2963_,
		_w5940_,
		_w5953_
	);
	LUT3 #(
		.INIT('h2a)
	) name5491 (
		\P2_reg1_reg[31]/NET0131 ,
		_w2661_,
		_w5950_,
		_w5954_
	);
	LUT4 #(
		.INIT('hffa8)
	) name5492 (
		_w4166_,
		_w5946_,
		_w5953_,
		_w5954_,
		_w5955_
	);
	LUT4 #(
		.INIT('h00f1)
	) name5493 (
		_w1491_,
		_w1493_,
		_w1496_,
		_w5948_,
		_w5956_
	);
	LUT4 #(
		.INIT('hef00)
	) name5494 (
		_w1491_,
		_w1493_,
		_w1496_,
		_w5830_,
		_w5957_
	);
	LUT3 #(
		.INIT('h08)
	) name5495 (
		\P1_state_reg[0]/NET0131 ,
		_w1489_,
		_w2086_,
		_w5958_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name5496 (
		\P2_reg2_reg[30]/NET0131 ,
		_w5957_,
		_w5956_,
		_w5958_,
		_w5959_
	);
	LUT4 #(
		.INIT('h0200)
	) name5497 (
		_w2039_,
		_w2604_,
		_w2605_,
		_w5924_,
		_w5960_
	);
	LUT3 #(
		.INIT('ha8)
	) name5498 (
		_w1497_,
		_w1509_,
		_w5922_,
		_w5961_
	);
	LUT4 #(
		.INIT('h5455)
	) name5499 (
		\P2_reg2_reg[30]/NET0131 ,
		_w1491_,
		_w1493_,
		_w1496_,
		_w5962_
	);
	LUT2 #(
		.INIT('h2)
	) name5500 (
		_w2084_,
		_w5962_,
		_w5963_
	);
	LUT2 #(
		.INIT('h4)
	) name5501 (
		_w5961_,
		_w5963_,
		_w5964_
	);
	LUT4 #(
		.INIT('hccc8)
	) name5502 (
		_w2677_,
		_w4166_,
		_w5960_,
		_w5964_,
		_w5965_
	);
	LUT2 #(
		.INIT('he)
	) name5503 (
		_w5959_,
		_w5965_,
		_w5966_
	);
	LUT4 #(
		.INIT('h2000)
	) name5504 (
		_w1497_,
		_w1509_,
		_w2084_,
		_w5940_,
		_w5967_
	);
	LUT4 #(
		.INIT('hccc8)
	) name5505 (
		_w2677_,
		_w4166_,
		_w5960_,
		_w5967_,
		_w5968_
	);
	LUT4 #(
		.INIT('h0100)
	) name5506 (
		_w2087_,
		_w5957_,
		_w5956_,
		_w5958_,
		_w5969_
	);
	LUT2 #(
		.INIT('h2)
	) name5507 (
		\P2_reg2_reg[31]/NET0131 ,
		_w5969_,
		_w5970_
	);
	LUT2 #(
		.INIT('he)
	) name5508 (
		_w5968_,
		_w5970_,
		_w5971_
	);
	LUT2 #(
		.INIT('h8)
	) name5509 (
		\P1_state_reg[0]/NET0131 ,
		_w540_,
		_w5972_
	);
	LUT3 #(
		.INIT('hf1)
	) name5510 (
		\P1_state_reg[0]/NET0131 ,
		_w1033_,
		_w5972_,
		_w5973_
	);
	LUT4 #(
		.INIT('h2228)
	) name5511 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[25]/NET0131 ,
		_w1476_,
		_w1480_,
		_w5974_
	);
	LUT4 #(
		.INIT('hff54)
	) name5512 (
		\P1_state_reg[0]/NET0131 ,
		_w1926_,
		_w1935_,
		_w5974_,
		_w5975_
	);
	LUT4 #(
		.INIT('h8828)
	) name5513 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[27]/NET0131 ,
		\P2_IR_reg[31]/NET0131 ,
		_w1504_,
		_w5976_
	);
	LUT3 #(
		.INIT('hf1)
	) name5514 (
		\P1_state_reg[0]/NET0131 ,
		_w1970_,
		_w5976_,
		_w5977_
	);
	LUT3 #(
		.INIT('h48)
	) name5515 (
		\P1_IR_reg[25]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w521_,
		_w5978_
	);
	LUT3 #(
		.INIT('hf1)
	) name5516 (
		\P1_state_reg[0]/NET0131 ,
		_w968_,
		_w5978_,
		_w5979_
	);
	LUT4 #(
		.INIT('h8884)
	) name5517 (
		\P1_IR_reg[26]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w513_,
		_w516_,
		_w5980_
	);
	LUT4 #(
		.INIT('h00fe)
	) name5518 (
		\P1_state_reg[0]/NET0131 ,
		_w980_,
		_w997_,
		_w5980_,
		_w5981_
	);
	LUT4 #(
		.INIT('h2228)
	) name5519 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[26]/NET0131 ,
		_w479_,
		_w1484_,
		_w5982_
	);
	LUT3 #(
		.INIT('hf1)
	) name5520 (
		\P1_state_reg[0]/NET0131 ,
		_w1984_,
		_w5982_,
		_w5983_
	);
	LUT3 #(
		.INIT('h20)
	) name5521 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[30]/NET0131 ,
		\P2_IR_reg[31]/NET0131 ,
		_w5984_
	);
	LUT2 #(
		.INIT('h8)
	) name5522 (
		_w485_,
		_w5984_,
		_w5985_
	);
	LUT2 #(
		.INIT('h8)
	) name5523 (
		_w1504_,
		_w5985_,
		_w5986_
	);
	LUT3 #(
		.INIT('hf4)
	) name5524 (
		\P1_state_reg[0]/NET0131 ,
		_w5940_,
		_w5986_,
		_w5987_
	);
	LUT4 #(
		.INIT('h2228)
	) name5525 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[10]/NET0131 ,
		_w1654_,
		_w1655_,
		_w5988_
	);
	LUT3 #(
		.INIT('hf1)
	) name5526 (
		\P1_state_reg[0]/NET0131 ,
		_w1653_,
		_w5988_,
		_w5989_
	);
	LUT4 #(
		.INIT('h8828)
	) name5527 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[11]/NET0131 ,
		\P2_IR_reg[31]/NET0131 ,
		_w476_,
		_w5990_
	);
	LUT4 #(
		.INIT('hff54)
	) name5528 (
		\P1_state_reg[0]/NET0131 ,
		_w1621_,
		_w1637_,
		_w5990_,
		_w5991_
	);
	LUT2 #(
		.INIT('h8)
	) name5529 (
		\P1_state_reg[0]/NET0131 ,
		_w1744_,
		_w5992_
	);
	LUT4 #(
		.INIT('hff54)
	) name5530 (
		\P1_state_reg[0]/NET0131 ,
		_w1737_,
		_w1743_,
		_w5992_,
		_w5993_
	);
	LUT2 #(
		.INIT('h8)
	) name5531 (
		\P1_state_reg[0]/NET0131 ,
		_w1759_,
		_w5994_
	);
	LUT4 #(
		.INIT('hff54)
	) name5532 (
		\P1_state_reg[0]/NET0131 ,
		_w1753_,
		_w1758_,
		_w5994_,
		_w5995_
	);
	LUT2 #(
		.INIT('h2)
	) name5533 (
		\P1_state_reg[0]/NET0131 ,
		_w1728_,
		_w5996_
	);
	LUT3 #(
		.INIT('hf1)
	) name5534 (
		\P1_state_reg[0]/NET0131 ,
		_w1727_,
		_w5996_,
		_w5997_
	);
	LUT3 #(
		.INIT('h82)
	) name5535 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[15]/NET0131 ,
		_w1712_,
		_w5998_
	);
	LUT3 #(
		.INIT('hf1)
	) name5536 (
		\P1_state_reg[0]/NET0131 ,
		_w1711_,
		_w5998_,
		_w5999_
	);
	LUT3 #(
		.INIT('h82)
	) name5537 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[16]/NET0131 ,
		_w1792_,
		_w6000_
	);
	LUT3 #(
		.INIT('hf1)
	) name5538 (
		\P1_state_reg[0]/NET0131 ,
		_w1790_,
		_w6000_,
		_w6001_
	);
	LUT3 #(
		.INIT('h82)
	) name5539 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[17]/NET0131 ,
		_w1773_,
		_w6002_
	);
	LUT3 #(
		.INIT('hf1)
	) name5540 (
		\P1_state_reg[0]/NET0131 ,
		_w1771_,
		_w6002_,
		_w6003_
	);
	LUT3 #(
		.INIT('h82)
	) name5541 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[18]/NET0131 ,
		_w1830_,
		_w6004_
	);
	LUT4 #(
		.INIT('hff54)
	) name5542 (
		\P1_state_reg[0]/NET0131 ,
		_w1822_,
		_w1828_,
		_w6004_,
		_w6005_
	);
	LUT3 #(
		.INIT('h82)
	) name5543 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[19]/NET0131 ,
		_w1810_,
		_w6006_
	);
	LUT4 #(
		.INIT('hff54)
	) name5544 (
		\P1_state_reg[0]/NET0131 ,
		_w1797_,
		_w1808_,
		_w6006_,
		_w6007_
	);
	LUT4 #(
		.INIT('h28a0)
	) name5545 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[0]/NET0131 ,
		\P2_IR_reg[1]/NET0131 ,
		\P2_IR_reg[31]/NET0131 ,
		_w6008_
	);
	LUT3 #(
		.INIT('hf4)
	) name5546 (
		\P1_state_reg[0]/NET0131 ,
		_w1572_,
		_w6008_,
		_w6009_
	);
	LUT4 #(
		.INIT('h8828)
	) name5547 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[20]/NET0131 ,
		\P2_IR_reg[31]/NET0131 ,
		_w2030_,
		_w6010_
	);
	LUT4 #(
		.INIT('hff54)
	) name5548 (
		\P1_state_reg[0]/NET0131 ,
		_w1858_,
		_w1865_,
		_w6010_,
		_w6011_
	);
	LUT4 #(
		.INIT('h8882)
	) name5549 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[21]/NET0131 ,
		_w2031_,
		_w2034_,
		_w6012_
	);
	LUT3 #(
		.INIT('h0b)
	) name5550 (
		\P1_state_reg[0]/NET0131 ,
		_w1882_,
		_w6012_,
		_w6013_
	);
	LUT4 #(
		.INIT('h8882)
	) name5551 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[22]/NET0131 ,
		_w2031_,
		_w2032_,
		_w6014_
	);
	LUT3 #(
		.INIT('h0b)
	) name5552 (
		\P1_state_reg[0]/NET0131 ,
		_w1916_,
		_w6014_,
		_w6015_
	);
	LUT3 #(
		.INIT('h23)
	) name5553 (
		\P1_state_reg[0]/NET0131 ,
		_w1478_,
		_w1903_,
		_w6016_
	);
	LUT3 #(
		.INIT('h82)
	) name5554 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[24]/NET0131 ,
		_w1482_,
		_w6017_
	);
	LUT3 #(
		.INIT('hf1)
	) name5555 (
		\P1_state_reg[0]/NET0131 ,
		_w1953_,
		_w6017_,
		_w6018_
	);
	LUT4 #(
		.INIT('h2228)
	) name5556 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[28]/NET0131 ,
		_w1484_,
		_w1507_,
		_w6019_
	);
	LUT3 #(
		.INIT('hf1)
	) name5557 (
		\P1_state_reg[0]/NET0131 ,
		_w2017_,
		_w6019_,
		_w6020_
	);
	LUT4 #(
		.INIT('h2228)
	) name5558 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[29]/NET0131 ,
		_w489_,
		_w493_,
		_w6021_
	);
	LUT3 #(
		.INIT('hf1)
	) name5559 (
		\P1_state_reg[0]/NET0131 ,
		_w2616_,
		_w6021_,
		_w6022_
	);
	LUT2 #(
		.INIT('h2)
	) name5560 (
		\P1_state_reg[0]/NET0131 ,
		_w1561_,
		_w6023_
	);
	LUT3 #(
		.INIT('hf4)
	) name5561 (
		\P1_state_reg[0]/NET0131 ,
		_w1563_,
		_w6023_,
		_w6024_
	);
	LUT4 #(
		.INIT('h2228)
	) name5562 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[30]/NET0131 ,
		_w479_,
		_w487_,
		_w6025_
	);
	LUT3 #(
		.INIT('hf1)
	) name5563 (
		\P1_state_reg[0]/NET0131 ,
		_w5922_,
		_w6025_,
		_w6026_
	);
	LUT3 #(
		.INIT('h28)
	) name5564 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[3]/NET0131 ,
		_w1553_,
		_w6027_
	);
	LUT3 #(
		.INIT('hf1)
	) name5565 (
		\P1_state_reg[0]/NET0131 ,
		_w1552_,
		_w6027_,
		_w6028_
	);
	LUT4 #(
		.INIT('ha028)
	) name5566 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[31]/NET0131 ,
		\P2_IR_reg[4]/NET0131 ,
		_w472_,
		_w6029_
	);
	LUT3 #(
		.INIT('hf4)
	) name5567 (
		\P1_state_reg[0]/NET0131 ,
		_w1603_,
		_w6029_,
		_w6030_
	);
	LUT2 #(
		.INIT('h2)
	) name5568 (
		\P1_state_reg[0]/NET0131 ,
		_w1592_,
		_w6031_
	);
	LUT4 #(
		.INIT('hff54)
	) name5569 (
		\P1_state_reg[0]/NET0131 ,
		_w1588_,
		_w1590_,
		_w6031_,
		_w6032_
	);
	LUT3 #(
		.INIT('h28)
	) name5570 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[6]/NET0131 ,
		_w1510_,
		_w6033_
	);
	LUT3 #(
		.INIT('hf4)
	) name5571 (
		\P1_state_reg[0]/NET0131 ,
		_w1526_,
		_w6033_,
		_w6034_
	);
	LUT4 #(
		.INIT('h2228)
	) name5572 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[7]/NET0131 ,
		_w1510_,
		_w1543_,
		_w6035_
	);
	LUT3 #(
		.INIT('hf1)
	) name5573 (
		\P1_state_reg[0]/NET0131 ,
		_w1542_,
		_w6035_,
		_w6036_
	);
	LUT4 #(
		.INIT('ha028)
	) name5574 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[31]/NET0131 ,
		\P2_IR_reg[8]/NET0131 ,
		_w474_,
		_w6037_
	);
	LUT3 #(
		.INIT('hf1)
	) name5575 (
		\P1_state_reg[0]/NET0131 ,
		_w1681_,
		_w6037_,
		_w6038_
	);
	LUT4 #(
		.INIT('h2228)
	) name5576 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[9]/NET0131 ,
		_w1654_,
		_w1669_,
		_w6039_
	);
	LUT3 #(
		.INIT('hf1)
	) name5577 (
		\P1_state_reg[0]/NET0131 ,
		_w1668_,
		_w6039_,
		_w6040_
	);
	LUT4 #(
		.INIT('ha060)
	) name5578 (
		\P1_IR_reg[10]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w503_,
		_w6041_
	);
	LUT4 #(
		.INIT('hff54)
	) name5579 (
		\P1_state_reg[0]/NET0131 ,
		_w821_,
		_w823_,
		_w6041_,
		_w6042_
	);
	LUT2 #(
		.INIT('h8)
	) name5580 (
		\P1_state_reg[0]/NET0131 ,
		_w802_,
		_w6043_
	);
	LUT3 #(
		.INIT('hf1)
	) name5581 (
		\P1_state_reg[0]/NET0131 ,
		_w801_,
		_w6043_,
		_w6044_
	);
	LUT2 #(
		.INIT('h8)
	) name5582 (
		\P1_state_reg[0]/NET0131 ,
		_w812_,
		_w6045_
	);
	LUT3 #(
		.INIT('hf1)
	) name5583 (
		\P1_state_reg[0]/NET0131 ,
		_w810_,
		_w6045_,
		_w6046_
	);
	LUT2 #(
		.INIT('h8)
	) name5584 (
		\P1_state_reg[0]/NET0131 ,
		_w756_,
		_w6047_
	);
	LUT3 #(
		.INIT('hf1)
	) name5585 (
		\P1_state_reg[0]/NET0131 ,
		_w754_,
		_w6047_,
		_w6048_
	);
	LUT2 #(
		.INIT('h2)
	) name5586 (
		\P1_state_reg[0]/NET0131 ,
		_w765_,
		_w6049_
	);
	LUT3 #(
		.INIT('hf1)
	) name5587 (
		\P1_state_reg[0]/NET0131 ,
		_w764_,
		_w6049_,
		_w6050_
	);
	LUT3 #(
		.INIT('h48)
	) name5588 (
		\P1_IR_reg[15]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w777_,
		_w6051_
	);
	LUT4 #(
		.INIT('hff54)
	) name5589 (
		\P1_state_reg[0]/NET0131 ,
		_w774_,
		_w776_,
		_w6051_,
		_w6052_
	);
	LUT4 #(
		.INIT('ha060)
	) name5590 (
		\P1_IR_reg[16]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w648_,
		_w6053_
	);
	LUT4 #(
		.INIT('hff54)
	) name5591 (
		\P1_state_reg[0]/NET0131 ,
		_w781_,
		_w783_,
		_w6053_,
		_w6054_
	);
	LUT2 #(
		.INIT('h8)
	) name5592 (
		\P1_state_reg[0]/NET0131 ,
		_w715_,
		_w6055_
	);
	LUT4 #(
		.INIT('hff54)
	) name5593 (
		\P1_state_reg[0]/NET0131 ,
		_w710_,
		_w714_,
		_w6055_,
		_w6056_
	);
	LUT4 #(
		.INIT('ha060)
	) name5594 (
		\P1_IR_reg[18]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w649_,
		_w6057_
	);
	LUT3 #(
		.INIT('hf1)
	) name5595 (
		\P1_state_reg[0]/NET0131 ,
		_w735_,
		_w6057_,
		_w6058_
	);
	LUT4 #(
		.INIT('h4448)
	) name5596 (
		\P1_IR_reg[19]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w650_,
		_w651_,
		_w6059_
	);
	LUT3 #(
		.INIT('hf1)
	) name5597 (
		\P1_state_reg[0]/NET0131 ,
		_w673_,
		_w6059_,
		_w6060_
	);
	LUT4 #(
		.INIT('h6c00)
	) name5598 (
		\P1_IR_reg[0]/NET0131 ,
		\P1_IR_reg[1]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w6061_
	);
	LUT3 #(
		.INIT('hf4)
	) name5599 (
		\P1_state_reg[0]/NET0131 ,
		_w860_,
		_w6061_,
		_w6062_
	);
	LUT4 #(
		.INIT('ha060)
	) name5600 (
		\P1_IR_reg[20]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w1105_,
		_w6063_
	);
	LUT3 #(
		.INIT('hf1)
	) name5601 (
		\P1_state_reg[0]/NET0131 ,
		_w701_,
		_w6063_,
		_w6064_
	);
	LUT2 #(
		.INIT('h2)
	) name5602 (
		\P1_state_reg[0]/NET0131 ,
		_w1106_,
		_w6065_
	);
	LUT3 #(
		.INIT('h0b)
	) name5603 (
		\P1_state_reg[0]/NET0131 ,
		_w1073_,
		_w6065_,
		_w6066_
	);
	LUT3 #(
		.INIT('h48)
	) name5604 (
		\P1_IR_reg[22]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w513_,
		_w6067_
	);
	LUT4 #(
		.INIT('hff54)
	) name5605 (
		\P1_state_reg[0]/NET0131 ,
		_w1062_,
		_w1065_,
		_w6067_,
		_w6068_
	);
	LUT3 #(
		.INIT('hf1)
	) name5606 (
		\P1_state_reg[0]/NET0131 ,
		_w1046_,
		_w1294_,
		_w6069_
	);
	LUT4 #(
		.INIT('h8884)
	) name5607 (
		\P1_IR_reg[24]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w513_,
		_w518_,
		_w6070_
	);
	LUT3 #(
		.INIT('h0b)
	) name5608 (
		\P1_state_reg[0]/NET0131 ,
		_w1054_,
		_w6070_,
		_w6071_
	);
	LUT4 #(
		.INIT('h4448)
	) name5609 (
		\P1_IR_reg[28]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w513_,
		_w536_,
		_w6072_
	);
	LUT4 #(
		.INIT('hff54)
	) name5610 (
		\P1_state_reg[0]/NET0131 ,
		_w1008_,
		_w1017_,
		_w6072_,
		_w6073_
	);
	LUT4 #(
		.INIT('h8884)
	) name5611 (
		\P1_IR_reg[29]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w521_,
		_w626_,
		_w6074_
	);
	LUT4 #(
		.INIT('h00fe)
	) name5612 (
		\P1_state_reg[0]/NET0131 ,
		_w543_,
		_w620_,
		_w6074_,
		_w6075_
	);
	LUT2 #(
		.INIT('h8)
	) name5613 (
		\P1_state_reg[0]/NET0131 ,
		_w852_,
		_w6076_
	);
	LUT3 #(
		.INIT('hf1)
	) name5614 (
		\P1_state_reg[0]/NET0131 ,
		_w851_,
		_w6076_,
		_w6077_
	);
	LUT4 #(
		.INIT('h4448)
	) name5615 (
		\P1_IR_reg[30]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w513_,
		_w623_,
		_w6078_
	);
	LUT3 #(
		.INIT('hf1)
	) name5616 (
		\P1_state_reg[0]/NET0131 ,
		_w1311_,
		_w6078_,
		_w6079_
	);
	LUT3 #(
		.INIT('h40)
	) name5617 (
		\P1_IR_reg[30]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w6080_
	);
	LUT3 #(
		.INIT('h80)
	) name5618 (
		_w538_,
		_w622_,
		_w6080_,
		_w6081_
	);
	LUT2 #(
		.INIT('h8)
	) name5619 (
		_w509_,
		_w6081_,
		_w6082_
	);
	LUT4 #(
		.INIT('hff14)
	) name5620 (
		\P1_state_reg[0]/NET0131 ,
		\P2_datao_reg[31]/NET0131 ,
		_w1303_,
		_w6082_,
		_w6083_
	);
	LUT3 #(
		.INIT('h48)
	) name5621 (
		\P1_IR_reg[3]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w878_,
		_w6084_
	);
	LUT3 #(
		.INIT('hf4)
	) name5622 (
		\P1_state_reg[0]/NET0131 ,
		_w880_,
		_w6084_,
		_w6085_
	);
	LUT4 #(
		.INIT('hc060)
	) name5623 (
		\P1_IR_reg[31]/NET0131 ,
		\P1_IR_reg[4]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w500_,
		_w6086_
	);
	LUT4 #(
		.INIT('hff01)
	) name5624 (
		\P1_state_reg[0]/NET0131 ,
		_w890_,
		_w892_,
		_w6086_,
		_w6087_
	);
	LUT2 #(
		.INIT('h8)
	) name5625 (
		\P1_state_reg[0]/NET0131 ,
		_w937_,
		_w6088_
	);
	LUT3 #(
		.INIT('hf1)
	) name5626 (
		\P1_state_reg[0]/NET0131 ,
		_w936_,
		_w6088_,
		_w6089_
	);
	LUT3 #(
		.INIT('h48)
	) name5627 (
		\P1_IR_reg[6]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w915_,
		_w6090_
	);
	LUT3 #(
		.INIT('hf4)
	) name5628 (
		\P1_state_reg[0]/NET0131 ,
		_w928_,
		_w6090_,
		_w6091_
	);
	LUT4 #(
		.INIT('h4448)
	) name5629 (
		\P1_IR_reg[7]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w915_,
		_w916_,
		_w6092_
	);
	LUT3 #(
		.INIT('hf1)
	) name5630 (
		\P1_state_reg[0]/NET0131 ,
		_w914_,
		_w6092_,
		_w6093_
	);
	LUT4 #(
		.INIT('hc060)
	) name5631 (
		\P1_IR_reg[31]/NET0131 ,
		\P1_IR_reg[8]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w839_,
		_w6094_
	);
	LUT3 #(
		.INIT('hf1)
	) name5632 (
		\P1_state_reg[0]/NET0131 ,
		_w905_,
		_w6094_,
		_w6095_
	);
	LUT2 #(
		.INIT('h8)
	) name5633 (
		\P1_state_reg[0]/NET0131 ,
		_w840_,
		_w6096_
	);
	LUT4 #(
		.INIT('hff54)
	) name5634 (
		\P1_state_reg[0]/NET0131 ,
		_w835_,
		_w837_,
		_w6096_,
		_w6097_
	);
	LUT3 #(
		.INIT('h21)
	) name5635 (
		\P2_IR_reg[18]/NET0131 ,
		\P2_reg1_reg[18]/NET0131 ,
		_w1830_,
		_w6098_
	);
	LUT3 #(
		.INIT('h48)
	) name5636 (
		\P2_IR_reg[18]/NET0131 ,
		\P2_reg1_reg[18]/NET0131 ,
		_w1830_,
		_w6099_
	);
	LUT3 #(
		.INIT('h96)
	) name5637 (
		\P2_IR_reg[18]/NET0131 ,
		\P2_reg1_reg[18]/NET0131 ,
		_w1830_,
		_w6100_
	);
	LUT3 #(
		.INIT('h48)
	) name5638 (
		\P2_IR_reg[17]/NET0131 ,
		\P2_reg1_reg[17]/NET0131 ,
		_w1773_,
		_w6101_
	);
	LUT3 #(
		.INIT('h48)
	) name5639 (
		\P2_IR_reg[16]/NET0131 ,
		\P2_reg1_reg[16]/NET0131 ,
		_w1792_,
		_w6102_
	);
	LUT3 #(
		.INIT('h48)
	) name5640 (
		\P2_IR_reg[15]/NET0131 ,
		\P2_reg1_reg[15]/NET0131 ,
		_w1712_,
		_w6103_
	);
	LUT3 #(
		.INIT('h21)
	) name5641 (
		\P2_IR_reg[15]/NET0131 ,
		\P2_reg1_reg[15]/NET0131 ,
		_w1712_,
		_w6104_
	);
	LUT2 #(
		.INIT('h1)
	) name5642 (
		\P2_reg1_reg[14]/NET0131 ,
		_w1728_,
		_w6105_
	);
	LUT2 #(
		.INIT('h1)
	) name5643 (
		_w6104_,
		_w6105_,
		_w6106_
	);
	LUT2 #(
		.INIT('h8)
	) name5644 (
		\P2_reg1_reg[14]/NET0131 ,
		_w1728_,
		_w6107_
	);
	LUT2 #(
		.INIT('h2)
	) name5645 (
		\P2_reg1_reg[13]/NET0131 ,
		_w1759_,
		_w6108_
	);
	LUT2 #(
		.INIT('h4)
	) name5646 (
		\P2_reg1_reg[12]/NET0131 ,
		_w1744_,
		_w6109_
	);
	LUT4 #(
		.INIT('h8caf)
	) name5647 (
		\P2_reg1_reg[12]/NET0131 ,
		\P2_reg1_reg[13]/NET0131 ,
		_w1744_,
		_w1759_,
		_w6110_
	);
	LUT2 #(
		.INIT('h2)
	) name5648 (
		\P2_reg1_reg[12]/NET0131 ,
		_w1744_,
		_w6111_
	);
	LUT4 #(
		.INIT('h5090)
	) name5649 (
		\P2_IR_reg[11]/NET0131 ,
		\P2_IR_reg[31]/NET0131 ,
		\P2_reg1_reg[11]/NET0131 ,
		_w476_,
		_w6112_
	);
	LUT4 #(
		.INIT('h8884)
	) name5650 (
		\P2_IR_reg[10]/NET0131 ,
		\P2_reg1_reg[10]/NET0131 ,
		_w1654_,
		_w1655_,
		_w6113_
	);
	LUT4 #(
		.INIT('h8884)
	) name5651 (
		\P2_IR_reg[9]/NET0131 ,
		\P2_reg1_reg[9]/NET0131 ,
		_w1654_,
		_w1669_,
		_w6114_
	);
	LUT4 #(
		.INIT('h1112)
	) name5652 (
		\P2_IR_reg[9]/NET0131 ,
		\P2_reg1_reg[9]/NET0131 ,
		_w1654_,
		_w1669_,
		_w6115_
	);
	LUT4 #(
		.INIT('h0c06)
	) name5653 (
		\P2_IR_reg[31]/NET0131 ,
		\P2_IR_reg[8]/NET0131 ,
		\P2_reg1_reg[8]/NET0131 ,
		_w474_,
		_w6116_
	);
	LUT2 #(
		.INIT('h1)
	) name5654 (
		_w6115_,
		_w6116_,
		_w6117_
	);
	LUT4 #(
		.INIT('h3090)
	) name5655 (
		\P2_IR_reg[31]/NET0131 ,
		\P2_IR_reg[8]/NET0131 ,
		\P2_reg1_reg[8]/NET0131 ,
		_w474_,
		_w6118_
	);
	LUT4 #(
		.INIT('h8884)
	) name5656 (
		\P2_IR_reg[7]/NET0131 ,
		\P2_reg1_reg[7]/NET0131 ,
		_w1510_,
		_w1543_,
		_w6119_
	);
	LUT4 #(
		.INIT('h1112)
	) name5657 (
		\P2_IR_reg[7]/NET0131 ,
		\P2_reg1_reg[7]/NET0131 ,
		_w1510_,
		_w1543_,
		_w6120_
	);
	LUT3 #(
		.INIT('h12)
	) name5658 (
		\P2_IR_reg[6]/NET0131 ,
		\P2_reg1_reg[6]/NET0131 ,
		_w1510_,
		_w6121_
	);
	LUT2 #(
		.INIT('h1)
	) name5659 (
		_w6120_,
		_w6121_,
		_w6122_
	);
	LUT3 #(
		.INIT('h84)
	) name5660 (
		\P2_IR_reg[6]/NET0131 ,
		\P2_reg1_reg[6]/NET0131 ,
		_w1510_,
		_w6123_
	);
	LUT2 #(
		.INIT('h1)
	) name5661 (
		\P2_reg1_reg[5]/NET0131 ,
		_w1592_,
		_w6124_
	);
	LUT2 #(
		.INIT('h8)
	) name5662 (
		\P2_reg1_reg[5]/NET0131 ,
		_w1592_,
		_w6125_
	);
	LUT4 #(
		.INIT('h3090)
	) name5663 (
		\P2_IR_reg[31]/NET0131 ,
		\P2_IR_reg[4]/NET0131 ,
		\P2_reg1_reg[4]/NET0131 ,
		_w472_,
		_w6126_
	);
	LUT4 #(
		.INIT('h0c06)
	) name5664 (
		\P2_IR_reg[31]/NET0131 ,
		\P2_IR_reg[4]/NET0131 ,
		\P2_reg1_reg[4]/NET0131 ,
		_w472_,
		_w6127_
	);
	LUT3 #(
		.INIT('h84)
	) name5665 (
		\P2_IR_reg[3]/NET0131 ,
		\P2_reg1_reg[3]/NET0131 ,
		_w1553_,
		_w6128_
	);
	LUT3 #(
		.INIT('h12)
	) name5666 (
		\P2_IR_reg[3]/NET0131 ,
		\P2_reg1_reg[3]/NET0131 ,
		_w1553_,
		_w6129_
	);
	LUT2 #(
		.INIT('h4)
	) name5667 (
		\P2_IR_reg[0]/NET0131 ,
		\P2_reg1_reg[0]/NET0131 ,
		_w6130_
	);
	LUT3 #(
		.INIT('he8)
	) name5668 (
		\P2_reg1_reg[1]/NET0131 ,
		_w1571_,
		_w6130_,
		_w6131_
	);
	LUT4 #(
		.INIT('h0e08)
	) name5669 (
		\P2_reg1_reg[2]/NET0131 ,
		_w1561_,
		_w6129_,
		_w6131_,
		_w6132_
	);
	LUT4 #(
		.INIT('h444d)
	) name5670 (
		\P2_reg1_reg[4]/NET0131 ,
		_w1601_,
		_w6128_,
		_w6132_,
		_w6133_
	);
	LUT4 #(
		.INIT('h0701)
	) name5671 (
		\P2_reg1_reg[5]/NET0131 ,
		_w1592_,
		_w6123_,
		_w6133_,
		_w6134_
	);
	LUT3 #(
		.INIT('h51)
	) name5672 (
		_w6119_,
		_w6122_,
		_w6134_,
		_w6135_
	);
	LUT4 #(
		.INIT('h1101)
	) name5673 (
		_w6118_,
		_w6119_,
		_w6122_,
		_w6134_,
		_w6136_
	);
	LUT4 #(
		.INIT('h1101)
	) name5674 (
		_w6113_,
		_w6114_,
		_w6117_,
		_w6136_,
		_w6137_
	);
	LUT4 #(
		.INIT('h0a06)
	) name5675 (
		\P2_IR_reg[11]/NET0131 ,
		\P2_IR_reg[31]/NET0131 ,
		\P2_reg1_reg[11]/NET0131 ,
		_w476_,
		_w6138_
	);
	LUT4 #(
		.INIT('h1112)
	) name5676 (
		\P2_IR_reg[10]/NET0131 ,
		\P2_reg1_reg[10]/NET0131 ,
		_w1654_,
		_w1655_,
		_w6139_
	);
	LUT2 #(
		.INIT('h1)
	) name5677 (
		_w6138_,
		_w6139_,
		_w6140_
	);
	LUT4 #(
		.INIT('h1011)
	) name5678 (
		_w6111_,
		_w6112_,
		_w6137_,
		_w6140_,
		_w6141_
	);
	LUT4 #(
		.INIT('h1101)
	) name5679 (
		_w6107_,
		_w6108_,
		_w6110_,
		_w6141_,
		_w6142_
	);
	LUT3 #(
		.INIT('h51)
	) name5680 (
		_w6103_,
		_w6106_,
		_w6142_,
		_w6143_
	);
	LUT4 #(
		.INIT('h1101)
	) name5681 (
		_w6102_,
		_w6103_,
		_w6106_,
		_w6142_,
		_w6144_
	);
	LUT3 #(
		.INIT('h21)
	) name5682 (
		\P2_IR_reg[17]/NET0131 ,
		\P2_reg1_reg[17]/NET0131 ,
		_w1773_,
		_w6145_
	);
	LUT3 #(
		.INIT('h21)
	) name5683 (
		\P2_IR_reg[16]/NET0131 ,
		\P2_reg1_reg[16]/NET0131 ,
		_w1792_,
		_w6146_
	);
	LUT2 #(
		.INIT('h1)
	) name5684 (
		_w6145_,
		_w6146_,
		_w6147_
	);
	LUT4 #(
		.INIT('h4544)
	) name5685 (
		_w6100_,
		_w6101_,
		_w6144_,
		_w6147_,
		_w6148_
	);
	LUT2 #(
		.INIT('h8)
	) name5686 (
		_w1505_,
		_w1508_,
		_w6149_
	);
	LUT4 #(
		.INIT('h2022)
	) name5687 (
		_w6100_,
		_w6101_,
		_w6144_,
		_w6147_,
		_w6150_
	);
	LUT3 #(
		.INIT('h02)
	) name5688 (
		_w6149_,
		_w6150_,
		_w6148_,
		_w6151_
	);
	LUT3 #(
		.INIT('h21)
	) name5689 (
		\P2_IR_reg[18]/NET0131 ,
		\P2_reg2_reg[18]/NET0131 ,
		_w1830_,
		_w6152_
	);
	LUT3 #(
		.INIT('h48)
	) name5690 (
		\P2_IR_reg[18]/NET0131 ,
		\P2_reg2_reg[18]/NET0131 ,
		_w1830_,
		_w6153_
	);
	LUT3 #(
		.INIT('h96)
	) name5691 (
		\P2_IR_reg[18]/NET0131 ,
		\P2_reg2_reg[18]/NET0131 ,
		_w1830_,
		_w6154_
	);
	LUT3 #(
		.INIT('h48)
	) name5692 (
		\P2_IR_reg[17]/NET0131 ,
		\P2_reg2_reg[17]/NET0131 ,
		_w1773_,
		_w6155_
	);
	LUT3 #(
		.INIT('h48)
	) name5693 (
		\P2_IR_reg[16]/NET0131 ,
		\P2_reg2_reg[16]/NET0131 ,
		_w1792_,
		_w6156_
	);
	LUT3 #(
		.INIT('h48)
	) name5694 (
		\P2_IR_reg[15]/NET0131 ,
		\P2_reg2_reg[15]/NET0131 ,
		_w1712_,
		_w6157_
	);
	LUT3 #(
		.INIT('h21)
	) name5695 (
		\P2_IR_reg[15]/NET0131 ,
		\P2_reg2_reg[15]/NET0131 ,
		_w1712_,
		_w6158_
	);
	LUT2 #(
		.INIT('h1)
	) name5696 (
		\P2_reg2_reg[14]/NET0131 ,
		_w1728_,
		_w6159_
	);
	LUT2 #(
		.INIT('h1)
	) name5697 (
		_w6158_,
		_w6159_,
		_w6160_
	);
	LUT2 #(
		.INIT('h8)
	) name5698 (
		\P2_reg2_reg[14]/NET0131 ,
		_w1728_,
		_w6161_
	);
	LUT2 #(
		.INIT('h2)
	) name5699 (
		\P2_reg2_reg[13]/NET0131 ,
		_w1759_,
		_w6162_
	);
	LUT2 #(
		.INIT('h4)
	) name5700 (
		\P2_reg2_reg[12]/NET0131 ,
		_w1744_,
		_w6163_
	);
	LUT4 #(
		.INIT('h8caf)
	) name5701 (
		\P2_reg2_reg[12]/NET0131 ,
		\P2_reg2_reg[13]/NET0131 ,
		_w1744_,
		_w1759_,
		_w6164_
	);
	LUT2 #(
		.INIT('h2)
	) name5702 (
		\P2_reg2_reg[12]/NET0131 ,
		_w1744_,
		_w6165_
	);
	LUT4 #(
		.INIT('h5090)
	) name5703 (
		\P2_IR_reg[11]/NET0131 ,
		\P2_IR_reg[31]/NET0131 ,
		\P2_reg2_reg[11]/NET0131 ,
		_w476_,
		_w6166_
	);
	LUT4 #(
		.INIT('h0a06)
	) name5704 (
		\P2_IR_reg[11]/NET0131 ,
		\P2_IR_reg[31]/NET0131 ,
		\P2_reg2_reg[11]/NET0131 ,
		_w476_,
		_w6167_
	);
	LUT4 #(
		.INIT('h1112)
	) name5705 (
		\P2_IR_reg[10]/NET0131 ,
		\P2_reg2_reg[10]/NET0131 ,
		_w1654_,
		_w1655_,
		_w6168_
	);
	LUT2 #(
		.INIT('h1)
	) name5706 (
		_w6167_,
		_w6168_,
		_w6169_
	);
	LUT4 #(
		.INIT('h8884)
	) name5707 (
		\P2_IR_reg[10]/NET0131 ,
		\P2_reg2_reg[10]/NET0131 ,
		_w1654_,
		_w1655_,
		_w6170_
	);
	LUT4 #(
		.INIT('h8884)
	) name5708 (
		\P2_IR_reg[9]/NET0131 ,
		\P2_reg2_reg[9]/NET0131 ,
		_w1654_,
		_w1669_,
		_w6171_
	);
	LUT4 #(
		.INIT('h1112)
	) name5709 (
		\P2_IR_reg[9]/NET0131 ,
		\P2_reg2_reg[9]/NET0131 ,
		_w1654_,
		_w1669_,
		_w6172_
	);
	LUT4 #(
		.INIT('h0c06)
	) name5710 (
		\P2_IR_reg[31]/NET0131 ,
		\P2_IR_reg[8]/NET0131 ,
		\P2_reg2_reg[8]/NET0131 ,
		_w474_,
		_w6173_
	);
	LUT2 #(
		.INIT('h1)
	) name5711 (
		_w6172_,
		_w6173_,
		_w6174_
	);
	LUT4 #(
		.INIT('h3090)
	) name5712 (
		\P2_IR_reg[31]/NET0131 ,
		\P2_IR_reg[8]/NET0131 ,
		\P2_reg2_reg[8]/NET0131 ,
		_w474_,
		_w6175_
	);
	LUT4 #(
		.INIT('h8884)
	) name5713 (
		\P2_IR_reg[7]/NET0131 ,
		\P2_reg2_reg[7]/NET0131 ,
		_w1510_,
		_w1543_,
		_w6176_
	);
	LUT4 #(
		.INIT('h1112)
	) name5714 (
		\P2_IR_reg[7]/NET0131 ,
		\P2_reg2_reg[7]/NET0131 ,
		_w1510_,
		_w1543_,
		_w6177_
	);
	LUT3 #(
		.INIT('h12)
	) name5715 (
		\P2_IR_reg[6]/NET0131 ,
		\P2_reg2_reg[6]/NET0131 ,
		_w1510_,
		_w6178_
	);
	LUT2 #(
		.INIT('h1)
	) name5716 (
		_w6177_,
		_w6178_,
		_w6179_
	);
	LUT3 #(
		.INIT('h84)
	) name5717 (
		\P2_IR_reg[6]/NET0131 ,
		\P2_reg2_reg[6]/NET0131 ,
		_w1510_,
		_w6180_
	);
	LUT2 #(
		.INIT('h1)
	) name5718 (
		\P2_reg2_reg[5]/NET0131 ,
		_w1592_,
		_w6181_
	);
	LUT2 #(
		.INIT('h8)
	) name5719 (
		\P2_reg2_reg[5]/NET0131 ,
		_w1592_,
		_w6182_
	);
	LUT3 #(
		.INIT('h84)
	) name5720 (
		\P2_IR_reg[3]/NET0131 ,
		\P2_reg2_reg[3]/NET0131 ,
		_w1553_,
		_w6183_
	);
	LUT3 #(
		.INIT('h12)
	) name5721 (
		\P2_IR_reg[3]/NET0131 ,
		\P2_reg2_reg[3]/NET0131 ,
		_w1553_,
		_w6184_
	);
	LUT2 #(
		.INIT('h4)
	) name5722 (
		\P2_IR_reg[0]/NET0131 ,
		\P2_reg2_reg[0]/NET0131 ,
		_w6185_
	);
	LUT3 #(
		.INIT('he8)
	) name5723 (
		\P2_reg2_reg[1]/NET0131 ,
		_w1571_,
		_w6185_,
		_w6186_
	);
	LUT4 #(
		.INIT('h0e08)
	) name5724 (
		\P2_reg2_reg[2]/NET0131 ,
		_w1561_,
		_w6184_,
		_w6186_,
		_w6187_
	);
	LUT4 #(
		.INIT('h444d)
	) name5725 (
		\P2_reg2_reg[4]/NET0131 ,
		_w1601_,
		_w6183_,
		_w6187_,
		_w6188_
	);
	LUT4 #(
		.INIT('h0701)
	) name5726 (
		\P2_reg2_reg[5]/NET0131 ,
		_w1592_,
		_w6180_,
		_w6188_,
		_w6189_
	);
	LUT4 #(
		.INIT('h1101)
	) name5727 (
		_w6175_,
		_w6176_,
		_w6179_,
		_w6189_,
		_w6190_
	);
	LUT3 #(
		.INIT('h51)
	) name5728 (
		_w6171_,
		_w6174_,
		_w6190_,
		_w6191_
	);
	LUT4 #(
		.INIT('h1101)
	) name5729 (
		_w6170_,
		_w6171_,
		_w6174_,
		_w6190_,
		_w6192_
	);
	LUT3 #(
		.INIT('h51)
	) name5730 (
		_w6166_,
		_w6169_,
		_w6192_,
		_w6193_
	);
	LUT4 #(
		.INIT('h1101)
	) name5731 (
		_w6165_,
		_w6166_,
		_w6169_,
		_w6192_,
		_w6194_
	);
	LUT3 #(
		.INIT('h51)
	) name5732 (
		_w6162_,
		_w6164_,
		_w6194_,
		_w6195_
	);
	LUT4 #(
		.INIT('h1101)
	) name5733 (
		_w6161_,
		_w6162_,
		_w6164_,
		_w6194_,
		_w6196_
	);
	LUT4 #(
		.INIT('h1101)
	) name5734 (
		_w6156_,
		_w6157_,
		_w6160_,
		_w6196_,
		_w6197_
	);
	LUT3 #(
		.INIT('h21)
	) name5735 (
		\P2_IR_reg[16]/NET0131 ,
		\P2_reg2_reg[16]/NET0131 ,
		_w1792_,
		_w6198_
	);
	LUT3 #(
		.INIT('h21)
	) name5736 (
		\P2_IR_reg[17]/NET0131 ,
		\P2_reg2_reg[17]/NET0131 ,
		_w1773_,
		_w6199_
	);
	LUT2 #(
		.INIT('h1)
	) name5737 (
		_w6198_,
		_w6199_,
		_w6200_
	);
	LUT3 #(
		.INIT('h45)
	) name5738 (
		_w6155_,
		_w6197_,
		_w6200_,
		_w6201_
	);
	LUT3 #(
		.INIT('ha8)
	) name5739 (
		_w1477_,
		_w1486_,
		_w2080_,
		_w6202_
	);
	LUT2 #(
		.INIT('h1)
	) name5740 (
		_w1505_,
		_w1508_,
		_w6203_
	);
	LUT4 #(
		.INIT('hf4f7)
	) name5741 (
		\P2_addr_reg[18]/NET0131 ,
		_w1505_,
		_w1508_,
		_w1831_,
		_w6204_
	);
	LUT4 #(
		.INIT('h5700)
	) name5742 (
		_w1477_,
		_w1486_,
		_w2080_,
		_w6204_,
		_w6205_
	);
	LUT4 #(
		.INIT('hd700)
	) name5743 (
		_w2041_,
		_w6154_,
		_w6201_,
		_w6205_,
		_w6206_
	);
	LUT2 #(
		.INIT('h2)
	) name5744 (
		\P2_IR_reg[0]/NET0131 ,
		\P2_reg1_reg[0]/NET0131 ,
		_w6207_
	);
	LUT3 #(
		.INIT('h8e)
	) name5745 (
		\P2_reg1_reg[1]/NET0131 ,
		_w1571_,
		_w6207_,
		_w6208_
	);
	LUT4 #(
		.INIT('h0107)
	) name5746 (
		\P2_reg1_reg[2]/NET0131 ,
		_w1561_,
		_w6128_,
		_w6208_,
		_w6209_
	);
	LUT3 #(
		.INIT('h0e)
	) name5747 (
		\P2_reg1_reg[5]/NET0131 ,
		_w1592_,
		_w6127_,
		_w6210_
	);
	LUT4 #(
		.INIT('hab00)
	) name5748 (
		_w6126_,
		_w6129_,
		_w6209_,
		_w6210_,
		_w6211_
	);
	LUT2 #(
		.INIT('h1)
	) name5749 (
		_w6123_,
		_w6125_,
		_w6212_
	);
	LUT4 #(
		.INIT('h1511)
	) name5750 (
		_w6119_,
		_w6122_,
		_w6211_,
		_w6212_,
		_w6213_
	);
	LUT4 #(
		.INIT('h1511)
	) name5751 (
		_w6114_,
		_w6117_,
		_w6118_,
		_w6213_,
		_w6214_
	);
	LUT4 #(
		.INIT('h020b)
	) name5752 (
		\P2_reg1_reg[10]/NET0131 ,
		_w1656_,
		_w6138_,
		_w6214_,
		_w6215_
	);
	LUT3 #(
		.INIT('h0d)
	) name5753 (
		\P2_reg1_reg[12]/NET0131 ,
		_w1744_,
		_w6112_,
		_w6216_
	);
	LUT4 #(
		.INIT('h3f15)
	) name5754 (
		\P2_reg1_reg[13]/NET0131 ,
		\P2_reg1_reg[14]/NET0131 ,
		_w1728_,
		_w1759_,
		_w6217_
	);
	LUT4 #(
		.INIT('h7500)
	) name5755 (
		_w6110_,
		_w6215_,
		_w6216_,
		_w6217_,
		_w6218_
	);
	LUT3 #(
		.INIT('h51)
	) name5756 (
		_w6103_,
		_w6106_,
		_w6218_,
		_w6219_
	);
	LUT4 #(
		.INIT('h4454)
	) name5757 (
		_w6146_,
		_w6103_,
		_w6106_,
		_w6218_,
		_w6220_
	);
	LUT2 #(
		.INIT('h1)
	) name5758 (
		_w6101_,
		_w6102_,
		_w6221_
	);
	LUT4 #(
		.INIT('h2022)
	) name5759 (
		_w6100_,
		_w6145_,
		_w6220_,
		_w6221_,
		_w6222_
	);
	LUT4 #(
		.INIT('h4544)
	) name5760 (
		_w6100_,
		_w6145_,
		_w6220_,
		_w6221_,
		_w6223_
	);
	LUT3 #(
		.INIT('h02)
	) name5761 (
		_w1509_,
		_w6223_,
		_w6222_,
		_w6224_
	);
	LUT2 #(
		.INIT('h2)
	) name5762 (
		\P2_IR_reg[0]/NET0131 ,
		\P2_reg2_reg[0]/NET0131 ,
		_w6225_
	);
	LUT3 #(
		.INIT('h8e)
	) name5763 (
		\P2_reg2_reg[1]/NET0131 ,
		_w1571_,
		_w6225_,
		_w6226_
	);
	LUT4 #(
		.INIT('h0107)
	) name5764 (
		\P2_reg2_reg[2]/NET0131 ,
		_w1561_,
		_w6183_,
		_w6226_,
		_w6227_
	);
	LUT4 #(
		.INIT('h222b)
	) name5765 (
		\P2_reg2_reg[4]/NET0131 ,
		_w1601_,
		_w6184_,
		_w6227_,
		_w6228_
	);
	LUT4 #(
		.INIT('h0107)
	) name5766 (
		\P2_reg2_reg[5]/NET0131 ,
		_w1592_,
		_w6180_,
		_w6228_,
		_w6229_
	);
	LUT3 #(
		.INIT('h51)
	) name5767 (
		_w6176_,
		_w6179_,
		_w6229_,
		_w6230_
	);
	LUT4 #(
		.INIT('h1101)
	) name5768 (
		_w6175_,
		_w6176_,
		_w6179_,
		_w6229_,
		_w6231_
	);
	LUT3 #(
		.INIT('h51)
	) name5769 (
		_w6171_,
		_w6174_,
		_w6231_,
		_w6232_
	);
	LUT4 #(
		.INIT('h88a8)
	) name5770 (
		_w6169_,
		_w6171_,
		_w6174_,
		_w6231_,
		_w6233_
	);
	LUT3 #(
		.INIT('h4d)
	) name5771 (
		\P2_reg2_reg[11]/NET0131 ,
		_w1639_,
		_w6170_,
		_w6234_
	);
	LUT4 #(
		.INIT('hf731)
	) name5772 (
		\P2_reg2_reg[12]/NET0131 ,
		\P2_reg2_reg[13]/NET0131 ,
		_w1744_,
		_w1759_,
		_w6235_
	);
	LUT4 #(
		.INIT('h7500)
	) name5773 (
		_w6164_,
		_w6233_,
		_w6234_,
		_w6235_,
		_w6236_
	);
	LUT3 #(
		.INIT('hb2)
	) name5774 (
		\P2_reg2_reg[15]/NET0131 ,
		_w1713_,
		_w6161_,
		_w6237_
	);
	LUT4 #(
		.INIT('h5504)
	) name5775 (
		_w6198_,
		_w6160_,
		_w6236_,
		_w6237_,
		_w6238_
	);
	LUT2 #(
		.INIT('h1)
	) name5776 (
		_w6155_,
		_w6156_,
		_w6239_
	);
	LUT3 #(
		.INIT('h45)
	) name5777 (
		_w6199_,
		_w6238_,
		_w6239_,
		_w6240_
	);
	LUT2 #(
		.INIT('h8)
	) name5778 (
		_w1508_,
		_w1831_,
		_w6241_
	);
	LUT2 #(
		.INIT('h2)
	) name5779 (
		_w1486_,
		_w6241_,
		_w6242_
	);
	LUT4 #(
		.INIT('hb700)
	) name5780 (
		_w6154_,
		_w6203_,
		_w6240_,
		_w6242_,
		_w6243_
	);
	LUT4 #(
		.INIT('h1555)
	) name5781 (
		\P2_addr_reg[18]/NET0131 ,
		_w1483_,
		_w1485_,
		_w1481_,
		_w6244_
	);
	LUT2 #(
		.INIT('h8)
	) name5782 (
		_w2080_,
		_w6244_,
		_w6245_
	);
	LUT4 #(
		.INIT('haa20)
	) name5783 (
		_w1477_,
		_w6224_,
		_w6243_,
		_w6245_,
		_w6246_
	);
	LUT4 #(
		.INIT('h008a)
	) name5784 (
		\P1_state_reg[0]/NET0131 ,
		_w6151_,
		_w6206_,
		_w6246_,
		_w6247_
	);
	LUT2 #(
		.INIT('he)
	) name5785 (
		_w2744_,
		_w6247_,
		_w6248_
	);
	LUT2 #(
		.INIT('h9)
	) name5786 (
		\P2_IR_reg[0]/NET0131 ,
		\P2_reg1_reg[0]/NET0131 ,
		_w6249_
	);
	LUT3 #(
		.INIT('h02)
	) name5787 (
		_w1505_,
		_w1508_,
		_w6249_,
		_w6250_
	);
	LUT2 #(
		.INIT('h9)
	) name5788 (
		\P2_IR_reg[0]/NET0131 ,
		\P2_reg2_reg[0]/NET0131 ,
		_w6251_
	);
	LUT3 #(
		.INIT('h01)
	) name5789 (
		_w1505_,
		_w1508_,
		_w6251_,
		_w6252_
	);
	LUT4 #(
		.INIT('h2228)
	) name5790 (
		\P2_IR_reg[0]/NET0131 ,
		\P2_IR_reg[28]/NET0131 ,
		_w1484_,
		_w1507_,
		_w6253_
	);
	LUT4 #(
		.INIT('h0080)
	) name5791 (
		_w1483_,
		_w1485_,
		_w1481_,
		_w6253_,
		_w6254_
	);
	LUT3 #(
		.INIT('h10)
	) name5792 (
		_w6252_,
		_w6250_,
		_w6254_,
		_w6255_
	);
	LUT4 #(
		.INIT('h1555)
	) name5793 (
		\P2_addr_reg[0]/NET0131 ,
		_w1483_,
		_w1485_,
		_w1481_,
		_w6256_
	);
	LUT2 #(
		.INIT('h8)
	) name5794 (
		_w2080_,
		_w6256_,
		_w6257_
	);
	LUT3 #(
		.INIT('ha8)
	) name5795 (
		_w1477_,
		_w6255_,
		_w6257_,
		_w6258_
	);
	LUT4 #(
		.INIT('hf737)
	) name5796 (
		\P2_addr_reg[0]/NET0131 ,
		_w1505_,
		_w1508_,
		_w6249_,
		_w6259_
	);
	LUT4 #(
		.INIT('hf9f5)
	) name5797 (
		\P2_IR_reg[0]/NET0131 ,
		\P2_reg2_reg[0]/NET0131 ,
		_w1505_,
		_w1508_,
		_w6260_
	);
	LUT2 #(
		.INIT('h8)
	) name5798 (
		_w6259_,
		_w6260_,
		_w6261_
	);
	LUT2 #(
		.INIT('h4)
	) name5799 (
		_w6202_,
		_w6261_,
		_w6262_
	);
	LUT4 #(
		.INIT('h444e)
	) name5800 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[0]/NET0131 ,
		_w6258_,
		_w6262_,
		_w6263_
	);
	LUT4 #(
		.INIT('h6669)
	) name5801 (
		\P2_IR_reg[10]/NET0131 ,
		\P2_reg2_reg[10]/NET0131 ,
		_w1654_,
		_w1655_,
		_w6264_
	);
	LUT4 #(
		.INIT('h5600)
	) name5802 (
		\P2_IR_reg[28]/NET0131 ,
		_w1484_,
		_w1507_,
		_w1656_,
		_w6265_
	);
	LUT4 #(
		.INIT('h6669)
	) name5803 (
		\P2_IR_reg[10]/NET0131 ,
		\P2_reg1_reg[10]/NET0131 ,
		_w1654_,
		_w1655_,
		_w6266_
	);
	LUT4 #(
		.INIT('h070d)
	) name5804 (
		_w1509_,
		_w6214_,
		_w6265_,
		_w6266_,
		_w6267_
	);
	LUT4 #(
		.INIT('h7d00)
	) name5805 (
		_w6203_,
		_w6232_,
		_w6264_,
		_w6267_,
		_w6268_
	);
	LUT4 #(
		.INIT('hc4c0)
	) name5806 (
		\P2_addr_reg[10]/NET0131 ,
		_w1477_,
		_w1486_,
		_w2080_,
		_w6269_
	);
	LUT3 #(
		.INIT('hd0)
	) name5807 (
		_w1486_,
		_w6268_,
		_w6269_,
		_w6270_
	);
	LUT4 #(
		.INIT('h5100)
	) name5808 (
		_w6114_,
		_w6117_,
		_w6136_,
		_w6266_,
		_w6271_
	);
	LUT4 #(
		.INIT('h00ae)
	) name5809 (
		_w6114_,
		_w6117_,
		_w6136_,
		_w6266_,
		_w6272_
	);
	LUT3 #(
		.INIT('h02)
	) name5810 (
		_w6149_,
		_w6272_,
		_w6271_,
		_w6273_
	);
	LUT4 #(
		.INIT('hf4f7)
	) name5811 (
		\P2_addr_reg[10]/NET0131 ,
		_w1505_,
		_w1508_,
		_w1656_,
		_w6274_
	);
	LUT4 #(
		.INIT('h5700)
	) name5812 (
		_w1477_,
		_w1486_,
		_w2080_,
		_w6274_,
		_w6275_
	);
	LUT4 #(
		.INIT('hd700)
	) name5813 (
		_w2041_,
		_w6191_,
		_w6264_,
		_w6275_,
		_w6276_
	);
	LUT3 #(
		.INIT('h8a)
	) name5814 (
		\P1_state_reg[0]/NET0131 ,
		_w6273_,
		_w6276_,
		_w6277_
	);
	LUT3 #(
		.INIT('hba)
	) name5815 (
		_w4162_,
		_w6270_,
		_w6277_,
		_w6278_
	);
	LUT4 #(
		.INIT('ha569)
	) name5816 (
		\P2_IR_reg[11]/NET0131 ,
		\P2_IR_reg[31]/NET0131 ,
		\P2_reg1_reg[11]/NET0131 ,
		_w476_,
		_w6279_
	);
	LUT2 #(
		.INIT('h1)
	) name5817 (
		_w6121_,
		_w6124_,
		_w6280_
	);
	LUT4 #(
		.INIT('h1055)
	) name5818 (
		_w6123_,
		_w6125_,
		_w6133_,
		_w6280_,
		_w6281_
	);
	LUT2 #(
		.INIT('h1)
	) name5819 (
		_w6116_,
		_w6120_,
		_w6282_
	);
	LUT4 #(
		.INIT('h1055)
	) name5820 (
		_w6118_,
		_w6119_,
		_w6281_,
		_w6282_,
		_w6283_
	);
	LUT2 #(
		.INIT('h1)
	) name5821 (
		_w6115_,
		_w6139_,
		_w6284_
	);
	LUT4 #(
		.INIT('h1055)
	) name5822 (
		_w6113_,
		_w6114_,
		_w6283_,
		_w6284_,
		_w6285_
	);
	LUT3 #(
		.INIT('h28)
	) name5823 (
		_w6149_,
		_w6279_,
		_w6285_,
		_w6286_
	);
	LUT4 #(
		.INIT('ha569)
	) name5824 (
		\P2_IR_reg[11]/NET0131 ,
		\P2_IR_reg[31]/NET0131 ,
		\P2_reg2_reg[11]/NET0131 ,
		_w476_,
		_w6287_
	);
	LUT2 #(
		.INIT('h1)
	) name5825 (
		_w6168_,
		_w6172_,
		_w6288_
	);
	LUT2 #(
		.INIT('h1)
	) name5826 (
		_w6178_,
		_w6181_,
		_w6289_
	);
	LUT4 #(
		.INIT('h1055)
	) name5827 (
		_w6180_,
		_w6182_,
		_w6188_,
		_w6289_,
		_w6290_
	);
	LUT2 #(
		.INIT('h1)
	) name5828 (
		_w6173_,
		_w6177_,
		_w6291_
	);
	LUT4 #(
		.INIT('h1055)
	) name5829 (
		_w6175_,
		_w6176_,
		_w6290_,
		_w6291_,
		_w6292_
	);
	LUT4 #(
		.INIT('h1505)
	) name5830 (
		_w6170_,
		_w6171_,
		_w6288_,
		_w6292_,
		_w6293_
	);
	LUT4 #(
		.INIT('hf4f7)
	) name5831 (
		\P2_addr_reg[11]/NET0131 ,
		_w1505_,
		_w1508_,
		_w1639_,
		_w6294_
	);
	LUT4 #(
		.INIT('h5700)
	) name5832 (
		_w1477_,
		_w1486_,
		_w2080_,
		_w6294_,
		_w6295_
	);
	LUT4 #(
		.INIT('hd700)
	) name5833 (
		_w2041_,
		_w6287_,
		_w6293_,
		_w6295_,
		_w6296_
	);
	LUT2 #(
		.INIT('h4)
	) name5834 (
		_w6286_,
		_w6296_,
		_w6297_
	);
	LUT4 #(
		.INIT('h00d4)
	) name5835 (
		\P2_reg1_reg[10]/NET0131 ,
		_w1656_,
		_w6214_,
		_w6279_,
		_w6298_
	);
	LUT4 #(
		.INIT('h2b00)
	) name5836 (
		\P2_reg1_reg[10]/NET0131 ,
		_w1656_,
		_w6214_,
		_w6279_,
		_w6299_
	);
	LUT3 #(
		.INIT('h02)
	) name5837 (
		_w1509_,
		_w6299_,
		_w6298_,
		_w6300_
	);
	LUT4 #(
		.INIT('h5600)
	) name5838 (
		\P2_IR_reg[28]/NET0131 ,
		_w1484_,
		_w1507_,
		_w1639_,
		_w6301_
	);
	LUT3 #(
		.INIT('h4d)
	) name5839 (
		\P2_reg2_reg[6]/NET0131 ,
		_w1511_,
		_w6182_,
		_w6302_
	);
	LUT4 #(
		.INIT('h4055)
	) name5840 (
		_w6177_,
		_w6228_,
		_w6289_,
		_w6302_,
		_w6303_
	);
	LUT2 #(
		.INIT('h1)
	) name5841 (
		_w6175_,
		_w6176_,
		_w6304_
	);
	LUT4 #(
		.INIT('h4044)
	) name5842 (
		_w6173_,
		_w6288_,
		_w6303_,
		_w6304_,
		_w6305_
	);
	LUT3 #(
		.INIT('h4d)
	) name5843 (
		\P2_reg2_reg[10]/NET0131 ,
		_w1656_,
		_w6171_,
		_w6306_
	);
	LUT4 #(
		.INIT('h2822)
	) name5844 (
		_w6203_,
		_w6287_,
		_w6305_,
		_w6306_,
		_w6307_
	);
	LUT2 #(
		.INIT('h1)
	) name5845 (
		_w6301_,
		_w6307_,
		_w6308_
	);
	LUT4 #(
		.INIT('hc4c0)
	) name5846 (
		\P2_addr_reg[11]/NET0131 ,
		_w1477_,
		_w1486_,
		_w2080_,
		_w6309_
	);
	LUT4 #(
		.INIT('h7500)
	) name5847 (
		_w1486_,
		_w6300_,
		_w6308_,
		_w6309_,
		_w6310_
	);
	LUT4 #(
		.INIT('h444e)
	) name5848 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[11]/NET0131 ,
		_w6310_,
		_w6297_,
		_w6311_
	);
	LUT2 #(
		.INIT('h9)
	) name5849 (
		\P2_reg2_reg[12]/NET0131 ,
		_w1744_,
		_w6312_
	);
	LUT4 #(
		.INIT('h208a)
	) name5850 (
		_w6203_,
		_w6233_,
		_w6234_,
		_w6312_,
		_w6313_
	);
	LUT4 #(
		.INIT('h5600)
	) name5851 (
		\P2_IR_reg[28]/NET0131 ,
		_w1484_,
		_w1507_,
		_w1744_,
		_w6314_
	);
	LUT2 #(
		.INIT('h9)
	) name5852 (
		\P2_reg1_reg[12]/NET0131 ,
		_w1744_,
		_w6315_
	);
	LUT4 #(
		.INIT('h02a8)
	) name5853 (
		_w1509_,
		_w6112_,
		_w6215_,
		_w6315_,
		_w6316_
	);
	LUT4 #(
		.INIT('haaa8)
	) name5854 (
		_w1486_,
		_w6314_,
		_w6316_,
		_w6313_,
		_w6317_
	);
	LUT4 #(
		.INIT('hc4c0)
	) name5855 (
		\P2_addr_reg[12]/NET0131 ,
		_w1477_,
		_w1486_,
		_w2080_,
		_w6318_
	);
	LUT2 #(
		.INIT('h4)
	) name5856 (
		_w6317_,
		_w6318_,
		_w6319_
	);
	LUT4 #(
		.INIT('h4500)
	) name5857 (
		_w6112_,
		_w6137_,
		_w6140_,
		_w6315_,
		_w6320_
	);
	LUT4 #(
		.INIT('h00ba)
	) name5858 (
		_w6112_,
		_w6137_,
		_w6140_,
		_w6315_,
		_w6321_
	);
	LUT3 #(
		.INIT('h02)
	) name5859 (
		_w6149_,
		_w6321_,
		_w6320_,
		_w6322_
	);
	LUT4 #(
		.INIT('hf4f7)
	) name5860 (
		\P2_addr_reg[12]/NET0131 ,
		_w1505_,
		_w1508_,
		_w1744_,
		_w6323_
	);
	LUT4 #(
		.INIT('h5700)
	) name5861 (
		_w1477_,
		_w1486_,
		_w2080_,
		_w6323_,
		_w6324_
	);
	LUT4 #(
		.INIT('hd700)
	) name5862 (
		_w2041_,
		_w6193_,
		_w6312_,
		_w6324_,
		_w6325_
	);
	LUT3 #(
		.INIT('h8a)
	) name5863 (
		\P1_state_reg[0]/NET0131 ,
		_w6322_,
		_w6325_,
		_w6326_
	);
	LUT3 #(
		.INIT('hba)
	) name5864 (
		_w4185_,
		_w6319_,
		_w6326_,
		_w6327_
	);
	LUT2 #(
		.INIT('h9)
	) name5865 (
		\P2_reg1_reg[13]/NET0131 ,
		_w1759_,
		_w6328_
	);
	LUT3 #(
		.INIT('h0b)
	) name5866 (
		\P2_reg1_reg[12]/NET0131 ,
		_w1744_,
		_w6138_,
		_w6329_
	);
	LUT4 #(
		.INIT('h1055)
	) name5867 (
		_w6111_,
		_w6112_,
		_w6285_,
		_w6329_,
		_w6330_
	);
	LUT3 #(
		.INIT('h28)
	) name5868 (
		_w6149_,
		_w6328_,
		_w6330_,
		_w6331_
	);
	LUT2 #(
		.INIT('h9)
	) name5869 (
		\P2_reg2_reg[13]/NET0131 ,
		_w1759_,
		_w6332_
	);
	LUT3 #(
		.INIT('h0b)
	) name5870 (
		\P2_reg2_reg[12]/NET0131 ,
		_w1744_,
		_w6167_,
		_w6333_
	);
	LUT4 #(
		.INIT('h1055)
	) name5871 (
		_w6165_,
		_w6166_,
		_w6293_,
		_w6333_,
		_w6334_
	);
	LUT4 #(
		.INIT('hf4f7)
	) name5872 (
		\P2_addr_reg[13]/NET0131 ,
		_w1505_,
		_w1508_,
		_w1759_,
		_w6335_
	);
	LUT4 #(
		.INIT('h5700)
	) name5873 (
		_w1477_,
		_w1486_,
		_w2080_,
		_w6335_,
		_w6336_
	);
	LUT4 #(
		.INIT('hd700)
	) name5874 (
		_w2041_,
		_w6332_,
		_w6334_,
		_w6336_,
		_w6337_
	);
	LUT2 #(
		.INIT('h4)
	) name5875 (
		_w6331_,
		_w6337_,
		_w6338_
	);
	LUT4 #(
		.INIT('h4500)
	) name5876 (
		_w6109_,
		_w6215_,
		_w6216_,
		_w6328_,
		_w6339_
	);
	LUT4 #(
		.INIT('h00ba)
	) name5877 (
		_w6109_,
		_w6215_,
		_w6216_,
		_w6328_,
		_w6340_
	);
	LUT3 #(
		.INIT('h02)
	) name5878 (
		_w1509_,
		_w6340_,
		_w6339_,
		_w6341_
	);
	LUT4 #(
		.INIT('h5600)
	) name5879 (
		\P2_IR_reg[28]/NET0131 ,
		_w1484_,
		_w1507_,
		_w1759_,
		_w6342_
	);
	LUT3 #(
		.INIT('h0d)
	) name5880 (
		\P2_reg2_reg[12]/NET0131 ,
		_w1744_,
		_w6166_,
		_w6343_
	);
	LUT4 #(
		.INIT('hba00)
	) name5881 (
		_w6167_,
		_w6305_,
		_w6306_,
		_w6343_,
		_w6344_
	);
	LUT4 #(
		.INIT('hc084)
	) name5882 (
		_w6163_,
		_w6203_,
		_w6332_,
		_w6344_,
		_w6345_
	);
	LUT2 #(
		.INIT('h1)
	) name5883 (
		_w6342_,
		_w6345_,
		_w6346_
	);
	LUT4 #(
		.INIT('hc4c0)
	) name5884 (
		\P2_addr_reg[13]/NET0131 ,
		_w1477_,
		_w1486_,
		_w2080_,
		_w6347_
	);
	LUT4 #(
		.INIT('h7500)
	) name5885 (
		_w1486_,
		_w6341_,
		_w6346_,
		_w6347_,
		_w6348_
	);
	LUT4 #(
		.INIT('h444e)
	) name5886 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[13]/NET0131 ,
		_w6348_,
		_w6338_,
		_w6349_
	);
	LUT2 #(
		.INIT('h6)
	) name5887 (
		\P2_reg1_reg[14]/NET0131 ,
		_w1728_,
		_w6350_
	);
	LUT4 #(
		.INIT('h00ae)
	) name5888 (
		_w6108_,
		_w6110_,
		_w6141_,
		_w6350_,
		_w6351_
	);
	LUT4 #(
		.INIT('h5100)
	) name5889 (
		_w6108_,
		_w6110_,
		_w6141_,
		_w6350_,
		_w6352_
	);
	LUT3 #(
		.INIT('h02)
	) name5890 (
		_w6149_,
		_w6352_,
		_w6351_,
		_w6353_
	);
	LUT2 #(
		.INIT('h6)
	) name5891 (
		\P2_reg2_reg[14]/NET0131 ,
		_w1728_,
		_w6354_
	);
	LUT4 #(
		.INIT('hf7f4)
	) name5892 (
		\P2_addr_reg[14]/NET0131 ,
		_w1505_,
		_w1508_,
		_w1728_,
		_w6355_
	);
	LUT4 #(
		.INIT('h5700)
	) name5893 (
		_w1477_,
		_w1486_,
		_w2080_,
		_w6355_,
		_w6356_
	);
	LUT4 #(
		.INIT('hd700)
	) name5894 (
		_w2041_,
		_w6195_,
		_w6354_,
		_w6356_,
		_w6357_
	);
	LUT3 #(
		.INIT('h82)
	) name5895 (
		_w6203_,
		_w6236_,
		_w6354_,
		_w6358_
	);
	LUT4 #(
		.INIT('h0056)
	) name5896 (
		\P2_IR_reg[28]/NET0131 ,
		_w1484_,
		_w1507_,
		_w1728_,
		_w6359_
	);
	LUT4 #(
		.INIT('h1511)
	) name5897 (
		_w6108_,
		_w6110_,
		_w6215_,
		_w6216_,
		_w6360_
	);
	LUT4 #(
		.INIT('h1331)
	) name5898 (
		_w1509_,
		_w6359_,
		_w6350_,
		_w6360_,
		_w6361_
	);
	LUT4 #(
		.INIT('hc4c0)
	) name5899 (
		\P2_addr_reg[14]/NET0131 ,
		_w1477_,
		_w1486_,
		_w2080_,
		_w6362_
	);
	LUT4 #(
		.INIT('h7500)
	) name5900 (
		_w1486_,
		_w6358_,
		_w6361_,
		_w6362_,
		_w6363_
	);
	LUT4 #(
		.INIT('h2022)
	) name5901 (
		\P1_state_reg[0]/NET0131 ,
		_w6363_,
		_w6353_,
		_w6357_,
		_w6364_
	);
	LUT2 #(
		.INIT('he)
	) name5902 (
		_w4511_,
		_w6364_,
		_w6365_
	);
	LUT3 #(
		.INIT('h96)
	) name5903 (
		\P2_IR_reg[15]/NET0131 ,
		\P2_reg2_reg[15]/NET0131 ,
		_w1712_,
		_w6366_
	);
	LUT4 #(
		.INIT('ha8fc)
	) name5904 (
		\P2_reg2_reg[13]/NET0131 ,
		\P2_reg2_reg[14]/NET0131 ,
		_w1728_,
		_w1759_,
		_w6367_
	);
	LUT4 #(
		.INIT('h1055)
	) name5905 (
		_w6161_,
		_w6162_,
		_w6334_,
		_w6367_,
		_w6368_
	);
	LUT3 #(
		.INIT('h28)
	) name5906 (
		_w2041_,
		_w6366_,
		_w6368_,
		_w6369_
	);
	LUT3 #(
		.INIT('h96)
	) name5907 (
		\P2_IR_reg[15]/NET0131 ,
		\P2_reg1_reg[15]/NET0131 ,
		_w1712_,
		_w6370_
	);
	LUT4 #(
		.INIT('ha8fc)
	) name5908 (
		\P2_reg1_reg[13]/NET0131 ,
		\P2_reg1_reg[14]/NET0131 ,
		_w1728_,
		_w1759_,
		_w6371_
	);
	LUT4 #(
		.INIT('h1055)
	) name5909 (
		_w6107_,
		_w6108_,
		_w6330_,
		_w6371_,
		_w6372_
	);
	LUT4 #(
		.INIT('hf4f7)
	) name5910 (
		\P2_addr_reg[15]/NET0131 ,
		_w1505_,
		_w1508_,
		_w1713_,
		_w6373_
	);
	LUT4 #(
		.INIT('h5700)
	) name5911 (
		_w1477_,
		_w1486_,
		_w2080_,
		_w6373_,
		_w6374_
	);
	LUT4 #(
		.INIT('hd700)
	) name5912 (
		_w6149_,
		_w6370_,
		_w6372_,
		_w6374_,
		_w6375_
	);
	LUT4 #(
		.INIT('ha802)
	) name5913 (
		_w1509_,
		_w6105_,
		_w6218_,
		_w6370_,
		_w6376_
	);
	LUT2 #(
		.INIT('h8)
	) name5914 (
		_w1508_,
		_w1713_,
		_w6377_
	);
	LUT4 #(
		.INIT('h3f17)
	) name5915 (
		\P2_reg2_reg[13]/NET0131 ,
		\P2_reg2_reg[14]/NET0131 ,
		_w1728_,
		_w1759_,
		_w6378_
	);
	LUT4 #(
		.INIT('hef00)
	) name5916 (
		_w6163_,
		_w6344_,
		_w6367_,
		_w6378_,
		_w6379_
	);
	LUT4 #(
		.INIT('h1331)
	) name5917 (
		_w6203_,
		_w6377_,
		_w6366_,
		_w6379_,
		_w6380_
	);
	LUT4 #(
		.INIT('hc4c0)
	) name5918 (
		\P2_addr_reg[15]/NET0131 ,
		_w1477_,
		_w1486_,
		_w2080_,
		_w6381_
	);
	LUT4 #(
		.INIT('h7500)
	) name5919 (
		_w1486_,
		_w6376_,
		_w6380_,
		_w6381_,
		_w6382_
	);
	LUT4 #(
		.INIT('h2022)
	) name5920 (
		\P1_state_reg[0]/NET0131 ,
		_w6382_,
		_w6369_,
		_w6375_,
		_w6383_
	);
	LUT2 #(
		.INIT('he)
	) name5921 (
		_w4533_,
		_w6383_,
		_w6384_
	);
	LUT2 #(
		.INIT('h4)
	) name5922 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[16]/NET0131 ,
		_w6385_
	);
	LUT3 #(
		.INIT('h96)
	) name5923 (
		\P2_IR_reg[16]/NET0131 ,
		\P2_reg2_reg[16]/NET0131 ,
		_w1792_,
		_w6386_
	);
	LUT4 #(
		.INIT('h00ae)
	) name5924 (
		_w6157_,
		_w6160_,
		_w6196_,
		_w6386_,
		_w6387_
	);
	LUT4 #(
		.INIT('h5100)
	) name5925 (
		_w6157_,
		_w6160_,
		_w6196_,
		_w6386_,
		_w6388_
	);
	LUT3 #(
		.INIT('h02)
	) name5926 (
		_w2041_,
		_w6388_,
		_w6387_,
		_w6389_
	);
	LUT3 #(
		.INIT('h96)
	) name5927 (
		\P2_IR_reg[16]/NET0131 ,
		\P2_reg1_reg[16]/NET0131 ,
		_w1792_,
		_w6390_
	);
	LUT4 #(
		.INIT('hf4f7)
	) name5928 (
		\P2_addr_reg[16]/NET0131 ,
		_w1505_,
		_w1508_,
		_w1793_,
		_w6391_
	);
	LUT4 #(
		.INIT('h5700)
	) name5929 (
		_w1477_,
		_w1486_,
		_w2080_,
		_w6391_,
		_w6392_
	);
	LUT4 #(
		.INIT('hd700)
	) name5930 (
		_w6149_,
		_w6143_,
		_w6390_,
		_w6392_,
		_w6393_
	);
	LUT4 #(
		.INIT('h000d)
	) name5931 (
		_w6160_,
		_w6236_,
		_w6237_,
		_w6386_,
		_w6394_
	);
	LUT4 #(
		.INIT('hf200)
	) name5932 (
		_w6160_,
		_w6236_,
		_w6237_,
		_w6386_,
		_w6395_
	);
	LUT3 #(
		.INIT('h02)
	) name5933 (
		_w6203_,
		_w6395_,
		_w6394_,
		_w6396_
	);
	LUT2 #(
		.INIT('h8)
	) name5934 (
		_w1508_,
		_w1793_,
		_w6397_
	);
	LUT4 #(
		.INIT('h070d)
	) name5935 (
		_w1509_,
		_w6219_,
		_w6397_,
		_w6390_,
		_w6398_
	);
	LUT4 #(
		.INIT('hc4c0)
	) name5936 (
		\P2_addr_reg[16]/NET0131 ,
		_w1477_,
		_w1486_,
		_w2080_,
		_w6399_
	);
	LUT4 #(
		.INIT('h7500)
	) name5937 (
		_w1486_,
		_w6396_,
		_w6398_,
		_w6399_,
		_w6400_
	);
	LUT4 #(
		.INIT('h2022)
	) name5938 (
		\P1_state_reg[0]/NET0131 ,
		_w6400_,
		_w6389_,
		_w6393_,
		_w6401_
	);
	LUT2 #(
		.INIT('he)
	) name5939 (
		_w6385_,
		_w6401_,
		_w6402_
	);
	LUT3 #(
		.INIT('h96)
	) name5940 (
		\P2_IR_reg[17]/NET0131 ,
		\P2_reg1_reg[17]/NET0131 ,
		_w1773_,
		_w6403_
	);
	LUT2 #(
		.INIT('h1)
	) name5941 (
		_w6102_,
		_w6103_,
		_w6404_
	);
	LUT4 #(
		.INIT('h0455)
	) name5942 (
		_w6146_,
		_w6106_,
		_w6218_,
		_w6404_,
		_w6405_
	);
	LUT3 #(
		.INIT('h28)
	) name5943 (
		_w1509_,
		_w6403_,
		_w6405_,
		_w6406_
	);
	LUT2 #(
		.INIT('h8)
	) name5944 (
		_w1508_,
		_w1774_,
		_w6407_
	);
	LUT3 #(
		.INIT('h96)
	) name5945 (
		\P2_IR_reg[17]/NET0131 ,
		\P2_reg2_reg[17]/NET0131 ,
		_w1773_,
		_w6408_
	);
	LUT2 #(
		.INIT('h1)
	) name5946 (
		_w6156_,
		_w6157_,
		_w6409_
	);
	LUT3 #(
		.INIT('hb2)
	) name5947 (
		\P2_reg2_reg[16]/NET0131 ,
		_w1793_,
		_w6157_,
		_w6410_
	);
	LUT2 #(
		.INIT('h1)
	) name5948 (
		_w6198_,
		_w6158_,
		_w6411_
	);
	LUT3 #(
		.INIT('h23)
	) name5949 (
		_w6379_,
		_w6410_,
		_w6411_,
		_w6412_
	);
	LUT4 #(
		.INIT('h1331)
	) name5950 (
		_w6203_,
		_w6407_,
		_w6408_,
		_w6412_,
		_w6413_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name5951 (
		\P2_addr_reg[17]/NET0131 ,
		_w1483_,
		_w1485_,
		_w1481_,
		_w6414_
	);
	LUT2 #(
		.INIT('h8)
	) name5952 (
		_w2080_,
		_w6414_,
		_w6415_
	);
	LUT4 #(
		.INIT('h0075)
	) name5953 (
		_w1486_,
		_w6406_,
		_w6413_,
		_w6415_,
		_w6416_
	);
	LUT2 #(
		.INIT('h2)
	) name5954 (
		_w1477_,
		_w6416_,
		_w6417_
	);
	LUT4 #(
		.INIT('hc4c0)
	) name5955 (
		\P2_addr_reg[17]/NET0131 ,
		_w1477_,
		_w1486_,
		_w2080_,
		_w6418_
	);
	LUT3 #(
		.INIT('hd4)
	) name5956 (
		\P2_reg2_reg[16]/NET0131 ,
		_w1793_,
		_w6158_,
		_w6419_
	);
	LUT4 #(
		.INIT('h0013)
	) name5957 (
		_w6368_,
		_w6408_,
		_w6409_,
		_w6419_,
		_w6420_
	);
	LUT4 #(
		.INIT('hcc80)
	) name5958 (
		_w6368_,
		_w6408_,
		_w6409_,
		_w6419_,
		_w6421_
	);
	LUT3 #(
		.INIT('h02)
	) name5959 (
		_w2041_,
		_w6421_,
		_w6420_,
		_w6422_
	);
	LUT3 #(
		.INIT('hd4)
	) name5960 (
		\P2_reg1_reg[16]/NET0131 ,
		_w1793_,
		_w6104_,
		_w6423_
	);
	LUT3 #(
		.INIT('h07)
	) name5961 (
		_w6372_,
		_w6404_,
		_w6423_,
		_w6424_
	);
	LUT4 #(
		.INIT('hf4f7)
	) name5962 (
		\P2_addr_reg[17]/NET0131 ,
		_w1505_,
		_w1508_,
		_w1774_,
		_w6425_
	);
	LUT4 #(
		.INIT('h7d00)
	) name5963 (
		_w6149_,
		_w6403_,
		_w6424_,
		_w6425_,
		_w6426_
	);
	LUT3 #(
		.INIT('h45)
	) name5964 (
		_w6418_,
		_w6422_,
		_w6426_,
		_w6427_
	);
	LUT4 #(
		.INIT('heee4)
	) name5965 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[17]/NET0131 ,
		_w6417_,
		_w6427_,
		_w6428_
	);
	LUT2 #(
		.INIT('h1)
	) name5966 (
		_w6098_,
		_w6145_,
		_w6429_
	);
	LUT4 #(
		.INIT('h5540)
	) name5967 (
		_w6101_,
		_w6372_,
		_w6404_,
		_w6423_,
		_w6430_
	);
	LUT3 #(
		.INIT('h69)
	) name5968 (
		\P2_IR_reg[19]/NET0131 ,
		\P2_reg1_reg[19]/NET0131 ,
		_w1810_,
		_w6431_
	);
	LUT4 #(
		.INIT('h0051)
	) name5969 (
		_w6099_,
		_w6429_,
		_w6430_,
		_w6431_,
		_w6432_
	);
	LUT4 #(
		.INIT('hae00)
	) name5970 (
		_w6099_,
		_w6429_,
		_w6430_,
		_w6431_,
		_w6433_
	);
	LUT3 #(
		.INIT('h02)
	) name5971 (
		_w6149_,
		_w6433_,
		_w6432_,
		_w6434_
	);
	LUT2 #(
		.INIT('h1)
	) name5972 (
		_w6152_,
		_w6199_,
		_w6435_
	);
	LUT4 #(
		.INIT('h0d04)
	) name5973 (
		\P2_reg2_reg[16]/NET0131 ,
		_w1793_,
		_w6155_,
		_w6158_,
		_w6436_
	);
	LUT2 #(
		.INIT('h2)
	) name5974 (
		_w6435_,
		_w6436_,
		_w6437_
	);
	LUT4 #(
		.INIT('hbf00)
	) name5975 (
		_w6155_,
		_w6368_,
		_w6409_,
		_w6437_,
		_w6438_
	);
	LUT3 #(
		.INIT('h69)
	) name5976 (
		\P2_IR_reg[19]/NET0131 ,
		\P2_reg2_reg[19]/NET0131 ,
		_w1810_,
		_w6439_
	);
	LUT4 #(
		.INIT('h02a8)
	) name5977 (
		_w2041_,
		_w6153_,
		_w6438_,
		_w6439_,
		_w6440_
	);
	LUT4 #(
		.INIT('hf4f7)
	) name5978 (
		\P2_addr_reg[19]/NET0131 ,
		_w1505_,
		_w1508_,
		_w1811_,
		_w6441_
	);
	LUT2 #(
		.INIT('h4)
	) name5979 (
		_w6440_,
		_w6441_,
		_w6442_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name5980 (
		\P2_addr_reg[19]/NET0131 ,
		_w1483_,
		_w1485_,
		_w1481_,
		_w6443_
	);
	LUT4 #(
		.INIT('hc4c0)
	) name5981 (
		\P2_addr_reg[19]/NET0131 ,
		_w1477_,
		_w1486_,
		_w2080_,
		_w6444_
	);
	LUT3 #(
		.INIT('h0b)
	) name5982 (
		_w6434_,
		_w6442_,
		_w6444_,
		_w6445_
	);
	LUT2 #(
		.INIT('h8)
	) name5983 (
		_w2080_,
		_w6443_,
		_w6446_
	);
	LUT4 #(
		.INIT('h0155)
	) name5984 (
		_w6099_,
		_w6101_,
		_w6405_,
		_w6429_,
		_w6447_
	);
	LUT3 #(
		.INIT('h28)
	) name5985 (
		_w1509_,
		_w6431_,
		_w6447_,
		_w6448_
	);
	LUT2 #(
		.INIT('h8)
	) name5986 (
		_w1508_,
		_w1811_,
		_w6449_
	);
	LUT4 #(
		.INIT('h0405)
	) name5987 (
		_w6155_,
		_w6379_,
		_w6410_,
		_w6411_,
		_w6450_
	);
	LUT3 #(
		.INIT('h51)
	) name5988 (
		_w6153_,
		_w6435_,
		_w6450_,
		_w6451_
	);
	LUT4 #(
		.INIT('h0d07)
	) name5989 (
		_w6203_,
		_w6439_,
		_w6449_,
		_w6451_,
		_w6452_
	);
	LUT4 #(
		.INIT('h1311)
	) name5990 (
		_w1486_,
		_w6446_,
		_w6448_,
		_w6452_,
		_w6453_
	);
	LUT2 #(
		.INIT('h2)
	) name5991 (
		_w1477_,
		_w6453_,
		_w6454_
	);
	LUT4 #(
		.INIT('heee4)
	) name5992 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[19]/NET0131 ,
		_w6445_,
		_w6454_,
		_w6455_
	);
	LUT4 #(
		.INIT('h6c93)
	) name5993 (
		\P2_IR_reg[0]/NET0131 ,
		\P2_IR_reg[1]/NET0131 ,
		\P2_IR_reg[31]/NET0131 ,
		\P2_reg1_reg[1]/NET0131 ,
		_w6456_
	);
	LUT2 #(
		.INIT('h9)
	) name5994 (
		_w6207_,
		_w6456_,
		_w6457_
	);
	LUT3 #(
		.INIT('h20)
	) name5995 (
		_w1505_,
		_w1508_,
		_w6457_,
		_w6458_
	);
	LUT4 #(
		.INIT('h6c93)
	) name5996 (
		\P2_IR_reg[0]/NET0131 ,
		\P2_IR_reg[1]/NET0131 ,
		\P2_IR_reg[31]/NET0131 ,
		\P2_reg2_reg[1]/NET0131 ,
		_w6459_
	);
	LUT2 #(
		.INIT('h9)
	) name5997 (
		_w6225_,
		_w6459_,
		_w6460_
	);
	LUT3 #(
		.INIT('h10)
	) name5998 (
		_w1505_,
		_w1508_,
		_w6460_,
		_w6461_
	);
	LUT4 #(
		.INIT('h0056)
	) name5999 (
		\P2_IR_reg[28]/NET0131 ,
		_w1484_,
		_w1507_,
		_w1571_,
		_w6462_
	);
	LUT4 #(
		.INIT('h0080)
	) name6000 (
		_w1483_,
		_w1485_,
		_w1481_,
		_w6462_,
		_w6463_
	);
	LUT3 #(
		.INIT('h10)
	) name6001 (
		_w6461_,
		_w6458_,
		_w6463_,
		_w6464_
	);
	LUT4 #(
		.INIT('h1555)
	) name6002 (
		\P2_addr_reg[1]/NET0131 ,
		_w1483_,
		_w1485_,
		_w1481_,
		_w6465_
	);
	LUT2 #(
		.INIT('h8)
	) name6003 (
		_w2080_,
		_w6465_,
		_w6466_
	);
	LUT3 #(
		.INIT('ha8)
	) name6004 (
		_w1477_,
		_w6464_,
		_w6466_,
		_w6467_
	);
	LUT2 #(
		.INIT('h9)
	) name6005 (
		_w6185_,
		_w6459_,
		_w6468_
	);
	LUT4 #(
		.INIT('hc7f7)
	) name6006 (
		\P2_addr_reg[1]/NET0131 ,
		_w1505_,
		_w1508_,
		_w6468_,
		_w6469_
	);
	LUT2 #(
		.INIT('h9)
	) name6007 (
		_w6130_,
		_w6456_,
		_w6470_
	);
	LUT4 #(
		.INIT('h76fe)
	) name6008 (
		_w1505_,
		_w1508_,
		_w1571_,
		_w6470_,
		_w6471_
	);
	LUT2 #(
		.INIT('h8)
	) name6009 (
		_w6469_,
		_w6471_,
		_w6472_
	);
	LUT2 #(
		.INIT('h4)
	) name6010 (
		_w6202_,
		_w6472_,
		_w6473_
	);
	LUT4 #(
		.INIT('h444e)
	) name6011 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[1]/NET0131 ,
		_w6467_,
		_w6473_,
		_w6474_
	);
	LUT2 #(
		.INIT('h6)
	) name6012 (
		\P2_reg2_reg[2]/NET0131 ,
		_w1561_,
		_w6475_
	);
	LUT2 #(
		.INIT('h6)
	) name6013 (
		_w6226_,
		_w6475_,
		_w6476_
	);
	LUT3 #(
		.INIT('h10)
	) name6014 (
		_w1505_,
		_w1508_,
		_w6476_,
		_w6477_
	);
	LUT2 #(
		.INIT('h6)
	) name6015 (
		\P2_reg1_reg[2]/NET0131 ,
		_w1561_,
		_w6478_
	);
	LUT2 #(
		.INIT('h6)
	) name6016 (
		_w6208_,
		_w6478_,
		_w6479_
	);
	LUT3 #(
		.INIT('h20)
	) name6017 (
		_w1505_,
		_w1508_,
		_w6479_,
		_w6480_
	);
	LUT4 #(
		.INIT('h0056)
	) name6018 (
		\P2_IR_reg[28]/NET0131 ,
		_w1484_,
		_w1507_,
		_w1561_,
		_w6481_
	);
	LUT4 #(
		.INIT('h0080)
	) name6019 (
		_w1483_,
		_w1485_,
		_w1481_,
		_w6481_,
		_w6482_
	);
	LUT3 #(
		.INIT('h10)
	) name6020 (
		_w6480_,
		_w6477_,
		_w6482_,
		_w6483_
	);
	LUT4 #(
		.INIT('h1555)
	) name6021 (
		\P2_addr_reg[2]/NET0131 ,
		_w1483_,
		_w1485_,
		_w1481_,
		_w6484_
	);
	LUT2 #(
		.INIT('h8)
	) name6022 (
		_w2080_,
		_w6484_,
		_w6485_
	);
	LUT3 #(
		.INIT('ha8)
	) name6023 (
		_w1477_,
		_w6483_,
		_w6485_,
		_w6486_
	);
	LUT2 #(
		.INIT('h9)
	) name6024 (
		_w6131_,
		_w6478_,
		_w6487_
	);
	LUT4 #(
		.INIT('h37f7)
	) name6025 (
		\P2_addr_reg[2]/NET0131 ,
		_w1505_,
		_w1508_,
		_w6487_,
		_w6488_
	);
	LUT2 #(
		.INIT('h9)
	) name6026 (
		_w6186_,
		_w6475_,
		_w6489_
	);
	LUT4 #(
		.INIT('hbafe)
	) name6027 (
		_w1505_,
		_w1508_,
		_w1561_,
		_w6489_,
		_w6490_
	);
	LUT2 #(
		.INIT('h8)
	) name6028 (
		_w6488_,
		_w6490_,
		_w6491_
	);
	LUT2 #(
		.INIT('h4)
	) name6029 (
		_w6202_,
		_w6491_,
		_w6492_
	);
	LUT4 #(
		.INIT('h444e)
	) name6030 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[2]/NET0131 ,
		_w6486_,
		_w6492_,
		_w6493_
	);
	LUT3 #(
		.INIT('h69)
	) name6031 (
		\P2_IR_reg[3]/NET0131 ,
		\P2_reg1_reg[3]/NET0131 ,
		_w1553_,
		_w6494_
	);
	LUT4 #(
		.INIT('h17e8)
	) name6032 (
		\P2_reg1_reg[2]/NET0131 ,
		_w1561_,
		_w6208_,
		_w6494_,
		_w6495_
	);
	LUT3 #(
		.INIT('h20)
	) name6033 (
		_w1505_,
		_w1508_,
		_w6495_,
		_w6496_
	);
	LUT3 #(
		.INIT('h69)
	) name6034 (
		\P2_IR_reg[3]/NET0131 ,
		\P2_reg2_reg[3]/NET0131 ,
		_w1553_,
		_w6497_
	);
	LUT4 #(
		.INIT('h17e8)
	) name6035 (
		\P2_reg2_reg[2]/NET0131 ,
		_w1561_,
		_w6226_,
		_w6497_,
		_w6498_
	);
	LUT3 #(
		.INIT('h10)
	) name6036 (
		_w1505_,
		_w1508_,
		_w6498_,
		_w6499_
	);
	LUT4 #(
		.INIT('h5600)
	) name6037 (
		\P2_IR_reg[28]/NET0131 ,
		_w1484_,
		_w1507_,
		_w1554_,
		_w6500_
	);
	LUT4 #(
		.INIT('h0080)
	) name6038 (
		_w1483_,
		_w1485_,
		_w1481_,
		_w6500_,
		_w6501_
	);
	LUT3 #(
		.INIT('h10)
	) name6039 (
		_w6499_,
		_w6496_,
		_w6501_,
		_w6502_
	);
	LUT4 #(
		.INIT('h1555)
	) name6040 (
		\P2_addr_reg[3]/NET0131 ,
		_w1483_,
		_w1485_,
		_w1481_,
		_w6503_
	);
	LUT2 #(
		.INIT('h8)
	) name6041 (
		_w2080_,
		_w6503_,
		_w6504_
	);
	LUT3 #(
		.INIT('ha8)
	) name6042 (
		_w1477_,
		_w6502_,
		_w6504_,
		_w6505_
	);
	LUT4 #(
		.INIT('he817)
	) name6043 (
		\P2_reg1_reg[2]/NET0131 ,
		_w1561_,
		_w6131_,
		_w6494_,
		_w6506_
	);
	LUT4 #(
		.INIT('h67ef)
	) name6044 (
		_w1505_,
		_w1508_,
		_w1554_,
		_w6506_,
		_w6507_
	);
	LUT4 #(
		.INIT('he817)
	) name6045 (
		\P2_reg2_reg[2]/NET0131 ,
		_w1561_,
		_w6186_,
		_w6497_,
		_w6508_
	);
	LUT4 #(
		.INIT('hc7f7)
	) name6046 (
		\P2_addr_reg[3]/NET0131 ,
		_w1505_,
		_w1508_,
		_w6508_,
		_w6509_
	);
	LUT2 #(
		.INIT('h8)
	) name6047 (
		_w6507_,
		_w6509_,
		_w6510_
	);
	LUT3 #(
		.INIT('h8a)
	) name6048 (
		\P1_state_reg[0]/NET0131 ,
		_w6202_,
		_w6510_,
		_w6511_
	);
	LUT3 #(
		.INIT('hba)
	) name6049 (
		_w5544_,
		_w6505_,
		_w6511_,
		_w6512_
	);
	LUT4 #(
		.INIT('hc369)
	) name6050 (
		\P2_IR_reg[31]/NET0131 ,
		\P2_IR_reg[4]/NET0131 ,
		\P2_reg1_reg[4]/NET0131 ,
		_w472_,
		_w6513_
	);
	LUT3 #(
		.INIT('he1)
	) name6051 (
		_w6129_,
		_w6209_,
		_w6513_,
		_w6514_
	);
	LUT3 #(
		.INIT('h20)
	) name6052 (
		_w1505_,
		_w1508_,
		_w6514_,
		_w6515_
	);
	LUT4 #(
		.INIT('hc369)
	) name6053 (
		\P2_IR_reg[31]/NET0131 ,
		\P2_IR_reg[4]/NET0131 ,
		\P2_reg2_reg[4]/NET0131 ,
		_w472_,
		_w6516_
	);
	LUT3 #(
		.INIT('he1)
	) name6054 (
		_w6184_,
		_w6227_,
		_w6516_,
		_w6517_
	);
	LUT3 #(
		.INIT('h10)
	) name6055 (
		_w1505_,
		_w1508_,
		_w6517_,
		_w6518_
	);
	LUT4 #(
		.INIT('h5600)
	) name6056 (
		\P2_IR_reg[28]/NET0131 ,
		_w1484_,
		_w1507_,
		_w1601_,
		_w6519_
	);
	LUT4 #(
		.INIT('h0080)
	) name6057 (
		_w1483_,
		_w1485_,
		_w1481_,
		_w6519_,
		_w6520_
	);
	LUT3 #(
		.INIT('h10)
	) name6058 (
		_w6518_,
		_w6515_,
		_w6520_,
		_w6521_
	);
	LUT4 #(
		.INIT('h1555)
	) name6059 (
		\P2_addr_reg[4]/NET0131 ,
		_w1483_,
		_w1485_,
		_w1481_,
		_w6522_
	);
	LUT2 #(
		.INIT('h8)
	) name6060 (
		_w2080_,
		_w6522_,
		_w6523_
	);
	LUT3 #(
		.INIT('ha8)
	) name6061 (
		_w1477_,
		_w6521_,
		_w6523_,
		_w6524_
	);
	LUT4 #(
		.INIT('hf4f7)
	) name6062 (
		\P2_addr_reg[4]/NET0131 ,
		_w1505_,
		_w1508_,
		_w1601_,
		_w6525_
	);
	LUT3 #(
		.INIT('he1)
	) name6063 (
		_w6128_,
		_w6132_,
		_w6513_,
		_w6526_
	);
	LUT3 #(
		.INIT('he1)
	) name6064 (
		_w6183_,
		_w6187_,
		_w6516_,
		_w6527_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name6065 (
		_w1505_,
		_w1508_,
		_w6526_,
		_w6527_,
		_w6528_
	);
	LUT2 #(
		.INIT('h8)
	) name6066 (
		_w6525_,
		_w6528_,
		_w6529_
	);
	LUT3 #(
		.INIT('h8a)
	) name6067 (
		\P1_state_reg[0]/NET0131 ,
		_w6202_,
		_w6529_,
		_w6530_
	);
	LUT3 #(
		.INIT('hba)
	) name6068 (
		_w5279_,
		_w6524_,
		_w6530_,
		_w6531_
	);
	LUT3 #(
		.INIT('h69)
	) name6069 (
		\P2_IR_reg[6]/NET0131 ,
		\P2_reg2_reg[6]/NET0131 ,
		_w1510_,
		_w6532_
	);
	LUT4 #(
		.INIT('he800)
	) name6070 (
		\P2_reg2_reg[5]/NET0131 ,
		_w1592_,
		_w6228_,
		_w6532_,
		_w6533_
	);
	LUT4 #(
		.INIT('h0017)
	) name6071 (
		\P2_reg2_reg[5]/NET0131 ,
		_w1592_,
		_w6228_,
		_w6532_,
		_w6534_
	);
	LUT3 #(
		.INIT('h02)
	) name6072 (
		_w6203_,
		_w6534_,
		_w6533_,
		_w6535_
	);
	LUT4 #(
		.INIT('h5600)
	) name6073 (
		\P2_IR_reg[28]/NET0131 ,
		_w1484_,
		_w1507_,
		_w1511_,
		_w6536_
	);
	LUT3 #(
		.INIT('h69)
	) name6074 (
		\P2_IR_reg[6]/NET0131 ,
		\P2_reg1_reg[6]/NET0131 ,
		_w1510_,
		_w6537_
	);
	LUT2 #(
		.INIT('h1)
	) name6075 (
		_w6125_,
		_w6211_,
		_w6538_
	);
	LUT4 #(
		.INIT('h070d)
	) name6076 (
		_w1509_,
		_w6537_,
		_w6536_,
		_w6538_,
		_w6539_
	);
	LUT4 #(
		.INIT('hc4c0)
	) name6077 (
		\P2_addr_reg[6]/NET0131 ,
		_w1477_,
		_w1486_,
		_w2080_,
		_w6540_
	);
	LUT4 #(
		.INIT('h7500)
	) name6078 (
		_w1486_,
		_w6535_,
		_w6539_,
		_w6540_,
		_w6541_
	);
	LUT4 #(
		.INIT('h008e)
	) name6079 (
		\P2_reg1_reg[5]/NET0131 ,
		_w1592_,
		_w6133_,
		_w6537_,
		_w6542_
	);
	LUT4 #(
		.INIT('h7100)
	) name6080 (
		\P2_reg1_reg[5]/NET0131 ,
		_w1592_,
		_w6133_,
		_w6537_,
		_w6543_
	);
	LUT3 #(
		.INIT('h02)
	) name6081 (
		_w6149_,
		_w6543_,
		_w6542_,
		_w6544_
	);
	LUT4 #(
		.INIT('h7100)
	) name6082 (
		\P2_reg2_reg[5]/NET0131 ,
		_w1592_,
		_w6188_,
		_w6532_,
		_w6545_
	);
	LUT4 #(
		.INIT('h008e)
	) name6083 (
		\P2_reg2_reg[5]/NET0131 ,
		_w1592_,
		_w6188_,
		_w6532_,
		_w6546_
	);
	LUT3 #(
		.INIT('h02)
	) name6084 (
		_w2041_,
		_w6546_,
		_w6545_,
		_w6547_
	);
	LUT4 #(
		.INIT('hf4f7)
	) name6085 (
		\P2_addr_reg[6]/NET0131 ,
		_w1505_,
		_w1508_,
		_w1511_,
		_w6548_
	);
	LUT4 #(
		.INIT('h5700)
	) name6086 (
		_w1477_,
		_w1486_,
		_w2080_,
		_w6548_,
		_w6549_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name6087 (
		\P1_state_reg[0]/NET0131 ,
		_w6547_,
		_w6544_,
		_w6549_,
		_w6550_
	);
	LUT3 #(
		.INIT('hba)
	) name6088 (
		_w4977_,
		_w6541_,
		_w6550_,
		_w6551_
	);
	LUT4 #(
		.INIT('h6669)
	) name6089 (
		\P2_IR_reg[7]/NET0131 ,
		\P2_reg2_reg[7]/NET0131 ,
		_w1510_,
		_w1543_,
		_w6552_
	);
	LUT4 #(
		.INIT('h8f00)
	) name6090 (
		_w6228_,
		_w6289_,
		_w6302_,
		_w6552_,
		_w6553_
	);
	LUT4 #(
		.INIT('h0070)
	) name6091 (
		_w6228_,
		_w6289_,
		_w6302_,
		_w6552_,
		_w6554_
	);
	LUT3 #(
		.INIT('h02)
	) name6092 (
		_w6203_,
		_w6554_,
		_w6553_,
		_w6555_
	);
	LUT4 #(
		.INIT('h6669)
	) name6093 (
		\P2_IR_reg[7]/NET0131 ,
		\P2_reg1_reg[7]/NET0131 ,
		_w1510_,
		_w1543_,
		_w6556_
	);
	LUT4 #(
		.INIT('h00ba)
	) name6094 (
		_w6121_,
		_w6211_,
		_w6212_,
		_w6556_,
		_w6557_
	);
	LUT4 #(
		.INIT('h4044)
	) name6095 (
		_w6119_,
		_w6122_,
		_w6211_,
		_w6212_,
		_w6558_
	);
	LUT4 #(
		.INIT('h5600)
	) name6096 (
		\P2_IR_reg[28]/NET0131 ,
		_w1484_,
		_w1507_,
		_w1544_,
		_w6559_
	);
	LUT4 #(
		.INIT('h0080)
	) name6097 (
		_w1483_,
		_w1485_,
		_w1481_,
		_w6559_,
		_w6560_
	);
	LUT4 #(
		.INIT('hfd00)
	) name6098 (
		_w1509_,
		_w6558_,
		_w6557_,
		_w6560_,
		_w6561_
	);
	LUT4 #(
		.INIT('h1555)
	) name6099 (
		\P2_addr_reg[7]/NET0131 ,
		_w1483_,
		_w1485_,
		_w1481_,
		_w6562_
	);
	LUT2 #(
		.INIT('h8)
	) name6100 (
		_w2080_,
		_w6562_,
		_w6563_
	);
	LUT4 #(
		.INIT('haa20)
	) name6101 (
		_w1477_,
		_w6555_,
		_w6561_,
		_w6563_,
		_w6564_
	);
	LUT3 #(
		.INIT('h28)
	) name6102 (
		_w6149_,
		_w6281_,
		_w6556_,
		_w6565_
	);
	LUT3 #(
		.INIT('h28)
	) name6103 (
		_w2041_,
		_w6290_,
		_w6552_,
		_w6566_
	);
	LUT4 #(
		.INIT('hf4f7)
	) name6104 (
		\P2_addr_reg[7]/NET0131 ,
		_w1505_,
		_w1508_,
		_w1544_,
		_w6567_
	);
	LUT4 #(
		.INIT('h5700)
	) name6105 (
		_w1477_,
		_w1486_,
		_w2080_,
		_w6567_,
		_w6568_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name6106 (
		\P1_state_reg[0]/NET0131 ,
		_w6566_,
		_w6565_,
		_w6568_,
		_w6569_
	);
	LUT3 #(
		.INIT('hba)
	) name6107 (
		_w5018_,
		_w6564_,
		_w6569_,
		_w6570_
	);
	LUT4 #(
		.INIT('hc369)
	) name6108 (
		\P2_IR_reg[31]/NET0131 ,
		\P2_IR_reg[8]/NET0131 ,
		\P2_reg2_reg[8]/NET0131 ,
		_w474_,
		_w6571_
	);
	LUT4 #(
		.INIT('h5600)
	) name6109 (
		\P2_IR_reg[28]/NET0131 ,
		_w1484_,
		_w1507_,
		_w1682_,
		_w6572_
	);
	LUT4 #(
		.INIT('hc369)
	) name6110 (
		\P2_IR_reg[31]/NET0131 ,
		\P2_IR_reg[8]/NET0131 ,
		\P2_reg1_reg[8]/NET0131 ,
		_w474_,
		_w6573_
	);
	LUT4 #(
		.INIT('h070d)
	) name6111 (
		_w1509_,
		_w6213_,
		_w6572_,
		_w6573_,
		_w6574_
	);
	LUT4 #(
		.INIT('h7d00)
	) name6112 (
		_w6203_,
		_w6230_,
		_w6571_,
		_w6574_,
		_w6575_
	);
	LUT4 #(
		.INIT('hc4c0)
	) name6113 (
		\P2_addr_reg[8]/NET0131 ,
		_w1477_,
		_w1486_,
		_w2080_,
		_w6576_
	);
	LUT3 #(
		.INIT('hd0)
	) name6114 (
		_w1486_,
		_w6575_,
		_w6576_,
		_w6577_
	);
	LUT4 #(
		.INIT('h5100)
	) name6115 (
		_w6176_,
		_w6179_,
		_w6189_,
		_w6571_,
		_w6578_
	);
	LUT4 #(
		.INIT('h00ae)
	) name6116 (
		_w6176_,
		_w6179_,
		_w6189_,
		_w6571_,
		_w6579_
	);
	LUT3 #(
		.INIT('h02)
	) name6117 (
		_w2041_,
		_w6579_,
		_w6578_,
		_w6580_
	);
	LUT4 #(
		.INIT('hf4f7)
	) name6118 (
		\P2_addr_reg[8]/NET0131 ,
		_w1505_,
		_w1508_,
		_w1682_,
		_w6581_
	);
	LUT4 #(
		.INIT('h5700)
	) name6119 (
		_w1477_,
		_w1486_,
		_w2080_,
		_w6581_,
		_w6582_
	);
	LUT4 #(
		.INIT('hd700)
	) name6120 (
		_w6149_,
		_w6135_,
		_w6573_,
		_w6582_,
		_w6583_
	);
	LUT3 #(
		.INIT('h8a)
	) name6121 (
		\P1_state_reg[0]/NET0131 ,
		_w6580_,
		_w6583_,
		_w6584_
	);
	LUT3 #(
		.INIT('hba)
	) name6122 (
		_w4571_,
		_w6577_,
		_w6584_,
		_w6585_
	);
	LUT4 #(
		.INIT('h6669)
	) name6123 (
		\P2_IR_reg[9]/NET0131 ,
		\P2_reg2_reg[9]/NET0131 ,
		_w1654_,
		_w1669_,
		_w6586_
	);
	LUT4 #(
		.INIT('h00ba)
	) name6124 (
		_w6173_,
		_w6303_,
		_w6304_,
		_w6586_,
		_w6587_
	);
	LUT4 #(
		.INIT('h4500)
	) name6125 (
		_w6173_,
		_w6303_,
		_w6304_,
		_w6586_,
		_w6588_
	);
	LUT3 #(
		.INIT('h02)
	) name6126 (
		_w6203_,
		_w6588_,
		_w6587_,
		_w6589_
	);
	LUT4 #(
		.INIT('h4044)
	) name6127 (
		_w6114_,
		_w6117_,
		_w6118_,
		_w6213_,
		_w6590_
	);
	LUT4 #(
		.INIT('h6669)
	) name6128 (
		\P2_IR_reg[9]/NET0131 ,
		\P2_reg1_reg[9]/NET0131 ,
		_w1654_,
		_w1669_,
		_w6591_
	);
	LUT4 #(
		.INIT('h00d4)
	) name6129 (
		\P2_reg1_reg[8]/NET0131 ,
		_w1682_,
		_w6213_,
		_w6591_,
		_w6592_
	);
	LUT4 #(
		.INIT('h5600)
	) name6130 (
		\P2_IR_reg[28]/NET0131 ,
		_w1484_,
		_w1507_,
		_w1670_,
		_w6593_
	);
	LUT4 #(
		.INIT('h0080)
	) name6131 (
		_w1483_,
		_w1485_,
		_w1481_,
		_w6593_,
		_w6594_
	);
	LUT4 #(
		.INIT('hfd00)
	) name6132 (
		_w1509_,
		_w6592_,
		_w6590_,
		_w6594_,
		_w6595_
	);
	LUT4 #(
		.INIT('h1555)
	) name6133 (
		\P2_addr_reg[9]/NET0131 ,
		_w1483_,
		_w1485_,
		_w1481_,
		_w6596_
	);
	LUT2 #(
		.INIT('h8)
	) name6134 (
		_w2080_,
		_w6596_,
		_w6597_
	);
	LUT4 #(
		.INIT('haa20)
	) name6135 (
		_w1477_,
		_w6589_,
		_w6595_,
		_w6597_,
		_w6598_
	);
	LUT3 #(
		.INIT('h28)
	) name6136 (
		_w2041_,
		_w6292_,
		_w6586_,
		_w6599_
	);
	LUT4 #(
		.INIT('hf4f7)
	) name6137 (
		\P2_addr_reg[9]/NET0131 ,
		_w1505_,
		_w1508_,
		_w1670_,
		_w6600_
	);
	LUT4 #(
		.INIT('h5700)
	) name6138 (
		_w1477_,
		_w1486_,
		_w2080_,
		_w6600_,
		_w6601_
	);
	LUT4 #(
		.INIT('hd700)
	) name6139 (
		_w6149_,
		_w6283_,
		_w6591_,
		_w6601_,
		_w6602_
	);
	LUT3 #(
		.INIT('h8a)
	) name6140 (
		\P1_state_reg[0]/NET0131 ,
		_w6599_,
		_w6602_,
		_w6603_
	);
	LUT3 #(
		.INIT('hba)
	) name6141 (
		_w4243_,
		_w6598_,
		_w6603_,
		_w6604_
	);
	LUT4 #(
		.INIT('h1555)
	) name6142 (
		\P2_addr_reg[5]/NET0131 ,
		_w1483_,
		_w1485_,
		_w1481_,
		_w6605_
	);
	LUT2 #(
		.INIT('h6)
	) name6143 (
		\P2_reg2_reg[5]/NET0131 ,
		_w1592_,
		_w6606_
	);
	LUT4 #(
		.INIT('h0110)
	) name6144 (
		_w1505_,
		_w1508_,
		_w6228_,
		_w6606_,
		_w6607_
	);
	LUT2 #(
		.INIT('h4)
	) name6145 (
		_w6125_,
		_w6211_,
		_w6608_
	);
	LUT2 #(
		.INIT('h6)
	) name6146 (
		\P2_reg1_reg[5]/NET0131 ,
		_w1592_,
		_w6609_
	);
	LUT4 #(
		.INIT('h222b)
	) name6147 (
		\P2_reg1_reg[4]/NET0131 ,
		_w1601_,
		_w6129_,
		_w6209_,
		_w6610_
	);
	LUT4 #(
		.INIT('h2220)
	) name6148 (
		_w1505_,
		_w1508_,
		_w6609_,
		_w6610_,
		_w6611_
	);
	LUT4 #(
		.INIT('h0056)
	) name6149 (
		\P2_IR_reg[28]/NET0131 ,
		_w1484_,
		_w1507_,
		_w1592_,
		_w6612_
	);
	LUT4 #(
		.INIT('h0080)
	) name6150 (
		_w1483_,
		_w1485_,
		_w1481_,
		_w6612_,
		_w6613_
	);
	LUT4 #(
		.INIT('h0b00)
	) name6151 (
		_w6608_,
		_w6611_,
		_w6607_,
		_w6613_,
		_w6614_
	);
	LUT3 #(
		.INIT('ha8)
	) name6152 (
		_w6202_,
		_w6605_,
		_w6614_,
		_w6615_
	);
	LUT4 #(
		.INIT('h0440)
	) name6153 (
		_w1505_,
		_w1508_,
		_w6188_,
		_w6606_,
		_w6616_
	);
	LUT4 #(
		.INIT('h0880)
	) name6154 (
		_w1505_,
		_w1508_,
		_w6133_,
		_w6609_,
		_w6617_
	);
	LUT4 #(
		.INIT('hf7f4)
	) name6155 (
		\P2_addr_reg[5]/NET0131 ,
		_w1505_,
		_w1508_,
		_w1592_,
		_w6618_
	);
	LUT4 #(
		.INIT('h5700)
	) name6156 (
		_w1477_,
		_w1486_,
		_w2080_,
		_w6618_,
		_w6619_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name6157 (
		\P1_state_reg[0]/NET0131 ,
		_w6617_,
		_w6616_,
		_w6619_,
		_w6620_
	);
	LUT3 #(
		.INIT('hba)
	) name6158 (
		_w4973_,
		_w6615_,
		_w6620_,
		_w6621_
	);
	LUT2 #(
		.INIT('h2)
	) name6159 (
		_w537_,
		_w540_,
		_w6622_
	);
	LUT2 #(
		.INIT('h8)
	) name6160 (
		\P1_IR_reg[0]/NET0131 ,
		\P1_reg1_reg[0]/NET0131 ,
		_w6623_
	);
	LUT2 #(
		.INIT('h6)
	) name6161 (
		\P1_IR_reg[0]/NET0131 ,
		\P1_reg1_reg[0]/NET0131 ,
		_w6624_
	);
	LUT2 #(
		.INIT('h8)
	) name6162 (
		\P1_IR_reg[0]/NET0131 ,
		\P1_reg2_reg[0]/NET0131 ,
		_w6625_
	);
	LUT2 #(
		.INIT('h6)
	) name6163 (
		\P1_IR_reg[0]/NET0131 ,
		\P1_reg2_reg[0]/NET0131 ,
		_w6626_
	);
	LUT4 #(
		.INIT('h57df)
	) name6164 (
		_w537_,
		_w540_,
		_w6624_,
		_w6626_,
		_w6627_
	);
	LUT4 #(
		.INIT('h8882)
	) name6165 (
		\P1_IR_reg[0]/NET0131 ,
		\P1_IR_reg[28]/NET0131 ,
		_w513_,
		_w536_,
		_w6628_
	);
	LUT4 #(
		.INIT('h0080)
	) name6166 (
		_w519_,
		_w522_,
		_w517_,
		_w6628_,
		_w6629_
	);
	LUT2 #(
		.INIT('h8)
	) name6167 (
		_w6627_,
		_w6629_,
		_w6630_
	);
	LUT4 #(
		.INIT('h1555)
	) name6168 (
		\P1_addr_reg[2]/NET0131 ,
		_w519_,
		_w522_,
		_w517_,
		_w6631_
	);
	LUT3 #(
		.INIT('h80)
	) name6169 (
		_w1104_,
		_w1106_,
		_w6631_,
		_w6632_
	);
	LUT3 #(
		.INIT('h54)
	) name6170 (
		_w510_,
		_w6630_,
		_w6632_,
		_w6633_
	);
	LUT4 #(
		.INIT('h2333)
	) name6171 (
		_w510_,
		_w524_,
		_w1104_,
		_w1106_,
		_w6634_
	);
	LUT2 #(
		.INIT('h6)
	) name6172 (
		\P1_reg2_reg[2]/NET0131 ,
		_w852_,
		_w6635_
	);
	LUT3 #(
		.INIT('hb2)
	) name6173 (
		\P1_reg2_reg[1]/NET0131 ,
		_w859_,
		_w6625_,
		_w6636_
	);
	LUT2 #(
		.INIT('h6)
	) name6174 (
		_w6635_,
		_w6636_,
		_w6637_
	);
	LUT4 #(
		.INIT('h3dfd)
	) name6175 (
		\P1_addr_reg[2]/NET0131 ,
		_w537_,
		_w540_,
		_w6637_,
		_w6638_
	);
	LUT2 #(
		.INIT('h6)
	) name6176 (
		\P1_reg1_reg[2]/NET0131 ,
		_w852_,
		_w6639_
	);
	LUT3 #(
		.INIT('hb2)
	) name6177 (
		\P1_reg1_reg[1]/NET0131 ,
		_w859_,
		_w6623_,
		_w6640_
	);
	LUT2 #(
		.INIT('h6)
	) name6178 (
		_w6639_,
		_w6640_,
		_w6641_
	);
	LUT2 #(
		.INIT('h4)
	) name6179 (
		_w537_,
		_w540_,
		_w6642_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name6180 (
		_w537_,
		_w540_,
		_w852_,
		_w6641_,
		_w6643_
	);
	LUT2 #(
		.INIT('h8)
	) name6181 (
		_w6638_,
		_w6643_,
		_w6644_
	);
	LUT2 #(
		.INIT('h8)
	) name6182 (
		_w6634_,
		_w6644_,
		_w6645_
	);
	LUT4 #(
		.INIT('h222e)
	) name6183 (
		\P1_reg3_reg[2]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w6633_,
		_w6645_,
		_w6646_
	);
	LUT4 #(
		.INIT('h1555)
	) name6184 (
		\P1_addr_reg[4]/NET0131 ,
		_w519_,
		_w522_,
		_w517_,
		_w6647_
	);
	LUT3 #(
		.INIT('h80)
	) name6185 (
		_w1104_,
		_w1106_,
		_w6647_,
		_w6648_
	);
	LUT3 #(
		.INIT('h54)
	) name6186 (
		_w510_,
		_w6630_,
		_w6648_,
		_w6649_
	);
	LUT4 #(
		.INIT('h3c96)
	) name6187 (
		\P1_IR_reg[31]/NET0131 ,
		\P1_IR_reg[4]/NET0131 ,
		\P1_reg1_reg[4]/NET0131 ,
		_w500_,
		_w6650_
	);
	LUT3 #(
		.INIT('h21)
	) name6188 (
		\P1_IR_reg[3]/NET0131 ,
		\P1_reg1_reg[3]/NET0131 ,
		_w878_,
		_w6651_
	);
	LUT3 #(
		.INIT('h48)
	) name6189 (
		\P1_IR_reg[3]/NET0131 ,
		\P1_reg1_reg[3]/NET0131 ,
		_w878_,
		_w6652_
	);
	LUT4 #(
		.INIT('h0017)
	) name6190 (
		\P1_reg1_reg[2]/NET0131 ,
		_w852_,
		_w6640_,
		_w6652_,
		_w6653_
	);
	LUT3 #(
		.INIT('ha9)
	) name6191 (
		_w6650_,
		_w6651_,
		_w6653_,
		_w6654_
	);
	LUT4 #(
		.INIT('hf1fd)
	) name6192 (
		\P1_addr_reg[4]/NET0131 ,
		_w537_,
		_w540_,
		_w6654_,
		_w6655_
	);
	LUT4 #(
		.INIT('h3c96)
	) name6193 (
		\P1_IR_reg[31]/NET0131 ,
		\P1_IR_reg[4]/NET0131 ,
		\P1_reg2_reg[4]/NET0131 ,
		_w500_,
		_w6656_
	);
	LUT3 #(
		.INIT('h21)
	) name6194 (
		\P1_IR_reg[3]/NET0131 ,
		\P1_reg2_reg[3]/NET0131 ,
		_w878_,
		_w6657_
	);
	LUT3 #(
		.INIT('h48)
	) name6195 (
		\P1_IR_reg[3]/NET0131 ,
		\P1_reg2_reg[3]/NET0131 ,
		_w878_,
		_w6658_
	);
	LUT4 #(
		.INIT('h0017)
	) name6196 (
		\P1_reg2_reg[2]/NET0131 ,
		_w852_,
		_w6636_,
		_w6658_,
		_w6659_
	);
	LUT3 #(
		.INIT('ha9)
	) name6197 (
		_w6656_,
		_w6657_,
		_w6659_,
		_w6660_
	);
	LUT4 #(
		.INIT('h73fb)
	) name6198 (
		_w537_,
		_w540_,
		_w889_,
		_w6660_,
		_w6661_
	);
	LUT2 #(
		.INIT('h8)
	) name6199 (
		_w6655_,
		_w6661_,
		_w6662_
	);
	LUT2 #(
		.INIT('h8)
	) name6200 (
		_w6634_,
		_w6662_,
		_w6663_
	);
	LUT4 #(
		.INIT('h222e)
	) name6201 (
		\P1_reg3_reg[4]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w6649_,
		_w6663_,
		_w6664_
	);
	LUT3 #(
		.INIT('h75)
	) name6202 (
		\P1_state_reg[0]/NET0131 ,
		_w541_,
		_w6634_,
		_w6665_
	);
	LUT4 #(
		.INIT('h0507)
	) name6203 (
		_w1477_,
		_w1486_,
		_w1509_,
		_w2080_,
		_w6666_
	);
	LUT2 #(
		.INIT('hd)
	) name6204 (
		\P1_state_reg[0]/NET0131 ,
		_w6666_,
		_w6667_
	);
	LUT2 #(
		.INIT('h8)
	) name6205 (
		\P1_state_reg[0]/NET0131 ,
		_w6634_,
		_w6668_
	);
	LUT2 #(
		.INIT('h1)
	) name6206 (
		\P1_reg2_reg[11]/NET0131 ,
		_w802_,
		_w6669_
	);
	LUT2 #(
		.INIT('h8)
	) name6207 (
		\P1_reg2_reg[11]/NET0131 ,
		_w802_,
		_w6670_
	);
	LUT2 #(
		.INIT('h6)
	) name6208 (
		\P1_reg2_reg[11]/NET0131 ,
		_w802_,
		_w6671_
	);
	LUT4 #(
		.INIT('ha060)
	) name6209 (
		\P1_IR_reg[10]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		\P1_reg2_reg[10]/NET0131 ,
		_w503_,
		_w6672_
	);
	LUT2 #(
		.INIT('h8)
	) name6210 (
		\P1_reg2_reg[9]/NET0131 ,
		_w840_,
		_w6673_
	);
	LUT3 #(
		.INIT('h21)
	) name6211 (
		\P1_IR_reg[6]/NET0131 ,
		\P1_reg2_reg[6]/NET0131 ,
		_w915_,
		_w6674_
	);
	LUT3 #(
		.INIT('h48)
	) name6212 (
		\P1_IR_reg[6]/NET0131 ,
		\P1_reg2_reg[6]/NET0131 ,
		_w915_,
		_w6675_
	);
	LUT4 #(
		.INIT('h222b)
	) name6213 (
		\P1_reg2_reg[4]/NET0131 ,
		_w889_,
		_w6657_,
		_w6659_,
		_w6676_
	);
	LUT3 #(
		.INIT('he8)
	) name6214 (
		\P1_reg2_reg[5]/NET0131 ,
		_w937_,
		_w6676_,
		_w6677_
	);
	LUT4 #(
		.INIT('h0107)
	) name6215 (
		\P1_reg2_reg[5]/NET0131 ,
		_w937_,
		_w6675_,
		_w6676_,
		_w6678_
	);
	LUT4 #(
		.INIT('h888e)
	) name6216 (
		\P1_reg2_reg[7]/NET0131 ,
		_w917_,
		_w6674_,
		_w6678_,
		_w6679_
	);
	LUT4 #(
		.INIT('h0107)
	) name6217 (
		\P1_reg2_reg[8]/NET0131 ,
		_w906_,
		_w6673_,
		_w6679_,
		_w6680_
	);
	LUT4 #(
		.INIT('h0509)
	) name6218 (
		\P1_IR_reg[10]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		\P1_reg2_reg[10]/NET0131 ,
		_w503_,
		_w6681_
	);
	LUT2 #(
		.INIT('h1)
	) name6219 (
		\P1_reg2_reg[9]/NET0131 ,
		_w840_,
		_w6682_
	);
	LUT3 #(
		.INIT('h0e)
	) name6220 (
		\P1_reg2_reg[9]/NET0131 ,
		_w840_,
		_w6681_,
		_w6683_
	);
	LUT4 #(
		.INIT('h1011)
	) name6221 (
		_w6671_,
		_w6672_,
		_w6680_,
		_w6683_,
		_w6684_
	);
	LUT4 #(
		.INIT('h8a88)
	) name6222 (
		_w6671_,
		_w6672_,
		_w6680_,
		_w6683_,
		_w6685_
	);
	LUT3 #(
		.INIT('h02)
	) name6223 (
		_w1290_,
		_w6685_,
		_w6684_,
		_w6686_
	);
	LUT2 #(
		.INIT('h1)
	) name6224 (
		\P1_reg1_reg[11]/NET0131 ,
		_w802_,
		_w6687_
	);
	LUT2 #(
		.INIT('h6)
	) name6225 (
		\P1_reg1_reg[11]/NET0131 ,
		_w802_,
		_w6688_
	);
	LUT4 #(
		.INIT('ha060)
	) name6226 (
		\P1_IR_reg[10]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		\P1_reg1_reg[10]/NET0131 ,
		_w503_,
		_w6689_
	);
	LUT4 #(
		.INIT('h0509)
	) name6227 (
		\P1_IR_reg[10]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		\P1_reg1_reg[10]/NET0131 ,
		_w503_,
		_w6690_
	);
	LUT4 #(
		.INIT('h0309)
	) name6228 (
		\P1_IR_reg[31]/NET0131 ,
		\P1_IR_reg[8]/NET0131 ,
		\P1_reg1_reg[8]/NET0131 ,
		_w839_,
		_w6691_
	);
	LUT4 #(
		.INIT('hc060)
	) name6229 (
		\P1_IR_reg[31]/NET0131 ,
		\P1_IR_reg[8]/NET0131 ,
		\P1_reg1_reg[8]/NET0131 ,
		_w839_,
		_w6692_
	);
	LUT4 #(
		.INIT('h2221)
	) name6230 (
		\P1_IR_reg[7]/NET0131 ,
		\P1_reg1_reg[7]/NET0131 ,
		_w915_,
		_w916_,
		_w6693_
	);
	LUT3 #(
		.INIT('h21)
	) name6231 (
		\P1_IR_reg[6]/NET0131 ,
		\P1_reg1_reg[6]/NET0131 ,
		_w915_,
		_w6694_
	);
	LUT4 #(
		.INIT('h222b)
	) name6232 (
		\P1_reg1_reg[4]/NET0131 ,
		_w889_,
		_w6651_,
		_w6653_,
		_w6695_
	);
	LUT4 #(
		.INIT('h0e08)
	) name6233 (
		\P1_reg1_reg[5]/NET0131 ,
		_w937_,
		_w6694_,
		_w6695_,
		_w6696_
	);
	LUT4 #(
		.INIT('h4448)
	) name6234 (
		\P1_IR_reg[7]/NET0131 ,
		\P1_reg1_reg[7]/NET0131 ,
		_w915_,
		_w916_,
		_w6697_
	);
	LUT3 #(
		.INIT('h48)
	) name6235 (
		\P1_IR_reg[6]/NET0131 ,
		\P1_reg1_reg[6]/NET0131 ,
		_w915_,
		_w6698_
	);
	LUT2 #(
		.INIT('h1)
	) name6236 (
		_w6697_,
		_w6698_,
		_w6699_
	);
	LUT3 #(
		.INIT('h45)
	) name6237 (
		_w6693_,
		_w6696_,
		_w6699_,
		_w6700_
	);
	LUT4 #(
		.INIT('h4544)
	) name6238 (
		_w6692_,
		_w6693_,
		_w6696_,
		_w6699_,
		_w6701_
	);
	LUT4 #(
		.INIT('h888e)
	) name6239 (
		\P1_reg1_reg[9]/NET0131 ,
		_w840_,
		_w6691_,
		_w6701_,
		_w6702_
	);
	LUT3 #(
		.INIT('h17)
	) name6240 (
		\P1_reg1_reg[10]/NET0131 ,
		_w825_,
		_w6702_,
		_w6703_
	);
	LUT4 #(
		.INIT('hcdfd)
	) name6241 (
		\P1_addr_reg[11]/NET0131 ,
		_w537_,
		_w540_,
		_w802_,
		_w6704_
	);
	LUT4 #(
		.INIT('h7d00)
	) name6242 (
		_w6622_,
		_w6688_,
		_w6703_,
		_w6704_,
		_w6705_
	);
	LUT4 #(
		.INIT('h8000)
	) name6243 (
		\P1_addr_reg[11]/NET0131 ,
		_w1104_,
		_w1106_,
		_w3443_,
		_w6706_
	);
	LUT2 #(
		.INIT('h1)
	) name6244 (
		_w4451_,
		_w6706_,
		_w6707_
	);
	LUT4 #(
		.INIT('h8aff)
	) name6245 (
		_w6668_,
		_w6686_,
		_w6705_,
		_w6707_,
		_w6708_
	);
	LUT2 #(
		.INIT('h2)
	) name6246 (
		\P1_reg3_reg[0]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w6709_
	);
	LUT4 #(
		.INIT('hbf00)
	) name6247 (
		\P1_addr_reg[0]/NET0131 ,
		_w1104_,
		_w1106_,
		_w3443_,
		_w6710_
	);
	LUT2 #(
		.INIT('h1)
	) name6248 (
		_w1294_,
		_w6710_,
		_w6711_
	);
	LUT4 #(
		.INIT('h1555)
	) name6249 (
		_w541_,
		_w1104_,
		_w1106_,
		_w3443_,
		_w6712_
	);
	LUT2 #(
		.INIT('h8)
	) name6250 (
		_w540_,
		_w6628_,
		_w6713_
	);
	LUT2 #(
		.INIT('h2)
	) name6251 (
		_w6627_,
		_w6713_,
		_w6714_
	);
	LUT3 #(
		.INIT('hd0)
	) name6252 (
		\P1_addr_reg[0]/NET0131 ,
		_w6712_,
		_w6714_,
		_w6715_
	);
	LUT3 #(
		.INIT('hab)
	) name6253 (
		_w6709_,
		_w6711_,
		_w6715_,
		_w6716_
	);
	LUT4 #(
		.INIT('hbf00)
	) name6254 (
		\P1_addr_reg[10]/NET0131 ,
		_w1104_,
		_w1106_,
		_w3443_,
		_w6717_
	);
	LUT2 #(
		.INIT('h1)
	) name6255 (
		_w1294_,
		_w6717_,
		_w6718_
	);
	LUT3 #(
		.INIT('h10)
	) name6256 (
		_w6672_,
		_w6680_,
		_w6683_,
		_w6719_
	);
	LUT4 #(
		.INIT('h5a96)
	) name6257 (
		\P1_IR_reg[10]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		\P1_reg2_reg[10]/NET0131 ,
		_w503_,
		_w6720_
	);
	LUT4 #(
		.INIT('haa02)
	) name6258 (
		_w1290_,
		_w6680_,
		_w6682_,
		_w6720_,
		_w6721_
	);
	LUT4 #(
		.INIT('h5a96)
	) name6259 (
		\P1_IR_reg[10]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		\P1_reg1_reg[10]/NET0131 ,
		_w503_,
		_w6722_
	);
	LUT4 #(
		.INIT('hcdfd)
	) name6260 (
		\P1_addr_reg[10]/NET0131 ,
		_w537_,
		_w540_,
		_w825_,
		_w6723_
	);
	LUT4 #(
		.INIT('hd700)
	) name6261 (
		_w6622_,
		_w6702_,
		_w6722_,
		_w6723_,
		_w6724_
	);
	LUT4 #(
		.INIT('h1055)
	) name6262 (
		_w6718_,
		_w6719_,
		_w6721_,
		_w6724_,
		_w6725_
	);
	LUT4 #(
		.INIT('h8000)
	) name6263 (
		\P1_addr_reg[10]/NET0131 ,
		_w1104_,
		_w1106_,
		_w3443_,
		_w6726_
	);
	LUT2 #(
		.INIT('h1)
	) name6264 (
		_w4098_,
		_w6726_,
		_w6727_
	);
	LUT2 #(
		.INIT('hb)
	) name6265 (
		_w6725_,
		_w6727_,
		_w6728_
	);
	LUT4 #(
		.INIT('hbf00)
	) name6266 (
		\P1_addr_reg[12]/NET0131 ,
		_w1104_,
		_w1106_,
		_w3443_,
		_w6729_
	);
	LUT2 #(
		.INIT('h1)
	) name6267 (
		_w1294_,
		_w6729_,
		_w6730_
	);
	LUT2 #(
		.INIT('h1)
	) name6268 (
		\P1_reg2_reg[12]/NET0131 ,
		_w812_,
		_w6731_
	);
	LUT2 #(
		.INIT('h6)
	) name6269 (
		\P1_reg2_reg[12]/NET0131 ,
		_w812_,
		_w6732_
	);
	LUT4 #(
		.INIT('h4544)
	) name6270 (
		_w6669_,
		_w6672_,
		_w6680_,
		_w6683_,
		_w6733_
	);
	LUT4 #(
		.INIT('h0a28)
	) name6271 (
		_w1290_,
		_w6670_,
		_w6732_,
		_w6733_,
		_w6734_
	);
	LUT2 #(
		.INIT('h1)
	) name6272 (
		\P1_reg1_reg[12]/NET0131 ,
		_w812_,
		_w6735_
	);
	LUT2 #(
		.INIT('h6)
	) name6273 (
		\P1_reg1_reg[12]/NET0131 ,
		_w812_,
		_w6736_
	);
	LUT3 #(
		.INIT('h07)
	) name6274 (
		\P1_reg1_reg[11]/NET0131 ,
		_w802_,
		_w6689_,
		_w6737_
	);
	LUT4 #(
		.INIT('h1055)
	) name6275 (
		_w6687_,
		_w6690_,
		_w6702_,
		_w6737_,
		_w6738_
	);
	LUT3 #(
		.INIT('h40)
	) name6276 (
		_w537_,
		_w540_,
		_w812_,
		_w6739_
	);
	LUT3 #(
		.INIT('h0d)
	) name6277 (
		\P1_addr_reg[12]/NET0131 ,
		_w6712_,
		_w6739_,
		_w6740_
	);
	LUT4 #(
		.INIT('hd700)
	) name6278 (
		_w6622_,
		_w6736_,
		_w6738_,
		_w6740_,
		_w6741_
	);
	LUT4 #(
		.INIT('hbabb)
	) name6279 (
		_w3464_,
		_w6730_,
		_w6734_,
		_w6741_,
		_w6742_
	);
	LUT2 #(
		.INIT('h1)
	) name6280 (
		\P1_reg2_reg[13]/NET0131 ,
		_w756_,
		_w6743_
	);
	LUT2 #(
		.INIT('h6)
	) name6281 (
		\P1_reg2_reg[13]/NET0131 ,
		_w756_,
		_w6744_
	);
	LUT4 #(
		.INIT('h135f)
	) name6282 (
		\P1_reg2_reg[11]/NET0131 ,
		\P1_reg2_reg[12]/NET0131 ,
		_w802_,
		_w812_,
		_w6745_
	);
	LUT4 #(
		.INIT('h0b0a)
	) name6283 (
		_w6731_,
		_w6733_,
		_w6744_,
		_w6745_,
		_w6746_
	);
	LUT4 #(
		.INIT('h4050)
	) name6284 (
		_w6731_,
		_w6733_,
		_w6744_,
		_w6745_,
		_w6747_
	);
	LUT3 #(
		.INIT('h02)
	) name6285 (
		_w1290_,
		_w6747_,
		_w6746_,
		_w6748_
	);
	LUT2 #(
		.INIT('h8)
	) name6286 (
		\P1_reg1_reg[13]/NET0131 ,
		_w756_,
		_w6749_
	);
	LUT2 #(
		.INIT('h1)
	) name6287 (
		\P1_reg1_reg[13]/NET0131 ,
		_w756_,
		_w6750_
	);
	LUT2 #(
		.INIT('h6)
	) name6288 (
		\P1_reg1_reg[13]/NET0131 ,
		_w756_,
		_w6751_
	);
	LUT4 #(
		.INIT('h0e08)
	) name6289 (
		\P1_reg1_reg[10]/NET0131 ,
		_w825_,
		_w6687_,
		_w6702_,
		_w6752_
	);
	LUT4 #(
		.INIT('h135f)
	) name6290 (
		\P1_reg1_reg[11]/NET0131 ,
		\P1_reg1_reg[12]/NET0131 ,
		_w802_,
		_w812_,
		_w6753_
	);
	LUT3 #(
		.INIT('h45)
	) name6291 (
		_w6735_,
		_w6752_,
		_w6753_,
		_w6754_
	);
	LUT4 #(
		.INIT('hcdfd)
	) name6292 (
		\P1_addr_reg[13]/NET0131 ,
		_w537_,
		_w540_,
		_w756_,
		_w6755_
	);
	LUT4 #(
		.INIT('hd700)
	) name6293 (
		_w6622_,
		_w6751_,
		_w6754_,
		_w6755_,
		_w6756_
	);
	LUT4 #(
		.INIT('h8000)
	) name6294 (
		\P1_addr_reg[13]/NET0131 ,
		_w1104_,
		_w1106_,
		_w3443_,
		_w6757_
	);
	LUT2 #(
		.INIT('h1)
	) name6295 (
		_w4469_,
		_w6757_,
		_w6758_
	);
	LUT4 #(
		.INIT('h8aff)
	) name6296 (
		_w6668_,
		_w6748_,
		_w6756_,
		_w6758_,
		_w6759_
	);
	LUT4 #(
		.INIT('hbf00)
	) name6297 (
		\P1_addr_reg[14]/NET0131 ,
		_w1104_,
		_w1106_,
		_w3443_,
		_w6760_
	);
	LUT2 #(
		.INIT('h1)
	) name6298 (
		_w1294_,
		_w6760_,
		_w6761_
	);
	LUT4 #(
		.INIT('h153f)
	) name6299 (
		\P1_reg2_reg[12]/NET0131 ,
		\P1_reg2_reg[13]/NET0131 ,
		_w756_,
		_w812_,
		_w6762_
	);
	LUT4 #(
		.INIT('hcd00)
	) name6300 (
		_w6670_,
		_w6731_,
		_w6733_,
		_w6762_,
		_w6763_
	);
	LUT2 #(
		.INIT('h2)
	) name6301 (
		\P1_reg2_reg[14]/NET0131 ,
		_w765_,
		_w6764_
	);
	LUT2 #(
		.INIT('h4)
	) name6302 (
		\P1_reg2_reg[14]/NET0131 ,
		_w765_,
		_w6765_
	);
	LUT2 #(
		.INIT('h9)
	) name6303 (
		\P1_reg2_reg[14]/NET0131 ,
		_w765_,
		_w6766_
	);
	LUT4 #(
		.INIT('ha802)
	) name6304 (
		_w1290_,
		_w6743_,
		_w6763_,
		_w6766_,
		_w6767_
	);
	LUT4 #(
		.INIT('h153f)
	) name6305 (
		\P1_reg1_reg[12]/NET0131 ,
		\P1_reg1_reg[13]/NET0131 ,
		_w756_,
		_w812_,
		_w6768_
	);
	LUT4 #(
		.INIT('h040f)
	) name6306 (
		_w6735_,
		_w6738_,
		_w6750_,
		_w6768_,
		_w6769_
	);
	LUT2 #(
		.INIT('h2)
	) name6307 (
		\P1_reg1_reg[14]/NET0131 ,
		_w765_,
		_w6770_
	);
	LUT2 #(
		.INIT('h4)
	) name6308 (
		\P1_reg1_reg[14]/NET0131 ,
		_w765_,
		_w6771_
	);
	LUT2 #(
		.INIT('h9)
	) name6309 (
		\P1_reg1_reg[14]/NET0131 ,
		_w765_,
		_w6772_
	);
	LUT4 #(
		.INIT('hfdcd)
	) name6310 (
		\P1_addr_reg[14]/NET0131 ,
		_w537_,
		_w540_,
		_w765_,
		_w6773_
	);
	LUT4 #(
		.INIT('hd700)
	) name6311 (
		_w6622_,
		_w6769_,
		_w6772_,
		_w6773_,
		_w6774_
	);
	LUT4 #(
		.INIT('h8000)
	) name6312 (
		\P1_addr_reg[14]/NET0131 ,
		_w1104_,
		_w1106_,
		_w3443_,
		_w6775_
	);
	LUT2 #(
		.INIT('h1)
	) name6313 (
		_w4118_,
		_w6775_,
		_w6776_
	);
	LUT4 #(
		.INIT('h45ff)
	) name6314 (
		_w6761_,
		_w6767_,
		_w6774_,
		_w6776_,
		_w6777_
	);
	LUT4 #(
		.INIT('hbf00)
	) name6315 (
		\P1_addr_reg[15]/NET0131 ,
		_w1104_,
		_w1106_,
		_w3443_,
		_w6778_
	);
	LUT2 #(
		.INIT('h1)
	) name6316 (
		_w1294_,
		_w6778_,
		_w6779_
	);
	LUT3 #(
		.INIT('h48)
	) name6317 (
		\P1_IR_reg[15]/NET0131 ,
		\P1_reg1_reg[15]/NET0131 ,
		_w777_,
		_w6780_
	);
	LUT3 #(
		.INIT('h21)
	) name6318 (
		\P1_IR_reg[15]/NET0131 ,
		\P1_reg1_reg[15]/NET0131 ,
		_w777_,
		_w6781_
	);
	LUT3 #(
		.INIT('h96)
	) name6319 (
		\P1_IR_reg[15]/NET0131 ,
		\P1_reg1_reg[15]/NET0131 ,
		_w777_,
		_w6782_
	);
	LUT4 #(
		.INIT('h2322)
	) name6320 (
		_w6735_,
		_w6749_,
		_w6752_,
		_w6753_,
		_w6783_
	);
	LUT4 #(
		.INIT('hc8fa)
	) name6321 (
		\P1_reg1_reg[13]/NET0131 ,
		\P1_reg1_reg[14]/NET0131 ,
		_w756_,
		_w765_,
		_w6784_
	);
	LUT4 #(
		.INIT('h8c88)
	) name6322 (
		_w6770_,
		_w6782_,
		_w6783_,
		_w6784_,
		_w6785_
	);
	LUT4 #(
		.INIT('h1011)
	) name6323 (
		_w6770_,
		_w6782_,
		_w6783_,
		_w6784_,
		_w6786_
	);
	LUT3 #(
		.INIT('h02)
	) name6324 (
		_w6622_,
		_w6786_,
		_w6785_,
		_w6787_
	);
	LUT3 #(
		.INIT('h48)
	) name6325 (
		\P1_IR_reg[15]/NET0131 ,
		\P1_reg2_reg[15]/NET0131 ,
		_w777_,
		_w6788_
	);
	LUT3 #(
		.INIT('h21)
	) name6326 (
		\P1_IR_reg[15]/NET0131 ,
		\P1_reg2_reg[15]/NET0131 ,
		_w777_,
		_w6789_
	);
	LUT3 #(
		.INIT('h96)
	) name6327 (
		\P1_IR_reg[15]/NET0131 ,
		\P1_reg2_reg[15]/NET0131 ,
		_w777_,
		_w6790_
	);
	LUT4 #(
		.INIT('hc8fa)
	) name6328 (
		\P1_reg2_reg[13]/NET0131 ,
		\P1_reg2_reg[14]/NET0131 ,
		_w756_,
		_w765_,
		_w6791_
	);
	LUT4 #(
		.INIT('h4500)
	) name6329 (
		_w6731_,
		_w6733_,
		_w6745_,
		_w6791_,
		_w6792_
	);
	LUT4 #(
		.INIT('h7f13)
	) name6330 (
		\P1_reg2_reg[13]/NET0131 ,
		\P1_reg2_reg[14]/NET0131 ,
		_w756_,
		_w765_,
		_w6793_
	);
	LUT4 #(
		.INIT('h2822)
	) name6331 (
		_w1290_,
		_w6790_,
		_w6792_,
		_w6793_,
		_w6794_
	);
	LUT3 #(
		.INIT('h04)
	) name6332 (
		_w537_,
		_w540_,
		_w778_,
		_w6795_
	);
	LUT3 #(
		.INIT('h0d)
	) name6333 (
		\P1_addr_reg[15]/NET0131 ,
		_w6712_,
		_w6795_,
		_w6796_
	);
	LUT2 #(
		.INIT('h4)
	) name6334 (
		_w6794_,
		_w6796_,
		_w6797_
	);
	LUT4 #(
		.INIT('hbabb)
	) name6335 (
		_w4137_,
		_w6779_,
		_w6787_,
		_w6797_,
		_w6798_
	);
	LUT4 #(
		.INIT('hbf00)
	) name6336 (
		\P1_addr_reg[16]/NET0131 ,
		_w1104_,
		_w1106_,
		_w3443_,
		_w6799_
	);
	LUT2 #(
		.INIT('h1)
	) name6337 (
		_w1294_,
		_w6799_,
		_w6800_
	);
	LUT2 #(
		.INIT('h1)
	) name6338 (
		_w6764_,
		_w6788_,
		_w6801_
	);
	LUT4 #(
		.INIT('hfe00)
	) name6339 (
		_w6743_,
		_w6763_,
		_w6765_,
		_w6801_,
		_w6802_
	);
	LUT4 #(
		.INIT('ha060)
	) name6340 (
		\P1_IR_reg[16]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		\P1_reg2_reg[16]/NET0131 ,
		_w648_,
		_w6803_
	);
	LUT4 #(
		.INIT('h0509)
	) name6341 (
		\P1_IR_reg[16]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		\P1_reg2_reg[16]/NET0131 ,
		_w648_,
		_w6804_
	);
	LUT4 #(
		.INIT('h5a96)
	) name6342 (
		\P1_IR_reg[16]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		\P1_reg2_reg[16]/NET0131 ,
		_w648_,
		_w6805_
	);
	LUT4 #(
		.INIT('ha802)
	) name6343 (
		_w1290_,
		_w6789_,
		_w6802_,
		_w6805_,
		_w6806_
	);
	LUT2 #(
		.INIT('h1)
	) name6344 (
		_w6770_,
		_w6780_,
		_w6807_
	);
	LUT4 #(
		.INIT('h020f)
	) name6345 (
		_w6769_,
		_w6771_,
		_w6781_,
		_w6807_,
		_w6808_
	);
	LUT4 #(
		.INIT('ha060)
	) name6346 (
		\P1_IR_reg[16]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		\P1_reg1_reg[16]/NET0131 ,
		_w648_,
		_w6809_
	);
	LUT4 #(
		.INIT('h0509)
	) name6347 (
		\P1_IR_reg[16]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		\P1_reg1_reg[16]/NET0131 ,
		_w648_,
		_w6810_
	);
	LUT4 #(
		.INIT('h5a96)
	) name6348 (
		\P1_IR_reg[16]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		\P1_reg1_reg[16]/NET0131 ,
		_w648_,
		_w6811_
	);
	LUT4 #(
		.INIT('hcdfd)
	) name6349 (
		\P1_addr_reg[16]/NET0131 ,
		_w537_,
		_w540_,
		_w784_,
		_w6812_
	);
	LUT4 #(
		.INIT('hd700)
	) name6350 (
		_w6622_,
		_w6808_,
		_w6811_,
		_w6812_,
		_w6813_
	);
	LUT4 #(
		.INIT('h8000)
	) name6351 (
		\P1_addr_reg[16]/NET0131 ,
		_w1104_,
		_w1106_,
		_w3443_,
		_w6814_
	);
	LUT2 #(
		.INIT('h1)
	) name6352 (
		_w3125_,
		_w6814_,
		_w6815_
	);
	LUT4 #(
		.INIT('h45ff)
	) name6353 (
		_w6800_,
		_w6806_,
		_w6813_,
		_w6815_,
		_w6816_
	);
	LUT4 #(
		.INIT('hbf00)
	) name6354 (
		\P1_addr_reg[17]/NET0131 ,
		_w1104_,
		_w1106_,
		_w3443_,
		_w6817_
	);
	LUT2 #(
		.INIT('h1)
	) name6355 (
		_w1294_,
		_w6817_,
		_w6818_
	);
	LUT2 #(
		.INIT('h8)
	) name6356 (
		\P1_reg1_reg[17]/NET0131 ,
		_w715_,
		_w6819_
	);
	LUT2 #(
		.INIT('h1)
	) name6357 (
		\P1_reg1_reg[17]/NET0131 ,
		_w715_,
		_w6820_
	);
	LUT2 #(
		.INIT('h6)
	) name6358 (
		\P1_reg1_reg[17]/NET0131 ,
		_w715_,
		_w6821_
	);
	LUT2 #(
		.INIT('h1)
	) name6359 (
		_w6781_,
		_w6810_,
		_w6822_
	);
	LUT4 #(
		.INIT('hba00)
	) name6360 (
		_w6770_,
		_w6783_,
		_w6784_,
		_w6822_,
		_w6823_
	);
	LUT3 #(
		.INIT('h17)
	) name6361 (
		\P1_reg1_reg[16]/NET0131 ,
		_w784_,
		_w6780_,
		_w6824_
	);
	LUT4 #(
		.INIT('h2822)
	) name6362 (
		_w6622_,
		_w6821_,
		_w6823_,
		_w6824_,
		_w6825_
	);
	LUT2 #(
		.INIT('h8)
	) name6363 (
		\P1_reg2_reg[17]/NET0131 ,
		_w715_,
		_w6826_
	);
	LUT2 #(
		.INIT('h1)
	) name6364 (
		\P1_reg2_reg[17]/NET0131 ,
		_w715_,
		_w6827_
	);
	LUT2 #(
		.INIT('h6)
	) name6365 (
		\P1_reg2_reg[17]/NET0131 ,
		_w715_,
		_w6828_
	);
	LUT2 #(
		.INIT('h1)
	) name6366 (
		_w6789_,
		_w6804_,
		_w6829_
	);
	LUT3 #(
		.INIT('h17)
	) name6367 (
		\P1_reg2_reg[16]/NET0131 ,
		_w784_,
		_w6788_,
		_w6830_
	);
	LUT4 #(
		.INIT('h4f00)
	) name6368 (
		_w6792_,
		_w6793_,
		_w6829_,
		_w6830_,
		_w6831_
	);
	LUT3 #(
		.INIT('h40)
	) name6369 (
		_w537_,
		_w540_,
		_w715_,
		_w6832_
	);
	LUT3 #(
		.INIT('h0d)
	) name6370 (
		\P1_addr_reg[17]/NET0131 ,
		_w6712_,
		_w6832_,
		_w6833_
	);
	LUT4 #(
		.INIT('h7d00)
	) name6371 (
		_w1290_,
		_w6828_,
		_w6831_,
		_w6833_,
		_w6834_
	);
	LUT4 #(
		.INIT('hbabb)
	) name6372 (
		_w3504_,
		_w6818_,
		_w6825_,
		_w6834_,
		_w6835_
	);
	LUT4 #(
		.INIT('h0509)
	) name6373 (
		\P1_IR_reg[18]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		\P1_reg2_reg[18]/NET0131 ,
		_w649_,
		_w6836_
	);
	LUT4 #(
		.INIT('h5a96)
	) name6374 (
		\P1_IR_reg[18]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		\P1_reg2_reg[18]/NET0131 ,
		_w649_,
		_w6837_
	);
	LUT3 #(
		.INIT('h07)
	) name6375 (
		\P1_reg2_reg[17]/NET0131 ,
		_w715_,
		_w6803_,
		_w6838_
	);
	LUT4 #(
		.INIT('hfe00)
	) name6376 (
		_w6789_,
		_w6802_,
		_w6804_,
		_w6838_,
		_w6839_
	);
	LUT4 #(
		.INIT('ha082)
	) name6377 (
		_w1290_,
		_w6827_,
		_w6837_,
		_w6839_,
		_w6840_
	);
	LUT4 #(
		.INIT('h0509)
	) name6378 (
		\P1_IR_reg[18]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		\P1_reg1_reg[18]/NET0131 ,
		_w649_,
		_w6841_
	);
	LUT4 #(
		.INIT('h5a96)
	) name6379 (
		\P1_IR_reg[18]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		\P1_reg1_reg[18]/NET0131 ,
		_w649_,
		_w6842_
	);
	LUT3 #(
		.INIT('h07)
	) name6380 (
		\P1_reg1_reg[17]/NET0131 ,
		_w715_,
		_w6809_,
		_w6843_
	);
	LUT4 #(
		.INIT('h020f)
	) name6381 (
		_w6808_,
		_w6810_,
		_w6820_,
		_w6843_,
		_w6844_
	);
	LUT3 #(
		.INIT('h02)
	) name6382 (
		\P1_addr_reg[18]/NET0131 ,
		_w537_,
		_w540_,
		_w6845_
	);
	LUT3 #(
		.INIT('h07)
	) name6383 (
		_w736_,
		_w6642_,
		_w6845_,
		_w6846_
	);
	LUT4 #(
		.INIT('hd700)
	) name6384 (
		_w6622_,
		_w6842_,
		_w6844_,
		_w6846_,
		_w6847_
	);
	LUT4 #(
		.INIT('hbf00)
	) name6385 (
		\P1_addr_reg[18]/NET0131 ,
		_w1104_,
		_w1106_,
		_w3443_,
		_w6848_
	);
	LUT2 #(
		.INIT('h1)
	) name6386 (
		_w1294_,
		_w6848_,
		_w6849_
	);
	LUT4 #(
		.INIT('h8000)
	) name6387 (
		\P1_addr_reg[18]/NET0131 ,
		_w1104_,
		_w1106_,
		_w3443_,
		_w6850_
	);
	LUT2 #(
		.INIT('h1)
	) name6388 (
		_w3483_,
		_w6850_,
		_w6851_
	);
	LUT4 #(
		.INIT('h0bff)
	) name6389 (
		_w6840_,
		_w6847_,
		_w6849_,
		_w6851_,
		_w6852_
	);
	LUT4 #(
		.INIT('hbf00)
	) name6390 (
		\P1_addr_reg[19]/NET0131 ,
		_w1104_,
		_w1106_,
		_w3443_,
		_w6853_
	);
	LUT2 #(
		.INIT('h1)
	) name6391 (
		_w1294_,
		_w6853_,
		_w6854_
	);
	LUT2 #(
		.INIT('h1)
	) name6392 (
		_w6827_,
		_w6836_,
		_w6855_
	);
	LUT3 #(
		.INIT('h17)
	) name6393 (
		\P1_reg2_reg[18]/NET0131 ,
		_w736_,
		_w6826_,
		_w6856_
	);
	LUT4 #(
		.INIT('h9a55)
	) name6394 (
		\P1_reg2_reg[19]/NET0131 ,
		_w6831_,
		_w6855_,
		_w6856_,
		_w6857_
	);
	LUT3 #(
		.INIT('h48)
	) name6395 (
		_w652_,
		_w1290_,
		_w6857_,
		_w6858_
	);
	LUT2 #(
		.INIT('h1)
	) name6396 (
		_w6820_,
		_w6841_,
		_w6859_
	);
	LUT3 #(
		.INIT('h17)
	) name6397 (
		\P1_reg1_reg[18]/NET0131 ,
		_w736_,
		_w6819_,
		_w6860_
	);
	LUT4 #(
		.INIT('h4f00)
	) name6398 (
		_w6823_,
		_w6824_,
		_w6859_,
		_w6860_,
		_w6861_
	);
	LUT4 #(
		.INIT('h9996)
	) name6399 (
		\P1_IR_reg[19]/NET0131 ,
		\P1_reg1_reg[19]/NET0131 ,
		_w650_,
		_w651_,
		_w6862_
	);
	LUT3 #(
		.INIT('h02)
	) name6400 (
		\P1_addr_reg[19]/NET0131 ,
		_w537_,
		_w540_,
		_w6863_
	);
	LUT3 #(
		.INIT('h07)
	) name6401 (
		_w652_,
		_w6642_,
		_w6863_,
		_w6864_
	);
	LUT4 #(
		.INIT('h7d00)
	) name6402 (
		_w6622_,
		_w6861_,
		_w6862_,
		_w6864_,
		_w6865_
	);
	LUT4 #(
		.INIT('h8000)
	) name6403 (
		\P1_addr_reg[19]/NET0131 ,
		_w1104_,
		_w1106_,
		_w3443_,
		_w6866_
	);
	LUT2 #(
		.INIT('h1)
	) name6404 (
		_w3724_,
		_w6866_,
		_w6867_
	);
	LUT4 #(
		.INIT('h45ff)
	) name6405 (
		_w6854_,
		_w6858_,
		_w6865_,
		_w6867_,
		_w6868_
	);
	LUT2 #(
		.INIT('h2)
	) name6406 (
		\P1_reg3_reg[1]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w6869_
	);
	LUT4 #(
		.INIT('hbf00)
	) name6407 (
		\P1_addr_reg[1]/NET0131 ,
		_w1104_,
		_w1106_,
		_w3443_,
		_w6870_
	);
	LUT2 #(
		.INIT('h1)
	) name6408 (
		_w1294_,
		_w6870_,
		_w6871_
	);
	LUT4 #(
		.INIT('h936c)
	) name6409 (
		\P1_IR_reg[0]/NET0131 ,
		\P1_IR_reg[1]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		\P1_reg2_reg[1]/NET0131 ,
		_w6872_
	);
	LUT2 #(
		.INIT('h6)
	) name6410 (
		_w6625_,
		_w6872_,
		_w6873_
	);
	LUT3 #(
		.INIT('h80)
	) name6411 (
		_w537_,
		_w540_,
		_w6873_,
		_w6874_
	);
	LUT4 #(
		.INIT('h936c)
	) name6412 (
		\P1_IR_reg[0]/NET0131 ,
		\P1_IR_reg[1]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		\P1_reg1_reg[1]/NET0131 ,
		_w6875_
	);
	LUT2 #(
		.INIT('h6)
	) name6413 (
		_w6623_,
		_w6875_,
		_w6876_
	);
	LUT4 #(
		.INIT('hd9fb)
	) name6414 (
		_w537_,
		_w540_,
		_w859_,
		_w6876_,
		_w6877_
	);
	LUT2 #(
		.INIT('h4)
	) name6415 (
		_w6874_,
		_w6877_,
		_w6878_
	);
	LUT3 #(
		.INIT('hd0)
	) name6416 (
		\P1_addr_reg[1]/NET0131 ,
		_w6712_,
		_w6878_,
		_w6879_
	);
	LUT3 #(
		.INIT('hab)
	) name6417 (
		_w6869_,
		_w6871_,
		_w6879_,
		_w6880_
	);
	LUT4 #(
		.INIT('hbf00)
	) name6418 (
		\P1_addr_reg[3]/NET0131 ,
		_w1104_,
		_w1106_,
		_w3443_,
		_w6881_
	);
	LUT2 #(
		.INIT('h1)
	) name6419 (
		_w1294_,
		_w6881_,
		_w6882_
	);
	LUT3 #(
		.INIT('h96)
	) name6420 (
		\P1_IR_reg[3]/NET0131 ,
		\P1_reg2_reg[3]/NET0131 ,
		_w878_,
		_w6883_
	);
	LUT4 #(
		.INIT('h17e8)
	) name6421 (
		\P1_reg2_reg[2]/NET0131 ,
		_w852_,
		_w6636_,
		_w6883_,
		_w6884_
	);
	LUT3 #(
		.INIT('h80)
	) name6422 (
		_w537_,
		_w540_,
		_w6884_,
		_w6885_
	);
	LUT3 #(
		.INIT('h96)
	) name6423 (
		\P1_IR_reg[3]/NET0131 ,
		\P1_reg1_reg[3]/NET0131 ,
		_w878_,
		_w6886_
	);
	LUT4 #(
		.INIT('h17e8)
	) name6424 (
		\P1_reg1_reg[2]/NET0131 ,
		_w852_,
		_w6640_,
		_w6886_,
		_w6887_
	);
	LUT4 #(
		.INIT('hd9fb)
	) name6425 (
		_w537_,
		_w540_,
		_w879_,
		_w6887_,
		_w6888_
	);
	LUT2 #(
		.INIT('h4)
	) name6426 (
		_w6885_,
		_w6888_,
		_w6889_
	);
	LUT3 #(
		.INIT('hd0)
	) name6427 (
		\P1_addr_reg[3]/NET0131 ,
		_w6712_,
		_w6889_,
		_w6890_
	);
	LUT3 #(
		.INIT('hab)
	) name6428 (
		_w4931_,
		_w6882_,
		_w6890_,
		_w6891_
	);
	LUT4 #(
		.INIT('hbf00)
	) name6429 (
		\P1_addr_reg[5]/NET0131 ,
		_w1104_,
		_w1106_,
		_w3443_,
		_w6892_
	);
	LUT2 #(
		.INIT('h1)
	) name6430 (
		_w1294_,
		_w6892_,
		_w6893_
	);
	LUT2 #(
		.INIT('h6)
	) name6431 (
		\P1_reg1_reg[5]/NET0131 ,
		_w937_,
		_w6894_
	);
	LUT4 #(
		.INIT('h0220)
	) name6432 (
		_w537_,
		_w540_,
		_w6695_,
		_w6894_,
		_w6895_
	);
	LUT3 #(
		.INIT('h40)
	) name6433 (
		_w537_,
		_w540_,
		_w937_,
		_w6896_
	);
	LUT2 #(
		.INIT('h6)
	) name6434 (
		\P1_reg2_reg[5]/NET0131 ,
		_w937_,
		_w6897_
	);
	LUT4 #(
		.INIT('h0880)
	) name6435 (
		_w537_,
		_w540_,
		_w6676_,
		_w6897_,
		_w6898_
	);
	LUT3 #(
		.INIT('h01)
	) name6436 (
		_w6896_,
		_w6898_,
		_w6895_,
		_w6899_
	);
	LUT3 #(
		.INIT('hd0)
	) name6437 (
		\P1_addr_reg[5]/NET0131 ,
		_w6712_,
		_w6899_,
		_w6900_
	);
	LUT3 #(
		.INIT('hab)
	) name6438 (
		_w4568_,
		_w6893_,
		_w6900_,
		_w6901_
	);
	LUT3 #(
		.INIT('h96)
	) name6439 (
		\P1_IR_reg[6]/NET0131 ,
		\P1_reg1_reg[6]/NET0131 ,
		_w915_,
		_w6902_
	);
	LUT4 #(
		.INIT('h0017)
	) name6440 (
		\P1_reg1_reg[5]/NET0131 ,
		_w937_,
		_w6695_,
		_w6902_,
		_w6903_
	);
	LUT4 #(
		.INIT('he800)
	) name6441 (
		\P1_reg1_reg[5]/NET0131 ,
		_w937_,
		_w6695_,
		_w6902_,
		_w6904_
	);
	LUT3 #(
		.INIT('h02)
	) name6442 (
		_w6622_,
		_w6904_,
		_w6903_,
		_w6905_
	);
	LUT3 #(
		.INIT('h96)
	) name6443 (
		\P1_IR_reg[6]/NET0131 ,
		\P1_reg2_reg[6]/NET0131 ,
		_w915_,
		_w6906_
	);
	LUT4 #(
		.INIT('hfdcd)
	) name6444 (
		\P1_addr_reg[6]/NET0131 ,
		_w537_,
		_w540_,
		_w926_,
		_w6907_
	);
	LUT4 #(
		.INIT('hd700)
	) name6445 (
		_w1290_,
		_w6677_,
		_w6906_,
		_w6907_,
		_w6908_
	);
	LUT4 #(
		.INIT('h8088)
	) name6446 (
		\P1_state_reg[0]/NET0131 ,
		_w6634_,
		_w6905_,
		_w6908_,
		_w6909_
	);
	LUT4 #(
		.INIT('h8000)
	) name6447 (
		\P1_addr_reg[6]/NET0131 ,
		_w1104_,
		_w1106_,
		_w3443_,
		_w6910_
	);
	LUT2 #(
		.INIT('h1)
	) name6448 (
		_w5258_,
		_w6910_,
		_w6911_
	);
	LUT2 #(
		.INIT('hb)
	) name6449 (
		_w6909_,
		_w6911_,
		_w6912_
	);
	LUT4 #(
		.INIT('h9996)
	) name6450 (
		\P1_IR_reg[7]/NET0131 ,
		\P1_reg2_reg[7]/NET0131 ,
		_w915_,
		_w916_,
		_w6913_
	);
	LUT4 #(
		.INIT('ha802)
	) name6451 (
		_w1290_,
		_w6674_,
		_w6678_,
		_w6913_,
		_w6914_
	);
	LUT4 #(
		.INIT('h9996)
	) name6452 (
		\P1_IR_reg[7]/NET0131 ,
		\P1_reg1_reg[7]/NET0131 ,
		_w915_,
		_w916_,
		_w6915_
	);
	LUT4 #(
		.INIT('h02a8)
	) name6453 (
		_w6622_,
		_w6696_,
		_w6698_,
		_w6915_,
		_w6916_
	);
	LUT4 #(
		.INIT('hcdfd)
	) name6454 (
		\P1_addr_reg[7]/NET0131 ,
		_w537_,
		_w540_,
		_w917_,
		_w6917_
	);
	LUT3 #(
		.INIT('h10)
	) name6455 (
		_w6916_,
		_w6914_,
		_w6917_,
		_w6918_
	);
	LUT4 #(
		.INIT('h8000)
	) name6456 (
		\P1_addr_reg[7]/NET0131 ,
		_w1104_,
		_w1106_,
		_w3443_,
		_w6919_
	);
	LUT2 #(
		.INIT('h1)
	) name6457 (
		_w4949_,
		_w6919_,
		_w6920_
	);
	LUT3 #(
		.INIT('h2f)
	) name6458 (
		_w6668_,
		_w6918_,
		_w6920_,
		_w6921_
	);
	LUT4 #(
		.INIT('h3c96)
	) name6459 (
		\P1_IR_reg[31]/NET0131 ,
		\P1_IR_reg[8]/NET0131 ,
		\P1_reg2_reg[8]/NET0131 ,
		_w839_,
		_w6922_
	);
	LUT3 #(
		.INIT('h28)
	) name6460 (
		_w1290_,
		_w6679_,
		_w6922_,
		_w6923_
	);
	LUT4 #(
		.INIT('h3c96)
	) name6461 (
		\P1_IR_reg[31]/NET0131 ,
		\P1_IR_reg[8]/NET0131 ,
		\P1_reg1_reg[8]/NET0131 ,
		_w839_,
		_w6924_
	);
	LUT4 #(
		.INIT('hcdfd)
	) name6462 (
		\P1_addr_reg[8]/NET0131 ,
		_w537_,
		_w540_,
		_w906_,
		_w6925_
	);
	LUT4 #(
		.INIT('hd700)
	) name6463 (
		_w6622_,
		_w6700_,
		_w6924_,
		_w6925_,
		_w6926_
	);
	LUT4 #(
		.INIT('h8000)
	) name6464 (
		\P1_addr_reg[8]/NET0131 ,
		_w1104_,
		_w1106_,
		_w3443_,
		_w6927_
	);
	LUT2 #(
		.INIT('h1)
	) name6465 (
		_w3743_,
		_w6927_,
		_w6928_
	);
	LUT4 #(
		.INIT('h8aff)
	) name6466 (
		_w6668_,
		_w6923_,
		_w6926_,
		_w6928_,
		_w6929_
	);
	LUT2 #(
		.INIT('h6)
	) name6467 (
		\P1_reg2_reg[9]/NET0131 ,
		_w840_,
		_w6930_
	);
	LUT4 #(
		.INIT('he800)
	) name6468 (
		\P1_reg2_reg[8]/NET0131 ,
		_w906_,
		_w6679_,
		_w6930_,
		_w6931_
	);
	LUT4 #(
		.INIT('h0017)
	) name6469 (
		\P1_reg2_reg[8]/NET0131 ,
		_w906_,
		_w6679_,
		_w6930_,
		_w6932_
	);
	LUT3 #(
		.INIT('h02)
	) name6470 (
		_w1290_,
		_w6932_,
		_w6931_,
		_w6933_
	);
	LUT2 #(
		.INIT('h6)
	) name6471 (
		\P1_reg1_reg[9]/NET0131 ,
		_w840_,
		_w6934_
	);
	LUT4 #(
		.INIT('ha802)
	) name6472 (
		_w6622_,
		_w6691_,
		_w6701_,
		_w6934_,
		_w6935_
	);
	LUT4 #(
		.INIT('hcdfd)
	) name6473 (
		\P1_addr_reg[9]/NET0131 ,
		_w537_,
		_w540_,
		_w840_,
		_w6936_
	);
	LUT2 #(
		.INIT('h4)
	) name6474 (
		_w6935_,
		_w6936_,
		_w6937_
	);
	LUT4 #(
		.INIT('h8000)
	) name6475 (
		\P1_addr_reg[9]/NET0131 ,
		_w1104_,
		_w1106_,
		_w3443_,
		_w6938_
	);
	LUT2 #(
		.INIT('h1)
	) name6476 (
		_w4224_,
		_w6938_,
		_w6939_
	);
	LUT4 #(
		.INIT('h8aff)
	) name6477 (
		_w6668_,
		_w6933_,
		_w6937_,
		_w6939_,
		_w6940_
	);
	LUT4 #(
		.INIT('h8000)
	) name6478 (
		_w511_,
		_w519_,
		_w522_,
		_w517_,
		_w6941_
	);
	LUT4 #(
		.INIT('h8000)
	) name6479 (
		_w1478_,
		_w1483_,
		_w1485_,
		_w1481_,
		_w6942_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name6480 (
		_w1477_,
		_w1486_,
		_w2081_,
		_w6149_,
		_w6943_
	);
	LUT3 #(
		.INIT('hc4)
	) name6481 (
		\P1_state_reg[0]/NET0131 ,
		\P2_B_reg/NET0131 ,
		_w6943_,
		_w6944_
	);
	LUT4 #(
		.INIT('h2228)
	) name6482 (
		\P2_B_reg/NET0131 ,
		\P2_IR_reg[22]/NET0131 ,
		_w2031_,
		_w2032_,
		_w6945_
	);
	LUT3 #(
		.INIT('h23)
	) name6483 (
		_w1509_,
		_w2053_,
		_w5940_,
		_w6946_
	);
	LUT3 #(
		.INIT('h32)
	) name6484 (
		_w1509_,
		_w2602_,
		_w5922_,
		_w6947_
	);
	LUT3 #(
		.INIT('h40)
	) name6485 (
		_w1509_,
		_w2053_,
		_w5940_,
		_w6948_
	);
	LUT2 #(
		.INIT('h1)
	) name6486 (
		_w6947_,
		_w6948_,
		_w6949_
	);
	LUT3 #(
		.INIT('h04)
	) name6487 (
		_w1509_,
		_w2602_,
		_w5922_,
		_w6950_
	);
	LUT4 #(
		.INIT('h0071)
	) name6488 (
		_w2049_,
		_w2617_,
		_w2628_,
		_w6950_,
		_w6951_
	);
	LUT3 #(
		.INIT('h51)
	) name6489 (
		_w6946_,
		_w6949_,
		_w6951_,
		_w6952_
	);
	LUT4 #(
		.INIT('h30b0)
	) name6490 (
		_w2136_,
		_w2154_,
		_w2161_,
		_w4599_,
		_w6953_
	);
	LUT4 #(
		.INIT('h050d)
	) name6491 (
		_w2167_,
		_w2177_,
		_w2185_,
		_w6953_,
		_w6954_
	);
	LUT2 #(
		.INIT('h1)
	) name6492 (
		_w6946_,
		_w6950_,
		_w6955_
	);
	LUT3 #(
		.INIT('h10)
	) name6493 (
		_w2619_,
		_w2624_,
		_w6955_,
		_w6956_
	);
	LUT4 #(
		.INIT('h1011)
	) name6494 (
		_w6945_,
		_w6952_,
		_w6954_,
		_w6956_,
		_w6957_
	);
	LUT2 #(
		.INIT('h2)
	) name6495 (
		_w2275_,
		_w6957_,
		_w6958_
	);
	LUT4 #(
		.INIT('h00e8)
	) name6496 (
		_w1883_,
		_w1889_,
		_w2156_,
		_w2174_,
		_w6959_
	);
	LUT3 #(
		.INIT('h31)
	) name6497 (
		_w2160_,
		_w2175_,
		_w6959_,
		_w6960_
	);
	LUT3 #(
		.INIT('h07)
	) name6498 (
		_w2154_,
		_w2177_,
		_w6960_,
		_w6961_
	);
	LUT4 #(
		.INIT('h1311)
	) name6499 (
		_w2096_,
		_w2099_,
		_w2125_,
		_w2360_,
		_w6962_
	);
	LUT4 #(
		.INIT('h0705)
	) name6500 (
		_w2128_,
		_w2129_,
		_w2141_,
		_w2371_,
		_w6963_
	);
	LUT3 #(
		.INIT('ha8)
	) name6501 (
		_w2144_,
		_w6962_,
		_w6963_,
		_w6964_
	);
	LUT4 #(
		.INIT('h004c)
	) name6502 (
		_w2124_,
		_w2451_,
		_w2448_,
		_w6964_,
		_w6965_
	);
	LUT4 #(
		.INIT('h1113)
	) name6503 (
		_w2167_,
		_w2185_,
		_w6961_,
		_w6965_,
		_w6966_
	);
	LUT4 #(
		.INIT('h0777)
	) name6504 (
		_w2051_,
		_w2052_,
		_w2600_,
		_w2601_,
		_w6967_
	);
	LUT3 #(
		.INIT('h01)
	) name6505 (
		_w1509_,
		_w5922_,
		_w6967_,
		_w6968_
	);
	LUT2 #(
		.INIT('h1)
	) name6506 (
		_w6946_,
		_w6968_,
		_w6969_
	);
	LUT3 #(
		.INIT('h10)
	) name6507 (
		_w2619_,
		_w2624_,
		_w6969_,
		_w6970_
	);
	LUT4 #(
		.INIT('h7100)
	) name6508 (
		_w2049_,
		_w2617_,
		_w2628_,
		_w6969_,
		_w6971_
	);
	LUT4 #(
		.INIT('h3031)
	) name6509 (
		_w1509_,
		_w2053_,
		_w2602_,
		_w5922_,
		_w6972_
	);
	LUT2 #(
		.INIT('h2)
	) name6510 (
		_w5941_,
		_w6972_,
		_w6973_
	);
	LUT2 #(
		.INIT('h1)
	) name6511 (
		_w6971_,
		_w6973_,
		_w6974_
	);
	LUT4 #(
		.INIT('h65aa)
	) name6512 (
		_w1811_,
		_w6966_,
		_w6970_,
		_w6974_,
		_w6975_
	);
	LUT3 #(
		.INIT('h80)
	) name6513 (
		_w2033_,
		_w2035_,
		_w2036_,
		_w6976_
	);
	LUT3 #(
		.INIT('he0)
	) name6514 (
		\P2_B_reg/NET0131 ,
		_w6975_,
		_w6976_,
		_w6977_
	);
	LUT3 #(
		.INIT('h01)
	) name6515 (
		_w1811_,
		_w2035_,
		_w2036_,
		_w6978_
	);
	LUT4 #(
		.INIT('h4500)
	) name6516 (
		_w6952_,
		_w6954_,
		_w6956_,
		_w6978_,
		_w6979_
	);
	LUT2 #(
		.INIT('h8)
	) name6517 (
		_w2037_,
		_w6975_,
		_w6980_
	);
	LUT4 #(
		.INIT('h0203)
	) name6518 (
		_w2164_,
		_w2165_,
		_w2166_,
		_w2383_,
		_w6981_
	);
	LUT4 #(
		.INIT('he800)
	) name6519 (
		_w2049_,
		_w2617_,
		_w2624_,
		_w6949_,
		_w6982_
	);
	LUT3 #(
		.INIT('h32)
	) name6520 (
		_w6946_,
		_w6948_,
		_w6950_,
		_w6983_
	);
	LUT4 #(
		.INIT('h0032)
	) name6521 (
		_w2180_,
		_w6982_,
		_w6981_,
		_w6983_,
		_w6984_
	);
	LUT2 #(
		.INIT('h1)
	) name6522 (
		_w6952_,
		_w6984_,
		_w6985_
	);
	LUT4 #(
		.INIT('h00d4)
	) name6523 (
		_w1776_,
		_w1781_,
		_w2132_,
		_w2151_,
		_w6986_
	);
	LUT3 #(
		.INIT('h31)
	) name6524 (
		_w2135_,
		_w2150_,
		_w6986_,
		_w6987_
	);
	LUT3 #(
		.INIT('ha8)
	) name6525 (
		_w2177_,
		_w6960_,
		_w6987_,
		_w6988_
	);
	LUT4 #(
		.INIT('h020b)
	) name6526 (
		_w1569_,
		_w1573_,
		_w2115_,
		_w5813_,
		_w6989_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name6527 (
		_w2108_,
		_w2111_,
		_w2352_,
		_w6989_,
		_w6990_
	);
	LUT3 #(
		.INIT('h01)
	) name6528 (
		_w2099_,
		_w2100_,
		_w2121_,
		_w6991_
	);
	LUT4 #(
		.INIT('h8000)
	) name6529 (
		_w2097_,
		_w2139_,
		_w2142_,
		_w6991_,
		_w6992_
	);
	LUT4 #(
		.INIT('h5d00)
	) name6530 (
		_w2105_,
		_w2350_,
		_w6990_,
		_w6992_,
		_w6993_
	);
	LUT3 #(
		.INIT('h02)
	) name6531 (
		_w2152_,
		_w2174_,
		_w2175_,
		_w6994_
	);
	LUT3 #(
		.INIT('h80)
	) name6532 (
		_w2147_,
		_w2172_,
		_w6994_,
		_w6995_
	);
	LUT3 #(
		.INIT('he0)
	) name6533 (
		_w6964_,
		_w6993_,
		_w6995_,
		_w6996_
	);
	LUT3 #(
		.INIT('h10)
	) name6534 (
		_w2179_,
		_w2180_,
		_w2183_,
		_w6997_
	);
	LUT3 #(
		.INIT('h10)
	) name6535 (
		_w2618_,
		_w2628_,
		_w6949_,
		_w6998_
	);
	LUT2 #(
		.INIT('h8)
	) name6536 (
		_w6997_,
		_w6998_,
		_w6999_
	);
	LUT3 #(
		.INIT('he0)
	) name6537 (
		_w6988_,
		_w6996_,
		_w6999_,
		_w7000_
	);
	LUT4 #(
		.INIT('h4448)
	) name6538 (
		_w1811_,
		_w2191_,
		_w6985_,
		_w7000_,
		_w7001_
	);
	LUT4 #(
		.INIT('h0080)
	) name6539 (
		_w1811_,
		_w2033_,
		_w2035_,
		_w2036_,
		_w7002_
	);
	LUT4 #(
		.INIT('hab00)
	) name6540 (
		\P2_B_reg/NET0131 ,
		_w6985_,
		_w7000_,
		_w7002_,
		_w7003_
	);
	LUT3 #(
		.INIT('hd0)
	) name6541 (
		_w1811_,
		_w2036_,
		_w6945_,
		_w7004_
	);
	LUT3 #(
		.INIT('h01)
	) name6542 (
		_w4593_,
		_w6947_,
		_w6948_,
		_w7005_
	);
	LUT3 #(
		.INIT('h40)
	) name6543 (
		_w2437_,
		_w6955_,
		_w7005_,
		_w7006_
	);
	LUT2 #(
		.INIT('h4)
	) name6544 (
		_w2463_,
		_w2620_,
		_w7007_
	);
	LUT2 #(
		.INIT('h8)
	) name6545 (
		_w7006_,
		_w7007_,
		_w7008_
	);
	LUT3 #(
		.INIT('h01)
	) name6546 (
		_w2531_,
		_w2705_,
		_w3190_,
		_w7009_
	);
	LUT4 #(
		.INIT('h4000)
	) name6547 (
		_w5533_,
		_w5690_,
		_w5711_,
		_w5814_,
		_w7010_
	);
	LUT3 #(
		.INIT('h10)
	) name6548 (
		_w2749_,
		_w3511_,
		_w7010_,
		_w7011_
	);
	LUT4 #(
		.INIT('h9009)
	) name6549 (
		_w1697_,
		_w1715_,
		_w1720_,
		_w1730_,
		_w7012_
	);
	LUT4 #(
		.INIT('h0008)
	) name6550 (
		_w4959_,
		_w4984_,
		_w5002_,
		_w5263_,
		_w7013_
	);
	LUT4 #(
		.INIT('h0900)
	) name6551 (
		_w1663_,
		_w1672_,
		_w4142_,
		_w4474_,
		_w7014_
	);
	LUT4 #(
		.INIT('h8000)
	) name6552 (
		_w4573_,
		_w7013_,
		_w7014_,
		_w7012_,
		_w7015_
	);
	LUT2 #(
		.INIT('h1)
	) name6553 (
		_w2793_,
		_w3212_,
		_w7016_
	);
	LUT3 #(
		.INIT('h80)
	) name6554 (
		_w7011_,
		_w7015_,
		_w7016_,
		_w7017_
	);
	LUT4 #(
		.INIT('h9009)
	) name6555 (
		_w1735_,
		_w1746_,
		_w1833_,
		_w1838_,
		_w7018_
	);
	LUT2 #(
		.INIT('h8)
	) name6556 (
		_w4190_,
		_w7018_,
		_w7019_
	);
	LUT2 #(
		.INIT('h4)
	) name6557 (
		_w2301_,
		_w7019_,
		_w7020_
	);
	LUT4 #(
		.INIT('h4000)
	) name6558 (
		_w2027_,
		_w7017_,
		_w7020_,
		_w7009_,
		_w7021_
	);
	LUT4 #(
		.INIT('h4888)
	) name6559 (
		_w1811_,
		_w2036_,
		_w7008_,
		_w7021_,
		_w7022_
	);
	LUT3 #(
		.INIT('h54)
	) name6560 (
		_w2035_,
		_w7004_,
		_w7022_,
		_w7023_
	);
	LUT4 #(
		.INIT('hccc8)
	) name6561 (
		\P2_B_reg/NET0131 ,
		_w2081_,
		_w6985_,
		_w7000_,
		_w7024_
	);
	LUT4 #(
		.INIT('h0001)
	) name6562 (
		_w7001_,
		_w7023_,
		_w7024_,
		_w7003_,
		_w7025_
	);
	LUT4 #(
		.INIT('h0100)
	) name6563 (
		_w6979_,
		_w6977_,
		_w6980_,
		_w7025_,
		_w7026_
	);
	LUT4 #(
		.INIT('hecee)
	) name6564 (
		_w2293_,
		_w6944_,
		_w6958_,
		_w7026_,
		_w7027_
	);
	LUT4 #(
		.INIT('h70d0)
	) name6565 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg2_reg[17]/NET0131 ,
		_w1476_,
		_w7028_
	);
	LUT2 #(
		.INIT('h8)
	) name6566 (
		\P2_reg2_reg[17]/NET0131 ,
		_w1487_,
		_w7029_
	);
	LUT4 #(
		.INIT('h1dd1)
	) name6567 (
		\P2_reg2_reg[17]/NET0131 ,
		_w1497_,
		_w2705_,
		_w2706_,
		_w7030_
	);
	LUT2 #(
		.INIT('h2)
	) name6568 (
		_w2038_,
		_w7030_,
		_w7031_
	);
	LUT4 #(
		.INIT('hd11d)
	) name6569 (
		\P2_reg2_reg[17]/NET0131 ,
		_w1497_,
		_w2705_,
		_w2712_,
		_w7032_
	);
	LUT2 #(
		.INIT('h2)
	) name6570 (
		_w2193_,
		_w7032_,
		_w7033_
	);
	LUT4 #(
		.INIT('haa02)
	) name6571 (
		\P2_reg2_reg[17]/NET0131 ,
		_w1491_,
		_w1493_,
		_w1496_,
		_w7034_
	);
	LUT4 #(
		.INIT('hd11d)
	) name6572 (
		\P2_reg2_reg[17]/NET0131 ,
		_w2039_,
		_w2705_,
		_w2712_,
		_w7035_
	);
	LUT4 #(
		.INIT('h8a88)
	) name6573 (
		_w2039_,
		_w2714_,
		_w2715_,
		_w2716_,
		_w7036_
	);
	LUT4 #(
		.INIT('hf100)
	) name6574 (
		_w1509_,
		_w1771_,
		_w1775_,
		_w2085_,
		_w7037_
	);
	LUT2 #(
		.INIT('h4)
	) name6575 (
		_w1777_,
		_w2088_,
		_w7038_
	);
	LUT4 #(
		.INIT('h0057)
	) name6576 (
		\P2_reg2_reg[17]/NET0131 ,
		_w2086_,
		_w2087_,
		_w7038_,
		_w7039_
	);
	LUT2 #(
		.INIT('h4)
	) name6577 (
		_w7037_,
		_w7039_,
		_w7040_
	);
	LUT4 #(
		.INIT('h5700)
	) name6578 (
		_w2081_,
		_w7034_,
		_w7036_,
		_w7040_,
		_w7041_
	);
	LUT3 #(
		.INIT('hd0)
	) name6579 (
		_w2188_,
		_w7035_,
		_w7041_,
		_w7042_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name6580 (
		_w1489_,
		_w7033_,
		_w7031_,
		_w7042_,
		_w7043_
	);
	LUT4 #(
		.INIT('heeec)
	) name6581 (
		\P1_state_reg[0]/NET0131 ,
		_w7028_,
		_w7029_,
		_w7043_,
		_w7044_
	);
	LUT4 #(
		.INIT('h70d0)
	) name6582 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg0_reg[9]/NET0131 ,
		_w1476_,
		_w7045_
	);
	LUT2 #(
		.INIT('h8)
	) name6583 (
		\P2_reg0_reg[9]/NET0131 ,
		_w1487_,
		_w7046_
	);
	LUT4 #(
		.INIT('h3202)
	) name6584 (
		\P2_reg0_reg[9]/NET0131 ,
		_w2276_,
		_w2277_,
		_w4229_,
		_w7047_
	);
	LUT4 #(
		.INIT('h0232)
	) name6585 (
		\P2_reg0_reg[9]/NET0131 ,
		_w2192_,
		_w2277_,
		_w4231_,
		_w7048_
	);
	LUT2 #(
		.INIT('h8)
	) name6586 (
		_w2277_,
		_w4749_,
		_w7049_
	);
	LUT3 #(
		.INIT('ha2)
	) name6587 (
		\P2_reg0_reg[9]/NET0131 ,
		_w2633_,
		_w2634_,
		_w7050_
	);
	LUT2 #(
		.INIT('h1)
	) name6588 (
		_w7049_,
		_w7050_,
		_w7051_
	);
	LUT3 #(
		.INIT('h10)
	) name6589 (
		_w7047_,
		_w7048_,
		_w7051_,
		_w7052_
	);
	LUT4 #(
		.INIT('h08c8)
	) name6590 (
		\P2_reg0_reg[9]/NET0131 ,
		_w2081_,
		_w2272_,
		_w4238_,
		_w7053_
	);
	LUT4 #(
		.INIT('he020)
	) name6591 (
		\P2_reg0_reg[9]/NET0131 ,
		_w2272_,
		_w2290_,
		_w4229_,
		_w7054_
	);
	LUT2 #(
		.INIT('h1)
	) name6592 (
		_w7053_,
		_w7054_,
		_w7055_
	);
	LUT4 #(
		.INIT('h3111)
	) name6593 (
		_w1489_,
		_w7046_,
		_w7052_,
		_w7055_,
		_w7056_
	);
	LUT3 #(
		.INIT('hce)
	) name6594 (
		\P1_state_reg[0]/NET0131 ,
		_w7045_,
		_w7056_,
		_w7057_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name6595 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg2_reg[9]/NET0131 ,
		_w1489_,
		_w2086_,
		_w7058_
	);
	LUT4 #(
		.INIT('h20e0)
	) name6596 (
		\P2_reg2_reg[9]/NET0131 ,
		_w2039_,
		_w2188_,
		_w4231_,
		_w7059_
	);
	LUT4 #(
		.INIT('h20e0)
	) name6597 (
		\P2_reg2_reg[9]/NET0131 ,
		_w1497_,
		_w2193_,
		_w4231_,
		_w7060_
	);
	LUT2 #(
		.INIT('h4)
	) name6598 (
		_w1660_,
		_w2088_,
		_w7061_
	);
	LUT4 #(
		.INIT('h2e00)
	) name6599 (
		\P2_reg2_reg[9]/NET0131 ,
		_w1497_,
		_w1672_,
		_w2084_,
		_w7062_
	);
	LUT2 #(
		.INIT('h1)
	) name6600 (
		_w7061_,
		_w7062_,
		_w7063_
	);
	LUT3 #(
		.INIT('h10)
	) name6601 (
		_w7060_,
		_w7059_,
		_w7063_,
		_w7064_
	);
	LUT4 #(
		.INIT('he020)
	) name6602 (
		\P2_reg2_reg[9]/NET0131 ,
		_w1497_,
		_w2038_,
		_w4229_,
		_w7065_
	);
	LUT4 #(
		.INIT('h20e0)
	) name6603 (
		\P2_reg2_reg[9]/NET0131 ,
		_w2039_,
		_w2081_,
		_w4238_,
		_w7066_
	);
	LUT2 #(
		.INIT('h1)
	) name6604 (
		_w7065_,
		_w7066_,
		_w7067_
	);
	LUT4 #(
		.INIT('hceee)
	) name6605 (
		_w4166_,
		_w7058_,
		_w7064_,
		_w7067_,
		_w7068_
	);
	LUT2 #(
		.INIT('h4)
	) name6606 (
		_w471_,
		_w1487_,
		_w7069_
	);
	LUT4 #(
		.INIT('h5554)
	) name6607 (
		_w471_,
		_w1491_,
		_w1493_,
		_w1496_,
		_w7070_
	);
	LUT4 #(
		.INIT('h007d)
	) name6608 (
		_w2277_,
		_w4593_,
		_w4594_,
		_w7070_,
		_w7071_
	);
	LUT2 #(
		.INIT('h2)
	) name6609 (
		_w2290_,
		_w7071_,
		_w7072_
	);
	LUT4 #(
		.INIT('h0155)
	) name6610 (
		_w471_,
		_w1491_,
		_w1493_,
		_w1496_,
		_w7073_
	);
	LUT4 #(
		.INIT('h007d)
	) name6611 (
		_w2272_,
		_w4593_,
		_w4594_,
		_w7073_,
		_w7074_
	);
	LUT2 #(
		.INIT('h1)
	) name6612 (
		_w2276_,
		_w7074_,
		_w7075_
	);
	LUT4 #(
		.INIT('h00d7)
	) name6613 (
		_w2272_,
		_w4593_,
		_w4599_,
		_w7073_,
		_w7076_
	);
	LUT4 #(
		.INIT('hcc40)
	) name6614 (
		_w1781_,
		_w2277_,
		_w4524_,
		_w4602_,
		_w7077_
	);
	LUT3 #(
		.INIT('h54)
	) name6615 (
		_w471_,
		_w2086_,
		_w2280_,
		_w7078_
	);
	LUT3 #(
		.INIT('h0b)
	) name6616 (
		_w1795_,
		_w2283_,
		_w7078_,
		_w7079_
	);
	LUT4 #(
		.INIT('h5700)
	) name6617 (
		_w2081_,
		_w7070_,
		_w7077_,
		_w7079_,
		_w7080_
	);
	LUT3 #(
		.INIT('he0)
	) name6618 (
		_w2192_,
		_w7076_,
		_w7080_,
		_w7081_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name6619 (
		_w1489_,
		_w7075_,
		_w7072_,
		_w7081_,
		_w7082_
	);
	LUT4 #(
		.INIT('hf200)
	) name6620 (
		\P2_reg3_reg[16]/NET0131 ,
		_w468_,
		_w470_,
		_w2293_,
		_w7083_
	);
	LUT2 #(
		.INIT('h1)
	) name6621 (
		_w6385_,
		_w7083_,
		_w7084_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name6622 (
		\P1_state_reg[0]/NET0131 ,
		_w7069_,
		_w7082_,
		_w7084_,
		_w7085_
	);
	LUT3 #(
		.INIT('h8a)
	) name6623 (
		\P1_reg2_reg[25]/NET0131 ,
		_w1141_,
		_w3443_,
		_w7086_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name6624 (
		\P1_reg2_reg[25]/NET0131 ,
		_w528_,
		_w530_,
		_w533_,
		_w7087_
	);
	LUT4 #(
		.INIT('hd11d)
	) name6625 (
		\P1_reg2_reg[25]/NET0131 ,
		_w534_,
		_w1420_,
		_w3017_,
		_w7088_
	);
	LUT4 #(
		.INIT('h2822)
	) name6626 (
		_w534_,
		_w969_,
		_w1055_,
		_w1128_,
		_w7089_
	);
	LUT2 #(
		.INIT('h8)
	) name6627 (
		_w972_,
		_w1143_,
		_w7090_
	);
	LUT4 #(
		.INIT('hddd1)
	) name6628 (
		\P1_reg2_reg[25]/NET0131 ,
		_w534_,
		_w541_,
		_w968_,
		_w7091_
	);
	LUT3 #(
		.INIT('h31)
	) name6629 (
		_w1138_,
		_w7090_,
		_w7091_,
		_w7092_
	);
	LUT4 #(
		.INIT('h5700)
	) name6630 (
		_w1136_,
		_w7087_,
		_w7089_,
		_w7092_,
		_w7093_
	);
	LUT3 #(
		.INIT('hd0)
	) name6631 (
		_w1286_,
		_w7088_,
		_w7093_,
		_w7094_
	);
	LUT4 #(
		.INIT('h1dd1)
	) name6632 (
		\P1_reg2_reg[25]/NET0131 ,
		_w534_,
		_w1420_,
		_w3003_,
		_w7095_
	);
	LUT4 #(
		.INIT('h2a08)
	) name6633 (
		_w534_,
		_w537_,
		_w1059_,
		_w3011_,
		_w7096_
	);
	LUT3 #(
		.INIT('ha8)
	) name6634 (
		_w1183_,
		_w7087_,
		_w7096_,
		_w7097_
	);
	LUT3 #(
		.INIT('h0d)
	) name6635 (
		_w1114_,
		_w7095_,
		_w7097_,
		_w7098_
	);
	LUT4 #(
		.INIT('hceee)
	) name6636 (
		_w3443_,
		_w7086_,
		_w7094_,
		_w7098_,
		_w7099_
	);
	LUT2 #(
		.INIT('h2)
	) name6637 (
		_w972_,
		_w2197_,
		_w7100_
	);
	LUT4 #(
		.INIT('h00b7)
	) name6638 (
		_w1420_,
		_w2197_,
		_w3017_,
		_w7100_,
		_w7101_
	);
	LUT2 #(
		.INIT('h2)
	) name6639 (
		_w972_,
		_w2860_,
		_w7102_
	);
	LUT3 #(
		.INIT('h10)
	) name6640 (
		_w541_,
		_w968_,
		_w2261_,
		_w7103_
	);
	LUT2 #(
		.INIT('h1)
	) name6641 (
		_w7102_,
		_w7103_,
		_w7104_
	);
	LUT3 #(
		.INIT('h70)
	) name6642 (
		_w2197_,
		_w3008_,
		_w7104_,
		_w7105_
	);
	LUT3 #(
		.INIT('hd0)
	) name6643 (
		_w1286_,
		_w7101_,
		_w7105_,
		_w7106_
	);
	LUT4 #(
		.INIT('h007b)
	) name6644 (
		_w1420_,
		_w2197_,
		_w3003_,
		_w7100_,
		_w7107_
	);
	LUT4 #(
		.INIT('h7020)
	) name6645 (
		_w537_,
		_w1059_,
		_w2197_,
		_w3011_,
		_w7108_
	);
	LUT3 #(
		.INIT('ha8)
	) name6646 (
		_w1183_,
		_w7100_,
		_w7108_,
		_w7109_
	);
	LUT3 #(
		.INIT('h0d)
	) name6647 (
		_w1114_,
		_w7107_,
		_w7109_,
		_w7110_
	);
	LUT2 #(
		.INIT('h2)
	) name6648 (
		\P1_reg3_reg[25]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w7111_
	);
	LUT2 #(
		.INIT('h2)
	) name6649 (
		\P1_state_reg[0]/NET0131 ,
		_w526_,
		_w7112_
	);
	LUT3 #(
		.INIT('h13)
	) name6650 (
		_w972_,
		_w7111_,
		_w7112_,
		_w7113_
	);
	LUT4 #(
		.INIT('h2aff)
	) name6651 (
		_w3443_,
		_w7106_,
		_w7110_,
		_w7113_,
		_w7114_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name6652 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg2_reg[3]/NET0131 ,
		_w1489_,
		_w2086_,
		_w7115_
	);
	LUT4 #(
		.INIT('haa02)
	) name6653 (
		\P2_reg2_reg[3]/NET0131 ,
		_w1491_,
		_w1493_,
		_w1496_,
		_w7116_
	);
	LUT4 #(
		.INIT('h20e0)
	) name6654 (
		\P2_reg2_reg[3]/NET0131 ,
		_w2039_,
		_w2081_,
		_w5530_,
		_w7117_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name6655 (
		\P2_reg2_reg[3]/NET0131 ,
		_w1491_,
		_w1493_,
		_w1496_,
		_w7118_
	);
	LUT4 #(
		.INIT('ha802)
	) name6656 (
		_w1497_,
		_w1565_,
		_w1582_,
		_w5533_,
		_w7119_
	);
	LUT3 #(
		.INIT('ha8)
	) name6657 (
		_w2038_,
		_w7118_,
		_w7119_,
		_w7120_
	);
	LUT3 #(
		.INIT('ha8)
	) name6658 (
		_w2193_,
		_w5633_,
		_w7118_,
		_w7121_
	);
	LUT2 #(
		.INIT('h4)
	) name6659 (
		\P2_reg3_reg[3]/NET0131 ,
		_w2088_,
		_w7122_
	);
	LUT4 #(
		.INIT('h0010)
	) name6660 (
		_w1491_,
		_w1493_,
		_w1496_,
		_w1555_,
		_w7123_
	);
	LUT4 #(
		.INIT('h1113)
	) name6661 (
		_w2084_,
		_w7122_,
		_w7118_,
		_w7123_,
		_w7124_
	);
	LUT4 #(
		.INIT('h5700)
	) name6662 (
		_w2188_,
		_w5631_,
		_w7116_,
		_w7124_,
		_w7125_
	);
	LUT4 #(
		.INIT('h0100)
	) name6663 (
		_w7121_,
		_w7117_,
		_w7120_,
		_w7125_,
		_w7126_
	);
	LUT3 #(
		.INIT('hce)
	) name6664 (
		_w4166_,
		_w7115_,
		_w7126_,
		_w7127_
	);
	LUT4 #(
		.INIT('h70d0)
	) name6665 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg0_reg[2]/NET0131 ,
		_w1476_,
		_w7128_
	);
	LUT2 #(
		.INIT('h8)
	) name6666 (
		\P2_reg0_reg[2]/NET0131 ,
		_w1487_,
		_w7129_
	);
	LUT4 #(
		.INIT('h08c8)
	) name6667 (
		\P2_reg0_reg[2]/NET0131 ,
		_w2081_,
		_w2272_,
		_w5709_,
		_w7130_
	);
	LUT4 #(
		.INIT('h20e0)
	) name6668 (
		\P2_reg0_reg[2]/NET0131 ,
		_w2272_,
		_w2290_,
		_w5718_,
		_w7131_
	);
	LUT2 #(
		.INIT('h8)
	) name6669 (
		_w2277_,
		_w5714_,
		_w7132_
	);
	LUT3 #(
		.INIT('ha2)
	) name6670 (
		\P2_reg0_reg[2]/NET0131 ,
		_w2633_,
		_w2634_,
		_w7133_
	);
	LUT2 #(
		.INIT('h1)
	) name6671 (
		_w7132_,
		_w7133_,
		_w7134_
	);
	LUT4 #(
		.INIT('h3202)
	) name6672 (
		\P2_reg0_reg[2]/NET0131 ,
		_w2192_,
		_w2277_,
		_w5712_,
		_w7135_
	);
	LUT4 #(
		.INIT('h0232)
	) name6673 (
		\P2_reg0_reg[2]/NET0131 ,
		_w2276_,
		_w2277_,
		_w5718_,
		_w7136_
	);
	LUT4 #(
		.INIT('h0100)
	) name6674 (
		_w7131_,
		_w7135_,
		_w7136_,
		_w7134_,
		_w7137_
	);
	LUT4 #(
		.INIT('h1311)
	) name6675 (
		_w1489_,
		_w7129_,
		_w7130_,
		_w7137_,
		_w7138_
	);
	LUT3 #(
		.INIT('hce)
	) name6676 (
		\P1_state_reg[0]/NET0131 ,
		_w7128_,
		_w7138_,
		_w7139_
	);
	LUT4 #(
		.INIT('h70d0)
	) name6677 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg3_reg[2]/NET0131 ,
		_w1476_,
		_w7140_
	);
	LUT2 #(
		.INIT('h8)
	) name6678 (
		\P2_reg3_reg[2]/NET0131 ,
		_w1487_,
		_w7141_
	);
	LUT4 #(
		.INIT('h08c8)
	) name6679 (
		\P2_reg3_reg[2]/NET0131 ,
		_w2081_,
		_w2277_,
		_w5709_,
		_w7142_
	);
	LUT4 #(
		.INIT('h20e0)
	) name6680 (
		\P2_reg3_reg[2]/NET0131 ,
		_w2277_,
		_w2290_,
		_w5718_,
		_w7143_
	);
	LUT3 #(
		.INIT('ha8)
	) name6681 (
		\P2_reg3_reg[2]/NET0131 ,
		_w2086_,
		_w2280_,
		_w7144_
	);
	LUT3 #(
		.INIT('h04)
	) name6682 (
		_w1564_,
		_w2083_,
		_w2282_,
		_w7145_
	);
	LUT2 #(
		.INIT('h1)
	) name6683 (
		_w7144_,
		_w7145_,
		_w7146_
	);
	LUT4 #(
		.INIT('h020e)
	) name6684 (
		\P2_reg3_reg[2]/NET0131 ,
		_w2272_,
		_w2276_,
		_w5718_,
		_w7147_
	);
	LUT4 #(
		.INIT('h3202)
	) name6685 (
		\P2_reg3_reg[2]/NET0131 ,
		_w2192_,
		_w2272_,
		_w5712_,
		_w7148_
	);
	LUT4 #(
		.INIT('h0100)
	) name6686 (
		_w7143_,
		_w7147_,
		_w7148_,
		_w7146_,
		_w7149_
	);
	LUT4 #(
		.INIT('h1311)
	) name6687 (
		_w1489_,
		_w7141_,
		_w7142_,
		_w7149_,
		_w7150_
	);
	LUT3 #(
		.INIT('hce)
	) name6688 (
		\P1_state_reg[0]/NET0131 ,
		_w7140_,
		_w7150_,
		_w7151_
	);
	LUT2 #(
		.INIT('h9)
	) name6689 (
		\P1_rd_reg/NET0131 ,
		\P2_rd_reg/NET0131 ,
		_w7152_
	);
	LUT2 #(
		.INIT('h6)
	) name6690 (
		\P1_addr_reg[0]/NET0131 ,
		\P2_addr_reg[0]/NET0131 ,
		_w7153_
	);
	LUT2 #(
		.INIT('h6)
	) name6691 (
		\P1_addr_reg[10]/NET0131 ,
		\P2_addr_reg[10]/NET0131 ,
		_w7154_
	);
	LUT2 #(
		.INIT('h1)
	) name6692 (
		\P1_addr_reg[9]/NET0131 ,
		\P2_addr_reg[9]/NET0131 ,
		_w7155_
	);
	LUT2 #(
		.INIT('h8)
	) name6693 (
		\P1_addr_reg[9]/NET0131 ,
		\P2_addr_reg[9]/NET0131 ,
		_w7156_
	);
	LUT2 #(
		.INIT('h1)
	) name6694 (
		\P1_addr_reg[6]/NET0131 ,
		\P2_addr_reg[6]/NET0131 ,
		_w7157_
	);
	LUT2 #(
		.INIT('h8)
	) name6695 (
		\P1_addr_reg[6]/NET0131 ,
		\P2_addr_reg[6]/NET0131 ,
		_w7158_
	);
	LUT2 #(
		.INIT('h1)
	) name6696 (
		\P1_addr_reg[3]/NET0131 ,
		\P2_addr_reg[3]/NET0131 ,
		_w7159_
	);
	LUT2 #(
		.INIT('h8)
	) name6697 (
		\P1_addr_reg[3]/NET0131 ,
		\P2_addr_reg[3]/NET0131 ,
		_w7160_
	);
	LUT4 #(
		.INIT('hec80)
	) name6698 (
		\P1_addr_reg[0]/NET0131 ,
		\P1_addr_reg[1]/NET0131 ,
		\P2_addr_reg[0]/NET0131 ,
		\P2_addr_reg[1]/NET0131 ,
		_w7161_
	);
	LUT4 #(
		.INIT('h0107)
	) name6699 (
		\P1_addr_reg[2]/NET0131 ,
		\P2_addr_reg[2]/NET0131 ,
		_w7160_,
		_w7161_,
		_w7162_
	);
	LUT4 #(
		.INIT('h888e)
	) name6700 (
		\P1_addr_reg[4]/NET0131 ,
		\P2_addr_reg[4]/NET0131 ,
		_w7159_,
		_w7162_,
		_w7163_
	);
	LUT4 #(
		.INIT('h0107)
	) name6701 (
		\P1_addr_reg[5]/NET0131 ,
		\P2_addr_reg[5]/NET0131 ,
		_w7158_,
		_w7163_,
		_w7164_
	);
	LUT4 #(
		.INIT('h888e)
	) name6702 (
		\P1_addr_reg[7]/NET0131 ,
		\P2_addr_reg[7]/NET0131 ,
		_w7157_,
		_w7164_,
		_w7165_
	);
	LUT4 #(
		.INIT('h0107)
	) name6703 (
		\P1_addr_reg[8]/NET0131 ,
		\P2_addr_reg[8]/NET0131 ,
		_w7156_,
		_w7165_,
		_w7166_
	);
	LUT3 #(
		.INIT('ha9)
	) name6704 (
		_w7154_,
		_w7155_,
		_w7166_,
		_w7167_
	);
	LUT2 #(
		.INIT('h6)
	) name6705 (
		\P1_addr_reg[11]/NET0131 ,
		\P2_addr_reg[11]/NET0131 ,
		_w7168_
	);
	LUT4 #(
		.INIT('h888e)
	) name6706 (
		\P1_addr_reg[10]/NET0131 ,
		\P2_addr_reg[10]/NET0131 ,
		_w7155_,
		_w7166_,
		_w7169_
	);
	LUT2 #(
		.INIT('h6)
	) name6707 (
		_w7168_,
		_w7169_,
		_w7170_
	);
	LUT2 #(
		.INIT('h8)
	) name6708 (
		\P1_addr_reg[12]/NET0131 ,
		\P2_addr_reg[12]/NET0131 ,
		_w7171_
	);
	LUT2 #(
		.INIT('h1)
	) name6709 (
		\P1_addr_reg[12]/NET0131 ,
		\P2_addr_reg[12]/NET0131 ,
		_w7172_
	);
	LUT2 #(
		.INIT('h6)
	) name6710 (
		\P1_addr_reg[12]/NET0131 ,
		\P2_addr_reg[12]/NET0131 ,
		_w7173_
	);
	LUT4 #(
		.INIT('h17e8)
	) name6711 (
		\P1_addr_reg[11]/NET0131 ,
		\P2_addr_reg[11]/NET0131 ,
		_w7169_,
		_w7173_,
		_w7174_
	);
	LUT2 #(
		.INIT('h6)
	) name6712 (
		\P1_addr_reg[13]/NET0131 ,
		\P2_addr_reg[13]/NET0131 ,
		_w7175_
	);
	LUT4 #(
		.INIT('h0017)
	) name6713 (
		\P1_addr_reg[11]/NET0131 ,
		\P2_addr_reg[11]/NET0131 ,
		_w7169_,
		_w7171_,
		_w7176_
	);
	LUT3 #(
		.INIT('hc9)
	) name6714 (
		_w7172_,
		_w7175_,
		_w7176_,
		_w7177_
	);
	LUT2 #(
		.INIT('h6)
	) name6715 (
		\P1_addr_reg[14]/NET0131 ,
		\P2_addr_reg[14]/NET0131 ,
		_w7178_
	);
	LUT4 #(
		.INIT('h888e)
	) name6716 (
		\P1_addr_reg[13]/NET0131 ,
		\P2_addr_reg[13]/NET0131 ,
		_w7172_,
		_w7176_,
		_w7179_
	);
	LUT2 #(
		.INIT('h6)
	) name6717 (
		_w7178_,
		_w7179_,
		_w7180_
	);
	LUT2 #(
		.INIT('h8)
	) name6718 (
		\P1_addr_reg[15]/NET0131 ,
		\P2_addr_reg[15]/NET0131 ,
		_w7181_
	);
	LUT2 #(
		.INIT('h1)
	) name6719 (
		\P1_addr_reg[15]/NET0131 ,
		\P2_addr_reg[15]/NET0131 ,
		_w7182_
	);
	LUT2 #(
		.INIT('h6)
	) name6720 (
		\P1_addr_reg[15]/NET0131 ,
		\P2_addr_reg[15]/NET0131 ,
		_w7183_
	);
	LUT4 #(
		.INIT('h17e8)
	) name6721 (
		\P1_addr_reg[14]/NET0131 ,
		\P2_addr_reg[14]/NET0131 ,
		_w7179_,
		_w7183_,
		_w7184_
	);
	LUT2 #(
		.INIT('h6)
	) name6722 (
		\P1_addr_reg[16]/NET0131 ,
		\P2_addr_reg[16]/NET0131 ,
		_w7185_
	);
	LUT4 #(
		.INIT('h0017)
	) name6723 (
		\P1_addr_reg[14]/NET0131 ,
		\P2_addr_reg[14]/NET0131 ,
		_w7179_,
		_w7181_,
		_w7186_
	);
	LUT3 #(
		.INIT('hc9)
	) name6724 (
		_w7182_,
		_w7185_,
		_w7186_,
		_w7187_
	);
	LUT2 #(
		.INIT('h6)
	) name6725 (
		\P1_addr_reg[17]/NET0131 ,
		\P2_addr_reg[17]/NET0131 ,
		_w7188_
	);
	LUT4 #(
		.INIT('h888e)
	) name6726 (
		\P1_addr_reg[16]/NET0131 ,
		\P2_addr_reg[16]/NET0131 ,
		_w7182_,
		_w7186_,
		_w7189_
	);
	LUT2 #(
		.INIT('h6)
	) name6727 (
		_w7188_,
		_w7189_,
		_w7190_
	);
	LUT2 #(
		.INIT('h8)
	) name6728 (
		\P1_addr_reg[18]/NET0131 ,
		\P2_addr_reg[18]/NET0131 ,
		_w7191_
	);
	LUT2 #(
		.INIT('h1)
	) name6729 (
		\P1_addr_reg[18]/NET0131 ,
		\P2_addr_reg[18]/NET0131 ,
		_w7192_
	);
	LUT2 #(
		.INIT('h6)
	) name6730 (
		\P1_addr_reg[18]/NET0131 ,
		\P2_addr_reg[18]/NET0131 ,
		_w7193_
	);
	LUT4 #(
		.INIT('h17e8)
	) name6731 (
		\P1_addr_reg[17]/NET0131 ,
		\P2_addr_reg[17]/NET0131 ,
		_w7189_,
		_w7193_,
		_w7194_
	);
	LUT2 #(
		.INIT('h6)
	) name6732 (
		\P1_addr_reg[19]/NET0131 ,
		\P2_addr_reg[19]/NET0131 ,
		_w7195_
	);
	LUT4 #(
		.INIT('h0017)
	) name6733 (
		\P1_addr_reg[17]/NET0131 ,
		\P2_addr_reg[17]/NET0131 ,
		_w7189_,
		_w7191_,
		_w7196_
	);
	LUT3 #(
		.INIT('hc9)
	) name6734 (
		_w7192_,
		_w7195_,
		_w7196_,
		_w7197_
	);
	LUT4 #(
		.INIT('h936c)
	) name6735 (
		\P1_addr_reg[0]/NET0131 ,
		\P1_addr_reg[1]/NET0131 ,
		\P2_addr_reg[0]/NET0131 ,
		\P2_addr_reg[1]/NET0131 ,
		_w7198_
	);
	LUT2 #(
		.INIT('h6)
	) name6736 (
		\P1_addr_reg[2]/NET0131 ,
		\P2_addr_reg[2]/NET0131 ,
		_w7199_
	);
	LUT2 #(
		.INIT('h6)
	) name6737 (
		_w7161_,
		_w7199_,
		_w7200_
	);
	LUT2 #(
		.INIT('h6)
	) name6738 (
		\P1_addr_reg[3]/NET0131 ,
		\P2_addr_reg[3]/NET0131 ,
		_w7201_
	);
	LUT4 #(
		.INIT('h17e8)
	) name6739 (
		\P1_addr_reg[2]/NET0131 ,
		\P2_addr_reg[2]/NET0131 ,
		_w7161_,
		_w7201_,
		_w7202_
	);
	LUT2 #(
		.INIT('h6)
	) name6740 (
		\P1_addr_reg[4]/NET0131 ,
		\P2_addr_reg[4]/NET0131 ,
		_w7203_
	);
	LUT3 #(
		.INIT('he1)
	) name6741 (
		_w7159_,
		_w7162_,
		_w7203_,
		_w7204_
	);
	LUT2 #(
		.INIT('h6)
	) name6742 (
		\P1_addr_reg[5]/NET0131 ,
		\P2_addr_reg[5]/NET0131 ,
		_w7205_
	);
	LUT2 #(
		.INIT('h6)
	) name6743 (
		_w7163_,
		_w7205_,
		_w7206_
	);
	LUT2 #(
		.INIT('h6)
	) name6744 (
		\P1_addr_reg[6]/NET0131 ,
		\P2_addr_reg[6]/NET0131 ,
		_w7207_
	);
	LUT4 #(
		.INIT('h17e8)
	) name6745 (
		\P1_addr_reg[5]/NET0131 ,
		\P2_addr_reg[5]/NET0131 ,
		_w7163_,
		_w7207_,
		_w7208_
	);
	LUT2 #(
		.INIT('h6)
	) name6746 (
		\P1_addr_reg[7]/NET0131 ,
		\P2_addr_reg[7]/NET0131 ,
		_w7209_
	);
	LUT3 #(
		.INIT('he1)
	) name6747 (
		_w7157_,
		_w7164_,
		_w7209_,
		_w7210_
	);
	LUT2 #(
		.INIT('h6)
	) name6748 (
		\P1_addr_reg[8]/NET0131 ,
		\P2_addr_reg[8]/NET0131 ,
		_w7211_
	);
	LUT2 #(
		.INIT('h6)
	) name6749 (
		_w7165_,
		_w7211_,
		_w7212_
	);
	LUT2 #(
		.INIT('h6)
	) name6750 (
		\P1_addr_reg[9]/NET0131 ,
		\P2_addr_reg[9]/NET0131 ,
		_w7213_
	);
	LUT4 #(
		.INIT('h17e8)
	) name6751 (
		\P1_addr_reg[8]/NET0131 ,
		\P2_addr_reg[8]/NET0131 ,
		_w7165_,
		_w7213_,
		_w7214_
	);
	LUT2 #(
		.INIT('h9)
	) name6752 (
		\P1_wr_reg/NET0131 ,
		\P2_wr_reg/NET0131 ,
		_w7215_
	);
	assign \P1_state_reg[0]/NET0131_syn_2  = _w216_ ;
	assign \_al_n0  = 1'b0;
	assign \_al_n1  = 1'b1;
	assign \g21_dup/_0_  = _w499_ ;
	assign \g71037/_0_  = _w1289_ ;
	assign \g71048/_0_  = _w1475_ ;
	assign \g71049/_0_  = _w2196_ ;
	assign \g71050/_0_  = _w2270_ ;
	assign \g71052/_0_  = _w2297_ ;
	assign \g71053/_0_  = _w2401_ ;
	assign \g71054/_0_  = _w2418_ ;
	assign \g71055/_0_  = _w2435_ ;
	assign \g71080/_0_  = _w2460_ ;
	assign \g71081/_0_  = _w2514_ ;
	assign \g71082/_0_  = _w2527_ ;
	assign \g71084/_0_  = _w2581_ ;
	assign \g71085/_0_  = _w2596_ ;
	assign \g71086/_0_  = _w2654_ ;
	assign \g71087/_0_  = _w2670_ ;
	assign \g71088/_0_  = _w2685_ ;
	assign \g71089/_0_  = _w2702_ ;
	assign \g71121/_0_  = _w2725_ ;
	assign \g71122/_0_  = _w2746_ ;
	assign \g71123/_0_  = _w2765_ ;
	assign \g71130/_0_  = _w2790_ ;
	assign \g71131/_0_  = _w2821_ ;
	assign \g71132/_0_  = _w2837_ ;
	assign \g71135/_0_  = _w2893_ ;
	assign \g71136/_0_  = _w2910_ ;
	assign \g71137/_0_  = _w2926_ ;
	assign \g71138/_0_  = _w2942_ ;
	assign \g71139/_0_  = _w2955_ ;
	assign \g71141/_0_  = _w2970_ ;
	assign \g71142/_0_  = _w2984_ ;
	assign \g71143/_0_  = _w2996_ ;
	assign \g71144/_0_  = _w3021_ ;
	assign \g71145/_0_  = _w3035_ ;
	assign \g71146/_0_  = _w3091_ ;
	assign \g71147/_0_  = _w3103_ ;
	assign \g71179/_0_  = _w3127_ ;
	assign \g71186/_0_  = _w3150_ ;
	assign \g71194/_0_  = _w3169_ ;
	assign \g71195/_0_  = _w3186_ ;
	assign \g71196/_0_  = _w3208_ ;
	assign \g71197/_0_  = _w3230_ ;
	assign \g71200/_0_  = _w3245_ ;
	assign \g71201/_0_  = _w3263_ ;
	assign \g71202/_0_  = _w3279_ ;
	assign \g71203/_0_  = _w3295_ ;
	assign \g71204/_0_  = _w3310_ ;
	assign \g71205/_0_  = _w3322_ ;
	assign \g71206/_0_  = _w3336_ ;
	assign \g71207/_0_  = _w3356_ ;
	assign \g71208/_0_  = _w3365_ ;
	assign \g71209/_0_  = _w3382_ ;
	assign \g71210/_0_  = _w3394_ ;
	assign \g71211/_0_  = _w3409_ ;
	assign \g71212/_0_  = _w3423_ ;
	assign \g71213/_0_  = _w3430_ ;
	assign \g71214/_0_  = _w3442_ ;
	assign \g71215/_0_  = _w3452_ ;
	assign \g71262/_0_  = _w3466_ ;
	assign \g71263/_0_  = _w3485_ ;
	assign \g71264/_0_  = _w3507_ ;
	assign \g71291/_0_  = _w3537_ ;
	assign \g71294/_0_  = _w3558_ ;
	assign \g71295/_0_  = _w3574_ ;
	assign \g71296/_0_  = _w3588_ ;
	assign \g71297/_0_  = _w3601_ ;
	assign \g71298/_0_  = _w3610_ ;
	assign \g71299/_0_  = _w3625_ ;
	assign \g71300/_0_  = _w3637_ ;
	assign \g71302/_0_  = _w3650_ ;
	assign \g71303/_0_  = _w3661_ ;
	assign \g71304/_0_  = _w3669_ ;
	assign \g71305/_0_  = _w3681_ ;
	assign \g71306/_0_  = _w3691_ ;
	assign \g71307/_0_  = _w3696_ ;
	assign \g71308/_0_  = _w3707_ ;
	assign \g71354/_0_  = _w3726_ ;
	assign \g71359/_0_  = _w3745_ ;
	assign \g71400/_0_  = _w3772_ ;
	assign \g71401/_0_  = _w3795_ ;
	assign \g71402/_0_  = _w3814_ ;
	assign \g71403/_0_  = _w3830_ ;
	assign \g71404/_0_  = _w3845_ ;
	assign \g71405/_0_  = _w3859_ ;
	assign \g71406/_0_  = _w3876_ ;
	assign \g71407/_0_  = _w3892_ ;
	assign \g71408/_0_  = _w3908_ ;
	assign \g71409/_0_  = _w3924_ ;
	assign \g71410/_0_  = _w3937_ ;
	assign \g71411/_0_  = _w3942_ ;
	assign \g71412/_0_  = _w3959_ ;
	assign \g71413/_0_  = _w3970_ ;
	assign \g71414/_0_  = _w3986_ ;
	assign \g71415/_0_  = _w4002_ ;
	assign \g71416/_0_  = _w4018_ ;
	assign \g71417/_0_  = _w4034_ ;
	assign \g71418/_0_  = _w4050_ ;
	assign \g71420/_0_  = _w4053_ ;
	assign \g71421/_0_  = _w4060_ ;
	assign \g71422/_0_  = _w4072_ ;
	assign \g71423/_0_  = _w4077_ ;
	assign \g71424/_0_  = _w4081_ ;
	assign \g71484/_0_  = _w4100_ ;
	assign \g71485/_0_  = _w4120_ ;
	assign \g71486/_0_  = _w4139_ ;
	assign \g71488/_0_  = _w4165_ ;
	assign \g71489/_0_  = _w4187_ ;
	assign \g71490/_0_  = _w4209_ ;
	assign \g71492/_0_  = _w4226_ ;
	assign \g71493/_0_  = _w4246_ ;
	assign \g71537/_0_  = _w4252_ ;
	assign \g71538/_0_  = _w4258_ ;
	assign \g71539/_0_  = _w4272_ ;
	assign \g71540/_0_  = _w4280_ ;
	assign \g71541/_0_  = _w4292_ ;
	assign \g71542/_0_  = _w4306_ ;
	assign \g71543/_0_  = _w4312_ ;
	assign \g71544/_0_  = _w4325_ ;
	assign \g71545/_0_  = _w4340_ ;
	assign \g71546/_0_  = _w4354_ ;
	assign \g71547/_0_  = _w4360_ ;
	assign \g71548/_0_  = _w4370_ ;
	assign \g71549/_0_  = _w4374_ ;
	assign \g71550/_0_  = _w4379_ ;
	assign \g71551/_0_  = _w4392_ ;
	assign \g71552/_0_  = _w4407_ ;
	assign \g71553/_0_  = _w4413_ ;
	assign \g71554/_0_  = _w4426_ ;
	assign \g71555/_0_  = _w4436_ ;
	assign \g71608/_0_  = _w4453_ ;
	assign \g71609/_0_  = _w4471_ ;
	assign \g71613/_0_  = _w4493_ ;
	assign \g71615/_0_  = _w4513_ ;
	assign \g71617/_0_  = _w4535_ ;
	assign \g71619/_0_  = _w4552_ ;
	assign \g71620/_0_  = _w4570_ ;
	assign \g71621/_0_  = _w4589_ ;
	assign \g71690/_0_  = _w4610_ ;
	assign \g71691/_0_  = _w4627_ ;
	assign \g71692/_0_  = _w4637_ ;
	assign \g71693/_0_  = _w4652_ ;
	assign \g71694/_0_  = _w4668_ ;
	assign \g71696/_0_  = _w4687_ ;
	assign \g71697/_0_  = _w4702_ ;
	assign \g71698/_0_  = _w4720_ ;
	assign \g71699/_0_  = _w4736_ ;
	assign \g71700/_0_  = _w4744_ ;
	assign \g71701/_0_  = _w4758_ ;
	assign \g71702/_0_  = _w4775_ ;
	assign \g71703/_0_  = _w4791_ ;
	assign \g71704/_0_  = _w4808_ ;
	assign \g71705/_0_  = _w4825_ ;
	assign \g71707/_0_  = _w4834_ ;
	assign \g71708/_0_  = _w4849_ ;
	assign \g71709/_0_  = _w4855_ ;
	assign \g71710/_0_  = _w4872_ ;
	assign \g71711/_0_  = _w4887_ ;
	assign \g71712/_0_  = _w4903_ ;
	assign \g71713/_0_  = _w4917_ ;
	assign \g71788/_0_  = _w4933_ ;
	assign \g71789/_0_  = _w4951_ ;
	assign \g71792/_0_  = _w4976_ ;
	assign \g71793/_0_  = _w4999_ ;
	assign \g71794/_0_  = _w5021_ ;
	assign \g71859/_0_  = _w5029_ ;
	assign \g71860/_0_  = _w5038_ ;
	assign \g71861/_0_  = _w5055_ ;
	assign \g71862/_0_  = _w5070_ ;
	assign \g71863/_0_  = _w5085_ ;
	assign \g71864/_0_  = _w5101_ ;
	assign \g71865/_0_  = _w5106_ ;
	assign \g71866/_0_  = _w5123_ ;
	assign \g71867/_0_  = _w5138_ ;
	assign \g71868/_0_  = _w5153_ ;
	assign \g71869/_0_  = _w5155_ ;
	assign \g71870/_0_  = _w5164_ ;
	assign \g71871/_0_  = _w5169_ ;
	assign \g71872/_0_  = _w5171_ ;
	assign \g71873/_0_  = _w5187_ ;
	assign \g71874/_0_  = _w5189_ ;
	assign \g71875/_0_  = _w5195_ ;
	assign \g71876/_0_  = _w5210_ ;
	assign \g71877/_0_  = _w5224_ ;
	assign \g71878/_0_  = _w5238_ ;
	assign \g71879/_0_  = _w5240_ ;
	assign \g71918/_0_  = _w5260_ ;
	assign \g71921/_0_  = _w5282_ ;
	assign \g72042/_0_  = _w5287_ ;
	assign \g72045/_0_  = _w5303_ ;
	assign \g72046/_0_  = _w5319_ ;
	assign \g72047/_0_  = _w5335_ ;
	assign \g72048/_0_  = _w5349_ ;
	assign \g72049/_0_  = _w5359_ ;
	assign \g72050/_0_  = _w5363_ ;
	assign \g72051/_0_  = _w5380_ ;
	assign \g72052/_0_  = _w5385_ ;
	assign \g72053/_0_  = _w5400_ ;
	assign \g72054/_0_  = _w5417_ ;
	assign \g72055/_0_  = _w5434_ ;
	assign \g72056/_0_  = _w5447_ ;
	assign \g72059/_0_  = _w5463_ ;
	assign \g72060/_0_  = _w5479_ ;
	assign \g72061/_0_  = _w5495_ ;
	assign \g72062/_0_  = _w5509_ ;
	assign \g72063/_0_  = _w5518_ ;
	assign \g72064/_0_  = _w5521_ ;
	assign \g72065/_0_  = _w5527_ ;
	assign \g72185/_0_  = _w5546_ ;
	assign \g72302/_0_  = _w5562_ ;
	assign \g72304/_0_  = _w5578_ ;
	assign \g72468/_0_  = _w5593_ ;
	assign \g72577/_0_  = _w5609_ ;
	assign \g72578/_0_  = _w5623_ ;
	assign \g72579/_0_  = _w5640_ ;
	assign \g72580/_0_  = _w5654_ ;
	assign \g72585/_0_  = _w5669_ ;
	assign \g72742/_0_  = _w5683_ ;
	assign \g72758/_0_  = _w5701_ ;
	assign \g72947/_0_  = _w5705_ ;
	assign \g72948/_0_  = _w5723_ ;
	assign \g72952/_0_  = _w5736_ ;
	assign \g72954/_0_  = _w5739_ ;
	assign \g72955/_0_  = _w5741_ ;
	assign \g72956/_0_  = _w5744_ ;
	assign \g72957/_0_  = _w5749_ ;
	assign \g73346/_0_  = _w5764_ ;
	assign \g73349/_0_  = _w5776_ ;
	assign \g73350/_0_  = _w5791_ ;
	assign \g73357/_0_  = _w5806_ ;
	assign \g73618/_0_  = _w5823_ ;
	assign \g74419/_0_  = _w5838_ ;
	assign \g74422/_0_  = _w5852_ ;
	assign \g74426/_0_  = _w5866_ ;
	assign \g74671/_0_  = _w5878_ ;
	assign \g75421/_0_  = _w5889_ ;
	assign \g75424/_0_  = _w5900_ ;
	assign \g75430/_0_  = _w5911_ ;
	assign \g76173/_0_  = _w5931_ ;
	assign \g76175/_0_  = _w5944_ ;
	assign \g76177/_0_  = _w5952_ ;
	assign \g76178/_0_  = _w5955_ ;
	assign \g76179/_0_  = _w5966_ ;
	assign \g76506/_0_  = _w5971_ ;
	assign \g80645/_3_  = _w5973_ ;
	assign \g80646/_3_  = _w5975_ ;
	assign \g80647/_3_  = _w5977_ ;
	assign \g80648/_3_  = _w5979_ ;
	assign \g80649/_0_  = _w5981_ ;
	assign \g80650/_0_  = _w5983_ ;
	assign \g80952/_0_  = _w5987_ ;
	assign \g80956/_0_  = _w5989_ ;
	assign \g80957/_0_  = _w5991_ ;
	assign \g80958/_0_  = _w5993_ ;
	assign \g80959/_0_  = _w5995_ ;
	assign \g80960/_0_  = _w5997_ ;
	assign \g80961/_0_  = _w5999_ ;
	assign \g80962/_0_  = _w6001_ ;
	assign \g80963/_0_  = _w6003_ ;
	assign \g80964/_0_  = _w6005_ ;
	assign \g80965/_0_  = _w6007_ ;
	assign \g80966/_3_  = _w6009_ ;
	assign \g80967/_0_  = _w6011_ ;
	assign \g80968/_0_  = _w6013_ ;
	assign \g80969/_0_  = _w6015_ ;
	assign \g80970/_0_  = _w6016_ ;
	assign \g80971/_0_  = _w6018_ ;
	assign \g80972/_0_  = _w6020_ ;
	assign \g80973/_0_  = _w6022_ ;
	assign \g80974/_3_  = _w6024_ ;
	assign \g80975/_0_  = _w6026_ ;
	assign \g80976/_0_  = _w6028_ ;
	assign \g80977/_0_  = _w6030_ ;
	assign \g80978/_3_  = _w6032_ ;
	assign \g80979/_0_  = _w6034_ ;
	assign \g80980/_0_  = _w6036_ ;
	assign \g80981/_0_  = _w6038_ ;
	assign \g80982/_3_  = _w6040_ ;
	assign \g81025/_3_  = _w6042_ ;
	assign \g81026/_3_  = _w6044_ ;
	assign \g81027/_3_  = _w6046_ ;
	assign \g81028/_3_  = _w6048_ ;
	assign \g81029/_3_  = _w6050_ ;
	assign \g81030/_3_  = _w6052_ ;
	assign \g81031/_3_  = _w6054_ ;
	assign \g81032/_3_  = _w6056_ ;
	assign \g81033/_3_  = _w6058_ ;
	assign \g81034/_3_  = _w6060_ ;
	assign \g81035/_3_  = _w6062_ ;
	assign \g81036/_3_  = _w6064_ ;
	assign \g81037/_3_  = _w6066_ ;
	assign \g81038/_3_  = _w6068_ ;
	assign \g81039/_3_  = _w6069_ ;
	assign \g81040/_3_  = _w6071_ ;
	assign \g81041/_3_  = _w6073_ ;
	assign \g81042/_3_  = _w6075_ ;
	assign \g81043/_0_  = _w6077_ ;
	assign \g81044/_3_  = _w6079_ ;
	assign \g81045/_0_  = _w6083_ ;
	assign \g81046/_3_  = _w6085_ ;
	assign \g81047/_3_  = _w6087_ ;
	assign \g81048/_0_  = _w6089_ ;
	assign \g81049/_3_  = _w6091_ ;
	assign \g81050/_3_  = _w6093_ ;
	assign \g81051/_3_  = _w6095_ ;
	assign \g81052/_3_  = _w6097_ ;
	assign \g81524/_0_  = _w1579_ ;
	assign \g81534/_0_  = _w868_ ;
	assign \g82411/_0_  = _w6248_ ;
	assign \g82413/_0_  = _w6263_ ;
	assign \g82414/_0_  = _w6278_ ;
	assign \g82415/_0_  = _w6311_ ;
	assign \g82416/_0_  = _w6327_ ;
	assign \g82417/_0_  = _w6349_ ;
	assign \g82418/_0_  = _w6365_ ;
	assign \g82419/_0_  = _w6384_ ;
	assign \g82420/_0_  = _w6402_ ;
	assign \g82421/_0_  = _w6428_ ;
	assign \g82422/_0_  = _w6455_ ;
	assign \g82423/_0_  = _w6474_ ;
	assign \g82424/_0_  = _w6493_ ;
	assign \g82425/_0_  = _w6512_ ;
	assign \g82426/_0_  = _w6531_ ;
	assign \g82427/_0_  = _w6551_ ;
	assign \g82428/_0_  = _w6570_ ;
	assign \g82429/_0_  = _w6585_ ;
	assign \g82430/_0_  = _w6604_ ;
	assign \g82432/_0_  = _w6621_ ;
	assign \g82435/_0_  = _w6646_ ;
	assign \g82436/_0_  = _w6664_ ;
	assign \g83031/u3_syn_4  = _w3443_ ;
	assign \g83221/_0_  = _w6665_ ;
	assign \g83364/_0_  = _w6667_ ;
	assign \g83474/_0_  = _w6708_ ;
	assign \g83478/_0_  = _w6716_ ;
	assign \g83479/_0_  = _w6728_ ;
	assign \g83480/_0_  = _w6742_ ;
	assign \g83481/_0_  = _w6759_ ;
	assign \g83482/_0_  = _w6777_ ;
	assign \g83484/_0_  = _w6798_ ;
	assign \g83486/_0_  = _w6816_ ;
	assign \g83487/_0_  = _w6835_ ;
	assign \g83488/_0_  = _w6852_ ;
	assign \g83489/_0_  = _w6868_ ;
	assign \g83490/_0_  = _w6880_ ;
	assign \g83491/_0_  = _w6891_ ;
	assign \g83492/_0_  = _w6901_ ;
	assign \g83493/_0_  = _w6912_ ;
	assign \g83494/_0_  = _w6921_ ;
	assign \g83495/_0_  = _w6929_ ;
	assign \g83496/_0_  = _w6940_ ;
	assign \g83505/_0_  = _w1494_ ;
	assign \g83622/u3_syn_4  = _w4166_ ;
	assign \g83853/_0_  = _w533_ ;
	assign \g83905/_0_  = _w1496_ ;
	assign \g84145/u3_syn_4  = _w6941_ ;
	assign \g84148/u3_syn_4  = _w6942_ ;
	assign \g85427/_2_  = _w1976_ ;
	assign \g85433/_0_  = _w644_ ;
	assign \g85458/_0_  = _w1152_ ;
	assign \g85512/_0_  = _w1180_ ;
	assign \g85517/_0_  = _w2050_ ;
	assign \g85963/_0_  = _w1664_ ;
	assign \g85996/_0_  = _w978_ ;
	assign \g86064/_0_  = _w723_ ;
	assign \g86079/_0_  = _w707_ ;
	assign \g86088/_0_  = _w1560_ ;
	assign \g86096/_0_  = _w1079_ ;
	assign \g86107/_0_  = _w925_ ;
	assign \g86159/_0_  = _w1024_ ;
	assign \g86232_dup/_0_  = _w753_ ;
	assign \g86249/_0_  = _w792_ ;
	assign \g86258/_0_  = _w1961_ ;
	assign \g86268/_0_  = _w1944_ ;
	assign \g86278/_0_  = _w800_ ;
	assign \g86281/_0_  = _w1071_ ;
	assign \g86293/_0_  = _w2024_ ;
	assign \g86305/_0_  = _w820_ ;
	assign \g86313/_0_  = _w1922_ ;
	assign \g86329/_0_  = _w1721_ ;
	assign \g86338/_0_  = _w1698_ ;
	assign \g86355/_0_  = _w1752_ ;
	assign \g86362/_0_  = _w904_ ;
	assign \g86375/_0_  = _w1647_ ;
	assign \g86385/_0_  = _w1677_ ;
	assign \g86394/_0_  = _w1533_ ;
	assign \g86405/_0_  = _w1503_ ;
	assign \g86413/_0_  = _w1587_ ;
	assign \g86425/_0_  = _w834_ ;
	assign \g86433_dup/_0_  = _w1600_ ;
	assign \g86441/_0_  = _w1551_ ;
	assign \g86448/_0_  = _w1989_ ;
	assign \g86484/_0_  = _w1839_ ;
	assign \g86493/_0_  = _w1820_ ;
	assign \g86501/_0_  = _w913_ ;
	assign \g86509/_0_  = _w746_ ;
	assign \g86518/_0_  = _w888_ ;
	assign \g86527/_0_  = _w877_ ;
	assign \g86531/_0_  = _w850_ ;
	assign \g86541/_0_  = _w867_ ;
	assign \g86549/_0_  = _w858_ ;
	assign \g86577/_0_  = _w1005_ ;
	assign \g86598/_0_  = _w1570_ ;
	assign \g86607/_0_  = _w1060_ ;
	assign \g87968/_0_  = _w1478_ ;
	assign \g93740/_0_  = _w1782_ ;
	assign \g93779/_0_  = _w2603_ ;
	assign \g93782/_0_  = _w2054_ ;
	assign \g93859/_0_  = _w1908_ ;
	assign \g93950/_0_  = _w7027_ ;
	assign \g93972/_0_  = _w7044_ ;
	assign \g94026/_0_  = _w1873_ ;
	assign \g94078/_0_  = _w680_ ;
	assign \g94095/_0_  = _w1890_ ;
	assign \g94136/_0_  = _w1041_ ;
	assign \g94238/_0_  = _w7057_ ;
	assign \g94252/_0_  = _w935_ ;
	assign \g94278/_0_  = _w7068_ ;
	assign \g94380/_0_  = _w7085_ ;
	assign \g94545/_0_  = _w7099_ ;
	assign \g94586/_0_  = _w1052_ ;
	assign \g94640/_0_  = _w7114_ ;
	assign \g94710/_0_  = _w7127_ ;
	assign \g94743/_0_  = _w7139_ ;
	assign \g94877/_0_  = _w1736_ ;
	assign \g95093/_0_  = _w1578_ ;
	assign \g95139/_0_  = _w1620_ ;
	assign \g95161/_0_  = _w763_ ;
	assign \g95165/_0_  = _w773_ ;
	assign \g95204/_0_  = _w531_ ;
	assign \g95395/_0_  = _w809_ ;
	assign \g95447/_0_  = _w7151_ ;
	assign rd_pad = _w7152_ ;
	assign \so[0]_pad  = _w7153_ ;
	assign \so[10]_pad  = _w7167_ ;
	assign \so[11]_pad  = _w7170_ ;
	assign \so[12]_pad  = _w7174_ ;
	assign \so[13]_pad  = _w7177_ ;
	assign \so[14]_pad  = _w7180_ ;
	assign \so[15]_pad  = _w7184_ ;
	assign \so[16]_pad  = _w7187_ ;
	assign \so[17]_pad  = _w7190_ ;
	assign \so[18]_pad  = _w7194_ ;
	assign \so[19]_pad  = _w7197_ ;
	assign \so[1]_pad  = _w7198_ ;
	assign \so[2]_pad  = _w7200_ ;
	assign \so[3]_pad  = _w7202_ ;
	assign \so[4]_pad  = _w7204_ ;
	assign \so[5]_pad  = _w7206_ ;
	assign \so[6]_pad  = _w7208_ ;
	assign \so[7]_pad  = _w7210_ ;
	assign \so[8]_pad  = _w7212_ ;
	assign \so[9]_pad  = _w7214_ ;
	assign wr_pad = _w7215_ ;
endmodule;