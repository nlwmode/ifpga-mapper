module top( a_pad , b_pad , c_pad , d_pad , e_pad , f_pad , g_pad , h_pad , i_pad , j_pad , k_pad , l_pad , m_pad , n_pad );
  input a_pad ;
  input b_pad ;
  input c_pad ;
  input d_pad ;
  input e_pad ;
  input f_pad ;
  output g_pad ;
  output h_pad ;
  output i_pad ;
  output j_pad ;
  output k_pad ;
  output l_pad ;
  output m_pad ;
  output n_pad ;
  wire n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 ;
  assign n7 = d_pad & ~e_pad ;
  assign n8 = ~c_pad & ~f_pad ;
  assign n9 = n7 & n8 ;
  assign n10 = ~a_pad & ~b_pad ;
  assign n11 = n9 & n10 ;
  assign n12 = a_pad & ~b_pad ;
  assign n13 = n9 & n12 ;
  assign n14 = ~a_pad & b_pad ;
  assign n15 = n9 & n14 ;
  assign n16 = a_pad & b_pad ;
  assign n17 = n9 & n16 ;
  assign n18 = c_pad & ~f_pad ;
  assign n19 = n7 & n18 ;
  assign n20 = n10 & n19 ;
  assign n21 = n12 & n19 ;
  assign n22 = n14 & n19 ;
  assign n23 = n16 & n19 ;
  assign g_pad = ~n11 ;
  assign h_pad = ~n13 ;
  assign i_pad = ~n15 ;
  assign j_pad = ~n17 ;
  assign k_pad = ~n20 ;
  assign l_pad = ~n21 ;
  assign m_pad = ~n22 ;
  assign n_pad = ~n23 ;
endmodule
