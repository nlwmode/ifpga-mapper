module top (\a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] , \a[17] , \a[18] , \a[19] , \a[20] , \a[21] , \a[22] , \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[30] , \a[31] , \a[32] , \a[33] , \a[34] , \a[35] , \a[36] , \a[37] , \a[38] , \a[39] , \a[40] , \a[41] , \a[42] , \a[43] , \a[44] , \a[45] , \a[46] , \a[47] , \a[48] , \a[49] , \a[50] , \a[51] , \a[52] , \a[53] , \a[54] , \a[55] , \a[56] , \a[57] , \a[58] , \a[59] , \a[60] , \a[61] , \a[62] , \a[63] , \a[64] , \a[65] , \a[66] , \a[67] , \a[68] , \a[69] , \a[70] , \a[71] , \a[72] , \a[73] , \a[74] , \a[75] , \a[76] , \a[77] , \a[78] , \a[79] , \a[80] , \a[81] , \a[82] , \a[83] , \a[84] , \a[85] , \a[86] , \a[87] , \a[88] , \a[89] , \a[90] , \a[91] , \a[92] , \a[93] , \a[94] , \a[95] , \a[96] , \a[97] , \a[98] , \a[99] , \a[100] , \a[101] , \a[102] , \a[103] , \a[104] , \a[105] , \a[106] , \a[107] , \a[108] , \a[109] , \a[110] , \a[111] , \a[112] , \a[113] , \a[114] , \a[115] , \a[116] , \a[117] , \a[118] , \a[119] , \a[120] , \a[121] , \a[122] , \a[123] , \a[124] , \a[125] , \a[126] , \a[127] , \shift[0] , \shift[1] , \shift[2] , \shift[3] , \shift[4] , \shift[5] , \shift[6] , \result[0] , \result[1] , \result[2] , \result[3] , \result[4] , \result[5] , \result[6] , \result[7] , \result[8] , \result[9] , \result[10] , \result[11] , \result[12] , \result[13] , \result[14] , \result[15] , \result[16] , \result[17] , \result[18] , \result[19] , \result[20] , \result[21] , \result[22] , \result[23] , \result[24] , \result[25] , \result[26] , \result[27] , \result[28] , \result[29] , \result[30] , \result[31] , \result[32] , \result[33] , \result[34] , \result[35] , \result[36] , \result[37] , \result[38] , \result[39] , \result[40] , \result[41] , \result[42] , \result[43] , \result[44] , \result[45] , \result[46] , \result[47] , \result[48] , \result[49] , \result[50] , \result[51] , \result[52] , \result[53] , \result[54] , \result[55] , \result[56] , \result[57] , \result[58] , \result[59] , \result[60] , \result[61] , \result[62] , \result[63] , \result[64] , \result[65] , \result[66] , \result[67] , \result[68] , \result[69] , \result[70] , \result[71] , \result[72] , \result[73] , \result[74] , \result[75] , \result[76] , \result[77] , \result[78] , \result[79] , \result[80] , \result[81] , \result[82] , \result[83] , \result[84] , \result[85] , \result[86] , \result[87] , \result[88] , \result[89] , \result[90] , \result[91] , \result[92] , \result[93] , \result[94] , \result[95] , \result[96] , \result[97] , \result[98] , \result[99] , \result[100] , \result[101] , \result[102] , \result[103] , \result[104] , \result[105] , \result[106] , \result[107] , \result[108] , \result[109] , \result[110] , \result[111] , \result[112] , \result[113] , \result[114] , \result[115] , \result[116] , \result[117] , \result[118] , \result[119] , \result[120] , \result[121] , \result[122] , \result[123] , \result[124] , \result[125] , \result[126] , \result[127] );
	input \a[0]  ;
	input \a[1]  ;
	input \a[2]  ;
	input \a[3]  ;
	input \a[4]  ;
	input \a[5]  ;
	input \a[6]  ;
	input \a[7]  ;
	input \a[8]  ;
	input \a[9]  ;
	input \a[10]  ;
	input \a[11]  ;
	input \a[12]  ;
	input \a[13]  ;
	input \a[14]  ;
	input \a[15]  ;
	input \a[16]  ;
	input \a[17]  ;
	input \a[18]  ;
	input \a[19]  ;
	input \a[20]  ;
	input \a[21]  ;
	input \a[22]  ;
	input \a[23]  ;
	input \a[24]  ;
	input \a[25]  ;
	input \a[26]  ;
	input \a[27]  ;
	input \a[28]  ;
	input \a[29]  ;
	input \a[30]  ;
	input \a[31]  ;
	input \a[32]  ;
	input \a[33]  ;
	input \a[34]  ;
	input \a[35]  ;
	input \a[36]  ;
	input \a[37]  ;
	input \a[38]  ;
	input \a[39]  ;
	input \a[40]  ;
	input \a[41]  ;
	input \a[42]  ;
	input \a[43]  ;
	input \a[44]  ;
	input \a[45]  ;
	input \a[46]  ;
	input \a[47]  ;
	input \a[48]  ;
	input \a[49]  ;
	input \a[50]  ;
	input \a[51]  ;
	input \a[52]  ;
	input \a[53]  ;
	input \a[54]  ;
	input \a[55]  ;
	input \a[56]  ;
	input \a[57]  ;
	input \a[58]  ;
	input \a[59]  ;
	input \a[60]  ;
	input \a[61]  ;
	input \a[62]  ;
	input \a[63]  ;
	input \a[64]  ;
	input \a[65]  ;
	input \a[66]  ;
	input \a[67]  ;
	input \a[68]  ;
	input \a[69]  ;
	input \a[70]  ;
	input \a[71]  ;
	input \a[72]  ;
	input \a[73]  ;
	input \a[74]  ;
	input \a[75]  ;
	input \a[76]  ;
	input \a[77]  ;
	input \a[78]  ;
	input \a[79]  ;
	input \a[80]  ;
	input \a[81]  ;
	input \a[82]  ;
	input \a[83]  ;
	input \a[84]  ;
	input \a[85]  ;
	input \a[86]  ;
	input \a[87]  ;
	input \a[88]  ;
	input \a[89]  ;
	input \a[90]  ;
	input \a[91]  ;
	input \a[92]  ;
	input \a[93]  ;
	input \a[94]  ;
	input \a[95]  ;
	input \a[96]  ;
	input \a[97]  ;
	input \a[98]  ;
	input \a[99]  ;
	input \a[100]  ;
	input \a[101]  ;
	input \a[102]  ;
	input \a[103]  ;
	input \a[104]  ;
	input \a[105]  ;
	input \a[106]  ;
	input \a[107]  ;
	input \a[108]  ;
	input \a[109]  ;
	input \a[110]  ;
	input \a[111]  ;
	input \a[112]  ;
	input \a[113]  ;
	input \a[114]  ;
	input \a[115]  ;
	input \a[116]  ;
	input \a[117]  ;
	input \a[118]  ;
	input \a[119]  ;
	input \a[120]  ;
	input \a[121]  ;
	input \a[122]  ;
	input \a[123]  ;
	input \a[124]  ;
	input \a[125]  ;
	input \a[126]  ;
	input \a[127]  ;
	input \shift[0]  ;
	input \shift[1]  ;
	input \shift[2]  ;
	input \shift[3]  ;
	input \shift[4]  ;
	input \shift[5]  ;
	input \shift[6]  ;
	output \result[0]  ;
	output \result[1]  ;
	output \result[2]  ;
	output \result[3]  ;
	output \result[4]  ;
	output \result[5]  ;
	output \result[6]  ;
	output \result[7]  ;
	output \result[8]  ;
	output \result[9]  ;
	output \result[10]  ;
	output \result[11]  ;
	output \result[12]  ;
	output \result[13]  ;
	output \result[14]  ;
	output \result[15]  ;
	output \result[16]  ;
	output \result[17]  ;
	output \result[18]  ;
	output \result[19]  ;
	output \result[20]  ;
	output \result[21]  ;
	output \result[22]  ;
	output \result[23]  ;
	output \result[24]  ;
	output \result[25]  ;
	output \result[26]  ;
	output \result[27]  ;
	output \result[28]  ;
	output \result[29]  ;
	output \result[30]  ;
	output \result[31]  ;
	output \result[32]  ;
	output \result[33]  ;
	output \result[34]  ;
	output \result[35]  ;
	output \result[36]  ;
	output \result[37]  ;
	output \result[38]  ;
	output \result[39]  ;
	output \result[40]  ;
	output \result[41]  ;
	output \result[42]  ;
	output \result[43]  ;
	output \result[44]  ;
	output \result[45]  ;
	output \result[46]  ;
	output \result[47]  ;
	output \result[48]  ;
	output \result[49]  ;
	output \result[50]  ;
	output \result[51]  ;
	output \result[52]  ;
	output \result[53]  ;
	output \result[54]  ;
	output \result[55]  ;
	output \result[56]  ;
	output \result[57]  ;
	output \result[58]  ;
	output \result[59]  ;
	output \result[60]  ;
	output \result[61]  ;
	output \result[62]  ;
	output \result[63]  ;
	output \result[64]  ;
	output \result[65]  ;
	output \result[66]  ;
	output \result[67]  ;
	output \result[68]  ;
	output \result[69]  ;
	output \result[70]  ;
	output \result[71]  ;
	output \result[72]  ;
	output \result[73]  ;
	output \result[74]  ;
	output \result[75]  ;
	output \result[76]  ;
	output \result[77]  ;
	output \result[78]  ;
	output \result[79]  ;
	output \result[80]  ;
	output \result[81]  ;
	output \result[82]  ;
	output \result[83]  ;
	output \result[84]  ;
	output \result[85]  ;
	output \result[86]  ;
	output \result[87]  ;
	output \result[88]  ;
	output \result[89]  ;
	output \result[90]  ;
	output \result[91]  ;
	output \result[92]  ;
	output \result[93]  ;
	output \result[94]  ;
	output \result[95]  ;
	output \result[96]  ;
	output \result[97]  ;
	output \result[98]  ;
	output \result[99]  ;
	output \result[100]  ;
	output \result[101]  ;
	output \result[102]  ;
	output \result[103]  ;
	output \result[104]  ;
	output \result[105]  ;
	output \result[106]  ;
	output \result[107]  ;
	output \result[108]  ;
	output \result[109]  ;
	output \result[110]  ;
	output \result[111]  ;
	output \result[112]  ;
	output \result[113]  ;
	output \result[114]  ;
	output \result[115]  ;
	output \result[116]  ;
	output \result[117]  ;
	output \result[118]  ;
	output \result[119]  ;
	output \result[120]  ;
	output \result[121]  ;
	output \result[122]  ;
	output \result[123]  ;
	output \result[124]  ;
	output \result[125]  ;
	output \result[126]  ;
	output \result[127]  ;
	wire _w3276_ ;
	wire _w3275_ ;
	wire _w3274_ ;
	wire _w3273_ ;
	wire _w3272_ ;
	wire _w3271_ ;
	wire _w3270_ ;
	wire _w3269_ ;
	wire _w3268_ ;
	wire _w3267_ ;
	wire _w3266_ ;
	wire _w3265_ ;
	wire _w3264_ ;
	wire _w3263_ ;
	wire _w3262_ ;
	wire _w3261_ ;
	wire _w3260_ ;
	wire _w3259_ ;
	wire _w3258_ ;
	wire _w3257_ ;
	wire _w3256_ ;
	wire _w3255_ ;
	wire _w3254_ ;
	wire _w3253_ ;
	wire _w3252_ ;
	wire _w3251_ ;
	wire _w3250_ ;
	wire _w3249_ ;
	wire _w3248_ ;
	wire _w3247_ ;
	wire _w3246_ ;
	wire _w3245_ ;
	wire _w3244_ ;
	wire _w3243_ ;
	wire _w3242_ ;
	wire _w3241_ ;
	wire _w3240_ ;
	wire _w3239_ ;
	wire _w3238_ ;
	wire _w3237_ ;
	wire _w3236_ ;
	wire _w3235_ ;
	wire _w3234_ ;
	wire _w3233_ ;
	wire _w3232_ ;
	wire _w3231_ ;
	wire _w3230_ ;
	wire _w3229_ ;
	wire _w3228_ ;
	wire _w3227_ ;
	wire _w3226_ ;
	wire _w3225_ ;
	wire _w3224_ ;
	wire _w3223_ ;
	wire _w3222_ ;
	wire _w3221_ ;
	wire _w3220_ ;
	wire _w3219_ ;
	wire _w3218_ ;
	wire _w3217_ ;
	wire _w3216_ ;
	wire _w3215_ ;
	wire _w3214_ ;
	wire _w3213_ ;
	wire _w3212_ ;
	wire _w3211_ ;
	wire _w3210_ ;
	wire _w3209_ ;
	wire _w3208_ ;
	wire _w3207_ ;
	wire _w3206_ ;
	wire _w3205_ ;
	wire _w3204_ ;
	wire _w3203_ ;
	wire _w3202_ ;
	wire _w3201_ ;
	wire _w3200_ ;
	wire _w3199_ ;
	wire _w3198_ ;
	wire _w3197_ ;
	wire _w3196_ ;
	wire _w3195_ ;
	wire _w3194_ ;
	wire _w3193_ ;
	wire _w3192_ ;
	wire _w3191_ ;
	wire _w3190_ ;
	wire _w3189_ ;
	wire _w3188_ ;
	wire _w3187_ ;
	wire _w3186_ ;
	wire _w3185_ ;
	wire _w3184_ ;
	wire _w3183_ ;
	wire _w3182_ ;
	wire _w3181_ ;
	wire _w3180_ ;
	wire _w3179_ ;
	wire _w3178_ ;
	wire _w3177_ ;
	wire _w3176_ ;
	wire _w3175_ ;
	wire _w3174_ ;
	wire _w3173_ ;
	wire _w3172_ ;
	wire _w3171_ ;
	wire _w3170_ ;
	wire _w3169_ ;
	wire _w3168_ ;
	wire _w3167_ ;
	wire _w3166_ ;
	wire _w3165_ ;
	wire _w3164_ ;
	wire _w3163_ ;
	wire _w3162_ ;
	wire _w3161_ ;
	wire _w3160_ ;
	wire _w3159_ ;
	wire _w3158_ ;
	wire _w3157_ ;
	wire _w3156_ ;
	wire _w3155_ ;
	wire _w3154_ ;
	wire _w3153_ ;
	wire _w3152_ ;
	wire _w3151_ ;
	wire _w3150_ ;
	wire _w3149_ ;
	wire _w3148_ ;
	wire _w3147_ ;
	wire _w3146_ ;
	wire _w3145_ ;
	wire _w3144_ ;
	wire _w3143_ ;
	wire _w3142_ ;
	wire _w3141_ ;
	wire _w3140_ ;
	wire _w3139_ ;
	wire _w3138_ ;
	wire _w3137_ ;
	wire _w3136_ ;
	wire _w3135_ ;
	wire _w3134_ ;
	wire _w3133_ ;
	wire _w3132_ ;
	wire _w3131_ ;
	wire _w3130_ ;
	wire _w3129_ ;
	wire _w3128_ ;
	wire _w3127_ ;
	wire _w3126_ ;
	wire _w3125_ ;
	wire _w3124_ ;
	wire _w3123_ ;
	wire _w3122_ ;
	wire _w3121_ ;
	wire _w3120_ ;
	wire _w3119_ ;
	wire _w3118_ ;
	wire _w3117_ ;
	wire _w3116_ ;
	wire _w3115_ ;
	wire _w3114_ ;
	wire _w3113_ ;
	wire _w3112_ ;
	wire _w3111_ ;
	wire _w3110_ ;
	wire _w3109_ ;
	wire _w3108_ ;
	wire _w3107_ ;
	wire _w3106_ ;
	wire _w3105_ ;
	wire _w3104_ ;
	wire _w3103_ ;
	wire _w3102_ ;
	wire _w3101_ ;
	wire _w3100_ ;
	wire _w3099_ ;
	wire _w3098_ ;
	wire _w3097_ ;
	wire _w3096_ ;
	wire _w3095_ ;
	wire _w3094_ ;
	wire _w3093_ ;
	wire _w3092_ ;
	wire _w3091_ ;
	wire _w3090_ ;
	wire _w3089_ ;
	wire _w3088_ ;
	wire _w3087_ ;
	wire _w3086_ ;
	wire _w3085_ ;
	wire _w3084_ ;
	wire _w3083_ ;
	wire _w3082_ ;
	wire _w3081_ ;
	wire _w3080_ ;
	wire _w3079_ ;
	wire _w3078_ ;
	wire _w3077_ ;
	wire _w3076_ ;
	wire _w3075_ ;
	wire _w3074_ ;
	wire _w3073_ ;
	wire _w3072_ ;
	wire _w3071_ ;
	wire _w3070_ ;
	wire _w3069_ ;
	wire _w3068_ ;
	wire _w3067_ ;
	wire _w3066_ ;
	wire _w3065_ ;
	wire _w3064_ ;
	wire _w3063_ ;
	wire _w3062_ ;
	wire _w3061_ ;
	wire _w3060_ ;
	wire _w3059_ ;
	wire _w3058_ ;
	wire _w3057_ ;
	wire _w3056_ ;
	wire _w3055_ ;
	wire _w3054_ ;
	wire _w3053_ ;
	wire _w3052_ ;
	wire _w3051_ ;
	wire _w3050_ ;
	wire _w3049_ ;
	wire _w3048_ ;
	wire _w3047_ ;
	wire _w3046_ ;
	wire _w3045_ ;
	wire _w3044_ ;
	wire _w3043_ ;
	wire _w3042_ ;
	wire _w3041_ ;
	wire _w3040_ ;
	wire _w3039_ ;
	wire _w3038_ ;
	wire _w3037_ ;
	wire _w3036_ ;
	wire _w3035_ ;
	wire _w3034_ ;
	wire _w3033_ ;
	wire _w3032_ ;
	wire _w3031_ ;
	wire _w3030_ ;
	wire _w3029_ ;
	wire _w3028_ ;
	wire _w3027_ ;
	wire _w3026_ ;
	wire _w3025_ ;
	wire _w3024_ ;
	wire _w3023_ ;
	wire _w3022_ ;
	wire _w3021_ ;
	wire _w3020_ ;
	wire _w3019_ ;
	wire _w3018_ ;
	wire _w3017_ ;
	wire _w3016_ ;
	wire _w3015_ ;
	wire _w3014_ ;
	wire _w3013_ ;
	wire _w3012_ ;
	wire _w3011_ ;
	wire _w3010_ ;
	wire _w3009_ ;
	wire _w3008_ ;
	wire _w3007_ ;
	wire _w3006_ ;
	wire _w3005_ ;
	wire _w3004_ ;
	wire _w3003_ ;
	wire _w3002_ ;
	wire _w3001_ ;
	wire _w3000_ ;
	wire _w2999_ ;
	wire _w2998_ ;
	wire _w2997_ ;
	wire _w2996_ ;
	wire _w2995_ ;
	wire _w2994_ ;
	wire _w2993_ ;
	wire _w2992_ ;
	wire _w2991_ ;
	wire _w2990_ ;
	wire _w2989_ ;
	wire _w2988_ ;
	wire _w2987_ ;
	wire _w2986_ ;
	wire _w2985_ ;
	wire _w2984_ ;
	wire _w2983_ ;
	wire _w2982_ ;
	wire _w2981_ ;
	wire _w2980_ ;
	wire _w2979_ ;
	wire _w2978_ ;
	wire _w2977_ ;
	wire _w2976_ ;
	wire _w2975_ ;
	wire _w2974_ ;
	wire _w2973_ ;
	wire _w2972_ ;
	wire _w2971_ ;
	wire _w2970_ ;
	wire _w2969_ ;
	wire _w2968_ ;
	wire _w2967_ ;
	wire _w2966_ ;
	wire _w2965_ ;
	wire _w2964_ ;
	wire _w2963_ ;
	wire _w2962_ ;
	wire _w2961_ ;
	wire _w2960_ ;
	wire _w2959_ ;
	wire _w2958_ ;
	wire _w2957_ ;
	wire _w2956_ ;
	wire _w2955_ ;
	wire _w2954_ ;
	wire _w2953_ ;
	wire _w2952_ ;
	wire _w2951_ ;
	wire _w2950_ ;
	wire _w2949_ ;
	wire _w2948_ ;
	wire _w2947_ ;
	wire _w2946_ ;
	wire _w2945_ ;
	wire _w2944_ ;
	wire _w2943_ ;
	wire _w2942_ ;
	wire _w2941_ ;
	wire _w2940_ ;
	wire _w2939_ ;
	wire _w2938_ ;
	wire _w2937_ ;
	wire _w2936_ ;
	wire _w2935_ ;
	wire _w2934_ ;
	wire _w2933_ ;
	wire _w2932_ ;
	wire _w2931_ ;
	wire _w2930_ ;
	wire _w2929_ ;
	wire _w2928_ ;
	wire _w2927_ ;
	wire _w2926_ ;
	wire _w2925_ ;
	wire _w2924_ ;
	wire _w2923_ ;
	wire _w2922_ ;
	wire _w2921_ ;
	wire _w2920_ ;
	wire _w2919_ ;
	wire _w2918_ ;
	wire _w2917_ ;
	wire _w2916_ ;
	wire _w2915_ ;
	wire _w2914_ ;
	wire _w2913_ ;
	wire _w2912_ ;
	wire _w2911_ ;
	wire _w2910_ ;
	wire _w2909_ ;
	wire _w2908_ ;
	wire _w2907_ ;
	wire _w2906_ ;
	wire _w2905_ ;
	wire _w2904_ ;
	wire _w2903_ ;
	wire _w2902_ ;
	wire _w2901_ ;
	wire _w2900_ ;
	wire _w2899_ ;
	wire _w2898_ ;
	wire _w2897_ ;
	wire _w2896_ ;
	wire _w2895_ ;
	wire _w2894_ ;
	wire _w2893_ ;
	wire _w2892_ ;
	wire _w2891_ ;
	wire _w2890_ ;
	wire _w2889_ ;
	wire _w2888_ ;
	wire _w2887_ ;
	wire _w2886_ ;
	wire _w2885_ ;
	wire _w2884_ ;
	wire _w2883_ ;
	wire _w2882_ ;
	wire _w2881_ ;
	wire _w2880_ ;
	wire _w2879_ ;
	wire _w2878_ ;
	wire _w2877_ ;
	wire _w2876_ ;
	wire _w2875_ ;
	wire _w2874_ ;
	wire _w2873_ ;
	wire _w2872_ ;
	wire _w2871_ ;
	wire _w2870_ ;
	wire _w2869_ ;
	wire _w2868_ ;
	wire _w2867_ ;
	wire _w2866_ ;
	wire _w2865_ ;
	wire _w2864_ ;
	wire _w2863_ ;
	wire _w2862_ ;
	wire _w2861_ ;
	wire _w2860_ ;
	wire _w2859_ ;
	wire _w2858_ ;
	wire _w2857_ ;
	wire _w2856_ ;
	wire _w2855_ ;
	wire _w2854_ ;
	wire _w2853_ ;
	wire _w2852_ ;
	wire _w2851_ ;
	wire _w2850_ ;
	wire _w2849_ ;
	wire _w2848_ ;
	wire _w2847_ ;
	wire _w2846_ ;
	wire _w2845_ ;
	wire _w2844_ ;
	wire _w2843_ ;
	wire _w2842_ ;
	wire _w2841_ ;
	wire _w2840_ ;
	wire _w2839_ ;
	wire _w2838_ ;
	wire _w2837_ ;
	wire _w2836_ ;
	wire _w2835_ ;
	wire _w2834_ ;
	wire _w2833_ ;
	wire _w2832_ ;
	wire _w2831_ ;
	wire _w2830_ ;
	wire _w2829_ ;
	wire _w2828_ ;
	wire _w2827_ ;
	wire _w2826_ ;
	wire _w2825_ ;
	wire _w2824_ ;
	wire _w2823_ ;
	wire _w2822_ ;
	wire _w2821_ ;
	wire _w2820_ ;
	wire _w2819_ ;
	wire _w2818_ ;
	wire _w2817_ ;
	wire _w2816_ ;
	wire _w2815_ ;
	wire _w2814_ ;
	wire _w2813_ ;
	wire _w2812_ ;
	wire _w2811_ ;
	wire _w2810_ ;
	wire _w2809_ ;
	wire _w2808_ ;
	wire _w2807_ ;
	wire _w2806_ ;
	wire _w2805_ ;
	wire _w2804_ ;
	wire _w2803_ ;
	wire _w2802_ ;
	wire _w2801_ ;
	wire _w2800_ ;
	wire _w2799_ ;
	wire _w2798_ ;
	wire _w2797_ ;
	wire _w2796_ ;
	wire _w2795_ ;
	wire _w2794_ ;
	wire _w2793_ ;
	wire _w2792_ ;
	wire _w2791_ ;
	wire _w2790_ ;
	wire _w2789_ ;
	wire _w2788_ ;
	wire _w2787_ ;
	wire _w2786_ ;
	wire _w2785_ ;
	wire _w2784_ ;
	wire _w2783_ ;
	wire _w2782_ ;
	wire _w2781_ ;
	wire _w2780_ ;
	wire _w2779_ ;
	wire _w2778_ ;
	wire _w2777_ ;
	wire _w2776_ ;
	wire _w2775_ ;
	wire _w2774_ ;
	wire _w2773_ ;
	wire _w2772_ ;
	wire _w2771_ ;
	wire _w2770_ ;
	wire _w2769_ ;
	wire _w2768_ ;
	wire _w2767_ ;
	wire _w2766_ ;
	wire _w2765_ ;
	wire _w2764_ ;
	wire _w2763_ ;
	wire _w2762_ ;
	wire _w2761_ ;
	wire _w2760_ ;
	wire _w2759_ ;
	wire _w2758_ ;
	wire _w2757_ ;
	wire _w2756_ ;
	wire _w2755_ ;
	wire _w2754_ ;
	wire _w2753_ ;
	wire _w2752_ ;
	wire _w2751_ ;
	wire _w2750_ ;
	wire _w2749_ ;
	wire _w2748_ ;
	wire _w2747_ ;
	wire _w2746_ ;
	wire _w2745_ ;
	wire _w2744_ ;
	wire _w2743_ ;
	wire _w2742_ ;
	wire _w2741_ ;
	wire _w2740_ ;
	wire _w2739_ ;
	wire _w2738_ ;
	wire _w2737_ ;
	wire _w2736_ ;
	wire _w2735_ ;
	wire _w2734_ ;
	wire _w2733_ ;
	wire _w2732_ ;
	wire _w2731_ ;
	wire _w2730_ ;
	wire _w2729_ ;
	wire _w2728_ ;
	wire _w2727_ ;
	wire _w2726_ ;
	wire _w2725_ ;
	wire _w2724_ ;
	wire _w2723_ ;
	wire _w2722_ ;
	wire _w2721_ ;
	wire _w2720_ ;
	wire _w2719_ ;
	wire _w2718_ ;
	wire _w2717_ ;
	wire _w2716_ ;
	wire _w2715_ ;
	wire _w2714_ ;
	wire _w2713_ ;
	wire _w2712_ ;
	wire _w2711_ ;
	wire _w2710_ ;
	wire _w2709_ ;
	wire _w2708_ ;
	wire _w2707_ ;
	wire _w2706_ ;
	wire _w2705_ ;
	wire _w2704_ ;
	wire _w2703_ ;
	wire _w2702_ ;
	wire _w2701_ ;
	wire _w2700_ ;
	wire _w2699_ ;
	wire _w2698_ ;
	wire _w2697_ ;
	wire _w2696_ ;
	wire _w2695_ ;
	wire _w2694_ ;
	wire _w2693_ ;
	wire _w2692_ ;
	wire _w2691_ ;
	wire _w2690_ ;
	wire _w2689_ ;
	wire _w2688_ ;
	wire _w2687_ ;
	wire _w2686_ ;
	wire _w2685_ ;
	wire _w2684_ ;
	wire _w2683_ ;
	wire _w2682_ ;
	wire _w2681_ ;
	wire _w2680_ ;
	wire _w2679_ ;
	wire _w2678_ ;
	wire _w2677_ ;
	wire _w2676_ ;
	wire _w2675_ ;
	wire _w2674_ ;
	wire _w2673_ ;
	wire _w2672_ ;
	wire _w2671_ ;
	wire _w2670_ ;
	wire _w2669_ ;
	wire _w2668_ ;
	wire _w2667_ ;
	wire _w2666_ ;
	wire _w2665_ ;
	wire _w2664_ ;
	wire _w2663_ ;
	wire _w2662_ ;
	wire _w2661_ ;
	wire _w2660_ ;
	wire _w2659_ ;
	wire _w2658_ ;
	wire _w2657_ ;
	wire _w2656_ ;
	wire _w2655_ ;
	wire _w2654_ ;
	wire _w2653_ ;
	wire _w2652_ ;
	wire _w2651_ ;
	wire _w2650_ ;
	wire _w2649_ ;
	wire _w2648_ ;
	wire _w2647_ ;
	wire _w2646_ ;
	wire _w2645_ ;
	wire _w2644_ ;
	wire _w2643_ ;
	wire _w2642_ ;
	wire _w2641_ ;
	wire _w2640_ ;
	wire _w2639_ ;
	wire _w2638_ ;
	wire _w2637_ ;
	wire _w2636_ ;
	wire _w2635_ ;
	wire _w2634_ ;
	wire _w2633_ ;
	wire _w2632_ ;
	wire _w2631_ ;
	wire _w2630_ ;
	wire _w2629_ ;
	wire _w2628_ ;
	wire _w2627_ ;
	wire _w2626_ ;
	wire _w2625_ ;
	wire _w2624_ ;
	wire _w2623_ ;
	wire _w2622_ ;
	wire _w2621_ ;
	wire _w2620_ ;
	wire _w2619_ ;
	wire _w2618_ ;
	wire _w2617_ ;
	wire _w2616_ ;
	wire _w2615_ ;
	wire _w2614_ ;
	wire _w2613_ ;
	wire _w2612_ ;
	wire _w2611_ ;
	wire _w2610_ ;
	wire _w2609_ ;
	wire _w2608_ ;
	wire _w2607_ ;
	wire _w2606_ ;
	wire _w2605_ ;
	wire _w2604_ ;
	wire _w2603_ ;
	wire _w2602_ ;
	wire _w2601_ ;
	wire _w2600_ ;
	wire _w2599_ ;
	wire _w2598_ ;
	wire _w2597_ ;
	wire _w2596_ ;
	wire _w2595_ ;
	wire _w2594_ ;
	wire _w2593_ ;
	wire _w2592_ ;
	wire _w2591_ ;
	wire _w2590_ ;
	wire _w2589_ ;
	wire _w2588_ ;
	wire _w2587_ ;
	wire _w2586_ ;
	wire _w2585_ ;
	wire _w2584_ ;
	wire _w2583_ ;
	wire _w2582_ ;
	wire _w2581_ ;
	wire _w2580_ ;
	wire _w2579_ ;
	wire _w2578_ ;
	wire _w2577_ ;
	wire _w2576_ ;
	wire _w2575_ ;
	wire _w2574_ ;
	wire _w2573_ ;
	wire _w2572_ ;
	wire _w2571_ ;
	wire _w2570_ ;
	wire _w2569_ ;
	wire _w2568_ ;
	wire _w2567_ ;
	wire _w2566_ ;
	wire _w2565_ ;
	wire _w2564_ ;
	wire _w2563_ ;
	wire _w2562_ ;
	wire _w2561_ ;
	wire _w2560_ ;
	wire _w2559_ ;
	wire _w2558_ ;
	wire _w2557_ ;
	wire _w2556_ ;
	wire _w2555_ ;
	wire _w2554_ ;
	wire _w2553_ ;
	wire _w2552_ ;
	wire _w2551_ ;
	wire _w2550_ ;
	wire _w2549_ ;
	wire _w2548_ ;
	wire _w2547_ ;
	wire _w2546_ ;
	wire _w2545_ ;
	wire _w2544_ ;
	wire _w2543_ ;
	wire _w2542_ ;
	wire _w2541_ ;
	wire _w2540_ ;
	wire _w2539_ ;
	wire _w2538_ ;
	wire _w2537_ ;
	wire _w2536_ ;
	wire _w2535_ ;
	wire _w2534_ ;
	wire _w2533_ ;
	wire _w2532_ ;
	wire _w2531_ ;
	wire _w2530_ ;
	wire _w2529_ ;
	wire _w2528_ ;
	wire _w2527_ ;
	wire _w2526_ ;
	wire _w2525_ ;
	wire _w2524_ ;
	wire _w2523_ ;
	wire _w2522_ ;
	wire _w2521_ ;
	wire _w2520_ ;
	wire _w2519_ ;
	wire _w2518_ ;
	wire _w2517_ ;
	wire _w2516_ ;
	wire _w2515_ ;
	wire _w2514_ ;
	wire _w2513_ ;
	wire _w2512_ ;
	wire _w2511_ ;
	wire _w2510_ ;
	wire _w2509_ ;
	wire _w2508_ ;
	wire _w2507_ ;
	wire _w2506_ ;
	wire _w2505_ ;
	wire _w2504_ ;
	wire _w2503_ ;
	wire _w2502_ ;
	wire _w2501_ ;
	wire _w2500_ ;
	wire _w2499_ ;
	wire _w2498_ ;
	wire _w2497_ ;
	wire _w2496_ ;
	wire _w2495_ ;
	wire _w2494_ ;
	wire _w2493_ ;
	wire _w1244_ ;
	wire _w1243_ ;
	wire _w1242_ ;
	wire _w1241_ ;
	wire _w1240_ ;
	wire _w1239_ ;
	wire _w1238_ ;
	wire _w1237_ ;
	wire _w1236_ ;
	wire _w1235_ ;
	wire _w1234_ ;
	wire _w1233_ ;
	wire _w1232_ ;
	wire _w1231_ ;
	wire _w1230_ ;
	wire _w1229_ ;
	wire _w1228_ ;
	wire _w1227_ ;
	wire _w1226_ ;
	wire _w1225_ ;
	wire _w1224_ ;
	wire _w1223_ ;
	wire _w1222_ ;
	wire _w1221_ ;
	wire _w1220_ ;
	wire _w1219_ ;
	wire _w1218_ ;
	wire _w1217_ ;
	wire _w1216_ ;
	wire _w1215_ ;
	wire _w1214_ ;
	wire _w1213_ ;
	wire _w1212_ ;
	wire _w1211_ ;
	wire _w1210_ ;
	wire _w1209_ ;
	wire _w1208_ ;
	wire _w1207_ ;
	wire _w1206_ ;
	wire _w1205_ ;
	wire _w1204_ ;
	wire _w1203_ ;
	wire _w1202_ ;
	wire _w1201_ ;
	wire _w1200_ ;
	wire _w1199_ ;
	wire _w1198_ ;
	wire _w1197_ ;
	wire _w1196_ ;
	wire _w1195_ ;
	wire _w1194_ ;
	wire _w1193_ ;
	wire _w1192_ ;
	wire _w1191_ ;
	wire _w1190_ ;
	wire _w1189_ ;
	wire _w1188_ ;
	wire _w1187_ ;
	wire _w1186_ ;
	wire _w1185_ ;
	wire _w1184_ ;
	wire _w1183_ ;
	wire _w1182_ ;
	wire _w1181_ ;
	wire _w1180_ ;
	wire _w1179_ ;
	wire _w1178_ ;
	wire _w1177_ ;
	wire _w1176_ ;
	wire _w1175_ ;
	wire _w1174_ ;
	wire _w1173_ ;
	wire _w1172_ ;
	wire _w1171_ ;
	wire _w1170_ ;
	wire _w1169_ ;
	wire _w1168_ ;
	wire _w1167_ ;
	wire _w1166_ ;
	wire _w1165_ ;
	wire _w1164_ ;
	wire _w1163_ ;
	wire _w1162_ ;
	wire _w1161_ ;
	wire _w1160_ ;
	wire _w1159_ ;
	wire _w1158_ ;
	wire _w1157_ ;
	wire _w1156_ ;
	wire _w1155_ ;
	wire _w1154_ ;
	wire _w1153_ ;
	wire _w1152_ ;
	wire _w1151_ ;
	wire _w1150_ ;
	wire _w1149_ ;
	wire _w1148_ ;
	wire _w1147_ ;
	wire _w1146_ ;
	wire _w1145_ ;
	wire _w1144_ ;
	wire _w1143_ ;
	wire _w1142_ ;
	wire _w1141_ ;
	wire _w1140_ ;
	wire _w1139_ ;
	wire _w1138_ ;
	wire _w1137_ ;
	wire _w1136_ ;
	wire _w1135_ ;
	wire _w1134_ ;
	wire _w1133_ ;
	wire _w1132_ ;
	wire _w1131_ ;
	wire _w1130_ ;
	wire _w1129_ ;
	wire _w1128_ ;
	wire _w1127_ ;
	wire _w1126_ ;
	wire _w1125_ ;
	wire _w1124_ ;
	wire _w1123_ ;
	wire _w1122_ ;
	wire _w1121_ ;
	wire _w1120_ ;
	wire _w1119_ ;
	wire _w1118_ ;
	wire _w1117_ ;
	wire _w1116_ ;
	wire _w1115_ ;
	wire _w1114_ ;
	wire _w1113_ ;
	wire _w1112_ ;
	wire _w1111_ ;
	wire _w1110_ ;
	wire _w1109_ ;
	wire _w1108_ ;
	wire _w1107_ ;
	wire _w1106_ ;
	wire _w1105_ ;
	wire _w1104_ ;
	wire _w1103_ ;
	wire _w1102_ ;
	wire _w1101_ ;
	wire _w1100_ ;
	wire _w1099_ ;
	wire _w1098_ ;
	wire _w1097_ ;
	wire _w1096_ ;
	wire _w1095_ ;
	wire _w1094_ ;
	wire _w1093_ ;
	wire _w1092_ ;
	wire _w1091_ ;
	wire _w1090_ ;
	wire _w1089_ ;
	wire _w1088_ ;
	wire _w1087_ ;
	wire _w1086_ ;
	wire _w1085_ ;
	wire _w1084_ ;
	wire _w1083_ ;
	wire _w1082_ ;
	wire _w1081_ ;
	wire _w1080_ ;
	wire _w1079_ ;
	wire _w1078_ ;
	wire _w1077_ ;
	wire _w1076_ ;
	wire _w1075_ ;
	wire _w1074_ ;
	wire _w1073_ ;
	wire _w1072_ ;
	wire _w1071_ ;
	wire _w1070_ ;
	wire _w1069_ ;
	wire _w1068_ ;
	wire _w1067_ ;
	wire _w1066_ ;
	wire _w1065_ ;
	wire _w1064_ ;
	wire _w1063_ ;
	wire _w1062_ ;
	wire _w1061_ ;
	wire _w1060_ ;
	wire _w1059_ ;
	wire _w1058_ ;
	wire _w1057_ ;
	wire _w1056_ ;
	wire _w1055_ ;
	wire _w1054_ ;
	wire _w1053_ ;
	wire _w1052_ ;
	wire _w1051_ ;
	wire _w1050_ ;
	wire _w1049_ ;
	wire _w1048_ ;
	wire _w1047_ ;
	wire _w1046_ ;
	wire _w1045_ ;
	wire _w1044_ ;
	wire _w1043_ ;
	wire _w1042_ ;
	wire _w1041_ ;
	wire _w1040_ ;
	wire _w1039_ ;
	wire _w1038_ ;
	wire _w1037_ ;
	wire _w1036_ ;
	wire _w1035_ ;
	wire _w1034_ ;
	wire _w1033_ ;
	wire _w1032_ ;
	wire _w1031_ ;
	wire _w1030_ ;
	wire _w1029_ ;
	wire _w1028_ ;
	wire _w1027_ ;
	wire _w1026_ ;
	wire _w1025_ ;
	wire _w1024_ ;
	wire _w1023_ ;
	wire _w1022_ ;
	wire _w1021_ ;
	wire _w1020_ ;
	wire _w1019_ ;
	wire _w1018_ ;
	wire _w1017_ ;
	wire _w1016_ ;
	wire _w1015_ ;
	wire _w1014_ ;
	wire _w1013_ ;
	wire _w1012_ ;
	wire _w1011_ ;
	wire _w1010_ ;
	wire _w1009_ ;
	wire _w1008_ ;
	wire _w1007_ ;
	wire _w1006_ ;
	wire _w1005_ ;
	wire _w1004_ ;
	wire _w1003_ ;
	wire _w1002_ ;
	wire _w1001_ ;
	wire _w1000_ ;
	wire _w999_ ;
	wire _w998_ ;
	wire _w997_ ;
	wire _w996_ ;
	wire _w995_ ;
	wire _w994_ ;
	wire _w993_ ;
	wire _w992_ ;
	wire _w991_ ;
	wire _w990_ ;
	wire _w989_ ;
	wire _w988_ ;
	wire _w987_ ;
	wire _w986_ ;
	wire _w985_ ;
	wire _w984_ ;
	wire _w983_ ;
	wire _w982_ ;
	wire _w981_ ;
	wire _w980_ ;
	wire _w979_ ;
	wire _w978_ ;
	wire _w977_ ;
	wire _w976_ ;
	wire _w975_ ;
	wire _w974_ ;
	wire _w973_ ;
	wire _w972_ ;
	wire _w971_ ;
	wire _w970_ ;
	wire _w969_ ;
	wire _w968_ ;
	wire _w967_ ;
	wire _w966_ ;
	wire _w965_ ;
	wire _w964_ ;
	wire _w963_ ;
	wire _w962_ ;
	wire _w961_ ;
	wire _w960_ ;
	wire _w959_ ;
	wire _w958_ ;
	wire _w957_ ;
	wire _w956_ ;
	wire _w955_ ;
	wire _w954_ ;
	wire _w953_ ;
	wire _w952_ ;
	wire _w951_ ;
	wire _w950_ ;
	wire _w949_ ;
	wire _w948_ ;
	wire _w947_ ;
	wire _w946_ ;
	wire _w945_ ;
	wire _w944_ ;
	wire _w943_ ;
	wire _w942_ ;
	wire _w941_ ;
	wire _w940_ ;
	wire _w939_ ;
	wire _w938_ ;
	wire _w937_ ;
	wire _w936_ ;
	wire _w935_ ;
	wire _w934_ ;
	wire _w933_ ;
	wire _w932_ ;
	wire _w931_ ;
	wire _w930_ ;
	wire _w929_ ;
	wire _w928_ ;
	wire _w927_ ;
	wire _w926_ ;
	wire _w925_ ;
	wire _w924_ ;
	wire _w923_ ;
	wire _w922_ ;
	wire _w921_ ;
	wire _w920_ ;
	wire _w919_ ;
	wire _w918_ ;
	wire _w917_ ;
	wire _w916_ ;
	wire _w915_ ;
	wire _w914_ ;
	wire _w913_ ;
	wire _w912_ ;
	wire _w911_ ;
	wire _w910_ ;
	wire _w909_ ;
	wire _w908_ ;
	wire _w907_ ;
	wire _w906_ ;
	wire _w905_ ;
	wire _w904_ ;
	wire _w903_ ;
	wire _w902_ ;
	wire _w901_ ;
	wire _w900_ ;
	wire _w899_ ;
	wire _w898_ ;
	wire _w897_ ;
	wire _w896_ ;
	wire _w895_ ;
	wire _w894_ ;
	wire _w893_ ;
	wire _w892_ ;
	wire _w891_ ;
	wire _w890_ ;
	wire _w889_ ;
	wire _w888_ ;
	wire _w887_ ;
	wire _w886_ ;
	wire _w885_ ;
	wire _w884_ ;
	wire _w883_ ;
	wire _w882_ ;
	wire _w881_ ;
	wire _w880_ ;
	wire _w879_ ;
	wire _w878_ ;
	wire _w877_ ;
	wire _w876_ ;
	wire _w875_ ;
	wire _w874_ ;
	wire _w873_ ;
	wire _w872_ ;
	wire _w871_ ;
	wire _w870_ ;
	wire _w869_ ;
	wire _w868_ ;
	wire _w867_ ;
	wire _w866_ ;
	wire _w865_ ;
	wire _w864_ ;
	wire _w863_ ;
	wire _w862_ ;
	wire _w861_ ;
	wire _w860_ ;
	wire _w859_ ;
	wire _w858_ ;
	wire _w857_ ;
	wire _w856_ ;
	wire _w855_ ;
	wire _w854_ ;
	wire _w853_ ;
	wire _w852_ ;
	wire _w851_ ;
	wire _w850_ ;
	wire _w849_ ;
	wire _w848_ ;
	wire _w847_ ;
	wire _w846_ ;
	wire _w845_ ;
	wire _w844_ ;
	wire _w843_ ;
	wire _w842_ ;
	wire _w841_ ;
	wire _w840_ ;
	wire _w839_ ;
	wire _w838_ ;
	wire _w837_ ;
	wire _w836_ ;
	wire _w835_ ;
	wire _w834_ ;
	wire _w833_ ;
	wire _w832_ ;
	wire _w831_ ;
	wire _w830_ ;
	wire _w829_ ;
	wire _w828_ ;
	wire _w827_ ;
	wire _w826_ ;
	wire _w825_ ;
	wire _w824_ ;
	wire _w823_ ;
	wire _w822_ ;
	wire _w821_ ;
	wire _w820_ ;
	wire _w819_ ;
	wire _w818_ ;
	wire _w817_ ;
	wire _w816_ ;
	wire _w815_ ;
	wire _w814_ ;
	wire _w813_ ;
	wire _w812_ ;
	wire _w811_ ;
	wire _w810_ ;
	wire _w809_ ;
	wire _w808_ ;
	wire _w807_ ;
	wire _w806_ ;
	wire _w805_ ;
	wire _w804_ ;
	wire _w803_ ;
	wire _w802_ ;
	wire _w801_ ;
	wire _w800_ ;
	wire _w799_ ;
	wire _w798_ ;
	wire _w797_ ;
	wire _w796_ ;
	wire _w795_ ;
	wire _w794_ ;
	wire _w793_ ;
	wire _w792_ ;
	wire _w791_ ;
	wire _w790_ ;
	wire _w789_ ;
	wire _w788_ ;
	wire _w787_ ;
	wire _w786_ ;
	wire _w785_ ;
	wire _w784_ ;
	wire _w783_ ;
	wire _w782_ ;
	wire _w781_ ;
	wire _w780_ ;
	wire _w779_ ;
	wire _w778_ ;
	wire _w777_ ;
	wire _w776_ ;
	wire _w775_ ;
	wire _w774_ ;
	wire _w773_ ;
	wire _w772_ ;
	wire _w771_ ;
	wire _w770_ ;
	wire _w769_ ;
	wire _w768_ ;
	wire _w767_ ;
	wire _w766_ ;
	wire _w765_ ;
	wire _w764_ ;
	wire _w763_ ;
	wire _w762_ ;
	wire _w761_ ;
	wire _w760_ ;
	wire _w759_ ;
	wire _w758_ ;
	wire _w757_ ;
	wire _w756_ ;
	wire _w755_ ;
	wire _w754_ ;
	wire _w753_ ;
	wire _w752_ ;
	wire _w751_ ;
	wire _w750_ ;
	wire _w749_ ;
	wire _w748_ ;
	wire _w747_ ;
	wire _w746_ ;
	wire _w745_ ;
	wire _w744_ ;
	wire _w743_ ;
	wire _w742_ ;
	wire _w741_ ;
	wire _w740_ ;
	wire _w739_ ;
	wire _w738_ ;
	wire _w737_ ;
	wire _w736_ ;
	wire _w735_ ;
	wire _w734_ ;
	wire _w733_ ;
	wire _w732_ ;
	wire _w731_ ;
	wire _w730_ ;
	wire _w729_ ;
	wire _w728_ ;
	wire _w727_ ;
	wire _w726_ ;
	wire _w725_ ;
	wire _w724_ ;
	wire _w723_ ;
	wire _w722_ ;
	wire _w721_ ;
	wire _w720_ ;
	wire _w719_ ;
	wire _w718_ ;
	wire _w717_ ;
	wire _w716_ ;
	wire _w715_ ;
	wire _w714_ ;
	wire _w713_ ;
	wire _w712_ ;
	wire _w711_ ;
	wire _w710_ ;
	wire _w709_ ;
	wire _w708_ ;
	wire _w707_ ;
	wire _w706_ ;
	wire _w705_ ;
	wire _w704_ ;
	wire _w703_ ;
	wire _w702_ ;
	wire _w701_ ;
	wire _w700_ ;
	wire _w699_ ;
	wire _w698_ ;
	wire _w697_ ;
	wire _w696_ ;
	wire _w695_ ;
	wire _w694_ ;
	wire _w693_ ;
	wire _w692_ ;
	wire _w691_ ;
	wire _w690_ ;
	wire _w689_ ;
	wire _w688_ ;
	wire _w687_ ;
	wire _w686_ ;
	wire _w685_ ;
	wire _w684_ ;
	wire _w683_ ;
	wire _w682_ ;
	wire _w681_ ;
	wire _w680_ ;
	wire _w679_ ;
	wire _w678_ ;
	wire _w677_ ;
	wire _w392_ ;
	wire _w391_ ;
	wire _w390_ ;
	wire _w389_ ;
	wire _w388_ ;
	wire _w387_ ;
	wire _w386_ ;
	wire _w385_ ;
	wire _w384_ ;
	wire _w383_ ;
	wire _w382_ ;
	wire _w381_ ;
	wire _w380_ ;
	wire _w379_ ;
	wire _w378_ ;
	wire _w377_ ;
	wire _w376_ ;
	wire _w375_ ;
	wire _w374_ ;
	wire _w373_ ;
	wire _w372_ ;
	wire _w371_ ;
	wire _w370_ ;
	wire _w369_ ;
	wire _w368_ ;
	wire _w367_ ;
	wire _w366_ ;
	wire _w365_ ;
	wire _w364_ ;
	wire _w363_ ;
	wire _w362_ ;
	wire _w361_ ;
	wire _w360_ ;
	wire _w359_ ;
	wire _w358_ ;
	wire _w357_ ;
	wire _w356_ ;
	wire _w355_ ;
	wire _w354_ ;
	wire _w353_ ;
	wire _w352_ ;
	wire _w351_ ;
	wire _w350_ ;
	wire _w349_ ;
	wire _w348_ ;
	wire _w347_ ;
	wire _w346_ ;
	wire _w345_ ;
	wire _w344_ ;
	wire _w343_ ;
	wire _w342_ ;
	wire _w341_ ;
	wire _w340_ ;
	wire _w339_ ;
	wire _w338_ ;
	wire _w337_ ;
	wire _w336_ ;
	wire _w335_ ;
	wire _w334_ ;
	wire _w333_ ;
	wire _w332_ ;
	wire _w331_ ;
	wire _w330_ ;
	wire _w329_ ;
	wire _w328_ ;
	wire _w327_ ;
	wire _w326_ ;
	wire _w325_ ;
	wire _w324_ ;
	wire _w323_ ;
	wire _w322_ ;
	wire _w321_ ;
	wire _w320_ ;
	wire _w319_ ;
	wire _w318_ ;
	wire _w317_ ;
	wire _w316_ ;
	wire _w315_ ;
	wire _w314_ ;
	wire _w313_ ;
	wire _w312_ ;
	wire _w311_ ;
	wire _w310_ ;
	wire _w309_ ;
	wire _w308_ ;
	wire _w307_ ;
	wire _w306_ ;
	wire _w305_ ;
	wire _w304_ ;
	wire _w303_ ;
	wire _w302_ ;
	wire _w301_ ;
	wire _w300_ ;
	wire _w299_ ;
	wire _w298_ ;
	wire _w297_ ;
	wire _w296_ ;
	wire _w295_ ;
	wire _w294_ ;
	wire _w293_ ;
	wire _w292_ ;
	wire _w291_ ;
	wire _w290_ ;
	wire _w289_ ;
	wire _w288_ ;
	wire _w287_ ;
	wire _w286_ ;
	wire _w285_ ;
	wire _w284_ ;
	wire _w283_ ;
	wire _w282_ ;
	wire _w281_ ;
	wire _w280_ ;
	wire _w279_ ;
	wire _w278_ ;
	wire _w277_ ;
	wire _w276_ ;
	wire _w275_ ;
	wire _w274_ ;
	wire _w273_ ;
	wire _w272_ ;
	wire _w271_ ;
	wire _w270_ ;
	wire _w269_ ;
	wire _w268_ ;
	wire _w267_ ;
	wire _w266_ ;
	wire _w265_ ;
	wire _w264_ ;
	wire _w263_ ;
	wire _w194_ ;
	wire _w193_ ;
	wire _w192_ ;
	wire _w191_ ;
	wire _w190_ ;
	wire _w189_ ;
	wire _w188_ ;
	wire _w187_ ;
	wire _w186_ ;
	wire _w185_ ;
	wire _w184_ ;
	wire _w183_ ;
	wire _w182_ ;
	wire _w181_ ;
	wire _w180_ ;
	wire _w179_ ;
	wire _w178_ ;
	wire _w177_ ;
	wire _w176_ ;
	wire _w175_ ;
	wire _w174_ ;
	wire _w173_ ;
	wire _w172_ ;
	wire _w171_ ;
	wire _w170_ ;
	wire _w169_ ;
	wire _w168_ ;
	wire _w167_ ;
	wire _w166_ ;
	wire _w165_ ;
	wire _w148_ ;
	wire _w147_ ;
	wire _w146_ ;
	wire _w145_ ;
	wire _w144_ ;
	wire _w143_ ;
	wire _w142_ ;
	wire _w141_ ;
	wire _w140_ ;
	wire _w139_ ;
	wire _w138_ ;
	wire _w137_ ;
	wire _w136_ ;
	wire _w149_ ;
	wire _w150_ ;
	wire _w151_ ;
	wire _w152_ ;
	wire _w153_ ;
	wire _w154_ ;
	wire _w155_ ;
	wire _w156_ ;
	wire _w157_ ;
	wire _w158_ ;
	wire _w159_ ;
	wire _w160_ ;
	wire _w161_ ;
	wire _w162_ ;
	wire _w163_ ;
	wire _w164_ ;
	wire _w195_ ;
	wire _w196_ ;
	wire _w197_ ;
	wire _w198_ ;
	wire _w199_ ;
	wire _w200_ ;
	wire _w201_ ;
	wire _w202_ ;
	wire _w203_ ;
	wire _w204_ ;
	wire _w205_ ;
	wire _w206_ ;
	wire _w207_ ;
	wire _w208_ ;
	wire _w209_ ;
	wire _w210_ ;
	wire _w211_ ;
	wire _w212_ ;
	wire _w213_ ;
	wire _w214_ ;
	wire _w215_ ;
	wire _w216_ ;
	wire _w217_ ;
	wire _w218_ ;
	wire _w219_ ;
	wire _w220_ ;
	wire _w221_ ;
	wire _w222_ ;
	wire _w223_ ;
	wire _w224_ ;
	wire _w225_ ;
	wire _w226_ ;
	wire _w227_ ;
	wire _w228_ ;
	wire _w229_ ;
	wire _w230_ ;
	wire _w231_ ;
	wire _w232_ ;
	wire _w233_ ;
	wire _w234_ ;
	wire _w235_ ;
	wire _w236_ ;
	wire _w237_ ;
	wire _w238_ ;
	wire _w239_ ;
	wire _w240_ ;
	wire _w241_ ;
	wire _w242_ ;
	wire _w243_ ;
	wire _w244_ ;
	wire _w245_ ;
	wire _w246_ ;
	wire _w247_ ;
	wire _w248_ ;
	wire _w249_ ;
	wire _w250_ ;
	wire _w251_ ;
	wire _w252_ ;
	wire _w253_ ;
	wire _w254_ ;
	wire _w255_ ;
	wire _w256_ ;
	wire _w257_ ;
	wire _w258_ ;
	wire _w259_ ;
	wire _w260_ ;
	wire _w261_ ;
	wire _w262_ ;
	wire _w393_ ;
	wire _w394_ ;
	wire _w395_ ;
	wire _w396_ ;
	wire _w397_ ;
	wire _w398_ ;
	wire _w399_ ;
	wire _w400_ ;
	wire _w401_ ;
	wire _w402_ ;
	wire _w403_ ;
	wire _w404_ ;
	wire _w405_ ;
	wire _w406_ ;
	wire _w407_ ;
	wire _w408_ ;
	wire _w409_ ;
	wire _w410_ ;
	wire _w411_ ;
	wire _w412_ ;
	wire _w413_ ;
	wire _w414_ ;
	wire _w415_ ;
	wire _w416_ ;
	wire _w417_ ;
	wire _w418_ ;
	wire _w419_ ;
	wire _w420_ ;
	wire _w421_ ;
	wire _w422_ ;
	wire _w423_ ;
	wire _w424_ ;
	wire _w425_ ;
	wire _w426_ ;
	wire _w427_ ;
	wire _w428_ ;
	wire _w429_ ;
	wire _w430_ ;
	wire _w431_ ;
	wire _w432_ ;
	wire _w433_ ;
	wire _w434_ ;
	wire _w435_ ;
	wire _w436_ ;
	wire _w437_ ;
	wire _w438_ ;
	wire _w439_ ;
	wire _w440_ ;
	wire _w441_ ;
	wire _w442_ ;
	wire _w443_ ;
	wire _w444_ ;
	wire _w445_ ;
	wire _w446_ ;
	wire _w447_ ;
	wire _w448_ ;
	wire _w449_ ;
	wire _w450_ ;
	wire _w451_ ;
	wire _w452_ ;
	wire _w453_ ;
	wire _w454_ ;
	wire _w455_ ;
	wire _w456_ ;
	wire _w457_ ;
	wire _w458_ ;
	wire _w459_ ;
	wire _w460_ ;
	wire _w461_ ;
	wire _w462_ ;
	wire _w463_ ;
	wire _w464_ ;
	wire _w465_ ;
	wire _w466_ ;
	wire _w467_ ;
	wire _w468_ ;
	wire _w469_ ;
	wire _w470_ ;
	wire _w471_ ;
	wire _w472_ ;
	wire _w473_ ;
	wire _w474_ ;
	wire _w475_ ;
	wire _w476_ ;
	wire _w477_ ;
	wire _w478_ ;
	wire _w479_ ;
	wire _w480_ ;
	wire _w481_ ;
	wire _w482_ ;
	wire _w483_ ;
	wire _w484_ ;
	wire _w485_ ;
	wire _w486_ ;
	wire _w487_ ;
	wire _w488_ ;
	wire _w489_ ;
	wire _w490_ ;
	wire _w491_ ;
	wire _w492_ ;
	wire _w493_ ;
	wire _w494_ ;
	wire _w495_ ;
	wire _w496_ ;
	wire _w497_ ;
	wire _w498_ ;
	wire _w499_ ;
	wire _w500_ ;
	wire _w501_ ;
	wire _w502_ ;
	wire _w503_ ;
	wire _w504_ ;
	wire _w505_ ;
	wire _w506_ ;
	wire _w507_ ;
	wire _w508_ ;
	wire _w509_ ;
	wire _w510_ ;
	wire _w511_ ;
	wire _w512_ ;
	wire _w513_ ;
	wire _w514_ ;
	wire _w515_ ;
	wire _w516_ ;
	wire _w517_ ;
	wire _w518_ ;
	wire _w519_ ;
	wire _w520_ ;
	wire _w521_ ;
	wire _w522_ ;
	wire _w523_ ;
	wire _w524_ ;
	wire _w525_ ;
	wire _w526_ ;
	wire _w527_ ;
	wire _w528_ ;
	wire _w529_ ;
	wire _w530_ ;
	wire _w531_ ;
	wire _w532_ ;
	wire _w533_ ;
	wire _w534_ ;
	wire _w535_ ;
	wire _w536_ ;
	wire _w537_ ;
	wire _w538_ ;
	wire _w539_ ;
	wire _w540_ ;
	wire _w541_ ;
	wire _w542_ ;
	wire _w543_ ;
	wire _w544_ ;
	wire _w545_ ;
	wire _w546_ ;
	wire _w547_ ;
	wire _w548_ ;
	wire _w549_ ;
	wire _w550_ ;
	wire _w551_ ;
	wire _w552_ ;
	wire _w553_ ;
	wire _w554_ ;
	wire _w555_ ;
	wire _w556_ ;
	wire _w557_ ;
	wire _w558_ ;
	wire _w559_ ;
	wire _w560_ ;
	wire _w561_ ;
	wire _w562_ ;
	wire _w563_ ;
	wire _w564_ ;
	wire _w565_ ;
	wire _w566_ ;
	wire _w567_ ;
	wire _w568_ ;
	wire _w569_ ;
	wire _w570_ ;
	wire _w571_ ;
	wire _w572_ ;
	wire _w573_ ;
	wire _w574_ ;
	wire _w575_ ;
	wire _w576_ ;
	wire _w577_ ;
	wire _w578_ ;
	wire _w579_ ;
	wire _w580_ ;
	wire _w581_ ;
	wire _w582_ ;
	wire _w583_ ;
	wire _w584_ ;
	wire _w585_ ;
	wire _w586_ ;
	wire _w587_ ;
	wire _w588_ ;
	wire _w589_ ;
	wire _w590_ ;
	wire _w591_ ;
	wire _w592_ ;
	wire _w593_ ;
	wire _w594_ ;
	wire _w595_ ;
	wire _w596_ ;
	wire _w597_ ;
	wire _w598_ ;
	wire _w599_ ;
	wire _w600_ ;
	wire _w601_ ;
	wire _w602_ ;
	wire _w603_ ;
	wire _w604_ ;
	wire _w605_ ;
	wire _w606_ ;
	wire _w607_ ;
	wire _w608_ ;
	wire _w609_ ;
	wire _w610_ ;
	wire _w611_ ;
	wire _w612_ ;
	wire _w613_ ;
	wire _w614_ ;
	wire _w615_ ;
	wire _w616_ ;
	wire _w617_ ;
	wire _w618_ ;
	wire _w619_ ;
	wire _w620_ ;
	wire _w621_ ;
	wire _w622_ ;
	wire _w623_ ;
	wire _w624_ ;
	wire _w625_ ;
	wire _w626_ ;
	wire _w627_ ;
	wire _w628_ ;
	wire _w629_ ;
	wire _w630_ ;
	wire _w631_ ;
	wire _w632_ ;
	wire _w633_ ;
	wire _w634_ ;
	wire _w635_ ;
	wire _w636_ ;
	wire _w637_ ;
	wire _w638_ ;
	wire _w639_ ;
	wire _w640_ ;
	wire _w641_ ;
	wire _w642_ ;
	wire _w643_ ;
	wire _w644_ ;
	wire _w645_ ;
	wire _w646_ ;
	wire _w647_ ;
	wire _w648_ ;
	wire _w649_ ;
	wire _w650_ ;
	wire _w651_ ;
	wire _w652_ ;
	wire _w653_ ;
	wire _w654_ ;
	wire _w655_ ;
	wire _w656_ ;
	wire _w657_ ;
	wire _w658_ ;
	wire _w659_ ;
	wire _w660_ ;
	wire _w661_ ;
	wire _w662_ ;
	wire _w663_ ;
	wire _w664_ ;
	wire _w665_ ;
	wire _w666_ ;
	wire _w667_ ;
	wire _w668_ ;
	wire _w669_ ;
	wire _w670_ ;
	wire _w671_ ;
	wire _w672_ ;
	wire _w673_ ;
	wire _w674_ ;
	wire _w675_ ;
	wire _w676_ ;
	wire _w1245_ ;
	wire _w1246_ ;
	wire _w1247_ ;
	wire _w1248_ ;
	wire _w1249_ ;
	wire _w1250_ ;
	wire _w1251_ ;
	wire _w1252_ ;
	wire _w1253_ ;
	wire _w1254_ ;
	wire _w1255_ ;
	wire _w1256_ ;
	wire _w1257_ ;
	wire _w1258_ ;
	wire _w1259_ ;
	wire _w1260_ ;
	wire _w1261_ ;
	wire _w1262_ ;
	wire _w1263_ ;
	wire _w1264_ ;
	wire _w1265_ ;
	wire _w1266_ ;
	wire _w1267_ ;
	wire _w1268_ ;
	wire _w1269_ ;
	wire _w1270_ ;
	wire _w1271_ ;
	wire _w1272_ ;
	wire _w1273_ ;
	wire _w1274_ ;
	wire _w1275_ ;
	wire _w1276_ ;
	wire _w1277_ ;
	wire _w1278_ ;
	wire _w1279_ ;
	wire _w1280_ ;
	wire _w1281_ ;
	wire _w1282_ ;
	wire _w1283_ ;
	wire _w1284_ ;
	wire _w1285_ ;
	wire _w1286_ ;
	wire _w1287_ ;
	wire _w1288_ ;
	wire _w1289_ ;
	wire _w1290_ ;
	wire _w1291_ ;
	wire _w1292_ ;
	wire _w1293_ ;
	wire _w1294_ ;
	wire _w1295_ ;
	wire _w1296_ ;
	wire _w1297_ ;
	wire _w1298_ ;
	wire _w1299_ ;
	wire _w1300_ ;
	wire _w1301_ ;
	wire _w1302_ ;
	wire _w1303_ ;
	wire _w1304_ ;
	wire _w1305_ ;
	wire _w1306_ ;
	wire _w1307_ ;
	wire _w1308_ ;
	wire _w1309_ ;
	wire _w1310_ ;
	wire _w1311_ ;
	wire _w1312_ ;
	wire _w1313_ ;
	wire _w1314_ ;
	wire _w1315_ ;
	wire _w1316_ ;
	wire _w1317_ ;
	wire _w1318_ ;
	wire _w1319_ ;
	wire _w1320_ ;
	wire _w1321_ ;
	wire _w1322_ ;
	wire _w1323_ ;
	wire _w1324_ ;
	wire _w1325_ ;
	wire _w1326_ ;
	wire _w1327_ ;
	wire _w1328_ ;
	wire _w1329_ ;
	wire _w1330_ ;
	wire _w1331_ ;
	wire _w1332_ ;
	wire _w1333_ ;
	wire _w1334_ ;
	wire _w1335_ ;
	wire _w1336_ ;
	wire _w1337_ ;
	wire _w1338_ ;
	wire _w1339_ ;
	wire _w1340_ ;
	wire _w1341_ ;
	wire _w1342_ ;
	wire _w1343_ ;
	wire _w1344_ ;
	wire _w1345_ ;
	wire _w1346_ ;
	wire _w1347_ ;
	wire _w1348_ ;
	wire _w1349_ ;
	wire _w1350_ ;
	wire _w1351_ ;
	wire _w1352_ ;
	wire _w1353_ ;
	wire _w1354_ ;
	wire _w1355_ ;
	wire _w1356_ ;
	wire _w1357_ ;
	wire _w1358_ ;
	wire _w1359_ ;
	wire _w1360_ ;
	wire _w1361_ ;
	wire _w1362_ ;
	wire _w1363_ ;
	wire _w1364_ ;
	wire _w1365_ ;
	wire _w1366_ ;
	wire _w1367_ ;
	wire _w1368_ ;
	wire _w1369_ ;
	wire _w1370_ ;
	wire _w1371_ ;
	wire _w1372_ ;
	wire _w1373_ ;
	wire _w1374_ ;
	wire _w1375_ ;
	wire _w1376_ ;
	wire _w1377_ ;
	wire _w1378_ ;
	wire _w1379_ ;
	wire _w1380_ ;
	wire _w1381_ ;
	wire _w1382_ ;
	wire _w1383_ ;
	wire _w1384_ ;
	wire _w1385_ ;
	wire _w1386_ ;
	wire _w1387_ ;
	wire _w1388_ ;
	wire _w1389_ ;
	wire _w1390_ ;
	wire _w1391_ ;
	wire _w1392_ ;
	wire _w1393_ ;
	wire _w1394_ ;
	wire _w1395_ ;
	wire _w1396_ ;
	wire _w1397_ ;
	wire _w1398_ ;
	wire _w1399_ ;
	wire _w1400_ ;
	wire _w1401_ ;
	wire _w1402_ ;
	wire _w1403_ ;
	wire _w1404_ ;
	wire _w1405_ ;
	wire _w1406_ ;
	wire _w1407_ ;
	wire _w1408_ ;
	wire _w1409_ ;
	wire _w1410_ ;
	wire _w1411_ ;
	wire _w1412_ ;
	wire _w1413_ ;
	wire _w1414_ ;
	wire _w1415_ ;
	wire _w1416_ ;
	wire _w1417_ ;
	wire _w1418_ ;
	wire _w1419_ ;
	wire _w1420_ ;
	wire _w1421_ ;
	wire _w1422_ ;
	wire _w1423_ ;
	wire _w1424_ ;
	wire _w1425_ ;
	wire _w1426_ ;
	wire _w1427_ ;
	wire _w1428_ ;
	wire _w1429_ ;
	wire _w1430_ ;
	wire _w1431_ ;
	wire _w1432_ ;
	wire _w1433_ ;
	wire _w1434_ ;
	wire _w1435_ ;
	wire _w1436_ ;
	wire _w1437_ ;
	wire _w1438_ ;
	wire _w1439_ ;
	wire _w1440_ ;
	wire _w1441_ ;
	wire _w1442_ ;
	wire _w1443_ ;
	wire _w1444_ ;
	wire _w1445_ ;
	wire _w1446_ ;
	wire _w1447_ ;
	wire _w1448_ ;
	wire _w1449_ ;
	wire _w1450_ ;
	wire _w1451_ ;
	wire _w1452_ ;
	wire _w1453_ ;
	wire _w1454_ ;
	wire _w1455_ ;
	wire _w1456_ ;
	wire _w1457_ ;
	wire _w1458_ ;
	wire _w1459_ ;
	wire _w1460_ ;
	wire _w1461_ ;
	wire _w1462_ ;
	wire _w1463_ ;
	wire _w1464_ ;
	wire _w1465_ ;
	wire _w1466_ ;
	wire _w1467_ ;
	wire _w1468_ ;
	wire _w1469_ ;
	wire _w1470_ ;
	wire _w1471_ ;
	wire _w1472_ ;
	wire _w1473_ ;
	wire _w1474_ ;
	wire _w1475_ ;
	wire _w1476_ ;
	wire _w1477_ ;
	wire _w1478_ ;
	wire _w1479_ ;
	wire _w1480_ ;
	wire _w1481_ ;
	wire _w1482_ ;
	wire _w1483_ ;
	wire _w1484_ ;
	wire _w1485_ ;
	wire _w1486_ ;
	wire _w1487_ ;
	wire _w1488_ ;
	wire _w1489_ ;
	wire _w1490_ ;
	wire _w1491_ ;
	wire _w1492_ ;
	wire _w1493_ ;
	wire _w1494_ ;
	wire _w1495_ ;
	wire _w1496_ ;
	wire _w1497_ ;
	wire _w1498_ ;
	wire _w1499_ ;
	wire _w1500_ ;
	wire _w1501_ ;
	wire _w1502_ ;
	wire _w1503_ ;
	wire _w1504_ ;
	wire _w1505_ ;
	wire _w1506_ ;
	wire _w1507_ ;
	wire _w1508_ ;
	wire _w1509_ ;
	wire _w1510_ ;
	wire _w1511_ ;
	wire _w1512_ ;
	wire _w1513_ ;
	wire _w1514_ ;
	wire _w1515_ ;
	wire _w1516_ ;
	wire _w1517_ ;
	wire _w1518_ ;
	wire _w1519_ ;
	wire _w1520_ ;
	wire _w1521_ ;
	wire _w1522_ ;
	wire _w1523_ ;
	wire _w1524_ ;
	wire _w1525_ ;
	wire _w1526_ ;
	wire _w1527_ ;
	wire _w1528_ ;
	wire _w1529_ ;
	wire _w1530_ ;
	wire _w1531_ ;
	wire _w1532_ ;
	wire _w1533_ ;
	wire _w1534_ ;
	wire _w1535_ ;
	wire _w1536_ ;
	wire _w1537_ ;
	wire _w1538_ ;
	wire _w1539_ ;
	wire _w1540_ ;
	wire _w1541_ ;
	wire _w1542_ ;
	wire _w1543_ ;
	wire _w1544_ ;
	wire _w1545_ ;
	wire _w1546_ ;
	wire _w1547_ ;
	wire _w1548_ ;
	wire _w1549_ ;
	wire _w1550_ ;
	wire _w1551_ ;
	wire _w1552_ ;
	wire _w1553_ ;
	wire _w1554_ ;
	wire _w1555_ ;
	wire _w1556_ ;
	wire _w1557_ ;
	wire _w1558_ ;
	wire _w1559_ ;
	wire _w1560_ ;
	wire _w1561_ ;
	wire _w1562_ ;
	wire _w1563_ ;
	wire _w1564_ ;
	wire _w1565_ ;
	wire _w1566_ ;
	wire _w1567_ ;
	wire _w1568_ ;
	wire _w1569_ ;
	wire _w1570_ ;
	wire _w1571_ ;
	wire _w1572_ ;
	wire _w1573_ ;
	wire _w1574_ ;
	wire _w1575_ ;
	wire _w1576_ ;
	wire _w1577_ ;
	wire _w1578_ ;
	wire _w1579_ ;
	wire _w1580_ ;
	wire _w1581_ ;
	wire _w1582_ ;
	wire _w1583_ ;
	wire _w1584_ ;
	wire _w1585_ ;
	wire _w1586_ ;
	wire _w1587_ ;
	wire _w1588_ ;
	wire _w1589_ ;
	wire _w1590_ ;
	wire _w1591_ ;
	wire _w1592_ ;
	wire _w1593_ ;
	wire _w1594_ ;
	wire _w1595_ ;
	wire _w1596_ ;
	wire _w1597_ ;
	wire _w1598_ ;
	wire _w1599_ ;
	wire _w1600_ ;
	wire _w1601_ ;
	wire _w1602_ ;
	wire _w1603_ ;
	wire _w1604_ ;
	wire _w1605_ ;
	wire _w1606_ ;
	wire _w1607_ ;
	wire _w1608_ ;
	wire _w1609_ ;
	wire _w1610_ ;
	wire _w1611_ ;
	wire _w1612_ ;
	wire _w1613_ ;
	wire _w1614_ ;
	wire _w1615_ ;
	wire _w1616_ ;
	wire _w1617_ ;
	wire _w1618_ ;
	wire _w1619_ ;
	wire _w1620_ ;
	wire _w1621_ ;
	wire _w1622_ ;
	wire _w1623_ ;
	wire _w1624_ ;
	wire _w1625_ ;
	wire _w1626_ ;
	wire _w1627_ ;
	wire _w1628_ ;
	wire _w1629_ ;
	wire _w1630_ ;
	wire _w1631_ ;
	wire _w1632_ ;
	wire _w1633_ ;
	wire _w1634_ ;
	wire _w1635_ ;
	wire _w1636_ ;
	wire _w1637_ ;
	wire _w1638_ ;
	wire _w1639_ ;
	wire _w1640_ ;
	wire _w1641_ ;
	wire _w1642_ ;
	wire _w1643_ ;
	wire _w1644_ ;
	wire _w1645_ ;
	wire _w1646_ ;
	wire _w1647_ ;
	wire _w1648_ ;
	wire _w1649_ ;
	wire _w1650_ ;
	wire _w1651_ ;
	wire _w1652_ ;
	wire _w1653_ ;
	wire _w1654_ ;
	wire _w1655_ ;
	wire _w1656_ ;
	wire _w1657_ ;
	wire _w1658_ ;
	wire _w1659_ ;
	wire _w1660_ ;
	wire _w1661_ ;
	wire _w1662_ ;
	wire _w1663_ ;
	wire _w1664_ ;
	wire _w1665_ ;
	wire _w1666_ ;
	wire _w1667_ ;
	wire _w1668_ ;
	wire _w1669_ ;
	wire _w1670_ ;
	wire _w1671_ ;
	wire _w1672_ ;
	wire _w1673_ ;
	wire _w1674_ ;
	wire _w1675_ ;
	wire _w1676_ ;
	wire _w1677_ ;
	wire _w1678_ ;
	wire _w1679_ ;
	wire _w1680_ ;
	wire _w1681_ ;
	wire _w1682_ ;
	wire _w1683_ ;
	wire _w1684_ ;
	wire _w1685_ ;
	wire _w1686_ ;
	wire _w1687_ ;
	wire _w1688_ ;
	wire _w1689_ ;
	wire _w1690_ ;
	wire _w1691_ ;
	wire _w1692_ ;
	wire _w1693_ ;
	wire _w1694_ ;
	wire _w1695_ ;
	wire _w1696_ ;
	wire _w1697_ ;
	wire _w1698_ ;
	wire _w1699_ ;
	wire _w1700_ ;
	wire _w1701_ ;
	wire _w1702_ ;
	wire _w1703_ ;
	wire _w1704_ ;
	wire _w1705_ ;
	wire _w1706_ ;
	wire _w1707_ ;
	wire _w1708_ ;
	wire _w1709_ ;
	wire _w1710_ ;
	wire _w1711_ ;
	wire _w1712_ ;
	wire _w1713_ ;
	wire _w1714_ ;
	wire _w1715_ ;
	wire _w1716_ ;
	wire _w1717_ ;
	wire _w1718_ ;
	wire _w1719_ ;
	wire _w1720_ ;
	wire _w1721_ ;
	wire _w1722_ ;
	wire _w1723_ ;
	wire _w1724_ ;
	wire _w1725_ ;
	wire _w1726_ ;
	wire _w1727_ ;
	wire _w1728_ ;
	wire _w1729_ ;
	wire _w1730_ ;
	wire _w1731_ ;
	wire _w1732_ ;
	wire _w1733_ ;
	wire _w1734_ ;
	wire _w1735_ ;
	wire _w1736_ ;
	wire _w1737_ ;
	wire _w1738_ ;
	wire _w1739_ ;
	wire _w1740_ ;
	wire _w1741_ ;
	wire _w1742_ ;
	wire _w1743_ ;
	wire _w1744_ ;
	wire _w1745_ ;
	wire _w1746_ ;
	wire _w1747_ ;
	wire _w1748_ ;
	wire _w1749_ ;
	wire _w1750_ ;
	wire _w1751_ ;
	wire _w1752_ ;
	wire _w1753_ ;
	wire _w1754_ ;
	wire _w1755_ ;
	wire _w1756_ ;
	wire _w1757_ ;
	wire _w1758_ ;
	wire _w1759_ ;
	wire _w1760_ ;
	wire _w1761_ ;
	wire _w1762_ ;
	wire _w1763_ ;
	wire _w1764_ ;
	wire _w1765_ ;
	wire _w1766_ ;
	wire _w1767_ ;
	wire _w1768_ ;
	wire _w1769_ ;
	wire _w1770_ ;
	wire _w1771_ ;
	wire _w1772_ ;
	wire _w1773_ ;
	wire _w1774_ ;
	wire _w1775_ ;
	wire _w1776_ ;
	wire _w1777_ ;
	wire _w1778_ ;
	wire _w1779_ ;
	wire _w1780_ ;
	wire _w1781_ ;
	wire _w1782_ ;
	wire _w1783_ ;
	wire _w1784_ ;
	wire _w1785_ ;
	wire _w1786_ ;
	wire _w1787_ ;
	wire _w1788_ ;
	wire _w1789_ ;
	wire _w1790_ ;
	wire _w1791_ ;
	wire _w1792_ ;
	wire _w1793_ ;
	wire _w1794_ ;
	wire _w1795_ ;
	wire _w1796_ ;
	wire _w1797_ ;
	wire _w1798_ ;
	wire _w1799_ ;
	wire _w1800_ ;
	wire _w1801_ ;
	wire _w1802_ ;
	wire _w1803_ ;
	wire _w1804_ ;
	wire _w1805_ ;
	wire _w1806_ ;
	wire _w1807_ ;
	wire _w1808_ ;
	wire _w1809_ ;
	wire _w1810_ ;
	wire _w1811_ ;
	wire _w1812_ ;
	wire _w1813_ ;
	wire _w1814_ ;
	wire _w1815_ ;
	wire _w1816_ ;
	wire _w1817_ ;
	wire _w1818_ ;
	wire _w1819_ ;
	wire _w1820_ ;
	wire _w1821_ ;
	wire _w1822_ ;
	wire _w1823_ ;
	wire _w1824_ ;
	wire _w1825_ ;
	wire _w1826_ ;
	wire _w1827_ ;
	wire _w1828_ ;
	wire _w1829_ ;
	wire _w1830_ ;
	wire _w1831_ ;
	wire _w1832_ ;
	wire _w1833_ ;
	wire _w1834_ ;
	wire _w1835_ ;
	wire _w1836_ ;
	wire _w1837_ ;
	wire _w1838_ ;
	wire _w1839_ ;
	wire _w1840_ ;
	wire _w1841_ ;
	wire _w1842_ ;
	wire _w1843_ ;
	wire _w1844_ ;
	wire _w1845_ ;
	wire _w1846_ ;
	wire _w1847_ ;
	wire _w1848_ ;
	wire _w1849_ ;
	wire _w1850_ ;
	wire _w1851_ ;
	wire _w1852_ ;
	wire _w1853_ ;
	wire _w1854_ ;
	wire _w1855_ ;
	wire _w1856_ ;
	wire _w1857_ ;
	wire _w1858_ ;
	wire _w1859_ ;
	wire _w1860_ ;
	wire _w1861_ ;
	wire _w1862_ ;
	wire _w1863_ ;
	wire _w1864_ ;
	wire _w1865_ ;
	wire _w1866_ ;
	wire _w1867_ ;
	wire _w1868_ ;
	wire _w1869_ ;
	wire _w1870_ ;
	wire _w1871_ ;
	wire _w1872_ ;
	wire _w1873_ ;
	wire _w1874_ ;
	wire _w1875_ ;
	wire _w1876_ ;
	wire _w1877_ ;
	wire _w1878_ ;
	wire _w1879_ ;
	wire _w1880_ ;
	wire _w1881_ ;
	wire _w1882_ ;
	wire _w1883_ ;
	wire _w1884_ ;
	wire _w1885_ ;
	wire _w1886_ ;
	wire _w1887_ ;
	wire _w1888_ ;
	wire _w1889_ ;
	wire _w1890_ ;
	wire _w1891_ ;
	wire _w1892_ ;
	wire _w1893_ ;
	wire _w1894_ ;
	wire _w1895_ ;
	wire _w1896_ ;
	wire _w1897_ ;
	wire _w1898_ ;
	wire _w1899_ ;
	wire _w1900_ ;
	wire _w1901_ ;
	wire _w1902_ ;
	wire _w1903_ ;
	wire _w1904_ ;
	wire _w1905_ ;
	wire _w1906_ ;
	wire _w1907_ ;
	wire _w1908_ ;
	wire _w1909_ ;
	wire _w1910_ ;
	wire _w1911_ ;
	wire _w1912_ ;
	wire _w1913_ ;
	wire _w1914_ ;
	wire _w1915_ ;
	wire _w1916_ ;
	wire _w1917_ ;
	wire _w1918_ ;
	wire _w1919_ ;
	wire _w1920_ ;
	wire _w1921_ ;
	wire _w1922_ ;
	wire _w1923_ ;
	wire _w1924_ ;
	wire _w1925_ ;
	wire _w1926_ ;
	wire _w1927_ ;
	wire _w1928_ ;
	wire _w1929_ ;
	wire _w1930_ ;
	wire _w1931_ ;
	wire _w1932_ ;
	wire _w1933_ ;
	wire _w1934_ ;
	wire _w1935_ ;
	wire _w1936_ ;
	wire _w1937_ ;
	wire _w1938_ ;
	wire _w1939_ ;
	wire _w1940_ ;
	wire _w1941_ ;
	wire _w1942_ ;
	wire _w1943_ ;
	wire _w1944_ ;
	wire _w1945_ ;
	wire _w1946_ ;
	wire _w1947_ ;
	wire _w1948_ ;
	wire _w1949_ ;
	wire _w1950_ ;
	wire _w1951_ ;
	wire _w1952_ ;
	wire _w1953_ ;
	wire _w1954_ ;
	wire _w1955_ ;
	wire _w1956_ ;
	wire _w1957_ ;
	wire _w1958_ ;
	wire _w1959_ ;
	wire _w1960_ ;
	wire _w1961_ ;
	wire _w1962_ ;
	wire _w1963_ ;
	wire _w1964_ ;
	wire _w1965_ ;
	wire _w1966_ ;
	wire _w1967_ ;
	wire _w1968_ ;
	wire _w1969_ ;
	wire _w1970_ ;
	wire _w1971_ ;
	wire _w1972_ ;
	wire _w1973_ ;
	wire _w1974_ ;
	wire _w1975_ ;
	wire _w1976_ ;
	wire _w1977_ ;
	wire _w1978_ ;
	wire _w1979_ ;
	wire _w1980_ ;
	wire _w1981_ ;
	wire _w1982_ ;
	wire _w1983_ ;
	wire _w1984_ ;
	wire _w1985_ ;
	wire _w1986_ ;
	wire _w1987_ ;
	wire _w1988_ ;
	wire _w1989_ ;
	wire _w1990_ ;
	wire _w1991_ ;
	wire _w1992_ ;
	wire _w1993_ ;
	wire _w1994_ ;
	wire _w1995_ ;
	wire _w1996_ ;
	wire _w1997_ ;
	wire _w1998_ ;
	wire _w1999_ ;
	wire _w2000_ ;
	wire _w2001_ ;
	wire _w2002_ ;
	wire _w2003_ ;
	wire _w2004_ ;
	wire _w2005_ ;
	wire _w2006_ ;
	wire _w2007_ ;
	wire _w2008_ ;
	wire _w2009_ ;
	wire _w2010_ ;
	wire _w2011_ ;
	wire _w2012_ ;
	wire _w2013_ ;
	wire _w2014_ ;
	wire _w2015_ ;
	wire _w2016_ ;
	wire _w2017_ ;
	wire _w2018_ ;
	wire _w2019_ ;
	wire _w2020_ ;
	wire _w2021_ ;
	wire _w2022_ ;
	wire _w2023_ ;
	wire _w2024_ ;
	wire _w2025_ ;
	wire _w2026_ ;
	wire _w2027_ ;
	wire _w2028_ ;
	wire _w2029_ ;
	wire _w2030_ ;
	wire _w2031_ ;
	wire _w2032_ ;
	wire _w2033_ ;
	wire _w2034_ ;
	wire _w2035_ ;
	wire _w2036_ ;
	wire _w2037_ ;
	wire _w2038_ ;
	wire _w2039_ ;
	wire _w2040_ ;
	wire _w2041_ ;
	wire _w2042_ ;
	wire _w2043_ ;
	wire _w2044_ ;
	wire _w2045_ ;
	wire _w2046_ ;
	wire _w2047_ ;
	wire _w2048_ ;
	wire _w2049_ ;
	wire _w2050_ ;
	wire _w2051_ ;
	wire _w2052_ ;
	wire _w2053_ ;
	wire _w2054_ ;
	wire _w2055_ ;
	wire _w2056_ ;
	wire _w2057_ ;
	wire _w2058_ ;
	wire _w2059_ ;
	wire _w2060_ ;
	wire _w2061_ ;
	wire _w2062_ ;
	wire _w2063_ ;
	wire _w2064_ ;
	wire _w2065_ ;
	wire _w2066_ ;
	wire _w2067_ ;
	wire _w2068_ ;
	wire _w2069_ ;
	wire _w2070_ ;
	wire _w2071_ ;
	wire _w2072_ ;
	wire _w2073_ ;
	wire _w2074_ ;
	wire _w2075_ ;
	wire _w2076_ ;
	wire _w2077_ ;
	wire _w2078_ ;
	wire _w2079_ ;
	wire _w2080_ ;
	wire _w2081_ ;
	wire _w2082_ ;
	wire _w2083_ ;
	wire _w2084_ ;
	wire _w2085_ ;
	wire _w2086_ ;
	wire _w2087_ ;
	wire _w2088_ ;
	wire _w2089_ ;
	wire _w2090_ ;
	wire _w2091_ ;
	wire _w2092_ ;
	wire _w2093_ ;
	wire _w2094_ ;
	wire _w2095_ ;
	wire _w2096_ ;
	wire _w2097_ ;
	wire _w2098_ ;
	wire _w2099_ ;
	wire _w2100_ ;
	wire _w2101_ ;
	wire _w2102_ ;
	wire _w2103_ ;
	wire _w2104_ ;
	wire _w2105_ ;
	wire _w2106_ ;
	wire _w2107_ ;
	wire _w2108_ ;
	wire _w2109_ ;
	wire _w2110_ ;
	wire _w2111_ ;
	wire _w2112_ ;
	wire _w2113_ ;
	wire _w2114_ ;
	wire _w2115_ ;
	wire _w2116_ ;
	wire _w2117_ ;
	wire _w2118_ ;
	wire _w2119_ ;
	wire _w2120_ ;
	wire _w2121_ ;
	wire _w2122_ ;
	wire _w2123_ ;
	wire _w2124_ ;
	wire _w2125_ ;
	wire _w2126_ ;
	wire _w2127_ ;
	wire _w2128_ ;
	wire _w2129_ ;
	wire _w2130_ ;
	wire _w2131_ ;
	wire _w2132_ ;
	wire _w2133_ ;
	wire _w2134_ ;
	wire _w2135_ ;
	wire _w2136_ ;
	wire _w2137_ ;
	wire _w2138_ ;
	wire _w2139_ ;
	wire _w2140_ ;
	wire _w2141_ ;
	wire _w2142_ ;
	wire _w2143_ ;
	wire _w2144_ ;
	wire _w2145_ ;
	wire _w2146_ ;
	wire _w2147_ ;
	wire _w2148_ ;
	wire _w2149_ ;
	wire _w2150_ ;
	wire _w2151_ ;
	wire _w2152_ ;
	wire _w2153_ ;
	wire _w2154_ ;
	wire _w2155_ ;
	wire _w2156_ ;
	wire _w2157_ ;
	wire _w2158_ ;
	wire _w2159_ ;
	wire _w2160_ ;
	wire _w2161_ ;
	wire _w2162_ ;
	wire _w2163_ ;
	wire _w2164_ ;
	wire _w2165_ ;
	wire _w2166_ ;
	wire _w2167_ ;
	wire _w2168_ ;
	wire _w2169_ ;
	wire _w2170_ ;
	wire _w2171_ ;
	wire _w2172_ ;
	wire _w2173_ ;
	wire _w2174_ ;
	wire _w2175_ ;
	wire _w2176_ ;
	wire _w2177_ ;
	wire _w2178_ ;
	wire _w2179_ ;
	wire _w2180_ ;
	wire _w2181_ ;
	wire _w2182_ ;
	wire _w2183_ ;
	wire _w2184_ ;
	wire _w2185_ ;
	wire _w2186_ ;
	wire _w2187_ ;
	wire _w2188_ ;
	wire _w2189_ ;
	wire _w2190_ ;
	wire _w2191_ ;
	wire _w2192_ ;
	wire _w2193_ ;
	wire _w2194_ ;
	wire _w2195_ ;
	wire _w2196_ ;
	wire _w2197_ ;
	wire _w2198_ ;
	wire _w2199_ ;
	wire _w2200_ ;
	wire _w2201_ ;
	wire _w2202_ ;
	wire _w2203_ ;
	wire _w2204_ ;
	wire _w2205_ ;
	wire _w2206_ ;
	wire _w2207_ ;
	wire _w2208_ ;
	wire _w2209_ ;
	wire _w2210_ ;
	wire _w2211_ ;
	wire _w2212_ ;
	wire _w2213_ ;
	wire _w2214_ ;
	wire _w2215_ ;
	wire _w2216_ ;
	wire _w2217_ ;
	wire _w2218_ ;
	wire _w2219_ ;
	wire _w2220_ ;
	wire _w2221_ ;
	wire _w2222_ ;
	wire _w2223_ ;
	wire _w2224_ ;
	wire _w2225_ ;
	wire _w2226_ ;
	wire _w2227_ ;
	wire _w2228_ ;
	wire _w2229_ ;
	wire _w2230_ ;
	wire _w2231_ ;
	wire _w2232_ ;
	wire _w2233_ ;
	wire _w2234_ ;
	wire _w2235_ ;
	wire _w2236_ ;
	wire _w2237_ ;
	wire _w2238_ ;
	wire _w2239_ ;
	wire _w2240_ ;
	wire _w2241_ ;
	wire _w2242_ ;
	wire _w2243_ ;
	wire _w2244_ ;
	wire _w2245_ ;
	wire _w2246_ ;
	wire _w2247_ ;
	wire _w2248_ ;
	wire _w2249_ ;
	wire _w2250_ ;
	wire _w2251_ ;
	wire _w2252_ ;
	wire _w2253_ ;
	wire _w2254_ ;
	wire _w2255_ ;
	wire _w2256_ ;
	wire _w2257_ ;
	wire _w2258_ ;
	wire _w2259_ ;
	wire _w2260_ ;
	wire _w2261_ ;
	wire _w2262_ ;
	wire _w2263_ ;
	wire _w2264_ ;
	wire _w2265_ ;
	wire _w2266_ ;
	wire _w2267_ ;
	wire _w2268_ ;
	wire _w2269_ ;
	wire _w2270_ ;
	wire _w2271_ ;
	wire _w2272_ ;
	wire _w2273_ ;
	wire _w2274_ ;
	wire _w2275_ ;
	wire _w2276_ ;
	wire _w2277_ ;
	wire _w2278_ ;
	wire _w2279_ ;
	wire _w2280_ ;
	wire _w2281_ ;
	wire _w2282_ ;
	wire _w2283_ ;
	wire _w2284_ ;
	wire _w2285_ ;
	wire _w2286_ ;
	wire _w2287_ ;
	wire _w2288_ ;
	wire _w2289_ ;
	wire _w2290_ ;
	wire _w2291_ ;
	wire _w2292_ ;
	wire _w2293_ ;
	wire _w2294_ ;
	wire _w2295_ ;
	wire _w2296_ ;
	wire _w2297_ ;
	wire _w2298_ ;
	wire _w2299_ ;
	wire _w2300_ ;
	wire _w2301_ ;
	wire _w2302_ ;
	wire _w2303_ ;
	wire _w2304_ ;
	wire _w2305_ ;
	wire _w2306_ ;
	wire _w2307_ ;
	wire _w2308_ ;
	wire _w2309_ ;
	wire _w2310_ ;
	wire _w2311_ ;
	wire _w2312_ ;
	wire _w2313_ ;
	wire _w2314_ ;
	wire _w2315_ ;
	wire _w2316_ ;
	wire _w2317_ ;
	wire _w2318_ ;
	wire _w2319_ ;
	wire _w2320_ ;
	wire _w2321_ ;
	wire _w2322_ ;
	wire _w2323_ ;
	wire _w2324_ ;
	wire _w2325_ ;
	wire _w2326_ ;
	wire _w2327_ ;
	wire _w2328_ ;
	wire _w2329_ ;
	wire _w2330_ ;
	wire _w2331_ ;
	wire _w2332_ ;
	wire _w2333_ ;
	wire _w2334_ ;
	wire _w2335_ ;
	wire _w2336_ ;
	wire _w2337_ ;
	wire _w2338_ ;
	wire _w2339_ ;
	wire _w2340_ ;
	wire _w2341_ ;
	wire _w2342_ ;
	wire _w2343_ ;
	wire _w2344_ ;
	wire _w2345_ ;
	wire _w2346_ ;
	wire _w2347_ ;
	wire _w2348_ ;
	wire _w2349_ ;
	wire _w2350_ ;
	wire _w2351_ ;
	wire _w2352_ ;
	wire _w2353_ ;
	wire _w2354_ ;
	wire _w2355_ ;
	wire _w2356_ ;
	wire _w2357_ ;
	wire _w2358_ ;
	wire _w2359_ ;
	wire _w2360_ ;
	wire _w2361_ ;
	wire _w2362_ ;
	wire _w2363_ ;
	wire _w2364_ ;
	wire _w2365_ ;
	wire _w2366_ ;
	wire _w2367_ ;
	wire _w2368_ ;
	wire _w2369_ ;
	wire _w2370_ ;
	wire _w2371_ ;
	wire _w2372_ ;
	wire _w2373_ ;
	wire _w2374_ ;
	wire _w2375_ ;
	wire _w2376_ ;
	wire _w2377_ ;
	wire _w2378_ ;
	wire _w2379_ ;
	wire _w2380_ ;
	wire _w2381_ ;
	wire _w2382_ ;
	wire _w2383_ ;
	wire _w2384_ ;
	wire _w2385_ ;
	wire _w2386_ ;
	wire _w2387_ ;
	wire _w2388_ ;
	wire _w2389_ ;
	wire _w2390_ ;
	wire _w2391_ ;
	wire _w2392_ ;
	wire _w2393_ ;
	wire _w2394_ ;
	wire _w2395_ ;
	wire _w2396_ ;
	wire _w2397_ ;
	wire _w2398_ ;
	wire _w2399_ ;
	wire _w2400_ ;
	wire _w2401_ ;
	wire _w2402_ ;
	wire _w2403_ ;
	wire _w2404_ ;
	wire _w2405_ ;
	wire _w2406_ ;
	wire _w2407_ ;
	wire _w2408_ ;
	wire _w2409_ ;
	wire _w2410_ ;
	wire _w2411_ ;
	wire _w2412_ ;
	wire _w2413_ ;
	wire _w2414_ ;
	wire _w2415_ ;
	wire _w2416_ ;
	wire _w2417_ ;
	wire _w2418_ ;
	wire _w2419_ ;
	wire _w2420_ ;
	wire _w2421_ ;
	wire _w2422_ ;
	wire _w2423_ ;
	wire _w2424_ ;
	wire _w2425_ ;
	wire _w2426_ ;
	wire _w2427_ ;
	wire _w2428_ ;
	wire _w2429_ ;
	wire _w2430_ ;
	wire _w2431_ ;
	wire _w2432_ ;
	wire _w2433_ ;
	wire _w2434_ ;
	wire _w2435_ ;
	wire _w2436_ ;
	wire _w2437_ ;
	wire _w2438_ ;
	wire _w2439_ ;
	wire _w2440_ ;
	wire _w2441_ ;
	wire _w2442_ ;
	wire _w2443_ ;
	wire _w2444_ ;
	wire _w2445_ ;
	wire _w2446_ ;
	wire _w2447_ ;
	wire _w2448_ ;
	wire _w2449_ ;
	wire _w2450_ ;
	wire _w2451_ ;
	wire _w2452_ ;
	wire _w2453_ ;
	wire _w2454_ ;
	wire _w2455_ ;
	wire _w2456_ ;
	wire _w2457_ ;
	wire _w2458_ ;
	wire _w2459_ ;
	wire _w2460_ ;
	wire _w2461_ ;
	wire _w2462_ ;
	wire _w2463_ ;
	wire _w2464_ ;
	wire _w2465_ ;
	wire _w2466_ ;
	wire _w2467_ ;
	wire _w2468_ ;
	wire _w2469_ ;
	wire _w2470_ ;
	wire _w2471_ ;
	wire _w2472_ ;
	wire _w2473_ ;
	wire _w2474_ ;
	wire _w2475_ ;
	wire _w2476_ ;
	wire _w2477_ ;
	wire _w2478_ ;
	wire _w2479_ ;
	wire _w2480_ ;
	wire _w2481_ ;
	wire _w2482_ ;
	wire _w2483_ ;
	wire _w2484_ ;
	wire _w2485_ ;
	wire _w2486_ ;
	wire _w2487_ ;
	wire _w2488_ ;
	wire _w2489_ ;
	wire _w2490_ ;
	wire _w2491_ ;
	wire _w2492_ ;
	LUT2 #(
		.INIT('h1)
	) name0 (
		\shift[2] ,
		\shift[3] ,
		_w136_
	);
	LUT2 #(
		.INIT('h8)
	) name1 (
		\a[77] ,
		\shift[0] ,
		_w137_
	);
	LUT2 #(
		.INIT('h2)
	) name2 (
		\a[78] ,
		\shift[0] ,
		_w138_
	);
	LUT2 #(
		.INIT('h1)
	) name3 (
		_w137_,
		_w138_,
		_w139_
	);
	LUT2 #(
		.INIT('h2)
	) name4 (
		\shift[1] ,
		_w139_,
		_w140_
	);
	LUT2 #(
		.INIT('h2)
	) name5 (
		\a[80] ,
		\shift[0] ,
		_w141_
	);
	LUT2 #(
		.INIT('h8)
	) name6 (
		\a[79] ,
		\shift[0] ,
		_w142_
	);
	LUT2 #(
		.INIT('h1)
	) name7 (
		_w141_,
		_w142_,
		_w143_
	);
	LUT2 #(
		.INIT('h1)
	) name8 (
		\shift[1] ,
		_w143_,
		_w144_
	);
	LUT2 #(
		.INIT('h1)
	) name9 (
		_w140_,
		_w144_,
		_w145_
	);
	LUT2 #(
		.INIT('h2)
	) name10 (
		_w136_,
		_w145_,
		_w146_
	);
	LUT2 #(
		.INIT('h2)
	) name11 (
		\shift[2] ,
		\shift[3] ,
		_w147_
	);
	LUT2 #(
		.INIT('h8)
	) name12 (
		\a[73] ,
		\shift[0] ,
		_w148_
	);
	LUT2 #(
		.INIT('h2)
	) name13 (
		\a[74] ,
		\shift[0] ,
		_w149_
	);
	LUT2 #(
		.INIT('h1)
	) name14 (
		_w148_,
		_w149_,
		_w150_
	);
	LUT2 #(
		.INIT('h2)
	) name15 (
		\shift[1] ,
		_w150_,
		_w151_
	);
	LUT2 #(
		.INIT('h2)
	) name16 (
		\a[76] ,
		\shift[0] ,
		_w152_
	);
	LUT2 #(
		.INIT('h8)
	) name17 (
		\a[75] ,
		\shift[0] ,
		_w153_
	);
	LUT2 #(
		.INIT('h1)
	) name18 (
		_w152_,
		_w153_,
		_w154_
	);
	LUT2 #(
		.INIT('h1)
	) name19 (
		\shift[1] ,
		_w154_,
		_w155_
	);
	LUT2 #(
		.INIT('h1)
	) name20 (
		_w151_,
		_w155_,
		_w156_
	);
	LUT2 #(
		.INIT('h2)
	) name21 (
		_w147_,
		_w156_,
		_w157_
	);
	LUT2 #(
		.INIT('h8)
	) name22 (
		\shift[2] ,
		\shift[3] ,
		_w158_
	);
	LUT2 #(
		.INIT('h8)
	) name23 (
		\a[65] ,
		\shift[0] ,
		_w159_
	);
	LUT2 #(
		.INIT('h2)
	) name24 (
		\a[66] ,
		\shift[0] ,
		_w160_
	);
	LUT2 #(
		.INIT('h1)
	) name25 (
		_w159_,
		_w160_,
		_w161_
	);
	LUT2 #(
		.INIT('h2)
	) name26 (
		\shift[1] ,
		_w161_,
		_w162_
	);
	LUT2 #(
		.INIT('h2)
	) name27 (
		\a[68] ,
		\shift[0] ,
		_w163_
	);
	LUT2 #(
		.INIT('h8)
	) name28 (
		\a[67] ,
		\shift[0] ,
		_w164_
	);
	LUT2 #(
		.INIT('h1)
	) name29 (
		_w163_,
		_w164_,
		_w165_
	);
	LUT2 #(
		.INIT('h1)
	) name30 (
		\shift[1] ,
		_w165_,
		_w166_
	);
	LUT2 #(
		.INIT('h1)
	) name31 (
		_w162_,
		_w166_,
		_w167_
	);
	LUT2 #(
		.INIT('h2)
	) name32 (
		_w158_,
		_w167_,
		_w168_
	);
	LUT2 #(
		.INIT('h4)
	) name33 (
		\shift[2] ,
		\shift[3] ,
		_w169_
	);
	LUT2 #(
		.INIT('h8)
	) name34 (
		\a[69] ,
		\shift[0] ,
		_w170_
	);
	LUT2 #(
		.INIT('h2)
	) name35 (
		\a[70] ,
		\shift[0] ,
		_w171_
	);
	LUT2 #(
		.INIT('h1)
	) name36 (
		_w170_,
		_w171_,
		_w172_
	);
	LUT2 #(
		.INIT('h2)
	) name37 (
		\shift[1] ,
		_w172_,
		_w173_
	);
	LUT2 #(
		.INIT('h2)
	) name38 (
		\a[72] ,
		\shift[0] ,
		_w174_
	);
	LUT2 #(
		.INIT('h8)
	) name39 (
		\a[71] ,
		\shift[0] ,
		_w175_
	);
	LUT2 #(
		.INIT('h1)
	) name40 (
		_w174_,
		_w175_,
		_w176_
	);
	LUT2 #(
		.INIT('h1)
	) name41 (
		\shift[1] ,
		_w176_,
		_w177_
	);
	LUT2 #(
		.INIT('h1)
	) name42 (
		_w173_,
		_w177_,
		_w178_
	);
	LUT2 #(
		.INIT('h2)
	) name43 (
		_w169_,
		_w178_,
		_w179_
	);
	LUT2 #(
		.INIT('h1)
	) name44 (
		_w146_,
		_w157_,
		_w180_
	);
	LUT2 #(
		.INIT('h1)
	) name45 (
		_w168_,
		_w179_,
		_w181_
	);
	LUT2 #(
		.INIT('h8)
	) name46 (
		_w180_,
		_w181_,
		_w182_
	);
	LUT2 #(
		.INIT('h8)
	) name47 (
		\shift[4] ,
		\shift[5] ,
		_w183_
	);
	LUT2 #(
		.INIT('h4)
	) name48 (
		_w182_,
		_w183_,
		_w184_
	);
	LUT2 #(
		.INIT('h8)
	) name49 (
		\a[93] ,
		\shift[0] ,
		_w185_
	);
	LUT2 #(
		.INIT('h2)
	) name50 (
		\a[94] ,
		\shift[0] ,
		_w186_
	);
	LUT2 #(
		.INIT('h1)
	) name51 (
		_w185_,
		_w186_,
		_w187_
	);
	LUT2 #(
		.INIT('h2)
	) name52 (
		\shift[1] ,
		_w187_,
		_w188_
	);
	LUT2 #(
		.INIT('h2)
	) name53 (
		\a[96] ,
		\shift[0] ,
		_w189_
	);
	LUT2 #(
		.INIT('h8)
	) name54 (
		\a[95] ,
		\shift[0] ,
		_w190_
	);
	LUT2 #(
		.INIT('h1)
	) name55 (
		_w189_,
		_w190_,
		_w191_
	);
	LUT2 #(
		.INIT('h1)
	) name56 (
		\shift[1] ,
		_w191_,
		_w192_
	);
	LUT2 #(
		.INIT('h1)
	) name57 (
		_w188_,
		_w192_,
		_w193_
	);
	LUT2 #(
		.INIT('h2)
	) name58 (
		_w136_,
		_w193_,
		_w194_
	);
	LUT2 #(
		.INIT('h8)
	) name59 (
		\a[89] ,
		\shift[0] ,
		_w195_
	);
	LUT2 #(
		.INIT('h2)
	) name60 (
		\a[90] ,
		\shift[0] ,
		_w196_
	);
	LUT2 #(
		.INIT('h1)
	) name61 (
		_w195_,
		_w196_,
		_w197_
	);
	LUT2 #(
		.INIT('h2)
	) name62 (
		\shift[1] ,
		_w197_,
		_w198_
	);
	LUT2 #(
		.INIT('h2)
	) name63 (
		\a[92] ,
		\shift[0] ,
		_w199_
	);
	LUT2 #(
		.INIT('h8)
	) name64 (
		\a[91] ,
		\shift[0] ,
		_w200_
	);
	LUT2 #(
		.INIT('h1)
	) name65 (
		_w199_,
		_w200_,
		_w201_
	);
	LUT2 #(
		.INIT('h1)
	) name66 (
		\shift[1] ,
		_w201_,
		_w202_
	);
	LUT2 #(
		.INIT('h1)
	) name67 (
		_w198_,
		_w202_,
		_w203_
	);
	LUT2 #(
		.INIT('h2)
	) name68 (
		_w147_,
		_w203_,
		_w204_
	);
	LUT2 #(
		.INIT('h8)
	) name69 (
		\a[81] ,
		\shift[0] ,
		_w205_
	);
	LUT2 #(
		.INIT('h2)
	) name70 (
		\a[82] ,
		\shift[0] ,
		_w206_
	);
	LUT2 #(
		.INIT('h1)
	) name71 (
		_w205_,
		_w206_,
		_w207_
	);
	LUT2 #(
		.INIT('h2)
	) name72 (
		\shift[1] ,
		_w207_,
		_w208_
	);
	LUT2 #(
		.INIT('h2)
	) name73 (
		\a[84] ,
		\shift[0] ,
		_w209_
	);
	LUT2 #(
		.INIT('h8)
	) name74 (
		\a[83] ,
		\shift[0] ,
		_w210_
	);
	LUT2 #(
		.INIT('h1)
	) name75 (
		_w209_,
		_w210_,
		_w211_
	);
	LUT2 #(
		.INIT('h1)
	) name76 (
		\shift[1] ,
		_w211_,
		_w212_
	);
	LUT2 #(
		.INIT('h1)
	) name77 (
		_w208_,
		_w212_,
		_w213_
	);
	LUT2 #(
		.INIT('h2)
	) name78 (
		_w158_,
		_w213_,
		_w214_
	);
	LUT2 #(
		.INIT('h8)
	) name79 (
		\a[85] ,
		\shift[0] ,
		_w215_
	);
	LUT2 #(
		.INIT('h2)
	) name80 (
		\a[86] ,
		\shift[0] ,
		_w216_
	);
	LUT2 #(
		.INIT('h1)
	) name81 (
		_w215_,
		_w216_,
		_w217_
	);
	LUT2 #(
		.INIT('h2)
	) name82 (
		\shift[1] ,
		_w217_,
		_w218_
	);
	LUT2 #(
		.INIT('h2)
	) name83 (
		\a[88] ,
		\shift[0] ,
		_w219_
	);
	LUT2 #(
		.INIT('h8)
	) name84 (
		\a[87] ,
		\shift[0] ,
		_w220_
	);
	LUT2 #(
		.INIT('h1)
	) name85 (
		_w219_,
		_w220_,
		_w221_
	);
	LUT2 #(
		.INIT('h1)
	) name86 (
		\shift[1] ,
		_w221_,
		_w222_
	);
	LUT2 #(
		.INIT('h1)
	) name87 (
		_w218_,
		_w222_,
		_w223_
	);
	LUT2 #(
		.INIT('h2)
	) name88 (
		_w169_,
		_w223_,
		_w224_
	);
	LUT2 #(
		.INIT('h1)
	) name89 (
		_w194_,
		_w204_,
		_w225_
	);
	LUT2 #(
		.INIT('h1)
	) name90 (
		_w214_,
		_w224_,
		_w226_
	);
	LUT2 #(
		.INIT('h8)
	) name91 (
		_w225_,
		_w226_,
		_w227_
	);
	LUT2 #(
		.INIT('h4)
	) name92 (
		\shift[4] ,
		\shift[5] ,
		_w228_
	);
	LUT2 #(
		.INIT('h4)
	) name93 (
		_w227_,
		_w228_,
		_w229_
	);
	LUT2 #(
		.INIT('h8)
	) name94 (
		\a[125] ,
		\shift[0] ,
		_w230_
	);
	LUT2 #(
		.INIT('h2)
	) name95 (
		\a[126] ,
		\shift[0] ,
		_w231_
	);
	LUT2 #(
		.INIT('h1)
	) name96 (
		_w230_,
		_w231_,
		_w232_
	);
	LUT2 #(
		.INIT('h2)
	) name97 (
		\shift[1] ,
		_w232_,
		_w233_
	);
	LUT2 #(
		.INIT('h2)
	) name98 (
		\a[0] ,
		\shift[0] ,
		_w234_
	);
	LUT2 #(
		.INIT('h8)
	) name99 (
		\a[127] ,
		\shift[0] ,
		_w235_
	);
	LUT2 #(
		.INIT('h1)
	) name100 (
		_w234_,
		_w235_,
		_w236_
	);
	LUT2 #(
		.INIT('h1)
	) name101 (
		\shift[1] ,
		_w236_,
		_w237_
	);
	LUT2 #(
		.INIT('h1)
	) name102 (
		_w233_,
		_w237_,
		_w238_
	);
	LUT2 #(
		.INIT('h2)
	) name103 (
		_w136_,
		_w238_,
		_w239_
	);
	LUT2 #(
		.INIT('h8)
	) name104 (
		\a[121] ,
		\shift[0] ,
		_w240_
	);
	LUT2 #(
		.INIT('h2)
	) name105 (
		\a[122] ,
		\shift[0] ,
		_w241_
	);
	LUT2 #(
		.INIT('h1)
	) name106 (
		_w240_,
		_w241_,
		_w242_
	);
	LUT2 #(
		.INIT('h2)
	) name107 (
		\shift[1] ,
		_w242_,
		_w243_
	);
	LUT2 #(
		.INIT('h2)
	) name108 (
		\a[124] ,
		\shift[0] ,
		_w244_
	);
	LUT2 #(
		.INIT('h8)
	) name109 (
		\a[123] ,
		\shift[0] ,
		_w245_
	);
	LUT2 #(
		.INIT('h1)
	) name110 (
		_w244_,
		_w245_,
		_w246_
	);
	LUT2 #(
		.INIT('h1)
	) name111 (
		\shift[1] ,
		_w246_,
		_w247_
	);
	LUT2 #(
		.INIT('h1)
	) name112 (
		_w243_,
		_w247_,
		_w248_
	);
	LUT2 #(
		.INIT('h2)
	) name113 (
		_w147_,
		_w248_,
		_w249_
	);
	LUT2 #(
		.INIT('h8)
	) name114 (
		\a[113] ,
		\shift[0] ,
		_w250_
	);
	LUT2 #(
		.INIT('h2)
	) name115 (
		\a[114] ,
		\shift[0] ,
		_w251_
	);
	LUT2 #(
		.INIT('h1)
	) name116 (
		_w250_,
		_w251_,
		_w252_
	);
	LUT2 #(
		.INIT('h2)
	) name117 (
		\shift[1] ,
		_w252_,
		_w253_
	);
	LUT2 #(
		.INIT('h2)
	) name118 (
		\a[116] ,
		\shift[0] ,
		_w254_
	);
	LUT2 #(
		.INIT('h8)
	) name119 (
		\a[115] ,
		\shift[0] ,
		_w255_
	);
	LUT2 #(
		.INIT('h1)
	) name120 (
		_w254_,
		_w255_,
		_w256_
	);
	LUT2 #(
		.INIT('h1)
	) name121 (
		\shift[1] ,
		_w256_,
		_w257_
	);
	LUT2 #(
		.INIT('h1)
	) name122 (
		_w253_,
		_w257_,
		_w258_
	);
	LUT2 #(
		.INIT('h2)
	) name123 (
		_w158_,
		_w258_,
		_w259_
	);
	LUT2 #(
		.INIT('h8)
	) name124 (
		\a[117] ,
		\shift[0] ,
		_w260_
	);
	LUT2 #(
		.INIT('h2)
	) name125 (
		\a[118] ,
		\shift[0] ,
		_w261_
	);
	LUT2 #(
		.INIT('h1)
	) name126 (
		_w260_,
		_w261_,
		_w262_
	);
	LUT2 #(
		.INIT('h2)
	) name127 (
		\shift[1] ,
		_w262_,
		_w263_
	);
	LUT2 #(
		.INIT('h2)
	) name128 (
		\a[120] ,
		\shift[0] ,
		_w264_
	);
	LUT2 #(
		.INIT('h8)
	) name129 (
		\a[119] ,
		\shift[0] ,
		_w265_
	);
	LUT2 #(
		.INIT('h1)
	) name130 (
		_w264_,
		_w265_,
		_w266_
	);
	LUT2 #(
		.INIT('h1)
	) name131 (
		\shift[1] ,
		_w266_,
		_w267_
	);
	LUT2 #(
		.INIT('h1)
	) name132 (
		_w263_,
		_w267_,
		_w268_
	);
	LUT2 #(
		.INIT('h2)
	) name133 (
		_w169_,
		_w268_,
		_w269_
	);
	LUT2 #(
		.INIT('h1)
	) name134 (
		_w239_,
		_w249_,
		_w270_
	);
	LUT2 #(
		.INIT('h1)
	) name135 (
		_w259_,
		_w269_,
		_w271_
	);
	LUT2 #(
		.INIT('h8)
	) name136 (
		_w270_,
		_w271_,
		_w272_
	);
	LUT2 #(
		.INIT('h1)
	) name137 (
		\shift[4] ,
		\shift[5] ,
		_w273_
	);
	LUT2 #(
		.INIT('h4)
	) name138 (
		_w272_,
		_w273_,
		_w274_
	);
	LUT2 #(
		.INIT('h8)
	) name139 (
		\a[109] ,
		\shift[0] ,
		_w275_
	);
	LUT2 #(
		.INIT('h2)
	) name140 (
		\a[110] ,
		\shift[0] ,
		_w276_
	);
	LUT2 #(
		.INIT('h1)
	) name141 (
		_w275_,
		_w276_,
		_w277_
	);
	LUT2 #(
		.INIT('h2)
	) name142 (
		\shift[1] ,
		_w277_,
		_w278_
	);
	LUT2 #(
		.INIT('h2)
	) name143 (
		\a[112] ,
		\shift[0] ,
		_w279_
	);
	LUT2 #(
		.INIT('h8)
	) name144 (
		\a[111] ,
		\shift[0] ,
		_w280_
	);
	LUT2 #(
		.INIT('h1)
	) name145 (
		_w279_,
		_w280_,
		_w281_
	);
	LUT2 #(
		.INIT('h1)
	) name146 (
		\shift[1] ,
		_w281_,
		_w282_
	);
	LUT2 #(
		.INIT('h1)
	) name147 (
		_w278_,
		_w282_,
		_w283_
	);
	LUT2 #(
		.INIT('h2)
	) name148 (
		_w136_,
		_w283_,
		_w284_
	);
	LUT2 #(
		.INIT('h8)
	) name149 (
		\a[105] ,
		\shift[0] ,
		_w285_
	);
	LUT2 #(
		.INIT('h2)
	) name150 (
		\a[106] ,
		\shift[0] ,
		_w286_
	);
	LUT2 #(
		.INIT('h1)
	) name151 (
		_w285_,
		_w286_,
		_w287_
	);
	LUT2 #(
		.INIT('h2)
	) name152 (
		\shift[1] ,
		_w287_,
		_w288_
	);
	LUT2 #(
		.INIT('h2)
	) name153 (
		\a[108] ,
		\shift[0] ,
		_w289_
	);
	LUT2 #(
		.INIT('h8)
	) name154 (
		\a[107] ,
		\shift[0] ,
		_w290_
	);
	LUT2 #(
		.INIT('h1)
	) name155 (
		_w289_,
		_w290_,
		_w291_
	);
	LUT2 #(
		.INIT('h1)
	) name156 (
		\shift[1] ,
		_w291_,
		_w292_
	);
	LUT2 #(
		.INIT('h1)
	) name157 (
		_w288_,
		_w292_,
		_w293_
	);
	LUT2 #(
		.INIT('h2)
	) name158 (
		_w147_,
		_w293_,
		_w294_
	);
	LUT2 #(
		.INIT('h8)
	) name159 (
		\a[97] ,
		\shift[0] ,
		_w295_
	);
	LUT2 #(
		.INIT('h2)
	) name160 (
		\a[98] ,
		\shift[0] ,
		_w296_
	);
	LUT2 #(
		.INIT('h1)
	) name161 (
		_w295_,
		_w296_,
		_w297_
	);
	LUT2 #(
		.INIT('h2)
	) name162 (
		\shift[1] ,
		_w297_,
		_w298_
	);
	LUT2 #(
		.INIT('h2)
	) name163 (
		\a[100] ,
		\shift[0] ,
		_w299_
	);
	LUT2 #(
		.INIT('h8)
	) name164 (
		\a[99] ,
		\shift[0] ,
		_w300_
	);
	LUT2 #(
		.INIT('h1)
	) name165 (
		_w299_,
		_w300_,
		_w301_
	);
	LUT2 #(
		.INIT('h1)
	) name166 (
		\shift[1] ,
		_w301_,
		_w302_
	);
	LUT2 #(
		.INIT('h1)
	) name167 (
		_w298_,
		_w302_,
		_w303_
	);
	LUT2 #(
		.INIT('h2)
	) name168 (
		_w158_,
		_w303_,
		_w304_
	);
	LUT2 #(
		.INIT('h8)
	) name169 (
		\a[101] ,
		\shift[0] ,
		_w305_
	);
	LUT2 #(
		.INIT('h2)
	) name170 (
		\a[102] ,
		\shift[0] ,
		_w306_
	);
	LUT2 #(
		.INIT('h1)
	) name171 (
		_w305_,
		_w306_,
		_w307_
	);
	LUT2 #(
		.INIT('h2)
	) name172 (
		\shift[1] ,
		_w307_,
		_w308_
	);
	LUT2 #(
		.INIT('h2)
	) name173 (
		\a[104] ,
		\shift[0] ,
		_w309_
	);
	LUT2 #(
		.INIT('h8)
	) name174 (
		\a[103] ,
		\shift[0] ,
		_w310_
	);
	LUT2 #(
		.INIT('h1)
	) name175 (
		_w309_,
		_w310_,
		_w311_
	);
	LUT2 #(
		.INIT('h1)
	) name176 (
		\shift[1] ,
		_w311_,
		_w312_
	);
	LUT2 #(
		.INIT('h1)
	) name177 (
		_w308_,
		_w312_,
		_w313_
	);
	LUT2 #(
		.INIT('h2)
	) name178 (
		_w169_,
		_w313_,
		_w314_
	);
	LUT2 #(
		.INIT('h1)
	) name179 (
		_w284_,
		_w294_,
		_w315_
	);
	LUT2 #(
		.INIT('h1)
	) name180 (
		_w304_,
		_w314_,
		_w316_
	);
	LUT2 #(
		.INIT('h8)
	) name181 (
		_w315_,
		_w316_,
		_w317_
	);
	LUT2 #(
		.INIT('h2)
	) name182 (
		\shift[4] ,
		\shift[5] ,
		_w318_
	);
	LUT2 #(
		.INIT('h4)
	) name183 (
		_w317_,
		_w318_,
		_w319_
	);
	LUT2 #(
		.INIT('h1)
	) name184 (
		_w184_,
		_w229_,
		_w320_
	);
	LUT2 #(
		.INIT('h1)
	) name185 (
		_w274_,
		_w319_,
		_w321_
	);
	LUT2 #(
		.INIT('h8)
	) name186 (
		_w320_,
		_w321_,
		_w322_
	);
	LUT2 #(
		.INIT('h1)
	) name187 (
		\shift[6] ,
		_w322_,
		_w323_
	);
	LUT2 #(
		.INIT('h8)
	) name188 (
		\a[13] ,
		\shift[0] ,
		_w324_
	);
	LUT2 #(
		.INIT('h2)
	) name189 (
		\a[14] ,
		\shift[0] ,
		_w325_
	);
	LUT2 #(
		.INIT('h1)
	) name190 (
		_w324_,
		_w325_,
		_w326_
	);
	LUT2 #(
		.INIT('h2)
	) name191 (
		\shift[1] ,
		_w326_,
		_w327_
	);
	LUT2 #(
		.INIT('h2)
	) name192 (
		\a[16] ,
		\shift[0] ,
		_w328_
	);
	LUT2 #(
		.INIT('h8)
	) name193 (
		\a[15] ,
		\shift[0] ,
		_w329_
	);
	LUT2 #(
		.INIT('h1)
	) name194 (
		_w328_,
		_w329_,
		_w330_
	);
	LUT2 #(
		.INIT('h1)
	) name195 (
		\shift[1] ,
		_w330_,
		_w331_
	);
	LUT2 #(
		.INIT('h1)
	) name196 (
		_w327_,
		_w331_,
		_w332_
	);
	LUT2 #(
		.INIT('h2)
	) name197 (
		_w136_,
		_w332_,
		_w333_
	);
	LUT2 #(
		.INIT('h8)
	) name198 (
		\a[9] ,
		\shift[0] ,
		_w334_
	);
	LUT2 #(
		.INIT('h2)
	) name199 (
		\a[10] ,
		\shift[0] ,
		_w335_
	);
	LUT2 #(
		.INIT('h1)
	) name200 (
		_w334_,
		_w335_,
		_w336_
	);
	LUT2 #(
		.INIT('h2)
	) name201 (
		\shift[1] ,
		_w336_,
		_w337_
	);
	LUT2 #(
		.INIT('h2)
	) name202 (
		\a[12] ,
		\shift[0] ,
		_w338_
	);
	LUT2 #(
		.INIT('h8)
	) name203 (
		\a[11] ,
		\shift[0] ,
		_w339_
	);
	LUT2 #(
		.INIT('h1)
	) name204 (
		_w338_,
		_w339_,
		_w340_
	);
	LUT2 #(
		.INIT('h1)
	) name205 (
		\shift[1] ,
		_w340_,
		_w341_
	);
	LUT2 #(
		.INIT('h1)
	) name206 (
		_w337_,
		_w341_,
		_w342_
	);
	LUT2 #(
		.INIT('h2)
	) name207 (
		_w147_,
		_w342_,
		_w343_
	);
	LUT2 #(
		.INIT('h8)
	) name208 (
		\a[1] ,
		\shift[0] ,
		_w344_
	);
	LUT2 #(
		.INIT('h2)
	) name209 (
		\a[2] ,
		\shift[0] ,
		_w345_
	);
	LUT2 #(
		.INIT('h1)
	) name210 (
		_w344_,
		_w345_,
		_w346_
	);
	LUT2 #(
		.INIT('h2)
	) name211 (
		\shift[1] ,
		_w346_,
		_w347_
	);
	LUT2 #(
		.INIT('h2)
	) name212 (
		\a[4] ,
		\shift[0] ,
		_w348_
	);
	LUT2 #(
		.INIT('h8)
	) name213 (
		\a[3] ,
		\shift[0] ,
		_w349_
	);
	LUT2 #(
		.INIT('h1)
	) name214 (
		_w348_,
		_w349_,
		_w350_
	);
	LUT2 #(
		.INIT('h1)
	) name215 (
		\shift[1] ,
		_w350_,
		_w351_
	);
	LUT2 #(
		.INIT('h1)
	) name216 (
		_w347_,
		_w351_,
		_w352_
	);
	LUT2 #(
		.INIT('h2)
	) name217 (
		_w158_,
		_w352_,
		_w353_
	);
	LUT2 #(
		.INIT('h8)
	) name218 (
		\a[5] ,
		\shift[0] ,
		_w354_
	);
	LUT2 #(
		.INIT('h2)
	) name219 (
		\a[6] ,
		\shift[0] ,
		_w355_
	);
	LUT2 #(
		.INIT('h1)
	) name220 (
		_w354_,
		_w355_,
		_w356_
	);
	LUT2 #(
		.INIT('h2)
	) name221 (
		\shift[1] ,
		_w356_,
		_w357_
	);
	LUT2 #(
		.INIT('h2)
	) name222 (
		\a[8] ,
		\shift[0] ,
		_w358_
	);
	LUT2 #(
		.INIT('h8)
	) name223 (
		\a[7] ,
		\shift[0] ,
		_w359_
	);
	LUT2 #(
		.INIT('h1)
	) name224 (
		_w358_,
		_w359_,
		_w360_
	);
	LUT2 #(
		.INIT('h1)
	) name225 (
		\shift[1] ,
		_w360_,
		_w361_
	);
	LUT2 #(
		.INIT('h1)
	) name226 (
		_w357_,
		_w361_,
		_w362_
	);
	LUT2 #(
		.INIT('h2)
	) name227 (
		_w169_,
		_w362_,
		_w363_
	);
	LUT2 #(
		.INIT('h1)
	) name228 (
		_w333_,
		_w343_,
		_w364_
	);
	LUT2 #(
		.INIT('h1)
	) name229 (
		_w353_,
		_w363_,
		_w365_
	);
	LUT2 #(
		.INIT('h8)
	) name230 (
		_w364_,
		_w365_,
		_w366_
	);
	LUT2 #(
		.INIT('h2)
	) name231 (
		_w183_,
		_w366_,
		_w367_
	);
	LUT2 #(
		.INIT('h8)
	) name232 (
		\a[29] ,
		\shift[0] ,
		_w368_
	);
	LUT2 #(
		.INIT('h2)
	) name233 (
		\a[30] ,
		\shift[0] ,
		_w369_
	);
	LUT2 #(
		.INIT('h1)
	) name234 (
		_w368_,
		_w369_,
		_w370_
	);
	LUT2 #(
		.INIT('h2)
	) name235 (
		\shift[1] ,
		_w370_,
		_w371_
	);
	LUT2 #(
		.INIT('h2)
	) name236 (
		\a[32] ,
		\shift[0] ,
		_w372_
	);
	LUT2 #(
		.INIT('h8)
	) name237 (
		\a[31] ,
		\shift[0] ,
		_w373_
	);
	LUT2 #(
		.INIT('h1)
	) name238 (
		_w372_,
		_w373_,
		_w374_
	);
	LUT2 #(
		.INIT('h1)
	) name239 (
		\shift[1] ,
		_w374_,
		_w375_
	);
	LUT2 #(
		.INIT('h1)
	) name240 (
		_w371_,
		_w375_,
		_w376_
	);
	LUT2 #(
		.INIT('h2)
	) name241 (
		_w136_,
		_w376_,
		_w377_
	);
	LUT2 #(
		.INIT('h8)
	) name242 (
		\a[25] ,
		\shift[0] ,
		_w378_
	);
	LUT2 #(
		.INIT('h2)
	) name243 (
		\a[26] ,
		\shift[0] ,
		_w379_
	);
	LUT2 #(
		.INIT('h1)
	) name244 (
		_w378_,
		_w379_,
		_w380_
	);
	LUT2 #(
		.INIT('h2)
	) name245 (
		\shift[1] ,
		_w380_,
		_w381_
	);
	LUT2 #(
		.INIT('h2)
	) name246 (
		\a[28] ,
		\shift[0] ,
		_w382_
	);
	LUT2 #(
		.INIT('h8)
	) name247 (
		\a[27] ,
		\shift[0] ,
		_w383_
	);
	LUT2 #(
		.INIT('h1)
	) name248 (
		_w382_,
		_w383_,
		_w384_
	);
	LUT2 #(
		.INIT('h1)
	) name249 (
		\shift[1] ,
		_w384_,
		_w385_
	);
	LUT2 #(
		.INIT('h1)
	) name250 (
		_w381_,
		_w385_,
		_w386_
	);
	LUT2 #(
		.INIT('h2)
	) name251 (
		_w147_,
		_w386_,
		_w387_
	);
	LUT2 #(
		.INIT('h8)
	) name252 (
		\a[17] ,
		\shift[0] ,
		_w388_
	);
	LUT2 #(
		.INIT('h2)
	) name253 (
		\a[18] ,
		\shift[0] ,
		_w389_
	);
	LUT2 #(
		.INIT('h1)
	) name254 (
		_w388_,
		_w389_,
		_w390_
	);
	LUT2 #(
		.INIT('h2)
	) name255 (
		\shift[1] ,
		_w390_,
		_w391_
	);
	LUT2 #(
		.INIT('h2)
	) name256 (
		\a[20] ,
		\shift[0] ,
		_w392_
	);
	LUT2 #(
		.INIT('h8)
	) name257 (
		\a[19] ,
		\shift[0] ,
		_w393_
	);
	LUT2 #(
		.INIT('h1)
	) name258 (
		_w392_,
		_w393_,
		_w394_
	);
	LUT2 #(
		.INIT('h1)
	) name259 (
		\shift[1] ,
		_w394_,
		_w395_
	);
	LUT2 #(
		.INIT('h1)
	) name260 (
		_w391_,
		_w395_,
		_w396_
	);
	LUT2 #(
		.INIT('h2)
	) name261 (
		_w158_,
		_w396_,
		_w397_
	);
	LUT2 #(
		.INIT('h8)
	) name262 (
		\a[21] ,
		\shift[0] ,
		_w398_
	);
	LUT2 #(
		.INIT('h2)
	) name263 (
		\a[22] ,
		\shift[0] ,
		_w399_
	);
	LUT2 #(
		.INIT('h1)
	) name264 (
		_w398_,
		_w399_,
		_w400_
	);
	LUT2 #(
		.INIT('h2)
	) name265 (
		\shift[1] ,
		_w400_,
		_w401_
	);
	LUT2 #(
		.INIT('h2)
	) name266 (
		\a[24] ,
		\shift[0] ,
		_w402_
	);
	LUT2 #(
		.INIT('h8)
	) name267 (
		\a[23] ,
		\shift[0] ,
		_w403_
	);
	LUT2 #(
		.INIT('h1)
	) name268 (
		_w402_,
		_w403_,
		_w404_
	);
	LUT2 #(
		.INIT('h1)
	) name269 (
		\shift[1] ,
		_w404_,
		_w405_
	);
	LUT2 #(
		.INIT('h1)
	) name270 (
		_w401_,
		_w405_,
		_w406_
	);
	LUT2 #(
		.INIT('h2)
	) name271 (
		_w169_,
		_w406_,
		_w407_
	);
	LUT2 #(
		.INIT('h1)
	) name272 (
		_w377_,
		_w387_,
		_w408_
	);
	LUT2 #(
		.INIT('h1)
	) name273 (
		_w397_,
		_w407_,
		_w409_
	);
	LUT2 #(
		.INIT('h8)
	) name274 (
		_w408_,
		_w409_,
		_w410_
	);
	LUT2 #(
		.INIT('h2)
	) name275 (
		_w228_,
		_w410_,
		_w411_
	);
	LUT2 #(
		.INIT('h8)
	) name276 (
		\a[61] ,
		\shift[0] ,
		_w412_
	);
	LUT2 #(
		.INIT('h2)
	) name277 (
		\a[62] ,
		\shift[0] ,
		_w413_
	);
	LUT2 #(
		.INIT('h1)
	) name278 (
		_w412_,
		_w413_,
		_w414_
	);
	LUT2 #(
		.INIT('h2)
	) name279 (
		\shift[1] ,
		_w414_,
		_w415_
	);
	LUT2 #(
		.INIT('h2)
	) name280 (
		\a[64] ,
		\shift[0] ,
		_w416_
	);
	LUT2 #(
		.INIT('h8)
	) name281 (
		\a[63] ,
		\shift[0] ,
		_w417_
	);
	LUT2 #(
		.INIT('h1)
	) name282 (
		_w416_,
		_w417_,
		_w418_
	);
	LUT2 #(
		.INIT('h1)
	) name283 (
		\shift[1] ,
		_w418_,
		_w419_
	);
	LUT2 #(
		.INIT('h1)
	) name284 (
		_w415_,
		_w419_,
		_w420_
	);
	LUT2 #(
		.INIT('h2)
	) name285 (
		_w136_,
		_w420_,
		_w421_
	);
	LUT2 #(
		.INIT('h8)
	) name286 (
		\a[57] ,
		\shift[0] ,
		_w422_
	);
	LUT2 #(
		.INIT('h2)
	) name287 (
		\a[58] ,
		\shift[0] ,
		_w423_
	);
	LUT2 #(
		.INIT('h1)
	) name288 (
		_w422_,
		_w423_,
		_w424_
	);
	LUT2 #(
		.INIT('h2)
	) name289 (
		\shift[1] ,
		_w424_,
		_w425_
	);
	LUT2 #(
		.INIT('h2)
	) name290 (
		\a[60] ,
		\shift[0] ,
		_w426_
	);
	LUT2 #(
		.INIT('h8)
	) name291 (
		\a[59] ,
		\shift[0] ,
		_w427_
	);
	LUT2 #(
		.INIT('h1)
	) name292 (
		_w426_,
		_w427_,
		_w428_
	);
	LUT2 #(
		.INIT('h1)
	) name293 (
		\shift[1] ,
		_w428_,
		_w429_
	);
	LUT2 #(
		.INIT('h1)
	) name294 (
		_w425_,
		_w429_,
		_w430_
	);
	LUT2 #(
		.INIT('h2)
	) name295 (
		_w147_,
		_w430_,
		_w431_
	);
	LUT2 #(
		.INIT('h8)
	) name296 (
		\a[49] ,
		\shift[0] ,
		_w432_
	);
	LUT2 #(
		.INIT('h2)
	) name297 (
		\a[50] ,
		\shift[0] ,
		_w433_
	);
	LUT2 #(
		.INIT('h1)
	) name298 (
		_w432_,
		_w433_,
		_w434_
	);
	LUT2 #(
		.INIT('h2)
	) name299 (
		\shift[1] ,
		_w434_,
		_w435_
	);
	LUT2 #(
		.INIT('h2)
	) name300 (
		\a[52] ,
		\shift[0] ,
		_w436_
	);
	LUT2 #(
		.INIT('h8)
	) name301 (
		\a[51] ,
		\shift[0] ,
		_w437_
	);
	LUT2 #(
		.INIT('h1)
	) name302 (
		_w436_,
		_w437_,
		_w438_
	);
	LUT2 #(
		.INIT('h1)
	) name303 (
		\shift[1] ,
		_w438_,
		_w439_
	);
	LUT2 #(
		.INIT('h1)
	) name304 (
		_w435_,
		_w439_,
		_w440_
	);
	LUT2 #(
		.INIT('h2)
	) name305 (
		_w158_,
		_w440_,
		_w441_
	);
	LUT2 #(
		.INIT('h8)
	) name306 (
		\a[53] ,
		\shift[0] ,
		_w442_
	);
	LUT2 #(
		.INIT('h2)
	) name307 (
		\a[54] ,
		\shift[0] ,
		_w443_
	);
	LUT2 #(
		.INIT('h1)
	) name308 (
		_w442_,
		_w443_,
		_w444_
	);
	LUT2 #(
		.INIT('h2)
	) name309 (
		\shift[1] ,
		_w444_,
		_w445_
	);
	LUT2 #(
		.INIT('h2)
	) name310 (
		\a[56] ,
		\shift[0] ,
		_w446_
	);
	LUT2 #(
		.INIT('h8)
	) name311 (
		\a[55] ,
		\shift[0] ,
		_w447_
	);
	LUT2 #(
		.INIT('h1)
	) name312 (
		_w446_,
		_w447_,
		_w448_
	);
	LUT2 #(
		.INIT('h1)
	) name313 (
		\shift[1] ,
		_w448_,
		_w449_
	);
	LUT2 #(
		.INIT('h1)
	) name314 (
		_w445_,
		_w449_,
		_w450_
	);
	LUT2 #(
		.INIT('h2)
	) name315 (
		_w169_,
		_w450_,
		_w451_
	);
	LUT2 #(
		.INIT('h1)
	) name316 (
		_w421_,
		_w431_,
		_w452_
	);
	LUT2 #(
		.INIT('h1)
	) name317 (
		_w441_,
		_w451_,
		_w453_
	);
	LUT2 #(
		.INIT('h8)
	) name318 (
		_w452_,
		_w453_,
		_w454_
	);
	LUT2 #(
		.INIT('h2)
	) name319 (
		_w273_,
		_w454_,
		_w455_
	);
	LUT2 #(
		.INIT('h8)
	) name320 (
		\a[45] ,
		\shift[0] ,
		_w456_
	);
	LUT2 #(
		.INIT('h2)
	) name321 (
		\a[46] ,
		\shift[0] ,
		_w457_
	);
	LUT2 #(
		.INIT('h1)
	) name322 (
		_w456_,
		_w457_,
		_w458_
	);
	LUT2 #(
		.INIT('h2)
	) name323 (
		\shift[1] ,
		_w458_,
		_w459_
	);
	LUT2 #(
		.INIT('h2)
	) name324 (
		\a[48] ,
		\shift[0] ,
		_w460_
	);
	LUT2 #(
		.INIT('h8)
	) name325 (
		\a[47] ,
		\shift[0] ,
		_w461_
	);
	LUT2 #(
		.INIT('h1)
	) name326 (
		_w460_,
		_w461_,
		_w462_
	);
	LUT2 #(
		.INIT('h1)
	) name327 (
		\shift[1] ,
		_w462_,
		_w463_
	);
	LUT2 #(
		.INIT('h1)
	) name328 (
		_w459_,
		_w463_,
		_w464_
	);
	LUT2 #(
		.INIT('h2)
	) name329 (
		_w136_,
		_w464_,
		_w465_
	);
	LUT2 #(
		.INIT('h8)
	) name330 (
		\a[41] ,
		\shift[0] ,
		_w466_
	);
	LUT2 #(
		.INIT('h2)
	) name331 (
		\a[42] ,
		\shift[0] ,
		_w467_
	);
	LUT2 #(
		.INIT('h1)
	) name332 (
		_w466_,
		_w467_,
		_w468_
	);
	LUT2 #(
		.INIT('h2)
	) name333 (
		\shift[1] ,
		_w468_,
		_w469_
	);
	LUT2 #(
		.INIT('h2)
	) name334 (
		\a[44] ,
		\shift[0] ,
		_w470_
	);
	LUT2 #(
		.INIT('h8)
	) name335 (
		\a[43] ,
		\shift[0] ,
		_w471_
	);
	LUT2 #(
		.INIT('h1)
	) name336 (
		_w470_,
		_w471_,
		_w472_
	);
	LUT2 #(
		.INIT('h1)
	) name337 (
		\shift[1] ,
		_w472_,
		_w473_
	);
	LUT2 #(
		.INIT('h1)
	) name338 (
		_w469_,
		_w473_,
		_w474_
	);
	LUT2 #(
		.INIT('h2)
	) name339 (
		_w147_,
		_w474_,
		_w475_
	);
	LUT2 #(
		.INIT('h8)
	) name340 (
		\a[33] ,
		\shift[0] ,
		_w476_
	);
	LUT2 #(
		.INIT('h2)
	) name341 (
		\a[34] ,
		\shift[0] ,
		_w477_
	);
	LUT2 #(
		.INIT('h1)
	) name342 (
		_w476_,
		_w477_,
		_w478_
	);
	LUT2 #(
		.INIT('h2)
	) name343 (
		\shift[1] ,
		_w478_,
		_w479_
	);
	LUT2 #(
		.INIT('h2)
	) name344 (
		\a[36] ,
		\shift[0] ,
		_w480_
	);
	LUT2 #(
		.INIT('h8)
	) name345 (
		\a[35] ,
		\shift[0] ,
		_w481_
	);
	LUT2 #(
		.INIT('h1)
	) name346 (
		_w480_,
		_w481_,
		_w482_
	);
	LUT2 #(
		.INIT('h1)
	) name347 (
		\shift[1] ,
		_w482_,
		_w483_
	);
	LUT2 #(
		.INIT('h1)
	) name348 (
		_w479_,
		_w483_,
		_w484_
	);
	LUT2 #(
		.INIT('h2)
	) name349 (
		_w158_,
		_w484_,
		_w485_
	);
	LUT2 #(
		.INIT('h2)
	) name350 (
		\a[40] ,
		\shift[0] ,
		_w486_
	);
	LUT2 #(
		.INIT('h1)
	) name351 (
		\shift[1] ,
		_w486_,
		_w487_
	);
	LUT2 #(
		.INIT('h8)
	) name352 (
		\a[37] ,
		\shift[0] ,
		_w488_
	);
	LUT2 #(
		.INIT('h2)
	) name353 (
		\shift[1] ,
		_w488_,
		_w489_
	);
	LUT2 #(
		.INIT('h1)
	) name354 (
		_w487_,
		_w489_,
		_w490_
	);
	LUT2 #(
		.INIT('h2)
	) name355 (
		\a[38] ,
		\shift[0] ,
		_w491_
	);
	LUT2 #(
		.INIT('h8)
	) name356 (
		\shift[1] ,
		_w491_,
		_w492_
	);
	LUT2 #(
		.INIT('h8)
	) name357 (
		\a[39] ,
		\shift[0] ,
		_w493_
	);
	LUT2 #(
		.INIT('h4)
	) name358 (
		\shift[1] ,
		_w493_,
		_w494_
	);
	LUT2 #(
		.INIT('h1)
	) name359 (
		_w492_,
		_w494_,
		_w495_
	);
	LUT2 #(
		.INIT('h4)
	) name360 (
		_w490_,
		_w495_,
		_w496_
	);
	LUT2 #(
		.INIT('h2)
	) name361 (
		_w169_,
		_w496_,
		_w497_
	);
	LUT2 #(
		.INIT('h1)
	) name362 (
		_w465_,
		_w475_,
		_w498_
	);
	LUT2 #(
		.INIT('h1)
	) name363 (
		_w485_,
		_w497_,
		_w499_
	);
	LUT2 #(
		.INIT('h8)
	) name364 (
		_w498_,
		_w499_,
		_w500_
	);
	LUT2 #(
		.INIT('h2)
	) name365 (
		_w318_,
		_w500_,
		_w501_
	);
	LUT2 #(
		.INIT('h1)
	) name366 (
		_w367_,
		_w411_,
		_w502_
	);
	LUT2 #(
		.INIT('h1)
	) name367 (
		_w455_,
		_w501_,
		_w503_
	);
	LUT2 #(
		.INIT('h8)
	) name368 (
		_w502_,
		_w503_,
		_w504_
	);
	LUT2 #(
		.INIT('h2)
	) name369 (
		\shift[6] ,
		_w504_,
		_w505_
	);
	LUT2 #(
		.INIT('h1)
	) name370 (
		_w323_,
		_w505_,
		_w506_
	);
	LUT2 #(
		.INIT('h2)
	) name371 (
		\a[81] ,
		\shift[0] ,
		_w507_
	);
	LUT2 #(
		.INIT('h1)
	) name372 (
		\shift[1] ,
		_w507_,
		_w508_
	);
	LUT2 #(
		.INIT('h8)
	) name373 (
		\a[78] ,
		\shift[0] ,
		_w509_
	);
	LUT2 #(
		.INIT('h2)
	) name374 (
		\shift[1] ,
		_w509_,
		_w510_
	);
	LUT2 #(
		.INIT('h1)
	) name375 (
		_w508_,
		_w510_,
		_w511_
	);
	LUT2 #(
		.INIT('h2)
	) name376 (
		\a[79] ,
		\shift[0] ,
		_w512_
	);
	LUT2 #(
		.INIT('h8)
	) name377 (
		\shift[1] ,
		_w512_,
		_w513_
	);
	LUT2 #(
		.INIT('h8)
	) name378 (
		\a[80] ,
		\shift[0] ,
		_w514_
	);
	LUT2 #(
		.INIT('h4)
	) name379 (
		\shift[1] ,
		_w514_,
		_w515_
	);
	LUT2 #(
		.INIT('h1)
	) name380 (
		_w513_,
		_w515_,
		_w516_
	);
	LUT2 #(
		.INIT('h4)
	) name381 (
		_w511_,
		_w516_,
		_w517_
	);
	LUT2 #(
		.INIT('h2)
	) name382 (
		_w136_,
		_w517_,
		_w518_
	);
	LUT2 #(
		.INIT('h2)
	) name383 (
		\a[77] ,
		\shift[0] ,
		_w519_
	);
	LUT2 #(
		.INIT('h1)
	) name384 (
		\shift[1] ,
		_w519_,
		_w520_
	);
	LUT2 #(
		.INIT('h8)
	) name385 (
		\a[74] ,
		\shift[0] ,
		_w521_
	);
	LUT2 #(
		.INIT('h2)
	) name386 (
		\shift[1] ,
		_w521_,
		_w522_
	);
	LUT2 #(
		.INIT('h1)
	) name387 (
		_w520_,
		_w522_,
		_w523_
	);
	LUT2 #(
		.INIT('h2)
	) name388 (
		\a[75] ,
		\shift[0] ,
		_w524_
	);
	LUT2 #(
		.INIT('h8)
	) name389 (
		\shift[1] ,
		_w524_,
		_w525_
	);
	LUT2 #(
		.INIT('h8)
	) name390 (
		\a[76] ,
		\shift[0] ,
		_w526_
	);
	LUT2 #(
		.INIT('h4)
	) name391 (
		\shift[1] ,
		_w526_,
		_w527_
	);
	LUT2 #(
		.INIT('h1)
	) name392 (
		_w525_,
		_w527_,
		_w528_
	);
	LUT2 #(
		.INIT('h4)
	) name393 (
		_w523_,
		_w528_,
		_w529_
	);
	LUT2 #(
		.INIT('h2)
	) name394 (
		_w147_,
		_w529_,
		_w530_
	);
	LUT2 #(
		.INIT('h2)
	) name395 (
		\a[69] ,
		\shift[0] ,
		_w531_
	);
	LUT2 #(
		.INIT('h1)
	) name396 (
		\shift[1] ,
		_w531_,
		_w532_
	);
	LUT2 #(
		.INIT('h8)
	) name397 (
		\a[66] ,
		\shift[0] ,
		_w533_
	);
	LUT2 #(
		.INIT('h2)
	) name398 (
		\shift[1] ,
		_w533_,
		_w534_
	);
	LUT2 #(
		.INIT('h1)
	) name399 (
		_w532_,
		_w534_,
		_w535_
	);
	LUT2 #(
		.INIT('h2)
	) name400 (
		\a[67] ,
		\shift[0] ,
		_w536_
	);
	LUT2 #(
		.INIT('h8)
	) name401 (
		\shift[1] ,
		_w536_,
		_w537_
	);
	LUT2 #(
		.INIT('h8)
	) name402 (
		\a[68] ,
		\shift[0] ,
		_w538_
	);
	LUT2 #(
		.INIT('h4)
	) name403 (
		\shift[1] ,
		_w538_,
		_w539_
	);
	LUT2 #(
		.INIT('h1)
	) name404 (
		_w537_,
		_w539_,
		_w540_
	);
	LUT2 #(
		.INIT('h4)
	) name405 (
		_w535_,
		_w540_,
		_w541_
	);
	LUT2 #(
		.INIT('h2)
	) name406 (
		_w158_,
		_w541_,
		_w542_
	);
	LUT2 #(
		.INIT('h2)
	) name407 (
		\a[73] ,
		\shift[0] ,
		_w543_
	);
	LUT2 #(
		.INIT('h1)
	) name408 (
		\shift[1] ,
		_w543_,
		_w544_
	);
	LUT2 #(
		.INIT('h8)
	) name409 (
		\a[70] ,
		\shift[0] ,
		_w545_
	);
	LUT2 #(
		.INIT('h2)
	) name410 (
		\shift[1] ,
		_w545_,
		_w546_
	);
	LUT2 #(
		.INIT('h1)
	) name411 (
		_w544_,
		_w546_,
		_w547_
	);
	LUT2 #(
		.INIT('h2)
	) name412 (
		\a[71] ,
		\shift[0] ,
		_w548_
	);
	LUT2 #(
		.INIT('h8)
	) name413 (
		\shift[1] ,
		_w548_,
		_w549_
	);
	LUT2 #(
		.INIT('h8)
	) name414 (
		\a[72] ,
		\shift[0] ,
		_w550_
	);
	LUT2 #(
		.INIT('h4)
	) name415 (
		\shift[1] ,
		_w550_,
		_w551_
	);
	LUT2 #(
		.INIT('h1)
	) name416 (
		_w549_,
		_w551_,
		_w552_
	);
	LUT2 #(
		.INIT('h4)
	) name417 (
		_w547_,
		_w552_,
		_w553_
	);
	LUT2 #(
		.INIT('h2)
	) name418 (
		_w169_,
		_w553_,
		_w554_
	);
	LUT2 #(
		.INIT('h1)
	) name419 (
		_w518_,
		_w530_,
		_w555_
	);
	LUT2 #(
		.INIT('h1)
	) name420 (
		_w542_,
		_w554_,
		_w556_
	);
	LUT2 #(
		.INIT('h8)
	) name421 (
		_w555_,
		_w556_,
		_w557_
	);
	LUT2 #(
		.INIT('h2)
	) name422 (
		_w183_,
		_w557_,
		_w558_
	);
	LUT2 #(
		.INIT('h2)
	) name423 (
		\a[97] ,
		\shift[0] ,
		_w559_
	);
	LUT2 #(
		.INIT('h1)
	) name424 (
		\shift[1] ,
		_w559_,
		_w560_
	);
	LUT2 #(
		.INIT('h8)
	) name425 (
		\a[94] ,
		\shift[0] ,
		_w561_
	);
	LUT2 #(
		.INIT('h2)
	) name426 (
		\shift[1] ,
		_w561_,
		_w562_
	);
	LUT2 #(
		.INIT('h1)
	) name427 (
		_w560_,
		_w562_,
		_w563_
	);
	LUT2 #(
		.INIT('h2)
	) name428 (
		\a[95] ,
		\shift[0] ,
		_w564_
	);
	LUT2 #(
		.INIT('h8)
	) name429 (
		\shift[1] ,
		_w564_,
		_w565_
	);
	LUT2 #(
		.INIT('h8)
	) name430 (
		\a[96] ,
		\shift[0] ,
		_w566_
	);
	LUT2 #(
		.INIT('h4)
	) name431 (
		\shift[1] ,
		_w566_,
		_w567_
	);
	LUT2 #(
		.INIT('h1)
	) name432 (
		_w565_,
		_w567_,
		_w568_
	);
	LUT2 #(
		.INIT('h4)
	) name433 (
		_w563_,
		_w568_,
		_w569_
	);
	LUT2 #(
		.INIT('h2)
	) name434 (
		_w136_,
		_w569_,
		_w570_
	);
	LUT2 #(
		.INIT('h2)
	) name435 (
		\a[93] ,
		\shift[0] ,
		_w571_
	);
	LUT2 #(
		.INIT('h1)
	) name436 (
		\shift[1] ,
		_w571_,
		_w572_
	);
	LUT2 #(
		.INIT('h8)
	) name437 (
		\a[90] ,
		\shift[0] ,
		_w573_
	);
	LUT2 #(
		.INIT('h2)
	) name438 (
		\shift[1] ,
		_w573_,
		_w574_
	);
	LUT2 #(
		.INIT('h1)
	) name439 (
		_w572_,
		_w574_,
		_w575_
	);
	LUT2 #(
		.INIT('h2)
	) name440 (
		\a[91] ,
		\shift[0] ,
		_w576_
	);
	LUT2 #(
		.INIT('h8)
	) name441 (
		\shift[1] ,
		_w576_,
		_w577_
	);
	LUT2 #(
		.INIT('h8)
	) name442 (
		\a[92] ,
		\shift[0] ,
		_w578_
	);
	LUT2 #(
		.INIT('h4)
	) name443 (
		\shift[1] ,
		_w578_,
		_w579_
	);
	LUT2 #(
		.INIT('h1)
	) name444 (
		_w577_,
		_w579_,
		_w580_
	);
	LUT2 #(
		.INIT('h4)
	) name445 (
		_w575_,
		_w580_,
		_w581_
	);
	LUT2 #(
		.INIT('h2)
	) name446 (
		_w147_,
		_w581_,
		_w582_
	);
	LUT2 #(
		.INIT('h2)
	) name447 (
		\a[85] ,
		\shift[0] ,
		_w583_
	);
	LUT2 #(
		.INIT('h1)
	) name448 (
		\shift[1] ,
		_w583_,
		_w584_
	);
	LUT2 #(
		.INIT('h8)
	) name449 (
		\a[82] ,
		\shift[0] ,
		_w585_
	);
	LUT2 #(
		.INIT('h2)
	) name450 (
		\shift[1] ,
		_w585_,
		_w586_
	);
	LUT2 #(
		.INIT('h1)
	) name451 (
		_w584_,
		_w586_,
		_w587_
	);
	LUT2 #(
		.INIT('h2)
	) name452 (
		\a[83] ,
		\shift[0] ,
		_w588_
	);
	LUT2 #(
		.INIT('h8)
	) name453 (
		\shift[1] ,
		_w588_,
		_w589_
	);
	LUT2 #(
		.INIT('h8)
	) name454 (
		\a[84] ,
		\shift[0] ,
		_w590_
	);
	LUT2 #(
		.INIT('h4)
	) name455 (
		\shift[1] ,
		_w590_,
		_w591_
	);
	LUT2 #(
		.INIT('h1)
	) name456 (
		_w589_,
		_w591_,
		_w592_
	);
	LUT2 #(
		.INIT('h4)
	) name457 (
		_w587_,
		_w592_,
		_w593_
	);
	LUT2 #(
		.INIT('h2)
	) name458 (
		_w158_,
		_w593_,
		_w594_
	);
	LUT2 #(
		.INIT('h2)
	) name459 (
		\a[89] ,
		\shift[0] ,
		_w595_
	);
	LUT2 #(
		.INIT('h1)
	) name460 (
		\shift[1] ,
		_w595_,
		_w596_
	);
	LUT2 #(
		.INIT('h8)
	) name461 (
		\a[86] ,
		\shift[0] ,
		_w597_
	);
	LUT2 #(
		.INIT('h2)
	) name462 (
		\shift[1] ,
		_w597_,
		_w598_
	);
	LUT2 #(
		.INIT('h1)
	) name463 (
		_w596_,
		_w598_,
		_w599_
	);
	LUT2 #(
		.INIT('h2)
	) name464 (
		\a[87] ,
		\shift[0] ,
		_w600_
	);
	LUT2 #(
		.INIT('h8)
	) name465 (
		\shift[1] ,
		_w600_,
		_w601_
	);
	LUT2 #(
		.INIT('h8)
	) name466 (
		\a[88] ,
		\shift[0] ,
		_w602_
	);
	LUT2 #(
		.INIT('h4)
	) name467 (
		\shift[1] ,
		_w602_,
		_w603_
	);
	LUT2 #(
		.INIT('h1)
	) name468 (
		_w601_,
		_w603_,
		_w604_
	);
	LUT2 #(
		.INIT('h4)
	) name469 (
		_w599_,
		_w604_,
		_w605_
	);
	LUT2 #(
		.INIT('h2)
	) name470 (
		_w169_,
		_w605_,
		_w606_
	);
	LUT2 #(
		.INIT('h1)
	) name471 (
		_w570_,
		_w582_,
		_w607_
	);
	LUT2 #(
		.INIT('h1)
	) name472 (
		_w594_,
		_w606_,
		_w608_
	);
	LUT2 #(
		.INIT('h8)
	) name473 (
		_w607_,
		_w608_,
		_w609_
	);
	LUT2 #(
		.INIT('h2)
	) name474 (
		_w228_,
		_w609_,
		_w610_
	);
	LUT2 #(
		.INIT('h2)
	) name475 (
		\a[1] ,
		\shift[0] ,
		_w611_
	);
	LUT2 #(
		.INIT('h1)
	) name476 (
		\shift[1] ,
		_w611_,
		_w612_
	);
	LUT2 #(
		.INIT('h8)
	) name477 (
		\a[126] ,
		\shift[0] ,
		_w613_
	);
	LUT2 #(
		.INIT('h2)
	) name478 (
		\shift[1] ,
		_w613_,
		_w614_
	);
	LUT2 #(
		.INIT('h1)
	) name479 (
		_w612_,
		_w614_,
		_w615_
	);
	LUT2 #(
		.INIT('h2)
	) name480 (
		\a[127] ,
		\shift[0] ,
		_w616_
	);
	LUT2 #(
		.INIT('h8)
	) name481 (
		\shift[1] ,
		_w616_,
		_w617_
	);
	LUT2 #(
		.INIT('h8)
	) name482 (
		\a[0] ,
		\shift[0] ,
		_w618_
	);
	LUT2 #(
		.INIT('h4)
	) name483 (
		\shift[1] ,
		_w618_,
		_w619_
	);
	LUT2 #(
		.INIT('h1)
	) name484 (
		_w617_,
		_w619_,
		_w620_
	);
	LUT2 #(
		.INIT('h4)
	) name485 (
		_w615_,
		_w620_,
		_w621_
	);
	LUT2 #(
		.INIT('h2)
	) name486 (
		_w136_,
		_w621_,
		_w622_
	);
	LUT2 #(
		.INIT('h2)
	) name487 (
		\a[125] ,
		\shift[0] ,
		_w623_
	);
	LUT2 #(
		.INIT('h1)
	) name488 (
		\shift[1] ,
		_w623_,
		_w624_
	);
	LUT2 #(
		.INIT('h8)
	) name489 (
		\a[122] ,
		\shift[0] ,
		_w625_
	);
	LUT2 #(
		.INIT('h2)
	) name490 (
		\shift[1] ,
		_w625_,
		_w626_
	);
	LUT2 #(
		.INIT('h1)
	) name491 (
		_w624_,
		_w626_,
		_w627_
	);
	LUT2 #(
		.INIT('h2)
	) name492 (
		\a[123] ,
		\shift[0] ,
		_w628_
	);
	LUT2 #(
		.INIT('h8)
	) name493 (
		\shift[1] ,
		_w628_,
		_w629_
	);
	LUT2 #(
		.INIT('h8)
	) name494 (
		\a[124] ,
		\shift[0] ,
		_w630_
	);
	LUT2 #(
		.INIT('h4)
	) name495 (
		\shift[1] ,
		_w630_,
		_w631_
	);
	LUT2 #(
		.INIT('h1)
	) name496 (
		_w629_,
		_w631_,
		_w632_
	);
	LUT2 #(
		.INIT('h4)
	) name497 (
		_w627_,
		_w632_,
		_w633_
	);
	LUT2 #(
		.INIT('h2)
	) name498 (
		_w147_,
		_w633_,
		_w634_
	);
	LUT2 #(
		.INIT('h2)
	) name499 (
		\a[117] ,
		\shift[0] ,
		_w635_
	);
	LUT2 #(
		.INIT('h1)
	) name500 (
		\shift[1] ,
		_w635_,
		_w636_
	);
	LUT2 #(
		.INIT('h8)
	) name501 (
		\a[114] ,
		\shift[0] ,
		_w637_
	);
	LUT2 #(
		.INIT('h2)
	) name502 (
		\shift[1] ,
		_w637_,
		_w638_
	);
	LUT2 #(
		.INIT('h1)
	) name503 (
		_w636_,
		_w638_,
		_w639_
	);
	LUT2 #(
		.INIT('h2)
	) name504 (
		\a[115] ,
		\shift[0] ,
		_w640_
	);
	LUT2 #(
		.INIT('h8)
	) name505 (
		\shift[1] ,
		_w640_,
		_w641_
	);
	LUT2 #(
		.INIT('h8)
	) name506 (
		\a[116] ,
		\shift[0] ,
		_w642_
	);
	LUT2 #(
		.INIT('h4)
	) name507 (
		\shift[1] ,
		_w642_,
		_w643_
	);
	LUT2 #(
		.INIT('h1)
	) name508 (
		_w641_,
		_w643_,
		_w644_
	);
	LUT2 #(
		.INIT('h4)
	) name509 (
		_w639_,
		_w644_,
		_w645_
	);
	LUT2 #(
		.INIT('h2)
	) name510 (
		_w158_,
		_w645_,
		_w646_
	);
	LUT2 #(
		.INIT('h2)
	) name511 (
		\a[121] ,
		\shift[0] ,
		_w647_
	);
	LUT2 #(
		.INIT('h1)
	) name512 (
		\shift[1] ,
		_w647_,
		_w648_
	);
	LUT2 #(
		.INIT('h8)
	) name513 (
		\a[118] ,
		\shift[0] ,
		_w649_
	);
	LUT2 #(
		.INIT('h2)
	) name514 (
		\shift[1] ,
		_w649_,
		_w650_
	);
	LUT2 #(
		.INIT('h1)
	) name515 (
		_w648_,
		_w650_,
		_w651_
	);
	LUT2 #(
		.INIT('h2)
	) name516 (
		\a[119] ,
		\shift[0] ,
		_w652_
	);
	LUT2 #(
		.INIT('h8)
	) name517 (
		\shift[1] ,
		_w652_,
		_w653_
	);
	LUT2 #(
		.INIT('h8)
	) name518 (
		\a[120] ,
		\shift[0] ,
		_w654_
	);
	LUT2 #(
		.INIT('h4)
	) name519 (
		\shift[1] ,
		_w654_,
		_w655_
	);
	LUT2 #(
		.INIT('h1)
	) name520 (
		_w653_,
		_w655_,
		_w656_
	);
	LUT2 #(
		.INIT('h4)
	) name521 (
		_w651_,
		_w656_,
		_w657_
	);
	LUT2 #(
		.INIT('h2)
	) name522 (
		_w169_,
		_w657_,
		_w658_
	);
	LUT2 #(
		.INIT('h1)
	) name523 (
		_w622_,
		_w634_,
		_w659_
	);
	LUT2 #(
		.INIT('h1)
	) name524 (
		_w646_,
		_w658_,
		_w660_
	);
	LUT2 #(
		.INIT('h8)
	) name525 (
		_w659_,
		_w660_,
		_w661_
	);
	LUT2 #(
		.INIT('h2)
	) name526 (
		_w273_,
		_w661_,
		_w662_
	);
	LUT2 #(
		.INIT('h2)
	) name527 (
		\a[113] ,
		\shift[0] ,
		_w663_
	);
	LUT2 #(
		.INIT('h1)
	) name528 (
		\shift[1] ,
		_w663_,
		_w664_
	);
	LUT2 #(
		.INIT('h8)
	) name529 (
		\a[110] ,
		\shift[0] ,
		_w665_
	);
	LUT2 #(
		.INIT('h2)
	) name530 (
		\shift[1] ,
		_w665_,
		_w666_
	);
	LUT2 #(
		.INIT('h1)
	) name531 (
		_w664_,
		_w666_,
		_w667_
	);
	LUT2 #(
		.INIT('h2)
	) name532 (
		\a[111] ,
		\shift[0] ,
		_w668_
	);
	LUT2 #(
		.INIT('h8)
	) name533 (
		\shift[1] ,
		_w668_,
		_w669_
	);
	LUT2 #(
		.INIT('h8)
	) name534 (
		\a[112] ,
		\shift[0] ,
		_w670_
	);
	LUT2 #(
		.INIT('h4)
	) name535 (
		\shift[1] ,
		_w670_,
		_w671_
	);
	LUT2 #(
		.INIT('h1)
	) name536 (
		_w669_,
		_w671_,
		_w672_
	);
	LUT2 #(
		.INIT('h4)
	) name537 (
		_w667_,
		_w672_,
		_w673_
	);
	LUT2 #(
		.INIT('h2)
	) name538 (
		_w136_,
		_w673_,
		_w674_
	);
	LUT2 #(
		.INIT('h2)
	) name539 (
		\a[109] ,
		\shift[0] ,
		_w675_
	);
	LUT2 #(
		.INIT('h1)
	) name540 (
		\shift[1] ,
		_w675_,
		_w676_
	);
	LUT2 #(
		.INIT('h8)
	) name541 (
		\a[106] ,
		\shift[0] ,
		_w677_
	);
	LUT2 #(
		.INIT('h2)
	) name542 (
		\shift[1] ,
		_w677_,
		_w678_
	);
	LUT2 #(
		.INIT('h1)
	) name543 (
		_w676_,
		_w678_,
		_w679_
	);
	LUT2 #(
		.INIT('h2)
	) name544 (
		\a[107] ,
		\shift[0] ,
		_w680_
	);
	LUT2 #(
		.INIT('h8)
	) name545 (
		\shift[1] ,
		_w680_,
		_w681_
	);
	LUT2 #(
		.INIT('h8)
	) name546 (
		\a[108] ,
		\shift[0] ,
		_w682_
	);
	LUT2 #(
		.INIT('h4)
	) name547 (
		\shift[1] ,
		_w682_,
		_w683_
	);
	LUT2 #(
		.INIT('h1)
	) name548 (
		_w681_,
		_w683_,
		_w684_
	);
	LUT2 #(
		.INIT('h4)
	) name549 (
		_w679_,
		_w684_,
		_w685_
	);
	LUT2 #(
		.INIT('h2)
	) name550 (
		_w147_,
		_w685_,
		_w686_
	);
	LUT2 #(
		.INIT('h2)
	) name551 (
		\a[101] ,
		\shift[0] ,
		_w687_
	);
	LUT2 #(
		.INIT('h1)
	) name552 (
		\shift[1] ,
		_w687_,
		_w688_
	);
	LUT2 #(
		.INIT('h8)
	) name553 (
		\a[98] ,
		\shift[0] ,
		_w689_
	);
	LUT2 #(
		.INIT('h2)
	) name554 (
		\shift[1] ,
		_w689_,
		_w690_
	);
	LUT2 #(
		.INIT('h1)
	) name555 (
		_w688_,
		_w690_,
		_w691_
	);
	LUT2 #(
		.INIT('h2)
	) name556 (
		\a[99] ,
		\shift[0] ,
		_w692_
	);
	LUT2 #(
		.INIT('h8)
	) name557 (
		\shift[1] ,
		_w692_,
		_w693_
	);
	LUT2 #(
		.INIT('h8)
	) name558 (
		\a[100] ,
		\shift[0] ,
		_w694_
	);
	LUT2 #(
		.INIT('h4)
	) name559 (
		\shift[1] ,
		_w694_,
		_w695_
	);
	LUT2 #(
		.INIT('h1)
	) name560 (
		_w693_,
		_w695_,
		_w696_
	);
	LUT2 #(
		.INIT('h4)
	) name561 (
		_w691_,
		_w696_,
		_w697_
	);
	LUT2 #(
		.INIT('h2)
	) name562 (
		_w158_,
		_w697_,
		_w698_
	);
	LUT2 #(
		.INIT('h2)
	) name563 (
		\a[105] ,
		\shift[0] ,
		_w699_
	);
	LUT2 #(
		.INIT('h1)
	) name564 (
		\shift[1] ,
		_w699_,
		_w700_
	);
	LUT2 #(
		.INIT('h8)
	) name565 (
		\a[102] ,
		\shift[0] ,
		_w701_
	);
	LUT2 #(
		.INIT('h2)
	) name566 (
		\shift[1] ,
		_w701_,
		_w702_
	);
	LUT2 #(
		.INIT('h1)
	) name567 (
		_w700_,
		_w702_,
		_w703_
	);
	LUT2 #(
		.INIT('h2)
	) name568 (
		\a[103] ,
		\shift[0] ,
		_w704_
	);
	LUT2 #(
		.INIT('h8)
	) name569 (
		\shift[1] ,
		_w704_,
		_w705_
	);
	LUT2 #(
		.INIT('h8)
	) name570 (
		\a[104] ,
		\shift[0] ,
		_w706_
	);
	LUT2 #(
		.INIT('h4)
	) name571 (
		\shift[1] ,
		_w706_,
		_w707_
	);
	LUT2 #(
		.INIT('h1)
	) name572 (
		_w705_,
		_w707_,
		_w708_
	);
	LUT2 #(
		.INIT('h4)
	) name573 (
		_w703_,
		_w708_,
		_w709_
	);
	LUT2 #(
		.INIT('h2)
	) name574 (
		_w169_,
		_w709_,
		_w710_
	);
	LUT2 #(
		.INIT('h1)
	) name575 (
		_w674_,
		_w686_,
		_w711_
	);
	LUT2 #(
		.INIT('h1)
	) name576 (
		_w698_,
		_w710_,
		_w712_
	);
	LUT2 #(
		.INIT('h8)
	) name577 (
		_w711_,
		_w712_,
		_w713_
	);
	LUT2 #(
		.INIT('h2)
	) name578 (
		_w318_,
		_w713_,
		_w714_
	);
	LUT2 #(
		.INIT('h1)
	) name579 (
		_w558_,
		_w610_,
		_w715_
	);
	LUT2 #(
		.INIT('h1)
	) name580 (
		_w662_,
		_w714_,
		_w716_
	);
	LUT2 #(
		.INIT('h8)
	) name581 (
		_w715_,
		_w716_,
		_w717_
	);
	LUT2 #(
		.INIT('h1)
	) name582 (
		\shift[6] ,
		_w717_,
		_w718_
	);
	LUT2 #(
		.INIT('h2)
	) name583 (
		\a[65] ,
		\shift[0] ,
		_w719_
	);
	LUT2 #(
		.INIT('h1)
	) name584 (
		\shift[1] ,
		_w719_,
		_w720_
	);
	LUT2 #(
		.INIT('h8)
	) name585 (
		\a[62] ,
		\shift[0] ,
		_w721_
	);
	LUT2 #(
		.INIT('h2)
	) name586 (
		\shift[1] ,
		_w721_,
		_w722_
	);
	LUT2 #(
		.INIT('h1)
	) name587 (
		_w720_,
		_w722_,
		_w723_
	);
	LUT2 #(
		.INIT('h2)
	) name588 (
		\a[63] ,
		\shift[0] ,
		_w724_
	);
	LUT2 #(
		.INIT('h8)
	) name589 (
		\shift[1] ,
		_w724_,
		_w725_
	);
	LUT2 #(
		.INIT('h8)
	) name590 (
		\a[64] ,
		\shift[0] ,
		_w726_
	);
	LUT2 #(
		.INIT('h4)
	) name591 (
		\shift[1] ,
		_w726_,
		_w727_
	);
	LUT2 #(
		.INIT('h1)
	) name592 (
		_w725_,
		_w727_,
		_w728_
	);
	LUT2 #(
		.INIT('h4)
	) name593 (
		_w723_,
		_w728_,
		_w729_
	);
	LUT2 #(
		.INIT('h2)
	) name594 (
		_w136_,
		_w729_,
		_w730_
	);
	LUT2 #(
		.INIT('h2)
	) name595 (
		\a[61] ,
		\shift[0] ,
		_w731_
	);
	LUT2 #(
		.INIT('h1)
	) name596 (
		\shift[1] ,
		_w731_,
		_w732_
	);
	LUT2 #(
		.INIT('h8)
	) name597 (
		\a[58] ,
		\shift[0] ,
		_w733_
	);
	LUT2 #(
		.INIT('h2)
	) name598 (
		\shift[1] ,
		_w733_,
		_w734_
	);
	LUT2 #(
		.INIT('h1)
	) name599 (
		_w732_,
		_w734_,
		_w735_
	);
	LUT2 #(
		.INIT('h2)
	) name600 (
		\a[59] ,
		\shift[0] ,
		_w736_
	);
	LUT2 #(
		.INIT('h8)
	) name601 (
		\shift[1] ,
		_w736_,
		_w737_
	);
	LUT2 #(
		.INIT('h8)
	) name602 (
		\a[60] ,
		\shift[0] ,
		_w738_
	);
	LUT2 #(
		.INIT('h4)
	) name603 (
		\shift[1] ,
		_w738_,
		_w739_
	);
	LUT2 #(
		.INIT('h1)
	) name604 (
		_w737_,
		_w739_,
		_w740_
	);
	LUT2 #(
		.INIT('h4)
	) name605 (
		_w735_,
		_w740_,
		_w741_
	);
	LUT2 #(
		.INIT('h2)
	) name606 (
		_w147_,
		_w741_,
		_w742_
	);
	LUT2 #(
		.INIT('h2)
	) name607 (
		\a[53] ,
		\shift[0] ,
		_w743_
	);
	LUT2 #(
		.INIT('h1)
	) name608 (
		\shift[1] ,
		_w743_,
		_w744_
	);
	LUT2 #(
		.INIT('h8)
	) name609 (
		\a[50] ,
		\shift[0] ,
		_w745_
	);
	LUT2 #(
		.INIT('h2)
	) name610 (
		\shift[1] ,
		_w745_,
		_w746_
	);
	LUT2 #(
		.INIT('h1)
	) name611 (
		_w744_,
		_w746_,
		_w747_
	);
	LUT2 #(
		.INIT('h2)
	) name612 (
		\a[51] ,
		\shift[0] ,
		_w748_
	);
	LUT2 #(
		.INIT('h8)
	) name613 (
		\shift[1] ,
		_w748_,
		_w749_
	);
	LUT2 #(
		.INIT('h8)
	) name614 (
		\a[52] ,
		\shift[0] ,
		_w750_
	);
	LUT2 #(
		.INIT('h4)
	) name615 (
		\shift[1] ,
		_w750_,
		_w751_
	);
	LUT2 #(
		.INIT('h1)
	) name616 (
		_w749_,
		_w751_,
		_w752_
	);
	LUT2 #(
		.INIT('h4)
	) name617 (
		_w747_,
		_w752_,
		_w753_
	);
	LUT2 #(
		.INIT('h2)
	) name618 (
		_w158_,
		_w753_,
		_w754_
	);
	LUT2 #(
		.INIT('h2)
	) name619 (
		\a[57] ,
		\shift[0] ,
		_w755_
	);
	LUT2 #(
		.INIT('h1)
	) name620 (
		\shift[1] ,
		_w755_,
		_w756_
	);
	LUT2 #(
		.INIT('h8)
	) name621 (
		\a[54] ,
		\shift[0] ,
		_w757_
	);
	LUT2 #(
		.INIT('h2)
	) name622 (
		\shift[1] ,
		_w757_,
		_w758_
	);
	LUT2 #(
		.INIT('h1)
	) name623 (
		_w756_,
		_w758_,
		_w759_
	);
	LUT2 #(
		.INIT('h2)
	) name624 (
		\a[55] ,
		\shift[0] ,
		_w760_
	);
	LUT2 #(
		.INIT('h8)
	) name625 (
		\shift[1] ,
		_w760_,
		_w761_
	);
	LUT2 #(
		.INIT('h8)
	) name626 (
		\a[56] ,
		\shift[0] ,
		_w762_
	);
	LUT2 #(
		.INIT('h4)
	) name627 (
		\shift[1] ,
		_w762_,
		_w763_
	);
	LUT2 #(
		.INIT('h1)
	) name628 (
		_w761_,
		_w763_,
		_w764_
	);
	LUT2 #(
		.INIT('h4)
	) name629 (
		_w759_,
		_w764_,
		_w765_
	);
	LUT2 #(
		.INIT('h2)
	) name630 (
		_w169_,
		_w765_,
		_w766_
	);
	LUT2 #(
		.INIT('h1)
	) name631 (
		_w730_,
		_w742_,
		_w767_
	);
	LUT2 #(
		.INIT('h1)
	) name632 (
		_w754_,
		_w766_,
		_w768_
	);
	LUT2 #(
		.INIT('h8)
	) name633 (
		_w767_,
		_w768_,
		_w769_
	);
	LUT2 #(
		.INIT('h2)
	) name634 (
		_w273_,
		_w769_,
		_w770_
	);
	LUT2 #(
		.INIT('h2)
	) name635 (
		\a[17] ,
		\shift[0] ,
		_w771_
	);
	LUT2 #(
		.INIT('h1)
	) name636 (
		\shift[1] ,
		_w771_,
		_w772_
	);
	LUT2 #(
		.INIT('h8)
	) name637 (
		\a[14] ,
		\shift[0] ,
		_w773_
	);
	LUT2 #(
		.INIT('h2)
	) name638 (
		\shift[1] ,
		_w773_,
		_w774_
	);
	LUT2 #(
		.INIT('h1)
	) name639 (
		_w772_,
		_w774_,
		_w775_
	);
	LUT2 #(
		.INIT('h2)
	) name640 (
		\a[15] ,
		\shift[0] ,
		_w776_
	);
	LUT2 #(
		.INIT('h8)
	) name641 (
		\shift[1] ,
		_w776_,
		_w777_
	);
	LUT2 #(
		.INIT('h8)
	) name642 (
		\a[16] ,
		\shift[0] ,
		_w778_
	);
	LUT2 #(
		.INIT('h4)
	) name643 (
		\shift[1] ,
		_w778_,
		_w779_
	);
	LUT2 #(
		.INIT('h1)
	) name644 (
		_w777_,
		_w779_,
		_w780_
	);
	LUT2 #(
		.INIT('h4)
	) name645 (
		_w775_,
		_w780_,
		_w781_
	);
	LUT2 #(
		.INIT('h2)
	) name646 (
		_w136_,
		_w781_,
		_w782_
	);
	LUT2 #(
		.INIT('h2)
	) name647 (
		\a[13] ,
		\shift[0] ,
		_w783_
	);
	LUT2 #(
		.INIT('h1)
	) name648 (
		\shift[1] ,
		_w783_,
		_w784_
	);
	LUT2 #(
		.INIT('h8)
	) name649 (
		\a[10] ,
		\shift[0] ,
		_w785_
	);
	LUT2 #(
		.INIT('h2)
	) name650 (
		\shift[1] ,
		_w785_,
		_w786_
	);
	LUT2 #(
		.INIT('h1)
	) name651 (
		_w784_,
		_w786_,
		_w787_
	);
	LUT2 #(
		.INIT('h2)
	) name652 (
		\a[11] ,
		\shift[0] ,
		_w788_
	);
	LUT2 #(
		.INIT('h8)
	) name653 (
		\shift[1] ,
		_w788_,
		_w789_
	);
	LUT2 #(
		.INIT('h8)
	) name654 (
		\a[12] ,
		\shift[0] ,
		_w790_
	);
	LUT2 #(
		.INIT('h4)
	) name655 (
		\shift[1] ,
		_w790_,
		_w791_
	);
	LUT2 #(
		.INIT('h1)
	) name656 (
		_w789_,
		_w791_,
		_w792_
	);
	LUT2 #(
		.INIT('h4)
	) name657 (
		_w787_,
		_w792_,
		_w793_
	);
	LUT2 #(
		.INIT('h2)
	) name658 (
		_w147_,
		_w793_,
		_w794_
	);
	LUT2 #(
		.INIT('h2)
	) name659 (
		\a[5] ,
		\shift[0] ,
		_w795_
	);
	LUT2 #(
		.INIT('h1)
	) name660 (
		\shift[1] ,
		_w795_,
		_w796_
	);
	LUT2 #(
		.INIT('h8)
	) name661 (
		\a[2] ,
		\shift[0] ,
		_w797_
	);
	LUT2 #(
		.INIT('h2)
	) name662 (
		\shift[1] ,
		_w797_,
		_w798_
	);
	LUT2 #(
		.INIT('h1)
	) name663 (
		_w796_,
		_w798_,
		_w799_
	);
	LUT2 #(
		.INIT('h2)
	) name664 (
		\a[3] ,
		\shift[0] ,
		_w800_
	);
	LUT2 #(
		.INIT('h8)
	) name665 (
		\shift[1] ,
		_w800_,
		_w801_
	);
	LUT2 #(
		.INIT('h8)
	) name666 (
		\a[4] ,
		\shift[0] ,
		_w802_
	);
	LUT2 #(
		.INIT('h4)
	) name667 (
		\shift[1] ,
		_w802_,
		_w803_
	);
	LUT2 #(
		.INIT('h1)
	) name668 (
		_w801_,
		_w803_,
		_w804_
	);
	LUT2 #(
		.INIT('h4)
	) name669 (
		_w799_,
		_w804_,
		_w805_
	);
	LUT2 #(
		.INIT('h2)
	) name670 (
		_w158_,
		_w805_,
		_w806_
	);
	LUT2 #(
		.INIT('h2)
	) name671 (
		\a[9] ,
		\shift[0] ,
		_w807_
	);
	LUT2 #(
		.INIT('h1)
	) name672 (
		\shift[1] ,
		_w807_,
		_w808_
	);
	LUT2 #(
		.INIT('h8)
	) name673 (
		\a[6] ,
		\shift[0] ,
		_w809_
	);
	LUT2 #(
		.INIT('h2)
	) name674 (
		\shift[1] ,
		_w809_,
		_w810_
	);
	LUT2 #(
		.INIT('h1)
	) name675 (
		_w808_,
		_w810_,
		_w811_
	);
	LUT2 #(
		.INIT('h2)
	) name676 (
		\a[7] ,
		\shift[0] ,
		_w812_
	);
	LUT2 #(
		.INIT('h8)
	) name677 (
		\shift[1] ,
		_w812_,
		_w813_
	);
	LUT2 #(
		.INIT('h8)
	) name678 (
		\a[8] ,
		\shift[0] ,
		_w814_
	);
	LUT2 #(
		.INIT('h4)
	) name679 (
		\shift[1] ,
		_w814_,
		_w815_
	);
	LUT2 #(
		.INIT('h1)
	) name680 (
		_w813_,
		_w815_,
		_w816_
	);
	LUT2 #(
		.INIT('h4)
	) name681 (
		_w811_,
		_w816_,
		_w817_
	);
	LUT2 #(
		.INIT('h2)
	) name682 (
		_w169_,
		_w817_,
		_w818_
	);
	LUT2 #(
		.INIT('h1)
	) name683 (
		_w782_,
		_w794_,
		_w819_
	);
	LUT2 #(
		.INIT('h1)
	) name684 (
		_w806_,
		_w818_,
		_w820_
	);
	LUT2 #(
		.INIT('h8)
	) name685 (
		_w819_,
		_w820_,
		_w821_
	);
	LUT2 #(
		.INIT('h2)
	) name686 (
		_w183_,
		_w821_,
		_w822_
	);
	LUT2 #(
		.INIT('h2)
	) name687 (
		\a[49] ,
		\shift[0] ,
		_w823_
	);
	LUT2 #(
		.INIT('h1)
	) name688 (
		\shift[1] ,
		_w823_,
		_w824_
	);
	LUT2 #(
		.INIT('h8)
	) name689 (
		\a[46] ,
		\shift[0] ,
		_w825_
	);
	LUT2 #(
		.INIT('h2)
	) name690 (
		\shift[1] ,
		_w825_,
		_w826_
	);
	LUT2 #(
		.INIT('h1)
	) name691 (
		_w824_,
		_w826_,
		_w827_
	);
	LUT2 #(
		.INIT('h2)
	) name692 (
		\a[47] ,
		\shift[0] ,
		_w828_
	);
	LUT2 #(
		.INIT('h8)
	) name693 (
		\shift[1] ,
		_w828_,
		_w829_
	);
	LUT2 #(
		.INIT('h8)
	) name694 (
		\a[48] ,
		\shift[0] ,
		_w830_
	);
	LUT2 #(
		.INIT('h4)
	) name695 (
		\shift[1] ,
		_w830_,
		_w831_
	);
	LUT2 #(
		.INIT('h1)
	) name696 (
		_w829_,
		_w831_,
		_w832_
	);
	LUT2 #(
		.INIT('h4)
	) name697 (
		_w827_,
		_w832_,
		_w833_
	);
	LUT2 #(
		.INIT('h2)
	) name698 (
		_w136_,
		_w833_,
		_w834_
	);
	LUT2 #(
		.INIT('h8)
	) name699 (
		\a[42] ,
		\shift[0] ,
		_w835_
	);
	LUT2 #(
		.INIT('h2)
	) name700 (
		\a[43] ,
		\shift[0] ,
		_w836_
	);
	LUT2 #(
		.INIT('h1)
	) name701 (
		_w835_,
		_w836_,
		_w837_
	);
	LUT2 #(
		.INIT('h2)
	) name702 (
		\shift[1] ,
		_w837_,
		_w838_
	);
	LUT2 #(
		.INIT('h2)
	) name703 (
		\a[45] ,
		\shift[0] ,
		_w839_
	);
	LUT2 #(
		.INIT('h8)
	) name704 (
		\a[44] ,
		\shift[0] ,
		_w840_
	);
	LUT2 #(
		.INIT('h1)
	) name705 (
		_w839_,
		_w840_,
		_w841_
	);
	LUT2 #(
		.INIT('h1)
	) name706 (
		\shift[1] ,
		_w841_,
		_w842_
	);
	LUT2 #(
		.INIT('h1)
	) name707 (
		_w838_,
		_w842_,
		_w843_
	);
	LUT2 #(
		.INIT('h2)
	) name708 (
		_w147_,
		_w843_,
		_w844_
	);
	LUT2 #(
		.INIT('h2)
	) name709 (
		\a[37] ,
		\shift[0] ,
		_w845_
	);
	LUT2 #(
		.INIT('h1)
	) name710 (
		\shift[1] ,
		_w845_,
		_w846_
	);
	LUT2 #(
		.INIT('h8)
	) name711 (
		\a[34] ,
		\shift[0] ,
		_w847_
	);
	LUT2 #(
		.INIT('h2)
	) name712 (
		\shift[1] ,
		_w847_,
		_w848_
	);
	LUT2 #(
		.INIT('h1)
	) name713 (
		_w846_,
		_w848_,
		_w849_
	);
	LUT2 #(
		.INIT('h2)
	) name714 (
		\a[35] ,
		\shift[0] ,
		_w850_
	);
	LUT2 #(
		.INIT('h8)
	) name715 (
		\shift[1] ,
		_w850_,
		_w851_
	);
	LUT2 #(
		.INIT('h8)
	) name716 (
		\a[36] ,
		\shift[0] ,
		_w852_
	);
	LUT2 #(
		.INIT('h4)
	) name717 (
		\shift[1] ,
		_w852_,
		_w853_
	);
	LUT2 #(
		.INIT('h1)
	) name718 (
		_w851_,
		_w853_,
		_w854_
	);
	LUT2 #(
		.INIT('h4)
	) name719 (
		_w849_,
		_w854_,
		_w855_
	);
	LUT2 #(
		.INIT('h2)
	) name720 (
		_w158_,
		_w855_,
		_w856_
	);
	LUT2 #(
		.INIT('h2)
	) name721 (
		\a[41] ,
		\shift[0] ,
		_w857_
	);
	LUT2 #(
		.INIT('h8)
	) name722 (
		\a[40] ,
		\shift[0] ,
		_w858_
	);
	LUT2 #(
		.INIT('h1)
	) name723 (
		_w857_,
		_w858_,
		_w859_
	);
	LUT2 #(
		.INIT('h1)
	) name724 (
		\shift[1] ,
		_w859_,
		_w860_
	);
	LUT2 #(
		.INIT('h2)
	) name725 (
		\a[39] ,
		\shift[0] ,
		_w861_
	);
	LUT2 #(
		.INIT('h8)
	) name726 (
		\a[38] ,
		\shift[0] ,
		_w862_
	);
	LUT2 #(
		.INIT('h1)
	) name727 (
		_w861_,
		_w862_,
		_w863_
	);
	LUT2 #(
		.INIT('h2)
	) name728 (
		\shift[1] ,
		_w863_,
		_w864_
	);
	LUT2 #(
		.INIT('h1)
	) name729 (
		_w860_,
		_w864_,
		_w865_
	);
	LUT2 #(
		.INIT('h2)
	) name730 (
		_w169_,
		_w865_,
		_w866_
	);
	LUT2 #(
		.INIT('h1)
	) name731 (
		_w834_,
		_w844_,
		_w867_
	);
	LUT2 #(
		.INIT('h1)
	) name732 (
		_w856_,
		_w866_,
		_w868_
	);
	LUT2 #(
		.INIT('h8)
	) name733 (
		_w867_,
		_w868_,
		_w869_
	);
	LUT2 #(
		.INIT('h2)
	) name734 (
		_w318_,
		_w869_,
		_w870_
	);
	LUT2 #(
		.INIT('h2)
	) name735 (
		\a[33] ,
		\shift[0] ,
		_w871_
	);
	LUT2 #(
		.INIT('h1)
	) name736 (
		\shift[1] ,
		_w871_,
		_w872_
	);
	LUT2 #(
		.INIT('h8)
	) name737 (
		\a[30] ,
		\shift[0] ,
		_w873_
	);
	LUT2 #(
		.INIT('h2)
	) name738 (
		\shift[1] ,
		_w873_,
		_w874_
	);
	LUT2 #(
		.INIT('h1)
	) name739 (
		_w872_,
		_w874_,
		_w875_
	);
	LUT2 #(
		.INIT('h2)
	) name740 (
		\a[31] ,
		\shift[0] ,
		_w876_
	);
	LUT2 #(
		.INIT('h8)
	) name741 (
		\shift[1] ,
		_w876_,
		_w877_
	);
	LUT2 #(
		.INIT('h8)
	) name742 (
		\a[32] ,
		\shift[0] ,
		_w878_
	);
	LUT2 #(
		.INIT('h4)
	) name743 (
		\shift[1] ,
		_w878_,
		_w879_
	);
	LUT2 #(
		.INIT('h1)
	) name744 (
		_w877_,
		_w879_,
		_w880_
	);
	LUT2 #(
		.INIT('h4)
	) name745 (
		_w875_,
		_w880_,
		_w881_
	);
	LUT2 #(
		.INIT('h2)
	) name746 (
		_w136_,
		_w881_,
		_w882_
	);
	LUT2 #(
		.INIT('h2)
	) name747 (
		\a[29] ,
		\shift[0] ,
		_w883_
	);
	LUT2 #(
		.INIT('h1)
	) name748 (
		\shift[1] ,
		_w883_,
		_w884_
	);
	LUT2 #(
		.INIT('h8)
	) name749 (
		\a[26] ,
		\shift[0] ,
		_w885_
	);
	LUT2 #(
		.INIT('h2)
	) name750 (
		\shift[1] ,
		_w885_,
		_w886_
	);
	LUT2 #(
		.INIT('h1)
	) name751 (
		_w884_,
		_w886_,
		_w887_
	);
	LUT2 #(
		.INIT('h2)
	) name752 (
		\a[27] ,
		\shift[0] ,
		_w888_
	);
	LUT2 #(
		.INIT('h8)
	) name753 (
		\shift[1] ,
		_w888_,
		_w889_
	);
	LUT2 #(
		.INIT('h8)
	) name754 (
		\a[28] ,
		\shift[0] ,
		_w890_
	);
	LUT2 #(
		.INIT('h4)
	) name755 (
		\shift[1] ,
		_w890_,
		_w891_
	);
	LUT2 #(
		.INIT('h1)
	) name756 (
		_w889_,
		_w891_,
		_w892_
	);
	LUT2 #(
		.INIT('h4)
	) name757 (
		_w887_,
		_w892_,
		_w893_
	);
	LUT2 #(
		.INIT('h2)
	) name758 (
		_w147_,
		_w893_,
		_w894_
	);
	LUT2 #(
		.INIT('h2)
	) name759 (
		\a[21] ,
		\shift[0] ,
		_w895_
	);
	LUT2 #(
		.INIT('h1)
	) name760 (
		\shift[1] ,
		_w895_,
		_w896_
	);
	LUT2 #(
		.INIT('h8)
	) name761 (
		\a[18] ,
		\shift[0] ,
		_w897_
	);
	LUT2 #(
		.INIT('h2)
	) name762 (
		\shift[1] ,
		_w897_,
		_w898_
	);
	LUT2 #(
		.INIT('h1)
	) name763 (
		_w896_,
		_w898_,
		_w899_
	);
	LUT2 #(
		.INIT('h2)
	) name764 (
		\a[19] ,
		\shift[0] ,
		_w900_
	);
	LUT2 #(
		.INIT('h8)
	) name765 (
		\shift[1] ,
		_w900_,
		_w901_
	);
	LUT2 #(
		.INIT('h8)
	) name766 (
		\a[20] ,
		\shift[0] ,
		_w902_
	);
	LUT2 #(
		.INIT('h4)
	) name767 (
		\shift[1] ,
		_w902_,
		_w903_
	);
	LUT2 #(
		.INIT('h1)
	) name768 (
		_w901_,
		_w903_,
		_w904_
	);
	LUT2 #(
		.INIT('h4)
	) name769 (
		_w899_,
		_w904_,
		_w905_
	);
	LUT2 #(
		.INIT('h2)
	) name770 (
		_w158_,
		_w905_,
		_w906_
	);
	LUT2 #(
		.INIT('h2)
	) name771 (
		\a[25] ,
		\shift[0] ,
		_w907_
	);
	LUT2 #(
		.INIT('h1)
	) name772 (
		\shift[1] ,
		_w907_,
		_w908_
	);
	LUT2 #(
		.INIT('h8)
	) name773 (
		\a[22] ,
		\shift[0] ,
		_w909_
	);
	LUT2 #(
		.INIT('h2)
	) name774 (
		\shift[1] ,
		_w909_,
		_w910_
	);
	LUT2 #(
		.INIT('h1)
	) name775 (
		_w908_,
		_w910_,
		_w911_
	);
	LUT2 #(
		.INIT('h2)
	) name776 (
		\a[23] ,
		\shift[0] ,
		_w912_
	);
	LUT2 #(
		.INIT('h8)
	) name777 (
		\shift[1] ,
		_w912_,
		_w913_
	);
	LUT2 #(
		.INIT('h8)
	) name778 (
		\a[24] ,
		\shift[0] ,
		_w914_
	);
	LUT2 #(
		.INIT('h4)
	) name779 (
		\shift[1] ,
		_w914_,
		_w915_
	);
	LUT2 #(
		.INIT('h1)
	) name780 (
		_w913_,
		_w915_,
		_w916_
	);
	LUT2 #(
		.INIT('h4)
	) name781 (
		_w911_,
		_w916_,
		_w917_
	);
	LUT2 #(
		.INIT('h2)
	) name782 (
		_w169_,
		_w917_,
		_w918_
	);
	LUT2 #(
		.INIT('h1)
	) name783 (
		_w882_,
		_w894_,
		_w919_
	);
	LUT2 #(
		.INIT('h1)
	) name784 (
		_w906_,
		_w918_,
		_w920_
	);
	LUT2 #(
		.INIT('h8)
	) name785 (
		_w919_,
		_w920_,
		_w921_
	);
	LUT2 #(
		.INIT('h2)
	) name786 (
		_w228_,
		_w921_,
		_w922_
	);
	LUT2 #(
		.INIT('h1)
	) name787 (
		_w770_,
		_w822_,
		_w923_
	);
	LUT2 #(
		.INIT('h1)
	) name788 (
		_w870_,
		_w922_,
		_w924_
	);
	LUT2 #(
		.INIT('h8)
	) name789 (
		_w923_,
		_w924_,
		_w925_
	);
	LUT2 #(
		.INIT('h2)
	) name790 (
		\shift[6] ,
		_w925_,
		_w926_
	);
	LUT2 #(
		.INIT('h1)
	) name791 (
		_w718_,
		_w926_,
		_w927_
	);
	LUT2 #(
		.INIT('h2)
	) name792 (
		\shift[1] ,
		_w143_,
		_w928_
	);
	LUT2 #(
		.INIT('h1)
	) name793 (
		\shift[1] ,
		_w207_,
		_w929_
	);
	LUT2 #(
		.INIT('h1)
	) name794 (
		_w928_,
		_w929_,
		_w930_
	);
	LUT2 #(
		.INIT('h2)
	) name795 (
		_w136_,
		_w930_,
		_w931_
	);
	LUT2 #(
		.INIT('h2)
	) name796 (
		\shift[1] ,
		_w154_,
		_w932_
	);
	LUT2 #(
		.INIT('h1)
	) name797 (
		\shift[1] ,
		_w139_,
		_w933_
	);
	LUT2 #(
		.INIT('h1)
	) name798 (
		_w932_,
		_w933_,
		_w934_
	);
	LUT2 #(
		.INIT('h2)
	) name799 (
		_w147_,
		_w934_,
		_w935_
	);
	LUT2 #(
		.INIT('h2)
	) name800 (
		\shift[1] ,
		_w165_,
		_w936_
	);
	LUT2 #(
		.INIT('h1)
	) name801 (
		\shift[1] ,
		_w172_,
		_w937_
	);
	LUT2 #(
		.INIT('h1)
	) name802 (
		_w936_,
		_w937_,
		_w938_
	);
	LUT2 #(
		.INIT('h2)
	) name803 (
		_w158_,
		_w938_,
		_w939_
	);
	LUT2 #(
		.INIT('h2)
	) name804 (
		\shift[1] ,
		_w176_,
		_w940_
	);
	LUT2 #(
		.INIT('h1)
	) name805 (
		\shift[1] ,
		_w150_,
		_w941_
	);
	LUT2 #(
		.INIT('h1)
	) name806 (
		_w940_,
		_w941_,
		_w942_
	);
	LUT2 #(
		.INIT('h2)
	) name807 (
		_w169_,
		_w942_,
		_w943_
	);
	LUT2 #(
		.INIT('h1)
	) name808 (
		_w931_,
		_w935_,
		_w944_
	);
	LUT2 #(
		.INIT('h1)
	) name809 (
		_w939_,
		_w943_,
		_w945_
	);
	LUT2 #(
		.INIT('h8)
	) name810 (
		_w944_,
		_w945_,
		_w946_
	);
	LUT2 #(
		.INIT('h2)
	) name811 (
		_w183_,
		_w946_,
		_w947_
	);
	LUT2 #(
		.INIT('h2)
	) name812 (
		\shift[1] ,
		_w191_,
		_w948_
	);
	LUT2 #(
		.INIT('h1)
	) name813 (
		\shift[1] ,
		_w297_,
		_w949_
	);
	LUT2 #(
		.INIT('h1)
	) name814 (
		_w948_,
		_w949_,
		_w950_
	);
	LUT2 #(
		.INIT('h2)
	) name815 (
		_w136_,
		_w950_,
		_w951_
	);
	LUT2 #(
		.INIT('h2)
	) name816 (
		\shift[1] ,
		_w201_,
		_w952_
	);
	LUT2 #(
		.INIT('h1)
	) name817 (
		\shift[1] ,
		_w187_,
		_w953_
	);
	LUT2 #(
		.INIT('h1)
	) name818 (
		_w952_,
		_w953_,
		_w954_
	);
	LUT2 #(
		.INIT('h2)
	) name819 (
		_w147_,
		_w954_,
		_w955_
	);
	LUT2 #(
		.INIT('h2)
	) name820 (
		\shift[1] ,
		_w211_,
		_w956_
	);
	LUT2 #(
		.INIT('h1)
	) name821 (
		\shift[1] ,
		_w217_,
		_w957_
	);
	LUT2 #(
		.INIT('h1)
	) name822 (
		_w956_,
		_w957_,
		_w958_
	);
	LUT2 #(
		.INIT('h2)
	) name823 (
		_w158_,
		_w958_,
		_w959_
	);
	LUT2 #(
		.INIT('h2)
	) name824 (
		\shift[1] ,
		_w221_,
		_w960_
	);
	LUT2 #(
		.INIT('h1)
	) name825 (
		\shift[1] ,
		_w197_,
		_w961_
	);
	LUT2 #(
		.INIT('h1)
	) name826 (
		_w960_,
		_w961_,
		_w962_
	);
	LUT2 #(
		.INIT('h2)
	) name827 (
		_w169_,
		_w962_,
		_w963_
	);
	LUT2 #(
		.INIT('h1)
	) name828 (
		_w951_,
		_w955_,
		_w964_
	);
	LUT2 #(
		.INIT('h1)
	) name829 (
		_w959_,
		_w963_,
		_w965_
	);
	LUT2 #(
		.INIT('h8)
	) name830 (
		_w964_,
		_w965_,
		_w966_
	);
	LUT2 #(
		.INIT('h2)
	) name831 (
		_w228_,
		_w966_,
		_w967_
	);
	LUT2 #(
		.INIT('h2)
	) name832 (
		\shift[1] ,
		_w236_,
		_w968_
	);
	LUT2 #(
		.INIT('h1)
	) name833 (
		\shift[1] ,
		_w346_,
		_w969_
	);
	LUT2 #(
		.INIT('h1)
	) name834 (
		_w968_,
		_w969_,
		_w970_
	);
	LUT2 #(
		.INIT('h2)
	) name835 (
		_w136_,
		_w970_,
		_w971_
	);
	LUT2 #(
		.INIT('h2)
	) name836 (
		\shift[1] ,
		_w246_,
		_w972_
	);
	LUT2 #(
		.INIT('h1)
	) name837 (
		\shift[1] ,
		_w232_,
		_w973_
	);
	LUT2 #(
		.INIT('h1)
	) name838 (
		_w972_,
		_w973_,
		_w974_
	);
	LUT2 #(
		.INIT('h2)
	) name839 (
		_w147_,
		_w974_,
		_w975_
	);
	LUT2 #(
		.INIT('h2)
	) name840 (
		\shift[1] ,
		_w256_,
		_w976_
	);
	LUT2 #(
		.INIT('h1)
	) name841 (
		\shift[1] ,
		_w262_,
		_w977_
	);
	LUT2 #(
		.INIT('h1)
	) name842 (
		_w976_,
		_w977_,
		_w978_
	);
	LUT2 #(
		.INIT('h2)
	) name843 (
		_w158_,
		_w978_,
		_w979_
	);
	LUT2 #(
		.INIT('h2)
	) name844 (
		\shift[1] ,
		_w266_,
		_w980_
	);
	LUT2 #(
		.INIT('h1)
	) name845 (
		\shift[1] ,
		_w242_,
		_w981_
	);
	LUT2 #(
		.INIT('h1)
	) name846 (
		_w980_,
		_w981_,
		_w982_
	);
	LUT2 #(
		.INIT('h2)
	) name847 (
		_w169_,
		_w982_,
		_w983_
	);
	LUT2 #(
		.INIT('h1)
	) name848 (
		_w971_,
		_w975_,
		_w984_
	);
	LUT2 #(
		.INIT('h1)
	) name849 (
		_w979_,
		_w983_,
		_w985_
	);
	LUT2 #(
		.INIT('h8)
	) name850 (
		_w984_,
		_w985_,
		_w986_
	);
	LUT2 #(
		.INIT('h2)
	) name851 (
		_w273_,
		_w986_,
		_w987_
	);
	LUT2 #(
		.INIT('h2)
	) name852 (
		\shift[1] ,
		_w281_,
		_w988_
	);
	LUT2 #(
		.INIT('h1)
	) name853 (
		\shift[1] ,
		_w252_,
		_w989_
	);
	LUT2 #(
		.INIT('h1)
	) name854 (
		_w988_,
		_w989_,
		_w990_
	);
	LUT2 #(
		.INIT('h2)
	) name855 (
		_w136_,
		_w990_,
		_w991_
	);
	LUT2 #(
		.INIT('h2)
	) name856 (
		\shift[1] ,
		_w291_,
		_w992_
	);
	LUT2 #(
		.INIT('h1)
	) name857 (
		\shift[1] ,
		_w277_,
		_w993_
	);
	LUT2 #(
		.INIT('h1)
	) name858 (
		_w992_,
		_w993_,
		_w994_
	);
	LUT2 #(
		.INIT('h2)
	) name859 (
		_w147_,
		_w994_,
		_w995_
	);
	LUT2 #(
		.INIT('h2)
	) name860 (
		\shift[1] ,
		_w301_,
		_w996_
	);
	LUT2 #(
		.INIT('h1)
	) name861 (
		\shift[1] ,
		_w307_,
		_w997_
	);
	LUT2 #(
		.INIT('h1)
	) name862 (
		_w996_,
		_w997_,
		_w998_
	);
	LUT2 #(
		.INIT('h2)
	) name863 (
		_w158_,
		_w998_,
		_w999_
	);
	LUT2 #(
		.INIT('h2)
	) name864 (
		\shift[1] ,
		_w311_,
		_w1000_
	);
	LUT2 #(
		.INIT('h1)
	) name865 (
		\shift[1] ,
		_w287_,
		_w1001_
	);
	LUT2 #(
		.INIT('h1)
	) name866 (
		_w1000_,
		_w1001_,
		_w1002_
	);
	LUT2 #(
		.INIT('h2)
	) name867 (
		_w169_,
		_w1002_,
		_w1003_
	);
	LUT2 #(
		.INIT('h1)
	) name868 (
		_w991_,
		_w995_,
		_w1004_
	);
	LUT2 #(
		.INIT('h1)
	) name869 (
		_w999_,
		_w1003_,
		_w1005_
	);
	LUT2 #(
		.INIT('h8)
	) name870 (
		_w1004_,
		_w1005_,
		_w1006_
	);
	LUT2 #(
		.INIT('h2)
	) name871 (
		_w318_,
		_w1006_,
		_w1007_
	);
	LUT2 #(
		.INIT('h1)
	) name872 (
		_w947_,
		_w967_,
		_w1008_
	);
	LUT2 #(
		.INIT('h1)
	) name873 (
		_w987_,
		_w1007_,
		_w1009_
	);
	LUT2 #(
		.INIT('h8)
	) name874 (
		_w1008_,
		_w1009_,
		_w1010_
	);
	LUT2 #(
		.INIT('h1)
	) name875 (
		\shift[6] ,
		_w1010_,
		_w1011_
	);
	LUT2 #(
		.INIT('h2)
	) name876 (
		\shift[1] ,
		_w418_,
		_w1012_
	);
	LUT2 #(
		.INIT('h1)
	) name877 (
		\shift[1] ,
		_w161_,
		_w1013_
	);
	LUT2 #(
		.INIT('h1)
	) name878 (
		_w1012_,
		_w1013_,
		_w1014_
	);
	LUT2 #(
		.INIT('h2)
	) name879 (
		_w136_,
		_w1014_,
		_w1015_
	);
	LUT2 #(
		.INIT('h2)
	) name880 (
		\shift[1] ,
		_w428_,
		_w1016_
	);
	LUT2 #(
		.INIT('h1)
	) name881 (
		\shift[1] ,
		_w414_,
		_w1017_
	);
	LUT2 #(
		.INIT('h1)
	) name882 (
		_w1016_,
		_w1017_,
		_w1018_
	);
	LUT2 #(
		.INIT('h2)
	) name883 (
		_w147_,
		_w1018_,
		_w1019_
	);
	LUT2 #(
		.INIT('h2)
	) name884 (
		\shift[1] ,
		_w438_,
		_w1020_
	);
	LUT2 #(
		.INIT('h1)
	) name885 (
		\shift[1] ,
		_w444_,
		_w1021_
	);
	LUT2 #(
		.INIT('h1)
	) name886 (
		_w1020_,
		_w1021_,
		_w1022_
	);
	LUT2 #(
		.INIT('h2)
	) name887 (
		_w158_,
		_w1022_,
		_w1023_
	);
	LUT2 #(
		.INIT('h2)
	) name888 (
		\shift[1] ,
		_w448_,
		_w1024_
	);
	LUT2 #(
		.INIT('h1)
	) name889 (
		\shift[1] ,
		_w424_,
		_w1025_
	);
	LUT2 #(
		.INIT('h1)
	) name890 (
		_w1024_,
		_w1025_,
		_w1026_
	);
	LUT2 #(
		.INIT('h2)
	) name891 (
		_w169_,
		_w1026_,
		_w1027_
	);
	LUT2 #(
		.INIT('h1)
	) name892 (
		_w1015_,
		_w1019_,
		_w1028_
	);
	LUT2 #(
		.INIT('h1)
	) name893 (
		_w1023_,
		_w1027_,
		_w1029_
	);
	LUT2 #(
		.INIT('h8)
	) name894 (
		_w1028_,
		_w1029_,
		_w1030_
	);
	LUT2 #(
		.INIT('h2)
	) name895 (
		_w273_,
		_w1030_,
		_w1031_
	);
	LUT2 #(
		.INIT('h2)
	) name896 (
		\shift[1] ,
		_w330_,
		_w1032_
	);
	LUT2 #(
		.INIT('h1)
	) name897 (
		\shift[1] ,
		_w390_,
		_w1033_
	);
	LUT2 #(
		.INIT('h1)
	) name898 (
		_w1032_,
		_w1033_,
		_w1034_
	);
	LUT2 #(
		.INIT('h2)
	) name899 (
		_w136_,
		_w1034_,
		_w1035_
	);
	LUT2 #(
		.INIT('h2)
	) name900 (
		\shift[1] ,
		_w340_,
		_w1036_
	);
	LUT2 #(
		.INIT('h1)
	) name901 (
		\shift[1] ,
		_w326_,
		_w1037_
	);
	LUT2 #(
		.INIT('h1)
	) name902 (
		_w1036_,
		_w1037_,
		_w1038_
	);
	LUT2 #(
		.INIT('h2)
	) name903 (
		_w147_,
		_w1038_,
		_w1039_
	);
	LUT2 #(
		.INIT('h2)
	) name904 (
		\shift[1] ,
		_w350_,
		_w1040_
	);
	LUT2 #(
		.INIT('h1)
	) name905 (
		\shift[1] ,
		_w356_,
		_w1041_
	);
	LUT2 #(
		.INIT('h1)
	) name906 (
		_w1040_,
		_w1041_,
		_w1042_
	);
	LUT2 #(
		.INIT('h2)
	) name907 (
		_w158_,
		_w1042_,
		_w1043_
	);
	LUT2 #(
		.INIT('h2)
	) name908 (
		\shift[1] ,
		_w360_,
		_w1044_
	);
	LUT2 #(
		.INIT('h1)
	) name909 (
		\shift[1] ,
		_w336_,
		_w1045_
	);
	LUT2 #(
		.INIT('h1)
	) name910 (
		_w1044_,
		_w1045_,
		_w1046_
	);
	LUT2 #(
		.INIT('h2)
	) name911 (
		_w169_,
		_w1046_,
		_w1047_
	);
	LUT2 #(
		.INIT('h1)
	) name912 (
		_w1035_,
		_w1039_,
		_w1048_
	);
	LUT2 #(
		.INIT('h1)
	) name913 (
		_w1043_,
		_w1047_,
		_w1049_
	);
	LUT2 #(
		.INIT('h8)
	) name914 (
		_w1048_,
		_w1049_,
		_w1050_
	);
	LUT2 #(
		.INIT('h2)
	) name915 (
		_w183_,
		_w1050_,
		_w1051_
	);
	LUT2 #(
		.INIT('h2)
	) name916 (
		\shift[1] ,
		_w462_,
		_w1052_
	);
	LUT2 #(
		.INIT('h1)
	) name917 (
		\shift[1] ,
		_w434_,
		_w1053_
	);
	LUT2 #(
		.INIT('h1)
	) name918 (
		_w1052_,
		_w1053_,
		_w1054_
	);
	LUT2 #(
		.INIT('h2)
	) name919 (
		_w136_,
		_w1054_,
		_w1055_
	);
	LUT2 #(
		.INIT('h2)
	) name920 (
		\shift[1] ,
		_w472_,
		_w1056_
	);
	LUT2 #(
		.INIT('h1)
	) name921 (
		\shift[1] ,
		_w458_,
		_w1057_
	);
	LUT2 #(
		.INIT('h1)
	) name922 (
		_w1056_,
		_w1057_,
		_w1058_
	);
	LUT2 #(
		.INIT('h2)
	) name923 (
		_w147_,
		_w1058_,
		_w1059_
	);
	LUT2 #(
		.INIT('h1)
	) name924 (
		_w488_,
		_w491_,
		_w1060_
	);
	LUT2 #(
		.INIT('h1)
	) name925 (
		\shift[1] ,
		_w1060_,
		_w1061_
	);
	LUT2 #(
		.INIT('h2)
	) name926 (
		\shift[1] ,
		_w482_,
		_w1062_
	);
	LUT2 #(
		.INIT('h1)
	) name927 (
		_w1061_,
		_w1062_,
		_w1063_
	);
	LUT2 #(
		.INIT('h2)
	) name928 (
		_w158_,
		_w1063_,
		_w1064_
	);
	LUT2 #(
		.INIT('h1)
	) name929 (
		\shift[1] ,
		_w468_,
		_w1065_
	);
	LUT2 #(
		.INIT('h1)
	) name930 (
		_w486_,
		_w493_,
		_w1066_
	);
	LUT2 #(
		.INIT('h2)
	) name931 (
		\shift[1] ,
		_w1066_,
		_w1067_
	);
	LUT2 #(
		.INIT('h1)
	) name932 (
		_w1065_,
		_w1067_,
		_w1068_
	);
	LUT2 #(
		.INIT('h2)
	) name933 (
		_w169_,
		_w1068_,
		_w1069_
	);
	LUT2 #(
		.INIT('h1)
	) name934 (
		_w1055_,
		_w1059_,
		_w1070_
	);
	LUT2 #(
		.INIT('h1)
	) name935 (
		_w1064_,
		_w1069_,
		_w1071_
	);
	LUT2 #(
		.INIT('h8)
	) name936 (
		_w1070_,
		_w1071_,
		_w1072_
	);
	LUT2 #(
		.INIT('h2)
	) name937 (
		_w318_,
		_w1072_,
		_w1073_
	);
	LUT2 #(
		.INIT('h2)
	) name938 (
		\shift[1] ,
		_w374_,
		_w1074_
	);
	LUT2 #(
		.INIT('h1)
	) name939 (
		\shift[1] ,
		_w478_,
		_w1075_
	);
	LUT2 #(
		.INIT('h1)
	) name940 (
		_w1074_,
		_w1075_,
		_w1076_
	);
	LUT2 #(
		.INIT('h2)
	) name941 (
		_w136_,
		_w1076_,
		_w1077_
	);
	LUT2 #(
		.INIT('h2)
	) name942 (
		\shift[1] ,
		_w384_,
		_w1078_
	);
	LUT2 #(
		.INIT('h1)
	) name943 (
		\shift[1] ,
		_w370_,
		_w1079_
	);
	LUT2 #(
		.INIT('h1)
	) name944 (
		_w1078_,
		_w1079_,
		_w1080_
	);
	LUT2 #(
		.INIT('h2)
	) name945 (
		_w147_,
		_w1080_,
		_w1081_
	);
	LUT2 #(
		.INIT('h2)
	) name946 (
		\shift[1] ,
		_w394_,
		_w1082_
	);
	LUT2 #(
		.INIT('h1)
	) name947 (
		\shift[1] ,
		_w400_,
		_w1083_
	);
	LUT2 #(
		.INIT('h1)
	) name948 (
		_w1082_,
		_w1083_,
		_w1084_
	);
	LUT2 #(
		.INIT('h2)
	) name949 (
		_w158_,
		_w1084_,
		_w1085_
	);
	LUT2 #(
		.INIT('h2)
	) name950 (
		\shift[1] ,
		_w404_,
		_w1086_
	);
	LUT2 #(
		.INIT('h1)
	) name951 (
		\shift[1] ,
		_w380_,
		_w1087_
	);
	LUT2 #(
		.INIT('h1)
	) name952 (
		_w1086_,
		_w1087_,
		_w1088_
	);
	LUT2 #(
		.INIT('h2)
	) name953 (
		_w169_,
		_w1088_,
		_w1089_
	);
	LUT2 #(
		.INIT('h1)
	) name954 (
		_w1077_,
		_w1081_,
		_w1090_
	);
	LUT2 #(
		.INIT('h1)
	) name955 (
		_w1085_,
		_w1089_,
		_w1091_
	);
	LUT2 #(
		.INIT('h8)
	) name956 (
		_w1090_,
		_w1091_,
		_w1092_
	);
	LUT2 #(
		.INIT('h2)
	) name957 (
		_w228_,
		_w1092_,
		_w1093_
	);
	LUT2 #(
		.INIT('h1)
	) name958 (
		_w1031_,
		_w1051_,
		_w1094_
	);
	LUT2 #(
		.INIT('h1)
	) name959 (
		_w1073_,
		_w1093_,
		_w1095_
	);
	LUT2 #(
		.INIT('h8)
	) name960 (
		_w1094_,
		_w1095_,
		_w1096_
	);
	LUT2 #(
		.INIT('h2)
	) name961 (
		\shift[6] ,
		_w1096_,
		_w1097_
	);
	LUT2 #(
		.INIT('h1)
	) name962 (
		_w1011_,
		_w1097_,
		_w1098_
	);
	LUT2 #(
		.INIT('h1)
	) name963 (
		\shift[1] ,
		_w637_,
		_w1099_
	);
	LUT2 #(
		.INIT('h2)
	) name964 (
		\shift[1] ,
		_w663_,
		_w1100_
	);
	LUT2 #(
		.INIT('h1)
	) name965 (
		_w1099_,
		_w1100_,
		_w1101_
	);
	LUT2 #(
		.INIT('h8)
	) name966 (
		\shift[1] ,
		_w670_,
		_w1102_
	);
	LUT2 #(
		.INIT('h4)
	) name967 (
		\shift[1] ,
		_w640_,
		_w1103_
	);
	LUT2 #(
		.INIT('h1)
	) name968 (
		_w1102_,
		_w1103_,
		_w1104_
	);
	LUT2 #(
		.INIT('h4)
	) name969 (
		_w1101_,
		_w1104_,
		_w1105_
	);
	LUT2 #(
		.INIT('h2)
	) name970 (
		_w136_,
		_w1105_,
		_w1106_
	);
	LUT2 #(
		.INIT('h1)
	) name971 (
		\shift[1] ,
		_w665_,
		_w1107_
	);
	LUT2 #(
		.INIT('h2)
	) name972 (
		\shift[1] ,
		_w675_,
		_w1108_
	);
	LUT2 #(
		.INIT('h1)
	) name973 (
		_w1107_,
		_w1108_,
		_w1109_
	);
	LUT2 #(
		.INIT('h8)
	) name974 (
		\shift[1] ,
		_w682_,
		_w1110_
	);
	LUT2 #(
		.INIT('h4)
	) name975 (
		\shift[1] ,
		_w668_,
		_w1111_
	);
	LUT2 #(
		.INIT('h1)
	) name976 (
		_w1110_,
		_w1111_,
		_w1112_
	);
	LUT2 #(
		.INIT('h4)
	) name977 (
		_w1109_,
		_w1112_,
		_w1113_
	);
	LUT2 #(
		.INIT('h2)
	) name978 (
		_w147_,
		_w1113_,
		_w1114_
	);
	LUT2 #(
		.INIT('h1)
	) name979 (
		\shift[1] ,
		_w701_,
		_w1115_
	);
	LUT2 #(
		.INIT('h2)
	) name980 (
		\shift[1] ,
		_w687_,
		_w1116_
	);
	LUT2 #(
		.INIT('h1)
	) name981 (
		_w1115_,
		_w1116_,
		_w1117_
	);
	LUT2 #(
		.INIT('h8)
	) name982 (
		\shift[1] ,
		_w694_,
		_w1118_
	);
	LUT2 #(
		.INIT('h4)
	) name983 (
		\shift[1] ,
		_w704_,
		_w1119_
	);
	LUT2 #(
		.INIT('h1)
	) name984 (
		_w1118_,
		_w1119_,
		_w1120_
	);
	LUT2 #(
		.INIT('h4)
	) name985 (
		_w1117_,
		_w1120_,
		_w1121_
	);
	LUT2 #(
		.INIT('h2)
	) name986 (
		_w158_,
		_w1121_,
		_w1122_
	);
	LUT2 #(
		.INIT('h1)
	) name987 (
		\shift[1] ,
		_w677_,
		_w1123_
	);
	LUT2 #(
		.INIT('h2)
	) name988 (
		\shift[1] ,
		_w699_,
		_w1124_
	);
	LUT2 #(
		.INIT('h1)
	) name989 (
		_w1123_,
		_w1124_,
		_w1125_
	);
	LUT2 #(
		.INIT('h8)
	) name990 (
		\shift[1] ,
		_w706_,
		_w1126_
	);
	LUT2 #(
		.INIT('h4)
	) name991 (
		\shift[1] ,
		_w680_,
		_w1127_
	);
	LUT2 #(
		.INIT('h1)
	) name992 (
		_w1126_,
		_w1127_,
		_w1128_
	);
	LUT2 #(
		.INIT('h4)
	) name993 (
		_w1125_,
		_w1128_,
		_w1129_
	);
	LUT2 #(
		.INIT('h2)
	) name994 (
		_w169_,
		_w1129_,
		_w1130_
	);
	LUT2 #(
		.INIT('h1)
	) name995 (
		_w1106_,
		_w1114_,
		_w1131_
	);
	LUT2 #(
		.INIT('h1)
	) name996 (
		_w1122_,
		_w1130_,
		_w1132_
	);
	LUT2 #(
		.INIT('h8)
	) name997 (
		_w1131_,
		_w1132_,
		_w1133_
	);
	LUT2 #(
		.INIT('h2)
	) name998 (
		_w318_,
		_w1133_,
		_w1134_
	);
	LUT2 #(
		.INIT('h1)
	) name999 (
		\shift[1] ,
		_w689_,
		_w1135_
	);
	LUT2 #(
		.INIT('h2)
	) name1000 (
		\shift[1] ,
		_w559_,
		_w1136_
	);
	LUT2 #(
		.INIT('h1)
	) name1001 (
		_w1135_,
		_w1136_,
		_w1137_
	);
	LUT2 #(
		.INIT('h8)
	) name1002 (
		\shift[1] ,
		_w566_,
		_w1138_
	);
	LUT2 #(
		.INIT('h4)
	) name1003 (
		\shift[1] ,
		_w692_,
		_w1139_
	);
	LUT2 #(
		.INIT('h1)
	) name1004 (
		_w1138_,
		_w1139_,
		_w1140_
	);
	LUT2 #(
		.INIT('h4)
	) name1005 (
		_w1137_,
		_w1140_,
		_w1141_
	);
	LUT2 #(
		.INIT('h2)
	) name1006 (
		_w136_,
		_w1141_,
		_w1142_
	);
	LUT2 #(
		.INIT('h1)
	) name1007 (
		\shift[1] ,
		_w561_,
		_w1143_
	);
	LUT2 #(
		.INIT('h2)
	) name1008 (
		\shift[1] ,
		_w571_,
		_w1144_
	);
	LUT2 #(
		.INIT('h1)
	) name1009 (
		_w1143_,
		_w1144_,
		_w1145_
	);
	LUT2 #(
		.INIT('h8)
	) name1010 (
		\shift[1] ,
		_w578_,
		_w1146_
	);
	LUT2 #(
		.INIT('h4)
	) name1011 (
		\shift[1] ,
		_w564_,
		_w1147_
	);
	LUT2 #(
		.INIT('h1)
	) name1012 (
		_w1146_,
		_w1147_,
		_w1148_
	);
	LUT2 #(
		.INIT('h4)
	) name1013 (
		_w1145_,
		_w1148_,
		_w1149_
	);
	LUT2 #(
		.INIT('h2)
	) name1014 (
		_w147_,
		_w1149_,
		_w1150_
	);
	LUT2 #(
		.INIT('h1)
	) name1015 (
		\shift[1] ,
		_w597_,
		_w1151_
	);
	LUT2 #(
		.INIT('h2)
	) name1016 (
		\shift[1] ,
		_w583_,
		_w1152_
	);
	LUT2 #(
		.INIT('h1)
	) name1017 (
		_w1151_,
		_w1152_,
		_w1153_
	);
	LUT2 #(
		.INIT('h8)
	) name1018 (
		\shift[1] ,
		_w590_,
		_w1154_
	);
	LUT2 #(
		.INIT('h4)
	) name1019 (
		\shift[1] ,
		_w600_,
		_w1155_
	);
	LUT2 #(
		.INIT('h1)
	) name1020 (
		_w1154_,
		_w1155_,
		_w1156_
	);
	LUT2 #(
		.INIT('h4)
	) name1021 (
		_w1153_,
		_w1156_,
		_w1157_
	);
	LUT2 #(
		.INIT('h2)
	) name1022 (
		_w158_,
		_w1157_,
		_w1158_
	);
	LUT2 #(
		.INIT('h1)
	) name1023 (
		\shift[1] ,
		_w573_,
		_w1159_
	);
	LUT2 #(
		.INIT('h2)
	) name1024 (
		\shift[1] ,
		_w595_,
		_w1160_
	);
	LUT2 #(
		.INIT('h1)
	) name1025 (
		_w1159_,
		_w1160_,
		_w1161_
	);
	LUT2 #(
		.INIT('h8)
	) name1026 (
		\shift[1] ,
		_w602_,
		_w1162_
	);
	LUT2 #(
		.INIT('h4)
	) name1027 (
		\shift[1] ,
		_w576_,
		_w1163_
	);
	LUT2 #(
		.INIT('h1)
	) name1028 (
		_w1162_,
		_w1163_,
		_w1164_
	);
	LUT2 #(
		.INIT('h4)
	) name1029 (
		_w1161_,
		_w1164_,
		_w1165_
	);
	LUT2 #(
		.INIT('h2)
	) name1030 (
		_w169_,
		_w1165_,
		_w1166_
	);
	LUT2 #(
		.INIT('h1)
	) name1031 (
		_w1142_,
		_w1150_,
		_w1167_
	);
	LUT2 #(
		.INIT('h1)
	) name1032 (
		_w1158_,
		_w1166_,
		_w1168_
	);
	LUT2 #(
		.INIT('h8)
	) name1033 (
		_w1167_,
		_w1168_,
		_w1169_
	);
	LUT2 #(
		.INIT('h2)
	) name1034 (
		_w228_,
		_w1169_,
		_w1170_
	);
	LUT2 #(
		.INIT('h1)
	) name1035 (
		\shift[1] ,
		_w797_,
		_w1171_
	);
	LUT2 #(
		.INIT('h2)
	) name1036 (
		\shift[1] ,
		_w611_,
		_w1172_
	);
	LUT2 #(
		.INIT('h1)
	) name1037 (
		_w1171_,
		_w1172_,
		_w1173_
	);
	LUT2 #(
		.INIT('h8)
	) name1038 (
		\shift[1] ,
		_w618_,
		_w1174_
	);
	LUT2 #(
		.INIT('h4)
	) name1039 (
		\shift[1] ,
		_w800_,
		_w1175_
	);
	LUT2 #(
		.INIT('h1)
	) name1040 (
		_w1174_,
		_w1175_,
		_w1176_
	);
	LUT2 #(
		.INIT('h4)
	) name1041 (
		_w1173_,
		_w1176_,
		_w1177_
	);
	LUT2 #(
		.INIT('h2)
	) name1042 (
		_w136_,
		_w1177_,
		_w1178_
	);
	LUT2 #(
		.INIT('h1)
	) name1043 (
		\shift[1] ,
		_w613_,
		_w1179_
	);
	LUT2 #(
		.INIT('h2)
	) name1044 (
		\shift[1] ,
		_w623_,
		_w1180_
	);
	LUT2 #(
		.INIT('h1)
	) name1045 (
		_w1179_,
		_w1180_,
		_w1181_
	);
	LUT2 #(
		.INIT('h8)
	) name1046 (
		\shift[1] ,
		_w630_,
		_w1182_
	);
	LUT2 #(
		.INIT('h4)
	) name1047 (
		\shift[1] ,
		_w616_,
		_w1183_
	);
	LUT2 #(
		.INIT('h1)
	) name1048 (
		_w1182_,
		_w1183_,
		_w1184_
	);
	LUT2 #(
		.INIT('h4)
	) name1049 (
		_w1181_,
		_w1184_,
		_w1185_
	);
	LUT2 #(
		.INIT('h2)
	) name1050 (
		_w147_,
		_w1185_,
		_w1186_
	);
	LUT2 #(
		.INIT('h1)
	) name1051 (
		\shift[1] ,
		_w649_,
		_w1187_
	);
	LUT2 #(
		.INIT('h2)
	) name1052 (
		\shift[1] ,
		_w635_,
		_w1188_
	);
	LUT2 #(
		.INIT('h1)
	) name1053 (
		_w1187_,
		_w1188_,
		_w1189_
	);
	LUT2 #(
		.INIT('h8)
	) name1054 (
		\shift[1] ,
		_w642_,
		_w1190_
	);
	LUT2 #(
		.INIT('h4)
	) name1055 (
		\shift[1] ,
		_w652_,
		_w1191_
	);
	LUT2 #(
		.INIT('h1)
	) name1056 (
		_w1190_,
		_w1191_,
		_w1192_
	);
	LUT2 #(
		.INIT('h4)
	) name1057 (
		_w1189_,
		_w1192_,
		_w1193_
	);
	LUT2 #(
		.INIT('h2)
	) name1058 (
		_w158_,
		_w1193_,
		_w1194_
	);
	LUT2 #(
		.INIT('h1)
	) name1059 (
		\shift[1] ,
		_w625_,
		_w1195_
	);
	LUT2 #(
		.INIT('h2)
	) name1060 (
		\shift[1] ,
		_w647_,
		_w1196_
	);
	LUT2 #(
		.INIT('h1)
	) name1061 (
		_w1195_,
		_w1196_,
		_w1197_
	);
	LUT2 #(
		.INIT('h8)
	) name1062 (
		\shift[1] ,
		_w654_,
		_w1198_
	);
	LUT2 #(
		.INIT('h4)
	) name1063 (
		\shift[1] ,
		_w628_,
		_w1199_
	);
	LUT2 #(
		.INIT('h1)
	) name1064 (
		_w1198_,
		_w1199_,
		_w1200_
	);
	LUT2 #(
		.INIT('h4)
	) name1065 (
		_w1197_,
		_w1200_,
		_w1201_
	);
	LUT2 #(
		.INIT('h2)
	) name1066 (
		_w169_,
		_w1201_,
		_w1202_
	);
	LUT2 #(
		.INIT('h1)
	) name1067 (
		_w1178_,
		_w1186_,
		_w1203_
	);
	LUT2 #(
		.INIT('h1)
	) name1068 (
		_w1194_,
		_w1202_,
		_w1204_
	);
	LUT2 #(
		.INIT('h8)
	) name1069 (
		_w1203_,
		_w1204_,
		_w1205_
	);
	LUT2 #(
		.INIT('h2)
	) name1070 (
		_w273_,
		_w1205_,
		_w1206_
	);
	LUT2 #(
		.INIT('h1)
	) name1071 (
		\shift[1] ,
		_w585_,
		_w1207_
	);
	LUT2 #(
		.INIT('h2)
	) name1072 (
		\shift[1] ,
		_w507_,
		_w1208_
	);
	LUT2 #(
		.INIT('h1)
	) name1073 (
		_w1207_,
		_w1208_,
		_w1209_
	);
	LUT2 #(
		.INIT('h8)
	) name1074 (
		\shift[1] ,
		_w514_,
		_w1210_
	);
	LUT2 #(
		.INIT('h4)
	) name1075 (
		\shift[1] ,
		_w588_,
		_w1211_
	);
	LUT2 #(
		.INIT('h1)
	) name1076 (
		_w1210_,
		_w1211_,
		_w1212_
	);
	LUT2 #(
		.INIT('h4)
	) name1077 (
		_w1209_,
		_w1212_,
		_w1213_
	);
	LUT2 #(
		.INIT('h2)
	) name1078 (
		_w136_,
		_w1213_,
		_w1214_
	);
	LUT2 #(
		.INIT('h1)
	) name1079 (
		\shift[1] ,
		_w509_,
		_w1215_
	);
	LUT2 #(
		.INIT('h2)
	) name1080 (
		\shift[1] ,
		_w519_,
		_w1216_
	);
	LUT2 #(
		.INIT('h1)
	) name1081 (
		_w1215_,
		_w1216_,
		_w1217_
	);
	LUT2 #(
		.INIT('h8)
	) name1082 (
		\shift[1] ,
		_w526_,
		_w1218_
	);
	LUT2 #(
		.INIT('h4)
	) name1083 (
		\shift[1] ,
		_w512_,
		_w1219_
	);
	LUT2 #(
		.INIT('h1)
	) name1084 (
		_w1218_,
		_w1219_,
		_w1220_
	);
	LUT2 #(
		.INIT('h4)
	) name1085 (
		_w1217_,
		_w1220_,
		_w1221_
	);
	LUT2 #(
		.INIT('h2)
	) name1086 (
		_w147_,
		_w1221_,
		_w1222_
	);
	LUT2 #(
		.INIT('h1)
	) name1087 (
		\shift[1] ,
		_w545_,
		_w1223_
	);
	LUT2 #(
		.INIT('h2)
	) name1088 (
		\shift[1] ,
		_w531_,
		_w1224_
	);
	LUT2 #(
		.INIT('h1)
	) name1089 (
		_w1223_,
		_w1224_,
		_w1225_
	);
	LUT2 #(
		.INIT('h8)
	) name1090 (
		\shift[1] ,
		_w538_,
		_w1226_
	);
	LUT2 #(
		.INIT('h4)
	) name1091 (
		\shift[1] ,
		_w548_,
		_w1227_
	);
	LUT2 #(
		.INIT('h1)
	) name1092 (
		_w1226_,
		_w1227_,
		_w1228_
	);
	LUT2 #(
		.INIT('h4)
	) name1093 (
		_w1225_,
		_w1228_,
		_w1229_
	);
	LUT2 #(
		.INIT('h2)
	) name1094 (
		_w158_,
		_w1229_,
		_w1230_
	);
	LUT2 #(
		.INIT('h1)
	) name1095 (
		\shift[1] ,
		_w521_,
		_w1231_
	);
	LUT2 #(
		.INIT('h2)
	) name1096 (
		\shift[1] ,
		_w543_,
		_w1232_
	);
	LUT2 #(
		.INIT('h1)
	) name1097 (
		_w1231_,
		_w1232_,
		_w1233_
	);
	LUT2 #(
		.INIT('h8)
	) name1098 (
		\shift[1] ,
		_w550_,
		_w1234_
	);
	LUT2 #(
		.INIT('h4)
	) name1099 (
		\shift[1] ,
		_w524_,
		_w1235_
	);
	LUT2 #(
		.INIT('h1)
	) name1100 (
		_w1234_,
		_w1235_,
		_w1236_
	);
	LUT2 #(
		.INIT('h4)
	) name1101 (
		_w1233_,
		_w1236_,
		_w1237_
	);
	LUT2 #(
		.INIT('h2)
	) name1102 (
		_w169_,
		_w1237_,
		_w1238_
	);
	LUT2 #(
		.INIT('h1)
	) name1103 (
		_w1214_,
		_w1222_,
		_w1239_
	);
	LUT2 #(
		.INIT('h1)
	) name1104 (
		_w1230_,
		_w1238_,
		_w1240_
	);
	LUT2 #(
		.INIT('h8)
	) name1105 (
		_w1239_,
		_w1240_,
		_w1241_
	);
	LUT2 #(
		.INIT('h2)
	) name1106 (
		_w183_,
		_w1241_,
		_w1242_
	);
	LUT2 #(
		.INIT('h1)
	) name1107 (
		_w1134_,
		_w1170_,
		_w1243_
	);
	LUT2 #(
		.INIT('h1)
	) name1108 (
		_w1206_,
		_w1242_,
		_w1244_
	);
	LUT2 #(
		.INIT('h8)
	) name1109 (
		_w1243_,
		_w1244_,
		_w1245_
	);
	LUT2 #(
		.INIT('h1)
	) name1110 (
		\shift[6] ,
		_w1245_,
		_w1246_
	);
	LUT2 #(
		.INIT('h1)
	) name1111 (
		\shift[1] ,
		_w533_,
		_w1247_
	);
	LUT2 #(
		.INIT('h2)
	) name1112 (
		\shift[1] ,
		_w719_,
		_w1248_
	);
	LUT2 #(
		.INIT('h1)
	) name1113 (
		_w1247_,
		_w1248_,
		_w1249_
	);
	LUT2 #(
		.INIT('h8)
	) name1114 (
		\shift[1] ,
		_w726_,
		_w1250_
	);
	LUT2 #(
		.INIT('h4)
	) name1115 (
		\shift[1] ,
		_w536_,
		_w1251_
	);
	LUT2 #(
		.INIT('h1)
	) name1116 (
		_w1250_,
		_w1251_,
		_w1252_
	);
	LUT2 #(
		.INIT('h4)
	) name1117 (
		_w1249_,
		_w1252_,
		_w1253_
	);
	LUT2 #(
		.INIT('h2)
	) name1118 (
		_w136_,
		_w1253_,
		_w1254_
	);
	LUT2 #(
		.INIT('h1)
	) name1119 (
		\shift[1] ,
		_w721_,
		_w1255_
	);
	LUT2 #(
		.INIT('h2)
	) name1120 (
		\shift[1] ,
		_w731_,
		_w1256_
	);
	LUT2 #(
		.INIT('h1)
	) name1121 (
		_w1255_,
		_w1256_,
		_w1257_
	);
	LUT2 #(
		.INIT('h8)
	) name1122 (
		\shift[1] ,
		_w738_,
		_w1258_
	);
	LUT2 #(
		.INIT('h4)
	) name1123 (
		\shift[1] ,
		_w724_,
		_w1259_
	);
	LUT2 #(
		.INIT('h1)
	) name1124 (
		_w1258_,
		_w1259_,
		_w1260_
	);
	LUT2 #(
		.INIT('h4)
	) name1125 (
		_w1257_,
		_w1260_,
		_w1261_
	);
	LUT2 #(
		.INIT('h2)
	) name1126 (
		_w147_,
		_w1261_,
		_w1262_
	);
	LUT2 #(
		.INIT('h1)
	) name1127 (
		\shift[1] ,
		_w757_,
		_w1263_
	);
	LUT2 #(
		.INIT('h2)
	) name1128 (
		\shift[1] ,
		_w743_,
		_w1264_
	);
	LUT2 #(
		.INIT('h1)
	) name1129 (
		_w1263_,
		_w1264_,
		_w1265_
	);
	LUT2 #(
		.INIT('h8)
	) name1130 (
		\shift[1] ,
		_w750_,
		_w1266_
	);
	LUT2 #(
		.INIT('h4)
	) name1131 (
		\shift[1] ,
		_w760_,
		_w1267_
	);
	LUT2 #(
		.INIT('h1)
	) name1132 (
		_w1266_,
		_w1267_,
		_w1268_
	);
	LUT2 #(
		.INIT('h4)
	) name1133 (
		_w1265_,
		_w1268_,
		_w1269_
	);
	LUT2 #(
		.INIT('h2)
	) name1134 (
		_w158_,
		_w1269_,
		_w1270_
	);
	LUT2 #(
		.INIT('h1)
	) name1135 (
		\shift[1] ,
		_w733_,
		_w1271_
	);
	LUT2 #(
		.INIT('h2)
	) name1136 (
		\shift[1] ,
		_w755_,
		_w1272_
	);
	LUT2 #(
		.INIT('h1)
	) name1137 (
		_w1271_,
		_w1272_,
		_w1273_
	);
	LUT2 #(
		.INIT('h8)
	) name1138 (
		\shift[1] ,
		_w762_,
		_w1274_
	);
	LUT2 #(
		.INIT('h4)
	) name1139 (
		\shift[1] ,
		_w736_,
		_w1275_
	);
	LUT2 #(
		.INIT('h1)
	) name1140 (
		_w1274_,
		_w1275_,
		_w1276_
	);
	LUT2 #(
		.INIT('h4)
	) name1141 (
		_w1273_,
		_w1276_,
		_w1277_
	);
	LUT2 #(
		.INIT('h2)
	) name1142 (
		_w169_,
		_w1277_,
		_w1278_
	);
	LUT2 #(
		.INIT('h1)
	) name1143 (
		_w1254_,
		_w1262_,
		_w1279_
	);
	LUT2 #(
		.INIT('h1)
	) name1144 (
		_w1270_,
		_w1278_,
		_w1280_
	);
	LUT2 #(
		.INIT('h8)
	) name1145 (
		_w1279_,
		_w1280_,
		_w1281_
	);
	LUT2 #(
		.INIT('h2)
	) name1146 (
		_w273_,
		_w1281_,
		_w1282_
	);
	LUT2 #(
		.INIT('h1)
	) name1147 (
		\shift[1] ,
		_w745_,
		_w1283_
	);
	LUT2 #(
		.INIT('h2)
	) name1148 (
		\shift[1] ,
		_w823_,
		_w1284_
	);
	LUT2 #(
		.INIT('h1)
	) name1149 (
		_w1283_,
		_w1284_,
		_w1285_
	);
	LUT2 #(
		.INIT('h8)
	) name1150 (
		\shift[1] ,
		_w830_,
		_w1286_
	);
	LUT2 #(
		.INIT('h4)
	) name1151 (
		\shift[1] ,
		_w748_,
		_w1287_
	);
	LUT2 #(
		.INIT('h1)
	) name1152 (
		_w1286_,
		_w1287_,
		_w1288_
	);
	LUT2 #(
		.INIT('h4)
	) name1153 (
		_w1285_,
		_w1288_,
		_w1289_
	);
	LUT2 #(
		.INIT('h2)
	) name1154 (
		_w136_,
		_w1289_,
		_w1290_
	);
	LUT2 #(
		.INIT('h2)
	) name1155 (
		\shift[1] ,
		_w841_,
		_w1291_
	);
	LUT2 #(
		.INIT('h1)
	) name1156 (
		_w825_,
		_w828_,
		_w1292_
	);
	LUT2 #(
		.INIT('h1)
	) name1157 (
		\shift[1] ,
		_w1292_,
		_w1293_
	);
	LUT2 #(
		.INIT('h1)
	) name1158 (
		_w1291_,
		_w1293_,
		_w1294_
	);
	LUT2 #(
		.INIT('h2)
	) name1159 (
		_w147_,
		_w1294_,
		_w1295_
	);
	LUT2 #(
		.INIT('h1)
	) name1160 (
		\shift[1] ,
		_w862_,
		_w1296_
	);
	LUT2 #(
		.INIT('h2)
	) name1161 (
		\shift[1] ,
		_w845_,
		_w1297_
	);
	LUT2 #(
		.INIT('h1)
	) name1162 (
		_w1296_,
		_w1297_,
		_w1298_
	);
	LUT2 #(
		.INIT('h8)
	) name1163 (
		\shift[1] ,
		_w852_,
		_w1299_
	);
	LUT2 #(
		.INIT('h4)
	) name1164 (
		\shift[1] ,
		_w861_,
		_w1300_
	);
	LUT2 #(
		.INIT('h1)
	) name1165 (
		_w1299_,
		_w1300_,
		_w1301_
	);
	LUT2 #(
		.INIT('h4)
	) name1166 (
		_w1298_,
		_w1301_,
		_w1302_
	);
	LUT2 #(
		.INIT('h2)
	) name1167 (
		_w158_,
		_w1302_,
		_w1303_
	);
	LUT2 #(
		.INIT('h1)
	) name1168 (
		\shift[1] ,
		_w835_,
		_w1304_
	);
	LUT2 #(
		.INIT('h2)
	) name1169 (
		\shift[1] ,
		_w857_,
		_w1305_
	);
	LUT2 #(
		.INIT('h1)
	) name1170 (
		_w1304_,
		_w1305_,
		_w1306_
	);
	LUT2 #(
		.INIT('h8)
	) name1171 (
		\shift[1] ,
		_w858_,
		_w1307_
	);
	LUT2 #(
		.INIT('h4)
	) name1172 (
		\shift[1] ,
		_w836_,
		_w1308_
	);
	LUT2 #(
		.INIT('h1)
	) name1173 (
		_w1307_,
		_w1308_,
		_w1309_
	);
	LUT2 #(
		.INIT('h4)
	) name1174 (
		_w1306_,
		_w1309_,
		_w1310_
	);
	LUT2 #(
		.INIT('h2)
	) name1175 (
		_w169_,
		_w1310_,
		_w1311_
	);
	LUT2 #(
		.INIT('h1)
	) name1176 (
		_w1290_,
		_w1295_,
		_w1312_
	);
	LUT2 #(
		.INIT('h1)
	) name1177 (
		_w1303_,
		_w1311_,
		_w1313_
	);
	LUT2 #(
		.INIT('h8)
	) name1178 (
		_w1312_,
		_w1313_,
		_w1314_
	);
	LUT2 #(
		.INIT('h2)
	) name1179 (
		_w318_,
		_w1314_,
		_w1315_
	);
	LUT2 #(
		.INIT('h1)
	) name1180 (
		\shift[1] ,
		_w897_,
		_w1316_
	);
	LUT2 #(
		.INIT('h2)
	) name1181 (
		\shift[1] ,
		_w771_,
		_w1317_
	);
	LUT2 #(
		.INIT('h1)
	) name1182 (
		_w1316_,
		_w1317_,
		_w1318_
	);
	LUT2 #(
		.INIT('h8)
	) name1183 (
		\shift[1] ,
		_w778_,
		_w1319_
	);
	LUT2 #(
		.INIT('h4)
	) name1184 (
		\shift[1] ,
		_w900_,
		_w1320_
	);
	LUT2 #(
		.INIT('h1)
	) name1185 (
		_w1319_,
		_w1320_,
		_w1321_
	);
	LUT2 #(
		.INIT('h4)
	) name1186 (
		_w1318_,
		_w1321_,
		_w1322_
	);
	LUT2 #(
		.INIT('h2)
	) name1187 (
		_w136_,
		_w1322_,
		_w1323_
	);
	LUT2 #(
		.INIT('h1)
	) name1188 (
		\shift[1] ,
		_w773_,
		_w1324_
	);
	LUT2 #(
		.INIT('h2)
	) name1189 (
		\shift[1] ,
		_w783_,
		_w1325_
	);
	LUT2 #(
		.INIT('h1)
	) name1190 (
		_w1324_,
		_w1325_,
		_w1326_
	);
	LUT2 #(
		.INIT('h8)
	) name1191 (
		\shift[1] ,
		_w790_,
		_w1327_
	);
	LUT2 #(
		.INIT('h4)
	) name1192 (
		\shift[1] ,
		_w776_,
		_w1328_
	);
	LUT2 #(
		.INIT('h1)
	) name1193 (
		_w1327_,
		_w1328_,
		_w1329_
	);
	LUT2 #(
		.INIT('h4)
	) name1194 (
		_w1326_,
		_w1329_,
		_w1330_
	);
	LUT2 #(
		.INIT('h2)
	) name1195 (
		_w147_,
		_w1330_,
		_w1331_
	);
	LUT2 #(
		.INIT('h1)
	) name1196 (
		\shift[1] ,
		_w809_,
		_w1332_
	);
	LUT2 #(
		.INIT('h2)
	) name1197 (
		\shift[1] ,
		_w795_,
		_w1333_
	);
	LUT2 #(
		.INIT('h1)
	) name1198 (
		_w1332_,
		_w1333_,
		_w1334_
	);
	LUT2 #(
		.INIT('h8)
	) name1199 (
		\shift[1] ,
		_w802_,
		_w1335_
	);
	LUT2 #(
		.INIT('h4)
	) name1200 (
		\shift[1] ,
		_w812_,
		_w1336_
	);
	LUT2 #(
		.INIT('h1)
	) name1201 (
		_w1335_,
		_w1336_,
		_w1337_
	);
	LUT2 #(
		.INIT('h4)
	) name1202 (
		_w1334_,
		_w1337_,
		_w1338_
	);
	LUT2 #(
		.INIT('h2)
	) name1203 (
		_w158_,
		_w1338_,
		_w1339_
	);
	LUT2 #(
		.INIT('h1)
	) name1204 (
		\shift[1] ,
		_w785_,
		_w1340_
	);
	LUT2 #(
		.INIT('h2)
	) name1205 (
		\shift[1] ,
		_w807_,
		_w1341_
	);
	LUT2 #(
		.INIT('h1)
	) name1206 (
		_w1340_,
		_w1341_,
		_w1342_
	);
	LUT2 #(
		.INIT('h8)
	) name1207 (
		\shift[1] ,
		_w814_,
		_w1343_
	);
	LUT2 #(
		.INIT('h4)
	) name1208 (
		\shift[1] ,
		_w788_,
		_w1344_
	);
	LUT2 #(
		.INIT('h1)
	) name1209 (
		_w1343_,
		_w1344_,
		_w1345_
	);
	LUT2 #(
		.INIT('h4)
	) name1210 (
		_w1342_,
		_w1345_,
		_w1346_
	);
	LUT2 #(
		.INIT('h2)
	) name1211 (
		_w169_,
		_w1346_,
		_w1347_
	);
	LUT2 #(
		.INIT('h1)
	) name1212 (
		_w1323_,
		_w1331_,
		_w1348_
	);
	LUT2 #(
		.INIT('h1)
	) name1213 (
		_w1339_,
		_w1347_,
		_w1349_
	);
	LUT2 #(
		.INIT('h8)
	) name1214 (
		_w1348_,
		_w1349_,
		_w1350_
	);
	LUT2 #(
		.INIT('h2)
	) name1215 (
		_w183_,
		_w1350_,
		_w1351_
	);
	LUT2 #(
		.INIT('h1)
	) name1216 (
		\shift[1] ,
		_w847_,
		_w1352_
	);
	LUT2 #(
		.INIT('h2)
	) name1217 (
		\shift[1] ,
		_w871_,
		_w1353_
	);
	LUT2 #(
		.INIT('h1)
	) name1218 (
		_w1352_,
		_w1353_,
		_w1354_
	);
	LUT2 #(
		.INIT('h8)
	) name1219 (
		\shift[1] ,
		_w878_,
		_w1355_
	);
	LUT2 #(
		.INIT('h4)
	) name1220 (
		\shift[1] ,
		_w850_,
		_w1356_
	);
	LUT2 #(
		.INIT('h1)
	) name1221 (
		_w1355_,
		_w1356_,
		_w1357_
	);
	LUT2 #(
		.INIT('h4)
	) name1222 (
		_w1354_,
		_w1357_,
		_w1358_
	);
	LUT2 #(
		.INIT('h2)
	) name1223 (
		_w136_,
		_w1358_,
		_w1359_
	);
	LUT2 #(
		.INIT('h1)
	) name1224 (
		\shift[1] ,
		_w873_,
		_w1360_
	);
	LUT2 #(
		.INIT('h2)
	) name1225 (
		\shift[1] ,
		_w883_,
		_w1361_
	);
	LUT2 #(
		.INIT('h1)
	) name1226 (
		_w1360_,
		_w1361_,
		_w1362_
	);
	LUT2 #(
		.INIT('h8)
	) name1227 (
		\shift[1] ,
		_w890_,
		_w1363_
	);
	LUT2 #(
		.INIT('h4)
	) name1228 (
		\shift[1] ,
		_w876_,
		_w1364_
	);
	LUT2 #(
		.INIT('h1)
	) name1229 (
		_w1363_,
		_w1364_,
		_w1365_
	);
	LUT2 #(
		.INIT('h4)
	) name1230 (
		_w1362_,
		_w1365_,
		_w1366_
	);
	LUT2 #(
		.INIT('h2)
	) name1231 (
		_w147_,
		_w1366_,
		_w1367_
	);
	LUT2 #(
		.INIT('h1)
	) name1232 (
		\shift[1] ,
		_w909_,
		_w1368_
	);
	LUT2 #(
		.INIT('h2)
	) name1233 (
		\shift[1] ,
		_w895_,
		_w1369_
	);
	LUT2 #(
		.INIT('h1)
	) name1234 (
		_w1368_,
		_w1369_,
		_w1370_
	);
	LUT2 #(
		.INIT('h8)
	) name1235 (
		\shift[1] ,
		_w902_,
		_w1371_
	);
	LUT2 #(
		.INIT('h4)
	) name1236 (
		\shift[1] ,
		_w912_,
		_w1372_
	);
	LUT2 #(
		.INIT('h1)
	) name1237 (
		_w1371_,
		_w1372_,
		_w1373_
	);
	LUT2 #(
		.INIT('h4)
	) name1238 (
		_w1370_,
		_w1373_,
		_w1374_
	);
	LUT2 #(
		.INIT('h2)
	) name1239 (
		_w158_,
		_w1374_,
		_w1375_
	);
	LUT2 #(
		.INIT('h1)
	) name1240 (
		\shift[1] ,
		_w885_,
		_w1376_
	);
	LUT2 #(
		.INIT('h2)
	) name1241 (
		\shift[1] ,
		_w907_,
		_w1377_
	);
	LUT2 #(
		.INIT('h1)
	) name1242 (
		_w1376_,
		_w1377_,
		_w1378_
	);
	LUT2 #(
		.INIT('h8)
	) name1243 (
		\shift[1] ,
		_w914_,
		_w1379_
	);
	LUT2 #(
		.INIT('h4)
	) name1244 (
		\shift[1] ,
		_w888_,
		_w1380_
	);
	LUT2 #(
		.INIT('h1)
	) name1245 (
		_w1379_,
		_w1380_,
		_w1381_
	);
	LUT2 #(
		.INIT('h4)
	) name1246 (
		_w1378_,
		_w1381_,
		_w1382_
	);
	LUT2 #(
		.INIT('h2)
	) name1247 (
		_w169_,
		_w1382_,
		_w1383_
	);
	LUT2 #(
		.INIT('h1)
	) name1248 (
		_w1359_,
		_w1367_,
		_w1384_
	);
	LUT2 #(
		.INIT('h1)
	) name1249 (
		_w1375_,
		_w1383_,
		_w1385_
	);
	LUT2 #(
		.INIT('h8)
	) name1250 (
		_w1384_,
		_w1385_,
		_w1386_
	);
	LUT2 #(
		.INIT('h2)
	) name1251 (
		_w228_,
		_w1386_,
		_w1387_
	);
	LUT2 #(
		.INIT('h1)
	) name1252 (
		_w1282_,
		_w1315_,
		_w1388_
	);
	LUT2 #(
		.INIT('h1)
	) name1253 (
		_w1351_,
		_w1387_,
		_w1389_
	);
	LUT2 #(
		.INIT('h8)
	) name1254 (
		_w1388_,
		_w1389_,
		_w1390_
	);
	LUT2 #(
		.INIT('h2)
	) name1255 (
		\shift[6] ,
		_w1390_,
		_w1391_
	);
	LUT2 #(
		.INIT('h1)
	) name1256 (
		_w1246_,
		_w1391_,
		_w1392_
	);
	LUT2 #(
		.INIT('h2)
	) name1257 (
		_w136_,
		_w213_,
		_w1393_
	);
	LUT2 #(
		.INIT('h4)
	) name1258 (
		_w145_,
		_w147_,
		_w1394_
	);
	LUT2 #(
		.INIT('h2)
	) name1259 (
		_w158_,
		_w178_,
		_w1395_
	);
	LUT2 #(
		.INIT('h4)
	) name1260 (
		_w156_,
		_w169_,
		_w1396_
	);
	LUT2 #(
		.INIT('h1)
	) name1261 (
		_w1393_,
		_w1394_,
		_w1397_
	);
	LUT2 #(
		.INIT('h1)
	) name1262 (
		_w1395_,
		_w1396_,
		_w1398_
	);
	LUT2 #(
		.INIT('h8)
	) name1263 (
		_w1397_,
		_w1398_,
		_w1399_
	);
	LUT2 #(
		.INIT('h2)
	) name1264 (
		_w183_,
		_w1399_,
		_w1400_
	);
	LUT2 #(
		.INIT('h2)
	) name1265 (
		_w136_,
		_w303_,
		_w1401_
	);
	LUT2 #(
		.INIT('h2)
	) name1266 (
		_w147_,
		_w193_,
		_w1402_
	);
	LUT2 #(
		.INIT('h2)
	) name1267 (
		_w158_,
		_w223_,
		_w1403_
	);
	LUT2 #(
		.INIT('h2)
	) name1268 (
		_w169_,
		_w203_,
		_w1404_
	);
	LUT2 #(
		.INIT('h1)
	) name1269 (
		_w1401_,
		_w1402_,
		_w1405_
	);
	LUT2 #(
		.INIT('h1)
	) name1270 (
		_w1403_,
		_w1404_,
		_w1406_
	);
	LUT2 #(
		.INIT('h8)
	) name1271 (
		_w1405_,
		_w1406_,
		_w1407_
	);
	LUT2 #(
		.INIT('h2)
	) name1272 (
		_w228_,
		_w1407_,
		_w1408_
	);
	LUT2 #(
		.INIT('h2)
	) name1273 (
		_w136_,
		_w352_,
		_w1409_
	);
	LUT2 #(
		.INIT('h2)
	) name1274 (
		_w147_,
		_w238_,
		_w1410_
	);
	LUT2 #(
		.INIT('h2)
	) name1275 (
		_w158_,
		_w268_,
		_w1411_
	);
	LUT2 #(
		.INIT('h2)
	) name1276 (
		_w169_,
		_w248_,
		_w1412_
	);
	LUT2 #(
		.INIT('h1)
	) name1277 (
		_w1409_,
		_w1410_,
		_w1413_
	);
	LUT2 #(
		.INIT('h1)
	) name1278 (
		_w1411_,
		_w1412_,
		_w1414_
	);
	LUT2 #(
		.INIT('h8)
	) name1279 (
		_w1413_,
		_w1414_,
		_w1415_
	);
	LUT2 #(
		.INIT('h2)
	) name1280 (
		_w273_,
		_w1415_,
		_w1416_
	);
	LUT2 #(
		.INIT('h2)
	) name1281 (
		_w136_,
		_w258_,
		_w1417_
	);
	LUT2 #(
		.INIT('h2)
	) name1282 (
		_w147_,
		_w283_,
		_w1418_
	);
	LUT2 #(
		.INIT('h2)
	) name1283 (
		_w158_,
		_w313_,
		_w1419_
	);
	LUT2 #(
		.INIT('h2)
	) name1284 (
		_w169_,
		_w293_,
		_w1420_
	);
	LUT2 #(
		.INIT('h1)
	) name1285 (
		_w1417_,
		_w1418_,
		_w1421_
	);
	LUT2 #(
		.INIT('h1)
	) name1286 (
		_w1419_,
		_w1420_,
		_w1422_
	);
	LUT2 #(
		.INIT('h8)
	) name1287 (
		_w1421_,
		_w1422_,
		_w1423_
	);
	LUT2 #(
		.INIT('h2)
	) name1288 (
		_w318_,
		_w1423_,
		_w1424_
	);
	LUT2 #(
		.INIT('h1)
	) name1289 (
		_w1400_,
		_w1408_,
		_w1425_
	);
	LUT2 #(
		.INIT('h1)
	) name1290 (
		_w1416_,
		_w1424_,
		_w1426_
	);
	LUT2 #(
		.INIT('h8)
	) name1291 (
		_w1425_,
		_w1426_,
		_w1427_
	);
	LUT2 #(
		.INIT('h1)
	) name1292 (
		\shift[6] ,
		_w1427_,
		_w1428_
	);
	LUT2 #(
		.INIT('h2)
	) name1293 (
		_w136_,
		_w440_,
		_w1429_
	);
	LUT2 #(
		.INIT('h2)
	) name1294 (
		_w147_,
		_w464_,
		_w1430_
	);
	LUT2 #(
		.INIT('h2)
	) name1295 (
		_w158_,
		_w496_,
		_w1431_
	);
	LUT2 #(
		.INIT('h2)
	) name1296 (
		_w169_,
		_w474_,
		_w1432_
	);
	LUT2 #(
		.INIT('h1)
	) name1297 (
		_w1429_,
		_w1430_,
		_w1433_
	);
	LUT2 #(
		.INIT('h1)
	) name1298 (
		_w1431_,
		_w1432_,
		_w1434_
	);
	LUT2 #(
		.INIT('h8)
	) name1299 (
		_w1433_,
		_w1434_,
		_w1435_
	);
	LUT2 #(
		.INIT('h2)
	) name1300 (
		_w318_,
		_w1435_,
		_w1436_
	);
	LUT2 #(
		.INIT('h2)
	) name1301 (
		_w136_,
		_w167_,
		_w1437_
	);
	LUT2 #(
		.INIT('h2)
	) name1302 (
		_w147_,
		_w420_,
		_w1438_
	);
	LUT2 #(
		.INIT('h2)
	) name1303 (
		_w158_,
		_w450_,
		_w1439_
	);
	LUT2 #(
		.INIT('h2)
	) name1304 (
		_w169_,
		_w430_,
		_w1440_
	);
	LUT2 #(
		.INIT('h1)
	) name1305 (
		_w1437_,
		_w1438_,
		_w1441_
	);
	LUT2 #(
		.INIT('h1)
	) name1306 (
		_w1439_,
		_w1440_,
		_w1442_
	);
	LUT2 #(
		.INIT('h8)
	) name1307 (
		_w1441_,
		_w1442_,
		_w1443_
	);
	LUT2 #(
		.INIT('h2)
	) name1308 (
		_w273_,
		_w1443_,
		_w1444_
	);
	LUT2 #(
		.INIT('h2)
	) name1309 (
		_w136_,
		_w484_,
		_w1445_
	);
	LUT2 #(
		.INIT('h2)
	) name1310 (
		_w147_,
		_w376_,
		_w1446_
	);
	LUT2 #(
		.INIT('h2)
	) name1311 (
		_w158_,
		_w406_,
		_w1447_
	);
	LUT2 #(
		.INIT('h2)
	) name1312 (
		_w169_,
		_w386_,
		_w1448_
	);
	LUT2 #(
		.INIT('h1)
	) name1313 (
		_w1445_,
		_w1446_,
		_w1449_
	);
	LUT2 #(
		.INIT('h1)
	) name1314 (
		_w1447_,
		_w1448_,
		_w1450_
	);
	LUT2 #(
		.INIT('h8)
	) name1315 (
		_w1449_,
		_w1450_,
		_w1451_
	);
	LUT2 #(
		.INIT('h2)
	) name1316 (
		_w228_,
		_w1451_,
		_w1452_
	);
	LUT2 #(
		.INIT('h2)
	) name1317 (
		_w136_,
		_w396_,
		_w1453_
	);
	LUT2 #(
		.INIT('h2)
	) name1318 (
		_w147_,
		_w332_,
		_w1454_
	);
	LUT2 #(
		.INIT('h2)
	) name1319 (
		_w158_,
		_w362_,
		_w1455_
	);
	LUT2 #(
		.INIT('h2)
	) name1320 (
		_w169_,
		_w342_,
		_w1456_
	);
	LUT2 #(
		.INIT('h1)
	) name1321 (
		_w1453_,
		_w1454_,
		_w1457_
	);
	LUT2 #(
		.INIT('h1)
	) name1322 (
		_w1455_,
		_w1456_,
		_w1458_
	);
	LUT2 #(
		.INIT('h8)
	) name1323 (
		_w1457_,
		_w1458_,
		_w1459_
	);
	LUT2 #(
		.INIT('h2)
	) name1324 (
		_w183_,
		_w1459_,
		_w1460_
	);
	LUT2 #(
		.INIT('h1)
	) name1325 (
		_w1436_,
		_w1444_,
		_w1461_
	);
	LUT2 #(
		.INIT('h1)
	) name1326 (
		_w1452_,
		_w1460_,
		_w1462_
	);
	LUT2 #(
		.INIT('h8)
	) name1327 (
		_w1461_,
		_w1462_,
		_w1463_
	);
	LUT2 #(
		.INIT('h2)
	) name1328 (
		\shift[6] ,
		_w1463_,
		_w1464_
	);
	LUT2 #(
		.INIT('h1)
	) name1329 (
		_w1428_,
		_w1464_,
		_w1465_
	);
	LUT2 #(
		.INIT('h2)
	) name1330 (
		_w136_,
		_w593_,
		_w1466_
	);
	LUT2 #(
		.INIT('h2)
	) name1331 (
		_w147_,
		_w517_,
		_w1467_
	);
	LUT2 #(
		.INIT('h2)
	) name1332 (
		_w158_,
		_w553_,
		_w1468_
	);
	LUT2 #(
		.INIT('h2)
	) name1333 (
		_w169_,
		_w529_,
		_w1469_
	);
	LUT2 #(
		.INIT('h1)
	) name1334 (
		_w1466_,
		_w1467_,
		_w1470_
	);
	LUT2 #(
		.INIT('h1)
	) name1335 (
		_w1468_,
		_w1469_,
		_w1471_
	);
	LUT2 #(
		.INIT('h8)
	) name1336 (
		_w1470_,
		_w1471_,
		_w1472_
	);
	LUT2 #(
		.INIT('h2)
	) name1337 (
		_w183_,
		_w1472_,
		_w1473_
	);
	LUT2 #(
		.INIT('h2)
	) name1338 (
		_w136_,
		_w697_,
		_w1474_
	);
	LUT2 #(
		.INIT('h2)
	) name1339 (
		_w147_,
		_w569_,
		_w1475_
	);
	LUT2 #(
		.INIT('h2)
	) name1340 (
		_w158_,
		_w605_,
		_w1476_
	);
	LUT2 #(
		.INIT('h2)
	) name1341 (
		_w169_,
		_w581_,
		_w1477_
	);
	LUT2 #(
		.INIT('h1)
	) name1342 (
		_w1474_,
		_w1475_,
		_w1478_
	);
	LUT2 #(
		.INIT('h1)
	) name1343 (
		_w1476_,
		_w1477_,
		_w1479_
	);
	LUT2 #(
		.INIT('h8)
	) name1344 (
		_w1478_,
		_w1479_,
		_w1480_
	);
	LUT2 #(
		.INIT('h2)
	) name1345 (
		_w228_,
		_w1480_,
		_w1481_
	);
	LUT2 #(
		.INIT('h2)
	) name1346 (
		_w136_,
		_w805_,
		_w1482_
	);
	LUT2 #(
		.INIT('h2)
	) name1347 (
		_w147_,
		_w621_,
		_w1483_
	);
	LUT2 #(
		.INIT('h2)
	) name1348 (
		_w158_,
		_w657_,
		_w1484_
	);
	LUT2 #(
		.INIT('h2)
	) name1349 (
		_w169_,
		_w633_,
		_w1485_
	);
	LUT2 #(
		.INIT('h1)
	) name1350 (
		_w1482_,
		_w1483_,
		_w1486_
	);
	LUT2 #(
		.INIT('h1)
	) name1351 (
		_w1484_,
		_w1485_,
		_w1487_
	);
	LUT2 #(
		.INIT('h8)
	) name1352 (
		_w1486_,
		_w1487_,
		_w1488_
	);
	LUT2 #(
		.INIT('h2)
	) name1353 (
		_w273_,
		_w1488_,
		_w1489_
	);
	LUT2 #(
		.INIT('h2)
	) name1354 (
		_w136_,
		_w645_,
		_w1490_
	);
	LUT2 #(
		.INIT('h2)
	) name1355 (
		_w147_,
		_w673_,
		_w1491_
	);
	LUT2 #(
		.INIT('h2)
	) name1356 (
		_w158_,
		_w709_,
		_w1492_
	);
	LUT2 #(
		.INIT('h2)
	) name1357 (
		_w169_,
		_w685_,
		_w1493_
	);
	LUT2 #(
		.INIT('h1)
	) name1358 (
		_w1490_,
		_w1491_,
		_w1494_
	);
	LUT2 #(
		.INIT('h1)
	) name1359 (
		_w1492_,
		_w1493_,
		_w1495_
	);
	LUT2 #(
		.INIT('h8)
	) name1360 (
		_w1494_,
		_w1495_,
		_w1496_
	);
	LUT2 #(
		.INIT('h2)
	) name1361 (
		_w318_,
		_w1496_,
		_w1497_
	);
	LUT2 #(
		.INIT('h1)
	) name1362 (
		_w1473_,
		_w1481_,
		_w1498_
	);
	LUT2 #(
		.INIT('h1)
	) name1363 (
		_w1489_,
		_w1497_,
		_w1499_
	);
	LUT2 #(
		.INIT('h8)
	) name1364 (
		_w1498_,
		_w1499_,
		_w1500_
	);
	LUT2 #(
		.INIT('h1)
	) name1365 (
		\shift[6] ,
		_w1500_,
		_w1501_
	);
	LUT2 #(
		.INIT('h2)
	) name1366 (
		_w136_,
		_w753_,
		_w1502_
	);
	LUT2 #(
		.INIT('h2)
	) name1367 (
		_w147_,
		_w833_,
		_w1503_
	);
	LUT2 #(
		.INIT('h2)
	) name1368 (
		_w158_,
		_w865_,
		_w1504_
	);
	LUT2 #(
		.INIT('h2)
	) name1369 (
		_w169_,
		_w843_,
		_w1505_
	);
	LUT2 #(
		.INIT('h1)
	) name1370 (
		_w1502_,
		_w1503_,
		_w1506_
	);
	LUT2 #(
		.INIT('h1)
	) name1371 (
		_w1504_,
		_w1505_,
		_w1507_
	);
	LUT2 #(
		.INIT('h8)
	) name1372 (
		_w1506_,
		_w1507_,
		_w1508_
	);
	LUT2 #(
		.INIT('h2)
	) name1373 (
		_w318_,
		_w1508_,
		_w1509_
	);
	LUT2 #(
		.INIT('h2)
	) name1374 (
		_w136_,
		_w541_,
		_w1510_
	);
	LUT2 #(
		.INIT('h2)
	) name1375 (
		_w147_,
		_w729_,
		_w1511_
	);
	LUT2 #(
		.INIT('h2)
	) name1376 (
		_w158_,
		_w765_,
		_w1512_
	);
	LUT2 #(
		.INIT('h2)
	) name1377 (
		_w169_,
		_w741_,
		_w1513_
	);
	LUT2 #(
		.INIT('h1)
	) name1378 (
		_w1510_,
		_w1511_,
		_w1514_
	);
	LUT2 #(
		.INIT('h1)
	) name1379 (
		_w1512_,
		_w1513_,
		_w1515_
	);
	LUT2 #(
		.INIT('h8)
	) name1380 (
		_w1514_,
		_w1515_,
		_w1516_
	);
	LUT2 #(
		.INIT('h2)
	) name1381 (
		_w273_,
		_w1516_,
		_w1517_
	);
	LUT2 #(
		.INIT('h2)
	) name1382 (
		_w136_,
		_w855_,
		_w1518_
	);
	LUT2 #(
		.INIT('h2)
	) name1383 (
		_w147_,
		_w881_,
		_w1519_
	);
	LUT2 #(
		.INIT('h2)
	) name1384 (
		_w158_,
		_w917_,
		_w1520_
	);
	LUT2 #(
		.INIT('h2)
	) name1385 (
		_w169_,
		_w893_,
		_w1521_
	);
	LUT2 #(
		.INIT('h1)
	) name1386 (
		_w1518_,
		_w1519_,
		_w1522_
	);
	LUT2 #(
		.INIT('h1)
	) name1387 (
		_w1520_,
		_w1521_,
		_w1523_
	);
	LUT2 #(
		.INIT('h8)
	) name1388 (
		_w1522_,
		_w1523_,
		_w1524_
	);
	LUT2 #(
		.INIT('h2)
	) name1389 (
		_w228_,
		_w1524_,
		_w1525_
	);
	LUT2 #(
		.INIT('h2)
	) name1390 (
		_w136_,
		_w905_,
		_w1526_
	);
	LUT2 #(
		.INIT('h2)
	) name1391 (
		_w147_,
		_w781_,
		_w1527_
	);
	LUT2 #(
		.INIT('h2)
	) name1392 (
		_w158_,
		_w817_,
		_w1528_
	);
	LUT2 #(
		.INIT('h2)
	) name1393 (
		_w169_,
		_w793_,
		_w1529_
	);
	LUT2 #(
		.INIT('h1)
	) name1394 (
		_w1526_,
		_w1527_,
		_w1530_
	);
	LUT2 #(
		.INIT('h1)
	) name1395 (
		_w1528_,
		_w1529_,
		_w1531_
	);
	LUT2 #(
		.INIT('h8)
	) name1396 (
		_w1530_,
		_w1531_,
		_w1532_
	);
	LUT2 #(
		.INIT('h2)
	) name1397 (
		_w183_,
		_w1532_,
		_w1533_
	);
	LUT2 #(
		.INIT('h1)
	) name1398 (
		_w1509_,
		_w1517_,
		_w1534_
	);
	LUT2 #(
		.INIT('h1)
	) name1399 (
		_w1525_,
		_w1533_,
		_w1535_
	);
	LUT2 #(
		.INIT('h8)
	) name1400 (
		_w1534_,
		_w1535_,
		_w1536_
	);
	LUT2 #(
		.INIT('h2)
	) name1401 (
		\shift[6] ,
		_w1536_,
		_w1537_
	);
	LUT2 #(
		.INIT('h1)
	) name1402 (
		_w1501_,
		_w1537_,
		_w1538_
	);
	LUT2 #(
		.INIT('h2)
	) name1403 (
		_w136_,
		_w958_,
		_w1539_
	);
	LUT2 #(
		.INIT('h2)
	) name1404 (
		_w147_,
		_w930_,
		_w1540_
	);
	LUT2 #(
		.INIT('h2)
	) name1405 (
		_w158_,
		_w942_,
		_w1541_
	);
	LUT2 #(
		.INIT('h2)
	) name1406 (
		_w169_,
		_w934_,
		_w1542_
	);
	LUT2 #(
		.INIT('h1)
	) name1407 (
		_w1539_,
		_w1540_,
		_w1543_
	);
	LUT2 #(
		.INIT('h1)
	) name1408 (
		_w1541_,
		_w1542_,
		_w1544_
	);
	LUT2 #(
		.INIT('h8)
	) name1409 (
		_w1543_,
		_w1544_,
		_w1545_
	);
	LUT2 #(
		.INIT('h2)
	) name1410 (
		_w183_,
		_w1545_,
		_w1546_
	);
	LUT2 #(
		.INIT('h2)
	) name1411 (
		_w136_,
		_w998_,
		_w1547_
	);
	LUT2 #(
		.INIT('h2)
	) name1412 (
		_w147_,
		_w950_,
		_w1548_
	);
	LUT2 #(
		.INIT('h2)
	) name1413 (
		_w158_,
		_w962_,
		_w1549_
	);
	LUT2 #(
		.INIT('h2)
	) name1414 (
		_w169_,
		_w954_,
		_w1550_
	);
	LUT2 #(
		.INIT('h1)
	) name1415 (
		_w1547_,
		_w1548_,
		_w1551_
	);
	LUT2 #(
		.INIT('h1)
	) name1416 (
		_w1549_,
		_w1550_,
		_w1552_
	);
	LUT2 #(
		.INIT('h8)
	) name1417 (
		_w1551_,
		_w1552_,
		_w1553_
	);
	LUT2 #(
		.INIT('h2)
	) name1418 (
		_w228_,
		_w1553_,
		_w1554_
	);
	LUT2 #(
		.INIT('h2)
	) name1419 (
		_w136_,
		_w1042_,
		_w1555_
	);
	LUT2 #(
		.INIT('h2)
	) name1420 (
		_w147_,
		_w970_,
		_w1556_
	);
	LUT2 #(
		.INIT('h2)
	) name1421 (
		_w158_,
		_w982_,
		_w1557_
	);
	LUT2 #(
		.INIT('h2)
	) name1422 (
		_w169_,
		_w974_,
		_w1558_
	);
	LUT2 #(
		.INIT('h1)
	) name1423 (
		_w1555_,
		_w1556_,
		_w1559_
	);
	LUT2 #(
		.INIT('h1)
	) name1424 (
		_w1557_,
		_w1558_,
		_w1560_
	);
	LUT2 #(
		.INIT('h8)
	) name1425 (
		_w1559_,
		_w1560_,
		_w1561_
	);
	LUT2 #(
		.INIT('h2)
	) name1426 (
		_w273_,
		_w1561_,
		_w1562_
	);
	LUT2 #(
		.INIT('h2)
	) name1427 (
		_w136_,
		_w978_,
		_w1563_
	);
	LUT2 #(
		.INIT('h2)
	) name1428 (
		_w147_,
		_w990_,
		_w1564_
	);
	LUT2 #(
		.INIT('h2)
	) name1429 (
		_w158_,
		_w1002_,
		_w1565_
	);
	LUT2 #(
		.INIT('h2)
	) name1430 (
		_w169_,
		_w994_,
		_w1566_
	);
	LUT2 #(
		.INIT('h1)
	) name1431 (
		_w1563_,
		_w1564_,
		_w1567_
	);
	LUT2 #(
		.INIT('h1)
	) name1432 (
		_w1565_,
		_w1566_,
		_w1568_
	);
	LUT2 #(
		.INIT('h8)
	) name1433 (
		_w1567_,
		_w1568_,
		_w1569_
	);
	LUT2 #(
		.INIT('h2)
	) name1434 (
		_w318_,
		_w1569_,
		_w1570_
	);
	LUT2 #(
		.INIT('h1)
	) name1435 (
		_w1546_,
		_w1554_,
		_w1571_
	);
	LUT2 #(
		.INIT('h1)
	) name1436 (
		_w1562_,
		_w1570_,
		_w1572_
	);
	LUT2 #(
		.INIT('h8)
	) name1437 (
		_w1571_,
		_w1572_,
		_w1573_
	);
	LUT2 #(
		.INIT('h1)
	) name1438 (
		\shift[6] ,
		_w1573_,
		_w1574_
	);
	LUT2 #(
		.INIT('h2)
	) name1439 (
		_w136_,
		_w1022_,
		_w1575_
	);
	LUT2 #(
		.INIT('h2)
	) name1440 (
		_w147_,
		_w1054_,
		_w1576_
	);
	LUT2 #(
		.INIT('h2)
	) name1441 (
		_w158_,
		_w1068_,
		_w1577_
	);
	LUT2 #(
		.INIT('h2)
	) name1442 (
		_w169_,
		_w1058_,
		_w1578_
	);
	LUT2 #(
		.INIT('h1)
	) name1443 (
		_w1575_,
		_w1576_,
		_w1579_
	);
	LUT2 #(
		.INIT('h1)
	) name1444 (
		_w1577_,
		_w1578_,
		_w1580_
	);
	LUT2 #(
		.INIT('h8)
	) name1445 (
		_w1579_,
		_w1580_,
		_w1581_
	);
	LUT2 #(
		.INIT('h2)
	) name1446 (
		_w318_,
		_w1581_,
		_w1582_
	);
	LUT2 #(
		.INIT('h2)
	) name1447 (
		_w136_,
		_w938_,
		_w1583_
	);
	LUT2 #(
		.INIT('h2)
	) name1448 (
		_w147_,
		_w1014_,
		_w1584_
	);
	LUT2 #(
		.INIT('h2)
	) name1449 (
		_w158_,
		_w1026_,
		_w1585_
	);
	LUT2 #(
		.INIT('h2)
	) name1450 (
		_w169_,
		_w1018_,
		_w1586_
	);
	LUT2 #(
		.INIT('h1)
	) name1451 (
		_w1583_,
		_w1584_,
		_w1587_
	);
	LUT2 #(
		.INIT('h1)
	) name1452 (
		_w1585_,
		_w1586_,
		_w1588_
	);
	LUT2 #(
		.INIT('h8)
	) name1453 (
		_w1587_,
		_w1588_,
		_w1589_
	);
	LUT2 #(
		.INIT('h2)
	) name1454 (
		_w273_,
		_w1589_,
		_w1590_
	);
	LUT2 #(
		.INIT('h2)
	) name1455 (
		_w136_,
		_w1063_,
		_w1591_
	);
	LUT2 #(
		.INIT('h2)
	) name1456 (
		_w147_,
		_w1076_,
		_w1592_
	);
	LUT2 #(
		.INIT('h2)
	) name1457 (
		_w158_,
		_w1088_,
		_w1593_
	);
	LUT2 #(
		.INIT('h2)
	) name1458 (
		_w169_,
		_w1080_,
		_w1594_
	);
	LUT2 #(
		.INIT('h1)
	) name1459 (
		_w1591_,
		_w1592_,
		_w1595_
	);
	LUT2 #(
		.INIT('h1)
	) name1460 (
		_w1593_,
		_w1594_,
		_w1596_
	);
	LUT2 #(
		.INIT('h8)
	) name1461 (
		_w1595_,
		_w1596_,
		_w1597_
	);
	LUT2 #(
		.INIT('h2)
	) name1462 (
		_w228_,
		_w1597_,
		_w1598_
	);
	LUT2 #(
		.INIT('h2)
	) name1463 (
		_w136_,
		_w1084_,
		_w1599_
	);
	LUT2 #(
		.INIT('h2)
	) name1464 (
		_w147_,
		_w1034_,
		_w1600_
	);
	LUT2 #(
		.INIT('h2)
	) name1465 (
		_w158_,
		_w1046_,
		_w1601_
	);
	LUT2 #(
		.INIT('h2)
	) name1466 (
		_w169_,
		_w1038_,
		_w1602_
	);
	LUT2 #(
		.INIT('h1)
	) name1467 (
		_w1599_,
		_w1600_,
		_w1603_
	);
	LUT2 #(
		.INIT('h1)
	) name1468 (
		_w1601_,
		_w1602_,
		_w1604_
	);
	LUT2 #(
		.INIT('h8)
	) name1469 (
		_w1603_,
		_w1604_,
		_w1605_
	);
	LUT2 #(
		.INIT('h2)
	) name1470 (
		_w183_,
		_w1605_,
		_w1606_
	);
	LUT2 #(
		.INIT('h1)
	) name1471 (
		_w1582_,
		_w1590_,
		_w1607_
	);
	LUT2 #(
		.INIT('h1)
	) name1472 (
		_w1598_,
		_w1606_,
		_w1608_
	);
	LUT2 #(
		.INIT('h8)
	) name1473 (
		_w1607_,
		_w1608_,
		_w1609_
	);
	LUT2 #(
		.INIT('h2)
	) name1474 (
		\shift[6] ,
		_w1609_,
		_w1610_
	);
	LUT2 #(
		.INIT('h1)
	) name1475 (
		_w1574_,
		_w1610_,
		_w1611_
	);
	LUT2 #(
		.INIT('h2)
	) name1476 (
		_w136_,
		_w1157_,
		_w1612_
	);
	LUT2 #(
		.INIT('h2)
	) name1477 (
		_w147_,
		_w1213_,
		_w1613_
	);
	LUT2 #(
		.INIT('h2)
	) name1478 (
		_w158_,
		_w1237_,
		_w1614_
	);
	LUT2 #(
		.INIT('h2)
	) name1479 (
		_w169_,
		_w1221_,
		_w1615_
	);
	LUT2 #(
		.INIT('h1)
	) name1480 (
		_w1612_,
		_w1613_,
		_w1616_
	);
	LUT2 #(
		.INIT('h1)
	) name1481 (
		_w1614_,
		_w1615_,
		_w1617_
	);
	LUT2 #(
		.INIT('h8)
	) name1482 (
		_w1616_,
		_w1617_,
		_w1618_
	);
	LUT2 #(
		.INIT('h2)
	) name1483 (
		_w183_,
		_w1618_,
		_w1619_
	);
	LUT2 #(
		.INIT('h2)
	) name1484 (
		_w136_,
		_w1121_,
		_w1620_
	);
	LUT2 #(
		.INIT('h2)
	) name1485 (
		_w147_,
		_w1141_,
		_w1621_
	);
	LUT2 #(
		.INIT('h2)
	) name1486 (
		_w158_,
		_w1165_,
		_w1622_
	);
	LUT2 #(
		.INIT('h2)
	) name1487 (
		_w169_,
		_w1149_,
		_w1623_
	);
	LUT2 #(
		.INIT('h1)
	) name1488 (
		_w1620_,
		_w1621_,
		_w1624_
	);
	LUT2 #(
		.INIT('h1)
	) name1489 (
		_w1622_,
		_w1623_,
		_w1625_
	);
	LUT2 #(
		.INIT('h8)
	) name1490 (
		_w1624_,
		_w1625_,
		_w1626_
	);
	LUT2 #(
		.INIT('h2)
	) name1491 (
		_w228_,
		_w1626_,
		_w1627_
	);
	LUT2 #(
		.INIT('h2)
	) name1492 (
		_w136_,
		_w1338_,
		_w1628_
	);
	LUT2 #(
		.INIT('h2)
	) name1493 (
		_w147_,
		_w1177_,
		_w1629_
	);
	LUT2 #(
		.INIT('h2)
	) name1494 (
		_w158_,
		_w1201_,
		_w1630_
	);
	LUT2 #(
		.INIT('h2)
	) name1495 (
		_w169_,
		_w1185_,
		_w1631_
	);
	LUT2 #(
		.INIT('h1)
	) name1496 (
		_w1628_,
		_w1629_,
		_w1632_
	);
	LUT2 #(
		.INIT('h1)
	) name1497 (
		_w1630_,
		_w1631_,
		_w1633_
	);
	LUT2 #(
		.INIT('h8)
	) name1498 (
		_w1632_,
		_w1633_,
		_w1634_
	);
	LUT2 #(
		.INIT('h2)
	) name1499 (
		_w273_,
		_w1634_,
		_w1635_
	);
	LUT2 #(
		.INIT('h2)
	) name1500 (
		_w136_,
		_w1193_,
		_w1636_
	);
	LUT2 #(
		.INIT('h2)
	) name1501 (
		_w147_,
		_w1105_,
		_w1637_
	);
	LUT2 #(
		.INIT('h2)
	) name1502 (
		_w158_,
		_w1129_,
		_w1638_
	);
	LUT2 #(
		.INIT('h2)
	) name1503 (
		_w169_,
		_w1113_,
		_w1639_
	);
	LUT2 #(
		.INIT('h1)
	) name1504 (
		_w1636_,
		_w1637_,
		_w1640_
	);
	LUT2 #(
		.INIT('h1)
	) name1505 (
		_w1638_,
		_w1639_,
		_w1641_
	);
	LUT2 #(
		.INIT('h8)
	) name1506 (
		_w1640_,
		_w1641_,
		_w1642_
	);
	LUT2 #(
		.INIT('h2)
	) name1507 (
		_w318_,
		_w1642_,
		_w1643_
	);
	LUT2 #(
		.INIT('h1)
	) name1508 (
		_w1619_,
		_w1627_,
		_w1644_
	);
	LUT2 #(
		.INIT('h1)
	) name1509 (
		_w1635_,
		_w1643_,
		_w1645_
	);
	LUT2 #(
		.INIT('h8)
	) name1510 (
		_w1644_,
		_w1645_,
		_w1646_
	);
	LUT2 #(
		.INIT('h1)
	) name1511 (
		\shift[6] ,
		_w1646_,
		_w1647_
	);
	LUT2 #(
		.INIT('h2)
	) name1512 (
		_w147_,
		_w1289_,
		_w1648_
	);
	LUT2 #(
		.INIT('h2)
	) name1513 (
		_w169_,
		_w1294_,
		_w1649_
	);
	LUT2 #(
		.INIT('h2)
	) name1514 (
		_w158_,
		_w1310_,
		_w1650_
	);
	LUT2 #(
		.INIT('h2)
	) name1515 (
		_w136_,
		_w1269_,
		_w1651_
	);
	LUT2 #(
		.INIT('h1)
	) name1516 (
		_w1648_,
		_w1649_,
		_w1652_
	);
	LUT2 #(
		.INIT('h1)
	) name1517 (
		_w1650_,
		_w1651_,
		_w1653_
	);
	LUT2 #(
		.INIT('h8)
	) name1518 (
		_w1652_,
		_w1653_,
		_w1654_
	);
	LUT2 #(
		.INIT('h2)
	) name1519 (
		_w318_,
		_w1654_,
		_w1655_
	);
	LUT2 #(
		.INIT('h2)
	) name1520 (
		_w136_,
		_w1229_,
		_w1656_
	);
	LUT2 #(
		.INIT('h2)
	) name1521 (
		_w147_,
		_w1253_,
		_w1657_
	);
	LUT2 #(
		.INIT('h2)
	) name1522 (
		_w158_,
		_w1277_,
		_w1658_
	);
	LUT2 #(
		.INIT('h2)
	) name1523 (
		_w169_,
		_w1261_,
		_w1659_
	);
	LUT2 #(
		.INIT('h1)
	) name1524 (
		_w1656_,
		_w1657_,
		_w1660_
	);
	LUT2 #(
		.INIT('h1)
	) name1525 (
		_w1658_,
		_w1659_,
		_w1661_
	);
	LUT2 #(
		.INIT('h8)
	) name1526 (
		_w1660_,
		_w1661_,
		_w1662_
	);
	LUT2 #(
		.INIT('h2)
	) name1527 (
		_w273_,
		_w1662_,
		_w1663_
	);
	LUT2 #(
		.INIT('h2)
	) name1528 (
		_w136_,
		_w1302_,
		_w1664_
	);
	LUT2 #(
		.INIT('h2)
	) name1529 (
		_w147_,
		_w1358_,
		_w1665_
	);
	LUT2 #(
		.INIT('h2)
	) name1530 (
		_w158_,
		_w1382_,
		_w1666_
	);
	LUT2 #(
		.INIT('h2)
	) name1531 (
		_w169_,
		_w1366_,
		_w1667_
	);
	LUT2 #(
		.INIT('h1)
	) name1532 (
		_w1664_,
		_w1665_,
		_w1668_
	);
	LUT2 #(
		.INIT('h1)
	) name1533 (
		_w1666_,
		_w1667_,
		_w1669_
	);
	LUT2 #(
		.INIT('h8)
	) name1534 (
		_w1668_,
		_w1669_,
		_w1670_
	);
	LUT2 #(
		.INIT('h2)
	) name1535 (
		_w228_,
		_w1670_,
		_w1671_
	);
	LUT2 #(
		.INIT('h2)
	) name1536 (
		_w136_,
		_w1374_,
		_w1672_
	);
	LUT2 #(
		.INIT('h2)
	) name1537 (
		_w147_,
		_w1322_,
		_w1673_
	);
	LUT2 #(
		.INIT('h2)
	) name1538 (
		_w158_,
		_w1346_,
		_w1674_
	);
	LUT2 #(
		.INIT('h2)
	) name1539 (
		_w169_,
		_w1330_,
		_w1675_
	);
	LUT2 #(
		.INIT('h1)
	) name1540 (
		_w1672_,
		_w1673_,
		_w1676_
	);
	LUT2 #(
		.INIT('h1)
	) name1541 (
		_w1674_,
		_w1675_,
		_w1677_
	);
	LUT2 #(
		.INIT('h8)
	) name1542 (
		_w1676_,
		_w1677_,
		_w1678_
	);
	LUT2 #(
		.INIT('h2)
	) name1543 (
		_w183_,
		_w1678_,
		_w1679_
	);
	LUT2 #(
		.INIT('h1)
	) name1544 (
		_w1655_,
		_w1663_,
		_w1680_
	);
	LUT2 #(
		.INIT('h1)
	) name1545 (
		_w1671_,
		_w1679_,
		_w1681_
	);
	LUT2 #(
		.INIT('h8)
	) name1546 (
		_w1680_,
		_w1681_,
		_w1682_
	);
	LUT2 #(
		.INIT('h2)
	) name1547 (
		\shift[6] ,
		_w1682_,
		_w1683_
	);
	LUT2 #(
		.INIT('h1)
	) name1548 (
		_w1647_,
		_w1683_,
		_w1684_
	);
	LUT2 #(
		.INIT('h2)
	) name1549 (
		_w136_,
		_w223_,
		_w1685_
	);
	LUT2 #(
		.INIT('h2)
	) name1550 (
		_w147_,
		_w213_,
		_w1686_
	);
	LUT2 #(
		.INIT('h4)
	) name1551 (
		_w156_,
		_w158_,
		_w1687_
	);
	LUT2 #(
		.INIT('h4)
	) name1552 (
		_w145_,
		_w169_,
		_w1688_
	);
	LUT2 #(
		.INIT('h1)
	) name1553 (
		_w1685_,
		_w1686_,
		_w1689_
	);
	LUT2 #(
		.INIT('h1)
	) name1554 (
		_w1687_,
		_w1688_,
		_w1690_
	);
	LUT2 #(
		.INIT('h8)
	) name1555 (
		_w1689_,
		_w1690_,
		_w1691_
	);
	LUT2 #(
		.INIT('h2)
	) name1556 (
		_w183_,
		_w1691_,
		_w1692_
	);
	LUT2 #(
		.INIT('h2)
	) name1557 (
		_w136_,
		_w313_,
		_w1693_
	);
	LUT2 #(
		.INIT('h2)
	) name1558 (
		_w147_,
		_w303_,
		_w1694_
	);
	LUT2 #(
		.INIT('h2)
	) name1559 (
		_w158_,
		_w203_,
		_w1695_
	);
	LUT2 #(
		.INIT('h2)
	) name1560 (
		_w169_,
		_w193_,
		_w1696_
	);
	LUT2 #(
		.INIT('h1)
	) name1561 (
		_w1693_,
		_w1694_,
		_w1697_
	);
	LUT2 #(
		.INIT('h1)
	) name1562 (
		_w1695_,
		_w1696_,
		_w1698_
	);
	LUT2 #(
		.INIT('h8)
	) name1563 (
		_w1697_,
		_w1698_,
		_w1699_
	);
	LUT2 #(
		.INIT('h2)
	) name1564 (
		_w228_,
		_w1699_,
		_w1700_
	);
	LUT2 #(
		.INIT('h2)
	) name1565 (
		_w136_,
		_w362_,
		_w1701_
	);
	LUT2 #(
		.INIT('h2)
	) name1566 (
		_w147_,
		_w352_,
		_w1702_
	);
	LUT2 #(
		.INIT('h2)
	) name1567 (
		_w158_,
		_w248_,
		_w1703_
	);
	LUT2 #(
		.INIT('h2)
	) name1568 (
		_w169_,
		_w238_,
		_w1704_
	);
	LUT2 #(
		.INIT('h1)
	) name1569 (
		_w1701_,
		_w1702_,
		_w1705_
	);
	LUT2 #(
		.INIT('h1)
	) name1570 (
		_w1703_,
		_w1704_,
		_w1706_
	);
	LUT2 #(
		.INIT('h8)
	) name1571 (
		_w1705_,
		_w1706_,
		_w1707_
	);
	LUT2 #(
		.INIT('h2)
	) name1572 (
		_w273_,
		_w1707_,
		_w1708_
	);
	LUT2 #(
		.INIT('h2)
	) name1573 (
		_w136_,
		_w268_,
		_w1709_
	);
	LUT2 #(
		.INIT('h2)
	) name1574 (
		_w147_,
		_w258_,
		_w1710_
	);
	LUT2 #(
		.INIT('h2)
	) name1575 (
		_w158_,
		_w293_,
		_w1711_
	);
	LUT2 #(
		.INIT('h2)
	) name1576 (
		_w169_,
		_w283_,
		_w1712_
	);
	LUT2 #(
		.INIT('h1)
	) name1577 (
		_w1709_,
		_w1710_,
		_w1713_
	);
	LUT2 #(
		.INIT('h1)
	) name1578 (
		_w1711_,
		_w1712_,
		_w1714_
	);
	LUT2 #(
		.INIT('h8)
	) name1579 (
		_w1713_,
		_w1714_,
		_w1715_
	);
	LUT2 #(
		.INIT('h2)
	) name1580 (
		_w318_,
		_w1715_,
		_w1716_
	);
	LUT2 #(
		.INIT('h1)
	) name1581 (
		_w1692_,
		_w1700_,
		_w1717_
	);
	LUT2 #(
		.INIT('h1)
	) name1582 (
		_w1708_,
		_w1716_,
		_w1718_
	);
	LUT2 #(
		.INIT('h8)
	) name1583 (
		_w1717_,
		_w1718_,
		_w1719_
	);
	LUT2 #(
		.INIT('h1)
	) name1584 (
		\shift[6] ,
		_w1719_,
		_w1720_
	);
	LUT2 #(
		.INIT('h2)
	) name1585 (
		_w136_,
		_w450_,
		_w1721_
	);
	LUT2 #(
		.INIT('h2)
	) name1586 (
		_w147_,
		_w440_,
		_w1722_
	);
	LUT2 #(
		.INIT('h2)
	) name1587 (
		_w158_,
		_w474_,
		_w1723_
	);
	LUT2 #(
		.INIT('h2)
	) name1588 (
		_w169_,
		_w464_,
		_w1724_
	);
	LUT2 #(
		.INIT('h1)
	) name1589 (
		_w1721_,
		_w1722_,
		_w1725_
	);
	LUT2 #(
		.INIT('h1)
	) name1590 (
		_w1723_,
		_w1724_,
		_w1726_
	);
	LUT2 #(
		.INIT('h8)
	) name1591 (
		_w1725_,
		_w1726_,
		_w1727_
	);
	LUT2 #(
		.INIT('h2)
	) name1592 (
		_w318_,
		_w1727_,
		_w1728_
	);
	LUT2 #(
		.INIT('h2)
	) name1593 (
		_w136_,
		_w178_,
		_w1729_
	);
	LUT2 #(
		.INIT('h2)
	) name1594 (
		_w147_,
		_w167_,
		_w1730_
	);
	LUT2 #(
		.INIT('h2)
	) name1595 (
		_w158_,
		_w430_,
		_w1731_
	);
	LUT2 #(
		.INIT('h2)
	) name1596 (
		_w169_,
		_w420_,
		_w1732_
	);
	LUT2 #(
		.INIT('h1)
	) name1597 (
		_w1729_,
		_w1730_,
		_w1733_
	);
	LUT2 #(
		.INIT('h1)
	) name1598 (
		_w1731_,
		_w1732_,
		_w1734_
	);
	LUT2 #(
		.INIT('h8)
	) name1599 (
		_w1733_,
		_w1734_,
		_w1735_
	);
	LUT2 #(
		.INIT('h2)
	) name1600 (
		_w273_,
		_w1735_,
		_w1736_
	);
	LUT2 #(
		.INIT('h2)
	) name1601 (
		_w136_,
		_w496_,
		_w1737_
	);
	LUT2 #(
		.INIT('h2)
	) name1602 (
		_w147_,
		_w484_,
		_w1738_
	);
	LUT2 #(
		.INIT('h2)
	) name1603 (
		_w158_,
		_w386_,
		_w1739_
	);
	LUT2 #(
		.INIT('h2)
	) name1604 (
		_w169_,
		_w376_,
		_w1740_
	);
	LUT2 #(
		.INIT('h1)
	) name1605 (
		_w1737_,
		_w1738_,
		_w1741_
	);
	LUT2 #(
		.INIT('h1)
	) name1606 (
		_w1739_,
		_w1740_,
		_w1742_
	);
	LUT2 #(
		.INIT('h8)
	) name1607 (
		_w1741_,
		_w1742_,
		_w1743_
	);
	LUT2 #(
		.INIT('h2)
	) name1608 (
		_w228_,
		_w1743_,
		_w1744_
	);
	LUT2 #(
		.INIT('h2)
	) name1609 (
		_w136_,
		_w406_,
		_w1745_
	);
	LUT2 #(
		.INIT('h2)
	) name1610 (
		_w147_,
		_w396_,
		_w1746_
	);
	LUT2 #(
		.INIT('h2)
	) name1611 (
		_w158_,
		_w342_,
		_w1747_
	);
	LUT2 #(
		.INIT('h2)
	) name1612 (
		_w169_,
		_w332_,
		_w1748_
	);
	LUT2 #(
		.INIT('h1)
	) name1613 (
		_w1745_,
		_w1746_,
		_w1749_
	);
	LUT2 #(
		.INIT('h1)
	) name1614 (
		_w1747_,
		_w1748_,
		_w1750_
	);
	LUT2 #(
		.INIT('h8)
	) name1615 (
		_w1749_,
		_w1750_,
		_w1751_
	);
	LUT2 #(
		.INIT('h2)
	) name1616 (
		_w183_,
		_w1751_,
		_w1752_
	);
	LUT2 #(
		.INIT('h1)
	) name1617 (
		_w1728_,
		_w1736_,
		_w1753_
	);
	LUT2 #(
		.INIT('h1)
	) name1618 (
		_w1744_,
		_w1752_,
		_w1754_
	);
	LUT2 #(
		.INIT('h8)
	) name1619 (
		_w1753_,
		_w1754_,
		_w1755_
	);
	LUT2 #(
		.INIT('h2)
	) name1620 (
		\shift[6] ,
		_w1755_,
		_w1756_
	);
	LUT2 #(
		.INIT('h1)
	) name1621 (
		_w1720_,
		_w1756_,
		_w1757_
	);
	LUT2 #(
		.INIT('h2)
	) name1622 (
		_w136_,
		_w605_,
		_w1758_
	);
	LUT2 #(
		.INIT('h2)
	) name1623 (
		_w147_,
		_w593_,
		_w1759_
	);
	LUT2 #(
		.INIT('h2)
	) name1624 (
		_w158_,
		_w529_,
		_w1760_
	);
	LUT2 #(
		.INIT('h2)
	) name1625 (
		_w169_,
		_w517_,
		_w1761_
	);
	LUT2 #(
		.INIT('h1)
	) name1626 (
		_w1758_,
		_w1759_,
		_w1762_
	);
	LUT2 #(
		.INIT('h1)
	) name1627 (
		_w1760_,
		_w1761_,
		_w1763_
	);
	LUT2 #(
		.INIT('h8)
	) name1628 (
		_w1762_,
		_w1763_,
		_w1764_
	);
	LUT2 #(
		.INIT('h2)
	) name1629 (
		_w183_,
		_w1764_,
		_w1765_
	);
	LUT2 #(
		.INIT('h2)
	) name1630 (
		_w136_,
		_w709_,
		_w1766_
	);
	LUT2 #(
		.INIT('h2)
	) name1631 (
		_w147_,
		_w697_,
		_w1767_
	);
	LUT2 #(
		.INIT('h2)
	) name1632 (
		_w158_,
		_w581_,
		_w1768_
	);
	LUT2 #(
		.INIT('h2)
	) name1633 (
		_w169_,
		_w569_,
		_w1769_
	);
	LUT2 #(
		.INIT('h1)
	) name1634 (
		_w1766_,
		_w1767_,
		_w1770_
	);
	LUT2 #(
		.INIT('h1)
	) name1635 (
		_w1768_,
		_w1769_,
		_w1771_
	);
	LUT2 #(
		.INIT('h8)
	) name1636 (
		_w1770_,
		_w1771_,
		_w1772_
	);
	LUT2 #(
		.INIT('h2)
	) name1637 (
		_w228_,
		_w1772_,
		_w1773_
	);
	LUT2 #(
		.INIT('h2)
	) name1638 (
		_w136_,
		_w817_,
		_w1774_
	);
	LUT2 #(
		.INIT('h2)
	) name1639 (
		_w147_,
		_w805_,
		_w1775_
	);
	LUT2 #(
		.INIT('h2)
	) name1640 (
		_w158_,
		_w633_,
		_w1776_
	);
	LUT2 #(
		.INIT('h2)
	) name1641 (
		_w169_,
		_w621_,
		_w1777_
	);
	LUT2 #(
		.INIT('h1)
	) name1642 (
		_w1774_,
		_w1775_,
		_w1778_
	);
	LUT2 #(
		.INIT('h1)
	) name1643 (
		_w1776_,
		_w1777_,
		_w1779_
	);
	LUT2 #(
		.INIT('h8)
	) name1644 (
		_w1778_,
		_w1779_,
		_w1780_
	);
	LUT2 #(
		.INIT('h2)
	) name1645 (
		_w273_,
		_w1780_,
		_w1781_
	);
	LUT2 #(
		.INIT('h2)
	) name1646 (
		_w136_,
		_w657_,
		_w1782_
	);
	LUT2 #(
		.INIT('h2)
	) name1647 (
		_w147_,
		_w645_,
		_w1783_
	);
	LUT2 #(
		.INIT('h2)
	) name1648 (
		_w158_,
		_w685_,
		_w1784_
	);
	LUT2 #(
		.INIT('h2)
	) name1649 (
		_w169_,
		_w673_,
		_w1785_
	);
	LUT2 #(
		.INIT('h1)
	) name1650 (
		_w1782_,
		_w1783_,
		_w1786_
	);
	LUT2 #(
		.INIT('h1)
	) name1651 (
		_w1784_,
		_w1785_,
		_w1787_
	);
	LUT2 #(
		.INIT('h8)
	) name1652 (
		_w1786_,
		_w1787_,
		_w1788_
	);
	LUT2 #(
		.INIT('h2)
	) name1653 (
		_w318_,
		_w1788_,
		_w1789_
	);
	LUT2 #(
		.INIT('h1)
	) name1654 (
		_w1765_,
		_w1773_,
		_w1790_
	);
	LUT2 #(
		.INIT('h1)
	) name1655 (
		_w1781_,
		_w1789_,
		_w1791_
	);
	LUT2 #(
		.INIT('h8)
	) name1656 (
		_w1790_,
		_w1791_,
		_w1792_
	);
	LUT2 #(
		.INIT('h1)
	) name1657 (
		\shift[6] ,
		_w1792_,
		_w1793_
	);
	LUT2 #(
		.INIT('h2)
	) name1658 (
		_w136_,
		_w765_,
		_w1794_
	);
	LUT2 #(
		.INIT('h2)
	) name1659 (
		_w147_,
		_w753_,
		_w1795_
	);
	LUT2 #(
		.INIT('h2)
	) name1660 (
		_w158_,
		_w843_,
		_w1796_
	);
	LUT2 #(
		.INIT('h2)
	) name1661 (
		_w169_,
		_w833_,
		_w1797_
	);
	LUT2 #(
		.INIT('h1)
	) name1662 (
		_w1794_,
		_w1795_,
		_w1798_
	);
	LUT2 #(
		.INIT('h1)
	) name1663 (
		_w1796_,
		_w1797_,
		_w1799_
	);
	LUT2 #(
		.INIT('h8)
	) name1664 (
		_w1798_,
		_w1799_,
		_w1800_
	);
	LUT2 #(
		.INIT('h2)
	) name1665 (
		_w318_,
		_w1800_,
		_w1801_
	);
	LUT2 #(
		.INIT('h2)
	) name1666 (
		_w136_,
		_w553_,
		_w1802_
	);
	LUT2 #(
		.INIT('h2)
	) name1667 (
		_w147_,
		_w541_,
		_w1803_
	);
	LUT2 #(
		.INIT('h2)
	) name1668 (
		_w158_,
		_w741_,
		_w1804_
	);
	LUT2 #(
		.INIT('h2)
	) name1669 (
		_w169_,
		_w729_,
		_w1805_
	);
	LUT2 #(
		.INIT('h1)
	) name1670 (
		_w1802_,
		_w1803_,
		_w1806_
	);
	LUT2 #(
		.INIT('h1)
	) name1671 (
		_w1804_,
		_w1805_,
		_w1807_
	);
	LUT2 #(
		.INIT('h8)
	) name1672 (
		_w1806_,
		_w1807_,
		_w1808_
	);
	LUT2 #(
		.INIT('h2)
	) name1673 (
		_w273_,
		_w1808_,
		_w1809_
	);
	LUT2 #(
		.INIT('h2)
	) name1674 (
		_w136_,
		_w865_,
		_w1810_
	);
	LUT2 #(
		.INIT('h2)
	) name1675 (
		_w147_,
		_w855_,
		_w1811_
	);
	LUT2 #(
		.INIT('h2)
	) name1676 (
		_w158_,
		_w893_,
		_w1812_
	);
	LUT2 #(
		.INIT('h2)
	) name1677 (
		_w169_,
		_w881_,
		_w1813_
	);
	LUT2 #(
		.INIT('h1)
	) name1678 (
		_w1810_,
		_w1811_,
		_w1814_
	);
	LUT2 #(
		.INIT('h1)
	) name1679 (
		_w1812_,
		_w1813_,
		_w1815_
	);
	LUT2 #(
		.INIT('h8)
	) name1680 (
		_w1814_,
		_w1815_,
		_w1816_
	);
	LUT2 #(
		.INIT('h2)
	) name1681 (
		_w228_,
		_w1816_,
		_w1817_
	);
	LUT2 #(
		.INIT('h2)
	) name1682 (
		_w136_,
		_w917_,
		_w1818_
	);
	LUT2 #(
		.INIT('h2)
	) name1683 (
		_w147_,
		_w905_,
		_w1819_
	);
	LUT2 #(
		.INIT('h2)
	) name1684 (
		_w158_,
		_w793_,
		_w1820_
	);
	LUT2 #(
		.INIT('h2)
	) name1685 (
		_w169_,
		_w781_,
		_w1821_
	);
	LUT2 #(
		.INIT('h1)
	) name1686 (
		_w1818_,
		_w1819_,
		_w1822_
	);
	LUT2 #(
		.INIT('h1)
	) name1687 (
		_w1820_,
		_w1821_,
		_w1823_
	);
	LUT2 #(
		.INIT('h8)
	) name1688 (
		_w1822_,
		_w1823_,
		_w1824_
	);
	LUT2 #(
		.INIT('h2)
	) name1689 (
		_w183_,
		_w1824_,
		_w1825_
	);
	LUT2 #(
		.INIT('h1)
	) name1690 (
		_w1801_,
		_w1809_,
		_w1826_
	);
	LUT2 #(
		.INIT('h1)
	) name1691 (
		_w1817_,
		_w1825_,
		_w1827_
	);
	LUT2 #(
		.INIT('h8)
	) name1692 (
		_w1826_,
		_w1827_,
		_w1828_
	);
	LUT2 #(
		.INIT('h2)
	) name1693 (
		\shift[6] ,
		_w1828_,
		_w1829_
	);
	LUT2 #(
		.INIT('h1)
	) name1694 (
		_w1793_,
		_w1829_,
		_w1830_
	);
	LUT2 #(
		.INIT('h2)
	) name1695 (
		_w136_,
		_w962_,
		_w1831_
	);
	LUT2 #(
		.INIT('h2)
	) name1696 (
		_w147_,
		_w958_,
		_w1832_
	);
	LUT2 #(
		.INIT('h2)
	) name1697 (
		_w158_,
		_w934_,
		_w1833_
	);
	LUT2 #(
		.INIT('h2)
	) name1698 (
		_w169_,
		_w930_,
		_w1834_
	);
	LUT2 #(
		.INIT('h1)
	) name1699 (
		_w1831_,
		_w1832_,
		_w1835_
	);
	LUT2 #(
		.INIT('h1)
	) name1700 (
		_w1833_,
		_w1834_,
		_w1836_
	);
	LUT2 #(
		.INIT('h8)
	) name1701 (
		_w1835_,
		_w1836_,
		_w1837_
	);
	LUT2 #(
		.INIT('h2)
	) name1702 (
		_w183_,
		_w1837_,
		_w1838_
	);
	LUT2 #(
		.INIT('h2)
	) name1703 (
		_w136_,
		_w1002_,
		_w1839_
	);
	LUT2 #(
		.INIT('h2)
	) name1704 (
		_w147_,
		_w998_,
		_w1840_
	);
	LUT2 #(
		.INIT('h2)
	) name1705 (
		_w158_,
		_w954_,
		_w1841_
	);
	LUT2 #(
		.INIT('h2)
	) name1706 (
		_w169_,
		_w950_,
		_w1842_
	);
	LUT2 #(
		.INIT('h1)
	) name1707 (
		_w1839_,
		_w1840_,
		_w1843_
	);
	LUT2 #(
		.INIT('h1)
	) name1708 (
		_w1841_,
		_w1842_,
		_w1844_
	);
	LUT2 #(
		.INIT('h8)
	) name1709 (
		_w1843_,
		_w1844_,
		_w1845_
	);
	LUT2 #(
		.INIT('h2)
	) name1710 (
		_w228_,
		_w1845_,
		_w1846_
	);
	LUT2 #(
		.INIT('h2)
	) name1711 (
		_w136_,
		_w1046_,
		_w1847_
	);
	LUT2 #(
		.INIT('h2)
	) name1712 (
		_w147_,
		_w1042_,
		_w1848_
	);
	LUT2 #(
		.INIT('h2)
	) name1713 (
		_w158_,
		_w974_,
		_w1849_
	);
	LUT2 #(
		.INIT('h2)
	) name1714 (
		_w169_,
		_w970_,
		_w1850_
	);
	LUT2 #(
		.INIT('h1)
	) name1715 (
		_w1847_,
		_w1848_,
		_w1851_
	);
	LUT2 #(
		.INIT('h1)
	) name1716 (
		_w1849_,
		_w1850_,
		_w1852_
	);
	LUT2 #(
		.INIT('h8)
	) name1717 (
		_w1851_,
		_w1852_,
		_w1853_
	);
	LUT2 #(
		.INIT('h2)
	) name1718 (
		_w273_,
		_w1853_,
		_w1854_
	);
	LUT2 #(
		.INIT('h2)
	) name1719 (
		_w136_,
		_w982_,
		_w1855_
	);
	LUT2 #(
		.INIT('h2)
	) name1720 (
		_w147_,
		_w978_,
		_w1856_
	);
	LUT2 #(
		.INIT('h2)
	) name1721 (
		_w158_,
		_w994_,
		_w1857_
	);
	LUT2 #(
		.INIT('h2)
	) name1722 (
		_w169_,
		_w990_,
		_w1858_
	);
	LUT2 #(
		.INIT('h1)
	) name1723 (
		_w1855_,
		_w1856_,
		_w1859_
	);
	LUT2 #(
		.INIT('h1)
	) name1724 (
		_w1857_,
		_w1858_,
		_w1860_
	);
	LUT2 #(
		.INIT('h8)
	) name1725 (
		_w1859_,
		_w1860_,
		_w1861_
	);
	LUT2 #(
		.INIT('h2)
	) name1726 (
		_w318_,
		_w1861_,
		_w1862_
	);
	LUT2 #(
		.INIT('h1)
	) name1727 (
		_w1838_,
		_w1846_,
		_w1863_
	);
	LUT2 #(
		.INIT('h1)
	) name1728 (
		_w1854_,
		_w1862_,
		_w1864_
	);
	LUT2 #(
		.INIT('h8)
	) name1729 (
		_w1863_,
		_w1864_,
		_w1865_
	);
	LUT2 #(
		.INIT('h1)
	) name1730 (
		\shift[6] ,
		_w1865_,
		_w1866_
	);
	LUT2 #(
		.INIT('h2)
	) name1731 (
		_w136_,
		_w1026_,
		_w1867_
	);
	LUT2 #(
		.INIT('h2)
	) name1732 (
		_w147_,
		_w1022_,
		_w1868_
	);
	LUT2 #(
		.INIT('h2)
	) name1733 (
		_w158_,
		_w1058_,
		_w1869_
	);
	LUT2 #(
		.INIT('h2)
	) name1734 (
		_w169_,
		_w1054_,
		_w1870_
	);
	LUT2 #(
		.INIT('h1)
	) name1735 (
		_w1867_,
		_w1868_,
		_w1871_
	);
	LUT2 #(
		.INIT('h1)
	) name1736 (
		_w1869_,
		_w1870_,
		_w1872_
	);
	LUT2 #(
		.INIT('h8)
	) name1737 (
		_w1871_,
		_w1872_,
		_w1873_
	);
	LUT2 #(
		.INIT('h2)
	) name1738 (
		_w318_,
		_w1873_,
		_w1874_
	);
	LUT2 #(
		.INIT('h2)
	) name1739 (
		_w136_,
		_w942_,
		_w1875_
	);
	LUT2 #(
		.INIT('h2)
	) name1740 (
		_w147_,
		_w938_,
		_w1876_
	);
	LUT2 #(
		.INIT('h2)
	) name1741 (
		_w158_,
		_w1018_,
		_w1877_
	);
	LUT2 #(
		.INIT('h2)
	) name1742 (
		_w169_,
		_w1014_,
		_w1878_
	);
	LUT2 #(
		.INIT('h1)
	) name1743 (
		_w1875_,
		_w1876_,
		_w1879_
	);
	LUT2 #(
		.INIT('h1)
	) name1744 (
		_w1877_,
		_w1878_,
		_w1880_
	);
	LUT2 #(
		.INIT('h8)
	) name1745 (
		_w1879_,
		_w1880_,
		_w1881_
	);
	LUT2 #(
		.INIT('h2)
	) name1746 (
		_w273_,
		_w1881_,
		_w1882_
	);
	LUT2 #(
		.INIT('h2)
	) name1747 (
		_w136_,
		_w1068_,
		_w1883_
	);
	LUT2 #(
		.INIT('h2)
	) name1748 (
		_w147_,
		_w1063_,
		_w1884_
	);
	LUT2 #(
		.INIT('h2)
	) name1749 (
		_w158_,
		_w1080_,
		_w1885_
	);
	LUT2 #(
		.INIT('h2)
	) name1750 (
		_w169_,
		_w1076_,
		_w1886_
	);
	LUT2 #(
		.INIT('h1)
	) name1751 (
		_w1883_,
		_w1884_,
		_w1887_
	);
	LUT2 #(
		.INIT('h1)
	) name1752 (
		_w1885_,
		_w1886_,
		_w1888_
	);
	LUT2 #(
		.INIT('h8)
	) name1753 (
		_w1887_,
		_w1888_,
		_w1889_
	);
	LUT2 #(
		.INIT('h2)
	) name1754 (
		_w228_,
		_w1889_,
		_w1890_
	);
	LUT2 #(
		.INIT('h2)
	) name1755 (
		_w136_,
		_w1088_,
		_w1891_
	);
	LUT2 #(
		.INIT('h2)
	) name1756 (
		_w147_,
		_w1084_,
		_w1892_
	);
	LUT2 #(
		.INIT('h2)
	) name1757 (
		_w158_,
		_w1038_,
		_w1893_
	);
	LUT2 #(
		.INIT('h2)
	) name1758 (
		_w169_,
		_w1034_,
		_w1894_
	);
	LUT2 #(
		.INIT('h1)
	) name1759 (
		_w1891_,
		_w1892_,
		_w1895_
	);
	LUT2 #(
		.INIT('h1)
	) name1760 (
		_w1893_,
		_w1894_,
		_w1896_
	);
	LUT2 #(
		.INIT('h8)
	) name1761 (
		_w1895_,
		_w1896_,
		_w1897_
	);
	LUT2 #(
		.INIT('h2)
	) name1762 (
		_w183_,
		_w1897_,
		_w1898_
	);
	LUT2 #(
		.INIT('h1)
	) name1763 (
		_w1874_,
		_w1882_,
		_w1899_
	);
	LUT2 #(
		.INIT('h1)
	) name1764 (
		_w1890_,
		_w1898_,
		_w1900_
	);
	LUT2 #(
		.INIT('h8)
	) name1765 (
		_w1899_,
		_w1900_,
		_w1901_
	);
	LUT2 #(
		.INIT('h2)
	) name1766 (
		\shift[6] ,
		_w1901_,
		_w1902_
	);
	LUT2 #(
		.INIT('h1)
	) name1767 (
		_w1866_,
		_w1902_,
		_w1903_
	);
	LUT2 #(
		.INIT('h2)
	) name1768 (
		_w136_,
		_w1165_,
		_w1904_
	);
	LUT2 #(
		.INIT('h2)
	) name1769 (
		_w147_,
		_w1157_,
		_w1905_
	);
	LUT2 #(
		.INIT('h2)
	) name1770 (
		_w158_,
		_w1221_,
		_w1906_
	);
	LUT2 #(
		.INIT('h2)
	) name1771 (
		_w169_,
		_w1213_,
		_w1907_
	);
	LUT2 #(
		.INIT('h1)
	) name1772 (
		_w1904_,
		_w1905_,
		_w1908_
	);
	LUT2 #(
		.INIT('h1)
	) name1773 (
		_w1906_,
		_w1907_,
		_w1909_
	);
	LUT2 #(
		.INIT('h8)
	) name1774 (
		_w1908_,
		_w1909_,
		_w1910_
	);
	LUT2 #(
		.INIT('h2)
	) name1775 (
		_w183_,
		_w1910_,
		_w1911_
	);
	LUT2 #(
		.INIT('h2)
	) name1776 (
		_w136_,
		_w1129_,
		_w1912_
	);
	LUT2 #(
		.INIT('h2)
	) name1777 (
		_w147_,
		_w1121_,
		_w1913_
	);
	LUT2 #(
		.INIT('h2)
	) name1778 (
		_w158_,
		_w1149_,
		_w1914_
	);
	LUT2 #(
		.INIT('h2)
	) name1779 (
		_w169_,
		_w1141_,
		_w1915_
	);
	LUT2 #(
		.INIT('h1)
	) name1780 (
		_w1912_,
		_w1913_,
		_w1916_
	);
	LUT2 #(
		.INIT('h1)
	) name1781 (
		_w1914_,
		_w1915_,
		_w1917_
	);
	LUT2 #(
		.INIT('h8)
	) name1782 (
		_w1916_,
		_w1917_,
		_w1918_
	);
	LUT2 #(
		.INIT('h2)
	) name1783 (
		_w228_,
		_w1918_,
		_w1919_
	);
	LUT2 #(
		.INIT('h2)
	) name1784 (
		_w136_,
		_w1346_,
		_w1920_
	);
	LUT2 #(
		.INIT('h2)
	) name1785 (
		_w147_,
		_w1338_,
		_w1921_
	);
	LUT2 #(
		.INIT('h2)
	) name1786 (
		_w158_,
		_w1185_,
		_w1922_
	);
	LUT2 #(
		.INIT('h2)
	) name1787 (
		_w169_,
		_w1177_,
		_w1923_
	);
	LUT2 #(
		.INIT('h1)
	) name1788 (
		_w1920_,
		_w1921_,
		_w1924_
	);
	LUT2 #(
		.INIT('h1)
	) name1789 (
		_w1922_,
		_w1923_,
		_w1925_
	);
	LUT2 #(
		.INIT('h8)
	) name1790 (
		_w1924_,
		_w1925_,
		_w1926_
	);
	LUT2 #(
		.INIT('h2)
	) name1791 (
		_w273_,
		_w1926_,
		_w1927_
	);
	LUT2 #(
		.INIT('h2)
	) name1792 (
		_w136_,
		_w1201_,
		_w1928_
	);
	LUT2 #(
		.INIT('h2)
	) name1793 (
		_w147_,
		_w1193_,
		_w1929_
	);
	LUT2 #(
		.INIT('h2)
	) name1794 (
		_w158_,
		_w1113_,
		_w1930_
	);
	LUT2 #(
		.INIT('h2)
	) name1795 (
		_w169_,
		_w1105_,
		_w1931_
	);
	LUT2 #(
		.INIT('h1)
	) name1796 (
		_w1928_,
		_w1929_,
		_w1932_
	);
	LUT2 #(
		.INIT('h1)
	) name1797 (
		_w1930_,
		_w1931_,
		_w1933_
	);
	LUT2 #(
		.INIT('h8)
	) name1798 (
		_w1932_,
		_w1933_,
		_w1934_
	);
	LUT2 #(
		.INIT('h2)
	) name1799 (
		_w318_,
		_w1934_,
		_w1935_
	);
	LUT2 #(
		.INIT('h1)
	) name1800 (
		_w1911_,
		_w1919_,
		_w1936_
	);
	LUT2 #(
		.INIT('h1)
	) name1801 (
		_w1927_,
		_w1935_,
		_w1937_
	);
	LUT2 #(
		.INIT('h8)
	) name1802 (
		_w1936_,
		_w1937_,
		_w1938_
	);
	LUT2 #(
		.INIT('h1)
	) name1803 (
		\shift[6] ,
		_w1938_,
		_w1939_
	);
	LUT2 #(
		.INIT('h2)
	) name1804 (
		_w136_,
		_w1277_,
		_w1940_
	);
	LUT2 #(
		.INIT('h2)
	) name1805 (
		_w169_,
		_w1289_,
		_w1941_
	);
	LUT2 #(
		.INIT('h2)
	) name1806 (
		_w158_,
		_w1294_,
		_w1942_
	);
	LUT2 #(
		.INIT('h2)
	) name1807 (
		_w147_,
		_w1269_,
		_w1943_
	);
	LUT2 #(
		.INIT('h1)
	) name1808 (
		_w1940_,
		_w1941_,
		_w1944_
	);
	LUT2 #(
		.INIT('h1)
	) name1809 (
		_w1942_,
		_w1943_,
		_w1945_
	);
	LUT2 #(
		.INIT('h8)
	) name1810 (
		_w1944_,
		_w1945_,
		_w1946_
	);
	LUT2 #(
		.INIT('h2)
	) name1811 (
		_w318_,
		_w1946_,
		_w1947_
	);
	LUT2 #(
		.INIT('h2)
	) name1812 (
		_w136_,
		_w1237_,
		_w1948_
	);
	LUT2 #(
		.INIT('h2)
	) name1813 (
		_w147_,
		_w1229_,
		_w1949_
	);
	LUT2 #(
		.INIT('h2)
	) name1814 (
		_w158_,
		_w1261_,
		_w1950_
	);
	LUT2 #(
		.INIT('h2)
	) name1815 (
		_w169_,
		_w1253_,
		_w1951_
	);
	LUT2 #(
		.INIT('h1)
	) name1816 (
		_w1948_,
		_w1949_,
		_w1952_
	);
	LUT2 #(
		.INIT('h1)
	) name1817 (
		_w1950_,
		_w1951_,
		_w1953_
	);
	LUT2 #(
		.INIT('h8)
	) name1818 (
		_w1952_,
		_w1953_,
		_w1954_
	);
	LUT2 #(
		.INIT('h2)
	) name1819 (
		_w273_,
		_w1954_,
		_w1955_
	);
	LUT2 #(
		.INIT('h2)
	) name1820 (
		_w136_,
		_w1310_,
		_w1956_
	);
	LUT2 #(
		.INIT('h2)
	) name1821 (
		_w147_,
		_w1302_,
		_w1957_
	);
	LUT2 #(
		.INIT('h2)
	) name1822 (
		_w158_,
		_w1366_,
		_w1958_
	);
	LUT2 #(
		.INIT('h2)
	) name1823 (
		_w169_,
		_w1358_,
		_w1959_
	);
	LUT2 #(
		.INIT('h1)
	) name1824 (
		_w1956_,
		_w1957_,
		_w1960_
	);
	LUT2 #(
		.INIT('h1)
	) name1825 (
		_w1958_,
		_w1959_,
		_w1961_
	);
	LUT2 #(
		.INIT('h8)
	) name1826 (
		_w1960_,
		_w1961_,
		_w1962_
	);
	LUT2 #(
		.INIT('h2)
	) name1827 (
		_w228_,
		_w1962_,
		_w1963_
	);
	LUT2 #(
		.INIT('h2)
	) name1828 (
		_w136_,
		_w1382_,
		_w1964_
	);
	LUT2 #(
		.INIT('h2)
	) name1829 (
		_w147_,
		_w1374_,
		_w1965_
	);
	LUT2 #(
		.INIT('h2)
	) name1830 (
		_w158_,
		_w1330_,
		_w1966_
	);
	LUT2 #(
		.INIT('h2)
	) name1831 (
		_w169_,
		_w1322_,
		_w1967_
	);
	LUT2 #(
		.INIT('h1)
	) name1832 (
		_w1964_,
		_w1965_,
		_w1968_
	);
	LUT2 #(
		.INIT('h1)
	) name1833 (
		_w1966_,
		_w1967_,
		_w1969_
	);
	LUT2 #(
		.INIT('h8)
	) name1834 (
		_w1968_,
		_w1969_,
		_w1970_
	);
	LUT2 #(
		.INIT('h2)
	) name1835 (
		_w183_,
		_w1970_,
		_w1971_
	);
	LUT2 #(
		.INIT('h1)
	) name1836 (
		_w1947_,
		_w1955_,
		_w1972_
	);
	LUT2 #(
		.INIT('h1)
	) name1837 (
		_w1963_,
		_w1971_,
		_w1973_
	);
	LUT2 #(
		.INIT('h8)
	) name1838 (
		_w1972_,
		_w1973_,
		_w1974_
	);
	LUT2 #(
		.INIT('h2)
	) name1839 (
		\shift[6] ,
		_w1974_,
		_w1975_
	);
	LUT2 #(
		.INIT('h1)
	) name1840 (
		_w1939_,
		_w1975_,
		_w1976_
	);
	LUT2 #(
		.INIT('h2)
	) name1841 (
		_w136_,
		_w203_,
		_w1977_
	);
	LUT2 #(
		.INIT('h2)
	) name1842 (
		_w147_,
		_w223_,
		_w1978_
	);
	LUT2 #(
		.INIT('h4)
	) name1843 (
		_w145_,
		_w158_,
		_w1979_
	);
	LUT2 #(
		.INIT('h2)
	) name1844 (
		_w169_,
		_w213_,
		_w1980_
	);
	LUT2 #(
		.INIT('h1)
	) name1845 (
		_w1977_,
		_w1978_,
		_w1981_
	);
	LUT2 #(
		.INIT('h1)
	) name1846 (
		_w1979_,
		_w1980_,
		_w1982_
	);
	LUT2 #(
		.INIT('h8)
	) name1847 (
		_w1981_,
		_w1982_,
		_w1983_
	);
	LUT2 #(
		.INIT('h2)
	) name1848 (
		_w183_,
		_w1983_,
		_w1984_
	);
	LUT2 #(
		.INIT('h2)
	) name1849 (
		_w136_,
		_w293_,
		_w1985_
	);
	LUT2 #(
		.INIT('h2)
	) name1850 (
		_w147_,
		_w313_,
		_w1986_
	);
	LUT2 #(
		.INIT('h2)
	) name1851 (
		_w158_,
		_w193_,
		_w1987_
	);
	LUT2 #(
		.INIT('h2)
	) name1852 (
		_w169_,
		_w303_,
		_w1988_
	);
	LUT2 #(
		.INIT('h1)
	) name1853 (
		_w1985_,
		_w1986_,
		_w1989_
	);
	LUT2 #(
		.INIT('h1)
	) name1854 (
		_w1987_,
		_w1988_,
		_w1990_
	);
	LUT2 #(
		.INIT('h8)
	) name1855 (
		_w1989_,
		_w1990_,
		_w1991_
	);
	LUT2 #(
		.INIT('h2)
	) name1856 (
		_w228_,
		_w1991_,
		_w1992_
	);
	LUT2 #(
		.INIT('h2)
	) name1857 (
		_w136_,
		_w342_,
		_w1993_
	);
	LUT2 #(
		.INIT('h2)
	) name1858 (
		_w147_,
		_w362_,
		_w1994_
	);
	LUT2 #(
		.INIT('h2)
	) name1859 (
		_w158_,
		_w238_,
		_w1995_
	);
	LUT2 #(
		.INIT('h2)
	) name1860 (
		_w169_,
		_w352_,
		_w1996_
	);
	LUT2 #(
		.INIT('h1)
	) name1861 (
		_w1993_,
		_w1994_,
		_w1997_
	);
	LUT2 #(
		.INIT('h1)
	) name1862 (
		_w1995_,
		_w1996_,
		_w1998_
	);
	LUT2 #(
		.INIT('h8)
	) name1863 (
		_w1997_,
		_w1998_,
		_w1999_
	);
	LUT2 #(
		.INIT('h2)
	) name1864 (
		_w273_,
		_w1999_,
		_w2000_
	);
	LUT2 #(
		.INIT('h2)
	) name1865 (
		_w136_,
		_w248_,
		_w2001_
	);
	LUT2 #(
		.INIT('h2)
	) name1866 (
		_w147_,
		_w268_,
		_w2002_
	);
	LUT2 #(
		.INIT('h2)
	) name1867 (
		_w158_,
		_w283_,
		_w2003_
	);
	LUT2 #(
		.INIT('h2)
	) name1868 (
		_w169_,
		_w258_,
		_w2004_
	);
	LUT2 #(
		.INIT('h1)
	) name1869 (
		_w2001_,
		_w2002_,
		_w2005_
	);
	LUT2 #(
		.INIT('h1)
	) name1870 (
		_w2003_,
		_w2004_,
		_w2006_
	);
	LUT2 #(
		.INIT('h8)
	) name1871 (
		_w2005_,
		_w2006_,
		_w2007_
	);
	LUT2 #(
		.INIT('h2)
	) name1872 (
		_w318_,
		_w2007_,
		_w2008_
	);
	LUT2 #(
		.INIT('h1)
	) name1873 (
		_w1984_,
		_w1992_,
		_w2009_
	);
	LUT2 #(
		.INIT('h1)
	) name1874 (
		_w2000_,
		_w2008_,
		_w2010_
	);
	LUT2 #(
		.INIT('h8)
	) name1875 (
		_w2009_,
		_w2010_,
		_w2011_
	);
	LUT2 #(
		.INIT('h1)
	) name1876 (
		\shift[6] ,
		_w2011_,
		_w2012_
	);
	LUT2 #(
		.INIT('h2)
	) name1877 (
		_w136_,
		_w430_,
		_w2013_
	);
	LUT2 #(
		.INIT('h2)
	) name1878 (
		_w147_,
		_w450_,
		_w2014_
	);
	LUT2 #(
		.INIT('h2)
	) name1879 (
		_w158_,
		_w464_,
		_w2015_
	);
	LUT2 #(
		.INIT('h2)
	) name1880 (
		_w169_,
		_w440_,
		_w2016_
	);
	LUT2 #(
		.INIT('h1)
	) name1881 (
		_w2013_,
		_w2014_,
		_w2017_
	);
	LUT2 #(
		.INIT('h1)
	) name1882 (
		_w2015_,
		_w2016_,
		_w2018_
	);
	LUT2 #(
		.INIT('h8)
	) name1883 (
		_w2017_,
		_w2018_,
		_w2019_
	);
	LUT2 #(
		.INIT('h2)
	) name1884 (
		_w318_,
		_w2019_,
		_w2020_
	);
	LUT2 #(
		.INIT('h2)
	) name1885 (
		_w136_,
		_w156_,
		_w2021_
	);
	LUT2 #(
		.INIT('h2)
	) name1886 (
		_w147_,
		_w178_,
		_w2022_
	);
	LUT2 #(
		.INIT('h2)
	) name1887 (
		_w158_,
		_w420_,
		_w2023_
	);
	LUT2 #(
		.INIT('h4)
	) name1888 (
		_w167_,
		_w169_,
		_w2024_
	);
	LUT2 #(
		.INIT('h1)
	) name1889 (
		_w2021_,
		_w2022_,
		_w2025_
	);
	LUT2 #(
		.INIT('h1)
	) name1890 (
		_w2023_,
		_w2024_,
		_w2026_
	);
	LUT2 #(
		.INIT('h8)
	) name1891 (
		_w2025_,
		_w2026_,
		_w2027_
	);
	LUT2 #(
		.INIT('h2)
	) name1892 (
		_w273_,
		_w2027_,
		_w2028_
	);
	LUT2 #(
		.INIT('h2)
	) name1893 (
		_w136_,
		_w474_,
		_w2029_
	);
	LUT2 #(
		.INIT('h2)
	) name1894 (
		_w147_,
		_w496_,
		_w2030_
	);
	LUT2 #(
		.INIT('h2)
	) name1895 (
		_w158_,
		_w376_,
		_w2031_
	);
	LUT2 #(
		.INIT('h2)
	) name1896 (
		_w169_,
		_w484_,
		_w2032_
	);
	LUT2 #(
		.INIT('h1)
	) name1897 (
		_w2029_,
		_w2030_,
		_w2033_
	);
	LUT2 #(
		.INIT('h1)
	) name1898 (
		_w2031_,
		_w2032_,
		_w2034_
	);
	LUT2 #(
		.INIT('h8)
	) name1899 (
		_w2033_,
		_w2034_,
		_w2035_
	);
	LUT2 #(
		.INIT('h2)
	) name1900 (
		_w228_,
		_w2035_,
		_w2036_
	);
	LUT2 #(
		.INIT('h2)
	) name1901 (
		_w136_,
		_w386_,
		_w2037_
	);
	LUT2 #(
		.INIT('h2)
	) name1902 (
		_w147_,
		_w406_,
		_w2038_
	);
	LUT2 #(
		.INIT('h2)
	) name1903 (
		_w158_,
		_w332_,
		_w2039_
	);
	LUT2 #(
		.INIT('h2)
	) name1904 (
		_w169_,
		_w396_,
		_w2040_
	);
	LUT2 #(
		.INIT('h1)
	) name1905 (
		_w2037_,
		_w2038_,
		_w2041_
	);
	LUT2 #(
		.INIT('h1)
	) name1906 (
		_w2039_,
		_w2040_,
		_w2042_
	);
	LUT2 #(
		.INIT('h8)
	) name1907 (
		_w2041_,
		_w2042_,
		_w2043_
	);
	LUT2 #(
		.INIT('h2)
	) name1908 (
		_w183_,
		_w2043_,
		_w2044_
	);
	LUT2 #(
		.INIT('h1)
	) name1909 (
		_w2020_,
		_w2028_,
		_w2045_
	);
	LUT2 #(
		.INIT('h1)
	) name1910 (
		_w2036_,
		_w2044_,
		_w2046_
	);
	LUT2 #(
		.INIT('h8)
	) name1911 (
		_w2045_,
		_w2046_,
		_w2047_
	);
	LUT2 #(
		.INIT('h2)
	) name1912 (
		\shift[6] ,
		_w2047_,
		_w2048_
	);
	LUT2 #(
		.INIT('h1)
	) name1913 (
		_w2012_,
		_w2048_,
		_w2049_
	);
	LUT2 #(
		.INIT('h2)
	) name1914 (
		_w136_,
		_w581_,
		_w2050_
	);
	LUT2 #(
		.INIT('h2)
	) name1915 (
		_w147_,
		_w605_,
		_w2051_
	);
	LUT2 #(
		.INIT('h2)
	) name1916 (
		_w158_,
		_w517_,
		_w2052_
	);
	LUT2 #(
		.INIT('h2)
	) name1917 (
		_w169_,
		_w593_,
		_w2053_
	);
	LUT2 #(
		.INIT('h1)
	) name1918 (
		_w2050_,
		_w2051_,
		_w2054_
	);
	LUT2 #(
		.INIT('h1)
	) name1919 (
		_w2052_,
		_w2053_,
		_w2055_
	);
	LUT2 #(
		.INIT('h8)
	) name1920 (
		_w2054_,
		_w2055_,
		_w2056_
	);
	LUT2 #(
		.INIT('h2)
	) name1921 (
		_w183_,
		_w2056_,
		_w2057_
	);
	LUT2 #(
		.INIT('h2)
	) name1922 (
		_w136_,
		_w685_,
		_w2058_
	);
	LUT2 #(
		.INIT('h2)
	) name1923 (
		_w147_,
		_w709_,
		_w2059_
	);
	LUT2 #(
		.INIT('h2)
	) name1924 (
		_w158_,
		_w569_,
		_w2060_
	);
	LUT2 #(
		.INIT('h2)
	) name1925 (
		_w169_,
		_w697_,
		_w2061_
	);
	LUT2 #(
		.INIT('h1)
	) name1926 (
		_w2058_,
		_w2059_,
		_w2062_
	);
	LUT2 #(
		.INIT('h1)
	) name1927 (
		_w2060_,
		_w2061_,
		_w2063_
	);
	LUT2 #(
		.INIT('h8)
	) name1928 (
		_w2062_,
		_w2063_,
		_w2064_
	);
	LUT2 #(
		.INIT('h2)
	) name1929 (
		_w228_,
		_w2064_,
		_w2065_
	);
	LUT2 #(
		.INIT('h2)
	) name1930 (
		_w136_,
		_w793_,
		_w2066_
	);
	LUT2 #(
		.INIT('h2)
	) name1931 (
		_w147_,
		_w817_,
		_w2067_
	);
	LUT2 #(
		.INIT('h2)
	) name1932 (
		_w158_,
		_w621_,
		_w2068_
	);
	LUT2 #(
		.INIT('h2)
	) name1933 (
		_w169_,
		_w805_,
		_w2069_
	);
	LUT2 #(
		.INIT('h1)
	) name1934 (
		_w2066_,
		_w2067_,
		_w2070_
	);
	LUT2 #(
		.INIT('h1)
	) name1935 (
		_w2068_,
		_w2069_,
		_w2071_
	);
	LUT2 #(
		.INIT('h8)
	) name1936 (
		_w2070_,
		_w2071_,
		_w2072_
	);
	LUT2 #(
		.INIT('h2)
	) name1937 (
		_w273_,
		_w2072_,
		_w2073_
	);
	LUT2 #(
		.INIT('h2)
	) name1938 (
		_w136_,
		_w633_,
		_w2074_
	);
	LUT2 #(
		.INIT('h2)
	) name1939 (
		_w147_,
		_w657_,
		_w2075_
	);
	LUT2 #(
		.INIT('h2)
	) name1940 (
		_w158_,
		_w673_,
		_w2076_
	);
	LUT2 #(
		.INIT('h2)
	) name1941 (
		_w169_,
		_w645_,
		_w2077_
	);
	LUT2 #(
		.INIT('h1)
	) name1942 (
		_w2074_,
		_w2075_,
		_w2078_
	);
	LUT2 #(
		.INIT('h1)
	) name1943 (
		_w2076_,
		_w2077_,
		_w2079_
	);
	LUT2 #(
		.INIT('h8)
	) name1944 (
		_w2078_,
		_w2079_,
		_w2080_
	);
	LUT2 #(
		.INIT('h2)
	) name1945 (
		_w318_,
		_w2080_,
		_w2081_
	);
	LUT2 #(
		.INIT('h1)
	) name1946 (
		_w2057_,
		_w2065_,
		_w2082_
	);
	LUT2 #(
		.INIT('h1)
	) name1947 (
		_w2073_,
		_w2081_,
		_w2083_
	);
	LUT2 #(
		.INIT('h8)
	) name1948 (
		_w2082_,
		_w2083_,
		_w2084_
	);
	LUT2 #(
		.INIT('h1)
	) name1949 (
		\shift[6] ,
		_w2084_,
		_w2085_
	);
	LUT2 #(
		.INIT('h2)
	) name1950 (
		_w136_,
		_w741_,
		_w2086_
	);
	LUT2 #(
		.INIT('h2)
	) name1951 (
		_w147_,
		_w765_,
		_w2087_
	);
	LUT2 #(
		.INIT('h2)
	) name1952 (
		_w158_,
		_w833_,
		_w2088_
	);
	LUT2 #(
		.INIT('h2)
	) name1953 (
		_w169_,
		_w753_,
		_w2089_
	);
	LUT2 #(
		.INIT('h1)
	) name1954 (
		_w2086_,
		_w2087_,
		_w2090_
	);
	LUT2 #(
		.INIT('h1)
	) name1955 (
		_w2088_,
		_w2089_,
		_w2091_
	);
	LUT2 #(
		.INIT('h8)
	) name1956 (
		_w2090_,
		_w2091_,
		_w2092_
	);
	LUT2 #(
		.INIT('h2)
	) name1957 (
		_w318_,
		_w2092_,
		_w2093_
	);
	LUT2 #(
		.INIT('h2)
	) name1958 (
		_w136_,
		_w529_,
		_w2094_
	);
	LUT2 #(
		.INIT('h2)
	) name1959 (
		_w147_,
		_w553_,
		_w2095_
	);
	LUT2 #(
		.INIT('h2)
	) name1960 (
		_w158_,
		_w729_,
		_w2096_
	);
	LUT2 #(
		.INIT('h2)
	) name1961 (
		_w169_,
		_w541_,
		_w2097_
	);
	LUT2 #(
		.INIT('h1)
	) name1962 (
		_w2094_,
		_w2095_,
		_w2098_
	);
	LUT2 #(
		.INIT('h1)
	) name1963 (
		_w2096_,
		_w2097_,
		_w2099_
	);
	LUT2 #(
		.INIT('h8)
	) name1964 (
		_w2098_,
		_w2099_,
		_w2100_
	);
	LUT2 #(
		.INIT('h2)
	) name1965 (
		_w273_,
		_w2100_,
		_w2101_
	);
	LUT2 #(
		.INIT('h2)
	) name1966 (
		_w136_,
		_w843_,
		_w2102_
	);
	LUT2 #(
		.INIT('h2)
	) name1967 (
		_w147_,
		_w865_,
		_w2103_
	);
	LUT2 #(
		.INIT('h2)
	) name1968 (
		_w158_,
		_w881_,
		_w2104_
	);
	LUT2 #(
		.INIT('h2)
	) name1969 (
		_w169_,
		_w855_,
		_w2105_
	);
	LUT2 #(
		.INIT('h1)
	) name1970 (
		_w2102_,
		_w2103_,
		_w2106_
	);
	LUT2 #(
		.INIT('h1)
	) name1971 (
		_w2104_,
		_w2105_,
		_w2107_
	);
	LUT2 #(
		.INIT('h8)
	) name1972 (
		_w2106_,
		_w2107_,
		_w2108_
	);
	LUT2 #(
		.INIT('h2)
	) name1973 (
		_w228_,
		_w2108_,
		_w2109_
	);
	LUT2 #(
		.INIT('h2)
	) name1974 (
		_w136_,
		_w893_,
		_w2110_
	);
	LUT2 #(
		.INIT('h2)
	) name1975 (
		_w147_,
		_w917_,
		_w2111_
	);
	LUT2 #(
		.INIT('h2)
	) name1976 (
		_w158_,
		_w781_,
		_w2112_
	);
	LUT2 #(
		.INIT('h2)
	) name1977 (
		_w169_,
		_w905_,
		_w2113_
	);
	LUT2 #(
		.INIT('h1)
	) name1978 (
		_w2110_,
		_w2111_,
		_w2114_
	);
	LUT2 #(
		.INIT('h1)
	) name1979 (
		_w2112_,
		_w2113_,
		_w2115_
	);
	LUT2 #(
		.INIT('h8)
	) name1980 (
		_w2114_,
		_w2115_,
		_w2116_
	);
	LUT2 #(
		.INIT('h2)
	) name1981 (
		_w183_,
		_w2116_,
		_w2117_
	);
	LUT2 #(
		.INIT('h1)
	) name1982 (
		_w2093_,
		_w2101_,
		_w2118_
	);
	LUT2 #(
		.INIT('h1)
	) name1983 (
		_w2109_,
		_w2117_,
		_w2119_
	);
	LUT2 #(
		.INIT('h8)
	) name1984 (
		_w2118_,
		_w2119_,
		_w2120_
	);
	LUT2 #(
		.INIT('h2)
	) name1985 (
		\shift[6] ,
		_w2120_,
		_w2121_
	);
	LUT2 #(
		.INIT('h1)
	) name1986 (
		_w2085_,
		_w2121_,
		_w2122_
	);
	LUT2 #(
		.INIT('h2)
	) name1987 (
		_w136_,
		_w954_,
		_w2123_
	);
	LUT2 #(
		.INIT('h2)
	) name1988 (
		_w147_,
		_w962_,
		_w2124_
	);
	LUT2 #(
		.INIT('h2)
	) name1989 (
		_w158_,
		_w930_,
		_w2125_
	);
	LUT2 #(
		.INIT('h2)
	) name1990 (
		_w169_,
		_w958_,
		_w2126_
	);
	LUT2 #(
		.INIT('h1)
	) name1991 (
		_w2123_,
		_w2124_,
		_w2127_
	);
	LUT2 #(
		.INIT('h1)
	) name1992 (
		_w2125_,
		_w2126_,
		_w2128_
	);
	LUT2 #(
		.INIT('h8)
	) name1993 (
		_w2127_,
		_w2128_,
		_w2129_
	);
	LUT2 #(
		.INIT('h2)
	) name1994 (
		_w183_,
		_w2129_,
		_w2130_
	);
	LUT2 #(
		.INIT('h2)
	) name1995 (
		_w136_,
		_w994_,
		_w2131_
	);
	LUT2 #(
		.INIT('h2)
	) name1996 (
		_w147_,
		_w1002_,
		_w2132_
	);
	LUT2 #(
		.INIT('h2)
	) name1997 (
		_w158_,
		_w950_,
		_w2133_
	);
	LUT2 #(
		.INIT('h2)
	) name1998 (
		_w169_,
		_w998_,
		_w2134_
	);
	LUT2 #(
		.INIT('h1)
	) name1999 (
		_w2131_,
		_w2132_,
		_w2135_
	);
	LUT2 #(
		.INIT('h1)
	) name2000 (
		_w2133_,
		_w2134_,
		_w2136_
	);
	LUT2 #(
		.INIT('h8)
	) name2001 (
		_w2135_,
		_w2136_,
		_w2137_
	);
	LUT2 #(
		.INIT('h2)
	) name2002 (
		_w228_,
		_w2137_,
		_w2138_
	);
	LUT2 #(
		.INIT('h2)
	) name2003 (
		_w136_,
		_w1038_,
		_w2139_
	);
	LUT2 #(
		.INIT('h2)
	) name2004 (
		_w147_,
		_w1046_,
		_w2140_
	);
	LUT2 #(
		.INIT('h2)
	) name2005 (
		_w158_,
		_w970_,
		_w2141_
	);
	LUT2 #(
		.INIT('h2)
	) name2006 (
		_w169_,
		_w1042_,
		_w2142_
	);
	LUT2 #(
		.INIT('h1)
	) name2007 (
		_w2139_,
		_w2140_,
		_w2143_
	);
	LUT2 #(
		.INIT('h1)
	) name2008 (
		_w2141_,
		_w2142_,
		_w2144_
	);
	LUT2 #(
		.INIT('h8)
	) name2009 (
		_w2143_,
		_w2144_,
		_w2145_
	);
	LUT2 #(
		.INIT('h2)
	) name2010 (
		_w273_,
		_w2145_,
		_w2146_
	);
	LUT2 #(
		.INIT('h2)
	) name2011 (
		_w136_,
		_w974_,
		_w2147_
	);
	LUT2 #(
		.INIT('h2)
	) name2012 (
		_w147_,
		_w982_,
		_w2148_
	);
	LUT2 #(
		.INIT('h2)
	) name2013 (
		_w158_,
		_w990_,
		_w2149_
	);
	LUT2 #(
		.INIT('h2)
	) name2014 (
		_w169_,
		_w978_,
		_w2150_
	);
	LUT2 #(
		.INIT('h1)
	) name2015 (
		_w2147_,
		_w2148_,
		_w2151_
	);
	LUT2 #(
		.INIT('h1)
	) name2016 (
		_w2149_,
		_w2150_,
		_w2152_
	);
	LUT2 #(
		.INIT('h8)
	) name2017 (
		_w2151_,
		_w2152_,
		_w2153_
	);
	LUT2 #(
		.INIT('h2)
	) name2018 (
		_w318_,
		_w2153_,
		_w2154_
	);
	LUT2 #(
		.INIT('h1)
	) name2019 (
		_w2130_,
		_w2138_,
		_w2155_
	);
	LUT2 #(
		.INIT('h1)
	) name2020 (
		_w2146_,
		_w2154_,
		_w2156_
	);
	LUT2 #(
		.INIT('h8)
	) name2021 (
		_w2155_,
		_w2156_,
		_w2157_
	);
	LUT2 #(
		.INIT('h1)
	) name2022 (
		\shift[6] ,
		_w2157_,
		_w2158_
	);
	LUT2 #(
		.INIT('h2)
	) name2023 (
		_w136_,
		_w1018_,
		_w2159_
	);
	LUT2 #(
		.INIT('h2)
	) name2024 (
		_w147_,
		_w1026_,
		_w2160_
	);
	LUT2 #(
		.INIT('h2)
	) name2025 (
		_w158_,
		_w1054_,
		_w2161_
	);
	LUT2 #(
		.INIT('h2)
	) name2026 (
		_w169_,
		_w1022_,
		_w2162_
	);
	LUT2 #(
		.INIT('h1)
	) name2027 (
		_w2159_,
		_w2160_,
		_w2163_
	);
	LUT2 #(
		.INIT('h1)
	) name2028 (
		_w2161_,
		_w2162_,
		_w2164_
	);
	LUT2 #(
		.INIT('h8)
	) name2029 (
		_w2163_,
		_w2164_,
		_w2165_
	);
	LUT2 #(
		.INIT('h2)
	) name2030 (
		_w318_,
		_w2165_,
		_w2166_
	);
	LUT2 #(
		.INIT('h2)
	) name2031 (
		_w136_,
		_w934_,
		_w2167_
	);
	LUT2 #(
		.INIT('h2)
	) name2032 (
		_w147_,
		_w942_,
		_w2168_
	);
	LUT2 #(
		.INIT('h2)
	) name2033 (
		_w158_,
		_w1014_,
		_w2169_
	);
	LUT2 #(
		.INIT('h2)
	) name2034 (
		_w169_,
		_w938_,
		_w2170_
	);
	LUT2 #(
		.INIT('h1)
	) name2035 (
		_w2167_,
		_w2168_,
		_w2171_
	);
	LUT2 #(
		.INIT('h1)
	) name2036 (
		_w2169_,
		_w2170_,
		_w2172_
	);
	LUT2 #(
		.INIT('h8)
	) name2037 (
		_w2171_,
		_w2172_,
		_w2173_
	);
	LUT2 #(
		.INIT('h2)
	) name2038 (
		_w273_,
		_w2173_,
		_w2174_
	);
	LUT2 #(
		.INIT('h2)
	) name2039 (
		_w136_,
		_w1058_,
		_w2175_
	);
	LUT2 #(
		.INIT('h2)
	) name2040 (
		_w147_,
		_w1068_,
		_w2176_
	);
	LUT2 #(
		.INIT('h2)
	) name2041 (
		_w158_,
		_w1076_,
		_w2177_
	);
	LUT2 #(
		.INIT('h2)
	) name2042 (
		_w169_,
		_w1063_,
		_w2178_
	);
	LUT2 #(
		.INIT('h1)
	) name2043 (
		_w2175_,
		_w2176_,
		_w2179_
	);
	LUT2 #(
		.INIT('h1)
	) name2044 (
		_w2177_,
		_w2178_,
		_w2180_
	);
	LUT2 #(
		.INIT('h8)
	) name2045 (
		_w2179_,
		_w2180_,
		_w2181_
	);
	LUT2 #(
		.INIT('h2)
	) name2046 (
		_w228_,
		_w2181_,
		_w2182_
	);
	LUT2 #(
		.INIT('h2)
	) name2047 (
		_w136_,
		_w1080_,
		_w2183_
	);
	LUT2 #(
		.INIT('h2)
	) name2048 (
		_w147_,
		_w1088_,
		_w2184_
	);
	LUT2 #(
		.INIT('h2)
	) name2049 (
		_w158_,
		_w1034_,
		_w2185_
	);
	LUT2 #(
		.INIT('h2)
	) name2050 (
		_w169_,
		_w1084_,
		_w2186_
	);
	LUT2 #(
		.INIT('h1)
	) name2051 (
		_w2183_,
		_w2184_,
		_w2187_
	);
	LUT2 #(
		.INIT('h1)
	) name2052 (
		_w2185_,
		_w2186_,
		_w2188_
	);
	LUT2 #(
		.INIT('h8)
	) name2053 (
		_w2187_,
		_w2188_,
		_w2189_
	);
	LUT2 #(
		.INIT('h2)
	) name2054 (
		_w183_,
		_w2189_,
		_w2190_
	);
	LUT2 #(
		.INIT('h1)
	) name2055 (
		_w2166_,
		_w2174_,
		_w2191_
	);
	LUT2 #(
		.INIT('h1)
	) name2056 (
		_w2182_,
		_w2190_,
		_w2192_
	);
	LUT2 #(
		.INIT('h8)
	) name2057 (
		_w2191_,
		_w2192_,
		_w2193_
	);
	LUT2 #(
		.INIT('h2)
	) name2058 (
		\shift[6] ,
		_w2193_,
		_w2194_
	);
	LUT2 #(
		.INIT('h1)
	) name2059 (
		_w2158_,
		_w2194_,
		_w2195_
	);
	LUT2 #(
		.INIT('h2)
	) name2060 (
		_w136_,
		_w1149_,
		_w2196_
	);
	LUT2 #(
		.INIT('h2)
	) name2061 (
		_w147_,
		_w1165_,
		_w2197_
	);
	LUT2 #(
		.INIT('h2)
	) name2062 (
		_w158_,
		_w1213_,
		_w2198_
	);
	LUT2 #(
		.INIT('h2)
	) name2063 (
		_w169_,
		_w1157_,
		_w2199_
	);
	LUT2 #(
		.INIT('h1)
	) name2064 (
		_w2196_,
		_w2197_,
		_w2200_
	);
	LUT2 #(
		.INIT('h1)
	) name2065 (
		_w2198_,
		_w2199_,
		_w2201_
	);
	LUT2 #(
		.INIT('h8)
	) name2066 (
		_w2200_,
		_w2201_,
		_w2202_
	);
	LUT2 #(
		.INIT('h2)
	) name2067 (
		_w183_,
		_w2202_,
		_w2203_
	);
	LUT2 #(
		.INIT('h2)
	) name2068 (
		_w136_,
		_w1113_,
		_w2204_
	);
	LUT2 #(
		.INIT('h2)
	) name2069 (
		_w147_,
		_w1129_,
		_w2205_
	);
	LUT2 #(
		.INIT('h2)
	) name2070 (
		_w158_,
		_w1141_,
		_w2206_
	);
	LUT2 #(
		.INIT('h2)
	) name2071 (
		_w169_,
		_w1121_,
		_w2207_
	);
	LUT2 #(
		.INIT('h1)
	) name2072 (
		_w2204_,
		_w2205_,
		_w2208_
	);
	LUT2 #(
		.INIT('h1)
	) name2073 (
		_w2206_,
		_w2207_,
		_w2209_
	);
	LUT2 #(
		.INIT('h8)
	) name2074 (
		_w2208_,
		_w2209_,
		_w2210_
	);
	LUT2 #(
		.INIT('h2)
	) name2075 (
		_w228_,
		_w2210_,
		_w2211_
	);
	LUT2 #(
		.INIT('h2)
	) name2076 (
		_w136_,
		_w1330_,
		_w2212_
	);
	LUT2 #(
		.INIT('h2)
	) name2077 (
		_w147_,
		_w1346_,
		_w2213_
	);
	LUT2 #(
		.INIT('h2)
	) name2078 (
		_w158_,
		_w1177_,
		_w2214_
	);
	LUT2 #(
		.INIT('h2)
	) name2079 (
		_w169_,
		_w1338_,
		_w2215_
	);
	LUT2 #(
		.INIT('h1)
	) name2080 (
		_w2212_,
		_w2213_,
		_w2216_
	);
	LUT2 #(
		.INIT('h1)
	) name2081 (
		_w2214_,
		_w2215_,
		_w2217_
	);
	LUT2 #(
		.INIT('h8)
	) name2082 (
		_w2216_,
		_w2217_,
		_w2218_
	);
	LUT2 #(
		.INIT('h2)
	) name2083 (
		_w273_,
		_w2218_,
		_w2219_
	);
	LUT2 #(
		.INIT('h2)
	) name2084 (
		_w136_,
		_w1185_,
		_w2220_
	);
	LUT2 #(
		.INIT('h2)
	) name2085 (
		_w147_,
		_w1201_,
		_w2221_
	);
	LUT2 #(
		.INIT('h2)
	) name2086 (
		_w158_,
		_w1105_,
		_w2222_
	);
	LUT2 #(
		.INIT('h2)
	) name2087 (
		_w169_,
		_w1193_,
		_w2223_
	);
	LUT2 #(
		.INIT('h1)
	) name2088 (
		_w2220_,
		_w2221_,
		_w2224_
	);
	LUT2 #(
		.INIT('h1)
	) name2089 (
		_w2222_,
		_w2223_,
		_w2225_
	);
	LUT2 #(
		.INIT('h8)
	) name2090 (
		_w2224_,
		_w2225_,
		_w2226_
	);
	LUT2 #(
		.INIT('h2)
	) name2091 (
		_w318_,
		_w2226_,
		_w2227_
	);
	LUT2 #(
		.INIT('h1)
	) name2092 (
		_w2203_,
		_w2211_,
		_w2228_
	);
	LUT2 #(
		.INIT('h1)
	) name2093 (
		_w2219_,
		_w2227_,
		_w2229_
	);
	LUT2 #(
		.INIT('h8)
	) name2094 (
		_w2228_,
		_w2229_,
		_w2230_
	);
	LUT2 #(
		.INIT('h1)
	) name2095 (
		\shift[6] ,
		_w2230_,
		_w2231_
	);
	LUT2 #(
		.INIT('h2)
	) name2096 (
		_w136_,
		_w1261_,
		_w2232_
	);
	LUT2 #(
		.INIT('h2)
	) name2097 (
		_w147_,
		_w1277_,
		_w2233_
	);
	LUT2 #(
		.INIT('h2)
	) name2098 (
		_w158_,
		_w1289_,
		_w2234_
	);
	LUT2 #(
		.INIT('h2)
	) name2099 (
		_w169_,
		_w1269_,
		_w2235_
	);
	LUT2 #(
		.INIT('h1)
	) name2100 (
		_w2232_,
		_w2233_,
		_w2236_
	);
	LUT2 #(
		.INIT('h1)
	) name2101 (
		_w2234_,
		_w2235_,
		_w2237_
	);
	LUT2 #(
		.INIT('h8)
	) name2102 (
		_w2236_,
		_w2237_,
		_w2238_
	);
	LUT2 #(
		.INIT('h2)
	) name2103 (
		_w318_,
		_w2238_,
		_w2239_
	);
	LUT2 #(
		.INIT('h2)
	) name2104 (
		_w136_,
		_w1221_,
		_w2240_
	);
	LUT2 #(
		.INIT('h2)
	) name2105 (
		_w147_,
		_w1237_,
		_w2241_
	);
	LUT2 #(
		.INIT('h2)
	) name2106 (
		_w158_,
		_w1253_,
		_w2242_
	);
	LUT2 #(
		.INIT('h2)
	) name2107 (
		_w169_,
		_w1229_,
		_w2243_
	);
	LUT2 #(
		.INIT('h1)
	) name2108 (
		_w2240_,
		_w2241_,
		_w2244_
	);
	LUT2 #(
		.INIT('h1)
	) name2109 (
		_w2242_,
		_w2243_,
		_w2245_
	);
	LUT2 #(
		.INIT('h8)
	) name2110 (
		_w2244_,
		_w2245_,
		_w2246_
	);
	LUT2 #(
		.INIT('h2)
	) name2111 (
		_w273_,
		_w2246_,
		_w2247_
	);
	LUT2 #(
		.INIT('h2)
	) name2112 (
		_w136_,
		_w1294_,
		_w2248_
	);
	LUT2 #(
		.INIT('h2)
	) name2113 (
		_w147_,
		_w1310_,
		_w2249_
	);
	LUT2 #(
		.INIT('h2)
	) name2114 (
		_w158_,
		_w1358_,
		_w2250_
	);
	LUT2 #(
		.INIT('h2)
	) name2115 (
		_w169_,
		_w1302_,
		_w2251_
	);
	LUT2 #(
		.INIT('h1)
	) name2116 (
		_w2248_,
		_w2249_,
		_w2252_
	);
	LUT2 #(
		.INIT('h1)
	) name2117 (
		_w2250_,
		_w2251_,
		_w2253_
	);
	LUT2 #(
		.INIT('h8)
	) name2118 (
		_w2252_,
		_w2253_,
		_w2254_
	);
	LUT2 #(
		.INIT('h2)
	) name2119 (
		_w228_,
		_w2254_,
		_w2255_
	);
	LUT2 #(
		.INIT('h2)
	) name2120 (
		_w136_,
		_w1366_,
		_w2256_
	);
	LUT2 #(
		.INIT('h2)
	) name2121 (
		_w147_,
		_w1382_,
		_w2257_
	);
	LUT2 #(
		.INIT('h2)
	) name2122 (
		_w158_,
		_w1322_,
		_w2258_
	);
	LUT2 #(
		.INIT('h2)
	) name2123 (
		_w169_,
		_w1374_,
		_w2259_
	);
	LUT2 #(
		.INIT('h1)
	) name2124 (
		_w2256_,
		_w2257_,
		_w2260_
	);
	LUT2 #(
		.INIT('h1)
	) name2125 (
		_w2258_,
		_w2259_,
		_w2261_
	);
	LUT2 #(
		.INIT('h8)
	) name2126 (
		_w2260_,
		_w2261_,
		_w2262_
	);
	LUT2 #(
		.INIT('h2)
	) name2127 (
		_w183_,
		_w2262_,
		_w2263_
	);
	LUT2 #(
		.INIT('h1)
	) name2128 (
		_w2239_,
		_w2247_,
		_w2264_
	);
	LUT2 #(
		.INIT('h1)
	) name2129 (
		_w2255_,
		_w2263_,
		_w2265_
	);
	LUT2 #(
		.INIT('h8)
	) name2130 (
		_w2264_,
		_w2265_,
		_w2266_
	);
	LUT2 #(
		.INIT('h2)
	) name2131 (
		\shift[6] ,
		_w2266_,
		_w2267_
	);
	LUT2 #(
		.INIT('h1)
	) name2132 (
		_w2231_,
		_w2267_,
		_w2268_
	);
	LUT2 #(
		.INIT('h2)
	) name2133 (
		_w183_,
		_w227_,
		_w2269_
	);
	LUT2 #(
		.INIT('h2)
	) name2134 (
		_w228_,
		_w317_,
		_w2270_
	);
	LUT2 #(
		.INIT('h2)
	) name2135 (
		_w273_,
		_w366_,
		_w2271_
	);
	LUT2 #(
		.INIT('h4)
	) name2136 (
		_w272_,
		_w318_,
		_w2272_
	);
	LUT2 #(
		.INIT('h1)
	) name2137 (
		_w2269_,
		_w2270_,
		_w2273_
	);
	LUT2 #(
		.INIT('h1)
	) name2138 (
		_w2271_,
		_w2272_,
		_w2274_
	);
	LUT2 #(
		.INIT('h8)
	) name2139 (
		_w2273_,
		_w2274_,
		_w2275_
	);
	LUT2 #(
		.INIT('h1)
	) name2140 (
		\shift[6] ,
		_w2275_,
		_w2276_
	);
	LUT2 #(
		.INIT('h4)
	) name2141 (
		_w182_,
		_w273_,
		_w2277_
	);
	LUT2 #(
		.INIT('h2)
	) name2142 (
		_w183_,
		_w410_,
		_w2278_
	);
	LUT2 #(
		.INIT('h2)
	) name2143 (
		_w318_,
		_w454_,
		_w2279_
	);
	LUT2 #(
		.INIT('h2)
	) name2144 (
		_w228_,
		_w500_,
		_w2280_
	);
	LUT2 #(
		.INIT('h1)
	) name2145 (
		_w2277_,
		_w2278_,
		_w2281_
	);
	LUT2 #(
		.INIT('h1)
	) name2146 (
		_w2279_,
		_w2280_,
		_w2282_
	);
	LUT2 #(
		.INIT('h8)
	) name2147 (
		_w2281_,
		_w2282_,
		_w2283_
	);
	LUT2 #(
		.INIT('h2)
	) name2148 (
		\shift[6] ,
		_w2283_,
		_w2284_
	);
	LUT2 #(
		.INIT('h1)
	) name2149 (
		_w2276_,
		_w2284_,
		_w2285_
	);
	LUT2 #(
		.INIT('h2)
	) name2150 (
		_w183_,
		_w609_,
		_w2286_
	);
	LUT2 #(
		.INIT('h2)
	) name2151 (
		_w228_,
		_w713_,
		_w2287_
	);
	LUT2 #(
		.INIT('h2)
	) name2152 (
		_w273_,
		_w821_,
		_w2288_
	);
	LUT2 #(
		.INIT('h2)
	) name2153 (
		_w318_,
		_w661_,
		_w2289_
	);
	LUT2 #(
		.INIT('h1)
	) name2154 (
		_w2286_,
		_w2287_,
		_w2290_
	);
	LUT2 #(
		.INIT('h1)
	) name2155 (
		_w2288_,
		_w2289_,
		_w2291_
	);
	LUT2 #(
		.INIT('h8)
	) name2156 (
		_w2290_,
		_w2291_,
		_w2292_
	);
	LUT2 #(
		.INIT('h1)
	) name2157 (
		\shift[6] ,
		_w2292_,
		_w2293_
	);
	LUT2 #(
		.INIT('h2)
	) name2158 (
		_w318_,
		_w769_,
		_w2294_
	);
	LUT2 #(
		.INIT('h2)
	) name2159 (
		_w273_,
		_w557_,
		_w2295_
	);
	LUT2 #(
		.INIT('h2)
	) name2160 (
		_w228_,
		_w869_,
		_w2296_
	);
	LUT2 #(
		.INIT('h2)
	) name2161 (
		_w183_,
		_w921_,
		_w2297_
	);
	LUT2 #(
		.INIT('h1)
	) name2162 (
		_w2294_,
		_w2295_,
		_w2298_
	);
	LUT2 #(
		.INIT('h1)
	) name2163 (
		_w2296_,
		_w2297_,
		_w2299_
	);
	LUT2 #(
		.INIT('h8)
	) name2164 (
		_w2298_,
		_w2299_,
		_w2300_
	);
	LUT2 #(
		.INIT('h2)
	) name2165 (
		\shift[6] ,
		_w2300_,
		_w2301_
	);
	LUT2 #(
		.INIT('h1)
	) name2166 (
		_w2293_,
		_w2301_,
		_w2302_
	);
	LUT2 #(
		.INIT('h2)
	) name2167 (
		_w183_,
		_w966_,
		_w2303_
	);
	LUT2 #(
		.INIT('h2)
	) name2168 (
		_w228_,
		_w1006_,
		_w2304_
	);
	LUT2 #(
		.INIT('h2)
	) name2169 (
		_w273_,
		_w1050_,
		_w2305_
	);
	LUT2 #(
		.INIT('h2)
	) name2170 (
		_w318_,
		_w986_,
		_w2306_
	);
	LUT2 #(
		.INIT('h1)
	) name2171 (
		_w2303_,
		_w2304_,
		_w2307_
	);
	LUT2 #(
		.INIT('h1)
	) name2172 (
		_w2305_,
		_w2306_,
		_w2308_
	);
	LUT2 #(
		.INIT('h8)
	) name2173 (
		_w2307_,
		_w2308_,
		_w2309_
	);
	LUT2 #(
		.INIT('h1)
	) name2174 (
		\shift[6] ,
		_w2309_,
		_w2310_
	);
	LUT2 #(
		.INIT('h2)
	) name2175 (
		_w318_,
		_w1030_,
		_w2311_
	);
	LUT2 #(
		.INIT('h2)
	) name2176 (
		_w273_,
		_w946_,
		_w2312_
	);
	LUT2 #(
		.INIT('h2)
	) name2177 (
		_w228_,
		_w1072_,
		_w2313_
	);
	LUT2 #(
		.INIT('h2)
	) name2178 (
		_w183_,
		_w1092_,
		_w2314_
	);
	LUT2 #(
		.INIT('h1)
	) name2179 (
		_w2311_,
		_w2312_,
		_w2315_
	);
	LUT2 #(
		.INIT('h1)
	) name2180 (
		_w2313_,
		_w2314_,
		_w2316_
	);
	LUT2 #(
		.INIT('h8)
	) name2181 (
		_w2315_,
		_w2316_,
		_w2317_
	);
	LUT2 #(
		.INIT('h2)
	) name2182 (
		\shift[6] ,
		_w2317_,
		_w2318_
	);
	LUT2 #(
		.INIT('h1)
	) name2183 (
		_w2310_,
		_w2318_,
		_w2319_
	);
	LUT2 #(
		.INIT('h2)
	) name2184 (
		_w228_,
		_w1133_,
		_w2320_
	);
	LUT2 #(
		.INIT('h2)
	) name2185 (
		_w183_,
		_w1169_,
		_w2321_
	);
	LUT2 #(
		.INIT('h2)
	) name2186 (
		_w318_,
		_w1205_,
		_w2322_
	);
	LUT2 #(
		.INIT('h2)
	) name2187 (
		_w273_,
		_w1350_,
		_w2323_
	);
	LUT2 #(
		.INIT('h1)
	) name2188 (
		_w2320_,
		_w2321_,
		_w2324_
	);
	LUT2 #(
		.INIT('h1)
	) name2189 (
		_w2322_,
		_w2323_,
		_w2325_
	);
	LUT2 #(
		.INIT('h8)
	) name2190 (
		_w2324_,
		_w2325_,
		_w2326_
	);
	LUT2 #(
		.INIT('h1)
	) name2191 (
		\shift[6] ,
		_w2326_,
		_w2327_
	);
	LUT2 #(
		.INIT('h2)
	) name2192 (
		_w318_,
		_w1281_,
		_w2328_
	);
	LUT2 #(
		.INIT('h2)
	) name2193 (
		_w273_,
		_w1241_,
		_w2329_
	);
	LUT2 #(
		.INIT('h2)
	) name2194 (
		_w183_,
		_w1386_,
		_w2330_
	);
	LUT2 #(
		.INIT('h2)
	) name2195 (
		_w228_,
		_w1314_,
		_w2331_
	);
	LUT2 #(
		.INIT('h1)
	) name2196 (
		_w2328_,
		_w2329_,
		_w2332_
	);
	LUT2 #(
		.INIT('h1)
	) name2197 (
		_w2330_,
		_w2331_,
		_w2333_
	);
	LUT2 #(
		.INIT('h8)
	) name2198 (
		_w2332_,
		_w2333_,
		_w2334_
	);
	LUT2 #(
		.INIT('h2)
	) name2199 (
		\shift[6] ,
		_w2334_,
		_w2335_
	);
	LUT2 #(
		.INIT('h1)
	) name2200 (
		_w2327_,
		_w2335_,
		_w2336_
	);
	LUT2 #(
		.INIT('h2)
	) name2201 (
		_w183_,
		_w1407_,
		_w2337_
	);
	LUT2 #(
		.INIT('h2)
	) name2202 (
		_w228_,
		_w1423_,
		_w2338_
	);
	LUT2 #(
		.INIT('h2)
	) name2203 (
		_w273_,
		_w1459_,
		_w2339_
	);
	LUT2 #(
		.INIT('h2)
	) name2204 (
		_w318_,
		_w1415_,
		_w2340_
	);
	LUT2 #(
		.INIT('h1)
	) name2205 (
		_w2337_,
		_w2338_,
		_w2341_
	);
	LUT2 #(
		.INIT('h1)
	) name2206 (
		_w2339_,
		_w2340_,
		_w2342_
	);
	LUT2 #(
		.INIT('h8)
	) name2207 (
		_w2341_,
		_w2342_,
		_w2343_
	);
	LUT2 #(
		.INIT('h1)
	) name2208 (
		\shift[6] ,
		_w2343_,
		_w2344_
	);
	LUT2 #(
		.INIT('h2)
	) name2209 (
		_w273_,
		_w1399_,
		_w2345_
	);
	LUT2 #(
		.INIT('h2)
	) name2210 (
		_w228_,
		_w1435_,
		_w2346_
	);
	LUT2 #(
		.INIT('h2)
	) name2211 (
		_w183_,
		_w1451_,
		_w2347_
	);
	LUT2 #(
		.INIT('h2)
	) name2212 (
		_w318_,
		_w1443_,
		_w2348_
	);
	LUT2 #(
		.INIT('h1)
	) name2213 (
		_w2345_,
		_w2346_,
		_w2349_
	);
	LUT2 #(
		.INIT('h1)
	) name2214 (
		_w2347_,
		_w2348_,
		_w2350_
	);
	LUT2 #(
		.INIT('h8)
	) name2215 (
		_w2349_,
		_w2350_,
		_w2351_
	);
	LUT2 #(
		.INIT('h2)
	) name2216 (
		\shift[6] ,
		_w2351_,
		_w2352_
	);
	LUT2 #(
		.INIT('h1)
	) name2217 (
		_w2344_,
		_w2352_,
		_w2353_
	);
	LUT2 #(
		.INIT('h2)
	) name2218 (
		_w183_,
		_w1480_,
		_w2354_
	);
	LUT2 #(
		.INIT('h2)
	) name2219 (
		_w228_,
		_w1496_,
		_w2355_
	);
	LUT2 #(
		.INIT('h2)
	) name2220 (
		_w273_,
		_w1532_,
		_w2356_
	);
	LUT2 #(
		.INIT('h2)
	) name2221 (
		_w318_,
		_w1488_,
		_w2357_
	);
	LUT2 #(
		.INIT('h1)
	) name2222 (
		_w2354_,
		_w2355_,
		_w2358_
	);
	LUT2 #(
		.INIT('h1)
	) name2223 (
		_w2356_,
		_w2357_,
		_w2359_
	);
	LUT2 #(
		.INIT('h8)
	) name2224 (
		_w2358_,
		_w2359_,
		_w2360_
	);
	LUT2 #(
		.INIT('h1)
	) name2225 (
		\shift[6] ,
		_w2360_,
		_w2361_
	);
	LUT2 #(
		.INIT('h2)
	) name2226 (
		_w273_,
		_w1472_,
		_w2362_
	);
	LUT2 #(
		.INIT('h2)
	) name2227 (
		_w228_,
		_w1508_,
		_w2363_
	);
	LUT2 #(
		.INIT('h2)
	) name2228 (
		_w183_,
		_w1524_,
		_w2364_
	);
	LUT2 #(
		.INIT('h2)
	) name2229 (
		_w318_,
		_w1516_,
		_w2365_
	);
	LUT2 #(
		.INIT('h1)
	) name2230 (
		_w2362_,
		_w2363_,
		_w2366_
	);
	LUT2 #(
		.INIT('h1)
	) name2231 (
		_w2364_,
		_w2365_,
		_w2367_
	);
	LUT2 #(
		.INIT('h8)
	) name2232 (
		_w2366_,
		_w2367_,
		_w2368_
	);
	LUT2 #(
		.INIT('h2)
	) name2233 (
		\shift[6] ,
		_w2368_,
		_w2369_
	);
	LUT2 #(
		.INIT('h1)
	) name2234 (
		_w2361_,
		_w2369_,
		_w2370_
	);
	LUT2 #(
		.INIT('h2)
	) name2235 (
		_w183_,
		_w1553_,
		_w2371_
	);
	LUT2 #(
		.INIT('h2)
	) name2236 (
		_w228_,
		_w1569_,
		_w2372_
	);
	LUT2 #(
		.INIT('h2)
	) name2237 (
		_w273_,
		_w1605_,
		_w2373_
	);
	LUT2 #(
		.INIT('h2)
	) name2238 (
		_w318_,
		_w1561_,
		_w2374_
	);
	LUT2 #(
		.INIT('h1)
	) name2239 (
		_w2371_,
		_w2372_,
		_w2375_
	);
	LUT2 #(
		.INIT('h1)
	) name2240 (
		_w2373_,
		_w2374_,
		_w2376_
	);
	LUT2 #(
		.INIT('h8)
	) name2241 (
		_w2375_,
		_w2376_,
		_w2377_
	);
	LUT2 #(
		.INIT('h1)
	) name2242 (
		\shift[6] ,
		_w2377_,
		_w2378_
	);
	LUT2 #(
		.INIT('h2)
	) name2243 (
		_w273_,
		_w1545_,
		_w2379_
	);
	LUT2 #(
		.INIT('h2)
	) name2244 (
		_w228_,
		_w1581_,
		_w2380_
	);
	LUT2 #(
		.INIT('h2)
	) name2245 (
		_w183_,
		_w1597_,
		_w2381_
	);
	LUT2 #(
		.INIT('h2)
	) name2246 (
		_w318_,
		_w1589_,
		_w2382_
	);
	LUT2 #(
		.INIT('h1)
	) name2247 (
		_w2379_,
		_w2380_,
		_w2383_
	);
	LUT2 #(
		.INIT('h1)
	) name2248 (
		_w2381_,
		_w2382_,
		_w2384_
	);
	LUT2 #(
		.INIT('h8)
	) name2249 (
		_w2383_,
		_w2384_,
		_w2385_
	);
	LUT2 #(
		.INIT('h2)
	) name2250 (
		\shift[6] ,
		_w2385_,
		_w2386_
	);
	LUT2 #(
		.INIT('h1)
	) name2251 (
		_w2378_,
		_w2386_,
		_w2387_
	);
	LUT2 #(
		.INIT('h2)
	) name2252 (
		_w183_,
		_w1626_,
		_w2388_
	);
	LUT2 #(
		.INIT('h2)
	) name2253 (
		_w273_,
		_w1678_,
		_w2389_
	);
	LUT2 #(
		.INIT('h2)
	) name2254 (
		_w318_,
		_w1634_,
		_w2390_
	);
	LUT2 #(
		.INIT('h2)
	) name2255 (
		_w228_,
		_w1642_,
		_w2391_
	);
	LUT2 #(
		.INIT('h1)
	) name2256 (
		_w2388_,
		_w2389_,
		_w2392_
	);
	LUT2 #(
		.INIT('h1)
	) name2257 (
		_w2390_,
		_w2391_,
		_w2393_
	);
	LUT2 #(
		.INIT('h8)
	) name2258 (
		_w2392_,
		_w2393_,
		_w2394_
	);
	LUT2 #(
		.INIT('h1)
	) name2259 (
		\shift[6] ,
		_w2394_,
		_w2395_
	);
	LUT2 #(
		.INIT('h2)
	) name2260 (
		_w228_,
		_w1654_,
		_w2396_
	);
	LUT2 #(
		.INIT('h2)
	) name2261 (
		_w318_,
		_w1662_,
		_w2397_
	);
	LUT2 #(
		.INIT('h2)
	) name2262 (
		_w183_,
		_w1670_,
		_w2398_
	);
	LUT2 #(
		.INIT('h2)
	) name2263 (
		_w273_,
		_w1618_,
		_w2399_
	);
	LUT2 #(
		.INIT('h1)
	) name2264 (
		_w2396_,
		_w2397_,
		_w2400_
	);
	LUT2 #(
		.INIT('h1)
	) name2265 (
		_w2398_,
		_w2399_,
		_w2401_
	);
	LUT2 #(
		.INIT('h8)
	) name2266 (
		_w2400_,
		_w2401_,
		_w2402_
	);
	LUT2 #(
		.INIT('h2)
	) name2267 (
		\shift[6] ,
		_w2402_,
		_w2403_
	);
	LUT2 #(
		.INIT('h1)
	) name2268 (
		_w2395_,
		_w2403_,
		_w2404_
	);
	LUT2 #(
		.INIT('h2)
	) name2269 (
		_w183_,
		_w1699_,
		_w2405_
	);
	LUT2 #(
		.INIT('h2)
	) name2270 (
		_w273_,
		_w1751_,
		_w2406_
	);
	LUT2 #(
		.INIT('h2)
	) name2271 (
		_w318_,
		_w1707_,
		_w2407_
	);
	LUT2 #(
		.INIT('h2)
	) name2272 (
		_w228_,
		_w1715_,
		_w2408_
	);
	LUT2 #(
		.INIT('h1)
	) name2273 (
		_w2405_,
		_w2406_,
		_w2409_
	);
	LUT2 #(
		.INIT('h1)
	) name2274 (
		_w2407_,
		_w2408_,
		_w2410_
	);
	LUT2 #(
		.INIT('h8)
	) name2275 (
		_w2409_,
		_w2410_,
		_w2411_
	);
	LUT2 #(
		.INIT('h1)
	) name2276 (
		\shift[6] ,
		_w2411_,
		_w2412_
	);
	LUT2 #(
		.INIT('h2)
	) name2277 (
		_w228_,
		_w1727_,
		_w2413_
	);
	LUT2 #(
		.INIT('h2)
	) name2278 (
		_w318_,
		_w1735_,
		_w2414_
	);
	LUT2 #(
		.INIT('h2)
	) name2279 (
		_w183_,
		_w1743_,
		_w2415_
	);
	LUT2 #(
		.INIT('h2)
	) name2280 (
		_w273_,
		_w1691_,
		_w2416_
	);
	LUT2 #(
		.INIT('h1)
	) name2281 (
		_w2413_,
		_w2414_,
		_w2417_
	);
	LUT2 #(
		.INIT('h1)
	) name2282 (
		_w2415_,
		_w2416_,
		_w2418_
	);
	LUT2 #(
		.INIT('h8)
	) name2283 (
		_w2417_,
		_w2418_,
		_w2419_
	);
	LUT2 #(
		.INIT('h2)
	) name2284 (
		\shift[6] ,
		_w2419_,
		_w2420_
	);
	LUT2 #(
		.INIT('h1)
	) name2285 (
		_w2412_,
		_w2420_,
		_w2421_
	);
	LUT2 #(
		.INIT('h2)
	) name2286 (
		_w183_,
		_w1772_,
		_w2422_
	);
	LUT2 #(
		.INIT('h2)
	) name2287 (
		_w273_,
		_w1824_,
		_w2423_
	);
	LUT2 #(
		.INIT('h2)
	) name2288 (
		_w318_,
		_w1780_,
		_w2424_
	);
	LUT2 #(
		.INIT('h2)
	) name2289 (
		_w228_,
		_w1788_,
		_w2425_
	);
	LUT2 #(
		.INIT('h1)
	) name2290 (
		_w2422_,
		_w2423_,
		_w2426_
	);
	LUT2 #(
		.INIT('h1)
	) name2291 (
		_w2424_,
		_w2425_,
		_w2427_
	);
	LUT2 #(
		.INIT('h8)
	) name2292 (
		_w2426_,
		_w2427_,
		_w2428_
	);
	LUT2 #(
		.INIT('h1)
	) name2293 (
		\shift[6] ,
		_w2428_,
		_w2429_
	);
	LUT2 #(
		.INIT('h2)
	) name2294 (
		_w228_,
		_w1800_,
		_w2430_
	);
	LUT2 #(
		.INIT('h2)
	) name2295 (
		_w318_,
		_w1808_,
		_w2431_
	);
	LUT2 #(
		.INIT('h2)
	) name2296 (
		_w183_,
		_w1816_,
		_w2432_
	);
	LUT2 #(
		.INIT('h2)
	) name2297 (
		_w273_,
		_w1764_,
		_w2433_
	);
	LUT2 #(
		.INIT('h1)
	) name2298 (
		_w2430_,
		_w2431_,
		_w2434_
	);
	LUT2 #(
		.INIT('h1)
	) name2299 (
		_w2432_,
		_w2433_,
		_w2435_
	);
	LUT2 #(
		.INIT('h8)
	) name2300 (
		_w2434_,
		_w2435_,
		_w2436_
	);
	LUT2 #(
		.INIT('h2)
	) name2301 (
		\shift[6] ,
		_w2436_,
		_w2437_
	);
	LUT2 #(
		.INIT('h1)
	) name2302 (
		_w2429_,
		_w2437_,
		_w2438_
	);
	LUT2 #(
		.INIT('h2)
	) name2303 (
		_w183_,
		_w1845_,
		_w2439_
	);
	LUT2 #(
		.INIT('h2)
	) name2304 (
		_w228_,
		_w1861_,
		_w2440_
	);
	LUT2 #(
		.INIT('h2)
	) name2305 (
		_w273_,
		_w1897_,
		_w2441_
	);
	LUT2 #(
		.INIT('h2)
	) name2306 (
		_w318_,
		_w1853_,
		_w2442_
	);
	LUT2 #(
		.INIT('h1)
	) name2307 (
		_w2439_,
		_w2440_,
		_w2443_
	);
	LUT2 #(
		.INIT('h1)
	) name2308 (
		_w2441_,
		_w2442_,
		_w2444_
	);
	LUT2 #(
		.INIT('h8)
	) name2309 (
		_w2443_,
		_w2444_,
		_w2445_
	);
	LUT2 #(
		.INIT('h1)
	) name2310 (
		\shift[6] ,
		_w2445_,
		_w2446_
	);
	LUT2 #(
		.INIT('h2)
	) name2311 (
		_w228_,
		_w1873_,
		_w2447_
	);
	LUT2 #(
		.INIT('h2)
	) name2312 (
		_w318_,
		_w1881_,
		_w2448_
	);
	LUT2 #(
		.INIT('h2)
	) name2313 (
		_w183_,
		_w1889_,
		_w2449_
	);
	LUT2 #(
		.INIT('h2)
	) name2314 (
		_w273_,
		_w1837_,
		_w2450_
	);
	LUT2 #(
		.INIT('h1)
	) name2315 (
		_w2447_,
		_w2448_,
		_w2451_
	);
	LUT2 #(
		.INIT('h1)
	) name2316 (
		_w2449_,
		_w2450_,
		_w2452_
	);
	LUT2 #(
		.INIT('h8)
	) name2317 (
		_w2451_,
		_w2452_,
		_w2453_
	);
	LUT2 #(
		.INIT('h2)
	) name2318 (
		\shift[6] ,
		_w2453_,
		_w2454_
	);
	LUT2 #(
		.INIT('h1)
	) name2319 (
		_w2446_,
		_w2454_,
		_w2455_
	);
	LUT2 #(
		.INIT('h2)
	) name2320 (
		_w183_,
		_w1918_,
		_w2456_
	);
	LUT2 #(
		.INIT('h2)
	) name2321 (
		_w228_,
		_w1934_,
		_w2457_
	);
	LUT2 #(
		.INIT('h2)
	) name2322 (
		_w273_,
		_w1970_,
		_w2458_
	);
	LUT2 #(
		.INIT('h2)
	) name2323 (
		_w318_,
		_w1926_,
		_w2459_
	);
	LUT2 #(
		.INIT('h1)
	) name2324 (
		_w2456_,
		_w2457_,
		_w2460_
	);
	LUT2 #(
		.INIT('h1)
	) name2325 (
		_w2458_,
		_w2459_,
		_w2461_
	);
	LUT2 #(
		.INIT('h8)
	) name2326 (
		_w2460_,
		_w2461_,
		_w2462_
	);
	LUT2 #(
		.INIT('h1)
	) name2327 (
		\shift[6] ,
		_w2462_,
		_w2463_
	);
	LUT2 #(
		.INIT('h2)
	) name2328 (
		_w228_,
		_w1946_,
		_w2464_
	);
	LUT2 #(
		.INIT('h2)
	) name2329 (
		_w318_,
		_w1954_,
		_w2465_
	);
	LUT2 #(
		.INIT('h2)
	) name2330 (
		_w183_,
		_w1962_,
		_w2466_
	);
	LUT2 #(
		.INIT('h2)
	) name2331 (
		_w273_,
		_w1910_,
		_w2467_
	);
	LUT2 #(
		.INIT('h1)
	) name2332 (
		_w2464_,
		_w2465_,
		_w2468_
	);
	LUT2 #(
		.INIT('h1)
	) name2333 (
		_w2466_,
		_w2467_,
		_w2469_
	);
	LUT2 #(
		.INIT('h8)
	) name2334 (
		_w2468_,
		_w2469_,
		_w2470_
	);
	LUT2 #(
		.INIT('h2)
	) name2335 (
		\shift[6] ,
		_w2470_,
		_w2471_
	);
	LUT2 #(
		.INIT('h1)
	) name2336 (
		_w2463_,
		_w2471_,
		_w2472_
	);
	LUT2 #(
		.INIT('h2)
	) name2337 (
		_w183_,
		_w1991_,
		_w2473_
	);
	LUT2 #(
		.INIT('h2)
	) name2338 (
		_w228_,
		_w2007_,
		_w2474_
	);
	LUT2 #(
		.INIT('h2)
	) name2339 (
		_w273_,
		_w2043_,
		_w2475_
	);
	LUT2 #(
		.INIT('h2)
	) name2340 (
		_w318_,
		_w1999_,
		_w2476_
	);
	LUT2 #(
		.INIT('h1)
	) name2341 (
		_w2473_,
		_w2474_,
		_w2477_
	);
	LUT2 #(
		.INIT('h1)
	) name2342 (
		_w2475_,
		_w2476_,
		_w2478_
	);
	LUT2 #(
		.INIT('h8)
	) name2343 (
		_w2477_,
		_w2478_,
		_w2479_
	);
	LUT2 #(
		.INIT('h1)
	) name2344 (
		\shift[6] ,
		_w2479_,
		_w2480_
	);
	LUT2 #(
		.INIT('h2)
	) name2345 (
		_w228_,
		_w2019_,
		_w2481_
	);
	LUT2 #(
		.INIT('h2)
	) name2346 (
		_w318_,
		_w2027_,
		_w2482_
	);
	LUT2 #(
		.INIT('h2)
	) name2347 (
		_w183_,
		_w2035_,
		_w2483_
	);
	LUT2 #(
		.INIT('h2)
	) name2348 (
		_w273_,
		_w1983_,
		_w2484_
	);
	LUT2 #(
		.INIT('h1)
	) name2349 (
		_w2481_,
		_w2482_,
		_w2485_
	);
	LUT2 #(
		.INIT('h1)
	) name2350 (
		_w2483_,
		_w2484_,
		_w2486_
	);
	LUT2 #(
		.INIT('h8)
	) name2351 (
		_w2485_,
		_w2486_,
		_w2487_
	);
	LUT2 #(
		.INIT('h2)
	) name2352 (
		\shift[6] ,
		_w2487_,
		_w2488_
	);
	LUT2 #(
		.INIT('h1)
	) name2353 (
		_w2480_,
		_w2488_,
		_w2489_
	);
	LUT2 #(
		.INIT('h2)
	) name2354 (
		_w183_,
		_w2064_,
		_w2490_
	);
	LUT2 #(
		.INIT('h2)
	) name2355 (
		_w228_,
		_w2080_,
		_w2491_
	);
	LUT2 #(
		.INIT('h2)
	) name2356 (
		_w273_,
		_w2116_,
		_w2492_
	);
	LUT2 #(
		.INIT('h2)
	) name2357 (
		_w318_,
		_w2072_,
		_w2493_
	);
	LUT2 #(
		.INIT('h1)
	) name2358 (
		_w2490_,
		_w2491_,
		_w2494_
	);
	LUT2 #(
		.INIT('h1)
	) name2359 (
		_w2492_,
		_w2493_,
		_w2495_
	);
	LUT2 #(
		.INIT('h8)
	) name2360 (
		_w2494_,
		_w2495_,
		_w2496_
	);
	LUT2 #(
		.INIT('h1)
	) name2361 (
		\shift[6] ,
		_w2496_,
		_w2497_
	);
	LUT2 #(
		.INIT('h2)
	) name2362 (
		_w228_,
		_w2092_,
		_w2498_
	);
	LUT2 #(
		.INIT('h2)
	) name2363 (
		_w318_,
		_w2100_,
		_w2499_
	);
	LUT2 #(
		.INIT('h2)
	) name2364 (
		_w183_,
		_w2108_,
		_w2500_
	);
	LUT2 #(
		.INIT('h2)
	) name2365 (
		_w273_,
		_w2056_,
		_w2501_
	);
	LUT2 #(
		.INIT('h1)
	) name2366 (
		_w2498_,
		_w2499_,
		_w2502_
	);
	LUT2 #(
		.INIT('h1)
	) name2367 (
		_w2500_,
		_w2501_,
		_w2503_
	);
	LUT2 #(
		.INIT('h8)
	) name2368 (
		_w2502_,
		_w2503_,
		_w2504_
	);
	LUT2 #(
		.INIT('h2)
	) name2369 (
		\shift[6] ,
		_w2504_,
		_w2505_
	);
	LUT2 #(
		.INIT('h1)
	) name2370 (
		_w2497_,
		_w2505_,
		_w2506_
	);
	LUT2 #(
		.INIT('h2)
	) name2371 (
		_w183_,
		_w2137_,
		_w2507_
	);
	LUT2 #(
		.INIT('h2)
	) name2372 (
		_w228_,
		_w2153_,
		_w2508_
	);
	LUT2 #(
		.INIT('h2)
	) name2373 (
		_w273_,
		_w2189_,
		_w2509_
	);
	LUT2 #(
		.INIT('h2)
	) name2374 (
		_w318_,
		_w2145_,
		_w2510_
	);
	LUT2 #(
		.INIT('h1)
	) name2375 (
		_w2507_,
		_w2508_,
		_w2511_
	);
	LUT2 #(
		.INIT('h1)
	) name2376 (
		_w2509_,
		_w2510_,
		_w2512_
	);
	LUT2 #(
		.INIT('h8)
	) name2377 (
		_w2511_,
		_w2512_,
		_w2513_
	);
	LUT2 #(
		.INIT('h1)
	) name2378 (
		\shift[6] ,
		_w2513_,
		_w2514_
	);
	LUT2 #(
		.INIT('h2)
	) name2379 (
		_w228_,
		_w2165_,
		_w2515_
	);
	LUT2 #(
		.INIT('h2)
	) name2380 (
		_w318_,
		_w2173_,
		_w2516_
	);
	LUT2 #(
		.INIT('h2)
	) name2381 (
		_w183_,
		_w2181_,
		_w2517_
	);
	LUT2 #(
		.INIT('h2)
	) name2382 (
		_w273_,
		_w2129_,
		_w2518_
	);
	LUT2 #(
		.INIT('h1)
	) name2383 (
		_w2515_,
		_w2516_,
		_w2519_
	);
	LUT2 #(
		.INIT('h1)
	) name2384 (
		_w2517_,
		_w2518_,
		_w2520_
	);
	LUT2 #(
		.INIT('h8)
	) name2385 (
		_w2519_,
		_w2520_,
		_w2521_
	);
	LUT2 #(
		.INIT('h2)
	) name2386 (
		\shift[6] ,
		_w2521_,
		_w2522_
	);
	LUT2 #(
		.INIT('h1)
	) name2387 (
		_w2514_,
		_w2522_,
		_w2523_
	);
	LUT2 #(
		.INIT('h2)
	) name2388 (
		_w183_,
		_w2210_,
		_w2524_
	);
	LUT2 #(
		.INIT('h2)
	) name2389 (
		_w228_,
		_w2226_,
		_w2525_
	);
	LUT2 #(
		.INIT('h2)
	) name2390 (
		_w273_,
		_w2262_,
		_w2526_
	);
	LUT2 #(
		.INIT('h2)
	) name2391 (
		_w318_,
		_w2218_,
		_w2527_
	);
	LUT2 #(
		.INIT('h1)
	) name2392 (
		_w2524_,
		_w2525_,
		_w2528_
	);
	LUT2 #(
		.INIT('h1)
	) name2393 (
		_w2526_,
		_w2527_,
		_w2529_
	);
	LUT2 #(
		.INIT('h8)
	) name2394 (
		_w2528_,
		_w2529_,
		_w2530_
	);
	LUT2 #(
		.INIT('h1)
	) name2395 (
		\shift[6] ,
		_w2530_,
		_w2531_
	);
	LUT2 #(
		.INIT('h2)
	) name2396 (
		_w228_,
		_w2238_,
		_w2532_
	);
	LUT2 #(
		.INIT('h2)
	) name2397 (
		_w318_,
		_w2246_,
		_w2533_
	);
	LUT2 #(
		.INIT('h2)
	) name2398 (
		_w183_,
		_w2254_,
		_w2534_
	);
	LUT2 #(
		.INIT('h2)
	) name2399 (
		_w273_,
		_w2202_,
		_w2535_
	);
	LUT2 #(
		.INIT('h1)
	) name2400 (
		_w2532_,
		_w2533_,
		_w2536_
	);
	LUT2 #(
		.INIT('h1)
	) name2401 (
		_w2534_,
		_w2535_,
		_w2537_
	);
	LUT2 #(
		.INIT('h8)
	) name2402 (
		_w2536_,
		_w2537_,
		_w2538_
	);
	LUT2 #(
		.INIT('h2)
	) name2403 (
		\shift[6] ,
		_w2538_,
		_w2539_
	);
	LUT2 #(
		.INIT('h1)
	) name2404 (
		_w2531_,
		_w2539_,
		_w2540_
	);
	LUT2 #(
		.INIT('h2)
	) name2405 (
		_w183_,
		_w317_,
		_w2541_
	);
	LUT2 #(
		.INIT('h2)
	) name2406 (
		_w228_,
		_w272_,
		_w2542_
	);
	LUT2 #(
		.INIT('h2)
	) name2407 (
		_w273_,
		_w410_,
		_w2543_
	);
	LUT2 #(
		.INIT('h2)
	) name2408 (
		_w318_,
		_w366_,
		_w2544_
	);
	LUT2 #(
		.INIT('h1)
	) name2409 (
		_w2541_,
		_w2542_,
		_w2545_
	);
	LUT2 #(
		.INIT('h1)
	) name2410 (
		_w2543_,
		_w2544_,
		_w2546_
	);
	LUT2 #(
		.INIT('h8)
	) name2411 (
		_w2545_,
		_w2546_,
		_w2547_
	);
	LUT2 #(
		.INIT('h1)
	) name2412 (
		\shift[6] ,
		_w2547_,
		_w2548_
	);
	LUT2 #(
		.INIT('h4)
	) name2413 (
		_w182_,
		_w318_,
		_w2549_
	);
	LUT2 #(
		.INIT('h4)
	) name2414 (
		_w227_,
		_w273_,
		_w2550_
	);
	LUT2 #(
		.INIT('h2)
	) name2415 (
		_w228_,
		_w454_,
		_w2551_
	);
	LUT2 #(
		.INIT('h2)
	) name2416 (
		_w183_,
		_w500_,
		_w2552_
	);
	LUT2 #(
		.INIT('h1)
	) name2417 (
		_w2549_,
		_w2550_,
		_w2553_
	);
	LUT2 #(
		.INIT('h1)
	) name2418 (
		_w2551_,
		_w2552_,
		_w2554_
	);
	LUT2 #(
		.INIT('h8)
	) name2419 (
		_w2553_,
		_w2554_,
		_w2555_
	);
	LUT2 #(
		.INIT('h2)
	) name2420 (
		\shift[6] ,
		_w2555_,
		_w2556_
	);
	LUT2 #(
		.INIT('h1)
	) name2421 (
		_w2548_,
		_w2556_,
		_w2557_
	);
	LUT2 #(
		.INIT('h2)
	) name2422 (
		_w183_,
		_w713_,
		_w2558_
	);
	LUT2 #(
		.INIT('h2)
	) name2423 (
		_w228_,
		_w661_,
		_w2559_
	);
	LUT2 #(
		.INIT('h2)
	) name2424 (
		_w273_,
		_w921_,
		_w2560_
	);
	LUT2 #(
		.INIT('h2)
	) name2425 (
		_w318_,
		_w821_,
		_w2561_
	);
	LUT2 #(
		.INIT('h1)
	) name2426 (
		_w2558_,
		_w2559_,
		_w2562_
	);
	LUT2 #(
		.INIT('h1)
	) name2427 (
		_w2560_,
		_w2561_,
		_w2563_
	);
	LUT2 #(
		.INIT('h8)
	) name2428 (
		_w2562_,
		_w2563_,
		_w2564_
	);
	LUT2 #(
		.INIT('h1)
	) name2429 (
		\shift[6] ,
		_w2564_,
		_w2565_
	);
	LUT2 #(
		.INIT('h2)
	) name2430 (
		_w228_,
		_w769_,
		_w2566_
	);
	LUT2 #(
		.INIT('h2)
	) name2431 (
		_w318_,
		_w557_,
		_w2567_
	);
	LUT2 #(
		.INIT('h2)
	) name2432 (
		_w183_,
		_w869_,
		_w2568_
	);
	LUT2 #(
		.INIT('h2)
	) name2433 (
		_w273_,
		_w609_,
		_w2569_
	);
	LUT2 #(
		.INIT('h1)
	) name2434 (
		_w2566_,
		_w2567_,
		_w2570_
	);
	LUT2 #(
		.INIT('h1)
	) name2435 (
		_w2568_,
		_w2569_,
		_w2571_
	);
	LUT2 #(
		.INIT('h8)
	) name2436 (
		_w2570_,
		_w2571_,
		_w2572_
	);
	LUT2 #(
		.INIT('h2)
	) name2437 (
		\shift[6] ,
		_w2572_,
		_w2573_
	);
	LUT2 #(
		.INIT('h1)
	) name2438 (
		_w2565_,
		_w2573_,
		_w2574_
	);
	LUT2 #(
		.INIT('h2)
	) name2439 (
		_w183_,
		_w1006_,
		_w2575_
	);
	LUT2 #(
		.INIT('h2)
	) name2440 (
		_w228_,
		_w986_,
		_w2576_
	);
	LUT2 #(
		.INIT('h2)
	) name2441 (
		_w273_,
		_w1092_,
		_w2577_
	);
	LUT2 #(
		.INIT('h2)
	) name2442 (
		_w318_,
		_w1050_,
		_w2578_
	);
	LUT2 #(
		.INIT('h1)
	) name2443 (
		_w2575_,
		_w2576_,
		_w2579_
	);
	LUT2 #(
		.INIT('h1)
	) name2444 (
		_w2577_,
		_w2578_,
		_w2580_
	);
	LUT2 #(
		.INIT('h8)
	) name2445 (
		_w2579_,
		_w2580_,
		_w2581_
	);
	LUT2 #(
		.INIT('h1)
	) name2446 (
		\shift[6] ,
		_w2581_,
		_w2582_
	);
	LUT2 #(
		.INIT('h2)
	) name2447 (
		_w228_,
		_w1030_,
		_w2583_
	);
	LUT2 #(
		.INIT('h2)
	) name2448 (
		_w318_,
		_w946_,
		_w2584_
	);
	LUT2 #(
		.INIT('h2)
	) name2449 (
		_w183_,
		_w1072_,
		_w2585_
	);
	LUT2 #(
		.INIT('h2)
	) name2450 (
		_w273_,
		_w966_,
		_w2586_
	);
	LUT2 #(
		.INIT('h1)
	) name2451 (
		_w2583_,
		_w2584_,
		_w2587_
	);
	LUT2 #(
		.INIT('h1)
	) name2452 (
		_w2585_,
		_w2586_,
		_w2588_
	);
	LUT2 #(
		.INIT('h8)
	) name2453 (
		_w2587_,
		_w2588_,
		_w2589_
	);
	LUT2 #(
		.INIT('h2)
	) name2454 (
		\shift[6] ,
		_w2589_,
		_w2590_
	);
	LUT2 #(
		.INIT('h1)
	) name2455 (
		_w2582_,
		_w2590_,
		_w2591_
	);
	LUT2 #(
		.INIT('h2)
	) name2456 (
		_w183_,
		_w1133_,
		_w2592_
	);
	LUT2 #(
		.INIT('h2)
	) name2457 (
		_w273_,
		_w1386_,
		_w2593_
	);
	LUT2 #(
		.INIT('h2)
	) name2458 (
		_w228_,
		_w1205_,
		_w2594_
	);
	LUT2 #(
		.INIT('h2)
	) name2459 (
		_w318_,
		_w1350_,
		_w2595_
	);
	LUT2 #(
		.INIT('h1)
	) name2460 (
		_w2592_,
		_w2593_,
		_w2596_
	);
	LUT2 #(
		.INIT('h1)
	) name2461 (
		_w2594_,
		_w2595_,
		_w2597_
	);
	LUT2 #(
		.INIT('h8)
	) name2462 (
		_w2596_,
		_w2597_,
		_w2598_
	);
	LUT2 #(
		.INIT('h1)
	) name2463 (
		\shift[6] ,
		_w2598_,
		_w2599_
	);
	LUT2 #(
		.INIT('h2)
	) name2464 (
		_w228_,
		_w1281_,
		_w2600_
	);
	LUT2 #(
		.INIT('h2)
	) name2465 (
		_w273_,
		_w1169_,
		_w2601_
	);
	LUT2 #(
		.INIT('h2)
	) name2466 (
		_w183_,
		_w1314_,
		_w2602_
	);
	LUT2 #(
		.INIT('h2)
	) name2467 (
		_w318_,
		_w1241_,
		_w2603_
	);
	LUT2 #(
		.INIT('h1)
	) name2468 (
		_w2600_,
		_w2601_,
		_w2604_
	);
	LUT2 #(
		.INIT('h1)
	) name2469 (
		_w2602_,
		_w2603_,
		_w2605_
	);
	LUT2 #(
		.INIT('h8)
	) name2470 (
		_w2604_,
		_w2605_,
		_w2606_
	);
	LUT2 #(
		.INIT('h2)
	) name2471 (
		\shift[6] ,
		_w2606_,
		_w2607_
	);
	LUT2 #(
		.INIT('h1)
	) name2472 (
		_w2599_,
		_w2607_,
		_w2608_
	);
	LUT2 #(
		.INIT('h2)
	) name2473 (
		_w183_,
		_w1423_,
		_w2609_
	);
	LUT2 #(
		.INIT('h2)
	) name2474 (
		_w228_,
		_w1415_,
		_w2610_
	);
	LUT2 #(
		.INIT('h2)
	) name2475 (
		_w273_,
		_w1451_,
		_w2611_
	);
	LUT2 #(
		.INIT('h2)
	) name2476 (
		_w318_,
		_w1459_,
		_w2612_
	);
	LUT2 #(
		.INIT('h1)
	) name2477 (
		_w2609_,
		_w2610_,
		_w2613_
	);
	LUT2 #(
		.INIT('h1)
	) name2478 (
		_w2611_,
		_w2612_,
		_w2614_
	);
	LUT2 #(
		.INIT('h8)
	) name2479 (
		_w2613_,
		_w2614_,
		_w2615_
	);
	LUT2 #(
		.INIT('h1)
	) name2480 (
		\shift[6] ,
		_w2615_,
		_w2616_
	);
	LUT2 #(
		.INIT('h2)
	) name2481 (
		_w318_,
		_w1399_,
		_w2617_
	);
	LUT2 #(
		.INIT('h2)
	) name2482 (
		_w273_,
		_w1407_,
		_w2618_
	);
	LUT2 #(
		.INIT('h2)
	) name2483 (
		_w228_,
		_w1443_,
		_w2619_
	);
	LUT2 #(
		.INIT('h2)
	) name2484 (
		_w183_,
		_w1435_,
		_w2620_
	);
	LUT2 #(
		.INIT('h1)
	) name2485 (
		_w2617_,
		_w2618_,
		_w2621_
	);
	LUT2 #(
		.INIT('h1)
	) name2486 (
		_w2619_,
		_w2620_,
		_w2622_
	);
	LUT2 #(
		.INIT('h8)
	) name2487 (
		_w2621_,
		_w2622_,
		_w2623_
	);
	LUT2 #(
		.INIT('h2)
	) name2488 (
		\shift[6] ,
		_w2623_,
		_w2624_
	);
	LUT2 #(
		.INIT('h1)
	) name2489 (
		_w2616_,
		_w2624_,
		_w2625_
	);
	LUT2 #(
		.INIT('h2)
	) name2490 (
		_w183_,
		_w1496_,
		_w2626_
	);
	LUT2 #(
		.INIT('h2)
	) name2491 (
		_w228_,
		_w1488_,
		_w2627_
	);
	LUT2 #(
		.INIT('h2)
	) name2492 (
		_w273_,
		_w1524_,
		_w2628_
	);
	LUT2 #(
		.INIT('h2)
	) name2493 (
		_w318_,
		_w1532_,
		_w2629_
	);
	LUT2 #(
		.INIT('h1)
	) name2494 (
		_w2626_,
		_w2627_,
		_w2630_
	);
	LUT2 #(
		.INIT('h1)
	) name2495 (
		_w2628_,
		_w2629_,
		_w2631_
	);
	LUT2 #(
		.INIT('h8)
	) name2496 (
		_w2630_,
		_w2631_,
		_w2632_
	);
	LUT2 #(
		.INIT('h1)
	) name2497 (
		\shift[6] ,
		_w2632_,
		_w2633_
	);
	LUT2 #(
		.INIT('h2)
	) name2498 (
		_w318_,
		_w1472_,
		_w2634_
	);
	LUT2 #(
		.INIT('h2)
	) name2499 (
		_w273_,
		_w1480_,
		_w2635_
	);
	LUT2 #(
		.INIT('h2)
	) name2500 (
		_w228_,
		_w1516_,
		_w2636_
	);
	LUT2 #(
		.INIT('h2)
	) name2501 (
		_w183_,
		_w1508_,
		_w2637_
	);
	LUT2 #(
		.INIT('h1)
	) name2502 (
		_w2634_,
		_w2635_,
		_w2638_
	);
	LUT2 #(
		.INIT('h1)
	) name2503 (
		_w2636_,
		_w2637_,
		_w2639_
	);
	LUT2 #(
		.INIT('h8)
	) name2504 (
		_w2638_,
		_w2639_,
		_w2640_
	);
	LUT2 #(
		.INIT('h2)
	) name2505 (
		\shift[6] ,
		_w2640_,
		_w2641_
	);
	LUT2 #(
		.INIT('h1)
	) name2506 (
		_w2633_,
		_w2641_,
		_w2642_
	);
	LUT2 #(
		.INIT('h2)
	) name2507 (
		_w183_,
		_w1569_,
		_w2643_
	);
	LUT2 #(
		.INIT('h2)
	) name2508 (
		_w228_,
		_w1561_,
		_w2644_
	);
	LUT2 #(
		.INIT('h2)
	) name2509 (
		_w273_,
		_w1597_,
		_w2645_
	);
	LUT2 #(
		.INIT('h2)
	) name2510 (
		_w318_,
		_w1605_,
		_w2646_
	);
	LUT2 #(
		.INIT('h1)
	) name2511 (
		_w2643_,
		_w2644_,
		_w2647_
	);
	LUT2 #(
		.INIT('h1)
	) name2512 (
		_w2645_,
		_w2646_,
		_w2648_
	);
	LUT2 #(
		.INIT('h8)
	) name2513 (
		_w2647_,
		_w2648_,
		_w2649_
	);
	LUT2 #(
		.INIT('h1)
	) name2514 (
		\shift[6] ,
		_w2649_,
		_w2650_
	);
	LUT2 #(
		.INIT('h2)
	) name2515 (
		_w318_,
		_w1545_,
		_w2651_
	);
	LUT2 #(
		.INIT('h2)
	) name2516 (
		_w273_,
		_w1553_,
		_w2652_
	);
	LUT2 #(
		.INIT('h2)
	) name2517 (
		_w228_,
		_w1589_,
		_w2653_
	);
	LUT2 #(
		.INIT('h2)
	) name2518 (
		_w183_,
		_w1581_,
		_w2654_
	);
	LUT2 #(
		.INIT('h1)
	) name2519 (
		_w2651_,
		_w2652_,
		_w2655_
	);
	LUT2 #(
		.INIT('h1)
	) name2520 (
		_w2653_,
		_w2654_,
		_w2656_
	);
	LUT2 #(
		.INIT('h8)
	) name2521 (
		_w2655_,
		_w2656_,
		_w2657_
	);
	LUT2 #(
		.INIT('h2)
	) name2522 (
		\shift[6] ,
		_w2657_,
		_w2658_
	);
	LUT2 #(
		.INIT('h1)
	) name2523 (
		_w2650_,
		_w2658_,
		_w2659_
	);
	LUT2 #(
		.INIT('h2)
	) name2524 (
		_w318_,
		_w1678_,
		_w2660_
	);
	LUT2 #(
		.INIT('h2)
	) name2525 (
		_w273_,
		_w1670_,
		_w2661_
	);
	LUT2 #(
		.INIT('h2)
	) name2526 (
		_w228_,
		_w1634_,
		_w2662_
	);
	LUT2 #(
		.INIT('h2)
	) name2527 (
		_w183_,
		_w1642_,
		_w2663_
	);
	LUT2 #(
		.INIT('h1)
	) name2528 (
		_w2660_,
		_w2661_,
		_w2664_
	);
	LUT2 #(
		.INIT('h1)
	) name2529 (
		_w2662_,
		_w2663_,
		_w2665_
	);
	LUT2 #(
		.INIT('h8)
	) name2530 (
		_w2664_,
		_w2665_,
		_w2666_
	);
	LUT2 #(
		.INIT('h1)
	) name2531 (
		\shift[6] ,
		_w2666_,
		_w2667_
	);
	LUT2 #(
		.INIT('h2)
	) name2532 (
		_w183_,
		_w1654_,
		_w2668_
	);
	LUT2 #(
		.INIT('h2)
	) name2533 (
		_w228_,
		_w1662_,
		_w2669_
	);
	LUT2 #(
		.INIT('h2)
	) name2534 (
		_w273_,
		_w1626_,
		_w2670_
	);
	LUT2 #(
		.INIT('h2)
	) name2535 (
		_w318_,
		_w1618_,
		_w2671_
	);
	LUT2 #(
		.INIT('h1)
	) name2536 (
		_w2668_,
		_w2669_,
		_w2672_
	);
	LUT2 #(
		.INIT('h1)
	) name2537 (
		_w2670_,
		_w2671_,
		_w2673_
	);
	LUT2 #(
		.INIT('h8)
	) name2538 (
		_w2672_,
		_w2673_,
		_w2674_
	);
	LUT2 #(
		.INIT('h2)
	) name2539 (
		\shift[6] ,
		_w2674_,
		_w2675_
	);
	LUT2 #(
		.INIT('h1)
	) name2540 (
		_w2667_,
		_w2675_,
		_w2676_
	);
	LUT2 #(
		.INIT('h2)
	) name2541 (
		_w318_,
		_w1751_,
		_w2677_
	);
	LUT2 #(
		.INIT('h2)
	) name2542 (
		_w273_,
		_w1743_,
		_w2678_
	);
	LUT2 #(
		.INIT('h2)
	) name2543 (
		_w228_,
		_w1707_,
		_w2679_
	);
	LUT2 #(
		.INIT('h2)
	) name2544 (
		_w183_,
		_w1715_,
		_w2680_
	);
	LUT2 #(
		.INIT('h1)
	) name2545 (
		_w2677_,
		_w2678_,
		_w2681_
	);
	LUT2 #(
		.INIT('h1)
	) name2546 (
		_w2679_,
		_w2680_,
		_w2682_
	);
	LUT2 #(
		.INIT('h8)
	) name2547 (
		_w2681_,
		_w2682_,
		_w2683_
	);
	LUT2 #(
		.INIT('h1)
	) name2548 (
		\shift[6] ,
		_w2683_,
		_w2684_
	);
	LUT2 #(
		.INIT('h2)
	) name2549 (
		_w183_,
		_w1727_,
		_w2685_
	);
	LUT2 #(
		.INIT('h2)
	) name2550 (
		_w228_,
		_w1735_,
		_w2686_
	);
	LUT2 #(
		.INIT('h2)
	) name2551 (
		_w273_,
		_w1699_,
		_w2687_
	);
	LUT2 #(
		.INIT('h2)
	) name2552 (
		_w318_,
		_w1691_,
		_w2688_
	);
	LUT2 #(
		.INIT('h1)
	) name2553 (
		_w2685_,
		_w2686_,
		_w2689_
	);
	LUT2 #(
		.INIT('h1)
	) name2554 (
		_w2687_,
		_w2688_,
		_w2690_
	);
	LUT2 #(
		.INIT('h8)
	) name2555 (
		_w2689_,
		_w2690_,
		_w2691_
	);
	LUT2 #(
		.INIT('h2)
	) name2556 (
		\shift[6] ,
		_w2691_,
		_w2692_
	);
	LUT2 #(
		.INIT('h1)
	) name2557 (
		_w2684_,
		_w2692_,
		_w2693_
	);
	LUT2 #(
		.INIT('h2)
	) name2558 (
		_w318_,
		_w1824_,
		_w2694_
	);
	LUT2 #(
		.INIT('h2)
	) name2559 (
		_w273_,
		_w1816_,
		_w2695_
	);
	LUT2 #(
		.INIT('h2)
	) name2560 (
		_w228_,
		_w1780_,
		_w2696_
	);
	LUT2 #(
		.INIT('h2)
	) name2561 (
		_w183_,
		_w1788_,
		_w2697_
	);
	LUT2 #(
		.INIT('h1)
	) name2562 (
		_w2694_,
		_w2695_,
		_w2698_
	);
	LUT2 #(
		.INIT('h1)
	) name2563 (
		_w2696_,
		_w2697_,
		_w2699_
	);
	LUT2 #(
		.INIT('h8)
	) name2564 (
		_w2698_,
		_w2699_,
		_w2700_
	);
	LUT2 #(
		.INIT('h1)
	) name2565 (
		\shift[6] ,
		_w2700_,
		_w2701_
	);
	LUT2 #(
		.INIT('h2)
	) name2566 (
		_w183_,
		_w1800_,
		_w2702_
	);
	LUT2 #(
		.INIT('h2)
	) name2567 (
		_w228_,
		_w1808_,
		_w2703_
	);
	LUT2 #(
		.INIT('h2)
	) name2568 (
		_w273_,
		_w1772_,
		_w2704_
	);
	LUT2 #(
		.INIT('h2)
	) name2569 (
		_w318_,
		_w1764_,
		_w2705_
	);
	LUT2 #(
		.INIT('h1)
	) name2570 (
		_w2702_,
		_w2703_,
		_w2706_
	);
	LUT2 #(
		.INIT('h1)
	) name2571 (
		_w2704_,
		_w2705_,
		_w2707_
	);
	LUT2 #(
		.INIT('h8)
	) name2572 (
		_w2706_,
		_w2707_,
		_w2708_
	);
	LUT2 #(
		.INIT('h2)
	) name2573 (
		\shift[6] ,
		_w2708_,
		_w2709_
	);
	LUT2 #(
		.INIT('h1)
	) name2574 (
		_w2701_,
		_w2709_,
		_w2710_
	);
	LUT2 #(
		.INIT('h2)
	) name2575 (
		_w183_,
		_w1861_,
		_w2711_
	);
	LUT2 #(
		.INIT('h2)
	) name2576 (
		_w228_,
		_w1853_,
		_w2712_
	);
	LUT2 #(
		.INIT('h2)
	) name2577 (
		_w273_,
		_w1889_,
		_w2713_
	);
	LUT2 #(
		.INIT('h2)
	) name2578 (
		_w318_,
		_w1897_,
		_w2714_
	);
	LUT2 #(
		.INIT('h1)
	) name2579 (
		_w2711_,
		_w2712_,
		_w2715_
	);
	LUT2 #(
		.INIT('h1)
	) name2580 (
		_w2713_,
		_w2714_,
		_w2716_
	);
	LUT2 #(
		.INIT('h8)
	) name2581 (
		_w2715_,
		_w2716_,
		_w2717_
	);
	LUT2 #(
		.INIT('h1)
	) name2582 (
		\shift[6] ,
		_w2717_,
		_w2718_
	);
	LUT2 #(
		.INIT('h2)
	) name2583 (
		_w183_,
		_w1873_,
		_w2719_
	);
	LUT2 #(
		.INIT('h2)
	) name2584 (
		_w228_,
		_w1881_,
		_w2720_
	);
	LUT2 #(
		.INIT('h2)
	) name2585 (
		_w273_,
		_w1845_,
		_w2721_
	);
	LUT2 #(
		.INIT('h2)
	) name2586 (
		_w318_,
		_w1837_,
		_w2722_
	);
	LUT2 #(
		.INIT('h1)
	) name2587 (
		_w2719_,
		_w2720_,
		_w2723_
	);
	LUT2 #(
		.INIT('h1)
	) name2588 (
		_w2721_,
		_w2722_,
		_w2724_
	);
	LUT2 #(
		.INIT('h8)
	) name2589 (
		_w2723_,
		_w2724_,
		_w2725_
	);
	LUT2 #(
		.INIT('h2)
	) name2590 (
		\shift[6] ,
		_w2725_,
		_w2726_
	);
	LUT2 #(
		.INIT('h1)
	) name2591 (
		_w2718_,
		_w2726_,
		_w2727_
	);
	LUT2 #(
		.INIT('h2)
	) name2592 (
		_w183_,
		_w1934_,
		_w2728_
	);
	LUT2 #(
		.INIT('h2)
	) name2593 (
		_w228_,
		_w1926_,
		_w2729_
	);
	LUT2 #(
		.INIT('h2)
	) name2594 (
		_w273_,
		_w1962_,
		_w2730_
	);
	LUT2 #(
		.INIT('h2)
	) name2595 (
		_w318_,
		_w1970_,
		_w2731_
	);
	LUT2 #(
		.INIT('h1)
	) name2596 (
		_w2728_,
		_w2729_,
		_w2732_
	);
	LUT2 #(
		.INIT('h1)
	) name2597 (
		_w2730_,
		_w2731_,
		_w2733_
	);
	LUT2 #(
		.INIT('h8)
	) name2598 (
		_w2732_,
		_w2733_,
		_w2734_
	);
	LUT2 #(
		.INIT('h1)
	) name2599 (
		\shift[6] ,
		_w2734_,
		_w2735_
	);
	LUT2 #(
		.INIT('h2)
	) name2600 (
		_w183_,
		_w1946_,
		_w2736_
	);
	LUT2 #(
		.INIT('h2)
	) name2601 (
		_w228_,
		_w1954_,
		_w2737_
	);
	LUT2 #(
		.INIT('h2)
	) name2602 (
		_w273_,
		_w1918_,
		_w2738_
	);
	LUT2 #(
		.INIT('h2)
	) name2603 (
		_w318_,
		_w1910_,
		_w2739_
	);
	LUT2 #(
		.INIT('h1)
	) name2604 (
		_w2736_,
		_w2737_,
		_w2740_
	);
	LUT2 #(
		.INIT('h1)
	) name2605 (
		_w2738_,
		_w2739_,
		_w2741_
	);
	LUT2 #(
		.INIT('h8)
	) name2606 (
		_w2740_,
		_w2741_,
		_w2742_
	);
	LUT2 #(
		.INIT('h2)
	) name2607 (
		\shift[6] ,
		_w2742_,
		_w2743_
	);
	LUT2 #(
		.INIT('h1)
	) name2608 (
		_w2735_,
		_w2743_,
		_w2744_
	);
	LUT2 #(
		.INIT('h2)
	) name2609 (
		_w183_,
		_w2007_,
		_w2745_
	);
	LUT2 #(
		.INIT('h2)
	) name2610 (
		_w228_,
		_w1999_,
		_w2746_
	);
	LUT2 #(
		.INIT('h2)
	) name2611 (
		_w273_,
		_w2035_,
		_w2747_
	);
	LUT2 #(
		.INIT('h2)
	) name2612 (
		_w318_,
		_w2043_,
		_w2748_
	);
	LUT2 #(
		.INIT('h1)
	) name2613 (
		_w2745_,
		_w2746_,
		_w2749_
	);
	LUT2 #(
		.INIT('h1)
	) name2614 (
		_w2747_,
		_w2748_,
		_w2750_
	);
	LUT2 #(
		.INIT('h8)
	) name2615 (
		_w2749_,
		_w2750_,
		_w2751_
	);
	LUT2 #(
		.INIT('h1)
	) name2616 (
		\shift[6] ,
		_w2751_,
		_w2752_
	);
	LUT2 #(
		.INIT('h2)
	) name2617 (
		_w183_,
		_w2019_,
		_w2753_
	);
	LUT2 #(
		.INIT('h2)
	) name2618 (
		_w228_,
		_w2027_,
		_w2754_
	);
	LUT2 #(
		.INIT('h2)
	) name2619 (
		_w273_,
		_w1991_,
		_w2755_
	);
	LUT2 #(
		.INIT('h2)
	) name2620 (
		_w318_,
		_w1983_,
		_w2756_
	);
	LUT2 #(
		.INIT('h1)
	) name2621 (
		_w2753_,
		_w2754_,
		_w2757_
	);
	LUT2 #(
		.INIT('h1)
	) name2622 (
		_w2755_,
		_w2756_,
		_w2758_
	);
	LUT2 #(
		.INIT('h8)
	) name2623 (
		_w2757_,
		_w2758_,
		_w2759_
	);
	LUT2 #(
		.INIT('h2)
	) name2624 (
		\shift[6] ,
		_w2759_,
		_w2760_
	);
	LUT2 #(
		.INIT('h1)
	) name2625 (
		_w2752_,
		_w2760_,
		_w2761_
	);
	LUT2 #(
		.INIT('h2)
	) name2626 (
		_w183_,
		_w2080_,
		_w2762_
	);
	LUT2 #(
		.INIT('h2)
	) name2627 (
		_w228_,
		_w2072_,
		_w2763_
	);
	LUT2 #(
		.INIT('h2)
	) name2628 (
		_w273_,
		_w2108_,
		_w2764_
	);
	LUT2 #(
		.INIT('h2)
	) name2629 (
		_w318_,
		_w2116_,
		_w2765_
	);
	LUT2 #(
		.INIT('h1)
	) name2630 (
		_w2762_,
		_w2763_,
		_w2766_
	);
	LUT2 #(
		.INIT('h1)
	) name2631 (
		_w2764_,
		_w2765_,
		_w2767_
	);
	LUT2 #(
		.INIT('h8)
	) name2632 (
		_w2766_,
		_w2767_,
		_w2768_
	);
	LUT2 #(
		.INIT('h1)
	) name2633 (
		\shift[6] ,
		_w2768_,
		_w2769_
	);
	LUT2 #(
		.INIT('h2)
	) name2634 (
		_w183_,
		_w2092_,
		_w2770_
	);
	LUT2 #(
		.INIT('h2)
	) name2635 (
		_w228_,
		_w2100_,
		_w2771_
	);
	LUT2 #(
		.INIT('h2)
	) name2636 (
		_w273_,
		_w2064_,
		_w2772_
	);
	LUT2 #(
		.INIT('h2)
	) name2637 (
		_w318_,
		_w2056_,
		_w2773_
	);
	LUT2 #(
		.INIT('h1)
	) name2638 (
		_w2770_,
		_w2771_,
		_w2774_
	);
	LUT2 #(
		.INIT('h1)
	) name2639 (
		_w2772_,
		_w2773_,
		_w2775_
	);
	LUT2 #(
		.INIT('h8)
	) name2640 (
		_w2774_,
		_w2775_,
		_w2776_
	);
	LUT2 #(
		.INIT('h2)
	) name2641 (
		\shift[6] ,
		_w2776_,
		_w2777_
	);
	LUT2 #(
		.INIT('h1)
	) name2642 (
		_w2769_,
		_w2777_,
		_w2778_
	);
	LUT2 #(
		.INIT('h2)
	) name2643 (
		_w183_,
		_w2153_,
		_w2779_
	);
	LUT2 #(
		.INIT('h2)
	) name2644 (
		_w228_,
		_w2145_,
		_w2780_
	);
	LUT2 #(
		.INIT('h2)
	) name2645 (
		_w273_,
		_w2181_,
		_w2781_
	);
	LUT2 #(
		.INIT('h2)
	) name2646 (
		_w318_,
		_w2189_,
		_w2782_
	);
	LUT2 #(
		.INIT('h1)
	) name2647 (
		_w2779_,
		_w2780_,
		_w2783_
	);
	LUT2 #(
		.INIT('h1)
	) name2648 (
		_w2781_,
		_w2782_,
		_w2784_
	);
	LUT2 #(
		.INIT('h8)
	) name2649 (
		_w2783_,
		_w2784_,
		_w2785_
	);
	LUT2 #(
		.INIT('h1)
	) name2650 (
		\shift[6] ,
		_w2785_,
		_w2786_
	);
	LUT2 #(
		.INIT('h2)
	) name2651 (
		_w183_,
		_w2165_,
		_w2787_
	);
	LUT2 #(
		.INIT('h2)
	) name2652 (
		_w228_,
		_w2173_,
		_w2788_
	);
	LUT2 #(
		.INIT('h2)
	) name2653 (
		_w273_,
		_w2137_,
		_w2789_
	);
	LUT2 #(
		.INIT('h2)
	) name2654 (
		_w318_,
		_w2129_,
		_w2790_
	);
	LUT2 #(
		.INIT('h1)
	) name2655 (
		_w2787_,
		_w2788_,
		_w2791_
	);
	LUT2 #(
		.INIT('h1)
	) name2656 (
		_w2789_,
		_w2790_,
		_w2792_
	);
	LUT2 #(
		.INIT('h8)
	) name2657 (
		_w2791_,
		_w2792_,
		_w2793_
	);
	LUT2 #(
		.INIT('h2)
	) name2658 (
		\shift[6] ,
		_w2793_,
		_w2794_
	);
	LUT2 #(
		.INIT('h1)
	) name2659 (
		_w2786_,
		_w2794_,
		_w2795_
	);
	LUT2 #(
		.INIT('h2)
	) name2660 (
		_w183_,
		_w2226_,
		_w2796_
	);
	LUT2 #(
		.INIT('h2)
	) name2661 (
		_w228_,
		_w2218_,
		_w2797_
	);
	LUT2 #(
		.INIT('h2)
	) name2662 (
		_w273_,
		_w2254_,
		_w2798_
	);
	LUT2 #(
		.INIT('h2)
	) name2663 (
		_w318_,
		_w2262_,
		_w2799_
	);
	LUT2 #(
		.INIT('h1)
	) name2664 (
		_w2796_,
		_w2797_,
		_w2800_
	);
	LUT2 #(
		.INIT('h1)
	) name2665 (
		_w2798_,
		_w2799_,
		_w2801_
	);
	LUT2 #(
		.INIT('h8)
	) name2666 (
		_w2800_,
		_w2801_,
		_w2802_
	);
	LUT2 #(
		.INIT('h1)
	) name2667 (
		\shift[6] ,
		_w2802_,
		_w2803_
	);
	LUT2 #(
		.INIT('h2)
	) name2668 (
		_w183_,
		_w2238_,
		_w2804_
	);
	LUT2 #(
		.INIT('h2)
	) name2669 (
		_w228_,
		_w2246_,
		_w2805_
	);
	LUT2 #(
		.INIT('h2)
	) name2670 (
		_w273_,
		_w2210_,
		_w2806_
	);
	LUT2 #(
		.INIT('h2)
	) name2671 (
		_w318_,
		_w2202_,
		_w2807_
	);
	LUT2 #(
		.INIT('h1)
	) name2672 (
		_w2804_,
		_w2805_,
		_w2808_
	);
	LUT2 #(
		.INIT('h1)
	) name2673 (
		_w2806_,
		_w2807_,
		_w2809_
	);
	LUT2 #(
		.INIT('h8)
	) name2674 (
		_w2808_,
		_w2809_,
		_w2810_
	);
	LUT2 #(
		.INIT('h2)
	) name2675 (
		\shift[6] ,
		_w2810_,
		_w2811_
	);
	LUT2 #(
		.INIT('h1)
	) name2676 (
		_w2803_,
		_w2811_,
		_w2812_
	);
	LUT2 #(
		.INIT('h2)
	) name2677 (
		_w183_,
		_w272_,
		_w2813_
	);
	LUT2 #(
		.INIT('h2)
	) name2678 (
		_w228_,
		_w366_,
		_w2814_
	);
	LUT2 #(
		.INIT('h2)
	) name2679 (
		_w273_,
		_w500_,
		_w2815_
	);
	LUT2 #(
		.INIT('h2)
	) name2680 (
		_w318_,
		_w410_,
		_w2816_
	);
	LUT2 #(
		.INIT('h1)
	) name2681 (
		_w2813_,
		_w2814_,
		_w2817_
	);
	LUT2 #(
		.INIT('h1)
	) name2682 (
		_w2815_,
		_w2816_,
		_w2818_
	);
	LUT2 #(
		.INIT('h8)
	) name2683 (
		_w2817_,
		_w2818_,
		_w2819_
	);
	LUT2 #(
		.INIT('h1)
	) name2684 (
		\shift[6] ,
		_w2819_,
		_w2820_
	);
	LUT2 #(
		.INIT('h4)
	) name2685 (
		_w182_,
		_w228_,
		_w2821_
	);
	LUT2 #(
		.INIT('h4)
	) name2686 (
		_w227_,
		_w318_,
		_w2822_
	);
	LUT2 #(
		.INIT('h2)
	) name2687 (
		_w183_,
		_w454_,
		_w2823_
	);
	LUT2 #(
		.INIT('h2)
	) name2688 (
		_w273_,
		_w317_,
		_w2824_
	);
	LUT2 #(
		.INIT('h1)
	) name2689 (
		_w2821_,
		_w2822_,
		_w2825_
	);
	LUT2 #(
		.INIT('h1)
	) name2690 (
		_w2823_,
		_w2824_,
		_w2826_
	);
	LUT2 #(
		.INIT('h8)
	) name2691 (
		_w2825_,
		_w2826_,
		_w2827_
	);
	LUT2 #(
		.INIT('h2)
	) name2692 (
		\shift[6] ,
		_w2827_,
		_w2828_
	);
	LUT2 #(
		.INIT('h1)
	) name2693 (
		_w2820_,
		_w2828_,
		_w2829_
	);
	LUT2 #(
		.INIT('h2)
	) name2694 (
		_w183_,
		_w661_,
		_w2830_
	);
	LUT2 #(
		.INIT('h2)
	) name2695 (
		_w228_,
		_w821_,
		_w2831_
	);
	LUT2 #(
		.INIT('h2)
	) name2696 (
		_w273_,
		_w869_,
		_w2832_
	);
	LUT2 #(
		.INIT('h2)
	) name2697 (
		_w318_,
		_w921_,
		_w2833_
	);
	LUT2 #(
		.INIT('h1)
	) name2698 (
		_w2830_,
		_w2831_,
		_w2834_
	);
	LUT2 #(
		.INIT('h1)
	) name2699 (
		_w2832_,
		_w2833_,
		_w2835_
	);
	LUT2 #(
		.INIT('h8)
	) name2700 (
		_w2834_,
		_w2835_,
		_w2836_
	);
	LUT2 #(
		.INIT('h1)
	) name2701 (
		\shift[6] ,
		_w2836_,
		_w2837_
	);
	LUT2 #(
		.INIT('h2)
	) name2702 (
		_w183_,
		_w769_,
		_w2838_
	);
	LUT2 #(
		.INIT('h2)
	) name2703 (
		_w228_,
		_w557_,
		_w2839_
	);
	LUT2 #(
		.INIT('h2)
	) name2704 (
		_w273_,
		_w713_,
		_w2840_
	);
	LUT2 #(
		.INIT('h2)
	) name2705 (
		_w318_,
		_w609_,
		_w2841_
	);
	LUT2 #(
		.INIT('h1)
	) name2706 (
		_w2838_,
		_w2839_,
		_w2842_
	);
	LUT2 #(
		.INIT('h1)
	) name2707 (
		_w2840_,
		_w2841_,
		_w2843_
	);
	LUT2 #(
		.INIT('h8)
	) name2708 (
		_w2842_,
		_w2843_,
		_w2844_
	);
	LUT2 #(
		.INIT('h2)
	) name2709 (
		\shift[6] ,
		_w2844_,
		_w2845_
	);
	LUT2 #(
		.INIT('h1)
	) name2710 (
		_w2837_,
		_w2845_,
		_w2846_
	);
	LUT2 #(
		.INIT('h2)
	) name2711 (
		_w183_,
		_w986_,
		_w2847_
	);
	LUT2 #(
		.INIT('h2)
	) name2712 (
		_w228_,
		_w1050_,
		_w2848_
	);
	LUT2 #(
		.INIT('h2)
	) name2713 (
		_w273_,
		_w1072_,
		_w2849_
	);
	LUT2 #(
		.INIT('h2)
	) name2714 (
		_w318_,
		_w1092_,
		_w2850_
	);
	LUT2 #(
		.INIT('h1)
	) name2715 (
		_w2847_,
		_w2848_,
		_w2851_
	);
	LUT2 #(
		.INIT('h1)
	) name2716 (
		_w2849_,
		_w2850_,
		_w2852_
	);
	LUT2 #(
		.INIT('h8)
	) name2717 (
		_w2851_,
		_w2852_,
		_w2853_
	);
	LUT2 #(
		.INIT('h1)
	) name2718 (
		\shift[6] ,
		_w2853_,
		_w2854_
	);
	LUT2 #(
		.INIT('h2)
	) name2719 (
		_w183_,
		_w1030_,
		_w2855_
	);
	LUT2 #(
		.INIT('h2)
	) name2720 (
		_w228_,
		_w946_,
		_w2856_
	);
	LUT2 #(
		.INIT('h2)
	) name2721 (
		_w273_,
		_w1006_,
		_w2857_
	);
	LUT2 #(
		.INIT('h2)
	) name2722 (
		_w318_,
		_w966_,
		_w2858_
	);
	LUT2 #(
		.INIT('h1)
	) name2723 (
		_w2855_,
		_w2856_,
		_w2859_
	);
	LUT2 #(
		.INIT('h1)
	) name2724 (
		_w2857_,
		_w2858_,
		_w2860_
	);
	LUT2 #(
		.INIT('h8)
	) name2725 (
		_w2859_,
		_w2860_,
		_w2861_
	);
	LUT2 #(
		.INIT('h2)
	) name2726 (
		\shift[6] ,
		_w2861_,
		_w2862_
	);
	LUT2 #(
		.INIT('h1)
	) name2727 (
		_w2854_,
		_w2862_,
		_w2863_
	);
	LUT2 #(
		.INIT('h2)
	) name2728 (
		_w273_,
		_w1314_,
		_w2864_
	);
	LUT2 #(
		.INIT('h2)
	) name2729 (
		_w318_,
		_w1386_,
		_w2865_
	);
	LUT2 #(
		.INIT('h2)
	) name2730 (
		_w183_,
		_w1205_,
		_w2866_
	);
	LUT2 #(
		.INIT('h2)
	) name2731 (
		_w228_,
		_w1350_,
		_w2867_
	);
	LUT2 #(
		.INIT('h1)
	) name2732 (
		_w2864_,
		_w2865_,
		_w2868_
	);
	LUT2 #(
		.INIT('h1)
	) name2733 (
		_w2866_,
		_w2867_,
		_w2869_
	);
	LUT2 #(
		.INIT('h8)
	) name2734 (
		_w2868_,
		_w2869_,
		_w2870_
	);
	LUT2 #(
		.INIT('h1)
	) name2735 (
		\shift[6] ,
		_w2870_,
		_w2871_
	);
	LUT2 #(
		.INIT('h2)
	) name2736 (
		_w183_,
		_w1281_,
		_w2872_
	);
	LUT2 #(
		.INIT('h2)
	) name2737 (
		_w273_,
		_w1133_,
		_w2873_
	);
	LUT2 #(
		.INIT('h2)
	) name2738 (
		_w228_,
		_w1241_,
		_w2874_
	);
	LUT2 #(
		.INIT('h2)
	) name2739 (
		_w318_,
		_w1169_,
		_w2875_
	);
	LUT2 #(
		.INIT('h1)
	) name2740 (
		_w2872_,
		_w2873_,
		_w2876_
	);
	LUT2 #(
		.INIT('h1)
	) name2741 (
		_w2874_,
		_w2875_,
		_w2877_
	);
	LUT2 #(
		.INIT('h8)
	) name2742 (
		_w2876_,
		_w2877_,
		_w2878_
	);
	LUT2 #(
		.INIT('h2)
	) name2743 (
		\shift[6] ,
		_w2878_,
		_w2879_
	);
	LUT2 #(
		.INIT('h1)
	) name2744 (
		_w2871_,
		_w2879_,
		_w2880_
	);
	LUT2 #(
		.INIT('h2)
	) name2745 (
		_w273_,
		_w1435_,
		_w2881_
	);
	LUT2 #(
		.INIT('h2)
	) name2746 (
		_w183_,
		_w1415_,
		_w2882_
	);
	LUT2 #(
		.INIT('h2)
	) name2747 (
		_w318_,
		_w1451_,
		_w2883_
	);
	LUT2 #(
		.INIT('h2)
	) name2748 (
		_w228_,
		_w1459_,
		_w2884_
	);
	LUT2 #(
		.INIT('h1)
	) name2749 (
		_w2881_,
		_w2882_,
		_w2885_
	);
	LUT2 #(
		.INIT('h1)
	) name2750 (
		_w2883_,
		_w2884_,
		_w2886_
	);
	LUT2 #(
		.INIT('h8)
	) name2751 (
		_w2885_,
		_w2886_,
		_w2887_
	);
	LUT2 #(
		.INIT('h1)
	) name2752 (
		\shift[6] ,
		_w2887_,
		_w2888_
	);
	LUT2 #(
		.INIT('h2)
	) name2753 (
		_w228_,
		_w1399_,
		_w2889_
	);
	LUT2 #(
		.INIT('h2)
	) name2754 (
		_w318_,
		_w1407_,
		_w2890_
	);
	LUT2 #(
		.INIT('h2)
	) name2755 (
		_w273_,
		_w1423_,
		_w2891_
	);
	LUT2 #(
		.INIT('h2)
	) name2756 (
		_w183_,
		_w1443_,
		_w2892_
	);
	LUT2 #(
		.INIT('h1)
	) name2757 (
		_w2889_,
		_w2890_,
		_w2893_
	);
	LUT2 #(
		.INIT('h1)
	) name2758 (
		_w2891_,
		_w2892_,
		_w2894_
	);
	LUT2 #(
		.INIT('h8)
	) name2759 (
		_w2893_,
		_w2894_,
		_w2895_
	);
	LUT2 #(
		.INIT('h2)
	) name2760 (
		\shift[6] ,
		_w2895_,
		_w2896_
	);
	LUT2 #(
		.INIT('h1)
	) name2761 (
		_w2888_,
		_w2896_,
		_w2897_
	);
	LUT2 #(
		.INIT('h2)
	) name2762 (
		_w273_,
		_w1508_,
		_w2898_
	);
	LUT2 #(
		.INIT('h2)
	) name2763 (
		_w183_,
		_w1488_,
		_w2899_
	);
	LUT2 #(
		.INIT('h2)
	) name2764 (
		_w318_,
		_w1524_,
		_w2900_
	);
	LUT2 #(
		.INIT('h2)
	) name2765 (
		_w228_,
		_w1532_,
		_w2901_
	);
	LUT2 #(
		.INIT('h1)
	) name2766 (
		_w2898_,
		_w2899_,
		_w2902_
	);
	LUT2 #(
		.INIT('h1)
	) name2767 (
		_w2900_,
		_w2901_,
		_w2903_
	);
	LUT2 #(
		.INIT('h8)
	) name2768 (
		_w2902_,
		_w2903_,
		_w2904_
	);
	LUT2 #(
		.INIT('h1)
	) name2769 (
		\shift[6] ,
		_w2904_,
		_w2905_
	);
	LUT2 #(
		.INIT('h2)
	) name2770 (
		_w228_,
		_w1472_,
		_w2906_
	);
	LUT2 #(
		.INIT('h2)
	) name2771 (
		_w318_,
		_w1480_,
		_w2907_
	);
	LUT2 #(
		.INIT('h2)
	) name2772 (
		_w273_,
		_w1496_,
		_w2908_
	);
	LUT2 #(
		.INIT('h2)
	) name2773 (
		_w183_,
		_w1516_,
		_w2909_
	);
	LUT2 #(
		.INIT('h1)
	) name2774 (
		_w2906_,
		_w2907_,
		_w2910_
	);
	LUT2 #(
		.INIT('h1)
	) name2775 (
		_w2908_,
		_w2909_,
		_w2911_
	);
	LUT2 #(
		.INIT('h8)
	) name2776 (
		_w2910_,
		_w2911_,
		_w2912_
	);
	LUT2 #(
		.INIT('h2)
	) name2777 (
		\shift[6] ,
		_w2912_,
		_w2913_
	);
	LUT2 #(
		.INIT('h1)
	) name2778 (
		_w2905_,
		_w2913_,
		_w2914_
	);
	LUT2 #(
		.INIT('h2)
	) name2779 (
		_w273_,
		_w1581_,
		_w2915_
	);
	LUT2 #(
		.INIT('h2)
	) name2780 (
		_w183_,
		_w1561_,
		_w2916_
	);
	LUT2 #(
		.INIT('h2)
	) name2781 (
		_w318_,
		_w1597_,
		_w2917_
	);
	LUT2 #(
		.INIT('h2)
	) name2782 (
		_w228_,
		_w1605_,
		_w2918_
	);
	LUT2 #(
		.INIT('h1)
	) name2783 (
		_w2915_,
		_w2916_,
		_w2919_
	);
	LUT2 #(
		.INIT('h1)
	) name2784 (
		_w2917_,
		_w2918_,
		_w2920_
	);
	LUT2 #(
		.INIT('h8)
	) name2785 (
		_w2919_,
		_w2920_,
		_w2921_
	);
	LUT2 #(
		.INIT('h1)
	) name2786 (
		\shift[6] ,
		_w2921_,
		_w2922_
	);
	LUT2 #(
		.INIT('h2)
	) name2787 (
		_w228_,
		_w1545_,
		_w2923_
	);
	LUT2 #(
		.INIT('h2)
	) name2788 (
		_w318_,
		_w1553_,
		_w2924_
	);
	LUT2 #(
		.INIT('h2)
	) name2789 (
		_w273_,
		_w1569_,
		_w2925_
	);
	LUT2 #(
		.INIT('h2)
	) name2790 (
		_w183_,
		_w1589_,
		_w2926_
	);
	LUT2 #(
		.INIT('h1)
	) name2791 (
		_w2923_,
		_w2924_,
		_w2927_
	);
	LUT2 #(
		.INIT('h1)
	) name2792 (
		_w2925_,
		_w2926_,
		_w2928_
	);
	LUT2 #(
		.INIT('h8)
	) name2793 (
		_w2927_,
		_w2928_,
		_w2929_
	);
	LUT2 #(
		.INIT('h2)
	) name2794 (
		\shift[6] ,
		_w2929_,
		_w2930_
	);
	LUT2 #(
		.INIT('h1)
	) name2795 (
		_w2922_,
		_w2930_,
		_w2931_
	);
	LUT2 #(
		.INIT('h2)
	) name2796 (
		_w273_,
		_w1654_,
		_w2932_
	);
	LUT2 #(
		.INIT('h2)
	) name2797 (
		_w228_,
		_w1678_,
		_w2933_
	);
	LUT2 #(
		.INIT('h2)
	) name2798 (
		_w183_,
		_w1634_,
		_w2934_
	);
	LUT2 #(
		.INIT('h2)
	) name2799 (
		_w318_,
		_w1670_,
		_w2935_
	);
	LUT2 #(
		.INIT('h1)
	) name2800 (
		_w2932_,
		_w2933_,
		_w2936_
	);
	LUT2 #(
		.INIT('h1)
	) name2801 (
		_w2934_,
		_w2935_,
		_w2937_
	);
	LUT2 #(
		.INIT('h8)
	) name2802 (
		_w2936_,
		_w2937_,
		_w2938_
	);
	LUT2 #(
		.INIT('h1)
	) name2803 (
		\shift[6] ,
		_w2938_,
		_w2939_
	);
	LUT2 #(
		.INIT('h2)
	) name2804 (
		_w183_,
		_w1662_,
		_w2940_
	);
	LUT2 #(
		.INIT('h2)
	) name2805 (
		_w228_,
		_w1618_,
		_w2941_
	);
	LUT2 #(
		.INIT('h2)
	) name2806 (
		_w273_,
		_w1642_,
		_w2942_
	);
	LUT2 #(
		.INIT('h2)
	) name2807 (
		_w318_,
		_w1626_,
		_w2943_
	);
	LUT2 #(
		.INIT('h1)
	) name2808 (
		_w2940_,
		_w2941_,
		_w2944_
	);
	LUT2 #(
		.INIT('h1)
	) name2809 (
		_w2942_,
		_w2943_,
		_w2945_
	);
	LUT2 #(
		.INIT('h8)
	) name2810 (
		_w2944_,
		_w2945_,
		_w2946_
	);
	LUT2 #(
		.INIT('h2)
	) name2811 (
		\shift[6] ,
		_w2946_,
		_w2947_
	);
	LUT2 #(
		.INIT('h1)
	) name2812 (
		_w2939_,
		_w2947_,
		_w2948_
	);
	LUT2 #(
		.INIT('h2)
	) name2813 (
		_w273_,
		_w1727_,
		_w2949_
	);
	LUT2 #(
		.INIT('h2)
	) name2814 (
		_w228_,
		_w1751_,
		_w2950_
	);
	LUT2 #(
		.INIT('h2)
	) name2815 (
		_w183_,
		_w1707_,
		_w2951_
	);
	LUT2 #(
		.INIT('h2)
	) name2816 (
		_w318_,
		_w1743_,
		_w2952_
	);
	LUT2 #(
		.INIT('h1)
	) name2817 (
		_w2949_,
		_w2950_,
		_w2953_
	);
	LUT2 #(
		.INIT('h1)
	) name2818 (
		_w2951_,
		_w2952_,
		_w2954_
	);
	LUT2 #(
		.INIT('h8)
	) name2819 (
		_w2953_,
		_w2954_,
		_w2955_
	);
	LUT2 #(
		.INIT('h1)
	) name2820 (
		\shift[6] ,
		_w2955_,
		_w2956_
	);
	LUT2 #(
		.INIT('h2)
	) name2821 (
		_w183_,
		_w1735_,
		_w2957_
	);
	LUT2 #(
		.INIT('h2)
	) name2822 (
		_w228_,
		_w1691_,
		_w2958_
	);
	LUT2 #(
		.INIT('h2)
	) name2823 (
		_w273_,
		_w1715_,
		_w2959_
	);
	LUT2 #(
		.INIT('h2)
	) name2824 (
		_w318_,
		_w1699_,
		_w2960_
	);
	LUT2 #(
		.INIT('h1)
	) name2825 (
		_w2957_,
		_w2958_,
		_w2961_
	);
	LUT2 #(
		.INIT('h1)
	) name2826 (
		_w2959_,
		_w2960_,
		_w2962_
	);
	LUT2 #(
		.INIT('h8)
	) name2827 (
		_w2961_,
		_w2962_,
		_w2963_
	);
	LUT2 #(
		.INIT('h2)
	) name2828 (
		\shift[6] ,
		_w2963_,
		_w2964_
	);
	LUT2 #(
		.INIT('h1)
	) name2829 (
		_w2956_,
		_w2964_,
		_w2965_
	);
	LUT2 #(
		.INIT('h2)
	) name2830 (
		_w273_,
		_w1800_,
		_w2966_
	);
	LUT2 #(
		.INIT('h2)
	) name2831 (
		_w228_,
		_w1824_,
		_w2967_
	);
	LUT2 #(
		.INIT('h2)
	) name2832 (
		_w183_,
		_w1780_,
		_w2968_
	);
	LUT2 #(
		.INIT('h2)
	) name2833 (
		_w318_,
		_w1816_,
		_w2969_
	);
	LUT2 #(
		.INIT('h1)
	) name2834 (
		_w2966_,
		_w2967_,
		_w2970_
	);
	LUT2 #(
		.INIT('h1)
	) name2835 (
		_w2968_,
		_w2969_,
		_w2971_
	);
	LUT2 #(
		.INIT('h8)
	) name2836 (
		_w2970_,
		_w2971_,
		_w2972_
	);
	LUT2 #(
		.INIT('h1)
	) name2837 (
		\shift[6] ,
		_w2972_,
		_w2973_
	);
	LUT2 #(
		.INIT('h2)
	) name2838 (
		_w183_,
		_w1808_,
		_w2974_
	);
	LUT2 #(
		.INIT('h2)
	) name2839 (
		_w228_,
		_w1764_,
		_w2975_
	);
	LUT2 #(
		.INIT('h2)
	) name2840 (
		_w273_,
		_w1788_,
		_w2976_
	);
	LUT2 #(
		.INIT('h2)
	) name2841 (
		_w318_,
		_w1772_,
		_w2977_
	);
	LUT2 #(
		.INIT('h1)
	) name2842 (
		_w2974_,
		_w2975_,
		_w2978_
	);
	LUT2 #(
		.INIT('h1)
	) name2843 (
		_w2976_,
		_w2977_,
		_w2979_
	);
	LUT2 #(
		.INIT('h8)
	) name2844 (
		_w2978_,
		_w2979_,
		_w2980_
	);
	LUT2 #(
		.INIT('h2)
	) name2845 (
		\shift[6] ,
		_w2980_,
		_w2981_
	);
	LUT2 #(
		.INIT('h1)
	) name2846 (
		_w2973_,
		_w2981_,
		_w2982_
	);
	LUT2 #(
		.INIT('h2)
	) name2847 (
		_w273_,
		_w1873_,
		_w2983_
	);
	LUT2 #(
		.INIT('h2)
	) name2848 (
		_w183_,
		_w1853_,
		_w2984_
	);
	LUT2 #(
		.INIT('h2)
	) name2849 (
		_w318_,
		_w1889_,
		_w2985_
	);
	LUT2 #(
		.INIT('h2)
	) name2850 (
		_w228_,
		_w1897_,
		_w2986_
	);
	LUT2 #(
		.INIT('h1)
	) name2851 (
		_w2983_,
		_w2984_,
		_w2987_
	);
	LUT2 #(
		.INIT('h1)
	) name2852 (
		_w2985_,
		_w2986_,
		_w2988_
	);
	LUT2 #(
		.INIT('h8)
	) name2853 (
		_w2987_,
		_w2988_,
		_w2989_
	);
	LUT2 #(
		.INIT('h1)
	) name2854 (
		\shift[6] ,
		_w2989_,
		_w2990_
	);
	LUT2 #(
		.INIT('h2)
	) name2855 (
		_w183_,
		_w1881_,
		_w2991_
	);
	LUT2 #(
		.INIT('h2)
	) name2856 (
		_w228_,
		_w1837_,
		_w2992_
	);
	LUT2 #(
		.INIT('h2)
	) name2857 (
		_w273_,
		_w1861_,
		_w2993_
	);
	LUT2 #(
		.INIT('h2)
	) name2858 (
		_w318_,
		_w1845_,
		_w2994_
	);
	LUT2 #(
		.INIT('h1)
	) name2859 (
		_w2991_,
		_w2992_,
		_w2995_
	);
	LUT2 #(
		.INIT('h1)
	) name2860 (
		_w2993_,
		_w2994_,
		_w2996_
	);
	LUT2 #(
		.INIT('h8)
	) name2861 (
		_w2995_,
		_w2996_,
		_w2997_
	);
	LUT2 #(
		.INIT('h2)
	) name2862 (
		\shift[6] ,
		_w2997_,
		_w2998_
	);
	LUT2 #(
		.INIT('h1)
	) name2863 (
		_w2990_,
		_w2998_,
		_w2999_
	);
	LUT2 #(
		.INIT('h2)
	) name2864 (
		_w273_,
		_w1946_,
		_w3000_
	);
	LUT2 #(
		.INIT('h2)
	) name2865 (
		_w183_,
		_w1926_,
		_w3001_
	);
	LUT2 #(
		.INIT('h2)
	) name2866 (
		_w318_,
		_w1962_,
		_w3002_
	);
	LUT2 #(
		.INIT('h2)
	) name2867 (
		_w228_,
		_w1970_,
		_w3003_
	);
	LUT2 #(
		.INIT('h1)
	) name2868 (
		_w3000_,
		_w3001_,
		_w3004_
	);
	LUT2 #(
		.INIT('h1)
	) name2869 (
		_w3002_,
		_w3003_,
		_w3005_
	);
	LUT2 #(
		.INIT('h8)
	) name2870 (
		_w3004_,
		_w3005_,
		_w3006_
	);
	LUT2 #(
		.INIT('h1)
	) name2871 (
		\shift[6] ,
		_w3006_,
		_w3007_
	);
	LUT2 #(
		.INIT('h2)
	) name2872 (
		_w183_,
		_w1954_,
		_w3008_
	);
	LUT2 #(
		.INIT('h2)
	) name2873 (
		_w228_,
		_w1910_,
		_w3009_
	);
	LUT2 #(
		.INIT('h2)
	) name2874 (
		_w273_,
		_w1934_,
		_w3010_
	);
	LUT2 #(
		.INIT('h2)
	) name2875 (
		_w318_,
		_w1918_,
		_w3011_
	);
	LUT2 #(
		.INIT('h1)
	) name2876 (
		_w3008_,
		_w3009_,
		_w3012_
	);
	LUT2 #(
		.INIT('h1)
	) name2877 (
		_w3010_,
		_w3011_,
		_w3013_
	);
	LUT2 #(
		.INIT('h8)
	) name2878 (
		_w3012_,
		_w3013_,
		_w3014_
	);
	LUT2 #(
		.INIT('h2)
	) name2879 (
		\shift[6] ,
		_w3014_,
		_w3015_
	);
	LUT2 #(
		.INIT('h1)
	) name2880 (
		_w3007_,
		_w3015_,
		_w3016_
	);
	LUT2 #(
		.INIT('h2)
	) name2881 (
		_w273_,
		_w2019_,
		_w3017_
	);
	LUT2 #(
		.INIT('h2)
	) name2882 (
		_w183_,
		_w1999_,
		_w3018_
	);
	LUT2 #(
		.INIT('h2)
	) name2883 (
		_w318_,
		_w2035_,
		_w3019_
	);
	LUT2 #(
		.INIT('h2)
	) name2884 (
		_w228_,
		_w2043_,
		_w3020_
	);
	LUT2 #(
		.INIT('h1)
	) name2885 (
		_w3017_,
		_w3018_,
		_w3021_
	);
	LUT2 #(
		.INIT('h1)
	) name2886 (
		_w3019_,
		_w3020_,
		_w3022_
	);
	LUT2 #(
		.INIT('h8)
	) name2887 (
		_w3021_,
		_w3022_,
		_w3023_
	);
	LUT2 #(
		.INIT('h1)
	) name2888 (
		\shift[6] ,
		_w3023_,
		_w3024_
	);
	LUT2 #(
		.INIT('h2)
	) name2889 (
		_w183_,
		_w2027_,
		_w3025_
	);
	LUT2 #(
		.INIT('h2)
	) name2890 (
		_w228_,
		_w1983_,
		_w3026_
	);
	LUT2 #(
		.INIT('h2)
	) name2891 (
		_w273_,
		_w2007_,
		_w3027_
	);
	LUT2 #(
		.INIT('h2)
	) name2892 (
		_w318_,
		_w1991_,
		_w3028_
	);
	LUT2 #(
		.INIT('h1)
	) name2893 (
		_w3025_,
		_w3026_,
		_w3029_
	);
	LUT2 #(
		.INIT('h1)
	) name2894 (
		_w3027_,
		_w3028_,
		_w3030_
	);
	LUT2 #(
		.INIT('h8)
	) name2895 (
		_w3029_,
		_w3030_,
		_w3031_
	);
	LUT2 #(
		.INIT('h2)
	) name2896 (
		\shift[6] ,
		_w3031_,
		_w3032_
	);
	LUT2 #(
		.INIT('h1)
	) name2897 (
		_w3024_,
		_w3032_,
		_w3033_
	);
	LUT2 #(
		.INIT('h2)
	) name2898 (
		_w273_,
		_w2092_,
		_w3034_
	);
	LUT2 #(
		.INIT('h2)
	) name2899 (
		_w183_,
		_w2072_,
		_w3035_
	);
	LUT2 #(
		.INIT('h2)
	) name2900 (
		_w318_,
		_w2108_,
		_w3036_
	);
	LUT2 #(
		.INIT('h2)
	) name2901 (
		_w228_,
		_w2116_,
		_w3037_
	);
	LUT2 #(
		.INIT('h1)
	) name2902 (
		_w3034_,
		_w3035_,
		_w3038_
	);
	LUT2 #(
		.INIT('h1)
	) name2903 (
		_w3036_,
		_w3037_,
		_w3039_
	);
	LUT2 #(
		.INIT('h8)
	) name2904 (
		_w3038_,
		_w3039_,
		_w3040_
	);
	LUT2 #(
		.INIT('h1)
	) name2905 (
		\shift[6] ,
		_w3040_,
		_w3041_
	);
	LUT2 #(
		.INIT('h2)
	) name2906 (
		_w183_,
		_w2100_,
		_w3042_
	);
	LUT2 #(
		.INIT('h2)
	) name2907 (
		_w228_,
		_w2056_,
		_w3043_
	);
	LUT2 #(
		.INIT('h2)
	) name2908 (
		_w273_,
		_w2080_,
		_w3044_
	);
	LUT2 #(
		.INIT('h2)
	) name2909 (
		_w318_,
		_w2064_,
		_w3045_
	);
	LUT2 #(
		.INIT('h1)
	) name2910 (
		_w3042_,
		_w3043_,
		_w3046_
	);
	LUT2 #(
		.INIT('h1)
	) name2911 (
		_w3044_,
		_w3045_,
		_w3047_
	);
	LUT2 #(
		.INIT('h8)
	) name2912 (
		_w3046_,
		_w3047_,
		_w3048_
	);
	LUT2 #(
		.INIT('h2)
	) name2913 (
		\shift[6] ,
		_w3048_,
		_w3049_
	);
	LUT2 #(
		.INIT('h1)
	) name2914 (
		_w3041_,
		_w3049_,
		_w3050_
	);
	LUT2 #(
		.INIT('h2)
	) name2915 (
		_w273_,
		_w2165_,
		_w3051_
	);
	LUT2 #(
		.INIT('h2)
	) name2916 (
		_w183_,
		_w2145_,
		_w3052_
	);
	LUT2 #(
		.INIT('h2)
	) name2917 (
		_w318_,
		_w2181_,
		_w3053_
	);
	LUT2 #(
		.INIT('h2)
	) name2918 (
		_w228_,
		_w2189_,
		_w3054_
	);
	LUT2 #(
		.INIT('h1)
	) name2919 (
		_w3051_,
		_w3052_,
		_w3055_
	);
	LUT2 #(
		.INIT('h1)
	) name2920 (
		_w3053_,
		_w3054_,
		_w3056_
	);
	LUT2 #(
		.INIT('h8)
	) name2921 (
		_w3055_,
		_w3056_,
		_w3057_
	);
	LUT2 #(
		.INIT('h1)
	) name2922 (
		\shift[6] ,
		_w3057_,
		_w3058_
	);
	LUT2 #(
		.INIT('h2)
	) name2923 (
		_w183_,
		_w2173_,
		_w3059_
	);
	LUT2 #(
		.INIT('h2)
	) name2924 (
		_w228_,
		_w2129_,
		_w3060_
	);
	LUT2 #(
		.INIT('h2)
	) name2925 (
		_w273_,
		_w2153_,
		_w3061_
	);
	LUT2 #(
		.INIT('h2)
	) name2926 (
		_w318_,
		_w2137_,
		_w3062_
	);
	LUT2 #(
		.INIT('h1)
	) name2927 (
		_w3059_,
		_w3060_,
		_w3063_
	);
	LUT2 #(
		.INIT('h1)
	) name2928 (
		_w3061_,
		_w3062_,
		_w3064_
	);
	LUT2 #(
		.INIT('h8)
	) name2929 (
		_w3063_,
		_w3064_,
		_w3065_
	);
	LUT2 #(
		.INIT('h2)
	) name2930 (
		\shift[6] ,
		_w3065_,
		_w3066_
	);
	LUT2 #(
		.INIT('h1)
	) name2931 (
		_w3058_,
		_w3066_,
		_w3067_
	);
	LUT2 #(
		.INIT('h2)
	) name2932 (
		_w273_,
		_w2238_,
		_w3068_
	);
	LUT2 #(
		.INIT('h2)
	) name2933 (
		_w183_,
		_w2218_,
		_w3069_
	);
	LUT2 #(
		.INIT('h2)
	) name2934 (
		_w318_,
		_w2254_,
		_w3070_
	);
	LUT2 #(
		.INIT('h2)
	) name2935 (
		_w228_,
		_w2262_,
		_w3071_
	);
	LUT2 #(
		.INIT('h1)
	) name2936 (
		_w3068_,
		_w3069_,
		_w3072_
	);
	LUT2 #(
		.INIT('h1)
	) name2937 (
		_w3070_,
		_w3071_,
		_w3073_
	);
	LUT2 #(
		.INIT('h8)
	) name2938 (
		_w3072_,
		_w3073_,
		_w3074_
	);
	LUT2 #(
		.INIT('h1)
	) name2939 (
		\shift[6] ,
		_w3074_,
		_w3075_
	);
	LUT2 #(
		.INIT('h2)
	) name2940 (
		_w183_,
		_w2246_,
		_w3076_
	);
	LUT2 #(
		.INIT('h2)
	) name2941 (
		_w228_,
		_w2202_,
		_w3077_
	);
	LUT2 #(
		.INIT('h2)
	) name2942 (
		_w273_,
		_w2226_,
		_w3078_
	);
	LUT2 #(
		.INIT('h2)
	) name2943 (
		_w318_,
		_w2210_,
		_w3079_
	);
	LUT2 #(
		.INIT('h1)
	) name2944 (
		_w3076_,
		_w3077_,
		_w3080_
	);
	LUT2 #(
		.INIT('h1)
	) name2945 (
		_w3078_,
		_w3079_,
		_w3081_
	);
	LUT2 #(
		.INIT('h8)
	) name2946 (
		_w3080_,
		_w3081_,
		_w3082_
	);
	LUT2 #(
		.INIT('h2)
	) name2947 (
		\shift[6] ,
		_w3082_,
		_w3083_
	);
	LUT2 #(
		.INIT('h1)
	) name2948 (
		_w3075_,
		_w3083_,
		_w3084_
	);
	LUT2 #(
		.INIT('h1)
	) name2949 (
		\shift[6] ,
		_w504_,
		_w3085_
	);
	LUT2 #(
		.INIT('h2)
	) name2950 (
		\shift[6] ,
		_w322_,
		_w3086_
	);
	LUT2 #(
		.INIT('h1)
	) name2951 (
		_w3085_,
		_w3086_,
		_w3087_
	);
	LUT2 #(
		.INIT('h1)
	) name2952 (
		\shift[6] ,
		_w925_,
		_w3088_
	);
	LUT2 #(
		.INIT('h2)
	) name2953 (
		\shift[6] ,
		_w717_,
		_w3089_
	);
	LUT2 #(
		.INIT('h1)
	) name2954 (
		_w3088_,
		_w3089_,
		_w3090_
	);
	LUT2 #(
		.INIT('h1)
	) name2955 (
		\shift[6] ,
		_w1096_,
		_w3091_
	);
	LUT2 #(
		.INIT('h2)
	) name2956 (
		\shift[6] ,
		_w1010_,
		_w3092_
	);
	LUT2 #(
		.INIT('h1)
	) name2957 (
		_w3091_,
		_w3092_,
		_w3093_
	);
	LUT2 #(
		.INIT('h1)
	) name2958 (
		\shift[6] ,
		_w1390_,
		_w3094_
	);
	LUT2 #(
		.INIT('h2)
	) name2959 (
		\shift[6] ,
		_w1245_,
		_w3095_
	);
	LUT2 #(
		.INIT('h1)
	) name2960 (
		_w3094_,
		_w3095_,
		_w3096_
	);
	LUT2 #(
		.INIT('h1)
	) name2961 (
		\shift[6] ,
		_w1463_,
		_w3097_
	);
	LUT2 #(
		.INIT('h2)
	) name2962 (
		\shift[6] ,
		_w1427_,
		_w3098_
	);
	LUT2 #(
		.INIT('h1)
	) name2963 (
		_w3097_,
		_w3098_,
		_w3099_
	);
	LUT2 #(
		.INIT('h1)
	) name2964 (
		\shift[6] ,
		_w1536_,
		_w3100_
	);
	LUT2 #(
		.INIT('h2)
	) name2965 (
		\shift[6] ,
		_w1500_,
		_w3101_
	);
	LUT2 #(
		.INIT('h1)
	) name2966 (
		_w3100_,
		_w3101_,
		_w3102_
	);
	LUT2 #(
		.INIT('h1)
	) name2967 (
		\shift[6] ,
		_w1609_,
		_w3103_
	);
	LUT2 #(
		.INIT('h2)
	) name2968 (
		\shift[6] ,
		_w1573_,
		_w3104_
	);
	LUT2 #(
		.INIT('h1)
	) name2969 (
		_w3103_,
		_w3104_,
		_w3105_
	);
	LUT2 #(
		.INIT('h1)
	) name2970 (
		\shift[6] ,
		_w1682_,
		_w3106_
	);
	LUT2 #(
		.INIT('h2)
	) name2971 (
		\shift[6] ,
		_w1646_,
		_w3107_
	);
	LUT2 #(
		.INIT('h1)
	) name2972 (
		_w3106_,
		_w3107_,
		_w3108_
	);
	LUT2 #(
		.INIT('h1)
	) name2973 (
		\shift[6] ,
		_w1755_,
		_w3109_
	);
	LUT2 #(
		.INIT('h2)
	) name2974 (
		\shift[6] ,
		_w1719_,
		_w3110_
	);
	LUT2 #(
		.INIT('h1)
	) name2975 (
		_w3109_,
		_w3110_,
		_w3111_
	);
	LUT2 #(
		.INIT('h1)
	) name2976 (
		\shift[6] ,
		_w1828_,
		_w3112_
	);
	LUT2 #(
		.INIT('h2)
	) name2977 (
		\shift[6] ,
		_w1792_,
		_w3113_
	);
	LUT2 #(
		.INIT('h1)
	) name2978 (
		_w3112_,
		_w3113_,
		_w3114_
	);
	LUT2 #(
		.INIT('h1)
	) name2979 (
		\shift[6] ,
		_w1901_,
		_w3115_
	);
	LUT2 #(
		.INIT('h2)
	) name2980 (
		\shift[6] ,
		_w1865_,
		_w3116_
	);
	LUT2 #(
		.INIT('h1)
	) name2981 (
		_w3115_,
		_w3116_,
		_w3117_
	);
	LUT2 #(
		.INIT('h1)
	) name2982 (
		\shift[6] ,
		_w1974_,
		_w3118_
	);
	LUT2 #(
		.INIT('h2)
	) name2983 (
		\shift[6] ,
		_w1938_,
		_w3119_
	);
	LUT2 #(
		.INIT('h1)
	) name2984 (
		_w3118_,
		_w3119_,
		_w3120_
	);
	LUT2 #(
		.INIT('h1)
	) name2985 (
		\shift[6] ,
		_w2047_,
		_w3121_
	);
	LUT2 #(
		.INIT('h2)
	) name2986 (
		\shift[6] ,
		_w2011_,
		_w3122_
	);
	LUT2 #(
		.INIT('h1)
	) name2987 (
		_w3121_,
		_w3122_,
		_w3123_
	);
	LUT2 #(
		.INIT('h1)
	) name2988 (
		\shift[6] ,
		_w2120_,
		_w3124_
	);
	LUT2 #(
		.INIT('h2)
	) name2989 (
		\shift[6] ,
		_w2084_,
		_w3125_
	);
	LUT2 #(
		.INIT('h1)
	) name2990 (
		_w3124_,
		_w3125_,
		_w3126_
	);
	LUT2 #(
		.INIT('h1)
	) name2991 (
		\shift[6] ,
		_w2193_,
		_w3127_
	);
	LUT2 #(
		.INIT('h2)
	) name2992 (
		\shift[6] ,
		_w2157_,
		_w3128_
	);
	LUT2 #(
		.INIT('h1)
	) name2993 (
		_w3127_,
		_w3128_,
		_w3129_
	);
	LUT2 #(
		.INIT('h1)
	) name2994 (
		\shift[6] ,
		_w2266_,
		_w3130_
	);
	LUT2 #(
		.INIT('h2)
	) name2995 (
		\shift[6] ,
		_w2230_,
		_w3131_
	);
	LUT2 #(
		.INIT('h1)
	) name2996 (
		_w3130_,
		_w3131_,
		_w3132_
	);
	LUT2 #(
		.INIT('h1)
	) name2997 (
		\shift[6] ,
		_w2283_,
		_w3133_
	);
	LUT2 #(
		.INIT('h2)
	) name2998 (
		\shift[6] ,
		_w2275_,
		_w3134_
	);
	LUT2 #(
		.INIT('h1)
	) name2999 (
		_w3133_,
		_w3134_,
		_w3135_
	);
	LUT2 #(
		.INIT('h1)
	) name3000 (
		\shift[6] ,
		_w2300_,
		_w3136_
	);
	LUT2 #(
		.INIT('h2)
	) name3001 (
		\shift[6] ,
		_w2292_,
		_w3137_
	);
	LUT2 #(
		.INIT('h1)
	) name3002 (
		_w3136_,
		_w3137_,
		_w3138_
	);
	LUT2 #(
		.INIT('h1)
	) name3003 (
		\shift[6] ,
		_w2317_,
		_w3139_
	);
	LUT2 #(
		.INIT('h2)
	) name3004 (
		\shift[6] ,
		_w2309_,
		_w3140_
	);
	LUT2 #(
		.INIT('h1)
	) name3005 (
		_w3139_,
		_w3140_,
		_w3141_
	);
	LUT2 #(
		.INIT('h1)
	) name3006 (
		\shift[6] ,
		_w2334_,
		_w3142_
	);
	LUT2 #(
		.INIT('h2)
	) name3007 (
		\shift[6] ,
		_w2326_,
		_w3143_
	);
	LUT2 #(
		.INIT('h1)
	) name3008 (
		_w3142_,
		_w3143_,
		_w3144_
	);
	LUT2 #(
		.INIT('h1)
	) name3009 (
		\shift[6] ,
		_w2351_,
		_w3145_
	);
	LUT2 #(
		.INIT('h2)
	) name3010 (
		\shift[6] ,
		_w2343_,
		_w3146_
	);
	LUT2 #(
		.INIT('h1)
	) name3011 (
		_w3145_,
		_w3146_,
		_w3147_
	);
	LUT2 #(
		.INIT('h1)
	) name3012 (
		\shift[6] ,
		_w2368_,
		_w3148_
	);
	LUT2 #(
		.INIT('h2)
	) name3013 (
		\shift[6] ,
		_w2360_,
		_w3149_
	);
	LUT2 #(
		.INIT('h1)
	) name3014 (
		_w3148_,
		_w3149_,
		_w3150_
	);
	LUT2 #(
		.INIT('h1)
	) name3015 (
		\shift[6] ,
		_w2385_,
		_w3151_
	);
	LUT2 #(
		.INIT('h2)
	) name3016 (
		\shift[6] ,
		_w2377_,
		_w3152_
	);
	LUT2 #(
		.INIT('h1)
	) name3017 (
		_w3151_,
		_w3152_,
		_w3153_
	);
	LUT2 #(
		.INIT('h1)
	) name3018 (
		\shift[6] ,
		_w2402_,
		_w3154_
	);
	LUT2 #(
		.INIT('h2)
	) name3019 (
		\shift[6] ,
		_w2394_,
		_w3155_
	);
	LUT2 #(
		.INIT('h1)
	) name3020 (
		_w3154_,
		_w3155_,
		_w3156_
	);
	LUT2 #(
		.INIT('h1)
	) name3021 (
		\shift[6] ,
		_w2419_,
		_w3157_
	);
	LUT2 #(
		.INIT('h2)
	) name3022 (
		\shift[6] ,
		_w2411_,
		_w3158_
	);
	LUT2 #(
		.INIT('h1)
	) name3023 (
		_w3157_,
		_w3158_,
		_w3159_
	);
	LUT2 #(
		.INIT('h1)
	) name3024 (
		\shift[6] ,
		_w2436_,
		_w3160_
	);
	LUT2 #(
		.INIT('h2)
	) name3025 (
		\shift[6] ,
		_w2428_,
		_w3161_
	);
	LUT2 #(
		.INIT('h1)
	) name3026 (
		_w3160_,
		_w3161_,
		_w3162_
	);
	LUT2 #(
		.INIT('h1)
	) name3027 (
		\shift[6] ,
		_w2453_,
		_w3163_
	);
	LUT2 #(
		.INIT('h2)
	) name3028 (
		\shift[6] ,
		_w2445_,
		_w3164_
	);
	LUT2 #(
		.INIT('h1)
	) name3029 (
		_w3163_,
		_w3164_,
		_w3165_
	);
	LUT2 #(
		.INIT('h1)
	) name3030 (
		\shift[6] ,
		_w2470_,
		_w3166_
	);
	LUT2 #(
		.INIT('h2)
	) name3031 (
		\shift[6] ,
		_w2462_,
		_w3167_
	);
	LUT2 #(
		.INIT('h1)
	) name3032 (
		_w3166_,
		_w3167_,
		_w3168_
	);
	LUT2 #(
		.INIT('h1)
	) name3033 (
		\shift[6] ,
		_w2487_,
		_w3169_
	);
	LUT2 #(
		.INIT('h2)
	) name3034 (
		\shift[6] ,
		_w2479_,
		_w3170_
	);
	LUT2 #(
		.INIT('h1)
	) name3035 (
		_w3169_,
		_w3170_,
		_w3171_
	);
	LUT2 #(
		.INIT('h1)
	) name3036 (
		\shift[6] ,
		_w2504_,
		_w3172_
	);
	LUT2 #(
		.INIT('h2)
	) name3037 (
		\shift[6] ,
		_w2496_,
		_w3173_
	);
	LUT2 #(
		.INIT('h1)
	) name3038 (
		_w3172_,
		_w3173_,
		_w3174_
	);
	LUT2 #(
		.INIT('h1)
	) name3039 (
		\shift[6] ,
		_w2521_,
		_w3175_
	);
	LUT2 #(
		.INIT('h2)
	) name3040 (
		\shift[6] ,
		_w2513_,
		_w3176_
	);
	LUT2 #(
		.INIT('h1)
	) name3041 (
		_w3175_,
		_w3176_,
		_w3177_
	);
	LUT2 #(
		.INIT('h1)
	) name3042 (
		\shift[6] ,
		_w2538_,
		_w3178_
	);
	LUT2 #(
		.INIT('h2)
	) name3043 (
		\shift[6] ,
		_w2530_,
		_w3179_
	);
	LUT2 #(
		.INIT('h1)
	) name3044 (
		_w3178_,
		_w3179_,
		_w3180_
	);
	LUT2 #(
		.INIT('h1)
	) name3045 (
		\shift[6] ,
		_w2555_,
		_w3181_
	);
	LUT2 #(
		.INIT('h2)
	) name3046 (
		\shift[6] ,
		_w2547_,
		_w3182_
	);
	LUT2 #(
		.INIT('h1)
	) name3047 (
		_w3181_,
		_w3182_,
		_w3183_
	);
	LUT2 #(
		.INIT('h1)
	) name3048 (
		\shift[6] ,
		_w2572_,
		_w3184_
	);
	LUT2 #(
		.INIT('h2)
	) name3049 (
		\shift[6] ,
		_w2564_,
		_w3185_
	);
	LUT2 #(
		.INIT('h1)
	) name3050 (
		_w3184_,
		_w3185_,
		_w3186_
	);
	LUT2 #(
		.INIT('h1)
	) name3051 (
		\shift[6] ,
		_w2589_,
		_w3187_
	);
	LUT2 #(
		.INIT('h2)
	) name3052 (
		\shift[6] ,
		_w2581_,
		_w3188_
	);
	LUT2 #(
		.INIT('h1)
	) name3053 (
		_w3187_,
		_w3188_,
		_w3189_
	);
	LUT2 #(
		.INIT('h1)
	) name3054 (
		\shift[6] ,
		_w2606_,
		_w3190_
	);
	LUT2 #(
		.INIT('h2)
	) name3055 (
		\shift[6] ,
		_w2598_,
		_w3191_
	);
	LUT2 #(
		.INIT('h1)
	) name3056 (
		_w3190_,
		_w3191_,
		_w3192_
	);
	LUT2 #(
		.INIT('h1)
	) name3057 (
		\shift[6] ,
		_w2623_,
		_w3193_
	);
	LUT2 #(
		.INIT('h2)
	) name3058 (
		\shift[6] ,
		_w2615_,
		_w3194_
	);
	LUT2 #(
		.INIT('h1)
	) name3059 (
		_w3193_,
		_w3194_,
		_w3195_
	);
	LUT2 #(
		.INIT('h1)
	) name3060 (
		\shift[6] ,
		_w2640_,
		_w3196_
	);
	LUT2 #(
		.INIT('h2)
	) name3061 (
		\shift[6] ,
		_w2632_,
		_w3197_
	);
	LUT2 #(
		.INIT('h1)
	) name3062 (
		_w3196_,
		_w3197_,
		_w3198_
	);
	LUT2 #(
		.INIT('h1)
	) name3063 (
		\shift[6] ,
		_w2657_,
		_w3199_
	);
	LUT2 #(
		.INIT('h2)
	) name3064 (
		\shift[6] ,
		_w2649_,
		_w3200_
	);
	LUT2 #(
		.INIT('h1)
	) name3065 (
		_w3199_,
		_w3200_,
		_w3201_
	);
	LUT2 #(
		.INIT('h1)
	) name3066 (
		\shift[6] ,
		_w2674_,
		_w3202_
	);
	LUT2 #(
		.INIT('h2)
	) name3067 (
		\shift[6] ,
		_w2666_,
		_w3203_
	);
	LUT2 #(
		.INIT('h1)
	) name3068 (
		_w3202_,
		_w3203_,
		_w3204_
	);
	LUT2 #(
		.INIT('h1)
	) name3069 (
		\shift[6] ,
		_w2691_,
		_w3205_
	);
	LUT2 #(
		.INIT('h2)
	) name3070 (
		\shift[6] ,
		_w2683_,
		_w3206_
	);
	LUT2 #(
		.INIT('h1)
	) name3071 (
		_w3205_,
		_w3206_,
		_w3207_
	);
	LUT2 #(
		.INIT('h1)
	) name3072 (
		\shift[6] ,
		_w2708_,
		_w3208_
	);
	LUT2 #(
		.INIT('h2)
	) name3073 (
		\shift[6] ,
		_w2700_,
		_w3209_
	);
	LUT2 #(
		.INIT('h1)
	) name3074 (
		_w3208_,
		_w3209_,
		_w3210_
	);
	LUT2 #(
		.INIT('h1)
	) name3075 (
		\shift[6] ,
		_w2725_,
		_w3211_
	);
	LUT2 #(
		.INIT('h2)
	) name3076 (
		\shift[6] ,
		_w2717_,
		_w3212_
	);
	LUT2 #(
		.INIT('h1)
	) name3077 (
		_w3211_,
		_w3212_,
		_w3213_
	);
	LUT2 #(
		.INIT('h1)
	) name3078 (
		\shift[6] ,
		_w2742_,
		_w3214_
	);
	LUT2 #(
		.INIT('h2)
	) name3079 (
		\shift[6] ,
		_w2734_,
		_w3215_
	);
	LUT2 #(
		.INIT('h1)
	) name3080 (
		_w3214_,
		_w3215_,
		_w3216_
	);
	LUT2 #(
		.INIT('h1)
	) name3081 (
		\shift[6] ,
		_w2759_,
		_w3217_
	);
	LUT2 #(
		.INIT('h2)
	) name3082 (
		\shift[6] ,
		_w2751_,
		_w3218_
	);
	LUT2 #(
		.INIT('h1)
	) name3083 (
		_w3217_,
		_w3218_,
		_w3219_
	);
	LUT2 #(
		.INIT('h1)
	) name3084 (
		\shift[6] ,
		_w2776_,
		_w3220_
	);
	LUT2 #(
		.INIT('h2)
	) name3085 (
		\shift[6] ,
		_w2768_,
		_w3221_
	);
	LUT2 #(
		.INIT('h1)
	) name3086 (
		_w3220_,
		_w3221_,
		_w3222_
	);
	LUT2 #(
		.INIT('h1)
	) name3087 (
		\shift[6] ,
		_w2793_,
		_w3223_
	);
	LUT2 #(
		.INIT('h2)
	) name3088 (
		\shift[6] ,
		_w2785_,
		_w3224_
	);
	LUT2 #(
		.INIT('h1)
	) name3089 (
		_w3223_,
		_w3224_,
		_w3225_
	);
	LUT2 #(
		.INIT('h1)
	) name3090 (
		\shift[6] ,
		_w2810_,
		_w3226_
	);
	LUT2 #(
		.INIT('h2)
	) name3091 (
		\shift[6] ,
		_w2802_,
		_w3227_
	);
	LUT2 #(
		.INIT('h1)
	) name3092 (
		_w3226_,
		_w3227_,
		_w3228_
	);
	LUT2 #(
		.INIT('h1)
	) name3093 (
		\shift[6] ,
		_w2827_,
		_w3229_
	);
	LUT2 #(
		.INIT('h2)
	) name3094 (
		\shift[6] ,
		_w2819_,
		_w3230_
	);
	LUT2 #(
		.INIT('h1)
	) name3095 (
		_w3229_,
		_w3230_,
		_w3231_
	);
	LUT2 #(
		.INIT('h1)
	) name3096 (
		\shift[6] ,
		_w2844_,
		_w3232_
	);
	LUT2 #(
		.INIT('h2)
	) name3097 (
		\shift[6] ,
		_w2836_,
		_w3233_
	);
	LUT2 #(
		.INIT('h1)
	) name3098 (
		_w3232_,
		_w3233_,
		_w3234_
	);
	LUT2 #(
		.INIT('h1)
	) name3099 (
		\shift[6] ,
		_w2861_,
		_w3235_
	);
	LUT2 #(
		.INIT('h2)
	) name3100 (
		\shift[6] ,
		_w2853_,
		_w3236_
	);
	LUT2 #(
		.INIT('h1)
	) name3101 (
		_w3235_,
		_w3236_,
		_w3237_
	);
	LUT2 #(
		.INIT('h1)
	) name3102 (
		\shift[6] ,
		_w2878_,
		_w3238_
	);
	LUT2 #(
		.INIT('h2)
	) name3103 (
		\shift[6] ,
		_w2870_,
		_w3239_
	);
	LUT2 #(
		.INIT('h1)
	) name3104 (
		_w3238_,
		_w3239_,
		_w3240_
	);
	LUT2 #(
		.INIT('h1)
	) name3105 (
		\shift[6] ,
		_w2895_,
		_w3241_
	);
	LUT2 #(
		.INIT('h2)
	) name3106 (
		\shift[6] ,
		_w2887_,
		_w3242_
	);
	LUT2 #(
		.INIT('h1)
	) name3107 (
		_w3241_,
		_w3242_,
		_w3243_
	);
	LUT2 #(
		.INIT('h1)
	) name3108 (
		\shift[6] ,
		_w2912_,
		_w3244_
	);
	LUT2 #(
		.INIT('h2)
	) name3109 (
		\shift[6] ,
		_w2904_,
		_w3245_
	);
	LUT2 #(
		.INIT('h1)
	) name3110 (
		_w3244_,
		_w3245_,
		_w3246_
	);
	LUT2 #(
		.INIT('h1)
	) name3111 (
		\shift[6] ,
		_w2929_,
		_w3247_
	);
	LUT2 #(
		.INIT('h2)
	) name3112 (
		\shift[6] ,
		_w2921_,
		_w3248_
	);
	LUT2 #(
		.INIT('h1)
	) name3113 (
		_w3247_,
		_w3248_,
		_w3249_
	);
	LUT2 #(
		.INIT('h1)
	) name3114 (
		\shift[6] ,
		_w2946_,
		_w3250_
	);
	LUT2 #(
		.INIT('h2)
	) name3115 (
		\shift[6] ,
		_w2938_,
		_w3251_
	);
	LUT2 #(
		.INIT('h1)
	) name3116 (
		_w3250_,
		_w3251_,
		_w3252_
	);
	LUT2 #(
		.INIT('h1)
	) name3117 (
		\shift[6] ,
		_w2963_,
		_w3253_
	);
	LUT2 #(
		.INIT('h2)
	) name3118 (
		\shift[6] ,
		_w2955_,
		_w3254_
	);
	LUT2 #(
		.INIT('h1)
	) name3119 (
		_w3253_,
		_w3254_,
		_w3255_
	);
	LUT2 #(
		.INIT('h1)
	) name3120 (
		\shift[6] ,
		_w2980_,
		_w3256_
	);
	LUT2 #(
		.INIT('h2)
	) name3121 (
		\shift[6] ,
		_w2972_,
		_w3257_
	);
	LUT2 #(
		.INIT('h1)
	) name3122 (
		_w3256_,
		_w3257_,
		_w3258_
	);
	LUT2 #(
		.INIT('h1)
	) name3123 (
		\shift[6] ,
		_w2997_,
		_w3259_
	);
	LUT2 #(
		.INIT('h2)
	) name3124 (
		\shift[6] ,
		_w2989_,
		_w3260_
	);
	LUT2 #(
		.INIT('h1)
	) name3125 (
		_w3259_,
		_w3260_,
		_w3261_
	);
	LUT2 #(
		.INIT('h1)
	) name3126 (
		\shift[6] ,
		_w3014_,
		_w3262_
	);
	LUT2 #(
		.INIT('h2)
	) name3127 (
		\shift[6] ,
		_w3006_,
		_w3263_
	);
	LUT2 #(
		.INIT('h1)
	) name3128 (
		_w3262_,
		_w3263_,
		_w3264_
	);
	LUT2 #(
		.INIT('h1)
	) name3129 (
		\shift[6] ,
		_w3031_,
		_w3265_
	);
	LUT2 #(
		.INIT('h2)
	) name3130 (
		\shift[6] ,
		_w3023_,
		_w3266_
	);
	LUT2 #(
		.INIT('h1)
	) name3131 (
		_w3265_,
		_w3266_,
		_w3267_
	);
	LUT2 #(
		.INIT('h1)
	) name3132 (
		\shift[6] ,
		_w3048_,
		_w3268_
	);
	LUT2 #(
		.INIT('h2)
	) name3133 (
		\shift[6] ,
		_w3040_,
		_w3269_
	);
	LUT2 #(
		.INIT('h1)
	) name3134 (
		_w3268_,
		_w3269_,
		_w3270_
	);
	LUT2 #(
		.INIT('h1)
	) name3135 (
		\shift[6] ,
		_w3065_,
		_w3271_
	);
	LUT2 #(
		.INIT('h2)
	) name3136 (
		\shift[6] ,
		_w3057_,
		_w3272_
	);
	LUT2 #(
		.INIT('h1)
	) name3137 (
		_w3271_,
		_w3272_,
		_w3273_
	);
	LUT2 #(
		.INIT('h1)
	) name3138 (
		\shift[6] ,
		_w3082_,
		_w3274_
	);
	LUT2 #(
		.INIT('h2)
	) name3139 (
		\shift[6] ,
		_w3074_,
		_w3275_
	);
	LUT2 #(
		.INIT('h1)
	) name3140 (
		_w3274_,
		_w3275_,
		_w3276_
	);
	assign \result[0]  = _w506_ ;
	assign \result[1]  = _w927_ ;
	assign \result[2]  = _w1098_ ;
	assign \result[3]  = _w1392_ ;
	assign \result[4]  = _w1465_ ;
	assign \result[5]  = _w1538_ ;
	assign \result[6]  = _w1611_ ;
	assign \result[7]  = _w1684_ ;
	assign \result[8]  = _w1757_ ;
	assign \result[9]  = _w1830_ ;
	assign \result[10]  = _w1903_ ;
	assign \result[11]  = _w1976_ ;
	assign \result[12]  = _w2049_ ;
	assign \result[13]  = _w2122_ ;
	assign \result[14]  = _w2195_ ;
	assign \result[15]  = _w2268_ ;
	assign \result[16]  = _w2285_ ;
	assign \result[17]  = _w2302_ ;
	assign \result[18]  = _w2319_ ;
	assign \result[19]  = _w2336_ ;
	assign \result[20]  = _w2353_ ;
	assign \result[21]  = _w2370_ ;
	assign \result[22]  = _w2387_ ;
	assign \result[23]  = _w2404_ ;
	assign \result[24]  = _w2421_ ;
	assign \result[25]  = _w2438_ ;
	assign \result[26]  = _w2455_ ;
	assign \result[27]  = _w2472_ ;
	assign \result[28]  = _w2489_ ;
	assign \result[29]  = _w2506_ ;
	assign \result[30]  = _w2523_ ;
	assign \result[31]  = _w2540_ ;
	assign \result[32]  = _w2557_ ;
	assign \result[33]  = _w2574_ ;
	assign \result[34]  = _w2591_ ;
	assign \result[35]  = _w2608_ ;
	assign \result[36]  = _w2625_ ;
	assign \result[37]  = _w2642_ ;
	assign \result[38]  = _w2659_ ;
	assign \result[39]  = _w2676_ ;
	assign \result[40]  = _w2693_ ;
	assign \result[41]  = _w2710_ ;
	assign \result[42]  = _w2727_ ;
	assign \result[43]  = _w2744_ ;
	assign \result[44]  = _w2761_ ;
	assign \result[45]  = _w2778_ ;
	assign \result[46]  = _w2795_ ;
	assign \result[47]  = _w2812_ ;
	assign \result[48]  = _w2829_ ;
	assign \result[49]  = _w2846_ ;
	assign \result[50]  = _w2863_ ;
	assign \result[51]  = _w2880_ ;
	assign \result[52]  = _w2897_ ;
	assign \result[53]  = _w2914_ ;
	assign \result[54]  = _w2931_ ;
	assign \result[55]  = _w2948_ ;
	assign \result[56]  = _w2965_ ;
	assign \result[57]  = _w2982_ ;
	assign \result[58]  = _w2999_ ;
	assign \result[59]  = _w3016_ ;
	assign \result[60]  = _w3033_ ;
	assign \result[61]  = _w3050_ ;
	assign \result[62]  = _w3067_ ;
	assign \result[63]  = _w3084_ ;
	assign \result[64]  = _w3087_ ;
	assign \result[65]  = _w3090_ ;
	assign \result[66]  = _w3093_ ;
	assign \result[67]  = _w3096_ ;
	assign \result[68]  = _w3099_ ;
	assign \result[69]  = _w3102_ ;
	assign \result[70]  = _w3105_ ;
	assign \result[71]  = _w3108_ ;
	assign \result[72]  = _w3111_ ;
	assign \result[73]  = _w3114_ ;
	assign \result[74]  = _w3117_ ;
	assign \result[75]  = _w3120_ ;
	assign \result[76]  = _w3123_ ;
	assign \result[77]  = _w3126_ ;
	assign \result[78]  = _w3129_ ;
	assign \result[79]  = _w3132_ ;
	assign \result[80]  = _w3135_ ;
	assign \result[81]  = _w3138_ ;
	assign \result[82]  = _w3141_ ;
	assign \result[83]  = _w3144_ ;
	assign \result[84]  = _w3147_ ;
	assign \result[85]  = _w3150_ ;
	assign \result[86]  = _w3153_ ;
	assign \result[87]  = _w3156_ ;
	assign \result[88]  = _w3159_ ;
	assign \result[89]  = _w3162_ ;
	assign \result[90]  = _w3165_ ;
	assign \result[91]  = _w3168_ ;
	assign \result[92]  = _w3171_ ;
	assign \result[93]  = _w3174_ ;
	assign \result[94]  = _w3177_ ;
	assign \result[95]  = _w3180_ ;
	assign \result[96]  = _w3183_ ;
	assign \result[97]  = _w3186_ ;
	assign \result[98]  = _w3189_ ;
	assign \result[99]  = _w3192_ ;
	assign \result[100]  = _w3195_ ;
	assign \result[101]  = _w3198_ ;
	assign \result[102]  = _w3201_ ;
	assign \result[103]  = _w3204_ ;
	assign \result[104]  = _w3207_ ;
	assign \result[105]  = _w3210_ ;
	assign \result[106]  = _w3213_ ;
	assign \result[107]  = _w3216_ ;
	assign \result[108]  = _w3219_ ;
	assign \result[109]  = _w3222_ ;
	assign \result[110]  = _w3225_ ;
	assign \result[111]  = _w3228_ ;
	assign \result[112]  = _w3231_ ;
	assign \result[113]  = _w3234_ ;
	assign \result[114]  = _w3237_ ;
	assign \result[115]  = _w3240_ ;
	assign \result[116]  = _w3243_ ;
	assign \result[117]  = _w3246_ ;
	assign \result[118]  = _w3249_ ;
	assign \result[119]  = _w3252_ ;
	assign \result[120]  = _w3255_ ;
	assign \result[121]  = _w3258_ ;
	assign \result[122]  = _w3261_ ;
	assign \result[123]  = _w3264_ ;
	assign \result[124]  = _w3267_ ;
	assign \result[125]  = _w3270_ ;
	assign \result[126]  = _w3273_ ;
	assign \result[127]  = _w3276_ ;
endmodule;