module top (\1(0)_pad , \100(77)_pad , \101(78)_pad , \102(79)_pad , \103(80)_pad , \104(81)_pad , \105(82)_pad , \106(83)_pad , \107(84)_pad , \108(85)_pad , \11(8)_pad , \111(86)_pad , \112(87)_pad , \113(88)_pad , \114(89)_pad , \115(90)_pad , \116(91)_pad , \117(92)_pad , \118(93)_pad , \119(94)_pad , \120(95)_pad , \123(96)_pad , \124(97)_pad , \125(98)_pad , \126(99)_pad , \127(100)_pad , \128(101)_pad , \129(102)_pad , \130(103)_pad , \131(104)_pad , \132(105)_pad , \1341(200)_pad , \1348(201)_pad , \135(106)_pad , \136(107)_pad , \137(108)_pad , \138(109)_pad , \1384(202)_pad , \139(110)_pad , \14(9)_pad , \140(111)_pad , \141(112)_pad , \142(113)_pad , \15(10)_pad , \16(11)_pad , \19(12)_pad , \1956(203)_pad , \1961(204)_pad , \1966(205)_pad , \1971(206)_pad , \1976(207)_pad , \1981(208)_pad , \1986(209)_pad , \1991(210)_pad , \1996(211)_pad , \2(1)_pad , \20(13)_pad , \2067(213)_pad , \2072(214)_pad , \2078(215)_pad , \2084(216)_pad , \2090(217)_pad , \2096(218)_pad , \21(14)_pad , \2100(219)_pad , \2104(220)_pad , \2105(221)_pad , \2106(222)_pad , \22(15)_pad , \23(16)_pad , \24(17)_pad , \2427(223)_pad , \2430(224)_pad , \2435(225)_pad , \2438(226)_pad , \2443(227)_pad , \2446(228)_pad , \2451(229)_pad , \2454(230)_pad , \2474(231)_pad , \25(18)_pad , \26(19)_pad , \2678(232)_pad , \27(20)_pad , \28(21)_pad , \29(22)_pad , \3(2)_pad , \32(23)_pad , \33(24)_pad , \34(25)_pad , \35(26)_pad , \36(27)_pad , \37(28)_pad , \4(3)_pad , \40(29)_pad , \409(298)_pad , \43(30)_pad , \44(31)_pad , \47(32)_pad , \48(33)_pad , \483(191)_pad , \49(34)_pad , \5(4)_pad , \50(35)_pad , \51(36)_pad , \52(37)_pad , \53(38)_pad , \54(39)_pad , \543(192)_pad , \55(40)_pad , \559(193)_pad , \56(41)_pad , \567(194)_pad , \57(42)_pad , \6(5)_pad , \60(43)_pad , \61(44)_pad , \62(45)_pad , \63(46)_pad , \64(47)_pad , \65(48)_pad , \651(195)_pad , \66(49)_pad , \661(196)_pad , \67(50)_pad , \68(51)_pad , \69(52)_pad , \7(6)_pad , \72(53)_pad , \73(54)_pad , \74(55)_pad , \75(56)_pad , \76(57)_pad , \77(58)_pad , \78(59)_pad , \79(60)_pad , \8(7)_pad , \80(61)_pad , \81(62)_pad , \82(63)_pad , \85(64)_pad , \86(65)_pad , \860(197)_pad , \868(198)_pad , \87(66)_pad , \88(67)_pad , \89(68)_pad , \90(69)_pad , \91(70)_pad , \92(71)_pad , \93(72)_pad , \94(73)_pad , \95(74)_pad , \96(75)_pad , \99(76)_pad , \145(1358)_pad , \148(851)_pad , \150(1277)_pad , \153(671)_pad , \156(1046)_pad , \158(349)_pad , \160(609)_pad , \162(612)_pad , \164(607)_pad , \166(625)_pad , \168(623)_pad , \171(621)_pad , \173(389)_pad , \176(803)_pad , \188(761)_pad , \217(423)_pad , \218(311)_pad , \219(302)_pad , \220(306)_pad , \221(305)_pad , \223(413)_pad , \225(1424)_pad , \227(1179)_pad , \229(1180)_pad , \234(376)_pad , \235(307)_pad , \236(303)_pad , \237(309)_pad , \238(304)_pad , \259(414)_pad , \261(506)_pad , \282(922)_pad , \284(847)_pad , \286(696)_pad , \288(700)_pad , \290(704)_pad , \295(1400)_pad , \297(849)_pad , \299(692)_pad , \301(694)_pad , \303(698)_pad , \305(702)_pad , \325(507)_pad , \329(1414)_pad , \_al_n0 , \u1082_syn_3 , \u1396_syn_3 , \u1414_syn_3 , \u1447_syn_3 , \u538_syn_3 , \u539_syn_3 );
	input \1(0)_pad  ;
	input \100(77)_pad  ;
	input \101(78)_pad  ;
	input \102(79)_pad  ;
	input \103(80)_pad  ;
	input \104(81)_pad  ;
	input \105(82)_pad  ;
	input \106(83)_pad  ;
	input \107(84)_pad  ;
	input \108(85)_pad  ;
	input \11(8)_pad  ;
	input \111(86)_pad  ;
	input \112(87)_pad  ;
	input \113(88)_pad  ;
	input \114(89)_pad  ;
	input \115(90)_pad  ;
	input \116(91)_pad  ;
	input \117(92)_pad  ;
	input \118(93)_pad  ;
	input \119(94)_pad  ;
	input \120(95)_pad  ;
	input \123(96)_pad  ;
	input \124(97)_pad  ;
	input \125(98)_pad  ;
	input \126(99)_pad  ;
	input \127(100)_pad  ;
	input \128(101)_pad  ;
	input \129(102)_pad  ;
	input \130(103)_pad  ;
	input \131(104)_pad  ;
	input \132(105)_pad  ;
	input \1341(200)_pad  ;
	input \1348(201)_pad  ;
	input \135(106)_pad  ;
	input \136(107)_pad  ;
	input \137(108)_pad  ;
	input \138(109)_pad  ;
	input \1384(202)_pad  ;
	input \139(110)_pad  ;
	input \14(9)_pad  ;
	input \140(111)_pad  ;
	input \141(112)_pad  ;
	input \142(113)_pad  ;
	input \15(10)_pad  ;
	input \16(11)_pad  ;
	input \19(12)_pad  ;
	input \1956(203)_pad  ;
	input \1961(204)_pad  ;
	input \1966(205)_pad  ;
	input \1971(206)_pad  ;
	input \1976(207)_pad  ;
	input \1981(208)_pad  ;
	input \1986(209)_pad  ;
	input \1991(210)_pad  ;
	input \1996(211)_pad  ;
	input \2(1)_pad  ;
	input \20(13)_pad  ;
	input \2067(213)_pad  ;
	input \2072(214)_pad  ;
	input \2078(215)_pad  ;
	input \2084(216)_pad  ;
	input \2090(217)_pad  ;
	input \2096(218)_pad  ;
	input \21(14)_pad  ;
	input \2100(219)_pad  ;
	input \2104(220)_pad  ;
	input \2105(221)_pad  ;
	input \2106(222)_pad  ;
	input \22(15)_pad  ;
	input \23(16)_pad  ;
	input \24(17)_pad  ;
	input \2427(223)_pad  ;
	input \2430(224)_pad  ;
	input \2435(225)_pad  ;
	input \2438(226)_pad  ;
	input \2443(227)_pad  ;
	input \2446(228)_pad  ;
	input \2451(229)_pad  ;
	input \2454(230)_pad  ;
	input \2474(231)_pad  ;
	input \25(18)_pad  ;
	input \26(19)_pad  ;
	input \2678(232)_pad  ;
	input \27(20)_pad  ;
	input \28(21)_pad  ;
	input \29(22)_pad  ;
	input \3(2)_pad  ;
	input \32(23)_pad  ;
	input \33(24)_pad  ;
	input \34(25)_pad  ;
	input \35(26)_pad  ;
	input \36(27)_pad  ;
	input \37(28)_pad  ;
	input \4(3)_pad  ;
	input \40(29)_pad  ;
	input \409(298)_pad  ;
	input \43(30)_pad  ;
	input \44(31)_pad  ;
	input \47(32)_pad  ;
	input \48(33)_pad  ;
	input \483(191)_pad  ;
	input \49(34)_pad  ;
	input \5(4)_pad  ;
	input \50(35)_pad  ;
	input \51(36)_pad  ;
	input \52(37)_pad  ;
	input \53(38)_pad  ;
	input \54(39)_pad  ;
	input \543(192)_pad  ;
	input \55(40)_pad  ;
	input \559(193)_pad  ;
	input \56(41)_pad  ;
	input \567(194)_pad  ;
	input \57(42)_pad  ;
	input \6(5)_pad  ;
	input \60(43)_pad  ;
	input \61(44)_pad  ;
	input \62(45)_pad  ;
	input \63(46)_pad  ;
	input \64(47)_pad  ;
	input \65(48)_pad  ;
	input \651(195)_pad  ;
	input \66(49)_pad  ;
	input \661(196)_pad  ;
	input \67(50)_pad  ;
	input \68(51)_pad  ;
	input \69(52)_pad  ;
	input \7(6)_pad  ;
	input \72(53)_pad  ;
	input \73(54)_pad  ;
	input \74(55)_pad  ;
	input \75(56)_pad  ;
	input \76(57)_pad  ;
	input \77(58)_pad  ;
	input \78(59)_pad  ;
	input \79(60)_pad  ;
	input \8(7)_pad  ;
	input \80(61)_pad  ;
	input \81(62)_pad  ;
	input \82(63)_pad  ;
	input \85(64)_pad  ;
	input \86(65)_pad  ;
	input \860(197)_pad  ;
	input \868(198)_pad  ;
	input \87(66)_pad  ;
	input \88(67)_pad  ;
	input \89(68)_pad  ;
	input \90(69)_pad  ;
	input \91(70)_pad  ;
	input \92(71)_pad  ;
	input \93(72)_pad  ;
	input \94(73)_pad  ;
	input \95(74)_pad  ;
	input \96(75)_pad  ;
	input \99(76)_pad  ;
	output \145(1358)_pad  ;
	output \148(851)_pad  ;
	output \150(1277)_pad  ;
	output \153(671)_pad  ;
	output \156(1046)_pad  ;
	output \158(349)_pad  ;
	output \160(609)_pad  ;
	output \162(612)_pad  ;
	output \164(607)_pad  ;
	output \166(625)_pad  ;
	output \168(623)_pad  ;
	output \171(621)_pad  ;
	output \173(389)_pad  ;
	output \176(803)_pad  ;
	output \188(761)_pad  ;
	output \217(423)_pad  ;
	output \218(311)_pad  ;
	output \219(302)_pad  ;
	output \220(306)_pad  ;
	output \221(305)_pad  ;
	output \223(413)_pad  ;
	output \225(1424)_pad  ;
	output \227(1179)_pad  ;
	output \229(1180)_pad  ;
	output \234(376)_pad  ;
	output \235(307)_pad  ;
	output \236(303)_pad  ;
	output \237(309)_pad  ;
	output \238(304)_pad  ;
	output \259(414)_pad  ;
	output \261(506)_pad  ;
	output \282(922)_pad  ;
	output \284(847)_pad  ;
	output \286(696)_pad  ;
	output \288(700)_pad  ;
	output \290(704)_pad  ;
	output \295(1400)_pad  ;
	output \297(849)_pad  ;
	output \299(692)_pad  ;
	output \301(694)_pad  ;
	output \303(698)_pad  ;
	output \305(702)_pad  ;
	output \325(507)_pad  ;
	output \329(1414)_pad  ;
	output \_al_n0  ;
	output \u1082_syn_3  ;
	output \u1396_syn_3  ;
	output \u1414_syn_3  ;
	output \u1447_syn_3  ;
	output \u538_syn_3  ;
	output \u539_syn_3  ;
	wire _w688_ ;
	wire _w687_ ;
	wire _w686_ ;
	wire _w685_ ;
	wire _w684_ ;
	wire _w683_ ;
	wire _w682_ ;
	wire _w681_ ;
	wire _w680_ ;
	wire _w679_ ;
	wire _w678_ ;
	wire _w677_ ;
	wire _w676_ ;
	wire _w675_ ;
	wire _w674_ ;
	wire _w673_ ;
	wire _w672_ ;
	wire _w671_ ;
	wire _w670_ ;
	wire _w669_ ;
	wire _w668_ ;
	wire _w667_ ;
	wire _w666_ ;
	wire _w665_ ;
	wire _w664_ ;
	wire _w663_ ;
	wire _w662_ ;
	wire _w661_ ;
	wire _w660_ ;
	wire _w659_ ;
	wire _w658_ ;
	wire _w657_ ;
	wire _w656_ ;
	wire _w655_ ;
	wire _w654_ ;
	wire _w653_ ;
	wire _w652_ ;
	wire _w651_ ;
	wire _w650_ ;
	wire _w649_ ;
	wire _w648_ ;
	wire _w647_ ;
	wire _w646_ ;
	wire _w645_ ;
	wire _w644_ ;
	wire _w643_ ;
	wire _w642_ ;
	wire _w641_ ;
	wire _w640_ ;
	wire _w639_ ;
	wire _w638_ ;
	wire _w637_ ;
	wire _w636_ ;
	wire _w635_ ;
	wire _w634_ ;
	wire _w633_ ;
	wire _w632_ ;
	wire _w631_ ;
	wire _w630_ ;
	wire _w629_ ;
	wire _w628_ ;
	wire _w627_ ;
	wire _w626_ ;
	wire _w625_ ;
	wire _w624_ ;
	wire _w623_ ;
	wire _w622_ ;
	wire _w621_ ;
	wire _w620_ ;
	wire _w619_ ;
	wire _w618_ ;
	wire _w617_ ;
	wire _w616_ ;
	wire _w615_ ;
	wire _w614_ ;
	wire _w613_ ;
	wire _w612_ ;
	wire _w611_ ;
	wire _w610_ ;
	wire _w609_ ;
	wire _w608_ ;
	wire _w607_ ;
	wire _w606_ ;
	wire _w605_ ;
	wire _w604_ ;
	wire _w603_ ;
	wire _w602_ ;
	wire _w601_ ;
	wire _w600_ ;
	wire _w599_ ;
	wire _w598_ ;
	wire _w597_ ;
	wire _w596_ ;
	wire _w595_ ;
	wire _w594_ ;
	wire _w593_ ;
	wire _w592_ ;
	wire _w591_ ;
	wire _w590_ ;
	wire _w589_ ;
	wire _w588_ ;
	wire _w587_ ;
	wire _w586_ ;
	wire _w585_ ;
	wire _w584_ ;
	wire _w583_ ;
	wire _w582_ ;
	wire _w581_ ;
	wire _w580_ ;
	wire _w579_ ;
	wire _w578_ ;
	wire _w577_ ;
	wire _w576_ ;
	wire _w575_ ;
	wire _w574_ ;
	wire _w573_ ;
	wire _w572_ ;
	wire _w571_ ;
	wire _w570_ ;
	wire _w569_ ;
	wire _w568_ ;
	wire _w567_ ;
	wire _w566_ ;
	wire _w565_ ;
	wire _w564_ ;
	wire _w563_ ;
	wire _w562_ ;
	wire _w561_ ;
	wire _w560_ ;
	wire _w559_ ;
	wire _w558_ ;
	wire _w557_ ;
	wire _w556_ ;
	wire _w555_ ;
	wire _w554_ ;
	wire _w553_ ;
	wire _w552_ ;
	wire _w551_ ;
	wire _w550_ ;
	wire _w549_ ;
	wire _w548_ ;
	wire _w547_ ;
	wire _w546_ ;
	wire _w545_ ;
	wire _w544_ ;
	wire _w543_ ;
	wire _w542_ ;
	wire _w541_ ;
	wire _w540_ ;
	wire _w539_ ;
	wire _w538_ ;
	wire _w537_ ;
	wire _w536_ ;
	wire _w535_ ;
	wire _w534_ ;
	wire _w533_ ;
	wire _w532_ ;
	wire _w531_ ;
	wire _w530_ ;
	wire _w529_ ;
	wire _w528_ ;
	wire _w527_ ;
	wire _w526_ ;
	wire _w525_ ;
	wire _w524_ ;
	wire _w523_ ;
	wire _w522_ ;
	wire _w521_ ;
	wire _w520_ ;
	wire _w519_ ;
	wire _w518_ ;
	wire _w517_ ;
	wire _w516_ ;
	wire _w515_ ;
	wire _w514_ ;
	wire _w513_ ;
	wire _w512_ ;
	wire _w511_ ;
	wire _w510_ ;
	wire _w509_ ;
	wire _w508_ ;
	wire _w507_ ;
	wire _w506_ ;
	wire _w505_ ;
	wire _w504_ ;
	wire _w503_ ;
	wire _w502_ ;
	wire _w501_ ;
	wire _w500_ ;
	wire _w499_ ;
	wire _w498_ ;
	wire _w497_ ;
	wire _w496_ ;
	wire _w495_ ;
	wire _w494_ ;
	wire _w493_ ;
	wire _w492_ ;
	wire _w491_ ;
	wire _w490_ ;
	wire _w489_ ;
	wire _w488_ ;
	wire _w487_ ;
	wire _w486_ ;
	wire _w485_ ;
	wire _w484_ ;
	wire _w483_ ;
	wire _w482_ ;
	wire _w481_ ;
	wire _w480_ ;
	wire _w479_ ;
	wire _w478_ ;
	wire _w477_ ;
	wire _w476_ ;
	wire _w475_ ;
	wire _w474_ ;
	wire _w473_ ;
	wire _w472_ ;
	wire _w471_ ;
	wire _w470_ ;
	wire _w469_ ;
	wire _w468_ ;
	wire _w467_ ;
	wire _w466_ ;
	wire _w465_ ;
	wire _w464_ ;
	wire _w463_ ;
	wire _w462_ ;
	wire _w461_ ;
	wire _w460_ ;
	wire _w459_ ;
	wire _w458_ ;
	wire _w457_ ;
	wire _w456_ ;
	wire _w455_ ;
	wire _w454_ ;
	wire _w453_ ;
	wire _w452_ ;
	wire _w451_ ;
	wire _w450_ ;
	wire _w449_ ;
	wire _w448_ ;
	wire _w447_ ;
	wire _w446_ ;
	wire _w445_ ;
	wire _w444_ ;
	wire _w443_ ;
	wire _w442_ ;
	wire _w441_ ;
	wire _w440_ ;
	wire _w439_ ;
	wire _w438_ ;
	wire _w437_ ;
	wire _w436_ ;
	wire _w435_ ;
	wire _w434_ ;
	wire _w433_ ;
	wire _w432_ ;
	wire _w431_ ;
	wire _w430_ ;
	wire _w429_ ;
	wire _w428_ ;
	wire _w427_ ;
	wire _w426_ ;
	wire _w425_ ;
	wire _w424_ ;
	wire _w423_ ;
	wire _w422_ ;
	wire _w421_ ;
	wire _w420_ ;
	wire _w419_ ;
	wire _w418_ ;
	wire _w417_ ;
	wire _w416_ ;
	wire _w415_ ;
	wire _w414_ ;
	wire _w413_ ;
	wire _w282_ ;
	wire _w281_ ;
	wire _w280_ ;
	wire _w279_ ;
	wire _w278_ ;
	wire _w277_ ;
	wire _w276_ ;
	wire _w275_ ;
	wire _w274_ ;
	wire _w273_ ;
	wire _w272_ ;
	wire _w271_ ;
	wire _w270_ ;
	wire _w269_ ;
	wire _w268_ ;
	wire _w267_ ;
	wire _w266_ ;
	wire _w265_ ;
	wire _w264_ ;
	wire _w263_ ;
	wire _w262_ ;
	wire _w261_ ;
	wire _w260_ ;
	wire _w259_ ;
	wire _w258_ ;
	wire _w257_ ;
	wire _w256_ ;
	wire _w255_ ;
	wire _w254_ ;
	wire _w253_ ;
	wire _w252_ ;
	wire _w251_ ;
	wire _w250_ ;
	wire _w249_ ;
	wire _w248_ ;
	wire _w247_ ;
	wire _w246_ ;
	wire _w245_ ;
	wire _w244_ ;
	wire _w243_ ;
	wire _w242_ ;
	wire _w241_ ;
	wire _w240_ ;
	wire _w239_ ;
	wire _w238_ ;
	wire _w237_ ;
	wire _w236_ ;
	wire _w235_ ;
	wire _w234_ ;
	wire _w233_ ;
	wire _w232_ ;
	wire _w231_ ;
	wire _w230_ ;
	wire _w229_ ;
	wire _w228_ ;
	wire _w227_ ;
	wire _w226_ ;
	wire _w225_ ;
	wire _w224_ ;
	wire _w223_ ;
	wire _w222_ ;
	wire _w221_ ;
	wire _w220_ ;
	wire _w219_ ;
	wire _w218_ ;
	wire _w217_ ;
	wire _w216_ ;
	wire _w215_ ;
	wire _w184_ ;
	wire _w183_ ;
	wire _w182_ ;
	wire _w181_ ;
	wire _w180_ ;
	wire _w179_ ;
	wire _w178_ ;
	wire _w177_ ;
	wire _w176_ ;
	wire _w175_ ;
	wire _w174_ ;
	wire _w173_ ;
	wire _w172_ ;
	wire _w171_ ;
	wire _w170_ ;
	wire _w169_ ;
	wire _w156_ ;
	wire _w157_ ;
	wire _w158_ ;
	wire _w159_ ;
	wire _w160_ ;
	wire _w161_ ;
	wire _w162_ ;
	wire _w163_ ;
	wire _w164_ ;
	wire _w165_ ;
	wire _w166_ ;
	wire _w167_ ;
	wire _w168_ ;
	wire _w185_ ;
	wire _w186_ ;
	wire _w187_ ;
	wire _w188_ ;
	wire _w189_ ;
	wire _w190_ ;
	wire _w191_ ;
	wire _w192_ ;
	wire _w193_ ;
	wire _w194_ ;
	wire _w195_ ;
	wire _w196_ ;
	wire _w197_ ;
	wire _w198_ ;
	wire _w199_ ;
	wire _w200_ ;
	wire _w201_ ;
	wire _w202_ ;
	wire _w203_ ;
	wire _w204_ ;
	wire _w205_ ;
	wire _w206_ ;
	wire _w207_ ;
	wire _w208_ ;
	wire _w209_ ;
	wire _w210_ ;
	wire _w211_ ;
	wire _w212_ ;
	wire _w213_ ;
	wire _w214_ ;
	wire _w283_ ;
	wire _w284_ ;
	wire _w285_ ;
	wire _w286_ ;
	wire _w287_ ;
	wire _w288_ ;
	wire _w289_ ;
	wire _w290_ ;
	wire _w291_ ;
	wire _w292_ ;
	wire _w293_ ;
	wire _w294_ ;
	wire _w295_ ;
	wire _w296_ ;
	wire _w297_ ;
	wire _w298_ ;
	wire _w299_ ;
	wire _w300_ ;
	wire _w301_ ;
	wire _w302_ ;
	wire _w303_ ;
	wire _w304_ ;
	wire _w305_ ;
	wire _w306_ ;
	wire _w307_ ;
	wire _w308_ ;
	wire _w309_ ;
	wire _w310_ ;
	wire _w311_ ;
	wire _w312_ ;
	wire _w313_ ;
	wire _w314_ ;
	wire _w315_ ;
	wire _w316_ ;
	wire _w317_ ;
	wire _w318_ ;
	wire _w319_ ;
	wire _w320_ ;
	wire _w321_ ;
	wire _w322_ ;
	wire _w323_ ;
	wire _w324_ ;
	wire _w325_ ;
	wire _w326_ ;
	wire _w327_ ;
	wire _w328_ ;
	wire _w329_ ;
	wire _w330_ ;
	wire _w331_ ;
	wire _w332_ ;
	wire _w333_ ;
	wire _w334_ ;
	wire _w335_ ;
	wire _w336_ ;
	wire _w337_ ;
	wire _w338_ ;
	wire _w339_ ;
	wire _w340_ ;
	wire _w341_ ;
	wire _w342_ ;
	wire _w343_ ;
	wire _w344_ ;
	wire _w345_ ;
	wire _w346_ ;
	wire _w347_ ;
	wire _w348_ ;
	wire _w349_ ;
	wire _w350_ ;
	wire _w351_ ;
	wire _w352_ ;
	wire _w353_ ;
	wire _w354_ ;
	wire _w355_ ;
	wire _w356_ ;
	wire _w357_ ;
	wire _w358_ ;
	wire _w359_ ;
	wire _w360_ ;
	wire _w361_ ;
	wire _w362_ ;
	wire _w363_ ;
	wire _w364_ ;
	wire _w365_ ;
	wire _w366_ ;
	wire _w367_ ;
	wire _w368_ ;
	wire _w369_ ;
	wire _w370_ ;
	wire _w371_ ;
	wire _w372_ ;
	wire _w373_ ;
	wire _w374_ ;
	wire _w375_ ;
	wire _w376_ ;
	wire _w377_ ;
	wire _w378_ ;
	wire _w379_ ;
	wire _w380_ ;
	wire _w381_ ;
	wire _w382_ ;
	wire _w383_ ;
	wire _w384_ ;
	wire _w385_ ;
	wire _w386_ ;
	wire _w387_ ;
	wire _w388_ ;
	wire _w389_ ;
	wire _w390_ ;
	wire _w391_ ;
	wire _w392_ ;
	wire _w393_ ;
	wire _w394_ ;
	wire _w395_ ;
	wire _w396_ ;
	wire _w397_ ;
	wire _w398_ ;
	wire _w399_ ;
	wire _w400_ ;
	wire _w401_ ;
	wire _w402_ ;
	wire _w403_ ;
	wire _w404_ ;
	wire _w405_ ;
	wire _w406_ ;
	wire _w407_ ;
	wire _w408_ ;
	wire _w409_ ;
	wire _w410_ ;
	wire _w411_ ;
	wire _w412_ ;
	LUT2 #(
		.INIT('h2)
	) name0 (
		\543(192)_pad ,
		\651(195)_pad ,
		_w156_
	);
	LUT2 #(
		.INIT('h8)
	) name1 (
		\54(39)_pad ,
		_w156_,
		_w157_
	);
	LUT2 #(
		.INIT('h8)
	) name2 (
		\543(192)_pad ,
		\651(195)_pad ,
		_w158_
	);
	LUT2 #(
		.INIT('h8)
	) name3 (
		\79(60)_pad ,
		_w158_,
		_w159_
	);
	LUT2 #(
		.INIT('h4)
	) name4 (
		\543(192)_pad ,
		\651(195)_pad ,
		_w160_
	);
	LUT2 #(
		.INIT('h8)
	) name5 (
		\66(49)_pad ,
		_w160_,
		_w161_
	);
	LUT2 #(
		.INIT('h1)
	) name6 (
		\543(192)_pad ,
		\651(195)_pad ,
		_w162_
	);
	LUT2 #(
		.INIT('h8)
	) name7 (
		\92(71)_pad ,
		_w162_,
		_w163_
	);
	LUT2 #(
		.INIT('h1)
	) name8 (
		_w157_,
		_w159_,
		_w164_
	);
	LUT2 #(
		.INIT('h1)
	) name9 (
		_w161_,
		_w163_,
		_w165_
	);
	LUT2 #(
		.INIT('h8)
	) name10 (
		_w164_,
		_w165_,
		_w166_
	);
	LUT2 #(
		.INIT('h8)
	) name11 (
		\559(193)_pad ,
		_w166_,
		_w167_
	);
	LUT2 #(
		.INIT('h4)
	) name12 (
		\860(197)_pad ,
		_w167_,
		_w168_
	);
	LUT2 #(
		.INIT('h8)
	) name13 (
		\43(30)_pad ,
		_w156_,
		_w169_
	);
	LUT2 #(
		.INIT('h8)
	) name14 (
		\68(51)_pad ,
		_w158_,
		_w170_
	);
	LUT2 #(
		.INIT('h8)
	) name15 (
		\56(41)_pad ,
		_w160_,
		_w171_
	);
	LUT2 #(
		.INIT('h8)
	) name16 (
		\81(62)_pad ,
		_w162_,
		_w172_
	);
	LUT2 #(
		.INIT('h1)
	) name17 (
		_w169_,
		_w170_,
		_w173_
	);
	LUT2 #(
		.INIT('h1)
	) name18 (
		_w171_,
		_w172_,
		_w174_
	);
	LUT2 #(
		.INIT('h8)
	) name19 (
		_w173_,
		_w174_,
		_w175_
	);
	LUT2 #(
		.INIT('h8)
	) name20 (
		\860(197)_pad ,
		_w175_,
		_w176_
	);
	LUT2 #(
		.INIT('h1)
	) name21 (
		_w168_,
		_w176_,
		_w177_
	);
	LUT2 #(
		.INIT('h8)
	) name22 (
		\55(40)_pad ,
		_w156_,
		_w178_
	);
	LUT2 #(
		.INIT('h8)
	) name23 (
		\80(61)_pad ,
		_w158_,
		_w179_
	);
	LUT2 #(
		.INIT('h8)
	) name24 (
		\67(50)_pad ,
		_w160_,
		_w180_
	);
	LUT2 #(
		.INIT('h8)
	) name25 (
		\93(72)_pad ,
		_w162_,
		_w181_
	);
	LUT2 #(
		.INIT('h1)
	) name26 (
		_w178_,
		_w179_,
		_w182_
	);
	LUT2 #(
		.INIT('h1)
	) name27 (
		_w180_,
		_w181_,
		_w183_
	);
	LUT2 #(
		.INIT('h8)
	) name28 (
		_w182_,
		_w183_,
		_w184_
	);
	LUT2 #(
		.INIT('h2)
	) name29 (
		_w175_,
		_w184_,
		_w185_
	);
	LUT2 #(
		.INIT('h4)
	) name30 (
		_w175_,
		_w184_,
		_w186_
	);
	LUT2 #(
		.INIT('h1)
	) name31 (
		_w185_,
		_w186_,
		_w187_
	);
	LUT2 #(
		.INIT('h2)
	) name32 (
		_w177_,
		_w187_,
		_w188_
	);
	LUT2 #(
		.INIT('h4)
	) name33 (
		_w177_,
		_w187_,
		_w189_
	);
	LUT2 #(
		.INIT('h1)
	) name34 (
		_w188_,
		_w189_,
		_w190_
	);
	LUT2 #(
		.INIT('h2)
	) name35 (
		_w166_,
		_w168_,
		_w191_
	);
	LUT2 #(
		.INIT('h2)
	) name36 (
		\2104(220)_pad ,
		\2105(221)_pad ,
		_w192_
	);
	LUT2 #(
		.INIT('h8)
	) name37 (
		\100(77)_pad ,
		_w192_,
		_w193_
	);
	LUT2 #(
		.INIT('h8)
	) name38 (
		\2104(220)_pad ,
		\2105(221)_pad ,
		_w194_
	);
	LUT2 #(
		.INIT('h8)
	) name39 (
		\112(87)_pad ,
		_w194_,
		_w195_
	);
	LUT2 #(
		.INIT('h4)
	) name40 (
		\2104(220)_pad ,
		\2105(221)_pad ,
		_w196_
	);
	LUT2 #(
		.INIT('h8)
	) name41 (
		\124(97)_pad ,
		_w196_,
		_w197_
	);
	LUT2 #(
		.INIT('h1)
	) name42 (
		\2104(220)_pad ,
		\2105(221)_pad ,
		_w198_
	);
	LUT2 #(
		.INIT('h8)
	) name43 (
		\136(107)_pad ,
		_w198_,
		_w199_
	);
	LUT2 #(
		.INIT('h1)
	) name44 (
		_w193_,
		_w195_,
		_w200_
	);
	LUT2 #(
		.INIT('h1)
	) name45 (
		_w197_,
		_w199_,
		_w201_
	);
	LUT2 #(
		.INIT('h8)
	) name46 (
		_w200_,
		_w201_,
		_w202_
	);
	LUT2 #(
		.INIT('h2)
	) name47 (
		\29(22)_pad ,
		_w202_,
		_w203_
	);
	LUT2 #(
		.INIT('h4)
	) name48 (
		\29(22)_pad ,
		\35(26)_pad ,
		_w204_
	);
	LUT2 #(
		.INIT('h1)
	) name49 (
		_w203_,
		_w204_,
		_w205_
	);
	LUT2 #(
		.INIT('h1)
	) name50 (
		\2090(217)_pad ,
		_w205_,
		_w206_
	);
	LUT2 #(
		.INIT('h8)
	) name51 (
		\2090(217)_pad ,
		_w205_,
		_w207_
	);
	LUT2 #(
		.INIT('h1)
	) name52 (
		_w206_,
		_w207_,
		_w208_
	);
	LUT2 #(
		.INIT('h1)
	) name53 (
		\29(22)_pad ,
		\33(24)_pad ,
		_w209_
	);
	LUT2 #(
		.INIT('h8)
	) name54 (
		\103(80)_pad ,
		_w192_,
		_w210_
	);
	LUT2 #(
		.INIT('h8)
	) name55 (
		\115(90)_pad ,
		_w194_,
		_w211_
	);
	LUT2 #(
		.INIT('h8)
	) name56 (
		\127(100)_pad ,
		_w196_,
		_w212_
	);
	LUT2 #(
		.INIT('h8)
	) name57 (
		\139(110)_pad ,
		_w198_,
		_w213_
	);
	LUT2 #(
		.INIT('h1)
	) name58 (
		_w210_,
		_w211_,
		_w214_
	);
	LUT2 #(
		.INIT('h1)
	) name59 (
		_w212_,
		_w213_,
		_w215_
	);
	LUT2 #(
		.INIT('h8)
	) name60 (
		_w214_,
		_w215_,
		_w216_
	);
	LUT2 #(
		.INIT('h8)
	) name61 (
		\29(22)_pad ,
		_w216_,
		_w217_
	);
	LUT2 #(
		.INIT('h1)
	) name62 (
		_w209_,
		_w217_,
		_w218_
	);
	LUT2 #(
		.INIT('h1)
	) name63 (
		\2072(214)_pad ,
		_w218_,
		_w219_
	);
	LUT2 #(
		.INIT('h2)
	) name64 (
		\27(20)_pad ,
		\29(22)_pad ,
		_w220_
	);
	LUT2 #(
		.INIT('h8)
	) name65 (
		\102(79)_pad ,
		_w192_,
		_w221_
	);
	LUT2 #(
		.INIT('h8)
	) name66 (
		\114(89)_pad ,
		_w194_,
		_w222_
	);
	LUT2 #(
		.INIT('h8)
	) name67 (
		\126(99)_pad ,
		_w196_,
		_w223_
	);
	LUT2 #(
		.INIT('h8)
	) name68 (
		\138(109)_pad ,
		_w198_,
		_w224_
	);
	LUT2 #(
		.INIT('h1)
	) name69 (
		_w221_,
		_w222_,
		_w225_
	);
	LUT2 #(
		.INIT('h1)
	) name70 (
		_w223_,
		_w224_,
		_w226_
	);
	LUT2 #(
		.INIT('h8)
	) name71 (
		_w225_,
		_w226_,
		_w227_
	);
	LUT2 #(
		.INIT('h2)
	) name72 (
		\29(22)_pad ,
		_w227_,
		_w228_
	);
	LUT2 #(
		.INIT('h1)
	) name73 (
		_w220_,
		_w228_,
		_w229_
	);
	LUT2 #(
		.INIT('h4)
	) name74 (
		\2078(215)_pad ,
		_w229_,
		_w230_
	);
	LUT2 #(
		.INIT('h4)
	) name75 (
		\16(11)_pad ,
		\21(14)_pad ,
		_w231_
	);
	LUT2 #(
		.INIT('h8)
	) name76 (
		\51(36)_pad ,
		_w156_,
		_w232_
	);
	LUT2 #(
		.INIT('h8)
	) name77 (
		\76(57)_pad ,
		_w158_,
		_w233_
	);
	LUT2 #(
		.INIT('h8)
	) name78 (
		\63(46)_pad ,
		_w160_,
		_w234_
	);
	LUT2 #(
		.INIT('h8)
	) name79 (
		\89(68)_pad ,
		_w162_,
		_w235_
	);
	LUT2 #(
		.INIT('h1)
	) name80 (
		_w232_,
		_w233_,
		_w236_
	);
	LUT2 #(
		.INIT('h1)
	) name81 (
		_w234_,
		_w235_,
		_w237_
	);
	LUT2 #(
		.INIT('h8)
	) name82 (
		_w236_,
		_w237_,
		_w238_
	);
	LUT2 #(
		.INIT('h2)
	) name83 (
		\16(11)_pad ,
		_w238_,
		_w239_
	);
	LUT2 #(
		.INIT('h1)
	) name84 (
		_w231_,
		_w239_,
		_w240_
	);
	LUT2 #(
		.INIT('h4)
	) name85 (
		\1966(205)_pad ,
		_w240_,
		_w241_
	);
	LUT2 #(
		.INIT('h4)
	) name86 (
		\16(11)_pad ,
		\4(3)_pad ,
		_w242_
	);
	LUT2 #(
		.INIT('h2)
	) name87 (
		\16(11)_pad ,
		_w166_,
		_w243_
	);
	LUT2 #(
		.INIT('h1)
	) name88 (
		_w242_,
		_w243_,
		_w244_
	);
	LUT2 #(
		.INIT('h2)
	) name89 (
		\1348(201)_pad ,
		_w244_,
		_w245_
	);
	LUT2 #(
		.INIT('h8)
	) name90 (
		\48(33)_pad ,
		_w156_,
		_w246_
	);
	LUT2 #(
		.INIT('h8)
	) name91 (
		\73(54)_pad ,
		_w158_,
		_w247_
	);
	LUT2 #(
		.INIT('h8)
	) name92 (
		\61(44)_pad ,
		_w160_,
		_w248_
	);
	LUT2 #(
		.INIT('h8)
	) name93 (
		\86(65)_pad ,
		_w162_,
		_w249_
	);
	LUT2 #(
		.INIT('h1)
	) name94 (
		_w246_,
		_w247_,
		_w250_
	);
	LUT2 #(
		.INIT('h1)
	) name95 (
		_w248_,
		_w249_,
		_w251_
	);
	LUT2 #(
		.INIT('h8)
	) name96 (
		_w250_,
		_w251_,
		_w252_
	);
	LUT2 #(
		.INIT('h2)
	) name97 (
		\16(11)_pad ,
		_w252_,
		_w253_
	);
	LUT2 #(
		.INIT('h4)
	) name98 (
		\16(11)_pad ,
		\6(5)_pad ,
		_w254_
	);
	LUT2 #(
		.INIT('h1)
	) name99 (
		_w253_,
		_w254_,
		_w255_
	);
	LUT2 #(
		.INIT('h1)
	) name100 (
		\1981(208)_pad ,
		_w255_,
		_w256_
	);
	LUT2 #(
		.INIT('h8)
	) name101 (
		\1981(208)_pad ,
		_w255_,
		_w257_
	);
	LUT2 #(
		.INIT('h1)
	) name102 (
		_w256_,
		_w257_,
		_w258_
	);
	LUT2 #(
		.INIT('h8)
	) name103 (
		\99(76)_pad ,
		_w192_,
		_w259_
	);
	LUT2 #(
		.INIT('h8)
	) name104 (
		\111(86)_pad ,
		_w194_,
		_w260_
	);
	LUT2 #(
		.INIT('h8)
	) name105 (
		\123(96)_pad ,
		_w196_,
		_w261_
	);
	LUT2 #(
		.INIT('h8)
	) name106 (
		\135(106)_pad ,
		_w198_,
		_w262_
	);
	LUT2 #(
		.INIT('h1)
	) name107 (
		_w259_,
		_w260_,
		_w263_
	);
	LUT2 #(
		.INIT('h1)
	) name108 (
		_w261_,
		_w262_,
		_w264_
	);
	LUT2 #(
		.INIT('h8)
	) name109 (
		_w263_,
		_w264_,
		_w265_
	);
	LUT2 #(
		.INIT('h8)
	) name110 (
		\29(22)_pad ,
		_w265_,
		_w266_
	);
	LUT2 #(
		.INIT('h4)
	) name111 (
		\16(11)_pad ,
		\24(17)_pad ,
		_w267_
	);
	LUT2 #(
		.INIT('h8)
	) name112 (
		\47(32)_pad ,
		_w156_,
		_w268_
	);
	LUT2 #(
		.INIT('h8)
	) name113 (
		\72(53)_pad ,
		_w158_,
		_w269_
	);
	LUT2 #(
		.INIT('h8)
	) name114 (
		\60(43)_pad ,
		_w160_,
		_w270_
	);
	LUT2 #(
		.INIT('h8)
	) name115 (
		\85(64)_pad ,
		_w162_,
		_w271_
	);
	LUT2 #(
		.INIT('h1)
	) name116 (
		_w268_,
		_w269_,
		_w272_
	);
	LUT2 #(
		.INIT('h1)
	) name117 (
		_w270_,
		_w271_,
		_w273_
	);
	LUT2 #(
		.INIT('h8)
	) name118 (
		_w272_,
		_w273_,
		_w274_
	);
	LUT2 #(
		.INIT('h2)
	) name119 (
		\16(11)_pad ,
		_w274_,
		_w275_
	);
	LUT2 #(
		.INIT('h1)
	) name120 (
		_w267_,
		_w275_,
		_w276_
	);
	LUT2 #(
		.INIT('h4)
	) name121 (
		\1986(209)_pad ,
		_w276_,
		_w277_
	);
	LUT2 #(
		.INIT('h1)
	) name122 (
		\28(21)_pad ,
		\29(22)_pad ,
		_w278_
	);
	LUT2 #(
		.INIT('h4)
	) name123 (
		\1348(201)_pad ,
		_w244_,
		_w279_
	);
	LUT2 #(
		.INIT('h2)
	) name124 (
		\1986(209)_pad ,
		_w276_,
		_w280_
	);
	LUT2 #(
		.INIT('h2)
	) name125 (
		\25(18)_pad ,
		\29(22)_pad ,
		_w281_
	);
	LUT2 #(
		.INIT('h8)
	) name126 (
		\95(74)_pad ,
		_w192_,
		_w282_
	);
	LUT2 #(
		.INIT('h8)
	) name127 (
		\107(84)_pad ,
		_w194_,
		_w283_
	);
	LUT2 #(
		.INIT('h8)
	) name128 (
		\119(94)_pad ,
		_w196_,
		_w284_
	);
	LUT2 #(
		.INIT('h8)
	) name129 (
		\131(104)_pad ,
		_w198_,
		_w285_
	);
	LUT2 #(
		.INIT('h1)
	) name130 (
		_w282_,
		_w283_,
		_w286_
	);
	LUT2 #(
		.INIT('h1)
	) name131 (
		_w284_,
		_w285_,
		_w287_
	);
	LUT2 #(
		.INIT('h8)
	) name132 (
		_w286_,
		_w287_,
		_w288_
	);
	LUT2 #(
		.INIT('h2)
	) name133 (
		\29(22)_pad ,
		_w288_,
		_w289_
	);
	LUT2 #(
		.INIT('h1)
	) name134 (
		_w281_,
		_w289_,
		_w290_
	);
	LUT2 #(
		.INIT('h2)
	) name135 (
		\1991(210)_pad ,
		_w290_,
		_w291_
	);
	LUT2 #(
		.INIT('h1)
	) name136 (
		\29(22)_pad ,
		\34(25)_pad ,
		_w292_
	);
	LUT2 #(
		.INIT('h8)
	) name137 (
		\101(78)_pad ,
		_w192_,
		_w293_
	);
	LUT2 #(
		.INIT('h8)
	) name138 (
		\113(88)_pad ,
		_w194_,
		_w294_
	);
	LUT2 #(
		.INIT('h8)
	) name139 (
		\125(98)_pad ,
		_w196_,
		_w295_
	);
	LUT2 #(
		.INIT('h8)
	) name140 (
		\137(108)_pad ,
		_w198_,
		_w296_
	);
	LUT2 #(
		.INIT('h1)
	) name141 (
		_w293_,
		_w294_,
		_w297_
	);
	LUT2 #(
		.INIT('h1)
	) name142 (
		_w295_,
		_w296_,
		_w298_
	);
	LUT2 #(
		.INIT('h8)
	) name143 (
		_w297_,
		_w298_,
		_w299_
	);
	LUT2 #(
		.INIT('h8)
	) name144 (
		\29(22)_pad ,
		_w299_,
		_w300_
	);
	LUT2 #(
		.INIT('h1)
	) name145 (
		_w292_,
		_w300_,
		_w301_
	);
	LUT2 #(
		.INIT('h8)
	) name146 (
		\2084(216)_pad ,
		_w301_,
		_w302_
	);
	LUT2 #(
		.INIT('h4)
	) name147 (
		\16(11)_pad ,
		\20(13)_pad ,
		_w303_
	);
	LUT2 #(
		.INIT('h8)
	) name148 (
		\53(38)_pad ,
		_w156_,
		_w304_
	);
	LUT2 #(
		.INIT('h8)
	) name149 (
		\78(59)_pad ,
		_w158_,
		_w305_
	);
	LUT2 #(
		.INIT('h8)
	) name150 (
		\65(48)_pad ,
		_w160_,
		_w306_
	);
	LUT2 #(
		.INIT('h8)
	) name151 (
		\91(70)_pad ,
		_w162_,
		_w307_
	);
	LUT2 #(
		.INIT('h1)
	) name152 (
		_w304_,
		_w305_,
		_w308_
	);
	LUT2 #(
		.INIT('h1)
	) name153 (
		_w306_,
		_w307_,
		_w309_
	);
	LUT2 #(
		.INIT('h8)
	) name154 (
		_w308_,
		_w309_,
		_w310_
	);
	LUT2 #(
		.INIT('h2)
	) name155 (
		\16(11)_pad ,
		_w310_,
		_w311_
	);
	LUT2 #(
		.INIT('h1)
	) name156 (
		_w303_,
		_w311_,
		_w312_
	);
	LUT2 #(
		.INIT('h4)
	) name157 (
		\1956(203)_pad ,
		_w312_,
		_w313_
	);
	LUT2 #(
		.INIT('h2)
	) name158 (
		\1956(203)_pad ,
		_w312_,
		_w314_
	);
	LUT2 #(
		.INIT('h1)
	) name159 (
		\2084(216)_pad ,
		_w301_,
		_w315_
	);
	LUT2 #(
		.INIT('h1)
	) name160 (
		\26(19)_pad ,
		\29(22)_pad ,
		_w316_
	);
	LUT2 #(
		.INIT('h8)
	) name161 (
		\104(81)_pad ,
		_w192_,
		_w317_
	);
	LUT2 #(
		.INIT('h8)
	) name162 (
		\116(91)_pad ,
		_w194_,
		_w318_
	);
	LUT2 #(
		.INIT('h8)
	) name163 (
		\128(101)_pad ,
		_w196_,
		_w319_
	);
	LUT2 #(
		.INIT('h8)
	) name164 (
		\140(111)_pad ,
		_w198_,
		_w320_
	);
	LUT2 #(
		.INIT('h1)
	) name165 (
		_w317_,
		_w318_,
		_w321_
	);
	LUT2 #(
		.INIT('h1)
	) name166 (
		_w319_,
		_w320_,
		_w322_
	);
	LUT2 #(
		.INIT('h8)
	) name167 (
		_w321_,
		_w322_,
		_w323_
	);
	LUT2 #(
		.INIT('h8)
	) name168 (
		\29(22)_pad ,
		_w323_,
		_w324_
	);
	LUT2 #(
		.INIT('h1)
	) name169 (
		_w316_,
		_w324_,
		_w325_
	);
	LUT2 #(
		.INIT('h8)
	) name170 (
		\2067(213)_pad ,
		_w325_,
		_w326_
	);
	LUT2 #(
		.INIT('h4)
	) name171 (
		\1991(210)_pad ,
		_w290_,
		_w327_
	);
	LUT2 #(
		.INIT('h1)
	) name172 (
		\29(22)_pad ,
		\32(23)_pad ,
		_w328_
	);
	LUT2 #(
		.INIT('h8)
	) name173 (
		\105(82)_pad ,
		_w192_,
		_w329_
	);
	LUT2 #(
		.INIT('h8)
	) name174 (
		\117(92)_pad ,
		_w194_,
		_w330_
	);
	LUT2 #(
		.INIT('h8)
	) name175 (
		\129(102)_pad ,
		_w196_,
		_w331_
	);
	LUT2 #(
		.INIT('h8)
	) name176 (
		\141(112)_pad ,
		_w198_,
		_w332_
	);
	LUT2 #(
		.INIT('h1)
	) name177 (
		_w329_,
		_w330_,
		_w333_
	);
	LUT2 #(
		.INIT('h1)
	) name178 (
		_w331_,
		_w332_,
		_w334_
	);
	LUT2 #(
		.INIT('h8)
	) name179 (
		_w333_,
		_w334_,
		_w335_
	);
	LUT2 #(
		.INIT('h8)
	) name180 (
		\29(22)_pad ,
		_w335_,
		_w336_
	);
	LUT2 #(
		.INIT('h1)
	) name181 (
		_w328_,
		_w336_,
		_w337_
	);
	LUT2 #(
		.INIT('h1)
	) name182 (
		\1996(211)_pad ,
		_w337_,
		_w338_
	);
	LUT2 #(
		.INIT('h1)
	) name183 (
		\16(11)_pad ,
		\23(16)_pad ,
		_w339_
	);
	LUT2 #(
		.INIT('h8)
	) name184 (
		\87(66)_pad ,
		_w162_,
		_w340_
	);
	LUT2 #(
		.INIT('h8)
	) name185 (
		\74(55)_pad ,
		_w158_,
		_w341_
	);
	LUT2 #(
		.INIT('h8)
	) name186 (
		\49(34)_pad ,
		_w156_,
		_w342_
	);
	LUT2 #(
		.INIT('h1)
	) name187 (
		_w160_,
		_w340_,
		_w343_
	);
	LUT2 #(
		.INIT('h1)
	) name188 (
		_w341_,
		_w342_,
		_w344_
	);
	LUT2 #(
		.INIT('h8)
	) name189 (
		_w343_,
		_w344_,
		_w345_
	);
	LUT2 #(
		.INIT('h8)
	) name190 (
		\16(11)_pad ,
		_w345_,
		_w346_
	);
	LUT2 #(
		.INIT('h1)
	) name191 (
		_w339_,
		_w346_,
		_w347_
	);
	LUT2 #(
		.INIT('h8)
	) name192 (
		\1976(207)_pad ,
		_w347_,
		_w348_
	);
	LUT2 #(
		.INIT('h2)
	) name193 (
		\2078(215)_pad ,
		_w229_,
		_w349_
	);
	LUT2 #(
		.INIT('h1)
	) name194 (
		\16(11)_pad ,
		\22(15)_pad ,
		_w350_
	);
	LUT2 #(
		.INIT('h8)
	) name195 (
		\50(35)_pad ,
		_w156_,
		_w351_
	);
	LUT2 #(
		.INIT('h8)
	) name196 (
		\75(56)_pad ,
		_w158_,
		_w352_
	);
	LUT2 #(
		.INIT('h8)
	) name197 (
		\62(45)_pad ,
		_w160_,
		_w353_
	);
	LUT2 #(
		.INIT('h8)
	) name198 (
		\88(67)_pad ,
		_w162_,
		_w354_
	);
	LUT2 #(
		.INIT('h1)
	) name199 (
		_w351_,
		_w352_,
		_w355_
	);
	LUT2 #(
		.INIT('h1)
	) name200 (
		_w353_,
		_w354_,
		_w356_
	);
	LUT2 #(
		.INIT('h8)
	) name201 (
		_w355_,
		_w356_,
		_w357_
	);
	LUT2 #(
		.INIT('h8)
	) name202 (
		\16(11)_pad ,
		_w357_,
		_w358_
	);
	LUT2 #(
		.INIT('h1)
	) name203 (
		_w350_,
		_w358_,
		_w359_
	);
	LUT2 #(
		.INIT('h8)
	) name204 (
		\1971(206)_pad ,
		_w359_,
		_w360_
	);
	LUT2 #(
		.INIT('h8)
	) name205 (
		\1996(211)_pad ,
		_w337_,
		_w361_
	);
	LUT2 #(
		.INIT('h8)
	) name206 (
		\2072(214)_pad ,
		_w218_,
		_w362_
	);
	LUT2 #(
		.INIT('h1)
	) name207 (
		\2067(213)_pad ,
		_w325_,
		_w363_
	);
	LUT2 #(
		.INIT('h1)
	) name208 (
		\1971(206)_pad ,
		_w359_,
		_w364_
	);
	LUT2 #(
		.INIT('h2)
	) name209 (
		\1966(205)_pad ,
		_w240_,
		_w365_
	);
	LUT2 #(
		.INIT('h4)
	) name210 (
		\16(11)_pad ,
		\5(4)_pad ,
		_w366_
	);
	LUT2 #(
		.INIT('h8)
	) name211 (
		\52(37)_pad ,
		_w156_,
		_w367_
	);
	LUT2 #(
		.INIT('h8)
	) name212 (
		\77(58)_pad ,
		_w158_,
		_w368_
	);
	LUT2 #(
		.INIT('h8)
	) name213 (
		\64(47)_pad ,
		_w160_,
		_w369_
	);
	LUT2 #(
		.INIT('h8)
	) name214 (
		\90(69)_pad ,
		_w162_,
		_w370_
	);
	LUT2 #(
		.INIT('h1)
	) name215 (
		_w367_,
		_w368_,
		_w371_
	);
	LUT2 #(
		.INIT('h1)
	) name216 (
		_w369_,
		_w370_,
		_w372_
	);
	LUT2 #(
		.INIT('h8)
	) name217 (
		_w371_,
		_w372_,
		_w373_
	);
	LUT2 #(
		.INIT('h2)
	) name218 (
		\16(11)_pad ,
		_w373_,
		_w374_
	);
	LUT2 #(
		.INIT('h1)
	) name219 (
		_w366_,
		_w374_,
		_w375_
	);
	LUT2 #(
		.INIT('h4)
	) name220 (
		\1961(204)_pad ,
		_w375_,
		_w376_
	);
	LUT2 #(
		.INIT('h2)
	) name221 (
		\1961(204)_pad ,
		_w375_,
		_w377_
	);
	LUT2 #(
		.INIT('h1)
	) name222 (
		\1976(207)_pad ,
		_w347_,
		_w378_
	);
	LUT2 #(
		.INIT('h2)
	) name223 (
		\16(11)_pad ,
		_w175_,
		_w379_
	);
	LUT2 #(
		.INIT('h4)
	) name224 (
		\16(11)_pad ,
		\19(12)_pad ,
		_w380_
	);
	LUT2 #(
		.INIT('h1)
	) name225 (
		_w379_,
		_w380_,
		_w381_
	);
	LUT2 #(
		.INIT('h2)
	) name226 (
		\1341(200)_pad ,
		_w381_,
		_w382_
	);
	LUT2 #(
		.INIT('h4)
	) name227 (
		\1341(200)_pad ,
		_w381_,
		_w383_
	);
	LUT2 #(
		.INIT('h2)
	) name228 (
		\11(8)_pad ,
		_w278_,
		_w384_
	);
	LUT2 #(
		.INIT('h4)
	) name229 (
		_w266_,
		_w384_,
		_w385_
	);
	LUT2 #(
		.INIT('h4)
	) name230 (
		_w219_,
		_w385_,
		_w386_
	);
	LUT2 #(
		.INIT('h1)
	) name231 (
		_w230_,
		_w241_,
		_w387_
	);
	LUT2 #(
		.INIT('h1)
	) name232 (
		_w245_,
		_w277_,
		_w388_
	);
	LUT2 #(
		.INIT('h1)
	) name233 (
		_w279_,
		_w280_,
		_w389_
	);
	LUT2 #(
		.INIT('h1)
	) name234 (
		_w291_,
		_w302_,
		_w390_
	);
	LUT2 #(
		.INIT('h1)
	) name235 (
		_w313_,
		_w314_,
		_w391_
	);
	LUT2 #(
		.INIT('h1)
	) name236 (
		_w315_,
		_w326_,
		_w392_
	);
	LUT2 #(
		.INIT('h1)
	) name237 (
		_w327_,
		_w338_,
		_w393_
	);
	LUT2 #(
		.INIT('h1)
	) name238 (
		_w348_,
		_w349_,
		_w394_
	);
	LUT2 #(
		.INIT('h1)
	) name239 (
		_w360_,
		_w361_,
		_w395_
	);
	LUT2 #(
		.INIT('h1)
	) name240 (
		_w362_,
		_w363_,
		_w396_
	);
	LUT2 #(
		.INIT('h1)
	) name241 (
		_w364_,
		_w365_,
		_w397_
	);
	LUT2 #(
		.INIT('h1)
	) name242 (
		_w376_,
		_w377_,
		_w398_
	);
	LUT2 #(
		.INIT('h1)
	) name243 (
		_w378_,
		_w382_,
		_w399_
	);
	LUT2 #(
		.INIT('h4)
	) name244 (
		_w383_,
		_w399_,
		_w400_
	);
	LUT2 #(
		.INIT('h8)
	) name245 (
		_w397_,
		_w398_,
		_w401_
	);
	LUT2 #(
		.INIT('h8)
	) name246 (
		_w395_,
		_w396_,
		_w402_
	);
	LUT2 #(
		.INIT('h8)
	) name247 (
		_w393_,
		_w394_,
		_w403_
	);
	LUT2 #(
		.INIT('h8)
	) name248 (
		_w391_,
		_w392_,
		_w404_
	);
	LUT2 #(
		.INIT('h8)
	) name249 (
		_w389_,
		_w390_,
		_w405_
	);
	LUT2 #(
		.INIT('h8)
	) name250 (
		_w387_,
		_w388_,
		_w406_
	);
	LUT2 #(
		.INIT('h4)
	) name251 (
		_w208_,
		_w386_,
		_w407_
	);
	LUT2 #(
		.INIT('h4)
	) name252 (
		_w258_,
		_w407_,
		_w408_
	);
	LUT2 #(
		.INIT('h8)
	) name253 (
		_w405_,
		_w406_,
		_w409_
	);
	LUT2 #(
		.INIT('h8)
	) name254 (
		_w403_,
		_w404_,
		_w410_
	);
	LUT2 #(
		.INIT('h8)
	) name255 (
		_w401_,
		_w402_,
		_w411_
	);
	LUT2 #(
		.INIT('h8)
	) name256 (
		_w400_,
		_w411_,
		_w412_
	);
	LUT2 #(
		.INIT('h8)
	) name257 (
		_w409_,
		_w410_,
		_w413_
	);
	LUT2 #(
		.INIT('h8)
	) name258 (
		_w408_,
		_w413_,
		_w414_
	);
	LUT2 #(
		.INIT('h8)
	) name259 (
		_w412_,
		_w414_,
		_w415_
	);
	LUT2 #(
		.INIT('h2)
	) name260 (
		\2096(218)_pad ,
		_w265_,
		_w416_
	);
	LUT2 #(
		.INIT('h4)
	) name261 (
		\2096(218)_pad ,
		_w265_,
		_w417_
	);
	LUT2 #(
		.INIT('h1)
	) name262 (
		\2100(219)_pad ,
		_w416_,
		_w418_
	);
	LUT2 #(
		.INIT('h4)
	) name263 (
		_w417_,
		_w418_,
		_w419_
	);
	LUT2 #(
		.INIT('h8)
	) name264 (
		\2072(214)_pad ,
		\2078(215)_pad ,
		_w420_
	);
	LUT2 #(
		.INIT('h8)
	) name265 (
		\2084(216)_pad ,
		\2090(217)_pad ,
		_w421_
	);
	LUT2 #(
		.INIT('h8)
	) name266 (
		_w420_,
		_w421_,
		_w422_
	);
	LUT2 #(
		.INIT('h8)
	) name267 (
		\409(298)_pad ,
		\94(73)_pad ,
		_w423_
	);
	LUT2 #(
		.INIT('h8)
	) name268 (
		\108(85)_pad ,
		\120(95)_pad ,
		_w424_
	);
	LUT2 #(
		.INIT('h8)
	) name269 (
		\57(42)_pad ,
		\69(52)_pad ,
		_w425_
	);
	LUT2 #(
		.INIT('h8)
	) name270 (
		_w424_,
		_w425_,
		_w426_
	);
	LUT2 #(
		.INIT('h2)
	) name271 (
		\567(194)_pad ,
		_w426_,
		_w427_
	);
	LUT2 #(
		.INIT('h8)
	) name272 (
		\132(105)_pad ,
		\44(31)_pad ,
		_w428_
	);
	LUT2 #(
		.INIT('h8)
	) name273 (
		\82(63)_pad ,
		\96(75)_pad ,
		_w429_
	);
	LUT2 #(
		.INIT('h8)
	) name274 (
		_w428_,
		_w429_,
		_w430_
	);
	LUT2 #(
		.INIT('h2)
	) name275 (
		\2106(222)_pad ,
		_w430_,
		_w431_
	);
	LUT2 #(
		.INIT('h1)
	) name276 (
		_w427_,
		_w431_,
		_w432_
	);
	LUT2 #(
		.INIT('h8)
	) name277 (
		\483(191)_pad ,
		\661(196)_pad ,
		_w433_
	);
	LUT2 #(
		.INIT('h8)
	) name278 (
		\36(27)_pad ,
		_w433_,
		_w434_
	);
	LUT2 #(
		.INIT('h8)
	) name279 (
		_w432_,
		_w434_,
		_w435_
	);
	LUT2 #(
		.INIT('h8)
	) name280 (
		\1(0)_pad ,
		\3(2)_pad ,
		_w436_
	);
	LUT2 #(
		.INIT('h2)
	) name281 (
		_w433_,
		_w436_,
		_w437_
	);
	LUT2 #(
		.INIT('h8)
	) name282 (
		_w432_,
		_w437_,
		_w438_
	);
	LUT2 #(
		.INIT('h8)
	) name283 (
		\661(196)_pad ,
		\7(6)_pad ,
		_w439_
	);
	LUT2 #(
		.INIT('h8)
	) name284 (
		\2106(222)_pad ,
		_w439_,
		_w440_
	);
	LUT2 #(
		.INIT('h2)
	) name285 (
		_w310_,
		_w357_,
		_w441_
	);
	LUT2 #(
		.INIT('h4)
	) name286 (
		_w310_,
		_w357_,
		_w442_
	);
	LUT2 #(
		.INIT('h1)
	) name287 (
		_w441_,
		_w442_,
		_w443_
	);
	LUT2 #(
		.INIT('h2)
	) name288 (
		_w187_,
		_w252_,
		_w444_
	);
	LUT2 #(
		.INIT('h4)
	) name289 (
		_w187_,
		_w252_,
		_w445_
	);
	LUT2 #(
		.INIT('h1)
	) name290 (
		_w444_,
		_w445_,
		_w446_
	);
	LUT2 #(
		.INIT('h8)
	) name291 (
		_w274_,
		_w446_,
		_w447_
	);
	LUT2 #(
		.INIT('h1)
	) name292 (
		_w274_,
		_w446_,
		_w448_
	);
	LUT2 #(
		.INIT('h1)
	) name293 (
		_w447_,
		_w448_,
		_w449_
	);
	LUT2 #(
		.INIT('h2)
	) name294 (
		_w345_,
		_w449_,
		_w450_
	);
	LUT2 #(
		.INIT('h4)
	) name295 (
		_w345_,
		_w449_,
		_w451_
	);
	LUT2 #(
		.INIT('h1)
	) name296 (
		_w450_,
		_w451_,
		_w452_
	);
	LUT2 #(
		.INIT('h8)
	) name297 (
		_w443_,
		_w452_,
		_w453_
	);
	LUT2 #(
		.INIT('h1)
	) name298 (
		_w443_,
		_w452_,
		_w454_
	);
	LUT2 #(
		.INIT('h1)
	) name299 (
		_w453_,
		_w454_,
		_w455_
	);
	LUT2 #(
		.INIT('h2)
	) name300 (
		_w166_,
		_w373_,
		_w456_
	);
	LUT2 #(
		.INIT('h4)
	) name301 (
		_w166_,
		_w373_,
		_w457_
	);
	LUT2 #(
		.INIT('h1)
	) name302 (
		_w456_,
		_w457_,
		_w458_
	);
	LUT2 #(
		.INIT('h8)
	) name303 (
		_w238_,
		_w458_,
		_w459_
	);
	LUT2 #(
		.INIT('h1)
	) name304 (
		_w238_,
		_w458_,
		_w460_
	);
	LUT2 #(
		.INIT('h1)
	) name305 (
		_w459_,
		_w460_,
		_w461_
	);
	LUT2 #(
		.INIT('h8)
	) name306 (
		_w455_,
		_w461_,
		_w462_
	);
	LUT2 #(
		.INIT('h1)
	) name307 (
		_w455_,
		_w461_,
		_w463_
	);
	LUT2 #(
		.INIT('h1)
	) name308 (
		\37(28)_pad ,
		_w462_,
		_w464_
	);
	LUT2 #(
		.INIT('h4)
	) name309 (
		_w463_,
		_w464_,
		_w465_
	);
	LUT2 #(
		.INIT('h2)
	) name310 (
		\1341(200)_pad ,
		\1348(201)_pad ,
		_w466_
	);
	LUT2 #(
		.INIT('h4)
	) name311 (
		\1341(200)_pad ,
		\1348(201)_pad ,
		_w467_
	);
	LUT2 #(
		.INIT('h1)
	) name312 (
		_w466_,
		_w467_,
		_w468_
	);
	LUT2 #(
		.INIT('h1)
	) name313 (
		\2435(225)_pad ,
		\2438(226)_pad ,
		_w469_
	);
	LUT2 #(
		.INIT('h8)
	) name314 (
		\2435(225)_pad ,
		\2438(226)_pad ,
		_w470_
	);
	LUT2 #(
		.INIT('h1)
	) name315 (
		_w469_,
		_w470_,
		_w471_
	);
	LUT2 #(
		.INIT('h2)
	) name316 (
		_w468_,
		_w471_,
		_w472_
	);
	LUT2 #(
		.INIT('h4)
	) name317 (
		_w468_,
		_w471_,
		_w473_
	);
	LUT2 #(
		.INIT('h1)
	) name318 (
		_w472_,
		_w473_,
		_w474_
	);
	LUT2 #(
		.INIT('h1)
	) name319 (
		\2446(228)_pad ,
		\2454(230)_pad ,
		_w475_
	);
	LUT2 #(
		.INIT('h8)
	) name320 (
		\2446(228)_pad ,
		\2454(230)_pad ,
		_w476_
	);
	LUT2 #(
		.INIT('h1)
	) name321 (
		_w475_,
		_w476_,
		_w477_
	);
	LUT2 #(
		.INIT('h1)
	) name322 (
		\2427(223)_pad ,
		\2430(224)_pad ,
		_w478_
	);
	LUT2 #(
		.INIT('h8)
	) name323 (
		\2427(223)_pad ,
		\2430(224)_pad ,
		_w479_
	);
	LUT2 #(
		.INIT('h1)
	) name324 (
		_w478_,
		_w479_,
		_w480_
	);
	LUT2 #(
		.INIT('h2)
	) name325 (
		\2443(227)_pad ,
		\2451(229)_pad ,
		_w481_
	);
	LUT2 #(
		.INIT('h4)
	) name326 (
		\2443(227)_pad ,
		\2451(229)_pad ,
		_w482_
	);
	LUT2 #(
		.INIT('h1)
	) name327 (
		_w481_,
		_w482_,
		_w483_
	);
	LUT2 #(
		.INIT('h2)
	) name328 (
		_w480_,
		_w483_,
		_w484_
	);
	LUT2 #(
		.INIT('h4)
	) name329 (
		_w480_,
		_w483_,
		_w485_
	);
	LUT2 #(
		.INIT('h1)
	) name330 (
		_w484_,
		_w485_,
		_w486_
	);
	LUT2 #(
		.INIT('h4)
	) name331 (
		_w477_,
		_w486_,
		_w487_
	);
	LUT2 #(
		.INIT('h2)
	) name332 (
		_w477_,
		_w486_,
		_w488_
	);
	LUT2 #(
		.INIT('h1)
	) name333 (
		_w487_,
		_w488_,
		_w489_
	);
	LUT2 #(
		.INIT('h8)
	) name334 (
		_w474_,
		_w489_,
		_w490_
	);
	LUT2 #(
		.INIT('h1)
	) name335 (
		_w474_,
		_w489_,
		_w491_
	);
	LUT2 #(
		.INIT('h2)
	) name336 (
		\14(9)_pad ,
		_w490_,
		_w492_
	);
	LUT2 #(
		.INIT('h4)
	) name337 (
		_w491_,
		_w492_,
		_w493_
	);
	LUT2 #(
		.INIT('h4)
	) name338 (
		_w202_,
		_w265_,
		_w494_
	);
	LUT2 #(
		.INIT('h2)
	) name339 (
		_w202_,
		_w265_,
		_w495_
	);
	LUT2 #(
		.INIT('h1)
	) name340 (
		_w494_,
		_w495_,
		_w496_
	);
	LUT2 #(
		.INIT('h8)
	) name341 (
		_w299_,
		_w496_,
		_w497_
	);
	LUT2 #(
		.INIT('h1)
	) name342 (
		_w299_,
		_w496_,
		_w498_
	);
	LUT2 #(
		.INIT('h1)
	) name343 (
		_w497_,
		_w498_,
		_w499_
	);
	LUT2 #(
		.INIT('h8)
	) name344 (
		\106(83)_pad ,
		_w192_,
		_w500_
	);
	LUT2 #(
		.INIT('h8)
	) name345 (
		\118(93)_pad ,
		_w194_,
		_w501_
	);
	LUT2 #(
		.INIT('h8)
	) name346 (
		\130(103)_pad ,
		_w196_,
		_w502_
	);
	LUT2 #(
		.INIT('h8)
	) name347 (
		\142(113)_pad ,
		_w198_,
		_w503_
	);
	LUT2 #(
		.INIT('h1)
	) name348 (
		_w500_,
		_w501_,
		_w504_
	);
	LUT2 #(
		.INIT('h1)
	) name349 (
		_w502_,
		_w503_,
		_w505_
	);
	LUT2 #(
		.INIT('h8)
	) name350 (
		_w504_,
		_w505_,
		_w506_
	);
	LUT2 #(
		.INIT('h2)
	) name351 (
		_w227_,
		_w506_,
		_w507_
	);
	LUT2 #(
		.INIT('h4)
	) name352 (
		_w227_,
		_w506_,
		_w508_
	);
	LUT2 #(
		.INIT('h1)
	) name353 (
		_w507_,
		_w508_,
		_w509_
	);
	LUT2 #(
		.INIT('h2)
	) name354 (
		_w323_,
		_w335_,
		_w510_
	);
	LUT2 #(
		.INIT('h4)
	) name355 (
		_w323_,
		_w335_,
		_w511_
	);
	LUT2 #(
		.INIT('h1)
	) name356 (
		_w510_,
		_w511_,
		_w512_
	);
	LUT2 #(
		.INIT('h8)
	) name357 (
		_w216_,
		_w512_,
		_w513_
	);
	LUT2 #(
		.INIT('h1)
	) name358 (
		_w216_,
		_w512_,
		_w514_
	);
	LUT2 #(
		.INIT('h1)
	) name359 (
		_w513_,
		_w514_,
		_w515_
	);
	LUT2 #(
		.INIT('h2)
	) name360 (
		_w288_,
		_w515_,
		_w516_
	);
	LUT2 #(
		.INIT('h4)
	) name361 (
		_w288_,
		_w515_,
		_w517_
	);
	LUT2 #(
		.INIT('h1)
	) name362 (
		_w516_,
		_w517_,
		_w518_
	);
	LUT2 #(
		.INIT('h8)
	) name363 (
		_w509_,
		_w518_,
		_w519_
	);
	LUT2 #(
		.INIT('h1)
	) name364 (
		_w509_,
		_w518_,
		_w520_
	);
	LUT2 #(
		.INIT('h1)
	) name365 (
		_w519_,
		_w520_,
		_w521_
	);
	LUT2 #(
		.INIT('h4)
	) name366 (
		_w499_,
		_w521_,
		_w522_
	);
	LUT2 #(
		.INIT('h2)
	) name367 (
		_w499_,
		_w521_,
		_w523_
	);
	LUT2 #(
		.INIT('h1)
	) name368 (
		\37(28)_pad ,
		_w522_,
		_w524_
	);
	LUT2 #(
		.INIT('h4)
	) name369 (
		_w523_,
		_w524_,
		_w525_
	);
	LUT2 #(
		.INIT('h1)
	) name370 (
		\2072(214)_pad ,
		\2078(215)_pad ,
		_w526_
	);
	LUT2 #(
		.INIT('h1)
	) name371 (
		_w420_,
		_w526_,
		_w527_
	);
	LUT2 #(
		.INIT('h2)
	) name372 (
		\2096(218)_pad ,
		_w527_,
		_w528_
	);
	LUT2 #(
		.INIT('h4)
	) name373 (
		\2096(218)_pad ,
		_w527_,
		_w529_
	);
	LUT2 #(
		.INIT('h1)
	) name374 (
		_w528_,
		_w529_,
		_w530_
	);
	LUT2 #(
		.INIT('h2)
	) name375 (
		\2084(216)_pad ,
		_w530_,
		_w531_
	);
	LUT2 #(
		.INIT('h4)
	) name376 (
		\2084(216)_pad ,
		_w530_,
		_w532_
	);
	LUT2 #(
		.INIT('h1)
	) name377 (
		_w531_,
		_w532_,
		_w533_
	);
	LUT2 #(
		.INIT('h1)
	) name378 (
		\2090(217)_pad ,
		\2678(232)_pad ,
		_w534_
	);
	LUT2 #(
		.INIT('h8)
	) name379 (
		\2090(217)_pad ,
		\2678(232)_pad ,
		_w535_
	);
	LUT2 #(
		.INIT('h1)
	) name380 (
		_w534_,
		_w535_,
		_w536_
	);
	LUT2 #(
		.INIT('h8)
	) name381 (
		\2067(213)_pad ,
		_w536_,
		_w537_
	);
	LUT2 #(
		.INIT('h1)
	) name382 (
		\2067(213)_pad ,
		_w536_,
		_w538_
	);
	LUT2 #(
		.INIT('h1)
	) name383 (
		_w537_,
		_w538_,
		_w539_
	);
	LUT2 #(
		.INIT('h2)
	) name384 (
		\2100(219)_pad ,
		_w539_,
		_w540_
	);
	LUT2 #(
		.INIT('h4)
	) name385 (
		\2100(219)_pad ,
		_w539_,
		_w541_
	);
	LUT2 #(
		.INIT('h1)
	) name386 (
		_w540_,
		_w541_,
		_w542_
	);
	LUT2 #(
		.INIT('h8)
	) name387 (
		_w533_,
		_w542_,
		_w543_
	);
	LUT2 #(
		.INIT('h1)
	) name388 (
		_w533_,
		_w542_,
		_w544_
	);
	LUT2 #(
		.INIT('h1)
	) name389 (
		_w543_,
		_w544_,
		_w545_
	);
	LUT2 #(
		.INIT('h2)
	) name390 (
		\1971(206)_pad ,
		\1981(208)_pad ,
		_w546_
	);
	LUT2 #(
		.INIT('h4)
	) name391 (
		\1971(206)_pad ,
		\1981(208)_pad ,
		_w547_
	);
	LUT2 #(
		.INIT('h1)
	) name392 (
		_w546_,
		_w547_,
		_w548_
	);
	LUT2 #(
		.INIT('h1)
	) name393 (
		\1976(207)_pad ,
		\2474(231)_pad ,
		_w549_
	);
	LUT2 #(
		.INIT('h8)
	) name394 (
		\1976(207)_pad ,
		\2474(231)_pad ,
		_w550_
	);
	LUT2 #(
		.INIT('h1)
	) name395 (
		_w549_,
		_w550_,
		_w551_
	);
	LUT2 #(
		.INIT('h2)
	) name396 (
		_w548_,
		_w551_,
		_w552_
	);
	LUT2 #(
		.INIT('h4)
	) name397 (
		_w548_,
		_w551_,
		_w553_
	);
	LUT2 #(
		.INIT('h1)
	) name398 (
		_w552_,
		_w553_,
		_w554_
	);
	LUT2 #(
		.INIT('h1)
	) name399 (
		\1961(204)_pad ,
		\1986(209)_pad ,
		_w555_
	);
	LUT2 #(
		.INIT('h8)
	) name400 (
		\1961(204)_pad ,
		\1986(209)_pad ,
		_w556_
	);
	LUT2 #(
		.INIT('h1)
	) name401 (
		_w555_,
		_w556_,
		_w557_
	);
	LUT2 #(
		.INIT('h2)
	) name402 (
		\1966(205)_pad ,
		\1991(210)_pad ,
		_w558_
	);
	LUT2 #(
		.INIT('h4)
	) name403 (
		\1966(205)_pad ,
		\1991(210)_pad ,
		_w559_
	);
	LUT2 #(
		.INIT('h1)
	) name404 (
		_w558_,
		_w559_,
		_w560_
	);
	LUT2 #(
		.INIT('h8)
	) name405 (
		_w557_,
		_w560_,
		_w561_
	);
	LUT2 #(
		.INIT('h1)
	) name406 (
		_w557_,
		_w560_,
		_w562_
	);
	LUT2 #(
		.INIT('h1)
	) name407 (
		_w561_,
		_w562_,
		_w563_
	);
	LUT2 #(
		.INIT('h2)
	) name408 (
		\1956(203)_pad ,
		\1996(211)_pad ,
		_w564_
	);
	LUT2 #(
		.INIT('h4)
	) name409 (
		\1956(203)_pad ,
		\1996(211)_pad ,
		_w565_
	);
	LUT2 #(
		.INIT('h1)
	) name410 (
		_w564_,
		_w565_,
		_w566_
	);
	LUT2 #(
		.INIT('h2)
	) name411 (
		_w563_,
		_w566_,
		_w567_
	);
	LUT2 #(
		.INIT('h4)
	) name412 (
		_w563_,
		_w566_,
		_w568_
	);
	LUT2 #(
		.INIT('h1)
	) name413 (
		_w567_,
		_w568_,
		_w569_
	);
	LUT2 #(
		.INIT('h8)
	) name414 (
		_w554_,
		_w569_,
		_w570_
	);
	LUT2 #(
		.INIT('h1)
	) name415 (
		_w554_,
		_w569_,
		_w571_
	);
	LUT2 #(
		.INIT('h1)
	) name416 (
		_w570_,
		_w571_,
		_w572_
	);
	LUT2 #(
		.INIT('h2)
	) name417 (
		_w432_,
		_w545_,
		_w573_
	);
	LUT2 #(
		.INIT('h4)
	) name418 (
		_w572_,
		_w573_,
		_w574_
	);
	LUT2 #(
		.INIT('h4)
	) name419 (
		_w493_,
		_w574_,
		_w575_
	);
	LUT2 #(
		.INIT('h4)
	) name420 (
		_w525_,
		_w575_,
		_w576_
	);
	LUT2 #(
		.INIT('h4)
	) name421 (
		_w465_,
		_w576_,
		_w577_
	);
	LUT2 #(
		.INIT('h8)
	) name422 (
		\567(194)_pad ,
		_w439_,
		_w578_
	);
	LUT2 #(
		.INIT('h8)
	) name423 (
		\15(10)_pad ,
		\2(1)_pad ,
		_w579_
	);
	LUT2 #(
		.INIT('h8)
	) name424 (
		\661(196)_pad ,
		_w579_,
		_w580_
	);
	LUT2 #(
		.INIT('h8)
	) name425 (
		_w426_,
		_w430_,
		_w581_
	);
	LUT2 #(
		.INIT('h4)
	) name426 (
		\868(198)_pad ,
		_w175_,
		_w582_
	);
	LUT2 #(
		.INIT('h4)
	) name427 (
		\559(193)_pad ,
		\868(198)_pad ,
		_w583_
	);
	LUT2 #(
		.INIT('h8)
	) name428 (
		_w166_,
		_w583_,
		_w584_
	);
	LUT2 #(
		.INIT('h1)
	) name429 (
		_w582_,
		_w584_,
		_w585_
	);
	LUT2 #(
		.INIT('h2)
	) name430 (
		\868(198)_pad ,
		_w373_,
		_w586_
	);
	LUT2 #(
		.INIT('h1)
	) name431 (
		\868(198)_pad ,
		_w166_,
		_w587_
	);
	LUT2 #(
		.INIT('h1)
	) name432 (
		_w586_,
		_w587_,
		_w588_
	);
	LUT2 #(
		.INIT('h8)
	) name433 (
		_w167_,
		_w455_,
		_w589_
	);
	LUT2 #(
		.INIT('h1)
	) name434 (
		_w167_,
		_w455_,
		_w590_
	);
	LUT2 #(
		.INIT('h1)
	) name435 (
		_w589_,
		_w590_,
		_w591_
	);
	LUT2 #(
		.INIT('h2)
	) name436 (
		\868(198)_pad ,
		_w591_,
		_w592_
	);
	LUT2 #(
		.INIT('h1)
	) name437 (
		\868(198)_pad ,
		_w184_,
		_w593_
	);
	LUT2 #(
		.INIT('h1)
	) name438 (
		_w592_,
		_w593_,
		_w594_
	);
	LUT2 #(
		.INIT('h2)
	) name439 (
		\868(198)_pad ,
		_w238_,
		_w595_
	);
	LUT2 #(
		.INIT('h1)
	) name440 (
		\868(198)_pad ,
		_w310_,
		_w596_
	);
	LUT2 #(
		.INIT('h1)
	) name441 (
		_w595_,
		_w596_,
		_w597_
	);
	LUT2 #(
		.INIT('h1)
	) name442 (
		\1384(202)_pad ,
		_w227_,
		_w598_
	);
	LUT2 #(
		.INIT('h8)
	) name443 (
		\40(29)_pad ,
		_w299_,
		_w599_
	);
	LUT2 #(
		.INIT('h8)
	) name444 (
		_w598_,
		_w599_,
		_w600_
	);
	LUT2 #(
		.INIT('h2)
	) name445 (
		\1956(203)_pad ,
		_w600_,
		_w601_
	);
	LUT2 #(
		.INIT('h8)
	) name446 (
		\2072(214)_pad ,
		_w600_,
		_w602_
	);
	LUT2 #(
		.INIT('h1)
	) name447 (
		_w601_,
		_w602_,
		_w603_
	);
	LUT2 #(
		.INIT('h8)
	) name448 (
		_w310_,
		_w603_,
		_w604_
	);
	LUT2 #(
		.INIT('h2)
	) name449 (
		\1348(201)_pad ,
		_w600_,
		_w605_
	);
	LUT2 #(
		.INIT('h8)
	) name450 (
		\2067(213)_pad ,
		_w600_,
		_w606_
	);
	LUT2 #(
		.INIT('h1)
	) name451 (
		_w605_,
		_w606_,
		_w607_
	);
	LUT2 #(
		.INIT('h8)
	) name452 (
		_w166_,
		_w607_,
		_w608_
	);
	LUT2 #(
		.INIT('h8)
	) name453 (
		\1996(211)_pad ,
		_w600_,
		_w609_
	);
	LUT2 #(
		.INIT('h1)
	) name454 (
		_w166_,
		_w607_,
		_w610_
	);
	LUT2 #(
		.INIT('h2)
	) name455 (
		\1341(200)_pad ,
		_w600_,
		_w611_
	);
	LUT2 #(
		.INIT('h2)
	) name456 (
		_w175_,
		_w609_,
		_w612_
	);
	LUT2 #(
		.INIT('h4)
	) name457 (
		_w611_,
		_w612_,
		_w613_
	);
	LUT2 #(
		.INIT('h4)
	) name458 (
		_w610_,
		_w613_,
		_w614_
	);
	LUT2 #(
		.INIT('h1)
	) name459 (
		_w604_,
		_w608_,
		_w615_
	);
	LUT2 #(
		.INIT('h4)
	) name460 (
		_w614_,
		_w615_,
		_w616_
	);
	LUT2 #(
		.INIT('h8)
	) name461 (
		\2084(216)_pad ,
		_w600_,
		_w617_
	);
	LUT2 #(
		.INIT('h2)
	) name462 (
		\1966(205)_pad ,
		_w600_,
		_w618_
	);
	LUT2 #(
		.INIT('h2)
	) name463 (
		\8(7)_pad ,
		_w617_,
		_w619_
	);
	LUT2 #(
		.INIT('h4)
	) name464 (
		_w618_,
		_w619_,
		_w620_
	);
	LUT2 #(
		.INIT('h2)
	) name465 (
		\8(7)_pad ,
		_w238_,
		_w621_
	);
	LUT2 #(
		.INIT('h4)
	) name466 (
		_w620_,
		_w621_,
		_w622_
	);
	LUT2 #(
		.INIT('h1)
	) name467 (
		_w310_,
		_w603_,
		_w623_
	);
	LUT2 #(
		.INIT('h2)
	) name468 (
		\1961(204)_pad ,
		_w600_,
		_w624_
	);
	LUT2 #(
		.INIT('h8)
	) name469 (
		\2078(215)_pad ,
		_w600_,
		_w625_
	);
	LUT2 #(
		.INIT('h1)
	) name470 (
		_w624_,
		_w625_,
		_w626_
	);
	LUT2 #(
		.INIT('h8)
	) name471 (
		_w373_,
		_w626_,
		_w627_
	);
	LUT2 #(
		.INIT('h1)
	) name472 (
		_w373_,
		_w626_,
		_w628_
	);
	LUT2 #(
		.INIT('h8)
	) name473 (
		_w238_,
		_w620_,
		_w629_
	);
	LUT2 #(
		.INIT('h1)
	) name474 (
		_w623_,
		_w627_,
		_w630_
	);
	LUT2 #(
		.INIT('h4)
	) name475 (
		_w628_,
		_w630_,
		_w631_
	);
	LUT2 #(
		.INIT('h1)
	) name476 (
		_w622_,
		_w629_,
		_w632_
	);
	LUT2 #(
		.INIT('h8)
	) name477 (
		_w631_,
		_w632_,
		_w633_
	);
	LUT2 #(
		.INIT('h4)
	) name478 (
		_w616_,
		_w633_,
		_w634_
	);
	LUT2 #(
		.INIT('h4)
	) name479 (
		_w622_,
		_w627_,
		_w635_
	);
	LUT2 #(
		.INIT('h1)
	) name480 (
		_w629_,
		_w635_,
		_w636_
	);
	LUT2 #(
		.INIT('h4)
	) name481 (
		_w634_,
		_w636_,
		_w637_
	);
	LUT2 #(
		.INIT('h2)
	) name482 (
		\8(7)_pad ,
		_w600_,
		_w638_
	);
	LUT2 #(
		.INIT('h4)
	) name483 (
		\1976(207)_pad ,
		_w345_,
		_w639_
	);
	LUT2 #(
		.INIT('h8)
	) name484 (
		_w638_,
		_w639_,
		_w640_
	);
	LUT2 #(
		.INIT('h2)
	) name485 (
		\1981(208)_pad ,
		_w252_,
		_w641_
	);
	LUT2 #(
		.INIT('h8)
	) name486 (
		_w638_,
		_w641_,
		_w642_
	);
	LUT2 #(
		.INIT('h2)
	) name487 (
		\1976(207)_pad ,
		_w345_,
		_w643_
	);
	LUT2 #(
		.INIT('h8)
	) name488 (
		_w638_,
		_w643_,
		_w644_
	);
	LUT2 #(
		.INIT('h4)
	) name489 (
		\1981(208)_pad ,
		_w252_,
		_w645_
	);
	LUT2 #(
		.INIT('h8)
	) name490 (
		_w638_,
		_w645_,
		_w646_
	);
	LUT2 #(
		.INIT('h8)
	) name491 (
		\2090(217)_pad ,
		_w600_,
		_w647_
	);
	LUT2 #(
		.INIT('h2)
	) name492 (
		\1971(206)_pad ,
		_w600_,
		_w648_
	);
	LUT2 #(
		.INIT('h2)
	) name493 (
		\8(7)_pad ,
		_w647_,
		_w649_
	);
	LUT2 #(
		.INIT('h4)
	) name494 (
		_w648_,
		_w649_,
		_w650_
	);
	LUT2 #(
		.INIT('h8)
	) name495 (
		_w357_,
		_w650_,
		_w651_
	);
	LUT2 #(
		.INIT('h2)
	) name496 (
		\8(7)_pad ,
		_w357_,
		_w652_
	);
	LUT2 #(
		.INIT('h4)
	) name497 (
		_w650_,
		_w652_,
		_w653_
	);
	LUT2 #(
		.INIT('h1)
	) name498 (
		_w640_,
		_w642_,
		_w654_
	);
	LUT2 #(
		.INIT('h1)
	) name499 (
		_w644_,
		_w646_,
		_w655_
	);
	LUT2 #(
		.INIT('h8)
	) name500 (
		_w654_,
		_w655_,
		_w656_
	);
	LUT2 #(
		.INIT('h4)
	) name501 (
		_w651_,
		_w656_,
		_w657_
	);
	LUT2 #(
		.INIT('h4)
	) name502 (
		_w653_,
		_w657_,
		_w658_
	);
	LUT2 #(
		.INIT('h4)
	) name503 (
		_w637_,
		_w658_,
		_w659_
	);
	LUT2 #(
		.INIT('h4)
	) name504 (
		_w644_,
		_w651_,
		_w660_
	);
	LUT2 #(
		.INIT('h1)
	) name505 (
		_w640_,
		_w660_,
		_w661_
	);
	LUT2 #(
		.INIT('h1)
	) name506 (
		_w642_,
		_w661_,
		_w662_
	);
	LUT2 #(
		.INIT('h1)
	) name507 (
		_w646_,
		_w662_,
		_w663_
	);
	LUT2 #(
		.INIT('h4)
	) name508 (
		_w659_,
		_w663_,
		_w664_
	);
	LUT2 #(
		.INIT('h4)
	) name509 (
		_w598_,
		_w599_,
		_w665_
	);
	LUT2 #(
		.INIT('h4)
	) name510 (
		\2067(213)_pad ,
		_w323_,
		_w666_
	);
	LUT2 #(
		.INIT('h2)
	) name511 (
		\1986(209)_pad ,
		_w274_,
		_w667_
	);
	LUT2 #(
		.INIT('h2)
	) name512 (
		\1991(210)_pad ,
		_w288_,
		_w668_
	);
	LUT2 #(
		.INIT('h4)
	) name513 (
		\1986(209)_pad ,
		_w274_,
		_w669_
	);
	LUT2 #(
		.INIT('h2)
	) name514 (
		\2067(213)_pad ,
		_w323_,
		_w670_
	);
	LUT2 #(
		.INIT('h2)
	) name515 (
		\1996(211)_pad ,
		_w335_,
		_w671_
	);
	LUT2 #(
		.INIT('h1)
	) name516 (
		_w670_,
		_w671_,
		_w672_
	);
	LUT2 #(
		.INIT('h4)
	) name517 (
		\1991(210)_pad ,
		_w288_,
		_w673_
	);
	LUT2 #(
		.INIT('h4)
	) name518 (
		\1996(211)_pad ,
		_w335_,
		_w674_
	);
	LUT2 #(
		.INIT('h1)
	) name519 (
		_w673_,
		_w674_,
		_w675_
	);
	LUT2 #(
		.INIT('h1)
	) name520 (
		_w666_,
		_w667_,
		_w676_
	);
	LUT2 #(
		.INIT('h1)
	) name521 (
		_w668_,
		_w669_,
		_w677_
	);
	LUT2 #(
		.INIT('h8)
	) name522 (
		_w676_,
		_w677_,
		_w678_
	);
	LUT2 #(
		.INIT('h8)
	) name523 (
		_w672_,
		_w675_,
		_w679_
	);
	LUT2 #(
		.INIT('h8)
	) name524 (
		_w678_,
		_w679_,
		_w680_
	);
	LUT2 #(
		.INIT('h2)
	) name525 (
		_w665_,
		_w680_,
		_w681_
	);
	LUT2 #(
		.INIT('h1)
	) name526 (
		_w664_,
		_w681_,
		_w682_
	);
	LUT2 #(
		.INIT('h4)
	) name527 (
		_w668_,
		_w669_,
		_w683_
	);
	LUT2 #(
		.INIT('h2)
	) name528 (
		_w675_,
		_w683_,
		_w684_
	);
	LUT2 #(
		.INIT('h2)
	) name529 (
		_w672_,
		_w684_,
		_w685_
	);
	LUT2 #(
		.INIT('h1)
	) name530 (
		_w666_,
		_w685_,
		_w686_
	);
	LUT2 #(
		.INIT('h2)
	) name531 (
		_w665_,
		_w686_,
		_w687_
	);
	LUT2 #(
		.INIT('h1)
	) name532 (
		_w682_,
		_w687_,
		_w688_
	);
	assign \145(1358)_pad  = _w190_ ;
	assign \148(851)_pad  = _w191_ ;
	assign \150(1277)_pad  = _w415_ ;
	assign \153(671)_pad  = _w176_ ;
	assign \156(1046)_pad  = _w419_ ;
	assign \158(349)_pad  = _w422_ ;
	assign \160(609)_pad  = _w299_ ;
	assign \162(612)_pad  = _w202_ ;
	assign \164(607)_pad  = _w227_ ;
	assign \166(625)_pad  = _w357_ ;
	assign \168(623)_pad  = _w238_ ;
	assign \171(621)_pad  = _w373_ ;
	assign \173(389)_pad  = _w423_ ;
	assign \176(803)_pad  = _w435_ ;
	assign \188(761)_pad  = _w438_ ;
	assign \217(423)_pad  = _w440_ ;
	assign \218(311)_pad  = \44(31)_pad ;
	assign \219(302)_pad  = \132(105)_pad ;
	assign \220(306)_pad  = \82(63)_pad ;
	assign \221(305)_pad  = \96(75)_pad ;
	assign \223(413)_pad  = _w439_ ;
	assign \225(1424)_pad  = _w577_ ;
	assign \227(1179)_pad  = _w545_ ;
	assign \229(1180)_pad  = _w572_ ;
	assign \234(376)_pad  = _w578_ ;
	assign \235(307)_pad  = \69(52)_pad ;
	assign \236(303)_pad  = \120(95)_pad ;
	assign \237(309)_pad  = \57(42)_pad ;
	assign \238(304)_pad  = \108(85)_pad ;
	assign \259(414)_pad  = _w580_ ;
	assign \261(506)_pad  = _w581_ ;
	assign \282(922)_pad  = _w585_ ;
	assign \284(847)_pad  = _w588_ ;
	assign \286(696)_pad  = _w238_ ;
	assign \288(700)_pad  = _w345_ ;
	assign \290(704)_pad  = _w274_ ;
	assign \295(1400)_pad  = _w594_ ;
	assign \297(849)_pad  = _w597_ ;
	assign \299(692)_pad  = _w310_ ;
	assign \301(694)_pad  = _w373_ ;
	assign \303(698)_pad  = _w357_ ;
	assign \305(702)_pad  = _w252_ ;
	assign \325(507)_pad  = _w581_ ;
	assign \329(1414)_pad  = _w688_ ;
	assign \_al_n0  = 1'b0;
	assign \u1082_syn_3  = _w432_ ;
	assign \u1396_syn_3  = _w577_ ;
	assign \u1414_syn_3  = _w465_ ;
	assign \u1447_syn_3  = _w525_ ;
	assign \u538_syn_3  = _w415_ ;
	assign \u539_syn_3  = _w493_ ;
endmodule;