module top (a_pad, b_pad, c_pad, e_pad, f_pad, g_pad, h_pad, i_pad, j_pad, k_pad, l_pad, m_pad, n_pad, o_pad, p_pad, q_pad, r_pad, s_pad, t_pad, u_pad, v_pad, w_pad, x_pad, y_pad, \a0_pad , \b0_pad , \c0_pad , \d0_pad , \e0_pad , \f0_pad , \g0_pad , \h0_pad , \i0_pad , \j0_pad , \k0_pad , \l0_pad , \m0_pad , \n0_pad , \o0_pad , \p0_pad , \q0_pad , \r0_pad , \s0_pad , \t0_pad , z_pad);
	input a_pad ;
	input b_pad ;
	input c_pad ;
	input e_pad ;
	input f_pad ;
	input g_pad ;
	input h_pad ;
	input i_pad ;
	input j_pad ;
	input k_pad ;
	input l_pad ;
	input m_pad ;
	input n_pad ;
	input o_pad ;
	input p_pad ;
	input q_pad ;
	input r_pad ;
	input s_pad ;
	input t_pad ;
	input u_pad ;
	input v_pad ;
	input w_pad ;
	input x_pad ;
	input y_pad ;
	output \a0_pad  ;
	output \b0_pad  ;
	output \c0_pad  ;
	output \d0_pad  ;
	output \e0_pad  ;
	output \f0_pad  ;
	output \g0_pad  ;
	output \h0_pad  ;
	output \i0_pad  ;
	output \j0_pad  ;
	output \k0_pad  ;
	output \l0_pad  ;
	output \m0_pad  ;
	output \n0_pad  ;
	output \o0_pad  ;
	output \p0_pad  ;
	output \q0_pad  ;
	output \r0_pad  ;
	output \s0_pad  ;
	output \t0_pad  ;
	output z_pad ;
	wire _w160_ ;
	wire _w159_ ;
	wire _w158_ ;
	wire _w157_ ;
	wire _w156_ ;
	wire _w155_ ;
	wire _w154_ ;
	wire _w153_ ;
	wire _w152_ ;
	wire _w83_ ;
	wire _w82_ ;
	wire _w81_ ;
	wire _w80_ ;
	wire _w79_ ;
	wire _w78_ ;
	wire _w77_ ;
	wire _w76_ ;
	wire _w75_ ;
	wire _w74_ ;
	wire _w73_ ;
	wire _w72_ ;
	wire _w71_ ;
	wire _w70_ ;
	wire _w69_ ;
	wire _w68_ ;
	wire _w67_ ;
	wire _w66_ ;
	wire _w65_ ;
	wire _w64_ ;
	wire _w63_ ;
	wire _w62_ ;
	wire _w61_ ;
	wire _w60_ ;
	wire _w59_ ;
	wire _w58_ ;
	wire _w57_ ;
	wire _w56_ ;
	wire _w55_ ;
	wire _w54_ ;
	wire _w37_ ;
	wire _w36_ ;
	wire _w35_ ;
	wire _w34_ ;
	wire _w33_ ;
	wire _w32_ ;
	wire _w31_ ;
	wire _w30_ ;
	wire _w29_ ;
	wire _w28_ ;
	wire _w27_ ;
	wire _w26_ ;
	wire _w25_ ;
	wire _w38_ ;
	wire _w39_ ;
	wire _w40_ ;
	wire _w41_ ;
	wire _w42_ ;
	wire _w43_ ;
	wire _w44_ ;
	wire _w45_ ;
	wire _w46_ ;
	wire _w47_ ;
	wire _w48_ ;
	wire _w49_ ;
	wire _w50_ ;
	wire _w51_ ;
	wire _w52_ ;
	wire _w53_ ;
	wire _w84_ ;
	wire _w85_ ;
	wire _w86_ ;
	wire _w87_ ;
	wire _w88_ ;
	wire _w89_ ;
	wire _w90_ ;
	wire _w91_ ;
	wire _w92_ ;
	wire _w93_ ;
	wire _w94_ ;
	wire _w95_ ;
	wire _w96_ ;
	wire _w97_ ;
	wire _w98_ ;
	wire _w99_ ;
	wire _w100_ ;
	wire _w101_ ;
	wire _w102_ ;
	wire _w103_ ;
	wire _w104_ ;
	wire _w105_ ;
	wire _w106_ ;
	wire _w107_ ;
	wire _w108_ ;
	wire _w109_ ;
	wire _w110_ ;
	wire _w111_ ;
	wire _w112_ ;
	wire _w113_ ;
	wire _w114_ ;
	wire _w115_ ;
	wire _w116_ ;
	wire _w117_ ;
	wire _w118_ ;
	wire _w119_ ;
	wire _w120_ ;
	wire _w121_ ;
	wire _w122_ ;
	wire _w123_ ;
	wire _w124_ ;
	wire _w125_ ;
	wire _w126_ ;
	wire _w127_ ;
	wire _w128_ ;
	wire _w129_ ;
	wire _w130_ ;
	wire _w131_ ;
	wire _w132_ ;
	wire _w133_ ;
	wire _w134_ ;
	wire _w135_ ;
	wire _w136_ ;
	wire _w137_ ;
	wire _w138_ ;
	wire _w139_ ;
	wire _w140_ ;
	wire _w141_ ;
	wire _w142_ ;
	wire _w143_ ;
	wire _w144_ ;
	wire _w145_ ;
	wire _w146_ ;
	wire _w147_ ;
	wire _w148_ ;
	wire _w149_ ;
	wire _w150_ ;
	wire _w151_ ;
	LUT2 #(
		.INIT('h2)
	) name0 (
		v_pad,
		w_pad,
		_w25_
	);
	LUT2 #(
		.INIT('h2)
	) name1 (
		q_pad,
		_w25_,
		_w26_
	);
	LUT2 #(
		.INIT('h1)
	) name2 (
		v_pad,
		y_pad,
		_w27_
	);
	LUT2 #(
		.INIT('h2)
	) name3 (
		s_pad,
		t_pad,
		_w28_
	);
	LUT2 #(
		.INIT('h8)
	) name4 (
		_w27_,
		_w28_,
		_w29_
	);
	LUT2 #(
		.INIT('h8)
	) name5 (
		u_pad,
		_w29_,
		_w30_
	);
	LUT2 #(
		.INIT('h1)
	) name6 (
		s_pad,
		t_pad,
		_w31_
	);
	LUT2 #(
		.INIT('h4)
	) name7 (
		_w27_,
		_w31_,
		_w32_
	);
	LUT2 #(
		.INIT('h2)
	) name8 (
		u_pad,
		v_pad,
		_w33_
	);
	LUT2 #(
		.INIT('h4)
	) name9 (
		u_pad,
		v_pad,
		_w34_
	);
	LUT2 #(
		.INIT('h1)
	) name10 (
		_w33_,
		_w34_,
		_w35_
	);
	LUT2 #(
		.INIT('h2)
	) name11 (
		_w32_,
		_w35_,
		_w36_
	);
	LUT2 #(
		.INIT('h1)
	) name12 (
		t_pad,
		u_pad,
		_w37_
	);
	LUT2 #(
		.INIT('h2)
	) name13 (
		v_pad,
		_w37_,
		_w38_
	);
	LUT2 #(
		.INIT('h8)
	) name14 (
		f_pad,
		_w38_,
		_w39_
	);
	LUT2 #(
		.INIT('h1)
	) name15 (
		w_pad,
		_w36_,
		_w40_
	);
	LUT2 #(
		.INIT('h4)
	) name16 (
		_w39_,
		_w40_,
		_w41_
	);
	LUT2 #(
		.INIT('h1)
	) name17 (
		_w26_,
		_w30_,
		_w42_
	);
	LUT2 #(
		.INIT('h4)
	) name18 (
		_w41_,
		_w42_,
		_w43_
	);
	LUT2 #(
		.INIT('h2)
	) name19 (
		g_pad,
		_w37_,
		_w44_
	);
	LUT2 #(
		.INIT('h2)
	) name20 (
		v_pad,
		_w44_,
		_w45_
	);
	LUT2 #(
		.INIT('h8)
	) name21 (
		y_pad,
		_w31_,
		_w46_
	);
	LUT2 #(
		.INIT('h2)
	) name22 (
		u_pad,
		_w46_,
		_w47_
	);
	LUT2 #(
		.INIT('h1)
	) name23 (
		v_pad,
		_w47_,
		_w48_
	);
	LUT2 #(
		.INIT('h2)
	) name24 (
		w_pad,
		_w29_,
		_w49_
	);
	LUT2 #(
		.INIT('h1)
	) name25 (
		_w45_,
		_w49_,
		_w50_
	);
	LUT2 #(
		.INIT('h4)
	) name26 (
		_w48_,
		_w50_,
		_w51_
	);
	LUT2 #(
		.INIT('h8)
	) name27 (
		q_pad,
		_w32_,
		_w52_
	);
	LUT2 #(
		.INIT('h1)
	) name28 (
		u_pad,
		w_pad,
		_w53_
	);
	LUT2 #(
		.INIT('h1)
	) name29 (
		_w52_,
		_w53_,
		_w54_
	);
	LUT2 #(
		.INIT('h1)
	) name30 (
		v_pad,
		_w54_,
		_w55_
	);
	LUT2 #(
		.INIT('h1)
	) name31 (
		h_pad,
		_w33_,
		_w56_
	);
	LUT2 #(
		.INIT('h8)
	) name32 (
		_w30_,
		_w56_,
		_w57_
	);
	LUT2 #(
		.INIT('h2)
	) name33 (
		q_pad,
		_w57_,
		_w58_
	);
	LUT2 #(
		.INIT('h2)
	) name34 (
		w_pad,
		_w58_,
		_w59_
	);
	LUT2 #(
		.INIT('h4)
	) name35 (
		_w37_,
		_w56_,
		_w60_
	);
	LUT2 #(
		.INIT('h8)
	) name36 (
		s_pad,
		_w37_,
		_w61_
	);
	LUT2 #(
		.INIT('h1)
	) name37 (
		_w49_,
		_w61_,
		_w62_
	);
	LUT2 #(
		.INIT('h4)
	) name38 (
		_w60_,
		_w62_,
		_w63_
	);
	LUT2 #(
		.INIT('h1)
	) name39 (
		_w59_,
		_w63_,
		_w64_
	);
	LUT2 #(
		.INIT('h1)
	) name40 (
		_w55_,
		_w64_,
		_w65_
	);
	LUT2 #(
		.INIT('h2)
	) name41 (
		i_pad,
		_w37_,
		_w66_
	);
	LUT2 #(
		.INIT('h2)
	) name42 (
		v_pad,
		_w66_,
		_w67_
	);
	LUT2 #(
		.INIT('h2)
	) name43 (
		t_pad,
		u_pad,
		_w68_
	);
	LUT2 #(
		.INIT('h8)
	) name44 (
		s_pad,
		_w68_,
		_w69_
	);
	LUT2 #(
		.INIT('h1)
	) name45 (
		v_pad,
		_w69_,
		_w70_
	);
	LUT2 #(
		.INIT('h1)
	) name46 (
		w_pad,
		_w67_,
		_w71_
	);
	LUT2 #(
		.INIT('h4)
	) name47 (
		_w70_,
		_w71_,
		_w72_
	);
	LUT2 #(
		.INIT('h1)
	) name48 (
		s_pad,
		v_pad,
		_w73_
	);
	LUT2 #(
		.INIT('h1)
	) name49 (
		_w28_,
		_w73_,
		_w74_
	);
	LUT2 #(
		.INIT('h1)
	) name50 (
		u_pad,
		_w74_,
		_w75_
	);
	LUT2 #(
		.INIT('h8)
	) name51 (
		j_pad,
		_w38_,
		_w76_
	);
	LUT2 #(
		.INIT('h1)
	) name52 (
		_w75_,
		_w76_,
		_w77_
	);
	LUT2 #(
		.INIT('h1)
	) name53 (
		w_pad,
		_w77_,
		_w78_
	);
	LUT2 #(
		.INIT('h1)
	) name54 (
		a_pad,
		k_pad,
		_w79_
	);
	LUT2 #(
		.INIT('h8)
	) name55 (
		l_pad,
		_w79_,
		_w80_
	);
	LUT2 #(
		.INIT('h2)
	) name56 (
		k_pad,
		l_pad,
		_w81_
	);
	LUT2 #(
		.INIT('h4)
	) name57 (
		m_pad,
		n_pad,
		_w82_
	);
	LUT2 #(
		.INIT('h4)
	) name58 (
		a_pad,
		_w81_,
		_w83_
	);
	LUT2 #(
		.INIT('h4)
	) name59 (
		_w82_,
		_w83_,
		_w84_
	);
	LUT2 #(
		.INIT('h1)
	) name60 (
		_w80_,
		_w84_,
		_w85_
	);
	LUT2 #(
		.INIT('h8)
	) name61 (
		k_pad,
		l_pad,
		_w86_
	);
	LUT2 #(
		.INIT('h8)
	) name62 (
		m_pad,
		_w86_,
		_w87_
	);
	LUT2 #(
		.INIT('h1)
	) name63 (
		m_pad,
		_w86_,
		_w88_
	);
	LUT2 #(
		.INIT('h1)
	) name64 (
		a_pad,
		_w87_,
		_w89_
	);
	LUT2 #(
		.INIT('h4)
	) name65 (
		_w88_,
		_w89_,
		_w90_
	);
	LUT2 #(
		.INIT('h4)
	) name66 (
		m_pad,
		_w81_,
		_w91_
	);
	LUT2 #(
		.INIT('h8)
	) name67 (
		n_pad,
		_w87_,
		_w92_
	);
	LUT2 #(
		.INIT('h1)
	) name68 (
		n_pad,
		_w87_,
		_w93_
	);
	LUT2 #(
		.INIT('h1)
	) name69 (
		a_pad,
		_w91_,
		_w94_
	);
	LUT2 #(
		.INIT('h4)
	) name70 (
		_w92_,
		_w94_,
		_w95_
	);
	LUT2 #(
		.INIT('h4)
	) name71 (
		_w93_,
		_w95_,
		_w96_
	);
	LUT2 #(
		.INIT('h8)
	) name72 (
		_w81_,
		_w82_,
		_w97_
	);
	LUT2 #(
		.INIT('h1)
	) name73 (
		x_pad,
		_w97_,
		_w98_
	);
	LUT2 #(
		.INIT('h2)
	) name74 (
		o_pad,
		_w98_,
		_w99_
	);
	LUT2 #(
		.INIT('h4)
	) name75 (
		o_pad,
		_w98_,
		_w100_
	);
	LUT2 #(
		.INIT('h1)
	) name76 (
		a_pad,
		_w99_,
		_w101_
	);
	LUT2 #(
		.INIT('h4)
	) name77 (
		_w100_,
		_w101_,
		_w102_
	);
	LUT2 #(
		.INIT('h8)
	) name78 (
		p_pad,
		_w99_,
		_w103_
	);
	LUT2 #(
		.INIT('h4)
	) name79 (
		q_pad,
		r_pad,
		_w104_
	);
	LUT2 #(
		.INIT('h2)
	) name80 (
		_w99_,
		_w104_,
		_w105_
	);
	LUT2 #(
		.INIT('h1)
	) name81 (
		p_pad,
		_w105_,
		_w106_
	);
	LUT2 #(
		.INIT('h1)
	) name82 (
		a_pad,
		_w103_,
		_w107_
	);
	LUT2 #(
		.INIT('h4)
	) name83 (
		_w106_,
		_w107_,
		_w108_
	);
	LUT2 #(
		.INIT('h1)
	) name84 (
		q_pad,
		_w103_,
		_w109_
	);
	LUT2 #(
		.INIT('h8)
	) name85 (
		q_pad,
		_w103_,
		_w110_
	);
	LUT2 #(
		.INIT('h1)
	) name86 (
		a_pad,
		_w109_,
		_w111_
	);
	LUT2 #(
		.INIT('h4)
	) name87 (
		_w110_,
		_w111_,
		_w112_
	);
	LUT2 #(
		.INIT('h1)
	) name88 (
		p_pad,
		q_pad,
		_w113_
	);
	LUT2 #(
		.INIT('h8)
	) name89 (
		p_pad,
		q_pad,
		_w114_
	);
	LUT2 #(
		.INIT('h8)
	) name90 (
		r_pad,
		_w114_,
		_w115_
	);
	LUT2 #(
		.INIT('h1)
	) name91 (
		_w113_,
		_w115_,
		_w116_
	);
	LUT2 #(
		.INIT('h2)
	) name92 (
		_w99_,
		_w116_,
		_w117_
	);
	LUT2 #(
		.INIT('h1)
	) name93 (
		r_pad,
		_w110_,
		_w118_
	);
	LUT2 #(
		.INIT('h1)
	) name94 (
		a_pad,
		_w117_,
		_w119_
	);
	LUT2 #(
		.INIT('h4)
	) name95 (
		_w118_,
		_w119_,
		_w120_
	);
	LUT2 #(
		.INIT('h4)
	) name96 (
		p_pad,
		_w104_,
		_w121_
	);
	LUT2 #(
		.INIT('h8)
	) name97 (
		_w99_,
		_w121_,
		_w122_
	);
	LUT2 #(
		.INIT('h1)
	) name98 (
		s_pad,
		_w122_,
		_w123_
	);
	LUT2 #(
		.INIT('h8)
	) name99 (
		s_pad,
		_w122_,
		_w124_
	);
	LUT2 #(
		.INIT('h1)
	) name100 (
		a_pad,
		_w123_,
		_w125_
	);
	LUT2 #(
		.INIT('h4)
	) name101 (
		_w124_,
		_w125_,
		_w126_
	);
	LUT2 #(
		.INIT('h8)
	) name102 (
		t_pad,
		_w124_,
		_w127_
	);
	LUT2 #(
		.INIT('h4)
	) name103 (
		_w34_,
		_w124_,
		_w128_
	);
	LUT2 #(
		.INIT('h1)
	) name104 (
		t_pad,
		_w128_,
		_w129_
	);
	LUT2 #(
		.INIT('h1)
	) name105 (
		a_pad,
		_w127_,
		_w130_
	);
	LUT2 #(
		.INIT('h4)
	) name106 (
		_w129_,
		_w130_,
		_w131_
	);
	LUT2 #(
		.INIT('h2)
	) name107 (
		u_pad,
		_w127_,
		_w132_
	);
	LUT2 #(
		.INIT('h8)
	) name108 (
		_w69_,
		_w122_,
		_w133_
	);
	LUT2 #(
		.INIT('h1)
	) name109 (
		_w132_,
		_w133_,
		_w134_
	);
	LUT2 #(
		.INIT('h1)
	) name110 (
		a_pad,
		_w134_,
		_w135_
	);
	LUT2 #(
		.INIT('h4)
	) name111 (
		t_pad,
		u_pad,
		_w136_
	);
	LUT2 #(
		.INIT('h1)
	) name112 (
		_w68_,
		_w136_,
		_w137_
	);
	LUT2 #(
		.INIT('h8)
	) name113 (
		_w124_,
		_w137_,
		_w138_
	);
	LUT2 #(
		.INIT('h2)
	) name114 (
		v_pad,
		_w138_,
		_w139_
	);
	LUT2 #(
		.INIT('h8)
	) name115 (
		_w33_,
		_w127_,
		_w140_
	);
	LUT2 #(
		.INIT('h1)
	) name116 (
		_w139_,
		_w140_,
		_w141_
	);
	LUT2 #(
		.INIT('h1)
	) name117 (
		a_pad,
		_w141_,
		_w142_
	);
	LUT2 #(
		.INIT('h8)
	) name118 (
		y_pad,
		_w73_,
		_w143_
	);
	LUT2 #(
		.INIT('h8)
	) name119 (
		_w136_,
		_w143_,
		_w144_
	);
	LUT2 #(
		.INIT('h1)
	) name120 (
		w_pad,
		_w144_,
		_w145_
	);
	LUT2 #(
		.INIT('h1)
	) name121 (
		a_pad,
		_w30_,
		_w146_
	);
	LUT2 #(
		.INIT('h4)
	) name122 (
		_w145_,
		_w146_,
		_w147_
	);
	LUT2 #(
		.INIT('h2)
	) name123 (
		b_pad,
		x_pad,
		_w148_
	);
	LUT2 #(
		.INIT('h4)
	) name124 (
		b_pad,
		x_pad,
		_w149_
	);
	LUT2 #(
		.INIT('h1)
	) name125 (
		_w148_,
		_w149_,
		_w150_
	);
	LUT2 #(
		.INIT('h1)
	) name126 (
		a_pad,
		_w150_,
		_w151_
	);
	LUT2 #(
		.INIT('h2)
	) name127 (
		c_pad,
		y_pad,
		_w152_
	);
	LUT2 #(
		.INIT('h4)
	) name128 (
		c_pad,
		y_pad,
		_w153_
	);
	LUT2 #(
		.INIT('h1)
	) name129 (
		_w152_,
		_w153_,
		_w154_
	);
	LUT2 #(
		.INIT('h1)
	) name130 (
		a_pad,
		_w154_,
		_w155_
	);
	LUT2 #(
		.INIT('h2)
	) name131 (
		e_pad,
		_w37_,
		_w156_
	);
	LUT2 #(
		.INIT('h2)
	) name132 (
		v_pad,
		_w61_,
		_w157_
	);
	LUT2 #(
		.INIT('h4)
	) name133 (
		_w156_,
		_w157_,
		_w158_
	);
	LUT2 #(
		.INIT('h1)
	) name134 (
		w_pad,
		_w33_,
		_w159_
	);
	LUT2 #(
		.INIT('h4)
	) name135 (
		_w158_,
		_w159_,
		_w160_
	);
	assign \a0_pad  = _w43_ ;
	assign \b0_pad  = _w51_ ;
	assign \c0_pad  = _w65_ ;
	assign \d0_pad  = _w72_ ;
	assign \e0_pad  = _w78_ ;
	assign \f0_pad  = _w79_ ;
	assign \g0_pad  = _w85_ ;
	assign \h0_pad  = _w90_ ;
	assign \i0_pad  = _w96_ ;
	assign \j0_pad  = _w102_ ;
	assign \k0_pad  = _w108_ ;
	assign \l0_pad  = _w112_ ;
	assign \m0_pad  = _w120_ ;
	assign \n0_pad  = _w126_ ;
	assign \o0_pad  = _w131_ ;
	assign \p0_pad  = _w135_ ;
	assign \q0_pad  = _w142_ ;
	assign \r0_pad  = _w147_ ;
	assign \s0_pad  = _w151_ ;
	assign \t0_pad  = _w155_ ;
	assign z_pad = _w160_ ;
endmodule;