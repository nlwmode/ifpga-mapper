module top (\dest_x[0] , \dest_x[1] , \dest_x[2] , \dest_x[3] , \dest_x[4] , \dest_x[5] , \dest_x[6] , \dest_x[7] , \dest_x[8] , \dest_x[9] , \dest_x[10] , \dest_x[11] , \dest_x[12] , \dest_x[13] , \dest_x[14] , \dest_x[15] , \dest_x[16] , \dest_x[17] , \dest_x[18] , \dest_x[19] , \dest_x[20] , \dest_x[21] , \dest_x[22] , \dest_x[23] , \dest_x[24] , \dest_x[25] , \dest_x[26] , \dest_x[27] , \dest_x[28] , \dest_x[29] , \dest_y[0] , \dest_y[1] , \dest_y[2] , \dest_y[3] , \dest_y[4] , \dest_y[5] , \dest_y[6] , \dest_y[7] , \dest_y[8] , \dest_y[9] , \dest_y[10] , \dest_y[11] , \dest_y[12] , \dest_y[13] , \dest_y[14] , \dest_y[15] , \dest_y[16] , \dest_y[17] , \dest_y[18] , \dest_y[19] , \dest_y[20] , \dest_y[21] , \dest_y[22] , \dest_y[23] , \dest_y[24] , \dest_y[25] , \dest_y[26] , \dest_y[27] , \dest_y[28] , \dest_y[29] , \outport[0] , \outport[1] , \outport[2] , \outport[3] , \outport[4] , \outport[5] , \outport[6] , \outport[7] , \outport[8] , \outport[9] , \outport[10] , \outport[11] , \outport[12] , \outport[13] , \outport[14] , \outport[15] , \outport[16] , \outport[17] , \outport[18] , \outport[19] , \outport[20] , \outport[21] , \outport[22] , \outport[23] , \outport[24] , \outport[25] , \outport[26] , \outport[27] , \outport[28] , \outport[29] );
	input \dest_x[0]  ;
	input \dest_x[1]  ;
	input \dest_x[2]  ;
	input \dest_x[3]  ;
	input \dest_x[4]  ;
	input \dest_x[5]  ;
	input \dest_x[6]  ;
	input \dest_x[7]  ;
	input \dest_x[8]  ;
	input \dest_x[9]  ;
	input \dest_x[10]  ;
	input \dest_x[11]  ;
	input \dest_x[12]  ;
	input \dest_x[13]  ;
	input \dest_x[14]  ;
	input \dest_x[15]  ;
	input \dest_x[16]  ;
	input \dest_x[17]  ;
	input \dest_x[18]  ;
	input \dest_x[19]  ;
	input \dest_x[20]  ;
	input \dest_x[21]  ;
	input \dest_x[22]  ;
	input \dest_x[23]  ;
	input \dest_x[24]  ;
	input \dest_x[25]  ;
	input \dest_x[26]  ;
	input \dest_x[27]  ;
	input \dest_x[28]  ;
	input \dest_x[29]  ;
	input \dest_y[0]  ;
	input \dest_y[1]  ;
	input \dest_y[2]  ;
	input \dest_y[3]  ;
	input \dest_y[4]  ;
	input \dest_y[5]  ;
	input \dest_y[6]  ;
	input \dest_y[7]  ;
	input \dest_y[8]  ;
	input \dest_y[9]  ;
	input \dest_y[10]  ;
	input \dest_y[11]  ;
	input \dest_y[12]  ;
	input \dest_y[13]  ;
	input \dest_y[14]  ;
	input \dest_y[15]  ;
	input \dest_y[16]  ;
	input \dest_y[17]  ;
	input \dest_y[18]  ;
	input \dest_y[19]  ;
	input \dest_y[20]  ;
	input \dest_y[21]  ;
	input \dest_y[22]  ;
	input \dest_y[23]  ;
	input \dest_y[24]  ;
	input \dest_y[25]  ;
	input \dest_y[26]  ;
	input \dest_y[27]  ;
	input \dest_y[28]  ;
	input \dest_y[29]  ;
	output \outport[0]  ;
	output \outport[1]  ;
	output \outport[2]  ;
	output \outport[3]  ;
	output \outport[4]  ;
	output \outport[5]  ;
	output \outport[6]  ;
	output \outport[7]  ;
	output \outport[8]  ;
	output \outport[9]  ;
	output \outport[10]  ;
	output \outport[11]  ;
	output \outport[12]  ;
	output \outport[13]  ;
	output \outport[14]  ;
	output \outport[15]  ;
	output \outport[16]  ;
	output \outport[17]  ;
	output \outport[18]  ;
	output \outport[19]  ;
	output \outport[20]  ;
	output \outport[21]  ;
	output \outport[22]  ;
	output \outport[23]  ;
	output \outport[24]  ;
	output \outport[25]  ;
	output \outport[26]  ;
	output \outport[27]  ;
	output \outport[28]  ;
	output \outport[29]  ;
	wire _w183_ ;
	wire _w182_ ;
	wire _w181_ ;
	wire _w180_ ;
	wire _w179_ ;
	wire _w178_ ;
	wire _w177_ ;
	wire _w176_ ;
	wire _w175_ ;
	wire _w174_ ;
	wire _w173_ ;
	wire _w172_ ;
	wire _w171_ ;
	wire _w170_ ;
	wire _w169_ ;
	wire _w168_ ;
	wire _w167_ ;
	wire _w166_ ;
	wire _w165_ ;
	wire _w164_ ;
	wire _w163_ ;
	wire _w162_ ;
	wire _w161_ ;
	wire _w160_ ;
	wire _w159_ ;
	wire _w158_ ;
	wire _w157_ ;
	wire _w156_ ;
	wire _w155_ ;
	wire _w154_ ;
	wire _w153_ ;
	wire _w152_ ;
	wire _w151_ ;
	wire _w150_ ;
	wire _w149_ ;
	wire _w148_ ;
	wire _w147_ ;
	wire _w146_ ;
	wire _w145_ ;
	wire _w144_ ;
	wire _w143_ ;
	wire _w142_ ;
	wire _w141_ ;
	wire _w140_ ;
	wire _w139_ ;
	wire _w138_ ;
	wire _w137_ ;
	wire _w136_ ;
	wire _w135_ ;
	wire _w134_ ;
	wire _w133_ ;
	wire _w132_ ;
	wire _w131_ ;
	wire _w130_ ;
	wire _w129_ ;
	wire _w128_ ;
	wire _w127_ ;
	wire _w126_ ;
	wire _w125_ ;
	wire _w124_ ;
	wire _w123_ ;
	wire _w122_ ;
	wire _w121_ ;
	wire _w90_ ;
	wire _w89_ ;
	wire _w88_ ;
	wire _w87_ ;
	wire _w86_ ;
	wire _w85_ ;
	wire _w84_ ;
	wire _w83_ ;
	wire _w82_ ;
	wire _w81_ ;
	wire _w80_ ;
	wire _w79_ ;
	wire _w78_ ;
	wire _w77_ ;
	wire _w76_ ;
	wire _w75_ ;
	wire _w62_ ;
	wire _w63_ ;
	wire _w64_ ;
	wire _w65_ ;
	wire _w66_ ;
	wire _w67_ ;
	wire _w68_ ;
	wire _w69_ ;
	wire _w70_ ;
	wire _w71_ ;
	wire _w72_ ;
	wire _w73_ ;
	wire _w74_ ;
	wire _w91_ ;
	wire _w92_ ;
	wire _w93_ ;
	wire _w94_ ;
	wire _w95_ ;
	wire _w96_ ;
	wire _w97_ ;
	wire _w98_ ;
	wire _w99_ ;
	wire _w100_ ;
	wire _w101_ ;
	wire _w102_ ;
	wire _w103_ ;
	wire _w104_ ;
	wire _w105_ ;
	wire _w106_ ;
	wire _w107_ ;
	wire _w108_ ;
	wire _w109_ ;
	wire _w110_ ;
	wire _w111_ ;
	wire _w112_ ;
	wire _w113_ ;
	wire _w114_ ;
	wire _w115_ ;
	wire _w116_ ;
	wire _w117_ ;
	wire _w118_ ;
	wire _w119_ ;
	wire _w120_ ;
	LUT2 #(
		.INIT('h2)
	) name0 (
		\dest_x[22] ,
		\dest_x[23] ,
		_w62_
	);
	LUT4 #(
		.INIT('h0007)
	) name1 (
		\dest_x[14] ,
		\dest_x[15] ,
		\dest_x[16] ,
		\dest_x[18] ,
		_w63_
	);
	LUT3 #(
		.INIT('he0)
	) name2 (
		\dest_x[9] ,
		\dest_x[10] ,
		\dest_x[11] ,
		_w64_
	);
	LUT4 #(
		.INIT('h0001)
	) name3 (
		\dest_x[12] ,
		\dest_x[13] ,
		\dest_x[16] ,
		\dest_x[18] ,
		_w65_
	);
	LUT4 #(
		.INIT('he000)
	) name4 (
		\dest_x[17] ,
		\dest_x[18] ,
		\dest_x[19] ,
		\dest_x[20] ,
		_w66_
	);
	LUT4 #(
		.INIT('h4500)
	) name5 (
		_w63_,
		_w64_,
		_w65_,
		_w66_,
		_w67_
	);
	LUT2 #(
		.INIT('h1)
	) name6 (
		\dest_x[21] ,
		_w67_,
		_w68_
	);
	LUT4 #(
		.INIT('h8000)
	) name7 (
		\dest_x[6] ,
		\dest_x[7] ,
		\dest_x[8] ,
		\dest_x[11] ,
		_w69_
	);
	LUT4 #(
		.INIT('h8000)
	) name8 (
		\dest_x[2] ,
		\dest_x[3] ,
		\dest_x[4] ,
		\dest_x[5] ,
		_w70_
	);
	LUT2 #(
		.INIT('h2)
	) name9 (
		\dest_x[17] ,
		\dest_x[18] ,
		_w71_
	);
	LUT4 #(
		.INIT('h0008)
	) name10 (
		\dest_x[0] ,
		\dest_x[1] ,
		\dest_x[9] ,
		\dest_x[10] ,
		_w72_
	);
	LUT4 #(
		.INIT('h8000)
	) name11 (
		_w69_,
		_w70_,
		_w71_,
		_w72_,
		_w73_
	);
	LUT4 #(
		.INIT('h2000)
	) name12 (
		\dest_x[20] ,
		\dest_x[21] ,
		\dest_x[24] ,
		\dest_x[25] ,
		_w74_
	);
	LUT4 #(
		.INIT('h0040)
	) name13 (
		\dest_x[12] ,
		\dest_x[15] ,
		\dest_x[19] ,
		\dest_x[26] ,
		_w75_
	);
	LUT3 #(
		.INIT('h80)
	) name14 (
		\dest_x[27] ,
		\dest_x[28] ,
		\dest_x[29] ,
		_w76_
	);
	LUT3 #(
		.INIT('h80)
	) name15 (
		_w74_,
		_w75_,
		_w76_,
		_w77_
	);
	LUT3 #(
		.INIT('h07)
	) name16 (
		\dest_x[14] ,
		\dest_x[15] ,
		\dest_x[16] ,
		_w78_
	);
	LUT3 #(
		.INIT('h01)
	) name17 (
		\dest_x[12] ,
		\dest_x[13] ,
		\dest_x[16] ,
		_w79_
	);
	LUT3 #(
		.INIT('h23)
	) name18 (
		_w64_,
		_w78_,
		_w79_,
		_w80_
	);
	LUT3 #(
		.INIT('he0)
	) name19 (
		\dest_x[12] ,
		\dest_x[13] ,
		\dest_x[14] ,
		_w81_
	);
	LUT4 #(
		.INIT('he000)
	) name20 (
		\dest_x[9] ,
		\dest_x[10] ,
		\dest_x[11] ,
		\dest_x[14] ,
		_w82_
	);
	LUT4 #(
		.INIT('he000)
	) name21 (
		\dest_x[9] ,
		\dest_x[10] ,
		\dest_x[11] ,
		\dest_x[13] ,
		_w83_
	);
	LUT3 #(
		.INIT('h07)
	) name22 (
		\dest_x[12] ,
		\dest_x[13] ,
		\dest_x[14] ,
		_w84_
	);
	LUT4 #(
		.INIT('h1011)
	) name23 (
		_w81_,
		_w82_,
		_w83_,
		_w84_,
		_w85_
	);
	LUT4 #(
		.INIT('h0800)
	) name24 (
		_w73_,
		_w77_,
		_w80_,
		_w85_,
		_w86_
	);
	LUT3 #(
		.INIT('h10)
	) name25 (
		\dest_x[21] ,
		\dest_x[22] ,
		\dest_x[23] ,
		_w87_
	);
	LUT2 #(
		.INIT('h4)
	) name26 (
		_w67_,
		_w87_,
		_w88_
	);
	LUT4 #(
		.INIT('h0fdf)
	) name27 (
		_w62_,
		_w68_,
		_w86_,
		_w88_,
		_w89_
	);
	LUT4 #(
		.INIT('h007f)
	) name28 (
		\dest_x[23] ,
		\dest_x[24] ,
		\dest_x[25] ,
		\dest_x[26] ,
		_w90_
	);
	LUT2 #(
		.INIT('h1)
	) name29 (
		\dest_x[21] ,
		\dest_x[22] ,
		_w91_
	);
	LUT3 #(
		.INIT('h01)
	) name30 (
		\dest_x[21] ,
		\dest_x[22] ,
		\dest_x[26] ,
		_w92_
	);
	LUT4 #(
		.INIT('h080c)
	) name31 (
		_w67_,
		_w76_,
		_w90_,
		_w92_,
		_w93_
	);
	LUT3 #(
		.INIT('h8a)
	) name32 (
		\dest_x[23] ,
		_w67_,
		_w91_,
		_w94_
	);
	LUT3 #(
		.INIT('hc8)
	) name33 (
		\dest_x[21] ,
		\dest_x[22] ,
		_w67_,
		_w95_
	);
	LUT3 #(
		.INIT('h04)
	) name34 (
		\dest_x[7] ,
		\dest_x[9] ,
		\dest_x[10] ,
		_w96_
	);
	LUT4 #(
		.INIT('h0004)
	) name35 (
		\dest_x[8] ,
		\dest_x[11] ,
		\dest_x[12] ,
		\dest_x[13] ,
		_w97_
	);
	LUT3 #(
		.INIT('h80)
	) name36 (
		_w74_,
		_w96_,
		_w97_,
		_w98_
	);
	LUT4 #(
		.INIT('h0010)
	) name37 (
		\dest_x[1] ,
		\dest_x[2] ,
		\dest_x[17] ,
		\dest_x[18] ,
		_w99_
	);
	LUT4 #(
		.INIT('h0001)
	) name38 (
		\dest_x[3] ,
		\dest_x[4] ,
		\dest_x[5] ,
		\dest_x[6] ,
		_w100_
	);
	LUT2 #(
		.INIT('h8)
	) name39 (
		_w99_,
		_w100_,
		_w101_
	);
	LUT3 #(
		.INIT('h01)
	) name40 (
		\dest_x[12] ,
		\dest_x[14] ,
		\dest_x[15] ,
		_w102_
	);
	LUT3 #(
		.INIT('h8a)
	) name41 (
		\dest_x[16] ,
		_w64_,
		_w102_,
		_w103_
	);
	LUT4 #(
		.INIT('h0080)
	) name42 (
		_w80_,
		_w98_,
		_w101_,
		_w103_,
		_w104_
	);
	LUT3 #(
		.INIT('he0)
	) name43 (
		\dest_x[17] ,
		\dest_x[18] ,
		\dest_x[19] ,
		_w105_
	);
	LUT4 #(
		.INIT('h4500)
	) name44 (
		_w63_,
		_w64_,
		_w65_,
		_w105_,
		_w106_
	);
	LUT4 #(
		.INIT('h8000)
	) name45 (
		\dest_x[23] ,
		\dest_x[24] ,
		\dest_x[25] ,
		\dest_x[26] ,
		_w107_
	);
	LUT2 #(
		.INIT('h2)
	) name46 (
		_w106_,
		_w107_,
		_w108_
	);
	LUT4 #(
		.INIT('h2000)
	) name47 (
		_w94_,
		_w95_,
		_w104_,
		_w108_,
		_w109_
	);
	LUT2 #(
		.INIT('h2)
	) name48 (
		_w93_,
		_w109_,
		_w110_
	);
	LUT3 #(
		.INIT('hd1)
	) name49 (
		_w89_,
		_w93_,
		_w109_,
		_w111_
	);
	LUT3 #(
		.INIT('h2e)
	) name50 (
		_w89_,
		_w93_,
		_w109_,
		_w112_
	);
	LUT3 #(
		.INIT('h80)
	) name51 (
		\dest_y[23] ,
		\dest_y[24] ,
		\dest_y[25] ,
		_w113_
	);
	LUT4 #(
		.INIT('h007f)
	) name52 (
		\dest_y[23] ,
		\dest_y[24] ,
		\dest_y[25] ,
		\dest_y[26] ,
		_w114_
	);
	LUT4 #(
		.INIT('h0007)
	) name53 (
		\dest_y[14] ,
		\dest_y[15] ,
		\dest_y[16] ,
		\dest_y[18] ,
		_w115_
	);
	LUT3 #(
		.INIT('he0)
	) name54 (
		\dest_y[9] ,
		\dest_y[10] ,
		\dest_y[11] ,
		_w116_
	);
	LUT4 #(
		.INIT('h0001)
	) name55 (
		\dest_y[12] ,
		\dest_y[13] ,
		\dest_y[16] ,
		\dest_y[18] ,
		_w117_
	);
	LUT4 #(
		.INIT('he000)
	) name56 (
		\dest_y[17] ,
		\dest_y[18] ,
		\dest_y[19] ,
		\dest_y[20] ,
		_w118_
	);
	LUT4 #(
		.INIT('h4500)
	) name57 (
		_w115_,
		_w116_,
		_w117_,
		_w118_,
		_w119_
	);
	LUT2 #(
		.INIT('h1)
	) name58 (
		\dest_y[21] ,
		\dest_y[22] ,
		_w120_
	);
	LUT3 #(
		.INIT('h01)
	) name59 (
		\dest_y[21] ,
		\dest_y[22] ,
		\dest_y[26] ,
		_w121_
	);
	LUT3 #(
		.INIT('h80)
	) name60 (
		\dest_y[27] ,
		\dest_y[28] ,
		\dest_y[29] ,
		_w122_
	);
	LUT4 #(
		.INIT('h4500)
	) name61 (
		_w114_,
		_w119_,
		_w121_,
		_w122_,
		_w123_
	);
	LUT2 #(
		.INIT('h2)
	) name62 (
		\dest_x[0] ,
		_w123_,
		_w124_
	);
	LUT4 #(
		.INIT('hf322)
	) name63 (
		_w89_,
		_w93_,
		_w109_,
		_w124_,
		_w125_
	);
	LUT3 #(
		.INIT('he0)
	) name64 (
		\dest_y[17] ,
		\dest_y[18] ,
		\dest_y[19] ,
		_w126_
	);
	LUT4 #(
		.INIT('h4500)
	) name65 (
		_w115_,
		_w116_,
		_w117_,
		_w126_,
		_w127_
	);
	LUT2 #(
		.INIT('h8)
	) name66 (
		\dest_y[12] ,
		\dest_y[13] ,
		_w128_
	);
	LUT4 #(
		.INIT('he000)
	) name67 (
		\dest_y[9] ,
		\dest_y[10] ,
		\dest_y[11] ,
		\dest_y[13] ,
		_w129_
	);
	LUT4 #(
		.INIT('h0400)
	) name68 (
		\dest_y[18] ,
		\dest_y[19] ,
		\dest_y[22] ,
		\dest_y[23] ,
		_w130_
	);
	LUT4 #(
		.INIT('h0020)
	) name69 (
		\dest_y[11] ,
		\dest_y[12] ,
		\dest_y[15] ,
		\dest_y[16] ,
		_w131_
	);
	LUT4 #(
		.INIT('h1000)
	) name70 (
		_w128_,
		_w129_,
		_w130_,
		_w131_,
		_w132_
	);
	LUT4 #(
		.INIT('h0001)
	) name71 (
		\dest_y[5] ,
		\dest_y[6] ,
		\dest_y[7] ,
		\dest_y[8] ,
		_w133_
	);
	LUT4 #(
		.INIT('h0001)
	) name72 (
		\dest_y[1] ,
		\dest_y[2] ,
		\dest_y[3] ,
		\dest_y[4] ,
		_w134_
	);
	LUT3 #(
		.INIT('h20)
	) name73 (
		\dest_y[9] ,
		\dest_y[10] ,
		\dest_y[17] ,
		_w135_
	);
	LUT3 #(
		.INIT('h80)
	) name74 (
		_w133_,
		_w134_,
		_w135_,
		_w136_
	);
	LUT3 #(
		.INIT('he0)
	) name75 (
		\dest_y[12] ,
		\dest_y[13] ,
		\dest_y[14] ,
		_w137_
	);
	LUT4 #(
		.INIT('he000)
	) name76 (
		\dest_y[9] ,
		\dest_y[10] ,
		\dest_y[11] ,
		\dest_y[14] ,
		_w138_
	);
	LUT2 #(
		.INIT('h4)
	) name77 (
		\dest_y[20] ,
		\dest_y[21] ,
		_w139_
	);
	LUT3 #(
		.INIT('he0)
	) name78 (
		_w137_,
		_w138_,
		_w139_,
		_w140_
	);
	LUT4 #(
		.INIT('h4000)
	) name79 (
		_w127_,
		_w132_,
		_w136_,
		_w140_,
		_w141_
	);
	LUT3 #(
		.INIT('ha8)
	) name80 (
		\dest_y[20] ,
		_w137_,
		_w138_,
		_w142_
	);
	LUT3 #(
		.INIT('h80)
	) name81 (
		_w132_,
		_w136_,
		_w142_,
		_w143_
	);
	LUT2 #(
		.INIT('h4)
	) name82 (
		\dest_y[21] ,
		_w127_,
		_w144_
	);
	LUT4 #(
		.INIT('h9399)
	) name83 (
		\dest_y[23] ,
		\dest_y[24] ,
		_w119_,
		_w120_,
		_w145_
	);
	LUT4 #(
		.INIT('hea00)
	) name84 (
		_w141_,
		_w143_,
		_w144_,
		_w145_,
		_w146_
	);
	LUT4 #(
		.INIT('h8000)
	) name85 (
		\dest_y[23] ,
		\dest_y[24] ,
		\dest_y[25] ,
		\dest_y[26] ,
		_w147_
	);
	LUT2 #(
		.INIT('h1)
	) name86 (
		\dest_x[0] ,
		\dest_y[0] ,
		_w148_
	);
	LUT4 #(
		.INIT('h4f00)
	) name87 (
		_w119_,
		_w120_,
		_w147_,
		_w148_,
		_w149_
	);
	LUT3 #(
		.INIT('h8a)
	) name88 (
		_w113_,
		_w119_,
		_w120_,
		_w150_
	);
	LUT2 #(
		.INIT('h8)
	) name89 (
		\dest_y[23] ,
		\dest_y[24] ,
		_w151_
	);
	LUT3 #(
		.INIT('h07)
	) name90 (
		\dest_y[23] ,
		\dest_y[24] ,
		\dest_y[25] ,
		_w152_
	);
	LUT3 #(
		.INIT('h01)
	) name91 (
		\dest_y[21] ,
		\dest_y[22] ,
		\dest_y[25] ,
		_w153_
	);
	LUT3 #(
		.INIT('h23)
	) name92 (
		_w119_,
		_w152_,
		_w153_,
		_w154_
	);
	LUT3 #(
		.INIT('h8a)
	) name93 (
		_w149_,
		_w150_,
		_w154_,
		_w155_
	);
	LUT3 #(
		.INIT('h2a)
	) name94 (
		_w123_,
		_w146_,
		_w155_,
		_w156_
	);
	LUT4 #(
		.INIT('h1055)
	) name95 (
		\dest_y[27] ,
		_w119_,
		_w120_,
		_w147_,
		_w157_
	);
	LUT3 #(
		.INIT('hb0)
	) name96 (
		_w119_,
		_w120_,
		_w151_,
		_w158_
	);
	LUT2 #(
		.INIT('h1)
	) name97 (
		\dest_y[20] ,
		_w127_,
		_w159_
	);
	LUT2 #(
		.INIT('h1)
	) name98 (
		_w158_,
		_w159_,
		_w160_
	);
	LUT2 #(
		.INIT('h1)
	) name99 (
		\dest_y[23] ,
		\dest_y[24] ,
		_w161_
	);
	LUT3 #(
		.INIT('h01)
	) name100 (
		\dest_y[21] ,
		\dest_y[22] ,
		\dest_y[24] ,
		_w162_
	);
	LUT3 #(
		.INIT('h23)
	) name101 (
		_w119_,
		_w161_,
		_w162_,
		_w163_
	);
	LUT3 #(
		.INIT('h01)
	) name102 (
		\dest_y[17] ,
		_w137_,
		_w138_,
		_w164_
	);
	LUT4 #(
		.INIT('h1000)
	) name103 (
		\dest_y[9] ,
		\dest_y[10] ,
		\dest_y[28] ,
		\dest_y[29] ,
		_w165_
	);
	LUT4 #(
		.INIT('h0020)
	) name104 (
		\dest_y[8] ,
		\dest_y[13] ,
		\dest_y[14] ,
		\dest_y[21] ,
		_w166_
	);
	LUT4 #(
		.INIT('h8000)
	) name105 (
		\dest_y[4] ,
		\dest_y[5] ,
		\dest_y[6] ,
		\dest_y[7] ,
		_w167_
	);
	LUT3 #(
		.INIT('h80)
	) name106 (
		_w165_,
		_w166_,
		_w167_,
		_w168_
	);
	LUT4 #(
		.INIT('h8000)
	) name107 (
		\dest_y[0] ,
		\dest_y[1] ,
		\dest_y[2] ,
		\dest_y[3] ,
		_w169_
	);
	LUT3 #(
		.INIT('h80)
	) name108 (
		_w130_,
		_w131_,
		_w169_,
		_w170_
	);
	LUT3 #(
		.INIT('h40)
	) name109 (
		_w164_,
		_w168_,
		_w170_,
		_w171_
	);
	LUT3 #(
		.INIT('ha8)
	) name110 (
		\dest_y[17] ,
		_w137_,
		_w138_,
		_w172_
	);
	LUT2 #(
		.INIT('h1)
	) name111 (
		_w119_,
		_w172_,
		_w173_
	);
	LUT3 #(
		.INIT('h80)
	) name112 (
		_w163_,
		_w171_,
		_w173_,
		_w174_
	);
	LUT4 #(
		.INIT('h2022)
	) name113 (
		\dest_y[27] ,
		_w114_,
		_w119_,
		_w121_,
		_w175_
	);
	LUT3 #(
		.INIT('h04)
	) name114 (
		_w150_,
		_w154_,
		_w175_,
		_w176_
	);
	LUT4 #(
		.INIT('h4000)
	) name115 (
		_w157_,
		_w160_,
		_w174_,
		_w176_,
		_w177_
	);
	LUT4 #(
		.INIT('hcccd)
	) name116 (
		_w110_,
		_w125_,
		_w156_,
		_w177_,
		_w178_
	);
	LUT2 #(
		.INIT('h8)
	) name117 (
		\dest_x[0] ,
		\dest_y[0] ,
		_w179_
	);
	LUT4 #(
		.INIT('h004f)
	) name118 (
		_w119_,
		_w120_,
		_w147_,
		_w179_,
		_w180_
	);
	LUT3 #(
		.INIT('hb0)
	) name119 (
		_w150_,
		_w154_,
		_w180_,
		_w181_
	);
	LUT3 #(
		.INIT('h2a)
	) name120 (
		_w123_,
		_w146_,
		_w181_,
		_w182_
	);
	LUT2 #(
		.INIT('h8)
	) name121 (
		_w111_,
		_w182_,
		_w183_
	);
	assign \outport[0]  = _w112_ ;
	assign \outport[1]  = _w178_ ;
	assign \outport[2]  = _w183_ ;
	assign \outport[3]  = 1'b0;
	assign \outport[4]  = 1'b0;
	assign \outport[5]  = 1'b0;
	assign \outport[6]  = 1'b0;
	assign \outport[7]  = 1'b0;
	assign \outport[8]  = 1'b0;
	assign \outport[9]  = 1'b0;
	assign \outport[10]  = 1'b0;
	assign \outport[11]  = 1'b0;
	assign \outport[12]  = 1'b0;
	assign \outport[13]  = 1'b0;
	assign \outport[14]  = 1'b0;
	assign \outport[15]  = 1'b0;
	assign \outport[16]  = 1'b0;
	assign \outport[17]  = 1'b0;
	assign \outport[18]  = 1'b0;
	assign \outport[19]  = 1'b0;
	assign \outport[20]  = 1'b0;
	assign \outport[21]  = 1'b0;
	assign \outport[22]  = 1'b0;
	assign \outport[23]  = 1'b0;
	assign \outport[24]  = 1'b0;
	assign \outport[25]  = 1'b0;
	assign \outport[26]  = 1'b0;
	assign \outport[27]  = 1'b0;
	assign \outport[28]  = 1'b0;
	assign \outport[29]  = 1'b0;
endmodule;