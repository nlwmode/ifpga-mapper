module top( \a0_pad  , a_pad , \b0_pad  , b_pad , \c0_pad  , c_pad , \d0_pad  , d_pad , \e0_pad  , e_pad , \f0_pad  , f_pad , \g0_pad  , g_pad , h_pad , i_pad , j_pad , k_pad , l_pad , m_pad , n_pad , o_pad , p_pad , q_pad , r_pad , s_pad , t_pad , u_pad , v_pad , w_pad , x_pad , y_pad , z_pad , \h0_pad  , \i0_pad  , \j0_pad  , \k0_pad  , \l0_pad  , \m0_pad  , \n0_pad  , \o0_pad  , \p0_pad  , \q0_pad  , \r0_pad  , \s0_pad  , \t0_pad  , \u0_pad  , \v0_pad  , \w0_pad  , \x0_pad  );
  input \a0_pad  ;
  input a_pad ;
  input \b0_pad  ;
  input b_pad ;
  input \c0_pad  ;
  input c_pad ;
  input \d0_pad  ;
  input d_pad ;
  input \e0_pad  ;
  input e_pad ;
  input \f0_pad  ;
  input f_pad ;
  input \g0_pad  ;
  input g_pad ;
  input h_pad ;
  input i_pad ;
  input j_pad ;
  input k_pad ;
  input l_pad ;
  input m_pad ;
  input n_pad ;
  input o_pad ;
  input p_pad ;
  input q_pad ;
  input r_pad ;
  input s_pad ;
  input t_pad ;
  input u_pad ;
  input v_pad ;
  input w_pad ;
  input x_pad ;
  input y_pad ;
  input z_pad ;
  output \h0_pad  ;
  output \i0_pad  ;
  output \j0_pad  ;
  output \k0_pad  ;
  output \l0_pad  ;
  output \m0_pad  ;
  output \n0_pad  ;
  output \o0_pad  ;
  output \p0_pad  ;
  output \q0_pad  ;
  output \r0_pad  ;
  output \s0_pad  ;
  output \t0_pad  ;
  output \u0_pad  ;
  output \v0_pad  ;
  output \w0_pad  ;
  output \x0_pad  ;
  wire n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 ;
  assign n34 = ~c_pad & ~s_pad ;
  assign n35 = c_pad & s_pad ;
  assign n36 = d_pad & t_pad ;
  assign n37 = ~n35 & ~n36 ;
  assign n38 = ~n34 & ~n37 ;
  assign n39 = e_pad & u_pad ;
  assign n40 = ~f_pad & ~v_pad ;
  assign n41 = ~n39 & n40 ;
  assign n42 = ~g_pad & ~w_pad ;
  assign n43 = ~h_pad & ~x_pad ;
  assign n44 = ~n42 & ~n43 ;
  assign n45 = h_pad & x_pad ;
  assign n46 = n44 & n45 ;
  assign n47 = ~\c0_pad  & ~m_pad ;
  assign n48 = ~\d0_pad  & ~n_pad ;
  assign n49 = ~n47 & ~n48 ;
  assign n50 = \d0_pad  & n_pad ;
  assign n51 = n49 & n50 ;
  assign n52 = ~\f0_pad  & ~p_pad ;
  assign n53 = \g0_pad  & ~n52 ;
  assign n54 = \e0_pad  & o_pad ;
  assign n55 = \f0_pad  & p_pad ;
  assign n56 = ~n54 & ~n55 ;
  assign n57 = ~n53 & n56 ;
  assign n58 = ~\e0_pad  & ~o_pad ;
  assign n59 = n49 & ~n58 ;
  assign n60 = ~n57 & n59 ;
  assign n61 = ~n51 & ~n60 ;
  assign n62 = \b0_pad  & l_pad ;
  assign n63 = \c0_pad  & m_pad ;
  assign n64 = ~n62 & ~n63 ;
  assign n65 = n61 & n64 ;
  assign n66 = ~\b0_pad  & ~l_pad ;
  assign n67 = ~j_pad & ~z_pad ;
  assign n68 = ~\a0_pad  & ~k_pad ;
  assign n69 = ~n67 & ~n68 ;
  assign n70 = ~n66 & n69 ;
  assign n71 = ~n65 & n70 ;
  assign n72 = \a0_pad  & k_pad ;
  assign n73 = ~n67 & n72 ;
  assign n74 = i_pad & y_pad ;
  assign n75 = j_pad & z_pad ;
  assign n76 = ~n74 & ~n75 ;
  assign n77 = ~n73 & n76 ;
  assign n78 = ~n71 & n77 ;
  assign n79 = ~i_pad & ~y_pad ;
  assign n80 = n44 & ~n79 ;
  assign n81 = ~n78 & n80 ;
  assign n82 = ~n46 & ~n81 ;
  assign n83 = f_pad & v_pad ;
  assign n84 = g_pad & w_pad ;
  assign n85 = ~n83 & ~n84 ;
  assign n86 = ~n39 & n85 ;
  assign n87 = n82 & n86 ;
  assign n88 = ~n41 & ~n87 ;
  assign n89 = ~d_pad & ~t_pad ;
  assign n90 = ~e_pad & ~u_pad ;
  assign n91 = ~n89 & ~n90 ;
  assign n92 = ~n34 & n91 ;
  assign n93 = n88 & n92 ;
  assign n94 = ~n38 & ~n93 ;
  assign n95 = ~b_pad & ~r_pad ;
  assign n96 = ~n94 & ~n95 ;
  assign n97 = ~a_pad & ~q_pad ;
  assign n98 = a_pad & q_pad ;
  assign n99 = ~n97 & ~n98 ;
  assign n100 = b_pad & r_pad ;
  assign n101 = ~n99 & ~n100 ;
  assign n102 = ~n96 & n101 ;
  assign n103 = ~n95 & n99 ;
  assign n104 = ~n94 & n103 ;
  assign n105 = n99 & n100 ;
  assign n106 = ~n104 & ~n105 ;
  assign n107 = ~n102 & n106 ;
  assign n108 = ~n95 & ~n100 ;
  assign n109 = ~n94 & n108 ;
  assign n110 = n94 & ~n108 ;
  assign n111 = ~n109 & ~n110 ;
  assign n112 = ~n34 & ~n35 ;
  assign n113 = n36 & ~n112 ;
  assign n114 = n91 & ~n112 ;
  assign n115 = n88 & n114 ;
  assign n116 = ~n113 & ~n115 ;
  assign n117 = n88 & n91 ;
  assign n118 = ~n36 & n112 ;
  assign n119 = ~n117 & n118 ;
  assign n120 = n116 & ~n119 ;
  assign n121 = ~n36 & ~n89 ;
  assign n122 = ~n90 & n121 ;
  assign n123 = n88 & n122 ;
  assign n124 = n82 & n85 ;
  assign n125 = ~n40 & ~n90 ;
  assign n126 = ~n124 & n125 ;
  assign n127 = ~n39 & ~n121 ;
  assign n128 = ~n126 & n127 ;
  assign n129 = ~n123 & ~n128 ;
  assign n130 = ~n39 & ~n90 ;
  assign n131 = ~n40 & n130 ;
  assign n132 = ~n124 & n131 ;
  assign n133 = n40 & ~n130 ;
  assign n134 = n85 & ~n130 ;
  assign n135 = n82 & n134 ;
  assign n136 = ~n133 & ~n135 ;
  assign n137 = ~n132 & n136 ;
  assign n138 = n82 & ~n84 ;
  assign n139 = ~n40 & ~n83 ;
  assign n140 = ~n138 & ~n139 ;
  assign n141 = ~n84 & n139 ;
  assign n142 = n82 & n141 ;
  assign n143 = ~n140 & ~n142 ;
  assign n144 = ~n78 & ~n79 ;
  assign n145 = ~n45 & ~n144 ;
  assign n146 = ~n42 & ~n84 ;
  assign n147 = ~n43 & n146 ;
  assign n148 = ~n145 & n147 ;
  assign n149 = ~n43 & ~n79 ;
  assign n150 = ~n78 & n149 ;
  assign n151 = ~n45 & ~n146 ;
  assign n152 = ~n150 & n151 ;
  assign n153 = ~n148 & ~n152 ;
  assign n154 = ~n43 & ~n45 ;
  assign n155 = ~n79 & n154 ;
  assign n156 = ~n78 & n155 ;
  assign n157 = ~n144 & ~n154 ;
  assign n158 = ~n156 & ~n157 ;
  assign n159 = ~n73 & ~n75 ;
  assign n160 = ~n71 & n159 ;
  assign n161 = ~n74 & ~n79 ;
  assign n162 = ~n160 & ~n161 ;
  assign n163 = n159 & n161 ;
  assign n164 = ~n71 & n163 ;
  assign n165 = ~n162 & ~n164 ;
  assign n166 = ~n67 & ~n75 ;
  assign n167 = ~n68 & n166 ;
  assign n168 = n66 & ~n72 ;
  assign n169 = n64 & ~n72 ;
  assign n170 = n61 & n169 ;
  assign n171 = ~n168 & ~n170 ;
  assign n172 = n167 & n171 ;
  assign n173 = ~n66 & ~n68 ;
  assign n174 = ~n65 & n173 ;
  assign n175 = ~n72 & ~n166 ;
  assign n176 = ~n174 & n175 ;
  assign n177 = ~n172 & ~n176 ;
  assign n178 = ~n68 & ~n72 ;
  assign n179 = ~n66 & n178 ;
  assign n180 = ~n65 & n179 ;
  assign n181 = n66 & ~n178 ;
  assign n182 = n64 & ~n178 ;
  assign n183 = n61 & n182 ;
  assign n184 = ~n181 & ~n183 ;
  assign n185 = ~n180 & n184 ;
  assign n186 = n61 & ~n63 ;
  assign n187 = ~n62 & ~n66 ;
  assign n188 = ~n186 & ~n187 ;
  assign n189 = ~n63 & n187 ;
  assign n190 = n61 & n189 ;
  assign n191 = ~n188 & ~n190 ;
  assign n192 = ~n57 & ~n58 ;
  assign n193 = ~n50 & ~n192 ;
  assign n194 = ~n47 & ~n63 ;
  assign n195 = ~n48 & n194 ;
  assign n196 = ~n193 & n195 ;
  assign n197 = ~n48 & ~n58 ;
  assign n198 = ~n57 & n197 ;
  assign n199 = ~n50 & ~n194 ;
  assign n200 = ~n198 & n199 ;
  assign n201 = ~n196 & ~n200 ;
  assign n202 = ~n48 & ~n50 ;
  assign n203 = ~n58 & n202 ;
  assign n204 = ~n57 & n203 ;
  assign n205 = ~n192 & ~n202 ;
  assign n206 = ~n204 & ~n205 ;
  assign n207 = ~n53 & ~n55 ;
  assign n208 = ~n54 & ~n58 ;
  assign n209 = ~n207 & ~n208 ;
  assign n210 = n207 & n208 ;
  assign n211 = ~n209 & ~n210 ;
  assign n212 = ~n52 & ~n55 ;
  assign n213 = ~\g0_pad  & ~n212 ;
  assign n214 = \g0_pad  & n212 ;
  assign n215 = ~n213 & ~n214 ;
  assign n216 = ~n95 & ~n97 ;
  assign n217 = ~n98 & ~n216 ;
  assign n218 = ~n98 & ~n100 ;
  assign n219 = n94 & n218 ;
  assign n220 = ~n217 & ~n219 ;
  assign \h0_pad  = n107 ;
  assign \i0_pad  = n111 ;
  assign \j0_pad  = ~n120 ;
  assign \k0_pad  = n129 ;
  assign \l0_pad  = n137 ;
  assign \m0_pad  = ~n143 ;
  assign \n0_pad  = n153 ;
  assign \o0_pad  = n158 ;
  assign \p0_pad  = ~n165 ;
  assign \q0_pad  = n177 ;
  assign \r0_pad  = n185 ;
  assign \s0_pad  = ~n191 ;
  assign \t0_pad  = n201 ;
  assign \u0_pad  = n206 ;
  assign \v0_pad  = ~n211 ;
  assign \w0_pad  = n215 ;
  assign \x0_pad  = n220 ;
endmodule
