module top (\g1002_reg/NET0131 , \g1008_reg/NET0131 , \g10122_pad , \g1018_reg/NET0131 , \g1024_reg/NET0131 , \g10306_pad , \g1030_reg/NET0131 , \g1036_reg/NET0131 , \g1041_reg/NET0131 , \g1046_reg/NET0131 , \g10500_pad , \g10527_pad , \g1052_reg/NET0131 , \g1061_reg/NET0131 , \g1070_reg/NET0131 , \g1087_reg/NET0131 , \g1094_reg/NET0131 , \g1099_reg/NET0131 , \g1105_reg/NET0131 , \g1111_reg/NET0131 , \g1124_reg/NET0131 , \g1129_reg/NET0131 , \g1135_reg/NET0131 , \g1141_reg/NET0131 , \g11447_pad , \g1146_reg/NET0131 , \g1152_reg/NET0131 , \g1171_reg/NET0131 , \g11770_pad , \g1178_reg/NET0131 , \g1183_reg/NET0131 , \g1189_reg/NET0131 , \g1193_reg/NET0131 , \g1199_reg/NET0131 , \g1205_reg/NET0131 , \g1211_reg/NET0131 , \g1216_reg/NET0131 , \g12184_pad , \g1221_reg/NET0131 , \g1236_reg/NET0131 , \g1242_reg/NET0131 , \g1246_reg/NET0131 , \g12919_pad , \g12923_pad , \g1300_reg/NET0131 , \g13039_pad , \g1306_reg/NET0131 , \g1312_reg/NET0131 , \g1319_reg/NET0131 , \g1322_reg/NET0131 , \g13259_pad , \g13272_pad , \g1333_reg/NET0131 , \g1339_reg/NET0131 , \g1345_reg/NET0131 , \g1351_reg/NET0131 , \g1361_reg/NET0131 , \g1367_reg/NET0131 , \g1373_reg/NET0131 , \g1379_reg/NET0131 , \g1384_reg/NET0131 , \g13865_pad , \g13895_pad , \g1389_reg/NET0131 , \g1395_reg/NET0131 , \g1404_reg/NET0131 , \g14096_pad , \g14125_pad , \g1413_reg/NET0131 , \g14147_pad , \g14167_pad , \g14189_pad , \g14201_pad , \g14217_pad , \g142_reg/NET0131 , \g1430_reg/NET0131 , \g1437_reg/NET0131 , \g1442_reg/NET0131 , \g1448_reg/NET0131 , \g1454_reg/NET0131 , \g1467_reg/NET0131 , \g146_reg/NET0131 , \g1472_reg/NET0131 , \g1478_reg/NET0131 , \g1484_reg/NET0131 , \g1489_reg/NET0131 , \g1495_reg/NET0131 , \g150_reg/NET0131 , \g1514_reg/NET0131 , \g1521_reg/NET0131 , \g1526_reg/NET0131 , \g1532_reg/NET0131 , \g1536_reg/NET0131 , \g153_reg/NET0131 , \g1542_reg/NET0131 , \g1548_reg/NET0131 , \g1554_reg/NET0131 , \g1559_reg/NET0131 , \g1564_reg/NET0131 , \g1579_reg/NET0131 , \g157_reg/NET0131 , \g1585_reg/NET0131 , \g1589_reg/NET0131 , \g1592_reg/NET0131 , \g1600_reg/NET0131 , \g1604_reg/NET0131 , \g1608_reg/NET0131 , \g160_reg/NET0131 , \g1612_reg/NET0131 , \g1616_reg/NET0131 , \g1620_reg/NET0131 , \g1624_reg/NET0131 , \g1632_reg/NET0131 , \g1636_reg/NET0131 , \g1644_reg/NET0131 , \g1648_reg/NET0131 , \g164_reg/NET0131 , \g1657_reg/NET0131 , \g16603_pad , \g16624_pad , \g1664_reg/NET0131 , \g16686_pad , \g1668_reg/NET0131 , \g16718_pad , \g1677_reg/NET0131 , \g1682_reg/NET0131 , \g16874_pad , \g1687_reg/NET0131 , \g168_reg/NET0131 , \g1691_reg/NET0131 , \g1696_reg/NET0131 , \g1700_reg/NET0131 , \g1706_reg/NET0131 , \g1710_reg/NET0131 , \g1714_reg/NET0131 , \g1720_reg/NET0131 , \g1724_reg/NET0131 , \g1728_reg/NET0131 , \g17291_pad , \g17316_pad , \g17320_pad , \g1736_reg/NET0131 , \g17400_pad , \g17404_pad , \g1740_reg/NET0131 , \g17423_pad , \g1744_reg/NET0131 , \g1748_reg/NET0131 , \g174_reg/NET0131 , \g1752_reg/NET0131 , \g1756_reg/NET0131 , \g1760_reg/NET0131 , \g1768_reg/NET0131 , \g1772_reg/NET0131 , \g1779_reg/NET0131 , \g1783_reg/NET0131 , \g1792_reg/NET0131 , \g1798_reg/NET0131 , \g1802_reg/NET0131 , \g18094_pad , \g18095_pad , \g18096_pad , \g18098_pad , \g18099_pad , \g1811_reg/NET0131 , \g1816_reg/NET0131 , \g1821_reg/NET0131 , \g1825_reg/NET0131 , \g182_reg/NET0131 , \g1830_reg/NET0131 , \g1834_reg/NET0131 , \g1840_reg/NET0131 , \g1844_reg/NET0131 , \g1848_reg/NET0131 , \g1854_reg/NET0131 , \g1858_reg/NET0131 , \g1862_reg/NET0131 , \g1870_reg/NET0131 , \g1874_reg/NET0131 , \g1878_reg/NET0131 , \g1882_reg/NET0131 , \g1886_reg/NET0131 , \g1890_reg/NET0131 , \g1894_reg/NET0131 , \g1902_reg/NET0131 , \g1906_reg/NET0131 , \g1913_reg/NET0131 , \g1917_reg/NET0131 , \g191_reg/NET0131 , \g1926_reg/NET0131 , \g1932_reg/NET0131 , \g19334_pad , \g19357_pad , \g1936_reg/NET0131 , \g1945_reg/NET0131 , \g1950_reg/NET0131 , \g1955_reg/NET0131 , \g1959_reg/NET0131 , \g1964_reg/NET0131 , \g1968_reg/NET0131 , \g1974_reg/NET0131 , \g1978_reg/NET0131 , \g1982_reg/NET0131 , \g1988_reg/NET0131 , \g1992_reg/NET0131 , \g1996_reg/NET0131 , \g2004_reg/NET0131 , \g2008_reg/NET0131 , \g2012_reg/NET0131 , \g2016_reg/NET0131 , \g2020_reg/NET0131 , \g2024_reg/NET0131 , \g2028_reg/NET0131 , \g2036_reg/NET0131 , \g203_reg/NET0131 , \g2040_reg/NET0131 , \g2047_reg/NET0131 , \g2051_reg/NET0131 , \g2060_reg/NET0131 , \g2066_reg/NET0131 , \g2070_reg/NET0131 , \g2079_reg/NET0131 , \g2084_reg/NET0131 , \g2089_reg/NET0131 , \g2093_reg/NET0131 , \g2098_reg/NET0131 , \g209_reg/NET0131 , \g2102_reg/NET0131 , \g2108_reg/NET0131 , \g2112_reg/NET0131 , \g2116_reg/NET0131 , \g2122_reg/NET0131 , \g2126_reg/NET0131 , \g2153_reg/NET0131 , \g2161_reg/NET0131 , \g2165_reg/NET0131 , \g2169_reg/NET0131 , \g2173_reg/NET0131 , \g2177_reg/NET0131 , \g2181_reg/NET0131 , \g2185_reg/NET0131 , \g218_reg/NET0131 , \g2193_reg/NET0131 , \g2197_reg/NET0131 , \g2204_reg/NET0131 , \g2208_reg/NET0131 , \g2217_reg/NET0131 , \g2223_reg/NET0131 , \g2227_reg/NET0131 , \g222_reg/NET0131 , \g2236_reg/NET0131 , \g2241_reg/NET0131 , \g2246_reg/NET0131 , \g2250_reg/NET0131 , \g2255_reg/NET0131 , \g2259_reg/NET0131 , \g225_reg/NET0131 , \g2265_reg/NET0131 , \g2269_reg/NET0131 , \g2273_reg/NET0131 , \g2279_reg/NET0131 , \g2283_reg/NET0131 , \g2287_reg/NET0131 , \g2295_reg/NET0131 , \g2299_reg/NET0131 , \g2303_reg/NET0131 , \g2307_reg/NET0131 , \g2311_reg/NET0131 , \g2315_reg/NET0131 , \g2319_reg/NET0131 , \g2327_reg/NET0131 , \g232_reg/NET0131 , \g2331_reg/NET0131 , \g2338_reg/NET0131 , \g2342_reg/NET0131 , \g2351_reg/NET0131 , \g2357_reg/NET0131 , \g2361_reg/NET0131 , \g2370_reg/NET0131 , \g2375_reg/NET0131 , \g2380_reg/NET0131 , \g2384_reg/NET0131 , \g2389_reg/NET0131 , \g2393_reg/NET0131 , \g2399_reg/NET0131 , \g239_reg/NET0131 , \g2403_reg/NET0131 , \g2407_reg/NET0131 , \g2413_reg/NET0131 , \g2417_reg/NET0131 , \g2421_reg/NET0131 , \g2429_reg/NET0131 , \g2433_reg/NET0131 , \g2437_reg/NET0131 , \g2441_reg/NET0131 , \g2445_reg/NET0131 , \g2449_reg/NET0131 , \g2453_reg/NET0131 , \g2461_reg/NET0131 , \g2465_reg/NET0131 , \g246_reg/NET0131 , \g2472_reg/NET0131 , \g2476_reg/NET0131 , \g2485_reg/NET0131 , \g2491_reg/NET0131 , \g2495_reg/NET0131 , \g2504_reg/NET0131 , \g2509_reg/NET0131 , \g2514_reg/NET0131 , \g2518_reg/NET0131 , \g2523_reg/NET0131 , \g2527_reg/NET0131 , \g2533_reg/NET0131 , \g2537_reg/NET0131 , \g2541_reg/NET0131 , \g2547_reg/NET0131 , \g2551_reg/NET0131 , \g2555_reg/NET0131 , \g255_reg/NET0131 , \g2563_reg/NET0131 , \g2567_reg/NET0131 , \g2571_reg/NET0131 , \g2575_reg/NET0131 , \g2579_reg/NET0131 , \g2583_reg/NET0131 , \g2587_reg/NET0131 , \g2595_reg/NET0131 , \g2599_reg/NET0131 , \g2606_reg/NET0131 , \g2610_reg/NET0131 , \g2619_reg/NET0131 , \g2625_reg/NET0131 , \g2629_reg/NET0131 , \g262_reg/NET0131 , \g2638_reg/NET0131 , \g2643_reg/NET0131 , \g2648_reg/NET0131 , \g2652_reg/NET0131 , \g2657_reg/NET0131 , \g2661_reg/NET0131 , \g2667_reg/NET0131 , \g2671_reg/NET0131 , \g2675_reg/NET0131 , \g2681_reg/NET0131 , \g2685_reg/NET0131 , \g269_reg/NET0131 , \g2715_reg/NET0131 , \g2719_reg/NET0131 , \g2724_reg/NET0131 , \g2729_reg/NET0131 , \g2735_reg/NET0131 , \g2741_reg/NET0131 , \g2748_reg/NET0131 , \g2756_reg/NET0131 , \g2759_reg/NET0131 , \g2763_reg/NET0131 , \g2767_reg/NET0131 , \g2771_reg/NET0131 , \g2775_reg/NET0131 , \g2779_reg/NET0131 , \g2783_reg/NET0131 , \g2787_reg/NET0131 , \g278_reg/NET0131 , \g2791_reg/NET0131 , \g2795_reg/NET0131 , \g2799_reg/NET0131 , \g2803_reg/NET0131 , \g2807_reg/NET0131 , \g2811_reg/NET0131 , \g2815_reg/NET0131 , \g2819_reg/NET0131 , \g2823_reg/NET0131 , \g2827_reg/NET0131 , \g2831_reg/NET0131 , \g2834_reg/NET0131 , \g283_reg/NET0131 , \g2848_reg/NET0131 , \g2856_reg/NET0131 , \g2864_reg/NET0131 , \g2873_reg/NET0131 , \g2878_reg/NET0131 , \g287_reg/NET0131 , \g2882_reg/NET0131 , \g2886_reg/NET0131 , \g2898_reg/NET0131 , \g2902_reg/NET0131 , \g2907_reg/NET0131 , \g2912_reg/NET0131 , \g2917_reg/NET0131 , \g291_reg/NET0131 , \g29211_pad , \g29212_pad , \g29213_pad , \g29214_pad , \g29215_pad , \g29216_pad , \g29218_pad , \g29219_pad , \g29220_pad , \g29221_pad , \g2922_reg/NET0131 , \g2927_reg/NET0131 , \g2932_reg/NET0131 , \g2936_reg/NET0131 , \g2941_reg/NET0131 , \g2946_reg/NET0131 , \g294_reg/NET0131 , \g2950_reg/NET0131 , \g2955_reg/NET0131 , \g2960_reg/NET0131 , \g2965_reg/NET0131 , \g2970_reg/NET0131 , \g2975_reg/NET0131 , \g2980_reg/NET0131 , \g2984_reg/NET0131 , \g2988_reg/NET0131 , \g298_reg/NET0131 , \g2999_reg/NET0131 , \g3003_reg/NET0131 , \g301_reg/NET0131 , \g3050_reg/NET0131 , \g305_reg/NET0131 , \g3096_reg/NET0131 , \g3100_reg/NET0131 , \g3106_reg/NET0131 , \g3111_reg/NET0131 , \g3115_reg/NET0131 , \g3119_reg/NET0131 , \g311_reg/NET0131 , \g3125_reg/NET0131 , \g3129_reg/NET0131 , \g3133_reg/NET0131 , \g3139_reg/NET0131 , \g3143_reg/NET0131 , \g3147_reg/NET0131 , \g3155_reg/NET0131 , \g3161_reg/NET0131 , \g3167_reg/NET0131 , \g316_reg/NET0131 , \g3171_reg/NET0131 , \g3179_reg/NET0131 , \g3187_reg/NET0131 , \g3191_reg/NET0131 , \g3195_reg/NET0131 , \g3199_reg/NET0131 , \g319_reg/NET0131 , \g3203_reg/NET0131 , \g3207_reg/NET0131 , \g3211_reg/NET0131 , \g3215_reg/NET0131 , \g3219_reg/NET0131 , \g3223_reg/NET0131 , \g3227_reg/NET0131 , \g3231_reg/NET0131 , \g3235_reg/NET0131 , \g3239_reg/NET0131 , \g3243_reg/NET0131 , \g3247_reg/NET0131 , \g324_reg/NET0131 , \g3251_reg/NET0131 , \g3255_reg/NET0131 , \g3259_reg/NET0131 , \g3263_reg/NET0131 , \g3288_reg/NET0131 , \g329_reg/NET0131 , \g3303_reg/NET0131 , \g3329_reg/NET0131 , \g3333_reg/NET0131 , \g3338_reg/NET0131 , \g333_reg/NET0131 , \g3343_reg/NET0131 , \g3347_reg/NET0131 , \g3352_reg/NET0131 , \g336_reg/NET0131 , \g341_reg/NET0131 , \g3457_reg/NET0131 , \g3466_reg/NET0131 , \g3470_reg/NET0131 , \g3476_reg/NET0131 , \g347_reg/NET0131 , \g3480_reg/NET0131 , \g3484_reg/NET0131 , \g3490_reg/NET0131 , \g3494_reg/NET0131 , \g34_reg/NET0131 , \g351_reg/NET0131 , \g355_reg/NET0131 , \g358_reg/NET0131 , \g35_pad , \g3639_reg/NET0131 , \g3684_reg/NET0131 , \g3703_reg/NET0131 , \g370_reg/NET0131 , \g376_reg/NET0131 , \g37_reg/NET0131 , \g3808_reg/NET0131 , \g3817_reg/NET0131 , \g3821_reg/NET0131 , \g3827_reg/NET0131 , \g3831_reg/NET0131 , \g3835_reg/NET0131 , \g3841_reg/NET0131 , \g3845_reg/NET0131 , \g385_reg/NET0131 , \g392_reg/NET0131 , \g3990_reg/NET0131 , \g401_reg/NET0131 , \g4035_reg/NET0131 , \g4054_reg/NET0131 , \g4057_reg/NET0131 , \g405_reg/NET0131 , \g4064_reg/NET0131 , \g4072_reg/NET0131 , \g4076_reg/NET0131 , \g4082_reg/NET0131 , \g4087_reg/NET0131 , \g4093_reg/NET0131 , \g4098_reg/NET0131 , \g4104_reg/NET0131 , \g4108_reg/NET0131 , \g4112_reg/NET0131 , \g4116_reg/NET0131 , \g4119_reg/NET0131 , \g411_reg/NET0131 , \g4122_reg/NET0131 , \g4141_reg/NET0131 , \g4145_reg/NET0131 , \g4146_reg/NET0131 , \g4153_reg/NET0131 , \g4157_reg/NET0131 , \g4164_reg/NET0131 , \g4172_reg/NET0131 , \g4176_reg/NET0131 , \g417_reg/NET0131 , \g4180_reg/NET0131 , \g4235_reg/NET0131 , \g4239_reg/NET0131 , \g4242_reg/NET0131 , \g4245_reg/NET0131 , \g424_reg/NET0131 , \g4253_reg/NET0131 , \g4258_reg/NET0131 , \g4264_reg/NET0131 , \g4269_reg/NET0131 , \g4273_reg/NET0131 , \g4281_reg/NET0131 , \g4284_reg/NET0131 , \g4291_reg/NET0131 , \g4297_reg/NET0131 , \g4300_reg/NET0131 , \g4308_reg/NET0131 , \g4311_reg/NET0131 , \g4322_reg/NET0131 , \g4332_reg/NET0131 , \g433_reg/NET0131 , \g4340_reg/NET0131 , \g4349_reg/NET0131 , \g4358_reg/NET0131 , \g4366_reg/NET0131 , \g4369_reg/NET0131 , \g4372_reg/NET0131 , \g4375_reg/NET0131 , \g437_reg/NET0131 , \g4382_reg/NET0131 , \g4388_reg/NET0131 , \g4392_reg/NET0131 , \g4401_reg/NET0131 , \g4405_reg/NET0131 , \g4411_reg/NET0131 , \g4417_reg/NET0131 , \g441_reg/NET0131 , \g4420_reg/NET0131 , \g4423_reg/NET0131 , \g4427_reg/NET0131 , \g4430_reg/NET0131 , \g4434_reg/NET0131 , \g4438_reg/NET0131 , \g4443_reg/NET0131 , \g4452_reg/NET0131 , \g4455_reg/NET0131 , \g4459_reg/NET0131 , \g4462_reg/NET0131 , \g4467_reg/NET0131 , \g446_reg/NET0131 , \g4473_reg/NET0131 , \g4477_reg/NET0131 , \g4480_reg/NET0131 , \g4483_reg/NET0131 , \g4486_reg/NET0131 , \g4489_reg/NET0131 , \g4492_reg/NET0131 , \g4495_reg/NET0131 , \g4498_reg/NET0131 , \g4501_reg/NET0131 , \g4504_reg/NET0131 , \g4512_reg/NET0131 , \g4515_reg/NET0131 , \g4521_reg/NET0131 , \g4527_reg/NET0131 , \g452_reg/NET0131 , \g4531_reg/NET0131 , \g4534_reg/NET0131 , \g4540_reg/NET0131 , \g4543_reg/NET0131 , \g4546_reg/NET0131 , \g4549_reg/NET0131 , \g4552_reg/NET0131 , \g4555_reg/NET0131 , \g4558_reg/NET0131 , \g4561_reg/NET0131 , \g4564_reg/NET0131 , \g4567_reg/NET0131 , \g4572_reg/NET0131 , \g4575_reg/NET0131 , \g4581_reg/NET0131 , \g4584_reg/NET0131 , \g4593_reg/NET0131 , \g4601_reg/NET0131 , \g4608_reg/NET0131 , \g460_reg/NET0131 , \g4616_reg/NET0131 , \g4621_reg/NET0131 , \g4628_reg/NET0131 , \g4633_reg/NET0131 , \g4639_reg/NET0131 , \g4643_reg/NET0131 , \g4646_reg/NET0131 , \g4653_reg/NET0131 , \g4659_reg/NET0131 , \g4664_reg/NET0131 , \g4669_reg/NET0131 , \g4674_reg/NET0131 , \g4681_reg/NET0131 , \g4688_reg/NET0131 , \g4698_reg/NET0131 , \g4704_reg/NET0131 , \g4709_reg/NET0131 , \g4743_reg/NET0131 , \g4749_reg/NET0131 , \g4754_reg/NET0131 , \g475_reg/NET0131 , \g4760_reg/NET0131 , \g4765_reg/NET0131 , \g4771_reg/NET0131 , \g4776_reg/NET0131 , \g4785_reg/NET0131 , \g4793_reg/NET0131 , \g479_reg/NET0131 , \g4801_reg/NET0131 , \g482_reg/NET0131 , \g490_reg/NET0131 , \g496_reg/NET0131 , \g499_reg/NET0131 , \g5016_reg/NET0131 , \g5022_reg/NET0131 , \g5029_reg/NET0131 , \g5033_reg/NET0131 , \g5037_reg/NET0131 , \g5041_reg/NET0131 , \g5046_reg/NET0131 , \g504_reg/NET0131 , \g5052_reg/NET0131 , \g5057_reg/NET0131 , \g5069_reg/NET0131 , \g5073_reg/NET0131 , \g5077_reg/NET0131 , \g5080_reg/NET0131 , \g5084_reg/NET0131 , \g5092_reg/NET0131 , \g5097_reg/NET0131 , \g5101_reg/NET0131 , \g5112_reg/NET0131 , \g5115_reg/NET0131 , \g5124_reg/NET0131 , \g5128_reg/NET0131 , \g5134_reg/NET0131 , \g5138_reg/NET0131 , \g513_reg/NET0131 , \g5142_reg/NET0131 , \g5148_reg/NET0131 , \g5152_reg/NET0131 , \g518_reg/NET0131 , \g528_reg/NET0131 , \g5297_reg/NET0131 , \g534_reg/NET0131 , \g5357_reg/NET0131 , \g538_reg/NET0131 , \g542_reg/NET0131 , \g546_reg/NET0131 , \g550_reg/NET0131 , \g554_reg/NET0131 , \g645_reg/NET0131 , \g650_reg/NET0131 , \g655_reg/NET0131 , \g661_reg/NET0131 , \g667_reg/NET0131 , \g671_reg/NET0131 , \g676_reg/NET0131 , \g681_reg/NET0131 , \g686_reg/NET0131 , \g691_reg/NET0131 , \g699_reg/NET0131 , \g703_reg/NET0131 , \g714_reg/NET0131 , \g718_reg/NET0131 , \g723_reg/NET0131 , \g7243_pad , \g7245_pad , \g7257_pad , \g7260_pad , \g728_reg/NET0131 , \g732_reg/NET0131 , \g736_reg/NET0131 , \g739_reg/NET0131 , \g744_reg/NET0131 , \g749_reg/NET0131 , \g753_reg/NET0131 , \g7540_pad , \g758_reg/NET0131 , \g763_reg/NET0131 , \g767_reg/NET0131 , \g772_reg/NET0131 , \g776_reg/NET0131 , \g781_reg/NET0131 , \g785_reg/NET0131 , \g790_reg/NET0131 , \g7916_pad , \g7946_pad , \g794_reg/NET0131 , \g802_reg/NET0131 , \g807_reg/NET0131 , \g812_reg/NET0131 , \g817_reg/NET0131 , \g822_reg/NET0131 , \g827_reg/NET0131 , \g8291_pad , \g832_reg/NET0131 , \g8358_pad , \g837_reg/NET0131 , \g8416_pad , \g843_reg/NET0131 , \g8475_pad , \g847_reg/NET0131 , \g854_reg/NET0131 , \g862_reg/NET0131 , \g8719_pad , \g872_reg/NET0131 , \g8783_pad , \g8784_pad , \g8785_pad , \g8786_pad , \g8787_pad , \g8788_pad , \g8789_pad , \g8839_pad , \g8870_pad , \g890_reg/NET0131 , \g8915_pad , \g8916_pad , \g8917_pad , \g8918_pad , \g8919_pad , \g8920_pad , \g896_reg/NET0131 , \g9019_pad , \g9251_pad , \g956_reg/NET0131 , \g962_reg/NET0131 , \g969_reg/NET0131 , \g976_reg/NET0131 , \g979_reg/NET0131 , \g990_reg/NET0131 , \g996_reg/NET0131 , \g136_reg/P0001 , \g21727_pad , \g23190_pad , \g26875_pad , \g26876_pad , \g26877_pad , \g28041_pad , \g28042_pad , \g30327_pad , \g30330_pad , \g30331_pad , \g31793_pad , \g31860_pad , \g31862_pad , \g31863_pad , \g32185_pad , \g33079_pad , \g33435_pad , \g33959_pad , \g34435_pad , \g34788_pad , \g34956_pad , \g34_reg/P0001 , \g35_syn_2 , \g37/_0_ , \g41/_0_ , \g60853/_3_ , \g60856/_3_ , \g60879/_3_ , \g60882/_0_ , \g60888/_0_ , \g60891/_0_ , \g60896/_0_ , \g60899/_0_ , \g60900/_3_ , \g60909/_3_ , \g60911/_0_ , \g60915/_0_ , \g60918/_0_ , \g60919/_0_ , \g60928/_0_ , \g60929/_0_ , \g60936/_0_ , \g60937/_0_ , \g60939/_0_ , \g60940/_0_ , \g60941/_0_ , \g60942/_0_ , \g60943/_0_ , \g60944/_0_ , \g60952/_0_ , \g60954/_0_ , \g60958/_0_ , \g60962/_3_ , \g60972/_0_ , \g60980/_0_ , \g60984/_0_ , \g60986/_0_ , \g60989/_0_ , \g60991/_3_ , \g61006/_0_ , \g61008/_0_ , \g61013/_0_ , \g61014/_0_ , \g61015/_0_ , \g61016/_0_ , \g61017/_0_ , \g61026/_3_ , \g61027/_3_ , \g61030/_0_ , \g61031/_0_ , \g61037/_0_ , \g61038/_0_ , \g61042/_0_ , \g61044/_0_ , \g61045/_0_ , \g61046/_0_ , \g61050/_0_ , \g61051/_0_ , \g61052/_0_ , \g61078/_0_ , \g61131/_0_ , \g61137/_3_ , \g61142/_3_ , \g61143/_3_ , \g61151/_0_ , \g61152/_0_ , \g61161/_0_ , \g61168/_3_ , \g61169/_3_ , \g61170/_0_ , \g61171/_3_ , \g61172/_0_ , \g61173/_0_ , \g61174/_0_ , \g61175/_0_ , \g61176/_0_ , \g61177/_3_ , \g61178/_0_ , \g61179/_0_ , \g61180/_0_ , \g61181/_0_ , \g61182/_3_ , \g61183/_0_ , \g61184/_3_ , \g61185/_0_ , \g61186/_0_ , \g61187/_0_ , \g61188/_0_ , \g61189/_0_ , \g61190/_3_ , \g61191/_0_ , \g61192/_0_ , \g61193/_0_ , \g61194/_0_ , \g61221/_0_ , \g61222/_0_ , \g61223/_3_ , \g61224/_3_ , \g61261/_0_ , \g61295/_3_ , \g61308/_0_ , \g61316/_0_ , \g61327/_0_ , \g61329/_0_ , \g61330/_0_ , \g61331/_0_ , \g61332/_3_ , \g61333/_0_ , \g61334/_0_ , \g61335/_0_ , \g61336/_0_ , \g61337/_0_ , \g61338/_3_ , \g61339/_0_ , \g61340/_0_ , \g61341/_0_ , \g61342/_0_ , \g61343/_0_ , \g61344/_3_ , \g61345/_0_ , \g61346/_0_ , \g61347/_0_ , \g61348/_0_ , \g61349/_0_ , \g61350/_3_ , \g61351/_0_ , \g61352/_0_ , \g61353/_0_ , \g61354/_0_ , \g61367/_0_ , \g61372/_0_ , \g61373/_0_ , \g61375/_0_ , \g61382/_0_ , \g61385/_3_ , \g61386/_0_ , \g61399/_0_ , \g61400/_0_ , \g61402/_0_ , \g61405/_0_ , \g61435/_3_ , \g61449/_0_ , \g61468/_0_ , \g61475/_0_ , \g61480/_0_ , \g61482/_0_ , \g61483/_0_ , \g61484/_0_ , \g61486/_3_ , \g61494/_0_ , \g61496/_0_ , \g61497/_0_ , \g61514/_0_ , \g61517/_0_ , \g61519/_3_ , \g61520/_3_ , \g61527/_0_ , \g61541/_0_ , \g61544/_0_ , \g61550/_0_ , \g61551/_0_ , \g61554/_0_ , \g61556/_3_ , \g61567/_0_ , \g61571/_0_ , \g61574/_0_ , \g61587/_0_ , \g61592/_0_ , \g61632/_0_ , \g61634/_0_ , \g61635/_0_ , \g61639/_0_ , \g61644/_0_ , \g61652/_3_ , \g61709/_0_ , \g61714/_0_ , \g61720/_0_ , \g61721/_0_ , \g61723/_0_ , \g61725/_0_ , \g61726/_0_ , \g61734/_0_ , \g61739/_0_ , \g61744/_0_ , \g61746/_3_ , \g61747/_3_ , \g61748/_3_ , \g61750/u3_syn_7 , \g61802/_0_ , \g61804/_0_ , \g61808/_0_ , \g61811/_0_ , \g61816/_0_ , \g61818/_0_ , \g61820/_0_ , \g61823/_0_ , \g61824/_0_ , \g61841/_0_ , \g61842/_3_ , \g61844/_3_ , \g61845/_3_ , \g61846/_3_ , \g61847/u3_syn_7 , \g61848/_0_ , \g61849/_3_ , \g61850/_0_ , \g61851/u3_syn_7 , \g61852/_0_ , \g61853/_3_ , \g61854/_3_ , \g61855/_0_ , \g61856/u3_syn_7 , \g61857/_0_ , \g61858/_3_ , \g61859/_3_ , \g61860/u3_syn_7 , \g61861/_0_ , \g61862/_3_ , \g61863/_3_ , \g61864/u3_syn_7 , \g61865/_0_ , \g61866/_3_ , \g61867/_3_ , \g61868/u3_syn_7 , \g61869/_0_ , \g61870/_0_ , \g61871/_3_ , \g61872/_3_ , \g61873/u3_syn_7 , \g61874/_0_ , \g61875/_0_ , \g61877/_3_ , \g61878/_3_ , \g61879/u3_syn_7 , \g61880/_0_ , \g61881/_0_ , \g61882/_0_ , \g61883/_0_ , \g61884/_0_ , \g61914/_0_ , \g61915/_0_ , \g61917/_0_ , \g61918/_0_ , \g61922/_0_ , \g61923/_0_ , \g61924/_0_ , \g61932/_0_ , \g61936/_0_ , \g61945/_0_ , \g61947/_0_ , \g61959/_0_ , \g61960/_0_ , \g61962/_0_ , \g61973/_3_ , \g61974/u3_syn_7 , \g61975/_3_ , \g61976/u3_syn_7 , \g61977/_3_ , \g61978/_3_ , \g61979/u3_syn_7 , \g61980/_3_ , \g61981/_3_ , \g61982/_3_ , \g61983/u3_syn_7 , \g61984/_3_ , \g61985/_3_ , \g61986/u3_syn_7 , \g61987/_3_ , \g61988/_3_ , \g61989/u3_syn_7 , \g61990/_3_ , \g61991/_3_ , \g61992/u3_syn_7 , \g61993/_3_ , \g61994/u3_syn_7 , \g61995/_3_ , \g61996/_3_ , \g61997/_3_ , \g62022/_0_ , \g62028/_0_ , \g62029/_0_ , \g62031/_0_ , \g62033/_0_ , \g62038/_0_ , \g62042/_0_ , \g62046/_0_ , \g62048/_0_ , \g62049/_0_ , \g62051/_0_ , \g62053/_0_ , \g62085/_0_ , \g62101/_0_ , \g62102/_0_ , \g62103/_0_ , \g62105/_0_ , \g62108/_3_ , \g62112/_0_ , \g62137/_3_ , \g62207/_0_ , \g62239/_0_ , \g62240/_0_ , \g62267/_0_ , \g62273/_0_ , \g62284/_0_ , \g62291/_0_ , \g62293/_0_ , \g62298/_0_ , \g62303/_3_ , \g62322/_3_ , \g62323/_3_ , \g62324/_3_ , \g62325/_3_ , \g62583/_0_ , \g62598/_0_ , \g62609/_0_ , \g62636/_0_ , \g62646/_0_ , \g62649/_0_ , \g62658/_0_ , \g62663/_0_ , \g62664/_0_ , \g62667/_0_ , \g62676/_0_ , \g62677/_0_ , \g62678/_3_ , \g62679/_0_ , \g62687/u3_syn_7 , \g62688/u3_syn_7 , \g62689/_0_ , \g62690/_3_ , \g62691/_3_ , \g62693/_0_ , \g62694/_3_ , \g62695/_3_ , \g62696/_3_ , \g62697/_3_ , \g62698/_3_ , \g62699/_3_ , \g62700/_3_ , \g62701/_3_ , \g62702/_3_ , \g62703/_3_ , \g62704/u3_syn_7 , \g62705/_0_ , \g62706/_3_ , \g62707/_3_ , \g62708/u3_syn_7 , \g62709/_0_ , \g62710/_3_ , \g62711/_3_ , \g62712/u3_syn_7 , \g62713/_0_ , \g62714/_3_ , \g62715/_0_ , \g62716/u3_syn_7 , \g62717/_0_ , \g62718/_3_ , \g62719/_0_ , \g62720/u3_syn_7 , \g62721/_0_ , \g62722/_3_ , \g62723/_0_ , \g62724/u3_syn_7 , \g62725/_0_ , \g62726/_3_ , \g62728/_0_ , \g62790/_0_ , \g62791/_0_ , \g62793/_0_ , \g62794/_0_ , \g62795/_0_ , \g62796/_0_ , \g62797/_0_ , \g62807/_0_ , \g62823/_0_ , \g62824/_0_ , \g62833/_0_ , \g62846/_0_ , \g62859/_0_ , \g62860/_0_ , \g62897/_0_ , \g62898/_0_ , \g62922/_3_ , \g62923/_0_ , \g62927/_0_ , \g62938/_3_ , \g62939/_3_ , \g62940/_3_ , \g62941/u3_syn_7 , \g62942/_0_ , \g62943/_3_ , \g62987/_3_ , \g62991/_3_ , \g63015/u3_syn_7 , \g63016/_0_ , \g63017/_3_ , \g63018/_3_ , \g63019/_3_ , \g63020/_3_ , \g63021/_3_ , \g63022/_3_ , \g63025/_3_ , \g63026/_3_ , \g63027/_3_ , \g63029/_3_ , \g63030/_3_ , \g63031/_3_ , \g63033/_3_ , \g63034/_3_ , \g63043/_3_ , \g63044/_3_ , \g63051/_3_ , \g63057/_3_ , \g63068/_3_ , \g63070/_3_ , \g63073/_3_ , \g63081/_3_ , \g63082/_3_ , \g63083/u3_syn_7 , \g63084/_3_ , \g63085/_0_ , \g63086/_3_ , \g63107/_3_ , \g63108/u3_syn_7 , \g63109/u3_syn_7 , \g63110/_0_ , \g63111/_3_ , \g63132/_3_ , \g63133/_3_ , \g63134/_3_ , \g63135/_3_ , \g63136/_3_ , \g63137/_3_ , \g63138/_3_ , \g63139/u3_syn_7 , \g63140/_3_ , \g63141/_3_ , \g63142/_3_ , \g63143/_3_ , \g63144/_3_ , \g63145/_3_ , \g63146/u3_syn_7 , \g63198/_0_ , \g63205/_0_ , \g63208/_0_ , \g63212/_0_ , \g63215/_0_ , \g63219/_0_ , \g63244/_0_ , \g63246/_0_ , \g63254/_0_ , \g63255/_0_ , \g63272/_0_ , \g63276/_0_ , \g63278/_0_ , \g63279/_0_ , \g63280/_0_ , \g63327/_0_ , \g63345/_0_ , \g63346/_3_ , \g63347/_3_ , \g63354/_3_ , \g63358/_3_ , \g63359/u3_syn_7 , \g63361/_3_ , \g63365/_3_ , \g63366/_3_ , \g63367/_3_ , \g63368/_3_ , \g63370/_3_ , \g63479/_0_ , \g63484/_0_ , \g63499/_1_ , \g63520/_0_ , \g63523/_0_ , \g63526/_0_ , \g63538/_0_ , \g63539/_0_ , \g63541/_0_ , \g63555/_0_ , \g63642/_0_ , \g63645/_0_ , \g63648/_3_ , \g63777/_3_ , \g63778/_3_ , \g63781/_0_ , \g63786/u3_syn_7 , \g63787/_3_ , \g63788/_3_ , \g63790/_3_ , \g63791/_3_ , \g63792/u3_syn_7 , \g63794/_0_ , \g63795/_0_ , \g63796/_0_ , \g63798/_3_ , \g63800/_3_ , \g63804/_3_ , \g63805/_3_ , \g63806/_3_ , \g63807/_3_ , \g63808/_3_ , \g63809/_3_ , \g63870/_0_ , \g63883/_0_ , \g63934/_0_ , \g63936/_0_ , \g63938/_0_ , \g63939/_0_ , \g63966/_0_ , \g63970/_0_ , \g63999/_0_ , \g64039/_0_ , \g64040/_0_ , \g64043/_0_ , \g64062/_3_ , \g64078/_0_ , \g64091/_0_ , \g64095/_3_ , \g64096/_3_ , \g64097/u3_syn_7 , \g64098/u3_syn_7 , \g64099/u3_syn_7 , \g64100/u3_syn_7 , \g64134/_0_ , \g64135/_0_ , \g64153/_0_ , \g64155/_0_ , \g64179/_0_ , \g64229/_0_ , \g64235/_0_ , \g64236/_0_ , \g64280/_0_ , \g64315/_0_ , \g64365/_0_ , \g64426/_3_ , \g64438/_3_ , \g64442/u3_syn_7 , \g64445/_3_ , \g64447/_3_ , \g64449/_3_ , \g64451/_3_ , \g64453/_3_ , \g64454/_3_ , \g64460/_3_ , \g64461/_3_ , \g64510/_0_ , \g64527/_0_ , \g64528/_0_ , \g64544/_0_ , \g64549/_0_ , \g64566/_0_ , \g64576/_0_ , \g64602/_0_ , \g64691/_0_ , \g64697/_0_ , \g64707/_3_ , \g64778/_3_ , \g64790/_3_ , \g64791/_3_ , \g64792/_3_ , \g64793/_3_ , \g64794/_3_ , \g64795/_3_ , \g64796/_3_ , \g64797/_3_ , \g64877/_0_ , \g64912/_0_ , \g64973/_0_ , \g65047/_3_ , \g65081/_3_ , \g65088/_3_ , \g65097/_3_ , \g65100/_3_ , \g65101/_3_ , \g65104/_3_ , \g65105/_3_ , \g65107/_3_ , \g65110/_3_ , \g65111/_3_ , \g65113/_3_ , \g65114/_3_ , \g65266/_0_ , \g65267/_0_ , \g65294/_1_ , \g65328/_1_ , \g65495/_0_ , \g65499/_0_ , \g65503/_0_ , \g65529/_0_ , \g65530/_3_ , \g65531/_3_ , \g65532/_3_ , \g65533/_3_ , \g65624/_0_ , \g65625/_1_ , \g65641/_0_ , \g65701/_0_ , \g65704/_0_ , \g65853/_0_ , \g65891/_0_ , \g65901/_0_ , \g65986/_0_ , \g66029/_0_ , \g66066/_0_ , \g66067/_0_ , \g66068/_0_ , \g66154/_3_ , \g66362/_0_ , \g66369/_0_ , \g66398/_0_ , \g66409/_0_ , \g66419/_0_ , \g66439/_0_ , \g66443/_0_ , \g66464/_0_ , \g66471/_0_ , \g66512/_0_ , \g66528/_0_ , \g66541/_0_ , \g66558/_0_ , \g66644/_0_ , \g66684/_0_ , \g66697/_0_ , \g66698/_0_ , \g66701/_0_ , \g66714/_0_ , \g66715/_0_ , \g66745/_0_ , \g66750/_0_ , \g66751/_0_ , \g66810/_0_ , \g66844/_0_ , \g66853/_0_ , \g66897/_0_ , \g66905/_0_ , \g69743/_0_ , \g69750/_0_ , \g69773/_1_ , \g69792/_1_ , \g69858/_0_ , \g69938/_0_ , \g69949/_0_ , \g70167/_0_ , \g71190/_0_ , \g71198/_0_ , \g71284/_0_ , \g72369/_1_ , \g72467/_0_ , \g72476/_0_ , \g72477/_1_ , \g72648/_0_ , \g72741/_0_ , \g72772/_0_ , \g8132_pad );
	input \g1002_reg/NET0131  ;
	input \g1008_reg/NET0131  ;
	input \g10122_pad  ;
	input \g1018_reg/NET0131  ;
	input \g1024_reg/NET0131  ;
	input \g10306_pad  ;
	input \g1030_reg/NET0131  ;
	input \g1036_reg/NET0131  ;
	input \g1041_reg/NET0131  ;
	input \g1046_reg/NET0131  ;
	input \g10500_pad  ;
	input \g10527_pad  ;
	input \g1052_reg/NET0131  ;
	input \g1061_reg/NET0131  ;
	input \g1070_reg/NET0131  ;
	input \g1087_reg/NET0131  ;
	input \g1094_reg/NET0131  ;
	input \g1099_reg/NET0131  ;
	input \g1105_reg/NET0131  ;
	input \g1111_reg/NET0131  ;
	input \g1124_reg/NET0131  ;
	input \g1129_reg/NET0131  ;
	input \g1135_reg/NET0131  ;
	input \g1141_reg/NET0131  ;
	input \g11447_pad  ;
	input \g1146_reg/NET0131  ;
	input \g1152_reg/NET0131  ;
	input \g1171_reg/NET0131  ;
	input \g11770_pad  ;
	input \g1178_reg/NET0131  ;
	input \g1183_reg/NET0131  ;
	input \g1189_reg/NET0131  ;
	input \g1193_reg/NET0131  ;
	input \g1199_reg/NET0131  ;
	input \g1205_reg/NET0131  ;
	input \g1211_reg/NET0131  ;
	input \g1216_reg/NET0131  ;
	input \g12184_pad  ;
	input \g1221_reg/NET0131  ;
	input \g1236_reg/NET0131  ;
	input \g1242_reg/NET0131  ;
	input \g1246_reg/NET0131  ;
	input \g12919_pad  ;
	input \g12923_pad  ;
	input \g1300_reg/NET0131  ;
	input \g13039_pad  ;
	input \g1306_reg/NET0131  ;
	input \g1312_reg/NET0131  ;
	input \g1319_reg/NET0131  ;
	input \g1322_reg/NET0131  ;
	input \g13259_pad  ;
	input \g13272_pad  ;
	input \g1333_reg/NET0131  ;
	input \g1339_reg/NET0131  ;
	input \g1345_reg/NET0131  ;
	input \g1351_reg/NET0131  ;
	input \g1361_reg/NET0131  ;
	input \g1367_reg/NET0131  ;
	input \g1373_reg/NET0131  ;
	input \g1379_reg/NET0131  ;
	input \g1384_reg/NET0131  ;
	input \g13865_pad  ;
	input \g13895_pad  ;
	input \g1389_reg/NET0131  ;
	input \g1395_reg/NET0131  ;
	input \g1404_reg/NET0131  ;
	input \g14096_pad  ;
	input \g14125_pad  ;
	input \g1413_reg/NET0131  ;
	input \g14147_pad  ;
	input \g14167_pad  ;
	input \g14189_pad  ;
	input \g14201_pad  ;
	input \g14217_pad  ;
	input \g142_reg/NET0131  ;
	input \g1430_reg/NET0131  ;
	input \g1437_reg/NET0131  ;
	input \g1442_reg/NET0131  ;
	input \g1448_reg/NET0131  ;
	input \g1454_reg/NET0131  ;
	input \g1467_reg/NET0131  ;
	input \g146_reg/NET0131  ;
	input \g1472_reg/NET0131  ;
	input \g1478_reg/NET0131  ;
	input \g1484_reg/NET0131  ;
	input \g1489_reg/NET0131  ;
	input \g1495_reg/NET0131  ;
	input \g150_reg/NET0131  ;
	input \g1514_reg/NET0131  ;
	input \g1521_reg/NET0131  ;
	input \g1526_reg/NET0131  ;
	input \g1532_reg/NET0131  ;
	input \g1536_reg/NET0131  ;
	input \g153_reg/NET0131  ;
	input \g1542_reg/NET0131  ;
	input \g1548_reg/NET0131  ;
	input \g1554_reg/NET0131  ;
	input \g1559_reg/NET0131  ;
	input \g1564_reg/NET0131  ;
	input \g1579_reg/NET0131  ;
	input \g157_reg/NET0131  ;
	input \g1585_reg/NET0131  ;
	input \g1589_reg/NET0131  ;
	input \g1592_reg/NET0131  ;
	input \g1600_reg/NET0131  ;
	input \g1604_reg/NET0131  ;
	input \g1608_reg/NET0131  ;
	input \g160_reg/NET0131  ;
	input \g1612_reg/NET0131  ;
	input \g1616_reg/NET0131  ;
	input \g1620_reg/NET0131  ;
	input \g1624_reg/NET0131  ;
	input \g1632_reg/NET0131  ;
	input \g1636_reg/NET0131  ;
	input \g1644_reg/NET0131  ;
	input \g1648_reg/NET0131  ;
	input \g164_reg/NET0131  ;
	input \g1657_reg/NET0131  ;
	input \g16603_pad  ;
	input \g16624_pad  ;
	input \g1664_reg/NET0131  ;
	input \g16686_pad  ;
	input \g1668_reg/NET0131  ;
	input \g16718_pad  ;
	input \g1677_reg/NET0131  ;
	input \g1682_reg/NET0131  ;
	input \g16874_pad  ;
	input \g1687_reg/NET0131  ;
	input \g168_reg/NET0131  ;
	input \g1691_reg/NET0131  ;
	input \g1696_reg/NET0131  ;
	input \g1700_reg/NET0131  ;
	input \g1706_reg/NET0131  ;
	input \g1710_reg/NET0131  ;
	input \g1714_reg/NET0131  ;
	input \g1720_reg/NET0131  ;
	input \g1724_reg/NET0131  ;
	input \g1728_reg/NET0131  ;
	input \g17291_pad  ;
	input \g17316_pad  ;
	input \g17320_pad  ;
	input \g1736_reg/NET0131  ;
	input \g17400_pad  ;
	input \g17404_pad  ;
	input \g1740_reg/NET0131  ;
	input \g17423_pad  ;
	input \g1744_reg/NET0131  ;
	input \g1748_reg/NET0131  ;
	input \g174_reg/NET0131  ;
	input \g1752_reg/NET0131  ;
	input \g1756_reg/NET0131  ;
	input \g1760_reg/NET0131  ;
	input \g1768_reg/NET0131  ;
	input \g1772_reg/NET0131  ;
	input \g1779_reg/NET0131  ;
	input \g1783_reg/NET0131  ;
	input \g1792_reg/NET0131  ;
	input \g1798_reg/NET0131  ;
	input \g1802_reg/NET0131  ;
	input \g18094_pad  ;
	input \g18095_pad  ;
	input \g18096_pad  ;
	input \g18098_pad  ;
	input \g18099_pad  ;
	input \g1811_reg/NET0131  ;
	input \g1816_reg/NET0131  ;
	input \g1821_reg/NET0131  ;
	input \g1825_reg/NET0131  ;
	input \g182_reg/NET0131  ;
	input \g1830_reg/NET0131  ;
	input \g1834_reg/NET0131  ;
	input \g1840_reg/NET0131  ;
	input \g1844_reg/NET0131  ;
	input \g1848_reg/NET0131  ;
	input \g1854_reg/NET0131  ;
	input \g1858_reg/NET0131  ;
	input \g1862_reg/NET0131  ;
	input \g1870_reg/NET0131  ;
	input \g1874_reg/NET0131  ;
	input \g1878_reg/NET0131  ;
	input \g1882_reg/NET0131  ;
	input \g1886_reg/NET0131  ;
	input \g1890_reg/NET0131  ;
	input \g1894_reg/NET0131  ;
	input \g1902_reg/NET0131  ;
	input \g1906_reg/NET0131  ;
	input \g1913_reg/NET0131  ;
	input \g1917_reg/NET0131  ;
	input \g191_reg/NET0131  ;
	input \g1926_reg/NET0131  ;
	input \g1932_reg/NET0131  ;
	input \g19334_pad  ;
	input \g19357_pad  ;
	input \g1936_reg/NET0131  ;
	input \g1945_reg/NET0131  ;
	input \g1950_reg/NET0131  ;
	input \g1955_reg/NET0131  ;
	input \g1959_reg/NET0131  ;
	input \g1964_reg/NET0131  ;
	input \g1968_reg/NET0131  ;
	input \g1974_reg/NET0131  ;
	input \g1978_reg/NET0131  ;
	input \g1982_reg/NET0131  ;
	input \g1988_reg/NET0131  ;
	input \g1992_reg/NET0131  ;
	input \g1996_reg/NET0131  ;
	input \g2004_reg/NET0131  ;
	input \g2008_reg/NET0131  ;
	input \g2012_reg/NET0131  ;
	input \g2016_reg/NET0131  ;
	input \g2020_reg/NET0131  ;
	input \g2024_reg/NET0131  ;
	input \g2028_reg/NET0131  ;
	input \g2036_reg/NET0131  ;
	input \g203_reg/NET0131  ;
	input \g2040_reg/NET0131  ;
	input \g2047_reg/NET0131  ;
	input \g2051_reg/NET0131  ;
	input \g2060_reg/NET0131  ;
	input \g2066_reg/NET0131  ;
	input \g2070_reg/NET0131  ;
	input \g2079_reg/NET0131  ;
	input \g2084_reg/NET0131  ;
	input \g2089_reg/NET0131  ;
	input \g2093_reg/NET0131  ;
	input \g2098_reg/NET0131  ;
	input \g209_reg/NET0131  ;
	input \g2102_reg/NET0131  ;
	input \g2108_reg/NET0131  ;
	input \g2112_reg/NET0131  ;
	input \g2116_reg/NET0131  ;
	input \g2122_reg/NET0131  ;
	input \g2126_reg/NET0131  ;
	input \g2153_reg/NET0131  ;
	input \g2161_reg/NET0131  ;
	input \g2165_reg/NET0131  ;
	input \g2169_reg/NET0131  ;
	input \g2173_reg/NET0131  ;
	input \g2177_reg/NET0131  ;
	input \g2181_reg/NET0131  ;
	input \g2185_reg/NET0131  ;
	input \g218_reg/NET0131  ;
	input \g2193_reg/NET0131  ;
	input \g2197_reg/NET0131  ;
	input \g2204_reg/NET0131  ;
	input \g2208_reg/NET0131  ;
	input \g2217_reg/NET0131  ;
	input \g2223_reg/NET0131  ;
	input \g2227_reg/NET0131  ;
	input \g222_reg/NET0131  ;
	input \g2236_reg/NET0131  ;
	input \g2241_reg/NET0131  ;
	input \g2246_reg/NET0131  ;
	input \g2250_reg/NET0131  ;
	input \g2255_reg/NET0131  ;
	input \g2259_reg/NET0131  ;
	input \g225_reg/NET0131  ;
	input \g2265_reg/NET0131  ;
	input \g2269_reg/NET0131  ;
	input \g2273_reg/NET0131  ;
	input \g2279_reg/NET0131  ;
	input \g2283_reg/NET0131  ;
	input \g2287_reg/NET0131  ;
	input \g2295_reg/NET0131  ;
	input \g2299_reg/NET0131  ;
	input \g2303_reg/NET0131  ;
	input \g2307_reg/NET0131  ;
	input \g2311_reg/NET0131  ;
	input \g2315_reg/NET0131  ;
	input \g2319_reg/NET0131  ;
	input \g2327_reg/NET0131  ;
	input \g232_reg/NET0131  ;
	input \g2331_reg/NET0131  ;
	input \g2338_reg/NET0131  ;
	input \g2342_reg/NET0131  ;
	input \g2351_reg/NET0131  ;
	input \g2357_reg/NET0131  ;
	input \g2361_reg/NET0131  ;
	input \g2370_reg/NET0131  ;
	input \g2375_reg/NET0131  ;
	input \g2380_reg/NET0131  ;
	input \g2384_reg/NET0131  ;
	input \g2389_reg/NET0131  ;
	input \g2393_reg/NET0131  ;
	input \g2399_reg/NET0131  ;
	input \g239_reg/NET0131  ;
	input \g2403_reg/NET0131  ;
	input \g2407_reg/NET0131  ;
	input \g2413_reg/NET0131  ;
	input \g2417_reg/NET0131  ;
	input \g2421_reg/NET0131  ;
	input \g2429_reg/NET0131  ;
	input \g2433_reg/NET0131  ;
	input \g2437_reg/NET0131  ;
	input \g2441_reg/NET0131  ;
	input \g2445_reg/NET0131  ;
	input \g2449_reg/NET0131  ;
	input \g2453_reg/NET0131  ;
	input \g2461_reg/NET0131  ;
	input \g2465_reg/NET0131  ;
	input \g246_reg/NET0131  ;
	input \g2472_reg/NET0131  ;
	input \g2476_reg/NET0131  ;
	input \g2485_reg/NET0131  ;
	input \g2491_reg/NET0131  ;
	input \g2495_reg/NET0131  ;
	input \g2504_reg/NET0131  ;
	input \g2509_reg/NET0131  ;
	input \g2514_reg/NET0131  ;
	input \g2518_reg/NET0131  ;
	input \g2523_reg/NET0131  ;
	input \g2527_reg/NET0131  ;
	input \g2533_reg/NET0131  ;
	input \g2537_reg/NET0131  ;
	input \g2541_reg/NET0131  ;
	input \g2547_reg/NET0131  ;
	input \g2551_reg/NET0131  ;
	input \g2555_reg/NET0131  ;
	input \g255_reg/NET0131  ;
	input \g2563_reg/NET0131  ;
	input \g2567_reg/NET0131  ;
	input \g2571_reg/NET0131  ;
	input \g2575_reg/NET0131  ;
	input \g2579_reg/NET0131  ;
	input \g2583_reg/NET0131  ;
	input \g2587_reg/NET0131  ;
	input \g2595_reg/NET0131  ;
	input \g2599_reg/NET0131  ;
	input \g2606_reg/NET0131  ;
	input \g2610_reg/NET0131  ;
	input \g2619_reg/NET0131  ;
	input \g2625_reg/NET0131  ;
	input \g2629_reg/NET0131  ;
	input \g262_reg/NET0131  ;
	input \g2638_reg/NET0131  ;
	input \g2643_reg/NET0131  ;
	input \g2648_reg/NET0131  ;
	input \g2652_reg/NET0131  ;
	input \g2657_reg/NET0131  ;
	input \g2661_reg/NET0131  ;
	input \g2667_reg/NET0131  ;
	input \g2671_reg/NET0131  ;
	input \g2675_reg/NET0131  ;
	input \g2681_reg/NET0131  ;
	input \g2685_reg/NET0131  ;
	input \g269_reg/NET0131  ;
	input \g2715_reg/NET0131  ;
	input \g2719_reg/NET0131  ;
	input \g2724_reg/NET0131  ;
	input \g2729_reg/NET0131  ;
	input \g2735_reg/NET0131  ;
	input \g2741_reg/NET0131  ;
	input \g2748_reg/NET0131  ;
	input \g2756_reg/NET0131  ;
	input \g2759_reg/NET0131  ;
	input \g2763_reg/NET0131  ;
	input \g2767_reg/NET0131  ;
	input \g2771_reg/NET0131  ;
	input \g2775_reg/NET0131  ;
	input \g2779_reg/NET0131  ;
	input \g2783_reg/NET0131  ;
	input \g2787_reg/NET0131  ;
	input \g278_reg/NET0131  ;
	input \g2791_reg/NET0131  ;
	input \g2795_reg/NET0131  ;
	input \g2799_reg/NET0131  ;
	input \g2803_reg/NET0131  ;
	input \g2807_reg/NET0131  ;
	input \g2811_reg/NET0131  ;
	input \g2815_reg/NET0131  ;
	input \g2819_reg/NET0131  ;
	input \g2823_reg/NET0131  ;
	input \g2827_reg/NET0131  ;
	input \g2831_reg/NET0131  ;
	input \g2834_reg/NET0131  ;
	input \g283_reg/NET0131  ;
	input \g2848_reg/NET0131  ;
	input \g2856_reg/NET0131  ;
	input \g2864_reg/NET0131  ;
	input \g2873_reg/NET0131  ;
	input \g2878_reg/NET0131  ;
	input \g287_reg/NET0131  ;
	input \g2882_reg/NET0131  ;
	input \g2886_reg/NET0131  ;
	input \g2898_reg/NET0131  ;
	input \g2902_reg/NET0131  ;
	input \g2907_reg/NET0131  ;
	input \g2912_reg/NET0131  ;
	input \g2917_reg/NET0131  ;
	input \g291_reg/NET0131  ;
	input \g29211_pad  ;
	input \g29212_pad  ;
	input \g29213_pad  ;
	input \g29214_pad  ;
	input \g29215_pad  ;
	input \g29216_pad  ;
	input \g29218_pad  ;
	input \g29219_pad  ;
	input \g29220_pad  ;
	input \g29221_pad  ;
	input \g2922_reg/NET0131  ;
	input \g2927_reg/NET0131  ;
	input \g2932_reg/NET0131  ;
	input \g2936_reg/NET0131  ;
	input \g2941_reg/NET0131  ;
	input \g2946_reg/NET0131  ;
	input \g294_reg/NET0131  ;
	input \g2950_reg/NET0131  ;
	input \g2955_reg/NET0131  ;
	input \g2960_reg/NET0131  ;
	input \g2965_reg/NET0131  ;
	input \g2970_reg/NET0131  ;
	input \g2975_reg/NET0131  ;
	input \g2980_reg/NET0131  ;
	input \g2984_reg/NET0131  ;
	input \g2988_reg/NET0131  ;
	input \g298_reg/NET0131  ;
	input \g2999_reg/NET0131  ;
	input \g3003_reg/NET0131  ;
	input \g301_reg/NET0131  ;
	input \g3050_reg/NET0131  ;
	input \g305_reg/NET0131  ;
	input \g3096_reg/NET0131  ;
	input \g3100_reg/NET0131  ;
	input \g3106_reg/NET0131  ;
	input \g3111_reg/NET0131  ;
	input \g3115_reg/NET0131  ;
	input \g3119_reg/NET0131  ;
	input \g311_reg/NET0131  ;
	input \g3125_reg/NET0131  ;
	input \g3129_reg/NET0131  ;
	input \g3133_reg/NET0131  ;
	input \g3139_reg/NET0131  ;
	input \g3143_reg/NET0131  ;
	input \g3147_reg/NET0131  ;
	input \g3155_reg/NET0131  ;
	input \g3161_reg/NET0131  ;
	input \g3167_reg/NET0131  ;
	input \g316_reg/NET0131  ;
	input \g3171_reg/NET0131  ;
	input \g3179_reg/NET0131  ;
	input \g3187_reg/NET0131  ;
	input \g3191_reg/NET0131  ;
	input \g3195_reg/NET0131  ;
	input \g3199_reg/NET0131  ;
	input \g319_reg/NET0131  ;
	input \g3203_reg/NET0131  ;
	input \g3207_reg/NET0131  ;
	input \g3211_reg/NET0131  ;
	input \g3215_reg/NET0131  ;
	input \g3219_reg/NET0131  ;
	input \g3223_reg/NET0131  ;
	input \g3227_reg/NET0131  ;
	input \g3231_reg/NET0131  ;
	input \g3235_reg/NET0131  ;
	input \g3239_reg/NET0131  ;
	input \g3243_reg/NET0131  ;
	input \g3247_reg/NET0131  ;
	input \g324_reg/NET0131  ;
	input \g3251_reg/NET0131  ;
	input \g3255_reg/NET0131  ;
	input \g3259_reg/NET0131  ;
	input \g3263_reg/NET0131  ;
	input \g3288_reg/NET0131  ;
	input \g329_reg/NET0131  ;
	input \g3303_reg/NET0131  ;
	input \g3329_reg/NET0131  ;
	input \g3333_reg/NET0131  ;
	input \g3338_reg/NET0131  ;
	input \g333_reg/NET0131  ;
	input \g3343_reg/NET0131  ;
	input \g3347_reg/NET0131  ;
	input \g3352_reg/NET0131  ;
	input \g336_reg/NET0131  ;
	input \g341_reg/NET0131  ;
	input \g3457_reg/NET0131  ;
	input \g3466_reg/NET0131  ;
	input \g3470_reg/NET0131  ;
	input \g3476_reg/NET0131  ;
	input \g347_reg/NET0131  ;
	input \g3480_reg/NET0131  ;
	input \g3484_reg/NET0131  ;
	input \g3490_reg/NET0131  ;
	input \g3494_reg/NET0131  ;
	input \g34_reg/NET0131  ;
	input \g351_reg/NET0131  ;
	input \g355_reg/NET0131  ;
	input \g358_reg/NET0131  ;
	input \g35_pad  ;
	input \g3639_reg/NET0131  ;
	input \g3684_reg/NET0131  ;
	input \g3703_reg/NET0131  ;
	input \g370_reg/NET0131  ;
	input \g376_reg/NET0131  ;
	input \g37_reg/NET0131  ;
	input \g3808_reg/NET0131  ;
	input \g3817_reg/NET0131  ;
	input \g3821_reg/NET0131  ;
	input \g3827_reg/NET0131  ;
	input \g3831_reg/NET0131  ;
	input \g3835_reg/NET0131  ;
	input \g3841_reg/NET0131  ;
	input \g3845_reg/NET0131  ;
	input \g385_reg/NET0131  ;
	input \g392_reg/NET0131  ;
	input \g3990_reg/NET0131  ;
	input \g401_reg/NET0131  ;
	input \g4035_reg/NET0131  ;
	input \g4054_reg/NET0131  ;
	input \g4057_reg/NET0131  ;
	input \g405_reg/NET0131  ;
	input \g4064_reg/NET0131  ;
	input \g4072_reg/NET0131  ;
	input \g4076_reg/NET0131  ;
	input \g4082_reg/NET0131  ;
	input \g4087_reg/NET0131  ;
	input \g4093_reg/NET0131  ;
	input \g4098_reg/NET0131  ;
	input \g4104_reg/NET0131  ;
	input \g4108_reg/NET0131  ;
	input \g4112_reg/NET0131  ;
	input \g4116_reg/NET0131  ;
	input \g4119_reg/NET0131  ;
	input \g411_reg/NET0131  ;
	input \g4122_reg/NET0131  ;
	input \g4141_reg/NET0131  ;
	input \g4145_reg/NET0131  ;
	input \g4146_reg/NET0131  ;
	input \g4153_reg/NET0131  ;
	input \g4157_reg/NET0131  ;
	input \g4164_reg/NET0131  ;
	input \g4172_reg/NET0131  ;
	input \g4176_reg/NET0131  ;
	input \g417_reg/NET0131  ;
	input \g4180_reg/NET0131  ;
	input \g4235_reg/NET0131  ;
	input \g4239_reg/NET0131  ;
	input \g4242_reg/NET0131  ;
	input \g4245_reg/NET0131  ;
	input \g424_reg/NET0131  ;
	input \g4253_reg/NET0131  ;
	input \g4258_reg/NET0131  ;
	input \g4264_reg/NET0131  ;
	input \g4269_reg/NET0131  ;
	input \g4273_reg/NET0131  ;
	input \g4281_reg/NET0131  ;
	input \g4284_reg/NET0131  ;
	input \g4291_reg/NET0131  ;
	input \g4297_reg/NET0131  ;
	input \g4300_reg/NET0131  ;
	input \g4308_reg/NET0131  ;
	input \g4311_reg/NET0131  ;
	input \g4322_reg/NET0131  ;
	input \g4332_reg/NET0131  ;
	input \g433_reg/NET0131  ;
	input \g4340_reg/NET0131  ;
	input \g4349_reg/NET0131  ;
	input \g4358_reg/NET0131  ;
	input \g4366_reg/NET0131  ;
	input \g4369_reg/NET0131  ;
	input \g4372_reg/NET0131  ;
	input \g4375_reg/NET0131  ;
	input \g437_reg/NET0131  ;
	input \g4382_reg/NET0131  ;
	input \g4388_reg/NET0131  ;
	input \g4392_reg/NET0131  ;
	input \g4401_reg/NET0131  ;
	input \g4405_reg/NET0131  ;
	input \g4411_reg/NET0131  ;
	input \g4417_reg/NET0131  ;
	input \g441_reg/NET0131  ;
	input \g4420_reg/NET0131  ;
	input \g4423_reg/NET0131  ;
	input \g4427_reg/NET0131  ;
	input \g4430_reg/NET0131  ;
	input \g4434_reg/NET0131  ;
	input \g4438_reg/NET0131  ;
	input \g4443_reg/NET0131  ;
	input \g4452_reg/NET0131  ;
	input \g4455_reg/NET0131  ;
	input \g4459_reg/NET0131  ;
	input \g4462_reg/NET0131  ;
	input \g4467_reg/NET0131  ;
	input \g446_reg/NET0131  ;
	input \g4473_reg/NET0131  ;
	input \g4477_reg/NET0131  ;
	input \g4480_reg/NET0131  ;
	input \g4483_reg/NET0131  ;
	input \g4486_reg/NET0131  ;
	input \g4489_reg/NET0131  ;
	input \g4492_reg/NET0131  ;
	input \g4495_reg/NET0131  ;
	input \g4498_reg/NET0131  ;
	input \g4501_reg/NET0131  ;
	input \g4504_reg/NET0131  ;
	input \g4512_reg/NET0131  ;
	input \g4515_reg/NET0131  ;
	input \g4521_reg/NET0131  ;
	input \g4527_reg/NET0131  ;
	input \g452_reg/NET0131  ;
	input \g4531_reg/NET0131  ;
	input \g4534_reg/NET0131  ;
	input \g4540_reg/NET0131  ;
	input \g4543_reg/NET0131  ;
	input \g4546_reg/NET0131  ;
	input \g4549_reg/NET0131  ;
	input \g4552_reg/NET0131  ;
	input \g4555_reg/NET0131  ;
	input \g4558_reg/NET0131  ;
	input \g4561_reg/NET0131  ;
	input \g4564_reg/NET0131  ;
	input \g4567_reg/NET0131  ;
	input \g4572_reg/NET0131  ;
	input \g4575_reg/NET0131  ;
	input \g4581_reg/NET0131  ;
	input \g4584_reg/NET0131  ;
	input \g4593_reg/NET0131  ;
	input \g4601_reg/NET0131  ;
	input \g4608_reg/NET0131  ;
	input \g460_reg/NET0131  ;
	input \g4616_reg/NET0131  ;
	input \g4621_reg/NET0131  ;
	input \g4628_reg/NET0131  ;
	input \g4633_reg/NET0131  ;
	input \g4639_reg/NET0131  ;
	input \g4643_reg/NET0131  ;
	input \g4646_reg/NET0131  ;
	input \g4653_reg/NET0131  ;
	input \g4659_reg/NET0131  ;
	input \g4664_reg/NET0131  ;
	input \g4669_reg/NET0131  ;
	input \g4674_reg/NET0131  ;
	input \g4681_reg/NET0131  ;
	input \g4688_reg/NET0131  ;
	input \g4698_reg/NET0131  ;
	input \g4704_reg/NET0131  ;
	input \g4709_reg/NET0131  ;
	input \g4743_reg/NET0131  ;
	input \g4749_reg/NET0131  ;
	input \g4754_reg/NET0131  ;
	input \g475_reg/NET0131  ;
	input \g4760_reg/NET0131  ;
	input \g4765_reg/NET0131  ;
	input \g4771_reg/NET0131  ;
	input \g4776_reg/NET0131  ;
	input \g4785_reg/NET0131  ;
	input \g4793_reg/NET0131  ;
	input \g479_reg/NET0131  ;
	input \g4801_reg/NET0131  ;
	input \g482_reg/NET0131  ;
	input \g490_reg/NET0131  ;
	input \g496_reg/NET0131  ;
	input \g499_reg/NET0131  ;
	input \g5016_reg/NET0131  ;
	input \g5022_reg/NET0131  ;
	input \g5029_reg/NET0131  ;
	input \g5033_reg/NET0131  ;
	input \g5037_reg/NET0131  ;
	input \g5041_reg/NET0131  ;
	input \g5046_reg/NET0131  ;
	input \g504_reg/NET0131  ;
	input \g5052_reg/NET0131  ;
	input \g5057_reg/NET0131  ;
	input \g5069_reg/NET0131  ;
	input \g5073_reg/NET0131  ;
	input \g5077_reg/NET0131  ;
	input \g5080_reg/NET0131  ;
	input \g5084_reg/NET0131  ;
	input \g5092_reg/NET0131  ;
	input \g5097_reg/NET0131  ;
	input \g5101_reg/NET0131  ;
	input \g5112_reg/NET0131  ;
	input \g5115_reg/NET0131  ;
	input \g5124_reg/NET0131  ;
	input \g5128_reg/NET0131  ;
	input \g5134_reg/NET0131  ;
	input \g5138_reg/NET0131  ;
	input \g513_reg/NET0131  ;
	input \g5142_reg/NET0131  ;
	input \g5148_reg/NET0131  ;
	input \g5152_reg/NET0131  ;
	input \g518_reg/NET0131  ;
	input \g528_reg/NET0131  ;
	input \g5297_reg/NET0131  ;
	input \g534_reg/NET0131  ;
	input \g5357_reg/NET0131  ;
	input \g538_reg/NET0131  ;
	input \g542_reg/NET0131  ;
	input \g546_reg/NET0131  ;
	input \g550_reg/NET0131  ;
	input \g554_reg/NET0131  ;
	input \g645_reg/NET0131  ;
	input \g650_reg/NET0131  ;
	input \g655_reg/NET0131  ;
	input \g661_reg/NET0131  ;
	input \g667_reg/NET0131  ;
	input \g671_reg/NET0131  ;
	input \g676_reg/NET0131  ;
	input \g681_reg/NET0131  ;
	input \g686_reg/NET0131  ;
	input \g691_reg/NET0131  ;
	input \g699_reg/NET0131  ;
	input \g703_reg/NET0131  ;
	input \g714_reg/NET0131  ;
	input \g718_reg/NET0131  ;
	input \g723_reg/NET0131  ;
	input \g7243_pad  ;
	input \g7245_pad  ;
	input \g7257_pad  ;
	input \g7260_pad  ;
	input \g728_reg/NET0131  ;
	input \g732_reg/NET0131  ;
	input \g736_reg/NET0131  ;
	input \g739_reg/NET0131  ;
	input \g744_reg/NET0131  ;
	input \g749_reg/NET0131  ;
	input \g753_reg/NET0131  ;
	input \g7540_pad  ;
	input \g758_reg/NET0131  ;
	input \g763_reg/NET0131  ;
	input \g767_reg/NET0131  ;
	input \g772_reg/NET0131  ;
	input \g776_reg/NET0131  ;
	input \g781_reg/NET0131  ;
	input \g785_reg/NET0131  ;
	input \g790_reg/NET0131  ;
	input \g7916_pad  ;
	input \g7946_pad  ;
	input \g794_reg/NET0131  ;
	input \g802_reg/NET0131  ;
	input \g807_reg/NET0131  ;
	input \g812_reg/NET0131  ;
	input \g817_reg/NET0131  ;
	input \g822_reg/NET0131  ;
	input \g827_reg/NET0131  ;
	input \g8291_pad  ;
	input \g832_reg/NET0131  ;
	input \g8358_pad  ;
	input \g837_reg/NET0131  ;
	input \g8416_pad  ;
	input \g843_reg/NET0131  ;
	input \g8475_pad  ;
	input \g847_reg/NET0131  ;
	input \g854_reg/NET0131  ;
	input \g862_reg/NET0131  ;
	input \g8719_pad  ;
	input \g872_reg/NET0131  ;
	input \g8783_pad  ;
	input \g8784_pad  ;
	input \g8785_pad  ;
	input \g8786_pad  ;
	input \g8787_pad  ;
	input \g8788_pad  ;
	input \g8789_pad  ;
	input \g8839_pad  ;
	input \g8870_pad  ;
	input \g890_reg/NET0131  ;
	input \g8915_pad  ;
	input \g8916_pad  ;
	input \g8917_pad  ;
	input \g8918_pad  ;
	input \g8919_pad  ;
	input \g8920_pad  ;
	input \g896_reg/NET0131  ;
	input \g9019_pad  ;
	input \g9251_pad  ;
	input \g956_reg/NET0131  ;
	input \g962_reg/NET0131  ;
	input \g969_reg/NET0131  ;
	input \g976_reg/NET0131  ;
	input \g979_reg/NET0131  ;
	input \g990_reg/NET0131  ;
	input \g996_reg/NET0131  ;
	output \g136_reg/P0001  ;
	output \g21727_pad  ;
	output \g23190_pad  ;
	output \g26875_pad  ;
	output \g26876_pad  ;
	output \g26877_pad  ;
	output \g28041_pad  ;
	output \g28042_pad  ;
	output \g30327_pad  ;
	output \g30330_pad  ;
	output \g30331_pad  ;
	output \g31793_pad  ;
	output \g31860_pad  ;
	output \g31862_pad  ;
	output \g31863_pad  ;
	output \g32185_pad  ;
	output \g33079_pad  ;
	output \g33435_pad  ;
	output \g33959_pad  ;
	output \g34435_pad  ;
	output \g34788_pad  ;
	output \g34956_pad  ;
	output \g34_reg/P0001  ;
	output \g35_syn_2  ;
	output \g37/_0_  ;
	output \g41/_0_  ;
	output \g60853/_3_  ;
	output \g60856/_3_  ;
	output \g60879/_3_  ;
	output \g60882/_0_  ;
	output \g60888/_0_  ;
	output \g60891/_0_  ;
	output \g60896/_0_  ;
	output \g60899/_0_  ;
	output \g60900/_3_  ;
	output \g60909/_3_  ;
	output \g60911/_0_  ;
	output \g60915/_0_  ;
	output \g60918/_0_  ;
	output \g60919/_0_  ;
	output \g60928/_0_  ;
	output \g60929/_0_  ;
	output \g60936/_0_  ;
	output \g60937/_0_  ;
	output \g60939/_0_  ;
	output \g60940/_0_  ;
	output \g60941/_0_  ;
	output \g60942/_0_  ;
	output \g60943/_0_  ;
	output \g60944/_0_  ;
	output \g60952/_0_  ;
	output \g60954/_0_  ;
	output \g60958/_0_  ;
	output \g60962/_3_  ;
	output \g60972/_0_  ;
	output \g60980/_0_  ;
	output \g60984/_0_  ;
	output \g60986/_0_  ;
	output \g60989/_0_  ;
	output \g60991/_3_  ;
	output \g61006/_0_  ;
	output \g61008/_0_  ;
	output \g61013/_0_  ;
	output \g61014/_0_  ;
	output \g61015/_0_  ;
	output \g61016/_0_  ;
	output \g61017/_0_  ;
	output \g61026/_3_  ;
	output \g61027/_3_  ;
	output \g61030/_0_  ;
	output \g61031/_0_  ;
	output \g61037/_0_  ;
	output \g61038/_0_  ;
	output \g61042/_0_  ;
	output \g61044/_0_  ;
	output \g61045/_0_  ;
	output \g61046/_0_  ;
	output \g61050/_0_  ;
	output \g61051/_0_  ;
	output \g61052/_0_  ;
	output \g61078/_0_  ;
	output \g61131/_0_  ;
	output \g61137/_3_  ;
	output \g61142/_3_  ;
	output \g61143/_3_  ;
	output \g61151/_0_  ;
	output \g61152/_0_  ;
	output \g61161/_0_  ;
	output \g61168/_3_  ;
	output \g61169/_3_  ;
	output \g61170/_0_  ;
	output \g61171/_3_  ;
	output \g61172/_0_  ;
	output \g61173/_0_  ;
	output \g61174/_0_  ;
	output \g61175/_0_  ;
	output \g61176/_0_  ;
	output \g61177/_3_  ;
	output \g61178/_0_  ;
	output \g61179/_0_  ;
	output \g61180/_0_  ;
	output \g61181/_0_  ;
	output \g61182/_3_  ;
	output \g61183/_0_  ;
	output \g61184/_3_  ;
	output \g61185/_0_  ;
	output \g61186/_0_  ;
	output \g61187/_0_  ;
	output \g61188/_0_  ;
	output \g61189/_0_  ;
	output \g61190/_3_  ;
	output \g61191/_0_  ;
	output \g61192/_0_  ;
	output \g61193/_0_  ;
	output \g61194/_0_  ;
	output \g61221/_0_  ;
	output \g61222/_0_  ;
	output \g61223/_3_  ;
	output \g61224/_3_  ;
	output \g61261/_0_  ;
	output \g61295/_3_  ;
	output \g61308/_0_  ;
	output \g61316/_0_  ;
	output \g61327/_0_  ;
	output \g61329/_0_  ;
	output \g61330/_0_  ;
	output \g61331/_0_  ;
	output \g61332/_3_  ;
	output \g61333/_0_  ;
	output \g61334/_0_  ;
	output \g61335/_0_  ;
	output \g61336/_0_  ;
	output \g61337/_0_  ;
	output \g61338/_3_  ;
	output \g61339/_0_  ;
	output \g61340/_0_  ;
	output \g61341/_0_  ;
	output \g61342/_0_  ;
	output \g61343/_0_  ;
	output \g61344/_3_  ;
	output \g61345/_0_  ;
	output \g61346/_0_  ;
	output \g61347/_0_  ;
	output \g61348/_0_  ;
	output \g61349/_0_  ;
	output \g61350/_3_  ;
	output \g61351/_0_  ;
	output \g61352/_0_  ;
	output \g61353/_0_  ;
	output \g61354/_0_  ;
	output \g61367/_0_  ;
	output \g61372/_0_  ;
	output \g61373/_0_  ;
	output \g61375/_0_  ;
	output \g61382/_0_  ;
	output \g61385/_3_  ;
	output \g61386/_0_  ;
	output \g61399/_0_  ;
	output \g61400/_0_  ;
	output \g61402/_0_  ;
	output \g61405/_0_  ;
	output \g61435/_3_  ;
	output \g61449/_0_  ;
	output \g61468/_0_  ;
	output \g61475/_0_  ;
	output \g61480/_0_  ;
	output \g61482/_0_  ;
	output \g61483/_0_  ;
	output \g61484/_0_  ;
	output \g61486/_3_  ;
	output \g61494/_0_  ;
	output \g61496/_0_  ;
	output \g61497/_0_  ;
	output \g61514/_0_  ;
	output \g61517/_0_  ;
	output \g61519/_3_  ;
	output \g61520/_3_  ;
	output \g61527/_0_  ;
	output \g61541/_0_  ;
	output \g61544/_0_  ;
	output \g61550/_0_  ;
	output \g61551/_0_  ;
	output \g61554/_0_  ;
	output \g61556/_3_  ;
	output \g61567/_0_  ;
	output \g61571/_0_  ;
	output \g61574/_0_  ;
	output \g61587/_0_  ;
	output \g61592/_0_  ;
	output \g61632/_0_  ;
	output \g61634/_0_  ;
	output \g61635/_0_  ;
	output \g61639/_0_  ;
	output \g61644/_0_  ;
	output \g61652/_3_  ;
	output \g61709/_0_  ;
	output \g61714/_0_  ;
	output \g61720/_0_  ;
	output \g61721/_0_  ;
	output \g61723/_0_  ;
	output \g61725/_0_  ;
	output \g61726/_0_  ;
	output \g61734/_0_  ;
	output \g61739/_0_  ;
	output \g61744/_0_  ;
	output \g61746/_3_  ;
	output \g61747/_3_  ;
	output \g61748/_3_  ;
	output \g61750/u3_syn_7  ;
	output \g61802/_0_  ;
	output \g61804/_0_  ;
	output \g61808/_0_  ;
	output \g61811/_0_  ;
	output \g61816/_0_  ;
	output \g61818/_0_  ;
	output \g61820/_0_  ;
	output \g61823/_0_  ;
	output \g61824/_0_  ;
	output \g61841/_0_  ;
	output \g61842/_3_  ;
	output \g61844/_3_  ;
	output \g61845/_3_  ;
	output \g61846/_3_  ;
	output \g61847/u3_syn_7  ;
	output \g61848/_0_  ;
	output \g61849/_3_  ;
	output \g61850/_0_  ;
	output \g61851/u3_syn_7  ;
	output \g61852/_0_  ;
	output \g61853/_3_  ;
	output \g61854/_3_  ;
	output \g61855/_0_  ;
	output \g61856/u3_syn_7  ;
	output \g61857/_0_  ;
	output \g61858/_3_  ;
	output \g61859/_3_  ;
	output \g61860/u3_syn_7  ;
	output \g61861/_0_  ;
	output \g61862/_3_  ;
	output \g61863/_3_  ;
	output \g61864/u3_syn_7  ;
	output \g61865/_0_  ;
	output \g61866/_3_  ;
	output \g61867/_3_  ;
	output \g61868/u3_syn_7  ;
	output \g61869/_0_  ;
	output \g61870/_0_  ;
	output \g61871/_3_  ;
	output \g61872/_3_  ;
	output \g61873/u3_syn_7  ;
	output \g61874/_0_  ;
	output \g61875/_0_  ;
	output \g61877/_3_  ;
	output \g61878/_3_  ;
	output \g61879/u3_syn_7  ;
	output \g61880/_0_  ;
	output \g61881/_0_  ;
	output \g61882/_0_  ;
	output \g61883/_0_  ;
	output \g61884/_0_  ;
	output \g61914/_0_  ;
	output \g61915/_0_  ;
	output \g61917/_0_  ;
	output \g61918/_0_  ;
	output \g61922/_0_  ;
	output \g61923/_0_  ;
	output \g61924/_0_  ;
	output \g61932/_0_  ;
	output \g61936/_0_  ;
	output \g61945/_0_  ;
	output \g61947/_0_  ;
	output \g61959/_0_  ;
	output \g61960/_0_  ;
	output \g61962/_0_  ;
	output \g61973/_3_  ;
	output \g61974/u3_syn_7  ;
	output \g61975/_3_  ;
	output \g61976/u3_syn_7  ;
	output \g61977/_3_  ;
	output \g61978/_3_  ;
	output \g61979/u3_syn_7  ;
	output \g61980/_3_  ;
	output \g61981/_3_  ;
	output \g61982/_3_  ;
	output \g61983/u3_syn_7  ;
	output \g61984/_3_  ;
	output \g61985/_3_  ;
	output \g61986/u3_syn_7  ;
	output \g61987/_3_  ;
	output \g61988/_3_  ;
	output \g61989/u3_syn_7  ;
	output \g61990/_3_  ;
	output \g61991/_3_  ;
	output \g61992/u3_syn_7  ;
	output \g61993/_3_  ;
	output \g61994/u3_syn_7  ;
	output \g61995/_3_  ;
	output \g61996/_3_  ;
	output \g61997/_3_  ;
	output \g62022/_0_  ;
	output \g62028/_0_  ;
	output \g62029/_0_  ;
	output \g62031/_0_  ;
	output \g62033/_0_  ;
	output \g62038/_0_  ;
	output \g62042/_0_  ;
	output \g62046/_0_  ;
	output \g62048/_0_  ;
	output \g62049/_0_  ;
	output \g62051/_0_  ;
	output \g62053/_0_  ;
	output \g62085/_0_  ;
	output \g62101/_0_  ;
	output \g62102/_0_  ;
	output \g62103/_0_  ;
	output \g62105/_0_  ;
	output \g62108/_3_  ;
	output \g62112/_0_  ;
	output \g62137/_3_  ;
	output \g62207/_0_  ;
	output \g62239/_0_  ;
	output \g62240/_0_  ;
	output \g62267/_0_  ;
	output \g62273/_0_  ;
	output \g62284/_0_  ;
	output \g62291/_0_  ;
	output \g62293/_0_  ;
	output \g62298/_0_  ;
	output \g62303/_3_  ;
	output \g62322/_3_  ;
	output \g62323/_3_  ;
	output \g62324/_3_  ;
	output \g62325/_3_  ;
	output \g62583/_0_  ;
	output \g62598/_0_  ;
	output \g62609/_0_  ;
	output \g62636/_0_  ;
	output \g62646/_0_  ;
	output \g62649/_0_  ;
	output \g62658/_0_  ;
	output \g62663/_0_  ;
	output \g62664/_0_  ;
	output \g62667/_0_  ;
	output \g62676/_0_  ;
	output \g62677/_0_  ;
	output \g62678/_3_  ;
	output \g62679/_0_  ;
	output \g62687/u3_syn_7  ;
	output \g62688/u3_syn_7  ;
	output \g62689/_0_  ;
	output \g62690/_3_  ;
	output \g62691/_3_  ;
	output \g62693/_0_  ;
	output \g62694/_3_  ;
	output \g62695/_3_  ;
	output \g62696/_3_  ;
	output \g62697/_3_  ;
	output \g62698/_3_  ;
	output \g62699/_3_  ;
	output \g62700/_3_  ;
	output \g62701/_3_  ;
	output \g62702/_3_  ;
	output \g62703/_3_  ;
	output \g62704/u3_syn_7  ;
	output \g62705/_0_  ;
	output \g62706/_3_  ;
	output \g62707/_3_  ;
	output \g62708/u3_syn_7  ;
	output \g62709/_0_  ;
	output \g62710/_3_  ;
	output \g62711/_3_  ;
	output \g62712/u3_syn_7  ;
	output \g62713/_0_  ;
	output \g62714/_3_  ;
	output \g62715/_0_  ;
	output \g62716/u3_syn_7  ;
	output \g62717/_0_  ;
	output \g62718/_3_  ;
	output \g62719/_0_  ;
	output \g62720/u3_syn_7  ;
	output \g62721/_0_  ;
	output \g62722/_3_  ;
	output \g62723/_0_  ;
	output \g62724/u3_syn_7  ;
	output \g62725/_0_  ;
	output \g62726/_3_  ;
	output \g62728/_0_  ;
	output \g62790/_0_  ;
	output \g62791/_0_  ;
	output \g62793/_0_  ;
	output \g62794/_0_  ;
	output \g62795/_0_  ;
	output \g62796/_0_  ;
	output \g62797/_0_  ;
	output \g62807/_0_  ;
	output \g62823/_0_  ;
	output \g62824/_0_  ;
	output \g62833/_0_  ;
	output \g62846/_0_  ;
	output \g62859/_0_  ;
	output \g62860/_0_  ;
	output \g62897/_0_  ;
	output \g62898/_0_  ;
	output \g62922/_3_  ;
	output \g62923/_0_  ;
	output \g62927/_0_  ;
	output \g62938/_3_  ;
	output \g62939/_3_  ;
	output \g62940/_3_  ;
	output \g62941/u3_syn_7  ;
	output \g62942/_0_  ;
	output \g62943/_3_  ;
	output \g62987/_3_  ;
	output \g62991/_3_  ;
	output \g63015/u3_syn_7  ;
	output \g63016/_0_  ;
	output \g63017/_3_  ;
	output \g63018/_3_  ;
	output \g63019/_3_  ;
	output \g63020/_3_  ;
	output \g63021/_3_  ;
	output \g63022/_3_  ;
	output \g63025/_3_  ;
	output \g63026/_3_  ;
	output \g63027/_3_  ;
	output \g63029/_3_  ;
	output \g63030/_3_  ;
	output \g63031/_3_  ;
	output \g63033/_3_  ;
	output \g63034/_3_  ;
	output \g63043/_3_  ;
	output \g63044/_3_  ;
	output \g63051/_3_  ;
	output \g63057/_3_  ;
	output \g63068/_3_  ;
	output \g63070/_3_  ;
	output \g63073/_3_  ;
	output \g63081/_3_  ;
	output \g63082/_3_  ;
	output \g63083/u3_syn_7  ;
	output \g63084/_3_  ;
	output \g63085/_0_  ;
	output \g63086/_3_  ;
	output \g63107/_3_  ;
	output \g63108/u3_syn_7  ;
	output \g63109/u3_syn_7  ;
	output \g63110/_0_  ;
	output \g63111/_3_  ;
	output \g63132/_3_  ;
	output \g63133/_3_  ;
	output \g63134/_3_  ;
	output \g63135/_3_  ;
	output \g63136/_3_  ;
	output \g63137/_3_  ;
	output \g63138/_3_  ;
	output \g63139/u3_syn_7  ;
	output \g63140/_3_  ;
	output \g63141/_3_  ;
	output \g63142/_3_  ;
	output \g63143/_3_  ;
	output \g63144/_3_  ;
	output \g63145/_3_  ;
	output \g63146/u3_syn_7  ;
	output \g63198/_0_  ;
	output \g63205/_0_  ;
	output \g63208/_0_  ;
	output \g63212/_0_  ;
	output \g63215/_0_  ;
	output \g63219/_0_  ;
	output \g63244/_0_  ;
	output \g63246/_0_  ;
	output \g63254/_0_  ;
	output \g63255/_0_  ;
	output \g63272/_0_  ;
	output \g63276/_0_  ;
	output \g63278/_0_  ;
	output \g63279/_0_  ;
	output \g63280/_0_  ;
	output \g63327/_0_  ;
	output \g63345/_0_  ;
	output \g63346/_3_  ;
	output \g63347/_3_  ;
	output \g63354/_3_  ;
	output \g63358/_3_  ;
	output \g63359/u3_syn_7  ;
	output \g63361/_3_  ;
	output \g63365/_3_  ;
	output \g63366/_3_  ;
	output \g63367/_3_  ;
	output \g63368/_3_  ;
	output \g63370/_3_  ;
	output \g63479/_0_  ;
	output \g63484/_0_  ;
	output \g63499/_1_  ;
	output \g63520/_0_  ;
	output \g63523/_0_  ;
	output \g63526/_0_  ;
	output \g63538/_0_  ;
	output \g63539/_0_  ;
	output \g63541/_0_  ;
	output \g63555/_0_  ;
	output \g63642/_0_  ;
	output \g63645/_0_  ;
	output \g63648/_3_  ;
	output \g63777/_3_  ;
	output \g63778/_3_  ;
	output \g63781/_0_  ;
	output \g63786/u3_syn_7  ;
	output \g63787/_3_  ;
	output \g63788/_3_  ;
	output \g63790/_3_  ;
	output \g63791/_3_  ;
	output \g63792/u3_syn_7  ;
	output \g63794/_0_  ;
	output \g63795/_0_  ;
	output \g63796/_0_  ;
	output \g63798/_3_  ;
	output \g63800/_3_  ;
	output \g63804/_3_  ;
	output \g63805/_3_  ;
	output \g63806/_3_  ;
	output \g63807/_3_  ;
	output \g63808/_3_  ;
	output \g63809/_3_  ;
	output \g63870/_0_  ;
	output \g63883/_0_  ;
	output \g63934/_0_  ;
	output \g63936/_0_  ;
	output \g63938/_0_  ;
	output \g63939/_0_  ;
	output \g63966/_0_  ;
	output \g63970/_0_  ;
	output \g63999/_0_  ;
	output \g64039/_0_  ;
	output \g64040/_0_  ;
	output \g64043/_0_  ;
	output \g64062/_3_  ;
	output \g64078/_0_  ;
	output \g64091/_0_  ;
	output \g64095/_3_  ;
	output \g64096/_3_  ;
	output \g64097/u3_syn_7  ;
	output \g64098/u3_syn_7  ;
	output \g64099/u3_syn_7  ;
	output \g64100/u3_syn_7  ;
	output \g64134/_0_  ;
	output \g64135/_0_  ;
	output \g64153/_0_  ;
	output \g64155/_0_  ;
	output \g64179/_0_  ;
	output \g64229/_0_  ;
	output \g64235/_0_  ;
	output \g64236/_0_  ;
	output \g64280/_0_  ;
	output \g64315/_0_  ;
	output \g64365/_0_  ;
	output \g64426/_3_  ;
	output \g64438/_3_  ;
	output \g64442/u3_syn_7  ;
	output \g64445/_3_  ;
	output \g64447/_3_  ;
	output \g64449/_3_  ;
	output \g64451/_3_  ;
	output \g64453/_3_  ;
	output \g64454/_3_  ;
	output \g64460/_3_  ;
	output \g64461/_3_  ;
	output \g64510/_0_  ;
	output \g64527/_0_  ;
	output \g64528/_0_  ;
	output \g64544/_0_  ;
	output \g64549/_0_  ;
	output \g64566/_0_  ;
	output \g64576/_0_  ;
	output \g64602/_0_  ;
	output \g64691/_0_  ;
	output \g64697/_0_  ;
	output \g64707/_3_  ;
	output \g64778/_3_  ;
	output \g64790/_3_  ;
	output \g64791/_3_  ;
	output \g64792/_3_  ;
	output \g64793/_3_  ;
	output \g64794/_3_  ;
	output \g64795/_3_  ;
	output \g64796/_3_  ;
	output \g64797/_3_  ;
	output \g64877/_0_  ;
	output \g64912/_0_  ;
	output \g64973/_0_  ;
	output \g65047/_3_  ;
	output \g65081/_3_  ;
	output \g65088/_3_  ;
	output \g65097/_3_  ;
	output \g65100/_3_  ;
	output \g65101/_3_  ;
	output \g65104/_3_  ;
	output \g65105/_3_  ;
	output \g65107/_3_  ;
	output \g65110/_3_  ;
	output \g65111/_3_  ;
	output \g65113/_3_  ;
	output \g65114/_3_  ;
	output \g65266/_0_  ;
	output \g65267/_0_  ;
	output \g65294/_1_  ;
	output \g65328/_1_  ;
	output \g65495/_0_  ;
	output \g65499/_0_  ;
	output \g65503/_0_  ;
	output \g65529/_0_  ;
	output \g65530/_3_  ;
	output \g65531/_3_  ;
	output \g65532/_3_  ;
	output \g65533/_3_  ;
	output \g65624/_0_  ;
	output \g65625/_1_  ;
	output \g65641/_0_  ;
	output \g65701/_0_  ;
	output \g65704/_0_  ;
	output \g65853/_0_  ;
	output \g65891/_0_  ;
	output \g65901/_0_  ;
	output \g65986/_0_  ;
	output \g66029/_0_  ;
	output \g66066/_0_  ;
	output \g66067/_0_  ;
	output \g66068/_0_  ;
	output \g66154/_3_  ;
	output \g66362/_0_  ;
	output \g66369/_0_  ;
	output \g66398/_0_  ;
	output \g66409/_0_  ;
	output \g66419/_0_  ;
	output \g66439/_0_  ;
	output \g66443/_0_  ;
	output \g66464/_0_  ;
	output \g66471/_0_  ;
	output \g66512/_0_  ;
	output \g66528/_0_  ;
	output \g66541/_0_  ;
	output \g66558/_0_  ;
	output \g66644/_0_  ;
	output \g66684/_0_  ;
	output \g66697/_0_  ;
	output \g66698/_0_  ;
	output \g66701/_0_  ;
	output \g66714/_0_  ;
	output \g66715/_0_  ;
	output \g66745/_0_  ;
	output \g66750/_0_  ;
	output \g66751/_0_  ;
	output \g66810/_0_  ;
	output \g66844/_0_  ;
	output \g66853/_0_  ;
	output \g66897/_0_  ;
	output \g66905/_0_  ;
	output \g69743/_0_  ;
	output \g69750/_0_  ;
	output \g69773/_1_  ;
	output \g69792/_1_  ;
	output \g69858/_0_  ;
	output \g69938/_0_  ;
	output \g69949/_0_  ;
	output \g70167/_0_  ;
	output \g71190/_0_  ;
	output \g71198/_0_  ;
	output \g71284/_0_  ;
	output \g72369/_1_  ;
	output \g72467/_0_  ;
	output \g72476/_0_  ;
	output \g72477/_1_  ;
	output \g72648/_0_  ;
	output \g72741/_0_  ;
	output \g72772/_0_  ;
	output \g8132_pad  ;
	wire _w5177_ ;
	wire _w5176_ ;
	wire _w5175_ ;
	wire _w5174_ ;
	wire _w5173_ ;
	wire _w5172_ ;
	wire _w5171_ ;
	wire _w5170_ ;
	wire _w5169_ ;
	wire _w5168_ ;
	wire _w5167_ ;
	wire _w5166_ ;
	wire _w5165_ ;
	wire _w5164_ ;
	wire _w5163_ ;
	wire _w5162_ ;
	wire _w5161_ ;
	wire _w5160_ ;
	wire _w5159_ ;
	wire _w5158_ ;
	wire _w5157_ ;
	wire _w5156_ ;
	wire _w5155_ ;
	wire _w5154_ ;
	wire _w5153_ ;
	wire _w5152_ ;
	wire _w5151_ ;
	wire _w5150_ ;
	wire _w5149_ ;
	wire _w5148_ ;
	wire _w5147_ ;
	wire _w5146_ ;
	wire _w5145_ ;
	wire _w5144_ ;
	wire _w5143_ ;
	wire _w5142_ ;
	wire _w5141_ ;
	wire _w5140_ ;
	wire _w5139_ ;
	wire _w5138_ ;
	wire _w5137_ ;
	wire _w5136_ ;
	wire _w5135_ ;
	wire _w5134_ ;
	wire _w5133_ ;
	wire _w5132_ ;
	wire _w5131_ ;
	wire _w5130_ ;
	wire _w5129_ ;
	wire _w5128_ ;
	wire _w5127_ ;
	wire _w5126_ ;
	wire _w5125_ ;
	wire _w5124_ ;
	wire _w5123_ ;
	wire _w5122_ ;
	wire _w5121_ ;
	wire _w5120_ ;
	wire _w5119_ ;
	wire _w5118_ ;
	wire _w5117_ ;
	wire _w5116_ ;
	wire _w5115_ ;
	wire _w5114_ ;
	wire _w5113_ ;
	wire _w5112_ ;
	wire _w5111_ ;
	wire _w5110_ ;
	wire _w5109_ ;
	wire _w5108_ ;
	wire _w5107_ ;
	wire _w5106_ ;
	wire _w5105_ ;
	wire _w5104_ ;
	wire _w5103_ ;
	wire _w5102_ ;
	wire _w5101_ ;
	wire _w5100_ ;
	wire _w5099_ ;
	wire _w5098_ ;
	wire _w5097_ ;
	wire _w5096_ ;
	wire _w5095_ ;
	wire _w5094_ ;
	wire _w5093_ ;
	wire _w5092_ ;
	wire _w5091_ ;
	wire _w5090_ ;
	wire _w5089_ ;
	wire _w5088_ ;
	wire _w5087_ ;
	wire _w5086_ ;
	wire _w5085_ ;
	wire _w5084_ ;
	wire _w5083_ ;
	wire _w5082_ ;
	wire _w5081_ ;
	wire _w5080_ ;
	wire _w5079_ ;
	wire _w5078_ ;
	wire _w5077_ ;
	wire _w5076_ ;
	wire _w5075_ ;
	wire _w5074_ ;
	wire _w5073_ ;
	wire _w5072_ ;
	wire _w5071_ ;
	wire _w5070_ ;
	wire _w5069_ ;
	wire _w5068_ ;
	wire _w5067_ ;
	wire _w5066_ ;
	wire _w5065_ ;
	wire _w5064_ ;
	wire _w5063_ ;
	wire _w5062_ ;
	wire _w5061_ ;
	wire _w5060_ ;
	wire _w5059_ ;
	wire _w5058_ ;
	wire _w5057_ ;
	wire _w5056_ ;
	wire _w5055_ ;
	wire _w5054_ ;
	wire _w5053_ ;
	wire _w5052_ ;
	wire _w5051_ ;
	wire _w5050_ ;
	wire _w5049_ ;
	wire _w5048_ ;
	wire _w5047_ ;
	wire _w5046_ ;
	wire _w5045_ ;
	wire _w5044_ ;
	wire _w5043_ ;
	wire _w5042_ ;
	wire _w5041_ ;
	wire _w5040_ ;
	wire _w5039_ ;
	wire _w5038_ ;
	wire _w5037_ ;
	wire _w5036_ ;
	wire _w5035_ ;
	wire _w5034_ ;
	wire _w5033_ ;
	wire _w5032_ ;
	wire _w5031_ ;
	wire _w5030_ ;
	wire _w5029_ ;
	wire _w5028_ ;
	wire _w5027_ ;
	wire _w5026_ ;
	wire _w5025_ ;
	wire _w5024_ ;
	wire _w5023_ ;
	wire _w5022_ ;
	wire _w5021_ ;
	wire _w5020_ ;
	wire _w5019_ ;
	wire _w5018_ ;
	wire _w5017_ ;
	wire _w5016_ ;
	wire _w5015_ ;
	wire _w5014_ ;
	wire _w5013_ ;
	wire _w5012_ ;
	wire _w5011_ ;
	wire _w5010_ ;
	wire _w5009_ ;
	wire _w5008_ ;
	wire _w5007_ ;
	wire _w5006_ ;
	wire _w5005_ ;
	wire _w5004_ ;
	wire _w5003_ ;
	wire _w5002_ ;
	wire _w5001_ ;
	wire _w5000_ ;
	wire _w4999_ ;
	wire _w4998_ ;
	wire _w4997_ ;
	wire _w4996_ ;
	wire _w4995_ ;
	wire _w4994_ ;
	wire _w4993_ ;
	wire _w4992_ ;
	wire _w4991_ ;
	wire _w4990_ ;
	wire _w4989_ ;
	wire _w4988_ ;
	wire _w4987_ ;
	wire _w4986_ ;
	wire _w4985_ ;
	wire _w4984_ ;
	wire _w4983_ ;
	wire _w4982_ ;
	wire _w4981_ ;
	wire _w4980_ ;
	wire _w4979_ ;
	wire _w4978_ ;
	wire _w4977_ ;
	wire _w4976_ ;
	wire _w4975_ ;
	wire _w4974_ ;
	wire _w4973_ ;
	wire _w4972_ ;
	wire _w4971_ ;
	wire _w4970_ ;
	wire _w4969_ ;
	wire _w4968_ ;
	wire _w4967_ ;
	wire _w4966_ ;
	wire _w4965_ ;
	wire _w4964_ ;
	wire _w4963_ ;
	wire _w4962_ ;
	wire _w4961_ ;
	wire _w4960_ ;
	wire _w4959_ ;
	wire _w4958_ ;
	wire _w4957_ ;
	wire _w4956_ ;
	wire _w4955_ ;
	wire _w4954_ ;
	wire _w4953_ ;
	wire _w4952_ ;
	wire _w4951_ ;
	wire _w4950_ ;
	wire _w4949_ ;
	wire _w4948_ ;
	wire _w4947_ ;
	wire _w4946_ ;
	wire _w4945_ ;
	wire _w4944_ ;
	wire _w4943_ ;
	wire _w4942_ ;
	wire _w4941_ ;
	wire _w4940_ ;
	wire _w4939_ ;
	wire _w4938_ ;
	wire _w4937_ ;
	wire _w4936_ ;
	wire _w4935_ ;
	wire _w4934_ ;
	wire _w4933_ ;
	wire _w4932_ ;
	wire _w4931_ ;
	wire _w4930_ ;
	wire _w4929_ ;
	wire _w4928_ ;
	wire _w4927_ ;
	wire _w4926_ ;
	wire _w4925_ ;
	wire _w4924_ ;
	wire _w4923_ ;
	wire _w4922_ ;
	wire _w4921_ ;
	wire _w4920_ ;
	wire _w4919_ ;
	wire _w4918_ ;
	wire _w4917_ ;
	wire _w4916_ ;
	wire _w4915_ ;
	wire _w4914_ ;
	wire _w4913_ ;
	wire _w4912_ ;
	wire _w4911_ ;
	wire _w4910_ ;
	wire _w4909_ ;
	wire _w4908_ ;
	wire _w4907_ ;
	wire _w4906_ ;
	wire _w4905_ ;
	wire _w4904_ ;
	wire _w4903_ ;
	wire _w4902_ ;
	wire _w4901_ ;
	wire _w4900_ ;
	wire _w4899_ ;
	wire _w4898_ ;
	wire _w4897_ ;
	wire _w4896_ ;
	wire _w4895_ ;
	wire _w4894_ ;
	wire _w4893_ ;
	wire _w4892_ ;
	wire _w4891_ ;
	wire _w4890_ ;
	wire _w4889_ ;
	wire _w4888_ ;
	wire _w4887_ ;
	wire _w4886_ ;
	wire _w4885_ ;
	wire _w4884_ ;
	wire _w4883_ ;
	wire _w4882_ ;
	wire _w4881_ ;
	wire _w4880_ ;
	wire _w4879_ ;
	wire _w4878_ ;
	wire _w4877_ ;
	wire _w4876_ ;
	wire _w4875_ ;
	wire _w4874_ ;
	wire _w4873_ ;
	wire _w4872_ ;
	wire _w4871_ ;
	wire _w4870_ ;
	wire _w4869_ ;
	wire _w4868_ ;
	wire _w4867_ ;
	wire _w4866_ ;
	wire _w4865_ ;
	wire _w4864_ ;
	wire _w4863_ ;
	wire _w4862_ ;
	wire _w4861_ ;
	wire _w4860_ ;
	wire _w4859_ ;
	wire _w4858_ ;
	wire _w4857_ ;
	wire _w4856_ ;
	wire _w4855_ ;
	wire _w4854_ ;
	wire _w4853_ ;
	wire _w4852_ ;
	wire _w4851_ ;
	wire _w4850_ ;
	wire _w4849_ ;
	wire _w4848_ ;
	wire _w4847_ ;
	wire _w4846_ ;
	wire _w4845_ ;
	wire _w4844_ ;
	wire _w4843_ ;
	wire _w4842_ ;
	wire _w4841_ ;
	wire _w4840_ ;
	wire _w4839_ ;
	wire _w4838_ ;
	wire _w4837_ ;
	wire _w4836_ ;
	wire _w4835_ ;
	wire _w4834_ ;
	wire _w4833_ ;
	wire _w4832_ ;
	wire _w4831_ ;
	wire _w4830_ ;
	wire _w4829_ ;
	wire _w4828_ ;
	wire _w4827_ ;
	wire _w4826_ ;
	wire _w4825_ ;
	wire _w4824_ ;
	wire _w4823_ ;
	wire _w4822_ ;
	wire _w4821_ ;
	wire _w4820_ ;
	wire _w4819_ ;
	wire _w4818_ ;
	wire _w4817_ ;
	wire _w4816_ ;
	wire _w4815_ ;
	wire _w4814_ ;
	wire _w4813_ ;
	wire _w4812_ ;
	wire _w4811_ ;
	wire _w4810_ ;
	wire _w4809_ ;
	wire _w4808_ ;
	wire _w4807_ ;
	wire _w4806_ ;
	wire _w4805_ ;
	wire _w4804_ ;
	wire _w4803_ ;
	wire _w4802_ ;
	wire _w4801_ ;
	wire _w4800_ ;
	wire _w4799_ ;
	wire _w4798_ ;
	wire _w4797_ ;
	wire _w4796_ ;
	wire _w4795_ ;
	wire _w4794_ ;
	wire _w4793_ ;
	wire _w4792_ ;
	wire _w4791_ ;
	wire _w4790_ ;
	wire _w4789_ ;
	wire _w4788_ ;
	wire _w4787_ ;
	wire _w4786_ ;
	wire _w4785_ ;
	wire _w4784_ ;
	wire _w4783_ ;
	wire _w4782_ ;
	wire _w4781_ ;
	wire _w4780_ ;
	wire _w4779_ ;
	wire _w4778_ ;
	wire _w4777_ ;
	wire _w4776_ ;
	wire _w4775_ ;
	wire _w4774_ ;
	wire _w4773_ ;
	wire _w4772_ ;
	wire _w4771_ ;
	wire _w4770_ ;
	wire _w4769_ ;
	wire _w4768_ ;
	wire _w4767_ ;
	wire _w4766_ ;
	wire _w4765_ ;
	wire _w4764_ ;
	wire _w4763_ ;
	wire _w4762_ ;
	wire _w4761_ ;
	wire _w4760_ ;
	wire _w4759_ ;
	wire _w4758_ ;
	wire _w4757_ ;
	wire _w4756_ ;
	wire _w4755_ ;
	wire _w4754_ ;
	wire _w4753_ ;
	wire _w4752_ ;
	wire _w4751_ ;
	wire _w4750_ ;
	wire _w4749_ ;
	wire _w4748_ ;
	wire _w4747_ ;
	wire _w4746_ ;
	wire _w4745_ ;
	wire _w4744_ ;
	wire _w4743_ ;
	wire _w4742_ ;
	wire _w4741_ ;
	wire _w4740_ ;
	wire _w4739_ ;
	wire _w4738_ ;
	wire _w4737_ ;
	wire _w4736_ ;
	wire _w4735_ ;
	wire _w4734_ ;
	wire _w4733_ ;
	wire _w4732_ ;
	wire _w4731_ ;
	wire _w4730_ ;
	wire _w4729_ ;
	wire _w4728_ ;
	wire _w4727_ ;
	wire _w4726_ ;
	wire _w4725_ ;
	wire _w4724_ ;
	wire _w4723_ ;
	wire _w4722_ ;
	wire _w4721_ ;
	wire _w4720_ ;
	wire _w4719_ ;
	wire _w4718_ ;
	wire _w4717_ ;
	wire _w4716_ ;
	wire _w4715_ ;
	wire _w4714_ ;
	wire _w4713_ ;
	wire _w4712_ ;
	wire _w4711_ ;
	wire _w4710_ ;
	wire _w4709_ ;
	wire _w4708_ ;
	wire _w4707_ ;
	wire _w4706_ ;
	wire _w4705_ ;
	wire _w4704_ ;
	wire _w4703_ ;
	wire _w4702_ ;
	wire _w4701_ ;
	wire _w4700_ ;
	wire _w4699_ ;
	wire _w4698_ ;
	wire _w4697_ ;
	wire _w4696_ ;
	wire _w4695_ ;
	wire _w4694_ ;
	wire _w4693_ ;
	wire _w4692_ ;
	wire _w4691_ ;
	wire _w4690_ ;
	wire _w4689_ ;
	wire _w4688_ ;
	wire _w4687_ ;
	wire _w4686_ ;
	wire _w4685_ ;
	wire _w4684_ ;
	wire _w4683_ ;
	wire _w4682_ ;
	wire _w4681_ ;
	wire _w4680_ ;
	wire _w4679_ ;
	wire _w4678_ ;
	wire _w4677_ ;
	wire _w4676_ ;
	wire _w4675_ ;
	wire _w4674_ ;
	wire _w4673_ ;
	wire _w4672_ ;
	wire _w4671_ ;
	wire _w4670_ ;
	wire _w4669_ ;
	wire _w4668_ ;
	wire _w4667_ ;
	wire _w4666_ ;
	wire _w4665_ ;
	wire _w4664_ ;
	wire _w4663_ ;
	wire _w4662_ ;
	wire _w4661_ ;
	wire _w4660_ ;
	wire _w4659_ ;
	wire _w4658_ ;
	wire _w4657_ ;
	wire _w4656_ ;
	wire _w4655_ ;
	wire _w4654_ ;
	wire _w4653_ ;
	wire _w4652_ ;
	wire _w4651_ ;
	wire _w4650_ ;
	wire _w4649_ ;
	wire _w4648_ ;
	wire _w4647_ ;
	wire _w4646_ ;
	wire _w4645_ ;
	wire _w4644_ ;
	wire _w4643_ ;
	wire _w4642_ ;
	wire _w4641_ ;
	wire _w4640_ ;
	wire _w4639_ ;
	wire _w4638_ ;
	wire _w4637_ ;
	wire _w4636_ ;
	wire _w4635_ ;
	wire _w4634_ ;
	wire _w4633_ ;
	wire _w4632_ ;
	wire _w4631_ ;
	wire _w4630_ ;
	wire _w4629_ ;
	wire _w4628_ ;
	wire _w4627_ ;
	wire _w4626_ ;
	wire _w4625_ ;
	wire _w4624_ ;
	wire _w4623_ ;
	wire _w4622_ ;
	wire _w4621_ ;
	wire _w4620_ ;
	wire _w4619_ ;
	wire _w4618_ ;
	wire _w4617_ ;
	wire _w4616_ ;
	wire _w4615_ ;
	wire _w4614_ ;
	wire _w4613_ ;
	wire _w4612_ ;
	wire _w4611_ ;
	wire _w4610_ ;
	wire _w4609_ ;
	wire _w4608_ ;
	wire _w4607_ ;
	wire _w4606_ ;
	wire _w4605_ ;
	wire _w4604_ ;
	wire _w4603_ ;
	wire _w4602_ ;
	wire _w4601_ ;
	wire _w4600_ ;
	wire _w4599_ ;
	wire _w4598_ ;
	wire _w4597_ ;
	wire _w4596_ ;
	wire _w4595_ ;
	wire _w4594_ ;
	wire _w4593_ ;
	wire _w4592_ ;
	wire _w4591_ ;
	wire _w4590_ ;
	wire _w4589_ ;
	wire _w4588_ ;
	wire _w4587_ ;
	wire _w4586_ ;
	wire _w4585_ ;
	wire _w4584_ ;
	wire _w4583_ ;
	wire _w4582_ ;
	wire _w4581_ ;
	wire _w4580_ ;
	wire _w4579_ ;
	wire _w4578_ ;
	wire _w4577_ ;
	wire _w4576_ ;
	wire _w4575_ ;
	wire _w4574_ ;
	wire _w4573_ ;
	wire _w4572_ ;
	wire _w4571_ ;
	wire _w4570_ ;
	wire _w4569_ ;
	wire _w4568_ ;
	wire _w4567_ ;
	wire _w4566_ ;
	wire _w4565_ ;
	wire _w4564_ ;
	wire _w4563_ ;
	wire _w4562_ ;
	wire _w4561_ ;
	wire _w4560_ ;
	wire _w4559_ ;
	wire _w4558_ ;
	wire _w4557_ ;
	wire _w4556_ ;
	wire _w4555_ ;
	wire _w4554_ ;
	wire _w4553_ ;
	wire _w4552_ ;
	wire _w4551_ ;
	wire _w4550_ ;
	wire _w4549_ ;
	wire _w4548_ ;
	wire _w4547_ ;
	wire _w4546_ ;
	wire _w4545_ ;
	wire _w4544_ ;
	wire _w4543_ ;
	wire _w4542_ ;
	wire _w4541_ ;
	wire _w4540_ ;
	wire _w4539_ ;
	wire _w4538_ ;
	wire _w4537_ ;
	wire _w4536_ ;
	wire _w4535_ ;
	wire _w4534_ ;
	wire _w4533_ ;
	wire _w4532_ ;
	wire _w4531_ ;
	wire _w4530_ ;
	wire _w4529_ ;
	wire _w4528_ ;
	wire _w4527_ ;
	wire _w4526_ ;
	wire _w4525_ ;
	wire _w4524_ ;
	wire _w4523_ ;
	wire _w4522_ ;
	wire _w4521_ ;
	wire _w4520_ ;
	wire _w4519_ ;
	wire _w4518_ ;
	wire _w4517_ ;
	wire _w4516_ ;
	wire _w4515_ ;
	wire _w4514_ ;
	wire _w4513_ ;
	wire _w4512_ ;
	wire _w4511_ ;
	wire _w4510_ ;
	wire _w4509_ ;
	wire _w4508_ ;
	wire _w4507_ ;
	wire _w4506_ ;
	wire _w4505_ ;
	wire _w4504_ ;
	wire _w4503_ ;
	wire _w4502_ ;
	wire _w4501_ ;
	wire _w4500_ ;
	wire _w4499_ ;
	wire _w4498_ ;
	wire _w4497_ ;
	wire _w4496_ ;
	wire _w4495_ ;
	wire _w4494_ ;
	wire _w4493_ ;
	wire _w4492_ ;
	wire _w4491_ ;
	wire _w4490_ ;
	wire _w4489_ ;
	wire _w4488_ ;
	wire _w4487_ ;
	wire _w4486_ ;
	wire _w4485_ ;
	wire _w4484_ ;
	wire _w4483_ ;
	wire _w4482_ ;
	wire _w4481_ ;
	wire _w4480_ ;
	wire _w4479_ ;
	wire _w4478_ ;
	wire _w4477_ ;
	wire _w4476_ ;
	wire _w4475_ ;
	wire _w4474_ ;
	wire _w4473_ ;
	wire _w4472_ ;
	wire _w4471_ ;
	wire _w4470_ ;
	wire _w4469_ ;
	wire _w4468_ ;
	wire _w4467_ ;
	wire _w4466_ ;
	wire _w4465_ ;
	wire _w4464_ ;
	wire _w4463_ ;
	wire _w4462_ ;
	wire _w4461_ ;
	wire _w4460_ ;
	wire _w4459_ ;
	wire _w4458_ ;
	wire _w4457_ ;
	wire _w4456_ ;
	wire _w4455_ ;
	wire _w4454_ ;
	wire _w4453_ ;
	wire _w4452_ ;
	wire _w4451_ ;
	wire _w4450_ ;
	wire _w4449_ ;
	wire _w4448_ ;
	wire _w4447_ ;
	wire _w4446_ ;
	wire _w4445_ ;
	wire _w4444_ ;
	wire _w4443_ ;
	wire _w4442_ ;
	wire _w4441_ ;
	wire _w4440_ ;
	wire _w4439_ ;
	wire _w4438_ ;
	wire _w4437_ ;
	wire _w4436_ ;
	wire _w4435_ ;
	wire _w4434_ ;
	wire _w4433_ ;
	wire _w4432_ ;
	wire _w4431_ ;
	wire _w4430_ ;
	wire _w4429_ ;
	wire _w4428_ ;
	wire _w4427_ ;
	wire _w4426_ ;
	wire _w4425_ ;
	wire _w4424_ ;
	wire _w4423_ ;
	wire _w4422_ ;
	wire _w4421_ ;
	wire _w4420_ ;
	wire _w4419_ ;
	wire _w4418_ ;
	wire _w4417_ ;
	wire _w4416_ ;
	wire _w4415_ ;
	wire _w4414_ ;
	wire _w4413_ ;
	wire _w4412_ ;
	wire _w4411_ ;
	wire _w4410_ ;
	wire _w4409_ ;
	wire _w4408_ ;
	wire _w4407_ ;
	wire _w4406_ ;
	wire _w4405_ ;
	wire _w4404_ ;
	wire _w4403_ ;
	wire _w4402_ ;
	wire _w4401_ ;
	wire _w4400_ ;
	wire _w4399_ ;
	wire _w4398_ ;
	wire _w4397_ ;
	wire _w4396_ ;
	wire _w4395_ ;
	wire _w4394_ ;
	wire _w4393_ ;
	wire _w4392_ ;
	wire _w4391_ ;
	wire _w4390_ ;
	wire _w4389_ ;
	wire _w4388_ ;
	wire _w4387_ ;
	wire _w4386_ ;
	wire _w4385_ ;
	wire _w4384_ ;
	wire _w4383_ ;
	wire _w4382_ ;
	wire _w4381_ ;
	wire _w4380_ ;
	wire _w4379_ ;
	wire _w4378_ ;
	wire _w4377_ ;
	wire _w4376_ ;
	wire _w4375_ ;
	wire _w4374_ ;
	wire _w4373_ ;
	wire _w4372_ ;
	wire _w4371_ ;
	wire _w4370_ ;
	wire _w4369_ ;
	wire _w4368_ ;
	wire _w4367_ ;
	wire _w4366_ ;
	wire _w4365_ ;
	wire _w4364_ ;
	wire _w4363_ ;
	wire _w4362_ ;
	wire _w4361_ ;
	wire _w4360_ ;
	wire _w4359_ ;
	wire _w4358_ ;
	wire _w4357_ ;
	wire _w4356_ ;
	wire _w4355_ ;
	wire _w4354_ ;
	wire _w4353_ ;
	wire _w4352_ ;
	wire _w4351_ ;
	wire _w4350_ ;
	wire _w4349_ ;
	wire _w4348_ ;
	wire _w4347_ ;
	wire _w4346_ ;
	wire _w4345_ ;
	wire _w4344_ ;
	wire _w4343_ ;
	wire _w4342_ ;
	wire _w4341_ ;
	wire _w4340_ ;
	wire _w4339_ ;
	wire _w4338_ ;
	wire _w4337_ ;
	wire _w4336_ ;
	wire _w4335_ ;
	wire _w4334_ ;
	wire _w4333_ ;
	wire _w4332_ ;
	wire _w4331_ ;
	wire _w4330_ ;
	wire _w4329_ ;
	wire _w4328_ ;
	wire _w4327_ ;
	wire _w4326_ ;
	wire _w4325_ ;
	wire _w4324_ ;
	wire _w4323_ ;
	wire _w4322_ ;
	wire _w4321_ ;
	wire _w4320_ ;
	wire _w4319_ ;
	wire _w4318_ ;
	wire _w4317_ ;
	wire _w4316_ ;
	wire _w4315_ ;
	wire _w4314_ ;
	wire _w4313_ ;
	wire _w4312_ ;
	wire _w4311_ ;
	wire _w4310_ ;
	wire _w4309_ ;
	wire _w4308_ ;
	wire _w4307_ ;
	wire _w4306_ ;
	wire _w4305_ ;
	wire _w4304_ ;
	wire _w4303_ ;
	wire _w4302_ ;
	wire _w4301_ ;
	wire _w4300_ ;
	wire _w4299_ ;
	wire _w4298_ ;
	wire _w4297_ ;
	wire _w4296_ ;
	wire _w4295_ ;
	wire _w4294_ ;
	wire _w4293_ ;
	wire _w4292_ ;
	wire _w4291_ ;
	wire _w4290_ ;
	wire _w4289_ ;
	wire _w4288_ ;
	wire _w4287_ ;
	wire _w4286_ ;
	wire _w4285_ ;
	wire _w4284_ ;
	wire _w4283_ ;
	wire _w4282_ ;
	wire _w4281_ ;
	wire _w4280_ ;
	wire _w4279_ ;
	wire _w4278_ ;
	wire _w4277_ ;
	wire _w4276_ ;
	wire _w4275_ ;
	wire _w4274_ ;
	wire _w4273_ ;
	wire _w4272_ ;
	wire _w4271_ ;
	wire _w4270_ ;
	wire _w4269_ ;
	wire _w4268_ ;
	wire _w4267_ ;
	wire _w4266_ ;
	wire _w4265_ ;
	wire _w4264_ ;
	wire _w4263_ ;
	wire _w4262_ ;
	wire _w4261_ ;
	wire _w4260_ ;
	wire _w4259_ ;
	wire _w4258_ ;
	wire _w4257_ ;
	wire _w4256_ ;
	wire _w4255_ ;
	wire _w4254_ ;
	wire _w4253_ ;
	wire _w4252_ ;
	wire _w4251_ ;
	wire _w4250_ ;
	wire _w4249_ ;
	wire _w4248_ ;
	wire _w4247_ ;
	wire _w4246_ ;
	wire _w4245_ ;
	wire _w4244_ ;
	wire _w4243_ ;
	wire _w4242_ ;
	wire _w4241_ ;
	wire _w4240_ ;
	wire _w4239_ ;
	wire _w4238_ ;
	wire _w4237_ ;
	wire _w4236_ ;
	wire _w4235_ ;
	wire _w4234_ ;
	wire _w4233_ ;
	wire _w4232_ ;
	wire _w4231_ ;
	wire _w4230_ ;
	wire _w4229_ ;
	wire _w4228_ ;
	wire _w4227_ ;
	wire _w4226_ ;
	wire _w4225_ ;
	wire _w4224_ ;
	wire _w4223_ ;
	wire _w4222_ ;
	wire _w4221_ ;
	wire _w4220_ ;
	wire _w4219_ ;
	wire _w4218_ ;
	wire _w4217_ ;
	wire _w4216_ ;
	wire _w4215_ ;
	wire _w4214_ ;
	wire _w4213_ ;
	wire _w4212_ ;
	wire _w4211_ ;
	wire _w4210_ ;
	wire _w4209_ ;
	wire _w4208_ ;
	wire _w4207_ ;
	wire _w4206_ ;
	wire _w4205_ ;
	wire _w4204_ ;
	wire _w4203_ ;
	wire _w4202_ ;
	wire _w4201_ ;
	wire _w4200_ ;
	wire _w4199_ ;
	wire _w4198_ ;
	wire _w4197_ ;
	wire _w4196_ ;
	wire _w4195_ ;
	wire _w4194_ ;
	wire _w4193_ ;
	wire _w4192_ ;
	wire _w4191_ ;
	wire _w4190_ ;
	wire _w4189_ ;
	wire _w4188_ ;
	wire _w4187_ ;
	wire _w4186_ ;
	wire _w4185_ ;
	wire _w4184_ ;
	wire _w4183_ ;
	wire _w4182_ ;
	wire _w4181_ ;
	wire _w4180_ ;
	wire _w4179_ ;
	wire _w4178_ ;
	wire _w4177_ ;
	wire _w4176_ ;
	wire _w4175_ ;
	wire _w4174_ ;
	wire _w4173_ ;
	wire _w4172_ ;
	wire _w4171_ ;
	wire _w4170_ ;
	wire _w4169_ ;
	wire _w4168_ ;
	wire _w4167_ ;
	wire _w4166_ ;
	wire _w4165_ ;
	wire _w4164_ ;
	wire _w4163_ ;
	wire _w4162_ ;
	wire _w4161_ ;
	wire _w4160_ ;
	wire _w4159_ ;
	wire _w4158_ ;
	wire _w4157_ ;
	wire _w4156_ ;
	wire _w4155_ ;
	wire _w4154_ ;
	wire _w4153_ ;
	wire _w4152_ ;
	wire _w4151_ ;
	wire _w4150_ ;
	wire _w4149_ ;
	wire _w4148_ ;
	wire _w4147_ ;
	wire _w4146_ ;
	wire _w4145_ ;
	wire _w4144_ ;
	wire _w4143_ ;
	wire _w4142_ ;
	wire _w4141_ ;
	wire _w4140_ ;
	wire _w4139_ ;
	wire _w4138_ ;
	wire _w4137_ ;
	wire _w4136_ ;
	wire _w4135_ ;
	wire _w4134_ ;
	wire _w4133_ ;
	wire _w4132_ ;
	wire _w4131_ ;
	wire _w4130_ ;
	wire _w4129_ ;
	wire _w4128_ ;
	wire _w4127_ ;
	wire _w4126_ ;
	wire _w4125_ ;
	wire _w4124_ ;
	wire _w4123_ ;
	wire _w4122_ ;
	wire _w4121_ ;
	wire _w4120_ ;
	wire _w4119_ ;
	wire _w4118_ ;
	wire _w4117_ ;
	wire _w4116_ ;
	wire _w4115_ ;
	wire _w4114_ ;
	wire _w4113_ ;
	wire _w4112_ ;
	wire _w4111_ ;
	wire _w4110_ ;
	wire _w4109_ ;
	wire _w4108_ ;
	wire _w4107_ ;
	wire _w4106_ ;
	wire _w4105_ ;
	wire _w4104_ ;
	wire _w4103_ ;
	wire _w4102_ ;
	wire _w4101_ ;
	wire _w4100_ ;
	wire _w4099_ ;
	wire _w4098_ ;
	wire _w4097_ ;
	wire _w4096_ ;
	wire _w4095_ ;
	wire _w4094_ ;
	wire _w4093_ ;
	wire _w4092_ ;
	wire _w4091_ ;
	wire _w4090_ ;
	wire _w4089_ ;
	wire _w4088_ ;
	wire _w4087_ ;
	wire _w4086_ ;
	wire _w4085_ ;
	wire _w4084_ ;
	wire _w4083_ ;
	wire _w4082_ ;
	wire _w4081_ ;
	wire _w4080_ ;
	wire _w4079_ ;
	wire _w4078_ ;
	wire _w4077_ ;
	wire _w4076_ ;
	wire _w4075_ ;
	wire _w4074_ ;
	wire _w4073_ ;
	wire _w4072_ ;
	wire _w4071_ ;
	wire _w4070_ ;
	wire _w4069_ ;
	wire _w4068_ ;
	wire _w4067_ ;
	wire _w4066_ ;
	wire _w4065_ ;
	wire _w4064_ ;
	wire _w4063_ ;
	wire _w4062_ ;
	wire _w4061_ ;
	wire _w4060_ ;
	wire _w4059_ ;
	wire _w4058_ ;
	wire _w4057_ ;
	wire _w4056_ ;
	wire _w4055_ ;
	wire _w4054_ ;
	wire _w4053_ ;
	wire _w4052_ ;
	wire _w4051_ ;
	wire _w4050_ ;
	wire _w4049_ ;
	wire _w4048_ ;
	wire _w4047_ ;
	wire _w4046_ ;
	wire _w4045_ ;
	wire _w4044_ ;
	wire _w4043_ ;
	wire _w4042_ ;
	wire _w4041_ ;
	wire _w4040_ ;
	wire _w4039_ ;
	wire _w4038_ ;
	wire _w4037_ ;
	wire _w4036_ ;
	wire _w4035_ ;
	wire _w4034_ ;
	wire _w4033_ ;
	wire _w4032_ ;
	wire _w4031_ ;
	wire _w4030_ ;
	wire _w4029_ ;
	wire _w4028_ ;
	wire _w4027_ ;
	wire _w4026_ ;
	wire _w4025_ ;
	wire _w4024_ ;
	wire _w4023_ ;
	wire _w4022_ ;
	wire _w4021_ ;
	wire _w4020_ ;
	wire _w4019_ ;
	wire _w4018_ ;
	wire _w4017_ ;
	wire _w4016_ ;
	wire _w4015_ ;
	wire _w4014_ ;
	wire _w4013_ ;
	wire _w4012_ ;
	wire _w4011_ ;
	wire _w4010_ ;
	wire _w4009_ ;
	wire _w4008_ ;
	wire _w4007_ ;
	wire _w4006_ ;
	wire _w4005_ ;
	wire _w4004_ ;
	wire _w4003_ ;
	wire _w4002_ ;
	wire _w4001_ ;
	wire _w4000_ ;
	wire _w3999_ ;
	wire _w3998_ ;
	wire _w3997_ ;
	wire _w3996_ ;
	wire _w3995_ ;
	wire _w3994_ ;
	wire _w3993_ ;
	wire _w3992_ ;
	wire _w3991_ ;
	wire _w3990_ ;
	wire _w3989_ ;
	wire _w3988_ ;
	wire _w3987_ ;
	wire _w3986_ ;
	wire _w3985_ ;
	wire _w3984_ ;
	wire _w3983_ ;
	wire _w3982_ ;
	wire _w3981_ ;
	wire _w3980_ ;
	wire _w3979_ ;
	wire _w3978_ ;
	wire _w3977_ ;
	wire _w3976_ ;
	wire _w3975_ ;
	wire _w3974_ ;
	wire _w3973_ ;
	wire _w3972_ ;
	wire _w3971_ ;
	wire _w3970_ ;
	wire _w3969_ ;
	wire _w3968_ ;
	wire _w3967_ ;
	wire _w3966_ ;
	wire _w3965_ ;
	wire _w3964_ ;
	wire _w3963_ ;
	wire _w3962_ ;
	wire _w3961_ ;
	wire _w3960_ ;
	wire _w3959_ ;
	wire _w3958_ ;
	wire _w3957_ ;
	wire _w3956_ ;
	wire _w3955_ ;
	wire _w3954_ ;
	wire _w3953_ ;
	wire _w3952_ ;
	wire _w3951_ ;
	wire _w3950_ ;
	wire _w3949_ ;
	wire _w3948_ ;
	wire _w3947_ ;
	wire _w3946_ ;
	wire _w3945_ ;
	wire _w3944_ ;
	wire _w3943_ ;
	wire _w3942_ ;
	wire _w3941_ ;
	wire _w3940_ ;
	wire _w3939_ ;
	wire _w3938_ ;
	wire _w3937_ ;
	wire _w3936_ ;
	wire _w3935_ ;
	wire _w3934_ ;
	wire _w3933_ ;
	wire _w3932_ ;
	wire _w3931_ ;
	wire _w3930_ ;
	wire _w3929_ ;
	wire _w3928_ ;
	wire _w3927_ ;
	wire _w3926_ ;
	wire _w3925_ ;
	wire _w3924_ ;
	wire _w3923_ ;
	wire _w3922_ ;
	wire _w3921_ ;
	wire _w3920_ ;
	wire _w3919_ ;
	wire _w3918_ ;
	wire _w3917_ ;
	wire _w3916_ ;
	wire _w3915_ ;
	wire _w3914_ ;
	wire _w3913_ ;
	wire _w3912_ ;
	wire _w3911_ ;
	wire _w3910_ ;
	wire _w3909_ ;
	wire _w3908_ ;
	wire _w3907_ ;
	wire _w3906_ ;
	wire _w3905_ ;
	wire _w3904_ ;
	wire _w3903_ ;
	wire _w3902_ ;
	wire _w3901_ ;
	wire _w3900_ ;
	wire _w3899_ ;
	wire _w3898_ ;
	wire _w3897_ ;
	wire _w3896_ ;
	wire _w3895_ ;
	wire _w3894_ ;
	wire _w3893_ ;
	wire _w3892_ ;
	wire _w3891_ ;
	wire _w3890_ ;
	wire _w3889_ ;
	wire _w3888_ ;
	wire _w3887_ ;
	wire _w3886_ ;
	wire _w3885_ ;
	wire _w3884_ ;
	wire _w3883_ ;
	wire _w3882_ ;
	wire _w3881_ ;
	wire _w3880_ ;
	wire _w3879_ ;
	wire _w3878_ ;
	wire _w3877_ ;
	wire _w3876_ ;
	wire _w3875_ ;
	wire _w3874_ ;
	wire _w3873_ ;
	wire _w3872_ ;
	wire _w3871_ ;
	wire _w3870_ ;
	wire _w3869_ ;
	wire _w3868_ ;
	wire _w3867_ ;
	wire _w3866_ ;
	wire _w3865_ ;
	wire _w3864_ ;
	wire _w3863_ ;
	wire _w3862_ ;
	wire _w3861_ ;
	wire _w3860_ ;
	wire _w3859_ ;
	wire _w3858_ ;
	wire _w3857_ ;
	wire _w3856_ ;
	wire _w3855_ ;
	wire _w3854_ ;
	wire _w3853_ ;
	wire _w3852_ ;
	wire _w3851_ ;
	wire _w3850_ ;
	wire _w3849_ ;
	wire _w3848_ ;
	wire _w3847_ ;
	wire _w3846_ ;
	wire _w3845_ ;
	wire _w3844_ ;
	wire _w3843_ ;
	wire _w3842_ ;
	wire _w3841_ ;
	wire _w3840_ ;
	wire _w3839_ ;
	wire _w3838_ ;
	wire _w3837_ ;
	wire _w3836_ ;
	wire _w3835_ ;
	wire _w3834_ ;
	wire _w3833_ ;
	wire _w3832_ ;
	wire _w3831_ ;
	wire _w3830_ ;
	wire _w3829_ ;
	wire _w3828_ ;
	wire _w3827_ ;
	wire _w3826_ ;
	wire _w3825_ ;
	wire _w3824_ ;
	wire _w3823_ ;
	wire _w3822_ ;
	wire _w3821_ ;
	wire _w3820_ ;
	wire _w3819_ ;
	wire _w3818_ ;
	wire _w3817_ ;
	wire _w3816_ ;
	wire _w3815_ ;
	wire _w3814_ ;
	wire _w3813_ ;
	wire _w3812_ ;
	wire _w3811_ ;
	wire _w3810_ ;
	wire _w3809_ ;
	wire _w3808_ ;
	wire _w3807_ ;
	wire _w3806_ ;
	wire _w3805_ ;
	wire _w3804_ ;
	wire _w3803_ ;
	wire _w3802_ ;
	wire _w3801_ ;
	wire _w3800_ ;
	wire _w3799_ ;
	wire _w3798_ ;
	wire _w3797_ ;
	wire _w3796_ ;
	wire _w3795_ ;
	wire _w3794_ ;
	wire _w3793_ ;
	wire _w3792_ ;
	wire _w3791_ ;
	wire _w3790_ ;
	wire _w3789_ ;
	wire _w3788_ ;
	wire _w3787_ ;
	wire _w3786_ ;
	wire _w3785_ ;
	wire _w3784_ ;
	wire _w3783_ ;
	wire _w3782_ ;
	wire _w3781_ ;
	wire _w3780_ ;
	wire _w3779_ ;
	wire _w3778_ ;
	wire _w3777_ ;
	wire _w3776_ ;
	wire _w3775_ ;
	wire _w3774_ ;
	wire _w3773_ ;
	wire _w3772_ ;
	wire _w3771_ ;
	wire _w3770_ ;
	wire _w3769_ ;
	wire _w3768_ ;
	wire _w3767_ ;
	wire _w3766_ ;
	wire _w3765_ ;
	wire _w3764_ ;
	wire _w3763_ ;
	wire _w3762_ ;
	wire _w3761_ ;
	wire _w3760_ ;
	wire _w3759_ ;
	wire _w3758_ ;
	wire _w3757_ ;
	wire _w3756_ ;
	wire _w3755_ ;
	wire _w3754_ ;
	wire _w3753_ ;
	wire _w3752_ ;
	wire _w3751_ ;
	wire _w3750_ ;
	wire _w3749_ ;
	wire _w3748_ ;
	wire _w3747_ ;
	wire _w3746_ ;
	wire _w3745_ ;
	wire _w3744_ ;
	wire _w3743_ ;
	wire _w3742_ ;
	wire _w3741_ ;
	wire _w3740_ ;
	wire _w3739_ ;
	wire _w3738_ ;
	wire _w3737_ ;
	wire _w3736_ ;
	wire _w3735_ ;
	wire _w3734_ ;
	wire _w3733_ ;
	wire _w3732_ ;
	wire _w3731_ ;
	wire _w3730_ ;
	wire _w3729_ ;
	wire _w3728_ ;
	wire _w3727_ ;
	wire _w3726_ ;
	wire _w3725_ ;
	wire _w3724_ ;
	wire _w3723_ ;
	wire _w3722_ ;
	wire _w3721_ ;
	wire _w3720_ ;
	wire _w3719_ ;
	wire _w3718_ ;
	wire _w3717_ ;
	wire _w3716_ ;
	wire _w3715_ ;
	wire _w3714_ ;
	wire _w3713_ ;
	wire _w3712_ ;
	wire _w3711_ ;
	wire _w3710_ ;
	wire _w3709_ ;
	wire _w3708_ ;
	wire _w3707_ ;
	wire _w3706_ ;
	wire _w3705_ ;
	wire _w3704_ ;
	wire _w3703_ ;
	wire _w3702_ ;
	wire _w3701_ ;
	wire _w3700_ ;
	wire _w3699_ ;
	wire _w3698_ ;
	wire _w3697_ ;
	wire _w3696_ ;
	wire _w3695_ ;
	wire _w3694_ ;
	wire _w3693_ ;
	wire _w3692_ ;
	wire _w3691_ ;
	wire _w3690_ ;
	wire _w3689_ ;
	wire _w3688_ ;
	wire _w3687_ ;
	wire _w3686_ ;
	wire _w3685_ ;
	wire _w3684_ ;
	wire _w3683_ ;
	wire _w3682_ ;
	wire _w3681_ ;
	wire _w3680_ ;
	wire _w3679_ ;
	wire _w3678_ ;
	wire _w3677_ ;
	wire _w3676_ ;
	wire _w3675_ ;
	wire _w3674_ ;
	wire _w3673_ ;
	wire _w3672_ ;
	wire _w3671_ ;
	wire _w3670_ ;
	wire _w3669_ ;
	wire _w3668_ ;
	wire _w3667_ ;
	wire _w3666_ ;
	wire _w3665_ ;
	wire _w3664_ ;
	wire _w3663_ ;
	wire _w3662_ ;
	wire _w3661_ ;
	wire _w3660_ ;
	wire _w3659_ ;
	wire _w3658_ ;
	wire _w3657_ ;
	wire _w3656_ ;
	wire _w3655_ ;
	wire _w3654_ ;
	wire _w3653_ ;
	wire _w3652_ ;
	wire _w3651_ ;
	wire _w3650_ ;
	wire _w3649_ ;
	wire _w3648_ ;
	wire _w3647_ ;
	wire _w3646_ ;
	wire _w3645_ ;
	wire _w3644_ ;
	wire _w3643_ ;
	wire _w3642_ ;
	wire _w3641_ ;
	wire _w3640_ ;
	wire _w3639_ ;
	wire _w3638_ ;
	wire _w3637_ ;
	wire _w3636_ ;
	wire _w3635_ ;
	wire _w3634_ ;
	wire _w3633_ ;
	wire _w3632_ ;
	wire _w3631_ ;
	wire _w3630_ ;
	wire _w3629_ ;
	wire _w3628_ ;
	wire _w3627_ ;
	wire _w3626_ ;
	wire _w3625_ ;
	wire _w3624_ ;
	wire _w3623_ ;
	wire _w3622_ ;
	wire _w3621_ ;
	wire _w3620_ ;
	wire _w3619_ ;
	wire _w3618_ ;
	wire _w3617_ ;
	wire _w3616_ ;
	wire _w3615_ ;
	wire _w3614_ ;
	wire _w3613_ ;
	wire _w3612_ ;
	wire _w3611_ ;
	wire _w3610_ ;
	wire _w3609_ ;
	wire _w3608_ ;
	wire _w3607_ ;
	wire _w3606_ ;
	wire _w3605_ ;
	wire _w3604_ ;
	wire _w3603_ ;
	wire _w3602_ ;
	wire _w3601_ ;
	wire _w3600_ ;
	wire _w3599_ ;
	wire _w3598_ ;
	wire _w3597_ ;
	wire _w3596_ ;
	wire _w3595_ ;
	wire _w3594_ ;
	wire _w3593_ ;
	wire _w3592_ ;
	wire _w3591_ ;
	wire _w3590_ ;
	wire _w3589_ ;
	wire _w3588_ ;
	wire _w3587_ ;
	wire _w3586_ ;
	wire _w3585_ ;
	wire _w3584_ ;
	wire _w3583_ ;
	wire _w3582_ ;
	wire _w3581_ ;
	wire _w3580_ ;
	wire _w3579_ ;
	wire _w3578_ ;
	wire _w3577_ ;
	wire _w3576_ ;
	wire _w3575_ ;
	wire _w3574_ ;
	wire _w3573_ ;
	wire _w3572_ ;
	wire _w3571_ ;
	wire _w3570_ ;
	wire _w3569_ ;
	wire _w3568_ ;
	wire _w3567_ ;
	wire _w3566_ ;
	wire _w3565_ ;
	wire _w3564_ ;
	wire _w3563_ ;
	wire _w3562_ ;
	wire _w3561_ ;
	wire _w3560_ ;
	wire _w3559_ ;
	wire _w3558_ ;
	wire _w3557_ ;
	wire _w3556_ ;
	wire _w3555_ ;
	wire _w3554_ ;
	wire _w3553_ ;
	wire _w3552_ ;
	wire _w3551_ ;
	wire _w3550_ ;
	wire _w3549_ ;
	wire _w3548_ ;
	wire _w3547_ ;
	wire _w3546_ ;
	wire _w3545_ ;
	wire _w3544_ ;
	wire _w3543_ ;
	wire _w3542_ ;
	wire _w3541_ ;
	wire _w3540_ ;
	wire _w3539_ ;
	wire _w3538_ ;
	wire _w3537_ ;
	wire _w3536_ ;
	wire _w3535_ ;
	wire _w3534_ ;
	wire _w3533_ ;
	wire _w3532_ ;
	wire _w3531_ ;
	wire _w3530_ ;
	wire _w3529_ ;
	wire _w3528_ ;
	wire _w3527_ ;
	wire _w3526_ ;
	wire _w3525_ ;
	wire _w3524_ ;
	wire _w3523_ ;
	wire _w3522_ ;
	wire _w3521_ ;
	wire _w3520_ ;
	wire _w3519_ ;
	wire _w3518_ ;
	wire _w3517_ ;
	wire _w3516_ ;
	wire _w3515_ ;
	wire _w3514_ ;
	wire _w3513_ ;
	wire _w3512_ ;
	wire _w3511_ ;
	wire _w3510_ ;
	wire _w3509_ ;
	wire _w3508_ ;
	wire _w3507_ ;
	wire _w3506_ ;
	wire _w3505_ ;
	wire _w3504_ ;
	wire _w3503_ ;
	wire _w3502_ ;
	wire _w3501_ ;
	wire _w3500_ ;
	wire _w3499_ ;
	wire _w3498_ ;
	wire _w3497_ ;
	wire _w3496_ ;
	wire _w3495_ ;
	wire _w3494_ ;
	wire _w3493_ ;
	wire _w3492_ ;
	wire _w3491_ ;
	wire _w3490_ ;
	wire _w3489_ ;
	wire _w3488_ ;
	wire _w3487_ ;
	wire _w3486_ ;
	wire _w3485_ ;
	wire _w3484_ ;
	wire _w3483_ ;
	wire _w3482_ ;
	wire _w3481_ ;
	wire _w3480_ ;
	wire _w3479_ ;
	wire _w3478_ ;
	wire _w3477_ ;
	wire _w3476_ ;
	wire _w3475_ ;
	wire _w3474_ ;
	wire _w3473_ ;
	wire _w3472_ ;
	wire _w3471_ ;
	wire _w3470_ ;
	wire _w3469_ ;
	wire _w3468_ ;
	wire _w3467_ ;
	wire _w3466_ ;
	wire _w3465_ ;
	wire _w3464_ ;
	wire _w3463_ ;
	wire _w3462_ ;
	wire _w3461_ ;
	wire _w3460_ ;
	wire _w3459_ ;
	wire _w3458_ ;
	wire _w3457_ ;
	wire _w3456_ ;
	wire _w3455_ ;
	wire _w3454_ ;
	wire _w3453_ ;
	wire _w3452_ ;
	wire _w3451_ ;
	wire _w3450_ ;
	wire _w3449_ ;
	wire _w3448_ ;
	wire _w3447_ ;
	wire _w3446_ ;
	wire _w3445_ ;
	wire _w3444_ ;
	wire _w3443_ ;
	wire _w3442_ ;
	wire _w3441_ ;
	wire _w3440_ ;
	wire _w3439_ ;
	wire _w3438_ ;
	wire _w3437_ ;
	wire _w3436_ ;
	wire _w3435_ ;
	wire _w3434_ ;
	wire _w3433_ ;
	wire _w3432_ ;
	wire _w3431_ ;
	wire _w3430_ ;
	wire _w3429_ ;
	wire _w3428_ ;
	wire _w3427_ ;
	wire _w3426_ ;
	wire _w3425_ ;
	wire _w3424_ ;
	wire _w3423_ ;
	wire _w3422_ ;
	wire _w3421_ ;
	wire _w3420_ ;
	wire _w3419_ ;
	wire _w3418_ ;
	wire _w3417_ ;
	wire _w3416_ ;
	wire _w3415_ ;
	wire _w3414_ ;
	wire _w3413_ ;
	wire _w3412_ ;
	wire _w3411_ ;
	wire _w3410_ ;
	wire _w3409_ ;
	wire _w3408_ ;
	wire _w3407_ ;
	wire _w3406_ ;
	wire _w3405_ ;
	wire _w3404_ ;
	wire _w3403_ ;
	wire _w3402_ ;
	wire _w3401_ ;
	wire _w3400_ ;
	wire _w3399_ ;
	wire _w3398_ ;
	wire _w3397_ ;
	wire _w3396_ ;
	wire _w3395_ ;
	wire _w3394_ ;
	wire _w3393_ ;
	wire _w3392_ ;
	wire _w3391_ ;
	wire _w3390_ ;
	wire _w3389_ ;
	wire _w3388_ ;
	wire _w3387_ ;
	wire _w3386_ ;
	wire _w3385_ ;
	wire _w3384_ ;
	wire _w3383_ ;
	wire _w3382_ ;
	wire _w3381_ ;
	wire _w3380_ ;
	wire _w3379_ ;
	wire _w3378_ ;
	wire _w3377_ ;
	wire _w3376_ ;
	wire _w3375_ ;
	wire _w3374_ ;
	wire _w3373_ ;
	wire _w3372_ ;
	wire _w3371_ ;
	wire _w3370_ ;
	wire _w3369_ ;
	wire _w3368_ ;
	wire _w3367_ ;
	wire _w3366_ ;
	wire _w3365_ ;
	wire _w3364_ ;
	wire _w3363_ ;
	wire _w3362_ ;
	wire _w3361_ ;
	wire _w3360_ ;
	wire _w3359_ ;
	wire _w3358_ ;
	wire _w3357_ ;
	wire _w3356_ ;
	wire _w3355_ ;
	wire _w3354_ ;
	wire _w3353_ ;
	wire _w3352_ ;
	wire _w3351_ ;
	wire _w3350_ ;
	wire _w3349_ ;
	wire _w3348_ ;
	wire _w3347_ ;
	wire _w3346_ ;
	wire _w3345_ ;
	wire _w3344_ ;
	wire _w3343_ ;
	wire _w3342_ ;
	wire _w3341_ ;
	wire _w3340_ ;
	wire _w3339_ ;
	wire _w3338_ ;
	wire _w3337_ ;
	wire _w3336_ ;
	wire _w3335_ ;
	wire _w3334_ ;
	wire _w3333_ ;
	wire _w3332_ ;
	wire _w3331_ ;
	wire _w3330_ ;
	wire _w3329_ ;
	wire _w3328_ ;
	wire _w3327_ ;
	wire _w3326_ ;
	wire _w3325_ ;
	wire _w3324_ ;
	wire _w3323_ ;
	wire _w3322_ ;
	wire _w3321_ ;
	wire _w3320_ ;
	wire _w3319_ ;
	wire _w3318_ ;
	wire _w3317_ ;
	wire _w3316_ ;
	wire _w3315_ ;
	wire _w3314_ ;
	wire _w3313_ ;
	wire _w3312_ ;
	wire _w3311_ ;
	wire _w3310_ ;
	wire _w3309_ ;
	wire _w3308_ ;
	wire _w3307_ ;
	wire _w3306_ ;
	wire _w3305_ ;
	wire _w3304_ ;
	wire _w3303_ ;
	wire _w3302_ ;
	wire _w3301_ ;
	wire _w3300_ ;
	wire _w3299_ ;
	wire _w3298_ ;
	wire _w3297_ ;
	wire _w3296_ ;
	wire _w3295_ ;
	wire _w3294_ ;
	wire _w3293_ ;
	wire _w3292_ ;
	wire _w3291_ ;
	wire _w3290_ ;
	wire _w3289_ ;
	wire _w3288_ ;
	wire _w3287_ ;
	wire _w3286_ ;
	wire _w3285_ ;
	wire _w3284_ ;
	wire _w3283_ ;
	wire _w3282_ ;
	wire _w3281_ ;
	wire _w3280_ ;
	wire _w3279_ ;
	wire _w3278_ ;
	wire _w3277_ ;
	wire _w3276_ ;
	wire _w3275_ ;
	wire _w3274_ ;
	wire _w3273_ ;
	wire _w3272_ ;
	wire _w3271_ ;
	wire _w3270_ ;
	wire _w3269_ ;
	wire _w3268_ ;
	wire _w3267_ ;
	wire _w3266_ ;
	wire _w3265_ ;
	wire _w3264_ ;
	wire _w3263_ ;
	wire _w3262_ ;
	wire _w3261_ ;
	wire _w3260_ ;
	wire _w3259_ ;
	wire _w3258_ ;
	wire _w3257_ ;
	wire _w3256_ ;
	wire _w3255_ ;
	wire _w3254_ ;
	wire _w3253_ ;
	wire _w3252_ ;
	wire _w3251_ ;
	wire _w3250_ ;
	wire _w3249_ ;
	wire _w3248_ ;
	wire _w3247_ ;
	wire _w3246_ ;
	wire _w3245_ ;
	wire _w3244_ ;
	wire _w3243_ ;
	wire _w3242_ ;
	wire _w3241_ ;
	wire _w3240_ ;
	wire _w3239_ ;
	wire _w3238_ ;
	wire _w3237_ ;
	wire _w3236_ ;
	wire _w3235_ ;
	wire _w3234_ ;
	wire _w3233_ ;
	wire _w3232_ ;
	wire _w3231_ ;
	wire _w3230_ ;
	wire _w3229_ ;
	wire _w3228_ ;
	wire _w3227_ ;
	wire _w3226_ ;
	wire _w3225_ ;
	wire _w3224_ ;
	wire _w3223_ ;
	wire _w3222_ ;
	wire _w3221_ ;
	wire _w3220_ ;
	wire _w3219_ ;
	wire _w3218_ ;
	wire _w3217_ ;
	wire _w3216_ ;
	wire _w3215_ ;
	wire _w3214_ ;
	wire _w3213_ ;
	wire _w3212_ ;
	wire _w3211_ ;
	wire _w3210_ ;
	wire _w3209_ ;
	wire _w3208_ ;
	wire _w3207_ ;
	wire _w3206_ ;
	wire _w3205_ ;
	wire _w3204_ ;
	wire _w3203_ ;
	wire _w3202_ ;
	wire _w3201_ ;
	wire _w3200_ ;
	wire _w3199_ ;
	wire _w3198_ ;
	wire _w3197_ ;
	wire _w3196_ ;
	wire _w3195_ ;
	wire _w3194_ ;
	wire _w3193_ ;
	wire _w3192_ ;
	wire _w3191_ ;
	wire _w3190_ ;
	wire _w3189_ ;
	wire _w3188_ ;
	wire _w3187_ ;
	wire _w3186_ ;
	wire _w3185_ ;
	wire _w3184_ ;
	wire _w3183_ ;
	wire _w3182_ ;
	wire _w3181_ ;
	wire _w3180_ ;
	wire _w3179_ ;
	wire _w3178_ ;
	wire _w3177_ ;
	wire _w3176_ ;
	wire _w3175_ ;
	wire _w3174_ ;
	wire _w3173_ ;
	wire _w3172_ ;
	wire _w3171_ ;
	wire _w3170_ ;
	wire _w3169_ ;
	wire _w3168_ ;
	wire _w3167_ ;
	wire _w3166_ ;
	wire _w3165_ ;
	wire _w3164_ ;
	wire _w3163_ ;
	wire _w3162_ ;
	wire _w3161_ ;
	wire _w3160_ ;
	wire _w3159_ ;
	wire _w3158_ ;
	wire _w3157_ ;
	wire _w3156_ ;
	wire _w3155_ ;
	wire _w3154_ ;
	wire _w3153_ ;
	wire _w3152_ ;
	wire _w3151_ ;
	wire _w3150_ ;
	wire _w3149_ ;
	wire _w3148_ ;
	wire _w3147_ ;
	wire _w3146_ ;
	wire _w3145_ ;
	wire _w3144_ ;
	wire _w3143_ ;
	wire _w3142_ ;
	wire _w3141_ ;
	wire _w3140_ ;
	wire _w3139_ ;
	wire _w3138_ ;
	wire _w3137_ ;
	wire _w3136_ ;
	wire _w3135_ ;
	wire _w3134_ ;
	wire _w3133_ ;
	wire _w3132_ ;
	wire _w3131_ ;
	wire _w1882_ ;
	wire _w1881_ ;
	wire _w1880_ ;
	wire _w1879_ ;
	wire _w1878_ ;
	wire _w1877_ ;
	wire _w1876_ ;
	wire _w1875_ ;
	wire _w1874_ ;
	wire _w1873_ ;
	wire _w1872_ ;
	wire _w1871_ ;
	wire _w1870_ ;
	wire _w1869_ ;
	wire _w1868_ ;
	wire _w1867_ ;
	wire _w1866_ ;
	wire _w1865_ ;
	wire _w1864_ ;
	wire _w1863_ ;
	wire _w1862_ ;
	wire _w1861_ ;
	wire _w1860_ ;
	wire _w1859_ ;
	wire _w1858_ ;
	wire _w1857_ ;
	wire _w1856_ ;
	wire _w1855_ ;
	wire _w1854_ ;
	wire _w1853_ ;
	wire _w1852_ ;
	wire _w1851_ ;
	wire _w1850_ ;
	wire _w1849_ ;
	wire _w1848_ ;
	wire _w1847_ ;
	wire _w1846_ ;
	wire _w1845_ ;
	wire _w1844_ ;
	wire _w1843_ ;
	wire _w1842_ ;
	wire _w1841_ ;
	wire _w1840_ ;
	wire _w1839_ ;
	wire _w1838_ ;
	wire _w1837_ ;
	wire _w1836_ ;
	wire _w1835_ ;
	wire _w1834_ ;
	wire _w1833_ ;
	wire _w1832_ ;
	wire _w1831_ ;
	wire _w1830_ ;
	wire _w1829_ ;
	wire _w1828_ ;
	wire _w1827_ ;
	wire _w1826_ ;
	wire _w1825_ ;
	wire _w1824_ ;
	wire _w1823_ ;
	wire _w1822_ ;
	wire _w1821_ ;
	wire _w1820_ ;
	wire _w1819_ ;
	wire _w1818_ ;
	wire _w1817_ ;
	wire _w1816_ ;
	wire _w1815_ ;
	wire _w1814_ ;
	wire _w1813_ ;
	wire _w1812_ ;
	wire _w1811_ ;
	wire _w1810_ ;
	wire _w1809_ ;
	wire _w1808_ ;
	wire _w1807_ ;
	wire _w1806_ ;
	wire _w1805_ ;
	wire _w1804_ ;
	wire _w1803_ ;
	wire _w1802_ ;
	wire _w1801_ ;
	wire _w1800_ ;
	wire _w1799_ ;
	wire _w1798_ ;
	wire _w1797_ ;
	wire _w1796_ ;
	wire _w1795_ ;
	wire _w1794_ ;
	wire _w1793_ ;
	wire _w1792_ ;
	wire _w1791_ ;
	wire _w1790_ ;
	wire _w1789_ ;
	wire _w1788_ ;
	wire _w1787_ ;
	wire _w1786_ ;
	wire _w1785_ ;
	wire _w1784_ ;
	wire _w1783_ ;
	wire _w1782_ ;
	wire _w1781_ ;
	wire _w1780_ ;
	wire _w1779_ ;
	wire _w1778_ ;
	wire _w1777_ ;
	wire _w1776_ ;
	wire _w1775_ ;
	wire _w1774_ ;
	wire _w1773_ ;
	wire _w1772_ ;
	wire _w1771_ ;
	wire _w1770_ ;
	wire _w1769_ ;
	wire _w1768_ ;
	wire _w1767_ ;
	wire _w1766_ ;
	wire _w1765_ ;
	wire _w1764_ ;
	wire _w1763_ ;
	wire _w1762_ ;
	wire _w1761_ ;
	wire _w1760_ ;
	wire _w1759_ ;
	wire _w1758_ ;
	wire _w1757_ ;
	wire _w1756_ ;
	wire _w1755_ ;
	wire _w1754_ ;
	wire _w1753_ ;
	wire _w1752_ ;
	wire _w1751_ ;
	wire _w1750_ ;
	wire _w1749_ ;
	wire _w1748_ ;
	wire _w1747_ ;
	wire _w1746_ ;
	wire _w1745_ ;
	wire _w1744_ ;
	wire _w1743_ ;
	wire _w1742_ ;
	wire _w1741_ ;
	wire _w1740_ ;
	wire _w1739_ ;
	wire _w1738_ ;
	wire _w1737_ ;
	wire _w1736_ ;
	wire _w1735_ ;
	wire _w1734_ ;
	wire _w1733_ ;
	wire _w1732_ ;
	wire _w1731_ ;
	wire _w1730_ ;
	wire _w1729_ ;
	wire _w1728_ ;
	wire _w1727_ ;
	wire _w1726_ ;
	wire _w1725_ ;
	wire _w1724_ ;
	wire _w1723_ ;
	wire _w1722_ ;
	wire _w1721_ ;
	wire _w1720_ ;
	wire _w1719_ ;
	wire _w1718_ ;
	wire _w1717_ ;
	wire _w1716_ ;
	wire _w1715_ ;
	wire _w1714_ ;
	wire _w1713_ ;
	wire _w1712_ ;
	wire _w1711_ ;
	wire _w1710_ ;
	wire _w1709_ ;
	wire _w1708_ ;
	wire _w1707_ ;
	wire _w1706_ ;
	wire _w1705_ ;
	wire _w1704_ ;
	wire _w1703_ ;
	wire _w1702_ ;
	wire _w1701_ ;
	wire _w1700_ ;
	wire _w1699_ ;
	wire _w1698_ ;
	wire _w1697_ ;
	wire _w1696_ ;
	wire _w1695_ ;
	wire _w1694_ ;
	wire _w1693_ ;
	wire _w1692_ ;
	wire _w1691_ ;
	wire _w1690_ ;
	wire _w1689_ ;
	wire _w1688_ ;
	wire _w1687_ ;
	wire _w1686_ ;
	wire _w1685_ ;
	wire _w1684_ ;
	wire _w1683_ ;
	wire _w1682_ ;
	wire _w1681_ ;
	wire _w1680_ ;
	wire _w1679_ ;
	wire _w1678_ ;
	wire _w1677_ ;
	wire _w1676_ ;
	wire _w1675_ ;
	wire _w1674_ ;
	wire _w1673_ ;
	wire _w1672_ ;
	wire _w1671_ ;
	wire _w1670_ ;
	wire _w1669_ ;
	wire _w1668_ ;
	wire _w1667_ ;
	wire _w1666_ ;
	wire _w1665_ ;
	wire _w1664_ ;
	wire _w1663_ ;
	wire _w1662_ ;
	wire _w1661_ ;
	wire _w1660_ ;
	wire _w1659_ ;
	wire _w1658_ ;
	wire _w1657_ ;
	wire _w1656_ ;
	wire _w1655_ ;
	wire _w1654_ ;
	wire _w1653_ ;
	wire _w1652_ ;
	wire _w1651_ ;
	wire _w1650_ ;
	wire _w1649_ ;
	wire _w1648_ ;
	wire _w1647_ ;
	wire _w1646_ ;
	wire _w1645_ ;
	wire _w1644_ ;
	wire _w1643_ ;
	wire _w1642_ ;
	wire _w1641_ ;
	wire _w1640_ ;
	wire _w1639_ ;
	wire _w1638_ ;
	wire _w1637_ ;
	wire _w1636_ ;
	wire _w1635_ ;
	wire _w1634_ ;
	wire _w1633_ ;
	wire _w1632_ ;
	wire _w1631_ ;
	wire _w1630_ ;
	wire _w1629_ ;
	wire _w1628_ ;
	wire _w1627_ ;
	wire _w1626_ ;
	wire _w1625_ ;
	wire _w1624_ ;
	wire _w1623_ ;
	wire _w1622_ ;
	wire _w1621_ ;
	wire _w1620_ ;
	wire _w1619_ ;
	wire _w1618_ ;
	wire _w1617_ ;
	wire _w1616_ ;
	wire _w1615_ ;
	wire _w1614_ ;
	wire _w1613_ ;
	wire _w1612_ ;
	wire _w1611_ ;
	wire _w1610_ ;
	wire _w1609_ ;
	wire _w1608_ ;
	wire _w1607_ ;
	wire _w1606_ ;
	wire _w1605_ ;
	wire _w1604_ ;
	wire _w1603_ ;
	wire _w1602_ ;
	wire _w1601_ ;
	wire _w1600_ ;
	wire _w1599_ ;
	wire _w1598_ ;
	wire _w1597_ ;
	wire _w1596_ ;
	wire _w1595_ ;
	wire _w1594_ ;
	wire _w1593_ ;
	wire _w1592_ ;
	wire _w1591_ ;
	wire _w1590_ ;
	wire _w1589_ ;
	wire _w1588_ ;
	wire _w1587_ ;
	wire _w1586_ ;
	wire _w1585_ ;
	wire _w1584_ ;
	wire _w1583_ ;
	wire _w1582_ ;
	wire _w1581_ ;
	wire _w1580_ ;
	wire _w1579_ ;
	wire _w1578_ ;
	wire _w1577_ ;
	wire _w1576_ ;
	wire _w1575_ ;
	wire _w1574_ ;
	wire _w1573_ ;
	wire _w1572_ ;
	wire _w1571_ ;
	wire _w1570_ ;
	wire _w1569_ ;
	wire _w1568_ ;
	wire _w1567_ ;
	wire _w1566_ ;
	wire _w1565_ ;
	wire _w1564_ ;
	wire _w1563_ ;
	wire _w1562_ ;
	wire _w1561_ ;
	wire _w1560_ ;
	wire _w1559_ ;
	wire _w1558_ ;
	wire _w1557_ ;
	wire _w1556_ ;
	wire _w1555_ ;
	wire _w1554_ ;
	wire _w1553_ ;
	wire _w1552_ ;
	wire _w1551_ ;
	wire _w1550_ ;
	wire _w1549_ ;
	wire _w1548_ ;
	wire _w1547_ ;
	wire _w1546_ ;
	wire _w1545_ ;
	wire _w1544_ ;
	wire _w1543_ ;
	wire _w1542_ ;
	wire _w1541_ ;
	wire _w1540_ ;
	wire _w1539_ ;
	wire _w1538_ ;
	wire _w1537_ ;
	wire _w1536_ ;
	wire _w1535_ ;
	wire _w1534_ ;
	wire _w1533_ ;
	wire _w1532_ ;
	wire _w1531_ ;
	wire _w1530_ ;
	wire _w1529_ ;
	wire _w1528_ ;
	wire _w1527_ ;
	wire _w1526_ ;
	wire _w1525_ ;
	wire _w1524_ ;
	wire _w1523_ ;
	wire _w1522_ ;
	wire _w1521_ ;
	wire _w1520_ ;
	wire _w1519_ ;
	wire _w1518_ ;
	wire _w1517_ ;
	wire _w1516_ ;
	wire _w1515_ ;
	wire _w1514_ ;
	wire _w1513_ ;
	wire _w1512_ ;
	wire _w1511_ ;
	wire _w1510_ ;
	wire _w1509_ ;
	wire _w1508_ ;
	wire _w1507_ ;
	wire _w1506_ ;
	wire _w1505_ ;
	wire _w1504_ ;
	wire _w1503_ ;
	wire _w1502_ ;
	wire _w1501_ ;
	wire _w1500_ ;
	wire _w1499_ ;
	wire _w1498_ ;
	wire _w1497_ ;
	wire _w1496_ ;
	wire _w1495_ ;
	wire _w1494_ ;
	wire _w1493_ ;
	wire _w1492_ ;
	wire _w1491_ ;
	wire _w1490_ ;
	wire _w1489_ ;
	wire _w1488_ ;
	wire _w1487_ ;
	wire _w1486_ ;
	wire _w1485_ ;
	wire _w1484_ ;
	wire _w1483_ ;
	wire _w1482_ ;
	wire _w1481_ ;
	wire _w1480_ ;
	wire _w1479_ ;
	wire _w1478_ ;
	wire _w1477_ ;
	wire _w1476_ ;
	wire _w1475_ ;
	wire _w1474_ ;
	wire _w1473_ ;
	wire _w1472_ ;
	wire _w1471_ ;
	wire _w1470_ ;
	wire _w1469_ ;
	wire _w1468_ ;
	wire _w1467_ ;
	wire _w1466_ ;
	wire _w1465_ ;
	wire _w1464_ ;
	wire _w1463_ ;
	wire _w1462_ ;
	wire _w1461_ ;
	wire _w1460_ ;
	wire _w1459_ ;
	wire _w1458_ ;
	wire _w1457_ ;
	wire _w1456_ ;
	wire _w1455_ ;
	wire _w1454_ ;
	wire _w1453_ ;
	wire _w1452_ ;
	wire _w1451_ ;
	wire _w1450_ ;
	wire _w1449_ ;
	wire _w1448_ ;
	wire _w1447_ ;
	wire _w1446_ ;
	wire _w1445_ ;
	wire _w1444_ ;
	wire _w1443_ ;
	wire _w1442_ ;
	wire _w1441_ ;
	wire _w1440_ ;
	wire _w1439_ ;
	wire _w1438_ ;
	wire _w1437_ ;
	wire _w1436_ ;
	wire _w1435_ ;
	wire _w1434_ ;
	wire _w1433_ ;
	wire _w1432_ ;
	wire _w1431_ ;
	wire _w1430_ ;
	wire _w1429_ ;
	wire _w1428_ ;
	wire _w1427_ ;
	wire _w1426_ ;
	wire _w1425_ ;
	wire _w1424_ ;
	wire _w1423_ ;
	wire _w1422_ ;
	wire _w1421_ ;
	wire _w1420_ ;
	wire _w1419_ ;
	wire _w1418_ ;
	wire _w1417_ ;
	wire _w1416_ ;
	wire _w1415_ ;
	wire _w1414_ ;
	wire _w1413_ ;
	wire _w1412_ ;
	wire _w1411_ ;
	wire _w1410_ ;
	wire _w1409_ ;
	wire _w1408_ ;
	wire _w1407_ ;
	wire _w1406_ ;
	wire _w1405_ ;
	wire _w1404_ ;
	wire _w1403_ ;
	wire _w1402_ ;
	wire _w1401_ ;
	wire _w1400_ ;
	wire _w1399_ ;
	wire _w1398_ ;
	wire _w1397_ ;
	wire _w1396_ ;
	wire _w1395_ ;
	wire _w1394_ ;
	wire _w1393_ ;
	wire _w1392_ ;
	wire _w1391_ ;
	wire _w1390_ ;
	wire _w1389_ ;
	wire _w1388_ ;
	wire _w1387_ ;
	wire _w1386_ ;
	wire _w1385_ ;
	wire _w1384_ ;
	wire _w1383_ ;
	wire _w1382_ ;
	wire _w1381_ ;
	wire _w1380_ ;
	wire _w1379_ ;
	wire _w1378_ ;
	wire _w1377_ ;
	wire _w1376_ ;
	wire _w1375_ ;
	wire _w1374_ ;
	wire _w1373_ ;
	wire _w1372_ ;
	wire _w1371_ ;
	wire _w1370_ ;
	wire _w1369_ ;
	wire _w1368_ ;
	wire _w1367_ ;
	wire _w1366_ ;
	wire _w1365_ ;
	wire _w1364_ ;
	wire _w1363_ ;
	wire _w1362_ ;
	wire _w1361_ ;
	wire _w1360_ ;
	wire _w1359_ ;
	wire _w1358_ ;
	wire _w1357_ ;
	wire _w1356_ ;
	wire _w1355_ ;
	wire _w1354_ ;
	wire _w1353_ ;
	wire _w1352_ ;
	wire _w1351_ ;
	wire _w1350_ ;
	wire _w1349_ ;
	wire _w1348_ ;
	wire _w1347_ ;
	wire _w1346_ ;
	wire _w1345_ ;
	wire _w1344_ ;
	wire _w1343_ ;
	wire _w1342_ ;
	wire _w1341_ ;
	wire _w1340_ ;
	wire _w1339_ ;
	wire _w1338_ ;
	wire _w1337_ ;
	wire _w1336_ ;
	wire _w1335_ ;
	wire _w1334_ ;
	wire _w1333_ ;
	wire _w1332_ ;
	wire _w1331_ ;
	wire _w1330_ ;
	wire _w1329_ ;
	wire _w1328_ ;
	wire _w1327_ ;
	wire _w1326_ ;
	wire _w1325_ ;
	wire _w1324_ ;
	wire _w1323_ ;
	wire _w1322_ ;
	wire _w1321_ ;
	wire _w1320_ ;
	wire _w1319_ ;
	wire _w1318_ ;
	wire _w1317_ ;
	wire _w1316_ ;
	wire _w1315_ ;
	wire _w1030_ ;
	wire _w1029_ ;
	wire _w1028_ ;
	wire _w1027_ ;
	wire _w1026_ ;
	wire _w1025_ ;
	wire _w1024_ ;
	wire _w1023_ ;
	wire _w1022_ ;
	wire _w1021_ ;
	wire _w1020_ ;
	wire _w1019_ ;
	wire _w1018_ ;
	wire _w1017_ ;
	wire _w1016_ ;
	wire _w1015_ ;
	wire _w1014_ ;
	wire _w1013_ ;
	wire _w1012_ ;
	wire _w1011_ ;
	wire _w1010_ ;
	wire _w1009_ ;
	wire _w1008_ ;
	wire _w1007_ ;
	wire _w1006_ ;
	wire _w1005_ ;
	wire _w1004_ ;
	wire _w1003_ ;
	wire _w1002_ ;
	wire _w1001_ ;
	wire _w1000_ ;
	wire _w999_ ;
	wire _w998_ ;
	wire _w997_ ;
	wire _w996_ ;
	wire _w995_ ;
	wire _w994_ ;
	wire _w993_ ;
	wire _w992_ ;
	wire _w991_ ;
	wire _w990_ ;
	wire _w989_ ;
	wire _w988_ ;
	wire _w987_ ;
	wire _w986_ ;
	wire _w985_ ;
	wire _w984_ ;
	wire _w983_ ;
	wire _w982_ ;
	wire _w981_ ;
	wire _w980_ ;
	wire _w979_ ;
	wire _w978_ ;
	wire _w977_ ;
	wire _w976_ ;
	wire _w975_ ;
	wire _w974_ ;
	wire _w973_ ;
	wire _w972_ ;
	wire _w971_ ;
	wire _w970_ ;
	wire _w969_ ;
	wire _w968_ ;
	wire _w967_ ;
	wire _w966_ ;
	wire _w965_ ;
	wire _w964_ ;
	wire _w963_ ;
	wire _w962_ ;
	wire _w961_ ;
	wire _w960_ ;
	wire _w959_ ;
	wire _w958_ ;
	wire _w957_ ;
	wire _w956_ ;
	wire _w955_ ;
	wire _w954_ ;
	wire _w953_ ;
	wire _w952_ ;
	wire _w951_ ;
	wire _w950_ ;
	wire _w949_ ;
	wire _w948_ ;
	wire _w947_ ;
	wire _w946_ ;
	wire _w945_ ;
	wire _w944_ ;
	wire _w943_ ;
	wire _w942_ ;
	wire _w941_ ;
	wire _w940_ ;
	wire _w939_ ;
	wire _w938_ ;
	wire _w937_ ;
	wire _w936_ ;
	wire _w935_ ;
	wire _w934_ ;
	wire _w933_ ;
	wire _w932_ ;
	wire _w931_ ;
	wire _w930_ ;
	wire _w929_ ;
	wire _w928_ ;
	wire _w927_ ;
	wire _w926_ ;
	wire _w925_ ;
	wire _w924_ ;
	wire _w923_ ;
	wire _w922_ ;
	wire _w921_ ;
	wire _w920_ ;
	wire _w919_ ;
	wire _w918_ ;
	wire _w917_ ;
	wire _w916_ ;
	wire _w915_ ;
	wire _w914_ ;
	wire _w913_ ;
	wire _w912_ ;
	wire _w911_ ;
	wire _w910_ ;
	wire _w909_ ;
	wire _w908_ ;
	wire _w907_ ;
	wire _w906_ ;
	wire _w905_ ;
	wire _w904_ ;
	wire _w903_ ;
	wire _w902_ ;
	wire _w901_ ;
	wire _w832_ ;
	wire _w831_ ;
	wire _w830_ ;
	wire _w829_ ;
	wire _w828_ ;
	wire _w827_ ;
	wire _w826_ ;
	wire _w825_ ;
	wire _w824_ ;
	wire _w823_ ;
	wire _w822_ ;
	wire _w821_ ;
	wire _w820_ ;
	wire _w819_ ;
	wire _w818_ ;
	wire _w817_ ;
	wire _w816_ ;
	wire _w815_ ;
	wire _w814_ ;
	wire _w813_ ;
	wire _w812_ ;
	wire _w811_ ;
	wire _w810_ ;
	wire _w809_ ;
	wire _w808_ ;
	wire _w807_ ;
	wire _w806_ ;
	wire _w805_ ;
	wire _w804_ ;
	wire _w803_ ;
	wire _w786_ ;
	wire _w785_ ;
	wire _w784_ ;
	wire _w783_ ;
	wire _w782_ ;
	wire _w781_ ;
	wire _w780_ ;
	wire _w779_ ;
	wire _w778_ ;
	wire _w777_ ;
	wire _w776_ ;
	wire _w775_ ;
	wire _w774_ ;
	wire _w787_ ;
	wire _w788_ ;
	wire _w789_ ;
	wire _w790_ ;
	wire _w791_ ;
	wire _w792_ ;
	wire _w793_ ;
	wire _w794_ ;
	wire _w795_ ;
	wire _w796_ ;
	wire _w797_ ;
	wire _w798_ ;
	wire _w799_ ;
	wire _w800_ ;
	wire _w801_ ;
	wire _w802_ ;
	wire _w833_ ;
	wire _w834_ ;
	wire _w835_ ;
	wire _w836_ ;
	wire _w837_ ;
	wire _w838_ ;
	wire _w839_ ;
	wire _w840_ ;
	wire _w841_ ;
	wire _w842_ ;
	wire _w843_ ;
	wire _w844_ ;
	wire _w845_ ;
	wire _w846_ ;
	wire _w847_ ;
	wire _w848_ ;
	wire _w849_ ;
	wire _w850_ ;
	wire _w851_ ;
	wire _w852_ ;
	wire _w853_ ;
	wire _w854_ ;
	wire _w855_ ;
	wire _w856_ ;
	wire _w857_ ;
	wire _w858_ ;
	wire _w859_ ;
	wire _w860_ ;
	wire _w861_ ;
	wire _w862_ ;
	wire _w863_ ;
	wire _w864_ ;
	wire _w865_ ;
	wire _w866_ ;
	wire _w867_ ;
	wire _w868_ ;
	wire _w869_ ;
	wire _w870_ ;
	wire _w871_ ;
	wire _w872_ ;
	wire _w873_ ;
	wire _w874_ ;
	wire _w875_ ;
	wire _w876_ ;
	wire _w877_ ;
	wire _w878_ ;
	wire _w879_ ;
	wire _w880_ ;
	wire _w881_ ;
	wire _w882_ ;
	wire _w883_ ;
	wire _w884_ ;
	wire _w885_ ;
	wire _w886_ ;
	wire _w887_ ;
	wire _w888_ ;
	wire _w889_ ;
	wire _w890_ ;
	wire _w891_ ;
	wire _w892_ ;
	wire _w893_ ;
	wire _w894_ ;
	wire _w895_ ;
	wire _w896_ ;
	wire _w897_ ;
	wire _w898_ ;
	wire _w899_ ;
	wire _w900_ ;
	wire _w1031_ ;
	wire _w1032_ ;
	wire _w1033_ ;
	wire _w1034_ ;
	wire _w1035_ ;
	wire _w1036_ ;
	wire _w1037_ ;
	wire _w1038_ ;
	wire _w1039_ ;
	wire _w1040_ ;
	wire _w1041_ ;
	wire _w1042_ ;
	wire _w1043_ ;
	wire _w1044_ ;
	wire _w1045_ ;
	wire _w1046_ ;
	wire _w1047_ ;
	wire _w1048_ ;
	wire _w1049_ ;
	wire _w1050_ ;
	wire _w1051_ ;
	wire _w1052_ ;
	wire _w1053_ ;
	wire _w1054_ ;
	wire _w1055_ ;
	wire _w1056_ ;
	wire _w1057_ ;
	wire _w1058_ ;
	wire _w1059_ ;
	wire _w1060_ ;
	wire _w1061_ ;
	wire _w1062_ ;
	wire _w1063_ ;
	wire _w1064_ ;
	wire _w1065_ ;
	wire _w1066_ ;
	wire _w1067_ ;
	wire _w1068_ ;
	wire _w1069_ ;
	wire _w1070_ ;
	wire _w1071_ ;
	wire _w1072_ ;
	wire _w1073_ ;
	wire _w1074_ ;
	wire _w1075_ ;
	wire _w1076_ ;
	wire _w1077_ ;
	wire _w1078_ ;
	wire _w1079_ ;
	wire _w1080_ ;
	wire _w1081_ ;
	wire _w1082_ ;
	wire _w1083_ ;
	wire _w1084_ ;
	wire _w1085_ ;
	wire _w1086_ ;
	wire _w1087_ ;
	wire _w1088_ ;
	wire _w1089_ ;
	wire _w1090_ ;
	wire _w1091_ ;
	wire _w1092_ ;
	wire _w1093_ ;
	wire _w1094_ ;
	wire _w1095_ ;
	wire _w1096_ ;
	wire _w1097_ ;
	wire _w1098_ ;
	wire _w1099_ ;
	wire _w1100_ ;
	wire _w1101_ ;
	wire _w1102_ ;
	wire _w1103_ ;
	wire _w1104_ ;
	wire _w1105_ ;
	wire _w1106_ ;
	wire _w1107_ ;
	wire _w1108_ ;
	wire _w1109_ ;
	wire _w1110_ ;
	wire _w1111_ ;
	wire _w1112_ ;
	wire _w1113_ ;
	wire _w1114_ ;
	wire _w1115_ ;
	wire _w1116_ ;
	wire _w1117_ ;
	wire _w1118_ ;
	wire _w1119_ ;
	wire _w1120_ ;
	wire _w1121_ ;
	wire _w1122_ ;
	wire _w1123_ ;
	wire _w1124_ ;
	wire _w1125_ ;
	wire _w1126_ ;
	wire _w1127_ ;
	wire _w1128_ ;
	wire _w1129_ ;
	wire _w1130_ ;
	wire _w1131_ ;
	wire _w1132_ ;
	wire _w1133_ ;
	wire _w1134_ ;
	wire _w1135_ ;
	wire _w1136_ ;
	wire _w1137_ ;
	wire _w1138_ ;
	wire _w1139_ ;
	wire _w1140_ ;
	wire _w1141_ ;
	wire _w1142_ ;
	wire _w1143_ ;
	wire _w1144_ ;
	wire _w1145_ ;
	wire _w1146_ ;
	wire _w1147_ ;
	wire _w1148_ ;
	wire _w1149_ ;
	wire _w1150_ ;
	wire _w1151_ ;
	wire _w1152_ ;
	wire _w1153_ ;
	wire _w1154_ ;
	wire _w1155_ ;
	wire _w1156_ ;
	wire _w1157_ ;
	wire _w1158_ ;
	wire _w1159_ ;
	wire _w1160_ ;
	wire _w1161_ ;
	wire _w1162_ ;
	wire _w1163_ ;
	wire _w1164_ ;
	wire _w1165_ ;
	wire _w1166_ ;
	wire _w1167_ ;
	wire _w1168_ ;
	wire _w1169_ ;
	wire _w1170_ ;
	wire _w1171_ ;
	wire _w1172_ ;
	wire _w1173_ ;
	wire _w1174_ ;
	wire _w1175_ ;
	wire _w1176_ ;
	wire _w1177_ ;
	wire _w1178_ ;
	wire _w1179_ ;
	wire _w1180_ ;
	wire _w1181_ ;
	wire _w1182_ ;
	wire _w1183_ ;
	wire _w1184_ ;
	wire _w1185_ ;
	wire _w1186_ ;
	wire _w1187_ ;
	wire _w1188_ ;
	wire _w1189_ ;
	wire _w1190_ ;
	wire _w1191_ ;
	wire _w1192_ ;
	wire _w1193_ ;
	wire _w1194_ ;
	wire _w1195_ ;
	wire _w1196_ ;
	wire _w1197_ ;
	wire _w1198_ ;
	wire _w1199_ ;
	wire _w1200_ ;
	wire _w1201_ ;
	wire _w1202_ ;
	wire _w1203_ ;
	wire _w1204_ ;
	wire _w1205_ ;
	wire _w1206_ ;
	wire _w1207_ ;
	wire _w1208_ ;
	wire _w1209_ ;
	wire _w1210_ ;
	wire _w1211_ ;
	wire _w1212_ ;
	wire _w1213_ ;
	wire _w1214_ ;
	wire _w1215_ ;
	wire _w1216_ ;
	wire _w1217_ ;
	wire _w1218_ ;
	wire _w1219_ ;
	wire _w1220_ ;
	wire _w1221_ ;
	wire _w1222_ ;
	wire _w1223_ ;
	wire _w1224_ ;
	wire _w1225_ ;
	wire _w1226_ ;
	wire _w1227_ ;
	wire _w1228_ ;
	wire _w1229_ ;
	wire _w1230_ ;
	wire _w1231_ ;
	wire _w1232_ ;
	wire _w1233_ ;
	wire _w1234_ ;
	wire _w1235_ ;
	wire _w1236_ ;
	wire _w1237_ ;
	wire _w1238_ ;
	wire _w1239_ ;
	wire _w1240_ ;
	wire _w1241_ ;
	wire _w1242_ ;
	wire _w1243_ ;
	wire _w1244_ ;
	wire _w1245_ ;
	wire _w1246_ ;
	wire _w1247_ ;
	wire _w1248_ ;
	wire _w1249_ ;
	wire _w1250_ ;
	wire _w1251_ ;
	wire _w1252_ ;
	wire _w1253_ ;
	wire _w1254_ ;
	wire _w1255_ ;
	wire _w1256_ ;
	wire _w1257_ ;
	wire _w1258_ ;
	wire _w1259_ ;
	wire _w1260_ ;
	wire _w1261_ ;
	wire _w1262_ ;
	wire _w1263_ ;
	wire _w1264_ ;
	wire _w1265_ ;
	wire _w1266_ ;
	wire _w1267_ ;
	wire _w1268_ ;
	wire _w1269_ ;
	wire _w1270_ ;
	wire _w1271_ ;
	wire _w1272_ ;
	wire _w1273_ ;
	wire _w1274_ ;
	wire _w1275_ ;
	wire _w1276_ ;
	wire _w1277_ ;
	wire _w1278_ ;
	wire _w1279_ ;
	wire _w1280_ ;
	wire _w1281_ ;
	wire _w1282_ ;
	wire _w1283_ ;
	wire _w1284_ ;
	wire _w1285_ ;
	wire _w1286_ ;
	wire _w1287_ ;
	wire _w1288_ ;
	wire _w1289_ ;
	wire _w1290_ ;
	wire _w1291_ ;
	wire _w1292_ ;
	wire _w1293_ ;
	wire _w1294_ ;
	wire _w1295_ ;
	wire _w1296_ ;
	wire _w1297_ ;
	wire _w1298_ ;
	wire _w1299_ ;
	wire _w1300_ ;
	wire _w1301_ ;
	wire _w1302_ ;
	wire _w1303_ ;
	wire _w1304_ ;
	wire _w1305_ ;
	wire _w1306_ ;
	wire _w1307_ ;
	wire _w1308_ ;
	wire _w1309_ ;
	wire _w1310_ ;
	wire _w1311_ ;
	wire _w1312_ ;
	wire _w1313_ ;
	wire _w1314_ ;
	wire _w1883_ ;
	wire _w1884_ ;
	wire _w1885_ ;
	wire _w1886_ ;
	wire _w1887_ ;
	wire _w1888_ ;
	wire _w1889_ ;
	wire _w1890_ ;
	wire _w1891_ ;
	wire _w1892_ ;
	wire _w1893_ ;
	wire _w1894_ ;
	wire _w1895_ ;
	wire _w1896_ ;
	wire _w1897_ ;
	wire _w1898_ ;
	wire _w1899_ ;
	wire _w1900_ ;
	wire _w1901_ ;
	wire _w1902_ ;
	wire _w1903_ ;
	wire _w1904_ ;
	wire _w1905_ ;
	wire _w1906_ ;
	wire _w1907_ ;
	wire _w1908_ ;
	wire _w1909_ ;
	wire _w1910_ ;
	wire _w1911_ ;
	wire _w1912_ ;
	wire _w1913_ ;
	wire _w1914_ ;
	wire _w1915_ ;
	wire _w1916_ ;
	wire _w1917_ ;
	wire _w1918_ ;
	wire _w1919_ ;
	wire _w1920_ ;
	wire _w1921_ ;
	wire _w1922_ ;
	wire _w1923_ ;
	wire _w1924_ ;
	wire _w1925_ ;
	wire _w1926_ ;
	wire _w1927_ ;
	wire _w1928_ ;
	wire _w1929_ ;
	wire _w1930_ ;
	wire _w1931_ ;
	wire _w1932_ ;
	wire _w1933_ ;
	wire _w1934_ ;
	wire _w1935_ ;
	wire _w1936_ ;
	wire _w1937_ ;
	wire _w1938_ ;
	wire _w1939_ ;
	wire _w1940_ ;
	wire _w1941_ ;
	wire _w1942_ ;
	wire _w1943_ ;
	wire _w1944_ ;
	wire _w1945_ ;
	wire _w1946_ ;
	wire _w1947_ ;
	wire _w1948_ ;
	wire _w1949_ ;
	wire _w1950_ ;
	wire _w1951_ ;
	wire _w1952_ ;
	wire _w1953_ ;
	wire _w1954_ ;
	wire _w1955_ ;
	wire _w1956_ ;
	wire _w1957_ ;
	wire _w1958_ ;
	wire _w1959_ ;
	wire _w1960_ ;
	wire _w1961_ ;
	wire _w1962_ ;
	wire _w1963_ ;
	wire _w1964_ ;
	wire _w1965_ ;
	wire _w1966_ ;
	wire _w1967_ ;
	wire _w1968_ ;
	wire _w1969_ ;
	wire _w1970_ ;
	wire _w1971_ ;
	wire _w1972_ ;
	wire _w1973_ ;
	wire _w1974_ ;
	wire _w1975_ ;
	wire _w1976_ ;
	wire _w1977_ ;
	wire _w1978_ ;
	wire _w1979_ ;
	wire _w1980_ ;
	wire _w1981_ ;
	wire _w1982_ ;
	wire _w1983_ ;
	wire _w1984_ ;
	wire _w1985_ ;
	wire _w1986_ ;
	wire _w1987_ ;
	wire _w1988_ ;
	wire _w1989_ ;
	wire _w1990_ ;
	wire _w1991_ ;
	wire _w1992_ ;
	wire _w1993_ ;
	wire _w1994_ ;
	wire _w1995_ ;
	wire _w1996_ ;
	wire _w1997_ ;
	wire _w1998_ ;
	wire _w1999_ ;
	wire _w2000_ ;
	wire _w2001_ ;
	wire _w2002_ ;
	wire _w2003_ ;
	wire _w2004_ ;
	wire _w2005_ ;
	wire _w2006_ ;
	wire _w2007_ ;
	wire _w2008_ ;
	wire _w2009_ ;
	wire _w2010_ ;
	wire _w2011_ ;
	wire _w2012_ ;
	wire _w2013_ ;
	wire _w2014_ ;
	wire _w2015_ ;
	wire _w2016_ ;
	wire _w2017_ ;
	wire _w2018_ ;
	wire _w2019_ ;
	wire _w2020_ ;
	wire _w2021_ ;
	wire _w2022_ ;
	wire _w2023_ ;
	wire _w2024_ ;
	wire _w2025_ ;
	wire _w2026_ ;
	wire _w2027_ ;
	wire _w2028_ ;
	wire _w2029_ ;
	wire _w2030_ ;
	wire _w2031_ ;
	wire _w2032_ ;
	wire _w2033_ ;
	wire _w2034_ ;
	wire _w2035_ ;
	wire _w2036_ ;
	wire _w2037_ ;
	wire _w2038_ ;
	wire _w2039_ ;
	wire _w2040_ ;
	wire _w2041_ ;
	wire _w2042_ ;
	wire _w2043_ ;
	wire _w2044_ ;
	wire _w2045_ ;
	wire _w2046_ ;
	wire _w2047_ ;
	wire _w2048_ ;
	wire _w2049_ ;
	wire _w2050_ ;
	wire _w2051_ ;
	wire _w2052_ ;
	wire _w2053_ ;
	wire _w2054_ ;
	wire _w2055_ ;
	wire _w2056_ ;
	wire _w2057_ ;
	wire _w2058_ ;
	wire _w2059_ ;
	wire _w2060_ ;
	wire _w2061_ ;
	wire _w2062_ ;
	wire _w2063_ ;
	wire _w2064_ ;
	wire _w2065_ ;
	wire _w2066_ ;
	wire _w2067_ ;
	wire _w2068_ ;
	wire _w2069_ ;
	wire _w2070_ ;
	wire _w2071_ ;
	wire _w2072_ ;
	wire _w2073_ ;
	wire _w2074_ ;
	wire _w2075_ ;
	wire _w2076_ ;
	wire _w2077_ ;
	wire _w2078_ ;
	wire _w2079_ ;
	wire _w2080_ ;
	wire _w2081_ ;
	wire _w2082_ ;
	wire _w2083_ ;
	wire _w2084_ ;
	wire _w2085_ ;
	wire _w2086_ ;
	wire _w2087_ ;
	wire _w2088_ ;
	wire _w2089_ ;
	wire _w2090_ ;
	wire _w2091_ ;
	wire _w2092_ ;
	wire _w2093_ ;
	wire _w2094_ ;
	wire _w2095_ ;
	wire _w2096_ ;
	wire _w2097_ ;
	wire _w2098_ ;
	wire _w2099_ ;
	wire _w2100_ ;
	wire _w2101_ ;
	wire _w2102_ ;
	wire _w2103_ ;
	wire _w2104_ ;
	wire _w2105_ ;
	wire _w2106_ ;
	wire _w2107_ ;
	wire _w2108_ ;
	wire _w2109_ ;
	wire _w2110_ ;
	wire _w2111_ ;
	wire _w2112_ ;
	wire _w2113_ ;
	wire _w2114_ ;
	wire _w2115_ ;
	wire _w2116_ ;
	wire _w2117_ ;
	wire _w2118_ ;
	wire _w2119_ ;
	wire _w2120_ ;
	wire _w2121_ ;
	wire _w2122_ ;
	wire _w2123_ ;
	wire _w2124_ ;
	wire _w2125_ ;
	wire _w2126_ ;
	wire _w2127_ ;
	wire _w2128_ ;
	wire _w2129_ ;
	wire _w2130_ ;
	wire _w2131_ ;
	wire _w2132_ ;
	wire _w2133_ ;
	wire _w2134_ ;
	wire _w2135_ ;
	wire _w2136_ ;
	wire _w2137_ ;
	wire _w2138_ ;
	wire _w2139_ ;
	wire _w2140_ ;
	wire _w2141_ ;
	wire _w2142_ ;
	wire _w2143_ ;
	wire _w2144_ ;
	wire _w2145_ ;
	wire _w2146_ ;
	wire _w2147_ ;
	wire _w2148_ ;
	wire _w2149_ ;
	wire _w2150_ ;
	wire _w2151_ ;
	wire _w2152_ ;
	wire _w2153_ ;
	wire _w2154_ ;
	wire _w2155_ ;
	wire _w2156_ ;
	wire _w2157_ ;
	wire _w2158_ ;
	wire _w2159_ ;
	wire _w2160_ ;
	wire _w2161_ ;
	wire _w2162_ ;
	wire _w2163_ ;
	wire _w2164_ ;
	wire _w2165_ ;
	wire _w2166_ ;
	wire _w2167_ ;
	wire _w2168_ ;
	wire _w2169_ ;
	wire _w2170_ ;
	wire _w2171_ ;
	wire _w2172_ ;
	wire _w2173_ ;
	wire _w2174_ ;
	wire _w2175_ ;
	wire _w2176_ ;
	wire _w2177_ ;
	wire _w2178_ ;
	wire _w2179_ ;
	wire _w2180_ ;
	wire _w2181_ ;
	wire _w2182_ ;
	wire _w2183_ ;
	wire _w2184_ ;
	wire _w2185_ ;
	wire _w2186_ ;
	wire _w2187_ ;
	wire _w2188_ ;
	wire _w2189_ ;
	wire _w2190_ ;
	wire _w2191_ ;
	wire _w2192_ ;
	wire _w2193_ ;
	wire _w2194_ ;
	wire _w2195_ ;
	wire _w2196_ ;
	wire _w2197_ ;
	wire _w2198_ ;
	wire _w2199_ ;
	wire _w2200_ ;
	wire _w2201_ ;
	wire _w2202_ ;
	wire _w2203_ ;
	wire _w2204_ ;
	wire _w2205_ ;
	wire _w2206_ ;
	wire _w2207_ ;
	wire _w2208_ ;
	wire _w2209_ ;
	wire _w2210_ ;
	wire _w2211_ ;
	wire _w2212_ ;
	wire _w2213_ ;
	wire _w2214_ ;
	wire _w2215_ ;
	wire _w2216_ ;
	wire _w2217_ ;
	wire _w2218_ ;
	wire _w2219_ ;
	wire _w2220_ ;
	wire _w2221_ ;
	wire _w2222_ ;
	wire _w2223_ ;
	wire _w2224_ ;
	wire _w2225_ ;
	wire _w2226_ ;
	wire _w2227_ ;
	wire _w2228_ ;
	wire _w2229_ ;
	wire _w2230_ ;
	wire _w2231_ ;
	wire _w2232_ ;
	wire _w2233_ ;
	wire _w2234_ ;
	wire _w2235_ ;
	wire _w2236_ ;
	wire _w2237_ ;
	wire _w2238_ ;
	wire _w2239_ ;
	wire _w2240_ ;
	wire _w2241_ ;
	wire _w2242_ ;
	wire _w2243_ ;
	wire _w2244_ ;
	wire _w2245_ ;
	wire _w2246_ ;
	wire _w2247_ ;
	wire _w2248_ ;
	wire _w2249_ ;
	wire _w2250_ ;
	wire _w2251_ ;
	wire _w2252_ ;
	wire _w2253_ ;
	wire _w2254_ ;
	wire _w2255_ ;
	wire _w2256_ ;
	wire _w2257_ ;
	wire _w2258_ ;
	wire _w2259_ ;
	wire _w2260_ ;
	wire _w2261_ ;
	wire _w2262_ ;
	wire _w2263_ ;
	wire _w2264_ ;
	wire _w2265_ ;
	wire _w2266_ ;
	wire _w2267_ ;
	wire _w2268_ ;
	wire _w2269_ ;
	wire _w2270_ ;
	wire _w2271_ ;
	wire _w2272_ ;
	wire _w2273_ ;
	wire _w2274_ ;
	wire _w2275_ ;
	wire _w2276_ ;
	wire _w2277_ ;
	wire _w2278_ ;
	wire _w2279_ ;
	wire _w2280_ ;
	wire _w2281_ ;
	wire _w2282_ ;
	wire _w2283_ ;
	wire _w2284_ ;
	wire _w2285_ ;
	wire _w2286_ ;
	wire _w2287_ ;
	wire _w2288_ ;
	wire _w2289_ ;
	wire _w2290_ ;
	wire _w2291_ ;
	wire _w2292_ ;
	wire _w2293_ ;
	wire _w2294_ ;
	wire _w2295_ ;
	wire _w2296_ ;
	wire _w2297_ ;
	wire _w2298_ ;
	wire _w2299_ ;
	wire _w2300_ ;
	wire _w2301_ ;
	wire _w2302_ ;
	wire _w2303_ ;
	wire _w2304_ ;
	wire _w2305_ ;
	wire _w2306_ ;
	wire _w2307_ ;
	wire _w2308_ ;
	wire _w2309_ ;
	wire _w2310_ ;
	wire _w2311_ ;
	wire _w2312_ ;
	wire _w2313_ ;
	wire _w2314_ ;
	wire _w2315_ ;
	wire _w2316_ ;
	wire _w2317_ ;
	wire _w2318_ ;
	wire _w2319_ ;
	wire _w2320_ ;
	wire _w2321_ ;
	wire _w2322_ ;
	wire _w2323_ ;
	wire _w2324_ ;
	wire _w2325_ ;
	wire _w2326_ ;
	wire _w2327_ ;
	wire _w2328_ ;
	wire _w2329_ ;
	wire _w2330_ ;
	wire _w2331_ ;
	wire _w2332_ ;
	wire _w2333_ ;
	wire _w2334_ ;
	wire _w2335_ ;
	wire _w2336_ ;
	wire _w2337_ ;
	wire _w2338_ ;
	wire _w2339_ ;
	wire _w2340_ ;
	wire _w2341_ ;
	wire _w2342_ ;
	wire _w2343_ ;
	wire _w2344_ ;
	wire _w2345_ ;
	wire _w2346_ ;
	wire _w2347_ ;
	wire _w2348_ ;
	wire _w2349_ ;
	wire _w2350_ ;
	wire _w2351_ ;
	wire _w2352_ ;
	wire _w2353_ ;
	wire _w2354_ ;
	wire _w2355_ ;
	wire _w2356_ ;
	wire _w2357_ ;
	wire _w2358_ ;
	wire _w2359_ ;
	wire _w2360_ ;
	wire _w2361_ ;
	wire _w2362_ ;
	wire _w2363_ ;
	wire _w2364_ ;
	wire _w2365_ ;
	wire _w2366_ ;
	wire _w2367_ ;
	wire _w2368_ ;
	wire _w2369_ ;
	wire _w2370_ ;
	wire _w2371_ ;
	wire _w2372_ ;
	wire _w2373_ ;
	wire _w2374_ ;
	wire _w2375_ ;
	wire _w2376_ ;
	wire _w2377_ ;
	wire _w2378_ ;
	wire _w2379_ ;
	wire _w2380_ ;
	wire _w2381_ ;
	wire _w2382_ ;
	wire _w2383_ ;
	wire _w2384_ ;
	wire _w2385_ ;
	wire _w2386_ ;
	wire _w2387_ ;
	wire _w2388_ ;
	wire _w2389_ ;
	wire _w2390_ ;
	wire _w2391_ ;
	wire _w2392_ ;
	wire _w2393_ ;
	wire _w2394_ ;
	wire _w2395_ ;
	wire _w2396_ ;
	wire _w2397_ ;
	wire _w2398_ ;
	wire _w2399_ ;
	wire _w2400_ ;
	wire _w2401_ ;
	wire _w2402_ ;
	wire _w2403_ ;
	wire _w2404_ ;
	wire _w2405_ ;
	wire _w2406_ ;
	wire _w2407_ ;
	wire _w2408_ ;
	wire _w2409_ ;
	wire _w2410_ ;
	wire _w2411_ ;
	wire _w2412_ ;
	wire _w2413_ ;
	wire _w2414_ ;
	wire _w2415_ ;
	wire _w2416_ ;
	wire _w2417_ ;
	wire _w2418_ ;
	wire _w2419_ ;
	wire _w2420_ ;
	wire _w2421_ ;
	wire _w2422_ ;
	wire _w2423_ ;
	wire _w2424_ ;
	wire _w2425_ ;
	wire _w2426_ ;
	wire _w2427_ ;
	wire _w2428_ ;
	wire _w2429_ ;
	wire _w2430_ ;
	wire _w2431_ ;
	wire _w2432_ ;
	wire _w2433_ ;
	wire _w2434_ ;
	wire _w2435_ ;
	wire _w2436_ ;
	wire _w2437_ ;
	wire _w2438_ ;
	wire _w2439_ ;
	wire _w2440_ ;
	wire _w2441_ ;
	wire _w2442_ ;
	wire _w2443_ ;
	wire _w2444_ ;
	wire _w2445_ ;
	wire _w2446_ ;
	wire _w2447_ ;
	wire _w2448_ ;
	wire _w2449_ ;
	wire _w2450_ ;
	wire _w2451_ ;
	wire _w2452_ ;
	wire _w2453_ ;
	wire _w2454_ ;
	wire _w2455_ ;
	wire _w2456_ ;
	wire _w2457_ ;
	wire _w2458_ ;
	wire _w2459_ ;
	wire _w2460_ ;
	wire _w2461_ ;
	wire _w2462_ ;
	wire _w2463_ ;
	wire _w2464_ ;
	wire _w2465_ ;
	wire _w2466_ ;
	wire _w2467_ ;
	wire _w2468_ ;
	wire _w2469_ ;
	wire _w2470_ ;
	wire _w2471_ ;
	wire _w2472_ ;
	wire _w2473_ ;
	wire _w2474_ ;
	wire _w2475_ ;
	wire _w2476_ ;
	wire _w2477_ ;
	wire _w2478_ ;
	wire _w2479_ ;
	wire _w2480_ ;
	wire _w2481_ ;
	wire _w2482_ ;
	wire _w2483_ ;
	wire _w2484_ ;
	wire _w2485_ ;
	wire _w2486_ ;
	wire _w2487_ ;
	wire _w2488_ ;
	wire _w2489_ ;
	wire _w2490_ ;
	wire _w2491_ ;
	wire _w2492_ ;
	wire _w2493_ ;
	wire _w2494_ ;
	wire _w2495_ ;
	wire _w2496_ ;
	wire _w2497_ ;
	wire _w2498_ ;
	wire _w2499_ ;
	wire _w2500_ ;
	wire _w2501_ ;
	wire _w2502_ ;
	wire _w2503_ ;
	wire _w2504_ ;
	wire _w2505_ ;
	wire _w2506_ ;
	wire _w2507_ ;
	wire _w2508_ ;
	wire _w2509_ ;
	wire _w2510_ ;
	wire _w2511_ ;
	wire _w2512_ ;
	wire _w2513_ ;
	wire _w2514_ ;
	wire _w2515_ ;
	wire _w2516_ ;
	wire _w2517_ ;
	wire _w2518_ ;
	wire _w2519_ ;
	wire _w2520_ ;
	wire _w2521_ ;
	wire _w2522_ ;
	wire _w2523_ ;
	wire _w2524_ ;
	wire _w2525_ ;
	wire _w2526_ ;
	wire _w2527_ ;
	wire _w2528_ ;
	wire _w2529_ ;
	wire _w2530_ ;
	wire _w2531_ ;
	wire _w2532_ ;
	wire _w2533_ ;
	wire _w2534_ ;
	wire _w2535_ ;
	wire _w2536_ ;
	wire _w2537_ ;
	wire _w2538_ ;
	wire _w2539_ ;
	wire _w2540_ ;
	wire _w2541_ ;
	wire _w2542_ ;
	wire _w2543_ ;
	wire _w2544_ ;
	wire _w2545_ ;
	wire _w2546_ ;
	wire _w2547_ ;
	wire _w2548_ ;
	wire _w2549_ ;
	wire _w2550_ ;
	wire _w2551_ ;
	wire _w2552_ ;
	wire _w2553_ ;
	wire _w2554_ ;
	wire _w2555_ ;
	wire _w2556_ ;
	wire _w2557_ ;
	wire _w2558_ ;
	wire _w2559_ ;
	wire _w2560_ ;
	wire _w2561_ ;
	wire _w2562_ ;
	wire _w2563_ ;
	wire _w2564_ ;
	wire _w2565_ ;
	wire _w2566_ ;
	wire _w2567_ ;
	wire _w2568_ ;
	wire _w2569_ ;
	wire _w2570_ ;
	wire _w2571_ ;
	wire _w2572_ ;
	wire _w2573_ ;
	wire _w2574_ ;
	wire _w2575_ ;
	wire _w2576_ ;
	wire _w2577_ ;
	wire _w2578_ ;
	wire _w2579_ ;
	wire _w2580_ ;
	wire _w2581_ ;
	wire _w2582_ ;
	wire _w2583_ ;
	wire _w2584_ ;
	wire _w2585_ ;
	wire _w2586_ ;
	wire _w2587_ ;
	wire _w2588_ ;
	wire _w2589_ ;
	wire _w2590_ ;
	wire _w2591_ ;
	wire _w2592_ ;
	wire _w2593_ ;
	wire _w2594_ ;
	wire _w2595_ ;
	wire _w2596_ ;
	wire _w2597_ ;
	wire _w2598_ ;
	wire _w2599_ ;
	wire _w2600_ ;
	wire _w2601_ ;
	wire _w2602_ ;
	wire _w2603_ ;
	wire _w2604_ ;
	wire _w2605_ ;
	wire _w2606_ ;
	wire _w2607_ ;
	wire _w2608_ ;
	wire _w2609_ ;
	wire _w2610_ ;
	wire _w2611_ ;
	wire _w2612_ ;
	wire _w2613_ ;
	wire _w2614_ ;
	wire _w2615_ ;
	wire _w2616_ ;
	wire _w2617_ ;
	wire _w2618_ ;
	wire _w2619_ ;
	wire _w2620_ ;
	wire _w2621_ ;
	wire _w2622_ ;
	wire _w2623_ ;
	wire _w2624_ ;
	wire _w2625_ ;
	wire _w2626_ ;
	wire _w2627_ ;
	wire _w2628_ ;
	wire _w2629_ ;
	wire _w2630_ ;
	wire _w2631_ ;
	wire _w2632_ ;
	wire _w2633_ ;
	wire _w2634_ ;
	wire _w2635_ ;
	wire _w2636_ ;
	wire _w2637_ ;
	wire _w2638_ ;
	wire _w2639_ ;
	wire _w2640_ ;
	wire _w2641_ ;
	wire _w2642_ ;
	wire _w2643_ ;
	wire _w2644_ ;
	wire _w2645_ ;
	wire _w2646_ ;
	wire _w2647_ ;
	wire _w2648_ ;
	wire _w2649_ ;
	wire _w2650_ ;
	wire _w2651_ ;
	wire _w2652_ ;
	wire _w2653_ ;
	wire _w2654_ ;
	wire _w2655_ ;
	wire _w2656_ ;
	wire _w2657_ ;
	wire _w2658_ ;
	wire _w2659_ ;
	wire _w2660_ ;
	wire _w2661_ ;
	wire _w2662_ ;
	wire _w2663_ ;
	wire _w2664_ ;
	wire _w2665_ ;
	wire _w2666_ ;
	wire _w2667_ ;
	wire _w2668_ ;
	wire _w2669_ ;
	wire _w2670_ ;
	wire _w2671_ ;
	wire _w2672_ ;
	wire _w2673_ ;
	wire _w2674_ ;
	wire _w2675_ ;
	wire _w2676_ ;
	wire _w2677_ ;
	wire _w2678_ ;
	wire _w2679_ ;
	wire _w2680_ ;
	wire _w2681_ ;
	wire _w2682_ ;
	wire _w2683_ ;
	wire _w2684_ ;
	wire _w2685_ ;
	wire _w2686_ ;
	wire _w2687_ ;
	wire _w2688_ ;
	wire _w2689_ ;
	wire _w2690_ ;
	wire _w2691_ ;
	wire _w2692_ ;
	wire _w2693_ ;
	wire _w2694_ ;
	wire _w2695_ ;
	wire _w2696_ ;
	wire _w2697_ ;
	wire _w2698_ ;
	wire _w2699_ ;
	wire _w2700_ ;
	wire _w2701_ ;
	wire _w2702_ ;
	wire _w2703_ ;
	wire _w2704_ ;
	wire _w2705_ ;
	wire _w2706_ ;
	wire _w2707_ ;
	wire _w2708_ ;
	wire _w2709_ ;
	wire _w2710_ ;
	wire _w2711_ ;
	wire _w2712_ ;
	wire _w2713_ ;
	wire _w2714_ ;
	wire _w2715_ ;
	wire _w2716_ ;
	wire _w2717_ ;
	wire _w2718_ ;
	wire _w2719_ ;
	wire _w2720_ ;
	wire _w2721_ ;
	wire _w2722_ ;
	wire _w2723_ ;
	wire _w2724_ ;
	wire _w2725_ ;
	wire _w2726_ ;
	wire _w2727_ ;
	wire _w2728_ ;
	wire _w2729_ ;
	wire _w2730_ ;
	wire _w2731_ ;
	wire _w2732_ ;
	wire _w2733_ ;
	wire _w2734_ ;
	wire _w2735_ ;
	wire _w2736_ ;
	wire _w2737_ ;
	wire _w2738_ ;
	wire _w2739_ ;
	wire _w2740_ ;
	wire _w2741_ ;
	wire _w2742_ ;
	wire _w2743_ ;
	wire _w2744_ ;
	wire _w2745_ ;
	wire _w2746_ ;
	wire _w2747_ ;
	wire _w2748_ ;
	wire _w2749_ ;
	wire _w2750_ ;
	wire _w2751_ ;
	wire _w2752_ ;
	wire _w2753_ ;
	wire _w2754_ ;
	wire _w2755_ ;
	wire _w2756_ ;
	wire _w2757_ ;
	wire _w2758_ ;
	wire _w2759_ ;
	wire _w2760_ ;
	wire _w2761_ ;
	wire _w2762_ ;
	wire _w2763_ ;
	wire _w2764_ ;
	wire _w2765_ ;
	wire _w2766_ ;
	wire _w2767_ ;
	wire _w2768_ ;
	wire _w2769_ ;
	wire _w2770_ ;
	wire _w2771_ ;
	wire _w2772_ ;
	wire _w2773_ ;
	wire _w2774_ ;
	wire _w2775_ ;
	wire _w2776_ ;
	wire _w2777_ ;
	wire _w2778_ ;
	wire _w2779_ ;
	wire _w2780_ ;
	wire _w2781_ ;
	wire _w2782_ ;
	wire _w2783_ ;
	wire _w2784_ ;
	wire _w2785_ ;
	wire _w2786_ ;
	wire _w2787_ ;
	wire _w2788_ ;
	wire _w2789_ ;
	wire _w2790_ ;
	wire _w2791_ ;
	wire _w2792_ ;
	wire _w2793_ ;
	wire _w2794_ ;
	wire _w2795_ ;
	wire _w2796_ ;
	wire _w2797_ ;
	wire _w2798_ ;
	wire _w2799_ ;
	wire _w2800_ ;
	wire _w2801_ ;
	wire _w2802_ ;
	wire _w2803_ ;
	wire _w2804_ ;
	wire _w2805_ ;
	wire _w2806_ ;
	wire _w2807_ ;
	wire _w2808_ ;
	wire _w2809_ ;
	wire _w2810_ ;
	wire _w2811_ ;
	wire _w2812_ ;
	wire _w2813_ ;
	wire _w2814_ ;
	wire _w2815_ ;
	wire _w2816_ ;
	wire _w2817_ ;
	wire _w2818_ ;
	wire _w2819_ ;
	wire _w2820_ ;
	wire _w2821_ ;
	wire _w2822_ ;
	wire _w2823_ ;
	wire _w2824_ ;
	wire _w2825_ ;
	wire _w2826_ ;
	wire _w2827_ ;
	wire _w2828_ ;
	wire _w2829_ ;
	wire _w2830_ ;
	wire _w2831_ ;
	wire _w2832_ ;
	wire _w2833_ ;
	wire _w2834_ ;
	wire _w2835_ ;
	wire _w2836_ ;
	wire _w2837_ ;
	wire _w2838_ ;
	wire _w2839_ ;
	wire _w2840_ ;
	wire _w2841_ ;
	wire _w2842_ ;
	wire _w2843_ ;
	wire _w2844_ ;
	wire _w2845_ ;
	wire _w2846_ ;
	wire _w2847_ ;
	wire _w2848_ ;
	wire _w2849_ ;
	wire _w2850_ ;
	wire _w2851_ ;
	wire _w2852_ ;
	wire _w2853_ ;
	wire _w2854_ ;
	wire _w2855_ ;
	wire _w2856_ ;
	wire _w2857_ ;
	wire _w2858_ ;
	wire _w2859_ ;
	wire _w2860_ ;
	wire _w2861_ ;
	wire _w2862_ ;
	wire _w2863_ ;
	wire _w2864_ ;
	wire _w2865_ ;
	wire _w2866_ ;
	wire _w2867_ ;
	wire _w2868_ ;
	wire _w2869_ ;
	wire _w2870_ ;
	wire _w2871_ ;
	wire _w2872_ ;
	wire _w2873_ ;
	wire _w2874_ ;
	wire _w2875_ ;
	wire _w2876_ ;
	wire _w2877_ ;
	wire _w2878_ ;
	wire _w2879_ ;
	wire _w2880_ ;
	wire _w2881_ ;
	wire _w2882_ ;
	wire _w2883_ ;
	wire _w2884_ ;
	wire _w2885_ ;
	wire _w2886_ ;
	wire _w2887_ ;
	wire _w2888_ ;
	wire _w2889_ ;
	wire _w2890_ ;
	wire _w2891_ ;
	wire _w2892_ ;
	wire _w2893_ ;
	wire _w2894_ ;
	wire _w2895_ ;
	wire _w2896_ ;
	wire _w2897_ ;
	wire _w2898_ ;
	wire _w2899_ ;
	wire _w2900_ ;
	wire _w2901_ ;
	wire _w2902_ ;
	wire _w2903_ ;
	wire _w2904_ ;
	wire _w2905_ ;
	wire _w2906_ ;
	wire _w2907_ ;
	wire _w2908_ ;
	wire _w2909_ ;
	wire _w2910_ ;
	wire _w2911_ ;
	wire _w2912_ ;
	wire _w2913_ ;
	wire _w2914_ ;
	wire _w2915_ ;
	wire _w2916_ ;
	wire _w2917_ ;
	wire _w2918_ ;
	wire _w2919_ ;
	wire _w2920_ ;
	wire _w2921_ ;
	wire _w2922_ ;
	wire _w2923_ ;
	wire _w2924_ ;
	wire _w2925_ ;
	wire _w2926_ ;
	wire _w2927_ ;
	wire _w2928_ ;
	wire _w2929_ ;
	wire _w2930_ ;
	wire _w2931_ ;
	wire _w2932_ ;
	wire _w2933_ ;
	wire _w2934_ ;
	wire _w2935_ ;
	wire _w2936_ ;
	wire _w2937_ ;
	wire _w2938_ ;
	wire _w2939_ ;
	wire _w2940_ ;
	wire _w2941_ ;
	wire _w2942_ ;
	wire _w2943_ ;
	wire _w2944_ ;
	wire _w2945_ ;
	wire _w2946_ ;
	wire _w2947_ ;
	wire _w2948_ ;
	wire _w2949_ ;
	wire _w2950_ ;
	wire _w2951_ ;
	wire _w2952_ ;
	wire _w2953_ ;
	wire _w2954_ ;
	wire _w2955_ ;
	wire _w2956_ ;
	wire _w2957_ ;
	wire _w2958_ ;
	wire _w2959_ ;
	wire _w2960_ ;
	wire _w2961_ ;
	wire _w2962_ ;
	wire _w2963_ ;
	wire _w2964_ ;
	wire _w2965_ ;
	wire _w2966_ ;
	wire _w2967_ ;
	wire _w2968_ ;
	wire _w2969_ ;
	wire _w2970_ ;
	wire _w2971_ ;
	wire _w2972_ ;
	wire _w2973_ ;
	wire _w2974_ ;
	wire _w2975_ ;
	wire _w2976_ ;
	wire _w2977_ ;
	wire _w2978_ ;
	wire _w2979_ ;
	wire _w2980_ ;
	wire _w2981_ ;
	wire _w2982_ ;
	wire _w2983_ ;
	wire _w2984_ ;
	wire _w2985_ ;
	wire _w2986_ ;
	wire _w2987_ ;
	wire _w2988_ ;
	wire _w2989_ ;
	wire _w2990_ ;
	wire _w2991_ ;
	wire _w2992_ ;
	wire _w2993_ ;
	wire _w2994_ ;
	wire _w2995_ ;
	wire _w2996_ ;
	wire _w2997_ ;
	wire _w2998_ ;
	wire _w2999_ ;
	wire _w3000_ ;
	wire _w3001_ ;
	wire _w3002_ ;
	wire _w3003_ ;
	wire _w3004_ ;
	wire _w3005_ ;
	wire _w3006_ ;
	wire _w3007_ ;
	wire _w3008_ ;
	wire _w3009_ ;
	wire _w3010_ ;
	wire _w3011_ ;
	wire _w3012_ ;
	wire _w3013_ ;
	wire _w3014_ ;
	wire _w3015_ ;
	wire _w3016_ ;
	wire _w3017_ ;
	wire _w3018_ ;
	wire _w3019_ ;
	wire _w3020_ ;
	wire _w3021_ ;
	wire _w3022_ ;
	wire _w3023_ ;
	wire _w3024_ ;
	wire _w3025_ ;
	wire _w3026_ ;
	wire _w3027_ ;
	wire _w3028_ ;
	wire _w3029_ ;
	wire _w3030_ ;
	wire _w3031_ ;
	wire _w3032_ ;
	wire _w3033_ ;
	wire _w3034_ ;
	wire _w3035_ ;
	wire _w3036_ ;
	wire _w3037_ ;
	wire _w3038_ ;
	wire _w3039_ ;
	wire _w3040_ ;
	wire _w3041_ ;
	wire _w3042_ ;
	wire _w3043_ ;
	wire _w3044_ ;
	wire _w3045_ ;
	wire _w3046_ ;
	wire _w3047_ ;
	wire _w3048_ ;
	wire _w3049_ ;
	wire _w3050_ ;
	wire _w3051_ ;
	wire _w3052_ ;
	wire _w3053_ ;
	wire _w3054_ ;
	wire _w3055_ ;
	wire _w3056_ ;
	wire _w3057_ ;
	wire _w3058_ ;
	wire _w3059_ ;
	wire _w3060_ ;
	wire _w3061_ ;
	wire _w3062_ ;
	wire _w3063_ ;
	wire _w3064_ ;
	wire _w3065_ ;
	wire _w3066_ ;
	wire _w3067_ ;
	wire _w3068_ ;
	wire _w3069_ ;
	wire _w3070_ ;
	wire _w3071_ ;
	wire _w3072_ ;
	wire _w3073_ ;
	wire _w3074_ ;
	wire _w3075_ ;
	wire _w3076_ ;
	wire _w3077_ ;
	wire _w3078_ ;
	wire _w3079_ ;
	wire _w3080_ ;
	wire _w3081_ ;
	wire _w3082_ ;
	wire _w3083_ ;
	wire _w3084_ ;
	wire _w3085_ ;
	wire _w3086_ ;
	wire _w3087_ ;
	wire _w3088_ ;
	wire _w3089_ ;
	wire _w3090_ ;
	wire _w3091_ ;
	wire _w3092_ ;
	wire _w3093_ ;
	wire _w3094_ ;
	wire _w3095_ ;
	wire _w3096_ ;
	wire _w3097_ ;
	wire _w3098_ ;
	wire _w3099_ ;
	wire _w3100_ ;
	wire _w3101_ ;
	wire _w3102_ ;
	wire _w3103_ ;
	wire _w3104_ ;
	wire _w3105_ ;
	wire _w3106_ ;
	wire _w3107_ ;
	wire _w3108_ ;
	wire _w3109_ ;
	wire _w3110_ ;
	wire _w3111_ ;
	wire _w3112_ ;
	wire _w3113_ ;
	wire _w3114_ ;
	wire _w3115_ ;
	wire _w3116_ ;
	wire _w3117_ ;
	wire _w3118_ ;
	wire _w3119_ ;
	wire _w3120_ ;
	wire _w3121_ ;
	wire _w3122_ ;
	wire _w3123_ ;
	wire _w3124_ ;
	wire _w3125_ ;
	wire _w3126_ ;
	wire _w3127_ ;
	wire _w3128_ ;
	wire _w3129_ ;
	wire _w3130_ ;
	LUT2 #(
		.INIT('h2)
	) name0 (
		\g3003_reg/NET0131 ,
		\g35_pad ,
		_w774_
	);
	LUT2 #(
		.INIT('h1)
	) name1 (
		\g1696_reg/NET0131 ,
		\g1830_reg/NET0131 ,
		_w775_
	);
	LUT2 #(
		.INIT('h1)
	) name2 (
		\g1964_reg/NET0131 ,
		\g2098_reg/NET0131 ,
		_w776_
	);
	LUT2 #(
		.INIT('h8)
	) name3 (
		_w775_,
		_w776_,
		_w777_
	);
	LUT2 #(
		.INIT('h1)
	) name4 (
		\g2255_reg/NET0131 ,
		\g2389_reg/NET0131 ,
		_w778_
	);
	LUT2 #(
		.INIT('h1)
	) name5 (
		\g2523_reg/NET0131 ,
		\g2657_reg/NET0131 ,
		_w779_
	);
	LUT2 #(
		.INIT('h8)
	) name6 (
		_w778_,
		_w779_,
		_w780_
	);
	LUT2 #(
		.INIT('h2)
	) name7 (
		\g35_pad ,
		_w777_,
		_w781_
	);
	LUT2 #(
		.INIT('h4)
	) name8 (
		_w780_,
		_w781_,
		_w782_
	);
	LUT2 #(
		.INIT('h1)
	) name9 (
		\g1710_reg/NET0131 ,
		\g1724_reg/NET0131 ,
		_w783_
	);
	LUT2 #(
		.INIT('h1)
	) name10 (
		\g1844_reg/NET0131 ,
		\g1858_reg/NET0131 ,
		_w784_
	);
	LUT2 #(
		.INIT('h1)
	) name11 (
		\g1978_reg/NET0131 ,
		\g1992_reg/NET0131 ,
		_w785_
	);
	LUT2 #(
		.INIT('h1)
	) name12 (
		\g2112_reg/NET0131 ,
		\g2126_reg/NET0131 ,
		_w786_
	);
	LUT2 #(
		.INIT('h8)
	) name13 (
		_w785_,
		_w786_,
		_w787_
	);
	LUT2 #(
		.INIT('h8)
	) name14 (
		_w783_,
		_w784_,
		_w788_
	);
	LUT2 #(
		.INIT('h8)
	) name15 (
		_w787_,
		_w788_,
		_w789_
	);
	LUT2 #(
		.INIT('h2)
	) name16 (
		\g35_pad ,
		_w789_,
		_w790_
	);
	LUT2 #(
		.INIT('h1)
	) name17 (
		\g2269_reg/NET0131 ,
		\g2283_reg/NET0131 ,
		_w791_
	);
	LUT2 #(
		.INIT('h1)
	) name18 (
		\g2403_reg/NET0131 ,
		\g2417_reg/NET0131 ,
		_w792_
	);
	LUT2 #(
		.INIT('h1)
	) name19 (
		\g2537_reg/NET0131 ,
		\g2551_reg/NET0131 ,
		_w793_
	);
	LUT2 #(
		.INIT('h1)
	) name20 (
		\g2671_reg/NET0131 ,
		\g2685_reg/NET0131 ,
		_w794_
	);
	LUT2 #(
		.INIT('h8)
	) name21 (
		_w793_,
		_w794_,
		_w795_
	);
	LUT2 #(
		.INIT('h8)
	) name22 (
		_w791_,
		_w792_,
		_w796_
	);
	LUT2 #(
		.INIT('h8)
	) name23 (
		_w795_,
		_w796_,
		_w797_
	);
	LUT2 #(
		.INIT('h2)
	) name24 (
		_w790_,
		_w797_,
		_w798_
	);
	LUT2 #(
		.INIT('h1)
	) name25 (
		\g2204_reg/NET0131 ,
		\g2223_reg/NET0131 ,
		_w799_
	);
	LUT2 #(
		.INIT('h1)
	) name26 (
		\g2338_reg/NET0131 ,
		\g2357_reg/NET0131 ,
		_w800_
	);
	LUT2 #(
		.INIT('h1)
	) name27 (
		\g2472_reg/NET0131 ,
		\g2491_reg/NET0131 ,
		_w801_
	);
	LUT2 #(
		.INIT('h1)
	) name28 (
		\g2606_reg/NET0131 ,
		\g2625_reg/NET0131 ,
		_w802_
	);
	LUT2 #(
		.INIT('h8)
	) name29 (
		_w801_,
		_w802_,
		_w803_
	);
	LUT2 #(
		.INIT('h8)
	) name30 (
		_w799_,
		_w800_,
		_w804_
	);
	LUT2 #(
		.INIT('h8)
	) name31 (
		_w803_,
		_w804_,
		_w805_
	);
	LUT2 #(
		.INIT('h2)
	) name32 (
		\g35_pad ,
		_w805_,
		_w806_
	);
	LUT2 #(
		.INIT('h1)
	) name33 (
		\g1644_reg/NET0131 ,
		\g1664_reg/NET0131 ,
		_w807_
	);
	LUT2 #(
		.INIT('h1)
	) name34 (
		\g1779_reg/NET0131 ,
		\g1798_reg/NET0131 ,
		_w808_
	);
	LUT2 #(
		.INIT('h1)
	) name35 (
		\g1913_reg/NET0131 ,
		\g1932_reg/NET0131 ,
		_w809_
	);
	LUT2 #(
		.INIT('h1)
	) name36 (
		\g2047_reg/NET0131 ,
		\g2066_reg/NET0131 ,
		_w810_
	);
	LUT2 #(
		.INIT('h8)
	) name37 (
		_w809_,
		_w810_,
		_w811_
	);
	LUT2 #(
		.INIT('h8)
	) name38 (
		_w807_,
		_w808_,
		_w812_
	);
	LUT2 #(
		.INIT('h8)
	) name39 (
		_w811_,
		_w812_,
		_w813_
	);
	LUT2 #(
		.INIT('h2)
	) name40 (
		_w806_,
		_w813_,
		_w814_
	);
	LUT2 #(
		.INIT('h1)
	) name41 (
		\g1008_reg/NET0131 ,
		\g969_reg/NET0131 ,
		_w815_
	);
	LUT2 #(
		.INIT('h2)
	) name42 (
		\g1193_reg/NET0131 ,
		_w815_,
		_w816_
	);
	LUT2 #(
		.INIT('h1)
	) name43 (
		\g1312_reg/NET0131 ,
		\g1351_reg/NET0131 ,
		_w817_
	);
	LUT2 #(
		.INIT('h2)
	) name44 (
		\g1536_reg/NET0131 ,
		_w817_,
		_w818_
	);
	LUT2 #(
		.INIT('h2)
	) name45 (
		\g35_pad ,
		_w816_,
		_w819_
	);
	LUT2 #(
		.INIT('h4)
	) name46 (
		_w818_,
		_w819_,
		_w820_
	);
	LUT2 #(
		.INIT('h4)
	) name47 (
		\g1306_reg/NET0131 ,
		\g35_pad ,
		_w821_
	);
	LUT2 #(
		.INIT('h4)
	) name48 (
		\g962_reg/NET0131 ,
		_w821_,
		_w822_
	);
	LUT2 #(
		.INIT('h1)
	) name49 (
		\g3115_reg/NET0131 ,
		\g3466_reg/NET0131 ,
		_w823_
	);
	LUT2 #(
		.INIT('h1)
	) name50 (
		\g3817_reg/NET0131 ,
		\g5124_reg/NET0131 ,
		_w824_
	);
	LUT2 #(
		.INIT('h8)
	) name51 (
		_w823_,
		_w824_,
		_w825_
	);
	LUT2 #(
		.INIT('h2)
	) name52 (
		\g35_pad ,
		_w825_,
		_w826_
	);
	LUT2 #(
		.INIT('h8)
	) name53 (
		\g5297_reg/NET0131 ,
		\g5357_reg/NET0131 ,
		_w827_
	);
	LUT2 #(
		.INIT('h4)
	) name54 (
		\g1636_reg/NET0131 ,
		\g1668_reg/NET0131 ,
		_w828_
	);
	LUT2 #(
		.INIT('h2)
	) name55 (
		\g1648_reg/NET0131 ,
		\g1657_reg/NET0131 ,
		_w829_
	);
	LUT2 #(
		.INIT('h8)
	) name56 (
		\g2970_reg/NET0131 ,
		\g2975_reg/NET0131 ,
		_w830_
	);
	LUT2 #(
		.INIT('h8)
	) name57 (
		\g2960_reg/NET0131 ,
		\g2965_reg/NET0131 ,
		_w831_
	);
	LUT2 #(
		.INIT('h8)
	) name58 (
		\g2922_reg/NET0131 ,
		\g2927_reg/NET0131 ,
		_w832_
	);
	LUT2 #(
		.INIT('h8)
	) name59 (
		\g2950_reg/NET0131 ,
		\g2955_reg/NET0131 ,
		_w833_
	);
	LUT2 #(
		.INIT('h8)
	) name60 (
		\g2912_reg/NET0131 ,
		\g2917_reg/NET0131 ,
		_w834_
	);
	LUT2 #(
		.INIT('h8)
	) name61 (
		\g2936_reg/NET0131 ,
		\g2941_reg/NET0131 ,
		_w835_
	);
	LUT2 #(
		.INIT('h8)
	) name62 (
		\g2902_reg/NET0131 ,
		\g2907_reg/NET0131 ,
		_w836_
	);
	LUT2 #(
		.INIT('h1)
	) name63 (
		_w830_,
		_w831_,
		_w837_
	);
	LUT2 #(
		.INIT('h1)
	) name64 (
		_w832_,
		_w833_,
		_w838_
	);
	LUT2 #(
		.INIT('h1)
	) name65 (
		_w834_,
		_w835_,
		_w839_
	);
	LUT2 #(
		.INIT('h4)
	) name66 (
		_w836_,
		_w839_,
		_w840_
	);
	LUT2 #(
		.INIT('h8)
	) name67 (
		_w837_,
		_w838_,
		_w841_
	);
	LUT2 #(
		.INIT('h8)
	) name68 (
		_w840_,
		_w841_,
		_w842_
	);
	LUT2 #(
		.INIT('h4)
	) name69 (
		\g2724_reg/NET0131 ,
		\g2815_reg/NET0131 ,
		_w843_
	);
	LUT2 #(
		.INIT('h8)
	) name70 (
		\g2724_reg/NET0131 ,
		\g2819_reg/NET0131 ,
		_w844_
	);
	LUT2 #(
		.INIT('h2)
	) name71 (
		\g2729_reg/NET0131 ,
		_w843_,
		_w845_
	);
	LUT2 #(
		.INIT('h4)
	) name72 (
		_w844_,
		_w845_,
		_w846_
	);
	LUT2 #(
		.INIT('h4)
	) name73 (
		\g2724_reg/NET0131 ,
		\g2803_reg/NET0131 ,
		_w847_
	);
	LUT2 #(
		.INIT('h8)
	) name74 (
		\g2724_reg/NET0131 ,
		\g2807_reg/NET0131 ,
		_w848_
	);
	LUT2 #(
		.INIT('h1)
	) name75 (
		\g2729_reg/NET0131 ,
		_w847_,
		_w849_
	);
	LUT2 #(
		.INIT('h4)
	) name76 (
		_w848_,
		_w849_,
		_w850_
	);
	LUT2 #(
		.INIT('h1)
	) name77 (
		_w846_,
		_w850_,
		_w851_
	);
	LUT2 #(
		.INIT('h4)
	) name78 (
		\g2724_reg/NET0131 ,
		\g2783_reg/NET0131 ,
		_w852_
	);
	LUT2 #(
		.INIT('h8)
	) name79 (
		\g2724_reg/NET0131 ,
		\g2787_reg/NET0131 ,
		_w853_
	);
	LUT2 #(
		.INIT('h2)
	) name80 (
		\g2729_reg/NET0131 ,
		_w852_,
		_w854_
	);
	LUT2 #(
		.INIT('h4)
	) name81 (
		_w853_,
		_w854_,
		_w855_
	);
	LUT2 #(
		.INIT('h4)
	) name82 (
		\g2724_reg/NET0131 ,
		\g2771_reg/NET0131 ,
		_w856_
	);
	LUT2 #(
		.INIT('h8)
	) name83 (
		\g2724_reg/NET0131 ,
		\g2775_reg/NET0131 ,
		_w857_
	);
	LUT2 #(
		.INIT('h1)
	) name84 (
		\g2729_reg/NET0131 ,
		_w856_,
		_w858_
	);
	LUT2 #(
		.INIT('h4)
	) name85 (
		_w857_,
		_w858_,
		_w859_
	);
	LUT2 #(
		.INIT('h1)
	) name86 (
		_w855_,
		_w859_,
		_w860_
	);
	LUT2 #(
		.INIT('h1)
	) name87 (
		\g4709_reg/NET0131 ,
		\g4785_reg/NET0131 ,
		_w861_
	);
	LUT2 #(
		.INIT('h8)
	) name88 (
		\g4698_reg/NET0131 ,
		_w861_,
		_w862_
	);
	LUT2 #(
		.INIT('h2)
	) name89 (
		\g4776_reg/NET0131 ,
		\g4801_reg/NET0131 ,
		_w863_
	);
	LUT2 #(
		.INIT('h4)
	) name90 (
		\g4793_reg/NET0131 ,
		_w863_,
		_w864_
	);
	LUT2 #(
		.INIT('h8)
	) name91 (
		\g4659_reg/NET0131 ,
		\g4669_reg/NET0131 ,
		_w865_
	);
	LUT2 #(
		.INIT('h8)
	) name92 (
		\g4653_reg/NET0131 ,
		_w865_,
		_w866_
	);
	LUT2 #(
		.INIT('h8)
	) name93 (
		_w864_,
		_w866_,
		_w867_
	);
	LUT2 #(
		.INIT('h8)
	) name94 (
		_w862_,
		_w867_,
		_w868_
	);
	LUT2 #(
		.INIT('h2)
	) name95 (
		\g4646_reg/NET0131 ,
		_w868_,
		_w869_
	);
	LUT2 #(
		.INIT('h1)
	) name96 (
		\g4057_reg/NET0131 ,
		\g4064_reg/NET0131 ,
		_w870_
	);
	LUT2 #(
		.INIT('h1)
	) name97 (
		\g4082_reg/NET0131 ,
		\g4141_reg/NET0131 ,
		_w871_
	);
	LUT2 #(
		.INIT('h1)
	) name98 (
		\g4087_reg/NET0131 ,
		\g4093_reg/NET0131 ,
		_w872_
	);
	LUT2 #(
		.INIT('h4)
	) name99 (
		\g4098_reg/NET0131 ,
		_w872_,
		_w873_
	);
	LUT2 #(
		.INIT('h8)
	) name100 (
		\g4076_reg/NET0131 ,
		\g4112_reg/NET0131 ,
		_w874_
	);
	LUT2 #(
		.INIT('h8)
	) name101 (
		_w873_,
		_w874_,
		_w875_
	);
	LUT2 #(
		.INIT('h2)
	) name102 (
		_w871_,
		_w875_,
		_w876_
	);
	LUT2 #(
		.INIT('h2)
	) name103 (
		_w870_,
		_w876_,
		_w877_
	);
	LUT2 #(
		.INIT('h1)
	) name104 (
		\g482_reg/NET0131 ,
		\g490_reg/NET0131 ,
		_w878_
	);
	LUT2 #(
		.INIT('h4)
	) name105 (
		\g528_reg/NET0131 ,
		_w878_,
		_w879_
	);
	LUT2 #(
		.INIT('h8)
	) name106 (
		\g479_reg/NET0131 ,
		_w879_,
		_w880_
	);
	LUT2 #(
		.INIT('h2)
	) name107 (
		\g890_reg/NET0131 ,
		_w880_,
		_w881_
	);
	LUT2 #(
		.INIT('h1)
	) name108 (
		\g4311_reg/NET0131 ,
		\g4322_reg/NET0131 ,
		_w882_
	);
	LUT2 #(
		.INIT('h1)
	) name109 (
		\g4332_reg/NET0131 ,
		\g4366_reg/NET0131 ,
		_w883_
	);
	LUT2 #(
		.INIT('h8)
	) name110 (
		_w882_,
		_w883_,
		_w884_
	);
	LUT2 #(
		.INIT('h2)
	) name111 (
		\g4369_reg/NET0131 ,
		_w884_,
		_w885_
	);
	LUT2 #(
		.INIT('h2)
	) name112 (
		\g3111_reg/NET0131 ,
		\g35_pad ,
		_w886_
	);
	LUT2 #(
		.INIT('h8)
	) name113 (
		\g4709_reg/NET0131 ,
		\g4785_reg/NET0131 ,
		_w887_
	);
	LUT2 #(
		.INIT('h8)
	) name114 (
		\g4765_reg/NET0131 ,
		_w887_,
		_w888_
	);
	LUT2 #(
		.INIT('h8)
	) name115 (
		_w867_,
		_w888_,
		_w889_
	);
	LUT2 #(
		.INIT('h2)
	) name116 (
		\g4688_reg/NET0131 ,
		_w889_,
		_w890_
	);
	LUT2 #(
		.INIT('h2)
	) name117 (
		\g35_pad ,
		_w890_,
		_w891_
	);
	LUT2 #(
		.INIT('h8)
	) name118 (
		\g3808_reg/NET0131 ,
		_w891_,
		_w892_
	);
	LUT2 #(
		.INIT('h8)
	) name119 (
		\g35_pad ,
		_w890_,
		_w893_
	);
	LUT2 #(
		.INIT('h8)
	) name120 (
		\g16624_pad ,
		\g3338_reg/NET0131 ,
		_w894_
	);
	LUT2 #(
		.INIT('h8)
	) name121 (
		\g3990_reg/NET0131 ,
		_w894_,
		_w895_
	);
	LUT2 #(
		.INIT('h8)
	) name122 (
		\g4054_reg/NET0131 ,
		_w895_,
		_w896_
	);
	LUT2 #(
		.INIT('h2)
	) name123 (
		\g3808_reg/NET0131 ,
		_w896_,
		_w897_
	);
	LUT2 #(
		.INIT('h8)
	) name124 (
		\g3191_reg/NET0131 ,
		\g3303_reg/NET0131 ,
		_w898_
	);
	LUT2 #(
		.INIT('h8)
	) name125 (
		\g16874_pad ,
		\g3215_reg/NET0131 ,
		_w899_
	);
	LUT2 #(
		.INIT('h1)
	) name126 (
		_w898_,
		_w899_,
		_w900_
	);
	LUT2 #(
		.INIT('h2)
	) name127 (
		\g3338_reg/NET0131 ,
		_w900_,
		_w901_
	);
	LUT2 #(
		.INIT('h8)
	) name128 (
		\g16686_pad ,
		\g3255_reg/NET0131 ,
		_w902_
	);
	LUT2 #(
		.INIT('h8)
	) name129 (
		\g16624_pad ,
		\g3203_reg/NET0131 ,
		_w903_
	);
	LUT2 #(
		.INIT('h1)
	) name130 (
		_w902_,
		_w903_,
		_w904_
	);
	LUT2 #(
		.INIT('h1)
	) name131 (
		\g3338_reg/NET0131 ,
		_w904_,
		_w905_
	);
	LUT2 #(
		.INIT('h1)
	) name132 (
		\g3303_reg/NET0131 ,
		\g3338_reg/NET0131 ,
		_w906_
	);
	LUT2 #(
		.INIT('h8)
	) name133 (
		\g3303_reg/NET0131 ,
		\g3338_reg/NET0131 ,
		_w907_
	);
	LUT2 #(
		.INIT('h1)
	) name134 (
		_w906_,
		_w907_,
		_w908_
	);
	LUT2 #(
		.INIT('h8)
	) name135 (
		\g16718_pad ,
		\g3243_reg/NET0131 ,
		_w909_
	);
	LUT2 #(
		.INIT('h8)
	) name136 (
		_w908_,
		_w909_,
		_w910_
	);
	LUT2 #(
		.INIT('h1)
	) name137 (
		_w901_,
		_w905_,
		_w911_
	);
	LUT2 #(
		.INIT('h4)
	) name138 (
		_w910_,
		_w911_,
		_w912_
	);
	LUT2 #(
		.INIT('h4)
	) name139 (
		\g3990_reg/NET0131 ,
		_w912_,
		_w913_
	);
	LUT2 #(
		.INIT('h8)
	) name140 (
		\g16686_pad ,
		\g3247_reg/NET0131 ,
		_w914_
	);
	LUT2 #(
		.INIT('h8)
	) name141 (
		\g16624_pad ,
		\g3263_reg/NET0131 ,
		_w915_
	);
	LUT2 #(
		.INIT('h1)
	) name142 (
		_w914_,
		_w915_,
		_w916_
	);
	LUT2 #(
		.INIT('h2)
	) name143 (
		\g3338_reg/NET0131 ,
		_w916_,
		_w917_
	);
	LUT2 #(
		.INIT('h8)
	) name144 (
		\g16874_pad ,
		\g3223_reg/NET0131 ,
		_w918_
	);
	LUT2 #(
		.INIT('h8)
	) name145 (
		\g3207_reg/NET0131 ,
		\g3303_reg/NET0131 ,
		_w919_
	);
	LUT2 #(
		.INIT('h1)
	) name146 (
		_w918_,
		_w919_,
		_w920_
	);
	LUT2 #(
		.INIT('h1)
	) name147 (
		\g3338_reg/NET0131 ,
		_w920_,
		_w921_
	);
	LUT2 #(
		.INIT('h8)
	) name148 (
		\g16718_pad ,
		\g3235_reg/NET0131 ,
		_w922_
	);
	LUT2 #(
		.INIT('h4)
	) name149 (
		_w908_,
		_w922_,
		_w923_
	);
	LUT2 #(
		.INIT('h1)
	) name150 (
		_w917_,
		_w921_,
		_w924_
	);
	LUT2 #(
		.INIT('h4)
	) name151 (
		_w923_,
		_w924_,
		_w925_
	);
	LUT2 #(
		.INIT('h8)
	) name152 (
		\g3990_reg/NET0131 ,
		_w925_,
		_w926_
	);
	LUT2 #(
		.INIT('h2)
	) name153 (
		\g4054_reg/NET0131 ,
		_w913_,
		_w927_
	);
	LUT2 #(
		.INIT('h4)
	) name154 (
		_w926_,
		_w927_,
		_w928_
	);
	LUT2 #(
		.INIT('h8)
	) name155 (
		\g13039_pad ,
		\g3187_reg/NET0131 ,
		_w929_
	);
	LUT2 #(
		.INIT('h8)
	) name156 (
		\g3195_reg/NET0131 ,
		\g3329_reg/NET0131 ,
		_w930_
	);
	LUT2 #(
		.INIT('h1)
	) name157 (
		_w929_,
		_w930_,
		_w931_
	);
	LUT2 #(
		.INIT('h2)
	) name158 (
		\g3338_reg/NET0131 ,
		_w931_,
		_w932_
	);
	LUT2 #(
		.INIT('h8)
	) name159 (
		\g13865_pad ,
		\g3239_reg/NET0131 ,
		_w933_
	);
	LUT2 #(
		.INIT('h4)
	) name160 (
		\g3338_reg/NET0131 ,
		_w933_,
		_w934_
	);
	LUT2 #(
		.INIT('h8)
	) name161 (
		\g13895_pad ,
		\g3227_reg/NET0131 ,
		_w935_
	);
	LUT2 #(
		.INIT('h2)
	) name162 (
		_w908_,
		_w935_,
		_w936_
	);
	LUT2 #(
		.INIT('h8)
	) name163 (
		\g16603_pad ,
		\g3251_reg/NET0131 ,
		_w937_
	);
	LUT2 #(
		.INIT('h1)
	) name164 (
		_w908_,
		_w937_,
		_w938_
	);
	LUT2 #(
		.INIT('h1)
	) name165 (
		_w936_,
		_w938_,
		_w939_
	);
	LUT2 #(
		.INIT('h1)
	) name166 (
		_w932_,
		_w934_,
		_w940_
	);
	LUT2 #(
		.INIT('h4)
	) name167 (
		_w939_,
		_w940_,
		_w941_
	);
	LUT2 #(
		.INIT('h4)
	) name168 (
		\g3990_reg/NET0131 ,
		_w941_,
		_w942_
	);
	LUT2 #(
		.INIT('h8)
	) name169 (
		\g13039_pad ,
		\g3199_reg/NET0131 ,
		_w943_
	);
	LUT2 #(
		.INIT('h8)
	) name170 (
		\g3211_reg/NET0131 ,
		\g3329_reg/NET0131 ,
		_w944_
	);
	LUT2 #(
		.INIT('h1)
	) name171 (
		_w943_,
		_w944_,
		_w945_
	);
	LUT2 #(
		.INIT('h1)
	) name172 (
		\g3338_reg/NET0131 ,
		_w945_,
		_w946_
	);
	LUT2 #(
		.INIT('h8)
	) name173 (
		\g13865_pad ,
		\g3231_reg/NET0131 ,
		_w947_
	);
	LUT2 #(
		.INIT('h8)
	) name174 (
		\g3338_reg/NET0131 ,
		_w947_,
		_w948_
	);
	LUT2 #(
		.INIT('h8)
	) name175 (
		\g16603_pad ,
		\g3259_reg/NET0131 ,
		_w949_
	);
	LUT2 #(
		.INIT('h2)
	) name176 (
		_w908_,
		_w949_,
		_w950_
	);
	LUT2 #(
		.INIT('h8)
	) name177 (
		\g13895_pad ,
		\g3219_reg/NET0131 ,
		_w951_
	);
	LUT2 #(
		.INIT('h1)
	) name178 (
		_w908_,
		_w951_,
		_w952_
	);
	LUT2 #(
		.INIT('h1)
	) name179 (
		_w950_,
		_w952_,
		_w953_
	);
	LUT2 #(
		.INIT('h1)
	) name180 (
		_w946_,
		_w948_,
		_w954_
	);
	LUT2 #(
		.INIT('h4)
	) name181 (
		_w953_,
		_w954_,
		_w955_
	);
	LUT2 #(
		.INIT('h8)
	) name182 (
		\g3990_reg/NET0131 ,
		_w955_,
		_w956_
	);
	LUT2 #(
		.INIT('h1)
	) name183 (
		\g4054_reg/NET0131 ,
		_w942_,
		_w957_
	);
	LUT2 #(
		.INIT('h4)
	) name184 (
		_w956_,
		_w957_,
		_w958_
	);
	LUT2 #(
		.INIT('h1)
	) name185 (
		_w928_,
		_w958_,
		_w959_
	);
	LUT2 #(
		.INIT('h2)
	) name186 (
		_w897_,
		_w959_,
		_w960_
	);
	LUT2 #(
		.INIT('h4)
	) name187 (
		_w897_,
		_w959_,
		_w961_
	);
	LUT2 #(
		.INIT('h2)
	) name188 (
		_w893_,
		_w960_,
		_w962_
	);
	LUT2 #(
		.INIT('h4)
	) name189 (
		_w961_,
		_w962_,
		_w963_
	);
	LUT2 #(
		.INIT('h1)
	) name190 (
		_w886_,
		_w892_,
		_w964_
	);
	LUT2 #(
		.INIT('h4)
	) name191 (
		_w963_,
		_w964_,
		_w965_
	);
	LUT2 #(
		.INIT('h4)
	) name192 (
		\g736_reg/NET0131 ,
		\g802_reg/NET0131 ,
		_w966_
	);
	LUT2 #(
		.INIT('h2)
	) name193 (
		\g35_pad ,
		_w966_,
		_w967_
	);
	LUT2 #(
		.INIT('h8)
	) name194 (
		\g554_reg/NET0131 ,
		_w967_,
		_w968_
	);
	LUT2 #(
		.INIT('h4)
	) name195 (
		\g35_pad ,
		\g807_reg/NET0131 ,
		_w969_
	);
	LUT2 #(
		.INIT('h8)
	) name196 (
		\g807_reg/NET0131 ,
		_w967_,
		_w970_
	);
	LUT2 #(
		.INIT('h2)
	) name197 (
		\g772_reg/NET0131 ,
		_w966_,
		_w971_
	);
	LUT2 #(
		.INIT('h2)
	) name198 (
		\g12184_pad ,
		\g802_reg/NET0131 ,
		_w972_
	);
	LUT2 #(
		.INIT('h8)
	) name199 (
		\g655_reg/NET0131 ,
		\g718_reg/NET0131 ,
		_w973_
	);
	LUT2 #(
		.INIT('h8)
	) name200 (
		\g753_reg/NET0131 ,
		_w973_,
		_w974_
	);
	LUT2 #(
		.INIT('h4)
	) name201 (
		\g370_reg/NET0131 ,
		\g385_reg/NET0131 ,
		_w975_
	);
	LUT2 #(
		.INIT('h1)
	) name202 (
		\g655_reg/NET0131 ,
		\g718_reg/NET0131 ,
		_w976_
	);
	LUT2 #(
		.INIT('h4)
	) name203 (
		\g753_reg/NET0131 ,
		_w976_,
		_w977_
	);
	LUT2 #(
		.INIT('h4)
	) name204 (
		_w974_,
		_w975_,
		_w978_
	);
	LUT2 #(
		.INIT('h4)
	) name205 (
		_w977_,
		_w978_,
		_w979_
	);
	LUT2 #(
		.INIT('h4)
	) name206 (
		_w972_,
		_w979_,
		_w980_
	);
	LUT2 #(
		.INIT('h8)
	) name207 (
		\g554_reg/NET0131 ,
		\g807_reg/NET0131 ,
		_w981_
	);
	LUT2 #(
		.INIT('h1)
	) name208 (
		\g499_reg/NET0131 ,
		\g518_reg/NET0131 ,
		_w982_
	);
	LUT2 #(
		.INIT('h8)
	) name209 (
		_w879_,
		_w982_,
		_w983_
	);
	LUT2 #(
		.INIT('h4)
	) name210 (
		_w981_,
		_w983_,
		_w984_
	);
	LUT2 #(
		.INIT('h2)
	) name211 (
		\g749_reg/NET0131 ,
		_w966_,
		_w985_
	);
	LUT2 #(
		.INIT('h8)
	) name212 (
		\g758_reg/NET0131 ,
		_w985_,
		_w986_
	);
	LUT2 #(
		.INIT('h8)
	) name213 (
		\g358_reg/NET0131 ,
		\g376_reg/NET0131 ,
		_w987_
	);
	LUT2 #(
		.INIT('h8)
	) name214 (
		\g739_reg/NET0131 ,
		\g744_reg/NET0131 ,
		_w988_
	);
	LUT2 #(
		.INIT('h8)
	) name215 (
		\g763_reg/NET0131 ,
		\g767_reg/NET0131 ,
		_w989_
	);
	LUT2 #(
		.INIT('h8)
	) name216 (
		_w988_,
		_w989_,
		_w990_
	);
	LUT2 #(
		.INIT('h4)
	) name217 (
		_w966_,
		_w987_,
		_w991_
	);
	LUT2 #(
		.INIT('h8)
	) name218 (
		_w990_,
		_w991_,
		_w992_
	);
	LUT2 #(
		.INIT('h8)
	) name219 (
		_w986_,
		_w992_,
		_w993_
	);
	LUT2 #(
		.INIT('h8)
	) name220 (
		_w984_,
		_w993_,
		_w994_
	);
	LUT2 #(
		.INIT('h8)
	) name221 (
		_w980_,
		_w994_,
		_w995_
	);
	LUT2 #(
		.INIT('h8)
	) name222 (
		_w971_,
		_w995_,
		_w996_
	);
	LUT2 #(
		.INIT('h8)
	) name223 (
		\g776_reg/NET0131 ,
		_w996_,
		_w997_
	);
	LUT2 #(
		.INIT('h2)
	) name224 (
		\g785_reg/NET0131 ,
		_w966_,
		_w998_
	);
	LUT2 #(
		.INIT('h8)
	) name225 (
		\g781_reg/NET0131 ,
		\g790_reg/NET0131 ,
		_w999_
	);
	LUT2 #(
		.INIT('h8)
	) name226 (
		_w998_,
		_w999_,
		_w1000_
	);
	LUT2 #(
		.INIT('h8)
	) name227 (
		_w997_,
		_w1000_,
		_w1001_
	);
	LUT2 #(
		.INIT('h8)
	) name228 (
		\g794_reg/NET0131 ,
		_w1001_,
		_w1002_
	);
	LUT2 #(
		.INIT('h4)
	) name229 (
		\g554_reg/NET0131 ,
		_w970_,
		_w1003_
	);
	LUT2 #(
		.INIT('h8)
	) name230 (
		_w1002_,
		_w1003_,
		_w1004_
	);
	LUT2 #(
		.INIT('h1)
	) name231 (
		_w968_,
		_w969_,
		_w1005_
	);
	LUT2 #(
		.INIT('h4)
	) name232 (
		_w1004_,
		_w1005_,
		_w1006_
	);
	LUT2 #(
		.INIT('h1)
	) name233 (
		\g2941_reg/NET0131 ,
		\g35_pad ,
		_w1007_
	);
	LUT2 #(
		.INIT('h8)
	) name234 (
		\g35_pad ,
		_w777_,
		_w1008_
	);
	LUT2 #(
		.INIT('h8)
	) name235 (
		_w780_,
		_w1008_,
		_w1009_
	);
	LUT2 #(
		.INIT('h1)
	) name236 (
		\g3129_reg/NET0131 ,
		\g3143_reg/NET0131 ,
		_w1010_
	);
	LUT2 #(
		.INIT('h1)
	) name237 (
		\g3480_reg/NET0131 ,
		\g3494_reg/NET0131 ,
		_w1011_
	);
	LUT2 #(
		.INIT('h1)
	) name238 (
		\g3831_reg/NET0131 ,
		\g3845_reg/NET0131 ,
		_w1012_
	);
	LUT2 #(
		.INIT('h1)
	) name239 (
		\g5138_reg/NET0131 ,
		\g5152_reg/NET0131 ,
		_w1013_
	);
	LUT2 #(
		.INIT('h8)
	) name240 (
		_w1012_,
		_w1013_,
		_w1014_
	);
	LUT2 #(
		.INIT('h8)
	) name241 (
		_w1010_,
		_w1011_,
		_w1015_
	);
	LUT2 #(
		.INIT('h8)
	) name242 (
		_w1014_,
		_w1015_,
		_w1016_
	);
	LUT2 #(
		.INIT('h1)
	) name243 (
		\g4420_reg/NET0131 ,
		\g4427_reg/NET0131 ,
		_w1017_
	);
	LUT2 #(
		.INIT('h1)
	) name244 (
		\g2946_reg/NET0131 ,
		\g2955_reg/NET0131 ,
		_w1018_
	);
	LUT2 #(
		.INIT('h8)
	) name245 (
		_w1017_,
		_w1018_,
		_w1019_
	);
	LUT2 #(
		.INIT('h8)
	) name246 (
		_w825_,
		_w1019_,
		_w1020_
	);
	LUT2 #(
		.INIT('h8)
	) name247 (
		_w789_,
		_w1020_,
		_w1021_
	);
	LUT2 #(
		.INIT('h8)
	) name248 (
		_w797_,
		_w1016_,
		_w1022_
	);
	LUT2 #(
		.INIT('h8)
	) name249 (
		_w1021_,
		_w1022_,
		_w1023_
	);
	LUT2 #(
		.INIT('h8)
	) name250 (
		_w1009_,
		_w1023_,
		_w1024_
	);
	LUT2 #(
		.INIT('h1)
	) name251 (
		_w1007_,
		_w1024_,
		_w1025_
	);
	LUT2 #(
		.INIT('h1)
	) name252 (
		\g2856_reg/NET0131 ,
		\g35_pad ,
		_w1026_
	);
	LUT2 #(
		.INIT('h4)
	) name253 (
		\g2864_reg/NET0131 ,
		\g35_pad ,
		_w1027_
	);
	LUT2 #(
		.INIT('h8)
	) name254 (
		_w1017_,
		_w1027_,
		_w1028_
	);
	LUT2 #(
		.INIT('h8)
	) name255 (
		_w825_,
		_w1028_,
		_w1029_
	);
	LUT2 #(
		.INIT('h1)
	) name256 (
		_w1026_,
		_w1029_,
		_w1030_
	);
	LUT2 #(
		.INIT('h8)
	) name257 (
		\g10306_pad ,
		\g35_pad ,
		_w1031_
	);
	LUT2 #(
		.INIT('h1)
	) name258 (
		\g4534_reg/NET0131 ,
		_w1031_,
		_w1032_
	);
	LUT2 #(
		.INIT('h8)
	) name259 (
		\g4534_reg/NET0131 ,
		_w1031_,
		_w1033_
	);
	LUT2 #(
		.INIT('h1)
	) name260 (
		_w1032_,
		_w1033_,
		_w1034_
	);
	LUT2 #(
		.INIT('h8)
	) name261 (
		\g4555_reg/NET0131 ,
		\g4558_reg/NET0131 ,
		_w1035_
	);
	LUT2 #(
		.INIT('h8)
	) name262 (
		\g4561_reg/NET0131 ,
		_w1035_,
		_w1036_
	);
	LUT2 #(
		.INIT('h2)
	) name263 (
		\g35_pad ,
		_w1036_,
		_w1037_
	);
	LUT2 #(
		.INIT('h2)
	) name264 (
		\g4564_reg/NET0131 ,
		_w1037_,
		_w1038_
	);
	LUT2 #(
		.INIT('h8)
	) name265 (
		\g2988_reg/NET0131 ,
		\g35_pad ,
		_w1039_
	);
	LUT2 #(
		.INIT('h1)
	) name266 (
		_w1038_,
		_w1039_,
		_w1040_
	);
	LUT2 #(
		.INIT('h4)
	) name267 (
		\g35_pad ,
		\g4561_reg/NET0131 ,
		_w1041_
	);
	LUT2 #(
		.INIT('h8)
	) name268 (
		\g18096_pad ,
		\g35_pad ,
		_w1042_
	);
	LUT2 #(
		.INIT('h1)
	) name269 (
		_w1041_,
		_w1042_,
		_w1043_
	);
	LUT2 #(
		.INIT('h4)
	) name270 (
		\g35_pad ,
		\g4558_reg/NET0131 ,
		_w1044_
	);
	LUT2 #(
		.INIT('h8)
	) name271 (
		\g18095_pad ,
		\g35_pad ,
		_w1045_
	);
	LUT2 #(
		.INIT('h1)
	) name272 (
		_w1044_,
		_w1045_,
		_w1046_
	);
	LUT2 #(
		.INIT('h4)
	) name273 (
		\g35_pad ,
		\g4555_reg/NET0131 ,
		_w1047_
	);
	LUT2 #(
		.INIT('h8)
	) name274 (
		\g18094_pad ,
		\g35_pad ,
		_w1048_
	);
	LUT2 #(
		.INIT('h1)
	) name275 (
		_w1047_,
		_w1048_,
		_w1049_
	);
	LUT2 #(
		.INIT('h8)
	) name276 (
		\g4483_reg/NET0131 ,
		\g4486_reg/NET0131 ,
		_w1050_
	);
	LUT2 #(
		.INIT('h8)
	) name277 (
		\g4489_reg/NET0131 ,
		\g4492_reg/NET0131 ,
		_w1051_
	);
	LUT2 #(
		.INIT('h8)
	) name278 (
		_w1050_,
		_w1051_,
		_w1052_
	);
	LUT2 #(
		.INIT('h1)
	) name279 (
		\g4527_reg/NET0131 ,
		_w1052_,
		_w1053_
	);
	LUT2 #(
		.INIT('h8)
	) name280 (
		\g4527_reg/NET0131 ,
		_w1052_,
		_w1054_
	);
	LUT2 #(
		.INIT('h1)
	) name281 (
		_w1053_,
		_w1054_,
		_w1055_
	);
	LUT2 #(
		.INIT('h2)
	) name282 (
		\g35_pad ,
		_w1055_,
		_w1056_
	);
	LUT2 #(
		.INIT('h2)
	) name283 (
		\g4521_reg/NET0131 ,
		_w1056_,
		_w1057_
	);
	LUT2 #(
		.INIT('h4)
	) name284 (
		\g4584_reg/NET0131 ,
		\g4608_reg/NET0131 ,
		_w1058_
	);
	LUT2 #(
		.INIT('h2)
	) name285 (
		\g4593_reg/NET0131 ,
		\g4601_reg/NET0131 ,
		_w1059_
	);
	LUT2 #(
		.INIT('h1)
	) name286 (
		_w1058_,
		_w1059_,
		_w1060_
	);
	LUT2 #(
		.INIT('h2)
	) name287 (
		\g4584_reg/NET0131 ,
		\g4608_reg/NET0131 ,
		_w1061_
	);
	LUT2 #(
		.INIT('h2)
	) name288 (
		\g4593_reg/NET0131 ,
		_w1061_,
		_w1062_
	);
	LUT2 #(
		.INIT('h1)
	) name289 (
		_w1060_,
		_w1062_,
		_w1063_
	);
	LUT2 #(
		.INIT('h4)
	) name290 (
		\g4593_reg/NET0131 ,
		\g4601_reg/NET0131 ,
		_w1064_
	);
	LUT2 #(
		.INIT('h1)
	) name291 (
		\g4616_reg/NET0131 ,
		_w1061_,
		_w1065_
	);
	LUT2 #(
		.INIT('h4)
	) name292 (
		_w1064_,
		_w1065_,
		_w1066_
	);
	LUT2 #(
		.INIT('h8)
	) name293 (
		_w1060_,
		_w1066_,
		_w1067_
	);
	LUT2 #(
		.INIT('h1)
	) name294 (
		_w1063_,
		_w1067_,
		_w1068_
	);
	LUT2 #(
		.INIT('h2)
	) name295 (
		\g35_pad ,
		\g4521_reg/NET0131 ,
		_w1069_
	);
	LUT2 #(
		.INIT('h4)
	) name296 (
		_w1068_,
		_w1069_,
		_w1070_
	);
	LUT2 #(
		.INIT('h1)
	) name297 (
		_w1057_,
		_w1070_,
		_w1071_
	);
	LUT2 #(
		.INIT('h4)
	) name298 (
		\g4521_reg/NET0131 ,
		_w1055_,
		_w1072_
	);
	LUT2 #(
		.INIT('h8)
	) name299 (
		\g4515_reg/NET0131 ,
		\g4521_reg/NET0131 ,
		_w1073_
	);
	LUT2 #(
		.INIT('h1)
	) name300 (
		_w1072_,
		_w1073_,
		_w1074_
	);
	LUT2 #(
		.INIT('h2)
	) name301 (
		\g35_pad ,
		_w1074_,
		_w1075_
	);
	LUT2 #(
		.INIT('h4)
	) name302 (
		\g35_pad ,
		\g4527_reg/NET0131 ,
		_w1076_
	);
	LUT2 #(
		.INIT('h1)
	) name303 (
		_w1075_,
		_w1076_,
		_w1077_
	);
	LUT2 #(
		.INIT('h8)
	) name304 (
		\g35_pad ,
		\g4512_reg/NET0131 ,
		_w1078_
	);
	LUT2 #(
		.INIT('h4)
	) name305 (
		\g4581_reg/NET0131 ,
		_w1078_,
		_w1079_
	);
	LUT2 #(
		.INIT('h8)
	) name306 (
		\g35_pad ,
		\g4572_reg/NET0131 ,
		_w1080_
	);
	LUT2 #(
		.INIT('h8)
	) name307 (
		\g4581_reg/NET0131 ,
		_w1080_,
		_w1081_
	);
	LUT2 #(
		.INIT('h4)
	) name308 (
		\g35_pad ,
		\g4515_reg/NET0131 ,
		_w1082_
	);
	LUT2 #(
		.INIT('h1)
	) name309 (
		_w1079_,
		_w1082_,
		_w1083_
	);
	LUT2 #(
		.INIT('h4)
	) name310 (
		_w1081_,
		_w1083_,
		_w1084_
	);
	LUT2 #(
		.INIT('h8)
	) name311 (
		\g35_pad ,
		\g4581_reg/NET0131 ,
		_w1085_
	);
	LUT2 #(
		.INIT('h2)
	) name312 (
		\g4552_reg/NET0131 ,
		_w1085_,
		_w1086_
	);
	LUT2 #(
		.INIT('h8)
	) name313 (
		\g4575_reg/NET0131 ,
		_w1085_,
		_w1087_
	);
	LUT2 #(
		.INIT('h1)
	) name314 (
		_w1086_,
		_w1087_,
		_w1088_
	);
	LUT2 #(
		.INIT('h1)
	) name315 (
		\g35_pad ,
		\g4512_reg/NET0131 ,
		_w1089_
	);
	LUT2 #(
		.INIT('h8)
	) name316 (
		\g4531_reg/NET0131 ,
		_w1085_,
		_w1090_
	);
	LUT2 #(
		.INIT('h1)
	) name317 (
		_w1089_,
		_w1090_,
		_w1091_
	);
	LUT2 #(
		.INIT('h1)
	) name318 (
		\g1322_reg/NET0131 ,
		\g1333_reg/NET0131 ,
		_w1092_
	);
	LUT2 #(
		.INIT('h8)
	) name319 (
		\g1361_reg/NET0131 ,
		\g1373_reg/NET0131 ,
		_w1093_
	);
	LUT2 #(
		.INIT('h8)
	) name320 (
		\g1351_reg/NET0131 ,
		_w1093_,
		_w1094_
	);
	LUT2 #(
		.INIT('h1)
	) name321 (
		\g1322_reg/NET0131 ,
		\g1339_reg/NET0131 ,
		_w1095_
	);
	LUT2 #(
		.INIT('h8)
	) name322 (
		\g1322_reg/NET0131 ,
		\g1339_reg/NET0131 ,
		_w1096_
	);
	LUT2 #(
		.INIT('h1)
	) name323 (
		_w1095_,
		_w1096_,
		_w1097_
	);
	LUT2 #(
		.INIT('h2)
	) name324 (
		_w1094_,
		_w1097_,
		_w1098_
	);
	LUT2 #(
		.INIT('h2)
	) name325 (
		\g1351_reg/NET0131 ,
		\g1389_reg/NET0131 ,
		_w1099_
	);
	LUT2 #(
		.INIT('h2)
	) name326 (
		_w1097_,
		_w1099_,
		_w1100_
	);
	LUT2 #(
		.INIT('h1)
	) name327 (
		\g1312_reg/NET0131 ,
		_w1100_,
		_w1101_
	);
	LUT2 #(
		.INIT('h4)
	) name328 (
		_w1098_,
		_w1101_,
		_w1102_
	);
	LUT2 #(
		.INIT('h8)
	) name329 (
		\g1345_reg/NET0131 ,
		\g1361_reg/NET0131 ,
		_w1103_
	);
	LUT2 #(
		.INIT('h8)
	) name330 (
		\g1367_reg/NET0131 ,
		_w1103_,
		_w1104_
	);
	LUT2 #(
		.INIT('h2)
	) name331 (
		_w1102_,
		_w1104_,
		_w1105_
	);
	LUT2 #(
		.INIT('h1)
	) name332 (
		_w1092_,
		_w1105_,
		_w1106_
	);
	LUT2 #(
		.INIT('h4)
	) name333 (
		\g1373_reg/NET0131 ,
		_w1101_,
		_w1107_
	);
	LUT2 #(
		.INIT('h2)
	) name334 (
		_w1106_,
		_w1107_,
		_w1108_
	);
	LUT2 #(
		.INIT('h4)
	) name335 (
		\g1379_reg/NET0131 ,
		_w1102_,
		_w1109_
	);
	LUT2 #(
		.INIT('h2)
	) name336 (
		_w1108_,
		_w1109_,
		_w1110_
	);
	LUT2 #(
		.INIT('h1)
	) name337 (
		\g1379_reg/NET0131 ,
		_w1108_,
		_w1111_
	);
	LUT2 #(
		.INIT('h1)
	) name338 (
		_w1110_,
		_w1111_,
		_w1112_
	);
	LUT2 #(
		.INIT('h2)
	) name339 (
		\g35_pad ,
		_w1112_,
		_w1113_
	);
	LUT2 #(
		.INIT('h1)
	) name340 (
		\g1373_reg/NET0131 ,
		\g35_pad ,
		_w1114_
	);
	LUT2 #(
		.INIT('h1)
	) name341 (
		_w1113_,
		_w1114_,
		_w1115_
	);
	LUT2 #(
		.INIT('h4)
	) name342 (
		\g1514_reg/NET0131 ,
		\g1526_reg/NET0131 ,
		_w1116_
	);
	LUT2 #(
		.INIT('h2)
	) name343 (
		\g1536_reg/NET0131 ,
		_w1116_,
		_w1117_
	);
	LUT2 #(
		.INIT('h8)
	) name344 (
		\g1339_reg/NET0131 ,
		\g1521_reg/NET0131 ,
		_w1118_
	);
	LUT2 #(
		.INIT('h4)
	) name345 (
		\g1532_reg/NET0131 ,
		_w1118_,
		_w1119_
	);
	LUT2 #(
		.INIT('h8)
	) name346 (
		\g1345_reg/NET0131 ,
		\g1367_reg/NET0131 ,
		_w1120_
	);
	LUT2 #(
		.INIT('h8)
	) name347 (
		\g1379_reg/NET0131 ,
		_w1120_,
		_w1121_
	);
	LUT2 #(
		.INIT('h1)
	) name348 (
		_w1092_,
		_w1097_,
		_w1122_
	);
	LUT2 #(
		.INIT('h8)
	) name349 (
		_w1121_,
		_w1122_,
		_w1123_
	);
	LUT2 #(
		.INIT('h2)
	) name350 (
		_w817_,
		_w1123_,
		_w1124_
	);
	LUT2 #(
		.INIT('h8)
	) name351 (
		\g7946_pad ,
		_w1119_,
		_w1125_
	);
	LUT2 #(
		.INIT('h4)
	) name352 (
		_w1124_,
		_w1125_,
		_w1126_
	);
	LUT2 #(
		.INIT('h4)
	) name353 (
		_w1117_,
		_w1126_,
		_w1127_
	);
	LUT2 #(
		.INIT('h1)
	) name354 (
		\g1514_reg/NET0131 ,
		\g1526_reg/NET0131 ,
		_w1128_
	);
	LUT2 #(
		.INIT('h8)
	) name355 (
		\g1514_reg/NET0131 ,
		\g7946_pad ,
		_w1129_
	);
	LUT2 #(
		.INIT('h8)
	) name356 (
		\g1526_reg/NET0131 ,
		_w1129_,
		_w1130_
	);
	LUT2 #(
		.INIT('h1)
	) name357 (
		\g1526_reg/NET0131 ,
		\g7946_pad ,
		_w1131_
	);
	LUT2 #(
		.INIT('h1)
	) name358 (
		_w1130_,
		_w1131_,
		_w1132_
	);
	LUT2 #(
		.INIT('h2)
	) name359 (
		\g35_pad ,
		_w1132_,
		_w1133_
	);
	LUT2 #(
		.INIT('h1)
	) name360 (
		_w1128_,
		_w1133_,
		_w1134_
	);
	LUT2 #(
		.INIT('h1)
	) name361 (
		_w1127_,
		_w1134_,
		_w1135_
	);
	LUT2 #(
		.INIT('h1)
	) name362 (
		\g1514_reg/NET0131 ,
		\g35_pad ,
		_w1136_
	);
	LUT2 #(
		.INIT('h1)
	) name363 (
		_w1135_,
		_w1136_,
		_w1137_
	);
	LUT2 #(
		.INIT('h2)
	) name364 (
		\g1367_reg/NET0131 ,
		\g35_pad ,
		_w1138_
	);
	LUT2 #(
		.INIT('h1)
	) name365 (
		\g1373_reg/NET0131 ,
		_w1106_,
		_w1139_
	);
	LUT2 #(
		.INIT('h2)
	) name366 (
		\g35_pad ,
		_w1108_,
		_w1140_
	);
	LUT2 #(
		.INIT('h4)
	) name367 (
		_w1139_,
		_w1140_,
		_w1141_
	);
	LUT2 #(
		.INIT('h1)
	) name368 (
		_w1138_,
		_w1141_,
		_w1142_
	);
	LUT2 #(
		.INIT('h2)
	) name369 (
		\g4549_reg/NET0131 ,
		_w1085_,
		_w1143_
	);
	LUT2 #(
		.INIT('h1)
	) name370 (
		_w1087_,
		_w1143_,
		_w1144_
	);
	LUT2 #(
		.INIT('h1)
	) name371 (
		\g1514_reg/NET0131 ,
		\g7946_pad ,
		_w1145_
	);
	LUT2 #(
		.INIT('h1)
	) name372 (
		_w1129_,
		_w1145_,
		_w1146_
	);
	LUT2 #(
		.INIT('h1)
	) name373 (
		_w1127_,
		_w1146_,
		_w1147_
	);
	LUT2 #(
		.INIT('h2)
	) name374 (
		\g35_pad ,
		_w1147_,
		_w1148_
	);
	LUT2 #(
		.INIT('h4)
	) name375 (
		_w1092_,
		_w1102_,
		_w1149_
	);
	LUT2 #(
		.INIT('h2)
	) name376 (
		\g1345_reg/NET0131 ,
		\g1367_reg/NET0131 ,
		_w1150_
	);
	LUT2 #(
		.INIT('h8)
	) name377 (
		_w1149_,
		_w1150_,
		_w1151_
	);
	LUT2 #(
		.INIT('h2)
	) name378 (
		\g35_pad ,
		_w1151_,
		_w1152_
	);
	LUT2 #(
		.INIT('h2)
	) name379 (
		\g1361_reg/NET0131 ,
		_w1152_,
		_w1153_
	);
	LUT2 #(
		.INIT('h2)
	) name380 (
		_w1102_,
		_w1103_,
		_w1154_
	);
	LUT2 #(
		.INIT('h1)
	) name381 (
		_w1092_,
		_w1154_,
		_w1155_
	);
	LUT2 #(
		.INIT('h8)
	) name382 (
		\g1367_reg/NET0131 ,
		\g35_pad ,
		_w1156_
	);
	LUT2 #(
		.INIT('h4)
	) name383 (
		_w1155_,
		_w1156_,
		_w1157_
	);
	LUT2 #(
		.INIT('h1)
	) name384 (
		_w1153_,
		_w1157_,
		_w1158_
	);
	LUT2 #(
		.INIT('h8)
	) name385 (
		\g7946_pad ,
		_w1116_,
		_w1159_
	);
	LUT2 #(
		.INIT('h4)
	) name386 (
		_w1119_,
		_w1159_,
		_w1160_
	);
	LUT2 #(
		.INIT('h8)
	) name387 (
		\g1542_reg/NET0131 ,
		_w1160_,
		_w1161_
	);
	LUT2 #(
		.INIT('h2)
	) name388 (
		\g35_pad ,
		_w1161_,
		_w1162_
	);
	LUT2 #(
		.INIT('h4)
	) name389 (
		_w1127_,
		_w1162_,
		_w1163_
	);
	LUT2 #(
		.INIT('h8)
	) name390 (
		\g1413_reg/NET0131 ,
		_w1163_,
		_w1164_
	);
	LUT2 #(
		.INIT('h4)
	) name391 (
		\g1413_reg/NET0131 ,
		_w1160_,
		_w1165_
	);
	LUT2 #(
		.INIT('h2)
	) name392 (
		\g35_pad ,
		_w1165_,
		_w1166_
	);
	LUT2 #(
		.INIT('h2)
	) name393 (
		\g1542_reg/NET0131 ,
		_w1166_,
		_w1167_
	);
	LUT2 #(
		.INIT('h1)
	) name394 (
		_w1164_,
		_w1167_,
		_w1168_
	);
	LUT2 #(
		.INIT('h2)
	) name395 (
		\g1514_reg/NET0131 ,
		\g1526_reg/NET0131 ,
		_w1169_
	);
	LUT2 #(
		.INIT('h8)
	) name396 (
		\g13272_pad ,
		_w1169_,
		_w1170_
	);
	LUT2 #(
		.INIT('h1)
	) name397 (
		\g1442_reg/NET0131 ,
		\g1489_reg/NET0131 ,
		_w1171_
	);
	LUT2 #(
		.INIT('h8)
	) name398 (
		_w1170_,
		_w1171_,
		_w1172_
	);
	LUT2 #(
		.INIT('h1)
	) name399 (
		\g1437_reg/NET0131 ,
		_w1172_,
		_w1173_
	);
	LUT2 #(
		.INIT('h4)
	) name400 (
		\g1319_reg/NET0131 ,
		_w818_,
		_w1174_
	);
	LUT2 #(
		.INIT('h2)
	) name401 (
		\g1478_reg/NET0131 ,
		_w1174_,
		_w1175_
	);
	LUT2 #(
		.INIT('h4)
	) name402 (
		\g1478_reg/NET0131 ,
		_w1174_,
		_w1176_
	);
	LUT2 #(
		.INIT('h2)
	) name403 (
		_w1170_,
		_w1175_,
		_w1177_
	);
	LUT2 #(
		.INIT('h4)
	) name404 (
		_w1176_,
		_w1177_,
		_w1178_
	);
	LUT2 #(
		.INIT('h1)
	) name405 (
		_w1173_,
		_w1178_,
		_w1179_
	);
	LUT2 #(
		.INIT('h2)
	) name406 (
		\g35_pad ,
		_w1179_,
		_w1180_
	);
	LUT2 #(
		.INIT('h1)
	) name407 (
		\g1442_reg/NET0131 ,
		\g35_pad ,
		_w1181_
	);
	LUT2 #(
		.INIT('h1)
	) name408 (
		_w1180_,
		_w1181_,
		_w1182_
	);
	LUT2 #(
		.INIT('h8)
	) name409 (
		\g13272_pad ,
		_w1116_,
		_w1183_
	);
	LUT2 #(
		.INIT('h8)
	) name410 (
		_w1171_,
		_w1183_,
		_w1184_
	);
	LUT2 #(
		.INIT('h1)
	) name411 (
		\g1454_reg/NET0131 ,
		_w1184_,
		_w1185_
	);
	LUT2 #(
		.INIT('h2)
	) name412 (
		\g1448_reg/NET0131 ,
		_w1174_,
		_w1186_
	);
	LUT2 #(
		.INIT('h4)
	) name413 (
		\g1448_reg/NET0131 ,
		_w1174_,
		_w1187_
	);
	LUT2 #(
		.INIT('h2)
	) name414 (
		_w1183_,
		_w1186_,
		_w1188_
	);
	LUT2 #(
		.INIT('h4)
	) name415 (
		_w1187_,
		_w1188_,
		_w1189_
	);
	LUT2 #(
		.INIT('h1)
	) name416 (
		_w1185_,
		_w1189_,
		_w1190_
	);
	LUT2 #(
		.INIT('h2)
	) name417 (
		\g35_pad ,
		_w1190_,
		_w1191_
	);
	LUT2 #(
		.INIT('h1)
	) name418 (
		\g1478_reg/NET0131 ,
		\g35_pad ,
		_w1192_
	);
	LUT2 #(
		.INIT('h1)
	) name419 (
		_w1191_,
		_w1192_,
		_w1193_
	);
	LUT2 #(
		.INIT('h8)
	) name420 (
		\g1514_reg/NET0131 ,
		\g1526_reg/NET0131 ,
		_w1194_
	);
	LUT2 #(
		.INIT('h8)
	) name421 (
		\g13272_pad ,
		_w1194_,
		_w1195_
	);
	LUT2 #(
		.INIT('h8)
	) name422 (
		_w1171_,
		_w1195_,
		_w1196_
	);
	LUT2 #(
		.INIT('h1)
	) name423 (
		\g1467_reg/NET0131 ,
		_w1196_,
		_w1197_
	);
	LUT2 #(
		.INIT('h2)
	) name424 (
		\g1472_reg/NET0131 ,
		_w1174_,
		_w1198_
	);
	LUT2 #(
		.INIT('h4)
	) name425 (
		\g1472_reg/NET0131 ,
		_w1174_,
		_w1199_
	);
	LUT2 #(
		.INIT('h2)
	) name426 (
		_w1195_,
		_w1198_,
		_w1200_
	);
	LUT2 #(
		.INIT('h4)
	) name427 (
		_w1199_,
		_w1200_,
		_w1201_
	);
	LUT2 #(
		.INIT('h1)
	) name428 (
		_w1197_,
		_w1201_,
		_w1202_
	);
	LUT2 #(
		.INIT('h2)
	) name429 (
		\g35_pad ,
		_w1202_,
		_w1203_
	);
	LUT2 #(
		.INIT('h1)
	) name430 (
		\g1448_reg/NET0131 ,
		\g35_pad ,
		_w1204_
	);
	LUT2 #(
		.INIT('h1)
	) name431 (
		_w1203_,
		_w1204_,
		_w1205_
	);
	LUT2 #(
		.INIT('h8)
	) name432 (
		\g13272_pad ,
		_w1128_,
		_w1206_
	);
	LUT2 #(
		.INIT('h8)
	) name433 (
		_w1171_,
		_w1206_,
		_w1207_
	);
	LUT2 #(
		.INIT('h1)
	) name434 (
		\g1484_reg/NET0131 ,
		_w1207_,
		_w1208_
	);
	LUT2 #(
		.INIT('h2)
	) name435 (
		\g1300_reg/NET0131 ,
		_w1174_,
		_w1209_
	);
	LUT2 #(
		.INIT('h4)
	) name436 (
		\g1300_reg/NET0131 ,
		_w1174_,
		_w1210_
	);
	LUT2 #(
		.INIT('h2)
	) name437 (
		_w1206_,
		_w1209_,
		_w1211_
	);
	LUT2 #(
		.INIT('h4)
	) name438 (
		_w1210_,
		_w1211_,
		_w1212_
	);
	LUT2 #(
		.INIT('h1)
	) name439 (
		_w1208_,
		_w1212_,
		_w1213_
	);
	LUT2 #(
		.INIT('h2)
	) name440 (
		\g35_pad ,
		_w1213_,
		_w1214_
	);
	LUT2 #(
		.INIT('h1)
	) name441 (
		\g1472_reg/NET0131 ,
		\g35_pad ,
		_w1215_
	);
	LUT2 #(
		.INIT('h1)
	) name442 (
		_w1214_,
		_w1215_,
		_w1216_
	);
	LUT2 #(
		.INIT('h2)
	) name443 (
		\g4504_reg/NET0131 ,
		_w1085_,
		_w1217_
	);
	LUT2 #(
		.INIT('h1)
	) name444 (
		_w1081_,
		_w1217_,
		_w1218_
	);
	LUT2 #(
		.INIT('h4)
	) name445 (
		\g1345_reg/NET0131 ,
		_w1102_,
		_w1219_
	);
	LUT2 #(
		.INIT('h1)
	) name446 (
		_w1092_,
		_w1219_,
		_w1220_
	);
	LUT2 #(
		.INIT('h2)
	) name447 (
		\g35_pad ,
		_w1220_,
		_w1221_
	);
	LUT2 #(
		.INIT('h8)
	) name448 (
		\g1361_reg/NET0131 ,
		_w1221_,
		_w1222_
	);
	LUT2 #(
		.INIT('h4)
	) name449 (
		\g1361_reg/NET0131 ,
		_w1149_,
		_w1223_
	);
	LUT2 #(
		.INIT('h2)
	) name450 (
		\g35_pad ,
		_w1223_,
		_w1224_
	);
	LUT2 #(
		.INIT('h2)
	) name451 (
		\g1345_reg/NET0131 ,
		_w1224_,
		_w1225_
	);
	LUT2 #(
		.INIT('h1)
	) name452 (
		_w1222_,
		_w1225_,
		_w1226_
	);
	LUT2 #(
		.INIT('h1)
	) name453 (
		\g1532_reg/NET0131 ,
		\g35_pad ,
		_w1227_
	);
	LUT2 #(
		.INIT('h1)
	) name454 (
		\g1536_reg/NET0131 ,
		_w1126_,
		_w1228_
	);
	LUT2 #(
		.INIT('h8)
	) name455 (
		\g1413_reg/NET0131 ,
		\g1536_reg/NET0131 ,
		_w1229_
	);
	LUT2 #(
		.INIT('h8)
	) name456 (
		_w1161_,
		_w1229_,
		_w1230_
	);
	LUT2 #(
		.INIT('h1)
	) name457 (
		_w1228_,
		_w1230_,
		_w1231_
	);
	LUT2 #(
		.INIT('h2)
	) name458 (
		\g35_pad ,
		_w1231_,
		_w1232_
	);
	LUT2 #(
		.INIT('h1)
	) name459 (
		_w1227_,
		_w1232_,
		_w1233_
	);
	LUT2 #(
		.INIT('h2)
	) name460 (
		\g1536_reg/NET0131 ,
		\g35_pad ,
		_w1234_
	);
	LUT2 #(
		.INIT('h1)
	) name461 (
		\g1542_reg/NET0131 ,
		_w1160_,
		_w1235_
	);
	LUT2 #(
		.INIT('h2)
	) name462 (
		_w1163_,
		_w1235_,
		_w1236_
	);
	LUT2 #(
		.INIT('h1)
	) name463 (
		_w1234_,
		_w1236_,
		_w1237_
	);
	LUT2 #(
		.INIT('h4)
	) name464 (
		\g333_reg/NET0131 ,
		\g351_reg/NET0131 ,
		_w1238_
	);
	LUT2 #(
		.INIT('h2)
	) name465 (
		\g35_pad ,
		_w1238_,
		_w1239_
	);
	LUT2 #(
		.INIT('h1)
	) name466 (
		\g355_reg/NET0131 ,
		_w1239_,
		_w1240_
	);
	LUT2 #(
		.INIT('h1)
	) name467 (
		\g29211_pad ,
		\g351_reg/NET0131 ,
		_w1241_
	);
	LUT2 #(
		.INIT('h8)
	) name468 (
		\g35_pad ,
		_w1241_,
		_w1242_
	);
	LUT2 #(
		.INIT('h1)
	) name469 (
		_w1240_,
		_w1242_,
		_w1243_
	);
	LUT2 #(
		.INIT('h8)
	) name470 (
		\g1389_reg/NET0131 ,
		_w1097_,
		_w1244_
	);
	LUT2 #(
		.INIT('h2)
	) name471 (
		_w1094_,
		_w1244_,
		_w1245_
	);
	LUT2 #(
		.INIT('h1)
	) name472 (
		\g1351_reg/NET0131 ,
		_w1097_,
		_w1246_
	);
	LUT2 #(
		.INIT('h8)
	) name473 (
		_w1121_,
		_w1246_,
		_w1247_
	);
	LUT2 #(
		.INIT('h1)
	) name474 (
		_w1245_,
		_w1247_,
		_w1248_
	);
	LUT2 #(
		.INIT('h1)
	) name475 (
		_w1092_,
		_w1248_,
		_w1249_
	);
	LUT2 #(
		.INIT('h4)
	) name476 (
		_w1092_,
		_w1097_,
		_w1250_
	);
	LUT2 #(
		.INIT('h2)
	) name477 (
		\g1312_reg/NET0131 ,
		_w1250_,
		_w1251_
	);
	LUT2 #(
		.INIT('h1)
	) name478 (
		_w1249_,
		_w1251_,
		_w1252_
	);
	LUT2 #(
		.INIT('h2)
	) name479 (
		\g35_pad ,
		_w1252_,
		_w1253_
	);
	LUT2 #(
		.INIT('h2)
	) name480 (
		\g35_pad ,
		_w1250_,
		_w1254_
	);
	LUT2 #(
		.INIT('h2)
	) name481 (
		\g1312_reg/NET0131 ,
		_w1254_,
		_w1255_
	);
	LUT2 #(
		.INIT('h1)
	) name482 (
		_w1093_,
		_w1244_,
		_w1256_
	);
	LUT2 #(
		.INIT('h1)
	) name483 (
		_w1092_,
		_w1256_,
		_w1257_
	);
	LUT2 #(
		.INIT('h8)
	) name484 (
		\g1351_reg/NET0131 ,
		\g35_pad ,
		_w1258_
	);
	LUT2 #(
		.INIT('h4)
	) name485 (
		_w1257_,
		_w1258_,
		_w1259_
	);
	LUT2 #(
		.INIT('h1)
	) name486 (
		_w1255_,
		_w1259_,
		_w1260_
	);
	LUT2 #(
		.INIT('h1)
	) name487 (
		\g333_reg/NET0131 ,
		\g355_reg/NET0131 ,
		_w1261_
	);
	LUT2 #(
		.INIT('h2)
	) name488 (
		\g35_pad ,
		_w1261_,
		_w1262_
	);
	LUT2 #(
		.INIT('h1)
	) name489 (
		\g351_reg/NET0131 ,
		_w1262_,
		_w1263_
	);
	LUT2 #(
		.INIT('h8)
	) name490 (
		\g351_reg/NET0131 ,
		\g35_pad ,
		_w1264_
	);
	LUT2 #(
		.INIT('h1)
	) name491 (
		_w1263_,
		_w1264_,
		_w1265_
	);
	LUT2 #(
		.INIT('h1)
	) name492 (
		\g4546_reg/NET0131 ,
		_w1085_,
		_w1266_
	);
	LUT2 #(
		.INIT('h8)
	) name493 (
		_w817_,
		_w1250_,
		_w1267_
	);
	LUT2 #(
		.INIT('h2)
	) name494 (
		\g1322_reg/NET0131 ,
		\g1579_reg/NET0131 ,
		_w1268_
	);
	LUT2 #(
		.INIT('h4)
	) name495 (
		\g1322_reg/NET0131 ,
		\g1579_reg/NET0131 ,
		_w1269_
	);
	LUT2 #(
		.INIT('h1)
	) name496 (
		_w1268_,
		_w1269_,
		_w1270_
	);
	LUT2 #(
		.INIT('h2)
	) name497 (
		_w1267_,
		_w1270_,
		_w1271_
	);
	LUT2 #(
		.INIT('h1)
	) name498 (
		\g1333_reg/NET0131 ,
		\g19357_pad ,
		_w1272_
	);
	LUT2 #(
		.INIT('h4)
	) name499 (
		\g7946_pad ,
		_w1272_,
		_w1273_
	);
	LUT2 #(
		.INIT('h1)
	) name500 (
		\g13272_pad ,
		\g8475_pad ,
		_w1274_
	);
	LUT2 #(
		.INIT('h8)
	) name501 (
		_w1273_,
		_w1274_,
		_w1275_
	);
	LUT2 #(
		.INIT('h2)
	) name502 (
		_w1271_,
		_w1275_,
		_w1276_
	);
	LUT2 #(
		.INIT('h4)
	) name503 (
		_w1271_,
		_w1275_,
		_w1277_
	);
	LUT2 #(
		.INIT('h1)
	) name504 (
		_w1276_,
		_w1277_,
		_w1278_
	);
	LUT2 #(
		.INIT('h2)
	) name505 (
		\g35_pad ,
		_w1278_,
		_w1279_
	);
	LUT2 #(
		.INIT('h2)
	) name506 (
		\g1339_reg/NET0131 ,
		\g35_pad ,
		_w1280_
	);
	LUT2 #(
		.INIT('h1)
	) name507 (
		_w1279_,
		_w1280_,
		_w1281_
	);
	LUT2 #(
		.INIT('h8)
	) name508 (
		\g35_pad ,
		_w1271_,
		_w1282_
	);
	LUT2 #(
		.INIT('h1)
	) name509 (
		\g1333_reg/NET0131 ,
		_w1282_,
		_w1283_
	);
	LUT2 #(
		.INIT('h8)
	) name510 (
		\g1333_reg/NET0131 ,
		_w1282_,
		_w1284_
	);
	LUT2 #(
		.INIT('h1)
	) name511 (
		_w1283_,
		_w1284_,
		_w1285_
	);
	LUT2 #(
		.INIT('h2)
	) name512 (
		\g1351_reg/NET0131 ,
		\g35_pad ,
		_w1286_
	);
	LUT2 #(
		.INIT('h4)
	) name513 (
		\g1345_reg/NET0131 ,
		_w1092_,
		_w1287_
	);
	LUT2 #(
		.INIT('h2)
	) name514 (
		_w1221_,
		_w1287_,
		_w1288_
	);
	LUT2 #(
		.INIT('h1)
	) name515 (
		_w1286_,
		_w1288_,
		_w1289_
	);
	LUT2 #(
		.INIT('h2)
	) name516 (
		\g4375_reg/NET0131 ,
		\g4382_reg/NET0131 ,
		_w1290_
	);
	LUT2 #(
		.INIT('h4)
	) name517 (
		\g4375_reg/NET0131 ,
		\g4382_reg/NET0131 ,
		_w1291_
	);
	LUT2 #(
		.INIT('h1)
	) name518 (
		_w1290_,
		_w1291_,
		_w1292_
	);
	LUT2 #(
		.INIT('h1)
	) name519 (
		\g4375_reg/NET0131 ,
		\g4405_reg/NET0131 ,
		_w1293_
	);
	LUT2 #(
		.INIT('h1)
	) name520 (
		\g4411_reg/NET0131 ,
		\g7243_pad ,
		_w1294_
	);
	LUT2 #(
		.INIT('h4)
	) name521 (
		\g7257_pad ,
		_w1294_,
		_w1295_
	);
	LUT2 #(
		.INIT('h8)
	) name522 (
		_w1293_,
		_w1295_,
		_w1296_
	);
	LUT2 #(
		.INIT('h2)
	) name523 (
		\g35_pad ,
		_w1292_,
		_w1297_
	);
	LUT2 #(
		.INIT('h4)
	) name524 (
		_w1296_,
		_w1297_,
		_w1298_
	);
	LUT2 #(
		.INIT('h2)
	) name525 (
		\g35_pad ,
		\g4392_reg/NET0131 ,
		_w1299_
	);
	LUT2 #(
		.INIT('h8)
	) name526 (
		_w1296_,
		_w1299_,
		_w1300_
	);
	LUT2 #(
		.INIT('h4)
	) name527 (
		\g4417_reg/NET0131 ,
		_w1300_,
		_w1301_
	);
	LUT2 #(
		.INIT('h4)
	) name528 (
		\g35_pad ,
		\g4388_reg/NET0131 ,
		_w1302_
	);
	LUT2 #(
		.INIT('h1)
	) name529 (
		_w1298_,
		_w1302_,
		_w1303_
	);
	LUT2 #(
		.INIT('h4)
	) name530 (
		_w1301_,
		_w1303_,
		_w1304_
	);
	LUT2 #(
		.INIT('h2)
	) name531 (
		\g1171_reg/NET0131 ,
		\g1183_reg/NET0131 ,
		_w1305_
	);
	LUT2 #(
		.INIT('h8)
	) name532 (
		\g13259_pad ,
		_w1305_,
		_w1306_
	);
	LUT2 #(
		.INIT('h1)
	) name533 (
		\g1099_reg/NET0131 ,
		\g1146_reg/NET0131 ,
		_w1307_
	);
	LUT2 #(
		.INIT('h8)
	) name534 (
		_w1306_,
		_w1307_,
		_w1308_
	);
	LUT2 #(
		.INIT('h1)
	) name535 (
		\g1094_reg/NET0131 ,
		_w1308_,
		_w1309_
	);
	LUT2 #(
		.INIT('h4)
	) name536 (
		\g976_reg/NET0131 ,
		_w816_,
		_w1310_
	);
	LUT2 #(
		.INIT('h2)
	) name537 (
		\g1135_reg/NET0131 ,
		_w1310_,
		_w1311_
	);
	LUT2 #(
		.INIT('h4)
	) name538 (
		\g1135_reg/NET0131 ,
		_w1310_,
		_w1312_
	);
	LUT2 #(
		.INIT('h2)
	) name539 (
		_w1306_,
		_w1311_,
		_w1313_
	);
	LUT2 #(
		.INIT('h4)
	) name540 (
		_w1312_,
		_w1313_,
		_w1314_
	);
	LUT2 #(
		.INIT('h1)
	) name541 (
		_w1309_,
		_w1314_,
		_w1315_
	);
	LUT2 #(
		.INIT('h2)
	) name542 (
		\g35_pad ,
		_w1315_,
		_w1316_
	);
	LUT2 #(
		.INIT('h1)
	) name543 (
		\g1099_reg/NET0131 ,
		\g35_pad ,
		_w1317_
	);
	LUT2 #(
		.INIT('h1)
	) name544 (
		_w1316_,
		_w1317_,
		_w1318_
	);
	LUT2 #(
		.INIT('h4)
	) name545 (
		\g1171_reg/NET0131 ,
		\g1183_reg/NET0131 ,
		_w1319_
	);
	LUT2 #(
		.INIT('h8)
	) name546 (
		\g13259_pad ,
		_w1319_,
		_w1320_
	);
	LUT2 #(
		.INIT('h8)
	) name547 (
		_w1307_,
		_w1320_,
		_w1321_
	);
	LUT2 #(
		.INIT('h1)
	) name548 (
		\g1111_reg/NET0131 ,
		_w1321_,
		_w1322_
	);
	LUT2 #(
		.INIT('h2)
	) name549 (
		\g1105_reg/NET0131 ,
		_w1310_,
		_w1323_
	);
	LUT2 #(
		.INIT('h4)
	) name550 (
		\g1105_reg/NET0131 ,
		_w1310_,
		_w1324_
	);
	LUT2 #(
		.INIT('h2)
	) name551 (
		_w1320_,
		_w1323_,
		_w1325_
	);
	LUT2 #(
		.INIT('h4)
	) name552 (
		_w1324_,
		_w1325_,
		_w1326_
	);
	LUT2 #(
		.INIT('h1)
	) name553 (
		_w1322_,
		_w1326_,
		_w1327_
	);
	LUT2 #(
		.INIT('h2)
	) name554 (
		\g35_pad ,
		_w1327_,
		_w1328_
	);
	LUT2 #(
		.INIT('h1)
	) name555 (
		\g1135_reg/NET0131 ,
		\g35_pad ,
		_w1329_
	);
	LUT2 #(
		.INIT('h1)
	) name556 (
		_w1328_,
		_w1329_,
		_w1330_
	);
	LUT2 #(
		.INIT('h8)
	) name557 (
		\g1171_reg/NET0131 ,
		\g1183_reg/NET0131 ,
		_w1331_
	);
	LUT2 #(
		.INIT('h8)
	) name558 (
		\g13259_pad ,
		_w1331_,
		_w1332_
	);
	LUT2 #(
		.INIT('h8)
	) name559 (
		_w1307_,
		_w1332_,
		_w1333_
	);
	LUT2 #(
		.INIT('h1)
	) name560 (
		\g1124_reg/NET0131 ,
		_w1333_,
		_w1334_
	);
	LUT2 #(
		.INIT('h2)
	) name561 (
		\g1129_reg/NET0131 ,
		_w1310_,
		_w1335_
	);
	LUT2 #(
		.INIT('h4)
	) name562 (
		\g1129_reg/NET0131 ,
		_w1310_,
		_w1336_
	);
	LUT2 #(
		.INIT('h2)
	) name563 (
		_w1332_,
		_w1335_,
		_w1337_
	);
	LUT2 #(
		.INIT('h4)
	) name564 (
		_w1336_,
		_w1337_,
		_w1338_
	);
	LUT2 #(
		.INIT('h1)
	) name565 (
		_w1334_,
		_w1338_,
		_w1339_
	);
	LUT2 #(
		.INIT('h2)
	) name566 (
		\g35_pad ,
		_w1339_,
		_w1340_
	);
	LUT2 #(
		.INIT('h1)
	) name567 (
		\g1105_reg/NET0131 ,
		\g35_pad ,
		_w1341_
	);
	LUT2 #(
		.INIT('h1)
	) name568 (
		_w1340_,
		_w1341_,
		_w1342_
	);
	LUT2 #(
		.INIT('h1)
	) name569 (
		\g1171_reg/NET0131 ,
		\g1183_reg/NET0131 ,
		_w1343_
	);
	LUT2 #(
		.INIT('h8)
	) name570 (
		\g13259_pad ,
		_w1343_,
		_w1344_
	);
	LUT2 #(
		.INIT('h8)
	) name571 (
		_w1307_,
		_w1344_,
		_w1345_
	);
	LUT2 #(
		.INIT('h1)
	) name572 (
		\g1141_reg/NET0131 ,
		_w1345_,
		_w1346_
	);
	LUT2 #(
		.INIT('h2)
	) name573 (
		\g956_reg/NET0131 ,
		_w1310_,
		_w1347_
	);
	LUT2 #(
		.INIT('h4)
	) name574 (
		\g956_reg/NET0131 ,
		_w1310_,
		_w1348_
	);
	LUT2 #(
		.INIT('h2)
	) name575 (
		_w1344_,
		_w1347_,
		_w1349_
	);
	LUT2 #(
		.INIT('h4)
	) name576 (
		_w1348_,
		_w1349_,
		_w1350_
	);
	LUT2 #(
		.INIT('h1)
	) name577 (
		_w1346_,
		_w1350_,
		_w1351_
	);
	LUT2 #(
		.INIT('h2)
	) name578 (
		\g35_pad ,
		_w1351_,
		_w1352_
	);
	LUT2 #(
		.INIT('h1)
	) name579 (
		\g1129_reg/NET0131 ,
		\g35_pad ,
		_w1353_
	);
	LUT2 #(
		.INIT('h1)
	) name580 (
		_w1352_,
		_w1353_,
		_w1354_
	);
	LUT2 #(
		.INIT('h1)
	) name581 (
		\g4501_reg/NET0131 ,
		_w1085_,
		_w1355_
	);
	LUT2 #(
		.INIT('h8)
	) name582 (
		\g4392_reg/NET0131 ,
		_w1296_,
		_w1356_
	);
	LUT2 #(
		.INIT('h2)
	) name583 (
		\g35_pad ,
		_w1356_,
		_w1357_
	);
	LUT2 #(
		.INIT('h2)
	) name584 (
		\g4401_reg/NET0131 ,
		_w1357_,
		_w1358_
	);
	LUT2 #(
		.INIT('h8)
	) name585 (
		\g35_pad ,
		\g4411_reg/NET0131 ,
		_w1359_
	);
	LUT2 #(
		.INIT('h1)
	) name586 (
		_w1358_,
		_w1359_,
		_w1360_
	);
	LUT2 #(
		.INIT('h8)
	) name587 (
		\g4388_reg/NET0131 ,
		_w1300_,
		_w1361_
	);
	LUT2 #(
		.INIT('h1)
	) name588 (
		\g4405_reg/NET0131 ,
		_w1361_,
		_w1362_
	);
	LUT2 #(
		.INIT('h2)
	) name589 (
		\g35_pad ,
		\g4382_reg/NET0131 ,
		_w1363_
	);
	LUT2 #(
		.INIT('h2)
	) name590 (
		\g4375_reg/NET0131 ,
		_w1363_,
		_w1364_
	);
	LUT2 #(
		.INIT('h8)
	) name591 (
		\g35_pad ,
		\g4392_reg/NET0131 ,
		_w1365_
	);
	LUT2 #(
		.INIT('h8)
	) name592 (
		_w1296_,
		_w1365_,
		_w1366_
	);
	LUT2 #(
		.INIT('h1)
	) name593 (
		_w1364_,
		_w1366_,
		_w1367_
	);
	LUT2 #(
		.INIT('h4)
	) name594 (
		\g35_pad ,
		\g4455_reg/NET0131 ,
		_w1368_
	);
	LUT2 #(
		.INIT('h4)
	) name595 (
		_w1296_,
		_w1365_,
		_w1369_
	);
	LUT2 #(
		.INIT('h1)
	) name596 (
		_w1301_,
		_w1369_,
		_w1370_
	);
	LUT2 #(
		.INIT('h4)
	) name597 (
		_w1368_,
		_w1370_,
		_w1371_
	);
	LUT2 #(
		.INIT('h8)
	) name598 (
		_w1099_,
		_w1250_,
		_w1372_
	);
	LUT2 #(
		.INIT('h2)
	) name599 (
		\g35_pad ,
		_w1372_,
		_w1373_
	);
	LUT2 #(
		.INIT('h2)
	) name600 (
		\g1384_reg/NET0131 ,
		_w1373_,
		_w1374_
	);
	LUT2 #(
		.INIT('h2)
	) name601 (
		\g1351_reg/NET0131 ,
		\g1384_reg/NET0131 ,
		_w1375_
	);
	LUT2 #(
		.INIT('h2)
	) name602 (
		_w1250_,
		_w1375_,
		_w1376_
	);
	LUT2 #(
		.INIT('h2)
	) name603 (
		\g35_pad ,
		_w1376_,
		_w1377_
	);
	LUT2 #(
		.INIT('h8)
	) name604 (
		\g1389_reg/NET0131 ,
		_w1377_,
		_w1378_
	);
	LUT2 #(
		.INIT('h1)
	) name605 (
		_w1374_,
		_w1378_,
		_w1379_
	);
	LUT2 #(
		.INIT('h8)
	) name606 (
		\g1430_reg/NET0131 ,
		\g1548_reg/NET0131 ,
		_w1380_
	);
	LUT2 #(
		.INIT('h8)
	) name607 (
		\g1564_reg/NET0131 ,
		_w1380_,
		_w1381_
	);
	LUT2 #(
		.INIT('h8)
	) name608 (
		\g1554_reg/NET0131 ,
		_w1381_,
		_w1382_
	);
	LUT2 #(
		.INIT('h4)
	) name609 (
		_w1267_,
		_w1382_,
		_w1383_
	);
	LUT2 #(
		.INIT('h1)
	) name610 (
		\g17320_pad ,
		\g17404_pad ,
		_w1384_
	);
	LUT2 #(
		.INIT('h4)
	) name611 (
		\g17423_pad ,
		\g35_pad ,
		_w1385_
	);
	LUT2 #(
		.INIT('h8)
	) name612 (
		_w1384_,
		_w1385_,
		_w1386_
	);
	LUT2 #(
		.INIT('h4)
	) name613 (
		_w1383_,
		_w1386_,
		_w1387_
	);
	LUT2 #(
		.INIT('h4)
	) name614 (
		\g209_reg/NET0131 ,
		\g691_reg/NET0131 ,
		_w1388_
	);
	LUT2 #(
		.INIT('h8)
	) name615 (
		_w818_,
		_w1388_,
		_w1389_
	);
	LUT2 #(
		.INIT('h4)
	) name616 (
		\g1478_reg/NET0131 ,
		_w1389_,
		_w1390_
	);
	LUT2 #(
		.INIT('h8)
	) name617 (
		\g1322_reg/NET0131 ,
		\g1404_reg/NET0131 ,
		_w1391_
	);
	LUT2 #(
		.INIT('h1)
	) name618 (
		\g1548_reg/NET0131 ,
		\g1554_reg/NET0131 ,
		_w1392_
	);
	LUT2 #(
		.INIT('h1)
	) name619 (
		\g1559_reg/NET0131 ,
		\g1564_reg/NET0131 ,
		_w1393_
	);
	LUT2 #(
		.INIT('h8)
	) name620 (
		_w1392_,
		_w1393_,
		_w1394_
	);
	LUT2 #(
		.INIT('h8)
	) name621 (
		_w1391_,
		_w1394_,
		_w1395_
	);
	LUT2 #(
		.INIT('h8)
	) name622 (
		_w1169_,
		_w1395_,
		_w1396_
	);
	LUT2 #(
		.INIT('h2)
	) name623 (
		\g17320_pad ,
		_w1396_,
		_w1397_
	);
	LUT2 #(
		.INIT('h2)
	) name624 (
		_w1390_,
		_w1397_,
		_w1398_
	);
	LUT2 #(
		.INIT('h8)
	) name625 (
		\g35_pad ,
		_w1398_,
		_w1399_
	);
	LUT2 #(
		.INIT('h8)
	) name626 (
		\g2241_reg/NET0131 ,
		_w1399_,
		_w1400_
	);
	LUT2 #(
		.INIT('h2)
	) name627 (
		\g2227_reg/NET0131 ,
		\g35_pad ,
		_w1401_
	);
	LUT2 #(
		.INIT('h1)
	) name628 (
		\g2153_reg/NET0131 ,
		\g2227_reg/NET0131 ,
		_w1402_
	);
	LUT2 #(
		.INIT('h2)
	) name629 (
		\g2241_reg/NET0131 ,
		_w1402_,
		_w1403_
	);
	LUT2 #(
		.INIT('h4)
	) name630 (
		\g1589_reg/NET0131 ,
		_w1390_,
		_w1404_
	);
	LUT2 #(
		.INIT('h4)
	) name631 (
		_w1403_,
		_w1404_,
		_w1405_
	);
	LUT2 #(
		.INIT('h2)
	) name632 (
		_w1403_,
		_w1404_,
		_w1406_
	);
	LUT2 #(
		.INIT('h2)
	) name633 (
		\g35_pad ,
		_w1398_,
		_w1407_
	);
	LUT2 #(
		.INIT('h1)
	) name634 (
		_w1405_,
		_w1406_,
		_w1408_
	);
	LUT2 #(
		.INIT('h8)
	) name635 (
		_w1407_,
		_w1408_,
		_w1409_
	);
	LUT2 #(
		.INIT('h1)
	) name636 (
		_w1400_,
		_w1401_,
		_w1410_
	);
	LUT2 #(
		.INIT('h4)
	) name637 (
		_w1409_,
		_w1410_,
		_w1411_
	);
	LUT2 #(
		.INIT('h4)
	) name638 (
		\g1448_reg/NET0131 ,
		_w1389_,
		_w1412_
	);
	LUT2 #(
		.INIT('h8)
	) name639 (
		_w1116_,
		_w1395_,
		_w1413_
	);
	LUT2 #(
		.INIT('h2)
	) name640 (
		\g17404_pad ,
		_w1413_,
		_w1414_
	);
	LUT2 #(
		.INIT('h2)
	) name641 (
		_w1412_,
		_w1414_,
		_w1415_
	);
	LUT2 #(
		.INIT('h8)
	) name642 (
		\g35_pad ,
		_w1415_,
		_w1416_
	);
	LUT2 #(
		.INIT('h8)
	) name643 (
		\g2375_reg/NET0131 ,
		_w1416_,
		_w1417_
	);
	LUT2 #(
		.INIT('h2)
	) name644 (
		\g2361_reg/NET0131 ,
		\g35_pad ,
		_w1418_
	);
	LUT2 #(
		.INIT('h1)
	) name645 (
		\g2287_reg/NET0131 ,
		\g2361_reg/NET0131 ,
		_w1419_
	);
	LUT2 #(
		.INIT('h2)
	) name646 (
		\g2375_reg/NET0131 ,
		_w1419_,
		_w1420_
	);
	LUT2 #(
		.INIT('h8)
	) name647 (
		\g1589_reg/NET0131 ,
		_w1412_,
		_w1421_
	);
	LUT2 #(
		.INIT('h4)
	) name648 (
		_w1420_,
		_w1421_,
		_w1422_
	);
	LUT2 #(
		.INIT('h2)
	) name649 (
		_w1420_,
		_w1421_,
		_w1423_
	);
	LUT2 #(
		.INIT('h2)
	) name650 (
		\g35_pad ,
		_w1415_,
		_w1424_
	);
	LUT2 #(
		.INIT('h1)
	) name651 (
		_w1422_,
		_w1423_,
		_w1425_
	);
	LUT2 #(
		.INIT('h8)
	) name652 (
		_w1424_,
		_w1425_,
		_w1426_
	);
	LUT2 #(
		.INIT('h1)
	) name653 (
		_w1417_,
		_w1418_,
		_w1427_
	);
	LUT2 #(
		.INIT('h4)
	) name654 (
		_w1426_,
		_w1427_,
		_w1428_
	);
	LUT2 #(
		.INIT('h4)
	) name655 (
		\g1472_reg/NET0131 ,
		_w1389_,
		_w1429_
	);
	LUT2 #(
		.INIT('h8)
	) name656 (
		_w1194_,
		_w1395_,
		_w1430_
	);
	LUT2 #(
		.INIT('h2)
	) name657 (
		\g17423_pad ,
		_w1430_,
		_w1431_
	);
	LUT2 #(
		.INIT('h2)
	) name658 (
		_w1429_,
		_w1431_,
		_w1432_
	);
	LUT2 #(
		.INIT('h8)
	) name659 (
		\g35_pad ,
		_w1432_,
		_w1433_
	);
	LUT2 #(
		.INIT('h8)
	) name660 (
		\g2509_reg/NET0131 ,
		_w1433_,
		_w1434_
	);
	LUT2 #(
		.INIT('h2)
	) name661 (
		\g2495_reg/NET0131 ,
		\g35_pad ,
		_w1435_
	);
	LUT2 #(
		.INIT('h1)
	) name662 (
		\g2421_reg/NET0131 ,
		\g2495_reg/NET0131 ,
		_w1436_
	);
	LUT2 #(
		.INIT('h2)
	) name663 (
		\g2509_reg/NET0131 ,
		_w1436_,
		_w1437_
	);
	LUT2 #(
		.INIT('h4)
	) name664 (
		\g1589_reg/NET0131 ,
		_w1429_,
		_w1438_
	);
	LUT2 #(
		.INIT('h4)
	) name665 (
		_w1437_,
		_w1438_,
		_w1439_
	);
	LUT2 #(
		.INIT('h2)
	) name666 (
		_w1437_,
		_w1438_,
		_w1440_
	);
	LUT2 #(
		.INIT('h2)
	) name667 (
		\g35_pad ,
		_w1432_,
		_w1441_
	);
	LUT2 #(
		.INIT('h1)
	) name668 (
		_w1439_,
		_w1440_,
		_w1442_
	);
	LUT2 #(
		.INIT('h8)
	) name669 (
		_w1441_,
		_w1442_,
		_w1443_
	);
	LUT2 #(
		.INIT('h1)
	) name670 (
		_w1434_,
		_w1435_,
		_w1444_
	);
	LUT2 #(
		.INIT('h4)
	) name671 (
		_w1443_,
		_w1444_,
		_w1445_
	);
	LUT2 #(
		.INIT('h4)
	) name672 (
		\g1300_reg/NET0131 ,
		_w1389_,
		_w1446_
	);
	LUT2 #(
		.INIT('h8)
	) name673 (
		_w1128_,
		_w1395_,
		_w1447_
	);
	LUT2 #(
		.INIT('h2)
	) name674 (
		\g1430_reg/NET0131 ,
		_w1447_,
		_w1448_
	);
	LUT2 #(
		.INIT('h2)
	) name675 (
		_w1446_,
		_w1448_,
		_w1449_
	);
	LUT2 #(
		.INIT('h8)
	) name676 (
		\g35_pad ,
		_w1449_,
		_w1450_
	);
	LUT2 #(
		.INIT('h8)
	) name677 (
		\g2643_reg/NET0131 ,
		_w1450_,
		_w1451_
	);
	LUT2 #(
		.INIT('h2)
	) name678 (
		\g2629_reg/NET0131 ,
		\g35_pad ,
		_w1452_
	);
	LUT2 #(
		.INIT('h1)
	) name679 (
		\g2555_reg/NET0131 ,
		\g2629_reg/NET0131 ,
		_w1453_
	);
	LUT2 #(
		.INIT('h2)
	) name680 (
		\g2643_reg/NET0131 ,
		_w1453_,
		_w1454_
	);
	LUT2 #(
		.INIT('h8)
	) name681 (
		\g1589_reg/NET0131 ,
		_w1446_,
		_w1455_
	);
	LUT2 #(
		.INIT('h4)
	) name682 (
		_w1454_,
		_w1455_,
		_w1456_
	);
	LUT2 #(
		.INIT('h2)
	) name683 (
		_w1454_,
		_w1455_,
		_w1457_
	);
	LUT2 #(
		.INIT('h2)
	) name684 (
		\g35_pad ,
		_w1449_,
		_w1458_
	);
	LUT2 #(
		.INIT('h1)
	) name685 (
		_w1456_,
		_w1457_,
		_w1459_
	);
	LUT2 #(
		.INIT('h8)
	) name686 (
		_w1458_,
		_w1459_,
		_w1460_
	);
	LUT2 #(
		.INIT('h1)
	) name687 (
		_w1451_,
		_w1452_,
		_w1461_
	);
	LUT2 #(
		.INIT('h4)
	) name688 (
		_w1460_,
		_w1461_,
		_w1462_
	);
	LUT2 #(
		.INIT('h4)
	) name689 (
		\g35_pad ,
		\g4417_reg/NET0131 ,
		_w1463_
	);
	LUT2 #(
		.INIT('h2)
	) name690 (
		_w1370_,
		_w1463_,
		_w1464_
	);
	LUT2 #(
		.INIT('h4)
	) name691 (
		\g35_pad ,
		\g4411_reg/NET0131 ,
		_w1465_
	);
	LUT2 #(
		.INIT('h8)
	) name692 (
		\g35_pad ,
		_w1290_,
		_w1466_
	);
	LUT2 #(
		.INIT('h1)
	) name693 (
		_w1465_,
		_w1466_,
		_w1467_
	);
	LUT2 #(
		.INIT('h4)
	) name694 (
		_w1300_,
		_w1467_,
		_w1468_
	);
	LUT2 #(
		.INIT('h2)
	) name695 (
		\g1379_reg/NET0131 ,
		\g35_pad ,
		_w1469_
	);
	LUT2 #(
		.INIT('h1)
	) name696 (
		\g1384_reg/NET0131 ,
		_w1250_,
		_w1470_
	);
	LUT2 #(
		.INIT('h2)
	) name697 (
		_w1377_,
		_w1470_,
		_w1471_
	);
	LUT2 #(
		.INIT('h1)
	) name698 (
		_w1469_,
		_w1471_,
		_w1472_
	);
	LUT2 #(
		.INIT('h1)
	) name699 (
		\g4567_reg/NET0131 ,
		_w1085_,
		_w1473_
	);
	LUT2 #(
		.INIT('h1)
	) name700 (
		\g4498_reg/NET0131 ,
		_w1085_,
		_w1474_
	);
	LUT2 #(
		.INIT('h8)
	) name701 (
		\g218_reg/NET0131 ,
		\g8291_pad ,
		_w1475_
	);
	LUT2 #(
		.INIT('h2)
	) name702 (
		\g8358_pad ,
		_w1475_,
		_w1476_
	);
	LUT2 #(
		.INIT('h4)
	) name703 (
		\g191_reg/NET0131 ,
		_w1475_,
		_w1477_
	);
	LUT2 #(
		.INIT('h1)
	) name704 (
		_w1476_,
		_w1477_,
		_w1478_
	);
	LUT2 #(
		.INIT('h2)
	) name705 (
		\g35_pad ,
		_w1478_,
		_w1479_
	);
	LUT2 #(
		.INIT('h2)
	) name706 (
		\g222_reg/NET0131 ,
		\g35_pad ,
		_w1480_
	);
	LUT2 #(
		.INIT('h1)
	) name707 (
		_w1479_,
		_w1480_,
		_w1481_
	);
	LUT2 #(
		.INIT('h2)
	) name708 (
		\g347_reg/NET0131 ,
		\g35_pad ,
		_w1482_
	);
	LUT2 #(
		.INIT('h4)
	) name709 (
		\g347_reg/NET0131 ,
		\g35_pad ,
		_w1483_
	);
	LUT2 #(
		.INIT('h8)
	) name710 (
		\g7540_pad ,
		_w1483_,
		_w1484_
	);
	LUT2 #(
		.INIT('h1)
	) name711 (
		_w1482_,
		_w1484_,
		_w1485_
	);
	LUT2 #(
		.INIT('h1)
	) name712 (
		\g4242_reg/NET0131 ,
		\g4300_reg/NET0131 ,
		_w1486_
	);
	LUT2 #(
		.INIT('h2)
	) name713 (
		\g35_pad ,
		_w1486_,
		_w1487_
	);
	LUT2 #(
		.INIT('h4)
	) name714 (
		\g35_pad ,
		\g4297_reg/NET0131 ,
		_w1488_
	);
	LUT2 #(
		.INIT('h1)
	) name715 (
		_w1487_,
		_w1488_,
		_w1489_
	);
	LUT2 #(
		.INIT('h8)
	) name716 (
		_w816_,
		_w1388_,
		_w1490_
	);
	LUT2 #(
		.INIT('h4)
	) name717 (
		\g1105_reg/NET0131 ,
		_w1490_,
		_w1491_
	);
	LUT2 #(
		.INIT('h1)
	) name718 (
		\g1211_reg/NET0131 ,
		\g1216_reg/NET0131 ,
		_w1492_
	);
	LUT2 #(
		.INIT('h2)
	) name719 (
		\g1061_reg/NET0131 ,
		\g1205_reg/NET0131 ,
		_w1493_
	);
	LUT2 #(
		.INIT('h4)
	) name720 (
		\g1221_reg/NET0131 ,
		\g979_reg/NET0131 ,
		_w1494_
	);
	LUT2 #(
		.INIT('h8)
	) name721 (
		_w1493_,
		_w1494_,
		_w1495_
	);
	LUT2 #(
		.INIT('h8)
	) name722 (
		_w1492_,
		_w1495_,
		_w1496_
	);
	LUT2 #(
		.INIT('h8)
	) name723 (
		_w1319_,
		_w1496_,
		_w1497_
	);
	LUT2 #(
		.INIT('h2)
	) name724 (
		\g17316_pad ,
		_w1497_,
		_w1498_
	);
	LUT2 #(
		.INIT('h2)
	) name725 (
		_w1491_,
		_w1498_,
		_w1499_
	);
	LUT2 #(
		.INIT('h8)
	) name726 (
		\g35_pad ,
		_w1499_,
		_w1500_
	);
	LUT2 #(
		.INIT('h8)
	) name727 (
		\g1816_reg/NET0131 ,
		_w1500_,
		_w1501_
	);
	LUT2 #(
		.INIT('h2)
	) name728 (
		\g1802_reg/NET0131 ,
		\g35_pad ,
		_w1502_
	);
	LUT2 #(
		.INIT('h1)
	) name729 (
		\g1728_reg/NET0131 ,
		\g1802_reg/NET0131 ,
		_w1503_
	);
	LUT2 #(
		.INIT('h2)
	) name730 (
		\g1816_reg/NET0131 ,
		_w1503_,
		_w1504_
	);
	LUT2 #(
		.INIT('h8)
	) name731 (
		\g1246_reg/NET0131 ,
		_w1491_,
		_w1505_
	);
	LUT2 #(
		.INIT('h4)
	) name732 (
		_w1504_,
		_w1505_,
		_w1506_
	);
	LUT2 #(
		.INIT('h2)
	) name733 (
		_w1504_,
		_w1505_,
		_w1507_
	);
	LUT2 #(
		.INIT('h2)
	) name734 (
		\g35_pad ,
		_w1499_,
		_w1508_
	);
	LUT2 #(
		.INIT('h1)
	) name735 (
		_w1506_,
		_w1507_,
		_w1509_
	);
	LUT2 #(
		.INIT('h8)
	) name736 (
		_w1508_,
		_w1509_,
		_w1510_
	);
	LUT2 #(
		.INIT('h1)
	) name737 (
		_w1501_,
		_w1502_,
		_w1511_
	);
	LUT2 #(
		.INIT('h4)
	) name738 (
		_w1510_,
		_w1511_,
		_w1512_
	);
	LUT2 #(
		.INIT('h4)
	) name739 (
		\g1129_reg/NET0131 ,
		_w1490_,
		_w1513_
	);
	LUT2 #(
		.INIT('h8)
	) name740 (
		_w1331_,
		_w1496_,
		_w1514_
	);
	LUT2 #(
		.INIT('h2)
	) name741 (
		\g17400_pad ,
		_w1514_,
		_w1515_
	);
	LUT2 #(
		.INIT('h2)
	) name742 (
		_w1513_,
		_w1515_,
		_w1516_
	);
	LUT2 #(
		.INIT('h8)
	) name743 (
		\g35_pad ,
		_w1516_,
		_w1517_
	);
	LUT2 #(
		.INIT('h8)
	) name744 (
		\g1950_reg/NET0131 ,
		_w1517_,
		_w1518_
	);
	LUT2 #(
		.INIT('h2)
	) name745 (
		\g1936_reg/NET0131 ,
		\g35_pad ,
		_w1519_
	);
	LUT2 #(
		.INIT('h1)
	) name746 (
		\g1862_reg/NET0131 ,
		\g1936_reg/NET0131 ,
		_w1520_
	);
	LUT2 #(
		.INIT('h2)
	) name747 (
		\g1950_reg/NET0131 ,
		_w1520_,
		_w1521_
	);
	LUT2 #(
		.INIT('h4)
	) name748 (
		\g1246_reg/NET0131 ,
		_w1513_,
		_w1522_
	);
	LUT2 #(
		.INIT('h4)
	) name749 (
		_w1521_,
		_w1522_,
		_w1523_
	);
	LUT2 #(
		.INIT('h2)
	) name750 (
		_w1521_,
		_w1522_,
		_w1524_
	);
	LUT2 #(
		.INIT('h2)
	) name751 (
		\g35_pad ,
		_w1516_,
		_w1525_
	);
	LUT2 #(
		.INIT('h1)
	) name752 (
		_w1523_,
		_w1524_,
		_w1526_
	);
	LUT2 #(
		.INIT('h8)
	) name753 (
		_w1525_,
		_w1526_,
		_w1527_
	);
	LUT2 #(
		.INIT('h1)
	) name754 (
		_w1518_,
		_w1519_,
		_w1528_
	);
	LUT2 #(
		.INIT('h4)
	) name755 (
		_w1527_,
		_w1528_,
		_w1529_
	);
	LUT2 #(
		.INIT('h4)
	) name756 (
		\g956_reg/NET0131 ,
		_w1490_,
		_w1530_
	);
	LUT2 #(
		.INIT('h8)
	) name757 (
		_w1343_,
		_w1496_,
		_w1531_
	);
	LUT2 #(
		.INIT('h2)
	) name758 (
		\g1087_reg/NET0131 ,
		_w1531_,
		_w1532_
	);
	LUT2 #(
		.INIT('h2)
	) name759 (
		_w1530_,
		_w1532_,
		_w1533_
	);
	LUT2 #(
		.INIT('h8)
	) name760 (
		\g35_pad ,
		_w1533_,
		_w1534_
	);
	LUT2 #(
		.INIT('h8)
	) name761 (
		\g2084_reg/NET0131 ,
		_w1534_,
		_w1535_
	);
	LUT2 #(
		.INIT('h2)
	) name762 (
		\g2070_reg/NET0131 ,
		\g35_pad ,
		_w1536_
	);
	LUT2 #(
		.INIT('h1)
	) name763 (
		\g1996_reg/NET0131 ,
		\g2070_reg/NET0131 ,
		_w1537_
	);
	LUT2 #(
		.INIT('h2)
	) name764 (
		\g2084_reg/NET0131 ,
		_w1537_,
		_w1538_
	);
	LUT2 #(
		.INIT('h8)
	) name765 (
		\g1246_reg/NET0131 ,
		_w1530_,
		_w1539_
	);
	LUT2 #(
		.INIT('h4)
	) name766 (
		_w1538_,
		_w1539_,
		_w1540_
	);
	LUT2 #(
		.INIT('h2)
	) name767 (
		_w1538_,
		_w1539_,
		_w1541_
	);
	LUT2 #(
		.INIT('h2)
	) name768 (
		\g35_pad ,
		_w1533_,
		_w1542_
	);
	LUT2 #(
		.INIT('h1)
	) name769 (
		_w1540_,
		_w1541_,
		_w1543_
	);
	LUT2 #(
		.INIT('h8)
	) name770 (
		_w1542_,
		_w1543_,
		_w1544_
	);
	LUT2 #(
		.INIT('h1)
	) name771 (
		_w1535_,
		_w1536_,
		_w1545_
	);
	LUT2 #(
		.INIT('h4)
	) name772 (
		_w1544_,
		_w1545_,
		_w1546_
	);
	LUT2 #(
		.INIT('h1)
	) name773 (
		\g2970_reg/NET0131 ,
		\g35_pad ,
		_w1547_
	);
	LUT2 #(
		.INIT('h4)
	) name774 (
		\g301_reg/NET0131 ,
		\g35_pad ,
		_w1548_
	);
	LUT2 #(
		.INIT('h4)
	) name775 (
		\g2902_reg/NET0131 ,
		_w1388_,
		_w1549_
	);
	LUT2 #(
		.INIT('h8)
	) name776 (
		_w1548_,
		_w1549_,
		_w1550_
	);
	LUT2 #(
		.INIT('h1)
	) name777 (
		_w1547_,
		_w1550_,
		_w1551_
	);
	LUT2 #(
		.INIT('h2)
	) name778 (
		\g1306_reg/NET0131 ,
		_w1130_,
		_w1552_
	);
	LUT2 #(
		.INIT('h8)
	) name779 (
		\g1339_reg/NET0131 ,
		\g7946_pad ,
		_w1553_
	);
	LUT2 #(
		.INIT('h8)
	) name780 (
		_w1194_,
		_w1553_,
		_w1554_
	);
	LUT2 #(
		.INIT('h1)
	) name781 (
		_w1552_,
		_w1554_,
		_w1555_
	);
	LUT2 #(
		.INIT('h2)
	) name782 (
		\g35_pad ,
		_w1555_,
		_w1556_
	);
	LUT2 #(
		.INIT('h2)
	) name783 (
		\g1521_reg/NET0131 ,
		\g35_pad ,
		_w1557_
	);
	LUT2 #(
		.INIT('h1)
	) name784 (
		_w1556_,
		_w1557_,
		_w1558_
	);
	LUT2 #(
		.INIT('h4)
	) name785 (
		\g1585_reg/NET0131 ,
		_w1390_,
		_w1559_
	);
	LUT2 #(
		.INIT('h1)
	) name786 (
		\g2197_reg/NET0131 ,
		_w1398_,
		_w1560_
	);
	LUT2 #(
		.INIT('h8)
	) name787 (
		\g2153_reg/NET0131 ,
		_w1560_,
		_w1561_
	);
	LUT2 #(
		.INIT('h4)
	) name788 (
		_w1559_,
		_w1561_,
		_w1562_
	);
	LUT2 #(
		.INIT('h2)
	) name789 (
		\g2161_reg/NET0131 ,
		_w1561_,
		_w1563_
	);
	LUT2 #(
		.INIT('h1)
	) name790 (
		_w1562_,
		_w1563_,
		_w1564_
	);
	LUT2 #(
		.INIT('h2)
	) name791 (
		\g35_pad ,
		_w1564_,
		_w1565_
	);
	LUT2 #(
		.INIT('h2)
	) name792 (
		\g2165_reg/NET0131 ,
		\g35_pad ,
		_w1566_
	);
	LUT2 #(
		.INIT('h1)
	) name793 (
		_w1565_,
		_w1566_,
		_w1567_
	);
	LUT2 #(
		.INIT('h4)
	) name794 (
		_w1398_,
		_w1402_,
		_w1568_
	);
	LUT2 #(
		.INIT('h4)
	) name795 (
		_w1559_,
		_w1568_,
		_w1569_
	);
	LUT2 #(
		.INIT('h2)
	) name796 (
		\g2165_reg/NET0131 ,
		_w1568_,
		_w1570_
	);
	LUT2 #(
		.INIT('h1)
	) name797 (
		_w1569_,
		_w1570_,
		_w1571_
	);
	LUT2 #(
		.INIT('h2)
	) name798 (
		\g35_pad ,
		_w1571_,
		_w1572_
	);
	LUT2 #(
		.INIT('h2)
	) name799 (
		\g2246_reg/NET0131 ,
		\g35_pad ,
		_w1573_
	);
	LUT2 #(
		.INIT('h1)
	) name800 (
		_w1572_,
		_w1573_,
		_w1574_
	);
	LUT2 #(
		.INIT('h2)
	) name801 (
		\g2197_reg/NET0131 ,
		_w1398_,
		_w1575_
	);
	LUT2 #(
		.INIT('h4)
	) name802 (
		\g2227_reg/NET0131 ,
		_w1575_,
		_w1576_
	);
	LUT2 #(
		.INIT('h4)
	) name803 (
		_w1559_,
		_w1576_,
		_w1577_
	);
	LUT2 #(
		.INIT('h2)
	) name804 (
		\g2169_reg/NET0131 ,
		_w1576_,
		_w1578_
	);
	LUT2 #(
		.INIT('h1)
	) name805 (
		_w1577_,
		_w1578_,
		_w1579_
	);
	LUT2 #(
		.INIT('h2)
	) name806 (
		\g35_pad ,
		_w1579_,
		_w1580_
	);
	LUT2 #(
		.INIT('h2)
	) name807 (
		\g2161_reg/NET0131 ,
		\g35_pad ,
		_w1581_
	);
	LUT2 #(
		.INIT('h1)
	) name808 (
		_w1580_,
		_w1581_,
		_w1582_
	);
	LUT2 #(
		.INIT('h2)
	) name809 (
		\g2153_reg/NET0131 ,
		_w1398_,
		_w1583_
	);
	LUT2 #(
		.INIT('h8)
	) name810 (
		\g2227_reg/NET0131 ,
		_w1583_,
		_w1584_
	);
	LUT2 #(
		.INIT('h4)
	) name811 (
		_w1559_,
		_w1584_,
		_w1585_
	);
	LUT2 #(
		.INIT('h2)
	) name812 (
		\g2173_reg/NET0131 ,
		_w1584_,
		_w1586_
	);
	LUT2 #(
		.INIT('h1)
	) name813 (
		_w1585_,
		_w1586_,
		_w1587_
	);
	LUT2 #(
		.INIT('h2)
	) name814 (
		\g35_pad ,
		_w1587_,
		_w1588_
	);
	LUT2 #(
		.INIT('h2)
	) name815 (
		\g2177_reg/NET0131 ,
		\g35_pad ,
		_w1589_
	);
	LUT2 #(
		.INIT('h1)
	) name816 (
		_w1588_,
		_w1589_,
		_w1590_
	);
	LUT2 #(
		.INIT('h4)
	) name817 (
		\g2153_reg/NET0131 ,
		_w1575_,
		_w1591_
	);
	LUT2 #(
		.INIT('h4)
	) name818 (
		_w1559_,
		_w1591_,
		_w1592_
	);
	LUT2 #(
		.INIT('h2)
	) name819 (
		\g2177_reg/NET0131 ,
		_w1591_,
		_w1593_
	);
	LUT2 #(
		.INIT('h1)
	) name820 (
		_w1592_,
		_w1593_,
		_w1594_
	);
	LUT2 #(
		.INIT('h2)
	) name821 (
		\g35_pad ,
		_w1594_,
		_w1595_
	);
	LUT2 #(
		.INIT('h2)
	) name822 (
		\g2181_reg/NET0131 ,
		\g35_pad ,
		_w1596_
	);
	LUT2 #(
		.INIT('h1)
	) name823 (
		_w1595_,
		_w1596_,
		_w1597_
	);
	LUT2 #(
		.INIT('h8)
	) name824 (
		\g2227_reg/NET0131 ,
		_w1560_,
		_w1598_
	);
	LUT2 #(
		.INIT('h4)
	) name825 (
		_w1559_,
		_w1598_,
		_w1599_
	);
	LUT2 #(
		.INIT('h2)
	) name826 (
		\g2181_reg/NET0131 ,
		_w1598_,
		_w1600_
	);
	LUT2 #(
		.INIT('h1)
	) name827 (
		_w1599_,
		_w1600_,
		_w1601_
	);
	LUT2 #(
		.INIT('h2)
	) name828 (
		\g35_pad ,
		_w1601_,
		_w1602_
	);
	LUT2 #(
		.INIT('h2)
	) name829 (
		\g2169_reg/NET0131 ,
		\g35_pad ,
		_w1603_
	);
	LUT2 #(
		.INIT('h1)
	) name830 (
		_w1602_,
		_w1603_,
		_w1604_
	);
	LUT2 #(
		.INIT('h8)
	) name831 (
		\g1585_reg/NET0131 ,
		_w1412_,
		_w1605_
	);
	LUT2 #(
		.INIT('h1)
	) name832 (
		\g2331_reg/NET0131 ,
		_w1415_,
		_w1606_
	);
	LUT2 #(
		.INIT('h8)
	) name833 (
		\g2287_reg/NET0131 ,
		_w1606_,
		_w1607_
	);
	LUT2 #(
		.INIT('h4)
	) name834 (
		_w1605_,
		_w1607_,
		_w1608_
	);
	LUT2 #(
		.INIT('h2)
	) name835 (
		\g2295_reg/NET0131 ,
		_w1607_,
		_w1609_
	);
	LUT2 #(
		.INIT('h1)
	) name836 (
		_w1608_,
		_w1609_,
		_w1610_
	);
	LUT2 #(
		.INIT('h2)
	) name837 (
		\g35_pad ,
		_w1610_,
		_w1611_
	);
	LUT2 #(
		.INIT('h2)
	) name838 (
		\g2299_reg/NET0131 ,
		\g35_pad ,
		_w1612_
	);
	LUT2 #(
		.INIT('h1)
	) name839 (
		_w1611_,
		_w1612_,
		_w1613_
	);
	LUT2 #(
		.INIT('h4)
	) name840 (
		_w1415_,
		_w1419_,
		_w1614_
	);
	LUT2 #(
		.INIT('h4)
	) name841 (
		_w1605_,
		_w1614_,
		_w1615_
	);
	LUT2 #(
		.INIT('h2)
	) name842 (
		\g2299_reg/NET0131 ,
		_w1614_,
		_w1616_
	);
	LUT2 #(
		.INIT('h1)
	) name843 (
		_w1615_,
		_w1616_,
		_w1617_
	);
	LUT2 #(
		.INIT('h2)
	) name844 (
		\g35_pad ,
		_w1617_,
		_w1618_
	);
	LUT2 #(
		.INIT('h2)
	) name845 (
		\g2380_reg/NET0131 ,
		\g35_pad ,
		_w1619_
	);
	LUT2 #(
		.INIT('h1)
	) name846 (
		_w1618_,
		_w1619_,
		_w1620_
	);
	LUT2 #(
		.INIT('h2)
	) name847 (
		\g2331_reg/NET0131 ,
		_w1415_,
		_w1621_
	);
	LUT2 #(
		.INIT('h4)
	) name848 (
		\g2361_reg/NET0131 ,
		_w1621_,
		_w1622_
	);
	LUT2 #(
		.INIT('h4)
	) name849 (
		_w1605_,
		_w1622_,
		_w1623_
	);
	LUT2 #(
		.INIT('h2)
	) name850 (
		\g2303_reg/NET0131 ,
		_w1622_,
		_w1624_
	);
	LUT2 #(
		.INIT('h1)
	) name851 (
		_w1623_,
		_w1624_,
		_w1625_
	);
	LUT2 #(
		.INIT('h2)
	) name852 (
		\g35_pad ,
		_w1625_,
		_w1626_
	);
	LUT2 #(
		.INIT('h2)
	) name853 (
		\g2295_reg/NET0131 ,
		\g35_pad ,
		_w1627_
	);
	LUT2 #(
		.INIT('h1)
	) name854 (
		_w1626_,
		_w1627_,
		_w1628_
	);
	LUT2 #(
		.INIT('h2)
	) name855 (
		\g2287_reg/NET0131 ,
		_w1415_,
		_w1629_
	);
	LUT2 #(
		.INIT('h8)
	) name856 (
		\g2361_reg/NET0131 ,
		_w1629_,
		_w1630_
	);
	LUT2 #(
		.INIT('h4)
	) name857 (
		_w1605_,
		_w1630_,
		_w1631_
	);
	LUT2 #(
		.INIT('h2)
	) name858 (
		\g2307_reg/NET0131 ,
		_w1630_,
		_w1632_
	);
	LUT2 #(
		.INIT('h1)
	) name859 (
		_w1631_,
		_w1632_,
		_w1633_
	);
	LUT2 #(
		.INIT('h2)
	) name860 (
		\g35_pad ,
		_w1633_,
		_w1634_
	);
	LUT2 #(
		.INIT('h2)
	) name861 (
		\g2311_reg/NET0131 ,
		\g35_pad ,
		_w1635_
	);
	LUT2 #(
		.INIT('h1)
	) name862 (
		_w1634_,
		_w1635_,
		_w1636_
	);
	LUT2 #(
		.INIT('h4)
	) name863 (
		\g2287_reg/NET0131 ,
		_w1621_,
		_w1637_
	);
	LUT2 #(
		.INIT('h4)
	) name864 (
		_w1605_,
		_w1637_,
		_w1638_
	);
	LUT2 #(
		.INIT('h2)
	) name865 (
		\g2311_reg/NET0131 ,
		_w1637_,
		_w1639_
	);
	LUT2 #(
		.INIT('h1)
	) name866 (
		_w1638_,
		_w1639_,
		_w1640_
	);
	LUT2 #(
		.INIT('h2)
	) name867 (
		\g35_pad ,
		_w1640_,
		_w1641_
	);
	LUT2 #(
		.INIT('h2)
	) name868 (
		\g2315_reg/NET0131 ,
		\g35_pad ,
		_w1642_
	);
	LUT2 #(
		.INIT('h1)
	) name869 (
		_w1641_,
		_w1642_,
		_w1643_
	);
	LUT2 #(
		.INIT('h8)
	) name870 (
		\g2361_reg/NET0131 ,
		_w1606_,
		_w1644_
	);
	LUT2 #(
		.INIT('h4)
	) name871 (
		_w1605_,
		_w1644_,
		_w1645_
	);
	LUT2 #(
		.INIT('h2)
	) name872 (
		\g2315_reg/NET0131 ,
		_w1644_,
		_w1646_
	);
	LUT2 #(
		.INIT('h1)
	) name873 (
		_w1645_,
		_w1646_,
		_w1647_
	);
	LUT2 #(
		.INIT('h2)
	) name874 (
		\g35_pad ,
		_w1647_,
		_w1648_
	);
	LUT2 #(
		.INIT('h2)
	) name875 (
		\g2303_reg/NET0131 ,
		\g35_pad ,
		_w1649_
	);
	LUT2 #(
		.INIT('h1)
	) name876 (
		_w1648_,
		_w1649_,
		_w1650_
	);
	LUT2 #(
		.INIT('h2)
	) name877 (
		\g1521_reg/NET0131 ,
		\g7946_pad ,
		_w1651_
	);
	LUT2 #(
		.INIT('h1)
	) name878 (
		_w1553_,
		_w1651_,
		_w1652_
	);
	LUT2 #(
		.INIT('h2)
	) name879 (
		\g35_pad ,
		_w1652_,
		_w1653_
	);
	LUT2 #(
		.INIT('h2)
	) name880 (
		\g1526_reg/NET0131 ,
		\g35_pad ,
		_w1654_
	);
	LUT2 #(
		.INIT('h1)
	) name881 (
		_w1653_,
		_w1654_,
		_w1655_
	);
	LUT2 #(
		.INIT('h4)
	) name882 (
		\g1585_reg/NET0131 ,
		_w1429_,
		_w1656_
	);
	LUT2 #(
		.INIT('h1)
	) name883 (
		\g2465_reg/NET0131 ,
		_w1432_,
		_w1657_
	);
	LUT2 #(
		.INIT('h8)
	) name884 (
		\g2421_reg/NET0131 ,
		_w1657_,
		_w1658_
	);
	LUT2 #(
		.INIT('h4)
	) name885 (
		_w1656_,
		_w1658_,
		_w1659_
	);
	LUT2 #(
		.INIT('h2)
	) name886 (
		\g2429_reg/NET0131 ,
		_w1658_,
		_w1660_
	);
	LUT2 #(
		.INIT('h1)
	) name887 (
		_w1659_,
		_w1660_,
		_w1661_
	);
	LUT2 #(
		.INIT('h2)
	) name888 (
		\g35_pad ,
		_w1661_,
		_w1662_
	);
	LUT2 #(
		.INIT('h2)
	) name889 (
		\g2433_reg/NET0131 ,
		\g35_pad ,
		_w1663_
	);
	LUT2 #(
		.INIT('h1)
	) name890 (
		_w1662_,
		_w1663_,
		_w1664_
	);
	LUT2 #(
		.INIT('h4)
	) name891 (
		_w1432_,
		_w1436_,
		_w1665_
	);
	LUT2 #(
		.INIT('h4)
	) name892 (
		_w1656_,
		_w1665_,
		_w1666_
	);
	LUT2 #(
		.INIT('h2)
	) name893 (
		\g2433_reg/NET0131 ,
		_w1665_,
		_w1667_
	);
	LUT2 #(
		.INIT('h1)
	) name894 (
		_w1666_,
		_w1667_,
		_w1668_
	);
	LUT2 #(
		.INIT('h2)
	) name895 (
		\g35_pad ,
		_w1668_,
		_w1669_
	);
	LUT2 #(
		.INIT('h2)
	) name896 (
		\g2514_reg/NET0131 ,
		\g35_pad ,
		_w1670_
	);
	LUT2 #(
		.INIT('h1)
	) name897 (
		_w1669_,
		_w1670_,
		_w1671_
	);
	LUT2 #(
		.INIT('h2)
	) name898 (
		\g2465_reg/NET0131 ,
		_w1432_,
		_w1672_
	);
	LUT2 #(
		.INIT('h4)
	) name899 (
		\g2495_reg/NET0131 ,
		_w1672_,
		_w1673_
	);
	LUT2 #(
		.INIT('h4)
	) name900 (
		_w1656_,
		_w1673_,
		_w1674_
	);
	LUT2 #(
		.INIT('h2)
	) name901 (
		\g2437_reg/NET0131 ,
		_w1673_,
		_w1675_
	);
	LUT2 #(
		.INIT('h1)
	) name902 (
		_w1674_,
		_w1675_,
		_w1676_
	);
	LUT2 #(
		.INIT('h2)
	) name903 (
		\g35_pad ,
		_w1676_,
		_w1677_
	);
	LUT2 #(
		.INIT('h2)
	) name904 (
		\g2429_reg/NET0131 ,
		\g35_pad ,
		_w1678_
	);
	LUT2 #(
		.INIT('h1)
	) name905 (
		_w1677_,
		_w1678_,
		_w1679_
	);
	LUT2 #(
		.INIT('h2)
	) name906 (
		\g2421_reg/NET0131 ,
		_w1432_,
		_w1680_
	);
	LUT2 #(
		.INIT('h8)
	) name907 (
		\g2495_reg/NET0131 ,
		_w1680_,
		_w1681_
	);
	LUT2 #(
		.INIT('h4)
	) name908 (
		_w1656_,
		_w1681_,
		_w1682_
	);
	LUT2 #(
		.INIT('h2)
	) name909 (
		\g2441_reg/NET0131 ,
		_w1681_,
		_w1683_
	);
	LUT2 #(
		.INIT('h1)
	) name910 (
		_w1682_,
		_w1683_,
		_w1684_
	);
	LUT2 #(
		.INIT('h2)
	) name911 (
		\g35_pad ,
		_w1684_,
		_w1685_
	);
	LUT2 #(
		.INIT('h2)
	) name912 (
		\g2445_reg/NET0131 ,
		\g35_pad ,
		_w1686_
	);
	LUT2 #(
		.INIT('h1)
	) name913 (
		_w1685_,
		_w1686_,
		_w1687_
	);
	LUT2 #(
		.INIT('h4)
	) name914 (
		\g2421_reg/NET0131 ,
		_w1672_,
		_w1688_
	);
	LUT2 #(
		.INIT('h4)
	) name915 (
		_w1656_,
		_w1688_,
		_w1689_
	);
	LUT2 #(
		.INIT('h2)
	) name916 (
		\g2445_reg/NET0131 ,
		_w1688_,
		_w1690_
	);
	LUT2 #(
		.INIT('h1)
	) name917 (
		_w1689_,
		_w1690_,
		_w1691_
	);
	LUT2 #(
		.INIT('h2)
	) name918 (
		\g35_pad ,
		_w1691_,
		_w1692_
	);
	LUT2 #(
		.INIT('h2)
	) name919 (
		\g2449_reg/NET0131 ,
		\g35_pad ,
		_w1693_
	);
	LUT2 #(
		.INIT('h1)
	) name920 (
		_w1692_,
		_w1693_,
		_w1694_
	);
	LUT2 #(
		.INIT('h8)
	) name921 (
		\g2495_reg/NET0131 ,
		_w1657_,
		_w1695_
	);
	LUT2 #(
		.INIT('h4)
	) name922 (
		_w1656_,
		_w1695_,
		_w1696_
	);
	LUT2 #(
		.INIT('h2)
	) name923 (
		\g2449_reg/NET0131 ,
		_w1695_,
		_w1697_
	);
	LUT2 #(
		.INIT('h1)
	) name924 (
		_w1696_,
		_w1697_,
		_w1698_
	);
	LUT2 #(
		.INIT('h2)
	) name925 (
		\g35_pad ,
		_w1698_,
		_w1699_
	);
	LUT2 #(
		.INIT('h2)
	) name926 (
		\g2437_reg/NET0131 ,
		\g35_pad ,
		_w1700_
	);
	LUT2 #(
		.INIT('h1)
	) name927 (
		_w1699_,
		_w1700_,
		_w1701_
	);
	LUT2 #(
		.INIT('h8)
	) name928 (
		\g1585_reg/NET0131 ,
		_w1446_,
		_w1702_
	);
	LUT2 #(
		.INIT('h1)
	) name929 (
		\g2599_reg/NET0131 ,
		_w1449_,
		_w1703_
	);
	LUT2 #(
		.INIT('h8)
	) name930 (
		\g2555_reg/NET0131 ,
		_w1703_,
		_w1704_
	);
	LUT2 #(
		.INIT('h4)
	) name931 (
		_w1702_,
		_w1704_,
		_w1705_
	);
	LUT2 #(
		.INIT('h2)
	) name932 (
		\g2563_reg/NET0131 ,
		_w1704_,
		_w1706_
	);
	LUT2 #(
		.INIT('h1)
	) name933 (
		_w1705_,
		_w1706_,
		_w1707_
	);
	LUT2 #(
		.INIT('h2)
	) name934 (
		\g35_pad ,
		_w1707_,
		_w1708_
	);
	LUT2 #(
		.INIT('h2)
	) name935 (
		\g2567_reg/NET0131 ,
		\g35_pad ,
		_w1709_
	);
	LUT2 #(
		.INIT('h1)
	) name936 (
		_w1708_,
		_w1709_,
		_w1710_
	);
	LUT2 #(
		.INIT('h4)
	) name937 (
		_w1449_,
		_w1453_,
		_w1711_
	);
	LUT2 #(
		.INIT('h4)
	) name938 (
		_w1702_,
		_w1711_,
		_w1712_
	);
	LUT2 #(
		.INIT('h2)
	) name939 (
		\g2567_reg/NET0131 ,
		_w1711_,
		_w1713_
	);
	LUT2 #(
		.INIT('h1)
	) name940 (
		_w1712_,
		_w1713_,
		_w1714_
	);
	LUT2 #(
		.INIT('h2)
	) name941 (
		\g35_pad ,
		_w1714_,
		_w1715_
	);
	LUT2 #(
		.INIT('h2)
	) name942 (
		\g2648_reg/NET0131 ,
		\g35_pad ,
		_w1716_
	);
	LUT2 #(
		.INIT('h1)
	) name943 (
		_w1715_,
		_w1716_,
		_w1717_
	);
	LUT2 #(
		.INIT('h2)
	) name944 (
		\g2599_reg/NET0131 ,
		_w1449_,
		_w1718_
	);
	LUT2 #(
		.INIT('h4)
	) name945 (
		\g2629_reg/NET0131 ,
		_w1718_,
		_w1719_
	);
	LUT2 #(
		.INIT('h4)
	) name946 (
		_w1702_,
		_w1719_,
		_w1720_
	);
	LUT2 #(
		.INIT('h2)
	) name947 (
		\g2571_reg/NET0131 ,
		_w1719_,
		_w1721_
	);
	LUT2 #(
		.INIT('h1)
	) name948 (
		_w1720_,
		_w1721_,
		_w1722_
	);
	LUT2 #(
		.INIT('h2)
	) name949 (
		\g35_pad ,
		_w1722_,
		_w1723_
	);
	LUT2 #(
		.INIT('h2)
	) name950 (
		\g2563_reg/NET0131 ,
		\g35_pad ,
		_w1724_
	);
	LUT2 #(
		.INIT('h1)
	) name951 (
		_w1723_,
		_w1724_,
		_w1725_
	);
	LUT2 #(
		.INIT('h2)
	) name952 (
		\g2629_reg/NET0131 ,
		_w1449_,
		_w1726_
	);
	LUT2 #(
		.INIT('h8)
	) name953 (
		\g2555_reg/NET0131 ,
		_w1726_,
		_w1727_
	);
	LUT2 #(
		.INIT('h4)
	) name954 (
		_w1702_,
		_w1727_,
		_w1728_
	);
	LUT2 #(
		.INIT('h2)
	) name955 (
		\g2575_reg/NET0131 ,
		_w1727_,
		_w1729_
	);
	LUT2 #(
		.INIT('h1)
	) name956 (
		_w1728_,
		_w1729_,
		_w1730_
	);
	LUT2 #(
		.INIT('h2)
	) name957 (
		\g35_pad ,
		_w1730_,
		_w1731_
	);
	LUT2 #(
		.INIT('h2)
	) name958 (
		\g2579_reg/NET0131 ,
		\g35_pad ,
		_w1732_
	);
	LUT2 #(
		.INIT('h1)
	) name959 (
		_w1731_,
		_w1732_,
		_w1733_
	);
	LUT2 #(
		.INIT('h4)
	) name960 (
		\g2555_reg/NET0131 ,
		_w1718_,
		_w1734_
	);
	LUT2 #(
		.INIT('h4)
	) name961 (
		_w1702_,
		_w1734_,
		_w1735_
	);
	LUT2 #(
		.INIT('h2)
	) name962 (
		\g2579_reg/NET0131 ,
		_w1734_,
		_w1736_
	);
	LUT2 #(
		.INIT('h1)
	) name963 (
		_w1735_,
		_w1736_,
		_w1737_
	);
	LUT2 #(
		.INIT('h2)
	) name964 (
		\g35_pad ,
		_w1737_,
		_w1738_
	);
	LUT2 #(
		.INIT('h2)
	) name965 (
		\g2583_reg/NET0131 ,
		\g35_pad ,
		_w1739_
	);
	LUT2 #(
		.INIT('h1)
	) name966 (
		_w1738_,
		_w1739_,
		_w1740_
	);
	LUT2 #(
		.INIT('h8)
	) name967 (
		\g2629_reg/NET0131 ,
		_w1703_,
		_w1741_
	);
	LUT2 #(
		.INIT('h4)
	) name968 (
		_w1702_,
		_w1741_,
		_w1742_
	);
	LUT2 #(
		.INIT('h2)
	) name969 (
		\g2583_reg/NET0131 ,
		_w1741_,
		_w1743_
	);
	LUT2 #(
		.INIT('h1)
	) name970 (
		_w1742_,
		_w1743_,
		_w1744_
	);
	LUT2 #(
		.INIT('h2)
	) name971 (
		\g35_pad ,
		_w1744_,
		_w1745_
	);
	LUT2 #(
		.INIT('h2)
	) name972 (
		\g2571_reg/NET0131 ,
		\g35_pad ,
		_w1746_
	);
	LUT2 #(
		.INIT('h1)
	) name973 (
		_w1745_,
		_w1746_,
		_w1747_
	);
	LUT2 #(
		.INIT('h1)
	) name974 (
		\g4543_reg/NET0131 ,
		_w1085_,
		_w1748_
	);
	LUT2 #(
		.INIT('h2)
	) name975 (
		\g1395_reg/NET0131 ,
		\g35_pad ,
		_w1749_
	);
	LUT2 #(
		.INIT('h4)
	) name976 (
		\g1322_reg/NET0131 ,
		\g35_pad ,
		_w1750_
	);
	LUT2 #(
		.INIT('h2)
	) name977 (
		\g12923_pad ,
		_w1273_,
		_w1751_
	);
	LUT2 #(
		.INIT('h8)
	) name978 (
		\g1395_reg/NET0131 ,
		_w1751_,
		_w1752_
	);
	LUT2 #(
		.INIT('h8)
	) name979 (
		\g1404_reg/NET0131 ,
		_w1752_,
		_w1753_
	);
	LUT2 #(
		.INIT('h1)
	) name980 (
		\g1404_reg/NET0131 ,
		_w1752_,
		_w1754_
	);
	LUT2 #(
		.INIT('h2)
	) name981 (
		_w1750_,
		_w1753_,
		_w1755_
	);
	LUT2 #(
		.INIT('h4)
	) name982 (
		_w1754_,
		_w1755_,
		_w1756_
	);
	LUT2 #(
		.INIT('h1)
	) name983 (
		_w1749_,
		_w1756_,
		_w1757_
	);
	LUT2 #(
		.INIT('h2)
	) name984 (
		\g10527_pad ,
		\g17423_pad ,
		_w1758_
	);
	LUT2 #(
		.INIT('h8)
	) name985 (
		\g12923_pad ,
		\g17423_pad ,
		_w1759_
	);
	LUT2 #(
		.INIT('h1)
	) name986 (
		_w1758_,
		_w1759_,
		_w1760_
	);
	LUT2 #(
		.INIT('h2)
	) name987 (
		\g35_pad ,
		_w1760_,
		_w1761_
	);
	LUT2 #(
		.INIT('h2)
	) name988 (
		\g1589_reg/NET0131 ,
		\g35_pad ,
		_w1762_
	);
	LUT2 #(
		.INIT('h1)
	) name989 (
		_w1761_,
		_w1762_,
		_w1763_
	);
	LUT2 #(
		.INIT('h1)
	) name990 (
		\g35_pad ,
		\g542_reg/NET0131 ,
		_w1764_
	);
	LUT2 #(
		.INIT('h4)
	) name991 (
		\g534_reg/NET0131 ,
		_w1548_,
		_w1765_
	);
	LUT2 #(
		.INIT('h1)
	) name992 (
		_w1764_,
		_w1765_,
		_w1766_
	);
	LUT2 #(
		.INIT('h1)
	) name993 (
		\g4495_reg/NET0131 ,
		_w1085_,
		_w1767_
	);
	LUT2 #(
		.INIT('h2)
	) name994 (
		\g12923_pad ,
		\g1395_reg/NET0131 ,
		_w1768_
	);
	LUT2 #(
		.INIT('h8)
	) name995 (
		\g19357_pad ,
		_w1768_,
		_w1769_
	);
	LUT2 #(
		.INIT('h2)
	) name996 (
		\g35_pad ,
		_w1769_,
		_w1770_
	);
	LUT2 #(
		.INIT('h1)
	) name997 (
		\g1404_reg/NET0131 ,
		_w1770_,
		_w1771_
	);
	LUT2 #(
		.INIT('h4)
	) name998 (
		\g12923_pad ,
		\g1404_reg/NET0131 ,
		_w1772_
	);
	LUT2 #(
		.INIT('h8)
	) name999 (
		\g19357_pad ,
		\g35_pad ,
		_w1773_
	);
	LUT2 #(
		.INIT('h8)
	) name1000 (
		_w1772_,
		_w1773_,
		_w1774_
	);
	LUT2 #(
		.INIT('h1)
	) name1001 (
		_w1771_,
		_w1774_,
		_w1775_
	);
	LUT2 #(
		.INIT('h2)
	) name1002 (
		_w970_,
		_w1002_,
		_w1776_
	);
	LUT2 #(
		.INIT('h4)
	) name1003 (
		\g807_reg/NET0131 ,
		_w1001_,
		_w1777_
	);
	LUT2 #(
		.INIT('h2)
	) name1004 (
		\g35_pad ,
		_w1777_,
		_w1778_
	);
	LUT2 #(
		.INIT('h2)
	) name1005 (
		\g794_reg/NET0131 ,
		_w1778_,
		_w1779_
	);
	LUT2 #(
		.INIT('h1)
	) name1006 (
		_w1776_,
		_w1779_,
		_w1780_
	);
	LUT2 #(
		.INIT('h4)
	) name1007 (
		\g35_pad ,
		\g4427_reg/NET0131 ,
		_w1781_
	);
	LUT2 #(
		.INIT('h8)
	) name1008 (
		\g35_pad ,
		\g4423_reg/NET0131 ,
		_w1782_
	);
	LUT2 #(
		.INIT('h1)
	) name1009 (
		_w1781_,
		_w1782_,
		_w1783_
	);
	LUT2 #(
		.INIT('h1)
	) name1010 (
		\g1395_reg/NET0131 ,
		_w1751_,
		_w1784_
	);
	LUT2 #(
		.INIT('h2)
	) name1011 (
		_w1750_,
		_w1752_,
		_w1785_
	);
	LUT2 #(
		.INIT('h4)
	) name1012 (
		_w1784_,
		_w1785_,
		_w1786_
	);
	LUT2 #(
		.INIT('h4)
	) name1013 (
		\g4164_reg/NET0131 ,
		\g4253_reg/NET0131 ,
		_w1787_
	);
	LUT2 #(
		.INIT('h1)
	) name1014 (
		\g4145_reg/NET0131 ,
		\g4253_reg/NET0131 ,
		_w1788_
	);
	LUT2 #(
		.INIT('h1)
	) name1015 (
		_w1787_,
		_w1788_,
		_w1789_
	);
	LUT2 #(
		.INIT('h1)
	) name1016 (
		\g11770_pad ,
		\g8915_pad ,
		_w1790_
	);
	LUT2 #(
		.INIT('h1)
	) name1017 (
		\g8916_pad ,
		\g8917_pad ,
		_w1791_
	);
	LUT2 #(
		.INIT('h1)
	) name1018 (
		\g8918_pad ,
		\g8919_pad ,
		_w1792_
	);
	LUT2 #(
		.INIT('h4)
	) name1019 (
		\g8920_pad ,
		_w1792_,
		_w1793_
	);
	LUT2 #(
		.INIT('h8)
	) name1020 (
		_w1790_,
		_w1791_,
		_w1794_
	);
	LUT2 #(
		.INIT('h8)
	) name1021 (
		_w1793_,
		_w1794_,
		_w1795_
	);
	LUT2 #(
		.INIT('h1)
	) name1022 (
		\g8870_pad ,
		_w1795_,
		_w1796_
	);
	LUT2 #(
		.INIT('h1)
	) name1023 (
		\g4235_reg/NET0131 ,
		_w1796_,
		_w1797_
	);
	LUT2 #(
		.INIT('h2)
	) name1024 (
		\g4235_reg/NET0131 ,
		\g8870_pad ,
		_w1798_
	);
	LUT2 #(
		.INIT('h1)
	) name1025 (
		_w1797_,
		_w1798_,
		_w1799_
	);
	LUT2 #(
		.INIT('h2)
	) name1026 (
		_w1789_,
		_w1799_,
		_w1800_
	);
	LUT2 #(
		.INIT('h4)
	) name1027 (
		_w1789_,
		_w1799_,
		_w1801_
	);
	LUT2 #(
		.INIT('h1)
	) name1028 (
		_w1800_,
		_w1801_,
		_w1802_
	);
	LUT2 #(
		.INIT('h2)
	) name1029 (
		\g35_pad ,
		_w1802_,
		_w1803_
	);
	LUT2 #(
		.INIT('h4)
	) name1030 (
		\g35_pad ,
		\g4235_reg/NET0131 ,
		_w1804_
	);
	LUT2 #(
		.INIT('h1)
	) name1031 (
		_w1803_,
		_w1804_,
		_w1805_
	);
	LUT2 #(
		.INIT('h2)
	) name1032 (
		\g333_reg/NET0131 ,
		\g35_pad ,
		_w1806_
	);
	LUT2 #(
		.INIT('h1)
	) name1033 (
		_w1483_,
		_w1806_,
		_w1807_
	);
	LUT2 #(
		.INIT('h8)
	) name1034 (
		\g1242_reg/NET0131 ,
		_w1491_,
		_w1808_
	);
	LUT2 #(
		.INIT('h1)
	) name1035 (
		\g1772_reg/NET0131 ,
		_w1499_,
		_w1809_
	);
	LUT2 #(
		.INIT('h8)
	) name1036 (
		\g1728_reg/NET0131 ,
		_w1809_,
		_w1810_
	);
	LUT2 #(
		.INIT('h4)
	) name1037 (
		_w1808_,
		_w1810_,
		_w1811_
	);
	LUT2 #(
		.INIT('h2)
	) name1038 (
		\g1736_reg/NET0131 ,
		_w1810_,
		_w1812_
	);
	LUT2 #(
		.INIT('h1)
	) name1039 (
		_w1811_,
		_w1812_,
		_w1813_
	);
	LUT2 #(
		.INIT('h2)
	) name1040 (
		\g35_pad ,
		_w1813_,
		_w1814_
	);
	LUT2 #(
		.INIT('h2)
	) name1041 (
		\g1740_reg/NET0131 ,
		\g35_pad ,
		_w1815_
	);
	LUT2 #(
		.INIT('h1)
	) name1042 (
		_w1814_,
		_w1815_,
		_w1816_
	);
	LUT2 #(
		.INIT('h4)
	) name1043 (
		_w1499_,
		_w1503_,
		_w1817_
	);
	LUT2 #(
		.INIT('h4)
	) name1044 (
		_w1808_,
		_w1817_,
		_w1818_
	);
	LUT2 #(
		.INIT('h2)
	) name1045 (
		\g1740_reg/NET0131 ,
		_w1817_,
		_w1819_
	);
	LUT2 #(
		.INIT('h1)
	) name1046 (
		_w1818_,
		_w1819_,
		_w1820_
	);
	LUT2 #(
		.INIT('h2)
	) name1047 (
		\g35_pad ,
		_w1820_,
		_w1821_
	);
	LUT2 #(
		.INIT('h2)
	) name1048 (
		\g1821_reg/NET0131 ,
		\g35_pad ,
		_w1822_
	);
	LUT2 #(
		.INIT('h1)
	) name1049 (
		_w1821_,
		_w1822_,
		_w1823_
	);
	LUT2 #(
		.INIT('h2)
	) name1050 (
		\g1728_reg/NET0131 ,
		_w1499_,
		_w1824_
	);
	LUT2 #(
		.INIT('h8)
	) name1051 (
		\g1802_reg/NET0131 ,
		_w1824_,
		_w1825_
	);
	LUT2 #(
		.INIT('h4)
	) name1052 (
		_w1808_,
		_w1825_,
		_w1826_
	);
	LUT2 #(
		.INIT('h2)
	) name1053 (
		\g1748_reg/NET0131 ,
		_w1825_,
		_w1827_
	);
	LUT2 #(
		.INIT('h1)
	) name1054 (
		_w1826_,
		_w1827_,
		_w1828_
	);
	LUT2 #(
		.INIT('h2)
	) name1055 (
		\g35_pad ,
		_w1828_,
		_w1829_
	);
	LUT2 #(
		.INIT('h2)
	) name1056 (
		\g1752_reg/NET0131 ,
		\g35_pad ,
		_w1830_
	);
	LUT2 #(
		.INIT('h1)
	) name1057 (
		_w1829_,
		_w1830_,
		_w1831_
	);
	LUT2 #(
		.INIT('h2)
	) name1058 (
		\g1772_reg/NET0131 ,
		_w1499_,
		_w1832_
	);
	LUT2 #(
		.INIT('h4)
	) name1059 (
		\g1802_reg/NET0131 ,
		_w1832_,
		_w1833_
	);
	LUT2 #(
		.INIT('h4)
	) name1060 (
		_w1808_,
		_w1833_,
		_w1834_
	);
	LUT2 #(
		.INIT('h2)
	) name1061 (
		\g1744_reg/NET0131 ,
		_w1833_,
		_w1835_
	);
	LUT2 #(
		.INIT('h1)
	) name1062 (
		_w1834_,
		_w1835_,
		_w1836_
	);
	LUT2 #(
		.INIT('h2)
	) name1063 (
		\g35_pad ,
		_w1836_,
		_w1837_
	);
	LUT2 #(
		.INIT('h2)
	) name1064 (
		\g1736_reg/NET0131 ,
		\g35_pad ,
		_w1838_
	);
	LUT2 #(
		.INIT('h1)
	) name1065 (
		_w1837_,
		_w1838_,
		_w1839_
	);
	LUT2 #(
		.INIT('h4)
	) name1066 (
		\g1728_reg/NET0131 ,
		_w1832_,
		_w1840_
	);
	LUT2 #(
		.INIT('h4)
	) name1067 (
		_w1808_,
		_w1840_,
		_w1841_
	);
	LUT2 #(
		.INIT('h2)
	) name1068 (
		\g1752_reg/NET0131 ,
		_w1840_,
		_w1842_
	);
	LUT2 #(
		.INIT('h1)
	) name1069 (
		_w1841_,
		_w1842_,
		_w1843_
	);
	LUT2 #(
		.INIT('h2)
	) name1070 (
		\g35_pad ,
		_w1843_,
		_w1844_
	);
	LUT2 #(
		.INIT('h2)
	) name1071 (
		\g1756_reg/NET0131 ,
		\g35_pad ,
		_w1845_
	);
	LUT2 #(
		.INIT('h1)
	) name1072 (
		_w1844_,
		_w1845_,
		_w1846_
	);
	LUT2 #(
		.INIT('h8)
	) name1073 (
		\g1802_reg/NET0131 ,
		_w1809_,
		_w1847_
	);
	LUT2 #(
		.INIT('h4)
	) name1074 (
		_w1808_,
		_w1847_,
		_w1848_
	);
	LUT2 #(
		.INIT('h2)
	) name1075 (
		\g1756_reg/NET0131 ,
		_w1847_,
		_w1849_
	);
	LUT2 #(
		.INIT('h1)
	) name1076 (
		_w1848_,
		_w1849_,
		_w1850_
	);
	LUT2 #(
		.INIT('h2)
	) name1077 (
		\g35_pad ,
		_w1850_,
		_w1851_
	);
	LUT2 #(
		.INIT('h2)
	) name1078 (
		\g1744_reg/NET0131 ,
		\g35_pad ,
		_w1852_
	);
	LUT2 #(
		.INIT('h1)
	) name1079 (
		_w1851_,
		_w1852_,
		_w1853_
	);
	LUT2 #(
		.INIT('h4)
	) name1080 (
		\g1242_reg/NET0131 ,
		_w1513_,
		_w1854_
	);
	LUT2 #(
		.INIT('h1)
	) name1081 (
		\g1906_reg/NET0131 ,
		_w1516_,
		_w1855_
	);
	LUT2 #(
		.INIT('h8)
	) name1082 (
		\g1862_reg/NET0131 ,
		_w1855_,
		_w1856_
	);
	LUT2 #(
		.INIT('h4)
	) name1083 (
		_w1854_,
		_w1856_,
		_w1857_
	);
	LUT2 #(
		.INIT('h2)
	) name1084 (
		\g1870_reg/NET0131 ,
		_w1856_,
		_w1858_
	);
	LUT2 #(
		.INIT('h1)
	) name1085 (
		_w1857_,
		_w1858_,
		_w1859_
	);
	LUT2 #(
		.INIT('h2)
	) name1086 (
		\g35_pad ,
		_w1859_,
		_w1860_
	);
	LUT2 #(
		.INIT('h2)
	) name1087 (
		\g1874_reg/NET0131 ,
		\g35_pad ,
		_w1861_
	);
	LUT2 #(
		.INIT('h1)
	) name1088 (
		_w1860_,
		_w1861_,
		_w1862_
	);
	LUT2 #(
		.INIT('h4)
	) name1089 (
		_w1516_,
		_w1520_,
		_w1863_
	);
	LUT2 #(
		.INIT('h4)
	) name1090 (
		_w1854_,
		_w1863_,
		_w1864_
	);
	LUT2 #(
		.INIT('h2)
	) name1091 (
		\g1874_reg/NET0131 ,
		_w1863_,
		_w1865_
	);
	LUT2 #(
		.INIT('h1)
	) name1092 (
		_w1864_,
		_w1865_,
		_w1866_
	);
	LUT2 #(
		.INIT('h2)
	) name1093 (
		\g35_pad ,
		_w1866_,
		_w1867_
	);
	LUT2 #(
		.INIT('h2)
	) name1094 (
		\g1955_reg/NET0131 ,
		\g35_pad ,
		_w1868_
	);
	LUT2 #(
		.INIT('h1)
	) name1095 (
		_w1867_,
		_w1868_,
		_w1869_
	);
	LUT2 #(
		.INIT('h2)
	) name1096 (
		\g1906_reg/NET0131 ,
		_w1516_,
		_w1870_
	);
	LUT2 #(
		.INIT('h4)
	) name1097 (
		\g1936_reg/NET0131 ,
		_w1870_,
		_w1871_
	);
	LUT2 #(
		.INIT('h4)
	) name1098 (
		_w1854_,
		_w1871_,
		_w1872_
	);
	LUT2 #(
		.INIT('h2)
	) name1099 (
		\g1878_reg/NET0131 ,
		_w1871_,
		_w1873_
	);
	LUT2 #(
		.INIT('h1)
	) name1100 (
		_w1872_,
		_w1873_,
		_w1874_
	);
	LUT2 #(
		.INIT('h2)
	) name1101 (
		\g35_pad ,
		_w1874_,
		_w1875_
	);
	LUT2 #(
		.INIT('h2)
	) name1102 (
		\g1870_reg/NET0131 ,
		\g35_pad ,
		_w1876_
	);
	LUT2 #(
		.INIT('h1)
	) name1103 (
		_w1875_,
		_w1876_,
		_w1877_
	);
	LUT2 #(
		.INIT('h2)
	) name1104 (
		\g1862_reg/NET0131 ,
		_w1516_,
		_w1878_
	);
	LUT2 #(
		.INIT('h8)
	) name1105 (
		\g1936_reg/NET0131 ,
		_w1878_,
		_w1879_
	);
	LUT2 #(
		.INIT('h4)
	) name1106 (
		_w1854_,
		_w1879_,
		_w1880_
	);
	LUT2 #(
		.INIT('h2)
	) name1107 (
		\g1882_reg/NET0131 ,
		_w1879_,
		_w1881_
	);
	LUT2 #(
		.INIT('h1)
	) name1108 (
		_w1880_,
		_w1881_,
		_w1882_
	);
	LUT2 #(
		.INIT('h2)
	) name1109 (
		\g35_pad ,
		_w1882_,
		_w1883_
	);
	LUT2 #(
		.INIT('h2)
	) name1110 (
		\g1886_reg/NET0131 ,
		\g35_pad ,
		_w1884_
	);
	LUT2 #(
		.INIT('h1)
	) name1111 (
		_w1883_,
		_w1884_,
		_w1885_
	);
	LUT2 #(
		.INIT('h4)
	) name1112 (
		\g1862_reg/NET0131 ,
		_w1870_,
		_w1886_
	);
	LUT2 #(
		.INIT('h4)
	) name1113 (
		_w1854_,
		_w1886_,
		_w1887_
	);
	LUT2 #(
		.INIT('h2)
	) name1114 (
		\g1886_reg/NET0131 ,
		_w1886_,
		_w1888_
	);
	LUT2 #(
		.INIT('h1)
	) name1115 (
		_w1887_,
		_w1888_,
		_w1889_
	);
	LUT2 #(
		.INIT('h2)
	) name1116 (
		\g35_pad ,
		_w1889_,
		_w1890_
	);
	LUT2 #(
		.INIT('h2)
	) name1117 (
		\g1890_reg/NET0131 ,
		\g35_pad ,
		_w1891_
	);
	LUT2 #(
		.INIT('h1)
	) name1118 (
		_w1890_,
		_w1891_,
		_w1892_
	);
	LUT2 #(
		.INIT('h8)
	) name1119 (
		\g1936_reg/NET0131 ,
		_w1855_,
		_w1893_
	);
	LUT2 #(
		.INIT('h4)
	) name1120 (
		_w1854_,
		_w1893_,
		_w1894_
	);
	LUT2 #(
		.INIT('h2)
	) name1121 (
		\g1890_reg/NET0131 ,
		_w1893_,
		_w1895_
	);
	LUT2 #(
		.INIT('h1)
	) name1122 (
		_w1894_,
		_w1895_,
		_w1896_
	);
	LUT2 #(
		.INIT('h2)
	) name1123 (
		\g35_pad ,
		_w1896_,
		_w1897_
	);
	LUT2 #(
		.INIT('h2)
	) name1124 (
		\g1878_reg/NET0131 ,
		\g35_pad ,
		_w1898_
	);
	LUT2 #(
		.INIT('h1)
	) name1125 (
		_w1897_,
		_w1898_,
		_w1899_
	);
	LUT2 #(
		.INIT('h8)
	) name1126 (
		\g1242_reg/NET0131 ,
		_w1530_,
		_w1900_
	);
	LUT2 #(
		.INIT('h2)
	) name1127 (
		\g1996_reg/NET0131 ,
		_w1533_,
		_w1901_
	);
	LUT2 #(
		.INIT('h4)
	) name1128 (
		\g2040_reg/NET0131 ,
		_w1901_,
		_w1902_
	);
	LUT2 #(
		.INIT('h4)
	) name1129 (
		_w1900_,
		_w1902_,
		_w1903_
	);
	LUT2 #(
		.INIT('h2)
	) name1130 (
		\g2004_reg/NET0131 ,
		_w1902_,
		_w1904_
	);
	LUT2 #(
		.INIT('h1)
	) name1131 (
		_w1903_,
		_w1904_,
		_w1905_
	);
	LUT2 #(
		.INIT('h2)
	) name1132 (
		\g35_pad ,
		_w1905_,
		_w1906_
	);
	LUT2 #(
		.INIT('h2)
	) name1133 (
		\g2008_reg/NET0131 ,
		\g35_pad ,
		_w1907_
	);
	LUT2 #(
		.INIT('h1)
	) name1134 (
		_w1906_,
		_w1907_,
		_w1908_
	);
	LUT2 #(
		.INIT('h4)
	) name1135 (
		_w1533_,
		_w1537_,
		_w1909_
	);
	LUT2 #(
		.INIT('h4)
	) name1136 (
		_w1900_,
		_w1909_,
		_w1910_
	);
	LUT2 #(
		.INIT('h2)
	) name1137 (
		\g2008_reg/NET0131 ,
		_w1909_,
		_w1911_
	);
	LUT2 #(
		.INIT('h1)
	) name1138 (
		_w1910_,
		_w1911_,
		_w1912_
	);
	LUT2 #(
		.INIT('h2)
	) name1139 (
		\g35_pad ,
		_w1912_,
		_w1913_
	);
	LUT2 #(
		.INIT('h2)
	) name1140 (
		\g2089_reg/NET0131 ,
		\g35_pad ,
		_w1914_
	);
	LUT2 #(
		.INIT('h1)
	) name1141 (
		_w1913_,
		_w1914_,
		_w1915_
	);
	LUT2 #(
		.INIT('h2)
	) name1142 (
		\g2040_reg/NET0131 ,
		_w1533_,
		_w1916_
	);
	LUT2 #(
		.INIT('h4)
	) name1143 (
		\g2070_reg/NET0131 ,
		_w1916_,
		_w1917_
	);
	LUT2 #(
		.INIT('h4)
	) name1144 (
		_w1900_,
		_w1917_,
		_w1918_
	);
	LUT2 #(
		.INIT('h2)
	) name1145 (
		\g2012_reg/NET0131 ,
		_w1917_,
		_w1919_
	);
	LUT2 #(
		.INIT('h1)
	) name1146 (
		_w1918_,
		_w1919_,
		_w1920_
	);
	LUT2 #(
		.INIT('h2)
	) name1147 (
		\g35_pad ,
		_w1920_,
		_w1921_
	);
	LUT2 #(
		.INIT('h2)
	) name1148 (
		\g2004_reg/NET0131 ,
		\g35_pad ,
		_w1922_
	);
	LUT2 #(
		.INIT('h1)
	) name1149 (
		_w1921_,
		_w1922_,
		_w1923_
	);
	LUT2 #(
		.INIT('h8)
	) name1150 (
		\g2070_reg/NET0131 ,
		_w1901_,
		_w1924_
	);
	LUT2 #(
		.INIT('h4)
	) name1151 (
		_w1900_,
		_w1924_,
		_w1925_
	);
	LUT2 #(
		.INIT('h2)
	) name1152 (
		\g2016_reg/NET0131 ,
		_w1924_,
		_w1926_
	);
	LUT2 #(
		.INIT('h1)
	) name1153 (
		_w1925_,
		_w1926_,
		_w1927_
	);
	LUT2 #(
		.INIT('h2)
	) name1154 (
		\g35_pad ,
		_w1927_,
		_w1928_
	);
	LUT2 #(
		.INIT('h2)
	) name1155 (
		\g2020_reg/NET0131 ,
		\g35_pad ,
		_w1929_
	);
	LUT2 #(
		.INIT('h1)
	) name1156 (
		_w1928_,
		_w1929_,
		_w1930_
	);
	LUT2 #(
		.INIT('h4)
	) name1157 (
		\g1996_reg/NET0131 ,
		_w1916_,
		_w1931_
	);
	LUT2 #(
		.INIT('h4)
	) name1158 (
		_w1900_,
		_w1931_,
		_w1932_
	);
	LUT2 #(
		.INIT('h2)
	) name1159 (
		\g2020_reg/NET0131 ,
		_w1931_,
		_w1933_
	);
	LUT2 #(
		.INIT('h1)
	) name1160 (
		_w1932_,
		_w1933_,
		_w1934_
	);
	LUT2 #(
		.INIT('h2)
	) name1161 (
		\g35_pad ,
		_w1934_,
		_w1935_
	);
	LUT2 #(
		.INIT('h2)
	) name1162 (
		\g2024_reg/NET0131 ,
		\g35_pad ,
		_w1936_
	);
	LUT2 #(
		.INIT('h1)
	) name1163 (
		_w1935_,
		_w1936_,
		_w1937_
	);
	LUT2 #(
		.INIT('h1)
	) name1164 (
		\g2040_reg/NET0131 ,
		_w1533_,
		_w1938_
	);
	LUT2 #(
		.INIT('h8)
	) name1165 (
		\g2070_reg/NET0131 ,
		_w1938_,
		_w1939_
	);
	LUT2 #(
		.INIT('h4)
	) name1166 (
		_w1900_,
		_w1939_,
		_w1940_
	);
	LUT2 #(
		.INIT('h2)
	) name1167 (
		\g2024_reg/NET0131 ,
		_w1939_,
		_w1941_
	);
	LUT2 #(
		.INIT('h1)
	) name1168 (
		_w1940_,
		_w1941_,
		_w1942_
	);
	LUT2 #(
		.INIT('h2)
	) name1169 (
		\g35_pad ,
		_w1942_,
		_w1943_
	);
	LUT2 #(
		.INIT('h2)
	) name1170 (
		\g2012_reg/NET0131 ,
		\g35_pad ,
		_w1944_
	);
	LUT2 #(
		.INIT('h1)
	) name1171 (
		_w1943_,
		_w1944_,
		_w1945_
	);
	LUT2 #(
		.INIT('h4)
	) name1172 (
		\g1135_reg/NET0131 ,
		_w1490_,
		_w1946_
	);
	LUT2 #(
		.INIT('h4)
	) name1173 (
		\g1242_reg/NET0131 ,
		_w1946_,
		_w1947_
	);
	LUT2 #(
		.INIT('h8)
	) name1174 (
		_w1305_,
		_w1496_,
		_w1948_
	);
	LUT2 #(
		.INIT('h2)
	) name1175 (
		\g17291_pad ,
		_w1948_,
		_w1949_
	);
	LUT2 #(
		.INIT('h2)
	) name1176 (
		_w1946_,
		_w1949_,
		_w1950_
	);
	LUT2 #(
		.INIT('h2)
	) name1177 (
		\g1592_reg/NET0131 ,
		_w1950_,
		_w1951_
	);
	LUT2 #(
		.INIT('h4)
	) name1178 (
		\g1636_reg/NET0131 ,
		_w1951_,
		_w1952_
	);
	LUT2 #(
		.INIT('h4)
	) name1179 (
		_w1947_,
		_w1952_,
		_w1953_
	);
	LUT2 #(
		.INIT('h2)
	) name1180 (
		\g1600_reg/NET0131 ,
		_w1952_,
		_w1954_
	);
	LUT2 #(
		.INIT('h1)
	) name1181 (
		_w1953_,
		_w1954_,
		_w1955_
	);
	LUT2 #(
		.INIT('h2)
	) name1182 (
		\g35_pad ,
		_w1955_,
		_w1956_
	);
	LUT2 #(
		.INIT('h2)
	) name1183 (
		\g1604_reg/NET0131 ,
		\g35_pad ,
		_w1957_
	);
	LUT2 #(
		.INIT('h1)
	) name1184 (
		_w1956_,
		_w1957_,
		_w1958_
	);
	LUT2 #(
		.INIT('h1)
	) name1185 (
		\g1592_reg/NET0131 ,
		\g1668_reg/NET0131 ,
		_w1959_
	);
	LUT2 #(
		.INIT('h4)
	) name1186 (
		_w1950_,
		_w1959_,
		_w1960_
	);
	LUT2 #(
		.INIT('h4)
	) name1187 (
		_w1947_,
		_w1960_,
		_w1961_
	);
	LUT2 #(
		.INIT('h2)
	) name1188 (
		\g1604_reg/NET0131 ,
		_w1960_,
		_w1962_
	);
	LUT2 #(
		.INIT('h1)
	) name1189 (
		_w1961_,
		_w1962_,
		_w1963_
	);
	LUT2 #(
		.INIT('h2)
	) name1190 (
		\g35_pad ,
		_w1963_,
		_w1964_
	);
	LUT2 #(
		.INIT('h2)
	) name1191 (
		\g1687_reg/NET0131 ,
		\g35_pad ,
		_w1965_
	);
	LUT2 #(
		.INIT('h1)
	) name1192 (
		_w1964_,
		_w1965_,
		_w1966_
	);
	LUT2 #(
		.INIT('h2)
	) name1193 (
		\g1636_reg/NET0131 ,
		_w1950_,
		_w1967_
	);
	LUT2 #(
		.INIT('h4)
	) name1194 (
		\g1668_reg/NET0131 ,
		_w1967_,
		_w1968_
	);
	LUT2 #(
		.INIT('h4)
	) name1195 (
		_w1947_,
		_w1968_,
		_w1969_
	);
	LUT2 #(
		.INIT('h2)
	) name1196 (
		\g1608_reg/NET0131 ,
		_w1968_,
		_w1970_
	);
	LUT2 #(
		.INIT('h1)
	) name1197 (
		_w1969_,
		_w1970_,
		_w1971_
	);
	LUT2 #(
		.INIT('h2)
	) name1198 (
		\g35_pad ,
		_w1971_,
		_w1972_
	);
	LUT2 #(
		.INIT('h2)
	) name1199 (
		\g1600_reg/NET0131 ,
		\g35_pad ,
		_w1973_
	);
	LUT2 #(
		.INIT('h1)
	) name1200 (
		_w1972_,
		_w1973_,
		_w1974_
	);
	LUT2 #(
		.INIT('h8)
	) name1201 (
		\g1668_reg/NET0131 ,
		_w1951_,
		_w1975_
	);
	LUT2 #(
		.INIT('h4)
	) name1202 (
		_w1947_,
		_w1975_,
		_w1976_
	);
	LUT2 #(
		.INIT('h2)
	) name1203 (
		\g1612_reg/NET0131 ,
		_w1975_,
		_w1977_
	);
	LUT2 #(
		.INIT('h1)
	) name1204 (
		_w1976_,
		_w1977_,
		_w1978_
	);
	LUT2 #(
		.INIT('h2)
	) name1205 (
		\g35_pad ,
		_w1978_,
		_w1979_
	);
	LUT2 #(
		.INIT('h2)
	) name1206 (
		\g1616_reg/NET0131 ,
		\g35_pad ,
		_w1980_
	);
	LUT2 #(
		.INIT('h1)
	) name1207 (
		_w1979_,
		_w1980_,
		_w1981_
	);
	LUT2 #(
		.INIT('h4)
	) name1208 (
		\g1592_reg/NET0131 ,
		_w1967_,
		_w1982_
	);
	LUT2 #(
		.INIT('h4)
	) name1209 (
		_w1947_,
		_w1982_,
		_w1983_
	);
	LUT2 #(
		.INIT('h2)
	) name1210 (
		\g1616_reg/NET0131 ,
		_w1982_,
		_w1984_
	);
	LUT2 #(
		.INIT('h1)
	) name1211 (
		_w1983_,
		_w1984_,
		_w1985_
	);
	LUT2 #(
		.INIT('h2)
	) name1212 (
		\g35_pad ,
		_w1985_,
		_w1986_
	);
	LUT2 #(
		.INIT('h2)
	) name1213 (
		\g1620_reg/NET0131 ,
		\g35_pad ,
		_w1987_
	);
	LUT2 #(
		.INIT('h1)
	) name1214 (
		_w1986_,
		_w1987_,
		_w1988_
	);
	LUT2 #(
		.INIT('h2)
	) name1215 (
		_w828_,
		_w1950_,
		_w1989_
	);
	LUT2 #(
		.INIT('h4)
	) name1216 (
		_w1947_,
		_w1989_,
		_w1990_
	);
	LUT2 #(
		.INIT('h2)
	) name1217 (
		\g1620_reg/NET0131 ,
		_w1989_,
		_w1991_
	);
	LUT2 #(
		.INIT('h1)
	) name1218 (
		_w1990_,
		_w1991_,
		_w1992_
	);
	LUT2 #(
		.INIT('h2)
	) name1219 (
		\g35_pad ,
		_w1992_,
		_w1993_
	);
	LUT2 #(
		.INIT('h2)
	) name1220 (
		\g1608_reg/NET0131 ,
		\g35_pad ,
		_w1994_
	);
	LUT2 #(
		.INIT('h1)
	) name1221 (
		_w1993_,
		_w1994_,
		_w1995_
	);
	LUT2 #(
		.INIT('h4)
	) name1222 (
		\g35_pad ,
		\g790_reg/NET0131 ,
		_w1996_
	);
	LUT2 #(
		.INIT('h2)
	) name1223 (
		\g794_reg/NET0131 ,
		_w966_,
		_w1997_
	);
	LUT2 #(
		.INIT('h1)
	) name1224 (
		_w1001_,
		_w1997_,
		_w1998_
	);
	LUT2 #(
		.INIT('h2)
	) name1225 (
		\g35_pad ,
		_w1002_,
		_w1999_
	);
	LUT2 #(
		.INIT('h4)
	) name1226 (
		_w1998_,
		_w1999_,
		_w2000_
	);
	LUT2 #(
		.INIT('h1)
	) name1227 (
		_w1996_,
		_w2000_,
		_w2001_
	);
	LUT2 #(
		.INIT('h2)
	) name1228 (
		\g1585_reg/NET0131 ,
		\g35_pad ,
		_w2002_
	);
	LUT2 #(
		.INIT('h8)
	) name1229 (
		\g12923_pad ,
		\g35_pad ,
		_w2003_
	);
	LUT2 #(
		.INIT('h1)
	) name1230 (
		_w2002_,
		_w2003_,
		_w2004_
	);
	LUT2 #(
		.INIT('h4)
	) name1231 (
		\g513_reg/NET0131 ,
		\g518_reg/NET0131 ,
		_w2005_
	);
	LUT2 #(
		.INIT('h8)
	) name1232 (
		\g203_reg/NET0131 ,
		_w2005_,
		_w2006_
	);
	LUT2 #(
		.INIT('h1)
	) name1233 (
		\g174_reg/NET0131 ,
		\g182_reg/NET0131 ,
		_w2007_
	);
	LUT2 #(
		.INIT('h4)
	) name1234 (
		\g168_reg/NET0131 ,
		_w2007_,
		_w2008_
	);
	LUT2 #(
		.INIT('h2)
	) name1235 (
		_w2006_,
		_w2008_,
		_w2009_
	);
	LUT2 #(
		.INIT('h2)
	) name1236 (
		\g691_reg/NET0131 ,
		_w2009_,
		_w2010_
	);
	LUT2 #(
		.INIT('h8)
	) name1237 (
		\g146_reg/NET0131 ,
		_w2006_,
		_w2011_
	);
	LUT2 #(
		.INIT('h8)
	) name1238 (
		\g164_reg/NET0131 ,
		_w2011_,
		_w2012_
	);
	LUT2 #(
		.INIT('h8)
	) name1239 (
		_w2010_,
		_w2012_,
		_w2013_
	);
	LUT2 #(
		.INIT('h8)
	) name1240 (
		\g150_reg/NET0131 ,
		_w2013_,
		_w2014_
	);
	LUT2 #(
		.INIT('h8)
	) name1241 (
		_w984_,
		_w987_,
		_w2015_
	);
	LUT2 #(
		.INIT('h8)
	) name1242 (
		_w979_,
		_w2015_,
		_w2016_
	);
	LUT2 #(
		.INIT('h2)
	) name1243 (
		_w2010_,
		_w2016_,
		_w2017_
	);
	LUT2 #(
		.INIT('h8)
	) name1244 (
		\g153_reg/NET0131 ,
		_w2014_,
		_w2018_
	);
	LUT2 #(
		.INIT('h8)
	) name1245 (
		_w2017_,
		_w2018_,
		_w2019_
	);
	LUT2 #(
		.INIT('h4)
	) name1246 (
		\g160_reg/NET0131 ,
		_w2019_,
		_w2020_
	);
	LUT2 #(
		.INIT('h2)
	) name1247 (
		\g35_pad ,
		_w2020_,
		_w2021_
	);
	LUT2 #(
		.INIT('h2)
	) name1248 (
		\g157_reg/NET0131 ,
		_w2021_,
		_w2022_
	);
	LUT2 #(
		.INIT('h8)
	) name1249 (
		\g157_reg/NET0131 ,
		_w2019_,
		_w2023_
	);
	LUT2 #(
		.INIT('h8)
	) name1250 (
		\g35_pad ,
		_w2017_,
		_w2024_
	);
	LUT2 #(
		.INIT('h8)
	) name1251 (
		\g160_reg/NET0131 ,
		_w2024_,
		_w2025_
	);
	LUT2 #(
		.INIT('h4)
	) name1252 (
		_w2023_,
		_w2025_,
		_w2026_
	);
	LUT2 #(
		.INIT('h1)
	) name1253 (
		_w2022_,
		_w2026_,
		_w2027_
	);
	LUT2 #(
		.INIT('h2)
	) name1254 (
		\g246_reg/NET0131 ,
		\g269_reg/NET0131 ,
		_w2028_
	);
	LUT2 #(
		.INIT('h2)
	) name1255 (
		\g239_reg/NET0131 ,
		\g262_reg/NET0131 ,
		_w2029_
	);
	LUT2 #(
		.INIT('h2)
	) name1256 (
		\g232_reg/NET0131 ,
		\g255_reg/NET0131 ,
		_w2030_
	);
	LUT2 #(
		.INIT('h8)
	) name1257 (
		\g225_reg/NET0131 ,
		_w2028_,
		_w2031_
	);
	LUT2 #(
		.INIT('h8)
	) name1258 (
		_w2029_,
		_w2030_,
		_w2032_
	);
	LUT2 #(
		.INIT('h8)
	) name1259 (
		_w2031_,
		_w2032_,
		_w2033_
	);
	LUT2 #(
		.INIT('h2)
	) name1260 (
		\g278_reg/NET0131 ,
		_w2033_,
		_w2034_
	);
	LUT2 #(
		.INIT('h4)
	) name1261 (
		\g232_reg/NET0131 ,
		\g255_reg/NET0131 ,
		_w2035_
	);
	LUT2 #(
		.INIT('h4)
	) name1262 (
		\g239_reg/NET0131 ,
		\g262_reg/NET0131 ,
		_w2036_
	);
	LUT2 #(
		.INIT('h4)
	) name1263 (
		\g246_reg/NET0131 ,
		\g269_reg/NET0131 ,
		_w2037_
	);
	LUT2 #(
		.INIT('h4)
	) name1264 (
		\g225_reg/NET0131 ,
		_w2035_,
		_w2038_
	);
	LUT2 #(
		.INIT('h8)
	) name1265 (
		_w2036_,
		_w2037_,
		_w2039_
	);
	LUT2 #(
		.INIT('h8)
	) name1266 (
		_w2038_,
		_w2039_,
		_w2040_
	);
	LUT2 #(
		.INIT('h1)
	) name1267 (
		\g278_reg/NET0131 ,
		_w2040_,
		_w2041_
	);
	LUT2 #(
		.INIT('h2)
	) name1268 (
		\g691_reg/NET0131 ,
		_w2034_,
		_w2042_
	);
	LUT2 #(
		.INIT('h4)
	) name1269 (
		_w2041_,
		_w2042_,
		_w2043_
	);
	LUT2 #(
		.INIT('h4)
	) name1270 (
		_w2016_,
		_w2043_,
		_w2044_
	);
	LUT2 #(
		.INIT('h8)
	) name1271 (
		\g283_reg/NET0131 ,
		\g287_reg/NET0131 ,
		_w2045_
	);
	LUT2 #(
		.INIT('h8)
	) name1272 (
		_w2044_,
		_w2045_,
		_w2046_
	);
	LUT2 #(
		.INIT('h8)
	) name1273 (
		\g291_reg/NET0131 ,
		_w2046_,
		_w2047_
	);
	LUT2 #(
		.INIT('h8)
	) name1274 (
		\g294_reg/NET0131 ,
		\g298_reg/NET0131 ,
		_w2048_
	);
	LUT2 #(
		.INIT('h8)
	) name1275 (
		_w2047_,
		_w2048_,
		_w2049_
	);
	LUT2 #(
		.INIT('h4)
	) name1276 (
		\g142_reg/NET0131 ,
		\g35_pad ,
		_w2050_
	);
	LUT2 #(
		.INIT('h8)
	) name1277 (
		_w2049_,
		_w2050_,
		_w2051_
	);
	LUT2 #(
		.INIT('h2)
	) name1278 (
		\g298_reg/NET0131 ,
		\g35_pad ,
		_w2052_
	);
	LUT2 #(
		.INIT('h8)
	) name1279 (
		\g35_pad ,
		_w2044_,
		_w2053_
	);
	LUT2 #(
		.INIT('h8)
	) name1280 (
		\g142_reg/NET0131 ,
		_w2053_,
		_w2054_
	);
	LUT2 #(
		.INIT('h4)
	) name1281 (
		_w2049_,
		_w2054_,
		_w2055_
	);
	LUT2 #(
		.INIT('h1)
	) name1282 (
		_w2051_,
		_w2052_,
		_w2056_
	);
	LUT2 #(
		.INIT('h4)
	) name1283 (
		_w2055_,
		_w2056_,
		_w2057_
	);
	LUT2 #(
		.INIT('h1)
	) name1284 (
		\g4540_reg/NET0131 ,
		_w1085_,
		_w2058_
	);
	LUT2 #(
		.INIT('h2)
	) name1285 (
		\g10500_pad ,
		\g17400_pad ,
		_w2059_
	);
	LUT2 #(
		.INIT('h8)
	) name1286 (
		\g12919_pad ,
		\g17400_pad ,
		_w2060_
	);
	LUT2 #(
		.INIT('h1)
	) name1287 (
		_w2059_,
		_w2060_,
		_w2061_
	);
	LUT2 #(
		.INIT('h2)
	) name1288 (
		\g35_pad ,
		_w2061_,
		_w2062_
	);
	LUT2 #(
		.INIT('h2)
	) name1289 (
		\g1246_reg/NET0131 ,
		\g35_pad ,
		_w2063_
	);
	LUT2 #(
		.INIT('h1)
	) name1290 (
		_w2062_,
		_w2063_,
		_w2064_
	);
	LUT2 #(
		.INIT('h2)
	) name1291 (
		\g1052_reg/NET0131 ,
		\g35_pad ,
		_w2065_
	);
	LUT2 #(
		.INIT('h2)
	) name1292 (
		\g35_pad ,
		\g979_reg/NET0131 ,
		_w2066_
	);
	LUT2 #(
		.INIT('h1)
	) name1293 (
		\g19334_pad ,
		\g7916_pad ,
		_w2067_
	);
	LUT2 #(
		.INIT('h4)
	) name1294 (
		\g990_reg/NET0131 ,
		_w2067_,
		_w2068_
	);
	LUT2 #(
		.INIT('h2)
	) name1295 (
		\g12919_pad ,
		_w2068_,
		_w2069_
	);
	LUT2 #(
		.INIT('h8)
	) name1296 (
		\g1052_reg/NET0131 ,
		_w2069_,
		_w2070_
	);
	LUT2 #(
		.INIT('h8)
	) name1297 (
		\g1061_reg/NET0131 ,
		_w2070_,
		_w2071_
	);
	LUT2 #(
		.INIT('h1)
	) name1298 (
		\g1061_reg/NET0131 ,
		_w2070_,
		_w2072_
	);
	LUT2 #(
		.INIT('h2)
	) name1299 (
		_w2066_,
		_w2071_,
		_w2073_
	);
	LUT2 #(
		.INIT('h4)
	) name1300 (
		_w2072_,
		_w2073_,
		_w2074_
	);
	LUT2 #(
		.INIT('h1)
	) name1301 (
		_w2065_,
		_w2074_,
		_w2075_
	);
	LUT2 #(
		.INIT('h2)
	) name1302 (
		\g1579_reg/NET0131 ,
		\g35_pad ,
		_w2076_
	);
	LUT2 #(
		.INIT('h1)
	) name1303 (
		_w2003_,
		_w2076_,
		_w2077_
	);
	LUT2 #(
		.INIT('h2)
	) name1304 (
		\g781_reg/NET0131 ,
		_w966_,
		_w2078_
	);
	LUT2 #(
		.INIT('h8)
	) name1305 (
		_w997_,
		_w2078_,
		_w2079_
	);
	LUT2 #(
		.INIT('h4)
	) name1306 (
		\g790_reg/NET0131 ,
		_w2079_,
		_w2080_
	);
	LUT2 #(
		.INIT('h2)
	) name1307 (
		\g35_pad ,
		_w2080_,
		_w2081_
	);
	LUT2 #(
		.INIT('h2)
	) name1308 (
		\g785_reg/NET0131 ,
		_w2081_,
		_w2082_
	);
	LUT2 #(
		.INIT('h8)
	) name1309 (
		\g785_reg/NET0131 ,
		_w2079_,
		_w2083_
	);
	LUT2 #(
		.INIT('h8)
	) name1310 (
		\g790_reg/NET0131 ,
		_w967_,
		_w2084_
	);
	LUT2 #(
		.INIT('h4)
	) name1311 (
		_w2083_,
		_w2084_,
		_w2085_
	);
	LUT2 #(
		.INIT('h1)
	) name1312 (
		_w2082_,
		_w2085_,
		_w2086_
	);
	LUT2 #(
		.INIT('h2)
	) name1313 (
		\g35_pad ,
		_w2023_,
		_w2087_
	);
	LUT2 #(
		.INIT('h2)
	) name1314 (
		\g160_reg/NET0131 ,
		_w2087_,
		_w2088_
	);
	LUT2 #(
		.INIT('h1)
	) name1315 (
		\g4480_reg/NET0131 ,
		_w1085_,
		_w2089_
	);
	LUT2 #(
		.INIT('h4)
	) name1316 (
		\g1052_reg/NET0131 ,
		\g12919_pad ,
		_w2090_
	);
	LUT2 #(
		.INIT('h8)
	) name1317 (
		\g19334_pad ,
		_w2090_,
		_w2091_
	);
	LUT2 #(
		.INIT('h2)
	) name1318 (
		\g35_pad ,
		_w2091_,
		_w2092_
	);
	LUT2 #(
		.INIT('h1)
	) name1319 (
		\g1061_reg/NET0131 ,
		_w2092_,
		_w2093_
	);
	LUT2 #(
		.INIT('h2)
	) name1320 (
		\g1061_reg/NET0131 ,
		\g12919_pad ,
		_w2094_
	);
	LUT2 #(
		.INIT('h8)
	) name1321 (
		\g19334_pad ,
		\g35_pad ,
		_w2095_
	);
	LUT2 #(
		.INIT('h8)
	) name1322 (
		_w2094_,
		_w2095_,
		_w2096_
	);
	LUT2 #(
		.INIT('h1)
	) name1323 (
		_w2093_,
		_w2096_,
		_w2097_
	);
	LUT2 #(
		.INIT('h1)
	) name1324 (
		_w2030_,
		_w2035_,
		_w2098_
	);
	LUT2 #(
		.INIT('h8)
	) name1325 (
		\g225_reg/NET0131 ,
		_w2098_,
		_w2099_
	);
	LUT2 #(
		.INIT('h1)
	) name1326 (
		\g225_reg/NET0131 ,
		_w2098_,
		_w2100_
	);
	LUT2 #(
		.INIT('h1)
	) name1327 (
		_w2099_,
		_w2100_,
		_w2101_
	);
	LUT2 #(
		.INIT('h1)
	) name1328 (
		_w2028_,
		_w2037_,
		_w2102_
	);
	LUT2 #(
		.INIT('h8)
	) name1329 (
		_w2101_,
		_w2102_,
		_w2103_
	);
	LUT2 #(
		.INIT('h1)
	) name1330 (
		_w2101_,
		_w2102_,
		_w2104_
	);
	LUT2 #(
		.INIT('h1)
	) name1331 (
		_w2103_,
		_w2104_,
		_w2105_
	);
	LUT2 #(
		.INIT('h1)
	) name1332 (
		_w2029_,
		_w2036_,
		_w2106_
	);
	LUT2 #(
		.INIT('h8)
	) name1333 (
		_w975_,
		_w987_,
		_w2107_
	);
	LUT2 #(
		.INIT('h8)
	) name1334 (
		_w983_,
		_w2107_,
		_w2108_
	);
	LUT2 #(
		.INIT('h2)
	) name1335 (
		\g732_reg/NET0131 ,
		_w2108_,
		_w2109_
	);
	LUT2 #(
		.INIT('h8)
	) name1336 (
		_w2106_,
		_w2109_,
		_w2110_
	);
	LUT2 #(
		.INIT('h1)
	) name1337 (
		_w2106_,
		_w2109_,
		_w2111_
	);
	LUT2 #(
		.INIT('h1)
	) name1338 (
		_w2110_,
		_w2111_,
		_w2112_
	);
	LUT2 #(
		.INIT('h4)
	) name1339 (
		_w2105_,
		_w2112_,
		_w2113_
	);
	LUT2 #(
		.INIT('h2)
	) name1340 (
		_w2105_,
		_w2112_,
		_w2114_
	);
	LUT2 #(
		.INIT('h2)
	) name1341 (
		\g35_pad ,
		_w2113_,
		_w2115_
	);
	LUT2 #(
		.INIT('h4)
	) name1342 (
		_w2114_,
		_w2115_,
		_w2116_
	);
	LUT2 #(
		.INIT('h2)
	) name1343 (
		_w2014_,
		_w2016_,
		_w2117_
	);
	LUT2 #(
		.INIT('h4)
	) name1344 (
		\g157_reg/NET0131 ,
		_w2010_,
		_w2118_
	);
	LUT2 #(
		.INIT('h8)
	) name1345 (
		_w2117_,
		_w2118_,
		_w2119_
	);
	LUT2 #(
		.INIT('h2)
	) name1346 (
		\g35_pad ,
		_w2119_,
		_w2120_
	);
	LUT2 #(
		.INIT('h2)
	) name1347 (
		\g153_reg/NET0131 ,
		_w2120_,
		_w2121_
	);
	LUT2 #(
		.INIT('h2)
	) name1348 (
		\g157_reg/NET0131 ,
		_w2019_,
		_w2122_
	);
	LUT2 #(
		.INIT('h8)
	) name1349 (
		_w2024_,
		_w2122_,
		_w2123_
	);
	LUT2 #(
		.INIT('h1)
	) name1350 (
		_w2121_,
		_w2123_,
		_w2124_
	);
	LUT2 #(
		.INIT('h1)
	) name1351 (
		_w998_,
		_w2079_,
		_w2125_
	);
	LUT2 #(
		.INIT('h1)
	) name1352 (
		_w2083_,
		_w2125_,
		_w2126_
	);
	LUT2 #(
		.INIT('h2)
	) name1353 (
		\g35_pad ,
		_w2126_,
		_w2127_
	);
	LUT2 #(
		.INIT('h1)
	) name1354 (
		\g35_pad ,
		\g781_reg/NET0131 ,
		_w2128_
	);
	LUT2 #(
		.INIT('h1)
	) name1355 (
		_w2127_,
		_w2128_,
		_w2129_
	);
	LUT2 #(
		.INIT('h1)
	) name1356 (
		\g1052_reg/NET0131 ,
		_w2069_,
		_w2130_
	);
	LUT2 #(
		.INIT('h2)
	) name1357 (
		_w2066_,
		_w2070_,
		_w2131_
	);
	LUT2 #(
		.INIT('h4)
	) name1358 (
		_w2130_,
		_w2131_,
		_w2132_
	);
	LUT2 #(
		.INIT('h1)
	) name1359 (
		\g4438_reg/NET0131 ,
		\g4443_reg/NET0131 ,
		_w2133_
	);
	LUT2 #(
		.INIT('h1)
	) name1360 (
		\g4452_reg/NET0131 ,
		\g7245_pad ,
		_w2134_
	);
	LUT2 #(
		.INIT('h4)
	) name1361 (
		\g7260_pad ,
		_w2134_,
		_w2135_
	);
	LUT2 #(
		.INIT('h8)
	) name1362 (
		_w2133_,
		_w2135_,
		_w2136_
	);
	LUT2 #(
		.INIT('h8)
	) name1363 (
		\g4392_reg/NET0131 ,
		_w2136_,
		_w2137_
	);
	LUT2 #(
		.INIT('h2)
	) name1364 (
		\g35_pad ,
		_w2137_,
		_w2138_
	);
	LUT2 #(
		.INIT('h2)
	) name1365 (
		\g4434_reg/NET0131 ,
		_w2138_,
		_w2139_
	);
	LUT2 #(
		.INIT('h8)
	) name1366 (
		\g35_pad ,
		\g4443_reg/NET0131 ,
		_w2140_
	);
	LUT2 #(
		.INIT('h1)
	) name1367 (
		_w2139_,
		_w2140_,
		_w2141_
	);
	LUT2 #(
		.INIT('h2)
	) name1368 (
		\g329_reg/NET0131 ,
		\g35_pad ,
		_w2142_
	);
	LUT2 #(
		.INIT('h4)
	) name1369 (
		\g305_reg/NET0131 ,
		\g324_reg/NET0131 ,
		_w2143_
	);
	LUT2 #(
		.INIT('h1)
	) name1370 (
		\g311_reg/NET0131 ,
		\g324_reg/NET0131 ,
		_w2144_
	);
	LUT2 #(
		.INIT('h1)
	) name1371 (
		_w2143_,
		_w2144_,
		_w2145_
	);
	LUT2 #(
		.INIT('h2)
	) name1372 (
		\g311_reg/NET0131 ,
		\g336_reg/NET0131 ,
		_w2146_
	);
	LUT2 #(
		.INIT('h8)
	) name1373 (
		\g305_reg/NET0131 ,
		\g336_reg/NET0131 ,
		_w2147_
	);
	LUT2 #(
		.INIT('h1)
	) name1374 (
		\g319_reg/NET0131 ,
		_w2146_,
		_w2148_
	);
	LUT2 #(
		.INIT('h4)
	) name1375 (
		_w2147_,
		_w2148_,
		_w2149_
	);
	LUT2 #(
		.INIT('h2)
	) name1376 (
		_w2145_,
		_w2149_,
		_w2150_
	);
	LUT2 #(
		.INIT('h1)
	) name1377 (
		\g305_reg/NET0131 ,
		\g311_reg/NET0131 ,
		_w2151_
	);
	LUT2 #(
		.INIT('h1)
	) name1378 (
		\g319_reg/NET0131 ,
		\g329_reg/NET0131 ,
		_w2152_
	);
	LUT2 #(
		.INIT('h8)
	) name1379 (
		_w2151_,
		_w2152_,
		_w2153_
	);
	LUT2 #(
		.INIT('h1)
	) name1380 (
		_w2150_,
		_w2153_,
		_w2154_
	);
	LUT2 #(
		.INIT('h2)
	) name1381 (
		\g35_pad ,
		_w2154_,
		_w2155_
	);
	LUT2 #(
		.INIT('h1)
	) name1382 (
		_w2142_,
		_w2155_,
		_w2156_
	);
	LUT2 #(
		.INIT('h2)
	) name1383 (
		\g4621_reg/NET0131 ,
		\g4639_reg/NET0131 ,
		_w2157_
	);
	LUT2 #(
		.INIT('h8)
	) name1384 (
		\g4628_reg/NET0131 ,
		_w2157_,
		_w2158_
	);
	LUT2 #(
		.INIT('h8)
	) name1385 (
		\g4340_reg/NET0131 ,
		\g4349_reg/NET0131 ,
		_w2159_
	);
	LUT2 #(
		.INIT('h8)
	) name1386 (
		\g4358_reg/NET0131 ,
		_w2159_,
		_w2160_
	);
	LUT2 #(
		.INIT('h8)
	) name1387 (
		_w2158_,
		_w2160_,
		_w2161_
	);
	LUT2 #(
		.INIT('h8)
	) name1388 (
		\g4322_reg/NET0131 ,
		\g4332_reg/NET0131 ,
		_w2162_
	);
	LUT2 #(
		.INIT('h8)
	) name1389 (
		_w2161_,
		_w2162_,
		_w2163_
	);
	LUT2 #(
		.INIT('h8)
	) name1390 (
		\g4584_reg/NET0131 ,
		_w2163_,
		_w2164_
	);
	LUT2 #(
		.INIT('h8)
	) name1391 (
		\g4593_reg/NET0131 ,
		_w2164_,
		_w2165_
	);
	LUT2 #(
		.INIT('h8)
	) name1392 (
		\g4601_reg/NET0131 ,
		_w2165_,
		_w2166_
	);
	LUT2 #(
		.INIT('h8)
	) name1393 (
		\g4608_reg/NET0131 ,
		_w2166_,
		_w2167_
	);
	LUT2 #(
		.INIT('h8)
	) name1394 (
		\g4616_reg/NET0131 ,
		_w2164_,
		_w2168_
	);
	LUT2 #(
		.INIT('h2)
	) name1395 (
		\g35_pad ,
		_w2168_,
		_w2169_
	);
	LUT2 #(
		.INIT('h4)
	) name1396 (
		_w2167_,
		_w2169_,
		_w2170_
	);
	LUT2 #(
		.INIT('h8)
	) name1397 (
		\g4616_reg/NET0131 ,
		_w2170_,
		_w2171_
	);
	LUT2 #(
		.INIT('h4)
	) name1398 (
		\g4616_reg/NET0131 ,
		_w2166_,
		_w2172_
	);
	LUT2 #(
		.INIT('h2)
	) name1399 (
		\g35_pad ,
		_w2172_,
		_w2173_
	);
	LUT2 #(
		.INIT('h2)
	) name1400 (
		\g4608_reg/NET0131 ,
		_w2173_,
		_w2174_
	);
	LUT2 #(
		.INIT('h1)
	) name1401 (
		_w2171_,
		_w2174_,
		_w2175_
	);
	LUT2 #(
		.INIT('h8)
	) name1402 (
		\g35_pad ,
		\g4388_reg/NET0131 ,
		_w2176_
	);
	LUT2 #(
		.INIT('h2)
	) name1403 (
		\g4430_reg/NET0131 ,
		_w2176_,
		_w2177_
	);
	LUT2 #(
		.INIT('h4)
	) name1404 (
		\g4430_reg/NET0131 ,
		_w2176_,
		_w2178_
	);
	LUT2 #(
		.INIT('h2)
	) name1405 (
		\g4401_reg/NET0131 ,
		\g4434_reg/NET0131 ,
		_w2179_
	);
	LUT2 #(
		.INIT('h4)
	) name1406 (
		\g4401_reg/NET0131 ,
		\g4434_reg/NET0131 ,
		_w2180_
	);
	LUT2 #(
		.INIT('h1)
	) name1407 (
		_w2179_,
		_w2180_,
		_w2181_
	);
	LUT2 #(
		.INIT('h2)
	) name1408 (
		\g35_pad ,
		_w2181_,
		_w2182_
	);
	LUT2 #(
		.INIT('h1)
	) name1409 (
		_w2177_,
		_w2178_,
		_w2183_
	);
	LUT2 #(
		.INIT('h4)
	) name1410 (
		_w2182_,
		_w2183_,
		_w2184_
	);
	LUT2 #(
		.INIT('h2)
	) name1411 (
		\g1242_reg/NET0131 ,
		\g35_pad ,
		_w2185_
	);
	LUT2 #(
		.INIT('h8)
	) name1412 (
		\g12919_pad ,
		\g35_pad ,
		_w2186_
	);
	LUT2 #(
		.INIT('h1)
	) name1413 (
		_w2185_,
		_w2186_,
		_w2187_
	);
	LUT2 #(
		.INIT('h4)
	) name1414 (
		\g298_reg/NET0131 ,
		_w2047_,
		_w2188_
	);
	LUT2 #(
		.INIT('h2)
	) name1415 (
		\g35_pad ,
		_w2188_,
		_w2189_
	);
	LUT2 #(
		.INIT('h2)
	) name1416 (
		\g294_reg/NET0131 ,
		_w2189_,
		_w2190_
	);
	LUT2 #(
		.INIT('h8)
	) name1417 (
		\g294_reg/NET0131 ,
		_w2047_,
		_w2191_
	);
	LUT2 #(
		.INIT('h8)
	) name1418 (
		\g298_reg/NET0131 ,
		_w2053_,
		_w2192_
	);
	LUT2 #(
		.INIT('h4)
	) name1419 (
		_w2191_,
		_w2192_,
		_w2193_
	);
	LUT2 #(
		.INIT('h1)
	) name1420 (
		_w2190_,
		_w2193_,
		_w2194_
	);
	LUT2 #(
		.INIT('h4)
	) name1421 (
		\g781_reg/NET0131 ,
		_w996_,
		_w2195_
	);
	LUT2 #(
		.INIT('h2)
	) name1422 (
		\g35_pad ,
		_w2195_,
		_w2196_
	);
	LUT2 #(
		.INIT('h2)
	) name1423 (
		\g776_reg/NET0131 ,
		_w2196_,
		_w2197_
	);
	LUT2 #(
		.INIT('h8)
	) name1424 (
		\g35_pad ,
		_w2078_,
		_w2198_
	);
	LUT2 #(
		.INIT('h4)
	) name1425 (
		_w997_,
		_w2198_,
		_w2199_
	);
	LUT2 #(
		.INIT('h1)
	) name1426 (
		_w2197_,
		_w2199_,
		_w2200_
	);
	LUT2 #(
		.INIT('h4)
	) name1427 (
		\g35_pad ,
		\g4423_reg/NET0131 ,
		_w2201_
	);
	LUT2 #(
		.INIT('h1)
	) name1428 (
		\g4372_reg/NET0131 ,
		\g4581_reg/NET0131 ,
		_w2202_
	);
	LUT2 #(
		.INIT('h2)
	) name1429 (
		\g35_pad ,
		_w2202_,
		_w2203_
	);
	LUT2 #(
		.INIT('h1)
	) name1430 (
		_w2201_,
		_w2203_,
		_w2204_
	);
	LUT2 #(
		.INIT('h8)
	) name1431 (
		\g385_reg/NET0131 ,
		_w987_,
		_w2205_
	);
	LUT2 #(
		.INIT('h8)
	) name1432 (
		\g370_reg/NET0131 ,
		_w2205_,
		_w2206_
	);
	LUT2 #(
		.INIT('h8)
	) name1433 (
		\g817_reg/NET0131 ,
		_w2206_,
		_w2207_
	);
	LUT2 #(
		.INIT('h8)
	) name1434 (
		\g832_reg/NET0131 ,
		_w2207_,
		_w2208_
	);
	LUT2 #(
		.INIT('h8)
	) name1435 (
		\g822_reg/NET0131 ,
		_w2208_,
		_w2209_
	);
	LUT2 #(
		.INIT('h8)
	) name1436 (
		\g827_reg/NET0131 ,
		_w2209_,
		_w2210_
	);
	LUT2 #(
		.INIT('h4)
	) name1437 (
		\g812_reg/NET0131 ,
		\g837_reg/NET0131 ,
		_w2211_
	);
	LUT2 #(
		.INIT('h2)
	) name1438 (
		\g847_reg/NET0131 ,
		_w2211_,
		_w2212_
	);
	LUT2 #(
		.INIT('h2)
	) name1439 (
		\g35_pad ,
		_w2212_,
		_w2213_
	);
	LUT2 #(
		.INIT('h4)
	) name1440 (
		_w2210_,
		_w2213_,
		_w2214_
	);
	LUT2 #(
		.INIT('h8)
	) name1441 (
		\g723_reg/NET0131 ,
		_w2214_,
		_w2215_
	);
	LUT2 #(
		.INIT('h1)
	) name1442 (
		\g723_reg/NET0131 ,
		_w2212_,
		_w2216_
	);
	LUT2 #(
		.INIT('h8)
	) name1443 (
		_w2209_,
		_w2216_,
		_w2217_
	);
	LUT2 #(
		.INIT('h2)
	) name1444 (
		\g35_pad ,
		_w2217_,
		_w2218_
	);
	LUT2 #(
		.INIT('h2)
	) name1445 (
		\g827_reg/NET0131 ,
		_w2218_,
		_w2219_
	);
	LUT2 #(
		.INIT('h1)
	) name1446 (
		_w2215_,
		_w2219_,
		_w2220_
	);
	LUT2 #(
		.INIT('h2)
	) name1447 (
		\g3263_reg/NET0131 ,
		\g35_pad ,
		_w2221_
	);
	LUT2 #(
		.INIT('h4)
	) name1448 (
		\g4709_reg/NET0131 ,
		\g4785_reg/NET0131 ,
		_w2222_
	);
	LUT2 #(
		.INIT('h8)
	) name1449 (
		\g4743_reg/NET0131 ,
		_w2222_,
		_w2223_
	);
	LUT2 #(
		.INIT('h8)
	) name1450 (
		_w867_,
		_w2223_,
		_w2224_
	);
	LUT2 #(
		.INIT('h2)
	) name1451 (
		\g4674_reg/NET0131 ,
		_w2224_,
		_w2225_
	);
	LUT2 #(
		.INIT('h1)
	) name1452 (
		\g3333_reg/NET0131 ,
		_w2225_,
		_w2226_
	);
	LUT2 #(
		.INIT('h4)
	) name1453 (
		\g3288_reg/NET0131 ,
		_w912_,
		_w2227_
	);
	LUT2 #(
		.INIT('h8)
	) name1454 (
		\g3288_reg/NET0131 ,
		_w925_,
		_w2228_
	);
	LUT2 #(
		.INIT('h2)
	) name1455 (
		\g3352_reg/NET0131 ,
		_w2227_,
		_w2229_
	);
	LUT2 #(
		.INIT('h4)
	) name1456 (
		_w2228_,
		_w2229_,
		_w2230_
	);
	LUT2 #(
		.INIT('h4)
	) name1457 (
		\g3288_reg/NET0131 ,
		_w941_,
		_w2231_
	);
	LUT2 #(
		.INIT('h8)
	) name1458 (
		\g3288_reg/NET0131 ,
		_w955_,
		_w2232_
	);
	LUT2 #(
		.INIT('h1)
	) name1459 (
		\g3352_reg/NET0131 ,
		_w2231_,
		_w2233_
	);
	LUT2 #(
		.INIT('h4)
	) name1460 (
		_w2232_,
		_w2233_,
		_w2234_
	);
	LUT2 #(
		.INIT('h1)
	) name1461 (
		_w2230_,
		_w2234_,
		_w2235_
	);
	LUT2 #(
		.INIT('h8)
	) name1462 (
		_w2225_,
		_w2235_,
		_w2236_
	);
	LUT2 #(
		.INIT('h2)
	) name1463 (
		\g35_pad ,
		_w2226_,
		_w2237_
	);
	LUT2 #(
		.INIT('h4)
	) name1464 (
		_w2236_,
		_w2237_,
		_w2238_
	);
	LUT2 #(
		.INIT('h1)
	) name1465 (
		_w2221_,
		_w2238_,
		_w2239_
	);
	LUT2 #(
		.INIT('h2)
	) name1466 (
		\g4709_reg/NET0131 ,
		\g4785_reg/NET0131 ,
		_w2240_
	);
	LUT2 #(
		.INIT('h8)
	) name1467 (
		\g4754_reg/NET0131 ,
		_w2240_,
		_w2241_
	);
	LUT2 #(
		.INIT('h8)
	) name1468 (
		_w867_,
		_w2241_,
		_w2242_
	);
	LUT2 #(
		.INIT('h2)
	) name1469 (
		\g4681_reg/NET0131 ,
		_w2242_,
		_w2243_
	);
	LUT2 #(
		.INIT('h1)
	) name1470 (
		\g3684_reg/NET0131 ,
		_w2243_,
		_w2244_
	);
	LUT2 #(
		.INIT('h4)
	) name1471 (
		\g3703_reg/NET0131 ,
		_w955_,
		_w2245_
	);
	LUT2 #(
		.INIT('h8)
	) name1472 (
		\g3703_reg/NET0131 ,
		_w925_,
		_w2246_
	);
	LUT2 #(
		.INIT('h2)
	) name1473 (
		\g3639_reg/NET0131 ,
		_w2245_,
		_w2247_
	);
	LUT2 #(
		.INIT('h4)
	) name1474 (
		_w2246_,
		_w2247_,
		_w2248_
	);
	LUT2 #(
		.INIT('h4)
	) name1475 (
		\g3703_reg/NET0131 ,
		_w941_,
		_w2249_
	);
	LUT2 #(
		.INIT('h8)
	) name1476 (
		\g3703_reg/NET0131 ,
		_w912_,
		_w2250_
	);
	LUT2 #(
		.INIT('h1)
	) name1477 (
		\g3639_reg/NET0131 ,
		_w2249_,
		_w2251_
	);
	LUT2 #(
		.INIT('h4)
	) name1478 (
		_w2250_,
		_w2251_,
		_w2252_
	);
	LUT2 #(
		.INIT('h1)
	) name1479 (
		_w2248_,
		_w2252_,
		_w2253_
	);
	LUT2 #(
		.INIT('h8)
	) name1480 (
		_w2243_,
		_w2253_,
		_w2254_
	);
	LUT2 #(
		.INIT('h2)
	) name1481 (
		\g35_pad ,
		_w2244_,
		_w2255_
	);
	LUT2 #(
		.INIT('h4)
	) name1482 (
		_w2254_,
		_w2255_,
		_w2256_
	);
	LUT2 #(
		.INIT('h1)
	) name1483 (
		_w2221_,
		_w2256_,
		_w2257_
	);
	LUT2 #(
		.INIT('h4)
	) name1484 (
		\g35_pad ,
		\g4477_reg/NET0131 ,
		_w2258_
	);
	LUT2 #(
		.INIT('h1)
	) name1485 (
		_w2203_,
		_w2258_,
		_w2259_
	);
	LUT2 #(
		.INIT('h4)
	) name1486 (
		\g153_reg/NET0131 ,
		_w2012_,
		_w2260_
	);
	LUT2 #(
		.INIT('h8)
	) name1487 (
		_w2017_,
		_w2260_,
		_w2261_
	);
	LUT2 #(
		.INIT('h2)
	) name1488 (
		\g35_pad ,
		_w2261_,
		_w2262_
	);
	LUT2 #(
		.INIT('h2)
	) name1489 (
		\g150_reg/NET0131 ,
		_w2262_,
		_w2263_
	);
	LUT2 #(
		.INIT('h2)
	) name1490 (
		\g153_reg/NET0131 ,
		_w2117_,
		_w2264_
	);
	LUT2 #(
		.INIT('h8)
	) name1491 (
		_w2024_,
		_w2264_,
		_w2265_
	);
	LUT2 #(
		.INIT('h1)
	) name1492 (
		_w2263_,
		_w2265_,
		_w2266_
	);
	LUT2 #(
		.INIT('h1)
	) name1493 (
		\g776_reg/NET0131 ,
		_w966_,
		_w2267_
	);
	LUT2 #(
		.INIT('h8)
	) name1494 (
		_w995_,
		_w2267_,
		_w2268_
	);
	LUT2 #(
		.INIT('h2)
	) name1495 (
		\g35_pad ,
		_w2268_,
		_w2269_
	);
	LUT2 #(
		.INIT('h2)
	) name1496 (
		\g772_reg/NET0131 ,
		_w2269_,
		_w2270_
	);
	LUT2 #(
		.INIT('h8)
	) name1497 (
		\g776_reg/NET0131 ,
		_w967_,
		_w2271_
	);
	LUT2 #(
		.INIT('h4)
	) name1498 (
		_w996_,
		_w2271_,
		_w2272_
	);
	LUT2 #(
		.INIT('h1)
	) name1499 (
		_w2270_,
		_w2272_,
		_w2273_
	);
	LUT2 #(
		.INIT('h2)
	) name1500 (
		\g1236_reg/NET0131 ,
		\g35_pad ,
		_w2274_
	);
	LUT2 #(
		.INIT('h1)
	) name1501 (
		_w2186_,
		_w2274_,
		_w2275_
	);
	LUT2 #(
		.INIT('h2)
	) name1502 (
		\g1554_reg/NET0131 ,
		\g35_pad ,
		_w2276_
	);
	LUT2 #(
		.INIT('h8)
	) name1503 (
		\g35_pad ,
		\g496_reg/NET0131 ,
		_w2277_
	);
	LUT2 #(
		.INIT('h1)
	) name1504 (
		_w2276_,
		_w2277_,
		_w2278_
	);
	LUT2 #(
		.INIT('h4)
	) name1505 (
		\g35_pad ,
		\g4601_reg/NET0131 ,
		_w2279_
	);
	LUT2 #(
		.INIT('h1)
	) name1506 (
		\g4608_reg/NET0131 ,
		_w2166_,
		_w2280_
	);
	LUT2 #(
		.INIT('h2)
	) name1507 (
		_w2170_,
		_w2280_,
		_w2281_
	);
	LUT2 #(
		.INIT('h1)
	) name1508 (
		_w2279_,
		_w2281_,
		_w2282_
	);
	LUT2 #(
		.INIT('h1)
	) name1509 (
		\g4035_reg/NET0131 ,
		_w890_,
		_w2283_
	);
	LUT2 #(
		.INIT('h8)
	) name1510 (
		_w890_,
		_w959_,
		_w2284_
	);
	LUT2 #(
		.INIT('h2)
	) name1511 (
		\g35_pad ,
		_w2283_,
		_w2285_
	);
	LUT2 #(
		.INIT('h4)
	) name1512 (
		_w2284_,
		_w2285_,
		_w2286_
	);
	LUT2 #(
		.INIT('h1)
	) name1513 (
		_w2221_,
		_w2286_,
		_w2287_
	);
	LUT2 #(
		.INIT('h2)
	) name1514 (
		\g29219_pad ,
		\g35_pad ,
		_w2288_
	);
	LUT2 #(
		.INIT('h1)
	) name1515 (
		\g2748_reg/NET0131 ,
		\g2756_reg/NET0131 ,
		_w2289_
	);
	LUT2 #(
		.INIT('h8)
	) name1516 (
		\g2741_reg/NET0131 ,
		_w2289_,
		_w2290_
	);
	LUT2 #(
		.INIT('h2)
	) name1517 (
		\g35_pad ,
		_w2290_,
		_w2291_
	);
	LUT2 #(
		.INIT('h8)
	) name1518 (
		\g2735_reg/NET0131 ,
		\g2741_reg/NET0131 ,
		_w2292_
	);
	LUT2 #(
		.INIT('h8)
	) name1519 (
		\g2748_reg/NET0131 ,
		\g2756_reg/NET0131 ,
		_w2293_
	);
	LUT2 #(
		.INIT('h8)
	) name1520 (
		_w2292_,
		_w2293_,
		_w2294_
	);
	LUT2 #(
		.INIT('h1)
	) name1521 (
		_w2289_,
		_w2294_,
		_w2295_
	);
	LUT2 #(
		.INIT('h4)
	) name1522 (
		\g2193_reg/NET0131 ,
		_w2295_,
		_w2296_
	);
	LUT2 #(
		.INIT('h1)
	) name1523 (
		\g2799_reg/NET0131 ,
		_w2296_,
		_w2297_
	);
	LUT2 #(
		.INIT('h2)
	) name1524 (
		_w2291_,
		_w2297_,
		_w2298_
	);
	LUT2 #(
		.INIT('h1)
	) name1525 (
		_w2288_,
		_w2298_,
		_w2299_
	);
	LUT2 #(
		.INIT('h4)
	) name1526 (
		\g294_reg/NET0131 ,
		_w2046_,
		_w2300_
	);
	LUT2 #(
		.INIT('h2)
	) name1527 (
		\g35_pad ,
		_w2300_,
		_w2301_
	);
	LUT2 #(
		.INIT('h2)
	) name1528 (
		\g291_reg/NET0131 ,
		_w2301_,
		_w2302_
	);
	LUT2 #(
		.INIT('h8)
	) name1529 (
		\g294_reg/NET0131 ,
		_w2053_,
		_w2303_
	);
	LUT2 #(
		.INIT('h4)
	) name1530 (
		_w2047_,
		_w2303_,
		_w2304_
	);
	LUT2 #(
		.INIT('h1)
	) name1531 (
		_w2302_,
		_w2304_,
		_w2305_
	);
	LUT2 #(
		.INIT('h1)
	) name1532 (
		_w971_,
		_w995_,
		_w2306_
	);
	LUT2 #(
		.INIT('h8)
	) name1533 (
		\g772_reg/NET0131 ,
		_w995_,
		_w2307_
	);
	LUT2 #(
		.INIT('h1)
	) name1534 (
		_w2306_,
		_w2307_,
		_w2308_
	);
	LUT2 #(
		.INIT('h2)
	) name1535 (
		\g35_pad ,
		_w2308_,
		_w2309_
	);
	LUT2 #(
		.INIT('h1)
	) name1536 (
		\g35_pad ,
		\g767_reg/NET0131 ,
		_w2310_
	);
	LUT2 #(
		.INIT('h1)
	) name1537 (
		_w2309_,
		_w2310_,
		_w2311_
	);
	LUT2 #(
		.INIT('h2)
	) name1538 (
		\g29211_pad ,
		\g35_pad ,
		_w2312_
	);
	LUT2 #(
		.INIT('h2)
	) name1539 (
		\g35_pad ,
		_w2145_,
		_w2313_
	);
	LUT2 #(
		.INIT('h2)
	) name1540 (
		\g329_reg/NET0131 ,
		\g341_reg/NET0131 ,
		_w2314_
	);
	LUT2 #(
		.INIT('h8)
	) name1541 (
		_w2313_,
		_w2314_,
		_w2315_
	);
	LUT2 #(
		.INIT('h1)
	) name1542 (
		_w2312_,
		_w2315_,
		_w2316_
	);
	LUT2 #(
		.INIT('h4)
	) name1543 (
		\g35_pad ,
		\g822_reg/NET0131 ,
		_w2317_
	);
	LUT2 #(
		.INIT('h1)
	) name1544 (
		\g827_reg/NET0131 ,
		_w2209_,
		_w2318_
	);
	LUT2 #(
		.INIT('h2)
	) name1545 (
		_w2214_,
		_w2318_,
		_w2319_
	);
	LUT2 #(
		.INIT('h1)
	) name1546 (
		_w2317_,
		_w2319_,
		_w2320_
	);
	LUT2 #(
		.INIT('h2)
	) name1547 (
		\g164_reg/NET0131 ,
		\g35_pad ,
		_w2321_
	);
	LUT2 #(
		.INIT('h4)
	) name1548 (
		\g150_reg/NET0131 ,
		_w2013_,
		_w2322_
	);
	LUT2 #(
		.INIT('h2)
	) name1549 (
		\g150_reg/NET0131 ,
		_w2012_,
		_w2323_
	);
	LUT2 #(
		.INIT('h8)
	) name1550 (
		_w2017_,
		_w2323_,
		_w2324_
	);
	LUT2 #(
		.INIT('h1)
	) name1551 (
		_w2322_,
		_w2324_,
		_w2325_
	);
	LUT2 #(
		.INIT('h2)
	) name1552 (
		\g35_pad ,
		_w2325_,
		_w2326_
	);
	LUT2 #(
		.INIT('h1)
	) name1553 (
		_w2321_,
		_w2326_,
		_w2327_
	);
	LUT2 #(
		.INIT('h2)
	) name1554 (
		\g35_pad ,
		_w2225_,
		_w2328_
	);
	LUT2 #(
		.INIT('h8)
	) name1555 (
		\g4749_reg/NET0131 ,
		_w2328_,
		_w2329_
	);
	LUT2 #(
		.INIT('h8)
	) name1556 (
		\g4793_reg/NET0131 ,
		_w863_,
		_w2330_
	);
	LUT2 #(
		.INIT('h8)
	) name1557 (
		_w861_,
		_w2330_,
		_w2331_
	);
	LUT2 #(
		.INIT('h8)
	) name1558 (
		\g35_pad ,
		_w2225_,
		_w2332_
	);
	LUT2 #(
		.INIT('h2)
	) name1559 (
		\g3343_reg/NET0131 ,
		\g3352_reg/NET0131 ,
		_w2333_
	);
	LUT2 #(
		.INIT('h8)
	) name1560 (
		\g3347_reg/NET0131 ,
		\g3352_reg/NET0131 ,
		_w2334_
	);
	LUT2 #(
		.INIT('h1)
	) name1561 (
		_w2333_,
		_w2334_,
		_w2335_
	);
	LUT2 #(
		.INIT('h2)
	) name1562 (
		\g3288_reg/NET0131 ,
		_w2335_,
		_w2336_
	);
	LUT2 #(
		.INIT('h4)
	) name1563 (
		\g3288_reg/NET0131 ,
		_w2335_,
		_w2337_
	);
	LUT2 #(
		.INIT('h1)
	) name1564 (
		\g4749_reg/NET0131 ,
		_w2336_,
		_w2338_
	);
	LUT2 #(
		.INIT('h4)
	) name1565 (
		_w2337_,
		_w2338_,
		_w2339_
	);
	LUT2 #(
		.INIT('h2)
	) name1566 (
		_w2331_,
		_w2339_,
		_w2340_
	);
	LUT2 #(
		.INIT('h8)
	) name1567 (
		_w2332_,
		_w2340_,
		_w2341_
	);
	LUT2 #(
		.INIT('h1)
	) name1568 (
		_w2329_,
		_w2341_,
		_w2342_
	);
	LUT2 #(
		.INIT('h8)
	) name1569 (
		\g4771_reg/NET0131 ,
		_w891_,
		_w2343_
	);
	LUT2 #(
		.INIT('h8)
	) name1570 (
		_w2240_,
		_w2330_,
		_w2344_
	);
	LUT2 #(
		.INIT('h2)
	) name1571 (
		\g3343_reg/NET0131 ,
		\g4054_reg/NET0131 ,
		_w2345_
	);
	LUT2 #(
		.INIT('h8)
	) name1572 (
		\g3347_reg/NET0131 ,
		\g4054_reg/NET0131 ,
		_w2346_
	);
	LUT2 #(
		.INIT('h1)
	) name1573 (
		_w2345_,
		_w2346_,
		_w2347_
	);
	LUT2 #(
		.INIT('h2)
	) name1574 (
		\g3990_reg/NET0131 ,
		_w2347_,
		_w2348_
	);
	LUT2 #(
		.INIT('h4)
	) name1575 (
		\g3990_reg/NET0131 ,
		_w2347_,
		_w2349_
	);
	LUT2 #(
		.INIT('h1)
	) name1576 (
		\g4771_reg/NET0131 ,
		_w2348_,
		_w2350_
	);
	LUT2 #(
		.INIT('h4)
	) name1577 (
		_w2349_,
		_w2350_,
		_w2351_
	);
	LUT2 #(
		.INIT('h2)
	) name1578 (
		_w2344_,
		_w2351_,
		_w2352_
	);
	LUT2 #(
		.INIT('h8)
	) name1579 (
		_w893_,
		_w2352_,
		_w2353_
	);
	LUT2 #(
		.INIT('h1)
	) name1580 (
		_w2343_,
		_w2353_,
		_w2354_
	);
	LUT2 #(
		.INIT('h8)
	) name1581 (
		_w980_,
		_w2015_,
		_w2355_
	);
	LUT2 #(
		.INIT('h2)
	) name1582 (
		\g739_reg/NET0131 ,
		_w966_,
		_w2356_
	);
	LUT2 #(
		.INIT('h8)
	) name1583 (
		_w2355_,
		_w2356_,
		_w2357_
	);
	LUT2 #(
		.INIT('h8)
	) name1584 (
		\g744_reg/NET0131 ,
		_w2357_,
		_w2358_
	);
	LUT2 #(
		.INIT('h8)
	) name1585 (
		_w986_,
		_w2358_,
		_w2359_
	);
	LUT2 #(
		.INIT('h1)
	) name1586 (
		\g767_reg/NET0131 ,
		_w966_,
		_w2360_
	);
	LUT2 #(
		.INIT('h8)
	) name1587 (
		_w2359_,
		_w2360_,
		_w2361_
	);
	LUT2 #(
		.INIT('h2)
	) name1588 (
		\g35_pad ,
		_w2361_,
		_w2362_
	);
	LUT2 #(
		.INIT('h2)
	) name1589 (
		\g763_reg/NET0131 ,
		_w2362_,
		_w2363_
	);
	LUT2 #(
		.INIT('h8)
	) name1590 (
		\g763_reg/NET0131 ,
		_w2359_,
		_w2364_
	);
	LUT2 #(
		.INIT('h8)
	) name1591 (
		\g767_reg/NET0131 ,
		_w967_,
		_w2365_
	);
	LUT2 #(
		.INIT('h4)
	) name1592 (
		_w2364_,
		_w2365_,
		_w2366_
	);
	LUT2 #(
		.INIT('h1)
	) name1593 (
		_w2363_,
		_w2366_,
		_w2367_
	);
	LUT2 #(
		.INIT('h8)
	) name1594 (
		\g1152_reg/NET0131 ,
		_w1344_,
		_w2368_
	);
	LUT2 #(
		.INIT('h2)
	) name1595 (
		\g1146_reg/NET0131 ,
		_w2368_,
		_w2369_
	);
	LUT2 #(
		.INIT('h4)
	) name1596 (
		\g1099_reg/NET0131 ,
		_w1344_,
		_w2370_
	);
	LUT2 #(
		.INIT('h1)
	) name1597 (
		_w2369_,
		_w2370_,
		_w2371_
	);
	LUT2 #(
		.INIT('h2)
	) name1598 (
		\g35_pad ,
		_w2371_,
		_w2372_
	);
	LUT2 #(
		.INIT('h1)
	) name1599 (
		\g979_reg/NET0131 ,
		\g990_reg/NET0131 ,
		_w2373_
	);
	LUT2 #(
		.INIT('h2)
	) name1600 (
		\g979_reg/NET0131 ,
		\g996_reg/NET0131 ,
		_w2374_
	);
	LUT2 #(
		.INIT('h4)
	) name1601 (
		\g979_reg/NET0131 ,
		\g996_reg/NET0131 ,
		_w2375_
	);
	LUT2 #(
		.INIT('h1)
	) name1602 (
		_w2374_,
		_w2375_,
		_w2376_
	);
	LUT2 #(
		.INIT('h1)
	) name1603 (
		_w2373_,
		_w2376_,
		_w2377_
	);
	LUT2 #(
		.INIT('h8)
	) name1604 (
		_w815_,
		_w2377_,
		_w2378_
	);
	LUT2 #(
		.INIT('h2)
	) name1605 (
		\g1236_reg/NET0131 ,
		\g979_reg/NET0131 ,
		_w2379_
	);
	LUT2 #(
		.INIT('h4)
	) name1606 (
		\g1236_reg/NET0131 ,
		\g979_reg/NET0131 ,
		_w2380_
	);
	LUT2 #(
		.INIT('h1)
	) name1607 (
		_w2379_,
		_w2380_,
		_w2381_
	);
	LUT2 #(
		.INIT('h2)
	) name1608 (
		_w2378_,
		_w2381_,
		_w2382_
	);
	LUT2 #(
		.INIT('h1)
	) name1609 (
		\g13259_pad ,
		\g8416_pad ,
		_w2383_
	);
	LUT2 #(
		.INIT('h8)
	) name1610 (
		_w2067_,
		_w2383_,
		_w2384_
	);
	LUT2 #(
		.INIT('h2)
	) name1611 (
		_w2382_,
		_w2384_,
		_w2385_
	);
	LUT2 #(
		.INIT('h2)
	) name1612 (
		\g990_reg/NET0131 ,
		_w2382_,
		_w2386_
	);
	LUT2 #(
		.INIT('h4)
	) name1613 (
		\g990_reg/NET0131 ,
		_w2382_,
		_w2387_
	);
	LUT2 #(
		.INIT('h1)
	) name1614 (
		_w2386_,
		_w2387_,
		_w2388_
	);
	LUT2 #(
		.INIT('h8)
	) name1615 (
		_w2384_,
		_w2388_,
		_w2389_
	);
	LUT2 #(
		.INIT('h1)
	) name1616 (
		_w2385_,
		_w2389_,
		_w2390_
	);
	LUT2 #(
		.INIT('h2)
	) name1617 (
		\g35_pad ,
		_w2390_,
		_w2391_
	);
	LUT2 #(
		.INIT('h4)
	) name1618 (
		\g35_pad ,
		\g996_reg/NET0131 ,
		_w2392_
	);
	LUT2 #(
		.INIT('h1)
	) name1619 (
		_w2391_,
		_w2392_,
		_w2393_
	);
	LUT2 #(
		.INIT('h4)
	) name1620 (
		\g35_pad ,
		\g4664_reg/NET0131 ,
		_w2394_
	);
	LUT2 #(
		.INIT('h8)
	) name1621 (
		\g4653_reg/NET0131 ,
		\g4688_reg/NET0131 ,
		_w2395_
	);
	LUT2 #(
		.INIT('h8)
	) name1622 (
		_w865_,
		_w2395_,
		_w2396_
	);
	LUT2 #(
		.INIT('h2)
	) name1623 (
		\g35_pad ,
		_w2396_,
		_w2397_
	);
	LUT2 #(
		.INIT('h8)
	) name1624 (
		\g4659_reg/NET0131 ,
		_w2395_,
		_w2398_
	);
	LUT2 #(
		.INIT('h8)
	) name1625 (
		\g4664_reg/NET0131 ,
		_w2398_,
		_w2399_
	);
	LUT2 #(
		.INIT('h1)
	) name1626 (
		\g4669_reg/NET0131 ,
		_w2399_,
		_w2400_
	);
	LUT2 #(
		.INIT('h2)
	) name1627 (
		_w2397_,
		_w2400_,
		_w2401_
	);
	LUT2 #(
		.INIT('h1)
	) name1628 (
		_w2394_,
		_w2401_,
		_w2402_
	);
	LUT2 #(
		.INIT('h2)
	) name1629 (
		\g283_reg/NET0131 ,
		\g291_reg/NET0131 ,
		_w2403_
	);
	LUT2 #(
		.INIT('h8)
	) name1630 (
		_w2044_,
		_w2403_,
		_w2404_
	);
	LUT2 #(
		.INIT('h2)
	) name1631 (
		\g35_pad ,
		_w2404_,
		_w2405_
	);
	LUT2 #(
		.INIT('h2)
	) name1632 (
		\g287_reg/NET0131 ,
		_w2405_,
		_w2406_
	);
	LUT2 #(
		.INIT('h2)
	) name1633 (
		\g291_reg/NET0131 ,
		_w2046_,
		_w2407_
	);
	LUT2 #(
		.INIT('h8)
	) name1634 (
		_w2053_,
		_w2407_,
		_w2408_
	);
	LUT2 #(
		.INIT('h1)
	) name1635 (
		_w2406_,
		_w2408_,
		_w2409_
	);
	LUT2 #(
		.INIT('h2)
	) name1636 (
		\g763_reg/NET0131 ,
		_w966_,
		_w2410_
	);
	LUT2 #(
		.INIT('h1)
	) name1637 (
		_w2359_,
		_w2410_,
		_w2411_
	);
	LUT2 #(
		.INIT('h1)
	) name1638 (
		_w2364_,
		_w2411_,
		_w2412_
	);
	LUT2 #(
		.INIT('h2)
	) name1639 (
		\g35_pad ,
		_w2412_,
		_w2413_
	);
	LUT2 #(
		.INIT('h1)
	) name1640 (
		\g35_pad ,
		\g758_reg/NET0131 ,
		_w2414_
	);
	LUT2 #(
		.INIT('h1)
	) name1641 (
		_w2413_,
		_w2414_,
		_w2415_
	);
	LUT2 #(
		.INIT('h8)
	) name1642 (
		\g35_pad ,
		\g956_reg/NET0131 ,
		_w2416_
	);
	LUT2 #(
		.INIT('h2)
	) name1643 (
		\g1099_reg/NET0131 ,
		\g1152_reg/NET0131 ,
		_w2417_
	);
	LUT2 #(
		.INIT('h8)
	) name1644 (
		_w1344_,
		_w2417_,
		_w2418_
	);
	LUT2 #(
		.INIT('h2)
	) name1645 (
		\g35_pad ,
		_w2418_,
		_w2419_
	);
	LUT2 #(
		.INIT('h2)
	) name1646 (
		\g1141_reg/NET0131 ,
		_w2419_,
		_w2420_
	);
	LUT2 #(
		.INIT('h2)
	) name1647 (
		_w2416_,
		_w2420_,
		_w2421_
	);
	LUT2 #(
		.INIT('h4)
	) name1648 (
		_w2416_,
		_w2420_,
		_w2422_
	);
	LUT2 #(
		.INIT('h1)
	) name1649 (
		_w2421_,
		_w2422_,
		_w2423_
	);
	LUT2 #(
		.INIT('h8)
	) name1650 (
		\g1105_reg/NET0131 ,
		\g35_pad ,
		_w2424_
	);
	LUT2 #(
		.INIT('h8)
	) name1651 (
		_w1320_,
		_w2417_,
		_w2425_
	);
	LUT2 #(
		.INIT('h2)
	) name1652 (
		\g35_pad ,
		_w2425_,
		_w2426_
	);
	LUT2 #(
		.INIT('h2)
	) name1653 (
		\g1111_reg/NET0131 ,
		_w2426_,
		_w2427_
	);
	LUT2 #(
		.INIT('h2)
	) name1654 (
		_w2424_,
		_w2427_,
		_w2428_
	);
	LUT2 #(
		.INIT('h4)
	) name1655 (
		_w2424_,
		_w2427_,
		_w2429_
	);
	LUT2 #(
		.INIT('h1)
	) name1656 (
		_w2428_,
		_w2429_,
		_w2430_
	);
	LUT2 #(
		.INIT('h8)
	) name1657 (
		\g1129_reg/NET0131 ,
		\g35_pad ,
		_w2431_
	);
	LUT2 #(
		.INIT('h8)
	) name1658 (
		_w1332_,
		_w2417_,
		_w2432_
	);
	LUT2 #(
		.INIT('h2)
	) name1659 (
		\g35_pad ,
		_w2432_,
		_w2433_
	);
	LUT2 #(
		.INIT('h2)
	) name1660 (
		\g1124_reg/NET0131 ,
		_w2433_,
		_w2434_
	);
	LUT2 #(
		.INIT('h2)
	) name1661 (
		_w2431_,
		_w2434_,
		_w2435_
	);
	LUT2 #(
		.INIT('h4)
	) name1662 (
		_w2431_,
		_w2434_,
		_w2436_
	);
	LUT2 #(
		.INIT('h1)
	) name1663 (
		_w2435_,
		_w2436_,
		_w2437_
	);
	LUT2 #(
		.INIT('h8)
	) name1664 (
		\g1135_reg/NET0131 ,
		\g35_pad ,
		_w2438_
	);
	LUT2 #(
		.INIT('h8)
	) name1665 (
		_w1306_,
		_w2417_,
		_w2439_
	);
	LUT2 #(
		.INIT('h2)
	) name1666 (
		\g35_pad ,
		_w2439_,
		_w2440_
	);
	LUT2 #(
		.INIT('h2)
	) name1667 (
		\g1094_reg/NET0131 ,
		_w2440_,
		_w2441_
	);
	LUT2 #(
		.INIT('h2)
	) name1668 (
		_w2438_,
		_w2441_,
		_w2442_
	);
	LUT2 #(
		.INIT('h4)
	) name1669 (
		_w2438_,
		_w2441_,
		_w2443_
	);
	LUT2 #(
		.INIT('h1)
	) name1670 (
		_w2442_,
		_w2443_,
		_w2444_
	);
	LUT2 #(
		.INIT('h2)
	) name1671 (
		\g35_pad ,
		_w2243_,
		_w2445_
	);
	LUT2 #(
		.INIT('h8)
	) name1672 (
		\g4760_reg/NET0131 ,
		_w2445_,
		_w2446_
	);
	LUT2 #(
		.INIT('h8)
	) name1673 (
		_w2222_,
		_w2330_,
		_w2447_
	);
	LUT2 #(
		.INIT('h8)
	) name1674 (
		\g35_pad ,
		_w2243_,
		_w2448_
	);
	LUT2 #(
		.INIT('h2)
	) name1675 (
		\g3343_reg/NET0131 ,
		\g3703_reg/NET0131 ,
		_w2449_
	);
	LUT2 #(
		.INIT('h8)
	) name1676 (
		\g3347_reg/NET0131 ,
		\g3703_reg/NET0131 ,
		_w2450_
	);
	LUT2 #(
		.INIT('h1)
	) name1677 (
		_w2449_,
		_w2450_,
		_w2451_
	);
	LUT2 #(
		.INIT('h2)
	) name1678 (
		\g3639_reg/NET0131 ,
		_w2451_,
		_w2452_
	);
	LUT2 #(
		.INIT('h4)
	) name1679 (
		\g3639_reg/NET0131 ,
		_w2451_,
		_w2453_
	);
	LUT2 #(
		.INIT('h1)
	) name1680 (
		\g4760_reg/NET0131 ,
		_w2452_,
		_w2454_
	);
	LUT2 #(
		.INIT('h4)
	) name1681 (
		_w2453_,
		_w2454_,
		_w2455_
	);
	LUT2 #(
		.INIT('h2)
	) name1682 (
		_w2447_,
		_w2455_,
		_w2456_
	);
	LUT2 #(
		.INIT('h8)
	) name1683 (
		_w2448_,
		_w2456_,
		_w2457_
	);
	LUT2 #(
		.INIT('h1)
	) name1684 (
		_w2446_,
		_w2457_,
		_w2458_
	);
	LUT2 #(
		.INIT('h4)
	) name1685 (
		\g35_pad ,
		\g676_reg/NET0131 ,
		_w2459_
	);
	LUT2 #(
		.INIT('h8)
	) name1686 (
		\g482_reg/NET0131 ,
		\g490_reg/NET0131 ,
		_w2460_
	);
	LUT2 #(
		.INIT('h2)
	) name1687 (
		\g499_reg/NET0131 ,
		\g504_reg/NET0131 ,
		_w2461_
	);
	LUT2 #(
		.INIT('h4)
	) name1688 (
		\g528_reg/NET0131 ,
		_w2461_,
		_w2462_
	);
	LUT2 #(
		.INIT('h8)
	) name1689 (
		_w2460_,
		_w2462_,
		_w2463_
	);
	LUT2 #(
		.INIT('h8)
	) name1690 (
		_w2206_,
		_w2463_,
		_w2464_
	);
	LUT2 #(
		.INIT('h1)
	) name1691 (
		\g661_reg/NET0131 ,
		\g728_reg/NET0131 ,
		_w2465_
	);
	LUT2 #(
		.INIT('h8)
	) name1692 (
		\g661_reg/NET0131 ,
		\g728_reg/NET0131 ,
		_w2466_
	);
	LUT2 #(
		.INIT('h1)
	) name1693 (
		_w2465_,
		_w2466_,
		_w2467_
	);
	LUT2 #(
		.INIT('h1)
	) name1694 (
		_w973_,
		_w976_,
		_w2468_
	);
	LUT2 #(
		.INIT('h1)
	) name1695 (
		\g645_reg/NET0131 ,
		\g650_reg/NET0131 ,
		_w2469_
	);
	LUT2 #(
		.INIT('h8)
	) name1696 (
		\g681_reg/NET0131 ,
		\g699_reg/NET0131 ,
		_w2470_
	);
	LUT2 #(
		.INIT('h8)
	) name1697 (
		_w2469_,
		_w2470_,
		_w2471_
	);
	LUT2 #(
		.INIT('h4)
	) name1698 (
		_w2467_,
		_w2471_,
		_w2472_
	);
	LUT2 #(
		.INIT('h4)
	) name1699 (
		_w2468_,
		_w2472_,
		_w2473_
	);
	LUT2 #(
		.INIT('h8)
	) name1700 (
		_w2464_,
		_w2473_,
		_w2474_
	);
	LUT2 #(
		.INIT('h8)
	) name1701 (
		\g35_pad ,
		\g703_reg/NET0131 ,
		_w2475_
	);
	LUT2 #(
		.INIT('h4)
	) name1702 (
		_w2474_,
		_w2475_,
		_w2476_
	);
	LUT2 #(
		.INIT('h8)
	) name1703 (
		\g671_reg/NET0131 ,
		_w2464_,
		_w2477_
	);
	LUT2 #(
		.INIT('h8)
	) name1704 (
		\g676_reg/NET0131 ,
		_w2477_,
		_w2478_
	);
	LUT2 #(
		.INIT('h1)
	) name1705 (
		\g714_reg/NET0131 ,
		_w2478_,
		_w2479_
	);
	LUT2 #(
		.INIT('h8)
	) name1706 (
		\g714_reg/NET0131 ,
		_w2478_,
		_w2480_
	);
	LUT2 #(
		.INIT('h2)
	) name1707 (
		_w2476_,
		_w2479_,
		_w2481_
	);
	LUT2 #(
		.INIT('h4)
	) name1708 (
		_w2480_,
		_w2481_,
		_w2482_
	);
	LUT2 #(
		.INIT('h1)
	) name1709 (
		_w2459_,
		_w2482_,
		_w2483_
	);
	LUT2 #(
		.INIT('h4)
	) name1710 (
		\g35_pad ,
		\g4593_reg/NET0131 ,
		_w2484_
	);
	LUT2 #(
		.INIT('h1)
	) name1711 (
		\g4601_reg/NET0131 ,
		_w2165_,
		_w2485_
	);
	LUT2 #(
		.INIT('h4)
	) name1712 (
		_w2166_,
		_w2169_,
		_w2486_
	);
	LUT2 #(
		.INIT('h4)
	) name1713 (
		_w2485_,
		_w2486_,
		_w2487_
	);
	LUT2 #(
		.INIT('h1)
	) name1714 (
		_w2484_,
		_w2487_,
		_w2488_
	);
	LUT2 #(
		.INIT('h8)
	) name1715 (
		\g269_reg/NET0131 ,
		\g35_pad ,
		_w2489_
	);
	LUT2 #(
		.INIT('h2)
	) name1716 (
		\g29215_pad ,
		\g35_pad ,
		_w2490_
	);
	LUT2 #(
		.INIT('h1)
	) name1717 (
		_w2489_,
		_w2490_,
		_w2491_
	);
	LUT2 #(
		.INIT('h2)
	) name1718 (
		\g35_pad ,
		_w1344_,
		_w2492_
	);
	LUT2 #(
		.INIT('h2)
	) name1719 (
		\g1146_reg/NET0131 ,
		_w2492_,
		_w2493_
	);
	LUT2 #(
		.INIT('h8)
	) name1720 (
		\g1152_reg/NET0131 ,
		_w2492_,
		_w2494_
	);
	LUT2 #(
		.INIT('h1)
	) name1721 (
		_w2493_,
		_w2494_,
		_w2495_
	);
	LUT2 #(
		.INIT('h8)
	) name1722 (
		\g29215_pad ,
		\g35_pad ,
		_w2496_
	);
	LUT2 #(
		.INIT('h2)
	) name1723 (
		\g1211_reg/NET0131 ,
		\g35_pad ,
		_w2497_
	);
	LUT2 #(
		.INIT('h1)
	) name1724 (
		_w2496_,
		_w2497_,
		_w2498_
	);
	LUT2 #(
		.INIT('h4)
	) name1725 (
		\g1862_reg/NET0131 ,
		\g1906_reg/NET0131 ,
		_w2499_
	);
	LUT2 #(
		.INIT('h4)
	) name1726 (
		\g2715_reg/NET0131 ,
		\g2719_reg/NET0131 ,
		_w2500_
	);
	LUT2 #(
		.INIT('h1)
	) name1727 (
		\g2724_reg/NET0131 ,
		\g2729_reg/NET0131 ,
		_w2501_
	);
	LUT2 #(
		.INIT('h1)
	) name1728 (
		\g2741_reg/NET0131 ,
		\g2748_reg/NET0131 ,
		_w2502_
	);
	LUT2 #(
		.INIT('h4)
	) name1729 (
		\g2756_reg/NET0131 ,
		_w2502_,
		_w2503_
	);
	LUT2 #(
		.INIT('h8)
	) name1730 (
		\g2735_reg/NET0131 ,
		_w2503_,
		_w2504_
	);
	LUT2 #(
		.INIT('h4)
	) name1731 (
		\g2783_reg/NET0131 ,
		_w2504_,
		_w2505_
	);
	LUT2 #(
		.INIT('h2)
	) name1732 (
		_w2501_,
		_w2505_,
		_w2506_
	);
	LUT2 #(
		.INIT('h2)
	) name1733 (
		_w2500_,
		_w2506_,
		_w2507_
	);
	LUT2 #(
		.INIT('h2)
	) name1734 (
		\g1917_reg/NET0131 ,
		\g1926_reg/NET0131 ,
		_w2508_
	);
	LUT2 #(
		.INIT('h8)
	) name1735 (
		\g35_pad ,
		_w2508_,
		_w2509_
	);
	LUT2 #(
		.INIT('h8)
	) name1736 (
		_w2507_,
		_w2509_,
		_w2510_
	);
	LUT2 #(
		.INIT('h4)
	) name1737 (
		_w2499_,
		_w2510_,
		_w2511_
	);
	LUT2 #(
		.INIT('h1)
	) name1738 (
		\g1882_reg/NET0131 ,
		\g35_pad ,
		_w2512_
	);
	LUT2 #(
		.INIT('h4)
	) name1739 (
		\g1902_reg/NET0131 ,
		\g35_pad ,
		_w2513_
	);
	LUT2 #(
		.INIT('h1)
	) name1740 (
		_w2512_,
		_w2513_,
		_w2514_
	);
	LUT2 #(
		.INIT('h4)
	) name1741 (
		_w2510_,
		_w2514_,
		_w2515_
	);
	LUT2 #(
		.INIT('h1)
	) name1742 (
		_w2511_,
		_w2515_,
		_w2516_
	);
	LUT2 #(
		.INIT('h8)
	) name1743 (
		\g376_reg/NET0131 ,
		\g8719_pad ,
		_w2517_
	);
	LUT2 #(
		.INIT('h2)
	) name1744 (
		\g370_reg/NET0131 ,
		\g385_reg/NET0131 ,
		_w2518_
	);
	LUT2 #(
		.INIT('h8)
	) name1745 (
		_w2517_,
		_w2518_,
		_w2519_
	);
	LUT2 #(
		.INIT('h8)
	) name1746 (
		\g392_reg/NET0131 ,
		\g441_reg/NET0131 ,
		_w2520_
	);
	LUT2 #(
		.INIT('h4)
	) name1747 (
		\g392_reg/NET0131 ,
		\g411_reg/NET0131 ,
		_w2521_
	);
	LUT2 #(
		.INIT('h8)
	) name1748 (
		\g392_reg/NET0131 ,
		\g452_reg/NET0131 ,
		_w2522_
	);
	LUT2 #(
		.INIT('h2)
	) name1749 (
		\g174_reg/NET0131 ,
		\g392_reg/NET0131 ,
		_w2523_
	);
	LUT2 #(
		.INIT('h1)
	) name1750 (
		_w2522_,
		_w2523_,
		_w2524_
	);
	LUT2 #(
		.INIT('h2)
	) name1751 (
		\g182_reg/NET0131 ,
		_w2524_,
		_w2525_
	);
	LUT2 #(
		.INIT('h4)
	) name1752 (
		\g182_reg/NET0131 ,
		_w2524_,
		_w2526_
	);
	LUT2 #(
		.INIT('h1)
	) name1753 (
		\g417_reg/NET0131 ,
		\g691_reg/NET0131 ,
		_w2527_
	);
	LUT2 #(
		.INIT('h4)
	) name1754 (
		_w2520_,
		_w2527_,
		_w2528_
	);
	LUT2 #(
		.INIT('h4)
	) name1755 (
		_w2521_,
		_w2528_,
		_w2529_
	);
	LUT2 #(
		.INIT('h4)
	) name1756 (
		_w2525_,
		_w2529_,
		_w2530_
	);
	LUT2 #(
		.INIT('h4)
	) name1757 (
		_w2526_,
		_w2530_,
		_w2531_
	);
	LUT2 #(
		.INIT('h1)
	) name1758 (
		\g392_reg/NET0131 ,
		\g405_reg/NET0131 ,
		_w2532_
	);
	LUT2 #(
		.INIT('h8)
	) name1759 (
		\g392_reg/NET0131 ,
		\g405_reg/NET0131 ,
		_w2533_
	);
	LUT2 #(
		.INIT('h1)
	) name1760 (
		_w2532_,
		_w2533_,
		_w2534_
	);
	LUT2 #(
		.INIT('h4)
	) name1761 (
		\g437_reg/NET0131 ,
		_w2534_,
		_w2535_
	);
	LUT2 #(
		.INIT('h2)
	) name1762 (
		\g392_reg/NET0131 ,
		\g401_reg/NET0131 ,
		_w2536_
	);
	LUT2 #(
		.INIT('h1)
	) name1763 (
		\g392_reg/NET0131 ,
		\g424_reg/NET0131 ,
		_w2537_
	);
	LUT2 #(
		.INIT('h1)
	) name1764 (
		_w2536_,
		_w2537_,
		_w2538_
	);
	LUT2 #(
		.INIT('h1)
	) name1765 (
		_w2534_,
		_w2538_,
		_w2539_
	);
	LUT2 #(
		.INIT('h1)
	) name1766 (
		_w2535_,
		_w2539_,
		_w2540_
	);
	LUT2 #(
		.INIT('h1)
	) name1767 (
		\g417_reg/NET0131 ,
		_w2540_,
		_w2541_
	);
	LUT2 #(
		.INIT('h8)
	) name1768 (
		\g417_reg/NET0131 ,
		_w2540_,
		_w2542_
	);
	LUT2 #(
		.INIT('h1)
	) name1769 (
		_w2531_,
		_w2541_,
		_w2543_
	);
	LUT2 #(
		.INIT('h4)
	) name1770 (
		_w2542_,
		_w2543_,
		_w2544_
	);
	LUT2 #(
		.INIT('h2)
	) name1771 (
		_w2519_,
		_w2544_,
		_w2545_
	);
	LUT2 #(
		.INIT('h4)
	) name1772 (
		\g703_reg/NET0131 ,
		_w2545_,
		_w2546_
	);
	LUT2 #(
		.INIT('h8)
	) name1773 (
		\g385_reg/NET0131 ,
		_w2517_,
		_w2547_
	);
	LUT2 #(
		.INIT('h1)
	) name1774 (
		_w2546_,
		_w2547_,
		_w2548_
	);
	LUT2 #(
		.INIT('h2)
	) name1775 (
		\g896_reg/NET0131 ,
		_w2548_,
		_w2549_
	);
	LUT2 #(
		.INIT('h8)
	) name1776 (
		\g35_pad ,
		\g862_reg/NET0131 ,
		_w2550_
	);
	LUT2 #(
		.INIT('h4)
	) name1777 (
		_w2549_,
		_w2550_,
		_w2551_
	);
	LUT2 #(
		.INIT('h4)
	) name1778 (
		\g35_pad ,
		\g446_reg/NET0131 ,
		_w2552_
	);
	LUT2 #(
		.INIT('h8)
	) name1779 (
		\g35_pad ,
		\g890_reg/NET0131 ,
		_w2553_
	);
	LUT2 #(
		.INIT('h8)
	) name1780 (
		\g896_reg/NET0131 ,
		_w2553_,
		_w2554_
	);
	LUT2 #(
		.INIT('h1)
	) name1781 (
		_w2552_,
		_w2554_,
		_w2555_
	);
	LUT2 #(
		.INIT('h4)
	) name1782 (
		_w2551_,
		_w2555_,
		_w2556_
	);
	LUT2 #(
		.INIT('h4)
	) name1783 (
		\g2153_reg/NET0131 ,
		\g2197_reg/NET0131 ,
		_w2557_
	);
	LUT2 #(
		.INIT('h4)
	) name1784 (
		\g2803_reg/NET0131 ,
		_w2504_,
		_w2558_
	);
	LUT2 #(
		.INIT('h2)
	) name1785 (
		_w2501_,
		_w2558_,
		_w2559_
	);
	LUT2 #(
		.INIT('h1)
	) name1786 (
		\g2715_reg/NET0131 ,
		\g2719_reg/NET0131 ,
		_w2560_
	);
	LUT2 #(
		.INIT('h4)
	) name1787 (
		_w2559_,
		_w2560_,
		_w2561_
	);
	LUT2 #(
		.INIT('h2)
	) name1788 (
		\g2208_reg/NET0131 ,
		\g2217_reg/NET0131 ,
		_w2562_
	);
	LUT2 #(
		.INIT('h8)
	) name1789 (
		\g35_pad ,
		_w2562_,
		_w2563_
	);
	LUT2 #(
		.INIT('h8)
	) name1790 (
		_w2561_,
		_w2563_,
		_w2564_
	);
	LUT2 #(
		.INIT('h4)
	) name1791 (
		_w2557_,
		_w2564_,
		_w2565_
	);
	LUT2 #(
		.INIT('h1)
	) name1792 (
		\g2173_reg/NET0131 ,
		\g35_pad ,
		_w2566_
	);
	LUT2 #(
		.INIT('h4)
	) name1793 (
		\g2193_reg/NET0131 ,
		\g35_pad ,
		_w2567_
	);
	LUT2 #(
		.INIT('h1)
	) name1794 (
		_w2566_,
		_w2567_,
		_w2568_
	);
	LUT2 #(
		.INIT('h4)
	) name1795 (
		_w2564_,
		_w2568_,
		_w2569_
	);
	LUT2 #(
		.INIT('h1)
	) name1796 (
		_w2565_,
		_w2569_,
		_w2570_
	);
	LUT2 #(
		.INIT('h4)
	) name1797 (
		\g2287_reg/NET0131 ,
		\g2331_reg/NET0131 ,
		_w2571_
	);
	LUT2 #(
		.INIT('h2)
	) name1798 (
		\g2715_reg/NET0131 ,
		\g2807_reg/NET0131 ,
		_w2572_
	);
	LUT2 #(
		.INIT('h4)
	) name1799 (
		\g2719_reg/NET0131 ,
		_w2504_,
		_w2573_
	);
	LUT2 #(
		.INIT('h8)
	) name1800 (
		_w2572_,
		_w2573_,
		_w2574_
	);
	LUT2 #(
		.INIT('h2)
	) name1801 (
		\g2715_reg/NET0131 ,
		\g2719_reg/NET0131 ,
		_w2575_
	);
	LUT2 #(
		.INIT('h4)
	) name1802 (
		_w2501_,
		_w2575_,
		_w2576_
	);
	LUT2 #(
		.INIT('h1)
	) name1803 (
		_w2574_,
		_w2576_,
		_w2577_
	);
	LUT2 #(
		.INIT('h2)
	) name1804 (
		\g2342_reg/NET0131 ,
		\g2351_reg/NET0131 ,
		_w2578_
	);
	LUT2 #(
		.INIT('h8)
	) name1805 (
		\g35_pad ,
		_w2578_,
		_w2579_
	);
	LUT2 #(
		.INIT('h4)
	) name1806 (
		_w2577_,
		_w2579_,
		_w2580_
	);
	LUT2 #(
		.INIT('h4)
	) name1807 (
		_w2571_,
		_w2580_,
		_w2581_
	);
	LUT2 #(
		.INIT('h1)
	) name1808 (
		\g2307_reg/NET0131 ,
		\g35_pad ,
		_w2582_
	);
	LUT2 #(
		.INIT('h4)
	) name1809 (
		\g2327_reg/NET0131 ,
		\g35_pad ,
		_w2583_
	);
	LUT2 #(
		.INIT('h1)
	) name1810 (
		_w2582_,
		_w2583_,
		_w2584_
	);
	LUT2 #(
		.INIT('h4)
	) name1811 (
		_w2580_,
		_w2584_,
		_w2585_
	);
	LUT2 #(
		.INIT('h1)
	) name1812 (
		_w2581_,
		_w2585_,
		_w2586_
	);
	LUT2 #(
		.INIT('h2)
	) name1813 (
		\g35_pad ,
		_w869_,
		_w2587_
	);
	LUT2 #(
		.INIT('h8)
	) name1814 (
		\g4704_reg/NET0131 ,
		_w2587_,
		_w2588_
	);
	LUT2 #(
		.INIT('h8)
	) name1815 (
		_w887_,
		_w2330_,
		_w2589_
	);
	LUT2 #(
		.INIT('h8)
	) name1816 (
		\g35_pad ,
		_w869_,
		_w2590_
	);
	LUT2 #(
		.INIT('h2)
	) name1817 (
		\g3343_reg/NET0131 ,
		\g5357_reg/NET0131 ,
		_w2591_
	);
	LUT2 #(
		.INIT('h8)
	) name1818 (
		\g3347_reg/NET0131 ,
		\g5357_reg/NET0131 ,
		_w2592_
	);
	LUT2 #(
		.INIT('h1)
	) name1819 (
		_w2591_,
		_w2592_,
		_w2593_
	);
	LUT2 #(
		.INIT('h4)
	) name1820 (
		\g5297_reg/NET0131 ,
		_w2593_,
		_w2594_
	);
	LUT2 #(
		.INIT('h2)
	) name1821 (
		\g5297_reg/NET0131 ,
		_w2593_,
		_w2595_
	);
	LUT2 #(
		.INIT('h1)
	) name1822 (
		\g4704_reg/NET0131 ,
		_w2594_,
		_w2596_
	);
	LUT2 #(
		.INIT('h4)
	) name1823 (
		_w2595_,
		_w2596_,
		_w2597_
	);
	LUT2 #(
		.INIT('h2)
	) name1824 (
		_w2589_,
		_w2597_,
		_w2598_
	);
	LUT2 #(
		.INIT('h8)
	) name1825 (
		_w2590_,
		_w2598_,
		_w2599_
	);
	LUT2 #(
		.INIT('h1)
	) name1826 (
		_w2588_,
		_w2599_,
		_w2600_
	);
	LUT2 #(
		.INIT('h4)
	) name1827 (
		\g2421_reg/NET0131 ,
		\g2465_reg/NET0131 ,
		_w2601_
	);
	LUT2 #(
		.INIT('h4)
	) name1828 (
		\g2815_reg/NET0131 ,
		_w2504_,
		_w2602_
	);
	LUT2 #(
		.INIT('h2)
	) name1829 (
		_w2501_,
		_w2602_,
		_w2603_
	);
	LUT2 #(
		.INIT('h2)
	) name1830 (
		_w2500_,
		_w2603_,
		_w2604_
	);
	LUT2 #(
		.INIT('h2)
	) name1831 (
		\g2476_reg/NET0131 ,
		\g2485_reg/NET0131 ,
		_w2605_
	);
	LUT2 #(
		.INIT('h8)
	) name1832 (
		\g35_pad ,
		_w2605_,
		_w2606_
	);
	LUT2 #(
		.INIT('h8)
	) name1833 (
		_w2604_,
		_w2606_,
		_w2607_
	);
	LUT2 #(
		.INIT('h4)
	) name1834 (
		_w2601_,
		_w2607_,
		_w2608_
	);
	LUT2 #(
		.INIT('h1)
	) name1835 (
		\g2441_reg/NET0131 ,
		\g35_pad ,
		_w2609_
	);
	LUT2 #(
		.INIT('h4)
	) name1836 (
		\g2461_reg/NET0131 ,
		\g35_pad ,
		_w2610_
	);
	LUT2 #(
		.INIT('h1)
	) name1837 (
		_w2609_,
		_w2610_,
		_w2611_
	);
	LUT2 #(
		.INIT('h4)
	) name1838 (
		_w2607_,
		_w2611_,
		_w2612_
	);
	LUT2 #(
		.INIT('h1)
	) name1839 (
		_w2608_,
		_w2612_,
		_w2613_
	);
	LUT2 #(
		.INIT('h4)
	) name1840 (
		\g2771_reg/NET0131 ,
		_w2504_,
		_w2614_
	);
	LUT2 #(
		.INIT('h2)
	) name1841 (
		_w2501_,
		_w2614_,
		_w2615_
	);
	LUT2 #(
		.INIT('h2)
	) name1842 (
		_w2560_,
		_w2615_,
		_w2616_
	);
	LUT2 #(
		.INIT('h8)
	) name1843 (
		_w829_,
		_w2616_,
		_w2617_
	);
	LUT2 #(
		.INIT('h4)
	) name1844 (
		\g1592_reg/NET0131 ,
		\g1636_reg/NET0131 ,
		_w2618_
	);
	LUT2 #(
		.INIT('h2)
	) name1845 (
		_w2617_,
		_w2618_,
		_w2619_
	);
	LUT2 #(
		.INIT('h2)
	) name1846 (
		\g1632_reg/NET0131 ,
		_w2617_,
		_w2620_
	);
	LUT2 #(
		.INIT('h1)
	) name1847 (
		_w2619_,
		_w2620_,
		_w2621_
	);
	LUT2 #(
		.INIT('h2)
	) name1848 (
		\g35_pad ,
		_w2621_,
		_w2622_
	);
	LUT2 #(
		.INIT('h2)
	) name1849 (
		\g1612_reg/NET0131 ,
		\g35_pad ,
		_w2623_
	);
	LUT2 #(
		.INIT('h1)
	) name1850 (
		_w2622_,
		_w2623_,
		_w2624_
	);
	LUT2 #(
		.INIT('h2)
	) name1851 (
		\g146_reg/NET0131 ,
		\g35_pad ,
		_w2625_
	);
	LUT2 #(
		.INIT('h1)
	) name1852 (
		\g164_reg/NET0131 ,
		_w2011_,
		_w2626_
	);
	LUT2 #(
		.INIT('h1)
	) name1853 (
		_w2012_,
		_w2626_,
		_w2627_
	);
	LUT2 #(
		.INIT('h8)
	) name1854 (
		_w2024_,
		_w2627_,
		_w2628_
	);
	LUT2 #(
		.INIT('h1)
	) name1855 (
		_w2625_,
		_w2628_,
		_w2629_
	);
	LUT2 #(
		.INIT('h4)
	) name1856 (
		\g758_reg/NET0131 ,
		_w2358_,
		_w2630_
	);
	LUT2 #(
		.INIT('h2)
	) name1857 (
		\g35_pad ,
		_w2630_,
		_w2631_
	);
	LUT2 #(
		.INIT('h2)
	) name1858 (
		\g749_reg/NET0131 ,
		_w2631_,
		_w2632_
	);
	LUT2 #(
		.INIT('h8)
	) name1859 (
		\g749_reg/NET0131 ,
		_w2358_,
		_w2633_
	);
	LUT2 #(
		.INIT('h8)
	) name1860 (
		\g758_reg/NET0131 ,
		_w967_,
		_w2634_
	);
	LUT2 #(
		.INIT('h4)
	) name1861 (
		_w2633_,
		_w2634_,
		_w2635_
	);
	LUT2 #(
		.INIT('h1)
	) name1862 (
		_w2632_,
		_w2635_,
		_w2636_
	);
	LUT2 #(
		.INIT('h4)
	) name1863 (
		\g35_pad ,
		\g832_reg/NET0131 ,
		_w2637_
	);
	LUT2 #(
		.INIT('h1)
	) name1864 (
		\g822_reg/NET0131 ,
		_w2208_,
		_w2638_
	);
	LUT2 #(
		.INIT('h4)
	) name1865 (
		_w2209_,
		_w2213_,
		_w2639_
	);
	LUT2 #(
		.INIT('h4)
	) name1866 (
		_w2638_,
		_w2639_,
		_w2640_
	);
	LUT2 #(
		.INIT('h1)
	) name1867 (
		_w2637_,
		_w2640_,
		_w2641_
	);
	LUT2 #(
		.INIT('h8)
	) name1868 (
		_w1299_,
		_w2136_,
		_w2642_
	);
	LUT2 #(
		.INIT('h8)
	) name1869 (
		\g4430_reg/NET0131 ,
		_w2642_,
		_w2643_
	);
	LUT2 #(
		.INIT('h1)
	) name1870 (
		\g4452_reg/NET0131 ,
		_w2643_,
		_w2644_
	);
	LUT2 #(
		.INIT('h4)
	) name1871 (
		\g2819_reg/NET0131 ,
		_w2504_,
		_w2645_
	);
	LUT2 #(
		.INIT('h2)
	) name1872 (
		_w2501_,
		_w2645_,
		_w2646_
	);
	LUT2 #(
		.INIT('h8)
	) name1873 (
		\g2715_reg/NET0131 ,
		\g2719_reg/NET0131 ,
		_w2647_
	);
	LUT2 #(
		.INIT('h4)
	) name1874 (
		_w2646_,
		_w2647_,
		_w2648_
	);
	LUT2 #(
		.INIT('h4)
	) name1875 (
		\g2587_reg/NET0131 ,
		\g2610_reg/NET0131 ,
		_w2649_
	);
	LUT2 #(
		.INIT('h8)
	) name1876 (
		_w2648_,
		_w2649_,
		_w2650_
	);
	LUT2 #(
		.INIT('h2)
	) name1877 (
		\g2648_reg/NET0131 ,
		\g2652_reg/NET0131 ,
		_w2651_
	);
	LUT2 #(
		.INIT('h4)
	) name1878 (
		\g2648_reg/NET0131 ,
		\g2652_reg/NET0131 ,
		_w2652_
	);
	LUT2 #(
		.INIT('h1)
	) name1879 (
		_w2651_,
		_w2652_,
		_w2653_
	);
	LUT2 #(
		.INIT('h2)
	) name1880 (
		_w2650_,
		_w2653_,
		_w2654_
	);
	LUT2 #(
		.INIT('h2)
	) name1881 (
		\g2657_reg/NET0131 ,
		_w2650_,
		_w2655_
	);
	LUT2 #(
		.INIT('h1)
	) name1882 (
		_w2654_,
		_w2655_,
		_w2656_
	);
	LUT2 #(
		.INIT('h2)
	) name1883 (
		\g35_pad ,
		_w2656_,
		_w2657_
	);
	LUT2 #(
		.INIT('h2)
	) name1884 (
		\g2652_reg/NET0131 ,
		\g35_pad ,
		_w2658_
	);
	LUT2 #(
		.INIT('h1)
	) name1885 (
		_w2657_,
		_w2658_,
		_w2659_
	);
	LUT2 #(
		.INIT('h8)
	) name1886 (
		\g2619_reg/NET0131 ,
		_w2648_,
		_w2660_
	);
	LUT2 #(
		.INIT('h8)
	) name1887 (
		\g2587_reg/NET0131 ,
		_w2660_,
		_w2661_
	);
	LUT2 #(
		.INIT('h2)
	) name1888 (
		\g2661_reg/NET0131 ,
		_w2661_,
		_w2662_
	);
	LUT2 #(
		.INIT('h4)
	) name1889 (
		\g2661_reg/NET0131 ,
		_w2661_,
		_w2663_
	);
	LUT2 #(
		.INIT('h1)
	) name1890 (
		_w2662_,
		_w2663_,
		_w2664_
	);
	LUT2 #(
		.INIT('h2)
	) name1891 (
		\g35_pad ,
		_w2664_,
		_w2665_
	);
	LUT2 #(
		.INIT('h2)
	) name1892 (
		\g2657_reg/NET0131 ,
		\g35_pad ,
		_w2666_
	);
	LUT2 #(
		.INIT('h1)
	) name1893 (
		_w2665_,
		_w2666_,
		_w2667_
	);
	LUT2 #(
		.INIT('h4)
	) name1894 (
		\g1624_reg/NET0131 ,
		\g1648_reg/NET0131 ,
		_w2668_
	);
	LUT2 #(
		.INIT('h8)
	) name1895 (
		_w2616_,
		_w2668_,
		_w2669_
	);
	LUT2 #(
		.INIT('h2)
	) name1896 (
		\g1687_reg/NET0131 ,
		\g1691_reg/NET0131 ,
		_w2670_
	);
	LUT2 #(
		.INIT('h4)
	) name1897 (
		\g1687_reg/NET0131 ,
		\g1691_reg/NET0131 ,
		_w2671_
	);
	LUT2 #(
		.INIT('h1)
	) name1898 (
		_w2670_,
		_w2671_,
		_w2672_
	);
	LUT2 #(
		.INIT('h2)
	) name1899 (
		_w2669_,
		_w2672_,
		_w2673_
	);
	LUT2 #(
		.INIT('h2)
	) name1900 (
		\g1696_reg/NET0131 ,
		_w2669_,
		_w2674_
	);
	LUT2 #(
		.INIT('h1)
	) name1901 (
		_w2673_,
		_w2674_,
		_w2675_
	);
	LUT2 #(
		.INIT('h2)
	) name1902 (
		\g35_pad ,
		_w2675_,
		_w2676_
	);
	LUT2 #(
		.INIT('h2)
	) name1903 (
		\g1691_reg/NET0131 ,
		\g35_pad ,
		_w2677_
	);
	LUT2 #(
		.INIT('h1)
	) name1904 (
		_w2676_,
		_w2677_,
		_w2678_
	);
	LUT2 #(
		.INIT('h2)
	) name1905 (
		\g35_pad ,
		_w2661_,
		_w2679_
	);
	LUT2 #(
		.INIT('h8)
	) name1906 (
		\g2675_reg/NET0131 ,
		_w2661_,
		_w2680_
	);
	LUT2 #(
		.INIT('h2)
	) name1907 (
		\g35_pad ,
		_w2680_,
		_w2681_
	);
	LUT2 #(
		.INIT('h1)
	) name1908 (
		\g2681_reg/NET0131 ,
		_w2681_,
		_w2682_
	);
	LUT2 #(
		.INIT('h1)
	) name1909 (
		\g2685_reg/NET0131 ,
		_w2661_,
		_w2683_
	);
	LUT2 #(
		.INIT('h4)
	) name1910 (
		\g2675_reg/NET0131 ,
		\g2681_reg/NET0131 ,
		_w2684_
	);
	LUT2 #(
		.INIT('h8)
	) name1911 (
		_w2661_,
		_w2684_,
		_w2685_
	);
	LUT2 #(
		.INIT('h1)
	) name1912 (
		_w2683_,
		_w2685_,
		_w2686_
	);
	LUT2 #(
		.INIT('h2)
	) name1913 (
		\g35_pad ,
		_w2686_,
		_w2687_
	);
	LUT2 #(
		.INIT('h1)
	) name1914 (
		_w2682_,
		_w2687_,
		_w2688_
	);
	LUT2 #(
		.INIT('h8)
	) name1915 (
		\g1657_reg/NET0131 ,
		_w2616_,
		_w2689_
	);
	LUT2 #(
		.INIT('h8)
	) name1916 (
		\g1624_reg/NET0131 ,
		_w2689_,
		_w2690_
	);
	LUT2 #(
		.INIT('h2)
	) name1917 (
		\g1700_reg/NET0131 ,
		_w2690_,
		_w2691_
	);
	LUT2 #(
		.INIT('h4)
	) name1918 (
		\g1700_reg/NET0131 ,
		_w2690_,
		_w2692_
	);
	LUT2 #(
		.INIT('h1)
	) name1919 (
		_w2691_,
		_w2692_,
		_w2693_
	);
	LUT2 #(
		.INIT('h2)
	) name1920 (
		\g35_pad ,
		_w2693_,
		_w2694_
	);
	LUT2 #(
		.INIT('h2)
	) name1921 (
		\g1696_reg/NET0131 ,
		\g35_pad ,
		_w2695_
	);
	LUT2 #(
		.INIT('h1)
	) name1922 (
		_w2694_,
		_w2695_,
		_w2696_
	);
	LUT2 #(
		.INIT('h8)
	) name1923 (
		\g1714_reg/NET0131 ,
		_w2690_,
		_w2697_
	);
	LUT2 #(
		.INIT('h2)
	) name1924 (
		\g35_pad ,
		_w2697_,
		_w2698_
	);
	LUT2 #(
		.INIT('h1)
	) name1925 (
		\g1720_reg/NET0131 ,
		_w2698_,
		_w2699_
	);
	LUT2 #(
		.INIT('h1)
	) name1926 (
		\g1724_reg/NET0131 ,
		_w2690_,
		_w2700_
	);
	LUT2 #(
		.INIT('h4)
	) name1927 (
		\g1714_reg/NET0131 ,
		\g1720_reg/NET0131 ,
		_w2701_
	);
	LUT2 #(
		.INIT('h8)
	) name1928 (
		_w2690_,
		_w2701_,
		_w2702_
	);
	LUT2 #(
		.INIT('h1)
	) name1929 (
		_w2700_,
		_w2702_,
		_w2703_
	);
	LUT2 #(
		.INIT('h2)
	) name1930 (
		\g35_pad ,
		_w2703_,
		_w2704_
	);
	LUT2 #(
		.INIT('h1)
	) name1931 (
		_w2699_,
		_w2704_,
		_w2705_
	);
	LUT2 #(
		.INIT('h2)
	) name1932 (
		\g35_pad ,
		_w2690_,
		_w2706_
	);
	LUT2 #(
		.INIT('h2)
	) name1933 (
		\g2715_reg/NET0131 ,
		\g2775_reg/NET0131 ,
		_w2707_
	);
	LUT2 #(
		.INIT('h8)
	) name1934 (
		_w2573_,
		_w2707_,
		_w2708_
	);
	LUT2 #(
		.INIT('h1)
	) name1935 (
		_w2576_,
		_w2708_,
		_w2709_
	);
	LUT2 #(
		.INIT('h2)
	) name1936 (
		\g1792_reg/NET0131 ,
		_w2709_,
		_w2710_
	);
	LUT2 #(
		.INIT('h1)
	) name1937 (
		\g1783_reg/NET0131 ,
		_w2709_,
		_w2711_
	);
	LUT2 #(
		.INIT('h1)
	) name1938 (
		\g1760_reg/NET0131 ,
		_w2711_,
		_w2712_
	);
	LUT2 #(
		.INIT('h1)
	) name1939 (
		_w2710_,
		_w2712_,
		_w2713_
	);
	LUT2 #(
		.INIT('h2)
	) name1940 (
		\g35_pad ,
		_w2713_,
		_w2714_
	);
	LUT2 #(
		.INIT('h1)
	) name1941 (
		\g1768_reg/NET0131 ,
		\g35_pad ,
		_w2715_
	);
	LUT2 #(
		.INIT('h1)
	) name1942 (
		_w2714_,
		_w2715_,
		_w2716_
	);
	LUT2 #(
		.INIT('h2)
	) name1943 (
		\g1783_reg/NET0131 ,
		_w2709_,
		_w2717_
	);
	LUT2 #(
		.INIT('h4)
	) name1944 (
		\g1760_reg/NET0131 ,
		_w2717_,
		_w2718_
	);
	LUT2 #(
		.INIT('h2)
	) name1945 (
		\g1821_reg/NET0131 ,
		\g1825_reg/NET0131 ,
		_w2719_
	);
	LUT2 #(
		.INIT('h4)
	) name1946 (
		\g1821_reg/NET0131 ,
		\g1825_reg/NET0131 ,
		_w2720_
	);
	LUT2 #(
		.INIT('h1)
	) name1947 (
		_w2719_,
		_w2720_,
		_w2721_
	);
	LUT2 #(
		.INIT('h2)
	) name1948 (
		_w2718_,
		_w2721_,
		_w2722_
	);
	LUT2 #(
		.INIT('h2)
	) name1949 (
		\g1830_reg/NET0131 ,
		_w2718_,
		_w2723_
	);
	LUT2 #(
		.INIT('h1)
	) name1950 (
		_w2722_,
		_w2723_,
		_w2724_
	);
	LUT2 #(
		.INIT('h2)
	) name1951 (
		\g35_pad ,
		_w2724_,
		_w2725_
	);
	LUT2 #(
		.INIT('h2)
	) name1952 (
		\g1825_reg/NET0131 ,
		\g35_pad ,
		_w2726_
	);
	LUT2 #(
		.INIT('h1)
	) name1953 (
		_w2725_,
		_w2726_,
		_w2727_
	);
	LUT2 #(
		.INIT('h8)
	) name1954 (
		\g1760_reg/NET0131 ,
		_w2710_,
		_w2728_
	);
	LUT2 #(
		.INIT('h2)
	) name1955 (
		\g1834_reg/NET0131 ,
		_w2728_,
		_w2729_
	);
	LUT2 #(
		.INIT('h4)
	) name1956 (
		\g1834_reg/NET0131 ,
		_w2728_,
		_w2730_
	);
	LUT2 #(
		.INIT('h1)
	) name1957 (
		_w2729_,
		_w2730_,
		_w2731_
	);
	LUT2 #(
		.INIT('h2)
	) name1958 (
		\g35_pad ,
		_w2731_,
		_w2732_
	);
	LUT2 #(
		.INIT('h2)
	) name1959 (
		\g1830_reg/NET0131 ,
		\g35_pad ,
		_w2733_
	);
	LUT2 #(
		.INIT('h1)
	) name1960 (
		_w2732_,
		_w2733_,
		_w2734_
	);
	LUT2 #(
		.INIT('h8)
	) name1961 (
		\g1848_reg/NET0131 ,
		_w2728_,
		_w2735_
	);
	LUT2 #(
		.INIT('h2)
	) name1962 (
		\g35_pad ,
		_w2735_,
		_w2736_
	);
	LUT2 #(
		.INIT('h1)
	) name1963 (
		\g1854_reg/NET0131 ,
		_w2736_,
		_w2737_
	);
	LUT2 #(
		.INIT('h1)
	) name1964 (
		\g1858_reg/NET0131 ,
		_w2728_,
		_w2738_
	);
	LUT2 #(
		.INIT('h4)
	) name1965 (
		\g1848_reg/NET0131 ,
		\g1854_reg/NET0131 ,
		_w2739_
	);
	LUT2 #(
		.INIT('h8)
	) name1966 (
		_w2728_,
		_w2739_,
		_w2740_
	);
	LUT2 #(
		.INIT('h1)
	) name1967 (
		_w2738_,
		_w2740_,
		_w2741_
	);
	LUT2 #(
		.INIT('h2)
	) name1968 (
		\g35_pad ,
		_w2741_,
		_w2742_
	);
	LUT2 #(
		.INIT('h1)
	) name1969 (
		_w2737_,
		_w2742_,
		_w2743_
	);
	LUT2 #(
		.INIT('h2)
	) name1970 (
		\g35_pad ,
		_w2728_,
		_w2744_
	);
	LUT2 #(
		.INIT('h8)
	) name1971 (
		\g1926_reg/NET0131 ,
		_w2507_,
		_w2745_
	);
	LUT2 #(
		.INIT('h4)
	) name1972 (
		\g1917_reg/NET0131 ,
		_w2507_,
		_w2746_
	);
	LUT2 #(
		.INIT('h1)
	) name1973 (
		\g1894_reg/NET0131 ,
		_w2746_,
		_w2747_
	);
	LUT2 #(
		.INIT('h1)
	) name1974 (
		_w2745_,
		_w2747_,
		_w2748_
	);
	LUT2 #(
		.INIT('h2)
	) name1975 (
		\g35_pad ,
		_w2748_,
		_w2749_
	);
	LUT2 #(
		.INIT('h1)
	) name1976 (
		\g1902_reg/NET0131 ,
		\g35_pad ,
		_w2750_
	);
	LUT2 #(
		.INIT('h1)
	) name1977 (
		_w2749_,
		_w2750_,
		_w2751_
	);
	LUT2 #(
		.INIT('h4)
	) name1978 (
		\g1894_reg/NET0131 ,
		\g1917_reg/NET0131 ,
		_w2752_
	);
	LUT2 #(
		.INIT('h8)
	) name1979 (
		_w2507_,
		_w2752_,
		_w2753_
	);
	LUT2 #(
		.INIT('h2)
	) name1980 (
		\g1955_reg/NET0131 ,
		\g1959_reg/NET0131 ,
		_w2754_
	);
	LUT2 #(
		.INIT('h4)
	) name1981 (
		\g1955_reg/NET0131 ,
		\g1959_reg/NET0131 ,
		_w2755_
	);
	LUT2 #(
		.INIT('h1)
	) name1982 (
		_w2754_,
		_w2755_,
		_w2756_
	);
	LUT2 #(
		.INIT('h2)
	) name1983 (
		_w2753_,
		_w2756_,
		_w2757_
	);
	LUT2 #(
		.INIT('h2)
	) name1984 (
		\g1964_reg/NET0131 ,
		_w2753_,
		_w2758_
	);
	LUT2 #(
		.INIT('h1)
	) name1985 (
		_w2757_,
		_w2758_,
		_w2759_
	);
	LUT2 #(
		.INIT('h2)
	) name1986 (
		\g35_pad ,
		_w2759_,
		_w2760_
	);
	LUT2 #(
		.INIT('h2)
	) name1987 (
		\g1959_reg/NET0131 ,
		\g35_pad ,
		_w2761_
	);
	LUT2 #(
		.INIT('h1)
	) name1988 (
		_w2760_,
		_w2761_,
		_w2762_
	);
	LUT2 #(
		.INIT('h8)
	) name1989 (
		\g1894_reg/NET0131 ,
		_w2745_,
		_w2763_
	);
	LUT2 #(
		.INIT('h2)
	) name1990 (
		\g1968_reg/NET0131 ,
		_w2763_,
		_w2764_
	);
	LUT2 #(
		.INIT('h4)
	) name1991 (
		\g1968_reg/NET0131 ,
		_w2763_,
		_w2765_
	);
	LUT2 #(
		.INIT('h1)
	) name1992 (
		_w2764_,
		_w2765_,
		_w2766_
	);
	LUT2 #(
		.INIT('h2)
	) name1993 (
		\g35_pad ,
		_w2766_,
		_w2767_
	);
	LUT2 #(
		.INIT('h2)
	) name1994 (
		\g1964_reg/NET0131 ,
		\g35_pad ,
		_w2768_
	);
	LUT2 #(
		.INIT('h1)
	) name1995 (
		_w2767_,
		_w2768_,
		_w2769_
	);
	LUT2 #(
		.INIT('h2)
	) name1996 (
		\g35_pad ,
		_w2763_,
		_w2770_
	);
	LUT2 #(
		.INIT('h8)
	) name1997 (
		\g1982_reg/NET0131 ,
		_w2763_,
		_w2771_
	);
	LUT2 #(
		.INIT('h2)
	) name1998 (
		\g35_pad ,
		_w2771_,
		_w2772_
	);
	LUT2 #(
		.INIT('h1)
	) name1999 (
		\g1988_reg/NET0131 ,
		_w2772_,
		_w2773_
	);
	LUT2 #(
		.INIT('h1)
	) name2000 (
		\g1992_reg/NET0131 ,
		_w2763_,
		_w2774_
	);
	LUT2 #(
		.INIT('h4)
	) name2001 (
		\g1982_reg/NET0131 ,
		\g1988_reg/NET0131 ,
		_w2775_
	);
	LUT2 #(
		.INIT('h8)
	) name2002 (
		_w2763_,
		_w2775_,
		_w2776_
	);
	LUT2 #(
		.INIT('h1)
	) name2003 (
		_w2774_,
		_w2776_,
		_w2777_
	);
	LUT2 #(
		.INIT('h2)
	) name2004 (
		\g35_pad ,
		_w2777_,
		_w2778_
	);
	LUT2 #(
		.INIT('h1)
	) name2005 (
		_w2773_,
		_w2778_,
		_w2779_
	);
	LUT2 #(
		.INIT('h4)
	) name2006 (
		\g2787_reg/NET0131 ,
		_w2504_,
		_w2780_
	);
	LUT2 #(
		.INIT('h2)
	) name2007 (
		_w2501_,
		_w2780_,
		_w2781_
	);
	LUT2 #(
		.INIT('h2)
	) name2008 (
		_w2647_,
		_w2781_,
		_w2782_
	);
	LUT2 #(
		.INIT('h4)
	) name2009 (
		\g2028_reg/NET0131 ,
		\g2051_reg/NET0131 ,
		_w2783_
	);
	LUT2 #(
		.INIT('h8)
	) name2010 (
		_w2782_,
		_w2783_,
		_w2784_
	);
	LUT2 #(
		.INIT('h2)
	) name2011 (
		\g2089_reg/NET0131 ,
		\g2093_reg/NET0131 ,
		_w2785_
	);
	LUT2 #(
		.INIT('h4)
	) name2012 (
		\g2089_reg/NET0131 ,
		\g2093_reg/NET0131 ,
		_w2786_
	);
	LUT2 #(
		.INIT('h1)
	) name2013 (
		_w2785_,
		_w2786_,
		_w2787_
	);
	LUT2 #(
		.INIT('h2)
	) name2014 (
		_w2784_,
		_w2787_,
		_w2788_
	);
	LUT2 #(
		.INIT('h2)
	) name2015 (
		\g2098_reg/NET0131 ,
		_w2784_,
		_w2789_
	);
	LUT2 #(
		.INIT('h1)
	) name2016 (
		_w2788_,
		_w2789_,
		_w2790_
	);
	LUT2 #(
		.INIT('h2)
	) name2017 (
		\g35_pad ,
		_w2790_,
		_w2791_
	);
	LUT2 #(
		.INIT('h2)
	) name2018 (
		\g2093_reg/NET0131 ,
		\g35_pad ,
		_w2792_
	);
	LUT2 #(
		.INIT('h1)
	) name2019 (
		_w2791_,
		_w2792_,
		_w2793_
	);
	LUT2 #(
		.INIT('h8)
	) name2020 (
		\g2060_reg/NET0131 ,
		_w2782_,
		_w2794_
	);
	LUT2 #(
		.INIT('h8)
	) name2021 (
		\g2028_reg/NET0131 ,
		_w2794_,
		_w2795_
	);
	LUT2 #(
		.INIT('h2)
	) name2022 (
		\g2102_reg/NET0131 ,
		_w2795_,
		_w2796_
	);
	LUT2 #(
		.INIT('h4)
	) name2023 (
		\g2102_reg/NET0131 ,
		_w2795_,
		_w2797_
	);
	LUT2 #(
		.INIT('h1)
	) name2024 (
		_w2796_,
		_w2797_,
		_w2798_
	);
	LUT2 #(
		.INIT('h2)
	) name2025 (
		\g35_pad ,
		_w2798_,
		_w2799_
	);
	LUT2 #(
		.INIT('h2)
	) name2026 (
		\g2098_reg/NET0131 ,
		\g35_pad ,
		_w2800_
	);
	LUT2 #(
		.INIT('h1)
	) name2027 (
		_w2799_,
		_w2800_,
		_w2801_
	);
	LUT2 #(
		.INIT('h2)
	) name2028 (
		\g35_pad ,
		_w2795_,
		_w2802_
	);
	LUT2 #(
		.INIT('h8)
	) name2029 (
		\g2116_reg/NET0131 ,
		_w2795_,
		_w2803_
	);
	LUT2 #(
		.INIT('h2)
	) name2030 (
		\g35_pad ,
		_w2803_,
		_w2804_
	);
	LUT2 #(
		.INIT('h1)
	) name2031 (
		\g2122_reg/NET0131 ,
		_w2804_,
		_w2805_
	);
	LUT2 #(
		.INIT('h1)
	) name2032 (
		\g2126_reg/NET0131 ,
		_w2795_,
		_w2806_
	);
	LUT2 #(
		.INIT('h4)
	) name2033 (
		\g2116_reg/NET0131 ,
		\g2122_reg/NET0131 ,
		_w2807_
	);
	LUT2 #(
		.INIT('h8)
	) name2034 (
		_w2795_,
		_w2807_,
		_w2808_
	);
	LUT2 #(
		.INIT('h1)
	) name2035 (
		_w2806_,
		_w2808_,
		_w2809_
	);
	LUT2 #(
		.INIT('h2)
	) name2036 (
		\g35_pad ,
		_w2809_,
		_w2810_
	);
	LUT2 #(
		.INIT('h1)
	) name2037 (
		_w2805_,
		_w2810_,
		_w2811_
	);
	LUT2 #(
		.INIT('h4)
	) name2038 (
		\g2185_reg/NET0131 ,
		\g2208_reg/NET0131 ,
		_w2812_
	);
	LUT2 #(
		.INIT('h8)
	) name2039 (
		_w2561_,
		_w2812_,
		_w2813_
	);
	LUT2 #(
		.INIT('h2)
	) name2040 (
		\g2246_reg/NET0131 ,
		\g2250_reg/NET0131 ,
		_w2814_
	);
	LUT2 #(
		.INIT('h4)
	) name2041 (
		\g2246_reg/NET0131 ,
		\g2250_reg/NET0131 ,
		_w2815_
	);
	LUT2 #(
		.INIT('h1)
	) name2042 (
		_w2814_,
		_w2815_,
		_w2816_
	);
	LUT2 #(
		.INIT('h2)
	) name2043 (
		_w2813_,
		_w2816_,
		_w2817_
	);
	LUT2 #(
		.INIT('h2)
	) name2044 (
		\g2255_reg/NET0131 ,
		_w2813_,
		_w2818_
	);
	LUT2 #(
		.INIT('h1)
	) name2045 (
		_w2817_,
		_w2818_,
		_w2819_
	);
	LUT2 #(
		.INIT('h2)
	) name2046 (
		\g35_pad ,
		_w2819_,
		_w2820_
	);
	LUT2 #(
		.INIT('h2)
	) name2047 (
		\g2250_reg/NET0131 ,
		\g35_pad ,
		_w2821_
	);
	LUT2 #(
		.INIT('h1)
	) name2048 (
		_w2820_,
		_w2821_,
		_w2822_
	);
	LUT2 #(
		.INIT('h8)
	) name2049 (
		\g2217_reg/NET0131 ,
		_w2561_,
		_w2823_
	);
	LUT2 #(
		.INIT('h8)
	) name2050 (
		\g2185_reg/NET0131 ,
		_w2823_,
		_w2824_
	);
	LUT2 #(
		.INIT('h2)
	) name2051 (
		\g2259_reg/NET0131 ,
		_w2824_,
		_w2825_
	);
	LUT2 #(
		.INIT('h4)
	) name2052 (
		\g2259_reg/NET0131 ,
		_w2824_,
		_w2826_
	);
	LUT2 #(
		.INIT('h1)
	) name2053 (
		_w2825_,
		_w2826_,
		_w2827_
	);
	LUT2 #(
		.INIT('h2)
	) name2054 (
		\g35_pad ,
		_w2827_,
		_w2828_
	);
	LUT2 #(
		.INIT('h2)
	) name2055 (
		\g2255_reg/NET0131 ,
		\g35_pad ,
		_w2829_
	);
	LUT2 #(
		.INIT('h1)
	) name2056 (
		_w2828_,
		_w2829_,
		_w2830_
	);
	LUT2 #(
		.INIT('h2)
	) name2057 (
		\g35_pad ,
		_w2824_,
		_w2831_
	);
	LUT2 #(
		.INIT('h8)
	) name2058 (
		\g2273_reg/NET0131 ,
		_w2824_,
		_w2832_
	);
	LUT2 #(
		.INIT('h2)
	) name2059 (
		\g35_pad ,
		_w2832_,
		_w2833_
	);
	LUT2 #(
		.INIT('h1)
	) name2060 (
		\g2279_reg/NET0131 ,
		_w2833_,
		_w2834_
	);
	LUT2 #(
		.INIT('h1)
	) name2061 (
		\g2283_reg/NET0131 ,
		_w2824_,
		_w2835_
	);
	LUT2 #(
		.INIT('h4)
	) name2062 (
		\g2273_reg/NET0131 ,
		\g2279_reg/NET0131 ,
		_w2836_
	);
	LUT2 #(
		.INIT('h8)
	) name2063 (
		_w2824_,
		_w2836_,
		_w2837_
	);
	LUT2 #(
		.INIT('h1)
	) name2064 (
		_w2835_,
		_w2837_,
		_w2838_
	);
	LUT2 #(
		.INIT('h2)
	) name2065 (
		\g35_pad ,
		_w2838_,
		_w2839_
	);
	LUT2 #(
		.INIT('h1)
	) name2066 (
		_w2834_,
		_w2839_,
		_w2840_
	);
	LUT2 #(
		.INIT('h2)
	) name2067 (
		\g2351_reg/NET0131 ,
		_w2577_,
		_w2841_
	);
	LUT2 #(
		.INIT('h1)
	) name2068 (
		\g2342_reg/NET0131 ,
		_w2577_,
		_w2842_
	);
	LUT2 #(
		.INIT('h1)
	) name2069 (
		\g2319_reg/NET0131 ,
		_w2842_,
		_w2843_
	);
	LUT2 #(
		.INIT('h1)
	) name2070 (
		_w2841_,
		_w2843_,
		_w2844_
	);
	LUT2 #(
		.INIT('h2)
	) name2071 (
		\g35_pad ,
		_w2844_,
		_w2845_
	);
	LUT2 #(
		.INIT('h1)
	) name2072 (
		\g2327_reg/NET0131 ,
		\g35_pad ,
		_w2846_
	);
	LUT2 #(
		.INIT('h1)
	) name2073 (
		_w2845_,
		_w2846_,
		_w2847_
	);
	LUT2 #(
		.INIT('h4)
	) name2074 (
		\g2319_reg/NET0131 ,
		\g2342_reg/NET0131 ,
		_w2848_
	);
	LUT2 #(
		.INIT('h4)
	) name2075 (
		_w2577_,
		_w2848_,
		_w2849_
	);
	LUT2 #(
		.INIT('h2)
	) name2076 (
		\g2380_reg/NET0131 ,
		\g2384_reg/NET0131 ,
		_w2850_
	);
	LUT2 #(
		.INIT('h4)
	) name2077 (
		\g2380_reg/NET0131 ,
		\g2384_reg/NET0131 ,
		_w2851_
	);
	LUT2 #(
		.INIT('h1)
	) name2078 (
		_w2850_,
		_w2851_,
		_w2852_
	);
	LUT2 #(
		.INIT('h2)
	) name2079 (
		_w2849_,
		_w2852_,
		_w2853_
	);
	LUT2 #(
		.INIT('h2)
	) name2080 (
		\g2389_reg/NET0131 ,
		_w2849_,
		_w2854_
	);
	LUT2 #(
		.INIT('h1)
	) name2081 (
		_w2853_,
		_w2854_,
		_w2855_
	);
	LUT2 #(
		.INIT('h2)
	) name2082 (
		\g35_pad ,
		_w2855_,
		_w2856_
	);
	LUT2 #(
		.INIT('h2)
	) name2083 (
		\g2384_reg/NET0131 ,
		\g35_pad ,
		_w2857_
	);
	LUT2 #(
		.INIT('h1)
	) name2084 (
		_w2856_,
		_w2857_,
		_w2858_
	);
	LUT2 #(
		.INIT('h8)
	) name2085 (
		\g2319_reg/NET0131 ,
		_w2841_,
		_w2859_
	);
	LUT2 #(
		.INIT('h2)
	) name2086 (
		\g2393_reg/NET0131 ,
		_w2859_,
		_w2860_
	);
	LUT2 #(
		.INIT('h4)
	) name2087 (
		\g2393_reg/NET0131 ,
		_w2859_,
		_w2861_
	);
	LUT2 #(
		.INIT('h1)
	) name2088 (
		_w2860_,
		_w2861_,
		_w2862_
	);
	LUT2 #(
		.INIT('h2)
	) name2089 (
		\g35_pad ,
		_w2862_,
		_w2863_
	);
	LUT2 #(
		.INIT('h2)
	) name2090 (
		\g2389_reg/NET0131 ,
		\g35_pad ,
		_w2864_
	);
	LUT2 #(
		.INIT('h1)
	) name2091 (
		_w2863_,
		_w2864_,
		_w2865_
	);
	LUT2 #(
		.INIT('h2)
	) name2092 (
		\g35_pad ,
		_w2859_,
		_w2866_
	);
	LUT2 #(
		.INIT('h8)
	) name2093 (
		\g2407_reg/NET0131 ,
		_w2859_,
		_w2867_
	);
	LUT2 #(
		.INIT('h2)
	) name2094 (
		\g35_pad ,
		_w2867_,
		_w2868_
	);
	LUT2 #(
		.INIT('h1)
	) name2095 (
		\g2413_reg/NET0131 ,
		_w2868_,
		_w2869_
	);
	LUT2 #(
		.INIT('h1)
	) name2096 (
		\g2417_reg/NET0131 ,
		_w2859_,
		_w2870_
	);
	LUT2 #(
		.INIT('h4)
	) name2097 (
		\g2407_reg/NET0131 ,
		\g2413_reg/NET0131 ,
		_w2871_
	);
	LUT2 #(
		.INIT('h8)
	) name2098 (
		_w2859_,
		_w2871_,
		_w2872_
	);
	LUT2 #(
		.INIT('h1)
	) name2099 (
		_w2870_,
		_w2872_,
		_w2873_
	);
	LUT2 #(
		.INIT('h2)
	) name2100 (
		\g35_pad ,
		_w2873_,
		_w2874_
	);
	LUT2 #(
		.INIT('h1)
	) name2101 (
		_w2869_,
		_w2874_,
		_w2875_
	);
	LUT2 #(
		.INIT('h8)
	) name2102 (
		\g2485_reg/NET0131 ,
		_w2604_,
		_w2876_
	);
	LUT2 #(
		.INIT('h4)
	) name2103 (
		\g2476_reg/NET0131 ,
		_w2604_,
		_w2877_
	);
	LUT2 #(
		.INIT('h1)
	) name2104 (
		\g2453_reg/NET0131 ,
		_w2877_,
		_w2878_
	);
	LUT2 #(
		.INIT('h1)
	) name2105 (
		_w2876_,
		_w2878_,
		_w2879_
	);
	LUT2 #(
		.INIT('h2)
	) name2106 (
		\g35_pad ,
		_w2879_,
		_w2880_
	);
	LUT2 #(
		.INIT('h1)
	) name2107 (
		\g2461_reg/NET0131 ,
		\g35_pad ,
		_w2881_
	);
	LUT2 #(
		.INIT('h1)
	) name2108 (
		_w2880_,
		_w2881_,
		_w2882_
	);
	LUT2 #(
		.INIT('h4)
	) name2109 (
		\g2453_reg/NET0131 ,
		\g2476_reg/NET0131 ,
		_w2883_
	);
	LUT2 #(
		.INIT('h8)
	) name2110 (
		_w2604_,
		_w2883_,
		_w2884_
	);
	LUT2 #(
		.INIT('h2)
	) name2111 (
		\g2514_reg/NET0131 ,
		\g2518_reg/NET0131 ,
		_w2885_
	);
	LUT2 #(
		.INIT('h4)
	) name2112 (
		\g2514_reg/NET0131 ,
		\g2518_reg/NET0131 ,
		_w2886_
	);
	LUT2 #(
		.INIT('h1)
	) name2113 (
		_w2885_,
		_w2886_,
		_w2887_
	);
	LUT2 #(
		.INIT('h2)
	) name2114 (
		_w2884_,
		_w2887_,
		_w2888_
	);
	LUT2 #(
		.INIT('h2)
	) name2115 (
		\g2523_reg/NET0131 ,
		_w2884_,
		_w2889_
	);
	LUT2 #(
		.INIT('h1)
	) name2116 (
		_w2888_,
		_w2889_,
		_w2890_
	);
	LUT2 #(
		.INIT('h2)
	) name2117 (
		\g35_pad ,
		_w2890_,
		_w2891_
	);
	LUT2 #(
		.INIT('h2)
	) name2118 (
		\g2518_reg/NET0131 ,
		\g35_pad ,
		_w2892_
	);
	LUT2 #(
		.INIT('h1)
	) name2119 (
		_w2891_,
		_w2892_,
		_w2893_
	);
	LUT2 #(
		.INIT('h8)
	) name2120 (
		\g2453_reg/NET0131 ,
		_w2876_,
		_w2894_
	);
	LUT2 #(
		.INIT('h2)
	) name2121 (
		\g2527_reg/NET0131 ,
		_w2894_,
		_w2895_
	);
	LUT2 #(
		.INIT('h4)
	) name2122 (
		\g2527_reg/NET0131 ,
		_w2894_,
		_w2896_
	);
	LUT2 #(
		.INIT('h1)
	) name2123 (
		_w2895_,
		_w2896_,
		_w2897_
	);
	LUT2 #(
		.INIT('h2)
	) name2124 (
		\g35_pad ,
		_w2897_,
		_w2898_
	);
	LUT2 #(
		.INIT('h2)
	) name2125 (
		\g2523_reg/NET0131 ,
		\g35_pad ,
		_w2899_
	);
	LUT2 #(
		.INIT('h1)
	) name2126 (
		_w2898_,
		_w2899_,
		_w2900_
	);
	LUT2 #(
		.INIT('h2)
	) name2127 (
		\g35_pad ,
		_w2894_,
		_w2901_
	);
	LUT2 #(
		.INIT('h8)
	) name2128 (
		\g2541_reg/NET0131 ,
		_w2894_,
		_w2902_
	);
	LUT2 #(
		.INIT('h2)
	) name2129 (
		\g35_pad ,
		_w2902_,
		_w2903_
	);
	LUT2 #(
		.INIT('h1)
	) name2130 (
		\g2547_reg/NET0131 ,
		_w2903_,
		_w2904_
	);
	LUT2 #(
		.INIT('h1)
	) name2131 (
		\g2551_reg/NET0131 ,
		_w2894_,
		_w2905_
	);
	LUT2 #(
		.INIT('h4)
	) name2132 (
		\g2541_reg/NET0131 ,
		\g2547_reg/NET0131 ,
		_w2906_
	);
	LUT2 #(
		.INIT('h8)
	) name2133 (
		_w2894_,
		_w2906_,
		_w2907_
	);
	LUT2 #(
		.INIT('h1)
	) name2134 (
		_w2905_,
		_w2907_,
		_w2908_
	);
	LUT2 #(
		.INIT('h2)
	) name2135 (
		\g35_pad ,
		_w2908_,
		_w2909_
	);
	LUT2 #(
		.INIT('h1)
	) name2136 (
		_w2904_,
		_w2909_,
		_w2910_
	);
	LUT2 #(
		.INIT('h4)
	) name2137 (
		\g2051_reg/NET0131 ,
		_w2782_,
		_w2911_
	);
	LUT2 #(
		.INIT('h1)
	) name2138 (
		\g2028_reg/NET0131 ,
		_w2911_,
		_w2912_
	);
	LUT2 #(
		.INIT('h1)
	) name2139 (
		_w2794_,
		_w2912_,
		_w2913_
	);
	LUT2 #(
		.INIT('h2)
	) name2140 (
		\g35_pad ,
		_w2913_,
		_w2914_
	);
	LUT2 #(
		.INIT('h1)
	) name2141 (
		\g2036_reg/NET0131 ,
		\g35_pad ,
		_w2915_
	);
	LUT2 #(
		.INIT('h1)
	) name2142 (
		_w2914_,
		_w2915_,
		_w2916_
	);
	LUT2 #(
		.INIT('h4)
	) name2143 (
		\g2208_reg/NET0131 ,
		_w2561_,
		_w2917_
	);
	LUT2 #(
		.INIT('h1)
	) name2144 (
		\g2185_reg/NET0131 ,
		_w2917_,
		_w2918_
	);
	LUT2 #(
		.INIT('h1)
	) name2145 (
		_w2823_,
		_w2918_,
		_w2919_
	);
	LUT2 #(
		.INIT('h2)
	) name2146 (
		\g35_pad ,
		_w2919_,
		_w2920_
	);
	LUT2 #(
		.INIT('h1)
	) name2147 (
		\g2193_reg/NET0131 ,
		\g35_pad ,
		_w2921_
	);
	LUT2 #(
		.INIT('h1)
	) name2148 (
		_w2920_,
		_w2921_,
		_w2922_
	);
	LUT2 #(
		.INIT('h4)
	) name2149 (
		\g1648_reg/NET0131 ,
		_w2616_,
		_w2923_
	);
	LUT2 #(
		.INIT('h1)
	) name2150 (
		\g1624_reg/NET0131 ,
		_w2923_,
		_w2924_
	);
	LUT2 #(
		.INIT('h1)
	) name2151 (
		_w2689_,
		_w2924_,
		_w2925_
	);
	LUT2 #(
		.INIT('h2)
	) name2152 (
		\g35_pad ,
		_w2925_,
		_w2926_
	);
	LUT2 #(
		.INIT('h1)
	) name2153 (
		\g1632_reg/NET0131 ,
		\g35_pad ,
		_w2927_
	);
	LUT2 #(
		.INIT('h1)
	) name2154 (
		_w2926_,
		_w2927_,
		_w2928_
	);
	LUT2 #(
		.INIT('h4)
	) name2155 (
		\g2610_reg/NET0131 ,
		_w2648_,
		_w2929_
	);
	LUT2 #(
		.INIT('h1)
	) name2156 (
		\g2587_reg/NET0131 ,
		_w2929_,
		_w2930_
	);
	LUT2 #(
		.INIT('h1)
	) name2157 (
		_w2660_,
		_w2930_,
		_w2931_
	);
	LUT2 #(
		.INIT('h2)
	) name2158 (
		\g35_pad ,
		_w2931_,
		_w2932_
	);
	LUT2 #(
		.INIT('h1)
	) name2159 (
		\g2595_reg/NET0131 ,
		\g35_pad ,
		_w2933_
	);
	LUT2 #(
		.INIT('h1)
	) name2160 (
		_w2932_,
		_w2933_,
		_w2934_
	);
	LUT2 #(
		.INIT('h2)
	) name2161 (
		\g4438_reg/NET0131 ,
		_w1363_,
		_w2935_
	);
	LUT2 #(
		.INIT('h8)
	) name2162 (
		_w1365_,
		_w2136_,
		_w2936_
	);
	LUT2 #(
		.INIT('h1)
	) name2163 (
		_w2935_,
		_w2936_,
		_w2937_
	);
	LUT2 #(
		.INIT('h2)
	) name2164 (
		\g35_pad ,
		\g5084_reg/NET0131 ,
		_w2938_
	);
	LUT2 #(
		.INIT('h2)
	) name2165 (
		\g5080_reg/NET0131 ,
		_w2938_,
		_w2939_
	);
	LUT2 #(
		.INIT('h4)
	) name2166 (
		\g5073_reg/NET0131 ,
		\g5077_reg/NET0131 ,
		_w2940_
	);
	LUT2 #(
		.INIT('h4)
	) name2167 (
		\g5069_reg/NET0131 ,
		\g5077_reg/NET0131 ,
		_w2941_
	);
	LUT2 #(
		.INIT('h1)
	) name2168 (
		\g5080_reg/NET0131 ,
		\g5084_reg/NET0131 ,
		_w2942_
	);
	LUT2 #(
		.INIT('h4)
	) name2169 (
		_w2941_,
		_w2942_,
		_w2943_
	);
	LUT2 #(
		.INIT('h1)
	) name2170 (
		_w2940_,
		_w2943_,
		_w2944_
	);
	LUT2 #(
		.INIT('h2)
	) name2171 (
		\g35_pad ,
		_w2944_,
		_w2945_
	);
	LUT2 #(
		.INIT('h1)
	) name2172 (
		_w2939_,
		_w2945_,
		_w2946_
	);
	LUT2 #(
		.INIT('h2)
	) name2173 (
		\g2831_reg/NET0131 ,
		\g35_pad ,
		_w2947_
	);
	LUT2 #(
		.INIT('h2)
	) name2174 (
		\g1945_reg/NET0131 ,
		\g2715_reg/NET0131 ,
		_w2948_
	);
	LUT2 #(
		.INIT('h8)
	) name2175 (
		\g2079_reg/NET0131 ,
		\g2715_reg/NET0131 ,
		_w2949_
	);
	LUT2 #(
		.INIT('h2)
	) name2176 (
		\g2719_reg/NET0131 ,
		_w2948_,
		_w2950_
	);
	LUT2 #(
		.INIT('h4)
	) name2177 (
		_w2949_,
		_w2950_,
		_w2951_
	);
	LUT2 #(
		.INIT('h2)
	) name2178 (
		\g1677_reg/NET0131 ,
		\g2715_reg/NET0131 ,
		_w2952_
	);
	LUT2 #(
		.INIT('h8)
	) name2179 (
		\g1811_reg/NET0131 ,
		\g2715_reg/NET0131 ,
		_w2953_
	);
	LUT2 #(
		.INIT('h1)
	) name2180 (
		\g2719_reg/NET0131 ,
		_w2952_,
		_w2954_
	);
	LUT2 #(
		.INIT('h4)
	) name2181 (
		_w2953_,
		_w2954_,
		_w2955_
	);
	LUT2 #(
		.INIT('h1)
	) name2182 (
		_w2951_,
		_w2955_,
		_w2956_
	);
	LUT2 #(
		.INIT('h4)
	) name2183 (
		\g2735_reg/NET0131 ,
		_w2501_,
		_w2957_
	);
	LUT2 #(
		.INIT('h8)
	) name2184 (
		_w2503_,
		_w2957_,
		_w2958_
	);
	LUT2 #(
		.INIT('h1)
	) name2185 (
		_w2956_,
		_w2958_,
		_w2959_
	);
	LUT2 #(
		.INIT('h2)
	) name2186 (
		\g2715_reg/NET0131 ,
		\g2787_reg/NET0131 ,
		_w2960_
	);
	LUT2 #(
		.INIT('h1)
	) name2187 (
		\g2715_reg/NET0131 ,
		\g2783_reg/NET0131 ,
		_w2961_
	);
	LUT2 #(
		.INIT('h2)
	) name2188 (
		\g2719_reg/NET0131 ,
		_w2960_,
		_w2962_
	);
	LUT2 #(
		.INIT('h4)
	) name2189 (
		_w2961_,
		_w2962_,
		_w2963_
	);
	LUT2 #(
		.INIT('h1)
	) name2190 (
		\g2715_reg/NET0131 ,
		\g2771_reg/NET0131 ,
		_w2964_
	);
	LUT2 #(
		.INIT('h1)
	) name2191 (
		\g2719_reg/NET0131 ,
		_w2707_,
		_w2965_
	);
	LUT2 #(
		.INIT('h4)
	) name2192 (
		_w2964_,
		_w2965_,
		_w2966_
	);
	LUT2 #(
		.INIT('h1)
	) name2193 (
		_w2963_,
		_w2966_,
		_w2967_
	);
	LUT2 #(
		.INIT('h2)
	) name2194 (
		_w2958_,
		_w2967_,
		_w2968_
	);
	LUT2 #(
		.INIT('h2)
	) name2195 (
		\g35_pad ,
		_w2959_,
		_w2969_
	);
	LUT2 #(
		.INIT('h4)
	) name2196 (
		_w2968_,
		_w2969_,
		_w2970_
	);
	LUT2 #(
		.INIT('h1)
	) name2197 (
		_w2947_,
		_w2970_,
		_w2971_
	);
	LUT2 #(
		.INIT('h4)
	) name2198 (
		\g283_reg/NET0131 ,
		_w2053_,
		_w2972_
	);
	LUT2 #(
		.INIT('h8)
	) name2199 (
		\g287_reg/NET0131 ,
		_w2972_,
		_w2973_
	);
	LUT2 #(
		.INIT('h4)
	) name2200 (
		\g287_reg/NET0131 ,
		_w2044_,
		_w2974_
	);
	LUT2 #(
		.INIT('h2)
	) name2201 (
		\g35_pad ,
		_w2974_,
		_w2975_
	);
	LUT2 #(
		.INIT('h2)
	) name2202 (
		\g283_reg/NET0131 ,
		_w2975_,
		_w2976_
	);
	LUT2 #(
		.INIT('h1)
	) name2203 (
		_w2973_,
		_w2976_,
		_w2977_
	);
	LUT2 #(
		.INIT('h4)
	) name2204 (
		\g1728_reg/NET0131 ,
		\g1772_reg/NET0131 ,
		_w2978_
	);
	LUT2 #(
		.INIT('h4)
	) name2205 (
		\g1792_reg/NET0131 ,
		\g35_pad ,
		_w2979_
	);
	LUT2 #(
		.INIT('h8)
	) name2206 (
		_w2717_,
		_w2979_,
		_w2980_
	);
	LUT2 #(
		.INIT('h4)
	) name2207 (
		_w2978_,
		_w2980_,
		_w2981_
	);
	LUT2 #(
		.INIT('h1)
	) name2208 (
		\g1748_reg/NET0131 ,
		\g35_pad ,
		_w2982_
	);
	LUT2 #(
		.INIT('h4)
	) name2209 (
		\g1768_reg/NET0131 ,
		\g35_pad ,
		_w2983_
	);
	LUT2 #(
		.INIT('h1)
	) name2210 (
		_w2982_,
		_w2983_,
		_w2984_
	);
	LUT2 #(
		.INIT('h4)
	) name2211 (
		_w2980_,
		_w2984_,
		_w2985_
	);
	LUT2 #(
		.INIT('h1)
	) name2212 (
		_w2981_,
		_w2985_,
		_w2986_
	);
	LUT2 #(
		.INIT('h4)
	) name2213 (
		\g749_reg/NET0131 ,
		_w2357_,
		_w2987_
	);
	LUT2 #(
		.INIT('h2)
	) name2214 (
		\g35_pad ,
		_w2987_,
		_w2988_
	);
	LUT2 #(
		.INIT('h2)
	) name2215 (
		\g744_reg/NET0131 ,
		_w2988_,
		_w2989_
	);
	LUT2 #(
		.INIT('h2)
	) name2216 (
		\g35_pad ,
		_w2358_,
		_w2990_
	);
	LUT2 #(
		.INIT('h8)
	) name2217 (
		_w985_,
		_w2990_,
		_w2991_
	);
	LUT2 #(
		.INIT('h1)
	) name2218 (
		_w2989_,
		_w2991_,
		_w2992_
	);
	LUT2 #(
		.INIT('h2)
	) name2219 (
		\g2051_reg/NET0131 ,
		\g2060_reg/NET0131 ,
		_w2993_
	);
	LUT2 #(
		.INIT('h8)
	) name2220 (
		_w2782_,
		_w2993_,
		_w2994_
	);
	LUT2 #(
		.INIT('h1)
	) name2221 (
		\g2036_reg/NET0131 ,
		_w2994_,
		_w2995_
	);
	LUT2 #(
		.INIT('h4)
	) name2222 (
		\g1996_reg/NET0131 ,
		\g2040_reg/NET0131 ,
		_w2996_
	);
	LUT2 #(
		.INIT('h8)
	) name2223 (
		_w2994_,
		_w2996_,
		_w2997_
	);
	LUT2 #(
		.INIT('h1)
	) name2224 (
		_w2995_,
		_w2997_,
		_w2998_
	);
	LUT2 #(
		.INIT('h2)
	) name2225 (
		\g35_pad ,
		_w2998_,
		_w2999_
	);
	LUT2 #(
		.INIT('h1)
	) name2226 (
		\g2016_reg/NET0131 ,
		\g35_pad ,
		_w3000_
	);
	LUT2 #(
		.INIT('h1)
	) name2227 (
		_w2999_,
		_w3000_,
		_w3001_
	);
	LUT2 #(
		.INIT('h2)
	) name2228 (
		\g2834_reg/NET0131 ,
		\g35_pad ,
		_w3002_
	);
	LUT2 #(
		.INIT('h2)
	) name2229 (
		\g2504_reg/NET0131 ,
		\g2715_reg/NET0131 ,
		_w3003_
	);
	LUT2 #(
		.INIT('h8)
	) name2230 (
		\g2638_reg/NET0131 ,
		\g2715_reg/NET0131 ,
		_w3004_
	);
	LUT2 #(
		.INIT('h2)
	) name2231 (
		\g2719_reg/NET0131 ,
		_w3003_,
		_w3005_
	);
	LUT2 #(
		.INIT('h4)
	) name2232 (
		_w3004_,
		_w3005_,
		_w3006_
	);
	LUT2 #(
		.INIT('h2)
	) name2233 (
		\g2236_reg/NET0131 ,
		\g2715_reg/NET0131 ,
		_w3007_
	);
	LUT2 #(
		.INIT('h8)
	) name2234 (
		\g2370_reg/NET0131 ,
		\g2715_reg/NET0131 ,
		_w3008_
	);
	LUT2 #(
		.INIT('h1)
	) name2235 (
		\g2719_reg/NET0131 ,
		_w3007_,
		_w3009_
	);
	LUT2 #(
		.INIT('h4)
	) name2236 (
		_w3008_,
		_w3009_,
		_w3010_
	);
	LUT2 #(
		.INIT('h1)
	) name2237 (
		_w3006_,
		_w3010_,
		_w3011_
	);
	LUT2 #(
		.INIT('h1)
	) name2238 (
		_w2958_,
		_w3011_,
		_w3012_
	);
	LUT2 #(
		.INIT('h2)
	) name2239 (
		\g2715_reg/NET0131 ,
		\g2819_reg/NET0131 ,
		_w3013_
	);
	LUT2 #(
		.INIT('h1)
	) name2240 (
		\g2715_reg/NET0131 ,
		\g2815_reg/NET0131 ,
		_w3014_
	);
	LUT2 #(
		.INIT('h2)
	) name2241 (
		\g2719_reg/NET0131 ,
		_w3013_,
		_w3015_
	);
	LUT2 #(
		.INIT('h4)
	) name2242 (
		_w3014_,
		_w3015_,
		_w3016_
	);
	LUT2 #(
		.INIT('h1)
	) name2243 (
		\g2715_reg/NET0131 ,
		\g2803_reg/NET0131 ,
		_w3017_
	);
	LUT2 #(
		.INIT('h1)
	) name2244 (
		\g2719_reg/NET0131 ,
		_w2572_,
		_w3018_
	);
	LUT2 #(
		.INIT('h4)
	) name2245 (
		_w3017_,
		_w3018_,
		_w3019_
	);
	LUT2 #(
		.INIT('h1)
	) name2246 (
		_w3016_,
		_w3019_,
		_w3020_
	);
	LUT2 #(
		.INIT('h2)
	) name2247 (
		_w2958_,
		_w3020_,
		_w3021_
	);
	LUT2 #(
		.INIT('h2)
	) name2248 (
		\g35_pad ,
		_w3012_,
		_w3022_
	);
	LUT2 #(
		.INIT('h4)
	) name2249 (
		_w3021_,
		_w3022_,
		_w3023_
	);
	LUT2 #(
		.INIT('h1)
	) name2250 (
		_w3002_,
		_w3023_,
		_w3024_
	);
	LUT2 #(
		.INIT('h2)
	) name2251 (
		\g2610_reg/NET0131 ,
		\g2619_reg/NET0131 ,
		_w3025_
	);
	LUT2 #(
		.INIT('h8)
	) name2252 (
		_w2648_,
		_w3025_,
		_w3026_
	);
	LUT2 #(
		.INIT('h1)
	) name2253 (
		\g2595_reg/NET0131 ,
		_w3026_,
		_w3027_
	);
	LUT2 #(
		.INIT('h4)
	) name2254 (
		\g2555_reg/NET0131 ,
		\g2599_reg/NET0131 ,
		_w3028_
	);
	LUT2 #(
		.INIT('h8)
	) name2255 (
		_w3026_,
		_w3028_,
		_w3029_
	);
	LUT2 #(
		.INIT('h1)
	) name2256 (
		_w3027_,
		_w3029_,
		_w3030_
	);
	LUT2 #(
		.INIT('h2)
	) name2257 (
		\g35_pad ,
		_w3030_,
		_w3031_
	);
	LUT2 #(
		.INIT('h1)
	) name2258 (
		\g2575_reg/NET0131 ,
		\g35_pad ,
		_w3032_
	);
	LUT2 #(
		.INIT('h1)
	) name2259 (
		_w3031_,
		_w3032_,
		_w3033_
	);
	LUT2 #(
		.INIT('h2)
	) name2260 (
		\g142_reg/NET0131 ,
		\g35_pad ,
		_w3034_
	);
	LUT2 #(
		.INIT('h1)
	) name2261 (
		\g146_reg/NET0131 ,
		_w2006_,
		_w3035_
	);
	LUT2 #(
		.INIT('h1)
	) name2262 (
		_w2011_,
		_w3035_,
		_w3036_
	);
	LUT2 #(
		.INIT('h8)
	) name2263 (
		_w2024_,
		_w3036_,
		_w3037_
	);
	LUT2 #(
		.INIT('h1)
	) name2264 (
		_w3034_,
		_w3037_,
		_w3038_
	);
	LUT2 #(
		.INIT('h4)
	) name2265 (
		\g35_pad ,
		\g4443_reg/NET0131 ,
		_w3039_
	);
	LUT2 #(
		.INIT('h8)
	) name2266 (
		\g4438_reg/NET0131 ,
		_w1363_,
		_w3040_
	);
	LUT2 #(
		.INIT('h1)
	) name2267 (
		_w3039_,
		_w3040_,
		_w3041_
	);
	LUT2 #(
		.INIT('h4)
	) name2268 (
		_w2642_,
		_w3041_,
		_w3042_
	);
	LUT2 #(
		.INIT('h4)
	) name2269 (
		\g35_pad ,
		\g4801_reg/NET0131 ,
		_w3043_
	);
	LUT2 #(
		.INIT('h8)
	) name2270 (
		\g4793_reg/NET0131 ,
		_w2396_,
		_w3044_
	);
	LUT2 #(
		.INIT('h8)
	) name2271 (
		\g4776_reg/NET0131 ,
		_w3044_,
		_w3045_
	);
	LUT2 #(
		.INIT('h2)
	) name2272 (
		\g35_pad ,
		_w3045_,
		_w3046_
	);
	LUT2 #(
		.INIT('h8)
	) name2273 (
		\g4801_reg/NET0131 ,
		_w3044_,
		_w3047_
	);
	LUT2 #(
		.INIT('h1)
	) name2274 (
		\g4776_reg/NET0131 ,
		_w3047_,
		_w3048_
	);
	LUT2 #(
		.INIT('h2)
	) name2275 (
		_w3046_,
		_w3048_,
		_w3049_
	);
	LUT2 #(
		.INIT('h1)
	) name2276 (
		_w3043_,
		_w3049_,
		_w3050_
	);
	LUT2 #(
		.INIT('h4)
	) name2277 (
		\g35_pad ,
		\g671_reg/NET0131 ,
		_w3051_
	);
	LUT2 #(
		.INIT('h1)
	) name2278 (
		\g676_reg/NET0131 ,
		_w2477_,
		_w3052_
	);
	LUT2 #(
		.INIT('h2)
	) name2279 (
		_w2476_,
		_w2478_,
		_w3053_
	);
	LUT2 #(
		.INIT('h4)
	) name2280 (
		_w3052_,
		_w3053_,
		_w3054_
	);
	LUT2 #(
		.INIT('h1)
	) name2281 (
		_w3051_,
		_w3054_,
		_w3055_
	);
	LUT2 #(
		.INIT('h4)
	) name2282 (
		\g35_pad ,
		\g4659_reg/NET0131 ,
		_w3056_
	);
	LUT2 #(
		.INIT('h1)
	) name2283 (
		\g4664_reg/NET0131 ,
		_w2398_,
		_w3057_
	);
	LUT2 #(
		.INIT('h2)
	) name2284 (
		_w2397_,
		_w2399_,
		_w3058_
	);
	LUT2 #(
		.INIT('h4)
	) name2285 (
		_w3057_,
		_w3058_,
		_w3059_
	);
	LUT2 #(
		.INIT('h1)
	) name2286 (
		_w3056_,
		_w3059_,
		_w3060_
	);
	LUT2 #(
		.INIT('h2)
	) name2287 (
		\g1798_reg/NET0131 ,
		\g35_pad ,
		_w3061_
	);
	LUT2 #(
		.INIT('h4)
	) name2288 (
		\g1792_reg/NET0131 ,
		_w2709_,
		_w3062_
	);
	LUT2 #(
		.INIT('h2)
	) name2289 (
		\g35_pad ,
		_w2711_,
		_w3063_
	);
	LUT2 #(
		.INIT('h4)
	) name2290 (
		_w3062_,
		_w3063_,
		_w3064_
	);
	LUT2 #(
		.INIT('h1)
	) name2291 (
		_w3061_,
		_w3064_,
		_w3065_
	);
	LUT2 #(
		.INIT('h8)
	) name2292 (
		\g35_pad ,
		_w2709_,
		_w3066_
	);
	LUT2 #(
		.INIT('h4)
	) name2293 (
		\g1760_reg/NET0131 ,
		\g1783_reg/NET0131 ,
		_w3067_
	);
	LUT2 #(
		.INIT('h8)
	) name2294 (
		\g1736_reg/NET0131 ,
		_w3067_,
		_w3068_
	);
	LUT2 #(
		.INIT('h2)
	) name2295 (
		\g1748_reg/NET0131 ,
		\g1760_reg/NET0131 ,
		_w3069_
	);
	LUT2 #(
		.INIT('h8)
	) name2296 (
		\g1756_reg/NET0131 ,
		\g1783_reg/NET0131 ,
		_w3070_
	);
	LUT2 #(
		.INIT('h1)
	) name2297 (
		_w3069_,
		_w3070_,
		_w3071_
	);
	LUT2 #(
		.INIT('h1)
	) name2298 (
		\g1792_reg/NET0131 ,
		_w3071_,
		_w3072_
	);
	LUT2 #(
		.INIT('h8)
	) name2299 (
		\g1740_reg/NET0131 ,
		\g1792_reg/NET0131 ,
		_w3073_
	);
	LUT2 #(
		.INIT('h2)
	) name2300 (
		\g1752_reg/NET0131 ,
		\g1783_reg/NET0131 ,
		_w3074_
	);
	LUT2 #(
		.INIT('h1)
	) name2301 (
		_w3073_,
		_w3074_,
		_w3075_
	);
	LUT2 #(
		.INIT('h2)
	) name2302 (
		\g1760_reg/NET0131 ,
		_w3075_,
		_w3076_
	);
	LUT2 #(
		.INIT('h2)
	) name2303 (
		\g1744_reg/NET0131 ,
		\g1783_reg/NET0131 ,
		_w3077_
	);
	LUT2 #(
		.INIT('h8)
	) name2304 (
		\g1792_reg/NET0131 ,
		_w3077_,
		_w3078_
	);
	LUT2 #(
		.INIT('h1)
	) name2305 (
		_w3068_,
		_w3078_,
		_w3079_
	);
	LUT2 #(
		.INIT('h4)
	) name2306 (
		_w3072_,
		_w3079_,
		_w3080_
	);
	LUT2 #(
		.INIT('h4)
	) name2307 (
		_w3076_,
		_w3080_,
		_w3081_
	);
	LUT2 #(
		.INIT('h1)
	) name2308 (
		_w2709_,
		_w3081_,
		_w3082_
	);
	LUT2 #(
		.INIT('h8)
	) name2309 (
		\g1811_reg/NET0131 ,
		_w2709_,
		_w3083_
	);
	LUT2 #(
		.INIT('h1)
	) name2310 (
		_w3082_,
		_w3083_,
		_w3084_
	);
	LUT2 #(
		.INIT('h2)
	) name2311 (
		\g35_pad ,
		_w3084_,
		_w3085_
	);
	LUT2 #(
		.INIT('h2)
	) name2312 (
		\g1792_reg/NET0131 ,
		\g35_pad ,
		_w3086_
	);
	LUT2 #(
		.INIT('h1)
	) name2313 (
		_w3085_,
		_w3086_,
		_w3087_
	);
	LUT2 #(
		.INIT('h2)
	) name2314 (
		\g35_pad ,
		_w2507_,
		_w3088_
	);
	LUT2 #(
		.INIT('h1)
	) name2315 (
		\g1926_reg/NET0131 ,
		_w2507_,
		_w3089_
	);
	LUT2 #(
		.INIT('h1)
	) name2316 (
		_w2746_,
		_w3089_,
		_w3090_
	);
	LUT2 #(
		.INIT('h2)
	) name2317 (
		\g35_pad ,
		_w3090_,
		_w3091_
	);
	LUT2 #(
		.INIT('h1)
	) name2318 (
		\g1932_reg/NET0131 ,
		\g35_pad ,
		_w3092_
	);
	LUT2 #(
		.INIT('h1)
	) name2319 (
		_w3091_,
		_w3092_,
		_w3093_
	);
	LUT2 #(
		.INIT('h8)
	) name2320 (
		\g1870_reg/NET0131 ,
		_w2752_,
		_w3094_
	);
	LUT2 #(
		.INIT('h2)
	) name2321 (
		\g1882_reg/NET0131 ,
		\g1894_reg/NET0131 ,
		_w3095_
	);
	LUT2 #(
		.INIT('h8)
	) name2322 (
		\g1890_reg/NET0131 ,
		\g1917_reg/NET0131 ,
		_w3096_
	);
	LUT2 #(
		.INIT('h1)
	) name2323 (
		_w3095_,
		_w3096_,
		_w3097_
	);
	LUT2 #(
		.INIT('h1)
	) name2324 (
		\g1926_reg/NET0131 ,
		_w3097_,
		_w3098_
	);
	LUT2 #(
		.INIT('h8)
	) name2325 (
		\g1874_reg/NET0131 ,
		\g1926_reg/NET0131 ,
		_w3099_
	);
	LUT2 #(
		.INIT('h2)
	) name2326 (
		\g1886_reg/NET0131 ,
		\g1917_reg/NET0131 ,
		_w3100_
	);
	LUT2 #(
		.INIT('h1)
	) name2327 (
		_w3099_,
		_w3100_,
		_w3101_
	);
	LUT2 #(
		.INIT('h2)
	) name2328 (
		\g1894_reg/NET0131 ,
		_w3101_,
		_w3102_
	);
	LUT2 #(
		.INIT('h2)
	) name2329 (
		\g1878_reg/NET0131 ,
		\g1917_reg/NET0131 ,
		_w3103_
	);
	LUT2 #(
		.INIT('h8)
	) name2330 (
		\g1926_reg/NET0131 ,
		_w3103_,
		_w3104_
	);
	LUT2 #(
		.INIT('h1)
	) name2331 (
		_w3094_,
		_w3104_,
		_w3105_
	);
	LUT2 #(
		.INIT('h4)
	) name2332 (
		_w3098_,
		_w3105_,
		_w3106_
	);
	LUT2 #(
		.INIT('h4)
	) name2333 (
		_w3102_,
		_w3106_,
		_w3107_
	);
	LUT2 #(
		.INIT('h2)
	) name2334 (
		_w2507_,
		_w3107_,
		_w3108_
	);
	LUT2 #(
		.INIT('h2)
	) name2335 (
		\g1945_reg/NET0131 ,
		_w2507_,
		_w3109_
	);
	LUT2 #(
		.INIT('h1)
	) name2336 (
		_w3108_,
		_w3109_,
		_w3110_
	);
	LUT2 #(
		.INIT('h2)
	) name2337 (
		\g35_pad ,
		_w3110_,
		_w3111_
	);
	LUT2 #(
		.INIT('h2)
	) name2338 (
		\g1926_reg/NET0131 ,
		\g35_pad ,
		_w3112_
	);
	LUT2 #(
		.INIT('h1)
	) name2339 (
		_w3111_,
		_w3112_,
		_w3113_
	);
	LUT2 #(
		.INIT('h2)
	) name2340 (
		\g35_pad ,
		_w2782_,
		_w3114_
	);
	LUT2 #(
		.INIT('h2)
	) name2341 (
		\g2066_reg/NET0131 ,
		\g35_pad ,
		_w3115_
	);
	LUT2 #(
		.INIT('h1)
	) name2342 (
		\g2060_reg/NET0131 ,
		_w2782_,
		_w3116_
	);
	LUT2 #(
		.INIT('h2)
	) name2343 (
		\g35_pad ,
		_w2911_,
		_w3117_
	);
	LUT2 #(
		.INIT('h4)
	) name2344 (
		_w3116_,
		_w3117_,
		_w3118_
	);
	LUT2 #(
		.INIT('h1)
	) name2345 (
		_w3115_,
		_w3118_,
		_w3119_
	);
	LUT2 #(
		.INIT('h8)
	) name2346 (
		\g2004_reg/NET0131 ,
		_w2783_,
		_w3120_
	);
	LUT2 #(
		.INIT('h2)
	) name2347 (
		\g2016_reg/NET0131 ,
		\g2028_reg/NET0131 ,
		_w3121_
	);
	LUT2 #(
		.INIT('h8)
	) name2348 (
		\g2024_reg/NET0131 ,
		\g2051_reg/NET0131 ,
		_w3122_
	);
	LUT2 #(
		.INIT('h1)
	) name2349 (
		_w3121_,
		_w3122_,
		_w3123_
	);
	LUT2 #(
		.INIT('h1)
	) name2350 (
		\g2060_reg/NET0131 ,
		_w3123_,
		_w3124_
	);
	LUT2 #(
		.INIT('h8)
	) name2351 (
		\g2008_reg/NET0131 ,
		\g2060_reg/NET0131 ,
		_w3125_
	);
	LUT2 #(
		.INIT('h2)
	) name2352 (
		\g2020_reg/NET0131 ,
		\g2051_reg/NET0131 ,
		_w3126_
	);
	LUT2 #(
		.INIT('h1)
	) name2353 (
		_w3125_,
		_w3126_,
		_w3127_
	);
	LUT2 #(
		.INIT('h2)
	) name2354 (
		\g2028_reg/NET0131 ,
		_w3127_,
		_w3128_
	);
	LUT2 #(
		.INIT('h2)
	) name2355 (
		\g2012_reg/NET0131 ,
		\g2051_reg/NET0131 ,
		_w3129_
	);
	LUT2 #(
		.INIT('h8)
	) name2356 (
		\g2060_reg/NET0131 ,
		_w3129_,
		_w3130_
	);
	LUT2 #(
		.INIT('h1)
	) name2357 (
		_w3120_,
		_w3130_,
		_w3131_
	);
	LUT2 #(
		.INIT('h4)
	) name2358 (
		_w3124_,
		_w3131_,
		_w3132_
	);
	LUT2 #(
		.INIT('h4)
	) name2359 (
		_w3128_,
		_w3132_,
		_w3133_
	);
	LUT2 #(
		.INIT('h2)
	) name2360 (
		_w2782_,
		_w3133_,
		_w3134_
	);
	LUT2 #(
		.INIT('h2)
	) name2361 (
		\g2079_reg/NET0131 ,
		_w2782_,
		_w3135_
	);
	LUT2 #(
		.INIT('h1)
	) name2362 (
		_w3134_,
		_w3135_,
		_w3136_
	);
	LUT2 #(
		.INIT('h2)
	) name2363 (
		\g35_pad ,
		_w3136_,
		_w3137_
	);
	LUT2 #(
		.INIT('h2)
	) name2364 (
		\g2060_reg/NET0131 ,
		\g35_pad ,
		_w3138_
	);
	LUT2 #(
		.INIT('h1)
	) name2365 (
		_w3137_,
		_w3138_,
		_w3139_
	);
	LUT2 #(
		.INIT('h2)
	) name2366 (
		_w2206_,
		_w2540_,
		_w3140_
	);
	LUT2 #(
		.INIT('h2)
	) name2367 (
		\g411_reg/NET0131 ,
		_w2206_,
		_w3141_
	);
	LUT2 #(
		.INIT('h1)
	) name2368 (
		_w3140_,
		_w3141_,
		_w3142_
	);
	LUT2 #(
		.INIT('h2)
	) name2369 (
		\g35_pad ,
		_w3142_,
		_w3143_
	);
	LUT2 #(
		.INIT('h4)
	) name2370 (
		\g35_pad ,
		\g417_reg/NET0131 ,
		_w3144_
	);
	LUT2 #(
		.INIT('h1)
	) name2371 (
		_w3143_,
		_w3144_,
		_w3145_
	);
	LUT2 #(
		.INIT('h2)
	) name2372 (
		\g35_pad ,
		_w2561_,
		_w3146_
	);
	LUT2 #(
		.INIT('h1)
	) name2373 (
		\g2217_reg/NET0131 ,
		_w2561_,
		_w3147_
	);
	LUT2 #(
		.INIT('h1)
	) name2374 (
		_w2917_,
		_w3147_,
		_w3148_
	);
	LUT2 #(
		.INIT('h2)
	) name2375 (
		\g35_pad ,
		_w3148_,
		_w3149_
	);
	LUT2 #(
		.INIT('h1)
	) name2376 (
		\g2223_reg/NET0131 ,
		\g35_pad ,
		_w3150_
	);
	LUT2 #(
		.INIT('h1)
	) name2377 (
		_w3149_,
		_w3150_,
		_w3151_
	);
	LUT2 #(
		.INIT('h8)
	) name2378 (
		\g2181_reg/NET0131 ,
		_w2562_,
		_w3152_
	);
	LUT2 #(
		.INIT('h2)
	) name2379 (
		\g2173_reg/NET0131 ,
		\g2217_reg/NET0131 ,
		_w3153_
	);
	LUT2 #(
		.INIT('h8)
	) name2380 (
		\g2161_reg/NET0131 ,
		\g2208_reg/NET0131 ,
		_w3154_
	);
	LUT2 #(
		.INIT('h1)
	) name2381 (
		_w3153_,
		_w3154_,
		_w3155_
	);
	LUT2 #(
		.INIT('h1)
	) name2382 (
		\g2185_reg/NET0131 ,
		_w3155_,
		_w3156_
	);
	LUT2 #(
		.INIT('h2)
	) name2383 (
		\g2169_reg/NET0131 ,
		\g2208_reg/NET0131 ,
		_w3157_
	);
	LUT2 #(
		.INIT('h8)
	) name2384 (
		\g2165_reg/NET0131 ,
		\g2185_reg/NET0131 ,
		_w3158_
	);
	LUT2 #(
		.INIT('h1)
	) name2385 (
		_w3157_,
		_w3158_,
		_w3159_
	);
	LUT2 #(
		.INIT('h2)
	) name2386 (
		\g2217_reg/NET0131 ,
		_w3159_,
		_w3160_
	);
	LUT2 #(
		.INIT('h8)
	) name2387 (
		\g2177_reg/NET0131 ,
		\g2185_reg/NET0131 ,
		_w3161_
	);
	LUT2 #(
		.INIT('h4)
	) name2388 (
		\g2208_reg/NET0131 ,
		_w3161_,
		_w3162_
	);
	LUT2 #(
		.INIT('h1)
	) name2389 (
		_w3152_,
		_w3162_,
		_w3163_
	);
	LUT2 #(
		.INIT('h4)
	) name2390 (
		_w3156_,
		_w3163_,
		_w3164_
	);
	LUT2 #(
		.INIT('h4)
	) name2391 (
		_w3160_,
		_w3164_,
		_w3165_
	);
	LUT2 #(
		.INIT('h2)
	) name2392 (
		_w2561_,
		_w3165_,
		_w3166_
	);
	LUT2 #(
		.INIT('h2)
	) name2393 (
		\g2236_reg/NET0131 ,
		_w2561_,
		_w3167_
	);
	LUT2 #(
		.INIT('h1)
	) name2394 (
		_w3166_,
		_w3167_,
		_w3168_
	);
	LUT2 #(
		.INIT('h2)
	) name2395 (
		\g35_pad ,
		_w3168_,
		_w3169_
	);
	LUT2 #(
		.INIT('h2)
	) name2396 (
		\g2217_reg/NET0131 ,
		\g35_pad ,
		_w3170_
	);
	LUT2 #(
		.INIT('h1)
	) name2397 (
		_w3169_,
		_w3170_,
		_w3171_
	);
	LUT2 #(
		.INIT('h8)
	) name2398 (
		\g35_pad ,
		_w2577_,
		_w3172_
	);
	LUT2 #(
		.INIT('h4)
	) name2399 (
		\g2351_reg/NET0131 ,
		_w2577_,
		_w3173_
	);
	LUT2 #(
		.INIT('h1)
	) name2400 (
		_w2842_,
		_w3173_,
		_w3174_
	);
	LUT2 #(
		.INIT('h2)
	) name2401 (
		\g35_pad ,
		_w3174_,
		_w3175_
	);
	LUT2 #(
		.INIT('h1)
	) name2402 (
		\g2357_reg/NET0131 ,
		\g35_pad ,
		_w3176_
	);
	LUT2 #(
		.INIT('h1)
	) name2403 (
		_w3175_,
		_w3176_,
		_w3177_
	);
	LUT2 #(
		.INIT('h8)
	) name2404 (
		\g2315_reg/NET0131 ,
		_w2578_,
		_w3178_
	);
	LUT2 #(
		.INIT('h2)
	) name2405 (
		\g2307_reg/NET0131 ,
		\g2351_reg/NET0131 ,
		_w3179_
	);
	LUT2 #(
		.INIT('h8)
	) name2406 (
		\g2295_reg/NET0131 ,
		\g2342_reg/NET0131 ,
		_w3180_
	);
	LUT2 #(
		.INIT('h1)
	) name2407 (
		_w3179_,
		_w3180_,
		_w3181_
	);
	LUT2 #(
		.INIT('h1)
	) name2408 (
		\g2319_reg/NET0131 ,
		_w3181_,
		_w3182_
	);
	LUT2 #(
		.INIT('h2)
	) name2409 (
		\g2303_reg/NET0131 ,
		\g2342_reg/NET0131 ,
		_w3183_
	);
	LUT2 #(
		.INIT('h8)
	) name2410 (
		\g2299_reg/NET0131 ,
		\g2319_reg/NET0131 ,
		_w3184_
	);
	LUT2 #(
		.INIT('h1)
	) name2411 (
		_w3183_,
		_w3184_,
		_w3185_
	);
	LUT2 #(
		.INIT('h2)
	) name2412 (
		\g2351_reg/NET0131 ,
		_w3185_,
		_w3186_
	);
	LUT2 #(
		.INIT('h8)
	) name2413 (
		\g2311_reg/NET0131 ,
		\g2319_reg/NET0131 ,
		_w3187_
	);
	LUT2 #(
		.INIT('h4)
	) name2414 (
		\g2342_reg/NET0131 ,
		_w3187_,
		_w3188_
	);
	LUT2 #(
		.INIT('h1)
	) name2415 (
		_w3178_,
		_w3188_,
		_w3189_
	);
	LUT2 #(
		.INIT('h4)
	) name2416 (
		_w3182_,
		_w3189_,
		_w3190_
	);
	LUT2 #(
		.INIT('h4)
	) name2417 (
		_w3186_,
		_w3190_,
		_w3191_
	);
	LUT2 #(
		.INIT('h1)
	) name2418 (
		_w2577_,
		_w3191_,
		_w3192_
	);
	LUT2 #(
		.INIT('h8)
	) name2419 (
		\g2370_reg/NET0131 ,
		_w2577_,
		_w3193_
	);
	LUT2 #(
		.INIT('h1)
	) name2420 (
		_w3192_,
		_w3193_,
		_w3194_
	);
	LUT2 #(
		.INIT('h2)
	) name2421 (
		\g35_pad ,
		_w3194_,
		_w3195_
	);
	LUT2 #(
		.INIT('h2)
	) name2422 (
		\g2351_reg/NET0131 ,
		\g35_pad ,
		_w3196_
	);
	LUT2 #(
		.INIT('h1)
	) name2423 (
		_w3195_,
		_w3196_,
		_w3197_
	);
	LUT2 #(
		.INIT('h2)
	) name2424 (
		\g35_pad ,
		_w2604_,
		_w3198_
	);
	LUT2 #(
		.INIT('h1)
	) name2425 (
		\g2485_reg/NET0131 ,
		_w2604_,
		_w3199_
	);
	LUT2 #(
		.INIT('h1)
	) name2426 (
		_w2877_,
		_w3199_,
		_w3200_
	);
	LUT2 #(
		.INIT('h2)
	) name2427 (
		\g35_pad ,
		_w3200_,
		_w3201_
	);
	LUT2 #(
		.INIT('h1)
	) name2428 (
		\g2491_reg/NET0131 ,
		\g35_pad ,
		_w3202_
	);
	LUT2 #(
		.INIT('h1)
	) name2429 (
		_w3201_,
		_w3202_,
		_w3203_
	);
	LUT2 #(
		.INIT('h8)
	) name2430 (
		\g2449_reg/NET0131 ,
		_w2605_,
		_w3204_
	);
	LUT2 #(
		.INIT('h2)
	) name2431 (
		\g2441_reg/NET0131 ,
		\g2485_reg/NET0131 ,
		_w3205_
	);
	LUT2 #(
		.INIT('h8)
	) name2432 (
		\g2429_reg/NET0131 ,
		\g2476_reg/NET0131 ,
		_w3206_
	);
	LUT2 #(
		.INIT('h1)
	) name2433 (
		_w3205_,
		_w3206_,
		_w3207_
	);
	LUT2 #(
		.INIT('h1)
	) name2434 (
		\g2453_reg/NET0131 ,
		_w3207_,
		_w3208_
	);
	LUT2 #(
		.INIT('h2)
	) name2435 (
		\g2437_reg/NET0131 ,
		\g2476_reg/NET0131 ,
		_w3209_
	);
	LUT2 #(
		.INIT('h8)
	) name2436 (
		\g2433_reg/NET0131 ,
		\g2453_reg/NET0131 ,
		_w3210_
	);
	LUT2 #(
		.INIT('h1)
	) name2437 (
		_w3209_,
		_w3210_,
		_w3211_
	);
	LUT2 #(
		.INIT('h2)
	) name2438 (
		\g2485_reg/NET0131 ,
		_w3211_,
		_w3212_
	);
	LUT2 #(
		.INIT('h8)
	) name2439 (
		\g2445_reg/NET0131 ,
		\g2453_reg/NET0131 ,
		_w3213_
	);
	LUT2 #(
		.INIT('h4)
	) name2440 (
		\g2476_reg/NET0131 ,
		_w3213_,
		_w3214_
	);
	LUT2 #(
		.INIT('h1)
	) name2441 (
		_w3204_,
		_w3214_,
		_w3215_
	);
	LUT2 #(
		.INIT('h4)
	) name2442 (
		_w3208_,
		_w3215_,
		_w3216_
	);
	LUT2 #(
		.INIT('h4)
	) name2443 (
		_w3212_,
		_w3216_,
		_w3217_
	);
	LUT2 #(
		.INIT('h2)
	) name2444 (
		_w2604_,
		_w3217_,
		_w3218_
	);
	LUT2 #(
		.INIT('h2)
	) name2445 (
		\g2504_reg/NET0131 ,
		_w2604_,
		_w3219_
	);
	LUT2 #(
		.INIT('h1)
	) name2446 (
		_w3218_,
		_w3219_,
		_w3220_
	);
	LUT2 #(
		.INIT('h2)
	) name2447 (
		\g35_pad ,
		_w3220_,
		_w3221_
	);
	LUT2 #(
		.INIT('h2)
	) name2448 (
		\g2485_reg/NET0131 ,
		\g35_pad ,
		_w3222_
	);
	LUT2 #(
		.INIT('h1)
	) name2449 (
		_w3221_,
		_w3222_,
		_w3223_
	);
	LUT2 #(
		.INIT('h2)
	) name2450 (
		\g35_pad ,
		_w2616_,
		_w3224_
	);
	LUT2 #(
		.INIT('h1)
	) name2451 (
		\g1657_reg/NET0131 ,
		_w2616_,
		_w3225_
	);
	LUT2 #(
		.INIT('h1)
	) name2452 (
		_w2923_,
		_w3225_,
		_w3226_
	);
	LUT2 #(
		.INIT('h2)
	) name2453 (
		\g35_pad ,
		_w3226_,
		_w3227_
	);
	LUT2 #(
		.INIT('h1)
	) name2454 (
		\g1664_reg/NET0131 ,
		\g35_pad ,
		_w3228_
	);
	LUT2 #(
		.INIT('h1)
	) name2455 (
		_w3227_,
		_w3228_,
		_w3229_
	);
	LUT2 #(
		.INIT('h2)
	) name2456 (
		\g35_pad ,
		_w2648_,
		_w3230_
	);
	LUT2 #(
		.INIT('h8)
	) name2457 (
		\g1600_reg/NET0131 ,
		_w2668_,
		_w3231_
	);
	LUT2 #(
		.INIT('h2)
	) name2458 (
		\g1612_reg/NET0131 ,
		\g1624_reg/NET0131 ,
		_w3232_
	);
	LUT2 #(
		.INIT('h8)
	) name2459 (
		\g1620_reg/NET0131 ,
		\g1648_reg/NET0131 ,
		_w3233_
	);
	LUT2 #(
		.INIT('h1)
	) name2460 (
		_w3232_,
		_w3233_,
		_w3234_
	);
	LUT2 #(
		.INIT('h1)
	) name2461 (
		\g1657_reg/NET0131 ,
		_w3234_,
		_w3235_
	);
	LUT2 #(
		.INIT('h8)
	) name2462 (
		\g1604_reg/NET0131 ,
		\g1657_reg/NET0131 ,
		_w3236_
	);
	LUT2 #(
		.INIT('h2)
	) name2463 (
		\g1616_reg/NET0131 ,
		\g1648_reg/NET0131 ,
		_w3237_
	);
	LUT2 #(
		.INIT('h1)
	) name2464 (
		_w3236_,
		_w3237_,
		_w3238_
	);
	LUT2 #(
		.INIT('h2)
	) name2465 (
		\g1624_reg/NET0131 ,
		_w3238_,
		_w3239_
	);
	LUT2 #(
		.INIT('h2)
	) name2466 (
		\g1608_reg/NET0131 ,
		\g1648_reg/NET0131 ,
		_w3240_
	);
	LUT2 #(
		.INIT('h8)
	) name2467 (
		\g1657_reg/NET0131 ,
		_w3240_,
		_w3241_
	);
	LUT2 #(
		.INIT('h1)
	) name2468 (
		_w3231_,
		_w3241_,
		_w3242_
	);
	LUT2 #(
		.INIT('h4)
	) name2469 (
		_w3235_,
		_w3242_,
		_w3243_
	);
	LUT2 #(
		.INIT('h4)
	) name2470 (
		_w3239_,
		_w3243_,
		_w3244_
	);
	LUT2 #(
		.INIT('h2)
	) name2471 (
		_w2616_,
		_w3244_,
		_w3245_
	);
	LUT2 #(
		.INIT('h2)
	) name2472 (
		\g1677_reg/NET0131 ,
		_w2616_,
		_w3246_
	);
	LUT2 #(
		.INIT('h1)
	) name2473 (
		_w3245_,
		_w3246_,
		_w3247_
	);
	LUT2 #(
		.INIT('h2)
	) name2474 (
		\g35_pad ,
		_w3247_,
		_w3248_
	);
	LUT2 #(
		.INIT('h2)
	) name2475 (
		\g1657_reg/NET0131 ,
		\g35_pad ,
		_w3249_
	);
	LUT2 #(
		.INIT('h1)
	) name2476 (
		_w3248_,
		_w3249_,
		_w3250_
	);
	LUT2 #(
		.INIT('h2)
	) name2477 (
		\g2625_reg/NET0131 ,
		\g35_pad ,
		_w3251_
	);
	LUT2 #(
		.INIT('h1)
	) name2478 (
		\g2619_reg/NET0131 ,
		_w2648_,
		_w3252_
	);
	LUT2 #(
		.INIT('h2)
	) name2479 (
		\g35_pad ,
		_w2929_,
		_w3253_
	);
	LUT2 #(
		.INIT('h4)
	) name2480 (
		_w3252_,
		_w3253_,
		_w3254_
	);
	LUT2 #(
		.INIT('h1)
	) name2481 (
		_w3251_,
		_w3254_,
		_w3255_
	);
	LUT2 #(
		.INIT('h8)
	) name2482 (
		\g2563_reg/NET0131 ,
		_w2649_,
		_w3256_
	);
	LUT2 #(
		.INIT('h2)
	) name2483 (
		\g2575_reg/NET0131 ,
		\g2587_reg/NET0131 ,
		_w3257_
	);
	LUT2 #(
		.INIT('h8)
	) name2484 (
		\g2583_reg/NET0131 ,
		\g2610_reg/NET0131 ,
		_w3258_
	);
	LUT2 #(
		.INIT('h1)
	) name2485 (
		_w3257_,
		_w3258_,
		_w3259_
	);
	LUT2 #(
		.INIT('h1)
	) name2486 (
		\g2619_reg/NET0131 ,
		_w3259_,
		_w3260_
	);
	LUT2 #(
		.INIT('h8)
	) name2487 (
		\g2579_reg/NET0131 ,
		\g2587_reg/NET0131 ,
		_w3261_
	);
	LUT2 #(
		.INIT('h8)
	) name2488 (
		\g2571_reg/NET0131 ,
		\g2619_reg/NET0131 ,
		_w3262_
	);
	LUT2 #(
		.INIT('h1)
	) name2489 (
		_w3261_,
		_w3262_,
		_w3263_
	);
	LUT2 #(
		.INIT('h1)
	) name2490 (
		\g2610_reg/NET0131 ,
		_w3263_,
		_w3264_
	);
	LUT2 #(
		.INIT('h8)
	) name2491 (
		\g2567_reg/NET0131 ,
		\g2587_reg/NET0131 ,
		_w3265_
	);
	LUT2 #(
		.INIT('h8)
	) name2492 (
		\g2619_reg/NET0131 ,
		_w3265_,
		_w3266_
	);
	LUT2 #(
		.INIT('h1)
	) name2493 (
		_w3256_,
		_w3266_,
		_w3267_
	);
	LUT2 #(
		.INIT('h4)
	) name2494 (
		_w3260_,
		_w3267_,
		_w3268_
	);
	LUT2 #(
		.INIT('h4)
	) name2495 (
		_w3264_,
		_w3268_,
		_w3269_
	);
	LUT2 #(
		.INIT('h2)
	) name2496 (
		_w2648_,
		_w3269_,
		_w3270_
	);
	LUT2 #(
		.INIT('h2)
	) name2497 (
		\g2638_reg/NET0131 ,
		_w2648_,
		_w3271_
	);
	LUT2 #(
		.INIT('h1)
	) name2498 (
		_w3270_,
		_w3271_,
		_w3272_
	);
	LUT2 #(
		.INIT('h2)
	) name2499 (
		\g35_pad ,
		_w3272_,
		_w3273_
	);
	LUT2 #(
		.INIT('h2)
	) name2500 (
		\g2619_reg/NET0131 ,
		\g35_pad ,
		_w3274_
	);
	LUT2 #(
		.INIT('h1)
	) name2501 (
		_w3273_,
		_w3274_,
		_w3275_
	);
	LUT2 #(
		.INIT('h8)
	) name2502 (
		\g1691_reg/NET0131 ,
		\g35_pad ,
		_w3276_
	);
	LUT2 #(
		.INIT('h4)
	) name2503 (
		_w2616_,
		_w3276_,
		_w3277_
	);
	LUT2 #(
		.INIT('h4)
	) name2504 (
		_w2668_,
		_w3276_,
		_w3278_
	);
	LUT2 #(
		.INIT('h1)
	) name2505 (
		\g1677_reg/NET0131 ,
		_w3278_,
		_w3279_
	);
	LUT2 #(
		.INIT('h8)
	) name2506 (
		\g1677_reg/NET0131 ,
		_w3278_,
		_w3280_
	);
	LUT2 #(
		.INIT('h1)
	) name2507 (
		_w3279_,
		_w3280_,
		_w3281_
	);
	LUT2 #(
		.INIT('h4)
	) name2508 (
		_w3224_,
		_w3281_,
		_w3282_
	);
	LUT2 #(
		.INIT('h1)
	) name2509 (
		_w3277_,
		_w3282_,
		_w3283_
	);
	LUT2 #(
		.INIT('h8)
	) name2510 (
		\g1825_reg/NET0131 ,
		_w3066_,
		_w3284_
	);
	LUT2 #(
		.INIT('h8)
	) name2511 (
		\g1825_reg/NET0131 ,
		\g35_pad ,
		_w3285_
	);
	LUT2 #(
		.INIT('h4)
	) name2512 (
		_w3067_,
		_w3285_,
		_w3286_
	);
	LUT2 #(
		.INIT('h1)
	) name2513 (
		\g1811_reg/NET0131 ,
		_w3286_,
		_w3287_
	);
	LUT2 #(
		.INIT('h8)
	) name2514 (
		\g1811_reg/NET0131 ,
		_w3286_,
		_w3288_
	);
	LUT2 #(
		.INIT('h1)
	) name2515 (
		_w3287_,
		_w3288_,
		_w3289_
	);
	LUT2 #(
		.INIT('h4)
	) name2516 (
		_w3066_,
		_w3289_,
		_w3290_
	);
	LUT2 #(
		.INIT('h1)
	) name2517 (
		_w3284_,
		_w3290_,
		_w3291_
	);
	LUT2 #(
		.INIT('h2)
	) name2518 (
		\g35_pad ,
		_w2151_,
		_w3292_
	);
	LUT2 #(
		.INIT('h2)
	) name2519 (
		\g316_reg/NET0131 ,
		\g35_pad ,
		_w3293_
	);
	LUT2 #(
		.INIT('h1)
	) name2520 (
		_w3292_,
		_w3293_,
		_w3294_
	);
	LUT2 #(
		.INIT('h8)
	) name2521 (
		\g1018_reg/NET0131 ,
		\g1030_reg/NET0131 ,
		_w3295_
	);
	LUT2 #(
		.INIT('h8)
	) name2522 (
		\g1008_reg/NET0131 ,
		_w3295_,
		_w3296_
	);
	LUT2 #(
		.INIT('h8)
	) name2523 (
		_w2376_,
		_w3296_,
		_w3297_
	);
	LUT2 #(
		.INIT('h2)
	) name2524 (
		\g1008_reg/NET0131 ,
		\g1046_reg/NET0131 ,
		_w3298_
	);
	LUT2 #(
		.INIT('h1)
	) name2525 (
		_w2376_,
		_w3298_,
		_w3299_
	);
	LUT2 #(
		.INIT('h1)
	) name2526 (
		\g969_reg/NET0131 ,
		_w3299_,
		_w3300_
	);
	LUT2 #(
		.INIT('h4)
	) name2527 (
		_w3297_,
		_w3300_,
		_w3301_
	);
	LUT2 #(
		.INIT('h4)
	) name2528 (
		\g1024_reg/NET0131 ,
		_w3301_,
		_w3302_
	);
	LUT2 #(
		.INIT('h8)
	) name2529 (
		\g1002_reg/NET0131 ,
		\g1018_reg/NET0131 ,
		_w3303_
	);
	LUT2 #(
		.INIT('h2)
	) name2530 (
		_w3301_,
		_w3303_,
		_w3304_
	);
	LUT2 #(
		.INIT('h1)
	) name2531 (
		_w2373_,
		_w3304_,
		_w3305_
	);
	LUT2 #(
		.INIT('h4)
	) name2532 (
		_w3302_,
		_w3305_,
		_w3306_
	);
	LUT2 #(
		.INIT('h4)
	) name2533 (
		\g1030_reg/NET0131 ,
		_w3300_,
		_w3307_
	);
	LUT2 #(
		.INIT('h2)
	) name2534 (
		_w3306_,
		_w3307_,
		_w3308_
	);
	LUT2 #(
		.INIT('h4)
	) name2535 (
		\g1036_reg/NET0131 ,
		_w3301_,
		_w3309_
	);
	LUT2 #(
		.INIT('h2)
	) name2536 (
		_w3308_,
		_w3309_,
		_w3310_
	);
	LUT2 #(
		.INIT('h1)
	) name2537 (
		\g1036_reg/NET0131 ,
		_w3308_,
		_w3311_
	);
	LUT2 #(
		.INIT('h1)
	) name2538 (
		_w3310_,
		_w3311_,
		_w3312_
	);
	LUT2 #(
		.INIT('h2)
	) name2539 (
		\g35_pad ,
		_w3312_,
		_w3313_
	);
	LUT2 #(
		.INIT('h1)
	) name2540 (
		\g1030_reg/NET0131 ,
		\g35_pad ,
		_w3314_
	);
	LUT2 #(
		.INIT('h1)
	) name2541 (
		_w3313_,
		_w3314_,
		_w3315_
	);
	LUT2 #(
		.INIT('h8)
	) name2542 (
		\g1959_reg/NET0131 ,
		\g35_pad ,
		_w3316_
	);
	LUT2 #(
		.INIT('h4)
	) name2543 (
		_w2507_,
		_w3316_,
		_w3317_
	);
	LUT2 #(
		.INIT('h4)
	) name2544 (
		_w2752_,
		_w3316_,
		_w3318_
	);
	LUT2 #(
		.INIT('h1)
	) name2545 (
		\g1945_reg/NET0131 ,
		_w3318_,
		_w3319_
	);
	LUT2 #(
		.INIT('h8)
	) name2546 (
		\g1945_reg/NET0131 ,
		_w3318_,
		_w3320_
	);
	LUT2 #(
		.INIT('h1)
	) name2547 (
		_w3319_,
		_w3320_,
		_w3321_
	);
	LUT2 #(
		.INIT('h4)
	) name2548 (
		_w3088_,
		_w3321_,
		_w3322_
	);
	LUT2 #(
		.INIT('h1)
	) name2549 (
		_w3317_,
		_w3322_,
		_w3323_
	);
	LUT2 #(
		.INIT('h8)
	) name2550 (
		\g2250_reg/NET0131 ,
		_w3146_,
		_w3324_
	);
	LUT2 #(
		.INIT('h8)
	) name2551 (
		\g2250_reg/NET0131 ,
		\g35_pad ,
		_w3325_
	);
	LUT2 #(
		.INIT('h4)
	) name2552 (
		_w2812_,
		_w3325_,
		_w3326_
	);
	LUT2 #(
		.INIT('h1)
	) name2553 (
		\g2236_reg/NET0131 ,
		_w3326_,
		_w3327_
	);
	LUT2 #(
		.INIT('h8)
	) name2554 (
		\g2236_reg/NET0131 ,
		_w3326_,
		_w3328_
	);
	LUT2 #(
		.INIT('h1)
	) name2555 (
		_w3327_,
		_w3328_,
		_w3329_
	);
	LUT2 #(
		.INIT('h4)
	) name2556 (
		_w3146_,
		_w3329_,
		_w3330_
	);
	LUT2 #(
		.INIT('h1)
	) name2557 (
		_w3324_,
		_w3330_,
		_w3331_
	);
	LUT2 #(
		.INIT('h8)
	) name2558 (
		\g2384_reg/NET0131 ,
		_w3172_,
		_w3332_
	);
	LUT2 #(
		.INIT('h8)
	) name2559 (
		\g2384_reg/NET0131 ,
		\g35_pad ,
		_w3333_
	);
	LUT2 #(
		.INIT('h4)
	) name2560 (
		_w2848_,
		_w3333_,
		_w3334_
	);
	LUT2 #(
		.INIT('h1)
	) name2561 (
		\g2370_reg/NET0131 ,
		_w3334_,
		_w3335_
	);
	LUT2 #(
		.INIT('h8)
	) name2562 (
		\g2370_reg/NET0131 ,
		_w3334_,
		_w3336_
	);
	LUT2 #(
		.INIT('h1)
	) name2563 (
		_w3335_,
		_w3336_,
		_w3337_
	);
	LUT2 #(
		.INIT('h4)
	) name2564 (
		_w3172_,
		_w3337_,
		_w3338_
	);
	LUT2 #(
		.INIT('h1)
	) name2565 (
		_w3332_,
		_w3338_,
		_w3339_
	);
	LUT2 #(
		.INIT('h8)
	) name2566 (
		\g2518_reg/NET0131 ,
		_w3198_,
		_w3340_
	);
	LUT2 #(
		.INIT('h8)
	) name2567 (
		\g2518_reg/NET0131 ,
		\g35_pad ,
		_w3341_
	);
	LUT2 #(
		.INIT('h4)
	) name2568 (
		_w2883_,
		_w3341_,
		_w3342_
	);
	LUT2 #(
		.INIT('h1)
	) name2569 (
		\g2504_reg/NET0131 ,
		_w3342_,
		_w3343_
	);
	LUT2 #(
		.INIT('h8)
	) name2570 (
		\g2504_reg/NET0131 ,
		_w3342_,
		_w3344_
	);
	LUT2 #(
		.INIT('h1)
	) name2571 (
		_w3343_,
		_w3344_,
		_w3345_
	);
	LUT2 #(
		.INIT('h4)
	) name2572 (
		_w3198_,
		_w3345_,
		_w3346_
	);
	LUT2 #(
		.INIT('h1)
	) name2573 (
		_w3340_,
		_w3346_,
		_w3347_
	);
	LUT2 #(
		.INIT('h4)
	) name2574 (
		\g35_pad ,
		\g739_reg/NET0131 ,
		_w3348_
	);
	LUT2 #(
		.INIT('h8)
	) name2575 (
		\g739_reg/NET0131 ,
		_w2355_,
		_w3349_
	);
	LUT2 #(
		.INIT('h1)
	) name2576 (
		\g744_reg/NET0131 ,
		_w3349_,
		_w3350_
	);
	LUT2 #(
		.INIT('h1)
	) name2577 (
		_w966_,
		_w3350_,
		_w3351_
	);
	LUT2 #(
		.INIT('h8)
	) name2578 (
		_w2990_,
		_w3351_,
		_w3352_
	);
	LUT2 #(
		.INIT('h1)
	) name2579 (
		_w3348_,
		_w3352_,
		_w3353_
	);
	LUT2 #(
		.INIT('h8)
	) name2580 (
		\g2093_reg/NET0131 ,
		_w3114_,
		_w3354_
	);
	LUT2 #(
		.INIT('h8)
	) name2581 (
		\g2093_reg/NET0131 ,
		\g35_pad ,
		_w3355_
	);
	LUT2 #(
		.INIT('h4)
	) name2582 (
		_w2783_,
		_w3355_,
		_w3356_
	);
	LUT2 #(
		.INIT('h1)
	) name2583 (
		\g2079_reg/NET0131 ,
		_w3356_,
		_w3357_
	);
	LUT2 #(
		.INIT('h8)
	) name2584 (
		\g2079_reg/NET0131 ,
		_w3356_,
		_w3358_
	);
	LUT2 #(
		.INIT('h1)
	) name2585 (
		_w3357_,
		_w3358_,
		_w3359_
	);
	LUT2 #(
		.INIT('h4)
	) name2586 (
		_w3114_,
		_w3359_,
		_w3360_
	);
	LUT2 #(
		.INIT('h1)
	) name2587 (
		_w3354_,
		_w3360_,
		_w3361_
	);
	LUT2 #(
		.INIT('h8)
	) name2588 (
		\g2652_reg/NET0131 ,
		_w3230_,
		_w3362_
	);
	LUT2 #(
		.INIT('h8)
	) name2589 (
		\g2652_reg/NET0131 ,
		\g35_pad ,
		_w3363_
	);
	LUT2 #(
		.INIT('h4)
	) name2590 (
		_w2649_,
		_w3363_,
		_w3364_
	);
	LUT2 #(
		.INIT('h1)
	) name2591 (
		\g2638_reg/NET0131 ,
		_w3364_,
		_w3365_
	);
	LUT2 #(
		.INIT('h8)
	) name2592 (
		\g2638_reg/NET0131 ,
		_w3364_,
		_w3366_
	);
	LUT2 #(
		.INIT('h1)
	) name2593 (
		_w3365_,
		_w3366_,
		_w3367_
	);
	LUT2 #(
		.INIT('h4)
	) name2594 (
		_w3230_,
		_w3367_,
		_w3368_
	);
	LUT2 #(
		.INIT('h1)
	) name2595 (
		_w3362_,
		_w3368_,
		_w3369_
	);
	LUT2 #(
		.INIT('h2)
	) name2596 (
		\g358_reg/NET0131 ,
		\g376_reg/NET0131 ,
		_w3370_
	);
	LUT2 #(
		.INIT('h8)
	) name2597 (
		\g385_reg/NET0131 ,
		_w3370_,
		_w3371_
	);
	LUT2 #(
		.INIT('h8)
	) name2598 (
		_w2005_,
		_w3371_,
		_w3372_
	);
	LUT2 #(
		.INIT('h1)
	) name2599 (
		\g528_reg/NET0131 ,
		_w2460_,
		_w3373_
	);
	LUT2 #(
		.INIT('h2)
	) name2600 (
		_w3372_,
		_w3373_,
		_w3374_
	);
	LUT2 #(
		.INIT('h2)
	) name2601 (
		\g667_reg/NET0131 ,
		\g686_reg/NET0131 ,
		_w3375_
	);
	LUT2 #(
		.INIT('h2)
	) name2602 (
		\g490_reg/NET0131 ,
		_w3375_,
		_w3376_
	);
	LUT2 #(
		.INIT('h2)
	) name2603 (
		_w3374_,
		_w3376_,
		_w3377_
	);
	LUT2 #(
		.INIT('h2)
	) name2604 (
		\g35_pad ,
		_w3377_,
		_w3378_
	);
	LUT2 #(
		.INIT('h2)
	) name2605 (
		\g482_reg/NET0131 ,
		_w3378_,
		_w3379_
	);
	LUT2 #(
		.INIT('h1)
	) name2606 (
		\g490_reg/NET0131 ,
		_w3375_,
		_w3380_
	);
	LUT2 #(
		.INIT('h8)
	) name2607 (
		\g482_reg/NET0131 ,
		_w3374_,
		_w3381_
	);
	LUT2 #(
		.INIT('h2)
	) name2608 (
		\g35_pad ,
		_w3380_,
		_w3382_
	);
	LUT2 #(
		.INIT('h4)
	) name2609 (
		_w3381_,
		_w3382_,
		_w3383_
	);
	LUT2 #(
		.INIT('h1)
	) name2610 (
		_w3379_,
		_w3383_,
		_w3384_
	);
	LUT2 #(
		.INIT('h4)
	) name2611 (
		\g35_pad ,
		\g736_reg/NET0131 ,
		_w3385_
	);
	LUT2 #(
		.INIT('h1)
	) name2612 (
		\g739_reg/NET0131 ,
		_w2355_,
		_w3386_
	);
	LUT2 #(
		.INIT('h2)
	) name2613 (
		_w967_,
		_w3349_,
		_w3387_
	);
	LUT2 #(
		.INIT('h4)
	) name2614 (
		_w3386_,
		_w3387_,
		_w3388_
	);
	LUT2 #(
		.INIT('h1)
	) name2615 (
		_w3385_,
		_w3388_,
		_w3389_
	);
	LUT2 #(
		.INIT('h8)
	) name2616 (
		\g1087_reg/NET0131 ,
		\g1205_reg/NET0131 ,
		_w3390_
	);
	LUT2 #(
		.INIT('h8)
	) name2617 (
		\g1221_reg/NET0131 ,
		_w3390_,
		_w3391_
	);
	LUT2 #(
		.INIT('h2)
	) name2618 (
		\g35_pad ,
		_w3391_,
		_w3392_
	);
	LUT2 #(
		.INIT('h8)
	) name2619 (
		\g1211_reg/NET0131 ,
		_w3392_,
		_w3393_
	);
	LUT2 #(
		.INIT('h4)
	) name2620 (
		\g1211_reg/NET0131 ,
		_w3391_,
		_w3394_
	);
	LUT2 #(
		.INIT('h2)
	) name2621 (
		\g35_pad ,
		_w3394_,
		_w3395_
	);
	LUT2 #(
		.INIT('h2)
	) name2622 (
		\g1216_reg/NET0131 ,
		_w3395_,
		_w3396_
	);
	LUT2 #(
		.INIT('h1)
	) name2623 (
		_w3393_,
		_w3396_,
		_w3397_
	);
	LUT2 #(
		.INIT('h2)
	) name2624 (
		\g35_pad ,
		_w2163_,
		_w3398_
	);
	LUT2 #(
		.INIT('h8)
	) name2625 (
		\g4311_reg/NET0131 ,
		_w2161_,
		_w3399_
	);
	LUT2 #(
		.INIT('h8)
	) name2626 (
		\g4322_reg/NET0131 ,
		_w3399_,
		_w3400_
	);
	LUT2 #(
		.INIT('h2)
	) name2627 (
		_w3398_,
		_w3400_,
		_w3401_
	);
	LUT2 #(
		.INIT('h8)
	) name2628 (
		\g4332_reg/NET0131 ,
		_w3401_,
		_w3402_
	);
	LUT2 #(
		.INIT('h4)
	) name2629 (
		\g4332_reg/NET0131 ,
		_w3399_,
		_w3403_
	);
	LUT2 #(
		.INIT('h2)
	) name2630 (
		\g35_pad ,
		_w3403_,
		_w3404_
	);
	LUT2 #(
		.INIT('h2)
	) name2631 (
		\g4322_reg/NET0131 ,
		_w3404_,
		_w3405_
	);
	LUT2 #(
		.INIT('h1)
	) name2632 (
		_w3402_,
		_w3405_,
		_w3406_
	);
	LUT2 #(
		.INIT('h2)
	) name2633 (
		\g1559_reg/NET0131 ,
		\g35_pad ,
		_w3407_
	);
	LUT2 #(
		.INIT('h2)
	) name2634 (
		\g35_pad ,
		_w1382_,
		_w3408_
	);
	LUT2 #(
		.INIT('h8)
	) name2635 (
		\g1559_reg/NET0131 ,
		_w1381_,
		_w3409_
	);
	LUT2 #(
		.INIT('h1)
	) name2636 (
		\g1554_reg/NET0131 ,
		_w3409_,
		_w3410_
	);
	LUT2 #(
		.INIT('h2)
	) name2637 (
		_w3408_,
		_w3410_,
		_w3411_
	);
	LUT2 #(
		.INIT('h1)
	) name2638 (
		_w3407_,
		_w3411_,
		_w3412_
	);
	LUT2 #(
		.INIT('h1)
	) name2639 (
		\g5073_reg/NET0131 ,
		\g5084_reg/NET0131 ,
		_w3413_
	);
	LUT2 #(
		.INIT('h4)
	) name2640 (
		\g5069_reg/NET0131 ,
		\g5084_reg/NET0131 ,
		_w3414_
	);
	LUT2 #(
		.INIT('h2)
	) name2641 (
		\g35_pad ,
		_w3413_,
		_w3415_
	);
	LUT2 #(
		.INIT('h4)
	) name2642 (
		_w3414_,
		_w3415_,
		_w3416_
	);
	LUT2 #(
		.INIT('h2)
	) name2643 (
		\g5077_reg/NET0131 ,
		_w3416_,
		_w3417_
	);
	LUT2 #(
		.INIT('h8)
	) name2644 (
		\g246_reg/NET0131 ,
		\g35_pad ,
		_w3418_
	);
	LUT2 #(
		.INIT('h4)
	) name2645 (
		\g35_pad ,
		\g479_reg/NET0131 ,
		_w3419_
	);
	LUT2 #(
		.INIT('h1)
	) name2646 (
		_w3418_,
		_w3419_,
		_w3420_
	);
	LUT2 #(
		.INIT('h4)
	) name2647 (
		\g35_pad ,
		\g4584_reg/NET0131 ,
		_w3421_
	);
	LUT2 #(
		.INIT('h1)
	) name2648 (
		\g4593_reg/NET0131 ,
		_w2164_,
		_w3422_
	);
	LUT2 #(
		.INIT('h1)
	) name2649 (
		_w2165_,
		_w3422_,
		_w3423_
	);
	LUT2 #(
		.INIT('h8)
	) name2650 (
		_w2169_,
		_w3423_,
		_w3424_
	);
	LUT2 #(
		.INIT('h1)
	) name2651 (
		_w3421_,
		_w3424_,
		_w3425_
	);
	LUT2 #(
		.INIT('h4)
	) name2652 (
		\g862_reg/NET0131 ,
		\g890_reg/NET0131 ,
		_w3426_
	);
	LUT2 #(
		.INIT('h4)
	) name2653 (
		\g896_reg/NET0131 ,
		_w3426_,
		_w3427_
	);
	LUT2 #(
		.INIT('h2)
	) name2654 (
		\g446_reg/NET0131 ,
		_w3427_,
		_w3428_
	);
	LUT2 #(
		.INIT('h8)
	) name2655 (
		\g872_reg/NET0131 ,
		_w3427_,
		_w3429_
	);
	LUT2 #(
		.INIT('h1)
	) name2656 (
		_w3428_,
		_w3429_,
		_w3430_
	);
	LUT2 #(
		.INIT('h2)
	) name2657 (
		\g35_pad ,
		_w3430_,
		_w3431_
	);
	LUT2 #(
		.INIT('h2)
	) name2658 (
		\g246_reg/NET0131 ,
		\g35_pad ,
		_w3432_
	);
	LUT2 #(
		.INIT('h1)
	) name2659 (
		_w3431_,
		_w3432_,
		_w3433_
	);
	LUT2 #(
		.INIT('h2)
	) name2660 (
		\g854_reg/NET0131 ,
		_w2519_,
		_w3434_
	);
	LUT2 #(
		.INIT('h1)
	) name2661 (
		_w2545_,
		_w3434_,
		_w3435_
	);
	LUT2 #(
		.INIT('h2)
	) name2662 (
		\g35_pad ,
		_w3435_,
		_w3436_
	);
	LUT2 #(
		.INIT('h4)
	) name2663 (
		\g35_pad ,
		\g4366_reg/NET0131 ,
		_w3437_
	);
	LUT2 #(
		.INIT('h1)
	) name2664 (
		\g4340_reg/NET0131 ,
		_w1068_,
		_w3438_
	);
	LUT2 #(
		.INIT('h1)
	) name2665 (
		_w2159_,
		_w3438_,
		_w3439_
	);
	LUT2 #(
		.INIT('h8)
	) name2666 (
		\g35_pad ,
		\g4358_reg/NET0131 ,
		_w3440_
	);
	LUT2 #(
		.INIT('h4)
	) name2667 (
		_w3439_,
		_w3440_,
		_w3441_
	);
	LUT2 #(
		.INIT('h2)
	) name2668 (
		\g4349_reg/NET0131 ,
		_w3438_,
		_w3442_
	);
	LUT2 #(
		.INIT('h2)
	) name2669 (
		\g4322_reg/NET0131 ,
		\g4332_reg/NET0131 ,
		_w3443_
	);
	LUT2 #(
		.INIT('h4)
	) name2670 (
		\g4515_reg/NET0131 ,
		_w3443_,
		_w3444_
	);
	LUT2 #(
		.INIT('h2)
	) name2671 (
		\g4311_reg/NET0131 ,
		\g4322_reg/NET0131 ,
		_w3445_
	);
	LUT2 #(
		.INIT('h8)
	) name2672 (
		\g4332_reg/NET0131 ,
		_w3445_,
		_w3446_
	);
	LUT2 #(
		.INIT('h1)
	) name2673 (
		\g4340_reg/NET0131 ,
		\g4349_reg/NET0131 ,
		_w3447_
	);
	LUT2 #(
		.INIT('h4)
	) name2674 (
		_w3444_,
		_w3447_,
		_w3448_
	);
	LUT2 #(
		.INIT('h4)
	) name2675 (
		_w3446_,
		_w3448_,
		_w3449_
	);
	LUT2 #(
		.INIT('h2)
	) name2676 (
		\g35_pad ,
		\g4358_reg/NET0131 ,
		_w3450_
	);
	LUT2 #(
		.INIT('h4)
	) name2677 (
		_w3449_,
		_w3450_,
		_w3451_
	);
	LUT2 #(
		.INIT('h4)
	) name2678 (
		_w3442_,
		_w3451_,
		_w3452_
	);
	LUT2 #(
		.INIT('h1)
	) name2679 (
		_w3437_,
		_w3441_,
		_w3453_
	);
	LUT2 #(
		.INIT('h4)
	) name2680 (
		_w3452_,
		_w3453_,
		_w3454_
	);
	LUT2 #(
		.INIT('h2)
	) name2681 (
		\g1024_reg/NET0131 ,
		\g35_pad ,
		_w3455_
	);
	LUT2 #(
		.INIT('h1)
	) name2682 (
		\g1030_reg/NET0131 ,
		_w3306_,
		_w3456_
	);
	LUT2 #(
		.INIT('h2)
	) name2683 (
		\g35_pad ,
		_w3308_,
		_w3457_
	);
	LUT2 #(
		.INIT('h4)
	) name2684 (
		_w3456_,
		_w3457_,
		_w3458_
	);
	LUT2 #(
		.INIT('h1)
	) name2685 (
		_w3455_,
		_w3458_,
		_w3459_
	);
	LUT2 #(
		.INIT('h8)
	) name2686 (
		\g4785_reg/NET0131 ,
		_w3045_,
		_w3460_
	);
	LUT2 #(
		.INIT('h2)
	) name2687 (
		\g35_pad ,
		_w3460_,
		_w3461_
	);
	LUT2 #(
		.INIT('h8)
	) name2688 (
		\g4709_reg/NET0131 ,
		_w3461_,
		_w3462_
	);
	LUT2 #(
		.INIT('h8)
	) name2689 (
		\g35_pad ,
		\g4709_reg/NET0131 ,
		_w3463_
	);
	LUT2 #(
		.INIT('h2)
	) name2690 (
		\g4785_reg/NET0131 ,
		_w3463_,
		_w3464_
	);
	LUT2 #(
		.INIT('h4)
	) name2691 (
		_w3046_,
		_w3464_,
		_w3465_
	);
	LUT2 #(
		.INIT('h1)
	) name2692 (
		_w3462_,
		_w3465_,
		_w3466_
	);
	LUT2 #(
		.INIT('h1)
	) name2693 (
		\g35_pad ,
		\g843_reg/NET0131 ,
		_w3467_
	);
	LUT2 #(
		.INIT('h8)
	) name2694 (
		\g847_reg/NET0131 ,
		_w2206_,
		_w3468_
	);
	LUT2 #(
		.INIT('h8)
	) name2695 (
		\g843_reg/NET0131 ,
		_w3468_,
		_w3469_
	);
	LUT2 #(
		.INIT('h1)
	) name2696 (
		\g812_reg/NET0131 ,
		_w3469_,
		_w3470_
	);
	LUT2 #(
		.INIT('h8)
	) name2697 (
		\g812_reg/NET0131 ,
		_w3469_,
		_w3471_
	);
	LUT2 #(
		.INIT('h2)
	) name2698 (
		\g837_reg/NET0131 ,
		_w3470_,
		_w3472_
	);
	LUT2 #(
		.INIT('h4)
	) name2699 (
		_w3471_,
		_w3472_,
		_w3473_
	);
	LUT2 #(
		.INIT('h2)
	) name2700 (
		\g35_pad ,
		_w3473_,
		_w3474_
	);
	LUT2 #(
		.INIT('h1)
	) name2701 (
		_w3467_,
		_w3474_,
		_w3475_
	);
	LUT2 #(
		.INIT('h4)
	) name2702 (
		\g35_pad ,
		\g667_reg/NET0131 ,
		_w3476_
	);
	LUT2 #(
		.INIT('h1)
	) name2703 (
		\g671_reg/NET0131 ,
		_w2464_,
		_w3477_
	);
	LUT2 #(
		.INIT('h1)
	) name2704 (
		_w2477_,
		_w3477_,
		_w3478_
	);
	LUT2 #(
		.INIT('h8)
	) name2705 (
		_w2476_,
		_w3478_,
		_w3479_
	);
	LUT2 #(
		.INIT('h1)
	) name2706 (
		_w3476_,
		_w3479_,
		_w3480_
	);
	LUT2 #(
		.INIT('h2)
	) name2707 (
		\g278_reg/NET0131 ,
		\g35_pad ,
		_w3481_
	);
	LUT2 #(
		.INIT('h1)
	) name2708 (
		_w2972_,
		_w3481_,
		_w3482_
	);
	LUT2 #(
		.INIT('h4)
	) name2709 (
		\g35_pad ,
		\g817_reg/NET0131 ,
		_w3483_
	);
	LUT2 #(
		.INIT('h1)
	) name2710 (
		\g832_reg/NET0131 ,
		_w2207_,
		_w3484_
	);
	LUT2 #(
		.INIT('h4)
	) name2711 (
		_w2208_,
		_w2213_,
		_w3485_
	);
	LUT2 #(
		.INIT('h4)
	) name2712 (
		_w3484_,
		_w3485_,
		_w3486_
	);
	LUT2 #(
		.INIT('h1)
	) name2713 (
		_w3483_,
		_w3486_,
		_w3487_
	);
	LUT2 #(
		.INIT('h4)
	) name2714 (
		\g35_pad ,
		\g4793_reg/NET0131 ,
		_w3488_
	);
	LUT2 #(
		.INIT('h1)
	) name2715 (
		\g4801_reg/NET0131 ,
		_w3044_,
		_w3489_
	);
	LUT2 #(
		.INIT('h1)
	) name2716 (
		_w3047_,
		_w3489_,
		_w3490_
	);
	LUT2 #(
		.INIT('h8)
	) name2717 (
		_w3046_,
		_w3490_,
		_w3491_
	);
	LUT2 #(
		.INIT('h1)
	) name2718 (
		_w3488_,
		_w3491_,
		_w3492_
	);
	LUT2 #(
		.INIT('h4)
	) name2719 (
		\g5016_reg/NET0131 ,
		\g5022_reg/NET0131 ,
		_w3493_
	);
	LUT2 #(
		.INIT('h4)
	) name2720 (
		\g5029_reg/NET0131 ,
		_w3493_,
		_w3494_
	);
	LUT2 #(
		.INIT('h4)
	) name2721 (
		\g5033_reg/NET0131 ,
		_w3494_,
		_w3495_
	);
	LUT2 #(
		.INIT('h4)
	) name2722 (
		\g5037_reg/NET0131 ,
		_w3495_,
		_w3496_
	);
	LUT2 #(
		.INIT('h4)
	) name2723 (
		\g5041_reg/NET0131 ,
		_w3496_,
		_w3497_
	);
	LUT2 #(
		.INIT('h4)
	) name2724 (
		\g5046_reg/NET0131 ,
		_w3497_,
		_w3498_
	);
	LUT2 #(
		.INIT('h8)
	) name2725 (
		\g3050_reg/NET0131 ,
		\g5016_reg/NET0131 ,
		_w3499_
	);
	LUT2 #(
		.INIT('h8)
	) name2726 (
		\g5029_reg/NET0131 ,
		_w3499_,
		_w3500_
	);
	LUT2 #(
		.INIT('h8)
	) name2727 (
		\g5033_reg/NET0131 ,
		_w3500_,
		_w3501_
	);
	LUT2 #(
		.INIT('h8)
	) name2728 (
		\g5037_reg/NET0131 ,
		_w3501_,
		_w3502_
	);
	LUT2 #(
		.INIT('h8)
	) name2729 (
		\g5041_reg/NET0131 ,
		_w3502_,
		_w3503_
	);
	LUT2 #(
		.INIT('h8)
	) name2730 (
		\g5046_reg/NET0131 ,
		_w3503_,
		_w3504_
	);
	LUT2 #(
		.INIT('h1)
	) name2731 (
		_w3498_,
		_w3504_,
		_w3505_
	);
	LUT2 #(
		.INIT('h1)
	) name2732 (
		\g5052_reg/NET0131 ,
		_w3505_,
		_w3506_
	);
	LUT2 #(
		.INIT('h8)
	) name2733 (
		\g3050_reg/NET0131 ,
		\g5046_reg/NET0131 ,
		_w3507_
	);
	LUT2 #(
		.INIT('h2)
	) name2734 (
		\g5052_reg/NET0131 ,
		\g5057_reg/NET0131 ,
		_w3508_
	);
	LUT2 #(
		.INIT('h8)
	) name2735 (
		_w3507_,
		_w3508_,
		_w3509_
	);
	LUT2 #(
		.INIT('h2)
	) name2736 (
		\g5052_reg/NET0131 ,
		_w3509_,
		_w3510_
	);
	LUT2 #(
		.INIT('h8)
	) name2737 (
		_w3505_,
		_w3510_,
		_w3511_
	);
	LUT2 #(
		.INIT('h1)
	) name2738 (
		_w3506_,
		_w3511_,
		_w3512_
	);
	LUT2 #(
		.INIT('h2)
	) name2739 (
		\g35_pad ,
		_w3512_,
		_w3513_
	);
	LUT2 #(
		.INIT('h4)
	) name2740 (
		\g35_pad ,
		\g5046_reg/NET0131 ,
		_w3514_
	);
	LUT2 #(
		.INIT('h1)
	) name2741 (
		_w3513_,
		_w3514_,
		_w3515_
	);
	LUT2 #(
		.INIT('h4)
	) name2742 (
		\g691_reg/NET0131 ,
		\g703_reg/NET0131 ,
		_w3516_
	);
	LUT2 #(
		.INIT('h8)
	) name2743 (
		_w2473_,
		_w3516_,
		_w3517_
	);
	LUT2 #(
		.INIT('h2)
	) name2744 (
		_w3371_,
		_w3517_,
		_w3518_
	);
	LUT2 #(
		.INIT('h2)
	) name2745 (
		\g686_reg/NET0131 ,
		_w3371_,
		_w3519_
	);
	LUT2 #(
		.INIT('h1)
	) name2746 (
		_w3518_,
		_w3519_,
		_w3520_
	);
	LUT2 #(
		.INIT('h2)
	) name2747 (
		\g35_pad ,
		_w3520_,
		_w3521_
	);
	LUT2 #(
		.INIT('h4)
	) name2748 (
		\g35_pad ,
		\g691_reg/NET0131 ,
		_w3522_
	);
	LUT2 #(
		.INIT('h1)
	) name2749 (
		_w3521_,
		_w3522_,
		_w3523_
	);
	LUT2 #(
		.INIT('h8)
	) name2750 (
		\g316_reg/NET0131 ,
		\g35_pad ,
		_w3524_
	);
	LUT2 #(
		.INIT('h2)
	) name2751 (
		\g29216_pad ,
		\g35_pad ,
		_w3525_
	);
	LUT2 #(
		.INIT('h1)
	) name2752 (
		_w3524_,
		_w3525_,
		_w3526_
	);
	LUT2 #(
		.INIT('h4)
	) name2753 (
		\g35_pad ,
		\g4776_reg/NET0131 ,
		_w3527_
	);
	LUT2 #(
		.INIT('h1)
	) name2754 (
		\g4785_reg/NET0131 ,
		_w3045_,
		_w3528_
	);
	LUT2 #(
		.INIT('h2)
	) name2755 (
		_w3461_,
		_w3528_,
		_w3529_
	);
	LUT2 #(
		.INIT('h1)
	) name2756 (
		_w3527_,
		_w3529_,
		_w3530_
	);
	LUT2 #(
		.INIT('h2)
	) name2757 (
		\g246_reg/NET0131 ,
		_w3427_,
		_w3531_
	);
	LUT2 #(
		.INIT('h8)
	) name2758 (
		\g14167_pad ,
		_w3427_,
		_w3532_
	);
	LUT2 #(
		.INIT('h1)
	) name2759 (
		_w3531_,
		_w3532_,
		_w3533_
	);
	LUT2 #(
		.INIT('h2)
	) name2760 (
		\g35_pad ,
		_w3533_,
		_w3534_
	);
	LUT2 #(
		.INIT('h2)
	) name2761 (
		\g269_reg/NET0131 ,
		\g35_pad ,
		_w3535_
	);
	LUT2 #(
		.INIT('h1)
	) name2762 (
		_w3534_,
		_w3535_,
		_w3536_
	);
	LUT2 #(
		.INIT('h1)
	) name2763 (
		\g1171_reg/NET0131 ,
		\g7916_pad ,
		_w3537_
	);
	LUT2 #(
		.INIT('h8)
	) name2764 (
		\g1171_reg/NET0131 ,
		\g7916_pad ,
		_w3538_
	);
	LUT2 #(
		.INIT('h1)
	) name2765 (
		_w3537_,
		_w3538_,
		_w3539_
	);
	LUT2 #(
		.INIT('h2)
	) name2766 (
		\g1193_reg/NET0131 ,
		_w1319_,
		_w3540_
	);
	LUT2 #(
		.INIT('h2)
	) name2767 (
		\g1178_reg/NET0131 ,
		\g1189_reg/NET0131 ,
		_w3541_
	);
	LUT2 #(
		.INIT('h8)
	) name2768 (
		\g996_reg/NET0131 ,
		_w3541_,
		_w3542_
	);
	LUT2 #(
		.INIT('h8)
	) name2769 (
		\g1002_reg/NET0131 ,
		\g1024_reg/NET0131 ,
		_w3543_
	);
	LUT2 #(
		.INIT('h8)
	) name2770 (
		\g1036_reg/NET0131 ,
		_w3543_,
		_w3544_
	);
	LUT2 #(
		.INIT('h4)
	) name2771 (
		_w2373_,
		_w2376_,
		_w3545_
	);
	LUT2 #(
		.INIT('h8)
	) name2772 (
		_w3544_,
		_w3545_,
		_w3546_
	);
	LUT2 #(
		.INIT('h2)
	) name2773 (
		_w815_,
		_w3546_,
		_w3547_
	);
	LUT2 #(
		.INIT('h8)
	) name2774 (
		\g7916_pad ,
		_w3542_,
		_w3548_
	);
	LUT2 #(
		.INIT('h4)
	) name2775 (
		_w3547_,
		_w3548_,
		_w3549_
	);
	LUT2 #(
		.INIT('h4)
	) name2776 (
		_w3540_,
		_w3549_,
		_w3550_
	);
	LUT2 #(
		.INIT('h1)
	) name2777 (
		_w3539_,
		_w3550_,
		_w3551_
	);
	LUT2 #(
		.INIT('h2)
	) name2778 (
		\g35_pad ,
		_w3551_,
		_w3552_
	);
	LUT2 #(
		.INIT('h2)
	) name2779 (
		\g1018_reg/NET0131 ,
		\g35_pad ,
		_w3553_
	);
	LUT2 #(
		.INIT('h1)
	) name2780 (
		\g1024_reg/NET0131 ,
		_w3305_,
		_w3554_
	);
	LUT2 #(
		.INIT('h2)
	) name2781 (
		\g35_pad ,
		_w3306_,
		_w3555_
	);
	LUT2 #(
		.INIT('h4)
	) name2782 (
		_w3554_,
		_w3555_,
		_w3556_
	);
	LUT2 #(
		.INIT('h1)
	) name2783 (
		_w3553_,
		_w3556_,
		_w3557_
	);
	LUT2 #(
		.INIT('h8)
	) name2784 (
		\g7916_pad ,
		_w1319_,
		_w3558_
	);
	LUT2 #(
		.INIT('h4)
	) name2785 (
		_w3542_,
		_w3558_,
		_w3559_
	);
	LUT2 #(
		.INIT('h8)
	) name2786 (
		\g1199_reg/NET0131 ,
		_w3559_,
		_w3560_
	);
	LUT2 #(
		.INIT('h2)
	) name2787 (
		\g35_pad ,
		_w3560_,
		_w3561_
	);
	LUT2 #(
		.INIT('h4)
	) name2788 (
		_w3550_,
		_w3561_,
		_w3562_
	);
	LUT2 #(
		.INIT('h8)
	) name2789 (
		\g1070_reg/NET0131 ,
		_w3562_,
		_w3563_
	);
	LUT2 #(
		.INIT('h4)
	) name2790 (
		\g1070_reg/NET0131 ,
		_w3559_,
		_w3564_
	);
	LUT2 #(
		.INIT('h2)
	) name2791 (
		\g35_pad ,
		_w3564_,
		_w3565_
	);
	LUT2 #(
		.INIT('h2)
	) name2792 (
		\g1199_reg/NET0131 ,
		_w3565_,
		_w3566_
	);
	LUT2 #(
		.INIT('h1)
	) name2793 (
		_w3563_,
		_w3566_,
		_w3567_
	);
	LUT2 #(
		.INIT('h4)
	) name2794 (
		\g35_pad ,
		\g5052_reg/NET0131 ,
		_w3568_
	);
	LUT2 #(
		.INIT('h2)
	) name2795 (
		\g5022_reg/NET0131 ,
		\g5046_reg/NET0131 ,
		_w3569_
	);
	LUT2 #(
		.INIT('h4)
	) name2796 (
		\g5052_reg/NET0131 ,
		\g5057_reg/NET0131 ,
		_w3570_
	);
	LUT2 #(
		.INIT('h8)
	) name2797 (
		_w3569_,
		_w3570_,
		_w3571_
	);
	LUT2 #(
		.INIT('h2)
	) name2798 (
		\g35_pad ,
		_w3509_,
		_w3572_
	);
	LUT2 #(
		.INIT('h4)
	) name2799 (
		\g5052_reg/NET0131 ,
		_w3498_,
		_w3573_
	);
	LUT2 #(
		.INIT('h8)
	) name2800 (
		\g5052_reg/NET0131 ,
		_w3504_,
		_w3574_
	);
	LUT2 #(
		.INIT('h1)
	) name2801 (
		_w3573_,
		_w3574_,
		_w3575_
	);
	LUT2 #(
		.INIT('h2)
	) name2802 (
		\g5057_reg/NET0131 ,
		_w3571_,
		_w3576_
	);
	LUT2 #(
		.INIT('h8)
	) name2803 (
		_w3572_,
		_w3576_,
		_w3577_
	);
	LUT2 #(
		.INIT('h8)
	) name2804 (
		_w3575_,
		_w3577_,
		_w3578_
	);
	LUT2 #(
		.INIT('h2)
	) name2805 (
		\g35_pad ,
		\g5057_reg/NET0131 ,
		_w3579_
	);
	LUT2 #(
		.INIT('h4)
	) name2806 (
		_w3575_,
		_w3579_,
		_w3580_
	);
	LUT2 #(
		.INIT('h1)
	) name2807 (
		_w3568_,
		_w3578_,
		_w3581_
	);
	LUT2 #(
		.INIT('h4)
	) name2808 (
		_w3580_,
		_w3581_,
		_w3582_
	);
	LUT2 #(
		.INIT('h4)
	) name2809 (
		_w1492_,
		_w3391_,
		_w3583_
	);
	LUT2 #(
		.INIT('h1)
	) name2810 (
		\g1216_reg/NET0131 ,
		_w3391_,
		_w3584_
	);
	LUT2 #(
		.INIT('h1)
	) name2811 (
		_w3583_,
		_w3584_,
		_w3585_
	);
	LUT2 #(
		.INIT('h2)
	) name2812 (
		\g35_pad ,
		_w3585_,
		_w3586_
	);
	LUT2 #(
		.INIT('h1)
	) name2813 (
		\g1221_reg/NET0131 ,
		\g35_pad ,
		_w3587_
	);
	LUT2 #(
		.INIT('h1)
	) name2814 (
		_w3586_,
		_w3587_,
		_w3588_
	);
	LUT2 #(
		.INIT('h8)
	) name2815 (
		\g3338_reg/NET0131 ,
		\g35_pad ,
		_w3589_
	);
	LUT2 #(
		.INIT('h8)
	) name2816 (
		\g13895_pad ,
		\g3303_reg/NET0131 ,
		_w3590_
	);
	LUT2 #(
		.INIT('h8)
	) name2817 (
		\g16603_pad ,
		\g16718_pad ,
		_w3591_
	);
	LUT2 #(
		.INIT('h8)
	) name2818 (
		_w3590_,
		_w3591_,
		_w3592_
	);
	LUT2 #(
		.INIT('h8)
	) name2819 (
		_w3589_,
		_w3592_,
		_w3593_
	);
	LUT2 #(
		.INIT('h2)
	) name2820 (
		\g3343_reg/NET0131 ,
		_w3593_,
		_w3594_
	);
	LUT2 #(
		.INIT('h2)
	) name2821 (
		\g1564_reg/NET0131 ,
		\g35_pad ,
		_w3595_
	);
	LUT2 #(
		.INIT('h1)
	) name2822 (
		\g1559_reg/NET0131 ,
		_w1381_,
		_w3596_
	);
	LUT2 #(
		.INIT('h1)
	) name2823 (
		_w3409_,
		_w3596_,
		_w3597_
	);
	LUT2 #(
		.INIT('h8)
	) name2824 (
		_w3408_,
		_w3597_,
		_w3598_
	);
	LUT2 #(
		.INIT('h1)
	) name2825 (
		_w3595_,
		_w3598_,
		_w3599_
	);
	LUT2 #(
		.INIT('h2)
	) name2826 (
		\g2771_reg/NET0131 ,
		\g35_pad ,
		_w3600_
	);
	LUT2 #(
		.INIT('h1)
	) name2827 (
		_w2970_,
		_w3600_,
		_w3601_
	);
	LUT2 #(
		.INIT('h2)
	) name2828 (
		\g2803_reg/NET0131 ,
		\g35_pad ,
		_w3602_
	);
	LUT2 #(
		.INIT('h1)
	) name2829 (
		_w3023_,
		_w3602_,
		_w3603_
	);
	LUT2 #(
		.INIT('h8)
	) name2830 (
		_w2158_,
		_w2159_,
		_w3604_
	);
	LUT2 #(
		.INIT('h2)
	) name2831 (
		_w3440_,
		_w3604_,
		_w3605_
	);
	LUT2 #(
		.INIT('h8)
	) name2832 (
		\g4340_reg/NET0131 ,
		_w2158_,
		_w3606_
	);
	LUT2 #(
		.INIT('h2)
	) name2833 (
		\g35_pad ,
		_w3606_,
		_w3607_
	);
	LUT2 #(
		.INIT('h2)
	) name2834 (
		\g4349_reg/NET0131 ,
		_w3440_,
		_w3608_
	);
	LUT2 #(
		.INIT('h4)
	) name2835 (
		_w3607_,
		_w3608_,
		_w3609_
	);
	LUT2 #(
		.INIT('h1)
	) name2836 (
		_w3605_,
		_w3609_,
		_w3610_
	);
	LUT2 #(
		.INIT('h2)
	) name2837 (
		\g336_reg/NET0131 ,
		_w2145_,
		_w3611_
	);
	LUT2 #(
		.INIT('h2)
	) name2838 (
		\g305_reg/NET0131 ,
		_w2144_,
		_w3612_
	);
	LUT2 #(
		.INIT('h1)
	) name2839 (
		_w3611_,
		_w3612_,
		_w3613_
	);
	LUT2 #(
		.INIT('h2)
	) name2840 (
		\g35_pad ,
		_w3613_,
		_w3614_
	);
	LUT2 #(
		.INIT('h2)
	) name2841 (
		\g311_reg/NET0131 ,
		\g35_pad ,
		_w3615_
	);
	LUT2 #(
		.INIT('h1)
	) name2842 (
		_w3614_,
		_w3615_,
		_w3616_
	);
	LUT2 #(
		.INIT('h4)
	) name2843 (
		\g35_pad ,
		\g4311_reg/NET0131 ,
		_w3617_
	);
	LUT2 #(
		.INIT('h1)
	) name2844 (
		\g4322_reg/NET0131 ,
		_w3399_,
		_w3618_
	);
	LUT2 #(
		.INIT('h2)
	) name2845 (
		_w3401_,
		_w3618_,
		_w3619_
	);
	LUT2 #(
		.INIT('h1)
	) name2846 (
		_w3617_,
		_w3619_,
		_w3620_
	);
	LUT2 #(
		.INIT('h2)
	) name2847 (
		\g225_reg/NET0131 ,
		_w3427_,
		_w3621_
	);
	LUT2 #(
		.INIT('h8)
	) name2848 (
		\g14189_pad ,
		_w3427_,
		_w3622_
	);
	LUT2 #(
		.INIT('h1)
	) name2849 (
		_w3621_,
		_w3622_,
		_w3623_
	);
	LUT2 #(
		.INIT('h2)
	) name2850 (
		\g35_pad ,
		_w3623_,
		_w3624_
	);
	LUT2 #(
		.INIT('h4)
	) name2851 (
		\g35_pad ,
		\g872_reg/NET0131 ,
		_w3625_
	);
	LUT2 #(
		.INIT('h1)
	) name2852 (
		_w3624_,
		_w3625_,
		_w3626_
	);
	LUT2 #(
		.INIT('h4)
	) name2853 (
		\g35_pad ,
		\g4653_reg/NET0131 ,
		_w3627_
	);
	LUT2 #(
		.INIT('h1)
	) name2854 (
		\g4659_reg/NET0131 ,
		_w2395_,
		_w3628_
	);
	LUT2 #(
		.INIT('h1)
	) name2855 (
		_w2398_,
		_w3628_,
		_w3629_
	);
	LUT2 #(
		.INIT('h8)
	) name2856 (
		_w2397_,
		_w3629_,
		_w3630_
	);
	LUT2 #(
		.INIT('h1)
	) name2857 (
		_w3627_,
		_w3630_,
		_w3631_
	);
	LUT2 #(
		.INIT('h2)
	) name2858 (
		\g35_pad ,
		_w1960_,
		_w3632_
	);
	LUT2 #(
		.INIT('h2)
	) name2859 (
		\g35_pad ,
		_w1711_,
		_w3633_
	);
	LUT2 #(
		.INIT('h8)
	) name2860 (
		\g2661_reg/NET0131 ,
		_w1711_,
		_w3634_
	);
	LUT2 #(
		.INIT('h2)
	) name2861 (
		\g35_pad ,
		_w3634_,
		_w3635_
	);
	LUT2 #(
		.INIT('h1)
	) name2862 (
		\g2667_reg/NET0131 ,
		_w3635_,
		_w3636_
	);
	LUT2 #(
		.INIT('h1)
	) name2863 (
		\g2671_reg/NET0131 ,
		_w1711_,
		_w3637_
	);
	LUT2 #(
		.INIT('h4)
	) name2864 (
		\g2661_reg/NET0131 ,
		\g2667_reg/NET0131 ,
		_w3638_
	);
	LUT2 #(
		.INIT('h8)
	) name2865 (
		_w1711_,
		_w3638_,
		_w3639_
	);
	LUT2 #(
		.INIT('h1)
	) name2866 (
		_w3637_,
		_w3639_,
		_w3640_
	);
	LUT2 #(
		.INIT('h2)
	) name2867 (
		\g35_pad ,
		_w3640_,
		_w3641_
	);
	LUT2 #(
		.INIT('h1)
	) name2868 (
		_w3636_,
		_w3641_,
		_w3642_
	);
	LUT2 #(
		.INIT('h2)
	) name2869 (
		\g2675_reg/NET0131 ,
		_w1711_,
		_w3643_
	);
	LUT2 #(
		.INIT('h4)
	) name2870 (
		\g2675_reg/NET0131 ,
		_w1711_,
		_w3644_
	);
	LUT2 #(
		.INIT('h1)
	) name2871 (
		_w3643_,
		_w3644_,
		_w3645_
	);
	LUT2 #(
		.INIT('h2)
	) name2872 (
		\g35_pad ,
		_w3645_,
		_w3646_
	);
	LUT2 #(
		.INIT('h2)
	) name2873 (
		\g2671_reg/NET0131 ,
		\g35_pad ,
		_w3647_
	);
	LUT2 #(
		.INIT('h1)
	) name2874 (
		_w3646_,
		_w3647_,
		_w3648_
	);
	LUT2 #(
		.INIT('h2)
	) name2875 (
		\g269_reg/NET0131 ,
		_w3427_,
		_w3649_
	);
	LUT2 #(
		.INIT('h8)
	) name2876 (
		\g14147_pad ,
		_w3427_,
		_w3650_
	);
	LUT2 #(
		.INIT('h1)
	) name2877 (
		_w3649_,
		_w3650_,
		_w3651_
	);
	LUT2 #(
		.INIT('h2)
	) name2878 (
		\g35_pad ,
		_w3651_,
		_w3652_
	);
	LUT2 #(
		.INIT('h2)
	) name2879 (
		\g239_reg/NET0131 ,
		\g35_pad ,
		_w3653_
	);
	LUT2 #(
		.INIT('h1)
	) name2880 (
		_w3652_,
		_w3653_,
		_w3654_
	);
	LUT2 #(
		.INIT('h8)
	) name2881 (
		\g1700_reg/NET0131 ,
		_w1960_,
		_w3655_
	);
	LUT2 #(
		.INIT('h2)
	) name2882 (
		\g35_pad ,
		_w3655_,
		_w3656_
	);
	LUT2 #(
		.INIT('h1)
	) name2883 (
		\g1706_reg/NET0131 ,
		_w3656_,
		_w3657_
	);
	LUT2 #(
		.INIT('h1)
	) name2884 (
		\g1710_reg/NET0131 ,
		_w1960_,
		_w3658_
	);
	LUT2 #(
		.INIT('h4)
	) name2885 (
		\g1700_reg/NET0131 ,
		\g1706_reg/NET0131 ,
		_w3659_
	);
	LUT2 #(
		.INIT('h8)
	) name2886 (
		_w1960_,
		_w3659_,
		_w3660_
	);
	LUT2 #(
		.INIT('h1)
	) name2887 (
		_w3658_,
		_w3660_,
		_w3661_
	);
	LUT2 #(
		.INIT('h2)
	) name2888 (
		\g35_pad ,
		_w3661_,
		_w3662_
	);
	LUT2 #(
		.INIT('h1)
	) name2889 (
		_w3657_,
		_w3662_,
		_w3663_
	);
	LUT2 #(
		.INIT('h8)
	) name2890 (
		_w2294_,
		_w2501_,
		_w3664_
	);
	LUT2 #(
		.INIT('h2)
	) name2891 (
		\g2771_reg/NET0131 ,
		_w3664_,
		_w3665_
	);
	LUT2 #(
		.INIT('h4)
	) name2892 (
		\g2767_reg/NET0131 ,
		_w3664_,
		_w3666_
	);
	LUT2 #(
		.INIT('h1)
	) name2893 (
		_w3665_,
		_w3666_,
		_w3667_
	);
	LUT2 #(
		.INIT('h2)
	) name2894 (
		\g35_pad ,
		_w3667_,
		_w3668_
	);
	LUT2 #(
		.INIT('h2)
	) name2895 (
		\g2775_reg/NET0131 ,
		\g35_pad ,
		_w3669_
	);
	LUT2 #(
		.INIT('h1)
	) name2896 (
		_w3668_,
		_w3669_,
		_w3670_
	);
	LUT2 #(
		.INIT('h2)
	) name2897 (
		\g2724_reg/NET0131 ,
		\g2729_reg/NET0131 ,
		_w3671_
	);
	LUT2 #(
		.INIT('h8)
	) name2898 (
		_w2294_,
		_w3671_,
		_w3672_
	);
	LUT2 #(
		.INIT('h2)
	) name2899 (
		\g2775_reg/NET0131 ,
		_w3672_,
		_w3673_
	);
	LUT2 #(
		.INIT('h4)
	) name2900 (
		\g2779_reg/NET0131 ,
		_w3672_,
		_w3674_
	);
	LUT2 #(
		.INIT('h1)
	) name2901 (
		_w3673_,
		_w3674_,
		_w3675_
	);
	LUT2 #(
		.INIT('h2)
	) name2902 (
		\g35_pad ,
		_w3675_,
		_w3676_
	);
	LUT2 #(
		.INIT('h2)
	) name2903 (
		\g2783_reg/NET0131 ,
		\g35_pad ,
		_w3677_
	);
	LUT2 #(
		.INIT('h1)
	) name2904 (
		_w3676_,
		_w3677_,
		_w3678_
	);
	LUT2 #(
		.INIT('h8)
	) name2905 (
		\g2729_reg/NET0131 ,
		_w2294_,
		_w3679_
	);
	LUT2 #(
		.INIT('h4)
	) name2906 (
		\g2724_reg/NET0131 ,
		_w3679_,
		_w3680_
	);
	LUT2 #(
		.INIT('h2)
	) name2907 (
		\g2783_reg/NET0131 ,
		_w3680_,
		_w3681_
	);
	LUT2 #(
		.INIT('h4)
	) name2908 (
		\g2791_reg/NET0131 ,
		_w3680_,
		_w3682_
	);
	LUT2 #(
		.INIT('h1)
	) name2909 (
		_w3681_,
		_w3682_,
		_w3683_
	);
	LUT2 #(
		.INIT('h2)
	) name2910 (
		\g35_pad ,
		_w3683_,
		_w3684_
	);
	LUT2 #(
		.INIT('h2)
	) name2911 (
		\g2787_reg/NET0131 ,
		\g35_pad ,
		_w3685_
	);
	LUT2 #(
		.INIT('h1)
	) name2912 (
		_w3684_,
		_w3685_,
		_w3686_
	);
	LUT2 #(
		.INIT('h8)
	) name2913 (
		\g2724_reg/NET0131 ,
		_w3679_,
		_w3687_
	);
	LUT2 #(
		.INIT('h2)
	) name2914 (
		\g2787_reg/NET0131 ,
		_w3687_,
		_w3688_
	);
	LUT2 #(
		.INIT('h4)
	) name2915 (
		\g2795_reg/NET0131 ,
		_w3687_,
		_w3689_
	);
	LUT2 #(
		.INIT('h1)
	) name2916 (
		_w3688_,
		_w3689_,
		_w3690_
	);
	LUT2 #(
		.INIT('h2)
	) name2917 (
		\g35_pad ,
		_w3690_,
		_w3691_
	);
	LUT2 #(
		.INIT('h2)
	) name2918 (
		\g2795_reg/NET0131 ,
		\g35_pad ,
		_w3692_
	);
	LUT2 #(
		.INIT('h1)
	) name2919 (
		_w3691_,
		_w3692_,
		_w3693_
	);
	LUT2 #(
		.INIT('h2)
	) name2920 (
		\g1714_reg/NET0131 ,
		_w1960_,
		_w3694_
	);
	LUT2 #(
		.INIT('h4)
	) name2921 (
		\g1714_reg/NET0131 ,
		_w1960_,
		_w3695_
	);
	LUT2 #(
		.INIT('h1)
	) name2922 (
		_w3694_,
		_w3695_,
		_w3696_
	);
	LUT2 #(
		.INIT('h2)
	) name2923 (
		\g35_pad ,
		_w3696_,
		_w3697_
	);
	LUT2 #(
		.INIT('h2)
	) name2924 (
		\g1710_reg/NET0131 ,
		\g35_pad ,
		_w3698_
	);
	LUT2 #(
		.INIT('h1)
	) name2925 (
		_w3697_,
		_w3698_,
		_w3699_
	);
	LUT2 #(
		.INIT('h2)
	) name2926 (
		\g2803_reg/NET0131 ,
		_w3664_,
		_w3700_
	);
	LUT2 #(
		.INIT('h4)
	) name2927 (
		\g2799_reg/NET0131 ,
		_w3664_,
		_w3701_
	);
	LUT2 #(
		.INIT('h1)
	) name2928 (
		_w3700_,
		_w3701_,
		_w3702_
	);
	LUT2 #(
		.INIT('h2)
	) name2929 (
		\g35_pad ,
		_w3702_,
		_w3703_
	);
	LUT2 #(
		.INIT('h2)
	) name2930 (
		\g2807_reg/NET0131 ,
		\g35_pad ,
		_w3704_
	);
	LUT2 #(
		.INIT('h1)
	) name2931 (
		_w3703_,
		_w3704_,
		_w3705_
	);
	LUT2 #(
		.INIT('h2)
	) name2932 (
		\g2807_reg/NET0131 ,
		_w3672_,
		_w3706_
	);
	LUT2 #(
		.INIT('h4)
	) name2933 (
		\g2811_reg/NET0131 ,
		_w3672_,
		_w3707_
	);
	LUT2 #(
		.INIT('h1)
	) name2934 (
		_w3706_,
		_w3707_,
		_w3708_
	);
	LUT2 #(
		.INIT('h2)
	) name2935 (
		\g35_pad ,
		_w3708_,
		_w3709_
	);
	LUT2 #(
		.INIT('h2)
	) name2936 (
		\g2815_reg/NET0131 ,
		\g35_pad ,
		_w3710_
	);
	LUT2 #(
		.INIT('h1)
	) name2937 (
		_w3709_,
		_w3710_,
		_w3711_
	);
	LUT2 #(
		.INIT('h2)
	) name2938 (
		\g2815_reg/NET0131 ,
		_w3680_,
		_w3712_
	);
	LUT2 #(
		.INIT('h4)
	) name2939 (
		\g2823_reg/NET0131 ,
		_w3680_,
		_w3713_
	);
	LUT2 #(
		.INIT('h1)
	) name2940 (
		_w3712_,
		_w3713_,
		_w3714_
	);
	LUT2 #(
		.INIT('h2)
	) name2941 (
		\g35_pad ,
		_w3714_,
		_w3715_
	);
	LUT2 #(
		.INIT('h2)
	) name2942 (
		\g2819_reg/NET0131 ,
		\g35_pad ,
		_w3716_
	);
	LUT2 #(
		.INIT('h1)
	) name2943 (
		_w3715_,
		_w3716_,
		_w3717_
	);
	LUT2 #(
		.INIT('h2)
	) name2944 (
		\g2819_reg/NET0131 ,
		_w3687_,
		_w3718_
	);
	LUT2 #(
		.INIT('h4)
	) name2945 (
		\g2827_reg/NET0131 ,
		_w3687_,
		_w3719_
	);
	LUT2 #(
		.INIT('h1)
	) name2946 (
		_w3718_,
		_w3719_,
		_w3720_
	);
	LUT2 #(
		.INIT('h2)
	) name2947 (
		\g35_pad ,
		_w3720_,
		_w3721_
	);
	LUT2 #(
		.INIT('h2)
	) name2948 (
		\g2827_reg/NET0131 ,
		\g35_pad ,
		_w3722_
	);
	LUT2 #(
		.INIT('h1)
	) name2949 (
		_w3721_,
		_w3722_,
		_w3723_
	);
	LUT2 #(
		.INIT('h2)
	) name2950 (
		\g35_pad ,
		_w1817_,
		_w3724_
	);
	LUT2 #(
		.INIT('h2)
	) name2951 (
		\g1816_reg/NET0131 ,
		_w3724_,
		_w3725_
	);
	LUT2 #(
		.INIT('h8)
	) name2952 (
		\g1821_reg/NET0131 ,
		_w3724_,
		_w3726_
	);
	LUT2 #(
		.INIT('h1)
	) name2953 (
		_w3725_,
		_w3726_,
		_w3727_
	);
	LUT2 #(
		.INIT('h8)
	) name2954 (
		\g1834_reg/NET0131 ,
		_w1817_,
		_w3728_
	);
	LUT2 #(
		.INIT('h2)
	) name2955 (
		\g35_pad ,
		_w3728_,
		_w3729_
	);
	LUT2 #(
		.INIT('h1)
	) name2956 (
		\g1840_reg/NET0131 ,
		_w3729_,
		_w3730_
	);
	LUT2 #(
		.INIT('h1)
	) name2957 (
		\g1844_reg/NET0131 ,
		_w1817_,
		_w3731_
	);
	LUT2 #(
		.INIT('h4)
	) name2958 (
		\g1834_reg/NET0131 ,
		\g1840_reg/NET0131 ,
		_w3732_
	);
	LUT2 #(
		.INIT('h8)
	) name2959 (
		_w1817_,
		_w3732_,
		_w3733_
	);
	LUT2 #(
		.INIT('h1)
	) name2960 (
		_w3731_,
		_w3733_,
		_w3734_
	);
	LUT2 #(
		.INIT('h2)
	) name2961 (
		\g35_pad ,
		_w3734_,
		_w3735_
	);
	LUT2 #(
		.INIT('h1)
	) name2962 (
		_w3730_,
		_w3735_,
		_w3736_
	);
	LUT2 #(
		.INIT('h2)
	) name2963 (
		\g1848_reg/NET0131 ,
		_w1817_,
		_w3737_
	);
	LUT2 #(
		.INIT('h4)
	) name2964 (
		\g1848_reg/NET0131 ,
		_w1817_,
		_w3738_
	);
	LUT2 #(
		.INIT('h1)
	) name2965 (
		_w3737_,
		_w3738_,
		_w3739_
	);
	LUT2 #(
		.INIT('h2)
	) name2966 (
		\g35_pad ,
		_w3739_,
		_w3740_
	);
	LUT2 #(
		.INIT('h2)
	) name2967 (
		\g1844_reg/NET0131 ,
		\g35_pad ,
		_w3741_
	);
	LUT2 #(
		.INIT('h1)
	) name2968 (
		_w3740_,
		_w3741_,
		_w3742_
	);
	LUT2 #(
		.INIT('h2)
	) name2969 (
		\g35_pad ,
		_w1863_,
		_w3743_
	);
	LUT2 #(
		.INIT('h2)
	) name2970 (
		\g1950_reg/NET0131 ,
		_w3743_,
		_w3744_
	);
	LUT2 #(
		.INIT('h8)
	) name2971 (
		\g1955_reg/NET0131 ,
		_w3743_,
		_w3745_
	);
	LUT2 #(
		.INIT('h1)
	) name2972 (
		_w3744_,
		_w3745_,
		_w3746_
	);
	LUT2 #(
		.INIT('h8)
	) name2973 (
		\g1968_reg/NET0131 ,
		_w1863_,
		_w3747_
	);
	LUT2 #(
		.INIT('h2)
	) name2974 (
		\g35_pad ,
		_w3747_,
		_w3748_
	);
	LUT2 #(
		.INIT('h1)
	) name2975 (
		\g1974_reg/NET0131 ,
		_w3748_,
		_w3749_
	);
	LUT2 #(
		.INIT('h1)
	) name2976 (
		\g1978_reg/NET0131 ,
		_w1863_,
		_w3750_
	);
	LUT2 #(
		.INIT('h4)
	) name2977 (
		\g1968_reg/NET0131 ,
		\g1974_reg/NET0131 ,
		_w3751_
	);
	LUT2 #(
		.INIT('h8)
	) name2978 (
		_w1863_,
		_w3751_,
		_w3752_
	);
	LUT2 #(
		.INIT('h1)
	) name2979 (
		_w3750_,
		_w3752_,
		_w3753_
	);
	LUT2 #(
		.INIT('h2)
	) name2980 (
		\g35_pad ,
		_w3753_,
		_w3754_
	);
	LUT2 #(
		.INIT('h1)
	) name2981 (
		_w3749_,
		_w3754_,
		_w3755_
	);
	LUT2 #(
		.INIT('h2)
	) name2982 (
		\g1982_reg/NET0131 ,
		_w1863_,
		_w3756_
	);
	LUT2 #(
		.INIT('h4)
	) name2983 (
		\g1982_reg/NET0131 ,
		_w1863_,
		_w3757_
	);
	LUT2 #(
		.INIT('h1)
	) name2984 (
		_w3756_,
		_w3757_,
		_w3758_
	);
	LUT2 #(
		.INIT('h2)
	) name2985 (
		\g35_pad ,
		_w3758_,
		_w3759_
	);
	LUT2 #(
		.INIT('h2)
	) name2986 (
		\g1978_reg/NET0131 ,
		\g35_pad ,
		_w3760_
	);
	LUT2 #(
		.INIT('h1)
	) name2987 (
		_w3759_,
		_w3760_,
		_w3761_
	);
	LUT2 #(
		.INIT('h2)
	) name2988 (
		\g35_pad ,
		_w1909_,
		_w3762_
	);
	LUT2 #(
		.INIT('h2)
	) name2989 (
		\g2084_reg/NET0131 ,
		_w3762_,
		_w3763_
	);
	LUT2 #(
		.INIT('h8)
	) name2990 (
		\g2089_reg/NET0131 ,
		_w3762_,
		_w3764_
	);
	LUT2 #(
		.INIT('h1)
	) name2991 (
		_w3763_,
		_w3764_,
		_w3765_
	);
	LUT2 #(
		.INIT('h8)
	) name2992 (
		\g2102_reg/NET0131 ,
		_w1909_,
		_w3766_
	);
	LUT2 #(
		.INIT('h2)
	) name2993 (
		\g35_pad ,
		_w3766_,
		_w3767_
	);
	LUT2 #(
		.INIT('h1)
	) name2994 (
		\g2108_reg/NET0131 ,
		_w3767_,
		_w3768_
	);
	LUT2 #(
		.INIT('h1)
	) name2995 (
		\g2112_reg/NET0131 ,
		_w1909_,
		_w3769_
	);
	LUT2 #(
		.INIT('h4)
	) name2996 (
		\g2102_reg/NET0131 ,
		\g2108_reg/NET0131 ,
		_w3770_
	);
	LUT2 #(
		.INIT('h8)
	) name2997 (
		_w1909_,
		_w3770_,
		_w3771_
	);
	LUT2 #(
		.INIT('h1)
	) name2998 (
		_w3769_,
		_w3771_,
		_w3772_
	);
	LUT2 #(
		.INIT('h2)
	) name2999 (
		\g35_pad ,
		_w3772_,
		_w3773_
	);
	LUT2 #(
		.INIT('h1)
	) name3000 (
		_w3768_,
		_w3773_,
		_w3774_
	);
	LUT2 #(
		.INIT('h2)
	) name3001 (
		\g2116_reg/NET0131 ,
		_w1909_,
		_w3775_
	);
	LUT2 #(
		.INIT('h4)
	) name3002 (
		\g2116_reg/NET0131 ,
		_w1909_,
		_w3776_
	);
	LUT2 #(
		.INIT('h1)
	) name3003 (
		_w3775_,
		_w3776_,
		_w3777_
	);
	LUT2 #(
		.INIT('h2)
	) name3004 (
		\g35_pad ,
		_w3777_,
		_w3778_
	);
	LUT2 #(
		.INIT('h2)
	) name3005 (
		\g2112_reg/NET0131 ,
		\g35_pad ,
		_w3779_
	);
	LUT2 #(
		.INIT('h1)
	) name3006 (
		_w3778_,
		_w3779_,
		_w3780_
	);
	LUT2 #(
		.INIT('h2)
	) name3007 (
		\g35_pad ,
		_w1568_,
		_w3781_
	);
	LUT2 #(
		.INIT('h2)
	) name3008 (
		\g2241_reg/NET0131 ,
		_w3781_,
		_w3782_
	);
	LUT2 #(
		.INIT('h8)
	) name3009 (
		\g2246_reg/NET0131 ,
		_w3781_,
		_w3783_
	);
	LUT2 #(
		.INIT('h1)
	) name3010 (
		_w3782_,
		_w3783_,
		_w3784_
	);
	LUT2 #(
		.INIT('h8)
	) name3011 (
		\g2259_reg/NET0131 ,
		_w1568_,
		_w3785_
	);
	LUT2 #(
		.INIT('h2)
	) name3012 (
		\g35_pad ,
		_w3785_,
		_w3786_
	);
	LUT2 #(
		.INIT('h1)
	) name3013 (
		\g2265_reg/NET0131 ,
		_w3786_,
		_w3787_
	);
	LUT2 #(
		.INIT('h1)
	) name3014 (
		\g2269_reg/NET0131 ,
		_w1568_,
		_w3788_
	);
	LUT2 #(
		.INIT('h4)
	) name3015 (
		\g2259_reg/NET0131 ,
		\g2265_reg/NET0131 ,
		_w3789_
	);
	LUT2 #(
		.INIT('h8)
	) name3016 (
		_w1568_,
		_w3789_,
		_w3790_
	);
	LUT2 #(
		.INIT('h1)
	) name3017 (
		_w3788_,
		_w3790_,
		_w3791_
	);
	LUT2 #(
		.INIT('h2)
	) name3018 (
		\g35_pad ,
		_w3791_,
		_w3792_
	);
	LUT2 #(
		.INIT('h1)
	) name3019 (
		_w3787_,
		_w3792_,
		_w3793_
	);
	LUT2 #(
		.INIT('h2)
	) name3020 (
		\g2273_reg/NET0131 ,
		_w1568_,
		_w3794_
	);
	LUT2 #(
		.INIT('h4)
	) name3021 (
		\g2273_reg/NET0131 ,
		_w1568_,
		_w3795_
	);
	LUT2 #(
		.INIT('h1)
	) name3022 (
		_w3794_,
		_w3795_,
		_w3796_
	);
	LUT2 #(
		.INIT('h2)
	) name3023 (
		\g35_pad ,
		_w3796_,
		_w3797_
	);
	LUT2 #(
		.INIT('h2)
	) name3024 (
		\g2269_reg/NET0131 ,
		\g35_pad ,
		_w3798_
	);
	LUT2 #(
		.INIT('h1)
	) name3025 (
		_w3797_,
		_w3798_,
		_w3799_
	);
	LUT2 #(
		.INIT('h2)
	) name3026 (
		\g35_pad ,
		_w1614_,
		_w3800_
	);
	LUT2 #(
		.INIT('h2)
	) name3027 (
		\g2375_reg/NET0131 ,
		_w3800_,
		_w3801_
	);
	LUT2 #(
		.INIT('h8)
	) name3028 (
		\g2380_reg/NET0131 ,
		_w3800_,
		_w3802_
	);
	LUT2 #(
		.INIT('h1)
	) name3029 (
		_w3801_,
		_w3802_,
		_w3803_
	);
	LUT2 #(
		.INIT('h8)
	) name3030 (
		\g2393_reg/NET0131 ,
		_w1614_,
		_w3804_
	);
	LUT2 #(
		.INIT('h2)
	) name3031 (
		\g35_pad ,
		_w3804_,
		_w3805_
	);
	LUT2 #(
		.INIT('h1)
	) name3032 (
		\g2399_reg/NET0131 ,
		_w3805_,
		_w3806_
	);
	LUT2 #(
		.INIT('h1)
	) name3033 (
		\g2403_reg/NET0131 ,
		_w1614_,
		_w3807_
	);
	LUT2 #(
		.INIT('h4)
	) name3034 (
		\g2393_reg/NET0131 ,
		\g2399_reg/NET0131 ,
		_w3808_
	);
	LUT2 #(
		.INIT('h8)
	) name3035 (
		_w1614_,
		_w3808_,
		_w3809_
	);
	LUT2 #(
		.INIT('h1)
	) name3036 (
		_w3807_,
		_w3809_,
		_w3810_
	);
	LUT2 #(
		.INIT('h2)
	) name3037 (
		\g35_pad ,
		_w3810_,
		_w3811_
	);
	LUT2 #(
		.INIT('h1)
	) name3038 (
		_w3806_,
		_w3811_,
		_w3812_
	);
	LUT2 #(
		.INIT('h2)
	) name3039 (
		\g2407_reg/NET0131 ,
		_w1614_,
		_w3813_
	);
	LUT2 #(
		.INIT('h4)
	) name3040 (
		\g2407_reg/NET0131 ,
		_w1614_,
		_w3814_
	);
	LUT2 #(
		.INIT('h1)
	) name3041 (
		_w3813_,
		_w3814_,
		_w3815_
	);
	LUT2 #(
		.INIT('h2)
	) name3042 (
		\g35_pad ,
		_w3815_,
		_w3816_
	);
	LUT2 #(
		.INIT('h2)
	) name3043 (
		\g2403_reg/NET0131 ,
		\g35_pad ,
		_w3817_
	);
	LUT2 #(
		.INIT('h1)
	) name3044 (
		_w3816_,
		_w3817_,
		_w3818_
	);
	LUT2 #(
		.INIT('h2)
	) name3045 (
		\g35_pad ,
		_w1665_,
		_w3819_
	);
	LUT2 #(
		.INIT('h2)
	) name3046 (
		\g2509_reg/NET0131 ,
		_w3819_,
		_w3820_
	);
	LUT2 #(
		.INIT('h8)
	) name3047 (
		\g2514_reg/NET0131 ,
		_w3819_,
		_w3821_
	);
	LUT2 #(
		.INIT('h1)
	) name3048 (
		_w3820_,
		_w3821_,
		_w3822_
	);
	LUT2 #(
		.INIT('h8)
	) name3049 (
		\g2527_reg/NET0131 ,
		_w1665_,
		_w3823_
	);
	LUT2 #(
		.INIT('h2)
	) name3050 (
		\g35_pad ,
		_w3823_,
		_w3824_
	);
	LUT2 #(
		.INIT('h1)
	) name3051 (
		\g2533_reg/NET0131 ,
		_w3824_,
		_w3825_
	);
	LUT2 #(
		.INIT('h1)
	) name3052 (
		\g2537_reg/NET0131 ,
		_w1665_,
		_w3826_
	);
	LUT2 #(
		.INIT('h4)
	) name3053 (
		\g2527_reg/NET0131 ,
		\g2533_reg/NET0131 ,
		_w3827_
	);
	LUT2 #(
		.INIT('h8)
	) name3054 (
		_w1665_,
		_w3827_,
		_w3828_
	);
	LUT2 #(
		.INIT('h1)
	) name3055 (
		_w3826_,
		_w3828_,
		_w3829_
	);
	LUT2 #(
		.INIT('h2)
	) name3056 (
		\g35_pad ,
		_w3829_,
		_w3830_
	);
	LUT2 #(
		.INIT('h1)
	) name3057 (
		_w3825_,
		_w3830_,
		_w3831_
	);
	LUT2 #(
		.INIT('h2)
	) name3058 (
		\g2541_reg/NET0131 ,
		_w1665_,
		_w3832_
	);
	LUT2 #(
		.INIT('h4)
	) name3059 (
		\g2541_reg/NET0131 ,
		_w1665_,
		_w3833_
	);
	LUT2 #(
		.INIT('h1)
	) name3060 (
		_w3832_,
		_w3833_,
		_w3834_
	);
	LUT2 #(
		.INIT('h2)
	) name3061 (
		\g35_pad ,
		_w3834_,
		_w3835_
	);
	LUT2 #(
		.INIT('h2)
	) name3062 (
		\g2537_reg/NET0131 ,
		\g35_pad ,
		_w3836_
	);
	LUT2 #(
		.INIT('h1)
	) name3063 (
		_w3835_,
		_w3836_,
		_w3837_
	);
	LUT2 #(
		.INIT('h2)
	) name3064 (
		\g2643_reg/NET0131 ,
		_w3633_,
		_w3838_
	);
	LUT2 #(
		.INIT('h8)
	) name3065 (
		\g2648_reg/NET0131 ,
		_w3633_,
		_w3839_
	);
	LUT2 #(
		.INIT('h1)
	) name3066 (
		_w3838_,
		_w3839_,
		_w3840_
	);
	LUT2 #(
		.INIT('h2)
	) name3067 (
		\g1668_reg/NET0131 ,
		_w1950_,
		_w3841_
	);
	LUT2 #(
		.INIT('h1)
	) name3068 (
		\g1636_reg/NET0131 ,
		_w1950_,
		_w3842_
	);
	LUT2 #(
		.INIT('h1)
	) name3069 (
		\g1592_reg/NET0131 ,
		_w3842_,
		_w3843_
	);
	LUT2 #(
		.INIT('h2)
	) name3070 (
		\g35_pad ,
		_w3841_,
		_w3844_
	);
	LUT2 #(
		.INIT('h4)
	) name3071 (
		_w3843_,
		_w3844_,
		_w3845_
	);
	LUT2 #(
		.INIT('h2)
	) name3072 (
		\g1046_reg/NET0131 ,
		_w2376_,
		_w3846_
	);
	LUT2 #(
		.INIT('h2)
	) name3073 (
		_w3296_,
		_w3846_,
		_w3847_
	);
	LUT2 #(
		.INIT('h4)
	) name3074 (
		\g1008_reg/NET0131 ,
		_w2376_,
		_w3848_
	);
	LUT2 #(
		.INIT('h8)
	) name3075 (
		_w3544_,
		_w3848_,
		_w3849_
	);
	LUT2 #(
		.INIT('h1)
	) name3076 (
		_w3847_,
		_w3849_,
		_w3850_
	);
	LUT2 #(
		.INIT('h1)
	) name3077 (
		_w2373_,
		_w3850_,
		_w3851_
	);
	LUT2 #(
		.INIT('h2)
	) name3078 (
		\g969_reg/NET0131 ,
		_w2377_,
		_w3852_
	);
	LUT2 #(
		.INIT('h1)
	) name3079 (
		_w3851_,
		_w3852_,
		_w3853_
	);
	LUT2 #(
		.INIT('h2)
	) name3080 (
		\g35_pad ,
		_w3853_,
		_w3854_
	);
	LUT2 #(
		.INIT('h2)
	) name3081 (
		\g2763_reg/NET0131 ,
		\g35_pad ,
		_w3855_
	);
	LUT2 #(
		.INIT('h4)
	) name3082 (
		\g1632_reg/NET0131 ,
		_w2295_,
		_w3856_
	);
	LUT2 #(
		.INIT('h1)
	) name3083 (
		\g2767_reg/NET0131 ,
		_w3856_,
		_w3857_
	);
	LUT2 #(
		.INIT('h2)
	) name3084 (
		_w2291_,
		_w3857_,
		_w3858_
	);
	LUT2 #(
		.INIT('h1)
	) name3085 (
		_w3855_,
		_w3858_,
		_w3859_
	);
	LUT2 #(
		.INIT('h2)
	) name3086 (
		\g2767_reg/NET0131 ,
		\g35_pad ,
		_w3860_
	);
	LUT2 #(
		.INIT('h4)
	) name3087 (
		\g1768_reg/NET0131 ,
		_w2295_,
		_w3861_
	);
	LUT2 #(
		.INIT('h1)
	) name3088 (
		\g2779_reg/NET0131 ,
		_w3861_,
		_w3862_
	);
	LUT2 #(
		.INIT('h2)
	) name3089 (
		_w2291_,
		_w3862_,
		_w3863_
	);
	LUT2 #(
		.INIT('h1)
	) name3090 (
		_w3860_,
		_w3863_,
		_w3864_
	);
	LUT2 #(
		.INIT('h2)
	) name3091 (
		\g2779_reg/NET0131 ,
		\g35_pad ,
		_w3865_
	);
	LUT2 #(
		.INIT('h4)
	) name3092 (
		\g1902_reg/NET0131 ,
		_w2295_,
		_w3866_
	);
	LUT2 #(
		.INIT('h1)
	) name3093 (
		\g2791_reg/NET0131 ,
		_w3866_,
		_w3867_
	);
	LUT2 #(
		.INIT('h2)
	) name3094 (
		_w2291_,
		_w3867_,
		_w3868_
	);
	LUT2 #(
		.INIT('h1)
	) name3095 (
		_w3865_,
		_w3868_,
		_w3869_
	);
	LUT2 #(
		.INIT('h2)
	) name3096 (
		\g2791_reg/NET0131 ,
		\g35_pad ,
		_w3870_
	);
	LUT2 #(
		.INIT('h4)
	) name3097 (
		\g2036_reg/NET0131 ,
		_w2295_,
		_w3871_
	);
	LUT2 #(
		.INIT('h1)
	) name3098 (
		\g2795_reg/NET0131 ,
		_w3871_,
		_w3872_
	);
	LUT2 #(
		.INIT('h2)
	) name3099 (
		_w2291_,
		_w3872_,
		_w3873_
	);
	LUT2 #(
		.INIT('h1)
	) name3100 (
		_w3870_,
		_w3873_,
		_w3874_
	);
	LUT2 #(
		.INIT('h2)
	) name3101 (
		\g2799_reg/NET0131 ,
		\g35_pad ,
		_w3875_
	);
	LUT2 #(
		.INIT('h4)
	) name3102 (
		\g2327_reg/NET0131 ,
		_w2295_,
		_w3876_
	);
	LUT2 #(
		.INIT('h1)
	) name3103 (
		\g2811_reg/NET0131 ,
		_w3876_,
		_w3877_
	);
	LUT2 #(
		.INIT('h2)
	) name3104 (
		_w2291_,
		_w3877_,
		_w3878_
	);
	LUT2 #(
		.INIT('h1)
	) name3105 (
		_w3875_,
		_w3878_,
		_w3879_
	);
	LUT2 #(
		.INIT('h4)
	) name3106 (
		\g1002_reg/NET0131 ,
		_w3301_,
		_w3880_
	);
	LUT2 #(
		.INIT('h1)
	) name3107 (
		_w2373_,
		_w3880_,
		_w3881_
	);
	LUT2 #(
		.INIT('h2)
	) name3108 (
		\g35_pad ,
		_w3881_,
		_w3882_
	);
	LUT2 #(
		.INIT('h8)
	) name3109 (
		\g1018_reg/NET0131 ,
		_w3882_,
		_w3883_
	);
	LUT2 #(
		.INIT('h1)
	) name3110 (
		\g1018_reg/NET0131 ,
		_w2373_,
		_w3884_
	);
	LUT2 #(
		.INIT('h8)
	) name3111 (
		_w3301_,
		_w3884_,
		_w3885_
	);
	LUT2 #(
		.INIT('h2)
	) name3112 (
		\g35_pad ,
		_w3885_,
		_w3886_
	);
	LUT2 #(
		.INIT('h2)
	) name3113 (
		\g1002_reg/NET0131 ,
		_w3886_,
		_w3887_
	);
	LUT2 #(
		.INIT('h1)
	) name3114 (
		_w3883_,
		_w3887_,
		_w3888_
	);
	LUT2 #(
		.INIT('h1)
	) name3115 (
		\g4793_reg/NET0131 ,
		_w2396_,
		_w3889_
	);
	LUT2 #(
		.INIT('h1)
	) name3116 (
		_w3044_,
		_w3889_,
		_w3890_
	);
	LUT2 #(
		.INIT('h8)
	) name3117 (
		_w3046_,
		_w3890_,
		_w3891_
	);
	LUT2 #(
		.INIT('h8)
	) name3118 (
		\g174_reg/NET0131 ,
		\g182_reg/NET0131 ,
		_w3892_
	);
	LUT2 #(
		.INIT('h1)
	) name3119 (
		\g168_reg/NET0131 ,
		_w3892_,
		_w3893_
	);
	LUT2 #(
		.INIT('h2)
	) name3120 (
		\g35_pad ,
		_w2007_,
		_w3894_
	);
	LUT2 #(
		.INIT('h8)
	) name3121 (
		_w2006_,
		_w3894_,
		_w3895_
	);
	LUT2 #(
		.INIT('h4)
	) name3122 (
		_w3893_,
		_w3895_,
		_w3896_
	);
	LUT2 #(
		.INIT('h2)
	) name3123 (
		\g1189_reg/NET0131 ,
		\g35_pad ,
		_w3897_
	);
	LUT2 #(
		.INIT('h8)
	) name3124 (
		\g1070_reg/NET0131 ,
		_w3560_,
		_w3898_
	);
	LUT2 #(
		.INIT('h2)
	) name3125 (
		\g1193_reg/NET0131 ,
		_w3898_,
		_w3899_
	);
	LUT2 #(
		.INIT('h4)
	) name3126 (
		\g1193_reg/NET0131 ,
		_w3549_,
		_w3900_
	);
	LUT2 #(
		.INIT('h1)
	) name3127 (
		_w3899_,
		_w3900_,
		_w3901_
	);
	LUT2 #(
		.INIT('h2)
	) name3128 (
		\g35_pad ,
		_w3901_,
		_w3902_
	);
	LUT2 #(
		.INIT('h1)
	) name3129 (
		_w3897_,
		_w3902_,
		_w3903_
	);
	LUT2 #(
		.INIT('h2)
	) name3130 (
		\g29218_pad ,
		\g35_pad ,
		_w3904_
	);
	LUT2 #(
		.INIT('h1)
	) name3131 (
		\g4349_reg/NET0131 ,
		\g4358_reg/NET0131 ,
		_w3905_
	);
	LUT2 #(
		.INIT('h8)
	) name3132 (
		_w882_,
		_w3905_,
		_w3906_
	);
	LUT2 #(
		.INIT('h2)
	) name3133 (
		\g35_pad ,
		\g4332_reg/NET0131 ,
		_w3907_
	);
	LUT2 #(
		.INIT('h4)
	) name3134 (
		\g4340_reg/NET0131 ,
		\g4643_reg/NET0131 ,
		_w3908_
	);
	LUT2 #(
		.INIT('h8)
	) name3135 (
		_w3907_,
		_w3908_,
		_w3909_
	);
	LUT2 #(
		.INIT('h8)
	) name3136 (
		_w3906_,
		_w3909_,
		_w3910_
	);
	LUT2 #(
		.INIT('h1)
	) name3137 (
		_w3904_,
		_w3910_,
		_w3911_
	);
	LUT2 #(
		.INIT('h2)
	) name3138 (
		\g2811_reg/NET0131 ,
		\g35_pad ,
		_w3912_
	);
	LUT2 #(
		.INIT('h4)
	) name3139 (
		\g2461_reg/NET0131 ,
		_w2295_,
		_w3913_
	);
	LUT2 #(
		.INIT('h1)
	) name3140 (
		\g2823_reg/NET0131 ,
		_w3913_,
		_w3914_
	);
	LUT2 #(
		.INIT('h2)
	) name3141 (
		_w2291_,
		_w3914_,
		_w3915_
	);
	LUT2 #(
		.INIT('h1)
	) name3142 (
		_w3912_,
		_w3915_,
		_w3916_
	);
	LUT2 #(
		.INIT('h2)
	) name3143 (
		\g2823_reg/NET0131 ,
		\g35_pad ,
		_w3917_
	);
	LUT2 #(
		.INIT('h4)
	) name3144 (
		\g2595_reg/NET0131 ,
		_w2295_,
		_w3918_
	);
	LUT2 #(
		.INIT('h1)
	) name3145 (
		\g2827_reg/NET0131 ,
		_w3918_,
		_w3919_
	);
	LUT2 #(
		.INIT('h2)
	) name3146 (
		_w2291_,
		_w3919_,
		_w3920_
	);
	LUT2 #(
		.INIT('h1)
	) name3147 (
		_w3917_,
		_w3920_,
		_w3921_
	);
	LUT2 #(
		.INIT('h1)
	) name3148 (
		\g2927_reg/NET0131 ,
		\g35_pad ,
		_w3922_
	);
	LUT2 #(
		.INIT('h2)
	) name3149 (
		\g35_pad ,
		\g4072_reg/NET0131 ,
		_w3923_
	);
	LUT2 #(
		.INIT('h1)
	) name3150 (
		\g2941_reg/NET0131 ,
		\g4153_reg/NET0131 ,
		_w3924_
	);
	LUT2 #(
		.INIT('h8)
	) name3151 (
		_w3923_,
		_w3924_,
		_w3925_
	);
	LUT2 #(
		.INIT('h1)
	) name3152 (
		_w3922_,
		_w3925_,
		_w3926_
	);
	LUT2 #(
		.INIT('h2)
	) name3153 (
		\g1193_reg/NET0131 ,
		\g35_pad ,
		_w3927_
	);
	LUT2 #(
		.INIT('h1)
	) name3154 (
		\g1199_reg/NET0131 ,
		_w3559_,
		_w3928_
	);
	LUT2 #(
		.INIT('h2)
	) name3155 (
		_w3562_,
		_w3928_,
		_w3929_
	);
	LUT2 #(
		.INIT('h1)
	) name3156 (
		_w3927_,
		_w3929_,
		_w3930_
	);
	LUT2 #(
		.INIT('h2)
	) name3157 (
		\g3329_reg/NET0131 ,
		\g35_pad ,
		_w3931_
	);
	LUT2 #(
		.INIT('h1)
	) name3158 (
		\g3338_reg/NET0131 ,
		_w3592_,
		_w3932_
	);
	LUT2 #(
		.INIT('h8)
	) name3159 (
		\g3338_reg/NET0131 ,
		_w3592_,
		_w3933_
	);
	LUT2 #(
		.INIT('h2)
	) name3160 (
		\g35_pad ,
		_w3933_,
		_w3934_
	);
	LUT2 #(
		.INIT('h4)
	) name3161 (
		_w3932_,
		_w3934_,
		_w3935_
	);
	LUT2 #(
		.INIT('h1)
	) name3162 (
		_w3931_,
		_w3935_,
		_w3936_
	);
	LUT2 #(
		.INIT('h1)
	) name3163 (
		\g843_reg/NET0131 ,
		_w3468_,
		_w3937_
	);
	LUT2 #(
		.INIT('h1)
	) name3164 (
		_w3469_,
		_w3937_,
		_w3938_
	);
	LUT2 #(
		.INIT('h2)
	) name3165 (
		\g35_pad ,
		_w3938_,
		_w3939_
	);
	LUT2 #(
		.INIT('h2)
	) name3166 (
		\g837_reg/NET0131 ,
		_w3939_,
		_w3940_
	);
	LUT2 #(
		.INIT('h1)
	) name3167 (
		\g4584_reg/NET0131 ,
		_w2163_,
		_w3941_
	);
	LUT2 #(
		.INIT('h2)
	) name3168 (
		\g35_pad ,
		_w2164_,
		_w3942_
	);
	LUT2 #(
		.INIT('h4)
	) name3169 (
		_w3941_,
		_w3942_,
		_w3943_
	);
	LUT2 #(
		.INIT('h4)
	) name3170 (
		\g35_pad ,
		\g4332_reg/NET0131 ,
		_w3944_
	);
	LUT2 #(
		.INIT('h1)
	) name3171 (
		_w3943_,
		_w3944_,
		_w3945_
	);
	LUT2 #(
		.INIT('h2)
	) name3172 (
		\g2848_reg/NET0131 ,
		\g35_pad ,
		_w3946_
	);
	LUT2 #(
		.INIT('h4)
	) name3173 (
		\g2856_reg/NET0131 ,
		_w797_,
		_w3947_
	);
	LUT2 #(
		.INIT('h2)
	) name3174 (
		\g35_pad ,
		_w3947_,
		_w3948_
	);
	LUT2 #(
		.INIT('h1)
	) name3175 (
		_w790_,
		_w3946_,
		_w3949_
	);
	LUT2 #(
		.INIT('h4)
	) name3176 (
		_w3948_,
		_w3949_,
		_w3950_
	);
	LUT2 #(
		.INIT('h1)
	) name3177 (
		_w3496_,
		_w3502_,
		_w3951_
	);
	LUT2 #(
		.INIT('h1)
	) name3178 (
		\g5041_reg/NET0131 ,
		_w3951_,
		_w3952_
	);
	LUT2 #(
		.INIT('h1)
	) name3179 (
		_w3509_,
		_w3571_,
		_w3953_
	);
	LUT2 #(
		.INIT('h8)
	) name3180 (
		\g5041_reg/NET0131 ,
		_w3953_,
		_w3954_
	);
	LUT2 #(
		.INIT('h8)
	) name3181 (
		_w3951_,
		_w3954_,
		_w3955_
	);
	LUT2 #(
		.INIT('h1)
	) name3182 (
		_w3952_,
		_w3955_,
		_w3956_
	);
	LUT2 #(
		.INIT('h2)
	) name3183 (
		\g35_pad ,
		_w3956_,
		_w3957_
	);
	LUT2 #(
		.INIT('h4)
	) name3184 (
		\g35_pad ,
		\g5037_reg/NET0131 ,
		_w3958_
	);
	LUT2 #(
		.INIT('h1)
	) name3185 (
		_w3957_,
		_w3958_,
		_w3959_
	);
	LUT2 #(
		.INIT('h2)
	) name3186 (
		\g2898_reg/NET0131 ,
		\g35_pad ,
		_w3960_
	);
	LUT2 #(
		.INIT('h4)
	) name3187 (
		\g2882_reg/NET0131 ,
		_w813_,
		_w3961_
	);
	LUT2 #(
		.INIT('h2)
	) name3188 (
		\g35_pad ,
		_w3961_,
		_w3962_
	);
	LUT2 #(
		.INIT('h1)
	) name3189 (
		_w806_,
		_w3960_,
		_w3963_
	);
	LUT2 #(
		.INIT('h4)
	) name3190 (
		_w3962_,
		_w3963_,
		_w3964_
	);
	LUT2 #(
		.INIT('h8)
	) name3191 (
		_w827_,
		_w894_,
		_w3965_
	);
	LUT2 #(
		.INIT('h8)
	) name3192 (
		_w869_,
		_w3965_,
		_w3966_
	);
	LUT2 #(
		.INIT('h2)
	) name3193 (
		\g35_pad ,
		_w3966_,
		_w3967_
	);
	LUT2 #(
		.INIT('h8)
	) name3194 (
		\g5128_reg/NET0131 ,
		_w3966_,
		_w3968_
	);
	LUT2 #(
		.INIT('h2)
	) name3195 (
		\g35_pad ,
		_w3968_,
		_w3969_
	);
	LUT2 #(
		.INIT('h1)
	) name3196 (
		\g5134_reg/NET0131 ,
		_w3969_,
		_w3970_
	);
	LUT2 #(
		.INIT('h1)
	) name3197 (
		\g5138_reg/NET0131 ,
		_w3966_,
		_w3971_
	);
	LUT2 #(
		.INIT('h4)
	) name3198 (
		\g5128_reg/NET0131 ,
		\g5134_reg/NET0131 ,
		_w3972_
	);
	LUT2 #(
		.INIT('h8)
	) name3199 (
		_w3966_,
		_w3972_,
		_w3973_
	);
	LUT2 #(
		.INIT('h1)
	) name3200 (
		_w3971_,
		_w3973_,
		_w3974_
	);
	LUT2 #(
		.INIT('h2)
	) name3201 (
		\g35_pad ,
		_w3974_,
		_w3975_
	);
	LUT2 #(
		.INIT('h1)
	) name3202 (
		_w3970_,
		_w3975_,
		_w3976_
	);
	LUT2 #(
		.INIT('h2)
	) name3203 (
		\g5142_reg/NET0131 ,
		_w3966_,
		_w3977_
	);
	LUT2 #(
		.INIT('h4)
	) name3204 (
		\g5142_reg/NET0131 ,
		_w3966_,
		_w3978_
	);
	LUT2 #(
		.INIT('h1)
	) name3205 (
		_w3977_,
		_w3978_,
		_w3979_
	);
	LUT2 #(
		.INIT('h2)
	) name3206 (
		\g35_pad ,
		_w3979_,
		_w3980_
	);
	LUT2 #(
		.INIT('h4)
	) name3207 (
		\g35_pad ,
		\g5138_reg/NET0131 ,
		_w3981_
	);
	LUT2 #(
		.INIT('h1)
	) name3208 (
		_w3980_,
		_w3981_,
		_w3982_
	);
	LUT2 #(
		.INIT('h8)
	) name3209 (
		\g1772_reg/NET0131 ,
		_w1499_,
		_w3983_
	);
	LUT2 #(
		.INIT('h1)
	) name3210 (
		_w1824_,
		_w3983_,
		_w3984_
	);
	LUT2 #(
		.INIT('h2)
	) name3211 (
		\g35_pad ,
		_w3984_,
		_w3985_
	);
	LUT2 #(
		.INIT('h2)
	) name3212 (
		\g1779_reg/NET0131 ,
		\g35_pad ,
		_w3986_
	);
	LUT2 #(
		.INIT('h1)
	) name3213 (
		_w3985_,
		_w3986_,
		_w3987_
	);
	LUT2 #(
		.INIT('h2)
	) name3214 (
		\g1772_reg/NET0131 ,
		_w1500_,
		_w3988_
	);
	LUT2 #(
		.INIT('h8)
	) name3215 (
		\g1802_reg/NET0131 ,
		_w1500_,
		_w3989_
	);
	LUT2 #(
		.INIT('h1)
	) name3216 (
		_w3988_,
		_w3989_,
		_w3990_
	);
	LUT2 #(
		.INIT('h8)
	) name3217 (
		\g3352_reg/NET0131 ,
		_w2225_,
		_w3991_
	);
	LUT2 #(
		.INIT('h8)
	) name3218 (
		\g3288_reg/NET0131 ,
		_w894_,
		_w3992_
	);
	LUT2 #(
		.INIT('h8)
	) name3219 (
		_w3991_,
		_w3992_,
		_w3993_
	);
	LUT2 #(
		.INIT('h2)
	) name3220 (
		\g35_pad ,
		_w3993_,
		_w3994_
	);
	LUT2 #(
		.INIT('h8)
	) name3221 (
		\g3119_reg/NET0131 ,
		_w3993_,
		_w3995_
	);
	LUT2 #(
		.INIT('h2)
	) name3222 (
		\g35_pad ,
		_w3995_,
		_w3996_
	);
	LUT2 #(
		.INIT('h1)
	) name3223 (
		\g3125_reg/NET0131 ,
		_w3996_,
		_w3997_
	);
	LUT2 #(
		.INIT('h1)
	) name3224 (
		\g3129_reg/NET0131 ,
		_w3993_,
		_w3998_
	);
	LUT2 #(
		.INIT('h4)
	) name3225 (
		\g3119_reg/NET0131 ,
		\g3125_reg/NET0131 ,
		_w3999_
	);
	LUT2 #(
		.INIT('h8)
	) name3226 (
		_w3993_,
		_w3999_,
		_w4000_
	);
	LUT2 #(
		.INIT('h1)
	) name3227 (
		_w3998_,
		_w4000_,
		_w4001_
	);
	LUT2 #(
		.INIT('h2)
	) name3228 (
		\g35_pad ,
		_w4001_,
		_w4002_
	);
	LUT2 #(
		.INIT('h1)
	) name3229 (
		_w3997_,
		_w4002_,
		_w4003_
	);
	LUT2 #(
		.INIT('h1)
	) name3230 (
		\g3155_reg/NET0131 ,
		\g3161_reg/NET0131 ,
		_w4004_
	);
	LUT2 #(
		.INIT('h4)
	) name3231 (
		\g3167_reg/NET0131 ,
		_w4004_,
		_w4005_
	);
	LUT2 #(
		.INIT('h1)
	) name3232 (
		\g3171_reg/NET0131 ,
		\g3179_reg/NET0131 ,
		_w4006_
	);
	LUT2 #(
		.INIT('h8)
	) name3233 (
		_w4005_,
		_w4006_,
		_w4007_
	);
	LUT2 #(
		.INIT('h2)
	) name3234 (
		\g4180_reg/NET0131 ,
		\g4284_reg/NET0131 ,
		_w4008_
	);
	LUT2 #(
		.INIT('h2)
	) name3235 (
		_w4007_,
		_w4008_,
		_w4009_
	);
	LUT2 #(
		.INIT('h2)
	) name3236 (
		\g3187_reg/NET0131 ,
		_w4007_,
		_w4010_
	);
	LUT2 #(
		.INIT('h1)
	) name3237 (
		_w4009_,
		_w4010_,
		_w4011_
	);
	LUT2 #(
		.INIT('h2)
	) name3238 (
		\g35_pad ,
		_w4011_,
		_w4012_
	);
	LUT2 #(
		.INIT('h2)
	) name3239 (
		\g3179_reg/NET0131 ,
		\g35_pad ,
		_w4013_
	);
	LUT2 #(
		.INIT('h1)
	) name3240 (
		_w4012_,
		_w4013_,
		_w4014_
	);
	LUT2 #(
		.INIT('h2)
	) name3241 (
		\g3171_reg/NET0131 ,
		\g3179_reg/NET0131 ,
		_w4015_
	);
	LUT2 #(
		.INIT('h8)
	) name3242 (
		_w4005_,
		_w4015_,
		_w4016_
	);
	LUT2 #(
		.INIT('h4)
	) name3243 (
		_w4008_,
		_w4016_,
		_w4017_
	);
	LUT2 #(
		.INIT('h2)
	) name3244 (
		\g3191_reg/NET0131 ,
		_w4016_,
		_w4018_
	);
	LUT2 #(
		.INIT('h1)
	) name3245 (
		_w4017_,
		_w4018_,
		_w4019_
	);
	LUT2 #(
		.INIT('h2)
	) name3246 (
		\g35_pad ,
		_w4019_,
		_w4020_
	);
	LUT2 #(
		.INIT('h2)
	) name3247 (
		\g3195_reg/NET0131 ,
		\g35_pad ,
		_w4021_
	);
	LUT2 #(
		.INIT('h1)
	) name3248 (
		_w4020_,
		_w4021_,
		_w4022_
	);
	LUT2 #(
		.INIT('h2)
	) name3249 (
		\g3133_reg/NET0131 ,
		_w3993_,
		_w4023_
	);
	LUT2 #(
		.INIT('h4)
	) name3250 (
		\g3133_reg/NET0131 ,
		_w3993_,
		_w4024_
	);
	LUT2 #(
		.INIT('h1)
	) name3251 (
		_w4023_,
		_w4024_,
		_w4025_
	);
	LUT2 #(
		.INIT('h2)
	) name3252 (
		\g35_pad ,
		_w4025_,
		_w4026_
	);
	LUT2 #(
		.INIT('h2)
	) name3253 (
		\g3129_reg/NET0131 ,
		\g35_pad ,
		_w4027_
	);
	LUT2 #(
		.INIT('h1)
	) name3254 (
		_w4026_,
		_w4027_,
		_w4028_
	);
	LUT2 #(
		.INIT('h8)
	) name3255 (
		\g3167_reg/NET0131 ,
		_w4006_,
		_w4029_
	);
	LUT2 #(
		.INIT('h4)
	) name3256 (
		_w4008_,
		_w4029_,
		_w4030_
	);
	LUT2 #(
		.INIT('h2)
	) name3257 (
		\g3195_reg/NET0131 ,
		_w4029_,
		_w4031_
	);
	LUT2 #(
		.INIT('h1)
	) name3258 (
		_w4030_,
		_w4031_,
		_w4032_
	);
	LUT2 #(
		.INIT('h2)
	) name3259 (
		\g35_pad ,
		_w4032_,
		_w4033_
	);
	LUT2 #(
		.INIT('h2)
	) name3260 (
		\g3247_reg/NET0131 ,
		\g35_pad ,
		_w4034_
	);
	LUT2 #(
		.INIT('h1)
	) name3261 (
		_w4033_,
		_w4034_,
		_w4035_
	);
	LUT2 #(
		.INIT('h4)
	) name3262 (
		\g3171_reg/NET0131 ,
		\g3179_reg/NET0131 ,
		_w4036_
	);
	LUT2 #(
		.INIT('h8)
	) name3263 (
		_w4005_,
		_w4036_,
		_w4037_
	);
	LUT2 #(
		.INIT('h4)
	) name3264 (
		_w4008_,
		_w4037_,
		_w4038_
	);
	LUT2 #(
		.INIT('h2)
	) name3265 (
		\g3199_reg/NET0131 ,
		_w4037_,
		_w4039_
	);
	LUT2 #(
		.INIT('h1)
	) name3266 (
		_w4038_,
		_w4039_,
		_w4040_
	);
	LUT2 #(
		.INIT('h2)
	) name3267 (
		\g35_pad ,
		_w4040_,
		_w4041_
	);
	LUT2 #(
		.INIT('h2)
	) name3268 (
		\g3203_reg/NET0131 ,
		\g35_pad ,
		_w4042_
	);
	LUT2 #(
		.INIT('h1)
	) name3269 (
		_w4041_,
		_w4042_,
		_w4043_
	);
	LUT2 #(
		.INIT('h8)
	) name3270 (
		\g3167_reg/NET0131 ,
		_w4015_,
		_w4044_
	);
	LUT2 #(
		.INIT('h4)
	) name3271 (
		_w4008_,
		_w4044_,
		_w4045_
	);
	LUT2 #(
		.INIT('h2)
	) name3272 (
		\g3203_reg/NET0131 ,
		_w4044_,
		_w4046_
	);
	LUT2 #(
		.INIT('h1)
	) name3273 (
		_w4045_,
		_w4046_,
		_w4047_
	);
	LUT2 #(
		.INIT('h2)
	) name3274 (
		\g35_pad ,
		_w4047_,
		_w4048_
	);
	LUT2 #(
		.INIT('h2)
	) name3275 (
		\g3251_reg/NET0131 ,
		\g35_pad ,
		_w4049_
	);
	LUT2 #(
		.INIT('h1)
	) name3276 (
		_w4048_,
		_w4049_,
		_w4050_
	);
	LUT2 #(
		.INIT('h2)
	) name3277 (
		\g3155_reg/NET0131 ,
		\g3161_reg/NET0131 ,
		_w4051_
	);
	LUT2 #(
		.INIT('h8)
	) name3278 (
		_w4006_,
		_w4051_,
		_w4052_
	);
	LUT2 #(
		.INIT('h4)
	) name3279 (
		_w4008_,
		_w4052_,
		_w4053_
	);
	LUT2 #(
		.INIT('h2)
	) name3280 (
		\g3215_reg/NET0131 ,
		_w4052_,
		_w4054_
	);
	LUT2 #(
		.INIT('h1)
	) name3281 (
		_w4053_,
		_w4054_,
		_w4055_
	);
	LUT2 #(
		.INIT('h2)
	) name3282 (
		\g35_pad ,
		_w4055_,
		_w4056_
	);
	LUT2 #(
		.INIT('h2)
	) name3283 (
		\g3187_reg/NET0131 ,
		\g35_pad ,
		_w4057_
	);
	LUT2 #(
		.INIT('h1)
	) name3284 (
		_w4056_,
		_w4057_,
		_w4058_
	);
	LUT2 #(
		.INIT('h8)
	) name3285 (
		_w4015_,
		_w4051_,
		_w4059_
	);
	LUT2 #(
		.INIT('h4)
	) name3286 (
		_w4008_,
		_w4059_,
		_w4060_
	);
	LUT2 #(
		.INIT('h2)
	) name3287 (
		\g3219_reg/NET0131 ,
		_w4059_,
		_w4061_
	);
	LUT2 #(
		.INIT('h1)
	) name3288 (
		_w4060_,
		_w4061_,
		_w4062_
	);
	LUT2 #(
		.INIT('h2)
	) name3289 (
		\g35_pad ,
		_w4062_,
		_w4063_
	);
	LUT2 #(
		.INIT('h2)
	) name3290 (
		\g3191_reg/NET0131 ,
		\g35_pad ,
		_w4064_
	);
	LUT2 #(
		.INIT('h1)
	) name3291 (
		_w4063_,
		_w4064_,
		_w4065_
	);
	LUT2 #(
		.INIT('h8)
	) name3292 (
		_w4036_,
		_w4051_,
		_w4066_
	);
	LUT2 #(
		.INIT('h4)
	) name3293 (
		_w4008_,
		_w4066_,
		_w4067_
	);
	LUT2 #(
		.INIT('h2)
	) name3294 (
		\g3223_reg/NET0131 ,
		_w4066_,
		_w4068_
	);
	LUT2 #(
		.INIT('h1)
	) name3295 (
		_w4067_,
		_w4068_,
		_w4069_
	);
	LUT2 #(
		.INIT('h2)
	) name3296 (
		\g35_pad ,
		_w4069_,
		_w4070_
	);
	LUT2 #(
		.INIT('h2)
	) name3297 (
		\g3199_reg/NET0131 ,
		\g35_pad ,
		_w4071_
	);
	LUT2 #(
		.INIT('h1)
	) name3298 (
		_w4070_,
		_w4071_,
		_w4072_
	);
	LUT2 #(
		.INIT('h4)
	) name3299 (
		\g3155_reg/NET0131 ,
		\g3161_reg/NET0131 ,
		_w4073_
	);
	LUT2 #(
		.INIT('h8)
	) name3300 (
		_w4006_,
		_w4073_,
		_w4074_
	);
	LUT2 #(
		.INIT('h4)
	) name3301 (
		_w4008_,
		_w4074_,
		_w4075_
	);
	LUT2 #(
		.INIT('h2)
	) name3302 (
		\g3231_reg/NET0131 ,
		_w4074_,
		_w4076_
	);
	LUT2 #(
		.INIT('h1)
	) name3303 (
		_w4075_,
		_w4076_,
		_w4077_
	);
	LUT2 #(
		.INIT('h2)
	) name3304 (
		\g35_pad ,
		_w4077_,
		_w4078_
	);
	LUT2 #(
		.INIT('h2)
	) name3305 (
		\g3215_reg/NET0131 ,
		\g35_pad ,
		_w4079_
	);
	LUT2 #(
		.INIT('h1)
	) name3306 (
		_w4078_,
		_w4079_,
		_w4080_
	);
	LUT2 #(
		.INIT('h8)
	) name3307 (
		_w4015_,
		_w4073_,
		_w4081_
	);
	LUT2 #(
		.INIT('h4)
	) name3308 (
		_w4008_,
		_w4081_,
		_w4082_
	);
	LUT2 #(
		.INIT('h2)
	) name3309 (
		\g3235_reg/NET0131 ,
		_w4081_,
		_w4083_
	);
	LUT2 #(
		.INIT('h1)
	) name3310 (
		_w4082_,
		_w4083_,
		_w4084_
	);
	LUT2 #(
		.INIT('h2)
	) name3311 (
		\g35_pad ,
		_w4084_,
		_w4085_
	);
	LUT2 #(
		.INIT('h2)
	) name3312 (
		\g3219_reg/NET0131 ,
		\g35_pad ,
		_w4086_
	);
	LUT2 #(
		.INIT('h1)
	) name3313 (
		_w4085_,
		_w4086_,
		_w4087_
	);
	LUT2 #(
		.INIT('h8)
	) name3314 (
		_w4036_,
		_w4073_,
		_w4088_
	);
	LUT2 #(
		.INIT('h4)
	) name3315 (
		_w4008_,
		_w4088_,
		_w4089_
	);
	LUT2 #(
		.INIT('h2)
	) name3316 (
		\g3239_reg/NET0131 ,
		_w4088_,
		_w4090_
	);
	LUT2 #(
		.INIT('h1)
	) name3317 (
		_w4089_,
		_w4090_,
		_w4091_
	);
	LUT2 #(
		.INIT('h2)
	) name3318 (
		\g35_pad ,
		_w4091_,
		_w4092_
	);
	LUT2 #(
		.INIT('h2)
	) name3319 (
		\g3223_reg/NET0131 ,
		\g35_pad ,
		_w4093_
	);
	LUT2 #(
		.INIT('h1)
	) name3320 (
		_w4092_,
		_w4093_,
		_w4094_
	);
	LUT2 #(
		.INIT('h8)
	) name3321 (
		\g3155_reg/NET0131 ,
		\g3161_reg/NET0131 ,
		_w4095_
	);
	LUT2 #(
		.INIT('h8)
	) name3322 (
		_w4006_,
		_w4095_,
		_w4096_
	);
	LUT2 #(
		.INIT('h4)
	) name3323 (
		_w4008_,
		_w4096_,
		_w4097_
	);
	LUT2 #(
		.INIT('h2)
	) name3324 (
		\g3247_reg/NET0131 ,
		_w4096_,
		_w4098_
	);
	LUT2 #(
		.INIT('h1)
	) name3325 (
		_w4097_,
		_w4098_,
		_w4099_
	);
	LUT2 #(
		.INIT('h2)
	) name3326 (
		\g35_pad ,
		_w4099_,
		_w4100_
	);
	LUT2 #(
		.INIT('h2)
	) name3327 (
		\g3231_reg/NET0131 ,
		\g35_pad ,
		_w4101_
	);
	LUT2 #(
		.INIT('h1)
	) name3328 (
		_w4100_,
		_w4101_,
		_w4102_
	);
	LUT2 #(
		.INIT('h8)
	) name3329 (
		_w4015_,
		_w4095_,
		_w4103_
	);
	LUT2 #(
		.INIT('h4)
	) name3330 (
		_w4008_,
		_w4103_,
		_w4104_
	);
	LUT2 #(
		.INIT('h2)
	) name3331 (
		\g3251_reg/NET0131 ,
		_w4103_,
		_w4105_
	);
	LUT2 #(
		.INIT('h1)
	) name3332 (
		_w4104_,
		_w4105_,
		_w4106_
	);
	LUT2 #(
		.INIT('h2)
	) name3333 (
		\g35_pad ,
		_w4106_,
		_w4107_
	);
	LUT2 #(
		.INIT('h2)
	) name3334 (
		\g3235_reg/NET0131 ,
		\g35_pad ,
		_w4108_
	);
	LUT2 #(
		.INIT('h1)
	) name3335 (
		_w4107_,
		_w4108_,
		_w4109_
	);
	LUT2 #(
		.INIT('h8)
	) name3336 (
		\g3171_reg/NET0131 ,
		\g3179_reg/NET0131 ,
		_w4110_
	);
	LUT2 #(
		.INIT('h8)
	) name3337 (
		_w4005_,
		_w4110_,
		_w4111_
	);
	LUT2 #(
		.INIT('h4)
	) name3338 (
		_w4008_,
		_w4111_,
		_w4112_
	);
	LUT2 #(
		.INIT('h2)
	) name3339 (
		\g3207_reg/NET0131 ,
		_w4111_,
		_w4113_
	);
	LUT2 #(
		.INIT('h1)
	) name3340 (
		_w4112_,
		_w4113_,
		_w4114_
	);
	LUT2 #(
		.INIT('h2)
	) name3341 (
		\g35_pad ,
		_w4114_,
		_w4115_
	);
	LUT2 #(
		.INIT('h2)
	) name3342 (
		\g3211_reg/NET0131 ,
		\g35_pad ,
		_w4116_
	);
	LUT2 #(
		.INIT('h1)
	) name3343 (
		_w4115_,
		_w4116_,
		_w4117_
	);
	LUT2 #(
		.INIT('h8)
	) name3344 (
		\g3167_reg/NET0131 ,
		_w4036_,
		_w4118_
	);
	LUT2 #(
		.INIT('h4)
	) name3345 (
		_w4008_,
		_w4118_,
		_w4119_
	);
	LUT2 #(
		.INIT('h2)
	) name3346 (
		\g3211_reg/NET0131 ,
		_w4118_,
		_w4120_
	);
	LUT2 #(
		.INIT('h1)
	) name3347 (
		_w4119_,
		_w4120_,
		_w4121_
	);
	LUT2 #(
		.INIT('h2)
	) name3348 (
		\g35_pad ,
		_w4121_,
		_w4122_
	);
	LUT2 #(
		.INIT('h2)
	) name3349 (
		\g3255_reg/NET0131 ,
		\g35_pad ,
		_w4123_
	);
	LUT2 #(
		.INIT('h1)
	) name3350 (
		_w4122_,
		_w4123_,
		_w4124_
	);
	LUT2 #(
		.INIT('h8)
	) name3351 (
		_w4051_,
		_w4110_,
		_w4125_
	);
	LUT2 #(
		.INIT('h4)
	) name3352 (
		_w4008_,
		_w4125_,
		_w4126_
	);
	LUT2 #(
		.INIT('h2)
	) name3353 (
		\g3227_reg/NET0131 ,
		_w4125_,
		_w4127_
	);
	LUT2 #(
		.INIT('h1)
	) name3354 (
		_w4126_,
		_w4127_,
		_w4128_
	);
	LUT2 #(
		.INIT('h2)
	) name3355 (
		\g35_pad ,
		_w4128_,
		_w4129_
	);
	LUT2 #(
		.INIT('h2)
	) name3356 (
		\g3207_reg/NET0131 ,
		\g35_pad ,
		_w4130_
	);
	LUT2 #(
		.INIT('h1)
	) name3357 (
		_w4129_,
		_w4130_,
		_w4131_
	);
	LUT2 #(
		.INIT('h8)
	) name3358 (
		_w4073_,
		_w4110_,
		_w4132_
	);
	LUT2 #(
		.INIT('h4)
	) name3359 (
		_w4008_,
		_w4132_,
		_w4133_
	);
	LUT2 #(
		.INIT('h2)
	) name3360 (
		\g3243_reg/NET0131 ,
		_w4132_,
		_w4134_
	);
	LUT2 #(
		.INIT('h1)
	) name3361 (
		_w4133_,
		_w4134_,
		_w4135_
	);
	LUT2 #(
		.INIT('h2)
	) name3362 (
		\g35_pad ,
		_w4135_,
		_w4136_
	);
	LUT2 #(
		.INIT('h2)
	) name3363 (
		\g3227_reg/NET0131 ,
		\g35_pad ,
		_w4137_
	);
	LUT2 #(
		.INIT('h1)
	) name3364 (
		_w4136_,
		_w4137_,
		_w4138_
	);
	LUT2 #(
		.INIT('h8)
	) name3365 (
		_w4036_,
		_w4095_,
		_w4139_
	);
	LUT2 #(
		.INIT('h4)
	) name3366 (
		_w4008_,
		_w4139_,
		_w4140_
	);
	LUT2 #(
		.INIT('h2)
	) name3367 (
		\g3255_reg/NET0131 ,
		_w4139_,
		_w4141_
	);
	LUT2 #(
		.INIT('h1)
	) name3368 (
		_w4140_,
		_w4141_,
		_w4142_
	);
	LUT2 #(
		.INIT('h2)
	) name3369 (
		\g35_pad ,
		_w4142_,
		_w4143_
	);
	LUT2 #(
		.INIT('h2)
	) name3370 (
		\g3239_reg/NET0131 ,
		\g35_pad ,
		_w4144_
	);
	LUT2 #(
		.INIT('h1)
	) name3371 (
		_w4143_,
		_w4144_,
		_w4145_
	);
	LUT2 #(
		.INIT('h8)
	) name3372 (
		_w4095_,
		_w4110_,
		_w4146_
	);
	LUT2 #(
		.INIT('h4)
	) name3373 (
		_w4008_,
		_w4146_,
		_w4147_
	);
	LUT2 #(
		.INIT('h2)
	) name3374 (
		\g3259_reg/NET0131 ,
		_w4146_,
		_w4148_
	);
	LUT2 #(
		.INIT('h1)
	) name3375 (
		_w4147_,
		_w4148_,
		_w4149_
	);
	LUT2 #(
		.INIT('h2)
	) name3376 (
		\g35_pad ,
		_w4149_,
		_w4150_
	);
	LUT2 #(
		.INIT('h2)
	) name3377 (
		\g3243_reg/NET0131 ,
		\g35_pad ,
		_w4151_
	);
	LUT2 #(
		.INIT('h1)
	) name3378 (
		_w4150_,
		_w4151_,
		_w4152_
	);
	LUT2 #(
		.INIT('h8)
	) name3379 (
		\g3167_reg/NET0131 ,
		_w4110_,
		_w4153_
	);
	LUT2 #(
		.INIT('h4)
	) name3380 (
		_w4008_,
		_w4153_,
		_w4154_
	);
	LUT2 #(
		.INIT('h2)
	) name3381 (
		\g3263_reg/NET0131 ,
		_w4153_,
		_w4155_
	);
	LUT2 #(
		.INIT('h1)
	) name3382 (
		_w4154_,
		_w4155_,
		_w4156_
	);
	LUT2 #(
		.INIT('h2)
	) name3383 (
		\g35_pad ,
		_w4156_,
		_w4157_
	);
	LUT2 #(
		.INIT('h2)
	) name3384 (
		\g3259_reg/NET0131 ,
		\g35_pad ,
		_w4158_
	);
	LUT2 #(
		.INIT('h1)
	) name3385 (
		_w4157_,
		_w4158_,
		_w4159_
	);
	LUT2 #(
		.INIT('h8)
	) name3386 (
		\g1906_reg/NET0131 ,
		_w1516_,
		_w4160_
	);
	LUT2 #(
		.INIT('h1)
	) name3387 (
		_w1878_,
		_w4160_,
		_w4161_
	);
	LUT2 #(
		.INIT('h2)
	) name3388 (
		\g35_pad ,
		_w4161_,
		_w4162_
	);
	LUT2 #(
		.INIT('h2)
	) name3389 (
		\g1913_reg/NET0131 ,
		\g35_pad ,
		_w4163_
	);
	LUT2 #(
		.INIT('h1)
	) name3390 (
		_w4162_,
		_w4163_,
		_w4164_
	);
	LUT2 #(
		.INIT('h2)
	) name3391 (
		\g1906_reg/NET0131 ,
		_w1517_,
		_w4165_
	);
	LUT2 #(
		.INIT('h8)
	) name3392 (
		\g1936_reg/NET0131 ,
		_w1517_,
		_w4166_
	);
	LUT2 #(
		.INIT('h1)
	) name3393 (
		_w4165_,
		_w4166_,
		_w4167_
	);
	LUT2 #(
		.INIT('h2)
	) name3394 (
		\g35_pad ,
		_w2108_,
		_w4168_
	);
	LUT2 #(
		.INIT('h8)
	) name3395 (
		\g5084_reg/NET0131 ,
		\g5092_reg/NET0131 ,
		_w4169_
	);
	LUT2 #(
		.INIT('h2)
	) name3396 (
		\g35_pad ,
		_w4169_,
		_w4170_
	);
	LUT2 #(
		.INIT('h2)
	) name3397 (
		\g5097_reg/NET0131 ,
		_w4170_,
		_w4171_
	);
	LUT2 #(
		.INIT('h8)
	) name3398 (
		\g29213_pad ,
		\g35_pad ,
		_w4172_
	);
	LUT2 #(
		.INIT('h4)
	) name3399 (
		_w4171_,
		_w4172_,
		_w4173_
	);
	LUT2 #(
		.INIT('h2)
	) name3400 (
		_w4171_,
		_w4172_,
		_w4174_
	);
	LUT2 #(
		.INIT('h1)
	) name3401 (
		_w4173_,
		_w4174_,
		_w4175_
	);
	LUT2 #(
		.INIT('h8)
	) name3402 (
		\g3639_reg/NET0131 ,
		\g3703_reg/NET0131 ,
		_w4176_
	);
	LUT2 #(
		.INIT('h8)
	) name3403 (
		_w894_,
		_w4176_,
		_w4177_
	);
	LUT2 #(
		.INIT('h8)
	) name3404 (
		_w2243_,
		_w4177_,
		_w4178_
	);
	LUT2 #(
		.INIT('h8)
	) name3405 (
		\g3470_reg/NET0131 ,
		_w4178_,
		_w4179_
	);
	LUT2 #(
		.INIT('h2)
	) name3406 (
		\g35_pad ,
		_w4179_,
		_w4180_
	);
	LUT2 #(
		.INIT('h1)
	) name3407 (
		\g3476_reg/NET0131 ,
		_w4180_,
		_w4181_
	);
	LUT2 #(
		.INIT('h1)
	) name3408 (
		\g3480_reg/NET0131 ,
		_w4178_,
		_w4182_
	);
	LUT2 #(
		.INIT('h4)
	) name3409 (
		\g3470_reg/NET0131 ,
		\g3476_reg/NET0131 ,
		_w4183_
	);
	LUT2 #(
		.INIT('h8)
	) name3410 (
		_w4178_,
		_w4183_,
		_w4184_
	);
	LUT2 #(
		.INIT('h1)
	) name3411 (
		_w4182_,
		_w4184_,
		_w4185_
	);
	LUT2 #(
		.INIT('h2)
	) name3412 (
		\g35_pad ,
		_w4185_,
		_w4186_
	);
	LUT2 #(
		.INIT('h1)
	) name3413 (
		_w4181_,
		_w4186_,
		_w4187_
	);
	LUT2 #(
		.INIT('h2)
	) name3414 (
		\g3484_reg/NET0131 ,
		_w4178_,
		_w4188_
	);
	LUT2 #(
		.INIT('h4)
	) name3415 (
		\g3484_reg/NET0131 ,
		_w4178_,
		_w4189_
	);
	LUT2 #(
		.INIT('h1)
	) name3416 (
		_w4188_,
		_w4189_,
		_w4190_
	);
	LUT2 #(
		.INIT('h2)
	) name3417 (
		\g35_pad ,
		_w4190_,
		_w4191_
	);
	LUT2 #(
		.INIT('h2)
	) name3418 (
		\g3480_reg/NET0131 ,
		\g35_pad ,
		_w4192_
	);
	LUT2 #(
		.INIT('h1)
	) name3419 (
		_w4191_,
		_w4192_,
		_w4193_
	);
	LUT2 #(
		.INIT('h8)
	) name3420 (
		\g2040_reg/NET0131 ,
		_w1533_,
		_w4194_
	);
	LUT2 #(
		.INIT('h1)
	) name3421 (
		_w1901_,
		_w4194_,
		_w4195_
	);
	LUT2 #(
		.INIT('h2)
	) name3422 (
		\g35_pad ,
		_w4195_,
		_w4196_
	);
	LUT2 #(
		.INIT('h2)
	) name3423 (
		\g2047_reg/NET0131 ,
		\g35_pad ,
		_w4197_
	);
	LUT2 #(
		.INIT('h1)
	) name3424 (
		_w4196_,
		_w4197_,
		_w4198_
	);
	LUT2 #(
		.INIT('h8)
	) name3425 (
		\g4054_reg/NET0131 ,
		_w890_,
		_w4199_
	);
	LUT2 #(
		.INIT('h8)
	) name3426 (
		_w895_,
		_w4199_,
		_w4200_
	);
	LUT2 #(
		.INIT('h2)
	) name3427 (
		\g35_pad ,
		_w4200_,
		_w4201_
	);
	LUT2 #(
		.INIT('h8)
	) name3428 (
		\g3821_reg/NET0131 ,
		_w4200_,
		_w4202_
	);
	LUT2 #(
		.INIT('h2)
	) name3429 (
		\g35_pad ,
		_w4202_,
		_w4203_
	);
	LUT2 #(
		.INIT('h1)
	) name3430 (
		\g3827_reg/NET0131 ,
		_w4203_,
		_w4204_
	);
	LUT2 #(
		.INIT('h1)
	) name3431 (
		\g3831_reg/NET0131 ,
		_w4200_,
		_w4205_
	);
	LUT2 #(
		.INIT('h4)
	) name3432 (
		\g3821_reg/NET0131 ,
		\g3827_reg/NET0131 ,
		_w4206_
	);
	LUT2 #(
		.INIT('h8)
	) name3433 (
		_w4200_,
		_w4206_,
		_w4207_
	);
	LUT2 #(
		.INIT('h1)
	) name3434 (
		_w4205_,
		_w4207_,
		_w4208_
	);
	LUT2 #(
		.INIT('h2)
	) name3435 (
		\g35_pad ,
		_w4208_,
		_w4209_
	);
	LUT2 #(
		.INIT('h1)
	) name3436 (
		_w4204_,
		_w4209_,
		_w4210_
	);
	LUT2 #(
		.INIT('h2)
	) name3437 (
		\g3835_reg/NET0131 ,
		_w4200_,
		_w4211_
	);
	LUT2 #(
		.INIT('h4)
	) name3438 (
		\g3835_reg/NET0131 ,
		_w4200_,
		_w4212_
	);
	LUT2 #(
		.INIT('h1)
	) name3439 (
		_w4211_,
		_w4212_,
		_w4213_
	);
	LUT2 #(
		.INIT('h2)
	) name3440 (
		\g35_pad ,
		_w4213_,
		_w4214_
	);
	LUT2 #(
		.INIT('h4)
	) name3441 (
		\g35_pad ,
		\g3831_reg/NET0131 ,
		_w4215_
	);
	LUT2 #(
		.INIT('h1)
	) name3442 (
		_w4214_,
		_w4215_,
		_w4216_
	);
	LUT2 #(
		.INIT('h8)
	) name3443 (
		\g2197_reg/NET0131 ,
		_w1398_,
		_w4217_
	);
	LUT2 #(
		.INIT('h1)
	) name3444 (
		_w1583_,
		_w4217_,
		_w4218_
	);
	LUT2 #(
		.INIT('h2)
	) name3445 (
		\g35_pad ,
		_w4218_,
		_w4219_
	);
	LUT2 #(
		.INIT('h2)
	) name3446 (
		\g2204_reg/NET0131 ,
		\g35_pad ,
		_w4220_
	);
	LUT2 #(
		.INIT('h1)
	) name3447 (
		_w4219_,
		_w4220_,
		_w4221_
	);
	LUT2 #(
		.INIT('h2)
	) name3448 (
		\g2197_reg/NET0131 ,
		_w1399_,
		_w4222_
	);
	LUT2 #(
		.INIT('h8)
	) name3449 (
		\g2227_reg/NET0131 ,
		_w1399_,
		_w4223_
	);
	LUT2 #(
		.INIT('h1)
	) name3450 (
		_w4222_,
		_w4223_,
		_w4224_
	);
	LUT2 #(
		.INIT('h8)
	) name3451 (
		\g4258_reg/NET0131 ,
		\g4264_reg/NET0131 ,
		_w4225_
	);
	LUT2 #(
		.INIT('h2)
	) name3452 (
		\g35_pad ,
		_w4225_,
		_w4226_
	);
	LUT2 #(
		.INIT('h2)
	) name3453 (
		\g4269_reg/NET0131 ,
		_w4226_,
		_w4227_
	);
	LUT2 #(
		.INIT('h8)
	) name3454 (
		\g35_pad ,
		\g4273_reg/NET0131 ,
		_w4228_
	);
	LUT2 #(
		.INIT('h4)
	) name3455 (
		_w4227_,
		_w4228_,
		_w4229_
	);
	LUT2 #(
		.INIT('h2)
	) name3456 (
		_w4227_,
		_w4228_,
		_w4230_
	);
	LUT2 #(
		.INIT('h1)
	) name3457 (
		_w4229_,
		_w4230_,
		_w4231_
	);
	LUT2 #(
		.INIT('h4)
	) name3458 (
		\g35_pad ,
		\g4340_reg/NET0131 ,
		_w4232_
	);
	LUT2 #(
		.INIT('h1)
	) name3459 (
		\g4349_reg/NET0131 ,
		_w3606_,
		_w4233_
	);
	LUT2 #(
		.INIT('h2)
	) name3460 (
		\g35_pad ,
		_w3604_,
		_w4234_
	);
	LUT2 #(
		.INIT('h4)
	) name3461 (
		_w4233_,
		_w4234_,
		_w4235_
	);
	LUT2 #(
		.INIT('h1)
	) name3462 (
		_w4232_,
		_w4235_,
		_w4236_
	);
	LUT2 #(
		.INIT('h8)
	) name3463 (
		\g2331_reg/NET0131 ,
		_w1415_,
		_w4237_
	);
	LUT2 #(
		.INIT('h1)
	) name3464 (
		_w1629_,
		_w4237_,
		_w4238_
	);
	LUT2 #(
		.INIT('h2)
	) name3465 (
		\g35_pad ,
		_w4238_,
		_w4239_
	);
	LUT2 #(
		.INIT('h2)
	) name3466 (
		\g2338_reg/NET0131 ,
		\g35_pad ,
		_w4240_
	);
	LUT2 #(
		.INIT('h1)
	) name3467 (
		_w4239_,
		_w4240_,
		_w4241_
	);
	LUT2 #(
		.INIT('h2)
	) name3468 (
		\g2331_reg/NET0131 ,
		_w1416_,
		_w4242_
	);
	LUT2 #(
		.INIT('h8)
	) name3469 (
		\g2361_reg/NET0131 ,
		_w1416_,
		_w4243_
	);
	LUT2 #(
		.INIT('h1)
	) name3470 (
		_w4242_,
		_w4243_,
		_w4244_
	);
	LUT2 #(
		.INIT('h2)
	) name3471 (
		\g239_reg/NET0131 ,
		_w3427_,
		_w4245_
	);
	LUT2 #(
		.INIT('h8)
	) name3472 (
		\g14125_pad ,
		_w3427_,
		_w4246_
	);
	LUT2 #(
		.INIT('h1)
	) name3473 (
		_w4245_,
		_w4246_,
		_w4247_
	);
	LUT2 #(
		.INIT('h2)
	) name3474 (
		\g35_pad ,
		_w4247_,
		_w4248_
	);
	LUT2 #(
		.INIT('h2)
	) name3475 (
		\g262_reg/NET0131 ,
		\g35_pad ,
		_w4249_
	);
	LUT2 #(
		.INIT('h1)
	) name3476 (
		_w4248_,
		_w4249_,
		_w4250_
	);
	LUT2 #(
		.INIT('h2)
	) name3477 (
		\g35_pad ,
		_w4178_,
		_w4251_
	);
	LUT2 #(
		.INIT('h8)
	) name3478 (
		\g2465_reg/NET0131 ,
		_w1432_,
		_w4252_
	);
	LUT2 #(
		.INIT('h1)
	) name3479 (
		_w1680_,
		_w4252_,
		_w4253_
	);
	LUT2 #(
		.INIT('h2)
	) name3480 (
		\g35_pad ,
		_w4253_,
		_w4254_
	);
	LUT2 #(
		.INIT('h2)
	) name3481 (
		\g2472_reg/NET0131 ,
		\g35_pad ,
		_w4255_
	);
	LUT2 #(
		.INIT('h1)
	) name3482 (
		_w4254_,
		_w4255_,
		_w4256_
	);
	LUT2 #(
		.INIT('h2)
	) name3483 (
		\g2465_reg/NET0131 ,
		_w1433_,
		_w4257_
	);
	LUT2 #(
		.INIT('h8)
	) name3484 (
		\g2495_reg/NET0131 ,
		_w1433_,
		_w4258_
	);
	LUT2 #(
		.INIT('h1)
	) name3485 (
		_w4257_,
		_w4258_,
		_w4259_
	);
	LUT2 #(
		.INIT('h1)
	) name3486 (
		\g35_pad ,
		\g528_reg/NET0131 ,
		_w4260_
	);
	LUT2 #(
		.INIT('h1)
	) name3487 (
		\g482_reg/NET0131 ,
		_w3374_,
		_w4261_
	);
	LUT2 #(
		.INIT('h1)
	) name3488 (
		_w3381_,
		_w4261_,
		_w4262_
	);
	LUT2 #(
		.INIT('h2)
	) name3489 (
		\g35_pad ,
		_w3375_,
		_w4263_
	);
	LUT2 #(
		.INIT('h4)
	) name3490 (
		_w4262_,
		_w4263_,
		_w4264_
	);
	LUT2 #(
		.INIT('h1)
	) name3491 (
		_w4260_,
		_w4264_,
		_w4265_
	);
	LUT2 #(
		.INIT('h8)
	) name3492 (
		\g1636_reg/NET0131 ,
		_w1950_,
		_w4266_
	);
	LUT2 #(
		.INIT('h1)
	) name3493 (
		_w1951_,
		_w4266_,
		_w4267_
	);
	LUT2 #(
		.INIT('h2)
	) name3494 (
		\g35_pad ,
		_w4267_,
		_w4268_
	);
	LUT2 #(
		.INIT('h2)
	) name3495 (
		\g1644_reg/NET0131 ,
		\g35_pad ,
		_w4269_
	);
	LUT2 #(
		.INIT('h1)
	) name3496 (
		_w4268_,
		_w4269_,
		_w4270_
	);
	LUT2 #(
		.INIT('h1)
	) name3497 (
		\g2555_reg/NET0131 ,
		_w1449_,
		_w4271_
	);
	LUT2 #(
		.INIT('h4)
	) name3498 (
		\g2599_reg/NET0131 ,
		_w1449_,
		_w4272_
	);
	LUT2 #(
		.INIT('h1)
	) name3499 (
		_w4271_,
		_w4272_,
		_w4273_
	);
	LUT2 #(
		.INIT('h2)
	) name3500 (
		\g35_pad ,
		_w4273_,
		_w4274_
	);
	LUT2 #(
		.INIT('h1)
	) name3501 (
		\g2606_reg/NET0131 ,
		\g35_pad ,
		_w4275_
	);
	LUT2 #(
		.INIT('h1)
	) name3502 (
		_w4274_,
		_w4275_,
		_w4276_
	);
	LUT2 #(
		.INIT('h8)
	) name3503 (
		\g35_pad ,
		_w1950_,
		_w4277_
	);
	LUT2 #(
		.INIT('h2)
	) name3504 (
		\g1636_reg/NET0131 ,
		_w4277_,
		_w4278_
	);
	LUT2 #(
		.INIT('h8)
	) name3505 (
		\g1668_reg/NET0131 ,
		_w4277_,
		_w4279_
	);
	LUT2 #(
		.INIT('h1)
	) name3506 (
		_w4278_,
		_w4279_,
		_w4280_
	);
	LUT2 #(
		.INIT('h8)
	) name3507 (
		\g3111_reg/NET0131 ,
		\g35_pad ,
		_w4281_
	);
	LUT2 #(
		.INIT('h1)
	) name3508 (
		\g5115_reg/NET0131 ,
		_w4281_,
		_w4282_
	);
	LUT2 #(
		.INIT('h8)
	) name3509 (
		\g5115_reg/NET0131 ,
		_w4281_,
		_w4283_
	);
	LUT2 #(
		.INIT('h1)
	) name3510 (
		_w4282_,
		_w4283_,
		_w4284_
	);
	LUT2 #(
		.INIT('h1)
	) name3511 (
		_w3967_,
		_w4284_,
		_w4285_
	);
	LUT2 #(
		.INIT('h4)
	) name3512 (
		\g5124_reg/NET0131 ,
		_w3967_,
		_w4286_
	);
	LUT2 #(
		.INIT('h1)
	) name3513 (
		_w4285_,
		_w4286_,
		_w4287_
	);
	LUT2 #(
		.INIT('h1)
	) name3514 (
		\g3106_reg/NET0131 ,
		_w4281_,
		_w4288_
	);
	LUT2 #(
		.INIT('h8)
	) name3515 (
		\g3106_reg/NET0131 ,
		_w4281_,
		_w4289_
	);
	LUT2 #(
		.INIT('h1)
	) name3516 (
		_w4288_,
		_w4289_,
		_w4290_
	);
	LUT2 #(
		.INIT('h1)
	) name3517 (
		_w3994_,
		_w4290_,
		_w4291_
	);
	LUT2 #(
		.INIT('h4)
	) name3518 (
		\g3115_reg/NET0131 ,
		_w3994_,
		_w4292_
	);
	LUT2 #(
		.INIT('h1)
	) name3519 (
		_w4291_,
		_w4292_,
		_w4293_
	);
	LUT2 #(
		.INIT('h4)
	) name3520 (
		\g311_reg/NET0131 ,
		\g324_reg/NET0131 ,
		_w4294_
	);
	LUT2 #(
		.INIT('h1)
	) name3521 (
		\g305_reg/NET0131 ,
		_w4294_,
		_w4295_
	);
	LUT2 #(
		.INIT('h2)
	) name3522 (
		\g35_pad ,
		_w4295_,
		_w4296_
	);
	LUT2 #(
		.INIT('h2)
	) name3523 (
		\g336_reg/NET0131 ,
		\g35_pad ,
		_w4297_
	);
	LUT2 #(
		.INIT('h1)
	) name3524 (
		_w4296_,
		_w4297_,
		_w4298_
	);
	LUT2 #(
		.INIT('h4)
	) name3525 (
		\g661_reg/NET0131 ,
		_w2464_,
		_w4299_
	);
	LUT2 #(
		.INIT('h2)
	) name3526 (
		\g35_pad ,
		_w4299_,
		_w4300_
	);
	LUT2 #(
		.INIT('h1)
	) name3527 (
		\g728_reg/NET0131 ,
		_w4300_,
		_w4301_
	);
	LUT2 #(
		.INIT('h4)
	) name3528 (
		\g29212_pad ,
		\g35_pad ,
		_w4302_
	);
	LUT2 #(
		.INIT('h4)
	) name3529 (
		_w2464_,
		_w4302_,
		_w4303_
	);
	LUT2 #(
		.INIT('h1)
	) name3530 (
		_w4301_,
		_w4303_,
		_w4304_
	);
	LUT2 #(
		.INIT('h1)
	) name3531 (
		\g3457_reg/NET0131 ,
		_w4281_,
		_w4305_
	);
	LUT2 #(
		.INIT('h8)
	) name3532 (
		\g3457_reg/NET0131 ,
		_w4281_,
		_w4306_
	);
	LUT2 #(
		.INIT('h1)
	) name3533 (
		_w4305_,
		_w4306_,
		_w4307_
	);
	LUT2 #(
		.INIT('h1)
	) name3534 (
		_w4251_,
		_w4307_,
		_w4308_
	);
	LUT2 #(
		.INIT('h4)
	) name3535 (
		\g3466_reg/NET0131 ,
		_w4251_,
		_w4309_
	);
	LUT2 #(
		.INIT('h1)
	) name3536 (
		_w4308_,
		_w4309_,
		_w4310_
	);
	LUT2 #(
		.INIT('h1)
	) name3537 (
		\g3808_reg/NET0131 ,
		_w4281_,
		_w4311_
	);
	LUT2 #(
		.INIT('h8)
	) name3538 (
		\g3808_reg/NET0131 ,
		_w4281_,
		_w4312_
	);
	LUT2 #(
		.INIT('h1)
	) name3539 (
		_w4311_,
		_w4312_,
		_w4313_
	);
	LUT2 #(
		.INIT('h1)
	) name3540 (
		_w4201_,
		_w4313_,
		_w4314_
	);
	LUT2 #(
		.INIT('h4)
	) name3541 (
		\g3817_reg/NET0131 ,
		_w4201_,
		_w4315_
	);
	LUT2 #(
		.INIT('h1)
	) name3542 (
		_w4314_,
		_w4315_,
		_w4316_
	);
	LUT2 #(
		.INIT('h4)
	) name3543 (
		\g35_pad ,
		\g5041_reg/NET0131 ,
		_w4317_
	);
	LUT2 #(
		.INIT('h1)
	) name3544 (
		_w3497_,
		_w3503_,
		_w4318_
	);
	LUT2 #(
		.INIT('h8)
	) name3545 (
		\g5046_reg/NET0131 ,
		_w3572_,
		_w4319_
	);
	LUT2 #(
		.INIT('h8)
	) name3546 (
		_w4318_,
		_w4319_,
		_w4320_
	);
	LUT2 #(
		.INIT('h2)
	) name3547 (
		\g35_pad ,
		\g5046_reg/NET0131 ,
		_w4321_
	);
	LUT2 #(
		.INIT('h4)
	) name3548 (
		_w4318_,
		_w4321_,
		_w4322_
	);
	LUT2 #(
		.INIT('h1)
	) name3549 (
		_w4317_,
		_w4320_,
		_w4323_
	);
	LUT2 #(
		.INIT('h4)
	) name3550 (
		_w4322_,
		_w4323_,
		_w4324_
	);
	LUT2 #(
		.INIT('h2)
	) name3551 (
		\g35_pad ,
		\g5069_reg/NET0131 ,
		_w4325_
	);
	LUT2 #(
		.INIT('h2)
	) name3552 (
		\g5073_reg/NET0131 ,
		_w4325_,
		_w4326_
	);
	LUT2 #(
		.INIT('h2)
	) name3553 (
		\g3147_reg/NET0131 ,
		_w4153_,
		_w4327_
	);
	LUT2 #(
		.INIT('h2)
	) name3554 (
		_w4008_,
		_w4327_,
		_w4328_
	);
	LUT2 #(
		.INIT('h4)
	) name3555 (
		_w4008_,
		_w4327_,
		_w4329_
	);
	LUT2 #(
		.INIT('h2)
	) name3556 (
		\g35_pad ,
		_w4328_,
		_w4330_
	);
	LUT2 #(
		.INIT('h4)
	) name3557 (
		_w4329_,
		_w4330_,
		_w4331_
	);
	LUT2 #(
		.INIT('h2)
	) name3558 (
		\g35_pad ,
		_w2377_,
		_w4332_
	);
	LUT2 #(
		.INIT('h2)
	) name3559 (
		\g969_reg/NET0131 ,
		_w4332_,
		_w4333_
	);
	LUT2 #(
		.INIT('h1)
	) name3560 (
		_w3295_,
		_w3846_,
		_w4334_
	);
	LUT2 #(
		.INIT('h1)
	) name3561 (
		_w2373_,
		_w4334_,
		_w4335_
	);
	LUT2 #(
		.INIT('h8)
	) name3562 (
		\g1008_reg/NET0131 ,
		\g35_pad ,
		_w4336_
	);
	LUT2 #(
		.INIT('h4)
	) name3563 (
		_w4335_,
		_w4336_,
		_w4337_
	);
	LUT2 #(
		.INIT('h1)
	) name3564 (
		_w4333_,
		_w4337_,
		_w4338_
	);
	LUT2 #(
		.INIT('h8)
	) name3565 (
		\g5357_reg/NET0131 ,
		_w869_,
		_w4339_
	);
	LUT2 #(
		.INIT('h2)
	) name3566 (
		\g35_pad ,
		_w4339_,
		_w4340_
	);
	LUT2 #(
		.INIT('h8)
	) name3567 (
		\g5297_reg/NET0131 ,
		_w4340_,
		_w4341_
	);
	LUT2 #(
		.INIT('h8)
	) name3568 (
		\g35_pad ,
		\g5297_reg/NET0131 ,
		_w4342_
	);
	LUT2 #(
		.INIT('h2)
	) name3569 (
		\g5357_reg/NET0131 ,
		_w4342_,
		_w4343_
	);
	LUT2 #(
		.INIT('h4)
	) name3570 (
		_w2587_,
		_w4343_,
		_w4344_
	);
	LUT2 #(
		.INIT('h1)
	) name3571 (
		_w4341_,
		_w4344_,
		_w4345_
	);
	LUT2 #(
		.INIT('h2)
	) name3572 (
		\g3352_reg/NET0131 ,
		_w2328_,
		_w4346_
	);
	LUT2 #(
		.INIT('h8)
	) name3573 (
		\g3288_reg/NET0131 ,
		\g35_pad ,
		_w4347_
	);
	LUT2 #(
		.INIT('h4)
	) name3574 (
		_w4346_,
		_w4347_,
		_w4348_
	);
	LUT2 #(
		.INIT('h2)
	) name3575 (
		_w4346_,
		_w4347_,
		_w4349_
	);
	LUT2 #(
		.INIT('h1)
	) name3576 (
		_w4348_,
		_w4349_,
		_w4350_
	);
	LUT2 #(
		.INIT('h8)
	) name3577 (
		\g3703_reg/NET0131 ,
		_w2243_,
		_w4351_
	);
	LUT2 #(
		.INIT('h2)
	) name3578 (
		\g35_pad ,
		_w4351_,
		_w4352_
	);
	LUT2 #(
		.INIT('h8)
	) name3579 (
		\g3639_reg/NET0131 ,
		_w4352_,
		_w4353_
	);
	LUT2 #(
		.INIT('h8)
	) name3580 (
		\g35_pad ,
		\g3639_reg/NET0131 ,
		_w4354_
	);
	LUT2 #(
		.INIT('h2)
	) name3581 (
		\g3703_reg/NET0131 ,
		_w4354_,
		_w4355_
	);
	LUT2 #(
		.INIT('h4)
	) name3582 (
		_w2445_,
		_w4355_,
		_w4356_
	);
	LUT2 #(
		.INIT('h1)
	) name3583 (
		_w4353_,
		_w4356_,
		_w4357_
	);
	LUT2 #(
		.INIT('h2)
	) name3584 (
		\g35_pad ,
		_w4199_,
		_w4358_
	);
	LUT2 #(
		.INIT('h8)
	) name3585 (
		\g3990_reg/NET0131 ,
		_w4358_,
		_w4359_
	);
	LUT2 #(
		.INIT('h8)
	) name3586 (
		\g35_pad ,
		\g3990_reg/NET0131 ,
		_w4360_
	);
	LUT2 #(
		.INIT('h2)
	) name3587 (
		\g4054_reg/NET0131 ,
		_w4360_,
		_w4361_
	);
	LUT2 #(
		.INIT('h4)
	) name3588 (
		_w891_,
		_w4361_,
		_w4362_
	);
	LUT2 #(
		.INIT('h1)
	) name3589 (
		_w4359_,
		_w4362_,
		_w4363_
	);
	LUT2 #(
		.INIT('h2)
	) name3590 (
		\g3338_reg/NET0131 ,
		\g35_pad ,
		_w4364_
	);
	LUT2 #(
		.INIT('h4)
	) name3591 (
		\g3347_reg/NET0131 ,
		_w3934_,
		_w4365_
	);
	LUT2 #(
		.INIT('h1)
	) name3592 (
		_w4364_,
		_w4365_,
		_w4366_
	);
	LUT2 #(
		.INIT('h4)
	) name3593 (
		\g35_pad ,
		\g812_reg/NET0131 ,
		_w4367_
	);
	LUT2 #(
		.INIT('h1)
	) name3594 (
		\g817_reg/NET0131 ,
		_w2206_,
		_w4368_
	);
	LUT2 #(
		.INIT('h4)
	) name3595 (
		_w2207_,
		_w2213_,
		_w4369_
	);
	LUT2 #(
		.INIT('h4)
	) name3596 (
		_w4368_,
		_w4369_,
		_w4370_
	);
	LUT2 #(
		.INIT('h1)
	) name3597 (
		_w4367_,
		_w4370_,
		_w4371_
	);
	LUT2 #(
		.INIT('h1)
	) name3598 (
		\g2864_reg/NET0131 ,
		\g35_pad ,
		_w4372_
	);
	LUT2 #(
		.INIT('h4)
	) name3599 (
		\g2898_reg/NET0131 ,
		\g35_pad ,
		_w4373_
	);
	LUT2 #(
		.INIT('h8)
	) name3600 (
		_w1016_,
		_w4373_,
		_w4374_
	);
	LUT2 #(
		.INIT('h1)
	) name3601 (
		_w4372_,
		_w4374_,
		_w4375_
	);
	LUT2 #(
		.INIT('h1)
	) name3602 (
		\g35_pad ,
		\g4172_reg/NET0131 ,
		_w4376_
	);
	LUT2 #(
		.INIT('h4)
	) name3603 (
		\g4176_reg/NET0131 ,
		_w3923_,
		_w4377_
	);
	LUT2 #(
		.INIT('h1)
	) name3604 (
		_w4376_,
		_w4377_,
		_w4378_
	);
	LUT2 #(
		.INIT('h1)
	) name3605 (
		_w3494_,
		_w3500_,
		_w4379_
	);
	LUT2 #(
		.INIT('h1)
	) name3606 (
		\g5033_reg/NET0131 ,
		_w4379_,
		_w4380_
	);
	LUT2 #(
		.INIT('h8)
	) name3607 (
		\g5033_reg/NET0131 ,
		_w3953_,
		_w4381_
	);
	LUT2 #(
		.INIT('h8)
	) name3608 (
		_w4379_,
		_w4381_,
		_w4382_
	);
	LUT2 #(
		.INIT('h1)
	) name3609 (
		_w4380_,
		_w4382_,
		_w4383_
	);
	LUT2 #(
		.INIT('h2)
	) name3610 (
		\g35_pad ,
		_w4383_,
		_w4384_
	);
	LUT2 #(
		.INIT('h4)
	) name3611 (
		\g35_pad ,
		\g5029_reg/NET0131 ,
		_w4385_
	);
	LUT2 #(
		.INIT('h1)
	) name3612 (
		_w4384_,
		_w4385_,
		_w4386_
	);
	LUT2 #(
		.INIT('h2)
	) name3613 (
		\g3347_reg/NET0131 ,
		\g35_pad ,
		_w4387_
	);
	LUT2 #(
		.INIT('h1)
	) name3614 (
		\g5357_reg/NET0131 ,
		_w869_,
		_w4388_
	);
	LUT2 #(
		.INIT('h2)
	) name3615 (
		_w4340_,
		_w4388_,
		_w4389_
	);
	LUT2 #(
		.INIT('h1)
	) name3616 (
		_w4387_,
		_w4389_,
		_w4390_
	);
	LUT2 #(
		.INIT('h8)
	) name3617 (
		\g691_reg/NET0131 ,
		_w982_,
		_w4391_
	);
	LUT2 #(
		.INIT('h4)
	) name3618 (
		\g411_reg/NET0131 ,
		\g417_reg/NET0131 ,
		_w4392_
	);
	LUT2 #(
		.INIT('h1)
	) name3619 (
		\g424_reg/NET0131 ,
		\g691_reg/NET0131 ,
		_w4393_
	);
	LUT2 #(
		.INIT('h8)
	) name3620 (
		_w4392_,
		_w4393_,
		_w4394_
	);
	LUT2 #(
		.INIT('h1)
	) name3621 (
		_w4391_,
		_w4394_,
		_w4395_
	);
	LUT2 #(
		.INIT('h2)
	) name3622 (
		_w2107_,
		_w4395_,
		_w4396_
	);
	LUT2 #(
		.INIT('h2)
	) name3623 (
		\g650_reg/NET0131 ,
		_w4396_,
		_w4397_
	);
	LUT2 #(
		.INIT('h8)
	) name3624 (
		\g681_reg/NET0131 ,
		_w4396_,
		_w4398_
	);
	LUT2 #(
		.INIT('h1)
	) name3625 (
		_w4397_,
		_w4398_,
		_w4399_
	);
	LUT2 #(
		.INIT('h2)
	) name3626 (
		\g35_pad ,
		_w4399_,
		_w4400_
	);
	LUT2 #(
		.INIT('h4)
	) name3627 (
		\g35_pad ,
		\g699_reg/NET0131 ,
		_w4401_
	);
	LUT2 #(
		.INIT('h1)
	) name3628 (
		_w4400_,
		_w4401_,
		_w4402_
	);
	LUT2 #(
		.INIT('h2)
	) name3629 (
		\g35_pad ,
		_w4396_,
		_w4403_
	);
	LUT2 #(
		.INIT('h1)
	) name3630 (
		\g3352_reg/NET0131 ,
		_w2225_,
		_w4404_
	);
	LUT2 #(
		.INIT('h2)
	) name3631 (
		\g35_pad ,
		_w3991_,
		_w4405_
	);
	LUT2 #(
		.INIT('h4)
	) name3632 (
		_w4404_,
		_w4405_,
		_w4406_
	);
	LUT2 #(
		.INIT('h1)
	) name3633 (
		_w4387_,
		_w4406_,
		_w4407_
	);
	LUT2 #(
		.INIT('h2)
	) name3634 (
		\g35_pad ,
		_w2388_,
		_w4408_
	);
	LUT2 #(
		.INIT('h4)
	) name3635 (
		\g35_pad ,
		\g990_reg/NET0131 ,
		_w4409_
	);
	LUT2 #(
		.INIT('h1)
	) name3636 (
		_w4408_,
		_w4409_,
		_w4410_
	);
	LUT2 #(
		.INIT('h1)
	) name3637 (
		\g3703_reg/NET0131 ,
		_w2243_,
		_w4411_
	);
	LUT2 #(
		.INIT('h2)
	) name3638 (
		_w4352_,
		_w4411_,
		_w4412_
	);
	LUT2 #(
		.INIT('h1)
	) name3639 (
		_w4387_,
		_w4412_,
		_w4413_
	);
	LUT2 #(
		.INIT('h1)
	) name3640 (
		\g4054_reg/NET0131 ,
		_w890_,
		_w4414_
	);
	LUT2 #(
		.INIT('h2)
	) name3641 (
		_w4358_,
		_w4414_,
		_w4415_
	);
	LUT2 #(
		.INIT('h1)
	) name3642 (
		_w4387_,
		_w4415_,
		_w4416_
	);
	LUT2 #(
		.INIT('h1)
	) name3643 (
		\g324_reg/NET0131 ,
		\g35_pad ,
		_w4417_
	);
	LUT2 #(
		.INIT('h1)
	) name3644 (
		_w2313_,
		_w4417_,
		_w4418_
	);
	LUT2 #(
		.INIT('h2)
	) name3645 (
		\g262_reg/NET0131 ,
		_w3427_,
		_w4419_
	);
	LUT2 #(
		.INIT('h8)
	) name3646 (
		\g14096_pad ,
		_w3427_,
		_w4420_
	);
	LUT2 #(
		.INIT('h1)
	) name3647 (
		_w4419_,
		_w4420_,
		_w4421_
	);
	LUT2 #(
		.INIT('h2)
	) name3648 (
		\g35_pad ,
		_w4421_,
		_w4422_
	);
	LUT2 #(
		.INIT('h2)
	) name3649 (
		\g232_reg/NET0131 ,
		\g35_pad ,
		_w4423_
	);
	LUT2 #(
		.INIT('h1)
	) name3650 (
		_w4422_,
		_w4423_,
		_w4424_
	);
	LUT2 #(
		.INIT('h2)
	) name3651 (
		\g1008_reg/NET0131 ,
		\g35_pad ,
		_w4425_
	);
	LUT2 #(
		.INIT('h4)
	) name3652 (
		\g1002_reg/NET0131 ,
		_w2373_,
		_w4426_
	);
	LUT2 #(
		.INIT('h2)
	) name3653 (
		_w3882_,
		_w4426_,
		_w4427_
	);
	LUT2 #(
		.INIT('h1)
	) name3654 (
		_w4425_,
		_w4427_,
		_w4428_
	);
	LUT2 #(
		.INIT('h1)
	) name3655 (
		\g645_reg/NET0131 ,
		_w4396_,
		_w4429_
	);
	LUT2 #(
		.INIT('h4)
	) name3656 (
		\g446_reg/NET0131 ,
		_w4396_,
		_w4430_
	);
	LUT2 #(
		.INIT('h2)
	) name3657 (
		\g35_pad ,
		_w4429_,
		_w4431_
	);
	LUT2 #(
		.INIT('h4)
	) name3658 (
		_w4430_,
		_w4431_,
		_w4432_
	);
	LUT2 #(
		.INIT('h4)
	) name3659 (
		\g35_pad ,
		\g546_reg/NET0131 ,
		_w4433_
	);
	LUT2 #(
		.INIT('h4)
	) name3660 (
		\g542_reg/NET0131 ,
		\g691_reg/NET0131 ,
		_w4434_
	);
	LUT2 #(
		.INIT('h2)
	) name3661 (
		_w967_,
		_w4434_,
		_w4435_
	);
	LUT2 #(
		.INIT('h1)
	) name3662 (
		_w4433_,
		_w4435_,
		_w4436_
	);
	LUT2 #(
		.INIT('h1)
	) name3663 (
		\g13895_pad ,
		\g16718_pad ,
		_w4437_
	);
	LUT2 #(
		.INIT('h1)
	) name3664 (
		_w3590_,
		_w4437_,
		_w4438_
	);
	LUT2 #(
		.INIT('h1)
	) name3665 (
		\g13039_pad ,
		\g16603_pad ,
		_w4439_
	);
	LUT2 #(
		.INIT('h4)
	) name3666 (
		\g16624_pad ,
		\g35_pad ,
		_w4440_
	);
	LUT2 #(
		.INIT('h8)
	) name3667 (
		_w4439_,
		_w4440_,
		_w4441_
	);
	LUT2 #(
		.INIT('h4)
	) name3668 (
		_w4438_,
		_w4441_,
		_w4442_
	);
	LUT2 #(
		.INIT('h8)
	) name3669 (
		\g4633_reg/NET0131 ,
		_w2157_,
		_w4443_
	);
	LUT2 #(
		.INIT('h8)
	) name3670 (
		_w2160_,
		_w4443_,
		_w4444_
	);
	LUT2 #(
		.INIT('h4)
	) name3671 (
		_w1068_,
		_w4444_,
		_w4445_
	);
	LUT2 #(
		.INIT('h2)
	) name3672 (
		\g35_pad ,
		_w4445_,
		_w4446_
	);
	LUT2 #(
		.INIT('h8)
	) name3673 (
		\g35_pad ,
		\g4653_reg/NET0131 ,
		_w4447_
	);
	LUT2 #(
		.INIT('h4)
	) name3674 (
		\g4688_reg/NET0131 ,
		_w4447_,
		_w4448_
	);
	LUT2 #(
		.INIT('h2)
	) name3675 (
		\g4688_reg/NET0131 ,
		_w4447_,
		_w4449_
	);
	LUT2 #(
		.INIT('h1)
	) name3676 (
		_w4448_,
		_w4449_,
		_w4450_
	);
	LUT2 #(
		.INIT('h8)
	) name3677 (
		\g4621_reg/NET0131 ,
		\g4639_reg/NET0131 ,
		_w4451_
	);
	LUT2 #(
		.INIT('h8)
	) name3678 (
		\g4628_reg/NET0131 ,
		_w4451_,
		_w4452_
	);
	LUT2 #(
		.INIT('h2)
	) name3679 (
		\g35_pad ,
		\g4643_reg/NET0131 ,
		_w4453_
	);
	LUT2 #(
		.INIT('h4)
	) name3680 (
		_w4452_,
		_w4453_,
		_w4454_
	);
	LUT2 #(
		.INIT('h8)
	) name3681 (
		\g4633_reg/NET0131 ,
		_w4454_,
		_w4455_
	);
	LUT2 #(
		.INIT('h1)
	) name3682 (
		\g4633_reg/NET0131 ,
		\g4643_reg/NET0131 ,
		_w4456_
	);
	LUT2 #(
		.INIT('h8)
	) name3683 (
		_w4451_,
		_w4456_,
		_w4457_
	);
	LUT2 #(
		.INIT('h2)
	) name3684 (
		\g35_pad ,
		_w4457_,
		_w4458_
	);
	LUT2 #(
		.INIT('h2)
	) name3685 (
		\g4628_reg/NET0131 ,
		_w4458_,
		_w4459_
	);
	LUT2 #(
		.INIT('h1)
	) name3686 (
		_w4455_,
		_w4459_,
		_w4460_
	);
	LUT2 #(
		.INIT('h1)
	) name3687 (
		\g2878_reg/NET0131 ,
		\g35_pad ,
		_w4461_
	);
	LUT2 #(
		.INIT('h1)
	) name3688 (
		\g2886_reg/NET0131 ,
		\g2946_reg/NET0131 ,
		_w4462_
	);
	LUT2 #(
		.INIT('h8)
	) name3689 (
		\g35_pad ,
		_w4462_,
		_w4463_
	);
	LUT2 #(
		.INIT('h1)
	) name3690 (
		_w4461_,
		_w4463_,
		_w4464_
	);
	LUT2 #(
		.INIT('h1)
	) name3691 (
		\g11447_pad ,
		\g8783_pad ,
		_w4465_
	);
	LUT2 #(
		.INIT('h1)
	) name3692 (
		\g8784_pad ,
		\g8785_pad ,
		_w4466_
	);
	LUT2 #(
		.INIT('h1)
	) name3693 (
		\g8787_pad ,
		\g8788_pad ,
		_w4467_
	);
	LUT2 #(
		.INIT('h4)
	) name3694 (
		\g8789_pad ,
		_w4467_,
		_w4468_
	);
	LUT2 #(
		.INIT('h8)
	) name3695 (
		_w4465_,
		_w4466_,
		_w4469_
	);
	LUT2 #(
		.INIT('h8)
	) name3696 (
		_w4468_,
		_w4469_,
		_w4470_
	);
	LUT2 #(
		.INIT('h1)
	) name3697 (
		\g4180_reg/NET0131 ,
		\g8786_pad ,
		_w4471_
	);
	LUT2 #(
		.INIT('h4)
	) name3698 (
		_w4470_,
		_w4471_,
		_w4472_
	);
	LUT2 #(
		.INIT('h8)
	) name3699 (
		\g4180_reg/NET0131 ,
		\g8786_pad ,
		_w4473_
	);
	LUT2 #(
		.INIT('h1)
	) name3700 (
		_w4472_,
		_w4473_,
		_w4474_
	);
	LUT2 #(
		.INIT('h2)
	) name3701 (
		\g35_pad ,
		_w4474_,
		_w4475_
	);
	LUT2 #(
		.INIT('h1)
	) name3702 (
		\g2946_reg/NET0131 ,
		\g35_pad ,
		_w4476_
	);
	LUT2 #(
		.INIT('h1)
	) name3703 (
		_w4475_,
		_w4476_,
		_w4477_
	);
	LUT2 #(
		.INIT('h4)
	) name3704 (
		\g4076_reg/NET0131 ,
		_w871_,
		_w4478_
	);
	LUT2 #(
		.INIT('h8)
	) name3705 (
		_w873_,
		_w4478_,
		_w4479_
	);
	LUT2 #(
		.INIT('h8)
	) name3706 (
		_w870_,
		_w4479_,
		_w4480_
	);
	LUT2 #(
		.INIT('h2)
	) name3707 (
		\g35_pad ,
		_w4480_,
		_w4481_
	);
	LUT2 #(
		.INIT('h2)
	) name3708 (
		\g4145_reg/NET0131 ,
		_w4481_,
		_w4482_
	);
	LUT2 #(
		.INIT('h8)
	) name3709 (
		\g4112_reg/NET0131 ,
		_w4481_,
		_w4483_
	);
	LUT2 #(
		.INIT('h1)
	) name3710 (
		_w4482_,
		_w4483_,
		_w4484_
	);
	LUT2 #(
		.INIT('h4)
	) name3711 (
		\g35_pad ,
		\g4369_reg/NET0131 ,
		_w4485_
	);
	LUT2 #(
		.INIT('h4)
	) name3712 (
		\g4462_reg/NET0131 ,
		\g4473_reg/NET0131 ,
		_w4486_
	);
	LUT2 #(
		.INIT('h1)
	) name3713 (
		\g4459_reg/NET0131 ,
		_w4486_,
		_w4487_
	);
	LUT2 #(
		.INIT('h2)
	) name3714 (
		\g35_pad ,
		_w4487_,
		_w4488_
	);
	LUT2 #(
		.INIT('h1)
	) name3715 (
		_w4485_,
		_w4488_,
		_w4489_
	);
	LUT2 #(
		.INIT('h4)
	) name3716 (
		\g35_pad ,
		\g518_reg/NET0131 ,
		_w4490_
	);
	LUT2 #(
		.INIT('h1)
	) name3717 (
		\g528_reg/NET0131 ,
		_w3372_,
		_w4491_
	);
	LUT2 #(
		.INIT('h4)
	) name3718 (
		_w3374_,
		_w4263_,
		_w4492_
	);
	LUT2 #(
		.INIT('h4)
	) name3719 (
		_w4491_,
		_w4492_,
		_w4493_
	);
	LUT2 #(
		.INIT('h1)
	) name3720 (
		_w4490_,
		_w4493_,
		_w4494_
	);
	LUT2 #(
		.INIT('h2)
	) name3721 (
		\g699_reg/NET0131 ,
		_w2206_,
		_w4495_
	);
	LUT2 #(
		.INIT('h1)
	) name3722 (
		_w4396_,
		_w4495_,
		_w4496_
	);
	LUT2 #(
		.INIT('h2)
	) name3723 (
		\g35_pad ,
		_w4496_,
		_w4497_
	);
	LUT2 #(
		.INIT('h4)
	) name3724 (
		\g35_pad ,
		\g681_reg/NET0131 ,
		_w4498_
	);
	LUT2 #(
		.INIT('h1)
	) name3725 (
		_w4497_,
		_w4498_,
		_w4499_
	);
	LUT2 #(
		.INIT('h8)
	) name3726 (
		\g812_reg/NET0131 ,
		\g847_reg/NET0131 ,
		_w4500_
	);
	LUT2 #(
		.INIT('h8)
	) name3727 (
		\g837_reg/NET0131 ,
		_w4500_,
		_w4501_
	);
	LUT2 #(
		.INIT('h8)
	) name3728 (
		_w2206_,
		_w4501_,
		_w4502_
	);
	LUT2 #(
		.INIT('h2)
	) name3729 (
		\g703_reg/NET0131 ,
		_w4502_,
		_w4503_
	);
	LUT2 #(
		.INIT('h8)
	) name3730 (
		\g723_reg/NET0131 ,
		\g822_reg/NET0131 ,
		_w4504_
	);
	LUT2 #(
		.INIT('h4)
	) name3731 (
		\g847_reg/NET0131 ,
		_w4504_,
		_w4505_
	);
	LUT2 #(
		.INIT('h8)
	) name3732 (
		_w2207_,
		_w4505_,
		_w4506_
	);
	LUT2 #(
		.INIT('h1)
	) name3733 (
		_w4503_,
		_w4506_,
		_w4507_
	);
	LUT2 #(
		.INIT('h2)
	) name3734 (
		\g35_pad ,
		_w4507_,
		_w4508_
	);
	LUT2 #(
		.INIT('h4)
	) name3735 (
		\g35_pad ,
		\g847_reg/NET0131 ,
		_w4509_
	);
	LUT2 #(
		.INIT('h1)
	) name3736 (
		_w4508_,
		_w4509_,
		_w4510_
	);
	LUT2 #(
		.INIT('h2)
	) name3737 (
		\g35_pad ,
		_w2206_,
		_w4511_
	);
	LUT2 #(
		.INIT('h2)
	) name3738 (
		\g854_reg/NET0131 ,
		_w4511_,
		_w4512_
	);
	LUT2 #(
		.INIT('h8)
	) name3739 (
		\g847_reg/NET0131 ,
		_w4511_,
		_w4513_
	);
	LUT2 #(
		.INIT('h1)
	) name3740 (
		_w4512_,
		_w4513_,
		_w4514_
	);
	LUT2 #(
		.INIT('h2)
	) name3741 (
		\g35_pad ,
		_w2107_,
		_w4515_
	);
	LUT2 #(
		.INIT('h8)
	) name3742 (
		\g5097_reg/NET0131 ,
		_w4170_,
		_w4516_
	);
	LUT2 #(
		.INIT('h8)
	) name3743 (
		\g35_pad ,
		\g5097_reg/NET0131 ,
		_w4517_
	);
	LUT2 #(
		.INIT('h2)
	) name3744 (
		\g5092_reg/NET0131 ,
		_w2938_,
		_w4518_
	);
	LUT2 #(
		.INIT('h4)
	) name3745 (
		_w4517_,
		_w4518_,
		_w4519_
	);
	LUT2 #(
		.INIT('h1)
	) name3746 (
		_w4516_,
		_w4519_,
		_w4520_
	);
	LUT2 #(
		.INIT('h2)
	) name3747 (
		\g1205_reg/NET0131 ,
		\g35_pad ,
		_w4521_
	);
	LUT2 #(
		.INIT('h1)
	) name3748 (
		\g1221_reg/NET0131 ,
		_w3390_,
		_w4522_
	);
	LUT2 #(
		.INIT('h2)
	) name3749 (
		_w3392_,
		_w4522_,
		_w4523_
	);
	LUT2 #(
		.INIT('h1)
	) name3750 (
		_w4521_,
		_w4523_,
		_w4524_
	);
	LUT2 #(
		.INIT('h2)
	) name3751 (
		\g182_reg/NET0131 ,
		_w2107_,
		_w4525_
	);
	LUT2 #(
		.INIT('h8)
	) name3752 (
		\g446_reg/NET0131 ,
		_w2107_,
		_w4526_
	);
	LUT2 #(
		.INIT('h1)
	) name3753 (
		_w4525_,
		_w4526_,
		_w4527_
	);
	LUT2 #(
		.INIT('h2)
	) name3754 (
		\g35_pad ,
		_w4527_,
		_w4528_
	);
	LUT2 #(
		.INIT('h4)
	) name3755 (
		\g35_pad ,
		\g405_reg/NET0131 ,
		_w4529_
	);
	LUT2 #(
		.INIT('h1)
	) name3756 (
		_w4528_,
		_w4529_,
		_w4530_
	);
	LUT2 #(
		.INIT('h4)
	) name3757 (
		\g837_reg/NET0131 ,
		_w3468_,
		_w4531_
	);
	LUT2 #(
		.INIT('h2)
	) name3758 (
		\g35_pad ,
		_w4531_,
		_w4532_
	);
	LUT2 #(
		.INIT('h2)
	) name3759 (
		\g703_reg/NET0131 ,
		_w4532_,
		_w4533_
	);
	LUT2 #(
		.INIT('h8)
	) name3760 (
		\g827_reg/NET0131 ,
		\g832_reg/NET0131 ,
		_w4534_
	);
	LUT2 #(
		.INIT('h1)
	) name3761 (
		_w4500_,
		_w4534_,
		_w4535_
	);
	LUT2 #(
		.INIT('h2)
	) name3762 (
		_w2206_,
		_w4535_,
		_w4536_
	);
	LUT2 #(
		.INIT('h8)
	) name3763 (
		\g35_pad ,
		\g837_reg/NET0131 ,
		_w4537_
	);
	LUT2 #(
		.INIT('h4)
	) name3764 (
		_w4536_,
		_w4537_,
		_w4538_
	);
	LUT2 #(
		.INIT('h1)
	) name3765 (
		_w4533_,
		_w4538_,
		_w4539_
	);
	LUT2 #(
		.INIT('h8)
	) name3766 (
		\g4064_reg/NET0131 ,
		_w4479_,
		_w4540_
	);
	LUT2 #(
		.INIT('h4)
	) name3767 (
		\g4057_reg/NET0131 ,
		_w4540_,
		_w4541_
	);
	LUT2 #(
		.INIT('h2)
	) name3768 (
		\g4116_reg/NET0131 ,
		_w4541_,
		_w4542_
	);
	LUT2 #(
		.INIT('h8)
	) name3769 (
		\g4145_reg/NET0131 ,
		_w4541_,
		_w4543_
	);
	LUT2 #(
		.INIT('h1)
	) name3770 (
		_w4542_,
		_w4543_,
		_w4544_
	);
	LUT2 #(
		.INIT('h2)
	) name3771 (
		\g35_pad ,
		_w4544_,
		_w4545_
	);
	LUT2 #(
		.INIT('h4)
	) name3772 (
		\g35_pad ,
		\g4112_reg/NET0131 ,
		_w4546_
	);
	LUT2 #(
		.INIT('h1)
	) name3773 (
		_w4545_,
		_w4546_,
		_w4547_
	);
	LUT2 #(
		.INIT('h2)
	) name3774 (
		\g4057_reg/NET0131 ,
		\g4064_reg/NET0131 ,
		_w4548_
	);
	LUT2 #(
		.INIT('h8)
	) name3775 (
		_w4479_,
		_w4548_,
		_w4549_
	);
	LUT2 #(
		.INIT('h2)
	) name3776 (
		\g4119_reg/NET0131 ,
		_w4549_,
		_w4550_
	);
	LUT2 #(
		.INIT('h8)
	) name3777 (
		\g4145_reg/NET0131 ,
		_w4549_,
		_w4551_
	);
	LUT2 #(
		.INIT('h1)
	) name3778 (
		_w4550_,
		_w4551_,
		_w4552_
	);
	LUT2 #(
		.INIT('h2)
	) name3779 (
		\g35_pad ,
		_w4552_,
		_w4553_
	);
	LUT2 #(
		.INIT('h4)
	) name3780 (
		\g35_pad ,
		\g4116_reg/NET0131 ,
		_w4554_
	);
	LUT2 #(
		.INIT('h1)
	) name3781 (
		_w4553_,
		_w4554_,
		_w4555_
	);
	LUT2 #(
		.INIT('h8)
	) name3782 (
		\g4057_reg/NET0131 ,
		_w4540_,
		_w4556_
	);
	LUT2 #(
		.INIT('h2)
	) name3783 (
		\g4122_reg/NET0131 ,
		_w4556_,
		_w4557_
	);
	LUT2 #(
		.INIT('h8)
	) name3784 (
		\g4145_reg/NET0131 ,
		_w4556_,
		_w4558_
	);
	LUT2 #(
		.INIT('h1)
	) name3785 (
		_w4557_,
		_w4558_,
		_w4559_
	);
	LUT2 #(
		.INIT('h2)
	) name3786 (
		\g35_pad ,
		_w4559_,
		_w4560_
	);
	LUT2 #(
		.INIT('h4)
	) name3787 (
		\g35_pad ,
		\g4119_reg/NET0131 ,
		_w4561_
	);
	LUT2 #(
		.INIT('h1)
	) name3788 (
		_w4560_,
		_w4561_,
		_w4562_
	);
	LUT2 #(
		.INIT('h8)
	) name3789 (
		\g4269_reg/NET0131 ,
		_w4226_,
		_w4563_
	);
	LUT2 #(
		.INIT('h8)
	) name3790 (
		\g35_pad ,
		\g4269_reg/NET0131 ,
		_w4564_
	);
	LUT2 #(
		.INIT('h2)
	) name3791 (
		\g35_pad ,
		\g4258_reg/NET0131 ,
		_w4565_
	);
	LUT2 #(
		.INIT('h2)
	) name3792 (
		\g4264_reg/NET0131 ,
		_w4564_,
		_w4566_
	);
	LUT2 #(
		.INIT('h4)
	) name3793 (
		_w4565_,
		_w4566_,
		_w4567_
	);
	LUT2 #(
		.INIT('h1)
	) name3794 (
		_w4563_,
		_w4567_,
		_w4568_
	);
	LUT2 #(
		.INIT('h2)
	) name3795 (
		\g433_reg/NET0131 ,
		_w2206_,
		_w4569_
	);
	LUT2 #(
		.INIT('h8)
	) name3796 (
		\g269_reg/NET0131 ,
		_w2206_,
		_w4570_
	);
	LUT2 #(
		.INIT('h1)
	) name3797 (
		_w4569_,
		_w4570_,
		_w4571_
	);
	LUT2 #(
		.INIT('h2)
	) name3798 (
		\g35_pad ,
		_w4571_,
		_w4572_
	);
	LUT2 #(
		.INIT('h4)
	) name3799 (
		\g35_pad ,
		\g437_reg/NET0131 ,
		_w4573_
	);
	LUT2 #(
		.INIT('h1)
	) name3800 (
		_w4572_,
		_w4573_,
		_w4574_
	);
	LUT2 #(
		.INIT('h2)
	) name3801 (
		\g232_reg/NET0131 ,
		_w3427_,
		_w4575_
	);
	LUT2 #(
		.INIT('h8)
	) name3802 (
		\g14217_pad ,
		_w3427_,
		_w4576_
	);
	LUT2 #(
		.INIT('h1)
	) name3803 (
		_w4575_,
		_w4576_,
		_w4577_
	);
	LUT2 #(
		.INIT('h2)
	) name3804 (
		\g35_pad ,
		_w4577_,
		_w4578_
	);
	LUT2 #(
		.INIT('h2)
	) name3805 (
		\g255_reg/NET0131 ,
		\g35_pad ,
		_w4579_
	);
	LUT2 #(
		.INIT('h1)
	) name3806 (
		_w4578_,
		_w4579_,
		_w4580_
	);
	LUT2 #(
		.INIT('h2)
	) name3807 (
		\g460_reg/NET0131 ,
		_w2107_,
		_w4581_
	);
	LUT2 #(
		.INIT('h8)
	) name3808 (
		\g246_reg/NET0131 ,
		_w2107_,
		_w4582_
	);
	LUT2 #(
		.INIT('h1)
	) name3809 (
		_w4581_,
		_w4582_,
		_w4583_
	);
	LUT2 #(
		.INIT('h2)
	) name3810 (
		\g35_pad ,
		_w4583_,
		_w4584_
	);
	LUT2 #(
		.INIT('h2)
	) name3811 (
		\g168_reg/NET0131 ,
		\g35_pad ,
		_w4585_
	);
	LUT2 #(
		.INIT('h1)
	) name3812 (
		_w4584_,
		_w4585_,
		_w4586_
	);
	LUT2 #(
		.INIT('h2)
	) name3813 (
		\g1548_reg/NET0131 ,
		\g35_pad ,
		_w4587_
	);
	LUT2 #(
		.INIT('h1)
	) name3814 (
		\g1564_reg/NET0131 ,
		_w1380_,
		_w4588_
	);
	LUT2 #(
		.INIT('h2)
	) name3815 (
		\g35_pad ,
		_w1381_,
		_w4589_
	);
	LUT2 #(
		.INIT('h4)
	) name3816 (
		_w4588_,
		_w4589_,
		_w4590_
	);
	LUT2 #(
		.INIT('h1)
	) name3817 (
		_w4587_,
		_w4590_,
		_w4591_
	);
	LUT2 #(
		.INIT('h2)
	) name3818 (
		\g475_reg/NET0131 ,
		_w2206_,
		_w4592_
	);
	LUT2 #(
		.INIT('h8)
	) name3819 (
		\g246_reg/NET0131 ,
		_w2206_,
		_w4593_
	);
	LUT2 #(
		.INIT('h1)
	) name3820 (
		_w4592_,
		_w4593_,
		_w4594_
	);
	LUT2 #(
		.INIT('h2)
	) name3821 (
		\g35_pad ,
		_w4594_,
		_w4595_
	);
	LUT2 #(
		.INIT('h4)
	) name3822 (
		\g35_pad ,
		\g424_reg/NET0131 ,
		_w4596_
	);
	LUT2 #(
		.INIT('h1)
	) name3823 (
		_w4595_,
		_w4596_,
		_w4597_
	);
	LUT2 #(
		.INIT('h2)
	) name3824 (
		\g255_reg/NET0131 ,
		_w3427_,
		_w4598_
	);
	LUT2 #(
		.INIT('h8)
	) name3825 (
		\g14201_pad ,
		_w3427_,
		_w4599_
	);
	LUT2 #(
		.INIT('h1)
	) name3826 (
		_w4598_,
		_w4599_,
		_w4600_
	);
	LUT2 #(
		.INIT('h2)
	) name3827 (
		\g35_pad ,
		_w4600_,
		_w4601_
	);
	LUT2 #(
		.INIT('h2)
	) name3828 (
		\g225_reg/NET0131 ,
		\g35_pad ,
		_w4602_
	);
	LUT2 #(
		.INIT('h1)
	) name3829 (
		_w4601_,
		_w4602_,
		_w4603_
	);
	LUT2 #(
		.INIT('h1)
	) name3830 (
		\g3050_reg/NET0131 ,
		\g5022_reg/NET0131 ,
		_w4604_
	);
	LUT2 #(
		.INIT('h1)
	) name3831 (
		\g5016_reg/NET0131 ,
		_w4604_,
		_w4605_
	);
	LUT2 #(
		.INIT('h8)
	) name3832 (
		_w3953_,
		_w4605_,
		_w4606_
	);
	LUT2 #(
		.INIT('h8)
	) name3833 (
		\g5016_reg/NET0131 ,
		_w4604_,
		_w4607_
	);
	LUT2 #(
		.INIT('h1)
	) name3834 (
		_w4606_,
		_w4607_,
		_w4608_
	);
	LUT2 #(
		.INIT('h2)
	) name3835 (
		\g35_pad ,
		_w4608_,
		_w4609_
	);
	LUT2 #(
		.INIT('h4)
	) name3836 (
		\g35_pad ,
		\g5022_reg/NET0131 ,
		_w4610_
	);
	LUT2 #(
		.INIT('h1)
	) name3837 (
		_w4609_,
		_w4610_,
		_w4611_
	);
	LUT2 #(
		.INIT('h2)
	) name3838 (
		\g3100_reg/NET0131 ,
		\g35_pad ,
		_w4612_
	);
	LUT2 #(
		.INIT('h4)
	) name3839 (
		\g3100_reg/NET0131 ,
		\g5101_reg/NET0131 ,
		_w4613_
	);
	LUT2 #(
		.INIT('h1)
	) name3840 (
		\g3050_reg/NET0131 ,
		_w4613_,
		_w4614_
	);
	LUT2 #(
		.INIT('h4)
	) name3841 (
		\g3096_reg/NET0131 ,
		\g35_pad ,
		_w4615_
	);
	LUT2 #(
		.INIT('h4)
	) name3842 (
		_w4614_,
		_w4615_,
		_w4616_
	);
	LUT2 #(
		.INIT('h1)
	) name3843 (
		_w4612_,
		_w4616_,
		_w4617_
	);
	LUT2 #(
		.INIT('h1)
	) name3844 (
		\g2932_reg/NET0131 ,
		\g2999_reg/NET0131 ,
		_w4618_
	);
	LUT2 #(
		.INIT('h2)
	) name3845 (
		\g35_pad ,
		_w4618_,
		_w4619_
	);
	LUT2 #(
		.INIT('h8)
	) name3846 (
		\g1211_reg/NET0131 ,
		_w3391_,
		_w4620_
	);
	LUT2 #(
		.INIT('h4)
	) name3847 (
		_w2378_,
		_w4620_,
		_w4621_
	);
	LUT2 #(
		.INIT('h1)
	) name3848 (
		\g17291_pad ,
		\g17316_pad ,
		_w4622_
	);
	LUT2 #(
		.INIT('h4)
	) name3849 (
		\g17400_pad ,
		\g35_pad ,
		_w4623_
	);
	LUT2 #(
		.INIT('h8)
	) name3850 (
		_w4622_,
		_w4623_,
		_w4624_
	);
	LUT2 #(
		.INIT('h4)
	) name3851 (
		_w4621_,
		_w4624_,
		_w4625_
	);
	LUT2 #(
		.INIT('h1)
	) name3852 (
		\g35_pad ,
		\g4072_reg/NET0131 ,
		_w4626_
	);
	LUT2 #(
		.INIT('h1)
	) name3853 (
		\g417_reg/NET0131 ,
		_w2206_,
		_w4627_
	);
	LUT2 #(
		.INIT('h4)
	) name3854 (
		\g446_reg/NET0131 ,
		_w2206_,
		_w4628_
	);
	LUT2 #(
		.INIT('h2)
	) name3855 (
		\g35_pad ,
		_w4627_,
		_w4629_
	);
	LUT2 #(
		.INIT('h4)
	) name3856 (
		_w4628_,
		_w4629_,
		_w4630_
	);
	LUT2 #(
		.INIT('h1)
	) name3857 (
		\g4311_reg/NET0131 ,
		_w2161_,
		_w4631_
	);
	LUT2 #(
		.INIT('h1)
	) name3858 (
		_w3399_,
		_w4631_,
		_w4632_
	);
	LUT2 #(
		.INIT('h8)
	) name3859 (
		_w3398_,
		_w4632_,
		_w4633_
	);
	LUT2 #(
		.INIT('h4)
	) name3860 (
		\g35_pad ,
		\g5033_reg/NET0131 ,
		_w4634_
	);
	LUT2 #(
		.INIT('h1)
	) name3861 (
		_w3495_,
		_w3501_,
		_w4635_
	);
	LUT2 #(
		.INIT('h2)
	) name3862 (
		\g5037_reg/NET0131 ,
		_w3571_,
		_w4636_
	);
	LUT2 #(
		.INIT('h8)
	) name3863 (
		_w3572_,
		_w4636_,
		_w4637_
	);
	LUT2 #(
		.INIT('h8)
	) name3864 (
		_w4635_,
		_w4637_,
		_w4638_
	);
	LUT2 #(
		.INIT('h2)
	) name3865 (
		\g35_pad ,
		\g5037_reg/NET0131 ,
		_w4639_
	);
	LUT2 #(
		.INIT('h4)
	) name3866 (
		_w4635_,
		_w4639_,
		_w4640_
	);
	LUT2 #(
		.INIT('h1)
	) name3867 (
		_w4634_,
		_w4638_,
		_w4641_
	);
	LUT2 #(
		.INIT('h4)
	) name3868 (
		_w4640_,
		_w4641_,
		_w4642_
	);
	LUT2 #(
		.INIT('h8)
	) name3869 (
		_w2377_,
		_w3298_,
		_w4643_
	);
	LUT2 #(
		.INIT('h2)
	) name3870 (
		\g35_pad ,
		_w4643_,
		_w4644_
	);
	LUT2 #(
		.INIT('h2)
	) name3871 (
		\g1041_reg/NET0131 ,
		_w4644_,
		_w4645_
	);
	LUT2 #(
		.INIT('h2)
	) name3872 (
		\g1008_reg/NET0131 ,
		\g1041_reg/NET0131 ,
		_w4646_
	);
	LUT2 #(
		.INIT('h2)
	) name3873 (
		_w2377_,
		_w4646_,
		_w4647_
	);
	LUT2 #(
		.INIT('h2)
	) name3874 (
		\g35_pad ,
		_w4647_,
		_w4648_
	);
	LUT2 #(
		.INIT('h8)
	) name3875 (
		\g1046_reg/NET0131 ,
		_w4648_,
		_w4649_
	);
	LUT2 #(
		.INIT('h1)
	) name3876 (
		_w4645_,
		_w4649_,
		_w4650_
	);
	LUT2 #(
		.INIT('h1)
	) name3877 (
		\g392_reg/NET0131 ,
		_w2206_,
		_w4651_
	);
	LUT2 #(
		.INIT('h4)
	) name3878 (
		\g703_reg/NET0131 ,
		\g854_reg/NET0131 ,
		_w4652_
	);
	LUT2 #(
		.INIT('h2)
	) name3879 (
		_w2206_,
		_w4652_,
		_w4653_
	);
	LUT2 #(
		.INIT('h1)
	) name3880 (
		_w4651_,
		_w4653_,
		_w4654_
	);
	LUT2 #(
		.INIT('h2)
	) name3881 (
		\g35_pad ,
		_w4654_,
		_w4655_
	);
	LUT2 #(
		.INIT('h1)
	) name3882 (
		\g35_pad ,
		\g401_reg/NET0131 ,
		_w4656_
	);
	LUT2 #(
		.INIT('h1)
	) name3883 (
		_w4655_,
		_w4656_,
		_w4657_
	);
	LUT2 #(
		.INIT('h2)
	) name3884 (
		\g1036_reg/NET0131 ,
		\g35_pad ,
		_w4658_
	);
	LUT2 #(
		.INIT('h1)
	) name3885 (
		\g1041_reg/NET0131 ,
		_w2377_,
		_w4659_
	);
	LUT2 #(
		.INIT('h2)
	) name3886 (
		_w4648_,
		_w4659_,
		_w4660_
	);
	LUT2 #(
		.INIT('h1)
	) name3887 (
		_w4658_,
		_w4660_,
		_w4661_
	);
	LUT2 #(
		.INIT('h4)
	) name3888 (
		\g35_pad ,
		\g4358_reg/NET0131 ,
		_w4662_
	);
	LUT2 #(
		.INIT('h2)
	) name3889 (
		\g4340_reg/NET0131 ,
		\g4584_reg/NET0131 ,
		_w4663_
	);
	LUT2 #(
		.INIT('h1)
	) name3890 (
		\g4593_reg/NET0131 ,
		\g4601_reg/NET0131 ,
		_w4664_
	);
	LUT2 #(
		.INIT('h1)
	) name3891 (
		\g4608_reg/NET0131 ,
		\g4616_reg/NET0131 ,
		_w4665_
	);
	LUT2 #(
		.INIT('h8)
	) name3892 (
		_w4664_,
		_w4665_,
		_w4666_
	);
	LUT2 #(
		.INIT('h8)
	) name3893 (
		_w3907_,
		_w4663_,
		_w4667_
	);
	LUT2 #(
		.INIT('h8)
	) name3894 (
		_w4666_,
		_w4667_,
		_w4668_
	);
	LUT2 #(
		.INIT('h8)
	) name3895 (
		_w3906_,
		_w4443_,
		_w4669_
	);
	LUT2 #(
		.INIT('h8)
	) name3896 (
		_w4668_,
		_w4669_,
		_w4670_
	);
	LUT2 #(
		.INIT('h1)
	) name3897 (
		_w4662_,
		_w4670_,
		_w4671_
	);
	LUT2 #(
		.INIT('h4)
	) name3898 (
		\g35_pad ,
		\g376_reg/NET0131 ,
		_w4672_
	);
	LUT2 #(
		.INIT('h1)
	) name3899 (
		\g385_reg/NET0131 ,
		_w987_,
		_w4673_
	);
	LUT2 #(
		.INIT('h2)
	) name3900 (
		\g35_pad ,
		_w2205_,
		_w4674_
	);
	LUT2 #(
		.INIT('h4)
	) name3901 (
		_w4673_,
		_w4674_,
		_w4675_
	);
	LUT2 #(
		.INIT('h1)
	) name3902 (
		_w4672_,
		_w4675_,
		_w4676_
	);
	LUT2 #(
		.INIT('h4)
	) name3903 (
		\g35_pad ,
		\g5069_reg/NET0131 ,
		_w4677_
	);
	LUT2 #(
		.INIT('h1)
	) name3904 (
		_w3572_,
		_w4677_,
		_w4678_
	);
	LUT2 #(
		.INIT('h4)
	) name3905 (
		\g35_pad ,
		\g4284_reg/NET0131 ,
		_w4679_
	);
	LUT2 #(
		.INIT('h2)
	) name3906 (
		\g35_pad ,
		\g4291_reg/NET0131 ,
		_w4680_
	);
	LUT2 #(
		.INIT('h1)
	) name3907 (
		_w4679_,
		_w4680_,
		_w4681_
	);
	LUT2 #(
		.INIT('h1)
	) name3908 (
		\g2902_reg/NET0131 ,
		\g35_pad ,
		_w4682_
	);
	LUT2 #(
		.INIT('h4)
	) name3909 (
		\g2917_reg/NET0131 ,
		\g35_pad ,
		_w4683_
	);
	LUT2 #(
		.INIT('h8)
	) name3910 (
		_w816_,
		_w4683_,
		_w4684_
	);
	LUT2 #(
		.INIT('h8)
	) name3911 (
		_w818_,
		_w4684_,
		_w4685_
	);
	LUT2 #(
		.INIT('h1)
	) name3912 (
		_w4682_,
		_w4685_,
		_w4686_
	);
	LUT2 #(
		.INIT('h1)
	) name3913 (
		\g29214_pad ,
		\g35_pad ,
		_w4687_
	);
	LUT2 #(
		.INIT('h4)
	) name3914 (
		\g2848_reg/NET0131 ,
		_w1009_,
		_w4688_
	);
	LUT2 #(
		.INIT('h1)
	) name3915 (
		_w4687_,
		_w4688_,
		_w4689_
	);
	LUT2 #(
		.INIT('h4)
	) name3916 (
		\g35_pad ,
		\g4643_reg/NET0131 ,
		_w4690_
	);
	LUT2 #(
		.INIT('h1)
	) name3917 (
		\g4340_reg/NET0131 ,
		_w2158_,
		_w4691_
	);
	LUT2 #(
		.INIT('h2)
	) name3918 (
		_w3607_,
		_w4691_,
		_w4692_
	);
	LUT2 #(
		.INIT('h1)
	) name3919 (
		_w4690_,
		_w4692_,
		_w4693_
	);
	LUT2 #(
		.INIT('h2)
	) name3920 (
		\g35_pad ,
		_w2589_,
		_w4694_
	);
	LUT2 #(
		.INIT('h2)
	) name3921 (
		\g35_pad ,
		_w2331_,
		_w4695_
	);
	LUT2 #(
		.INIT('h2)
	) name3922 (
		\g35_pad ,
		_w2447_,
		_w4696_
	);
	LUT2 #(
		.INIT('h2)
	) name3923 (
		\g35_pad ,
		_w2344_,
		_w4697_
	);
	LUT2 #(
		.INIT('h8)
	) name3924 (
		\g513_reg/NET0131 ,
		_w3371_,
		_w4698_
	);
	LUT2 #(
		.INIT('h2)
	) name3925 (
		\g499_reg/NET0131 ,
		_w4698_,
		_w4699_
	);
	LUT2 #(
		.INIT('h2)
	) name3926 (
		\g518_reg/NET0131 ,
		_w3375_,
		_w4700_
	);
	LUT2 #(
		.INIT('h2)
	) name3927 (
		_w3371_,
		_w4700_,
		_w4701_
	);
	LUT2 #(
		.INIT('h1)
	) name3928 (
		_w4699_,
		_w4701_,
		_w4702_
	);
	LUT2 #(
		.INIT('h2)
	) name3929 (
		\g35_pad ,
		_w4702_,
		_w4703_
	);
	LUT2 #(
		.INIT('h4)
	) name3930 (
		\g35_pad ,
		\g5112_reg/NET0131 ,
		_w4704_
	);
	LUT2 #(
		.INIT('h2)
	) name3931 (
		\g3096_reg/NET0131 ,
		\g5112_reg/NET0131 ,
		_w4705_
	);
	LUT2 #(
		.INIT('h1)
	) name3932 (
		\g5022_reg/NET0131 ,
		_w4705_,
		_w4706_
	);
	LUT2 #(
		.INIT('h2)
	) name3933 (
		\g35_pad ,
		\g5101_reg/NET0131 ,
		_w4707_
	);
	LUT2 #(
		.INIT('h4)
	) name3934 (
		_w4706_,
		_w4707_,
		_w4708_
	);
	LUT2 #(
		.INIT('h1)
	) name3935 (
		_w4704_,
		_w4708_,
		_w4709_
	);
	LUT2 #(
		.INIT('h2)
	) name3936 (
		\g35_pad ,
		_w4153_,
		_w4710_
	);
	LUT2 #(
		.INIT('h8)
	) name3937 (
		\g5152_reg/NET0131 ,
		_w4710_,
		_w4711_
	);
	LUT2 #(
		.INIT('h2)
	) name3938 (
		\g35_pad ,
		\g5142_reg/NET0131 ,
		_w4712_
	);
	LUT2 #(
		.INIT('h1)
	) name3939 (
		\g5148_reg/NET0131 ,
		_w4712_,
		_w4713_
	);
	LUT2 #(
		.INIT('h8)
	) name3940 (
		\g5148_reg/NET0131 ,
		_w4712_,
		_w4714_
	);
	LUT2 #(
		.INIT('h1)
	) name3941 (
		_w4713_,
		_w4714_,
		_w4715_
	);
	LUT2 #(
		.INIT('h4)
	) name3942 (
		_w4710_,
		_w4715_,
		_w4716_
	);
	LUT2 #(
		.INIT('h1)
	) name3943 (
		_w4711_,
		_w4716_,
		_w4717_
	);
	LUT2 #(
		.INIT('h2)
	) name3944 (
		\g35_pad ,
		_w2033_,
		_w4718_
	);
	LUT2 #(
		.INIT('h4)
	) name3945 (
		_w2041_,
		_w4718_,
		_w4719_
	);
	LUT2 #(
		.INIT('h8)
	) name3946 (
		\g1300_reg/NET0131 ,
		\g35_pad ,
		_w4720_
	);
	LUT2 #(
		.INIT('h2)
	) name3947 (
		\g1442_reg/NET0131 ,
		\g1495_reg/NET0131 ,
		_w4721_
	);
	LUT2 #(
		.INIT('h8)
	) name3948 (
		_w1206_,
		_w4721_,
		_w4722_
	);
	LUT2 #(
		.INIT('h2)
	) name3949 (
		\g35_pad ,
		_w4722_,
		_w4723_
	);
	LUT2 #(
		.INIT('h2)
	) name3950 (
		\g1484_reg/NET0131 ,
		_w4723_,
		_w4724_
	);
	LUT2 #(
		.INIT('h2)
	) name3951 (
		_w4720_,
		_w4724_,
		_w4725_
	);
	LUT2 #(
		.INIT('h4)
	) name3952 (
		_w4720_,
		_w4724_,
		_w4726_
	);
	LUT2 #(
		.INIT('h1)
	) name3953 (
		_w4725_,
		_w4726_,
		_w4727_
	);
	LUT2 #(
		.INIT('h8)
	) name3954 (
		\g1448_reg/NET0131 ,
		\g35_pad ,
		_w4728_
	);
	LUT2 #(
		.INIT('h8)
	) name3955 (
		_w1183_,
		_w4721_,
		_w4729_
	);
	LUT2 #(
		.INIT('h2)
	) name3956 (
		\g35_pad ,
		_w4729_,
		_w4730_
	);
	LUT2 #(
		.INIT('h2)
	) name3957 (
		\g1454_reg/NET0131 ,
		_w4730_,
		_w4731_
	);
	LUT2 #(
		.INIT('h2)
	) name3958 (
		_w4728_,
		_w4731_,
		_w4732_
	);
	LUT2 #(
		.INIT('h4)
	) name3959 (
		_w4728_,
		_w4731_,
		_w4733_
	);
	LUT2 #(
		.INIT('h1)
	) name3960 (
		_w4732_,
		_w4733_,
		_w4734_
	);
	LUT2 #(
		.INIT('h8)
	) name3961 (
		\g1472_reg/NET0131 ,
		\g35_pad ,
		_w4735_
	);
	LUT2 #(
		.INIT('h8)
	) name3962 (
		_w1195_,
		_w4721_,
		_w4736_
	);
	LUT2 #(
		.INIT('h2)
	) name3963 (
		\g35_pad ,
		_w4736_,
		_w4737_
	);
	LUT2 #(
		.INIT('h2)
	) name3964 (
		\g1467_reg/NET0131 ,
		_w4737_,
		_w4738_
	);
	LUT2 #(
		.INIT('h2)
	) name3965 (
		_w4735_,
		_w4738_,
		_w4739_
	);
	LUT2 #(
		.INIT('h4)
	) name3966 (
		_w4735_,
		_w4738_,
		_w4740_
	);
	LUT2 #(
		.INIT('h1)
	) name3967 (
		_w4739_,
		_w4740_,
		_w4741_
	);
	LUT2 #(
		.INIT('h8)
	) name3968 (
		\g1478_reg/NET0131 ,
		\g35_pad ,
		_w4742_
	);
	LUT2 #(
		.INIT('h8)
	) name3969 (
		_w1170_,
		_w4721_,
		_w4743_
	);
	LUT2 #(
		.INIT('h2)
	) name3970 (
		\g35_pad ,
		_w4743_,
		_w4744_
	);
	LUT2 #(
		.INIT('h2)
	) name3971 (
		\g1437_reg/NET0131 ,
		_w4744_,
		_w4745_
	);
	LUT2 #(
		.INIT('h2)
	) name3972 (
		_w4742_,
		_w4745_,
		_w4746_
	);
	LUT2 #(
		.INIT('h4)
	) name3973 (
		_w4742_,
		_w4745_,
		_w4747_
	);
	LUT2 #(
		.INIT('h1)
	) name3974 (
		_w4746_,
		_w4747_,
		_w4748_
	);
	LUT2 #(
		.INIT('h4)
	) name3975 (
		\g35_pad ,
		\g5016_reg/NET0131 ,
		_w4749_
	);
	LUT2 #(
		.INIT('h1)
	) name3976 (
		_w3493_,
		_w3499_,
		_w4750_
	);
	LUT2 #(
		.INIT('h8)
	) name3977 (
		\g35_pad ,
		\g5029_reg/NET0131 ,
		_w4751_
	);
	LUT2 #(
		.INIT('h8)
	) name3978 (
		_w4750_,
		_w4751_,
		_w4752_
	);
	LUT2 #(
		.INIT('h8)
	) name3979 (
		_w3953_,
		_w4752_,
		_w4753_
	);
	LUT2 #(
		.INIT('h2)
	) name3980 (
		\g35_pad ,
		\g5029_reg/NET0131 ,
		_w4754_
	);
	LUT2 #(
		.INIT('h4)
	) name3981 (
		_w4750_,
		_w4754_,
		_w4755_
	);
	LUT2 #(
		.INIT('h1)
	) name3982 (
		_w4749_,
		_w4755_,
		_w4756_
	);
	LUT2 #(
		.INIT('h4)
	) name3983 (
		_w4753_,
		_w4756_,
		_w4757_
	);
	LUT2 #(
		.INIT('h1)
	) name3984 (
		\g4646_reg/NET0131 ,
		\g4674_reg/NET0131 ,
		_w4758_
	);
	LUT2 #(
		.INIT('h4)
	) name3985 (
		\g4681_reg/NET0131 ,
		_w4758_,
		_w4759_
	);
	LUT2 #(
		.INIT('h8)
	) name3986 (
		_w2397_,
		_w4759_,
		_w4760_
	);
	LUT2 #(
		.INIT('h4)
	) name3987 (
		\g35_pad ,
		\g4621_reg/NET0131 ,
		_w4761_
	);
	LUT2 #(
		.INIT('h1)
	) name3988 (
		\g4628_reg/NET0131 ,
		_w4451_,
		_w4762_
	);
	LUT2 #(
		.INIT('h2)
	) name3989 (
		_w4454_,
		_w4762_,
		_w4763_
	);
	LUT2 #(
		.INIT('h1)
	) name3990 (
		_w4761_,
		_w4763_,
		_w4764_
	);
	LUT2 #(
		.INIT('h2)
	) name3991 (
		\g5128_reg/NET0131 ,
		_w4153_,
		_w4765_
	);
	LUT2 #(
		.INIT('h4)
	) name3992 (
		\g5128_reg/NET0131 ,
		_w4153_,
		_w4766_
	);
	LUT2 #(
		.INIT('h1)
	) name3993 (
		_w4765_,
		_w4766_,
		_w4767_
	);
	LUT2 #(
		.INIT('h2)
	) name3994 (
		\g35_pad ,
		_w4767_,
		_w4768_
	);
	LUT2 #(
		.INIT('h4)
	) name3995 (
		\g35_pad ,
		\g5124_reg/NET0131 ,
		_w4769_
	);
	LUT2 #(
		.INIT('h1)
	) name3996 (
		_w4768_,
		_w4769_,
		_w4770_
	);
	LUT2 #(
		.INIT('h2)
	) name3997 (
		\g3119_reg/NET0131 ,
		_w4153_,
		_w4771_
	);
	LUT2 #(
		.INIT('h4)
	) name3998 (
		\g3119_reg/NET0131 ,
		_w4153_,
		_w4772_
	);
	LUT2 #(
		.INIT('h1)
	) name3999 (
		_w4771_,
		_w4772_,
		_w4773_
	);
	LUT2 #(
		.INIT('h2)
	) name4000 (
		\g35_pad ,
		_w4773_,
		_w4774_
	);
	LUT2 #(
		.INIT('h2)
	) name4001 (
		\g3115_reg/NET0131 ,
		\g35_pad ,
		_w4775_
	);
	LUT2 #(
		.INIT('h1)
	) name4002 (
		_w4774_,
		_w4775_,
		_w4776_
	);
	LUT2 #(
		.INIT('h2)
	) name4003 (
		\g35_pad ,
		_w3371_,
		_w4777_
	);
	LUT2 #(
		.INIT('h2)
	) name4004 (
		\g3470_reg/NET0131 ,
		_w4153_,
		_w4778_
	);
	LUT2 #(
		.INIT('h4)
	) name4005 (
		\g3470_reg/NET0131 ,
		_w4153_,
		_w4779_
	);
	LUT2 #(
		.INIT('h1)
	) name4006 (
		_w4778_,
		_w4779_,
		_w4780_
	);
	LUT2 #(
		.INIT('h2)
	) name4007 (
		\g35_pad ,
		_w4780_,
		_w4781_
	);
	LUT2 #(
		.INIT('h2)
	) name4008 (
		\g3466_reg/NET0131 ,
		\g35_pad ,
		_w4782_
	);
	LUT2 #(
		.INIT('h1)
	) name4009 (
		_w4781_,
		_w4782_,
		_w4783_
	);
	LUT2 #(
		.INIT('h2)
	) name4010 (
		\g370_reg/NET0131 ,
		_w2547_,
		_w4784_
	);
	LUT2 #(
		.INIT('h8)
	) name4011 (
		_w975_,
		_w2517_,
		_w4785_
	);
	LUT2 #(
		.INIT('h1)
	) name4012 (
		_w4784_,
		_w4785_,
		_w4786_
	);
	LUT2 #(
		.INIT('h2)
	) name4013 (
		\g35_pad ,
		_w4786_,
		_w4787_
	);
	LUT2 #(
		.INIT('h2)
	) name4014 (
		\g358_reg/NET0131 ,
		\g35_pad ,
		_w4788_
	);
	LUT2 #(
		.INIT('h1)
	) name4015 (
		_w4787_,
		_w4788_,
		_w4789_
	);
	LUT2 #(
		.INIT('h2)
	) name4016 (
		\g3821_reg/NET0131 ,
		_w4153_,
		_w4790_
	);
	LUT2 #(
		.INIT('h4)
	) name4017 (
		\g3821_reg/NET0131 ,
		_w4153_,
		_w4791_
	);
	LUT2 #(
		.INIT('h1)
	) name4018 (
		_w4790_,
		_w4791_,
		_w4792_
	);
	LUT2 #(
		.INIT('h2)
	) name4019 (
		\g35_pad ,
		_w4792_,
		_w4793_
	);
	LUT2 #(
		.INIT('h4)
	) name4020 (
		\g35_pad ,
		\g3817_reg/NET0131 ,
		_w4794_
	);
	LUT2 #(
		.INIT('h1)
	) name4021 (
		_w4793_,
		_w4794_,
		_w4795_
	);
	LUT2 #(
		.INIT('h2)
	) name4022 (
		\g209_reg/NET0131 ,
		_w1475_,
		_w4796_
	);
	LUT2 #(
		.INIT('h8)
	) name4023 (
		\g8358_pad ,
		_w1477_,
		_w4797_
	);
	LUT2 #(
		.INIT('h1)
	) name4024 (
		_w4796_,
		_w4797_,
		_w4798_
	);
	LUT2 #(
		.INIT('h2)
	) name4025 (
		\g35_pad ,
		_w4798_,
		_w4799_
	);
	LUT2 #(
		.INIT('h4)
	) name4026 (
		\g8358_pad ,
		_w1475_,
		_w4800_
	);
	LUT2 #(
		.INIT('h2)
	) name4027 (
		\g35_pad ,
		_w4800_,
		_w4801_
	);
	LUT2 #(
		.INIT('h2)
	) name4028 (
		\g191_reg/NET0131 ,
		_w4801_,
		_w4802_
	);
	LUT2 #(
		.INIT('h1)
	) name4029 (
		_w4799_,
		_w4802_,
		_w4803_
	);
	LUT2 #(
		.INIT('h4)
	) name4030 (
		\g35_pad ,
		\g4180_reg/NET0131 ,
		_w4804_
	);
	LUT2 #(
		.INIT('h2)
	) name4031 (
		\g35_pad ,
		_w1789_,
		_w4805_
	);
	LUT2 #(
		.INIT('h1)
	) name4032 (
		_w4804_,
		_w4805_,
		_w4806_
	);
	LUT2 #(
		.INIT('h2)
	) name4033 (
		\g35_pad ,
		\g4281_reg/NET0131 ,
		_w4807_
	);
	LUT2 #(
		.INIT('h4)
	) name4034 (
		\g35_pad ,
		\g4245_reg/NET0131 ,
		_w4808_
	);
	LUT2 #(
		.INIT('h1)
	) name4035 (
		_w4807_,
		_w4808_,
		_w4809_
	);
	LUT2 #(
		.INIT('h8)
	) name4036 (
		\g1183_reg/NET0131 ,
		_w3538_,
		_w4810_
	);
	LUT2 #(
		.INIT('h2)
	) name4037 (
		\g962_reg/NET0131 ,
		_w4810_,
		_w4811_
	);
	LUT2 #(
		.INIT('h8)
	) name4038 (
		\g996_reg/NET0131 ,
		_w4810_,
		_w4812_
	);
	LUT2 #(
		.INIT('h1)
	) name4039 (
		_w4811_,
		_w4812_,
		_w4813_
	);
	LUT2 #(
		.INIT('h2)
	) name4040 (
		\g35_pad ,
		_w4813_,
		_w4814_
	);
	LUT2 #(
		.INIT('h2)
	) name4041 (
		\g1178_reg/NET0131 ,
		\g35_pad ,
		_w4815_
	);
	LUT2 #(
		.INIT('h1)
	) name4042 (
		_w4814_,
		_w4815_,
		_w4816_
	);
	LUT2 #(
		.INIT('h2)
	) name4043 (
		_w3371_,
		_w3375_,
		_w4817_
	);
	LUT2 #(
		.INIT('h2)
	) name4044 (
		\g35_pad ,
		_w4817_,
		_w4818_
	);
	LUT2 #(
		.INIT('h1)
	) name4045 (
		\g499_reg/NET0131 ,
		_w4818_,
		_w4819_
	);
	LUT2 #(
		.INIT('h4)
	) name4046 (
		\g504_reg/NET0131 ,
		_w4777_,
		_w4820_
	);
	LUT2 #(
		.INIT('h1)
	) name4047 (
		_w4819_,
		_w4820_,
		_w4821_
	);
	LUT2 #(
		.INIT('h2)
	) name4048 (
		\g35_pad ,
		\g4308_reg/NET0131 ,
		_w4822_
	);
	LUT2 #(
		.INIT('h2)
	) name4049 (
		\g504_reg/NET0131 ,
		_w4818_,
		_w4823_
	);
	LUT2 #(
		.INIT('h8)
	) name4050 (
		\g513_reg/NET0131 ,
		_w4777_,
		_w4824_
	);
	LUT2 #(
		.INIT('h1)
	) name4051 (
		_w4823_,
		_w4824_,
		_w4825_
	);
	LUT2 #(
		.INIT('h1)
	) name4052 (
		\g2748_reg/NET0131 ,
		\g35_pad ,
		_w4826_
	);
	LUT2 #(
		.INIT('h8)
	) name4053 (
		\g3143_reg/NET0131 ,
		_w4710_,
		_w4827_
	);
	LUT2 #(
		.INIT('h4)
	) name4054 (
		\g3133_reg/NET0131 ,
		\g35_pad ,
		_w4828_
	);
	LUT2 #(
		.INIT('h1)
	) name4055 (
		\g3139_reg/NET0131 ,
		_w4828_,
		_w4829_
	);
	LUT2 #(
		.INIT('h8)
	) name4056 (
		\g3139_reg/NET0131 ,
		_w4828_,
		_w4830_
	);
	LUT2 #(
		.INIT('h1)
	) name4057 (
		_w4829_,
		_w4830_,
		_w4831_
	);
	LUT2 #(
		.INIT('h4)
	) name4058 (
		_w4710_,
		_w4831_,
		_w4832_
	);
	LUT2 #(
		.INIT('h1)
	) name4059 (
		_w4827_,
		_w4832_,
		_w4833_
	);
	LUT2 #(
		.INIT('h8)
	) name4060 (
		\g3494_reg/NET0131 ,
		_w4710_,
		_w4834_
	);
	LUT2 #(
		.INIT('h4)
	) name4061 (
		\g3484_reg/NET0131 ,
		\g35_pad ,
		_w4835_
	);
	LUT2 #(
		.INIT('h1)
	) name4062 (
		\g3490_reg/NET0131 ,
		_w4835_,
		_w4836_
	);
	LUT2 #(
		.INIT('h8)
	) name4063 (
		\g3490_reg/NET0131 ,
		_w4835_,
		_w4837_
	);
	LUT2 #(
		.INIT('h1)
	) name4064 (
		_w4836_,
		_w4837_,
		_w4838_
	);
	LUT2 #(
		.INIT('h4)
	) name4065 (
		_w4710_,
		_w4838_,
		_w4839_
	);
	LUT2 #(
		.INIT('h1)
	) name4066 (
		_w4834_,
		_w4839_,
		_w4840_
	);
	LUT2 #(
		.INIT('h8)
	) name4067 (
		\g3845_reg/NET0131 ,
		_w4710_,
		_w4841_
	);
	LUT2 #(
		.INIT('h2)
	) name4068 (
		\g35_pad ,
		\g3835_reg/NET0131 ,
		_w4842_
	);
	LUT2 #(
		.INIT('h1)
	) name4069 (
		\g3841_reg/NET0131 ,
		_w4842_,
		_w4843_
	);
	LUT2 #(
		.INIT('h8)
	) name4070 (
		\g3841_reg/NET0131 ,
		_w4842_,
		_w4844_
	);
	LUT2 #(
		.INIT('h1)
	) name4071 (
		_w4843_,
		_w4844_,
		_w4845_
	);
	LUT2 #(
		.INIT('h4)
	) name4072 (
		_w4710_,
		_w4845_,
		_w4846_
	);
	LUT2 #(
		.INIT('h1)
	) name4073 (
		_w4841_,
		_w4846_,
		_w4847_
	);
	LUT2 #(
		.INIT('h8)
	) name4074 (
		\g4076_reg/NET0131 ,
		\g4087_reg/NET0131 ,
		_w4848_
	);
	LUT2 #(
		.INIT('h4)
	) name4075 (
		\g4093_reg/NET0131 ,
		\g4098_reg/NET0131 ,
		_w4849_
	);
	LUT2 #(
		.INIT('h8)
	) name4076 (
		_w4848_,
		_w4849_,
		_w4850_
	);
	LUT2 #(
		.INIT('h8)
	) name4077 (
		_w870_,
		_w871_,
		_w4851_
	);
	LUT2 #(
		.INIT('h8)
	) name4078 (
		_w4850_,
		_w4851_,
		_w4852_
	);
	LUT2 #(
		.INIT('h2)
	) name4079 (
		\g35_pad ,
		_w4852_,
		_w4853_
	);
	LUT2 #(
		.INIT('h4)
	) name4080 (
		\g4643_reg/NET0131 ,
		_w2157_,
		_w4854_
	);
	LUT2 #(
		.INIT('h2)
	) name4081 (
		\g35_pad ,
		_w4854_,
		_w4855_
	);
	LUT2 #(
		.INIT('h1)
	) name4082 (
		\g35_pad ,
		\g4639_reg/NET0131 ,
		_w4856_
	);
	LUT2 #(
		.INIT('h1)
	) name4083 (
		_w4855_,
		_w4856_,
		_w4857_
	);
	LUT2 #(
		.INIT('h4)
	) name4084 (
		\g4621_reg/NET0131 ,
		\g4639_reg/NET0131 ,
		_w4858_
	);
	LUT2 #(
		.INIT('h8)
	) name4085 (
		_w4453_,
		_w4858_,
		_w4859_
	);
	LUT2 #(
		.INIT('h1)
	) name4086 (
		_w4857_,
		_w4859_,
		_w4860_
	);
	LUT2 #(
		.INIT('h1)
	) name4087 (
		\g2965_reg/NET0131 ,
		\g35_pad ,
		_w4861_
	);
	LUT2 #(
		.INIT('h2)
	) name4088 (
		\g1306_reg/NET0131 ,
		\g2975_reg/NET0131 ,
		_w4862_
	);
	LUT2 #(
		.INIT('h8)
	) name4089 (
		\g35_pad ,
		\g962_reg/NET0131 ,
		_w4863_
	);
	LUT2 #(
		.INIT('h8)
	) name4090 (
		_w4862_,
		_w4863_,
		_w4864_
	);
	LUT2 #(
		.INIT('h1)
	) name4091 (
		_w4861_,
		_w4864_,
		_w4865_
	);
	LUT2 #(
		.INIT('h8)
	) name4092 (
		\g518_reg/NET0131 ,
		_w4777_,
		_w4866_
	);
	LUT2 #(
		.INIT('h2)
	) name4093 (
		\g513_reg/NET0131 ,
		_w4818_,
		_w4867_
	);
	LUT2 #(
		.INIT('h1)
	) name4094 (
		_w4866_,
		_w4867_,
		_w4868_
	);
	LUT2 #(
		.INIT('h8)
	) name4095 (
		\g1495_reg/NET0131 ,
		_w1206_,
		_w4869_
	);
	LUT2 #(
		.INIT('h2)
	) name4096 (
		\g1489_reg/NET0131 ,
		_w4869_,
		_w4870_
	);
	LUT2 #(
		.INIT('h4)
	) name4097 (
		\g1442_reg/NET0131 ,
		_w1206_,
		_w4871_
	);
	LUT2 #(
		.INIT('h1)
	) name4098 (
		_w4870_,
		_w4871_,
		_w4872_
	);
	LUT2 #(
		.INIT('h2)
	) name4099 (
		\g35_pad ,
		_w4872_,
		_w4873_
	);
	LUT2 #(
		.INIT('h8)
	) name4100 (
		\g35_pad ,
		\g4473_reg/NET0131 ,
		_w4874_
	);
	LUT2 #(
		.INIT('h4)
	) name4101 (
		\g35_pad ,
		\g4459_reg/NET0131 ,
		_w4875_
	);
	LUT2 #(
		.INIT('h1)
	) name4102 (
		_w4874_,
		_w4875_,
		_w4876_
	);
	LUT2 #(
		.INIT('h1)
	) name4103 (
		\g35_pad ,
		\g4492_reg/NET0131 ,
		_w4877_
	);
	LUT2 #(
		.INIT('h4)
	) name4104 (
		\g2988_reg/NET0131 ,
		\g35_pad ,
		_w4878_
	);
	LUT2 #(
		.INIT('h4)
	) name4105 (
		_w1052_,
		_w4878_,
		_w4879_
	);
	LUT2 #(
		.INIT('h1)
	) name4106 (
		_w4877_,
		_w4879_,
		_w4880_
	);
	LUT2 #(
		.INIT('h2)
	) name4107 (
		\g35_pad ,
		\g4467_reg/NET0131 ,
		_w4881_
	);
	LUT2 #(
		.INIT('h8)
	) name4108 (
		\g4462_reg/NET0131 ,
		\g4643_reg/NET0131 ,
		_w4882_
	);
	LUT2 #(
		.INIT('h8)
	) name4109 (
		_w4881_,
		_w4882_,
		_w4883_
	);
	LUT2 #(
		.INIT('h2)
	) name4110 (
		\g4473_reg/NET0131 ,
		_w4883_,
		_w4884_
	);
	LUT2 #(
		.INIT('h8)
	) name4111 (
		\g35_pad ,
		\g5092_reg/NET0131 ,
		_w4885_
	);
	LUT2 #(
		.INIT('h1)
	) name4112 (
		\g5084_reg/NET0131 ,
		_w4885_,
		_w4886_
	);
	LUT2 #(
		.INIT('h8)
	) name4113 (
		\g35_pad ,
		_w4169_,
		_w4887_
	);
	LUT2 #(
		.INIT('h1)
	) name4114 (
		_w4886_,
		_w4887_,
		_w4888_
	);
	LUT2 #(
		.INIT('h8)
	) name4115 (
		\g1205_reg/NET0131 ,
		\g35_pad ,
		_w4889_
	);
	LUT2 #(
		.INIT('h1)
	) name4116 (
		\g1087_reg/NET0131 ,
		_w4889_,
		_w4890_
	);
	LUT2 #(
		.INIT('h8)
	) name4117 (
		\g35_pad ,
		_w3390_,
		_w4891_
	);
	LUT2 #(
		.INIT('h1)
	) name4118 (
		_w4890_,
		_w4891_,
		_w4892_
	);
	LUT2 #(
		.INIT('h4)
	) name4119 (
		\g35_pad ,
		\g370_reg/NET0131 ,
		_w4893_
	);
	LUT2 #(
		.INIT('h1)
	) name4120 (
		\g358_reg/NET0131 ,
		\g376_reg/NET0131 ,
		_w4894_
	);
	LUT2 #(
		.INIT('h2)
	) name4121 (
		\g35_pad ,
		_w987_,
		_w4895_
	);
	LUT2 #(
		.INIT('h4)
	) name4122 (
		_w4894_,
		_w4895_,
		_w4896_
	);
	LUT2 #(
		.INIT('h1)
	) name4123 (
		_w4893_,
		_w4896_,
		_w4897_
	);
	LUT2 #(
		.INIT('h8)
	) name4124 (
		\g35_pad ,
		\g4264_reg/NET0131 ,
		_w4898_
	);
	LUT2 #(
		.INIT('h1)
	) name4125 (
		\g4258_reg/NET0131 ,
		_w4898_,
		_w4899_
	);
	LUT2 #(
		.INIT('h8)
	) name4126 (
		\g35_pad ,
		_w4225_,
		_w4900_
	);
	LUT2 #(
		.INIT('h1)
	) name4127 (
		_w4899_,
		_w4900_,
		_w4901_
	);
	LUT2 #(
		.INIT('h2)
	) name4128 (
		\g35_pad ,
		\g890_reg/NET0131 ,
		_w4902_
	);
	LUT2 #(
		.INIT('h1)
	) name4129 (
		\g862_reg/NET0131 ,
		_w4902_,
		_w4903_
	);
	LUT2 #(
		.INIT('h4)
	) name4130 (
		\g890_reg/NET0131 ,
		_w2550_,
		_w4904_
	);
	LUT2 #(
		.INIT('h1)
	) name4131 (
		_w4903_,
		_w4904_,
		_w4905_
	);
	LUT2 #(
		.INIT('h8)
	) name4132 (
		\g1548_reg/NET0131 ,
		\g35_pad ,
		_w4906_
	);
	LUT2 #(
		.INIT('h1)
	) name4133 (
		\g1430_reg/NET0131 ,
		_w4906_,
		_w4907_
	);
	LUT2 #(
		.INIT('h8)
	) name4134 (
		\g35_pad ,
		_w1380_,
		_w4908_
	);
	LUT2 #(
		.INIT('h1)
	) name4135 (
		_w4907_,
		_w4908_,
		_w4909_
	);
	LUT2 #(
		.INIT('h2)
	) name4136 (
		\g35_pad ,
		_w1016_,
		_w4910_
	);
	LUT2 #(
		.INIT('h2)
	) name4137 (
		\g4633_reg/NET0131 ,
		_w4855_,
		_w4911_
	);
	LUT2 #(
		.INIT('h8)
	) name4138 (
		\g3179_reg/NET0131 ,
		\g35_pad ,
		_w4912_
	);
	LUT2 #(
		.INIT('h8)
	) name4139 (
		\g3167_reg/NET0131 ,
		\g3171_reg/NET0131 ,
		_w4913_
	);
	LUT2 #(
		.INIT('h2)
	) name4140 (
		_w4912_,
		_w4913_,
		_w4914_
	);
	LUT2 #(
		.INIT('h4)
	) name4141 (
		\g3167_reg/NET0131 ,
		\g35_pad ,
		_w4915_
	);
	LUT2 #(
		.INIT('h2)
	) name4142 (
		\g3171_reg/NET0131 ,
		_w4912_,
		_w4916_
	);
	LUT2 #(
		.INIT('h4)
	) name4143 (
		_w4915_,
		_w4916_,
		_w4917_
	);
	LUT2 #(
		.INIT('h1)
	) name4144 (
		_w4914_,
		_w4917_,
		_w4918_
	);
	LUT2 #(
		.INIT('h8)
	) name4145 (
		\g18098_pad ,
		\g35_pad ,
		_w4919_
	);
	LUT2 #(
		.INIT('h2)
	) name4146 (
		\g305_reg/NET0131 ,
		\g35_pad ,
		_w4920_
	);
	LUT2 #(
		.INIT('h1)
	) name4147 (
		_w4919_,
		_w4920_,
		_w4921_
	);
	LUT2 #(
		.INIT('h1)
	) name4148 (
		\g2886_reg/NET0131 ,
		\g35_pad ,
		_w4922_
	);
	LUT2 #(
		.INIT('h1)
	) name4149 (
		\g2980_reg/NET0131 ,
		\g34_reg/NET0131 ,
		_w4923_
	);
	LUT2 #(
		.INIT('h8)
	) name4150 (
		\g35_pad ,
		_w4923_,
		_w4924_
	);
	LUT2 #(
		.INIT('h1)
	) name4151 (
		_w4922_,
		_w4924_,
		_w4925_
	);
	LUT2 #(
		.INIT('h8)
	) name4152 (
		\g3161_reg/NET0131 ,
		\g35_pad ,
		_w4926_
	);
	LUT2 #(
		.INIT('h1)
	) name4153 (
		\g3155_reg/NET0131 ,
		_w4926_,
		_w4927_
	);
	LUT2 #(
		.INIT('h8)
	) name4154 (
		\g35_pad ,
		_w4095_,
		_w4928_
	);
	LUT2 #(
		.INIT('h1)
	) name4155 (
		_w4927_,
		_w4928_,
		_w4929_
	);
	LUT2 #(
		.INIT('h2)
	) name4156 (
		\g35_pad ,
		_w3571_,
		_w4930_
	);
	LUT2 #(
		.INIT('h4)
	) name4157 (
		\g35_pad ,
		\g5057_reg/NET0131 ,
		_w4931_
	);
	LUT2 #(
		.INIT('h1)
	) name4158 (
		_w4930_,
		_w4931_,
		_w4932_
	);
	LUT2 #(
		.INIT('h8)
	) name4159 (
		\g35_pad ,
		\g9251_pad ,
		_w4933_
	);
	LUT2 #(
		.INIT('h1)
	) name4160 (
		\g4308_reg/NET0131 ,
		_w4933_,
		_w4934_
	);
	LUT2 #(
		.INIT('h8)
	) name4161 (
		\g4308_reg/NET0131 ,
		_w4933_,
		_w4935_
	);
	LUT2 #(
		.INIT('h1)
	) name4162 (
		_w4934_,
		_w4935_,
		_w4936_
	);
	LUT2 #(
		.INIT('h8)
	) name4163 (
		\g3171_reg/NET0131 ,
		\g35_pad ,
		_w4937_
	);
	LUT2 #(
		.INIT('h1)
	) name4164 (
		\g3167_reg/NET0131 ,
		_w4937_,
		_w4938_
	);
	LUT2 #(
		.INIT('h8)
	) name4165 (
		\g35_pad ,
		_w4913_,
		_w4939_
	);
	LUT2 #(
		.INIT('h1)
	) name4166 (
		_w4938_,
		_w4939_,
		_w4940_
	);
	LUT2 #(
		.INIT('h1)
	) name4167 (
		\g35_pad ,
		\g890_reg/NET0131 ,
		_w4941_
	);
	LUT2 #(
		.INIT('h2)
	) name4168 (
		\g35_pad ,
		\g862_reg/NET0131 ,
		_w4942_
	);
	LUT2 #(
		.INIT('h4)
	) name4169 (
		\g896_reg/NET0131 ,
		_w4942_,
		_w4943_
	);
	LUT2 #(
		.INIT('h1)
	) name4170 (
		_w2554_,
		_w4941_,
		_w4944_
	);
	LUT2 #(
		.INIT('h4)
	) name4171 (
		_w4943_,
		_w4944_,
		_w4945_
	);
	LUT2 #(
		.INIT('h8)
	) name4172 (
		\g35_pad ,
		\g9019_pad ,
		_w4946_
	);
	LUT2 #(
		.INIT('h1)
	) name4173 (
		\g4291_reg/NET0131 ,
		_w4946_,
		_w4947_
	);
	LUT2 #(
		.INIT('h8)
	) name4174 (
		\g4291_reg/NET0131 ,
		_w4946_,
		_w4948_
	);
	LUT2 #(
		.INIT('h1)
	) name4175 (
		_w4947_,
		_w4948_,
		_w4949_
	);
	LUT2 #(
		.INIT('h2)
	) name4176 (
		\g35_pad ,
		_w2517_,
		_w4950_
	);
	LUT2 #(
		.INIT('h2)
	) name4177 (
		\g385_reg/NET0131 ,
		_w4950_,
		_w4951_
	);
	LUT2 #(
		.INIT('h8)
	) name4178 (
		\g35_pad ,
		\g8839_pad ,
		_w4952_
	);
	LUT2 #(
		.INIT('h1)
	) name4179 (
		\g4281_reg/NET0131 ,
		_w4952_,
		_w4953_
	);
	LUT2 #(
		.INIT('h8)
	) name4180 (
		\g4281_reg/NET0131 ,
		_w4952_,
		_w4954_
	);
	LUT2 #(
		.INIT('h1)
	) name4181 (
		_w4953_,
		_w4954_,
		_w4955_
	);
	LUT2 #(
		.INIT('h2)
	) name4182 (
		\g1532_reg/NET0131 ,
		\g7946_pad ,
		_w4956_
	);
	LUT2 #(
		.INIT('h8)
	) name4183 (
		\g1521_reg/NET0131 ,
		\g7946_pad ,
		_w4957_
	);
	LUT2 #(
		.INIT('h1)
	) name4184 (
		_w4956_,
		_w4957_,
		_w4958_
	);
	LUT2 #(
		.INIT('h2)
	) name4185 (
		\g35_pad ,
		_w4958_,
		_w4959_
	);
	LUT2 #(
		.INIT('h2)
	) name4186 (
		\g1306_reg/NET0131 ,
		\g35_pad ,
		_w4960_
	);
	LUT2 #(
		.INIT('h1)
	) name4187 (
		_w4959_,
		_w4960_,
		_w4961_
	);
	LUT2 #(
		.INIT('h2)
	) name4188 (
		\g1178_reg/NET0131 ,
		\g7916_pad ,
		_w4962_
	);
	LUT2 #(
		.INIT('h8)
	) name4189 (
		\g7916_pad ,
		\g996_reg/NET0131 ,
		_w4963_
	);
	LUT2 #(
		.INIT('h1)
	) name4190 (
		_w4962_,
		_w4963_,
		_w4964_
	);
	LUT2 #(
		.INIT('h2)
	) name4191 (
		\g35_pad ,
		_w4964_,
		_w4965_
	);
	LUT2 #(
		.INIT('h2)
	) name4192 (
		\g1183_reg/NET0131 ,
		\g35_pad ,
		_w4966_
	);
	LUT2 #(
		.INIT('h1)
	) name4193 (
		_w4965_,
		_w4966_,
		_w4967_
	);
	LUT2 #(
		.INIT('h2)
	) name4194 (
		\g1189_reg/NET0131 ,
		\g7916_pad ,
		_w4968_
	);
	LUT2 #(
		.INIT('h8)
	) name4195 (
		\g1178_reg/NET0131 ,
		\g7916_pad ,
		_w4969_
	);
	LUT2 #(
		.INIT('h1)
	) name4196 (
		_w4968_,
		_w4969_,
		_w4970_
	);
	LUT2 #(
		.INIT('h2)
	) name4197 (
		\g35_pad ,
		_w4970_,
		_w4971_
	);
	LUT2 #(
		.INIT('h4)
	) name4198 (
		\g35_pad ,
		\g962_reg/NET0131 ,
		_w4972_
	);
	LUT2 #(
		.INIT('h1)
	) name4199 (
		_w4971_,
		_w4972_,
		_w4973_
	);
	LUT2 #(
		.INIT('h1)
	) name4200 (
		\g2724_reg/NET0131 ,
		\g35_pad ,
		_w4974_
	);
	LUT2 #(
		.INIT('h2)
	) name4201 (
		\g2741_reg/NET0131 ,
		\g35_pad ,
		_w4975_
	);
	LUT2 #(
		.INIT('h2)
	) name4202 (
		\g35_pad ,
		_w1206_,
		_w4976_
	);
	LUT2 #(
		.INIT('h2)
	) name4203 (
		\g3155_reg/NET0131 ,
		\g3167_reg/NET0131 ,
		_w4977_
	);
	LUT2 #(
		.INIT('h2)
	) name4204 (
		\g35_pad ,
		_w4977_,
		_w4978_
	);
	LUT2 #(
		.INIT('h2)
	) name4205 (
		\g3161_reg/NET0131 ,
		_w4978_,
		_w4979_
	);
	LUT2 #(
		.INIT('h4)
	) name4206 (
		\g35_pad ,
		\g4239_reg/NET0131 ,
		_w4980_
	);
	LUT2 #(
		.INIT('h4)
	) name4207 (
		\g10122_pad ,
		\g35_pad ,
		_w4981_
	);
	LUT2 #(
		.INIT('h4)
	) name4208 (
		\g4297_reg/NET0131 ,
		_w4981_,
		_w4982_
	);
	LUT2 #(
		.INIT('h1)
	) name4209 (
		_w4980_,
		_w4982_,
		_w4983_
	);
	LUT2 #(
		.INIT('h4)
	) name4210 (
		\g35_pad ,
		\g4462_reg/NET0131 ,
		_w4984_
	);
	LUT2 #(
		.INIT('h4)
	) name4211 (
		\g4473_reg/NET0131 ,
		_w4881_,
		_w4985_
	);
	LUT2 #(
		.INIT('h1)
	) name4212 (
		_w4984_,
		_w4985_,
		_w4986_
	);
	LUT2 #(
		.INIT('h1)
	) name4213 (
		\g35_pad ,
		\g534_reg/NET0131 ,
		_w4987_
	);
	LUT2 #(
		.INIT('h8)
	) name4214 (
		\g29212_pad ,
		\g35_pad ,
		_w4988_
	);
	LUT2 #(
		.INIT('h4)
	) name4215 (
		\g550_reg/NET0131 ,
		_w4988_,
		_w4989_
	);
	LUT2 #(
		.INIT('h1)
	) name4216 (
		_w4987_,
		_w4989_,
		_w4990_
	);
	LUT2 #(
		.INIT('h1)
	) name4217 (
		\g2980_reg/NET0131 ,
		\g35_pad ,
		_w4991_
	);
	LUT2 #(
		.INIT('h4)
	) name4218 (
		\g2984_reg/NET0131 ,
		\g34_reg/NET0131 ,
		_w4992_
	);
	LUT2 #(
		.INIT('h8)
	) name4219 (
		\g35_pad ,
		_w4992_,
		_w4993_
	);
	LUT2 #(
		.INIT('h1)
	) name4220 (
		_w4991_,
		_w4993_,
		_w4994_
	);
	LUT2 #(
		.INIT('h1)
	) name4221 (
		\g35_pad ,
		\g538_reg/NET0131 ,
		_w4995_
	);
	LUT2 #(
		.INIT('h2)
	) name4222 (
		\g35_pad ,
		\g546_reg/NET0131 ,
		_w4996_
	);
	LUT2 #(
		.INIT('h8)
	) name4223 (
		\g691_reg/NET0131 ,
		_w4996_,
		_w4997_
	);
	LUT2 #(
		.INIT('h1)
	) name4224 (
		_w4995_,
		_w4997_,
		_w4998_
	);
	LUT2 #(
		.INIT('h4)
	) name4225 (
		\g218_reg/NET0131 ,
		\g35_pad ,
		_w4999_
	);
	LUT2 #(
		.INIT('h2)
	) name4226 (
		\g209_reg/NET0131 ,
		\g35_pad ,
		_w5000_
	);
	LUT2 #(
		.INIT('h1)
	) name4227 (
		_w4999_,
		_w5000_,
		_w5001_
	);
	LUT2 #(
		.INIT('h8)
	) name4228 (
		\g4146_reg/NET0131 ,
		\g4157_reg/NET0131 ,
		_w5002_
	);
	LUT2 #(
		.INIT('h2)
	) name4229 (
		\g35_pad ,
		_w5002_,
		_w5003_
	);
	LUT2 #(
		.INIT('h4)
	) name4230 (
		\g35_pad ,
		\g4122_reg/NET0131 ,
		_w5004_
	);
	LUT2 #(
		.INIT('h1)
	) name4231 (
		_w5003_,
		_w5004_,
		_w5005_
	);
	LUT2 #(
		.INIT('h1)
	) name4232 (
		\g209_reg/NET0131 ,
		\g538_reg/NET0131 ,
		_w5006_
	);
	LUT2 #(
		.INIT('h2)
	) name4233 (
		\g35_pad ,
		_w5006_,
		_w5007_
	);
	LUT2 #(
		.INIT('h1)
	) name4234 (
		\g4153_reg/NET0131 ,
		\g4172_reg/NET0131 ,
		_w5008_
	);
	LUT2 #(
		.INIT('h2)
	) name4235 (
		\g35_pad ,
		_w5008_,
		_w5009_
	);
	LUT2 #(
		.INIT('h8)
	) name4236 (
		\g4467_reg/NET0131 ,
		\g4473_reg/NET0131 ,
		_w5010_
	);
	LUT2 #(
		.INIT('h2)
	) name4237 (
		\g35_pad ,
		\g4462_reg/NET0131 ,
		_w5011_
	);
	LUT2 #(
		.INIT('h4)
	) name4238 (
		_w5010_,
		_w5011_,
		_w5012_
	);
	LUT2 #(
		.INIT('h4)
	) name4239 (
		\g3155_reg/NET0131 ,
		_w4915_,
		_w5013_
	);
	LUT2 #(
		.INIT('h1)
	) name4240 (
		\g2715_reg/NET0131 ,
		\g35_pad ,
		_w5014_
	);
	LUT2 #(
		.INIT('h4)
	) name4241 (
		\g4639_reg/NET0131 ,
		_w4453_,
		_w5015_
	);
	LUT2 #(
		.INIT('h4)
	) name4242 (
		\g358_reg/NET0131 ,
		\g35_pad ,
		_w5016_
	);
	LUT2 #(
		.INIT('h4)
	) name4243 (
		\g8719_pad ,
		_w5016_,
		_w5017_
	);
	LUT2 #(
		.INIT('h1)
	) name4244 (
		_w4881_,
		_w5011_,
		_w5018_
	);
	LUT2 #(
		.INIT('h2)
	) name4245 (
		\g3050_reg/NET0131 ,
		\g35_pad ,
		_w5019_
	);
	LUT2 #(
		.INIT('h1)
	) name4246 (
		_w3589_,
		_w5019_,
		_w5020_
	);
	LUT2 #(
		.INIT('h4)
	) name4247 (
		\g35_pad ,
		\g4483_reg/NET0131 ,
		_w5021_
	);
	LUT2 #(
		.INIT('h1)
	) name4248 (
		_w1048_,
		_w5021_,
		_w5022_
	);
	LUT2 #(
		.INIT('h4)
	) name4249 (
		\g35_pad ,
		\g4486_reg/NET0131 ,
		_w5023_
	);
	LUT2 #(
		.INIT('h1)
	) name4250 (
		_w1045_,
		_w5023_,
		_w5024_
	);
	LUT2 #(
		.INIT('h4)
	) name4251 (
		\g35_pad ,
		\g4489_reg/NET0131 ,
		_w5025_
	);
	LUT2 #(
		.INIT('h1)
	) name4252 (
		_w1042_,
		_w5025_,
		_w5026_
	);
	LUT2 #(
		.INIT('h2)
	) name4253 (
		\g35_pad ,
		\g4239_reg/NET0131 ,
		_w5027_
	);
	LUT2 #(
		.INIT('h4)
	) name4254 (
		\g35_pad ,
		\g4273_reg/NET0131 ,
		_w5028_
	);
	LUT2 #(
		.INIT('h1)
	) name4255 (
		_w5027_,
		_w5028_,
		_w5029_
	);
	LUT2 #(
		.INIT('h2)
	) name4256 (
		\g2735_reg/NET0131 ,
		\g35_pad ,
		_w5030_
	);
	LUT2 #(
		.INIT('h4)
	) name4257 (
		\g35_pad ,
		\g4382_reg/NET0131 ,
		_w5031_
	);
	LUT2 #(
		.INIT('h2)
	) name4258 (
		\g2719_reg/NET0131 ,
		\g35_pad ,
		_w5032_
	);
	LUT2 #(
		.INIT('h4)
	) name4259 (
		\g35_pad ,
		\g4392_reg/NET0131 ,
		_w5033_
	);
	LUT2 #(
		.INIT('h4)
	) name4260 (
		\g35_pad ,
		\g4153_reg/NET0131 ,
		_w5034_
	);
	LUT2 #(
		.INIT('h2)
	) name4261 (
		\g2975_reg/NET0131 ,
		\g35_pad ,
		_w5035_
	);
	LUT2 #(
		.INIT('h4)
	) name4262 (
		\g35_pad ,
		\g4104_reg/NET0131 ,
		_w5036_
	);
	LUT2 #(
		.INIT('h4)
	) name4263 (
		\g35_pad ,
		\g4087_reg/NET0131 ,
		_w5037_
	);
	LUT2 #(
		.INIT('h4)
	) name4264 (
		\g35_pad ,
		\g4057_reg/NET0131 ,
		_w5038_
	);
	LUT2 #(
		.INIT('h4)
	) name4265 (
		\g35_pad ,
		\g4076_reg/NET0131 ,
		_w5039_
	);
	LUT2 #(
		.INIT('h4)
	) name4266 (
		\g35_pad ,
		\g4064_reg/NET0131 ,
		_w5040_
	);
	LUT2 #(
		.INIT('h4)
	) name4267 (
		\g35_pad ,
		\g753_reg/NET0131 ,
		_w5041_
	);
	LUT2 #(
		.INIT('h1)
	) name4268 (
		\g2759_reg/NET0131 ,
		\g35_pad ,
		_w5042_
	);
	LUT2 #(
		.INIT('h1)
	) name4269 (
		\g35_pad ,
		\g4108_reg/NET0131 ,
		_w5043_
	);
	LUT2 #(
		.INIT('h1)
	) name4270 (
		\g2756_reg/NET0131 ,
		\g35_pad ,
		_w5044_
	);
	LUT2 #(
		.INIT('h1)
	) name4271 (
		\g2917_reg/NET0131 ,
		\g35_pad ,
		_w5045_
	);
	LUT2 #(
		.INIT('h8)
	) name4272 (
		\g18099_pad ,
		\g35_pad ,
		_w5046_
	);
	LUT2 #(
		.INIT('h1)
	) name4273 (
		\g2882_reg/NET0131 ,
		\g35_pad ,
		_w5047_
	);
	LUT2 #(
		.INIT('h1)
	) name4274 (
		\g35_pad ,
		\g4141_reg/NET0131 ,
		_w5048_
	);
	LUT2 #(
		.INIT('h1)
	) name4275 (
		\g35_pad ,
		\g4082_reg/NET0131 ,
		_w5049_
	);
	LUT2 #(
		.INIT('h8)
	) name4276 (
		\g29216_pad ,
		\g35_pad ,
		_w5050_
	);
	LUT2 #(
		.INIT('h1)
	) name4277 (
		\g2955_reg/NET0131 ,
		\g35_pad ,
		_w5051_
	);
	LUT2 #(
		.INIT('h1)
	) name4278 (
		\g35_pad ,
		\g4098_reg/NET0131 ,
		_w5052_
	);
	LUT2 #(
		.INIT('h1)
	) name4279 (
		\g35_pad ,
		\g4093_reg/NET0131 ,
		_w5053_
	);
	LUT2 #(
		.INIT('h1)
	) name4280 (
		\g2873_reg/NET0131 ,
		\g35_pad ,
		_w5054_
	);
	LUT2 #(
		.INIT('h1)
	) name4281 (
		\g2729_reg/NET0131 ,
		\g35_pad ,
		_w5055_
	);
	LUT2 #(
		.INIT('h2)
	) name4282 (
		\g2495_reg/NET0131 ,
		_w1432_,
		_w5056_
	);
	LUT2 #(
		.INIT('h1)
	) name4283 (
		\g2421_reg/NET0131 ,
		_w1657_,
		_w5057_
	);
	LUT2 #(
		.INIT('h2)
	) name4284 (
		\g35_pad ,
		_w5056_,
		_w5058_
	);
	LUT2 #(
		.INIT('h4)
	) name4285 (
		_w5057_,
		_w5058_,
		_w5059_
	);
	LUT2 #(
		.INIT('h2)
	) name4286 (
		\g2361_reg/NET0131 ,
		_w1415_,
		_w5060_
	);
	LUT2 #(
		.INIT('h1)
	) name4287 (
		\g2287_reg/NET0131 ,
		_w1606_,
		_w5061_
	);
	LUT2 #(
		.INIT('h2)
	) name4288 (
		\g35_pad ,
		_w5060_,
		_w5062_
	);
	LUT2 #(
		.INIT('h4)
	) name4289 (
		_w5061_,
		_w5062_,
		_w5063_
	);
	LUT2 #(
		.INIT('h1)
	) name4290 (
		\g2555_reg/NET0131 ,
		_w1703_,
		_w5064_
	);
	LUT2 #(
		.INIT('h2)
	) name4291 (
		\g35_pad ,
		_w1726_,
		_w5065_
	);
	LUT2 #(
		.INIT('h4)
	) name4292 (
		_w5064_,
		_w5065_,
		_w5066_
	);
	LUT2 #(
		.INIT('h2)
	) name4293 (
		\g1936_reg/NET0131 ,
		_w1516_,
		_w5067_
	);
	LUT2 #(
		.INIT('h1)
	) name4294 (
		\g1862_reg/NET0131 ,
		_w1855_,
		_w5068_
	);
	LUT2 #(
		.INIT('h2)
	) name4295 (
		\g35_pad ,
		_w5067_,
		_w5069_
	);
	LUT2 #(
		.INIT('h4)
	) name4296 (
		_w5068_,
		_w5069_,
		_w5070_
	);
	LUT2 #(
		.INIT('h2)
	) name4297 (
		\g2070_reg/NET0131 ,
		_w1533_,
		_w5071_
	);
	LUT2 #(
		.INIT('h1)
	) name4298 (
		\g1996_reg/NET0131 ,
		_w1938_,
		_w5072_
	);
	LUT2 #(
		.INIT('h2)
	) name4299 (
		\g35_pad ,
		_w5071_,
		_w5073_
	);
	LUT2 #(
		.INIT('h4)
	) name4300 (
		_w5072_,
		_w5073_,
		_w5074_
	);
	LUT2 #(
		.INIT('h8)
	) name4301 (
		\g1682_reg/NET0131 ,
		_w4277_,
		_w5075_
	);
	LUT2 #(
		.INIT('h2)
	) name4302 (
		\g1668_reg/NET0131 ,
		\g35_pad ,
		_w5076_
	);
	LUT2 #(
		.INIT('h2)
	) name4303 (
		\g1682_reg/NET0131 ,
		_w1959_,
		_w5077_
	);
	LUT2 #(
		.INIT('h4)
	) name4304 (
		\g1246_reg/NET0131 ,
		_w1946_,
		_w5078_
	);
	LUT2 #(
		.INIT('h4)
	) name4305 (
		_w5077_,
		_w5078_,
		_w5079_
	);
	LUT2 #(
		.INIT('h2)
	) name4306 (
		_w5077_,
		_w5078_,
		_w5080_
	);
	LUT2 #(
		.INIT('h2)
	) name4307 (
		\g35_pad ,
		_w1950_,
		_w5081_
	);
	LUT2 #(
		.INIT('h1)
	) name4308 (
		_w5079_,
		_w5080_,
		_w5082_
	);
	LUT2 #(
		.INIT('h8)
	) name4309 (
		_w5081_,
		_w5082_,
		_w5083_
	);
	LUT2 #(
		.INIT('h1)
	) name4310 (
		_w5075_,
		_w5076_,
		_w5084_
	);
	LUT2 #(
		.INIT('h4)
	) name4311 (
		_w5083_,
		_w5084_,
		_w5085_
	);
	LUT2 #(
		.INIT('h2)
	) name4312 (
		\g1802_reg/NET0131 ,
		_w1499_,
		_w5086_
	);
	LUT2 #(
		.INIT('h1)
	) name4313 (
		\g1728_reg/NET0131 ,
		_w1809_,
		_w5087_
	);
	LUT2 #(
		.INIT('h2)
	) name4314 (
		\g35_pad ,
		_w5086_,
		_w5088_
	);
	LUT2 #(
		.INIT('h4)
	) name4315 (
		_w5087_,
		_w5088_,
		_w5089_
	);
	LUT2 #(
		.INIT('h8)
	) name4316 (
		\g3457_reg/NET0131 ,
		_w2445_,
		_w5090_
	);
	LUT2 #(
		.INIT('h2)
	) name4317 (
		\g3457_reg/NET0131 ,
		_w4177_,
		_w5091_
	);
	LUT2 #(
		.INIT('h2)
	) name4318 (
		_w2253_,
		_w5091_,
		_w5092_
	);
	LUT2 #(
		.INIT('h4)
	) name4319 (
		_w2253_,
		_w5091_,
		_w5093_
	);
	LUT2 #(
		.INIT('h2)
	) name4320 (
		_w2448_,
		_w5092_,
		_w5094_
	);
	LUT2 #(
		.INIT('h4)
	) name4321 (
		_w5093_,
		_w5094_,
		_w5095_
	);
	LUT2 #(
		.INIT('h1)
	) name4322 (
		_w886_,
		_w5090_,
		_w5096_
	);
	LUT2 #(
		.INIT('h4)
	) name4323 (
		_w5095_,
		_w5096_,
		_w5097_
	);
	LUT2 #(
		.INIT('h8)
	) name4324 (
		\g3106_reg/NET0131 ,
		_w2328_,
		_w5098_
	);
	LUT2 #(
		.INIT('h8)
	) name4325 (
		\g3352_reg/NET0131 ,
		_w3992_,
		_w5099_
	);
	LUT2 #(
		.INIT('h2)
	) name4326 (
		\g3106_reg/NET0131 ,
		_w5099_,
		_w5100_
	);
	LUT2 #(
		.INIT('h2)
	) name4327 (
		_w2235_,
		_w5100_,
		_w5101_
	);
	LUT2 #(
		.INIT('h4)
	) name4328 (
		_w2235_,
		_w5100_,
		_w5102_
	);
	LUT2 #(
		.INIT('h2)
	) name4329 (
		_w2332_,
		_w5101_,
		_w5103_
	);
	LUT2 #(
		.INIT('h4)
	) name4330 (
		_w5102_,
		_w5103_,
		_w5104_
	);
	LUT2 #(
		.INIT('h1)
	) name4331 (
		_w886_,
		_w5098_,
		_w5105_
	);
	LUT2 #(
		.INIT('h4)
	) name4332 (
		_w5104_,
		_w5105_,
		_w5106_
	);
	LUT2 #(
		.INIT('h2)
	) name4333 (
		\g35_pad ,
		_w3900_,
		_w5107_
	);
	LUT2 #(
		.INIT('h2)
	) name4334 (
		\g1171_reg/NET0131 ,
		_w5107_,
		_w5108_
	);
	LUT2 #(
		.INIT('h4)
	) name4335 (
		\g1171_reg/NET0131 ,
		_w3550_,
		_w5109_
	);
	LUT2 #(
		.INIT('h1)
	) name4336 (
		\g1183_reg/NET0131 ,
		_w3538_,
		_w5110_
	);
	LUT2 #(
		.INIT('h1)
	) name4337 (
		_w4810_,
		_w5110_,
		_w5111_
	);
	LUT2 #(
		.INIT('h1)
	) name4338 (
		_w5109_,
		_w5111_,
		_w5112_
	);
	LUT2 #(
		.INIT('h2)
	) name4339 (
		\g35_pad ,
		_w5112_,
		_w5113_
	);
	LUT2 #(
		.INIT('h1)
	) name4340 (
		_w5108_,
		_w5113_,
		_w5114_
	);
	LUT2 #(
		.INIT('h8)
	) name4341 (
		\g5115_reg/NET0131 ,
		_w2587_,
		_w5115_
	);
	LUT2 #(
		.INIT('h2)
	) name4342 (
		\g5115_reg/NET0131 ,
		_w3965_,
		_w5116_
	);
	LUT2 #(
		.INIT('h4)
	) name4343 (
		\g5297_reg/NET0131 ,
		_w912_,
		_w5117_
	);
	LUT2 #(
		.INIT('h8)
	) name4344 (
		\g5297_reg/NET0131 ,
		_w925_,
		_w5118_
	);
	LUT2 #(
		.INIT('h2)
	) name4345 (
		\g5357_reg/NET0131 ,
		_w5117_,
		_w5119_
	);
	LUT2 #(
		.INIT('h4)
	) name4346 (
		_w5118_,
		_w5119_,
		_w5120_
	);
	LUT2 #(
		.INIT('h4)
	) name4347 (
		\g5297_reg/NET0131 ,
		_w941_,
		_w5121_
	);
	LUT2 #(
		.INIT('h8)
	) name4348 (
		\g5297_reg/NET0131 ,
		_w955_,
		_w5122_
	);
	LUT2 #(
		.INIT('h1)
	) name4349 (
		\g5357_reg/NET0131 ,
		_w5121_,
		_w5123_
	);
	LUT2 #(
		.INIT('h4)
	) name4350 (
		_w5122_,
		_w5123_,
		_w5124_
	);
	LUT2 #(
		.INIT('h1)
	) name4351 (
		_w5120_,
		_w5124_,
		_w5125_
	);
	LUT2 #(
		.INIT('h2)
	) name4352 (
		_w5116_,
		_w5125_,
		_w5126_
	);
	LUT2 #(
		.INIT('h4)
	) name4353 (
		_w5116_,
		_w5125_,
		_w5127_
	);
	LUT2 #(
		.INIT('h2)
	) name4354 (
		_w2590_,
		_w5126_,
		_w5128_
	);
	LUT2 #(
		.INIT('h4)
	) name4355 (
		_w5127_,
		_w5128_,
		_w5129_
	);
	LUT2 #(
		.INIT('h1)
	) name4356 (
		_w886_,
		_w5115_,
		_w5130_
	);
	LUT2 #(
		.INIT('h4)
	) name4357 (
		_w5129_,
		_w5130_,
		_w5131_
	);
	LUT2 #(
		.INIT('h2)
	) name4358 (
		\g2227_reg/NET0131 ,
		_w1398_,
		_w5132_
	);
	LUT2 #(
		.INIT('h1)
	) name4359 (
		\g2153_reg/NET0131 ,
		_w1560_,
		_w5133_
	);
	LUT2 #(
		.INIT('h2)
	) name4360 (
		\g35_pad ,
		_w5132_,
		_w5134_
	);
	LUT2 #(
		.INIT('h4)
	) name4361 (
		_w5133_,
		_w5134_,
		_w5135_
	);
	LUT2 #(
		.INIT('h4)
	) name4362 (
		\g35_pad ,
		\g4572_reg/NET0131 ,
		_w5136_
	);
	LUT2 #(
		.INIT('h8)
	) name4363 (
		\g3684_reg/NET0131 ,
		\g4681_reg/NET0131 ,
		_w5137_
	);
	LUT2 #(
		.INIT('h4)
	) name4364 (
		\g4035_reg/NET0131 ,
		\g4688_reg/NET0131 ,
		_w5138_
	);
	LUT2 #(
		.INIT('h8)
	) name4365 (
		\g29220_pad ,
		\g4646_reg/NET0131 ,
		_w5139_
	);
	LUT2 #(
		.INIT('h4)
	) name4366 (
		\g3333_reg/NET0131 ,
		\g4674_reg/NET0131 ,
		_w5140_
	);
	LUT2 #(
		.INIT('h1)
	) name4367 (
		\g4776_reg/NET0131 ,
		\g4793_reg/NET0131 ,
		_w5141_
	);
	LUT2 #(
		.INIT('h4)
	) name4368 (
		\g4801_reg/NET0131 ,
		_w5141_,
		_w5142_
	);
	LUT2 #(
		.INIT('h4)
	) name4369 (
		_w861_,
		_w5142_,
		_w5143_
	);
	LUT2 #(
		.INIT('h4)
	) name4370 (
		\g4776_reg/NET0131 ,
		\g4793_reg/NET0131 ,
		_w5144_
	);
	LUT2 #(
		.INIT('h1)
	) name4371 (
		_w864_,
		_w5144_,
		_w5145_
	);
	LUT2 #(
		.INIT('h1)
	) name4372 (
		_w862_,
		_w888_,
		_w5146_
	);
	LUT2 #(
		.INIT('h1)
	) name4373 (
		_w2223_,
		_w2241_,
		_w5147_
	);
	LUT2 #(
		.INIT('h8)
	) name4374 (
		_w5146_,
		_w5147_,
		_w5148_
	);
	LUT2 #(
		.INIT('h1)
	) name4375 (
		_w5145_,
		_w5148_,
		_w5149_
	);
	LUT2 #(
		.INIT('h1)
	) name4376 (
		_w2330_,
		_w5143_,
		_w5150_
	);
	LUT2 #(
		.INIT('h4)
	) name4377 (
		_w5149_,
		_w5150_,
		_w5151_
	);
	LUT2 #(
		.INIT('h4)
	) name4378 (
		\g4688_reg/NET0131 ,
		_w4759_,
		_w5152_
	);
	LUT2 #(
		.INIT('h4)
	) name4379 (
		_w5151_,
		_w5152_,
		_w5153_
	);
	LUT2 #(
		.INIT('h1)
	) name4380 (
		_w5137_,
		_w5138_,
		_w5154_
	);
	LUT2 #(
		.INIT('h1)
	) name4381 (
		_w5139_,
		_w5140_,
		_w5155_
	);
	LUT2 #(
		.INIT('h8)
	) name4382 (
		_w5154_,
		_w5155_,
		_w5156_
	);
	LUT2 #(
		.INIT('h4)
	) name4383 (
		_w5153_,
		_w5156_,
		_w5157_
	);
	LUT2 #(
		.INIT('h2)
	) name4384 (
		\g35_pad ,
		_w5157_,
		_w5158_
	);
	LUT2 #(
		.INIT('h1)
	) name4385 (
		_w5136_,
		_w5158_,
		_w5159_
	);
	LUT2 #(
		.INIT('h8)
	) name4386 (
		\g691_reg/NET0131 ,
		_w4777_,
		_w5160_
	);
	LUT2 #(
		.INIT('h2)
	) name4387 (
		\g29212_pad ,
		\g35_pad ,
		_w5161_
	);
	LUT2 #(
		.INIT('h8)
	) name4388 (
		\g691_reg/NET0131 ,
		\g703_reg/NET0131 ,
		_w5162_
	);
	LUT2 #(
		.INIT('h4)
	) name4389 (
		\g714_reg/NET0131 ,
		_w5162_,
		_w5163_
	);
	LUT2 #(
		.INIT('h1)
	) name4390 (
		_w3517_,
		_w5163_,
		_w5164_
	);
	LUT2 #(
		.INIT('h8)
	) name4391 (
		\g35_pad ,
		_w3371_,
		_w5165_
	);
	LUT2 #(
		.INIT('h4)
	) name4392 (
		_w5164_,
		_w5165_,
		_w5166_
	);
	LUT2 #(
		.INIT('h1)
	) name4393 (
		_w5160_,
		_w5161_,
		_w5167_
	);
	LUT2 #(
		.INIT('h4)
	) name4394 (
		_w5166_,
		_w5167_,
		_w5168_
	);
	LUT2 #(
		.INIT('h1)
	) name4395 (
		\g29220_pad ,
		_w869_,
		_w5169_
	);
	LUT2 #(
		.INIT('h8)
	) name4396 (
		_w869_,
		_w5125_,
		_w5170_
	);
	LUT2 #(
		.INIT('h2)
	) name4397 (
		\g35_pad ,
		_w5169_,
		_w5171_
	);
	LUT2 #(
		.INIT('h4)
	) name4398 (
		_w5170_,
		_w5171_,
		_w5172_
	);
	LUT2 #(
		.INIT('h1)
	) name4399 (
		_w2221_,
		_w5172_,
		_w5173_
	);
	LUT2 #(
		.INIT('h2)
	) name4400 (
		\g301_reg/NET0131 ,
		\g35_pad ,
		_w5174_
	);
	LUT2 #(
		.INIT('h8)
	) name4401 (
		\g142_reg/NET0131 ,
		\g35_pad ,
		_w5175_
	);
	LUT2 #(
		.INIT('h8)
	) name4402 (
		_w2049_,
		_w5175_,
		_w5176_
	);
	LUT2 #(
		.INIT('h1)
	) name4403 (
		_w5174_,
		_w5176_,
		_w5177_
	);
	assign \g136_reg/P0001  = \g29221_pad ;
	assign \g21727_pad  = _w774_ ;
	assign \g23190_pad  = 1'b0;
	assign \g26875_pad  = _w782_ ;
	assign \g26876_pad  = _w798_ ;
	assign \g26877_pad  = _w814_ ;
	assign \g28041_pad  = _w820_ ;
	assign \g28042_pad  = _w822_ ;
	assign \g30327_pad  = \g37_reg/NET0131 ;
	assign \g30330_pad  = \g2834_reg/NET0131 ;
	assign \g30331_pad  = \g2831_reg/NET0131 ;
	assign \g31793_pad  = _w826_ ;
	assign \g31860_pad  = _w827_ ;
	assign \g31862_pad  = _w828_ ;
	assign \g31863_pad  = _w829_ ;
	assign \g32185_pad  = _w842_ ;
	assign \g33079_pad  = _w851_ ;
	assign \g33435_pad  = _w860_ ;
	assign \g33959_pad  = _w869_ ;
	assign \g34435_pad  = _w877_ ;
	assign \g34788_pad  = _w881_ ;
	assign \g34956_pad  = _w885_ ;
	assign \g34_reg/P0001  = \g34_reg/NET0131 ;
	assign \g35_syn_2  = \g35_pad ;
	assign \g37/_0_  = _w965_ ;
	assign \g41/_0_  = _w1006_ ;
	assign \g60853/_3_  = _w1025_ ;
	assign \g60856/_3_  = _w1030_ ;
	assign \g60879/_3_  = _w1034_ ;
	assign \g60882/_0_  = _w1040_ ;
	assign \g60888/_0_  = _w1043_ ;
	assign \g60891/_0_  = _w1046_ ;
	assign \g60896/_0_  = _w1049_ ;
	assign \g60899/_0_  = _w1071_ ;
	assign \g60900/_3_  = _w1077_ ;
	assign \g60909/_3_  = _w1084_ ;
	assign \g60911/_0_  = _w1088_ ;
	assign \g60915/_0_  = _w1091_ ;
	assign \g60918/_0_  = _w1115_ ;
	assign \g60919/_0_  = _w1137_ ;
	assign \g60928/_0_  = _w1142_ ;
	assign \g60929/_0_  = _w1144_ ;
	assign \g60936/_0_  = _w1148_ ;
	assign \g60937/_0_  = _w1158_ ;
	assign \g60939/_0_  = _w1168_ ;
	assign \g60940/_0_  = _w1182_ ;
	assign \g60941/_0_  = _w1193_ ;
	assign \g60942/_0_  = _w1205_ ;
	assign \g60943/_0_  = _w1216_ ;
	assign \g60944/_0_  = _w1218_ ;
	assign \g60952/_0_  = _w1226_ ;
	assign \g60954/_0_  = _w1233_ ;
	assign \g60958/_0_  = _w1237_ ;
	assign \g60962/_3_  = _w1243_ ;
	assign \g60972/_0_  = _w1253_ ;
	assign \g60980/_0_  = _w1260_ ;
	assign \g60984/_0_  = _w1265_ ;
	assign \g60986/_0_  = _w1266_ ;
	assign \g60989/_0_  = _w1281_ ;
	assign \g60991/_3_  = _w1285_ ;
	assign \g61006/_0_  = _w1289_ ;
	assign \g61008/_0_  = _w1304_ ;
	assign \g61013/_0_  = _w1318_ ;
	assign \g61014/_0_  = _w1330_ ;
	assign \g61015/_0_  = _w1342_ ;
	assign \g61016/_0_  = _w1354_ ;
	assign \g61017/_0_  = _w1355_ ;
	assign \g61026/_3_  = _w1360_ ;
	assign \g61027/_3_  = _w1362_ ;
	assign \g61030/_0_  = _w1367_ ;
	assign \g61031/_0_  = _w1371_ ;
	assign \g61037/_0_  = _w1379_ ;
	assign \g61038/_0_  = _w1387_ ;
	assign \g61042/_0_  = _w1411_ ;
	assign \g61044/_0_  = _w1428_ ;
	assign \g61045/_0_  = _w1445_ ;
	assign \g61046/_0_  = _w1462_ ;
	assign \g61050/_0_  = _w1464_ ;
	assign \g61051/_0_  = _w1468_ ;
	assign \g61052/_0_  = _w1472_ ;
	assign \g61078/_0_  = _w1473_ ;
	assign \g61131/_0_  = _w1474_ ;
	assign \g61137/_3_  = _w1481_ ;
	assign \g61142/_3_  = _w1485_ ;
	assign \g61143/_3_  = _w1489_ ;
	assign \g61151/_0_  = _w1512_ ;
	assign \g61152/_0_  = _w1529_ ;
	assign \g61161/_0_  = _w1546_ ;
	assign \g61168/_3_  = _w1551_ ;
	assign \g61169/_3_  = _w1558_ ;
	assign \g61170/_0_  = _w1567_ ;
	assign \g61171/_3_  = _w1574_ ;
	assign \g61172/_0_  = _w1582_ ;
	assign \g61173/_0_  = _w1590_ ;
	assign \g61174/_0_  = _w1597_ ;
	assign \g61175/_0_  = _w1604_ ;
	assign \g61176/_0_  = _w1613_ ;
	assign \g61177/_3_  = _w1620_ ;
	assign \g61178/_0_  = _w1628_ ;
	assign \g61179/_0_  = _w1636_ ;
	assign \g61180/_0_  = _w1643_ ;
	assign \g61181/_0_  = _w1650_ ;
	assign \g61182/_3_  = _w1655_ ;
	assign \g61183/_0_  = _w1664_ ;
	assign \g61184/_3_  = _w1671_ ;
	assign \g61185/_0_  = _w1679_ ;
	assign \g61186/_0_  = _w1687_ ;
	assign \g61187/_0_  = _w1694_ ;
	assign \g61188/_0_  = _w1701_ ;
	assign \g61189/_0_  = _w1710_ ;
	assign \g61190/_3_  = _w1717_ ;
	assign \g61191/_0_  = _w1725_ ;
	assign \g61192/_0_  = _w1733_ ;
	assign \g61193/_0_  = _w1740_ ;
	assign \g61194/_0_  = _w1747_ ;
	assign \g61221/_0_  = _w1748_ ;
	assign \g61222/_0_  = _w1757_ ;
	assign \g61223/_3_  = _w1763_ ;
	assign \g61224/_3_  = _w1766_ ;
	assign \g61261/_0_  = _w1767_ ;
	assign \g61295/_3_  = _w1775_ ;
	assign \g61308/_0_  = _w1780_ ;
	assign \g61316/_0_  = _w1783_ ;
	assign \g61327/_0_  = _w1786_ ;
	assign \g61329/_0_  = _w1805_ ;
	assign \g61330/_0_  = _w1807_ ;
	assign \g61331/_0_  = _w1816_ ;
	assign \g61332/_3_  = _w1823_ ;
	assign \g61333/_0_  = _w1831_ ;
	assign \g61334/_0_  = _w1839_ ;
	assign \g61335/_0_  = _w1846_ ;
	assign \g61336/_0_  = _w1853_ ;
	assign \g61337/_0_  = _w1862_ ;
	assign \g61338/_3_  = _w1869_ ;
	assign \g61339/_0_  = _w1877_ ;
	assign \g61340/_0_  = _w1885_ ;
	assign \g61341/_0_  = _w1892_ ;
	assign \g61342/_0_  = _w1899_ ;
	assign \g61343/_0_  = _w1908_ ;
	assign \g61344/_3_  = _w1915_ ;
	assign \g61345/_0_  = _w1923_ ;
	assign \g61346/_0_  = _w1930_ ;
	assign \g61347/_0_  = _w1937_ ;
	assign \g61348/_0_  = _w1945_ ;
	assign \g61349/_0_  = _w1958_ ;
	assign \g61350/_3_  = _w1966_ ;
	assign \g61351/_0_  = _w1974_ ;
	assign \g61352/_0_  = _w1981_ ;
	assign \g61353/_0_  = _w1988_ ;
	assign \g61354/_0_  = _w1995_ ;
	assign \g61367/_0_  = _w2001_ ;
	assign \g61372/_0_  = _w2004_ ;
	assign \g61373/_0_  = _w2027_ ;
	assign \g61375/_0_  = _w2057_ ;
	assign \g61382/_0_  = _w2058_ ;
	assign \g61385/_3_  = _w2064_ ;
	assign \g61386/_0_  = _w2075_ ;
	assign \g61399/_0_  = _w2077_ ;
	assign \g61400/_0_  = _w2086_ ;
	assign \g61402/_0_  = _w2088_ ;
	assign \g61405/_0_  = _w2089_ ;
	assign \g61435/_3_  = _w2097_ ;
	assign \g61449/_0_  = _w2116_ ;
	assign \g61468/_0_  = _w2124_ ;
	assign \g61475/_0_  = _w2129_ ;
	assign \g61480/_0_  = _w2132_ ;
	assign \g61482/_0_  = _w2141_ ;
	assign \g61483/_0_  = _w2156_ ;
	assign \g61484/_0_  = _w2175_ ;
	assign \g61486/_3_  = _w2184_ ;
	assign \g61494/_0_  = _w2187_ ;
	assign \g61496/_0_  = _w2194_ ;
	assign \g61497/_0_  = _w2200_ ;
	assign \g61514/_0_  = _w2204_ ;
	assign \g61517/_0_  = _w2220_ ;
	assign \g61519/_3_  = _w2239_ ;
	assign \g61520/_3_  = _w2257_ ;
	assign \g61527/_0_  = _w2259_ ;
	assign \g61541/_0_  = _w2266_ ;
	assign \g61544/_0_  = _w2273_ ;
	assign \g61550/_0_  = _w2275_ ;
	assign \g61551/_0_  = _w2278_ ;
	assign \g61554/_0_  = _w2282_ ;
	assign \g61556/_3_  = _w2287_ ;
	assign \g61567/_0_  = _w2299_ ;
	assign \g61571/_0_  = _w2305_ ;
	assign \g61574/_0_  = _w2311_ ;
	assign \g61587/_0_  = _w2316_ ;
	assign \g61592/_0_  = _w2320_ ;
	assign \g61632/_0_  = _w2327_ ;
	assign \g61634/_0_  = _w2342_ ;
	assign \g61635/_0_  = _w2354_ ;
	assign \g61639/_0_  = _w2367_ ;
	assign \g61644/_0_  = _w2372_ ;
	assign \g61652/_3_  = _w2393_ ;
	assign \g61709/_0_  = _w2402_ ;
	assign \g61714/_0_  = _w2409_ ;
	assign \g61720/_0_  = _w2415_ ;
	assign \g61721/_0_  = _w2423_ ;
	assign \g61723/_0_  = _w2430_ ;
	assign \g61725/_0_  = _w2437_ ;
	assign \g61726/_0_  = _w2444_ ;
	assign \g61734/_0_  = _w2458_ ;
	assign \g61739/_0_  = _w2483_ ;
	assign \g61744/_0_  = _w2488_ ;
	assign \g61746/_3_  = _w2491_ ;
	assign \g61747/_3_  = _w2495_ ;
	assign \g61748/_3_  = _w2498_ ;
	assign \g61750/u3_syn_7  = _w2492_ ;
	assign \g61802/_0_  = _w2516_ ;
	assign \g61804/_0_  = _w2556_ ;
	assign \g61808/_0_  = _w2570_ ;
	assign \g61811/_0_  = _w2586_ ;
	assign \g61816/_0_  = _w2600_ ;
	assign \g61818/_0_  = _w2613_ ;
	assign \g61820/_0_  = _w2624_ ;
	assign \g61823/_0_  = _w2629_ ;
	assign \g61824/_0_  = _w2636_ ;
	assign \g61841/_0_  = _w2641_ ;
	assign \g61842/_3_  = _w2644_ ;
	assign \g61844/_3_  = _w2659_ ;
	assign \g61845/_3_  = _w2667_ ;
	assign \g61846/_3_  = _w2678_ ;
	assign \g61847/u3_syn_7  = _w2679_ ;
	assign \g61848/_0_  = _w2688_ ;
	assign \g61849/_3_  = _w2696_ ;
	assign \g61850/_0_  = _w2705_ ;
	assign \g61851/u3_syn_7  = _w2706_ ;
	assign \g61852/_0_  = _w2716_ ;
	assign \g61853/_3_  = _w2727_ ;
	assign \g61854/_3_  = _w2734_ ;
	assign \g61855/_0_  = _w2743_ ;
	assign \g61856/u3_syn_7  = _w2744_ ;
	assign \g61857/_0_  = _w2751_ ;
	assign \g61858/_3_  = _w2762_ ;
	assign \g61859/_3_  = _w2769_ ;
	assign \g61860/u3_syn_7  = _w2770_ ;
	assign \g61861/_0_  = _w2779_ ;
	assign \g61862/_3_  = _w2793_ ;
	assign \g61863/_3_  = _w2801_ ;
	assign \g61864/u3_syn_7  = _w2802_ ;
	assign \g61865/_0_  = _w2811_ ;
	assign \g61866/_3_  = _w2822_ ;
	assign \g61867/_3_  = _w2830_ ;
	assign \g61868/u3_syn_7  = _w2831_ ;
	assign \g61869/_0_  = _w2840_ ;
	assign \g61870/_0_  = _w2847_ ;
	assign \g61871/_3_  = _w2858_ ;
	assign \g61872/_3_  = _w2865_ ;
	assign \g61873/u3_syn_7  = _w2866_ ;
	assign \g61874/_0_  = _w2875_ ;
	assign \g61875/_0_  = _w2882_ ;
	assign \g61877/_3_  = _w2893_ ;
	assign \g61878/_3_  = _w2900_ ;
	assign \g61879/u3_syn_7  = _w2901_ ;
	assign \g61880/_0_  = _w2910_ ;
	assign \g61881/_0_  = _w2916_ ;
	assign \g61882/_0_  = _w2922_ ;
	assign \g61883/_0_  = _w2928_ ;
	assign \g61884/_0_  = _w2934_ ;
	assign \g61914/_0_  = _w2937_ ;
	assign \g61915/_0_  = _w2946_ ;
	assign \g61917/_0_  = _w2971_ ;
	assign \g61918/_0_  = _w2977_ ;
	assign \g61922/_0_  = _w2986_ ;
	assign \g61923/_0_  = _w2992_ ;
	assign \g61924/_0_  = _w3001_ ;
	assign \g61932/_0_  = _w3024_ ;
	assign \g61936/_0_  = _w3033_ ;
	assign \g61945/_0_  = _w3038_ ;
	assign \g61947/_0_  = _w3042_ ;
	assign \g61959/_0_  = _w3050_ ;
	assign \g61960/_0_  = _w3055_ ;
	assign \g61962/_0_  = _w3060_ ;
	assign \g61973/_3_  = _w3065_ ;
	assign \g61974/u3_syn_7  = _w3066_ ;
	assign \g61975/_3_  = _w3087_ ;
	assign \g61976/u3_syn_7  = _w3088_ ;
	assign \g61977/_3_  = _w3093_ ;
	assign \g61978/_3_  = _w3113_ ;
	assign \g61979/u3_syn_7  = _w3114_ ;
	assign \g61980/_3_  = _w3119_ ;
	assign \g61981/_3_  = _w3139_ ;
	assign \g61982/_3_  = _w3145_ ;
	assign \g61983/u3_syn_7  = _w3146_ ;
	assign \g61984/_3_  = _w3151_ ;
	assign \g61985/_3_  = _w3171_ ;
	assign \g61986/u3_syn_7  = _w3172_ ;
	assign \g61987/_3_  = _w3177_ ;
	assign \g61988/_3_  = _w3197_ ;
	assign \g61989/u3_syn_7  = _w3198_ ;
	assign \g61990/_3_  = _w3203_ ;
	assign \g61991/_3_  = _w3223_ ;
	assign \g61992/u3_syn_7  = _w3224_ ;
	assign \g61993/_3_  = _w3229_ ;
	assign \g61994/u3_syn_7  = _w3230_ ;
	assign \g61995/_3_  = _w3250_ ;
	assign \g61996/_3_  = _w3255_ ;
	assign \g61997/_3_  = _w3275_ ;
	assign \g62022/_0_  = _w3283_ ;
	assign \g62028/_0_  = _w3291_ ;
	assign \g62029/_0_  = _w3294_ ;
	assign \g62031/_0_  = _w3315_ ;
	assign \g62033/_0_  = _w3323_ ;
	assign \g62038/_0_  = _w3331_ ;
	assign \g62042/_0_  = _w3339_ ;
	assign \g62046/_0_  = _w3347_ ;
	assign \g62048/_0_  = _w3353_ ;
	assign \g62049/_0_  = _w3361_ ;
	assign \g62051/_0_  = _w3369_ ;
	assign \g62053/_0_  = _w3384_ ;
	assign \g62085/_0_  = _w3389_ ;
	assign \g62101/_0_  = _w3397_ ;
	assign \g62102/_0_  = _w3406_ ;
	assign \g62103/_0_  = _w3412_ ;
	assign \g62105/_0_  = _w3417_ ;
	assign \g62108/_3_  = _w3420_ ;
	assign \g62112/_0_  = _w3425_ ;
	assign \g62137/_3_  = _w3433_ ;
	assign \g62207/_0_  = _w3436_ ;
	assign \g62239/_0_  = _w3454_ ;
	assign \g62240/_0_  = _w3459_ ;
	assign \g62267/_0_  = _w3466_ ;
	assign \g62273/_0_  = _w3475_ ;
	assign \g62284/_0_  = _w3480_ ;
	assign \g62291/_0_  = _w3482_ ;
	assign \g62293/_0_  = _w3487_ ;
	assign \g62298/_0_  = _w3492_ ;
	assign \g62303/_3_  = _w3515_ ;
	assign \g62322/_3_  = _w3523_ ;
	assign \g62323/_3_  = _w3526_ ;
	assign \g62324/_3_  = _w3530_ ;
	assign \g62325/_3_  = _w3536_ ;
	assign \g62583/_0_  = _w3552_ ;
	assign \g62598/_0_  = _w3557_ ;
	assign \g62609/_0_  = _w3567_ ;
	assign \g62636/_0_  = _w3582_ ;
	assign \g62646/_0_  = _w3588_ ;
	assign \g62649/_0_  = _w3594_ ;
	assign \g62658/_0_  = _w3599_ ;
	assign \g62663/_0_  = _w3601_ ;
	assign \g62664/_0_  = _w3603_ ;
	assign \g62667/_0_  = _w3610_ ;
	assign \g62676/_0_  = _w3616_ ;
	assign \g62677/_0_  = _w3620_ ;
	assign \g62678/_3_  = _w3626_ ;
	assign \g62679/_0_  = _w3631_ ;
	assign \g62687/u3_syn_7  = _w3632_ ;
	assign \g62688/u3_syn_7  = _w3633_ ;
	assign \g62689/_0_  = _w3642_ ;
	assign \g62690/_3_  = _w3648_ ;
	assign \g62691/_3_  = _w3654_ ;
	assign \g62693/_0_  = _w3663_ ;
	assign \g62694/_3_  = _w3670_ ;
	assign \g62695/_3_  = _w3678_ ;
	assign \g62696/_3_  = _w3686_ ;
	assign \g62697/_3_  = _w3693_ ;
	assign \g62698/_3_  = _w3699_ ;
	assign \g62699/_3_  = _w3705_ ;
	assign \g62700/_3_  = _w3711_ ;
	assign \g62701/_3_  = _w3717_ ;
	assign \g62702/_3_  = _w3723_ ;
	assign \g62703/_3_  = _w3727_ ;
	assign \g62704/u3_syn_7  = _w3724_ ;
	assign \g62705/_0_  = _w3736_ ;
	assign \g62706/_3_  = _w3742_ ;
	assign \g62707/_3_  = _w3746_ ;
	assign \g62708/u3_syn_7  = _w3743_ ;
	assign \g62709/_0_  = _w3755_ ;
	assign \g62710/_3_  = _w3761_ ;
	assign \g62711/_3_  = _w3765_ ;
	assign \g62712/u3_syn_7  = _w3762_ ;
	assign \g62713/_0_  = _w3774_ ;
	assign \g62714/_3_  = _w3780_ ;
	assign \g62715/_0_  = _w3784_ ;
	assign \g62716/u3_syn_7  = _w3781_ ;
	assign \g62717/_0_  = _w3793_ ;
	assign \g62718/_3_  = _w3799_ ;
	assign \g62719/_0_  = _w3803_ ;
	assign \g62720/u3_syn_7  = _w3800_ ;
	assign \g62721/_0_  = _w3812_ ;
	assign \g62722/_3_  = _w3818_ ;
	assign \g62723/_0_  = _w3822_ ;
	assign \g62724/u3_syn_7  = _w3819_ ;
	assign \g62725/_0_  = _w3831_ ;
	assign \g62726/_3_  = _w3837_ ;
	assign \g62728/_0_  = _w3840_ ;
	assign \g62790/_0_  = _w3845_ ;
	assign \g62791/_0_  = _w3854_ ;
	assign \g62793/_0_  = _w3859_ ;
	assign \g62794/_0_  = _w3864_ ;
	assign \g62795/_0_  = _w3869_ ;
	assign \g62796/_0_  = _w3874_ ;
	assign \g62797/_0_  = _w3879_ ;
	assign \g62807/_0_  = _w3888_ ;
	assign \g62823/_0_  = _w3891_ ;
	assign \g62824/_0_  = _w3896_ ;
	assign \g62833/_0_  = _w3903_ ;
	assign \g62846/_0_  = _w3911_ ;
	assign \g62859/_0_  = _w3916_ ;
	assign \g62860/_0_  = _w3921_ ;
	assign \g62897/_0_  = _w3926_ ;
	assign \g62898/_0_  = _w3930_ ;
	assign \g62922/_3_  = _w3936_ ;
	assign \g62923/_0_  = _w3940_ ;
	assign \g62927/_0_  = _w3945_ ;
	assign \g62938/_3_  = _w3950_ ;
	assign \g62939/_3_  = _w3959_ ;
	assign \g62940/_3_  = _w3964_ ;
	assign \g62941/u3_syn_7  = _w3967_ ;
	assign \g62942/_0_  = _w3976_ ;
	assign \g62943/_3_  = _w3982_ ;
	assign \g62987/_3_  = _w3987_ ;
	assign \g62991/_3_  = _w3990_ ;
	assign \g63015/u3_syn_7  = _w3994_ ;
	assign \g63016/_0_  = _w4003_ ;
	assign \g63017/_3_  = _w4014_ ;
	assign \g63018/_3_  = _w4022_ ;
	assign \g63019/_3_  = _w4028_ ;
	assign \g63020/_3_  = _w4035_ ;
	assign \g63021/_3_  = _w4043_ ;
	assign \g63022/_3_  = _w4050_ ;
	assign \g63025/_3_  = _w4058_ ;
	assign \g63026/_3_  = _w4065_ ;
	assign \g63027/_3_  = _w4072_ ;
	assign \g63029/_3_  = _w4080_ ;
	assign \g63030/_3_  = _w4087_ ;
	assign \g63031/_3_  = _w4094_ ;
	assign \g63033/_3_  = _w4102_ ;
	assign \g63034/_3_  = _w4109_ ;
	assign \g63043/_3_  = _w4117_ ;
	assign \g63044/_3_  = _w4124_ ;
	assign \g63051/_3_  = _w4131_ ;
	assign \g63057/_3_  = _w4138_ ;
	assign \g63068/_3_  = _w4145_ ;
	assign \g63070/_3_  = _w4152_ ;
	assign \g63073/_3_  = _w4159_ ;
	assign \g63081/_3_  = _w4164_ ;
	assign \g63082/_3_  = _w4167_ ;
	assign \g63083/u3_syn_7  = _w4168_ ;
	assign \g63084/_3_  = _w4175_ ;
	assign \g63085/_0_  = _w4187_ ;
	assign \g63086/_3_  = _w4193_ ;
	assign \g63107/_3_  = _w4198_ ;
	assign \g63108/u3_syn_7  = _w1534_ ;
	assign \g63109/u3_syn_7  = _w4201_ ;
	assign \g63110/_0_  = _w4210_ ;
	assign \g63111/_3_  = _w4216_ ;
	assign \g63132/_3_  = _w4221_ ;
	assign \g63133/_3_  = _w4224_ ;
	assign \g63134/_3_  = _w4231_ ;
	assign \g63135/_3_  = _w4236_ ;
	assign \g63136/_3_  = _w4241_ ;
	assign \g63137/_3_  = _w4244_ ;
	assign \g63138/_3_  = _w4250_ ;
	assign \g63139/u3_syn_7  = _w4251_ ;
	assign \g63140/_3_  = _w4256_ ;
	assign \g63141/_3_  = _w4259_ ;
	assign \g63142/_3_  = _w4265_ ;
	assign \g63143/_3_  = _w4270_ ;
	assign \g63144/_3_  = _w4276_ ;
	assign \g63145/_3_  = _w4280_ ;
	assign \g63146/u3_syn_7  = _w1450_ ;
	assign \g63198/_0_  = _w4287_ ;
	assign \g63205/_0_  = _w4293_ ;
	assign \g63208/_0_  = _w4298_ ;
	assign \g63212/_0_  = _w4304_ ;
	assign \g63215/_0_  = _w4310_ ;
	assign \g63219/_0_  = _w4316_ ;
	assign \g63244/_0_  = _w4324_ ;
	assign \g63246/_0_  = _w4326_ ;
	assign \g63254/_0_  = _w4331_ ;
	assign \g63255/_0_  = _w4338_ ;
	assign \g63272/_0_  = _w4345_ ;
	assign \g63276/_0_  = _w4350_ ;
	assign \g63278/_0_  = _w4357_ ;
	assign \g63279/_0_  = _w4363_ ;
	assign \g63280/_0_  = _w4366_ ;
	assign \g63327/_0_  = _w4371_ ;
	assign \g63345/_0_  = _w4375_ ;
	assign \g63346/_3_  = _w4378_ ;
	assign \g63347/_3_  = _w4386_ ;
	assign \g63354/_3_  = _w4390_ ;
	assign \g63358/_3_  = _w4402_ ;
	assign \g63359/u3_syn_7  = _w4403_ ;
	assign \g63361/_3_  = _w4407_ ;
	assign \g63365/_3_  = _w4410_ ;
	assign \g63366/_3_  = _w4413_ ;
	assign \g63367/_3_  = _w4416_ ;
	assign \g63368/_3_  = _w4418_ ;
	assign \g63370/_3_  = _w4424_ ;
	assign \g63479/_0_  = _w4428_ ;
	assign \g63484/_0_  = _w4432_ ;
	assign \g63499/_1_  = _w1782_ ;
	assign \g63520/_0_  = _w4436_ ;
	assign \g63523/_0_  = _w4442_ ;
	assign \g63526/_0_  = _w4446_ ;
	assign \g63538/_0_  = _w4450_ ;
	assign \g63539/_0_  = _w4460_ ;
	assign \g63541/_0_  = _w4464_ ;
	assign \g63555/_0_  = _w4477_ ;
	assign \g63642/_0_  = _w4484_ ;
	assign \g63645/_0_  = _w4489_ ;
	assign \g63648/_3_  = _w4494_ ;
	assign \g63777/_3_  = _w4499_ ;
	assign \g63778/_3_  = _w4510_ ;
	assign \g63781/_0_  = _w4514_ ;
	assign \g63786/u3_syn_7  = _w4515_ ;
	assign \g63787/_3_  = _w4520_ ;
	assign \g63788/_3_  = _w4524_ ;
	assign \g63790/_3_  = _w4530_ ;
	assign \g63791/_3_  = _w4539_ ;
	assign \g63792/u3_syn_7  = _w4511_ ;
	assign \g63794/_0_  = _w4547_ ;
	assign \g63795/_0_  = _w4555_ ;
	assign \g63796/_0_  = _w4562_ ;
	assign \g63798/_3_  = _w4568_ ;
	assign \g63800/_3_  = _w4574_ ;
	assign \g63804/_3_  = _w4580_ ;
	assign \g63805/_3_  = _w4586_ ;
	assign \g63806/_3_  = _w4591_ ;
	assign \g63807/_3_  = _w4597_ ;
	assign \g63808/_3_  = _w4603_ ;
	assign \g63809/_3_  = _w4611_ ;
	assign \g63870/_0_  = _w4617_ ;
	assign \g63883/_0_  = _w4619_ ;
	assign \g63934/_0_  = _w4625_ ;
	assign \g63936/_0_  = _w4626_ ;
	assign \g63938/_0_  = _w4630_ ;
	assign \g63939/_0_  = _w4633_ ;
	assign \g63966/_0_  = _w4642_ ;
	assign \g63970/_0_  = _w4650_ ;
	assign \g63999/_0_  = _w4657_ ;
	assign \g64039/_0_  = _w4661_ ;
	assign \g64040/_0_  = _w4671_ ;
	assign \g64043/_0_  = _w4676_ ;
	assign \g64062/_3_  = _w4678_ ;
	assign \g64078/_0_  = _w4681_ ;
	assign \g64091/_0_  = _w4686_ ;
	assign \g64095/_3_  = _w4689_ ;
	assign \g64096/_3_  = _w4693_ ;
	assign \g64097/u3_syn_7  = _w4694_ ;
	assign \g64098/u3_syn_7  = _w4695_ ;
	assign \g64099/u3_syn_7  = _w4696_ ;
	assign \g64100/u3_syn_7  = _w4697_ ;
	assign \g64134/_0_  = _w4703_ ;
	assign \g64135/_0_  = _w4709_ ;
	assign \g64153/_0_  = _w4717_ ;
	assign \g64155/_0_  = _w4719_ ;
	assign \g64179/_0_  = _w4727_ ;
	assign \g64229/_0_  = _w4734_ ;
	assign \g64235/_0_  = _w4741_ ;
	assign \g64236/_0_  = _w4748_ ;
	assign \g64280/_0_  = _w4757_ ;
	assign \g64315/_0_  = _w4760_ ;
	assign \g64365/_0_  = _w4764_ ;
	assign \g64426/_3_  = _w4770_ ;
	assign \g64438/_3_  = _w4776_ ;
	assign \g64442/u3_syn_7  = _w4777_ ;
	assign \g64445/_3_  = _w4783_ ;
	assign \g64447/_3_  = _w4789_ ;
	assign \g64449/_3_  = _w4795_ ;
	assign \g64451/_3_  = _w4803_ ;
	assign \g64453/_3_  = _w4806_ ;
	assign \g64454/_3_  = _w4809_ ;
	assign \g64460/_3_  = _w4816_ ;
	assign \g64461/_3_  = _w4821_ ;
	assign \g64510/_0_  = _w4822_ ;
	assign \g64527/_0_  = _w4825_ ;
	assign \g64528/_0_  = _w4826_ ;
	assign \g64544/_0_  = _w4833_ ;
	assign \g64549/_0_  = _w4840_ ;
	assign \g64566/_0_  = _w4847_ ;
	assign \g64576/_0_  = _w4853_ ;
	assign \g64602/_0_  = _w4860_ ;
	assign \g64691/_0_  = _w4865_ ;
	assign \g64697/_0_  = _w4868_ ;
	assign \g64707/_3_  = _w4873_ ;
	assign \g64778/_3_  = _w4876_ ;
	assign \g64790/_3_  = _w4880_ ;
	assign \g64791/_3_  = _w4884_ ;
	assign \g64792/_3_  = _w4888_ ;
	assign \g64793/_3_  = _w4892_ ;
	assign \g64794/_3_  = _w4897_ ;
	assign \g64795/_3_  = _w4901_ ;
	assign \g64796/_3_  = _w4905_ ;
	assign \g64797/_3_  = _w4909_ ;
	assign \g64877/_0_  = _w4910_ ;
	assign \g64912/_0_  = _w4911_ ;
	assign \g64973/_0_  = _w4918_ ;
	assign \g65047/_3_  = _w4921_ ;
	assign \g65081/_3_  = _w4925_ ;
	assign \g65088/_3_  = _w4929_ ;
	assign \g65097/_3_  = _w4932_ ;
	assign \g65100/_3_  = _w4936_ ;
	assign \g65101/_3_  = _w4940_ ;
	assign \g65104/_3_  = _w4945_ ;
	assign \g65105/_3_  = _w4949_ ;
	assign \g65107/_3_  = _w4951_ ;
	assign \g65110/_3_  = _w4955_ ;
	assign \g65111/_3_  = _w4961_ ;
	assign \g65113/_3_  = _w4967_ ;
	assign \g65114/_3_  = _w4973_ ;
	assign \g65266/_0_  = _w4974_ ;
	assign \g65267/_0_  = _w4975_ ;
	assign \g65294/_1_  = _w4710_ ;
	assign \g65328/_1_  = _w4976_ ;
	assign \g65495/_0_  = _w4979_ ;
	assign \g65499/_0_  = _w4983_ ;
	assign \g65503/_0_  = _w4986_ ;
	assign \g65529/_0_  = _w4990_ ;
	assign \g65530/_3_  = _w4994_ ;
	assign \g65531/_3_  = _w4998_ ;
	assign \g65532/_3_  = _w5001_ ;
	assign \g65533/_3_  = _w5005_ ;
	assign \g65624/_0_  = _w5007_ ;
	assign \g65625/_1_  = _w4153_ ;
	assign \g65641/_0_  = _w5009_ ;
	assign \g65701/_0_  = _w5012_ ;
	assign \g65704/_0_  = _w5013_ ;
	assign \g65853/_0_  = _w5014_ ;
	assign \g65891/_0_  = _w5015_ ;
	assign \g65901/_0_  = _w5017_ ;
	assign \g65986/_0_  = _w5018_ ;
	assign \g66029/_0_  = _w5020_ ;
	assign \g66066/_0_  = _w5022_ ;
	assign \g66067/_0_  = _w5024_ ;
	assign \g66068/_0_  = _w5026_ ;
	assign \g66154/_3_  = _w5029_ ;
	assign \g66362/_0_  = _w5030_ ;
	assign \g66369/_0_  = _w5031_ ;
	assign \g66398/_0_  = _w5032_ ;
	assign \g66409/_0_  = _w5033_ ;
	assign \g66419/_0_  = _w5034_ ;
	assign \g66439/_0_  = _w5035_ ;
	assign \g66443/_0_  = _w5036_ ;
	assign \g66464/_0_  = _w5037_ ;
	assign \g66471/_0_  = _w5038_ ;
	assign \g66512/_0_  = _w5039_ ;
	assign \g66528/_0_  = _w5040_ ;
	assign \g66541/_0_  = _w4565_ ;
	assign \g66558/_0_  = _w5041_ ;
	assign \g66644/_0_  = _w5042_ ;
	assign \g66684/_0_  = _w5043_ ;
	assign \g66697/_0_  = _w5044_ ;
	assign \g66698/_0_  = _w4912_ ;
	assign \g66701/_0_  = _w5045_ ;
	assign \g66714/_0_  = _w5046_ ;
	assign \g66715/_0_  = _w5047_ ;
	assign \g66745/_0_  = _w5048_ ;
	assign \g66750/_0_  = _w5049_ ;
	assign \g66751/_0_  = _w5050_ ;
	assign \g66810/_0_  = _w5051_ ;
	assign \g66844/_0_  = _w5052_ ;
	assign \g66853/_0_  = _w5053_ ;
	assign \g66897/_0_  = _w5054_ ;
	assign \g66905/_0_  = _w5055_ ;
	assign \g69743/_0_  = _w5059_ ;
	assign \g69750/_0_  = _w5063_ ;
	assign \g69773/_1_  = _w5066_ ;
	assign \g69792/_1_  = _w5070_ ;
	assign \g69858/_0_  = _w5074_ ;
	assign \g69938/_0_  = _w5085_ ;
	assign \g69949/_0_  = _w5089_ ;
	assign \g70167/_0_  = _w5097_ ;
	assign \g71190/_0_  = _w5106_ ;
	assign \g71198/_0_  = _w5114_ ;
	assign \g71284/_0_  = _w5131_ ;
	assign \g72369/_1_  = _w1949_ ;
	assign \g72467/_0_  = _w5135_ ;
	assign \g72476/_0_  = _w5159_ ;
	assign \g72477/_1_  = _w5158_ ;
	assign \g72648/_0_  = _w5168_ ;
	assign \g72741/_0_  = _w5173_ ;
	assign \g72772/_0_  = _w5177_ ;
	assign \g8132_pad  = 1'b0;
endmodule;