module top (\a0_pad , a_pad, \b0_pad , b_pad, \c0_pad , c_pad, \d0_pad , d_pad, \e0_pad , e_pad, \f0_pad , f_pad, g_pad, h_pad, i_pad, j_pad, k_pad, l_pad, m_pad, n_pad, o_pad, p_pad, q_pad, r_pad, s_pad, t_pad, u_pad, v_pad, w_pad, x_pad, y_pad, z_pad, \g0_pad , \h0_pad , \i0_pad );
	input \a0_pad  ;
	input a_pad ;
	input \b0_pad  ;
	input b_pad ;
	input \c0_pad  ;
	input c_pad ;
	input \d0_pad  ;
	input d_pad ;
	input \e0_pad  ;
	input e_pad ;
	input \f0_pad  ;
	input f_pad ;
	input g_pad ;
	input h_pad ;
	input i_pad ;
	input j_pad ;
	input k_pad ;
	input l_pad ;
	input m_pad ;
	input n_pad ;
	input o_pad ;
	input p_pad ;
	input q_pad ;
	input r_pad ;
	input s_pad ;
	input t_pad ;
	input u_pad ;
	input v_pad ;
	input w_pad ;
	input x_pad ;
	input y_pad ;
	input z_pad ;
	output \g0_pad  ;
	output \h0_pad  ;
	output \i0_pad  ;
	wire _w116_ ;
	wire _w115_ ;
	wire _w114_ ;
	wire _w113_ ;
	wire _w112_ ;
	wire _w111_ ;
	wire _w110_ ;
	wire _w109_ ;
	wire _w108_ ;
	wire _w107_ ;
	wire _w106_ ;
	wire _w105_ ;
	wire _w104_ ;
	wire _w103_ ;
	wire _w102_ ;
	wire _w101_ ;
	wire _w100_ ;
	wire _w99_ ;
	wire _w98_ ;
	wire _w97_ ;
	wire _w96_ ;
	wire _w95_ ;
	wire _w94_ ;
	wire _w93_ ;
	wire _w92_ ;
	wire _w61_ ;
	wire _w60_ ;
	wire _w59_ ;
	wire _w58_ ;
	wire _w57_ ;
	wire _w56_ ;
	wire _w55_ ;
	wire _w54_ ;
	wire _w53_ ;
	wire _w52_ ;
	wire _w51_ ;
	wire _w50_ ;
	wire _w49_ ;
	wire _w48_ ;
	wire _w47_ ;
	wire _w46_ ;
	wire _w33_ ;
	wire _w34_ ;
	wire _w35_ ;
	wire _w36_ ;
	wire _w37_ ;
	wire _w38_ ;
	wire _w39_ ;
	wire _w40_ ;
	wire _w41_ ;
	wire _w42_ ;
	wire _w43_ ;
	wire _w44_ ;
	wire _w45_ ;
	wire _w62_ ;
	wire _w63_ ;
	wire _w64_ ;
	wire _w65_ ;
	wire _w66_ ;
	wire _w67_ ;
	wire _w68_ ;
	wire _w69_ ;
	wire _w70_ ;
	wire _w71_ ;
	wire _w72_ ;
	wire _w73_ ;
	wire _w74_ ;
	wire _w75_ ;
	wire _w76_ ;
	wire _w77_ ;
	wire _w78_ ;
	wire _w79_ ;
	wire _w80_ ;
	wire _w81_ ;
	wire _w82_ ;
	wire _w83_ ;
	wire _w84_ ;
	wire _w85_ ;
	wire _w86_ ;
	wire _w87_ ;
	wire _w88_ ;
	wire _w89_ ;
	wire _w90_ ;
	wire _w91_ ;
	LUT2 #(
		.INIT('h2)
	) name0 (
		j_pad,
		z_pad,
		_w33_
	);
	LUT2 #(
		.INIT('h2)
	) name1 (
		i_pad,
		y_pad,
		_w34_
	);
	LUT2 #(
		.INIT('h1)
	) name2 (
		_w33_,
		_w34_,
		_w35_
	);
	LUT2 #(
		.INIT('h2)
	) name3 (
		\b0_pad ,
		l_pad,
		_w36_
	);
	LUT2 #(
		.INIT('h2)
	) name4 (
		\c0_pad ,
		m_pad,
		_w37_
	);
	LUT2 #(
		.INIT('h4)
	) name5 (
		i_pad,
		y_pad,
		_w38_
	);
	LUT2 #(
		.INIT('h2)
	) name6 (
		\a0_pad ,
		k_pad,
		_w39_
	);
	LUT2 #(
		.INIT('h4)
	) name7 (
		j_pad,
		z_pad,
		_w40_
	);
	LUT2 #(
		.INIT('h1)
	) name8 (
		_w39_,
		_w40_,
		_w41_
	);
	LUT2 #(
		.INIT('h4)
	) name9 (
		\a0_pad ,
		k_pad,
		_w42_
	);
	LUT2 #(
		.INIT('h4)
	) name10 (
		\b0_pad ,
		l_pad,
		_w43_
	);
	LUT2 #(
		.INIT('h1)
	) name11 (
		_w42_,
		_w43_,
		_w44_
	);
	LUT2 #(
		.INIT('h1)
	) name12 (
		_w36_,
		_w37_,
		_w45_
	);
	LUT2 #(
		.INIT('h4)
	) name13 (
		_w38_,
		_w45_,
		_w46_
	);
	LUT2 #(
		.INIT('h8)
	) name14 (
		_w35_,
		_w41_,
		_w47_
	);
	LUT2 #(
		.INIT('h8)
	) name15 (
		_w44_,
		_w47_,
		_w48_
	);
	LUT2 #(
		.INIT('h8)
	) name16 (
		_w46_,
		_w48_,
		_w49_
	);
	LUT2 #(
		.INIT('h4)
	) name17 (
		\c0_pad ,
		m_pad,
		_w50_
	);
	LUT2 #(
		.INIT('h4)
	) name18 (
		\e0_pad ,
		o_pad,
		_w51_
	);
	LUT2 #(
		.INIT('h4)
	) name19 (
		\f0_pad ,
		p_pad,
		_w52_
	);
	LUT2 #(
		.INIT('h1)
	) name20 (
		_w51_,
		_w52_,
		_w53_
	);
	LUT2 #(
		.INIT('h2)
	) name21 (
		\e0_pad ,
		o_pad,
		_w54_
	);
	LUT2 #(
		.INIT('h2)
	) name22 (
		\d0_pad ,
		n_pad,
		_w55_
	);
	LUT2 #(
		.INIT('h1)
	) name23 (
		_w54_,
		_w55_,
		_w56_
	);
	LUT2 #(
		.INIT('h4)
	) name24 (
		_w53_,
		_w56_,
		_w57_
	);
	LUT2 #(
		.INIT('h4)
	) name25 (
		\d0_pad ,
		n_pad,
		_w58_
	);
	LUT2 #(
		.INIT('h1)
	) name26 (
		_w50_,
		_w58_,
		_w59_
	);
	LUT2 #(
		.INIT('h4)
	) name27 (
		_w57_,
		_w59_,
		_w60_
	);
	LUT2 #(
		.INIT('h2)
	) name28 (
		_w49_,
		_w60_,
		_w61_
	);
	LUT2 #(
		.INIT('h2)
	) name29 (
		_w41_,
		_w44_,
		_w62_
	);
	LUT2 #(
		.INIT('h2)
	) name30 (
		_w35_,
		_w62_,
		_w63_
	);
	LUT2 #(
		.INIT('h1)
	) name31 (
		_w38_,
		_w63_,
		_w64_
	);
	LUT2 #(
		.INIT('h1)
	) name32 (
		_w61_,
		_w64_,
		_w65_
	);
	LUT2 #(
		.INIT('h4)
	) name33 (
		e_pad,
		u_pad,
		_w66_
	);
	LUT2 #(
		.INIT('h2)
	) name34 (
		e_pad,
		u_pad,
		_w67_
	);
	LUT2 #(
		.INIT('h2)
	) name35 (
		f_pad,
		v_pad,
		_w68_
	);
	LUT2 #(
		.INIT('h1)
	) name36 (
		_w67_,
		_w68_,
		_w69_
	);
	LUT2 #(
		.INIT('h2)
	) name37 (
		g_pad,
		w_pad,
		_w70_
	);
	LUT2 #(
		.INIT('h2)
	) name38 (
		h_pad,
		x_pad,
		_w71_
	);
	LUT2 #(
		.INIT('h1)
	) name39 (
		_w70_,
		_w71_,
		_w72_
	);
	LUT2 #(
		.INIT('h4)
	) name40 (
		f_pad,
		v_pad,
		_w73_
	);
	LUT2 #(
		.INIT('h4)
	) name41 (
		g_pad,
		w_pad,
		_w74_
	);
	LUT2 #(
		.INIT('h1)
	) name42 (
		_w73_,
		_w74_,
		_w75_
	);
	LUT2 #(
		.INIT('h4)
	) name43 (
		_w72_,
		_w75_,
		_w76_
	);
	LUT2 #(
		.INIT('h2)
	) name44 (
		_w69_,
		_w76_,
		_w77_
	);
	LUT2 #(
		.INIT('h1)
	) name45 (
		_w66_,
		_w77_,
		_w78_
	);
	LUT2 #(
		.INIT('h2)
	) name46 (
		b_pad,
		r_pad,
		_w79_
	);
	LUT2 #(
		.INIT('h2)
	) name47 (
		a_pad,
		q_pad,
		_w80_
	);
	LUT2 #(
		.INIT('h1)
	) name48 (
		_w79_,
		_w80_,
		_w81_
	);
	LUT2 #(
		.INIT('h4)
	) name49 (
		a_pad,
		q_pad,
		_w82_
	);
	LUT2 #(
		.INIT('h4)
	) name50 (
		d_pad,
		t_pad,
		_w83_
	);
	LUT2 #(
		.INIT('h2)
	) name51 (
		c_pad,
		s_pad,
		_w84_
	);
	LUT2 #(
		.INIT('h2)
	) name52 (
		d_pad,
		t_pad,
		_w85_
	);
	LUT2 #(
		.INIT('h1)
	) name53 (
		_w84_,
		_w85_,
		_w86_
	);
	LUT2 #(
		.INIT('h4)
	) name54 (
		c_pad,
		s_pad,
		_w87_
	);
	LUT2 #(
		.INIT('h4)
	) name55 (
		b_pad,
		r_pad,
		_w88_
	);
	LUT2 #(
		.INIT('h1)
	) name56 (
		_w87_,
		_w88_,
		_w89_
	);
	LUT2 #(
		.INIT('h1)
	) name57 (
		_w82_,
		_w83_,
		_w90_
	);
	LUT2 #(
		.INIT('h8)
	) name58 (
		_w81_,
		_w90_,
		_w91_
	);
	LUT2 #(
		.INIT('h8)
	) name59 (
		_w86_,
		_w89_,
		_w92_
	);
	LUT2 #(
		.INIT('h8)
	) name60 (
		_w91_,
		_w92_,
		_w93_
	);
	LUT2 #(
		.INIT('h4)
	) name61 (
		_w86_,
		_w89_,
		_w94_
	);
	LUT2 #(
		.INIT('h2)
	) name62 (
		_w81_,
		_w94_,
		_w95_
	);
	LUT2 #(
		.INIT('h1)
	) name63 (
		_w82_,
		_w95_,
		_w96_
	);
	LUT2 #(
		.INIT('h4)
	) name64 (
		h_pad,
		x_pad,
		_w97_
	);
	LUT2 #(
		.INIT('h1)
	) name65 (
		_w66_,
		_w97_,
		_w98_
	);
	LUT2 #(
		.INIT('h8)
	) name66 (
		_w69_,
		_w98_,
		_w99_
	);
	LUT2 #(
		.INIT('h8)
	) name67 (
		_w72_,
		_w75_,
		_w100_
	);
	LUT2 #(
		.INIT('h8)
	) name68 (
		_w99_,
		_w100_,
		_w101_
	);
	LUT2 #(
		.INIT('h8)
	) name69 (
		_w93_,
		_w101_,
		_w102_
	);
	LUT2 #(
		.INIT('h4)
	) name70 (
		_w78_,
		_w102_,
		_w103_
	);
	LUT2 #(
		.INIT('h4)
	) name71 (
		_w96_,
		_w103_,
		_w104_
	);
	LUT2 #(
		.INIT('h4)
	) name72 (
		_w65_,
		_w104_,
		_w105_
	);
	LUT2 #(
		.INIT('h8)
	) name73 (
		_w78_,
		_w93_,
		_w106_
	);
	LUT2 #(
		.INIT('h1)
	) name74 (
		_w96_,
		_w106_,
		_w107_
	);
	LUT2 #(
		.INIT('h4)
	) name75 (
		_w105_,
		_w107_,
		_w108_
	);
	LUT2 #(
		.INIT('h2)
	) name76 (
		\f0_pad ,
		p_pad,
		_w109_
	);
	LUT2 #(
		.INIT('h2)
	) name77 (
		_w53_,
		_w109_,
		_w110_
	);
	LUT2 #(
		.INIT('h8)
	) name78 (
		_w56_,
		_w110_,
		_w111_
	);
	LUT2 #(
		.INIT('h8)
	) name79 (
		_w60_,
		_w111_,
		_w112_
	);
	LUT2 #(
		.INIT('h8)
	) name80 (
		_w49_,
		_w112_,
		_w113_
	);
	LUT2 #(
		.INIT('h4)
	) name81 (
		_w64_,
		_w113_,
		_w114_
	);
	LUT2 #(
		.INIT('h8)
	) name82 (
		_w104_,
		_w114_,
		_w115_
	);
	LUT2 #(
		.INIT('h2)
	) name83 (
		_w108_,
		_w115_,
		_w116_
	);
	assign \g0_pad  = _w116_ ;
	assign \h0_pad  = _w115_ ;
	assign \i0_pad  = _w108_ ;
endmodule;