module top (\d_in_reg[0]/NET0131 , \d_in_reg[1]/NET0131 , \d_in_reg[2]/NET0131 , \d_in_reg[3]/NET0131 , \d_in_reg[4]/NET0131 , \d_in_reg[5]/NET0131 , \d_in_reg[6]/NET0131 , \d_in_reg[7]/NET0131 , \d_in_reg[8]/NET0131 , \d_out_reg[0]/NET0131 , \d_out_reg[1]/NET0131 , \d_out_reg[2]/NET0131 , \d_out_reg[3]/NET0131 , \d_out_reg[4]/NET0131 , \d_out_reg[5]/NET0131 , \d_out_reg[6]/NET0131 , \d_out_reg[7]/NET0131 , \old_reg[0]/NET0131 , \old_reg[1]/NET0131 , \old_reg[2]/NET0131 , \old_reg[3]/NET0131 , \old_reg[4]/NET0131 , \old_reg[5]/NET0131 , \old_reg[6]/NET0131 , \old_reg[7]/NET0131 , \stato_reg[0]/NET0131 , \stato_reg[1]/NET0131 , x_pad, y_pad, \_al_n0 , \_al_n1 , \g1026/_0_ , \g1035/_0_ , \g41/_0_ , \g708/_0_ , \g709/_0_ , \g711/_0_ , \g712/_0_ , \g714/_0_ , \g716/_0_ , \g718/_0_ , \g728/_0_ , \g770/_0_ , \g771/_0_ , \g772/_0_ , \g773/_0_ , \g774/_0_ , \g775/_0_ , \g776/_0_ , \g777/_0_ , \g782/_0_ , \g783/_0_ , \g784/_0_ , \g785/_0_ , \g786/_0_ , \g787/_0_ , \g788/_0_ , \g789/_0_ , \g806/_0_ );
	input \d_in_reg[0]/NET0131  ;
	input \d_in_reg[1]/NET0131  ;
	input \d_in_reg[2]/NET0131  ;
	input \d_in_reg[3]/NET0131  ;
	input \d_in_reg[4]/NET0131  ;
	input \d_in_reg[5]/NET0131  ;
	input \d_in_reg[6]/NET0131  ;
	input \d_in_reg[7]/NET0131  ;
	input \d_in_reg[8]/NET0131  ;
	input \d_out_reg[0]/NET0131  ;
	input \d_out_reg[1]/NET0131  ;
	input \d_out_reg[2]/NET0131  ;
	input \d_out_reg[3]/NET0131  ;
	input \d_out_reg[4]/NET0131  ;
	input \d_out_reg[5]/NET0131  ;
	input \d_out_reg[6]/NET0131  ;
	input \d_out_reg[7]/NET0131  ;
	input \old_reg[0]/NET0131  ;
	input \old_reg[1]/NET0131  ;
	input \old_reg[2]/NET0131  ;
	input \old_reg[3]/NET0131  ;
	input \old_reg[4]/NET0131  ;
	input \old_reg[5]/NET0131  ;
	input \old_reg[6]/NET0131  ;
	input \old_reg[7]/NET0131  ;
	input \stato_reg[0]/NET0131  ;
	input \stato_reg[1]/NET0131  ;
	input x_pad ;
	input y_pad ;
	output \_al_n0  ;
	output \_al_n1  ;
	output \g1026/_0_  ;
	output \g1035/_0_  ;
	output \g41/_0_  ;
	output \g708/_0_  ;
	output \g709/_0_  ;
	output \g711/_0_  ;
	output \g712/_0_  ;
	output \g714/_0_  ;
	output \g716/_0_  ;
	output \g718/_0_  ;
	output \g728/_0_  ;
	output \g770/_0_  ;
	output \g771/_0_  ;
	output \g772/_0_  ;
	output \g773/_0_  ;
	output \g774/_0_  ;
	output \g775/_0_  ;
	output \g776/_0_  ;
	output \g777/_0_  ;
	output \g782/_0_  ;
	output \g783/_0_  ;
	output \g784/_0_  ;
	output \g785/_0_  ;
	output \g786/_0_  ;
	output \g787/_0_  ;
	output \g788/_0_  ;
	output \g789/_0_  ;
	output \g806/_0_  ;
	wire _w135_ ;
	wire _w134_ ;
	wire _w133_ ;
	wire _w132_ ;
	wire _w131_ ;
	wire _w130_ ;
	wire _w129_ ;
	wire _w128_ ;
	wire _w127_ ;
	wire _w126_ ;
	wire _w125_ ;
	wire _w124_ ;
	wire _w123_ ;
	wire _w122_ ;
	wire _w121_ ;
	wire _w120_ ;
	wire _w119_ ;
	wire _w118_ ;
	wire _w117_ ;
	wire _w116_ ;
	wire _w115_ ;
	wire _w114_ ;
	wire _w113_ ;
	wire _w112_ ;
	wire _w111_ ;
	wire _w110_ ;
	wire _w109_ ;
	wire _w108_ ;
	wire _w107_ ;
	wire _w106_ ;
	wire _w105_ ;
	wire _w104_ ;
	wire _w103_ ;
	wire _w102_ ;
	wire _w101_ ;
	wire _w100_ ;
	wire _w99_ ;
	wire _w98_ ;
	wire _w97_ ;
	wire _w96_ ;
	wire _w95_ ;
	wire _w94_ ;
	wire _w93_ ;
	wire _w92_ ;
	wire _w91_ ;
	wire _w90_ ;
	wire _w59_ ;
	wire _w58_ ;
	wire _w57_ ;
	wire _w56_ ;
	wire _w55_ ;
	wire _w54_ ;
	wire _w53_ ;
	wire _w52_ ;
	wire _w51_ ;
	wire _w50_ ;
	wire _w49_ ;
	wire _w48_ ;
	wire _w47_ ;
	wire _w46_ ;
	wire _w45_ ;
	wire _w44_ ;
	wire _w31_ ;
	wire _w32_ ;
	wire _w33_ ;
	wire _w34_ ;
	wire _w35_ ;
	wire _w36_ ;
	wire _w37_ ;
	wire _w38_ ;
	wire _w39_ ;
	wire _w40_ ;
	wire _w41_ ;
	wire _w42_ ;
	wire _w43_ ;
	wire _w60_ ;
	wire _w61_ ;
	wire _w62_ ;
	wire _w63_ ;
	wire _w64_ ;
	wire _w65_ ;
	wire _w66_ ;
	wire _w67_ ;
	wire _w68_ ;
	wire _w69_ ;
	wire _w70_ ;
	wire _w71_ ;
	wire _w72_ ;
	wire _w73_ ;
	wire _w74_ ;
	wire _w75_ ;
	wire _w76_ ;
	wire _w77_ ;
	wire _w78_ ;
	wire _w79_ ;
	wire _w80_ ;
	wire _w81_ ;
	wire _w82_ ;
	wire _w83_ ;
	wire _w84_ ;
	wire _w85_ ;
	wire _w86_ ;
	wire _w87_ ;
	wire _w88_ ;
	wire _w89_ ;
	LUT4 #(
		.INIT('h8421)
	) name0 (
		\d_in_reg[4]/NET0131 ,
		\d_in_reg[5]/NET0131 ,
		\old_reg[3]/NET0131 ,
		\old_reg[4]/NET0131 ,
		_w31_
	);
	LUT4 #(
		.INIT('h8421)
	) name1 (
		\d_in_reg[7]/NET0131 ,
		\d_in_reg[8]/NET0131 ,
		\old_reg[6]/NET0131 ,
		\old_reg[7]/NET0131 ,
		_w32_
	);
	LUT4 #(
		.INIT('h8421)
	) name2 (
		\d_in_reg[3]/NET0131 ,
		\d_in_reg[6]/NET0131 ,
		\old_reg[2]/NET0131 ,
		\old_reg[5]/NET0131 ,
		_w33_
	);
	LUT4 #(
		.INIT('h8421)
	) name3 (
		\d_in_reg[1]/NET0131 ,
		\d_in_reg[2]/NET0131 ,
		\old_reg[0]/NET0131 ,
		\old_reg[1]/NET0131 ,
		_w34_
	);
	LUT4 #(
		.INIT('h8000)
	) name4 (
		_w31_,
		_w32_,
		_w33_,
		_w34_,
		_w35_
	);
	LUT3 #(
		.INIT('h80)
	) name5 (
		\d_in_reg[0]/NET0131 ,
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		_w36_
	);
	LUT4 #(
		.INIT('h8000)
	) name6 (
		\d_in_reg[0]/NET0131 ,
		\d_in_reg[1]/NET0131 ,
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		_w37_
	);
	LUT4 #(
		.INIT('h8000)
	) name7 (
		\d_in_reg[0]/NET0131 ,
		\d_out_reg[0]/NET0131 ,
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		_w38_
	);
	LUT4 #(
		.INIT('hb7bf)
	) name8 (
		\d_in_reg[0]/NET0131 ,
		\d_out_reg[0]/NET0131 ,
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		_w39_
	);
	LUT2 #(
		.INIT('h2)
	) name9 (
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		_w40_
	);
	LUT4 #(
		.INIT('h0080)
	) name10 (
		\d_in_reg[0]/NET0131 ,
		\d_in_reg[1]/NET0131 ,
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		_w41_
	);
	LUT4 #(
		.INIT('h0400)
	) name11 (
		\d_in_reg[0]/NET0131 ,
		\d_out_reg[1]/NET0131 ,
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		_w42_
	);
	LUT3 #(
		.INIT('h02)
	) name12 (
		_w39_,
		_w41_,
		_w42_,
		_w43_
	);
	LUT4 #(
		.INIT('he4ff)
	) name13 (
		_w35_,
		_w37_,
		_w38_,
		_w43_,
		_w44_
	);
	LUT4 #(
		.INIT('h8000)
	) name14 (
		\d_in_reg[0]/NET0131 ,
		\d_in_reg[2]/NET0131 ,
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		_w45_
	);
	LUT4 #(
		.INIT('h8000)
	) name15 (
		\d_in_reg[0]/NET0131 ,
		\d_out_reg[1]/NET0131 ,
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		_w46_
	);
	LUT4 #(
		.INIT('hb7bf)
	) name16 (
		\d_in_reg[0]/NET0131 ,
		\d_out_reg[1]/NET0131 ,
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		_w47_
	);
	LUT4 #(
		.INIT('h0080)
	) name17 (
		\d_in_reg[0]/NET0131 ,
		\d_in_reg[2]/NET0131 ,
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		_w48_
	);
	LUT4 #(
		.INIT('h0400)
	) name18 (
		\d_in_reg[0]/NET0131 ,
		\d_out_reg[2]/NET0131 ,
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		_w49_
	);
	LUT3 #(
		.INIT('h02)
	) name19 (
		_w47_,
		_w48_,
		_w49_,
		_w50_
	);
	LUT4 #(
		.INIT('he4ff)
	) name20 (
		_w35_,
		_w45_,
		_w46_,
		_w50_,
		_w51_
	);
	LUT4 #(
		.INIT('h8000)
	) name21 (
		\d_in_reg[0]/NET0131 ,
		\d_in_reg[8]/NET0131 ,
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		_w52_
	);
	LUT4 #(
		.INIT('h8000)
	) name22 (
		\d_in_reg[0]/NET0131 ,
		\d_out_reg[7]/NET0131 ,
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		_w53_
	);
	LUT4 #(
		.INIT('hb7bf)
	) name23 (
		\d_in_reg[0]/NET0131 ,
		\d_out_reg[7]/NET0131 ,
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		_w54_
	);
	LUT4 #(
		.INIT('h0080)
	) name24 (
		\d_in_reg[0]/NET0131 ,
		\d_in_reg[8]/NET0131 ,
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		_w55_
	);
	LUT2 #(
		.INIT('h2)
	) name25 (
		_w54_,
		_w55_,
		_w56_
	);
	LUT4 #(
		.INIT('he4ff)
	) name26 (
		_w35_,
		_w52_,
		_w53_,
		_w56_,
		_w57_
	);
	LUT4 #(
		.INIT('h0377)
	) name27 (
		\d_in_reg[0]/NET0131 ,
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		x_pad,
		_w58_
	);
	LUT4 #(
		.INIT('h80f0)
	) name28 (
		\d_in_reg[0]/NET0131 ,
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		x_pad,
		_w59_
	);
	LUT3 #(
		.INIT('h13)
	) name29 (
		_w35_,
		_w58_,
		_w59_,
		_w60_
	);
	LUT4 #(
		.INIT('h8000)
	) name30 (
		\d_in_reg[0]/NET0131 ,
		\d_in_reg[4]/NET0131 ,
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		_w61_
	);
	LUT4 #(
		.INIT('h8000)
	) name31 (
		\d_in_reg[0]/NET0131 ,
		\d_out_reg[3]/NET0131 ,
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		_w62_
	);
	LUT4 #(
		.INIT('hb7ff)
	) name32 (
		\d_in_reg[0]/NET0131 ,
		\d_out_reg[3]/NET0131 ,
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		_w63_
	);
	LUT3 #(
		.INIT('h27)
	) name33 (
		\d_in_reg[0]/NET0131 ,
		\d_in_reg[4]/NET0131 ,
		\d_out_reg[3]/NET0131 ,
		_w64_
	);
	LUT4 #(
		.INIT('h0400)
	) name34 (
		\d_in_reg[0]/NET0131 ,
		\d_out_reg[4]/NET0131 ,
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		_w65_
	);
	LUT4 #(
		.INIT('h00c4)
	) name35 (
		_w40_,
		_w63_,
		_w64_,
		_w65_,
		_w66_
	);
	LUT4 #(
		.INIT('he4ff)
	) name36 (
		_w35_,
		_w61_,
		_w62_,
		_w66_,
		_w67_
	);
	LUT4 #(
		.INIT('h8000)
	) name37 (
		\d_in_reg[0]/NET0131 ,
		\d_in_reg[5]/NET0131 ,
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		_w68_
	);
	LUT4 #(
		.INIT('h8000)
	) name38 (
		\d_in_reg[0]/NET0131 ,
		\d_out_reg[4]/NET0131 ,
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		_w69_
	);
	LUT4 #(
		.INIT('hb7bf)
	) name39 (
		\d_in_reg[0]/NET0131 ,
		\d_out_reg[4]/NET0131 ,
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		_w70_
	);
	LUT4 #(
		.INIT('h0080)
	) name40 (
		\d_in_reg[0]/NET0131 ,
		\d_in_reg[5]/NET0131 ,
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		_w71_
	);
	LUT4 #(
		.INIT('h0400)
	) name41 (
		\d_in_reg[0]/NET0131 ,
		\d_out_reg[5]/NET0131 ,
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		_w72_
	);
	LUT3 #(
		.INIT('h02)
	) name42 (
		_w70_,
		_w71_,
		_w72_,
		_w73_
	);
	LUT4 #(
		.INIT('he4ff)
	) name43 (
		_w35_,
		_w68_,
		_w69_,
		_w73_,
		_w74_
	);
	LUT4 #(
		.INIT('h8000)
	) name44 (
		\d_in_reg[0]/NET0131 ,
		\d_in_reg[6]/NET0131 ,
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		_w75_
	);
	LUT4 #(
		.INIT('h8000)
	) name45 (
		\d_in_reg[0]/NET0131 ,
		\d_out_reg[5]/NET0131 ,
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		_w76_
	);
	LUT4 #(
		.INIT('hb7bf)
	) name46 (
		\d_in_reg[0]/NET0131 ,
		\d_out_reg[5]/NET0131 ,
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		_w77_
	);
	LUT4 #(
		.INIT('h0080)
	) name47 (
		\d_in_reg[0]/NET0131 ,
		\d_in_reg[6]/NET0131 ,
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		_w78_
	);
	LUT4 #(
		.INIT('h0400)
	) name48 (
		\d_in_reg[0]/NET0131 ,
		\d_out_reg[6]/NET0131 ,
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		_w79_
	);
	LUT3 #(
		.INIT('h02)
	) name49 (
		_w77_,
		_w78_,
		_w79_,
		_w80_
	);
	LUT4 #(
		.INIT('he4ff)
	) name50 (
		_w35_,
		_w75_,
		_w76_,
		_w80_,
		_w81_
	);
	LUT4 #(
		.INIT('h8000)
	) name51 (
		\d_in_reg[0]/NET0131 ,
		\d_in_reg[7]/NET0131 ,
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		_w82_
	);
	LUT4 #(
		.INIT('h8000)
	) name52 (
		\d_in_reg[0]/NET0131 ,
		\d_out_reg[6]/NET0131 ,
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		_w83_
	);
	LUT4 #(
		.INIT('hb7bf)
	) name53 (
		\d_in_reg[0]/NET0131 ,
		\d_out_reg[6]/NET0131 ,
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		_w84_
	);
	LUT4 #(
		.INIT('h0080)
	) name54 (
		\d_in_reg[0]/NET0131 ,
		\d_in_reg[7]/NET0131 ,
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		_w85_
	);
	LUT4 #(
		.INIT('h0400)
	) name55 (
		\d_in_reg[0]/NET0131 ,
		\d_out_reg[7]/NET0131 ,
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		_w86_
	);
	LUT3 #(
		.INIT('h02)
	) name56 (
		_w84_,
		_w85_,
		_w86_,
		_w87_
	);
	LUT4 #(
		.INIT('he4ff)
	) name57 (
		_w35_,
		_w82_,
		_w83_,
		_w87_,
		_w88_
	);
	LUT4 #(
		.INIT('h8000)
	) name58 (
		\d_in_reg[0]/NET0131 ,
		\d_in_reg[3]/NET0131 ,
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		_w89_
	);
	LUT4 #(
		.INIT('h8000)
	) name59 (
		\d_in_reg[0]/NET0131 ,
		\d_out_reg[2]/NET0131 ,
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		_w90_
	);
	LUT4 #(
		.INIT('hb7bf)
	) name60 (
		\d_in_reg[0]/NET0131 ,
		\d_out_reg[2]/NET0131 ,
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		_w91_
	);
	LUT4 #(
		.INIT('h0400)
	) name61 (
		\d_in_reg[0]/NET0131 ,
		\d_out_reg[3]/NET0131 ,
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		_w92_
	);
	LUT4 #(
		.INIT('h0080)
	) name62 (
		\d_in_reg[0]/NET0131 ,
		\d_in_reg[3]/NET0131 ,
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		_w93_
	);
	LUT3 #(
		.INIT('h02)
	) name63 (
		_w91_,
		_w92_,
		_w93_,
		_w94_
	);
	LUT4 #(
		.INIT('he4ff)
	) name64 (
		_w35_,
		_w89_,
		_w90_,
		_w94_,
		_w95_
	);
	LUT3 #(
		.INIT('h67)
	) name65 (
		\d_in_reg[0]/NET0131 ,
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		_w96_
	);
	LUT3 #(
		.INIT('he0)
	) name66 (
		\d_in_reg[0]/NET0131 ,
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		_w97_
	);
	LUT3 #(
		.INIT('hec)
	) name67 (
		_w35_,
		_w96_,
		_w97_,
		_w98_
	);
	LUT4 #(
		.INIT('h0c08)
	) name68 (
		\d_in_reg[0]/NET0131 ,
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		y_pad,
		_w99_
	);
	LUT4 #(
		.INIT('h0400)
	) name69 (
		\d_in_reg[0]/NET0131 ,
		\d_out_reg[0]/NET0131 ,
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		_w100_
	);
	LUT2 #(
		.INIT('h1)
	) name70 (
		_w99_,
		_w100_,
		_w101_
	);
	LUT3 #(
		.INIT('h4f)
	) name71 (
		_w35_,
		_w36_,
		_w101_,
		_w102_
	);
	LUT4 #(
		.INIT('h4c40)
	) name72 (
		\d_in_reg[0]/NET0131 ,
		\d_in_reg[2]/NET0131 ,
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		_w103_
	);
	LUT4 #(
		.INIT('h4c40)
	) name73 (
		\d_in_reg[0]/NET0131 ,
		\d_in_reg[7]/NET0131 ,
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		_w104_
	);
	LUT4 #(
		.INIT('h4c40)
	) name74 (
		\d_in_reg[0]/NET0131 ,
		\d_in_reg[8]/NET0131 ,
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		_w105_
	);
	LUT4 #(
		.INIT('h4c40)
	) name75 (
		\d_in_reg[0]/NET0131 ,
		\d_in_reg[1]/NET0131 ,
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		_w106_
	);
	LUT4 #(
		.INIT('h4c40)
	) name76 (
		\d_in_reg[0]/NET0131 ,
		\d_in_reg[6]/NET0131 ,
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		_w107_
	);
	LUT4 #(
		.INIT('h4c40)
	) name77 (
		\d_in_reg[0]/NET0131 ,
		\d_in_reg[3]/NET0131 ,
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		_w108_
	);
	LUT4 #(
		.INIT('h4c40)
	) name78 (
		\d_in_reg[0]/NET0131 ,
		\d_in_reg[4]/NET0131 ,
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		_w109_
	);
	LUT4 #(
		.INIT('h4c40)
	) name79 (
		\d_in_reg[0]/NET0131 ,
		\d_in_reg[5]/NET0131 ,
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		_w110_
	);
	LUT4 #(
		.INIT('hd800)
	) name80 (
		\d_in_reg[0]/NET0131 ,
		\d_in_reg[6]/NET0131 ,
		\old_reg[5]/NET0131 ,
		\stato_reg[0]/NET0131 ,
		_w111_
	);
	LUT3 #(
		.INIT('h20)
	) name81 (
		\old_reg[5]/NET0131 ,
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		_w112_
	);
	LUT2 #(
		.INIT('he)
	) name82 (
		_w111_,
		_w112_,
		_w113_
	);
	LUT4 #(
		.INIT('hd800)
	) name83 (
		\d_in_reg[0]/NET0131 ,
		\d_in_reg[7]/NET0131 ,
		\old_reg[6]/NET0131 ,
		\stato_reg[0]/NET0131 ,
		_w114_
	);
	LUT3 #(
		.INIT('h20)
	) name84 (
		\old_reg[6]/NET0131 ,
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		_w115_
	);
	LUT2 #(
		.INIT('he)
	) name85 (
		_w114_,
		_w115_,
		_w116_
	);
	LUT4 #(
		.INIT('hd800)
	) name86 (
		\d_in_reg[0]/NET0131 ,
		\d_in_reg[8]/NET0131 ,
		\old_reg[7]/NET0131 ,
		\stato_reg[0]/NET0131 ,
		_w117_
	);
	LUT3 #(
		.INIT('h20)
	) name87 (
		\old_reg[7]/NET0131 ,
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		_w118_
	);
	LUT2 #(
		.INIT('he)
	) name88 (
		_w117_,
		_w118_,
		_w119_
	);
	LUT4 #(
		.INIT('hd800)
	) name89 (
		\d_in_reg[0]/NET0131 ,
		\d_in_reg[1]/NET0131 ,
		\old_reg[0]/NET0131 ,
		\stato_reg[0]/NET0131 ,
		_w120_
	);
	LUT3 #(
		.INIT('h20)
	) name90 (
		\old_reg[0]/NET0131 ,
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		_w121_
	);
	LUT2 #(
		.INIT('he)
	) name91 (
		_w120_,
		_w121_,
		_w122_
	);
	LUT4 #(
		.INIT('hd800)
	) name92 (
		\d_in_reg[0]/NET0131 ,
		\d_in_reg[2]/NET0131 ,
		\old_reg[1]/NET0131 ,
		\stato_reg[0]/NET0131 ,
		_w123_
	);
	LUT3 #(
		.INIT('h20)
	) name93 (
		\old_reg[1]/NET0131 ,
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		_w124_
	);
	LUT2 #(
		.INIT('he)
	) name94 (
		_w123_,
		_w124_,
		_w125_
	);
	LUT3 #(
		.INIT('h80)
	) name95 (
		\d_in_reg[0]/NET0131 ,
		\d_in_reg[3]/NET0131 ,
		\stato_reg[0]/NET0131 ,
		_w126_
	);
	LUT4 #(
		.INIT('h4c40)
	) name96 (
		\d_in_reg[0]/NET0131 ,
		\old_reg[2]/NET0131 ,
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		_w127_
	);
	LUT2 #(
		.INIT('he)
	) name97 (
		_w126_,
		_w127_,
		_w128_
	);
	LUT4 #(
		.INIT('hd800)
	) name98 (
		\d_in_reg[0]/NET0131 ,
		\d_in_reg[4]/NET0131 ,
		\old_reg[3]/NET0131 ,
		\stato_reg[0]/NET0131 ,
		_w129_
	);
	LUT3 #(
		.INIT('h20)
	) name99 (
		\old_reg[3]/NET0131 ,
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		_w130_
	);
	LUT2 #(
		.INIT('he)
	) name100 (
		_w129_,
		_w130_,
		_w131_
	);
	LUT4 #(
		.INIT('hd800)
	) name101 (
		\d_in_reg[0]/NET0131 ,
		\d_in_reg[5]/NET0131 ,
		\old_reg[4]/NET0131 ,
		\stato_reg[0]/NET0131 ,
		_w132_
	);
	LUT3 #(
		.INIT('h20)
	) name102 (
		\old_reg[4]/NET0131 ,
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		_w133_
	);
	LUT2 #(
		.INIT('he)
	) name103 (
		_w132_,
		_w133_,
		_w134_
	);
	LUT3 #(
		.INIT('hf8)
	) name104 (
		\d_in_reg[0]/NET0131 ,
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		_w135_
	);
	assign \_al_n0  = 1'b0;
	assign \_al_n1  = 1'b1;
	assign \g1026/_0_  = _w44_ ;
	assign \g1035/_0_  = _w51_ ;
	assign \g41/_0_  = _w57_ ;
	assign \g708/_0_  = _w60_ ;
	assign \g709/_0_  = _w67_ ;
	assign \g711/_0_  = _w74_ ;
	assign \g712/_0_  = _w81_ ;
	assign \g714/_0_  = _w88_ ;
	assign \g716/_0_  = _w95_ ;
	assign \g718/_0_  = _w98_ ;
	assign \g728/_0_  = _w102_ ;
	assign \g770/_0_  = _w103_ ;
	assign \g771/_0_  = _w104_ ;
	assign \g772/_0_  = _w105_ ;
	assign \g773/_0_  = _w106_ ;
	assign \g774/_0_  = _w107_ ;
	assign \g775/_0_  = _w108_ ;
	assign \g776/_0_  = _w109_ ;
	assign \g777/_0_  = _w110_ ;
	assign \g782/_0_  = _w113_ ;
	assign \g783/_0_  = _w116_ ;
	assign \g784/_0_  = _w119_ ;
	assign \g785/_0_  = _w122_ ;
	assign \g786/_0_  = _w125_ ;
	assign \g787/_0_  = _w128_ ;
	assign \g788/_0_  = _w131_ ;
	assign \g789/_0_  = _w134_ ;
	assign \g806/_0_  = _w135_ ;
endmodule;