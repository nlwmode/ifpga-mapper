module top( \1_pad  , \2_pad  , \3_pad  , \4_pad  , \5_pad  , \6_pad  , \7_pad  , \8_pad  , \44_pad  , \45_pad  , \46_pad  , \47_pad  , \48_pad  , \49_pad  , \50_pad  , \51_pad  );
  input \1_pad  ;
  input \2_pad  ;
  input \3_pad  ;
  input \4_pad  ;
  input \5_pad  ;
  input \6_pad  ;
  input \7_pad  ;
  input \8_pad  ;
  output \44_pad  ;
  output \45_pad  ;
  output \46_pad  ;
  output \47_pad  ;
  output \48_pad  ;
  output \49_pad  ;
  output \50_pad  ;
  output \51_pad  ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 ;
  assign n9 = \7_pad  & \8_pad  ;
  assign n10 = ~\1_pad  & \3_pad  ;
  assign n11 = \1_pad  & ~\3_pad  ;
  assign n12 = ~n10 & ~n11 ;
  assign n13 = ~\4_pad  & ~n12 ;
  assign n16 = ~n9 & ~n13 ;
  assign n17 = ~\1_pad  & ~\2_pad  ;
  assign n18 = \1_pad  & \2_pad  ;
  assign n19 = ~n17 & ~n18 ;
  assign n20 = \3_pad  & n19 ;
  assign n21 = ~\1_pad  & ~\3_pad  ;
  assign n22 = ~\4_pad  & ~n21 ;
  assign n23 = ~n20 & n22 ;
  assign n24 = \6_pad  & n23 ;
  assign n25 = n9 & ~n24 ;
  assign n26 = ~n16 & ~n25 ;
  assign n14 = n9 & ~n13 ;
  assign n15 = ~\6_pad  & ~n14 ;
  assign n27 = ~\3_pad  & ~n19 ;
  assign n28 = \4_pad  & ~n10 ;
  assign n29 = ~n27 & n28 ;
  assign n30 = ~n15 & ~n29 ;
  assign n31 = ~n26 & n30 ;
  assign n32 = ~n20 & ~n27 ;
  assign n33 = \4_pad  & n32 ;
  assign n34 = ~\6_pad  & n16 ;
  assign n35 = ~n33 & n34 ;
  assign n36 = ~n31 & ~n35 ;
  assign n37 = ~\5_pad  & ~n36 ;
  assign n38 = \4_pad  & n12 ;
  assign n41 = ~\4_pad  & n32 ;
  assign n42 = \8_pad  & n41 ;
  assign n39 = ~\7_pad  & ~n23 ;
  assign n40 = ~\8_pad  & ~n39 ;
  assign n43 = \6_pad  & ~n40 ;
  assign n44 = ~n42 & n43 ;
  assign n46 = \6_pad  & n41 ;
  assign n45 = ~\6_pad  & n23 ;
  assign n47 = \7_pad  & ~n45 ;
  assign n48 = ~n46 & n47 ;
  assign n49 = ~n44 & ~n48 ;
  assign n50 = ~n38 & ~n49 ;
  assign n51 = ~\6_pad  & ~n29 ;
  assign n52 = n39 & n51 ;
  assign n53 = ~n50 & ~n52 ;
  assign n54 = \5_pad  & ~n53 ;
  assign n55 = ~n37 & ~n54 ;
  assign n57 = \3_pad  & \5_pad  ;
  assign n60 = \3_pad  & \8_pad  ;
  assign n61 = ~\5_pad  & ~n60 ;
  assign n62 = \7_pad  & ~n61 ;
  assign n68 = ~n57 & ~n62 ;
  assign n69 = \4_pad  & ~n68 ;
  assign n56 = ~\3_pad  & ~\5_pad  ;
  assign n74 = ~\8_pad  & ~n56 ;
  assign n73 = ~\3_pad  & \7_pad  ;
  assign n75 = ~n57 & ~n73 ;
  assign n76 = n74 & n75 ;
  assign n70 = \4_pad  & \5_pad  ;
  assign n71 = \3_pad  & ~\5_pad  ;
  assign n72 = ~\7_pad  & n71 ;
  assign n77 = ~n70 & ~n72 ;
  assign n78 = ~n76 & n77 ;
  assign n79 = \6_pad  & ~n78 ;
  assign n80 = ~n69 & ~n79 ;
  assign n81 = ~\2_pad  & ~n80 ;
  assign n63 = \2_pad  & ~n62 ;
  assign n64 = \4_pad  & ~n63 ;
  assign n58 = ~\6_pad  & ~n57 ;
  assign n59 = ~n56 & ~n58 ;
  assign n65 = \2_pad  & ~\4_pad  ;
  assign n66 = ~n59 & ~n65 ;
  assign n67 = ~n64 & n66 ;
  assign n82 = ~\3_pad  & ~\8_pad  ;
  assign n83 = \5_pad  & ~n82 ;
  assign n84 = ~n62 & ~n83 ;
  assign n85 = ~n58 & n65 ;
  assign n86 = ~n84 & n85 ;
  assign n87 = ~n67 & ~n86 ;
  assign n88 = ~n81 & n87 ;
  assign n98 = ~\7_pad  & \8_pad  ;
  assign n99 = ~\4_pad  & n98 ;
  assign n100 = ~n70 & ~n99 ;
  assign n101 = ~\3_pad  & ~n100 ;
  assign n102 = \4_pad  & n71 ;
  assign n103 = ~n101 & ~n102 ;
  assign n104 = \6_pad  & ~n103 ;
  assign n89 = ~\4_pad  & ~\8_pad  ;
  assign n90 = \6_pad  & ~n89 ;
  assign n91 = \4_pad  & n9 ;
  assign n92 = n56 & ~n91 ;
  assign n93 = ~\4_pad  & ~\6_pad  ;
  assign n94 = \7_pad  & ~n93 ;
  assign n95 = n57 & ~n94 ;
  assign n96 = ~n92 & ~n95 ;
  assign n97 = ~n90 & ~n96 ;
  assign n105 = ~n57 & ~n93 ;
  assign n106 = n62 & n105 ;
  assign n107 = ~n97 & ~n106 ;
  assign n108 = ~n104 & n107 ;
  assign n109 = \4_pad  & \6_pad  ;
  assign n110 = ~\7_pad  & ~n93 ;
  assign n111 = ~n109 & n110 ;
  assign n112 = ~\4_pad  & ~\5_pad  ;
  assign n113 = ~n70 & ~n112 ;
  assign n115 = ~\6_pad  & ~n113 ;
  assign n114 = \6_pad  & n113 ;
  assign n116 = \7_pad  & ~n114 ;
  assign n117 = ~n115 & n116 ;
  assign n118 = ~n111 & ~n117 ;
  assign n119 = ~\8_pad  & ~n118 ;
  assign n120 = ~n93 & ~n109 ;
  assign n121 = \7_pad  & ~n120 ;
  assign n122 = n110 & ~n114 ;
  assign n123 = ~n121 & ~n122 ;
  assign n124 = \8_pad  & ~n123 ;
  assign n125 = ~n119 & ~n124 ;
  assign n126 = \7_pad  & ~\8_pad  ;
  assign n127 = \6_pad  & n98 ;
  assign n128 = ~n126 & ~n127 ;
  assign n129 = \5_pad  & ~n128 ;
  assign n130 = ~\5_pad  & n128 ;
  assign n131 = ~n129 & ~n130 ;
  assign n132 = ~\6_pad  & ~n98 ;
  assign n133 = ~n127 & ~n132 ;
  assign n134 = ~n98 & ~n126 ;
  assign \44_pad  = n55 ;
  assign \45_pad  = n88 ;
  assign \46_pad  = n108 ;
  assign \47_pad  = ~n125 ;
  assign \48_pad  = n131 ;
  assign \49_pad  = n133 ;
  assign \50_pad  = ~n134 ;
  assign \51_pad  = ~\8_pad  ;
endmodule
