module top( \a0_pad  , \a1_pad  , \a2_pad  , \a3_pad  , \a4_pad  , \b0_pad  , \b1_pad  , \b2_pad  , \b3_pad  , \b4_pad  , b_pad , \c0_pad  , \c1_pad  , \c2_pad  , \c3_pad  , \c4_pad  , c_pad , \d0_pad  , \d1_pad  , \d2_pad  , \d3_pad  , \d4_pad  , d_pad , \e0_pad  , \e1_pad  , \e2_pad  , \e3_pad  , \e4_pad  , e_pad , \f0_pad  , \f1_pad  , \f2_pad  , \f3_pad  , \f4_pad  , f_pad , \g0_pad  , \g1_pad  , \g2_pad  , \g3_pad  , \g4_pad  , g_pad , \h0_pad  , \h1_pad  , \h2_pad  , \h3_pad  , \h4_pad  , h_pad , \i0_pad  , \i1_pad  , \i2_pad  , \i3_pad  , i_pad , \j0_pad  , \j1_pad  , \j2_pad  , \j3_pad  , j_pad , \k0_pad  , \k1_pad  , \k2_pad  , \k3_pad  , k_pad , \l0_pad  , \l1_pad  , \l2_pad  , \l3_pad  , l_pad , \m0_pad  , \m1_pad  , \m2_pad  , \m3_pad  , m_pad , \n0_pad  , \n1_pad  , \n2_pad  , \n3_pad  , n_pad , \o0_pad  , \o1_pad  , \o2_pad  , \o3_pad  , o_pad , \p1_pad  , \p2_pad  , \p3_pad  , p_pad , \q1_pad  , \q2_pad  , \q3_pad  , q_pad , \r0_pad  , \r1_pad  , \r2_pad  , \r3_pad  , r_pad , \s0_pad  , \s1_pad  , \s2_pad  , \s3_pad  , s_pad , \t0_pad  , \t1_pad  , \t2_pad  , \t3_pad  , t_pad , \u0_pad  , \u1_pad  , \u2_pad  , \u3_pad  , u_pad , \v0_pad  , \v1_pad  , \v2_pad  , \v3_pad  , v_pad , \w0_pad  , \w1_pad  , \w2_pad  , \w3_pad  , w_pad , \x0_pad  , \x1_pad  , \x2_pad  , \x3_pad  , x_pad , \y0_pad  , \y1_pad  , \y2_pad  , \y3_pad  , y_pad , \z0_pad  , \z1_pad  , \z2_pad  , \z3_pad  , z_pad , \a5_pad  , \a6_pad  , \a7_pad  , \a8_pad  , \b5_pad  , \b6_pad  , \b7_pad  , \b8_pad  , \c5_pad  , \c6_pad  , \c7_pad  , \c8_pad  , \d5_pad  , \d6_pad  , \d7_pad  , \e5_pad  , \e6_pad  , \e7_pad  , \f5_pad  , \f6_pad  , \f7_pad  , \g5_pad  , \g6_pad  , \g7_pad  , \h5_pad  , \h6_pad  , \h7_pad  , \i4_pad  , \i5_pad  , \i6_pad  , \i7_pad  , \j4_pad  , \j5_pad  , \j6_pad  , \j7_pad  , \k4_pad  , \k5_pad  , \k6_pad  , \k7_pad  , \l4_pad  , \l5_pad  , \l6_pad  , \l7_pad  , \m4_pad  , \m5_pad  , \m6_pad  , \m7_pad  , \n4_pad  , \n5_pad  , \n6_pad  , \n7_pad  , \o4_pad  , \o5_pad  , \o6_pad  , \o7_pad  , \p4_pad  , \p5_pad  , \p6_pad  , \p7_pad  , \q4_pad  , \q5_pad  , \q6_pad  , \q7_pad  , \r4_pad  , \r5_pad  , \r6_pad  , \r7_pad  , \s4_pad  , \s5_pad  , \s6_pad  , \s7_pad  , \t4_pad  , \t5_pad  , \t6_pad  , \t7_pad  , \u4_pad  , \u5_pad  , \u6_pad  , \u7_pad  , \v4_pad  , \v5_pad  , \v6_pad  , \v7_pad  , \w4_pad  , \w5_pad  , \w6_pad  , \w7_pad  , \x4_pad  , \x5_pad  , \x6_pad  , \x7_pad  , \y4_pad  , \y5_pad  , \y6_pad  , \y7_pad  , \z4_pad  , \z5_pad  , \z6_pad  , \z7_pad  );
  input \a0_pad  ;
  input \a1_pad  ;
  input \a2_pad  ;
  input \a3_pad  ;
  input \a4_pad  ;
  input \b0_pad  ;
  input \b1_pad  ;
  input \b2_pad  ;
  input \b3_pad  ;
  input \b4_pad  ;
  input b_pad ;
  input \c0_pad  ;
  input \c1_pad  ;
  input \c2_pad  ;
  input \c3_pad  ;
  input \c4_pad  ;
  input c_pad ;
  input \d0_pad  ;
  input \d1_pad  ;
  input \d2_pad  ;
  input \d3_pad  ;
  input \d4_pad  ;
  input d_pad ;
  input \e0_pad  ;
  input \e1_pad  ;
  input \e2_pad  ;
  input \e3_pad  ;
  input \e4_pad  ;
  input e_pad ;
  input \f0_pad  ;
  input \f1_pad  ;
  input \f2_pad  ;
  input \f3_pad  ;
  input \f4_pad  ;
  input f_pad ;
  input \g0_pad  ;
  input \g1_pad  ;
  input \g2_pad  ;
  input \g3_pad  ;
  input \g4_pad  ;
  input g_pad ;
  input \h0_pad  ;
  input \h1_pad  ;
  input \h2_pad  ;
  input \h3_pad  ;
  input \h4_pad  ;
  input h_pad ;
  input \i0_pad  ;
  input \i1_pad  ;
  input \i2_pad  ;
  input \i3_pad  ;
  input i_pad ;
  input \j0_pad  ;
  input \j1_pad  ;
  input \j2_pad  ;
  input \j3_pad  ;
  input j_pad ;
  input \k0_pad  ;
  input \k1_pad  ;
  input \k2_pad  ;
  input \k3_pad  ;
  input k_pad ;
  input \l0_pad  ;
  input \l1_pad  ;
  input \l2_pad  ;
  input \l3_pad  ;
  input l_pad ;
  input \m0_pad  ;
  input \m1_pad  ;
  input \m2_pad  ;
  input \m3_pad  ;
  input m_pad ;
  input \n0_pad  ;
  input \n1_pad  ;
  input \n2_pad  ;
  input \n3_pad  ;
  input n_pad ;
  input \o0_pad  ;
  input \o1_pad  ;
  input \o2_pad  ;
  input \o3_pad  ;
  input o_pad ;
  input \p1_pad  ;
  input \p2_pad  ;
  input \p3_pad  ;
  input p_pad ;
  input \q1_pad  ;
  input \q2_pad  ;
  input \q3_pad  ;
  input q_pad ;
  input \r0_pad  ;
  input \r1_pad  ;
  input \r2_pad  ;
  input \r3_pad  ;
  input r_pad ;
  input \s0_pad  ;
  input \s1_pad  ;
  input \s2_pad  ;
  input \s3_pad  ;
  input s_pad ;
  input \t0_pad  ;
  input \t1_pad  ;
  input \t2_pad  ;
  input \t3_pad  ;
  input t_pad ;
  input \u0_pad  ;
  input \u1_pad  ;
  input \u2_pad  ;
  input \u3_pad  ;
  input u_pad ;
  input \v0_pad  ;
  input \v1_pad  ;
  input \v2_pad  ;
  input \v3_pad  ;
  input v_pad ;
  input \w0_pad  ;
  input \w1_pad  ;
  input \w2_pad  ;
  input \w3_pad  ;
  input w_pad ;
  input \x0_pad  ;
  input \x1_pad  ;
  input \x2_pad  ;
  input \x3_pad  ;
  input x_pad ;
  input \y0_pad  ;
  input \y1_pad  ;
  input \y2_pad  ;
  input \y3_pad  ;
  input y_pad ;
  input \z0_pad  ;
  input \z1_pad  ;
  input \z2_pad  ;
  input \z3_pad  ;
  input z_pad ;
  output \a5_pad  ;
  output \a6_pad  ;
  output \a7_pad  ;
  output \a8_pad  ;
  output \b5_pad  ;
  output \b6_pad  ;
  output \b7_pad  ;
  output \b8_pad  ;
  output \c5_pad  ;
  output \c6_pad  ;
  output \c7_pad  ;
  output \c8_pad  ;
  output \d5_pad  ;
  output \d6_pad  ;
  output \d7_pad  ;
  output \e5_pad  ;
  output \e6_pad  ;
  output \e7_pad  ;
  output \f5_pad  ;
  output \f6_pad  ;
  output \f7_pad  ;
  output \g5_pad  ;
  output \g6_pad  ;
  output \g7_pad  ;
  output \h5_pad  ;
  output \h6_pad  ;
  output \h7_pad  ;
  output \i4_pad  ;
  output \i5_pad  ;
  output \i6_pad  ;
  output \i7_pad  ;
  output \j4_pad  ;
  output \j5_pad  ;
  output \j6_pad  ;
  output \j7_pad  ;
  output \k4_pad  ;
  output \k5_pad  ;
  output \k6_pad  ;
  output \k7_pad  ;
  output \l4_pad  ;
  output \l5_pad  ;
  output \l6_pad  ;
  output \l7_pad  ;
  output \m4_pad  ;
  output \m5_pad  ;
  output \m6_pad  ;
  output \m7_pad  ;
  output \n4_pad  ;
  output \n5_pad  ;
  output \n6_pad  ;
  output \n7_pad  ;
  output \o4_pad  ;
  output \o5_pad  ;
  output \o6_pad  ;
  output \o7_pad  ;
  output \p4_pad  ;
  output \p5_pad  ;
  output \p6_pad  ;
  output \p7_pad  ;
  output \q4_pad  ;
  output \q5_pad  ;
  output \q6_pad  ;
  output \q7_pad  ;
  output \r4_pad  ;
  output \r5_pad  ;
  output \r6_pad  ;
  output \r7_pad  ;
  output \s4_pad  ;
  output \s5_pad  ;
  output \s6_pad  ;
  output \s7_pad  ;
  output \t4_pad  ;
  output \t5_pad  ;
  output \t6_pad  ;
  output \t7_pad  ;
  output \u4_pad  ;
  output \u5_pad  ;
  output \u6_pad  ;
  output \u7_pad  ;
  output \v4_pad  ;
  output \v5_pad  ;
  output \v6_pad  ;
  output \v7_pad  ;
  output \w4_pad  ;
  output \w5_pad  ;
  output \w6_pad  ;
  output \w7_pad  ;
  output \x4_pad  ;
  output \x5_pad  ;
  output \x6_pad  ;
  output \x7_pad  ;
  output \y4_pad  ;
  output \y5_pad  ;
  output \y6_pad  ;
  output \y7_pad  ;
  output \z4_pad  ;
  output \z5_pad  ;
  output \z6_pad  ;
  output \z7_pad  ;
  wire n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 ;
  assign n136 = i_pad & r_pad ;
  assign n138 = ~p_pad & n136 ;
  assign n137 = ~\f1_pad  & ~n136 ;
  assign n139 = ~\y1_pad  & ~n137 ;
  assign n140 = ~n138 & n139 ;
  assign n141 = \a4_pad  & \y3_pad  ;
  assign n142 = \z3_pad  & n141 ;
  assign n143 = \b4_pad  & n142 ;
  assign n144 = \c4_pad  & n143 ;
  assign n148 = ~\f4_pad  & \j0_pad  ;
  assign n146 = ~\d4_pad  & ~\h0_pad  ;
  assign n147 = \d4_pad  & \h0_pad  ;
  assign n156 = ~n146 & ~n147 ;
  assign n157 = ~n148 & n156 ;
  assign n152 = ~\g4_pad  & ~\k0_pad  ;
  assign n153 = \g4_pad  & \k0_pad  ;
  assign n154 = ~n152 & ~n153 ;
  assign n149 = ~\e4_pad  & ~\i0_pad  ;
  assign n150 = \e4_pad  & \i0_pad  ;
  assign n151 = ~n149 & ~n150 ;
  assign n145 = \f4_pad  & ~\j0_pad  ;
  assign n155 = \h4_pad  & ~n145 ;
  assign n158 = ~n151 & n155 ;
  assign n159 = ~n154 & n158 ;
  assign n160 = n157 & n159 ;
  assign n161 = n144 & n160 ;
  assign n162 = \d2_pad  & \l0_pad  ;
  assign n163 = ~\h0_pad  & ~\i0_pad  ;
  assign n164 = ~\j0_pad  & ~\k0_pad  ;
  assign n165 = n163 & n164 ;
  assign n166 = n162 & n165 ;
  assign n167 = ~n161 & ~n166 ;
  assign n168 = ~\a2_pad  & n167 ;
  assign n169 = \e2_pad  & ~n168 ;
  assign n171 = \f2_pad  & n169 ;
  assign n170 = ~\f2_pad  & ~n169 ;
  assign n172 = ~\n0_pad  & ~n170 ;
  assign n173 = ~n171 & n172 ;
  assign n174 = f_pad & h_pad ;
  assign n176 = ~\g3_pad  & n174 ;
  assign n175 = ~\f3_pad  & ~n174 ;
  assign n177 = ~\y1_pad  & ~n175 ;
  assign n178 = ~n176 & n177 ;
  assign n180 = ~\d4_pad  & n144 ;
  assign n181 = \e4_pad  & n180 ;
  assign n183 = \f4_pad  & n181 ;
  assign n179 = ~\l0_pad  & ~\n0_pad  ;
  assign n182 = ~\f4_pad  & ~n181 ;
  assign n184 = n179 & ~n182 ;
  assign n185 = ~n183 & n184 ;
  assign n187 = ~q_pad & n136 ;
  assign n186 = ~\g1_pad  & ~n136 ;
  assign n188 = ~\y1_pad  & ~n186 ;
  assign n189 = ~n187 & n188 ;
  assign n190 = \h2_pad  & ~\n0_pad  ;
  assign n192 = ~\h3_pad  & n174 ;
  assign n191 = ~\g3_pad  & ~n174 ;
  assign n193 = ~\y1_pad  & ~n191 ;
  assign n194 = ~n192 & n193 ;
  assign n196 = \g4_pad  & n183 ;
  assign n195 = ~\g4_pad  & ~n183 ;
  assign n197 = n179 & ~n195 ;
  assign n198 = ~n196 & n197 ;
  assign n199 = ~\b0_pad  & s_pad ;
  assign n201 = ~t_pad & n199 ;
  assign n200 = ~\h1_pad  & ~n199 ;
  assign n202 = ~\y1_pad  & ~n200 ;
  assign n203 = ~n201 & n202 ;
  assign n204 = \l0_pad  & ~\n0_pad  ;
  assign n206 = ~g_pad & n174 ;
  assign n205 = ~\h3_pad  & ~n174 ;
  assign n207 = ~\y1_pad  & ~n205 ;
  assign n208 = ~n206 & n207 ;
  assign n209 = ~\h4_pad  & ~n162 ;
  assign n210 = \g2_pad  & \h2_pad  ;
  assign n211 = b_pad & ~\n0_pad  ;
  assign n212 = ~n210 & n211 ;
  assign n213 = ~n209 & n212 ;
  assign n215 = ~u_pad & n199 ;
  assign n214 = ~\i1_pad  & ~n199 ;
  assign n216 = ~\y1_pad  & ~n214 ;
  assign n217 = ~n215 & n216 ;
  assign n222 = ~\o2_pad  & ~\p2_pad  ;
  assign n223 = \g0_pad  & n222 ;
  assign n218 = \j2_pad  & ~\p2_pad  ;
  assign n219 = \o2_pad  & ~n218 ;
  assign n220 = \l2_pad  & ~\m2_pad  ;
  assign n221 = \n2_pad  & n220 ;
  assign n224 = ~n219 & n221 ;
  assign n225 = ~n223 & n224 ;
  assign n226 = ~\x1_pad  & n225 ;
  assign n227 = ~\i2_pad  & ~n226 ;
  assign n228 = ~\y1_pad  & ~n227 ;
  assign n231 = ~\j2_pad  & ~\k2_pad  ;
  assign n232 = ~\x1_pad  & ~n231 ;
  assign n236 = \i3_pad  & ~n232 ;
  assign n233 = \j3_pad  & n232 ;
  assign n234 = ~c_pad & ~d_pad ;
  assign n235 = ~e_pad & n234 ;
  assign n237 = ~n233 & n235 ;
  assign n238 = ~n236 & n237 ;
  assign n240 = c_pad & ~d_pad ;
  assign n241 = ~e_pad & n240 ;
  assign n242 = ~\s2_pad  & n241 ;
  assign n229 = d_pad & ~e_pad ;
  assign n230 = ~\r0_pad  & n229 ;
  assign n239 = e_pad & ~\h1_pad  ;
  assign n243 = ~\y1_pad  & ~n239 ;
  assign n244 = ~n230 & n243 ;
  assign n245 = ~n242 & n244 ;
  assign n246 = ~n238 & n245 ;
  assign n248 = ~v_pad & n199 ;
  assign n247 = ~\j1_pad  & ~n199 ;
  assign n249 = ~\y1_pad  & ~n247 ;
  assign n250 = ~n248 & n249 ;
  assign n252 = ~\e0_pad  & ~\f0_pad  ;
  assign n253 = \g0_pad  & ~n252 ;
  assign n254 = ~\o2_pad  & ~n253 ;
  assign n255 = ~\p2_pad  & ~\x1_pad  ;
  assign n256 = n221 & n255 ;
  assign n257 = ~n254 & n256 ;
  assign n259 = ~\j2_pad  & ~n257 ;
  assign n251 = ~\j2_pad  & ~\o2_pad  ;
  assign n258 = ~n251 & n257 ;
  assign n260 = ~\y1_pad  & ~n258 ;
  assign n261 = ~n259 & n260 ;
  assign n264 = \j3_pad  & ~n232 ;
  assign n263 = \k3_pad  & n232 ;
  assign n265 = n235 & ~n263 ;
  assign n266 = ~n264 & n265 ;
  assign n268 = ~\t2_pad  & n241 ;
  assign n262 = ~\s0_pad  & n229 ;
  assign n267 = e_pad & ~\i1_pad  ;
  assign n269 = ~\y1_pad  & ~n267 ;
  assign n270 = ~n262 & n269 ;
  assign n271 = ~n268 & n270 ;
  assign n272 = ~n266 & n271 ;
  assign n274 = ~w_pad & n199 ;
  assign n273 = ~\k1_pad  & ~n199 ;
  assign n275 = ~\y1_pad  & ~n273 ;
  assign n276 = ~n274 & n275 ;
  assign n277 = \g0_pad  & n252 ;
  assign n278 = ~\p2_pad  & ~n277 ;
  assign n279 = ~\o2_pad  & ~\x1_pad  ;
  assign n280 = n221 & n279 ;
  assign n281 = ~n278 & n280 ;
  assign n283 = \k2_pad  & n281 ;
  assign n282 = ~\k2_pad  & ~n281 ;
  assign n284 = ~\y1_pad  & ~n282 ;
  assign n285 = ~n283 & n284 ;
  assign n288 = \k3_pad  & ~n232 ;
  assign n287 = \l3_pad  & n232 ;
  assign n289 = n235 & ~n287 ;
  assign n290 = ~n288 & n289 ;
  assign n292 = ~\u2_pad  & n241 ;
  assign n286 = ~\t0_pad  & n229 ;
  assign n291 = e_pad & ~\j1_pad  ;
  assign n293 = ~\y1_pad  & ~n291 ;
  assign n294 = ~n286 & n293 ;
  assign n295 = ~n292 & n294 ;
  assign n296 = ~n290 & n295 ;
  assign n298 = ~x_pad & n199 ;
  assign n297 = ~\l1_pad  & ~n199 ;
  assign n299 = ~\y1_pad  & ~n297 ;
  assign n300 = ~n298 & n299 ;
  assign n301 = \x1_pad  & n235 ;
  assign n303 = ~\l2_pad  & n301 ;
  assign n302 = \l2_pad  & ~n301 ;
  assign n304 = ~\y1_pad  & ~n302 ;
  assign n305 = ~n303 & n304 ;
  assign n308 = \l3_pad  & ~n232 ;
  assign n307 = \m3_pad  & n232 ;
  assign n309 = n235 & ~n307 ;
  assign n310 = ~n308 & n309 ;
  assign n312 = ~\v2_pad  & n241 ;
  assign n306 = ~\u0_pad  & n229 ;
  assign n311 = e_pad & ~\k1_pad  ;
  assign n313 = ~\y1_pad  & ~n311 ;
  assign n314 = ~n306 & n313 ;
  assign n315 = ~n312 & n314 ;
  assign n316 = ~n310 & n315 ;
  assign n318 = ~y_pad & n199 ;
  assign n317 = ~\m1_pad  & ~n199 ;
  assign n319 = ~\y1_pad  & ~n317 ;
  assign n320 = ~n318 & n319 ;
  assign n322 = \m2_pad  & n302 ;
  assign n321 = ~\m2_pad  & ~n302 ;
  assign n323 = ~\y1_pad  & ~n321 ;
  assign n324 = ~n322 & n323 ;
  assign n327 = \m3_pad  & ~n232 ;
  assign n326 = \n3_pad  & n232 ;
  assign n328 = n235 & ~n326 ;
  assign n329 = ~n327 & n328 ;
  assign n331 = ~\w2_pad  & n241 ;
  assign n325 = ~\v0_pad  & n229 ;
  assign n330 = e_pad & ~\l1_pad  ;
  assign n332 = ~\y1_pad  & ~n330 ;
  assign n333 = ~n325 & n332 ;
  assign n334 = ~n331 & n333 ;
  assign n335 = ~n329 & n334 ;
  assign n336 = ~\a2_pad  & \x1_pad  ;
  assign n338 = ~z_pad & n199 ;
  assign n337 = ~\n1_pad  & ~n199 ;
  assign n339 = ~\y1_pad  & ~n337 ;
  assign n340 = ~n338 & n339 ;
  assign n342 = \n2_pad  & n322 ;
  assign n341 = ~\n2_pad  & ~n322 ;
  assign n343 = ~\y1_pad  & ~n341 ;
  assign n344 = ~n342 & n343 ;
  assign n347 = \n3_pad  & ~n232 ;
  assign n346 = \o3_pad  & n232 ;
  assign n348 = n235 & ~n346 ;
  assign n349 = ~n347 & n348 ;
  assign n351 = ~\x2_pad  & n241 ;
  assign n345 = ~\w0_pad  & n229 ;
  assign n350 = e_pad & ~\m1_pad  ;
  assign n352 = ~\y1_pad  & ~n350 ;
  assign n353 = ~n345 & n352 ;
  assign n354 = ~n351 & n353 ;
  assign n355 = ~n349 & n354 ;
  assign n356 = \i2_pad  & \r2_pad  ;
  assign n357 = \q2_pad  & ~\x1_pad  ;
  assign n358 = n356 & n357 ;
  assign n359 = ~\o0_pad  & ~n358 ;
  assign n360 = n235 & ~n359 ;
  assign n361 = ~\y1_pad  & ~n360 ;
  assign n363 = ~\a0_pad  & n199 ;
  assign n362 = ~\o1_pad  & ~n199 ;
  assign n364 = ~\y1_pad  & ~n362 ;
  assign n365 = ~n363 & n364 ;
  assign n367 = \o2_pad  & n342 ;
  assign n366 = ~\o2_pad  & ~n342 ;
  assign n368 = ~\y1_pad  & ~n366 ;
  assign n369 = ~n367 & n368 ;
  assign n372 = \o3_pad  & ~n232 ;
  assign n371 = \p3_pad  & n232 ;
  assign n373 = n235 & ~n371 ;
  assign n374 = ~n372 & n373 ;
  assign n376 = ~\y2_pad  & n241 ;
  assign n370 = ~\x0_pad  & n229 ;
  assign n375 = e_pad & ~\n1_pad  ;
  assign n377 = ~\y1_pad  & ~n375 ;
  assign n378 = ~n370 & n377 ;
  assign n379 = ~n376 & n378 ;
  assign n380 = ~n374 & n379 ;
  assign n381 = ~\q2_pad  & ~\r2_pad  ;
  assign n382 = \i2_pad  & ~n381 ;
  assign n383 = n231 & ~n382 ;
  assign n384 = ~\x1_pad  & ~n383 ;
  assign n403 = ~\j0_pad  & \l2_pad  ;
  assign n402 = ~\k0_pad  & ~\l2_pad  ;
  assign n404 = ~\n2_pad  & ~n402 ;
  assign n405 = ~n403 & n404 ;
  assign n406 = \m2_pad  & ~n405 ;
  assign n398 = ~\h0_pad  & \l2_pad  ;
  assign n397 = ~\i0_pad  & ~\l2_pad  ;
  assign n399 = \n2_pad  & ~n397 ;
  assign n400 = ~n398 & n399 ;
  assign n401 = ~\m2_pad  & ~n400 ;
  assign n407 = n222 & ~n401 ;
  assign n408 = ~n406 & n407 ;
  assign n409 = ~n384 & ~n408 ;
  assign n385 = \d0_pad  & \r2_pad  ;
  assign n386 = ~\q2_pad  & ~n385 ;
  assign n387 = \i2_pad  & ~n386 ;
  assign n388 = \i3_pad  & ~n356 ;
  assign n389 = ~n387 & ~n388 ;
  assign n391 = ~\c0_pad  & ~\r2_pad  ;
  assign n390 = \r2_pad  & ~\z1_pad  ;
  assign n392 = \i2_pad  & \q2_pad  ;
  assign n393 = ~n390 & n392 ;
  assign n394 = ~n391 & n393 ;
  assign n395 = ~n389 & ~n394 ;
  assign n396 = n384 & ~n395 ;
  assign n410 = ~\a2_pad  & ~\y1_pad  ;
  assign n411 = ~n396 & n410 ;
  assign n412 = ~n409 & n411 ;
  assign n414 = \e2_pad  & \f2_pad  ;
  assign n415 = \a2_pad  & ~n414 ;
  assign n416 = ~\d0_pad  & ~\e2_pad  ;
  assign n413 = \d0_pad  & ~\f2_pad  ;
  assign n417 = \m0_pad  & ~\y1_pad  ;
  assign n418 = ~n413 & n417 ;
  assign n419 = ~n416 & n418 ;
  assign n420 = n415 & n419 ;
  assign n421 = ~n412 & ~n420 ;
  assign n422 = \b0_pad  & s_pad ;
  assign n424 = ~t_pad & n422 ;
  assign n423 = ~\p1_pad  & ~n422 ;
  assign n425 = ~\y1_pad  & ~n423 ;
  assign n426 = ~n424 & n425 ;
  assign n428 = \p2_pad  & n367 ;
  assign n427 = ~\p2_pad  & ~n367 ;
  assign n429 = ~\y1_pad  & ~n427 ;
  assign n430 = ~n428 & n429 ;
  assign n433 = \p3_pad  & ~n232 ;
  assign n432 = \q3_pad  & n232 ;
  assign n434 = n235 & ~n432 ;
  assign n435 = ~n433 & n434 ;
  assign n437 = ~\z2_pad  & n241 ;
  assign n431 = ~\y0_pad  & n229 ;
  assign n436 = e_pad & ~\o1_pad  ;
  assign n438 = ~\y1_pad  & ~n436 ;
  assign n439 = ~n431 & n438 ;
  assign n440 = ~n437 & n439 ;
  assign n441 = ~n435 & n440 ;
  assign n442 = ~\c2_pad  & ~n210 ;
  assign n443 = ~\n0_pad  & ~n442 ;
  assign n445 = ~u_pad & n422 ;
  assign n444 = ~\q1_pad  & ~n422 ;
  assign n446 = ~\y1_pad  & ~n444 ;
  assign n447 = ~n445 & n446 ;
  assign n448 = ~\i2_pad  & ~n225 ;
  assign n449 = ~\x1_pad  & ~n448 ;
  assign n451 = ~\q2_pad  & ~n449 ;
  assign n450 = \q2_pad  & n449 ;
  assign n452 = ~\y1_pad  & ~n450 ;
  assign n453 = ~n451 & n452 ;
  assign n456 = \q3_pad  & ~n232 ;
  assign n455 = \r3_pad  & n232 ;
  assign n457 = n235 & ~n455 ;
  assign n458 = ~n456 & n457 ;
  assign n460 = ~\a3_pad  & n241 ;
  assign n454 = ~\z0_pad  & n229 ;
  assign n459 = e_pad & ~\p1_pad  ;
  assign n461 = ~\y1_pad  & ~n459 ;
  assign n462 = ~n454 & n461 ;
  assign n463 = ~n460 & n462 ;
  assign n464 = ~n458 & n463 ;
  assign n465 = i_pad & ~r_pad ;
  assign n467 = ~j_pad & n465 ;
  assign n466 = ~\r0_pad  & ~n465 ;
  assign n468 = ~\y1_pad  & ~n466 ;
  assign n469 = ~n467 & n468 ;
  assign n471 = ~v_pad & n422 ;
  assign n470 = ~\r1_pad  & ~n422 ;
  assign n472 = ~\y1_pad  & ~n470 ;
  assign n473 = ~n471 & n472 ;
  assign n475 = \r2_pad  & n450 ;
  assign n474 = ~\r2_pad  & ~n450 ;
  assign n476 = ~\y1_pad  & ~n474 ;
  assign n477 = ~n475 & n476 ;
  assign n480 = \r3_pad  & ~n232 ;
  assign n479 = \s3_pad  & n232 ;
  assign n481 = n235 & ~n479 ;
  assign n482 = ~n480 & n481 ;
  assign n484 = ~\b3_pad  & n241 ;
  assign n478 = ~\a1_pad  & n229 ;
  assign n483 = e_pad & ~\q1_pad  ;
  assign n485 = ~\y1_pad  & ~n483 ;
  assign n486 = ~n478 & n485 ;
  assign n487 = ~n484 & n486 ;
  assign n488 = ~n482 & n487 ;
  assign n490 = ~k_pad & n465 ;
  assign n489 = ~\s0_pad  & ~n465 ;
  assign n491 = ~\y1_pad  & ~n489 ;
  assign n492 = ~n490 & n491 ;
  assign n494 = ~w_pad & n422 ;
  assign n493 = ~\s1_pad  & ~n422 ;
  assign n495 = ~\y1_pad  & ~n493 ;
  assign n496 = ~n494 & n495 ;
  assign n497 = f_pad & ~h_pad ;
  assign n499 = ~\t2_pad  & n497 ;
  assign n498 = ~\s2_pad  & ~n497 ;
  assign n500 = ~\y1_pad  & ~n498 ;
  assign n501 = ~n499 & n500 ;
  assign n504 = \s3_pad  & ~n232 ;
  assign n503 = \t3_pad  & n232 ;
  assign n505 = n235 & ~n503 ;
  assign n506 = ~n504 & n505 ;
  assign n508 = ~\c3_pad  & n241 ;
  assign n502 = ~\b1_pad  & n229 ;
  assign n507 = e_pad & ~\r1_pad  ;
  assign n509 = ~\y1_pad  & ~n507 ;
  assign n510 = ~n502 & n509 ;
  assign n511 = ~n508 & n510 ;
  assign n512 = ~n506 & n511 ;
  assign n514 = ~l_pad & n465 ;
  assign n513 = ~\t0_pad  & ~n465 ;
  assign n515 = ~\y1_pad  & ~n513 ;
  assign n516 = ~n514 & n515 ;
  assign n518 = ~x_pad & n422 ;
  assign n517 = ~\t1_pad  & ~n422 ;
  assign n519 = ~\y1_pad  & ~n517 ;
  assign n520 = ~n518 & n519 ;
  assign n522 = ~\u2_pad  & n497 ;
  assign n521 = ~\t2_pad  & ~n497 ;
  assign n523 = ~\y1_pad  & ~n521 ;
  assign n524 = ~n522 & n523 ;
  assign n527 = \t3_pad  & ~n232 ;
  assign n526 = \u3_pad  & n232 ;
  assign n528 = n235 & ~n526 ;
  assign n529 = ~n527 & n528 ;
  assign n531 = ~\d3_pad  & n241 ;
  assign n525 = ~\c1_pad  & n229 ;
  assign n530 = e_pad & ~\s1_pad  ;
  assign n532 = ~\y1_pad  & ~n530 ;
  assign n533 = ~n525 & n532 ;
  assign n534 = ~n531 & n533 ;
  assign n535 = ~n529 & n534 ;
  assign n537 = ~m_pad & n465 ;
  assign n536 = ~\u0_pad  & ~n465 ;
  assign n538 = ~\y1_pad  & ~n536 ;
  assign n539 = ~n537 & n538 ;
  assign n541 = ~y_pad & n422 ;
  assign n540 = ~\u1_pad  & ~n422 ;
  assign n542 = ~\y1_pad  & ~n540 ;
  assign n543 = ~n541 & n542 ;
  assign n545 = ~\v2_pad  & n497 ;
  assign n544 = ~\u2_pad  & ~n497 ;
  assign n546 = ~\y1_pad  & ~n544 ;
  assign n547 = ~n545 & n546 ;
  assign n550 = \u3_pad  & ~n232 ;
  assign n549 = \v3_pad  & n232 ;
  assign n551 = n235 & ~n549 ;
  assign n552 = ~n550 & n551 ;
  assign n554 = ~\e3_pad  & n241 ;
  assign n548 = ~\d1_pad  & n229 ;
  assign n553 = e_pad & ~\t1_pad  ;
  assign n555 = ~\y1_pad  & ~n553 ;
  assign n556 = ~n548 & n555 ;
  assign n557 = ~n554 & n556 ;
  assign n558 = ~n552 & n557 ;
  assign n560 = ~n_pad & n465 ;
  assign n559 = ~\v0_pad  & ~n465 ;
  assign n561 = ~\y1_pad  & ~n559 ;
  assign n562 = ~n560 & n561 ;
  assign n564 = ~z_pad & n422 ;
  assign n563 = ~\v1_pad  & ~n422 ;
  assign n565 = ~\y1_pad  & ~n563 ;
  assign n566 = ~n564 & n565 ;
  assign n568 = ~\w2_pad  & n497 ;
  assign n567 = ~\v2_pad  & ~n497 ;
  assign n569 = ~\y1_pad  & ~n567 ;
  assign n570 = ~n568 & n569 ;
  assign n573 = \v3_pad  & ~n232 ;
  assign n572 = \w3_pad  & n232 ;
  assign n574 = n235 & ~n572 ;
  assign n575 = ~n573 & n574 ;
  assign n577 = ~\f3_pad  & n241 ;
  assign n571 = ~\e1_pad  & n229 ;
  assign n576 = e_pad & ~\u1_pad  ;
  assign n578 = ~\y1_pad  & ~n576 ;
  assign n579 = ~n571 & n578 ;
  assign n580 = ~n577 & n579 ;
  assign n581 = ~n575 & n580 ;
  assign n583 = ~o_pad & n465 ;
  assign n582 = ~\w0_pad  & ~n465 ;
  assign n584 = ~\y1_pad  & ~n582 ;
  assign n585 = ~n583 & n584 ;
  assign n587 = ~\a0_pad  & n422 ;
  assign n586 = ~\w1_pad  & ~n422 ;
  assign n588 = ~\y1_pad  & ~n586 ;
  assign n589 = ~n587 & n588 ;
  assign n591 = ~\x2_pad  & n497 ;
  assign n590 = ~\w2_pad  & ~n497 ;
  assign n592 = ~\y1_pad  & ~n590 ;
  assign n593 = ~n591 & n592 ;
  assign n596 = \w3_pad  & ~n232 ;
  assign n595 = \x3_pad  & n232 ;
  assign n597 = n235 & ~n595 ;
  assign n598 = ~n596 & n597 ;
  assign n600 = ~\g3_pad  & n241 ;
  assign n594 = ~\f1_pad  & n229 ;
  assign n599 = e_pad & ~\v1_pad  ;
  assign n601 = ~\y1_pad  & ~n599 ;
  assign n602 = ~n594 & n601 ;
  assign n603 = ~n600 & n602 ;
  assign n604 = ~n598 & n603 ;
  assign n606 = ~p_pad & n465 ;
  assign n605 = ~\x0_pad  & ~n465 ;
  assign n607 = ~\y1_pad  & ~n605 ;
  assign n608 = ~n606 & n607 ;
  assign n609 = ~\y1_pad  & ~n301 ;
  assign n611 = ~\y2_pad  & n497 ;
  assign n610 = ~\x2_pad  & ~n497 ;
  assign n612 = ~\y1_pad  & ~n610 ;
  assign n613 = ~n611 & n612 ;
  assign n615 = \x3_pad  & ~n232 ;
  assign n616 = n235 & ~n615 ;
  assign n617 = ~\h3_pad  & n241 ;
  assign n618 = ~\g1_pad  & n229 ;
  assign n614 = e_pad & ~\w1_pad  ;
  assign n619 = ~\y1_pad  & ~n614 ;
  assign n620 = ~n618 & n619 ;
  assign n621 = ~n617 & n620 ;
  assign n622 = ~n616 & n621 ;
  assign n624 = ~q_pad & n465 ;
  assign n623 = ~\y0_pad  & ~n465 ;
  assign n625 = ~\y1_pad  & ~n623 ;
  assign n626 = ~n624 & n625 ;
  assign n627 = ~\n0_pad  & ~n358 ;
  assign n629 = ~\z2_pad  & n497 ;
  assign n628 = ~\y2_pad  & ~n497 ;
  assign n630 = ~\y1_pad  & ~n628 ;
  assign n631 = ~n629 & n630 ;
  assign n632 = ~\y3_pad  & n179 ;
  assign n634 = ~j_pad & n136 ;
  assign n633 = ~\z0_pad  & ~n136 ;
  assign n635 = ~\y1_pad  & ~n633 ;
  assign n636 = ~n634 & n635 ;
  assign n637 = n383 & ~n408 ;
  assign n642 = ~n231 & ~n382 ;
  assign n643 = ~\i3_pad  & n642 ;
  assign n638 = ~\d0_pad  & \r2_pad  ;
  assign n639 = \c0_pad  & \q2_pad  ;
  assign n640 = ~n638 & ~n639 ;
  assign n641 = \i2_pad  & ~n640 ;
  assign n644 = ~\x1_pad  & ~n641 ;
  assign n645 = ~n643 & n644 ;
  assign n646 = ~n637 & n645 ;
  assign n647 = \z1_pad  & ~n646 ;
  assign n648 = ~n358 & ~n647 ;
  assign n649 = ~\y1_pad  & ~n648 ;
  assign n651 = n383 & n408 ;
  assign n650 = \i3_pad  & n642 ;
  assign n652 = \c0_pad  & ~n385 ;
  assign n653 = n387 & ~n652 ;
  assign n654 = ~n650 & ~n653 ;
  assign n655 = ~n651 & n654 ;
  assign n656 = ~\x1_pad  & ~\y1_pad  ;
  assign n657 = ~\z1_pad  & n656 ;
  assign n658 = ~n655 & n657 ;
  assign n659 = ~n649 & ~n658 ;
  assign n661 = ~g_pad & n497 ;
  assign n660 = ~\z2_pad  & ~n497 ;
  assign n662 = ~\y1_pad  & ~n660 ;
  assign n663 = ~n661 & n662 ;
  assign n665 = ~\y3_pad  & ~\z3_pad  ;
  assign n664 = \y3_pad  & \z3_pad  ;
  assign n666 = n179 & ~n664 ;
  assign n667 = ~n665 & n666 ;
  assign n669 = ~k_pad & n136 ;
  assign n668 = ~\a1_pad  & ~n136 ;
  assign n670 = ~\y1_pad  & ~n668 ;
  assign n671 = ~n669 & n670 ;
  assign n672 = n167 & ~n415 ;
  assign n673 = ~\y1_pad  & ~n672 ;
  assign n675 = ~\b3_pad  & n174 ;
  assign n674 = ~\a3_pad  & ~n174 ;
  assign n676 = ~\y1_pad  & ~n674 ;
  assign n677 = ~n675 & n676 ;
  assign n678 = ~\a4_pad  & ~n664 ;
  assign n679 = ~n142 & n179 ;
  assign n680 = ~n678 & n679 ;
  assign n682 = ~l_pad & n136 ;
  assign n681 = ~\b1_pad  & ~n136 ;
  assign n683 = ~\y1_pad  & ~n681 ;
  assign n684 = ~n682 & n683 ;
  assign n685 = \d4_pad  & n144 ;
  assign n686 = ~\e4_pad  & ~\f4_pad  ;
  assign n687 = ~\g4_pad  & n686 ;
  assign n688 = n685 & n687 ;
  assign n690 = ~\b2_pad  & ~n688 ;
  assign n689 = \b2_pad  & n688 ;
  assign n691 = n179 & ~n689 ;
  assign n692 = ~n690 & n691 ;
  assign n694 = ~\c3_pad  & n174 ;
  assign n693 = ~\b3_pad  & ~n174 ;
  assign n695 = ~\y1_pad  & ~n693 ;
  assign n696 = ~n694 & n695 ;
  assign n697 = ~\b4_pad  & ~n142 ;
  assign n698 = ~n143 & n179 ;
  assign n699 = ~n697 & n698 ;
  assign n701 = ~m_pad & n136 ;
  assign n700 = ~\c1_pad  & ~n136 ;
  assign n702 = ~\y1_pad  & ~n700 ;
  assign n703 = ~n701 & n702 ;
  assign n705 = \c2_pad  & n689 ;
  assign n704 = ~\c2_pad  & ~n689 ;
  assign n706 = n179 & ~n704 ;
  assign n707 = ~n705 & n706 ;
  assign n709 = ~\d3_pad  & n174 ;
  assign n708 = ~\c3_pad  & ~n174 ;
  assign n710 = ~\y1_pad  & ~n708 ;
  assign n711 = ~n709 & n710 ;
  assign n712 = ~\c4_pad  & ~n143 ;
  assign n713 = ~n144 & n179 ;
  assign n714 = ~n712 & n713 ;
  assign n716 = ~n_pad & n136 ;
  assign n715 = ~\d1_pad  & ~n136 ;
  assign n717 = ~\y1_pad  & ~n715 ;
  assign n718 = ~n716 & n717 ;
  assign n719 = ~\d2_pad  & ~\l0_pad  ;
  assign n720 = n212 & ~n719 ;
  assign n722 = ~\e3_pad  & n174 ;
  assign n721 = ~\d3_pad  & ~n174 ;
  assign n723 = ~\y1_pad  & ~n721 ;
  assign n724 = ~n722 & n723 ;
  assign n725 = ~\d4_pad  & ~n144 ;
  assign n726 = n179 & ~n685 ;
  assign n727 = ~n725 & n726 ;
  assign n729 = ~o_pad & n136 ;
  assign n728 = ~\e1_pad  & ~n136 ;
  assign n730 = ~\y1_pad  & ~n728 ;
  assign n731 = ~n729 & n730 ;
  assign n732 = ~\e2_pad  & n168 ;
  assign n733 = ~\n0_pad  & ~n169 ;
  assign n734 = ~n732 & n733 ;
  assign n736 = ~\f3_pad  & n174 ;
  assign n735 = ~\e3_pad  & ~n174 ;
  assign n737 = ~\y1_pad  & ~n735 ;
  assign n738 = ~n736 & n737 ;
  assign n739 = ~\e4_pad  & ~n180 ;
  assign n740 = n179 & ~n181 ;
  assign n741 = ~n739 & n740 ;
  assign \a5_pad  = n140 ;
  assign \a6_pad  = n173 ;
  assign \a7_pad  = n178 ;
  assign \a8_pad  = n185 ;
  assign \b5_pad  = n189 ;
  assign \b6_pad  = n190 ;
  assign \b7_pad  = n194 ;
  assign \b8_pad  = n198 ;
  assign \c5_pad  = n203 ;
  assign \c6_pad  = n204 ;
  assign \c7_pad  = n208 ;
  assign \c8_pad  = n213 ;
  assign \d5_pad  = n217 ;
  assign \d6_pad  = n228 ;
  assign \d7_pad  = n246 ;
  assign \e5_pad  = n250 ;
  assign \e6_pad  = n261 ;
  assign \e7_pad  = n272 ;
  assign \f5_pad  = n276 ;
  assign \f6_pad  = n285 ;
  assign \f7_pad  = n296 ;
  assign \g5_pad  = n300 ;
  assign \g6_pad  = n305 ;
  assign \g7_pad  = n316 ;
  assign \h5_pad  = n320 ;
  assign \h6_pad  = n324 ;
  assign \h7_pad  = n335 ;
  assign \i4_pad  = ~n336 ;
  assign \i5_pad  = n340 ;
  assign \i6_pad  = n344 ;
  assign \i7_pad  = n355 ;
  assign \j4_pad  = ~n361 ;
  assign \j5_pad  = n365 ;
  assign \j6_pad  = n369 ;
  assign \j7_pad  = n380 ;
  assign \k4_pad  = ~n421 ;
  assign \k5_pad  = n426 ;
  assign \k6_pad  = n430 ;
  assign \k7_pad  = n441 ;
  assign \l4_pad  = n443 ;
  assign \l5_pad  = n447 ;
  assign \l6_pad  = n453 ;
  assign \l7_pad  = n464 ;
  assign \m4_pad  = n469 ;
  assign \m5_pad  = n473 ;
  assign \m6_pad  = n477 ;
  assign \m7_pad  = n488 ;
  assign \n4_pad  = n492 ;
  assign \n5_pad  = n496 ;
  assign \n6_pad  = n501 ;
  assign \n7_pad  = n512 ;
  assign \o4_pad  = n516 ;
  assign \o5_pad  = n520 ;
  assign \o6_pad  = n524 ;
  assign \o7_pad  = n535 ;
  assign \p4_pad  = n539 ;
  assign \p5_pad  = n543 ;
  assign \p6_pad  = n547 ;
  assign \p7_pad  = n558 ;
  assign \q4_pad  = n562 ;
  assign \q5_pad  = n566 ;
  assign \q6_pad  = n570 ;
  assign \q7_pad  = n581 ;
  assign \r4_pad  = n585 ;
  assign \r5_pad  = n589 ;
  assign \r6_pad  = n593 ;
  assign \r7_pad  = n604 ;
  assign \s4_pad  = n608 ;
  assign \s5_pad  = ~n609 ;
  assign \s6_pad  = n613 ;
  assign \s7_pad  = n622 ;
  assign \t4_pad  = n626 ;
  assign \t5_pad  = ~n627 ;
  assign \t6_pad  = n631 ;
  assign \t7_pad  = n632 ;
  assign \u4_pad  = n636 ;
  assign \u5_pad  = ~n659 ;
  assign \u6_pad  = n663 ;
  assign \u7_pad  = n667 ;
  assign \v4_pad  = n671 ;
  assign \v5_pad  = n673 ;
  assign \v6_pad  = n677 ;
  assign \v7_pad  = n680 ;
  assign \w4_pad  = n684 ;
  assign \w5_pad  = n692 ;
  assign \w6_pad  = n696 ;
  assign \w7_pad  = n699 ;
  assign \x4_pad  = n703 ;
  assign \x5_pad  = n707 ;
  assign \x6_pad  = n711 ;
  assign \x7_pad  = n714 ;
  assign \y4_pad  = n718 ;
  assign \y5_pad  = n720 ;
  assign \y6_pad  = n724 ;
  assign \y7_pad  = n727 ;
  assign \z4_pad  = n731 ;
  assign \z5_pad  = n734 ;
  assign \z6_pad  = n738 ;
  assign \z7_pad  = n741 ;
endmodule
