module top (\C_0_pad , \C_10_pad , \C_11_pad , \C_12_pad , \C_13_pad , \C_14_pad , \C_15_pad , \C_16_pad , \C_1_pad , \C_2_pad , \C_3_pad , \C_4_pad , \C_5_pad , \C_6_pad , \C_7_pad , \C_8_pad , \C_9_pad , \P_0_pad , \X_10_reg/NET0131 , \X_11_reg/NET0131 , \X_12_reg/NET0131 , \X_13_reg/NET0131 , \X_14_reg/NET0131 , \X_15_reg/NET0131 , \X_16_reg/P0002 , \X_1_reg/NET0131 , \X_2_reg/NET0131 , \X_3_reg/NET0131 , \X_4_reg/NET0131 , \X_5_reg/NET0131 , \X_6_reg/NET0131 , \X_7_reg/NET0131 , \X_8_reg/NET0131 , \X_9_reg/NET0131 , \X_12_reg/P0001 , \X_13_reg/P0001 , \X_14_reg/P0001 , \X_15_reg/P0001 , \X_16_reg/P0000 , \X_9_reg/P0001 , Z_pad, \_al_n0 , \_al_n1 , \g1160/_3_ , \g1169/_0_ , \g1185/_0_ , \g1212/_2_ , \g1218/_0_ , \g1234/_0_ , \g16/_1_ , \g17/_0_ , \g27/_2_ , \g29/_3_ , \g669/_1__syn_2 , \g714/_0_ , \g721/_0_ , \g734/_0_ , \g743/_0_ , \g763/_0_ );
	input \C_0_pad  ;
	input \C_10_pad  ;
	input \C_11_pad  ;
	input \C_12_pad  ;
	input \C_13_pad  ;
	input \C_14_pad  ;
	input \C_15_pad  ;
	input \C_16_pad  ;
	input \C_1_pad  ;
	input \C_2_pad  ;
	input \C_3_pad  ;
	input \C_4_pad  ;
	input \C_5_pad  ;
	input \C_6_pad  ;
	input \C_7_pad  ;
	input \C_8_pad  ;
	input \C_9_pad  ;
	input \P_0_pad  ;
	input \X_10_reg/NET0131  ;
	input \X_11_reg/NET0131  ;
	input \X_12_reg/NET0131  ;
	input \X_13_reg/NET0131  ;
	input \X_14_reg/NET0131  ;
	input \X_15_reg/NET0131  ;
	input \X_16_reg/P0002  ;
	input \X_1_reg/NET0131  ;
	input \X_2_reg/NET0131  ;
	input \X_3_reg/NET0131  ;
	input \X_4_reg/NET0131  ;
	input \X_5_reg/NET0131  ;
	input \X_6_reg/NET0131  ;
	input \X_7_reg/NET0131  ;
	input \X_8_reg/NET0131  ;
	input \X_9_reg/NET0131  ;
	output \X_12_reg/P0001  ;
	output \X_13_reg/P0001  ;
	output \X_14_reg/P0001  ;
	output \X_15_reg/P0001  ;
	output \X_16_reg/P0000  ;
	output \X_9_reg/P0001  ;
	output Z_pad ;
	output \_al_n0  ;
	output \_al_n1  ;
	output \g1160/_3_  ;
	output \g1169/_0_  ;
	output \g1185/_0_  ;
	output \g1212/_2_  ;
	output \g1218/_0_  ;
	output \g1234/_0_  ;
	output \g16/_1_  ;
	output \g17/_0_  ;
	output \g27/_2_  ;
	output \g29/_3_  ;
	output \g669/_1__syn_2  ;
	output \g714/_0_  ;
	output \g721/_0_  ;
	output \g734/_0_  ;
	output \g743/_0_  ;
	output \g763/_0_  ;
	wire _w94_ ;
	wire _w93_ ;
	wire _w92_ ;
	wire _w91_ ;
	wire _w89_ ;
	wire _w87_ ;
	wire _w85_ ;
	wire _w83_ ;
	wire _w81_ ;
	wire _w80_ ;
	wire _w79_ ;
	wire _w78_ ;
	wire _w77_ ;
	wire _w76_ ;
	wire _w75_ ;
	wire _w74_ ;
	wire _w73_ ;
	wire _w72_ ;
	wire _w71_ ;
	wire _w70_ ;
	wire _w69_ ;
	wire _w68_ ;
	wire _w67_ ;
	wire _w66_ ;
	wire _w65_ ;
	wire _w48_ ;
	wire _w47_ ;
	wire _w46_ ;
	wire _w45_ ;
	wire _w43_ ;
	wire _w41_ ;
	wire _w44_ ;
	wire _w90_ ;
	wire _w31_ ;
	wire _w60_ ;
	wire _w42_ ;
	wire _w88_ ;
	wire _w29_ ;
	wire _w58_ ;
	wire _w86_ ;
	wire _w27_ ;
	wire _w56_ ;
	wire _w84_ ;
	wire _w25_ ;
	wire _w54_ ;
	wire _w82_ ;
	wire _w23_ ;
	wire _w52_ ;
	wire _w49_ ;
	wire _w50_ ;
	wire _w51_ ;
	wire _w53_ ;
	wire _w55_ ;
	wire _w57_ ;
	wire _w59_ ;
	wire _w61_ ;
	wire _w62_ ;
	wire _w63_ ;
	wire _w64_ ;
	LUT1 #(
		.INIT('h1)
	) name0 (
		\X_12_reg/NET0131 ,
		_w23_
	);
	LUT1 #(
		.INIT('h1)
	) name1 (
		\X_13_reg/NET0131 ,
		_w25_
	);
	LUT1 #(
		.INIT('h1)
	) name2 (
		\X_14_reg/NET0131 ,
		_w27_
	);
	LUT1 #(
		.INIT('h1)
	) name3 (
		\X_15_reg/NET0131 ,
		_w29_
	);
	LUT1 #(
		.INIT('h1)
	) name4 (
		\X_16_reg/P0002 ,
		_w31_
	);
	LUT1 #(
		.INIT('h1)
	) name5 (
		\X_9_reg/NET0131 ,
		_w41_
	);
	LUT4 #(
		.INIT('h535f)
	) name6 (
		\C_13_pad ,
		\C_14_pad ,
		\X_13_reg/NET0131 ,
		\X_14_reg/NET0131 ,
		_w42_
	);
	LUT4 #(
		.INIT('h535f)
	) name7 (
		\C_15_pad ,
		\C_16_pad ,
		\X_15_reg/NET0131 ,
		\X_16_reg/P0002 ,
		_w43_
	);
	LUT3 #(
		.INIT('h02)
	) name8 (
		\P_0_pad ,
		\X_13_reg/NET0131 ,
		\X_14_reg/NET0131 ,
		_w44_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name9 (
		\P_0_pad ,
		_w42_,
		_w43_,
		_w44_,
		_w45_
	);
	LUT4 #(
		.INIT('h0001)
	) name10 (
		\X_10_reg/NET0131 ,
		\X_11_reg/NET0131 ,
		\X_12_reg/NET0131 ,
		\X_9_reg/NET0131 ,
		_w46_
	);
	LUT3 #(
		.INIT('h02)
	) name11 (
		\P_0_pad ,
		\X_10_reg/NET0131 ,
		\X_9_reg/NET0131 ,
		_w47_
	);
	LUT2 #(
		.INIT('h8)
	) name12 (
		\C_11_pad ,
		\X_11_reg/NET0131 ,
		_w48_
	);
	LUT4 #(
		.INIT('h0080)
	) name13 (
		\C_10_pad ,
		\P_0_pad ,
		\X_10_reg/NET0131 ,
		\X_9_reg/NET0131 ,
		_w49_
	);
	LUT3 #(
		.INIT('h07)
	) name14 (
		_w47_,
		_w48_,
		_w49_,
		_w50_
	);
	LUT2 #(
		.INIT('h1)
	) name15 (
		\X_1_reg/NET0131 ,
		\X_2_reg/NET0131 ,
		_w51_
	);
	LUT4 #(
		.INIT('h0001)
	) name16 (
		\X_1_reg/NET0131 ,
		\X_2_reg/NET0131 ,
		\X_3_reg/NET0131 ,
		\X_4_reg/NET0131 ,
		_w52_
	);
	LUT3 #(
		.INIT('h01)
	) name17 (
		\X_5_reg/NET0131 ,
		\X_7_reg/NET0131 ,
		\X_8_reg/NET0131 ,
		_w53_
	);
	LUT3 #(
		.INIT('h40)
	) name18 (
		\X_6_reg/NET0131 ,
		_w52_,
		_w53_,
		_w54_
	);
	LUT4 #(
		.INIT('h4f00)
	) name19 (
		_w45_,
		_w46_,
		_w50_,
		_w54_,
		_w55_
	);
	LUT4 #(
		.INIT('h535f)
	) name20 (
		\C_3_pad ,
		\C_4_pad ,
		\X_3_reg/NET0131 ,
		\X_4_reg/NET0131 ,
		_w56_
	);
	LUT2 #(
		.INIT('h2)
	) name21 (
		_w51_,
		_w56_,
		_w57_
	);
	LUT4 #(
		.INIT('h535f)
	) name22 (
		\C_5_pad ,
		\C_6_pad ,
		\X_5_reg/NET0131 ,
		\X_6_reg/NET0131 ,
		_w58_
	);
	LUT3 #(
		.INIT('h20)
	) name23 (
		\C_2_pad ,
		\X_1_reg/NET0131 ,
		\X_2_reg/NET0131 ,
		_w59_
	);
	LUT3 #(
		.INIT('h15)
	) name24 (
		\C_0_pad ,
		\C_1_pad ,
		\X_1_reg/NET0131 ,
		_w60_
	);
	LUT4 #(
		.INIT('h0d00)
	) name25 (
		_w52_,
		_w58_,
		_w59_,
		_w60_,
		_w61_
	);
	LUT3 #(
		.INIT('h8a)
	) name26 (
		\P_0_pad ,
		_w57_,
		_w61_,
		_w62_
	);
	LUT3 #(
		.INIT('h80)
	) name27 (
		\C_9_pad ,
		\P_0_pad ,
		\X_9_reg/NET0131 ,
		_w63_
	);
	LUT3 #(
		.INIT('h20)
	) name28 (
		\C_12_pad ,
		\X_11_reg/NET0131 ,
		\X_12_reg/NET0131 ,
		_w64_
	);
	LUT3 #(
		.INIT('h13)
	) name29 (
		_w47_,
		_w63_,
		_w64_,
		_w65_
	);
	LUT4 #(
		.INIT('h535f)
	) name30 (
		\C_7_pad ,
		\C_8_pad ,
		\X_7_reg/NET0131 ,
		\X_8_reg/NET0131 ,
		_w66_
	);
	LUT2 #(
		.INIT('h2)
	) name31 (
		\P_0_pad ,
		\X_5_reg/NET0131 ,
		_w67_
	);
	LUT4 #(
		.INIT('h0400)
	) name32 (
		\X_6_reg/NET0131 ,
		_w52_,
		_w66_,
		_w67_,
		_w68_
	);
	LUT3 #(
		.INIT('h0d)
	) name33 (
		_w54_,
		_w65_,
		_w68_,
		_w69_
	);
	LUT3 #(
		.INIT('hef)
	) name34 (
		_w55_,
		_w62_,
		_w69_,
		_w70_
	);
	LUT2 #(
		.INIT('h8)
	) name35 (
		\X_7_reg/NET0131 ,
		\X_8_reg/NET0131 ,
		_w71_
	);
	LUT4 #(
		.INIT('h8000)
	) name36 (
		\P_0_pad ,
		\X_1_reg/NET0131 ,
		\X_2_reg/NET0131 ,
		\X_3_reg/NET0131 ,
		_w72_
	);
	LUT2 #(
		.INIT('h8)
	) name37 (
		\X_5_reg/NET0131 ,
		\X_6_reg/NET0131 ,
		_w73_
	);
	LUT4 #(
		.INIT('h8000)
	) name38 (
		\X_4_reg/NET0131 ,
		_w71_,
		_w72_,
		_w73_,
		_w74_
	);
	LUT3 #(
		.INIT('h80)
	) name39 (
		\X_10_reg/NET0131 ,
		\X_4_reg/NET0131 ,
		\X_9_reg/NET0131 ,
		_w75_
	);
	LUT4 #(
		.INIT('h8000)
	) name40 (
		\X_5_reg/NET0131 ,
		\X_6_reg/NET0131 ,
		\X_7_reg/NET0131 ,
		\X_8_reg/NET0131 ,
		_w76_
	);
	LUT3 #(
		.INIT('h80)
	) name41 (
		_w72_,
		_w75_,
		_w76_,
		_w77_
	);
	LUT4 #(
		.INIT('h8000)
	) name42 (
		\X_11_reg/NET0131 ,
		_w72_,
		_w75_,
		_w76_,
		_w78_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name43 (
		\X_11_reg/NET0131 ,
		_w72_,
		_w75_,
		_w76_,
		_w79_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name44 (
		\X_4_reg/NET0131 ,
		\X_7_reg/NET0131 ,
		_w72_,
		_w73_,
		_w80_
	);
	LUT2 #(
		.INIT('h6)
	) name45 (
		\X_7_reg/NET0131 ,
		\X_8_reg/NET0131 ,
		_w81_
	);
	LUT2 #(
		.INIT('h6)
	) name46 (
		_w80_,
		_w81_,
		_w82_
	);
	LUT2 #(
		.INIT('h8)
	) name47 (
		\X_12_reg/NET0131 ,
		_w78_,
		_w83_
	);
	LUT3 #(
		.INIT('h80)
	) name48 (
		\X_12_reg/NET0131 ,
		\X_13_reg/NET0131 ,
		_w78_,
		_w84_
	);
	LUT3 #(
		.INIT('h78)
	) name49 (
		\P_0_pad ,
		\X_1_reg/NET0131 ,
		\X_2_reg/NET0131 ,
		_w85_
	);
	LUT4 #(
		.INIT('h00ea)
	) name50 (
		\X_10_reg/NET0131 ,
		\X_9_reg/NET0131 ,
		_w74_,
		_w77_,
		_w86_
	);
	LUT4 #(
		.INIT('h8000)
	) name51 (
		\X_12_reg/NET0131 ,
		\X_13_reg/NET0131 ,
		\X_14_reg/NET0131 ,
		_w78_,
		_w87_
	);
	LUT4 #(
		.INIT('h78f0)
	) name52 (
		\X_4_reg/NET0131 ,
		\X_5_reg/NET0131 ,
		\X_6_reg/NET0131 ,
		_w72_,
		_w88_
	);
	LUT2 #(
		.INIT('h8)
	) name53 (
		\X_15_reg/NET0131 ,
		_w87_,
		_w89_
	);
	LUT2 #(
		.INIT('h6)
	) name54 (
		\X_4_reg/NET0131 ,
		_w72_,
		_w90_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name55 (
		\X_4_reg/NET0131 ,
		\X_7_reg/NET0131 ,
		_w72_,
		_w73_,
		_w91_
	);
	LUT3 #(
		.INIT('h6c)
	) name56 (
		\X_4_reg/NET0131 ,
		\X_5_reg/NET0131 ,
		_w72_,
		_w92_
	);
	LUT4 #(
		.INIT('h7f80)
	) name57 (
		\P_0_pad ,
		\X_1_reg/NET0131 ,
		\X_2_reg/NET0131 ,
		\X_3_reg/NET0131 ,
		_w93_
	);
	LUT2 #(
		.INIT('h6)
	) name58 (
		\P_0_pad ,
		\X_1_reg/NET0131 ,
		_w94_
	);
	assign \X_12_reg/P0001  = _w23_ ;
	assign \X_13_reg/P0001  = _w25_ ;
	assign \X_14_reg/P0001  = _w27_ ;
	assign \X_15_reg/P0001  = _w29_ ;
	assign \X_16_reg/P0000  = _w31_ ;
	assign \X_9_reg/P0001  = _w41_ ;
	assign Z_pad = _w70_ ;
	assign \_al_n0  = 1'b0;
	assign \_al_n1  = 1'b1;
	assign \g1160/_3_  = _w74_ ;
	assign \g1169/_0_  = _w79_ ;
	assign \g1185/_0_  = _w82_ ;
	assign \g1212/_2_  = _w84_ ;
	assign \g1218/_0_  = _w85_ ;
	assign \g1234/_0_  = _w86_ ;
	assign \g16/_1_  = _w87_ ;
	assign \g17/_0_  = _w88_ ;
	assign \g27/_2_  = _w83_ ;
	assign \g29/_3_  = _w78_ ;
	assign \g669/_1__syn_2  = _w89_ ;
	assign \g714/_0_  = _w90_ ;
	assign \g721/_0_  = _w91_ ;
	assign \g734/_0_  = _w92_ ;
	assign \g743/_0_  = _w93_ ;
	assign \g763/_0_  = _w94_ ;
endmodule;