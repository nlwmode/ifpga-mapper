module top (\G0_pad , \G10_pad , \G11_pad , \G12_pad , \G13_pad , \G1_pad , \G29_reg/NET0131 , \G2_pad , \G30_reg/NET0131 , \G31_reg/NET0131 , \G32_reg/NET0131 , \G33_reg/NET0131 , \G34_reg/NET0131 , \G35_reg/NET0131 , \G36_reg/NET0131 , \G37_reg/NET0131 , \G38_reg/NET0131 , \G39_reg/NET0131 , \G3_pad , \G40_reg/NET0131 , \G41_reg/NET0131 , \G42_reg/NET0131 , \G43_reg/NET0131 , \G44_reg/NET0131 , \G46_reg/NET0131 , \G4_pad , \G5_pad , \G6_pad , \G7_pad , \G8_pad , \G9_pad , \G530_pad , \G532_pad , \G542_pad , \G546_pad , \G547_pad , \G548_pad , \G549_pad , \G550_pad , \G551_pad , \G552_pad , \_al_n0 , \_al_n1 , \g1594/_3_ , \g1613/_0_ , \g1618/_0_ , \g1620/_2_ , \g1692/_0_ , \g1727/_0_ , \g1740/_0_ , \g1742/_0_ , \g1760/_0_ , \g1769/_3_ , \g1771/_0_ , \g1780/_0_ , \g1799/_0_ , \g1867/_0_ , \g1873/_0_ , \g1900/_0_ , \g1930/_0_ , \g1936/_0_ , \g2340/_2_ , \g2396/_1_ , \g2408/_0_ );
	input \G0_pad  ;
	input \G10_pad  ;
	input \G11_pad  ;
	input \G12_pad  ;
	input \G13_pad  ;
	input \G1_pad  ;
	input \G29_reg/NET0131  ;
	input \G2_pad  ;
	input \G30_reg/NET0131  ;
	input \G31_reg/NET0131  ;
	input \G32_reg/NET0131  ;
	input \G33_reg/NET0131  ;
	input \G34_reg/NET0131  ;
	input \G35_reg/NET0131  ;
	input \G36_reg/NET0131  ;
	input \G37_reg/NET0131  ;
	input \G38_reg/NET0131  ;
	input \G39_reg/NET0131  ;
	input \G3_pad  ;
	input \G40_reg/NET0131  ;
	input \G41_reg/NET0131  ;
	input \G42_reg/NET0131  ;
	input \G43_reg/NET0131  ;
	input \G44_reg/NET0131  ;
	input \G46_reg/NET0131  ;
	input \G4_pad  ;
	input \G5_pad  ;
	input \G6_pad  ;
	input \G7_pad  ;
	input \G8_pad  ;
	input \G9_pad  ;
	output \G530_pad  ;
	output \G532_pad  ;
	output \G542_pad  ;
	output \G546_pad  ;
	output \G547_pad  ;
	output \G548_pad  ;
	output \G549_pad  ;
	output \G550_pad  ;
	output \G551_pad  ;
	output \G552_pad  ;
	output \_al_n0  ;
	output \_al_n1  ;
	output \g1594/_3_  ;
	output \g1613/_0_  ;
	output \g1618/_0_  ;
	output \g1620/_2_  ;
	output \g1692/_0_  ;
	output \g1727/_0_  ;
	output \g1740/_0_  ;
	output \g1742/_0_  ;
	output \g1760/_0_  ;
	output \g1769/_3_  ;
	output \g1771/_0_  ;
	output \g1780/_0_  ;
	output \g1799/_0_  ;
	output \g1867/_0_  ;
	output \g1873/_0_  ;
	output \g1900/_0_  ;
	output \g1930/_0_  ;
	output \g1936/_0_  ;
	output \g2340/_2_  ;
	output \g2396/_1_  ;
	output \g2408/_0_  ;
	wire _w337_ ;
	wire _w336_ ;
	wire _w335_ ;
	wire _w334_ ;
	wire _w333_ ;
	wire _w332_ ;
	wire _w331_ ;
	wire _w330_ ;
	wire _w329_ ;
	wire _w328_ ;
	wire _w327_ ;
	wire _w326_ ;
	wire _w325_ ;
	wire _w324_ ;
	wire _w323_ ;
	wire _w322_ ;
	wire _w321_ ;
	wire _w320_ ;
	wire _w319_ ;
	wire _w318_ ;
	wire _w317_ ;
	wire _w316_ ;
	wire _w315_ ;
	wire _w314_ ;
	wire _w313_ ;
	wire _w312_ ;
	wire _w311_ ;
	wire _w310_ ;
	wire _w309_ ;
	wire _w308_ ;
	wire _w307_ ;
	wire _w306_ ;
	wire _w305_ ;
	wire _w304_ ;
	wire _w303_ ;
	wire _w302_ ;
	wire _w301_ ;
	wire _w300_ ;
	wire _w299_ ;
	wire _w298_ ;
	wire _w297_ ;
	wire _w296_ ;
	wire _w295_ ;
	wire _w294_ ;
	wire _w293_ ;
	wire _w292_ ;
	wire _w291_ ;
	wire _w290_ ;
	wire _w159_ ;
	wire _w158_ ;
	wire _w157_ ;
	wire _w156_ ;
	wire _w155_ ;
	wire _w154_ ;
	wire _w153_ ;
	wire _w152_ ;
	wire _w151_ ;
	wire _w149_ ;
	wire _w148_ ;
	wire _w147_ ;
	wire _w146_ ;
	wire _w145_ ;
	wire _w144_ ;
	wire _w143_ ;
	wire _w142_ ;
	wire _w141_ ;
	wire _w140_ ;
	wire _w139_ ;
	wire _w138_ ;
	wire _w137_ ;
	wire _w136_ ;
	wire _w135_ ;
	wire _w134_ ;
	wire _w133_ ;
	wire _w132_ ;
	wire _w131_ ;
	wire _w130_ ;
	wire _w129_ ;
	wire _w128_ ;
	wire _w127_ ;
	wire _w126_ ;
	wire _w125_ ;
	wire _w124_ ;
	wire _w123_ ;
	wire _w122_ ;
	wire _w121_ ;
	wire _w120_ ;
	wire _w119_ ;
	wire _w118_ ;
	wire _w117_ ;
	wire _w116_ ;
	wire _w115_ ;
	wire _w114_ ;
	wire _w113_ ;
	wire _w112_ ;
	wire _w111_ ;
	wire _w110_ ;
	wire _w109_ ;
	wire _w108_ ;
	wire _w107_ ;
	wire _w106_ ;
	wire _w105_ ;
	wire _w104_ ;
	wire _w103_ ;
	wire _w102_ ;
	wire _w101_ ;
	wire _w100_ ;
	wire _w99_ ;
	wire _w98_ ;
	wire _w97_ ;
	wire _w96_ ;
	wire _w95_ ;
	wire _w94_ ;
	wire _w93_ ;
	wire _w92_ ;
	wire _w61_ ;
	wire _w60_ ;
	wire _w59_ ;
	wire _w58_ ;
	wire _w57_ ;
	wire _w56_ ;
	wire _w55_ ;
	wire _w54_ ;
	wire _w53_ ;
	wire _w51_ ;
	wire _w50_ ;
	wire _w49_ ;
	wire _w48_ ;
	wire _w47_ ;
	wire _w46_ ;
	wire _w52_ ;
	wire _w150_ ;
	wire _w23_ ;
	wire _w280_ ;
	wire _w82_ ;
	wire _w36_ ;
	wire _w34_ ;
	wire _w35_ ;
	wire _w37_ ;
	wire _w38_ ;
	wire _w39_ ;
	wire _w40_ ;
	wire _w41_ ;
	wire _w42_ ;
	wire _w43_ ;
	wire _w44_ ;
	wire _w45_ ;
	wire _w62_ ;
	wire _w63_ ;
	wire _w64_ ;
	wire _w65_ ;
	wire _w66_ ;
	wire _w67_ ;
	wire _w68_ ;
	wire _w69_ ;
	wire _w70_ ;
	wire _w71_ ;
	wire _w72_ ;
	wire _w73_ ;
	wire _w74_ ;
	wire _w75_ ;
	wire _w76_ ;
	wire _w77_ ;
	wire _w78_ ;
	wire _w79_ ;
	wire _w80_ ;
	wire _w81_ ;
	wire _w83_ ;
	wire _w84_ ;
	wire _w85_ ;
	wire _w86_ ;
	wire _w87_ ;
	wire _w88_ ;
	wire _w89_ ;
	wire _w90_ ;
	wire _w91_ ;
	wire _w160_ ;
	wire _w161_ ;
	wire _w162_ ;
	wire _w163_ ;
	wire _w164_ ;
	wire _w165_ ;
	wire _w166_ ;
	wire _w167_ ;
	wire _w168_ ;
	wire _w169_ ;
	wire _w170_ ;
	wire _w171_ ;
	wire _w172_ ;
	wire _w173_ ;
	wire _w174_ ;
	wire _w175_ ;
	wire _w176_ ;
	wire _w177_ ;
	wire _w178_ ;
	wire _w179_ ;
	wire _w180_ ;
	wire _w181_ ;
	wire _w182_ ;
	wire _w183_ ;
	wire _w184_ ;
	wire _w185_ ;
	wire _w186_ ;
	wire _w187_ ;
	wire _w188_ ;
	wire _w189_ ;
	wire _w190_ ;
	wire _w191_ ;
	wire _w192_ ;
	wire _w193_ ;
	wire _w194_ ;
	wire _w195_ ;
	wire _w196_ ;
	wire _w197_ ;
	wire _w198_ ;
	wire _w199_ ;
	wire _w200_ ;
	wire _w201_ ;
	wire _w202_ ;
	wire _w203_ ;
	wire _w204_ ;
	wire _w205_ ;
	wire _w206_ ;
	wire _w207_ ;
	wire _w208_ ;
	wire _w209_ ;
	wire _w210_ ;
	wire _w211_ ;
	wire _w212_ ;
	wire _w213_ ;
	wire _w214_ ;
	wire _w215_ ;
	wire _w216_ ;
	wire _w217_ ;
	wire _w218_ ;
	wire _w219_ ;
	wire _w220_ ;
	wire _w221_ ;
	wire _w222_ ;
	wire _w223_ ;
	wire _w224_ ;
	wire _w225_ ;
	wire _w226_ ;
	wire _w227_ ;
	wire _w228_ ;
	wire _w229_ ;
	wire _w230_ ;
	wire _w231_ ;
	wire _w232_ ;
	wire _w233_ ;
	wire _w234_ ;
	wire _w235_ ;
	wire _w236_ ;
	wire _w237_ ;
	wire _w238_ ;
	wire _w239_ ;
	wire _w240_ ;
	wire _w241_ ;
	wire _w242_ ;
	wire _w243_ ;
	wire _w244_ ;
	wire _w245_ ;
	wire _w246_ ;
	wire _w247_ ;
	wire _w248_ ;
	wire _w249_ ;
	wire _w250_ ;
	wire _w251_ ;
	wire _w252_ ;
	wire _w253_ ;
	wire _w254_ ;
	wire _w255_ ;
	wire _w256_ ;
	wire _w257_ ;
	wire _w258_ ;
	wire _w259_ ;
	wire _w260_ ;
	wire _w261_ ;
	wire _w262_ ;
	wire _w263_ ;
	wire _w264_ ;
	wire _w265_ ;
	wire _w266_ ;
	wire _w267_ ;
	wire _w268_ ;
	wire _w269_ ;
	wire _w270_ ;
	wire _w271_ ;
	wire _w272_ ;
	wire _w273_ ;
	wire _w274_ ;
	wire _w275_ ;
	wire _w276_ ;
	wire _w277_ ;
	wire _w278_ ;
	wire _w279_ ;
	wire _w281_ ;
	wire _w282_ ;
	wire _w283_ ;
	wire _w284_ ;
	wire _w285_ ;
	wire _w286_ ;
	wire _w287_ ;
	wire _w288_ ;
	wire _w289_ ;
	LUT1 #(
		.INIT('h1)
	) name0 (
		\G41_reg/NET0131 ,
		_w23_
	);
	LUT2 #(
		.INIT('h2)
	) name1 (
		\G3_pad ,
		\G4_pad ,
		_w34_
	);
	LUT2 #(
		.INIT('h2)
	) name2 (
		\G11_pad ,
		\G5_pad ,
		_w35_
	);
	LUT3 #(
		.INIT('h08)
	) name3 (
		\G11_pad ,
		\G35_reg/NET0131 ,
		\G5_pad ,
		_w36_
	);
	LUT3 #(
		.INIT('h80)
	) name4 (
		\G2_pad ,
		_w34_,
		_w36_,
		_w37_
	);
	LUT2 #(
		.INIT('h1)
	) name5 (
		\G7_pad ,
		\G8_pad ,
		_w38_
	);
	LUT4 #(
		.INIT('h0001)
	) name6 (
		\G10_pad ,
		\G11_pad ,
		\G7_pad ,
		\G8_pad ,
		_w39_
	);
	LUT2 #(
		.INIT('h8)
	) name7 (
		\G10_pad ,
		\G7_pad ,
		_w40_
	);
	LUT3 #(
		.INIT('h80)
	) name8 (
		\G11_pad ,
		\G8_pad ,
		\G9_pad ,
		_w41_
	);
	LUT4 #(
		.INIT('h0777)
	) name9 (
		\G9_pad ,
		_w39_,
		_w40_,
		_w41_,
		_w42_
	);
	LUT2 #(
		.INIT('h8)
	) name10 (
		\G3_pad ,
		\G5_pad ,
		_w43_
	);
	LUT4 #(
		.INIT('h8000)
	) name11 (
		\G3_pad ,
		\G4_pad ,
		\G5_pad ,
		\G6_pad ,
		_w44_
	);
	LUT2 #(
		.INIT('h8)
	) name12 (
		\G2_pad ,
		_w44_,
		_w45_
	);
	LUT3 #(
		.INIT('h45)
	) name13 (
		_w37_,
		_w42_,
		_w45_,
		_w46_
	);
	LUT2 #(
		.INIT('h8)
	) name14 (
		\G10_pad ,
		\G9_pad ,
		_w47_
	);
	LUT4 #(
		.INIT('h0240)
	) name15 (
		\G10_pad ,
		\G7_pad ,
		\G8_pad ,
		\G9_pad ,
		_w48_
	);
	LUT4 #(
		.INIT('h8000)
	) name16 (
		\G11_pad ,
		\G4_pad ,
		\G5_pad ,
		\G6_pad ,
		_w49_
	);
	LUT3 #(
		.INIT('h02)
	) name17 (
		\G36_reg/NET0131 ,
		\G3_pad ,
		\G6_pad ,
		_w50_
	);
	LUT4 #(
		.INIT('h00bf)
	) name18 (
		\G3_pad ,
		_w48_,
		_w49_,
		_w50_,
		_w51_
	);
	LUT4 #(
		.INIT('hedbf)
	) name19 (
		\G10_pad ,
		\G7_pad ,
		\G8_pad ,
		\G9_pad ,
		_w52_
	);
	LUT3 #(
		.INIT('h80)
	) name20 (
		\G3_pad ,
		\G4_pad ,
		\G6_pad ,
		_w53_
	);
	LUT3 #(
		.INIT('h20)
	) name21 (
		_w35_,
		_w52_,
		_w53_,
		_w54_
	);
	LUT3 #(
		.INIT('h51)
	) name22 (
		\G2_pad ,
		_w51_,
		_w54_,
		_w55_
	);
	LUT3 #(
		.INIT('h40)
	) name23 (
		\G10_pad ,
		\G7_pad ,
		\G9_pad ,
		_w56_
	);
	LUT3 #(
		.INIT('h20)
	) name24 (
		\G30_reg/NET0131 ,
		\G7_pad ,
		\G8_pad ,
		_w57_
	);
	LUT4 #(
		.INIT('h000d)
	) name25 (
		_w40_,
		_w41_,
		_w56_,
		_w57_,
		_w58_
	);
	LUT3 #(
		.INIT('h51)
	) name26 (
		\G13_pad ,
		\G32_reg/NET0131 ,
		_w58_,
		_w59_
	);
	LUT2 #(
		.INIT('h1)
	) name27 (
		\G12_pad ,
		_w51_,
		_w60_
	);
	LUT4 #(
		.INIT('hd000)
	) name28 (
		_w46_,
		_w55_,
		_w59_,
		_w60_,
		_w61_
	);
	LUT2 #(
		.INIT('h8)
	) name29 (
		\G11_pad ,
		\G8_pad ,
		_w62_
	);
	LUT3 #(
		.INIT('h2e)
	) name30 (
		\G10_pad ,
		\G11_pad ,
		\G8_pad ,
		_w63_
	);
	LUT3 #(
		.INIT('h20)
	) name31 (
		\G30_reg/NET0131 ,
		\G6_pad ,
		\G7_pad ,
		_w64_
	);
	LUT2 #(
		.INIT('h8)
	) name32 (
		\G31_reg/NET0131 ,
		\G8_pad ,
		_w65_
	);
	LUT4 #(
		.INIT('h2a3f)
	) name33 (
		\G10_pad ,
		\G31_reg/NET0131 ,
		\G8_pad ,
		\G9_pad ,
		_w66_
	);
	LUT3 #(
		.INIT('h10)
	) name34 (
		_w63_,
		_w64_,
		_w66_,
		_w67_
	);
	LUT3 #(
		.INIT('h20)
	) name35 (
		\G10_pad ,
		\G8_pad ,
		\G9_pad ,
		_w68_
	);
	LUT4 #(
		.INIT('hc5ff)
	) name36 (
		\G10_pad ,
		\G31_reg/NET0131 ,
		\G8_pad ,
		\G9_pad ,
		_w69_
	);
	LUT2 #(
		.INIT('h1)
	) name37 (
		\G11_pad ,
		\G7_pad ,
		_w70_
	);
	LUT2 #(
		.INIT('h4)
	) name38 (
		_w69_,
		_w70_,
		_w71_
	);
	LUT4 #(
		.INIT('h0407)
	) name39 (
		\G0_pad ,
		\G3_pad ,
		\G4_pad ,
		\G5_pad ,
		_w72_
	);
	LUT2 #(
		.INIT('h2)
	) name40 (
		\G46_reg/NET0131 ,
		_w72_,
		_w73_
	);
	LUT2 #(
		.INIT('h2)
	) name41 (
		\G12_pad ,
		\G13_pad ,
		_w74_
	);
	LUT3 #(
		.INIT('h02)
	) name42 (
		\G11_pad ,
		\G30_reg/NET0131 ,
		\G6_pad ,
		_w75_
	);
	LUT2 #(
		.INIT('h2)
	) name43 (
		\G11_pad ,
		\G9_pad ,
		_w76_
	);
	LUT4 #(
		.INIT('h0002)
	) name44 (
		\G11_pad ,
		\G7_pad ,
		\G8_pad ,
		\G9_pad ,
		_w77_
	);
	LUT3 #(
		.INIT('h02)
	) name45 (
		_w74_,
		_w75_,
		_w77_,
		_w78_
	);
	LUT4 #(
		.INIT('h1000)
	) name46 (
		_w67_,
		_w71_,
		_w73_,
		_w78_,
		_w79_
	);
	LUT4 #(
		.INIT('h44c4)
	) name47 (
		\G0_pad ,
		\G1_pad ,
		\G3_pad ,
		\G4_pad ,
		_w80_
	);
	LUT3 #(
		.INIT('h4c)
	) name48 (
		\G3_pad ,
		\G4_pad ,
		\G5_pad ,
		_w81_
	);
	LUT4 #(
		.INIT('h8a0f)
	) name49 (
		\G1_pad ,
		\G3_pad ,
		\G4_pad ,
		\G5_pad ,
		_w82_
	);
	LUT3 #(
		.INIT('he0)
	) name50 (
		\G0_pad ,
		\G1_pad ,
		\G2_pad ,
		_w83_
	);
	LUT3 #(
		.INIT('hb0)
	) name51 (
		_w80_,
		_w82_,
		_w83_,
		_w84_
	);
	LUT2 #(
		.INIT('h8)
	) name52 (
		_w79_,
		_w84_,
		_w85_
	);
	LUT2 #(
		.INIT('he)
	) name53 (
		_w61_,
		_w85_,
		_w86_
	);
	LUT2 #(
		.INIT('h8)
	) name54 (
		\G1_pad ,
		\G3_pad ,
		_w87_
	);
	LUT3 #(
		.INIT('h80)
	) name55 (
		\G1_pad ,
		\G3_pad ,
		\G5_pad ,
		_w88_
	);
	LUT3 #(
		.INIT('h80)
	) name56 (
		\G2_pad ,
		\G4_pad ,
		\G6_pad ,
		_w89_
	);
	LUT2 #(
		.INIT('h8)
	) name57 (
		_w88_,
		_w89_,
		_w90_
	);
	LUT2 #(
		.INIT('h4)
	) name58 (
		_w42_,
		_w90_,
		_w91_
	);
	LUT3 #(
		.INIT('h20)
	) name59 (
		\G13_pad ,
		_w42_,
		_w90_,
		_w92_
	);
	LUT4 #(
		.INIT('h4000)
	) name60 (
		\G1_pad ,
		\G3_pad ,
		\G4_pad ,
		\G6_pad ,
		_w93_
	);
	LUT2 #(
		.INIT('h4)
	) name61 (
		\G4_pad ,
		\G6_pad ,
		_w94_
	);
	LUT4 #(
		.INIT('hb7ff)
	) name62 (
		\G1_pad ,
		\G3_pad ,
		\G4_pad ,
		\G6_pad ,
		_w95_
	);
	LUT3 #(
		.INIT('h04)
	) name63 (
		\G10_pad ,
		\G7_pad ,
		\G9_pad ,
		_w96_
	);
	LUT2 #(
		.INIT('h2)
	) name64 (
		\G11_pad ,
		\G7_pad ,
		_w97_
	);
	LUT4 #(
		.INIT('h135f)
	) name65 (
		_w62_,
		_w68_,
		_w96_,
		_w97_,
		_w98_
	);
	LUT4 #(
		.INIT('h4000)
	) name66 (
		\G10_pad ,
		\G11_pad ,
		\G8_pad ,
		\G9_pad ,
		_w99_
	);
	LUT3 #(
		.INIT('h40)
	) name67 (
		\G7_pad ,
		_w93_,
		_w99_,
		_w100_
	);
	LUT3 #(
		.INIT('h04)
	) name68 (
		\G10_pad ,
		\G7_pad ,
		\G8_pad ,
		_w101_
	);
	LUT2 #(
		.INIT('h1)
	) name69 (
		\G4_pad ,
		\G6_pad ,
		_w102_
	);
	LUT4 #(
		.INIT('h0004)
	) name70 (
		\G1_pad ,
		\G3_pad ,
		\G4_pad ,
		\G6_pad ,
		_w103_
	);
	LUT3 #(
		.INIT('h80)
	) name71 (
		_w76_,
		_w101_,
		_w103_,
		_w104_
	);
	LUT4 #(
		.INIT('h000e)
	) name72 (
		_w95_,
		_w98_,
		_w100_,
		_w104_,
		_w105_
	);
	LUT2 #(
		.INIT('h2)
	) name73 (
		\G2_pad ,
		\G5_pad ,
		_w106_
	);
	LUT3 #(
		.INIT('h08)
	) name74 (
		\G13_pad ,
		\G2_pad ,
		\G5_pad ,
		_w107_
	);
	LUT4 #(
		.INIT('h1011)
	) name75 (
		_w53_,
		_w92_,
		_w105_,
		_w107_,
		_w108_
	);
	LUT4 #(
		.INIT('h0800)
	) name76 (
		\G10_pad ,
		\G11_pad ,
		\G8_pad ,
		\G9_pad ,
		_w109_
	);
	LUT4 #(
		.INIT('hba00)
	) name77 (
		_w92_,
		_w105_,
		_w107_,
		_w109_,
		_w110_
	);
	LUT4 #(
		.INIT('h5100)
	) name78 (
		\G13_pad ,
		\G32_reg/NET0131 ,
		_w58_,
		_w109_,
		_w111_
	);
	LUT3 #(
		.INIT('hd0)
	) name79 (
		_w46_,
		_w55_,
		_w111_,
		_w112_
	);
	LUT3 #(
		.INIT('h54)
	) name80 (
		_w108_,
		_w110_,
		_w112_,
		_w113_
	);
	LUT2 #(
		.INIT('h8)
	) name81 (
		\G5_pad ,
		\G9_pad ,
		_w114_
	);
	LUT3 #(
		.INIT('h80)
	) name82 (
		\G6_pad ,
		_w39_,
		_w114_,
		_w115_
	);
	LUT2 #(
		.INIT('h8)
	) name83 (
		_w48_,
		_w94_,
		_w116_
	);
	LUT2 #(
		.INIT('h1)
	) name84 (
		_w115_,
		_w116_,
		_w117_
	);
	LUT4 #(
		.INIT('h00ba)
	) name85 (
		_w92_,
		_w105_,
		_w107_,
		_w117_,
		_w118_
	);
	LUT4 #(
		.INIT('h00d0)
	) name86 (
		_w46_,
		_w55_,
		_w59_,
		_w117_,
		_w119_
	);
	LUT3 #(
		.INIT('h23)
	) name87 (
		\G4_pad ,
		\G5_pad ,
		\G6_pad ,
		_w120_
	);
	LUT2 #(
		.INIT('h4)
	) name88 (
		\G1_pad ,
		\G2_pad ,
		_w121_
	);
	LUT2 #(
		.INIT('h4)
	) name89 (
		_w120_,
		_w121_,
		_w122_
	);
	LUT2 #(
		.INIT('h4)
	) name90 (
		_w58_,
		_w122_,
		_w123_
	);
	LUT4 #(
		.INIT('h20a0)
	) name91 (
		\G3_pad ,
		\G4_pad ,
		\G5_pad ,
		\G6_pad ,
		_w124_
	);
	LUT2 #(
		.INIT('h4)
	) name92 (
		\G2_pad ,
		\G3_pad ,
		_w125_
	);
	LUT3 #(
		.INIT('h40)
	) name93 (
		\G2_pad ,
		\G3_pad ,
		\G6_pad ,
		_w126_
	);
	LUT2 #(
		.INIT('h2)
	) name94 (
		\G4_pad ,
		\G5_pad ,
		_w127_
	);
	LUT3 #(
		.INIT('h04)
	) name95 (
		\G3_pad ,
		\G4_pad ,
		\G5_pad ,
		_w128_
	);
	LUT3 #(
		.INIT('h01)
	) name96 (
		_w124_,
		_w126_,
		_w128_,
		_w129_
	);
	LUT3 #(
		.INIT('h20)
	) name97 (
		\G2_pad ,
		\G3_pad ,
		\G6_pad ,
		_w130_
	);
	LUT4 #(
		.INIT('h4c00)
	) name98 (
		\G3_pad ,
		\G4_pad ,
		\G5_pad ,
		\G6_pad ,
		_w131_
	);
	LUT4 #(
		.INIT('h00b8)
	) name99 (
		\G2_pad ,
		\G4_pad ,
		\G5_pad ,
		\G6_pad ,
		_w132_
	);
	LUT3 #(
		.INIT('h01)
	) name100 (
		_w130_,
		_w131_,
		_w132_,
		_w133_
	);
	LUT4 #(
		.INIT('h0222)
	) name101 (
		\G1_pad ,
		_w58_,
		_w129_,
		_w133_,
		_w134_
	);
	LUT2 #(
		.INIT('h2)
	) name102 (
		\G13_pad ,
		\G43_reg/NET0131 ,
		_w135_
	);
	LUT3 #(
		.INIT('he0)
	) name103 (
		_w123_,
		_w134_,
		_w135_,
		_w136_
	);
	LUT4 #(
		.INIT('h5540)
	) name104 (
		\G3_pad ,
		_w49_,
		_w96_,
		_w102_,
		_w137_
	);
	LUT4 #(
		.INIT('h5100)
	) name105 (
		\G13_pad ,
		\G32_reg/NET0131 ,
		_w58_,
		_w137_,
		_w138_
	);
	LUT3 #(
		.INIT('hd0)
	) name106 (
		_w46_,
		_w55_,
		_w138_,
		_w139_
	);
	LUT4 #(
		.INIT('h0001)
	) name107 (
		_w118_,
		_w119_,
		_w136_,
		_w139_,
		_w140_
	);
	LUT3 #(
		.INIT('h40)
	) name108 (
		\G2_pad ,
		\G3_pad ,
		\G5_pad ,
		_w141_
	);
	LUT4 #(
		.INIT('h4000)
	) name109 (
		\G2_pad ,
		\G3_pad ,
		\G4_pad ,
		\G5_pad ,
		_w142_
	);
	LUT3 #(
		.INIT('h54)
	) name110 (
		\G2_pad ,
		\G3_pad ,
		\G5_pad ,
		_w143_
	);
	LUT3 #(
		.INIT('h70)
	) name111 (
		\G1_pad ,
		\G3_pad ,
		\G4_pad ,
		_w144_
	);
	LUT4 #(
		.INIT('h02a2)
	) name112 (
		\G1_pad ,
		\G2_pad ,
		\G3_pad ,
		\G4_pad ,
		_w145_
	);
	LUT4 #(
		.INIT('h0045)
	) name113 (
		_w142_,
		_w143_,
		_w144_,
		_w145_,
		_w146_
	);
	LUT2 #(
		.INIT('h2)
	) name114 (
		\G0_pad ,
		_w146_,
		_w147_
	);
	LUT2 #(
		.INIT('h8)
	) name115 (
		_w79_,
		_w147_,
		_w148_
	);
	LUT4 #(
		.INIT('hff45)
	) name116 (
		\G12_pad ,
		_w113_,
		_w140_,
		_w148_,
		_w149_
	);
	LUT2 #(
		.INIT('h8)
	) name117 (
		\G34_reg/NET0131 ,
		\G8_pad ,
		_w150_
	);
	LUT2 #(
		.INIT('h8)
	) name118 (
		_w56_,
		_w150_,
		_w151_
	);
	LUT4 #(
		.INIT('h4000)
	) name119 (
		\G10_pad ,
		\G6_pad ,
		\G7_pad ,
		\G9_pad ,
		_w152_
	);
	LUT3 #(
		.INIT('h13)
	) name120 (
		_w79_,
		_w151_,
		_w152_,
		_w153_
	);
	LUT3 #(
		.INIT('h2a)
	) name121 (
		\G34_reg/NET0131 ,
		\G8_pad ,
		\G9_pad ,
		_w154_
	);
	LUT2 #(
		.INIT('h8)
	) name122 (
		_w40_,
		_w154_,
		_w155_
	);
	LUT4 #(
		.INIT('h00ae)
	) name123 (
		\G10_pad ,
		\G7_pad ,
		\G8_pad ,
		\G9_pad ,
		_w156_
	);
	LUT4 #(
		.INIT('h20a0)
	) name124 (
		\G10_pad ,
		\G7_pad ,
		\G8_pad ,
		\G9_pad ,
		_w157_
	);
	LUT4 #(
		.INIT('haaa8)
	) name125 (
		\G6_pad ,
		_w109_,
		_w156_,
		_w157_,
		_w158_
	);
	LUT3 #(
		.INIT('h13)
	) name126 (
		_w79_,
		_w155_,
		_w158_,
		_w159_
	);
	LUT2 #(
		.INIT('h7)
	) name127 (
		_w153_,
		_w159_,
		_w160_
	);
	LUT4 #(
		.INIT('h2000)
	) name128 (
		\G10_pad ,
		\G6_pad ,
		\G7_pad ,
		\G9_pad ,
		_w161_
	);
	LUT2 #(
		.INIT('h2)
	) name129 (
		\G10_pad ,
		\G9_pad ,
		_w162_
	);
	LUT4 #(
		.INIT('h0e00)
	) name130 (
		\G10_pad ,
		\G11_pad ,
		\G7_pad ,
		\G8_pad ,
		_w163_
	);
	LUT3 #(
		.INIT('h20)
	) name131 (
		\G11_pad ,
		\G8_pad ,
		\G9_pad ,
		_w164_
	);
	LUT4 #(
		.INIT('h4500)
	) name132 (
		\G10_pad ,
		\G7_pad ,
		\G8_pad ,
		\G9_pad ,
		_w165_
	);
	LUT4 #(
		.INIT('h000b)
	) name133 (
		_w162_,
		_w163_,
		_w164_,
		_w165_,
		_w166_
	);
	LUT3 #(
		.INIT('h31)
	) name134 (
		\G6_pad ,
		_w161_,
		_w166_,
		_w167_
	);
	LUT3 #(
		.INIT('h13)
	) name135 (
		\G10_pad ,
		\G7_pad ,
		\G8_pad ,
		_w168_
	);
	LUT3 #(
		.INIT('h80)
	) name136 (
		\G10_pad ,
		\G7_pad ,
		\G8_pad ,
		_w169_
	);
	LUT2 #(
		.INIT('h8)
	) name137 (
		\G34_reg/NET0131 ,
		\G9_pad ,
		_w170_
	);
	LUT3 #(
		.INIT('h10)
	) name138 (
		_w168_,
		_w169_,
		_w170_,
		_w171_
	);
	LUT3 #(
		.INIT('hf2)
	) name139 (
		_w79_,
		_w167_,
		_w171_,
		_w172_
	);
	LUT4 #(
		.INIT('h6cb8)
	) name140 (
		\G10_pad ,
		\G7_pad ,
		\G8_pad ,
		\G9_pad ,
		_w173_
	);
	LUT2 #(
		.INIT('h8)
	) name141 (
		\G11_pad ,
		\G34_reg/NET0131 ,
		_w174_
	);
	LUT2 #(
		.INIT('h8)
	) name142 (
		_w173_,
		_w174_,
		_w175_
	);
	LUT3 #(
		.INIT('hf4)
	) name143 (
		\G42_reg/NET0131 ,
		_w79_,
		_w175_,
		_w176_
	);
	LUT2 #(
		.INIT('h4)
	) name144 (
		\G12_pad ,
		\G13_pad ,
		_w177_
	);
	LUT4 #(
		.INIT('h4000)
	) name145 (
		\G3_pad ,
		\G4_pad ,
		\G5_pad ,
		\G6_pad ,
		_w178_
	);
	LUT4 #(
		.INIT('hf05d)
	) name146 (
		\G2_pad ,
		\G3_pad ,
		\G4_pad ,
		\G5_pad ,
		_w179_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name147 (
		\G1_pad ,
		_w141_,
		_w178_,
		_w179_,
		_w180_
	);
	LUT2 #(
		.INIT('h8)
	) name148 (
		_w177_,
		_w180_,
		_w181_
	);
	LUT3 #(
		.INIT('he0)
	) name149 (
		_w123_,
		_w134_,
		_w181_,
		_w182_
	);
	LUT4 #(
		.INIT('h4c00)
	) name150 (
		\G0_pad ,
		\G1_pad ,
		\G3_pad ,
		\G4_pad ,
		_w183_
	);
	LUT3 #(
		.INIT('h10)
	) name151 (
		\G13_pad ,
		\G33_reg/NET0131 ,
		\G3_pad ,
		_w184_
	);
	LUT2 #(
		.INIT('h4)
	) name152 (
		\G12_pad ,
		\G32_reg/NET0131 ,
		_w185_
	);
	LUT3 #(
		.INIT('h10)
	) name153 (
		\G12_pad ,
		\G13_pad ,
		\G32_reg/NET0131 ,
		_w186_
	);
	LUT2 #(
		.INIT('h4)
	) name154 (
		_w58_,
		_w186_,
		_w187_
	);
	LUT2 #(
		.INIT('h8)
	) name155 (
		\G2_pad ,
		\G5_pad ,
		_w188_
	);
	LUT4 #(
		.INIT('h2a00)
	) name156 (
		\G2_pad ,
		\G3_pad ,
		\G4_pad ,
		\G5_pad ,
		_w189_
	);
	LUT4 #(
		.INIT('h2333)
	) name157 (
		_w58_,
		_w184_,
		_w186_,
		_w189_,
		_w190_
	);
	LUT3 #(
		.INIT('h70)
	) name158 (
		_w79_,
		_w183_,
		_w190_,
		_w191_
	);
	LUT2 #(
		.INIT('hb)
	) name159 (
		_w182_,
		_w191_,
		_w192_
	);
	LUT4 #(
		.INIT('hb37f)
	) name160 (
		\G1_pad ,
		\G2_pad ,
		\G4_pad ,
		\G5_pad ,
		_w193_
	);
	LUT2 #(
		.INIT('h2)
	) name161 (
		_w177_,
		_w193_,
		_w194_
	);
	LUT3 #(
		.INIT('he0)
	) name162 (
		_w123_,
		_w134_,
		_w194_,
		_w195_
	);
	LUT4 #(
		.INIT('h4000)
	) name163 (
		\G0_pad ,
		\G1_pad ,
		\G3_pad ,
		\G4_pad ,
		_w196_
	);
	LUT2 #(
		.INIT('h2)
	) name164 (
		\G0_pad ,
		\G29_reg/NET0131 ,
		_w197_
	);
	LUT2 #(
		.INIT('h1)
	) name165 (
		_w196_,
		_w197_,
		_w198_
	);
	LUT4 #(
		.INIT('h4c00)
	) name166 (
		\G2_pad ,
		\G3_pad ,
		\G4_pad ,
		\G5_pad ,
		_w199_
	);
	LUT4 #(
		.INIT('h2333)
	) name167 (
		_w58_,
		_w184_,
		_w186_,
		_w199_,
		_w200_
	);
	LUT3 #(
		.INIT('hd0)
	) name168 (
		_w79_,
		_w198_,
		_w200_,
		_w201_
	);
	LUT2 #(
		.INIT('hb)
	) name169 (
		_w195_,
		_w201_,
		_w202_
	);
	LUT3 #(
		.INIT('h40)
	) name170 (
		\G3_pad ,
		\G4_pad ,
		\G6_pad ,
		_w203_
	);
	LUT3 #(
		.INIT('ha2)
	) name171 (
		\G1_pad ,
		\G4_pad ,
		\G5_pad ,
		_w204_
	);
	LUT4 #(
		.INIT('h0400)
	) name172 (
		\G2_pad ,
		\G3_pad ,
		\G5_pad ,
		\G6_pad ,
		_w205_
	);
	LUT3 #(
		.INIT('h40)
	) name173 (
		\G2_pad ,
		\G3_pad ,
		\G4_pad ,
		_w206_
	);
	LUT4 #(
		.INIT('h0004)
	) name174 (
		_w203_,
		_w204_,
		_w205_,
		_w206_,
		_w207_
	);
	LUT3 #(
		.INIT('h15)
	) name175 (
		\G1_pad ,
		\G2_pad ,
		\G4_pad ,
		_w208_
	);
	LUT3 #(
		.INIT('h02)
	) name176 (
		_w177_,
		_w207_,
		_w208_,
		_w209_
	);
	LUT3 #(
		.INIT('he0)
	) name177 (
		_w123_,
		_w134_,
		_w209_,
		_w210_
	);
	LUT2 #(
		.INIT('h8)
	) name178 (
		\G39_reg/NET0131 ,
		\G4_pad ,
		_w211_
	);
	LUT3 #(
		.INIT('h40)
	) name179 (
		_w58_,
		_w186_,
		_w211_,
		_w212_
	);
	LUT4 #(
		.INIT('h9b5f)
	) name180 (
		\G0_pad ,
		\G1_pad ,
		\G3_pad ,
		\G4_pad ,
		_w213_
	);
	LUT4 #(
		.INIT('h13b3)
	) name181 (
		\G0_pad ,
		\G1_pad ,
		\G2_pad ,
		\G4_pad ,
		_w214_
	);
	LUT4 #(
		.INIT('hf3b3)
	) name182 (
		\G3_pad ,
		\G5_pad ,
		_w213_,
		_w214_,
		_w215_
	);
	LUT3 #(
		.INIT('h31)
	) name183 (
		_w79_,
		_w212_,
		_w215_,
		_w216_
	);
	LUT2 #(
		.INIT('hb)
	) name184 (
		_w210_,
		_w216_,
		_w217_
	);
	LUT3 #(
		.INIT('h23)
	) name185 (
		\G40_reg/NET0131 ,
		\G6_pad ,
		_w79_,
		_w218_
	);
	LUT3 #(
		.INIT('h4c)
	) name186 (
		\G2_pad ,
		\G4_pad ,
		\G5_pad ,
		_w219_
	);
	LUT3 #(
		.INIT('h4c)
	) name187 (
		\G1_pad ,
		\G2_pad ,
		\G4_pad ,
		_w220_
	);
	LUT4 #(
		.INIT('hccc8)
	) name188 (
		_w43_,
		_w177_,
		_w219_,
		_w220_,
		_w221_
	);
	LUT3 #(
		.INIT('he0)
	) name189 (
		_w123_,
		_w134_,
		_w221_,
		_w222_
	);
	LUT4 #(
		.INIT('h4404)
	) name190 (
		\G2_pad ,
		\G3_pad ,
		\G4_pad ,
		\G5_pad ,
		_w223_
	);
	LUT4 #(
		.INIT('h915b)
	) name191 (
		\G2_pad ,
		\G3_pad ,
		\G4_pad ,
		\G5_pad ,
		_w224_
	);
	LUT3 #(
		.INIT('h04)
	) name192 (
		_w58_,
		_w186_,
		_w224_,
		_w225_
	);
	LUT3 #(
		.INIT('h0b)
	) name193 (
		\G40_reg/NET0131 ,
		_w79_,
		_w225_,
		_w226_
	);
	LUT3 #(
		.INIT('h45)
	) name194 (
		_w218_,
		_w222_,
		_w226_,
		_w227_
	);
	LUT4 #(
		.INIT('h0008)
	) name195 (
		\G10_pad ,
		\G11_pad ,
		\G7_pad ,
		\G8_pad ,
		_w228_
	);
	LUT2 #(
		.INIT('h2)
	) name196 (
		\G6_pad ,
		\G9_pad ,
		_w229_
	);
	LUT4 #(
		.INIT('h0001)
	) name197 (
		\G0_pad ,
		\G3_pad ,
		\G4_pad ,
		\G5_pad ,
		_w230_
	);
	LUT3 #(
		.INIT('h80)
	) name198 (
		_w228_,
		_w229_,
		_w230_,
		_w231_
	);
	LUT4 #(
		.INIT('h0100)
	) name199 (
		\G0_pad ,
		\G10_pad ,
		\G4_pad ,
		\G7_pad ,
		_w232_
	);
	LUT3 #(
		.INIT('h80)
	) name200 (
		\G37_reg/NET0131 ,
		\G3_pad ,
		\G5_pad ,
		_w233_
	);
	LUT3 #(
		.INIT('h80)
	) name201 (
		_w62_,
		_w232_,
		_w233_,
		_w234_
	);
	LUT4 #(
		.INIT('h8000)
	) name202 (
		\G0_pad ,
		_w40_,
		_w41_,
		_w44_,
		_w235_
	);
	LUT2 #(
		.INIT('h8)
	) name203 (
		\G1_pad ,
		\G2_pad ,
		_w236_
	);
	LUT4 #(
		.INIT('hfe00)
	) name204 (
		_w231_,
		_w234_,
		_w235_,
		_w236_,
		_w237_
	);
	LUT4 #(
		.INIT('h0002)
	) name205 (
		\G46_reg/NET0131 ,
		_w72_,
		_w75_,
		_w77_,
		_w238_
	);
	LUT2 #(
		.INIT('h8)
	) name206 (
		_w74_,
		_w88_,
		_w239_
	);
	LUT4 #(
		.INIT('hef00)
	) name207 (
		_w67_,
		_w71_,
		_w238_,
		_w239_,
		_w240_
	);
	LUT3 #(
		.INIT('h08)
	) name208 (
		\G38_reg/NET0131 ,
		\G6_pad ,
		\G9_pad ,
		_w241_
	);
	LUT2 #(
		.INIT('h1)
	) name209 (
		_w40_,
		_w241_,
		_w242_
	);
	LUT3 #(
		.INIT('h08)
	) name210 (
		_w237_,
		_w240_,
		_w242_,
		_w243_
	);
	LUT4 #(
		.INIT('haa2a)
	) name211 (
		\G12_pad ,
		_w237_,
		_w240_,
		_w242_,
		_w244_
	);
	LUT4 #(
		.INIT('h0040)
	) name212 (
		\G10_pad ,
		\G6_pad ,
		\G7_pad ,
		\G9_pad ,
		_w245_
	);
	LUT3 #(
		.INIT('ha8)
	) name213 (
		\G8_pad ,
		_w43_,
		_w245_,
		_w246_
	);
	LUT4 #(
		.INIT('hba00)
	) name214 (
		_w92_,
		_w105_,
		_w107_,
		_w246_,
		_w247_
	);
	LUT4 #(
		.INIT('h5100)
	) name215 (
		\G13_pad ,
		\G32_reg/NET0131 ,
		_w58_,
		_w246_,
		_w248_
	);
	LUT3 #(
		.INIT('hd0)
	) name216 (
		_w46_,
		_w55_,
		_w248_,
		_w249_
	);
	LUT2 #(
		.INIT('h8)
	) name217 (
		_w48_,
		_w53_,
		_w250_
	);
	LUT4 #(
		.INIT('hba00)
	) name218 (
		_w92_,
		_w105_,
		_w107_,
		_w250_,
		_w251_
	);
	LUT4 #(
		.INIT('h0001)
	) name219 (
		_w243_,
		_w247_,
		_w249_,
		_w251_,
		_w252_
	);
	LUT4 #(
		.INIT('h1101)
	) name220 (
		\G12_pad ,
		\G13_pad ,
		\G32_reg/NET0131 ,
		_w58_,
		_w253_
	);
	LUT3 #(
		.INIT('h01)
	) name221 (
		\G10_pad ,
		\G11_pad ,
		\G5_pad ,
		_w254_
	);
	LUT4 #(
		.INIT('h0777)
	) name222 (
		_w47_,
		_w49_,
		_w102_,
		_w254_,
		_w255_
	);
	LUT3 #(
		.INIT('h02)
	) name223 (
		\G4_pad ,
		\G5_pad ,
		\G6_pad ,
		_w256_
	);
	LUT3 #(
		.INIT('h80)
	) name224 (
		_w40_,
		_w41_,
		_w256_,
		_w257_
	);
	LUT4 #(
		.INIT('h0031)
	) name225 (
		_w38_,
		_w250_,
		_w255_,
		_w257_,
		_w258_
	);
	LUT4 #(
		.INIT('h00d0)
	) name226 (
		_w46_,
		_w55_,
		_w253_,
		_w258_,
		_w259_
	);
	LUT4 #(
		.INIT('hff02)
	) name227 (
		\G2_pad ,
		_w244_,
		_w252_,
		_w259_,
		_w260_
	);
	LUT3 #(
		.INIT('h08)
	) name228 (
		\G2_pad ,
		\G4_pad ,
		\G5_pad ,
		_w261_
	);
	LUT2 #(
		.INIT('h8)
	) name229 (
		_w185_,
		_w261_,
		_w262_
	);
	LUT2 #(
		.INIT('h4)
	) name230 (
		_w58_,
		_w262_,
		_w263_
	);
	LUT4 #(
		.INIT('h0080)
	) name231 (
		\G0_pad ,
		\G12_pad ,
		\G1_pad ,
		\G4_pad ,
		_w264_
	);
	LUT3 #(
		.INIT('h10)
	) name232 (
		_w75_,
		_w77_,
		_w264_,
		_w265_
	);
	LUT4 #(
		.INIT('h1000)
	) name233 (
		_w67_,
		_w71_,
		_w73_,
		_w265_,
		_w266_
	);
	LUT2 #(
		.INIT('h1)
	) name234 (
		_w263_,
		_w266_,
		_w267_
	);
	LUT3 #(
		.INIT('h45)
	) name235 (
		_w91_,
		_w105_,
		_w106_,
		_w268_
	);
	LUT3 #(
		.INIT('h10)
	) name236 (
		_w123_,
		_w134_,
		_w177_,
		_w269_
	);
	LUT3 #(
		.INIT('hd0)
	) name237 (
		_w46_,
		_w55_,
		_w253_,
		_w270_
	);
	LUT4 #(
		.INIT('he0f0)
	) name238 (
		_w67_,
		_w71_,
		_w74_,
		_w238_,
		_w271_
	);
	LUT2 #(
		.INIT('h8)
	) name239 (
		_w237_,
		_w271_,
		_w272_
	);
	LUT4 #(
		.INIT('hfff4)
	) name240 (
		_w268_,
		_w269_,
		_w270_,
		_w272_,
		_w273_
	);
	LUT2 #(
		.INIT('h4)
	) name241 (
		_w237_,
		_w271_,
		_w274_
	);
	LUT2 #(
		.INIT('h1)
	) name242 (
		\G12_pad ,
		\G13_pad ,
		_w275_
	);
	LUT3 #(
		.INIT('hd0)
	) name243 (
		\G32_reg/NET0131 ,
		_w58_,
		_w275_,
		_w276_
	);
	LUT3 #(
		.INIT('h20)
	) name244 (
		_w46_,
		_w55_,
		_w276_,
		_w277_
	);
	LUT4 #(
		.INIT('hfff8)
	) name245 (
		_w268_,
		_w269_,
		_w274_,
		_w277_,
		_w278_
	);
	LUT4 #(
		.INIT('heebe)
	) name246 (
		\G2_pad ,
		\G3_pad ,
		\G4_pad ,
		\G5_pad ,
		_w279_
	);
	LUT3 #(
		.INIT('h13)
	) name247 (
		\G0_pad ,
		\G1_pad ,
		_w279_,
		_w280_
	);
	LUT3 #(
		.INIT('h8c)
	) name248 (
		\G1_pad ,
		\G2_pad ,
		\G5_pad ,
		_w281_
	);
	LUT4 #(
		.INIT('h010f)
	) name249 (
		\G10_pad ,
		\G30_reg/NET0131 ,
		\G6_pad ,
		\G7_pad ,
		_w282_
	);
	LUT4 #(
		.INIT('h00ef)
	) name250 (
		_w80_,
		_w81_,
		_w281_,
		_w282_,
		_w283_
	);
	LUT2 #(
		.INIT('h4)
	) name251 (
		_w280_,
		_w283_,
		_w284_
	);
	LUT4 #(
		.INIT('h4000)
	) name252 (
		\G11_pad ,
		\G6_pad ,
		\G7_pad ,
		\G9_pad ,
		_w285_
	);
	LUT3 #(
		.INIT('ha8)
	) name253 (
		\G8_pad ,
		_w64_,
		_w285_,
		_w286_
	);
	LUT3 #(
		.INIT('ha8)
	) name254 (
		\G6_pad ,
		_w65_,
		_w99_,
		_w287_
	);
	LUT2 #(
		.INIT('h1)
	) name255 (
		_w286_,
		_w287_,
		_w288_
	);
	LUT3 #(
		.INIT('h02)
	) name256 (
		\G7_pad ,
		\G8_pad ,
		\G9_pad ,
		_w289_
	);
	LUT4 #(
		.INIT('h0080)
	) name257 (
		\G10_pad ,
		\G6_pad ,
		\G8_pad ,
		\G9_pad ,
		_w290_
	);
	LUT4 #(
		.INIT('h93cf)
	) name258 (
		\G10_pad ,
		\G6_pad ,
		\G7_pad ,
		\G9_pad ,
		_w291_
	);
	LUT4 #(
		.INIT('h5755)
	) name259 (
		\G11_pad ,
		_w289_,
		_w290_,
		_w291_,
		_w292_
	);
	LUT4 #(
		.INIT('hf377)
	) name260 (
		\G2_pad ,
		\G4_pad ,
		\G5_pad ,
		\G6_pad ,
		_w293_
	);
	LUT2 #(
		.INIT('h2)
	) name261 (
		_w87_,
		_w293_,
		_w294_
	);
	LUT3 #(
		.INIT('ha8)
	) name262 (
		\G1_pad ,
		_w124_,
		_w126_,
		_w295_
	);
	LUT3 #(
		.INIT('h40)
	) name263 (
		\G1_pad ,
		\G2_pad ,
		\G3_pad ,
		_w296_
	);
	LUT2 #(
		.INIT('h4)
	) name264 (
		_w120_,
		_w296_,
		_w297_
	);
	LUT3 #(
		.INIT('h01)
	) name265 (
		_w294_,
		_w295_,
		_w297_,
		_w298_
	);
	LUT4 #(
		.INIT('h0200)
	) name266 (
		\G10_pad ,
		\G7_pad ,
		\G8_pad ,
		\G9_pad ,
		_w299_
	);
	LUT2 #(
		.INIT('h8)
	) name267 (
		_w49_,
		_w299_,
		_w300_
	);
	LUT3 #(
		.INIT('h20)
	) name268 (
		\G10_pad ,
		\G4_pad ,
		\G7_pad ,
		_w301_
	);
	LUT4 #(
		.INIT('h0bbb)
	) name269 (
		\G9_pad ,
		_w39_,
		_w41_,
		_w301_,
		_w302_
	);
	LUT2 #(
		.INIT('h1)
	) name270 (
		\G5_pad ,
		\G6_pad ,
		_w303_
	);
	LUT3 #(
		.INIT('h45)
	) name271 (
		_w300_,
		_w302_,
		_w303_,
		_w304_
	);
	LUT4 #(
		.INIT('hb1a0)
	) name272 (
		\G6_pad ,
		\G9_pad ,
		_w48_,
		_w101_,
		_w305_
	);
	LUT4 #(
		.INIT('h5444)
	) name273 (
		\G5_pad ,
		_w39_,
		_w40_,
		_w41_,
		_w306_
	);
	LUT2 #(
		.INIT('h4)
	) name274 (
		_w53_,
		_w188_,
		_w307_
	);
	LUT3 #(
		.INIT('h0b)
	) name275 (
		_w120_,
		_w125_,
		_w261_,
		_w308_
	);
	LUT2 #(
		.INIT('hb)
	) name276 (
		_w307_,
		_w308_,
		_w309_
	);
	LUT3 #(
		.INIT('h47)
	) name277 (
		\G3_pad ,
		\G4_pad ,
		\G5_pad ,
		_w310_
	);
	LUT3 #(
		.INIT('h31)
	) name278 (
		_w121_,
		_w223_,
		_w310_,
		_w311_
	);
	LUT3 #(
		.INIT('h6a)
	) name279 (
		\G2_pad ,
		\G3_pad ,
		\G5_pad ,
		_w312_
	);
	LUT4 #(
		.INIT('h2eae)
	) name280 (
		\G10_pad ,
		\G11_pad ,
		\G7_pad ,
		\G9_pad ,
		_w313_
	);
	LUT3 #(
		.INIT('hae)
	) name281 (
		\G10_pad ,
		\G11_pad ,
		\G9_pad ,
		_w314_
	);
	LUT2 #(
		.INIT('h6)
	) name282 (
		\G6_pad ,
		\G9_pad ,
		_w315_
	);
	LUT4 #(
		.INIT('h20a0)
	) name283 (
		\G10_pad ,
		\G6_pad ,
		\G7_pad ,
		\G9_pad ,
		_w316_
	);
	LUT2 #(
		.INIT('h8)
	) name284 (
		\G34_reg/NET0131 ,
		_w157_,
		_w317_
	);
	LUT3 #(
		.INIT('h07)
	) name285 (
		_w79_,
		_w316_,
		_w317_,
		_w318_
	);
	LUT2 #(
		.INIT('h8)
	) name286 (
		_w153_,
		_w318_,
		_w319_
	);
	LUT2 #(
		.INIT('h4)
	) name287 (
		\G4_pad ,
		_w48_,
		_w320_
	);
	LUT4 #(
		.INIT('hba00)
	) name288 (
		_w92_,
		_w105_,
		_w107_,
		_w320_,
		_w321_
	);
	LUT4 #(
		.INIT('h5100)
	) name289 (
		\G13_pad ,
		\G32_reg/NET0131 ,
		_w58_,
		_w320_,
		_w322_
	);
	LUT3 #(
		.INIT('hd0)
	) name290 (
		_w46_,
		_w55_,
		_w322_,
		_w323_
	);
	LUT3 #(
		.INIT('h54)
	) name291 (
		\G10_pad ,
		\G7_pad ,
		\G9_pad ,
		_w324_
	);
	LUT2 #(
		.INIT('h8)
	) name292 (
		_w127_,
		_w324_,
		_w325_
	);
	LUT4 #(
		.INIT('hba00)
	) name293 (
		_w92_,
		_w105_,
		_w107_,
		_w325_,
		_w326_
	);
	LUT2 #(
		.INIT('h4)
	) name294 (
		\G12_pad ,
		\G6_pad ,
		_w327_
	);
	LUT4 #(
		.INIT('hfe00)
	) name295 (
		_w321_,
		_w323_,
		_w326_,
		_w327_,
		_w328_
	);
	LUT2 #(
		.INIT('h1)
	) name296 (
		\G3_pad ,
		\G44_reg/NET0131 ,
		_w329_
	);
	LUT4 #(
		.INIT('h007f)
	) name297 (
		_w35_,
		_w53_,
		_w324_,
		_w329_,
		_w330_
	);
	LUT2 #(
		.INIT('h1)
	) name298 (
		\G12_pad ,
		_w330_,
		_w331_
	);
	LUT4 #(
		.INIT('hd000)
	) name299 (
		_w46_,
		_w55_,
		_w59_,
		_w331_,
		_w332_
	);
	LUT2 #(
		.INIT('h8)
	) name300 (
		\G37_reg/NET0131 ,
		\G38_reg/NET0131 ,
		_w333_
	);
	LUT3 #(
		.INIT('h80)
	) name301 (
		_w237_,
		_w240_,
		_w333_,
		_w334_
	);
	LUT2 #(
		.INIT('h1)
	) name302 (
		_w332_,
		_w334_,
		_w335_
	);
	LUT2 #(
		.INIT('hb)
	) name303 (
		_w328_,
		_w335_,
		_w336_
	);
	LUT4 #(
		.INIT('hffe0)
	) name304 (
		_w123_,
		_w134_,
		_w177_,
		_w187_,
		_w337_
	);
	assign \G530_pad  = _w86_ ;
	assign \G532_pad  = _w149_ ;
	assign \G542_pad  = _w160_ ;
	assign \G546_pad  = _w23_ ;
	assign \G547_pad  = _w172_ ;
	assign \G548_pad  = _w176_ ;
	assign \G549_pad  = _w192_ ;
	assign \G550_pad  = _w202_ ;
	assign \G551_pad  = _w217_ ;
	assign \G552_pad  = _w227_ ;
	assign \_al_n0  = 1'b0;
	assign \_al_n1  = 1'b1;
	assign \g1594/_3_  = _w260_ ;
	assign \g1613/_0_  = _w267_ ;
	assign \g1618/_0_  = _w273_ ;
	assign \g1620/_2_  = _w278_ ;
	assign \g1692/_0_  = _w284_ ;
	assign \g1727/_0_  = _w288_ ;
	assign \g1740/_0_  = _w292_ ;
	assign \g1742/_0_  = _w298_ ;
	assign \g1760/_0_  = _w304_ ;
	assign \g1769/_3_  = _w305_ ;
	assign \g1771/_0_  = _w306_ ;
	assign \g1780/_0_  = _w309_ ;
	assign \g1799/_0_  = _w311_ ;
	assign \g1867/_0_  = _w312_ ;
	assign \g1873/_0_  = _w313_ ;
	assign \g1900/_0_  = _w232_ ;
	assign \g1930/_0_  = _w314_ ;
	assign \g1936/_0_  = _w315_ ;
	assign \g2340/_2_  = _w319_ ;
	assign \g2396/_1_  = _w336_ ;
	assign \g2408/_0_  = _w337_ ;
endmodule;