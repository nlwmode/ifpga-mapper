module top( \G0_pad  , \G1_pad  , \G2_pad  , \G3_pad  , \G5_reg/NET0131  , \G6_reg/NET0131  , \G7_reg/NET0131  , \G17_pad  , \_al_n0  , \_al_n1  , \g17/_1_  , \g70/_1_  , \g74/_0_  );
  input \G0_pad  ;
  input \G1_pad  ;
  input \G2_pad  ;
  input \G3_pad  ;
  input \G5_reg/NET0131  ;
  input \G6_reg/NET0131  ;
  input \G7_reg/NET0131  ;
  output \G17_pad  ;
  output \_al_n0  ;
  output \_al_n1  ;
  output \g17/_1_  ;
  output \g70/_1_  ;
  output \g74/_0_  ;
  wire n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 ;
  assign n8 = ~\G0_pad  & \G6_reg/NET0131  ;
  assign n9 = ~\G5_reg/NET0131  & n8 ;
  assign n10 = ~\G1_pad  & ~\G7_reg/NET0131  ;
  assign n11 = \G3_pad  & ~\G5_reg/NET0131  ;
  assign n12 = n10 & n11 ;
  assign n13 = ~n9 & ~n12 ;
  assign n14 = \G0_pad  & n13 ;
  assign n15 = ~\G2_pad  & ~n10 ;
  assign \G17_pad  = n13 ;
  assign \_al_n0  = 1'b0 ;
  assign \_al_n1  = ~1'b0 ;
  assign \g17/_1_  = ~n13 ;
  assign \g70/_1_  = n14 ;
  assign \g74/_0_  = n15 ;
endmodule
