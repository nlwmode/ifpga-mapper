module top (\address_reg[0]/NET0131 , \address_reg[1]/NET0131 , \address_reg[2]/NET0131 , \address_reg[3]/NET0131 , \address_reg[4]/NET0131 , \count_reg[0]/NET0131 , \count_reg[0]1198/NET0131 , \count_reg[1]/NET0131 , \count_reg[1]1200/NET0131 , \count_reg[2]/NET0131 , \count_reg[3]/NET0131 , \count_reg[4]/NET0131 , \count_reg[5]/NET0131 , \counter_reg[0]/NET0131 , \counter_reg[1]/NET0131 , \counter_reg[2]/NET0131 , \data_in_reg[0]/NET0131 , \data_in_reg[1]/NET0131 , \data_out_reg[0]/NET0131 , \data_out_reg[1]/NET0131 , \gamma_reg[0]/NET0131 , \gamma_reg[1]/NET0131 , \gamma_reg[2]/NET0131 , \gamma_reg[3]/NET0131 , \gamma_reg[4]/NET0131 , \ind_reg[0]/NET0131 , \ind_reg[1]/NET0131 , \k[0]_pad , \k[1]_pad , \k[2]_pad , \k[3]_pad , \max_reg[0]/NET0131 , \max_reg[1]/NET0131 , \max_reg[2]/NET0131 , \max_reg[3]/NET0131 , \max_reg[4]/NET0131 , \memory_reg[0][0]/NET0131 , \memory_reg[0][1]/NET0131 , \memory_reg[10][0]/NET0131 , \memory_reg[10][1]/NET0131 , \memory_reg[11][0]/NET0131 , \memory_reg[11][1]/NET0131 , \memory_reg[12][0]/NET0131 , \memory_reg[12][1]/NET0131 , \memory_reg[13][0]/NET0131 , \memory_reg[13][1]/NET0131 , \memory_reg[14][0]/NET0131 , \memory_reg[14][1]/NET0131 , \memory_reg[15][0]/NET0131 , \memory_reg[15][1]/NET0131 , \memory_reg[16][0]/NET0131 , \memory_reg[16][1]/NET0131 , \memory_reg[17][0]/NET0131 , \memory_reg[17][1]/NET0131 , \memory_reg[18][0]/NET0131 , \memory_reg[18][1]/NET0131 , \memory_reg[19][0]/NET0131 , \memory_reg[19][1]/NET0131 , \memory_reg[1][0]/NET0131 , \memory_reg[1][1]/NET0131 , \memory_reg[20][0]/NET0131 , \memory_reg[20][1]/NET0131 , \memory_reg[21][0]/NET0131 , \memory_reg[21][1]/NET0131 , \memory_reg[22][0]/NET0131 , \memory_reg[22][1]/NET0131 , \memory_reg[23][0]/NET0131 , \memory_reg[23][1]/NET0131 , \memory_reg[24][0]/NET0131 , \memory_reg[24][1]/NET0131 , \memory_reg[25][0]/NET0131 , \memory_reg[25][1]/NET0131 , \memory_reg[26][0]/NET0131 , \memory_reg[26][1]/NET0131 , \memory_reg[27][0]/NET0131 , \memory_reg[27][1]/NET0131 , \memory_reg[28][0]/NET0131 , \memory_reg[28][1]/NET0131 , \memory_reg[29][0]/NET0131 , \memory_reg[29][1]/NET0131 , \memory_reg[2][0]/NET0131 , \memory_reg[2][1]/NET0131 , \memory_reg[30][0]/NET0131 , \memory_reg[30][1]/NET0131 , \memory_reg[31][0]/NET0131 , \memory_reg[31][1]/NET0131 , \memory_reg[3][0]/NET0131 , \memory_reg[3][1]/NET0131 , \memory_reg[4][0]/NET0131 , \memory_reg[4][1]/NET0131 , \memory_reg[5][0]/NET0131 , \memory_reg[5][1]/NET0131 , \memory_reg[6][0]/NET0131 , \memory_reg[6][1]/NET0131 , \memory_reg[7][0]/NET0131 , \memory_reg[7][1]/NET0131 , \memory_reg[8][0]/NET0131 , \memory_reg[8][1]/NET0131 , \memory_reg[9][0]/NET0131 , \memory_reg[9][1]/NET0131 , \nl[0]_pad , \nl[2]_pad , \nl[3]_pad , \nl_reg[1]/NET0131 , nloss_pad, \play_reg/NET0131 , \s_reg/NET0131 , \scan_reg[0]/NET0131 , \scan_reg[1]/NET0131 , \scan_reg[2]/NET0131 , \scan_reg[3]/NET0131 , \scan_reg[4]/NET0131 , \sound_reg[0]/NET0131 , \sound_reg[1]/NET0131 , \sound_reg[2]/NET0131 , speaker_pad, start_pad, \timebase_reg[0]/NET0131 , \timebase_reg[1]/NET0131 , \timebase_reg[2]/NET0131 , \timebase_reg[3]/NET0131 , \timebase_reg[4]/NET0131 , \timebase_reg[5]/NET0131 , \wr_reg/NET0131 , \_al_n0 , \_al_n1 , \count_reg[0]/P0001 , \g10376/_0_ , \g11078/_0_ , \g11102/_0_ , \g11126/_0_ , \g11156/_0_ , \g11299/_0_ , \g11308/_0_ , \g11318/_0_ , \g11346/_0_ , \g11378/_0_ , \g11516/_0_ , \g63/_0_ , \g8501/_0_ , \g8516/_0_ , \g8517/_0_ , \g8519/_0_ , \g8520/_0_ , \g8522/_0_ , \g8526/_0_ , \g8529/_2_ , \g8545/_0_ , \g8546/_0_ , \g8547/_0_ , \g8555/_0_ , \g8556/_0_ , \g8557/_0_ , \g8558/_0_ , \g8559/_0_ , \g8560/_0_ , \g8562/_0_ , \g8563/_0_ , \g8581/_0_ , \g8586/_0_ , \g8591/_0_ , \g8594/_0_ , \g8606/_0_ , \g8608/_0_ , \g8647/_0_ , \g8659/_0_ , \g8695/_0_ , \g8784/_0_ , \g8797/_0_ , \g8854/_2_ , \g8869/_0_ , \g8871/_0_ , \g8889/_0_ , \g8891/_0_ , \g8892/_0_ , \g8894/_0_ , \g8970/_0_ , \g8975/_0_ , \g8992/_0_ , \g9180/_0_ , \g9183/_0_ , \g9511/u3_syn_4 , \g9513/u3_syn_4 , \g9515/u3_syn_4 , \g9517/u3_syn_4 , \g9519/u3_syn_4 , \g9521/u3_syn_4 , \g9523/u3_syn_4 , \g9525/u3_syn_4 , \g9527/u3_syn_4 , \g9529/u3_syn_4 , \g9531/u3_syn_4 , \g9533/u3_syn_4 , \g9535/u3_syn_4 , \g9537/u3_syn_4 , \g9539/u3_syn_4 , \g9541/u3_syn_4 , \g9543/u3_syn_4 , \g9545/u3_syn_4 , \g9547/u3_syn_4 , \g9549/u3_syn_4 , \g9551/u3_syn_4 , \g9553/u3_syn_4 , \g9555/u3_syn_4 , \g9557/u3_syn_4 , \g9559/u3_syn_4 , \g9560/u3_syn_4 , \g9562/u3_syn_4 , \g9564/u3_syn_4 , \g9566/u3_syn_4 , \g9568/u3_syn_4 , \g9570/u3_syn_4 , \g9572/u3_syn_4 );
	input \address_reg[0]/NET0131  ;
	input \address_reg[1]/NET0131  ;
	input \address_reg[2]/NET0131  ;
	input \address_reg[3]/NET0131  ;
	input \address_reg[4]/NET0131  ;
	input \count_reg[0]/NET0131  ;
	input \count_reg[0]1198/NET0131  ;
	input \count_reg[1]/NET0131  ;
	input \count_reg[1]1200/NET0131  ;
	input \count_reg[2]/NET0131  ;
	input \count_reg[3]/NET0131  ;
	input \count_reg[4]/NET0131  ;
	input \count_reg[5]/NET0131  ;
	input \counter_reg[0]/NET0131  ;
	input \counter_reg[1]/NET0131  ;
	input \counter_reg[2]/NET0131  ;
	input \data_in_reg[0]/NET0131  ;
	input \data_in_reg[1]/NET0131  ;
	input \data_out_reg[0]/NET0131  ;
	input \data_out_reg[1]/NET0131  ;
	input \gamma_reg[0]/NET0131  ;
	input \gamma_reg[1]/NET0131  ;
	input \gamma_reg[2]/NET0131  ;
	input \gamma_reg[3]/NET0131  ;
	input \gamma_reg[4]/NET0131  ;
	input \ind_reg[0]/NET0131  ;
	input \ind_reg[1]/NET0131  ;
	input \k[0]_pad  ;
	input \k[1]_pad  ;
	input \k[2]_pad  ;
	input \k[3]_pad  ;
	input \max_reg[0]/NET0131  ;
	input \max_reg[1]/NET0131  ;
	input \max_reg[2]/NET0131  ;
	input \max_reg[3]/NET0131  ;
	input \max_reg[4]/NET0131  ;
	input \memory_reg[0][0]/NET0131  ;
	input \memory_reg[0][1]/NET0131  ;
	input \memory_reg[10][0]/NET0131  ;
	input \memory_reg[10][1]/NET0131  ;
	input \memory_reg[11][0]/NET0131  ;
	input \memory_reg[11][1]/NET0131  ;
	input \memory_reg[12][0]/NET0131  ;
	input \memory_reg[12][1]/NET0131  ;
	input \memory_reg[13][0]/NET0131  ;
	input \memory_reg[13][1]/NET0131  ;
	input \memory_reg[14][0]/NET0131  ;
	input \memory_reg[14][1]/NET0131  ;
	input \memory_reg[15][0]/NET0131  ;
	input \memory_reg[15][1]/NET0131  ;
	input \memory_reg[16][0]/NET0131  ;
	input \memory_reg[16][1]/NET0131  ;
	input \memory_reg[17][0]/NET0131  ;
	input \memory_reg[17][1]/NET0131  ;
	input \memory_reg[18][0]/NET0131  ;
	input \memory_reg[18][1]/NET0131  ;
	input \memory_reg[19][0]/NET0131  ;
	input \memory_reg[19][1]/NET0131  ;
	input \memory_reg[1][0]/NET0131  ;
	input \memory_reg[1][1]/NET0131  ;
	input \memory_reg[20][0]/NET0131  ;
	input \memory_reg[20][1]/NET0131  ;
	input \memory_reg[21][0]/NET0131  ;
	input \memory_reg[21][1]/NET0131  ;
	input \memory_reg[22][0]/NET0131  ;
	input \memory_reg[22][1]/NET0131  ;
	input \memory_reg[23][0]/NET0131  ;
	input \memory_reg[23][1]/NET0131  ;
	input \memory_reg[24][0]/NET0131  ;
	input \memory_reg[24][1]/NET0131  ;
	input \memory_reg[25][0]/NET0131  ;
	input \memory_reg[25][1]/NET0131  ;
	input \memory_reg[26][0]/NET0131  ;
	input \memory_reg[26][1]/NET0131  ;
	input \memory_reg[27][0]/NET0131  ;
	input \memory_reg[27][1]/NET0131  ;
	input \memory_reg[28][0]/NET0131  ;
	input \memory_reg[28][1]/NET0131  ;
	input \memory_reg[29][0]/NET0131  ;
	input \memory_reg[29][1]/NET0131  ;
	input \memory_reg[2][0]/NET0131  ;
	input \memory_reg[2][1]/NET0131  ;
	input \memory_reg[30][0]/NET0131  ;
	input \memory_reg[30][1]/NET0131  ;
	input \memory_reg[31][0]/NET0131  ;
	input \memory_reg[31][1]/NET0131  ;
	input \memory_reg[3][0]/NET0131  ;
	input \memory_reg[3][1]/NET0131  ;
	input \memory_reg[4][0]/NET0131  ;
	input \memory_reg[4][1]/NET0131  ;
	input \memory_reg[5][0]/NET0131  ;
	input \memory_reg[5][1]/NET0131  ;
	input \memory_reg[6][0]/NET0131  ;
	input \memory_reg[6][1]/NET0131  ;
	input \memory_reg[7][0]/NET0131  ;
	input \memory_reg[7][1]/NET0131  ;
	input \memory_reg[8][0]/NET0131  ;
	input \memory_reg[8][1]/NET0131  ;
	input \memory_reg[9][0]/NET0131  ;
	input \memory_reg[9][1]/NET0131  ;
	input \nl[0]_pad  ;
	input \nl[2]_pad  ;
	input \nl[3]_pad  ;
	input \nl_reg[1]/NET0131  ;
	input nloss_pad ;
	input \play_reg/NET0131  ;
	input \s_reg/NET0131  ;
	input \scan_reg[0]/NET0131  ;
	input \scan_reg[1]/NET0131  ;
	input \scan_reg[2]/NET0131  ;
	input \scan_reg[3]/NET0131  ;
	input \scan_reg[4]/NET0131  ;
	input \sound_reg[0]/NET0131  ;
	input \sound_reg[1]/NET0131  ;
	input \sound_reg[2]/NET0131  ;
	input speaker_pad ;
	input start_pad ;
	input \timebase_reg[0]/NET0131  ;
	input \timebase_reg[1]/NET0131  ;
	input \timebase_reg[2]/NET0131  ;
	input \timebase_reg[3]/NET0131  ;
	input \timebase_reg[4]/NET0131  ;
	input \timebase_reg[5]/NET0131  ;
	input \wr_reg/NET0131  ;
	output \_al_n0  ;
	output \_al_n1  ;
	output \count_reg[0]/P0001  ;
	output \g10376/_0_  ;
	output \g11078/_0_  ;
	output \g11102/_0_  ;
	output \g11126/_0_  ;
	output \g11156/_0_  ;
	output \g11299/_0_  ;
	output \g11308/_0_  ;
	output \g11318/_0_  ;
	output \g11346/_0_  ;
	output \g11378/_0_  ;
	output \g11516/_0_  ;
	output \g63/_0_  ;
	output \g8501/_0_  ;
	output \g8516/_0_  ;
	output \g8517/_0_  ;
	output \g8519/_0_  ;
	output \g8520/_0_  ;
	output \g8522/_0_  ;
	output \g8526/_0_  ;
	output \g8529/_2_  ;
	output \g8545/_0_  ;
	output \g8546/_0_  ;
	output \g8547/_0_  ;
	output \g8555/_0_  ;
	output \g8556/_0_  ;
	output \g8557/_0_  ;
	output \g8558/_0_  ;
	output \g8559/_0_  ;
	output \g8560/_0_  ;
	output \g8562/_0_  ;
	output \g8563/_0_  ;
	output \g8581/_0_  ;
	output \g8586/_0_  ;
	output \g8591/_0_  ;
	output \g8594/_0_  ;
	output \g8606/_0_  ;
	output \g8608/_0_  ;
	output \g8647/_0_  ;
	output \g8659/_0_  ;
	output \g8695/_0_  ;
	output \g8784/_0_  ;
	output \g8797/_0_  ;
	output \g8854/_2_  ;
	output \g8869/_0_  ;
	output \g8871/_0_  ;
	output \g8889/_0_  ;
	output \g8891/_0_  ;
	output \g8892/_0_  ;
	output \g8894/_0_  ;
	output \g8970/_0_  ;
	output \g8975/_0_  ;
	output \g8992/_0_  ;
	output \g9180/_0_  ;
	output \g9183/_0_  ;
	output \g9511/u3_syn_4  ;
	output \g9513/u3_syn_4  ;
	output \g9515/u3_syn_4  ;
	output \g9517/u3_syn_4  ;
	output \g9519/u3_syn_4  ;
	output \g9521/u3_syn_4  ;
	output \g9523/u3_syn_4  ;
	output \g9525/u3_syn_4  ;
	output \g9527/u3_syn_4  ;
	output \g9529/u3_syn_4  ;
	output \g9531/u3_syn_4  ;
	output \g9533/u3_syn_4  ;
	output \g9535/u3_syn_4  ;
	output \g9537/u3_syn_4  ;
	output \g9539/u3_syn_4  ;
	output \g9541/u3_syn_4  ;
	output \g9543/u3_syn_4  ;
	output \g9545/u3_syn_4  ;
	output \g9547/u3_syn_4  ;
	output \g9549/u3_syn_4  ;
	output \g9551/u3_syn_4  ;
	output \g9553/u3_syn_4  ;
	output \g9555/u3_syn_4  ;
	output \g9557/u3_syn_4  ;
	output \g9559/u3_syn_4  ;
	output \g9560/u3_syn_4  ;
	output \g9562/u3_syn_4  ;
	output \g9564/u3_syn_4  ;
	output \g9566/u3_syn_4  ;
	output \g9568/u3_syn_4  ;
	output \g9570/u3_syn_4  ;
	output \g9572/u3_syn_4  ;
	wire _w1198_ ;
	wire _w1197_ ;
	wire _w1196_ ;
	wire _w1195_ ;
	wire _w1194_ ;
	wire _w1193_ ;
	wire _w1192_ ;
	wire _w1191_ ;
	wire _w1190_ ;
	wire _w1189_ ;
	wire _w1188_ ;
	wire _w1187_ ;
	wire _w1186_ ;
	wire _w1185_ ;
	wire _w1184_ ;
	wire _w1183_ ;
	wire _w1182_ ;
	wire _w1181_ ;
	wire _w1180_ ;
	wire _w1179_ ;
	wire _w1178_ ;
	wire _w1177_ ;
	wire _w1176_ ;
	wire _w1175_ ;
	wire _w1174_ ;
	wire _w1173_ ;
	wire _w1172_ ;
	wire _w1171_ ;
	wire _w1170_ ;
	wire _w1169_ ;
	wire _w1168_ ;
	wire _w1167_ ;
	wire _w1166_ ;
	wire _w1165_ ;
	wire _w1164_ ;
	wire _w1163_ ;
	wire _w1162_ ;
	wire _w1161_ ;
	wire _w1160_ ;
	wire _w1159_ ;
	wire _w1158_ ;
	wire _w1157_ ;
	wire _w1156_ ;
	wire _w1155_ ;
	wire _w1154_ ;
	wire _w1153_ ;
	wire _w1152_ ;
	wire _w1151_ ;
	wire _w1150_ ;
	wire _w1149_ ;
	wire _w1148_ ;
	wire _w1147_ ;
	wire _w1146_ ;
	wire _w1145_ ;
	wire _w1144_ ;
	wire _w1143_ ;
	wire _w1142_ ;
	wire _w1141_ ;
	wire _w1140_ ;
	wire _w1139_ ;
	wire _w1138_ ;
	wire _w1137_ ;
	wire _w1136_ ;
	wire _w1135_ ;
	wire _w1134_ ;
	wire _w1133_ ;
	wire _w1132_ ;
	wire _w1131_ ;
	wire _w1130_ ;
	wire _w1129_ ;
	wire _w1128_ ;
	wire _w1127_ ;
	wire _w1126_ ;
	wire _w1125_ ;
	wire _w1124_ ;
	wire _w1123_ ;
	wire _w1122_ ;
	wire _w1121_ ;
	wire _w1120_ ;
	wire _w1119_ ;
	wire _w1118_ ;
	wire _w1117_ ;
	wire _w1116_ ;
	wire _w1115_ ;
	wire _w1114_ ;
	wire _w1113_ ;
	wire _w1112_ ;
	wire _w1111_ ;
	wire _w1110_ ;
	wire _w1109_ ;
	wire _w1108_ ;
	wire _w1107_ ;
	wire _w1106_ ;
	wire _w1105_ ;
	wire _w1104_ ;
	wire _w1103_ ;
	wire _w1102_ ;
	wire _w1101_ ;
	wire _w1100_ ;
	wire _w1099_ ;
	wire _w1098_ ;
	wire _w1097_ ;
	wire _w1096_ ;
	wire _w1095_ ;
	wire _w1094_ ;
	wire _w1093_ ;
	wire _w1092_ ;
	wire _w1091_ ;
	wire _w1090_ ;
	wire _w1089_ ;
	wire _w1088_ ;
	wire _w1087_ ;
	wire _w1086_ ;
	wire _w1085_ ;
	wire _w1084_ ;
	wire _w1083_ ;
	wire _w1082_ ;
	wire _w1081_ ;
	wire _w1080_ ;
	wire _w1079_ ;
	wire _w1078_ ;
	wire _w1077_ ;
	wire _w1076_ ;
	wire _w1075_ ;
	wire _w1074_ ;
	wire _w1073_ ;
	wire _w1072_ ;
	wire _w1071_ ;
	wire _w1070_ ;
	wire _w1069_ ;
	wire _w1068_ ;
	wire _w1067_ ;
	wire _w1066_ ;
	wire _w1065_ ;
	wire _w1064_ ;
	wire _w1063_ ;
	wire _w1062_ ;
	wire _w1061_ ;
	wire _w1060_ ;
	wire _w1059_ ;
	wire _w1058_ ;
	wire _w1057_ ;
	wire _w1056_ ;
	wire _w1055_ ;
	wire _w1054_ ;
	wire _w1053_ ;
	wire _w1052_ ;
	wire _w1051_ ;
	wire _w1050_ ;
	wire _w1049_ ;
	wire _w1048_ ;
	wire _w1047_ ;
	wire _w1046_ ;
	wire _w1045_ ;
	wire _w1044_ ;
	wire _w1043_ ;
	wire _w1042_ ;
	wire _w1041_ ;
	wire _w1040_ ;
	wire _w1039_ ;
	wire _w1038_ ;
	wire _w1037_ ;
	wire _w1036_ ;
	wire _w1035_ ;
	wire _w1034_ ;
	wire _w1033_ ;
	wire _w1032_ ;
	wire _w1031_ ;
	wire _w1030_ ;
	wire _w1029_ ;
	wire _w1028_ ;
	wire _w1027_ ;
	wire _w1026_ ;
	wire _w1025_ ;
	wire _w1024_ ;
	wire _w1023_ ;
	wire _w1022_ ;
	wire _w1021_ ;
	wire _w1020_ ;
	wire _w1019_ ;
	wire _w1018_ ;
	wire _w1017_ ;
	wire _w1016_ ;
	wire _w1015_ ;
	wire _w1014_ ;
	wire _w1013_ ;
	wire _w1012_ ;
	wire _w1011_ ;
	wire _w1010_ ;
	wire _w1009_ ;
	wire _w1008_ ;
	wire _w1007_ ;
	wire _w1006_ ;
	wire _w1005_ ;
	wire _w1004_ ;
	wire _w1003_ ;
	wire _w1002_ ;
	wire _w1001_ ;
	wire _w1000_ ;
	wire _w999_ ;
	wire _w998_ ;
	wire _w997_ ;
	wire _w996_ ;
	wire _w995_ ;
	wire _w994_ ;
	wire _w993_ ;
	wire _w992_ ;
	wire _w991_ ;
	wire _w990_ ;
	wire _w989_ ;
	wire _w988_ ;
	wire _w987_ ;
	wire _w986_ ;
	wire _w985_ ;
	wire _w984_ ;
	wire _w983_ ;
	wire _w982_ ;
	wire _w981_ ;
	wire _w980_ ;
	wire _w979_ ;
	wire _w978_ ;
	wire _w977_ ;
	wire _w976_ ;
	wire _w975_ ;
	wire _w974_ ;
	wire _w973_ ;
	wire _w972_ ;
	wire _w971_ ;
	wire _w970_ ;
	wire _w969_ ;
	wire _w968_ ;
	wire _w967_ ;
	wire _w966_ ;
	wire _w965_ ;
	wire _w964_ ;
	wire _w963_ ;
	wire _w962_ ;
	wire _w961_ ;
	wire _w960_ ;
	wire _w959_ ;
	wire _w958_ ;
	wire _w957_ ;
	wire _w956_ ;
	wire _w955_ ;
	wire _w954_ ;
	wire _w953_ ;
	wire _w952_ ;
	wire _w951_ ;
	wire _w950_ ;
	wire _w949_ ;
	wire _w948_ ;
	wire _w947_ ;
	wire _w946_ ;
	wire _w945_ ;
	wire _w944_ ;
	wire _w943_ ;
	wire _w942_ ;
	wire _w941_ ;
	wire _w940_ ;
	wire _w939_ ;
	wire _w938_ ;
	wire _w937_ ;
	wire _w936_ ;
	wire _w935_ ;
	wire _w934_ ;
	wire _w933_ ;
	wire _w932_ ;
	wire _w931_ ;
	wire _w930_ ;
	wire _w929_ ;
	wire _w928_ ;
	wire _w927_ ;
	wire _w926_ ;
	wire _w925_ ;
	wire _w924_ ;
	wire _w923_ ;
	wire _w922_ ;
	wire _w921_ ;
	wire _w920_ ;
	wire _w919_ ;
	wire _w918_ ;
	wire _w917_ ;
	wire _w916_ ;
	wire _w915_ ;
	wire _w914_ ;
	wire _w913_ ;
	wire _w912_ ;
	wire _w911_ ;
	wire _w910_ ;
	wire _w909_ ;
	wire _w908_ ;
	wire _w907_ ;
	wire _w906_ ;
	wire _w905_ ;
	wire _w904_ ;
	wire _w903_ ;
	wire _w902_ ;
	wire _w901_ ;
	wire _w900_ ;
	wire _w899_ ;
	wire _w898_ ;
	wire _w897_ ;
	wire _w896_ ;
	wire _w895_ ;
	wire _w894_ ;
	wire _w893_ ;
	wire _w892_ ;
	wire _w891_ ;
	wire _w890_ ;
	wire _w889_ ;
	wire _w888_ ;
	wire _w887_ ;
	wire _w886_ ;
	wire _w885_ ;
	wire _w884_ ;
	wire _w883_ ;
	wire _w882_ ;
	wire _w881_ ;
	wire _w880_ ;
	wire _w879_ ;
	wire _w878_ ;
	wire _w877_ ;
	wire _w876_ ;
	wire _w875_ ;
	wire _w874_ ;
	wire _w873_ ;
	wire _w872_ ;
	wire _w871_ ;
	wire _w870_ ;
	wire _w869_ ;
	wire _w868_ ;
	wire _w867_ ;
	wire _w866_ ;
	wire _w865_ ;
	wire _w864_ ;
	wire _w863_ ;
	wire _w862_ ;
	wire _w861_ ;
	wire _w860_ ;
	wire _w859_ ;
	wire _w858_ ;
	wire _w857_ ;
	wire _w856_ ;
	wire _w855_ ;
	wire _w854_ ;
	wire _w853_ ;
	wire _w852_ ;
	wire _w851_ ;
	wire _w850_ ;
	wire _w849_ ;
	wire _w848_ ;
	wire _w847_ ;
	wire _w846_ ;
	wire _w845_ ;
	wire _w844_ ;
	wire _w843_ ;
	wire _w842_ ;
	wire _w841_ ;
	wire _w840_ ;
	wire _w839_ ;
	wire _w838_ ;
	wire _w837_ ;
	wire _w836_ ;
	wire _w835_ ;
	wire _w834_ ;
	wire _w833_ ;
	wire _w832_ ;
	wire _w831_ ;
	wire _w830_ ;
	wire _w829_ ;
	wire _w828_ ;
	wire _w827_ ;
	wire _w826_ ;
	wire _w825_ ;
	wire _w824_ ;
	wire _w823_ ;
	wire _w822_ ;
	wire _w821_ ;
	wire _w820_ ;
	wire _w819_ ;
	wire _w818_ ;
	wire _w817_ ;
	wire _w816_ ;
	wire _w815_ ;
	wire _w814_ ;
	wire _w813_ ;
	wire _w812_ ;
	wire _w811_ ;
	wire _w810_ ;
	wire _w809_ ;
	wire _w808_ ;
	wire _w807_ ;
	wire _w806_ ;
	wire _w805_ ;
	wire _w804_ ;
	wire _w803_ ;
	wire _w802_ ;
	wire _w801_ ;
	wire _w800_ ;
	wire _w799_ ;
	wire _w798_ ;
	wire _w797_ ;
	wire _w796_ ;
	wire _w795_ ;
	wire _w794_ ;
	wire _w793_ ;
	wire _w792_ ;
	wire _w791_ ;
	wire _w790_ ;
	wire _w789_ ;
	wire _w788_ ;
	wire _w787_ ;
	wire _w786_ ;
	wire _w785_ ;
	wire _w784_ ;
	wire _w783_ ;
	wire _w782_ ;
	wire _w781_ ;
	wire _w780_ ;
	wire _w779_ ;
	wire _w778_ ;
	wire _w777_ ;
	wire _w776_ ;
	wire _w775_ ;
	wire _w774_ ;
	wire _w773_ ;
	wire _w772_ ;
	wire _w771_ ;
	wire _w770_ ;
	wire _w769_ ;
	wire _w768_ ;
	wire _w767_ ;
	wire _w766_ ;
	wire _w765_ ;
	wire _w764_ ;
	wire _w763_ ;
	wire _w762_ ;
	wire _w761_ ;
	wire _w760_ ;
	wire _w759_ ;
	wire _w758_ ;
	wire _w757_ ;
	wire _w756_ ;
	wire _w755_ ;
	wire _w754_ ;
	wire _w753_ ;
	wire _w752_ ;
	wire _w751_ ;
	wire _w750_ ;
	wire _w749_ ;
	wire _w748_ ;
	wire _w747_ ;
	wire _w746_ ;
	wire _w745_ ;
	wire _w744_ ;
	wire _w743_ ;
	wire _w742_ ;
	wire _w741_ ;
	wire _w740_ ;
	wire _w739_ ;
	wire _w738_ ;
	wire _w737_ ;
	wire _w736_ ;
	wire _w735_ ;
	wire _w734_ ;
	wire _w733_ ;
	wire _w732_ ;
	wire _w731_ ;
	wire _w730_ ;
	wire _w729_ ;
	wire _w728_ ;
	wire _w727_ ;
	wire _w726_ ;
	wire _w725_ ;
	wire _w724_ ;
	wire _w723_ ;
	wire _w722_ ;
	wire _w721_ ;
	wire _w720_ ;
	wire _w719_ ;
	wire _w718_ ;
	wire _w717_ ;
	wire _w716_ ;
	wire _w715_ ;
	wire _w714_ ;
	wire _w713_ ;
	wire _w712_ ;
	wire _w711_ ;
	wire _w710_ ;
	wire _w709_ ;
	wire _w708_ ;
	wire _w707_ ;
	wire _w706_ ;
	wire _w705_ ;
	wire _w704_ ;
	wire _w703_ ;
	wire _w702_ ;
	wire _w701_ ;
	wire _w700_ ;
	wire _w699_ ;
	wire _w698_ ;
	wire _w697_ ;
	wire _w696_ ;
	wire _w695_ ;
	wire _w694_ ;
	wire _w693_ ;
	wire _w692_ ;
	wire _w691_ ;
	wire _w690_ ;
	wire _w689_ ;
	wire _w688_ ;
	wire _w687_ ;
	wire _w686_ ;
	wire _w685_ ;
	wire _w684_ ;
	wire _w683_ ;
	wire _w682_ ;
	wire _w681_ ;
	wire _w680_ ;
	wire _w679_ ;
	wire _w678_ ;
	wire _w677_ ;
	wire _w676_ ;
	wire _w675_ ;
	wire _w674_ ;
	wire _w673_ ;
	wire _w672_ ;
	wire _w671_ ;
	wire _w670_ ;
	wire _w669_ ;
	wire _w668_ ;
	wire _w667_ ;
	wire _w666_ ;
	wire _w381_ ;
	wire _w380_ ;
	wire _w379_ ;
	wire _w378_ ;
	wire _w377_ ;
	wire _w376_ ;
	wire _w375_ ;
	wire _w374_ ;
	wire _w373_ ;
	wire _w372_ ;
	wire _w371_ ;
	wire _w370_ ;
	wire _w369_ ;
	wire _w368_ ;
	wire _w367_ ;
	wire _w366_ ;
	wire _w365_ ;
	wire _w364_ ;
	wire _w363_ ;
	wire _w362_ ;
	wire _w361_ ;
	wire _w360_ ;
	wire _w359_ ;
	wire _w358_ ;
	wire _w357_ ;
	wire _w356_ ;
	wire _w355_ ;
	wire _w354_ ;
	wire _w353_ ;
	wire _w352_ ;
	wire _w351_ ;
	wire _w350_ ;
	wire _w349_ ;
	wire _w348_ ;
	wire _w347_ ;
	wire _w346_ ;
	wire _w345_ ;
	wire _w344_ ;
	wire _w343_ ;
	wire _w342_ ;
	wire _w341_ ;
	wire _w340_ ;
	wire _w339_ ;
	wire _w338_ ;
	wire _w337_ ;
	wire _w336_ ;
	wire _w335_ ;
	wire _w334_ ;
	wire _w333_ ;
	wire _w332_ ;
	wire _w331_ ;
	wire _w330_ ;
	wire _w329_ ;
	wire _w328_ ;
	wire _w327_ ;
	wire _w326_ ;
	wire _w325_ ;
	wire _w324_ ;
	wire _w323_ ;
	wire _w322_ ;
	wire _w321_ ;
	wire _w320_ ;
	wire _w319_ ;
	wire _w318_ ;
	wire _w317_ ;
	wire _w316_ ;
	wire _w315_ ;
	wire _w314_ ;
	wire _w313_ ;
	wire _w312_ ;
	wire _w311_ ;
	wire _w310_ ;
	wire _w309_ ;
	wire _w308_ ;
	wire _w307_ ;
	wire _w306_ ;
	wire _w305_ ;
	wire _w304_ ;
	wire _w303_ ;
	wire _w302_ ;
	wire _w301_ ;
	wire _w300_ ;
	wire _w299_ ;
	wire _w298_ ;
	wire _w297_ ;
	wire _w296_ ;
	wire _w295_ ;
	wire _w294_ ;
	wire _w293_ ;
	wire _w292_ ;
	wire _w291_ ;
	wire _w290_ ;
	wire _w289_ ;
	wire _w288_ ;
	wire _w287_ ;
	wire _w286_ ;
	wire _w285_ ;
	wire _w284_ ;
	wire _w283_ ;
	wire _w282_ ;
	wire _w281_ ;
	wire _w280_ ;
	wire _w279_ ;
	wire _w278_ ;
	wire _w277_ ;
	wire _w276_ ;
	wire _w275_ ;
	wire _w274_ ;
	wire _w273_ ;
	wire _w272_ ;
	wire _w271_ ;
	wire _w270_ ;
	wire _w269_ ;
	wire _w268_ ;
	wire _w267_ ;
	wire _w266_ ;
	wire _w265_ ;
	wire _w264_ ;
	wire _w263_ ;
	wire _w262_ ;
	wire _w261_ ;
	wire _w260_ ;
	wire _w259_ ;
	wire _w258_ ;
	wire _w257_ ;
	wire _w256_ ;
	wire _w255_ ;
	wire _w254_ ;
	wire _w253_ ;
	wire _w252_ ;
	wire _w183_ ;
	wire _w182_ ;
	wire _w181_ ;
	wire _w180_ ;
	wire _w179_ ;
	wire _w178_ ;
	wire _w177_ ;
	wire _w176_ ;
	wire _w175_ ;
	wire _w174_ ;
	wire _w173_ ;
	wire _w172_ ;
	wire _w171_ ;
	wire _w170_ ;
	wire _w169_ ;
	wire _w168_ ;
	wire _w167_ ;
	wire _w166_ ;
	wire _w165_ ;
	wire _w164_ ;
	wire _w163_ ;
	wire _w162_ ;
	wire _w161_ ;
	wire _w160_ ;
	wire _w159_ ;
	wire _w158_ ;
	wire _w157_ ;
	wire _w156_ ;
	wire _w155_ ;
	wire _w154_ ;
	wire _w137_ ;
	wire _w136_ ;
	wire _w135_ ;
	wire _w134_ ;
	wire _w133_ ;
	wire _w132_ ;
	wire _w131_ ;
	wire _w130_ ;
	wire _w129_ ;
	wire _w128_ ;
	wire _w127_ ;
	wire _w126_ ;
	wire _w125_ ;
	wire _w138_ ;
	wire _w139_ ;
	wire _w140_ ;
	wire _w141_ ;
	wire _w142_ ;
	wire _w143_ ;
	wire _w144_ ;
	wire _w145_ ;
	wire _w146_ ;
	wire _w147_ ;
	wire _w148_ ;
	wire _w149_ ;
	wire _w150_ ;
	wire _w151_ ;
	wire _w152_ ;
	wire _w153_ ;
	wire _w184_ ;
	wire _w185_ ;
	wire _w186_ ;
	wire _w187_ ;
	wire _w188_ ;
	wire _w189_ ;
	wire _w190_ ;
	wire _w191_ ;
	wire _w192_ ;
	wire _w193_ ;
	wire _w194_ ;
	wire _w195_ ;
	wire _w196_ ;
	wire _w197_ ;
	wire _w198_ ;
	wire _w199_ ;
	wire _w200_ ;
	wire _w201_ ;
	wire _w202_ ;
	wire _w203_ ;
	wire _w204_ ;
	wire _w205_ ;
	wire _w206_ ;
	wire _w207_ ;
	wire _w208_ ;
	wire _w209_ ;
	wire _w210_ ;
	wire _w211_ ;
	wire _w212_ ;
	wire _w213_ ;
	wire _w214_ ;
	wire _w215_ ;
	wire _w216_ ;
	wire _w217_ ;
	wire _w218_ ;
	wire _w219_ ;
	wire _w220_ ;
	wire _w221_ ;
	wire _w222_ ;
	wire _w223_ ;
	wire _w224_ ;
	wire _w225_ ;
	wire _w226_ ;
	wire _w227_ ;
	wire _w228_ ;
	wire _w229_ ;
	wire _w230_ ;
	wire _w231_ ;
	wire _w232_ ;
	wire _w233_ ;
	wire _w234_ ;
	wire _w235_ ;
	wire _w236_ ;
	wire _w237_ ;
	wire _w238_ ;
	wire _w239_ ;
	wire _w240_ ;
	wire _w241_ ;
	wire _w242_ ;
	wire _w243_ ;
	wire _w244_ ;
	wire _w245_ ;
	wire _w246_ ;
	wire _w247_ ;
	wire _w248_ ;
	wire _w249_ ;
	wire _w250_ ;
	wire _w251_ ;
	wire _w382_ ;
	wire _w383_ ;
	wire _w384_ ;
	wire _w385_ ;
	wire _w386_ ;
	wire _w387_ ;
	wire _w388_ ;
	wire _w389_ ;
	wire _w390_ ;
	wire _w391_ ;
	wire _w392_ ;
	wire _w393_ ;
	wire _w394_ ;
	wire _w395_ ;
	wire _w396_ ;
	wire _w397_ ;
	wire _w398_ ;
	wire _w399_ ;
	wire _w400_ ;
	wire _w401_ ;
	wire _w402_ ;
	wire _w403_ ;
	wire _w404_ ;
	wire _w405_ ;
	wire _w406_ ;
	wire _w407_ ;
	wire _w408_ ;
	wire _w409_ ;
	wire _w410_ ;
	wire _w411_ ;
	wire _w412_ ;
	wire _w413_ ;
	wire _w414_ ;
	wire _w415_ ;
	wire _w416_ ;
	wire _w417_ ;
	wire _w418_ ;
	wire _w419_ ;
	wire _w420_ ;
	wire _w421_ ;
	wire _w422_ ;
	wire _w423_ ;
	wire _w424_ ;
	wire _w425_ ;
	wire _w426_ ;
	wire _w427_ ;
	wire _w428_ ;
	wire _w429_ ;
	wire _w430_ ;
	wire _w431_ ;
	wire _w432_ ;
	wire _w433_ ;
	wire _w434_ ;
	wire _w435_ ;
	wire _w436_ ;
	wire _w437_ ;
	wire _w438_ ;
	wire _w439_ ;
	wire _w440_ ;
	wire _w441_ ;
	wire _w442_ ;
	wire _w443_ ;
	wire _w444_ ;
	wire _w445_ ;
	wire _w446_ ;
	wire _w447_ ;
	wire _w448_ ;
	wire _w449_ ;
	wire _w450_ ;
	wire _w451_ ;
	wire _w452_ ;
	wire _w453_ ;
	wire _w454_ ;
	wire _w455_ ;
	wire _w456_ ;
	wire _w457_ ;
	wire _w458_ ;
	wire _w459_ ;
	wire _w460_ ;
	wire _w461_ ;
	wire _w462_ ;
	wire _w463_ ;
	wire _w464_ ;
	wire _w465_ ;
	wire _w466_ ;
	wire _w467_ ;
	wire _w468_ ;
	wire _w469_ ;
	wire _w470_ ;
	wire _w471_ ;
	wire _w472_ ;
	wire _w473_ ;
	wire _w474_ ;
	wire _w475_ ;
	wire _w476_ ;
	wire _w477_ ;
	wire _w478_ ;
	wire _w479_ ;
	wire _w480_ ;
	wire _w481_ ;
	wire _w482_ ;
	wire _w483_ ;
	wire _w484_ ;
	wire _w485_ ;
	wire _w486_ ;
	wire _w487_ ;
	wire _w488_ ;
	wire _w489_ ;
	wire _w490_ ;
	wire _w491_ ;
	wire _w492_ ;
	wire _w493_ ;
	wire _w494_ ;
	wire _w495_ ;
	wire _w496_ ;
	wire _w497_ ;
	wire _w498_ ;
	wire _w499_ ;
	wire _w500_ ;
	wire _w501_ ;
	wire _w502_ ;
	wire _w503_ ;
	wire _w504_ ;
	wire _w505_ ;
	wire _w506_ ;
	wire _w507_ ;
	wire _w508_ ;
	wire _w509_ ;
	wire _w510_ ;
	wire _w511_ ;
	wire _w512_ ;
	wire _w513_ ;
	wire _w514_ ;
	wire _w515_ ;
	wire _w516_ ;
	wire _w517_ ;
	wire _w518_ ;
	wire _w519_ ;
	wire _w520_ ;
	wire _w521_ ;
	wire _w522_ ;
	wire _w523_ ;
	wire _w524_ ;
	wire _w525_ ;
	wire _w526_ ;
	wire _w527_ ;
	wire _w528_ ;
	wire _w529_ ;
	wire _w530_ ;
	wire _w531_ ;
	wire _w532_ ;
	wire _w533_ ;
	wire _w534_ ;
	wire _w535_ ;
	wire _w536_ ;
	wire _w537_ ;
	wire _w538_ ;
	wire _w539_ ;
	wire _w540_ ;
	wire _w541_ ;
	wire _w542_ ;
	wire _w543_ ;
	wire _w544_ ;
	wire _w545_ ;
	wire _w546_ ;
	wire _w547_ ;
	wire _w548_ ;
	wire _w549_ ;
	wire _w550_ ;
	wire _w551_ ;
	wire _w552_ ;
	wire _w553_ ;
	wire _w554_ ;
	wire _w555_ ;
	wire _w556_ ;
	wire _w557_ ;
	wire _w558_ ;
	wire _w559_ ;
	wire _w560_ ;
	wire _w561_ ;
	wire _w562_ ;
	wire _w563_ ;
	wire _w564_ ;
	wire _w565_ ;
	wire _w566_ ;
	wire _w567_ ;
	wire _w568_ ;
	wire _w569_ ;
	wire _w570_ ;
	wire _w571_ ;
	wire _w572_ ;
	wire _w573_ ;
	wire _w574_ ;
	wire _w575_ ;
	wire _w576_ ;
	wire _w577_ ;
	wire _w578_ ;
	wire _w579_ ;
	wire _w580_ ;
	wire _w581_ ;
	wire _w582_ ;
	wire _w583_ ;
	wire _w584_ ;
	wire _w585_ ;
	wire _w586_ ;
	wire _w587_ ;
	wire _w588_ ;
	wire _w589_ ;
	wire _w590_ ;
	wire _w591_ ;
	wire _w592_ ;
	wire _w593_ ;
	wire _w594_ ;
	wire _w595_ ;
	wire _w596_ ;
	wire _w597_ ;
	wire _w598_ ;
	wire _w599_ ;
	wire _w600_ ;
	wire _w601_ ;
	wire _w602_ ;
	wire _w603_ ;
	wire _w604_ ;
	wire _w605_ ;
	wire _w606_ ;
	wire _w607_ ;
	wire _w608_ ;
	wire _w609_ ;
	wire _w610_ ;
	wire _w611_ ;
	wire _w612_ ;
	wire _w613_ ;
	wire _w614_ ;
	wire _w615_ ;
	wire _w616_ ;
	wire _w617_ ;
	wire _w618_ ;
	wire _w619_ ;
	wire _w620_ ;
	wire _w621_ ;
	wire _w622_ ;
	wire _w623_ ;
	wire _w624_ ;
	wire _w625_ ;
	wire _w626_ ;
	wire _w627_ ;
	wire _w628_ ;
	wire _w629_ ;
	wire _w630_ ;
	wire _w631_ ;
	wire _w632_ ;
	wire _w633_ ;
	wire _w634_ ;
	wire _w635_ ;
	wire _w636_ ;
	wire _w637_ ;
	wire _w638_ ;
	wire _w639_ ;
	wire _w640_ ;
	wire _w641_ ;
	wire _w642_ ;
	wire _w643_ ;
	wire _w644_ ;
	wire _w645_ ;
	wire _w646_ ;
	wire _w647_ ;
	wire _w648_ ;
	wire _w649_ ;
	wire _w650_ ;
	wire _w651_ ;
	wire _w652_ ;
	wire _w653_ ;
	wire _w654_ ;
	wire _w655_ ;
	wire _w656_ ;
	wire _w657_ ;
	wire _w658_ ;
	wire _w659_ ;
	wire _w660_ ;
	wire _w661_ ;
	wire _w662_ ;
	wire _w663_ ;
	wire _w664_ ;
	wire _w665_ ;
	LUT2 #(
		.INIT('h2)
	) name0 (
		\count_reg[0]/NET0131 ,
		\count_reg[1]/NET0131 ,
		_w125_
	);
	LUT2 #(
		.INIT('h4)
	) name1 (
		\count_reg[0]/NET0131 ,
		\count_reg[1]/NET0131 ,
		_w126_
	);
	LUT2 #(
		.INIT('h1)
	) name2 (
		_w125_,
		_w126_,
		_w127_
	);
	LUT2 #(
		.INIT('h8)
	) name3 (
		\max_reg[3]/NET0131 ,
		\scan_reg[3]/NET0131 ,
		_w128_
	);
	LUT2 #(
		.INIT('h1)
	) name4 (
		\max_reg[3]/NET0131 ,
		\scan_reg[3]/NET0131 ,
		_w129_
	);
	LUT2 #(
		.INIT('h1)
	) name5 (
		_w128_,
		_w129_,
		_w130_
	);
	LUT2 #(
		.INIT('h2)
	) name6 (
		\max_reg[1]/NET0131 ,
		\scan_reg[1]/NET0131 ,
		_w131_
	);
	LUT2 #(
		.INIT('h4)
	) name7 (
		\max_reg[1]/NET0131 ,
		\scan_reg[1]/NET0131 ,
		_w132_
	);
	LUT2 #(
		.INIT('h1)
	) name8 (
		\max_reg[4]/NET0131 ,
		\scan_reg[4]/NET0131 ,
		_w133_
	);
	LUT2 #(
		.INIT('h8)
	) name9 (
		\max_reg[4]/NET0131 ,
		\scan_reg[4]/NET0131 ,
		_w134_
	);
	LUT2 #(
		.INIT('h1)
	) name10 (
		_w133_,
		_w134_,
		_w135_
	);
	LUT2 #(
		.INIT('h1)
	) name11 (
		\max_reg[2]/NET0131 ,
		\scan_reg[2]/NET0131 ,
		_w136_
	);
	LUT2 #(
		.INIT('h8)
	) name12 (
		\max_reg[2]/NET0131 ,
		\scan_reg[2]/NET0131 ,
		_w137_
	);
	LUT2 #(
		.INIT('h1)
	) name13 (
		_w136_,
		_w137_,
		_w138_
	);
	LUT2 #(
		.INIT('h1)
	) name14 (
		\max_reg[0]/NET0131 ,
		\scan_reg[0]/NET0131 ,
		_w139_
	);
	LUT2 #(
		.INIT('h8)
	) name15 (
		\max_reg[0]/NET0131 ,
		\scan_reg[0]/NET0131 ,
		_w140_
	);
	LUT2 #(
		.INIT('h1)
	) name16 (
		_w139_,
		_w140_,
		_w141_
	);
	LUT2 #(
		.INIT('h1)
	) name17 (
		_w131_,
		_w132_,
		_w142_
	);
	LUT2 #(
		.INIT('h4)
	) name18 (
		_w135_,
		_w142_,
		_w143_
	);
	LUT2 #(
		.INIT('h1)
	) name19 (
		_w138_,
		_w141_,
		_w144_
	);
	LUT2 #(
		.INIT('h8)
	) name20 (
		_w143_,
		_w144_,
		_w145_
	);
	LUT2 #(
		.INIT('h4)
	) name21 (
		_w130_,
		_w145_,
		_w146_
	);
	LUT2 #(
		.INIT('h4)
	) name22 (
		\scan_reg[1]/NET0131 ,
		_w146_,
		_w147_
	);
	LUT2 #(
		.INIT('h8)
	) name23 (
		\scan_reg[0]/NET0131 ,
		\scan_reg[1]/NET0131 ,
		_w148_
	);
	LUT2 #(
		.INIT('h1)
	) name24 (
		\scan_reg[0]/NET0131 ,
		\scan_reg[1]/NET0131 ,
		_w149_
	);
	LUT2 #(
		.INIT('h1)
	) name25 (
		_w148_,
		_w149_,
		_w150_
	);
	LUT2 #(
		.INIT('h1)
	) name26 (
		_w146_,
		_w150_,
		_w151_
	);
	LUT2 #(
		.INIT('h1)
	) name27 (
		\gamma_reg[0]/NET0131 ,
		start_pad,
		_w152_
	);
	LUT2 #(
		.INIT('h2)
	) name28 (
		\gamma_reg[2]/NET0131 ,
		start_pad,
		_w153_
	);
	LUT2 #(
		.INIT('h2)
	) name29 (
		\gamma_reg[1]/NET0131 ,
		start_pad,
		_w154_
	);
	LUT2 #(
		.INIT('h2)
	) name30 (
		_w153_,
		_w154_,
		_w155_
	);
	LUT2 #(
		.INIT('h2)
	) name31 (
		\gamma_reg[4]/NET0131 ,
		start_pad,
		_w156_
	);
	LUT2 #(
		.INIT('h2)
	) name32 (
		\gamma_reg[3]/NET0131 ,
		start_pad,
		_w157_
	);
	LUT2 #(
		.INIT('h4)
	) name33 (
		_w156_,
		_w157_,
		_w158_
	);
	LUT2 #(
		.INIT('h8)
	) name34 (
		_w155_,
		_w158_,
		_w159_
	);
	LUT2 #(
		.INIT('h4)
	) name35 (
		_w152_,
		_w159_,
		_w160_
	);
	LUT2 #(
		.INIT('h1)
	) name36 (
		\count_reg[0]1198/NET0131 ,
		\count_reg[1]1200/NET0131 ,
		_w161_
	);
	LUT2 #(
		.INIT('h4)
	) name37 (
		\count_reg[2]/NET0131 ,
		_w161_,
		_w162_
	);
	LUT2 #(
		.INIT('h1)
	) name38 (
		\count_reg[3]/NET0131 ,
		\count_reg[4]/NET0131 ,
		_w163_
	);
	LUT2 #(
		.INIT('h8)
	) name39 (
		_w162_,
		_w163_,
		_w164_
	);
	LUT2 #(
		.INIT('h4)
	) name40 (
		\count_reg[5]/NET0131 ,
		_w164_,
		_w165_
	);
	LUT2 #(
		.INIT('h8)
	) name41 (
		_w160_,
		_w165_,
		_w166_
	);
	LUT2 #(
		.INIT('h4)
	) name42 (
		_w147_,
		_w166_,
		_w167_
	);
	LUT2 #(
		.INIT('h4)
	) name43 (
		_w151_,
		_w167_,
		_w168_
	);
	LUT2 #(
		.INIT('h1)
	) name44 (
		_w156_,
		_w157_,
		_w169_
	);
	LUT2 #(
		.INIT('h8)
	) name45 (
		_w155_,
		_w169_,
		_w170_
	);
	LUT2 #(
		.INIT('h2)
	) name46 (
		_w156_,
		_w157_,
		_w171_
	);
	LUT2 #(
		.INIT('h8)
	) name47 (
		_w153_,
		_w154_,
		_w172_
	);
	LUT2 #(
		.INIT('h8)
	) name48 (
		_w171_,
		_w172_,
		_w173_
	);
	LUT2 #(
		.INIT('h1)
	) name49 (
		_w170_,
		_w173_,
		_w174_
	);
	LUT2 #(
		.INIT('h4)
	) name50 (
		_w153_,
		_w154_,
		_w175_
	);
	LUT2 #(
		.INIT('h8)
	) name51 (
		_w158_,
		_w175_,
		_w176_
	);
	LUT2 #(
		.INIT('h4)
	) name52 (
		_w152_,
		_w176_,
		_w177_
	);
	LUT2 #(
		.INIT('h8)
	) name53 (
		_w169_,
		_w172_,
		_w178_
	);
	LUT2 #(
		.INIT('h4)
	) name54 (
		\gamma_reg[0]/NET0131 ,
		_w178_,
		_w179_
	);
	LUT2 #(
		.INIT('h1)
	) name55 (
		_w177_,
		_w179_,
		_w180_
	);
	LUT2 #(
		.INIT('h2)
	) name56 (
		_w160_,
		_w165_,
		_w181_
	);
	LUT2 #(
		.INIT('h8)
	) name57 (
		_w169_,
		_w175_,
		_w182_
	);
	LUT2 #(
		.INIT('h4)
	) name58 (
		_w152_,
		_w182_,
		_w183_
	);
	LUT2 #(
		.INIT('h2)
	) name59 (
		_w174_,
		_w183_,
		_w184_
	);
	LUT2 #(
		.INIT('h8)
	) name60 (
		_w180_,
		_w184_,
		_w185_
	);
	LUT2 #(
		.INIT('h4)
	) name61 (
		_w181_,
		_w185_,
		_w186_
	);
	LUT2 #(
		.INIT('h1)
	) name62 (
		_w153_,
		_w154_,
		_w187_
	);
	LUT2 #(
		.INIT('h4)
	) name63 (
		_w171_,
		_w187_,
		_w188_
	);
	LUT2 #(
		.INIT('h8)
	) name64 (
		_w152_,
		_w159_,
		_w189_
	);
	LUT2 #(
		.INIT('h8)
	) name65 (
		_w158_,
		_w172_,
		_w190_
	);
	LUT2 #(
		.INIT('h4)
	) name66 (
		\gamma_reg[0]/NET0131 ,
		_w190_,
		_w191_
	);
	LUT2 #(
		.INIT('h1)
	) name67 (
		_w189_,
		_w191_,
		_w192_
	);
	LUT2 #(
		.INIT('h4)
	) name68 (
		\gamma_reg[0]/NET0131 ,
		_w171_,
		_w193_
	);
	LUT2 #(
		.INIT('h8)
	) name69 (
		_w155_,
		_w193_,
		_w194_
	);
	LUT2 #(
		.INIT('h8)
	) name70 (
		\gamma_reg[0]/NET0131 ,
		_w190_,
		_w195_
	);
	LUT2 #(
		.INIT('h1)
	) name71 (
		_w194_,
		_w195_,
		_w196_
	);
	LUT2 #(
		.INIT('h8)
	) name72 (
		\gamma_reg[0]/NET0131 ,
		_w171_,
		_w197_
	);
	LUT2 #(
		.INIT('h4)
	) name73 (
		_w153_,
		_w197_,
		_w198_
	);
	LUT2 #(
		.INIT('h2)
	) name74 (
		_w196_,
		_w198_,
		_w199_
	);
	LUT2 #(
		.INIT('h8)
	) name75 (
		_w175_,
		_w193_,
		_w200_
	);
	LUT2 #(
		.INIT('h8)
	) name76 (
		_w155_,
		_w197_,
		_w201_
	);
	LUT2 #(
		.INIT('h1)
	) name77 (
		_w200_,
		_w201_,
		_w202_
	);
	LUT2 #(
		.INIT('h8)
	) name78 (
		_w152_,
		_w176_,
		_w203_
	);
	LUT2 #(
		.INIT('h8)
	) name79 (
		_w187_,
		_w193_,
		_w204_
	);
	LUT2 #(
		.INIT('h1)
	) name80 (
		_w203_,
		_w204_,
		_w205_
	);
	LUT2 #(
		.INIT('h4)
	) name81 (
		_w188_,
		_w192_,
		_w206_
	);
	LUT2 #(
		.INIT('h8)
	) name82 (
		_w202_,
		_w205_,
		_w207_
	);
	LUT2 #(
		.INIT('h8)
	) name83 (
		_w206_,
		_w207_,
		_w208_
	);
	LUT2 #(
		.INIT('h8)
	) name84 (
		_w199_,
		_w208_,
		_w209_
	);
	LUT2 #(
		.INIT('h8)
	) name85 (
		_w186_,
		_w209_,
		_w210_
	);
	LUT2 #(
		.INIT('h2)
	) name86 (
		\scan_reg[1]/NET0131 ,
		_w210_,
		_w211_
	);
	LUT2 #(
		.INIT('h2)
	) name87 (
		\scan_reg[1]/NET0131 ,
		_w165_,
		_w212_
	);
	LUT2 #(
		.INIT('h4)
	) name88 (
		_w146_,
		_w165_,
		_w213_
	);
	LUT2 #(
		.INIT('h8)
	) name89 (
		_w150_,
		_w213_,
		_w214_
	);
	LUT2 #(
		.INIT('h1)
	) name90 (
		_w212_,
		_w214_,
		_w215_
	);
	LUT2 #(
		.INIT('h8)
	) name91 (
		\gamma_reg[0]/NET0131 ,
		_w178_,
		_w216_
	);
	LUT2 #(
		.INIT('h4)
	) name92 (
		_w215_,
		_w216_,
		_w217_
	);
	LUT2 #(
		.INIT('h1)
	) name93 (
		_w168_,
		_w217_,
		_w218_
	);
	LUT2 #(
		.INIT('h4)
	) name94 (
		_w211_,
		_w218_,
		_w219_
	);
	LUT2 #(
		.INIT('h8)
	) name95 (
		_w158_,
		_w187_,
		_w220_
	);
	LUT2 #(
		.INIT('h8)
	) name96 (
		_w152_,
		_w220_,
		_w221_
	);
	LUT2 #(
		.INIT('h1)
	) name97 (
		_w183_,
		_w221_,
		_w222_
	);
	LUT2 #(
		.INIT('h2)
	) name98 (
		\scan_reg[0]/NET0131 ,
		_w222_,
		_w223_
	);
	LUT2 #(
		.INIT('h8)
	) name99 (
		_w187_,
		_w197_,
		_w224_
	);
	LUT2 #(
		.INIT('h8)
	) name100 (
		_w152_,
		_w182_,
		_w225_
	);
	LUT2 #(
		.INIT('h1)
	) name101 (
		_w224_,
		_w225_,
		_w226_
	);
	LUT2 #(
		.INIT('h2)
	) name102 (
		\max_reg[0]/NET0131 ,
		_w226_,
		_w227_
	);
	LUT2 #(
		.INIT('h8)
	) name103 (
		_w169_,
		_w187_,
		_w228_
	);
	LUT2 #(
		.INIT('h4)
	) name104 (
		_w152_,
		_w228_,
		_w229_
	);
	LUT2 #(
		.INIT('h8)
	) name105 (
		_w152_,
		_w170_,
		_w230_
	);
	LUT2 #(
		.INIT('h8)
	) name106 (
		_w175_,
		_w197_,
		_w231_
	);
	LUT2 #(
		.INIT('h4)
	) name107 (
		_w153_,
		_w193_,
		_w232_
	);
	LUT2 #(
		.INIT('h1)
	) name108 (
		_w160_,
		_w232_,
		_w233_
	);
	LUT2 #(
		.INIT('h1)
	) name109 (
		_w190_,
		_w216_,
		_w234_
	);
	LUT2 #(
		.INIT('h8)
	) name110 (
		\gamma_reg[3]/NET0131 ,
		_w156_,
		_w235_
	);
	LUT2 #(
		.INIT('h8)
	) name111 (
		_w187_,
		_w235_,
		_w236_
	);
	LUT2 #(
		.INIT('h8)
	) name112 (
		_w152_,
		_w236_,
		_w237_
	);
	LUT2 #(
		.INIT('h1)
	) name113 (
		_w201_,
		_w203_,
		_w238_
	);
	LUT2 #(
		.INIT('h4)
	) name114 (
		_w237_,
		_w238_,
		_w239_
	);
	LUT2 #(
		.INIT('h1)
	) name115 (
		_w179_,
		_w189_,
		_w240_
	);
	LUT2 #(
		.INIT('h8)
	) name116 (
		_w152_,
		_w228_,
		_w241_
	);
	LUT2 #(
		.INIT('h1)
	) name117 (
		_w177_,
		_w241_,
		_w242_
	);
	LUT2 #(
		.INIT('h8)
	) name118 (
		_w240_,
		_w242_,
		_w243_
	);
	LUT2 #(
		.INIT('h8)
	) name119 (
		\gamma_reg[0]/NET0131 ,
		_w170_,
		_w244_
	);
	LUT2 #(
		.INIT('h4)
	) name120 (
		_w152_,
		_w220_,
		_w245_
	);
	LUT2 #(
		.INIT('h1)
	) name121 (
		_w244_,
		_w245_,
		_w246_
	);
	LUT2 #(
		.INIT('h8)
	) name122 (
		_w152_,
		_w173_,
		_w247_
	);
	LUT2 #(
		.INIT('h1)
	) name123 (
		_w194_,
		_w247_,
		_w248_
	);
	LUT2 #(
		.INIT('h1)
	) name124 (
		_w173_,
		_w236_,
		_w249_
	);
	LUT2 #(
		.INIT('h1)
	) name125 (
		_w152_,
		_w249_,
		_w250_
	);
	LUT2 #(
		.INIT('h2)
	) name126 (
		_w248_,
		_w250_,
		_w251_
	);
	LUT2 #(
		.INIT('h1)
	) name127 (
		_w229_,
		_w230_,
		_w252_
	);
	LUT2 #(
		.INIT('h4)
	) name128 (
		_w231_,
		_w252_,
		_w253_
	);
	LUT2 #(
		.INIT('h8)
	) name129 (
		_w233_,
		_w234_,
		_w254_
	);
	LUT2 #(
		.INIT('h8)
	) name130 (
		_w246_,
		_w254_,
		_w255_
	);
	LUT2 #(
		.INIT('h8)
	) name131 (
		_w239_,
		_w253_,
		_w256_
	);
	LUT2 #(
		.INIT('h8)
	) name132 (
		_w243_,
		_w251_,
		_w257_
	);
	LUT2 #(
		.INIT('h8)
	) name133 (
		_w256_,
		_w257_,
		_w258_
	);
	LUT2 #(
		.INIT('h8)
	) name134 (
		_w255_,
		_w258_,
		_w259_
	);
	LUT2 #(
		.INIT('h2)
	) name135 (
		\address_reg[0]/NET0131 ,
		_w259_,
		_w260_
	);
	LUT2 #(
		.INIT('h1)
	) name136 (
		_w223_,
		_w227_,
		_w261_
	);
	LUT2 #(
		.INIT('h4)
	) name137 (
		_w260_,
		_w261_,
		_w262_
	);
	LUT2 #(
		.INIT('h4)
	) name138 (
		\count_reg[5]/NET0131 ,
		_w163_,
		_w263_
	);
	LUT2 #(
		.INIT('h2)
	) name139 (
		\count_reg[3]/NET0131 ,
		_w162_,
		_w264_
	);
	LUT2 #(
		.INIT('h4)
	) name140 (
		\count_reg[3]/NET0131 ,
		_w162_,
		_w265_
	);
	LUT2 #(
		.INIT('h1)
	) name141 (
		_w264_,
		_w265_,
		_w266_
	);
	LUT2 #(
		.INIT('h1)
	) name142 (
		_w263_,
		_w266_,
		_w267_
	);
	LUT2 #(
		.INIT('h8)
	) name143 (
		_w146_,
		_w165_,
		_w268_
	);
	LUT2 #(
		.INIT('h8)
	) name144 (
		\max_reg[0]/NET0131 ,
		\max_reg[1]/NET0131 ,
		_w269_
	);
	LUT2 #(
		.INIT('h8)
	) name145 (
		\max_reg[2]/NET0131 ,
		_w269_,
		_w270_
	);
	LUT2 #(
		.INIT('h8)
	) name146 (
		\max_reg[3]/NET0131 ,
		_w270_,
		_w271_
	);
	LUT2 #(
		.INIT('h8)
	) name147 (
		\max_reg[4]/NET0131 ,
		_w271_,
		_w272_
	);
	LUT2 #(
		.INIT('h1)
	) name148 (
		\count_reg[3]/NET0131 ,
		_w272_,
		_w273_
	);
	LUT2 #(
		.INIT('h2)
	) name149 (
		_w268_,
		_w273_,
		_w274_
	);
	LUT2 #(
		.INIT('h1)
	) name150 (
		_w267_,
		_w274_,
		_w275_
	);
	LUT2 #(
		.INIT('h2)
	) name151 (
		_w160_,
		_w275_,
		_w276_
	);
	LUT2 #(
		.INIT('h1)
	) name152 (
		_w177_,
		_w191_,
		_w277_
	);
	LUT2 #(
		.INIT('h1)
	) name153 (
		_w183_,
		_w229_,
		_w278_
	);
	LUT2 #(
		.INIT('h1)
	) name154 (
		_w200_,
		_w230_,
		_w279_
	);
	LUT2 #(
		.INIT('h8)
	) name155 (
		_w278_,
		_w279_,
		_w280_
	);
	LUT2 #(
		.INIT('h4)
	) name156 (
		_w245_,
		_w277_,
		_w281_
	);
	LUT2 #(
		.INIT('h8)
	) name157 (
		_w280_,
		_w281_,
		_w282_
	);
	LUT2 #(
		.INIT('h2)
	) name158 (
		\count_reg[3]/NET0131 ,
		_w282_,
		_w283_
	);
	LUT2 #(
		.INIT('h4)
	) name159 (
		_w165_,
		_w216_,
		_w284_
	);
	LUT2 #(
		.INIT('h1)
	) name160 (
		_w201_,
		_w204_,
		_w285_
	);
	LUT2 #(
		.INIT('h1)
	) name161 (
		_w263_,
		_w285_,
		_w286_
	);
	LUT2 #(
		.INIT('h2)
	) name162 (
		_w249_,
		_w284_,
		_w287_
	);
	LUT2 #(
		.INIT('h4)
	) name163 (
		_w286_,
		_w287_,
		_w288_
	);
	LUT2 #(
		.INIT('h1)
	) name164 (
		_w266_,
		_w288_,
		_w289_
	);
	LUT2 #(
		.INIT('h1)
	) name165 (
		_w231_,
		_w244_,
		_w290_
	);
	LUT2 #(
		.INIT('h2)
	) name166 (
		\timebase_reg[3]/NET0131 ,
		_w290_,
		_w291_
	);
	LUT2 #(
		.INIT('h1)
	) name167 (
		_w225_,
		_w241_,
		_w292_
	);
	LUT2 #(
		.INIT('h4)
	) name168 (
		_w224_,
		_w292_,
		_w293_
	);
	LUT2 #(
		.INIT('h2)
	) name169 (
		\count_reg[3]/NET0131 ,
		_w293_,
		_w294_
	);
	LUT2 #(
		.INIT('h8)
	) name170 (
		_w165_,
		_w201_,
		_w295_
	);
	LUT2 #(
		.INIT('h8)
	) name171 (
		_w146_,
		_w295_,
		_w296_
	);
	LUT2 #(
		.INIT('h8)
	) name172 (
		\timebase_reg[3]/NET0131 ,
		_w165_,
		_w297_
	);
	LUT2 #(
		.INIT('h1)
	) name173 (
		_w267_,
		_w297_,
		_w298_
	);
	LUT2 #(
		.INIT('h8)
	) name174 (
		_w196_,
		_w240_,
		_w299_
	);
	LUT2 #(
		.INIT('h1)
	) name175 (
		_w298_,
		_w299_,
		_w300_
	);
	LUT2 #(
		.INIT('h4)
	) name176 (
		_w165_,
		_w203_,
		_w301_
	);
	LUT2 #(
		.INIT('h1)
	) name177 (
		\k[0]_pad ,
		\k[1]_pad ,
		_w302_
	);
	LUT2 #(
		.INIT('h1)
	) name178 (
		\k[2]_pad ,
		\k[3]_pad ,
		_w303_
	);
	LUT2 #(
		.INIT('h8)
	) name179 (
		_w302_,
		_w303_,
		_w304_
	);
	LUT2 #(
		.INIT('h1)
	) name180 (
		\timebase_reg[3]/NET0131 ,
		_w304_,
		_w305_
	);
	LUT2 #(
		.INIT('h8)
	) name181 (
		_w266_,
		_w304_,
		_w306_
	);
	LUT2 #(
		.INIT('h2)
	) name182 (
		_w301_,
		_w305_,
		_w307_
	);
	LUT2 #(
		.INIT('h4)
	) name183 (
		_w306_,
		_w307_,
		_w308_
	);
	LUT2 #(
		.INIT('h1)
	) name184 (
		_w291_,
		_w296_,
		_w309_
	);
	LUT2 #(
		.INIT('h4)
	) name185 (
		_w294_,
		_w309_,
		_w310_
	);
	LUT2 #(
		.INIT('h1)
	) name186 (
		_w300_,
		_w308_,
		_w311_
	);
	LUT2 #(
		.INIT('h8)
	) name187 (
		_w310_,
		_w311_,
		_w312_
	);
	LUT2 #(
		.INIT('h1)
	) name188 (
		_w283_,
		_w289_,
		_w313_
	);
	LUT2 #(
		.INIT('h8)
	) name189 (
		_w312_,
		_w313_,
		_w314_
	);
	LUT2 #(
		.INIT('h4)
	) name190 (
		_w276_,
		_w314_,
		_w315_
	);
	LUT2 #(
		.INIT('h2)
	) name191 (
		_w216_,
		_w268_,
		_w316_
	);
	LUT2 #(
		.INIT('h2)
	) name192 (
		_w146_,
		_w272_,
		_w317_
	);
	LUT2 #(
		.INIT('h8)
	) name193 (
		_w166_,
		_w317_,
		_w318_
	);
	LUT2 #(
		.INIT('h1)
	) name194 (
		_w179_,
		_w229_,
		_w319_
	);
	LUT2 #(
		.INIT('h1)
	) name195 (
		_w195_,
		_w203_,
		_w320_
	);
	LUT2 #(
		.INIT('h1)
	) name196 (
		_w165_,
		_w320_,
		_w321_
	);
	LUT2 #(
		.INIT('h1)
	) name197 (
		_w173_,
		_w191_,
		_w322_
	);
	LUT2 #(
		.INIT('h4)
	) name198 (
		_w200_,
		_w322_,
		_w323_
	);
	LUT2 #(
		.INIT('h8)
	) name199 (
		_w226_,
		_w246_,
		_w324_
	);
	LUT2 #(
		.INIT('h8)
	) name200 (
		_w319_,
		_w324_,
		_w325_
	);
	LUT2 #(
		.INIT('h4)
	) name201 (
		_w296_,
		_w323_,
		_w326_
	);
	LUT2 #(
		.INIT('h4)
	) name202 (
		_w321_,
		_w326_,
		_w327_
	);
	LUT2 #(
		.INIT('h4)
	) name203 (
		_w316_,
		_w325_,
		_w328_
	);
	LUT2 #(
		.INIT('h4)
	) name204 (
		_w318_,
		_w328_,
		_w329_
	);
	LUT2 #(
		.INIT('h8)
	) name205 (
		_w327_,
		_w329_,
		_w330_
	);
	LUT2 #(
		.INIT('h1)
	) name206 (
		\k[0]_pad ,
		\k[2]_pad ,
		_w331_
	);
	LUT2 #(
		.INIT('h1)
	) name207 (
		_w165_,
		_w331_,
		_w332_
	);
	LUT2 #(
		.INIT('h2)
	) name208 (
		\k[3]_pad ,
		_w165_,
		_w333_
	);
	LUT2 #(
		.INIT('h1)
	) name209 (
		\sound_reg[0]/NET0131 ,
		_w333_,
		_w334_
	);
	LUT2 #(
		.INIT('h1)
	) name210 (
		_w332_,
		_w334_,
		_w335_
	);
	LUT2 #(
		.INIT('h4)
	) name211 (
		\k[0]_pad ,
		\k[1]_pad ,
		_w336_
	);
	LUT2 #(
		.INIT('h4)
	) name212 (
		_w165_,
		_w336_,
		_w337_
	);
	LUT2 #(
		.INIT('h1)
	) name213 (
		_w335_,
		_w337_,
		_w338_
	);
	LUT2 #(
		.INIT('h2)
	) name214 (
		_w203_,
		_w338_,
		_w339_
	);
	LUT2 #(
		.INIT('h2)
	) name215 (
		\data_out_reg[0]/NET0131 ,
		_w290_,
		_w340_
	);
	LUT2 #(
		.INIT('h4)
	) name216 (
		_w152_,
		_w173_,
		_w341_
	);
	LUT2 #(
		.INIT('h8)
	) name217 (
		_w165_,
		_w341_,
		_w342_
	);
	LUT2 #(
		.INIT('h1)
	) name218 (
		_w296_,
		_w342_,
		_w343_
	);
	LUT2 #(
		.INIT('h1)
	) name219 (
		_w204_,
		_w237_,
		_w344_
	);
	LUT2 #(
		.INIT('h8)
	) name220 (
		_w279_,
		_w344_,
		_w345_
	);
	LUT2 #(
		.INIT('h4)
	) name221 (
		_w152_,
		_w236_,
		_w346_
	);
	LUT2 #(
		.INIT('h4)
	) name222 (
		_w165_,
		_w346_,
		_w347_
	);
	LUT2 #(
		.INIT('h1)
	) name223 (
		_w241_,
		_w347_,
		_w348_
	);
	LUT2 #(
		.INIT('h1)
	) name224 (
		_w177_,
		_w201_,
		_w349_
	);
	LUT2 #(
		.INIT('h4)
	) name225 (
		_w247_,
		_w349_,
		_w350_
	);
	LUT2 #(
		.INIT('h4)
	) name226 (
		_w181_,
		_w350_,
		_w351_
	);
	LUT2 #(
		.INIT('h8)
	) name227 (
		_w345_,
		_w348_,
		_w352_
	);
	LUT2 #(
		.INIT('h8)
	) name228 (
		_w351_,
		_w352_,
		_w353_
	);
	LUT2 #(
		.INIT('h2)
	) name229 (
		\sound_reg[0]/NET0131 ,
		_w353_,
		_w354_
	);
	LUT2 #(
		.INIT('h1)
	) name230 (
		_w189_,
		_w224_,
		_w355_
	);
	LUT2 #(
		.INIT('h1)
	) name231 (
		_w190_,
		_w194_,
		_w356_
	);
	LUT2 #(
		.INIT('h8)
	) name232 (
		_w355_,
		_w356_,
		_w357_
	);
	LUT2 #(
		.INIT('h8)
	) name233 (
		_w128_,
		_w145_,
		_w358_
	);
	LUT2 #(
		.INIT('h8)
	) name234 (
		_w270_,
		_w358_,
		_w359_
	);
	LUT2 #(
		.INIT('h8)
	) name235 (
		\max_reg[4]/NET0131 ,
		_w359_,
		_w360_
	);
	LUT2 #(
		.INIT('h2)
	) name236 (
		_w166_,
		_w360_,
		_w361_
	);
	LUT2 #(
		.INIT('h4)
	) name237 (
		_w182_,
		_w319_,
		_w362_
	);
	LUT2 #(
		.INIT('h1)
	) name238 (
		_w216_,
		_w220_,
		_w363_
	);
	LUT2 #(
		.INIT('h4)
	) name239 (
		_w341_,
		_w363_,
		_w364_
	);
	LUT2 #(
		.INIT('h8)
	) name240 (
		_w357_,
		_w364_,
		_w365_
	);
	LUT2 #(
		.INIT('h8)
	) name241 (
		_w362_,
		_w365_,
		_w366_
	);
	LUT2 #(
		.INIT('h4)
	) name242 (
		_w361_,
		_w366_,
		_w367_
	);
	LUT2 #(
		.INIT('h2)
	) name243 (
		\sound_reg[0]/NET0131 ,
		_w367_,
		_w368_
	);
	LUT2 #(
		.INIT('h4)
	) name244 (
		_w340_,
		_w343_,
		_w369_
	);
	LUT2 #(
		.INIT('h4)
	) name245 (
		_w339_,
		_w369_,
		_w370_
	);
	LUT2 #(
		.INIT('h4)
	) name246 (
		_w354_,
		_w370_,
		_w371_
	);
	LUT2 #(
		.INIT('h4)
	) name247 (
		_w368_,
		_w371_,
		_w372_
	);
	LUT2 #(
		.INIT('h8)
	) name248 (
		_w282_,
		_w293_,
		_w373_
	);
	LUT2 #(
		.INIT('h2)
	) name249 (
		\count_reg[4]/NET0131 ,
		_w373_,
		_w374_
	);
	LUT2 #(
		.INIT('h2)
	) name250 (
		\count_reg[4]/NET0131 ,
		_w265_,
		_w375_
	);
	LUT2 #(
		.INIT('h1)
	) name251 (
		_w164_,
		_w375_,
		_w376_
	);
	LUT2 #(
		.INIT('h1)
	) name252 (
		_w165_,
		_w376_,
		_w377_
	);
	LUT2 #(
		.INIT('h2)
	) name253 (
		_w165_,
		_w299_,
		_w378_
	);
	LUT2 #(
		.INIT('h8)
	) name254 (
		\timebase_reg[4]/NET0131 ,
		_w378_,
		_w379_
	);
	LUT2 #(
		.INIT('h1)
	) name255 (
		_w377_,
		_w379_,
		_w380_
	);
	LUT2 #(
		.INIT('h1)
	) name256 (
		_w201_,
		_w216_,
		_w381_
	);
	LUT2 #(
		.INIT('h1)
	) name257 (
		_w160_,
		_w341_,
		_w382_
	);
	LUT2 #(
		.INIT('h4)
	) name258 (
		_w237_,
		_w381_,
		_w383_
	);
	LUT2 #(
		.INIT('h8)
	) name259 (
		_w382_,
		_w383_,
		_w384_
	);
	LUT2 #(
		.INIT('h4)
	) name260 (
		_w204_,
		_w384_,
		_w385_
	);
	LUT2 #(
		.INIT('h1)
	) name261 (
		_w247_,
		_w346_,
		_w386_
	);
	LUT2 #(
		.INIT('h8)
	) name262 (
		_w240_,
		_w386_,
		_w387_
	);
	LUT2 #(
		.INIT('h8)
	) name263 (
		_w196_,
		_w387_,
		_w388_
	);
	LUT2 #(
		.INIT('h8)
	) name264 (
		_w385_,
		_w388_,
		_w389_
	);
	LUT2 #(
		.INIT('h1)
	) name265 (
		_w380_,
		_w389_,
		_w390_
	);
	LUT2 #(
		.INIT('h8)
	) name266 (
		_w301_,
		_w304_,
		_w391_
	);
	LUT2 #(
		.INIT('h4)
	) name267 (
		_w376_,
		_w391_,
		_w392_
	);
	LUT2 #(
		.INIT('h2)
	) name268 (
		_w301_,
		_w304_,
		_w393_
	);
	LUT2 #(
		.INIT('h2)
	) name269 (
		_w290_,
		_w393_,
		_w394_
	);
	LUT2 #(
		.INIT('h2)
	) name270 (
		\timebase_reg[4]/NET0131 ,
		_w394_,
		_w395_
	);
	LUT2 #(
		.INIT('h1)
	) name271 (
		_w392_,
		_w395_,
		_w396_
	);
	LUT2 #(
		.INIT('h4)
	) name272 (
		_w374_,
		_w396_,
		_w397_
	);
	LUT2 #(
		.INIT('h4)
	) name273 (
		_w390_,
		_w397_,
		_w398_
	);
	LUT2 #(
		.INIT('h1)
	) name274 (
		_w164_,
		_w386_,
		_w399_
	);
	LUT2 #(
		.INIT('h4)
	) name275 (
		_w220_,
		_w277_,
		_w400_
	);
	LUT2 #(
		.INIT('h8)
	) name276 (
		_w280_,
		_w400_,
		_w401_
	);
	LUT2 #(
		.INIT('h8)
	) name277 (
		_w293_,
		_w401_,
		_w402_
	);
	LUT2 #(
		.INIT('h4)
	) name278 (
		_w399_,
		_w402_,
		_w403_
	);
	LUT2 #(
		.INIT('h2)
	) name279 (
		\count_reg[5]/NET0131 ,
		_w403_,
		_w404_
	);
	LUT2 #(
		.INIT('h2)
	) name280 (
		\count_reg[5]/NET0131 ,
		_w164_,
		_w405_
	);
	LUT2 #(
		.INIT('h2)
	) name281 (
		_w385_,
		_w391_,
		_w406_
	);
	LUT2 #(
		.INIT('h2)
	) name282 (
		_w405_,
		_w406_,
		_w407_
	);
	LUT2 #(
		.INIT('h4)
	) name283 (
		_w378_,
		_w394_,
		_w408_
	);
	LUT2 #(
		.INIT('h2)
	) name284 (
		\timebase_reg[5]/NET0131 ,
		_w408_,
		_w409_
	);
	LUT2 #(
		.INIT('h4)
	) name285 (
		_w299_,
		_w405_,
		_w410_
	);
	LUT2 #(
		.INIT('h1)
	) name286 (
		_w221_,
		_w410_,
		_w411_
	);
	LUT2 #(
		.INIT('h4)
	) name287 (
		_w409_,
		_w411_,
		_w412_
	);
	LUT2 #(
		.INIT('h4)
	) name288 (
		_w404_,
		_w412_,
		_w413_
	);
	LUT2 #(
		.INIT('h4)
	) name289 (
		_w407_,
		_w413_,
		_w414_
	);
	LUT2 #(
		.INIT('h1)
	) name290 (
		_w165_,
		_w388_,
		_w415_
	);
	LUT2 #(
		.INIT('h1)
	) name291 (
		_w224_,
		_w415_,
		_w416_
	);
	LUT2 #(
		.INIT('h2)
	) name292 (
		_w205_,
		_w341_,
		_w417_
	);
	LUT2 #(
		.INIT('h4)
	) name293 (
		_w165_,
		_w201_,
		_w418_
	);
	LUT2 #(
		.INIT('h1)
	) name294 (
		_w200_,
		_w418_,
		_w419_
	);
	LUT2 #(
		.INIT('h8)
	) name295 (
		_w292_,
		_w417_,
		_w420_
	);
	LUT2 #(
		.INIT('h8)
	) name296 (
		_w419_,
		_w420_,
		_w421_
	);
	LUT2 #(
		.INIT('h8)
	) name297 (
		_w416_,
		_w421_,
		_w422_
	);
	LUT2 #(
		.INIT('h2)
	) name298 (
		\nl_reg[1]/NET0131 ,
		_w422_,
		_w423_
	);
	LUT2 #(
		.INIT('h4)
	) name299 (
		_w160_,
		_w277_,
		_w424_
	);
	LUT2 #(
		.INIT('h4)
	) name300 (
		_w237_,
		_w424_,
		_w425_
	);
	LUT2 #(
		.INIT('h2)
	) name301 (
		\ind_reg[0]/NET0131 ,
		\ind_reg[1]/NET0131 ,
		_w426_
	);
	LUT2 #(
		.INIT('h4)
	) name302 (
		_w277_,
		_w426_,
		_w427_
	);
	LUT2 #(
		.INIT('h1)
	) name303 (
		\nl_reg[1]/NET0131 ,
		_w427_,
		_w428_
	);
	LUT2 #(
		.INIT('h1)
	) name304 (
		_w425_,
		_w428_,
		_w429_
	);
	LUT2 #(
		.INIT('h2)
	) name305 (
		\data_out_reg[0]/NET0131 ,
		\data_out_reg[1]/NET0131 ,
		_w430_
	);
	LUT2 #(
		.INIT('h8)
	) name306 (
		_w290_,
		_w343_,
		_w431_
	);
	LUT2 #(
		.INIT('h2)
	) name307 (
		_w430_,
		_w431_,
		_w432_
	);
	LUT2 #(
		.INIT('h1)
	) name308 (
		_w183_,
		_w230_,
		_w433_
	);
	LUT2 #(
		.INIT('h8)
	) name309 (
		_w363_,
		_w433_,
		_w434_
	);
	LUT2 #(
		.INIT('h2)
	) name310 (
		_w290_,
		_w295_,
		_w435_
	);
	LUT2 #(
		.INIT('h8)
	) name311 (
		_w434_,
		_w435_,
		_w436_
	);
	LUT2 #(
		.INIT('h2)
	) name312 (
		\nl_reg[1]/NET0131 ,
		_w436_,
		_w437_
	);
	LUT2 #(
		.INIT('h8)
	) name313 (
		_w165_,
		_w237_,
		_w438_
	);
	LUT2 #(
		.INIT('h1)
	) name314 (
		_w429_,
		_w438_,
		_w439_
	);
	LUT2 #(
		.INIT('h4)
	) name315 (
		_w437_,
		_w439_,
		_w440_
	);
	LUT2 #(
		.INIT('h4)
	) name316 (
		_w432_,
		_w440_,
		_w441_
	);
	LUT2 #(
		.INIT('h4)
	) name317 (
		_w423_,
		_w441_,
		_w442_
	);
	LUT2 #(
		.INIT('h8)
	) name318 (
		_w216_,
		_w268_,
		_w443_
	);
	LUT2 #(
		.INIT('h8)
	) name319 (
		_w157_,
		_w187_,
		_w444_
	);
	LUT2 #(
		.INIT('h2)
	) name320 (
		_w268_,
		_w272_,
		_w445_
	);
	LUT2 #(
		.INIT('h2)
	) name321 (
		_w160_,
		_w445_,
		_w446_
	);
	LUT2 #(
		.INIT('h1)
	) name322 (
		_w189_,
		_w444_,
		_w447_
	);
	LUT2 #(
		.INIT('h8)
	) name323 (
		_w277_,
		_w447_,
		_w448_
	);
	LUT2 #(
		.INIT('h4)
	) name324 (
		_w321_,
		_w448_,
		_w449_
	);
	LUT2 #(
		.INIT('h4)
	) name325 (
		_w443_,
		_w449_,
		_w450_
	);
	LUT2 #(
		.INIT('h4)
	) name326 (
		_w446_,
		_w450_,
		_w451_
	);
	LUT2 #(
		.INIT('h1)
	) name327 (
		_w165_,
		_w303_,
		_w452_
	);
	LUT2 #(
		.INIT('h1)
	) name328 (
		_w165_,
		_w302_,
		_w453_
	);
	LUT2 #(
		.INIT('h2)
	) name329 (
		_w203_,
		_w453_,
		_w454_
	);
	LUT2 #(
		.INIT('h4)
	) name330 (
		_w452_,
		_w454_,
		_w455_
	);
	LUT2 #(
		.INIT('h4)
	) name331 (
		_w221_,
		_w345_,
		_w456_
	);
	LUT2 #(
		.INIT('h2)
	) name332 (
		_w242_,
		_w341_,
		_w457_
	);
	LUT2 #(
		.INIT('h4)
	) name333 (
		_w160_,
		_w386_,
		_w458_
	);
	LUT2 #(
		.INIT('h8)
	) name334 (
		_w357_,
		_w458_,
		_w459_
	);
	LUT2 #(
		.INIT('h8)
	) name335 (
		_w457_,
		_w459_,
		_w460_
	);
	LUT2 #(
		.INIT('h4)
	) name336 (
		_w455_,
		_w456_,
		_w461_
	);
	LUT2 #(
		.INIT('h8)
	) name337 (
		_w460_,
		_w461_,
		_w462_
	);
	LUT2 #(
		.INIT('h2)
	) name338 (
		\sound_reg[2]/NET0131 ,
		_w462_,
		_w463_
	);
	LUT2 #(
		.INIT('h8)
	) name339 (
		_w166_,
		_w360_,
		_w464_
	);
	LUT2 #(
		.INIT('h8)
	) name340 (
		_w165_,
		_w250_,
		_w465_
	);
	LUT2 #(
		.INIT('h1)
	) name341 (
		\sound_reg[2]/NET0131 ,
		_w296_,
		_w466_
	);
	LUT2 #(
		.INIT('h4)
	) name342 (
		_w245_,
		_w362_,
		_w467_
	);
	LUT2 #(
		.INIT('h8)
	) name343 (
		_w381_,
		_w467_,
		_w468_
	);
	LUT2 #(
		.INIT('h1)
	) name344 (
		_w466_,
		_w468_,
		_w469_
	);
	LUT2 #(
		.INIT('h1)
	) name345 (
		_w464_,
		_w465_,
		_w470_
	);
	LUT2 #(
		.INIT('h4)
	) name346 (
		_w469_,
		_w470_,
		_w471_
	);
	LUT2 #(
		.INIT('h4)
	) name347 (
		_w463_,
		_w471_,
		_w472_
	);
	LUT2 #(
		.INIT('h2)
	) name348 (
		_w202_,
		_w241_,
		_w473_
	);
	LUT2 #(
		.INIT('h8)
	) name349 (
		_w344_,
		_w473_,
		_w474_
	);
	LUT2 #(
		.INIT('h4)
	) name350 (
		\gamma_reg[4]/NET0131 ,
		_w155_,
		_w475_
	);
	LUT2 #(
		.INIT('h1)
	) name351 (
		_w190_,
		_w475_,
		_w476_
	);
	LUT2 #(
		.INIT('h4)
	) name352 (
		_w198_,
		_w476_,
		_w477_
	);
	LUT2 #(
		.INIT('h8)
	) name353 (
		_w180_,
		_w477_,
		_w478_
	);
	LUT2 #(
		.INIT('h8)
	) name354 (
		_w363_,
		_w478_,
		_w479_
	);
	LUT2 #(
		.INIT('h8)
	) name355 (
		_w251_,
		_w479_,
		_w480_
	);
	LUT2 #(
		.INIT('h4)
	) name356 (
		_w182_,
		_w474_,
		_w481_
	);
	LUT2 #(
		.INIT('h8)
	) name357 (
		_w480_,
		_w481_,
		_w482_
	);
	LUT2 #(
		.INIT('h2)
	) name358 (
		nloss_pad,
		_w482_,
		_w483_
	);
	LUT2 #(
		.INIT('h2)
	) name359 (
		\k[1]_pad ,
		_w430_,
		_w484_
	);
	LUT2 #(
		.INIT('h4)
	) name360 (
		\data_out_reg[0]/NET0131 ,
		\data_out_reg[1]/NET0131 ,
		_w485_
	);
	LUT2 #(
		.INIT('h8)
	) name361 (
		\k[2]_pad ,
		_w485_,
		_w486_
	);
	LUT2 #(
		.INIT('h8)
	) name362 (
		\data_out_reg[0]/NET0131 ,
		\data_out_reg[1]/NET0131 ,
		_w487_
	);
	LUT2 #(
		.INIT('h4)
	) name363 (
		\k[2]_pad ,
		_w487_,
		_w488_
	);
	LUT2 #(
		.INIT('h1)
	) name364 (
		\k[1]_pad ,
		_w303_,
		_w489_
	);
	LUT2 #(
		.INIT('h4)
	) name365 (
		_w486_,
		_w489_,
		_w490_
	);
	LUT2 #(
		.INIT('h4)
	) name366 (
		_w488_,
		_w490_,
		_w491_
	);
	LUT2 #(
		.INIT('h1)
	) name367 (
		_w484_,
		_w491_,
		_w492_
	);
	LUT2 #(
		.INIT('h1)
	) name368 (
		\k[0]_pad ,
		_w492_,
		_w493_
	);
	LUT2 #(
		.INIT('h1)
	) name369 (
		\data_out_reg[0]/NET0131 ,
		\data_out_reg[1]/NET0131 ,
		_w494_
	);
	LUT2 #(
		.INIT('h2)
	) name370 (
		\k[0]_pad ,
		_w494_,
		_w495_
	);
	LUT2 #(
		.INIT('h1)
	) name371 (
		_w493_,
		_w495_,
		_w496_
	);
	LUT2 #(
		.INIT('h1)
	) name372 (
		nloss_pad,
		_w165_,
		_w497_
	);
	LUT2 #(
		.INIT('h8)
	) name373 (
		_w496_,
		_w497_,
		_w498_
	);
	LUT2 #(
		.INIT('h2)
	) name374 (
		_w203_,
		_w498_,
		_w499_
	);
	LUT2 #(
		.INIT('h1)
	) name375 (
		_w483_,
		_w499_,
		_w500_
	);
	LUT2 #(
		.INIT('h8)
	) name376 (
		\k[3]_pad ,
		_w488_,
		_w501_
	);
	LUT2 #(
		.INIT('h1)
	) name377 (
		_w486_,
		_w501_,
		_w502_
	);
	LUT2 #(
		.INIT('h2)
	) name378 (
		_w302_,
		_w502_,
		_w503_
	);
	LUT2 #(
		.INIT('h1)
	) name379 (
		\k[0]_pad ,
		_w430_,
		_w504_
	);
	LUT2 #(
		.INIT('h1)
	) name380 (
		_w302_,
		_w495_,
		_w505_
	);
	LUT2 #(
		.INIT('h4)
	) name381 (
		_w504_,
		_w505_,
		_w506_
	);
	LUT2 #(
		.INIT('h1)
	) name382 (
		_w503_,
		_w506_,
		_w507_
	);
	LUT2 #(
		.INIT('h2)
	) name383 (
		_w203_,
		_w507_,
		_w508_
	);
	LUT2 #(
		.INIT('h4)
	) name384 (
		_w203_,
		_w240_,
		_w509_
	);
	LUT2 #(
		.INIT('h8)
	) name385 (
		_w248_,
		_w344_,
		_w510_
	);
	LUT2 #(
		.INIT('h8)
	) name386 (
		_w509_,
		_w510_,
		_w511_
	);
	LUT2 #(
		.INIT('h2)
	) name387 (
		_w165_,
		_w511_,
		_w512_
	);
	LUT2 #(
		.INIT('h4)
	) name388 (
		_w165_,
		_w195_,
		_w513_
	);
	LUT2 #(
		.INIT('h1)
	) name389 (
		_w165_,
		_w382_,
		_w514_
	);
	LUT2 #(
		.INIT('h2)
	) name390 (
		_w201_,
		_w268_,
		_w515_
	);
	LUT2 #(
		.INIT('h1)
	) name391 (
		_w191_,
		_w221_,
		_w516_
	);
	LUT2 #(
		.INIT('h4)
	) name392 (
		_w225_,
		_w516_,
		_w517_
	);
	LUT2 #(
		.INIT('h2)
	) name393 (
		_w279_,
		_w347_,
		_w518_
	);
	LUT2 #(
		.INIT('h4)
	) name394 (
		_w513_,
		_w518_,
		_w519_
	);
	LUT2 #(
		.INIT('h4)
	) name395 (
		_w514_,
		_w517_,
		_w520_
	);
	LUT2 #(
		.INIT('h8)
	) name396 (
		_w519_,
		_w520_,
		_w521_
	);
	LUT2 #(
		.INIT('h1)
	) name397 (
		_w316_,
		_w508_,
		_w522_
	);
	LUT2 #(
		.INIT('h4)
	) name398 (
		_w515_,
		_w522_,
		_w523_
	);
	LUT2 #(
		.INIT('h4)
	) name399 (
		_w512_,
		_w521_,
		_w524_
	);
	LUT2 #(
		.INIT('h8)
	) name400 (
		_w523_,
		_w524_,
		_w525_
	);
	LUT2 #(
		.INIT('h1)
	) name401 (
		_w194_,
		_w231_,
		_w526_
	);
	LUT2 #(
		.INIT('h2)
	) name402 (
		_w301_,
		_w496_,
		_w527_
	);
	LUT2 #(
		.INIT('h2)
	) name403 (
		_w201_,
		_w213_,
		_w528_
	);
	LUT2 #(
		.INIT('h2)
	) name404 (
		_w192_,
		_w284_,
		_w529_
	);
	LUT2 #(
		.INIT('h4)
	) name405 (
		_w513_,
		_w526_,
		_w530_
	);
	LUT2 #(
		.INIT('h8)
	) name406 (
		_w529_,
		_w530_,
		_w531_
	);
	LUT2 #(
		.INIT('h8)
	) name407 (
		_w186_,
		_w531_,
		_w532_
	);
	LUT2 #(
		.INIT('h4)
	) name408 (
		_w528_,
		_w532_,
		_w533_
	);
	LUT2 #(
		.INIT('h4)
	) name409 (
		_w527_,
		_w533_,
		_w534_
	);
	LUT2 #(
		.INIT('h2)
	) name410 (
		_w290_,
		_w415_,
		_w535_
	);
	LUT2 #(
		.INIT('h2)
	) name411 (
		\nl[0]_pad ,
		_w535_,
		_w536_
	);
	LUT2 #(
		.INIT('h4)
	) name412 (
		_w237_,
		_w434_,
		_w537_
	);
	LUT2 #(
		.INIT('h8)
	) name413 (
		_w202_,
		_w292_,
		_w538_
	);
	LUT2 #(
		.INIT('h8)
	) name414 (
		_w537_,
		_w538_,
		_w539_
	);
	LUT2 #(
		.INIT('h8)
	) name415 (
		_w417_,
		_w539_,
		_w540_
	);
	LUT2 #(
		.INIT('h2)
	) name416 (
		\nl[0]_pad ,
		_w540_,
		_w541_
	);
	LUT2 #(
		.INIT('h4)
	) name417 (
		_w431_,
		_w494_,
		_w542_
	);
	LUT2 #(
		.INIT('h1)
	) name418 (
		\ind_reg[0]/NET0131 ,
		\ind_reg[1]/NET0131 ,
		_w543_
	);
	LUT2 #(
		.INIT('h4)
	) name419 (
		_w277_,
		_w543_,
		_w544_
	);
	LUT2 #(
		.INIT('h1)
	) name420 (
		\nl[0]_pad ,
		_w544_,
		_w545_
	);
	LUT2 #(
		.INIT('h4)
	) name421 (
		_w224_,
		_w424_,
		_w546_
	);
	LUT2 #(
		.INIT('h1)
	) name422 (
		_w545_,
		_w546_,
		_w547_
	);
	LUT2 #(
		.INIT('h1)
	) name423 (
		_w438_,
		_w547_,
		_w548_
	);
	LUT2 #(
		.INIT('h4)
	) name424 (
		_w542_,
		_w548_,
		_w549_
	);
	LUT2 #(
		.INIT('h4)
	) name425 (
		_w536_,
		_w549_,
		_w550_
	);
	LUT2 #(
		.INIT('h4)
	) name426 (
		_w541_,
		_w550_,
		_w551_
	);
	LUT2 #(
		.INIT('h8)
	) name427 (
		_w146_,
		_w485_,
		_w552_
	);
	LUT2 #(
		.INIT('h1)
	) name428 (
		\nl[2]_pad ,
		_w552_,
		_w553_
	);
	LUT2 #(
		.INIT('h2)
	) name429 (
		_w295_,
		_w553_,
		_w554_
	);
	LUT2 #(
		.INIT('h4)
	) name430 (
		\ind_reg[0]/NET0131 ,
		\ind_reg[1]/NET0131 ,
		_w555_
	);
	LUT2 #(
		.INIT('h1)
	) name431 (
		\nl[2]_pad ,
		_w555_,
		_w556_
	);
	LUT2 #(
		.INIT('h1)
	) name432 (
		_w277_,
		_w556_,
		_w557_
	);
	LUT2 #(
		.INIT('h1)
	) name433 (
		\nl[2]_pad ,
		_w485_,
		_w558_
	);
	LUT2 #(
		.INIT('h1)
	) name434 (
		\nl[2]_pad ,
		_w165_,
		_w559_
	);
	LUT2 #(
		.INIT('h2)
	) name435 (
		_w341_,
		_w559_,
		_w560_
	);
	LUT2 #(
		.INIT('h2)
	) name436 (
		_w290_,
		_w560_,
		_w561_
	);
	LUT2 #(
		.INIT('h1)
	) name437 (
		_w558_,
		_w561_,
		_w562_
	);
	LUT2 #(
		.INIT('h4)
	) name438 (
		_w160_,
		_w205_,
		_w563_
	);
	LUT2 #(
		.INIT('h8)
	) name439 (
		_w293_,
		_w563_,
		_w564_
	);
	LUT2 #(
		.INIT('h8)
	) name440 (
		_w419_,
		_w564_,
		_w565_
	);
	LUT2 #(
		.INIT('h8)
	) name441 (
		_w537_,
		_w565_,
		_w566_
	);
	LUT2 #(
		.INIT('h4)
	) name442 (
		_w415_,
		_w566_,
		_w567_
	);
	LUT2 #(
		.INIT('h2)
	) name443 (
		\nl[2]_pad ,
		_w567_,
		_w568_
	);
	LUT2 #(
		.INIT('h1)
	) name444 (
		_w438_,
		_w557_,
		_w569_
	);
	LUT2 #(
		.INIT('h4)
	) name445 (
		_w554_,
		_w569_,
		_w570_
	);
	LUT2 #(
		.INIT('h4)
	) name446 (
		_w562_,
		_w570_,
		_w571_
	);
	LUT2 #(
		.INIT('h4)
	) name447 (
		_w568_,
		_w571_,
		_w572_
	);
	LUT2 #(
		.INIT('h8)
	) name448 (
		_w416_,
		_w539_,
		_w573_
	);
	LUT2 #(
		.INIT('h2)
	) name449 (
		\nl[3]_pad ,
		_w573_,
		_w574_
	);
	LUT2 #(
		.INIT('h2)
	) name450 (
		\nl[3]_pad ,
		_w290_,
		_w575_
	);
	LUT2 #(
		.INIT('h1)
	) name451 (
		_w487_,
		_w575_,
		_w576_
	);
	LUT2 #(
		.INIT('h1)
	) name452 (
		_w431_,
		_w576_,
		_w577_
	);
	LUT2 #(
		.INIT('h8)
	) name453 (
		_w417_,
		_w424_,
		_w578_
	);
	LUT2 #(
		.INIT('h8)
	) name454 (
		\ind_reg[0]/NET0131 ,
		\ind_reg[1]/NET0131 ,
		_w579_
	);
	LUT2 #(
		.INIT('h4)
	) name455 (
		_w277_,
		_w579_,
		_w580_
	);
	LUT2 #(
		.INIT('h1)
	) name456 (
		\nl[3]_pad ,
		_w580_,
		_w581_
	);
	LUT2 #(
		.INIT('h1)
	) name457 (
		_w578_,
		_w581_,
		_w582_
	);
	LUT2 #(
		.INIT('h1)
	) name458 (
		_w438_,
		_w582_,
		_w583_
	);
	LUT2 #(
		.INIT('h4)
	) name459 (
		_w577_,
		_w583_,
		_w584_
	);
	LUT2 #(
		.INIT('h4)
	) name460 (
		_w574_,
		_w584_,
		_w585_
	);
	LUT2 #(
		.INIT('h1)
	) name461 (
		_w173_,
		_w195_,
		_w586_
	);
	LUT2 #(
		.INIT('h8)
	) name462 (
		_w180_,
		_w586_,
		_w587_
	);
	LUT2 #(
		.INIT('h8)
	) name463 (
		_w293_,
		_w587_,
		_w588_
	);
	LUT2 #(
		.INIT('h4)
	) name464 (
		_w165_,
		_w204_,
		_w589_
	);
	LUT2 #(
		.INIT('h1)
	) name465 (
		_w183_,
		_w236_,
		_w590_
	);
	LUT2 #(
		.INIT('h4)
	) name466 (
		_w244_,
		_w590_,
		_w591_
	);
	LUT2 #(
		.INIT('h4)
	) name467 (
		_w181_,
		_w192_,
		_w592_
	);
	LUT2 #(
		.INIT('h2)
	) name468 (
		_w279_,
		_w301_,
		_w593_
	);
	LUT2 #(
		.INIT('h2)
	) name469 (
		_w363_,
		_w418_,
		_w594_
	);
	LUT2 #(
		.INIT('h2)
	) name470 (
		_w526_,
		_w589_,
		_w595_
	);
	LUT2 #(
		.INIT('h8)
	) name471 (
		_w594_,
		_w595_,
		_w596_
	);
	LUT2 #(
		.INIT('h8)
	) name472 (
		_w592_,
		_w593_,
		_w597_
	);
	LUT2 #(
		.INIT('h8)
	) name473 (
		_w591_,
		_w597_,
		_w598_
	);
	LUT2 #(
		.INIT('h8)
	) name474 (
		_w588_,
		_w596_,
		_w599_
	);
	LUT2 #(
		.INIT('h8)
	) name475 (
		_w598_,
		_w599_,
		_w600_
	);
	LUT2 #(
		.INIT('h2)
	) name476 (
		\max_reg[4]/NET0131 ,
		_w600_,
		_w601_
	);
	LUT2 #(
		.INIT('h1)
	) name477 (
		\max_reg[4]/NET0131 ,
		_w359_,
		_w602_
	);
	LUT2 #(
		.INIT('h2)
	) name478 (
		_w166_,
		_w602_,
		_w603_
	);
	LUT2 #(
		.INIT('h8)
	) name479 (
		\scan_reg[4]/NET0131 ,
		_w146_,
		_w604_
	);
	LUT2 #(
		.INIT('h1)
	) name480 (
		\max_reg[4]/NET0131 ,
		_w271_,
		_w605_
	);
	LUT2 #(
		.INIT('h1)
	) name481 (
		_w272_,
		_w605_,
		_w606_
	);
	LUT2 #(
		.INIT('h4)
	) name482 (
		_w146_,
		_w606_,
		_w607_
	);
	LUT2 #(
		.INIT('h1)
	) name483 (
		_w604_,
		_w607_,
		_w608_
	);
	LUT2 #(
		.INIT('h2)
	) name484 (
		_w295_,
		_w608_,
		_w609_
	);
	LUT2 #(
		.INIT('h1)
	) name485 (
		_w603_,
		_w609_,
		_w610_
	);
	LUT2 #(
		.INIT('h4)
	) name486 (
		_w601_,
		_w610_,
		_w611_
	);
	LUT2 #(
		.INIT('h8)
	) name487 (
		_w165_,
		_w360_,
		_w612_
	);
	LUT2 #(
		.INIT('h1)
	) name488 (
		\play_reg/NET0131 ,
		_w612_,
		_w613_
	);
	LUT2 #(
		.INIT('h2)
	) name489 (
		_w160_,
		_w613_,
		_w614_
	);
	LUT2 #(
		.INIT('h1)
	) name490 (
		_w165_,
		_w299_,
		_w615_
	);
	LUT2 #(
		.INIT('h2)
	) name491 (
		_w226_,
		_w615_,
		_w616_
	);
	LUT2 #(
		.INIT('h2)
	) name492 (
		\play_reg/NET0131 ,
		_w616_,
		_w617_
	);
	LUT2 #(
		.INIT('h1)
	) name493 (
		\play_reg/NET0131 ,
		_w296_,
		_w618_
	);
	LUT2 #(
		.INIT('h4)
	) name494 (
		_w232_,
		_w238_,
		_w619_
	);
	LUT2 #(
		.INIT('h8)
	) name495 (
		_w434_,
		_w619_,
		_w620_
	);
	LUT2 #(
		.INIT('h1)
	) name496 (
		_w618_,
		_w620_,
		_w621_
	);
	LUT2 #(
		.INIT('h2)
	) name497 (
		\play_reg/NET0131 ,
		_w165_,
		_w622_
	);
	LUT2 #(
		.INIT('h8)
	) name498 (
		_w237_,
		_w622_,
		_w623_
	);
	LUT2 #(
		.INIT('h4)
	) name499 (
		_w165_,
		_w247_,
		_w624_
	);
	LUT2 #(
		.INIT('h1)
	) name500 (
		_w191_,
		_w346_,
		_w625_
	);
	LUT2 #(
		.INIT('h4)
	) name501 (
		_w624_,
		_w625_,
		_w626_
	);
	LUT2 #(
		.INIT('h8)
	) name502 (
		_w457_,
		_w626_,
		_w627_
	);
	LUT2 #(
		.INIT('h2)
	) name503 (
		\play_reg/NET0131 ,
		_w627_,
		_w628_
	);
	LUT2 #(
		.INIT('h1)
	) name504 (
		_w465_,
		_w623_,
		_w629_
	);
	LUT2 #(
		.INIT('h8)
	) name505 (
		_w394_,
		_w629_,
		_w630_
	);
	LUT2 #(
		.INIT('h4)
	) name506 (
		_w621_,
		_w630_,
		_w631_
	);
	LUT2 #(
		.INIT('h4)
	) name507 (
		_w628_,
		_w631_,
		_w632_
	);
	LUT2 #(
		.INIT('h4)
	) name508 (
		_w617_,
		_w632_,
		_w633_
	);
	LUT2 #(
		.INIT('h4)
	) name509 (
		_w614_,
		_w633_,
		_w634_
	);
	LUT2 #(
		.INIT('h8)
	) name510 (
		_w385_,
		_w387_,
		_w635_
	);
	LUT2 #(
		.INIT('h1)
	) name511 (
		\count_reg[0]1198/NET0131 ,
		_w165_,
		_w636_
	);
	LUT2 #(
		.INIT('h4)
	) name512 (
		_w635_,
		_w636_,
		_w637_
	);
	LUT2 #(
		.INIT('h2)
	) name513 (
		_w165_,
		_w240_,
		_w638_
	);
	LUT2 #(
		.INIT('h2)
	) name514 (
		_w290_,
		_w638_,
		_w639_
	);
	LUT2 #(
		.INIT('h2)
	) name515 (
		\timebase_reg[0]/NET0131 ,
		_w639_,
		_w640_
	);
	LUT2 #(
		.INIT('h2)
	) name516 (
		\count_reg[0]1198/NET0131 ,
		_w402_,
		_w641_
	);
	LUT2 #(
		.INIT('h1)
	) name517 (
		\timebase_reg[0]/NET0131 ,
		_w304_,
		_w642_
	);
	LUT2 #(
		.INIT('h8)
	) name518 (
		\count_reg[0]1198/NET0131 ,
		_w304_,
		_w643_
	);
	LUT2 #(
		.INIT('h1)
	) name519 (
		_w642_,
		_w643_,
		_w644_
	);
	LUT2 #(
		.INIT('h8)
	) name520 (
		_w301_,
		_w644_,
		_w645_
	);
	LUT2 #(
		.INIT('h8)
	) name521 (
		\timebase_reg[0]/NET0131 ,
		_w165_,
		_w646_
	);
	LUT2 #(
		.INIT('h1)
	) name522 (
		_w636_,
		_w646_,
		_w647_
	);
	LUT2 #(
		.INIT('h1)
	) name523 (
		_w196_,
		_w647_,
		_w648_
	);
	LUT2 #(
		.INIT('h1)
	) name524 (
		_w221_,
		_w645_,
		_w649_
	);
	LUT2 #(
		.INIT('h4)
	) name525 (
		_w648_,
		_w649_,
		_w650_
	);
	LUT2 #(
		.INIT('h4)
	) name526 (
		_w640_,
		_w650_,
		_w651_
	);
	LUT2 #(
		.INIT('h4)
	) name527 (
		_w641_,
		_w651_,
		_w652_
	);
	LUT2 #(
		.INIT('h4)
	) name528 (
		_w637_,
		_w652_,
		_w653_
	);
	LUT2 #(
		.INIT('h2)
	) name529 (
		\count_reg[2]/NET0131 ,
		_w373_,
		_w654_
	);
	LUT2 #(
		.INIT('h2)
	) name530 (
		\count_reg[2]/NET0131 ,
		_w161_,
		_w655_
	);
	LUT2 #(
		.INIT('h1)
	) name531 (
		_w162_,
		_w655_,
		_w656_
	);
	LUT2 #(
		.INIT('h1)
	) name532 (
		_w165_,
		_w656_,
		_w657_
	);
	LUT2 #(
		.INIT('h8)
	) name533 (
		\timebase_reg[2]/NET0131 ,
		_w378_,
		_w658_
	);
	LUT2 #(
		.INIT('h1)
	) name534 (
		_w657_,
		_w658_,
		_w659_
	);
	LUT2 #(
		.INIT('h8)
	) name535 (
		_w384_,
		_w388_,
		_w660_
	);
	LUT2 #(
		.INIT('h1)
	) name536 (
		_w659_,
		_w660_,
		_w661_
	);
	LUT2 #(
		.INIT('h2)
	) name537 (
		\timebase_reg[2]/NET0131 ,
		_w394_,
		_w662_
	);
	LUT2 #(
		.INIT('h1)
	) name538 (
		_w391_,
		_w589_,
		_w663_
	);
	LUT2 #(
		.INIT('h1)
	) name539 (
		_w656_,
		_w663_,
		_w664_
	);
	LUT2 #(
		.INIT('h1)
	) name540 (
		_w662_,
		_w664_,
		_w665_
	);
	LUT2 #(
		.INIT('h4)
	) name541 (
		_w654_,
		_w665_,
		_w666_
	);
	LUT2 #(
		.INIT('h4)
	) name542 (
		_w661_,
		_w666_,
		_w667_
	);
	LUT2 #(
		.INIT('h1)
	) name543 (
		\timebase_reg[0]/NET0131 ,
		\timebase_reg[1]/NET0131 ,
		_w668_
	);
	LUT2 #(
		.INIT('h4)
	) name544 (
		_w272_,
		_w668_,
		_w669_
	);
	LUT2 #(
		.INIT('h4)
	) name545 (
		\timebase_reg[2]/NET0131 ,
		_w669_,
		_w670_
	);
	LUT2 #(
		.INIT('h8)
	) name546 (
		_w268_,
		_w670_,
		_w671_
	);
	LUT2 #(
		.INIT('h4)
	) name547 (
		\timebase_reg[3]/NET0131 ,
		_w671_,
		_w672_
	);
	LUT2 #(
		.INIT('h4)
	) name548 (
		\timebase_reg[4]/NET0131 ,
		_w672_,
		_w673_
	);
	LUT2 #(
		.INIT('h1)
	) name549 (
		\timebase_reg[5]/NET0131 ,
		_w673_,
		_w674_
	);
	LUT2 #(
		.INIT('h4)
	) name550 (
		\timebase_reg[4]/NET0131 ,
		\timebase_reg[5]/NET0131 ,
		_w675_
	);
	LUT2 #(
		.INIT('h8)
	) name551 (
		_w672_,
		_w675_,
		_w676_
	);
	LUT2 #(
		.INIT('h2)
	) name552 (
		_w160_,
		_w676_,
		_w677_
	);
	LUT2 #(
		.INIT('h4)
	) name553 (
		_w674_,
		_w677_,
		_w678_
	);
	LUT2 #(
		.INIT('h4)
	) name554 (
		_w172_,
		_w193_,
		_w679_
	);
	LUT2 #(
		.INIT('h8)
	) name555 (
		_w239_,
		_w363_,
		_w680_
	);
	LUT2 #(
		.INIT('h2)
	) name556 (
		_w192_,
		_w679_,
		_w681_
	);
	LUT2 #(
		.INIT('h8)
	) name557 (
		_w433_,
		_w681_,
		_w682_
	);
	LUT2 #(
		.INIT('h8)
	) name558 (
		_w588_,
		_w682_,
		_w683_
	);
	LUT2 #(
		.INIT('h8)
	) name559 (
		_w680_,
		_w683_,
		_w684_
	);
	LUT2 #(
		.INIT('h2)
	) name560 (
		\timebase_reg[5]/NET0131 ,
		_w684_,
		_w685_
	);
	LUT2 #(
		.INIT('h2)
	) name561 (
		_w290_,
		_w346_,
		_w686_
	);
	LUT2 #(
		.INIT('h2)
	) name562 (
		\timebase_reg[5]/NET0131 ,
		_w686_,
		_w687_
	);
	LUT2 #(
		.INIT('h1)
	) name563 (
		_w229_,
		_w687_,
		_w688_
	);
	LUT2 #(
		.INIT('h4)
	) name564 (
		_w685_,
		_w688_,
		_w689_
	);
	LUT2 #(
		.INIT('h4)
	) name565 (
		_w678_,
		_w689_,
		_w690_
	);
	LUT2 #(
		.INIT('h2)
	) name566 (
		\max_reg[3]/NET0131 ,
		_w600_,
		_w691_
	);
	LUT2 #(
		.INIT('h2)
	) name567 (
		\max_reg[3]/NET0131 ,
		_w317_,
		_w692_
	);
	LUT2 #(
		.INIT('h1)
	) name568 (
		\max_reg[3]/NET0131 ,
		_w270_,
		_w693_
	);
	LUT2 #(
		.INIT('h1)
	) name569 (
		_w271_,
		_w693_,
		_w694_
	);
	LUT2 #(
		.INIT('h8)
	) name570 (
		_w146_,
		_w694_,
		_w695_
	);
	LUT2 #(
		.INIT('h1)
	) name571 (
		_w692_,
		_w695_,
		_w696_
	);
	LUT2 #(
		.INIT('h2)
	) name572 (
		_w166_,
		_w696_,
		_w697_
	);
	LUT2 #(
		.INIT('h4)
	) name573 (
		_w146_,
		_w694_,
		_w698_
	);
	LUT2 #(
		.INIT('h1)
	) name574 (
		_w358_,
		_w698_,
		_w699_
	);
	LUT2 #(
		.INIT('h2)
	) name575 (
		_w295_,
		_w699_,
		_w700_
	);
	LUT2 #(
		.INIT('h1)
	) name576 (
		_w697_,
		_w700_,
		_w701_
	);
	LUT2 #(
		.INIT('h4)
	) name577 (
		_w691_,
		_w701_,
		_w702_
	);
	LUT2 #(
		.INIT('h2)
	) name578 (
		\timebase_reg[3]/NET0131 ,
		_w671_,
		_w703_
	);
	LUT2 #(
		.INIT('h1)
	) name579 (
		_w672_,
		_w703_,
		_w704_
	);
	LUT2 #(
		.INIT('h2)
	) name580 (
		_w160_,
		_w704_,
		_w705_
	);
	LUT2 #(
		.INIT('h8)
	) name581 (
		_w684_,
		_w686_,
		_w706_
	);
	LUT2 #(
		.INIT('h2)
	) name582 (
		\timebase_reg[3]/NET0131 ,
		_w706_,
		_w707_
	);
	LUT2 #(
		.INIT('h1)
	) name583 (
		_w705_,
		_w707_,
		_w708_
	);
	LUT2 #(
		.INIT('h2)
	) name584 (
		\count_reg[1]1200/NET0131 ,
		_w373_,
		_w709_
	);
	LUT2 #(
		.INIT('h8)
	) name585 (
		\count_reg[0]1198/NET0131 ,
		\count_reg[1]1200/NET0131 ,
		_w710_
	);
	LUT2 #(
		.INIT('h1)
	) name586 (
		_w161_,
		_w710_,
		_w711_
	);
	LUT2 #(
		.INIT('h1)
	) name587 (
		_w165_,
		_w711_,
		_w712_
	);
	LUT2 #(
		.INIT('h8)
	) name588 (
		\timebase_reg[1]/NET0131 ,
		_w378_,
		_w713_
	);
	LUT2 #(
		.INIT('h1)
	) name589 (
		_w712_,
		_w713_,
		_w714_
	);
	LUT2 #(
		.INIT('h1)
	) name590 (
		_w389_,
		_w714_,
		_w715_
	);
	LUT2 #(
		.INIT('h2)
	) name591 (
		_w391_,
		_w711_,
		_w716_
	);
	LUT2 #(
		.INIT('h2)
	) name592 (
		\timebase_reg[1]/NET0131 ,
		_w394_,
		_w717_
	);
	LUT2 #(
		.INIT('h1)
	) name593 (
		_w716_,
		_w717_,
		_w718_
	);
	LUT2 #(
		.INIT('h4)
	) name594 (
		_w709_,
		_w718_,
		_w719_
	);
	LUT2 #(
		.INIT('h4)
	) name595 (
		_w715_,
		_w719_,
		_w720_
	);
	LUT2 #(
		.INIT('h2)
	) name596 (
		\scan_reg[3]/NET0131 ,
		_w165_,
		_w721_
	);
	LUT2 #(
		.INIT('h8)
	) name597 (
		\scan_reg[2]/NET0131 ,
		_w148_,
		_w722_
	);
	LUT2 #(
		.INIT('h8)
	) name598 (
		\scan_reg[3]/NET0131 ,
		_w722_,
		_w723_
	);
	LUT2 #(
		.INIT('h1)
	) name599 (
		\scan_reg[3]/NET0131 ,
		_w722_,
		_w724_
	);
	LUT2 #(
		.INIT('h1)
	) name600 (
		_w723_,
		_w724_,
		_w725_
	);
	LUT2 #(
		.INIT('h8)
	) name601 (
		_w213_,
		_w725_,
		_w726_
	);
	LUT2 #(
		.INIT('h1)
	) name602 (
		_w721_,
		_w726_,
		_w727_
	);
	LUT2 #(
		.INIT('h2)
	) name603 (
		_w216_,
		_w727_,
		_w728_
	);
	LUT2 #(
		.INIT('h2)
	) name604 (
		\scan_reg[3]/NET0131 ,
		_w210_,
		_w729_
	);
	LUT2 #(
		.INIT('h4)
	) name605 (
		_w146_,
		_w725_,
		_w730_
	);
	LUT2 #(
		.INIT('h1)
	) name606 (
		_w358_,
		_w730_,
		_w731_
	);
	LUT2 #(
		.INIT('h2)
	) name607 (
		_w166_,
		_w731_,
		_w732_
	);
	LUT2 #(
		.INIT('h1)
	) name608 (
		_w728_,
		_w732_,
		_w733_
	);
	LUT2 #(
		.INIT('h4)
	) name609 (
		_w729_,
		_w733_,
		_w734_
	);
	LUT2 #(
		.INIT('h2)
	) name610 (
		\scan_reg[4]/NET0131 ,
		_w165_,
		_w735_
	);
	LUT2 #(
		.INIT('h2)
	) name611 (
		\scan_reg[4]/NET0131 ,
		_w723_,
		_w736_
	);
	LUT2 #(
		.INIT('h4)
	) name612 (
		\scan_reg[4]/NET0131 ,
		_w723_,
		_w737_
	);
	LUT2 #(
		.INIT('h1)
	) name613 (
		_w736_,
		_w737_,
		_w738_
	);
	LUT2 #(
		.INIT('h2)
	) name614 (
		_w213_,
		_w738_,
		_w739_
	);
	LUT2 #(
		.INIT('h1)
	) name615 (
		_w735_,
		_w739_,
		_w740_
	);
	LUT2 #(
		.INIT('h2)
	) name616 (
		_w216_,
		_w740_,
		_w741_
	);
	LUT2 #(
		.INIT('h2)
	) name617 (
		\scan_reg[4]/NET0131 ,
		_w210_,
		_w742_
	);
	LUT2 #(
		.INIT('h1)
	) name618 (
		_w146_,
		_w738_,
		_w743_
	);
	LUT2 #(
		.INIT('h1)
	) name619 (
		_w604_,
		_w743_,
		_w744_
	);
	LUT2 #(
		.INIT('h2)
	) name620 (
		_w166_,
		_w744_,
		_w745_
	);
	LUT2 #(
		.INIT('h1)
	) name621 (
		_w741_,
		_w745_,
		_w746_
	);
	LUT2 #(
		.INIT('h4)
	) name622 (
		_w742_,
		_w746_,
		_w747_
	);
	LUT2 #(
		.INIT('h1)
	) name623 (
		\sound_reg[1]/NET0131 ,
		_w452_,
		_w748_
	);
	LUT2 #(
		.INIT('h2)
	) name624 (
		_w454_,
		_w748_,
		_w749_
	);
	LUT2 #(
		.INIT('h2)
	) name625 (
		\data_out_reg[1]/NET0131 ,
		_w290_,
		_w750_
	);
	LUT2 #(
		.INIT('h8)
	) name626 (
		_w248_,
		_w348_,
		_w751_
	);
	LUT2 #(
		.INIT('h4)
	) name627 (
		_w514_,
		_w751_,
		_w752_
	);
	LUT2 #(
		.INIT('h2)
	) name628 (
		\sound_reg[1]/NET0131 ,
		_w752_,
		_w753_
	);
	LUT2 #(
		.INIT('h4)
	) name629 (
		_w177_,
		_w355_,
		_w754_
	);
	LUT2 #(
		.INIT('h8)
	) name630 (
		_w467_,
		_w754_,
		_w755_
	);
	LUT2 #(
		.INIT('h4)
	) name631 (
		_w515_,
		_w755_,
		_w756_
	);
	LUT2 #(
		.INIT('h2)
	) name632 (
		\sound_reg[1]/NET0131 ,
		_w756_,
		_w757_
	);
	LUT2 #(
		.INIT('h8)
	) name633 (
		_w234_,
		_w456_,
		_w758_
	);
	LUT2 #(
		.INIT('h4)
	) name634 (
		_w361_,
		_w758_,
		_w759_
	);
	LUT2 #(
		.INIT('h2)
	) name635 (
		\sound_reg[1]/NET0131 ,
		_w759_,
		_w760_
	);
	LUT2 #(
		.INIT('h1)
	) name636 (
		_w749_,
		_w750_,
		_w761_
	);
	LUT2 #(
		.INIT('h4)
	) name637 (
		_w753_,
		_w761_,
		_w762_
	);
	LUT2 #(
		.INIT('h4)
	) name638 (
		_w757_,
		_w762_,
		_w763_
	);
	LUT2 #(
		.INIT('h4)
	) name639 (
		_w760_,
		_w763_,
		_w764_
	);
	LUT2 #(
		.INIT('h2)
	) name640 (
		\timebase_reg[1]/NET0131 ,
		_w706_,
		_w765_
	);
	LUT2 #(
		.INIT('h4)
	) name641 (
		\timebase_reg[0]/NET0131 ,
		_w445_,
		_w766_
	);
	LUT2 #(
		.INIT('h2)
	) name642 (
		\timebase_reg[1]/NET0131 ,
		_w766_,
		_w767_
	);
	LUT2 #(
		.INIT('h8)
	) name643 (
		_w268_,
		_w669_,
		_w768_
	);
	LUT2 #(
		.INIT('h1)
	) name644 (
		_w767_,
		_w768_,
		_w769_
	);
	LUT2 #(
		.INIT('h2)
	) name645 (
		_w160_,
		_w769_,
		_w770_
	);
	LUT2 #(
		.INIT('h1)
	) name646 (
		_w765_,
		_w770_,
		_w771_
	);
	LUT2 #(
		.INIT('h2)
	) name647 (
		\timebase_reg[2]/NET0131 ,
		_w768_,
		_w772_
	);
	LUT2 #(
		.INIT('h1)
	) name648 (
		_w671_,
		_w772_,
		_w773_
	);
	LUT2 #(
		.INIT('h2)
	) name649 (
		_w160_,
		_w773_,
		_w774_
	);
	LUT2 #(
		.INIT('h2)
	) name650 (
		\timebase_reg[2]/NET0131 ,
		_w706_,
		_w775_
	);
	LUT2 #(
		.INIT('h1)
	) name651 (
		_w774_,
		_w775_,
		_w776_
	);
	LUT2 #(
		.INIT('h2)
	) name652 (
		\timebase_reg[4]/NET0131 ,
		_w706_,
		_w777_
	);
	LUT2 #(
		.INIT('h2)
	) name653 (
		\timebase_reg[4]/NET0131 ,
		_w672_,
		_w778_
	);
	LUT2 #(
		.INIT('h1)
	) name654 (
		_w673_,
		_w778_,
		_w779_
	);
	LUT2 #(
		.INIT('h2)
	) name655 (
		_w160_,
		_w779_,
		_w780_
	);
	LUT2 #(
		.INIT('h1)
	) name656 (
		_w777_,
		_w780_,
		_w781_
	);
	LUT2 #(
		.INIT('h2)
	) name657 (
		\timebase_reg[0]/NET0131 ,
		_w445_,
		_w782_
	);
	LUT2 #(
		.INIT('h1)
	) name658 (
		_w766_,
		_w782_,
		_w783_
	);
	LUT2 #(
		.INIT('h2)
	) name659 (
		_w160_,
		_w783_,
		_w784_
	);
	LUT2 #(
		.INIT('h2)
	) name660 (
		\timebase_reg[0]/NET0131 ,
		_w684_,
		_w785_
	);
	LUT2 #(
		.INIT('h2)
	) name661 (
		\timebase_reg[0]/NET0131 ,
		_w686_,
		_w786_
	);
	LUT2 #(
		.INIT('h1)
	) name662 (
		_w229_,
		_w786_,
		_w787_
	);
	LUT2 #(
		.INIT('h4)
	) name663 (
		_w784_,
		_w787_,
		_w788_
	);
	LUT2 #(
		.INIT('h4)
	) name664 (
		_w785_,
		_w788_,
		_w789_
	);
	LUT2 #(
		.INIT('h2)
	) name665 (
		\max_reg[2]/NET0131 ,
		_w600_,
		_w790_
	);
	LUT2 #(
		.INIT('h1)
	) name666 (
		\max_reg[2]/NET0131 ,
		_w269_,
		_w791_
	);
	LUT2 #(
		.INIT('h1)
	) name667 (
		_w270_,
		_w791_,
		_w792_
	);
	LUT2 #(
		.INIT('h2)
	) name668 (
		_w317_,
		_w792_,
		_w793_
	);
	LUT2 #(
		.INIT('h1)
	) name669 (
		\max_reg[2]/NET0131 ,
		_w317_,
		_w794_
	);
	LUT2 #(
		.INIT('h2)
	) name670 (
		_w166_,
		_w793_,
		_w795_
	);
	LUT2 #(
		.INIT('h4)
	) name671 (
		_w794_,
		_w795_,
		_w796_
	);
	LUT2 #(
		.INIT('h1)
	) name672 (
		_w146_,
		_w792_,
		_w797_
	);
	LUT2 #(
		.INIT('h4)
	) name673 (
		\max_reg[2]/NET0131 ,
		_w146_,
		_w798_
	);
	LUT2 #(
		.INIT('h2)
	) name674 (
		_w295_,
		_w797_,
		_w799_
	);
	LUT2 #(
		.INIT('h4)
	) name675 (
		_w798_,
		_w799_,
		_w800_
	);
	LUT2 #(
		.INIT('h1)
	) name676 (
		_w796_,
		_w800_,
		_w801_
	);
	LUT2 #(
		.INIT('h4)
	) name677 (
		_w790_,
		_w801_,
		_w802_
	);
	LUT2 #(
		.INIT('h2)
	) name678 (
		\max_reg[0]/NET0131 ,
		_w600_,
		_w803_
	);
	LUT2 #(
		.INIT('h1)
	) name679 (
		\max_reg[0]/NET0131 ,
		_w146_,
		_w804_
	);
	LUT2 #(
		.INIT('h8)
	) name680 (
		\max_reg[0]/NET0131 ,
		_w146_,
		_w805_
	);
	LUT2 #(
		.INIT('h1)
	) name681 (
		_w804_,
		_w805_,
		_w806_
	);
	LUT2 #(
		.INIT('h1)
	) name682 (
		_w360_,
		_w806_,
		_w807_
	);
	LUT2 #(
		.INIT('h2)
	) name683 (
		_w166_,
		_w807_,
		_w808_
	);
	LUT2 #(
		.INIT('h2)
	) name684 (
		_w295_,
		_w806_,
		_w809_
	);
	LUT2 #(
		.INIT('h1)
	) name685 (
		_w808_,
		_w809_,
		_w810_
	);
	LUT2 #(
		.INIT('h4)
	) name686 (
		_w803_,
		_w810_,
		_w811_
	);
	LUT2 #(
		.INIT('h2)
	) name687 (
		\max_reg[1]/NET0131 ,
		_w600_,
		_w812_
	);
	LUT2 #(
		.INIT('h1)
	) name688 (
		\max_reg[0]/NET0131 ,
		\max_reg[1]/NET0131 ,
		_w813_
	);
	LUT2 #(
		.INIT('h1)
	) name689 (
		_w269_,
		_w813_,
		_w814_
	);
	LUT2 #(
		.INIT('h2)
	) name690 (
		_w317_,
		_w814_,
		_w815_
	);
	LUT2 #(
		.INIT('h1)
	) name691 (
		\max_reg[1]/NET0131 ,
		_w317_,
		_w816_
	);
	LUT2 #(
		.INIT('h2)
	) name692 (
		_w166_,
		_w815_,
		_w817_
	);
	LUT2 #(
		.INIT('h4)
	) name693 (
		_w816_,
		_w817_,
		_w818_
	);
	LUT2 #(
		.INIT('h1)
	) name694 (
		_w146_,
		_w814_,
		_w819_
	);
	LUT2 #(
		.INIT('h4)
	) name695 (
		\max_reg[1]/NET0131 ,
		_w146_,
		_w820_
	);
	LUT2 #(
		.INIT('h2)
	) name696 (
		_w295_,
		_w819_,
		_w821_
	);
	LUT2 #(
		.INIT('h4)
	) name697 (
		_w820_,
		_w821_,
		_w822_
	);
	LUT2 #(
		.INIT('h1)
	) name698 (
		_w818_,
		_w822_,
		_w823_
	);
	LUT2 #(
		.INIT('h4)
	) name699 (
		_w812_,
		_w823_,
		_w824_
	);
	LUT2 #(
		.INIT('h8)
	) name700 (
		_w146_,
		_w166_,
		_w825_
	);
	LUT2 #(
		.INIT('h1)
	) name701 (
		_w284_,
		_w825_,
		_w826_
	);
	LUT2 #(
		.INIT('h8)
	) name702 (
		_w210_,
		_w826_,
		_w827_
	);
	LUT2 #(
		.INIT('h2)
	) name703 (
		\scan_reg[0]/NET0131 ,
		_w827_,
		_w828_
	);
	LUT2 #(
		.INIT('h1)
	) name704 (
		_w160_,
		_w216_,
		_w829_
	);
	LUT2 #(
		.INIT('h1)
	) name705 (
		\scan_reg[0]/NET0131 ,
		_w829_,
		_w830_
	);
	LUT2 #(
		.INIT('h8)
	) name706 (
		_w213_,
		_w830_,
		_w831_
	);
	LUT2 #(
		.INIT('h1)
	) name707 (
		_w828_,
		_w831_,
		_w832_
	);
	LUT2 #(
		.INIT('h1)
	) name708 (
		\scan_reg[2]/NET0131 ,
		_w165_,
		_w833_
	);
	LUT2 #(
		.INIT('h1)
	) name709 (
		\scan_reg[2]/NET0131 ,
		_w148_,
		_w834_
	);
	LUT2 #(
		.INIT('h1)
	) name710 (
		_w722_,
		_w834_,
		_w835_
	);
	LUT2 #(
		.INIT('h4)
	) name711 (
		_w146_,
		_w835_,
		_w836_
	);
	LUT2 #(
		.INIT('h2)
	) name712 (
		_w165_,
		_w836_,
		_w837_
	);
	LUT2 #(
		.INIT('h2)
	) name713 (
		_w216_,
		_w833_,
		_w838_
	);
	LUT2 #(
		.INIT('h4)
	) name714 (
		_w837_,
		_w838_,
		_w839_
	);
	LUT2 #(
		.INIT('h2)
	) name715 (
		\scan_reg[2]/NET0131 ,
		_w210_,
		_w840_
	);
	LUT2 #(
		.INIT('h8)
	) name716 (
		\scan_reg[2]/NET0131 ,
		_w146_,
		_w841_
	);
	LUT2 #(
		.INIT('h1)
	) name717 (
		_w836_,
		_w841_,
		_w842_
	);
	LUT2 #(
		.INIT('h2)
	) name718 (
		_w166_,
		_w842_,
		_w843_
	);
	LUT2 #(
		.INIT('h1)
	) name719 (
		_w839_,
		_w843_,
		_w844_
	);
	LUT2 #(
		.INIT('h4)
	) name720 (
		_w840_,
		_w844_,
		_w845_
	);
	LUT2 #(
		.INIT('h2)
	) name721 (
		_w165_,
		_w320_,
		_w846_
	);
	LUT2 #(
		.INIT('h1)
	) name722 (
		_w171_,
		_w236_,
		_w847_
	);
	LUT2 #(
		.INIT('h4)
	) name723 (
		_w846_,
		_w847_,
		_w848_
	);
	LUT2 #(
		.INIT('h4)
	) name724 (
		_w464_,
		_w848_,
		_w849_
	);
	LUT2 #(
		.INIT('h4)
	) name725 (
		_w229_,
		_w482_,
		_w850_
	);
	LUT2 #(
		.INIT('h2)
	) name726 (
		\ind_reg[0]/NET0131 ,
		_w850_,
		_w851_
	);
	LUT2 #(
		.INIT('h8)
	) name727 (
		\ind_reg[0]/NET0131 ,
		_w165_,
		_w852_
	);
	LUT2 #(
		.INIT('h1)
	) name728 (
		\ind_reg[0]/NET0131 ,
		\k[3]_pad ,
		_w853_
	);
	LUT2 #(
		.INIT('h2)
	) name729 (
		_w331_,
		_w853_,
		_w854_
	);
	LUT2 #(
		.INIT('h4)
	) name730 (
		_w165_,
		_w854_,
		_w855_
	);
	LUT2 #(
		.INIT('h1)
	) name731 (
		_w337_,
		_w852_,
		_w856_
	);
	LUT2 #(
		.INIT('h4)
	) name732 (
		_w855_,
		_w856_,
		_w857_
	);
	LUT2 #(
		.INIT('h2)
	) name733 (
		_w203_,
		_w857_,
		_w858_
	);
	LUT2 #(
		.INIT('h1)
	) name734 (
		_w851_,
		_w858_,
		_w859_
	);
	LUT2 #(
		.INIT('h2)
	) name735 (
		\ind_reg[1]/NET0131 ,
		_w850_,
		_w860_
	);
	LUT2 #(
		.INIT('h1)
	) name736 (
		\ind_reg[1]/NET0131 ,
		_w452_,
		_w861_
	);
	LUT2 #(
		.INIT('h2)
	) name737 (
		_w454_,
		_w861_,
		_w862_
	);
	LUT2 #(
		.INIT('h1)
	) name738 (
		_w860_,
		_w862_,
		_w863_
	);
	LUT2 #(
		.INIT('h4)
	) name739 (
		\sound_reg[1]/NET0131 ,
		\sound_reg[2]/NET0131 ,
		_w864_
	);
	LUT2 #(
		.INIT('h8)
	) name740 (
		\sound_reg[0]/NET0131 ,
		_w864_,
		_w865_
	);
	LUT2 #(
		.INIT('h1)
	) name741 (
		\counter_reg[1]/NET0131 ,
		\counter_reg[2]/NET0131 ,
		_w866_
	);
	LUT2 #(
		.INIT('h1)
	) name742 (
		\s_reg/NET0131 ,
		_w866_,
		_w867_
	);
	LUT2 #(
		.INIT('h8)
	) name743 (
		speaker_pad,
		_w866_,
		_w868_
	);
	LUT2 #(
		.INIT('h1)
	) name744 (
		_w867_,
		_w868_,
		_w869_
	);
	LUT2 #(
		.INIT('h2)
	) name745 (
		_w865_,
		_w869_,
		_w870_
	);
	LUT2 #(
		.INIT('h8)
	) name746 (
		\counter_reg[1]/NET0131 ,
		\counter_reg[2]/NET0131 ,
		_w871_
	);
	LUT2 #(
		.INIT('h2)
	) name747 (
		speaker_pad,
		_w871_,
		_w872_
	);
	LUT2 #(
		.INIT('h4)
	) name748 (
		\s_reg/NET0131 ,
		_w871_,
		_w873_
	);
	LUT2 #(
		.INIT('h1)
	) name749 (
		_w872_,
		_w873_,
		_w874_
	);
	LUT2 #(
		.INIT('h2)
	) name750 (
		\sound_reg[1]/NET0131 ,
		\sound_reg[2]/NET0131 ,
		_w875_
	);
	LUT2 #(
		.INIT('h8)
	) name751 (
		\sound_reg[0]/NET0131 ,
		_w875_,
		_w876_
	);
	LUT2 #(
		.INIT('h4)
	) name752 (
		_w874_,
		_w876_,
		_w877_
	);
	LUT2 #(
		.INIT('h1)
	) name753 (
		\sound_reg[1]/NET0131 ,
		\sound_reg[2]/NET0131 ,
		_w878_
	);
	LUT2 #(
		.INIT('h8)
	) name754 (
		\sound_reg[0]/NET0131 ,
		_w878_,
		_w879_
	);
	LUT2 #(
		.INIT('h4)
	) name755 (
		\counter_reg[2]/NET0131 ,
		speaker_pad,
		_w880_
	);
	LUT2 #(
		.INIT('h2)
	) name756 (
		\counter_reg[2]/NET0131 ,
		\s_reg/NET0131 ,
		_w881_
	);
	LUT2 #(
		.INIT('h1)
	) name757 (
		_w880_,
		_w881_,
		_w882_
	);
	LUT2 #(
		.INIT('h2)
	) name758 (
		_w879_,
		_w882_,
		_w883_
	);
	LUT2 #(
		.INIT('h4)
	) name759 (
		\sound_reg[0]/NET0131 ,
		_w878_,
		_w884_
	);
	LUT2 #(
		.INIT('h8)
	) name760 (
		\counter_reg[0]/NET0131 ,
		\counter_reg[1]/NET0131 ,
		_w885_
	);
	LUT2 #(
		.INIT('h1)
	) name761 (
		\counter_reg[2]/NET0131 ,
		_w885_,
		_w886_
	);
	LUT2 #(
		.INIT('h2)
	) name762 (
		_w884_,
		_w886_,
		_w887_
	);
	LUT2 #(
		.INIT('h4)
	) name763 (
		\sound_reg[0]/NET0131 ,
		_w864_,
		_w888_
	);
	LUT2 #(
		.INIT('h8)
	) name764 (
		\counter_reg[2]/NET0131 ,
		_w885_,
		_w889_
	);
	LUT2 #(
		.INIT('h8)
	) name765 (
		_w888_,
		_w889_,
		_w890_
	);
	LUT2 #(
		.INIT('h1)
	) name766 (
		_w887_,
		_w890_,
		_w891_
	);
	LUT2 #(
		.INIT('h1)
	) name767 (
		\s_reg/NET0131 ,
		_w891_,
		_w892_
	);
	LUT2 #(
		.INIT('h1)
	) name768 (
		_w864_,
		_w875_,
		_w893_
	);
	LUT2 #(
		.INIT('h4)
	) name769 (
		_w878_,
		_w893_,
		_w894_
	);
	LUT2 #(
		.INIT('h8)
	) name770 (
		_w884_,
		_w886_,
		_w895_
	);
	LUT2 #(
		.INIT('h2)
	) name771 (
		_w888_,
		_w889_,
		_w896_
	);
	LUT2 #(
		.INIT('h1)
	) name772 (
		_w895_,
		_w896_,
		_w897_
	);
	LUT2 #(
		.INIT('h4)
	) name773 (
		_w894_,
		_w897_,
		_w898_
	);
	LUT2 #(
		.INIT('h2)
	) name774 (
		speaker_pad,
		_w898_,
		_w899_
	);
	LUT2 #(
		.INIT('h4)
	) name775 (
		\sound_reg[0]/NET0131 ,
		_w875_,
		_w900_
	);
	LUT2 #(
		.INIT('h1)
	) name776 (
		\counter_reg[0]/NET0131 ,
		\counter_reg[1]/NET0131 ,
		_w901_
	);
	LUT2 #(
		.INIT('h2)
	) name777 (
		\counter_reg[2]/NET0131 ,
		_w901_,
		_w902_
	);
	LUT2 #(
		.INIT('h2)
	) name778 (
		speaker_pad,
		_w902_,
		_w903_
	);
	LUT2 #(
		.INIT('h2)
	) name779 (
		_w881_,
		_w901_,
		_w904_
	);
	LUT2 #(
		.INIT('h1)
	) name780 (
		_w903_,
		_w904_,
		_w905_
	);
	LUT2 #(
		.INIT('h2)
	) name781 (
		_w900_,
		_w905_,
		_w906_
	);
	LUT2 #(
		.INIT('h1)
	) name782 (
		_w870_,
		_w883_,
		_w907_
	);
	LUT2 #(
		.INIT('h4)
	) name783 (
		_w877_,
		_w907_,
		_w908_
	);
	LUT2 #(
		.INIT('h1)
	) name784 (
		_w892_,
		_w906_,
		_w909_
	);
	LUT2 #(
		.INIT('h8)
	) name785 (
		_w908_,
		_w909_,
		_w910_
	);
	LUT2 #(
		.INIT('h4)
	) name786 (
		_w899_,
		_w910_,
		_w911_
	);
	LUT2 #(
		.INIT('h2)
	) name787 (
		\play_reg/NET0131 ,
		_w911_,
		_w912_
	);
	LUT2 #(
		.INIT('h4)
	) name788 (
		_w203_,
		_w474_,
		_w913_
	);
	LUT2 #(
		.INIT('h8)
	) name789 (
		_w480_,
		_w913_,
		_w914_
	);
	LUT2 #(
		.INIT('h2)
	) name790 (
		\wr_reg/NET0131 ,
		_w914_,
		_w915_
	);
	LUT2 #(
		.INIT('h1)
	) name791 (
		_w225_,
		_w915_,
		_w916_
	);
	LUT2 #(
		.INIT('h8)
	) name792 (
		_w865_,
		_w867_,
		_w917_
	);
	LUT2 #(
		.INIT('h4)
	) name793 (
		\counter_reg[2]/NET0131 ,
		\s_reg/NET0131 ,
		_w918_
	);
	LUT2 #(
		.INIT('h1)
	) name794 (
		_w881_,
		_w918_,
		_w919_
	);
	LUT2 #(
		.INIT('h2)
	) name795 (
		_w879_,
		_w919_,
		_w920_
	);
	LUT2 #(
		.INIT('h2)
	) name796 (
		\s_reg/NET0131 ,
		_w871_,
		_w921_
	);
	LUT2 #(
		.INIT('h1)
	) name797 (
		_w873_,
		_w921_,
		_w922_
	);
	LUT2 #(
		.INIT('h2)
	) name798 (
		_w876_,
		_w922_,
		_w923_
	);
	LUT2 #(
		.INIT('h2)
	) name799 (
		_w900_,
		_w902_,
		_w924_
	);
	LUT2 #(
		.INIT('h8)
	) name800 (
		_w865_,
		_w866_,
		_w925_
	);
	LUT2 #(
		.INIT('h1)
	) name801 (
		_w924_,
		_w925_,
		_w926_
	);
	LUT2 #(
		.INIT('h8)
	) name802 (
		_w897_,
		_w926_,
		_w927_
	);
	LUT2 #(
		.INIT('h2)
	) name803 (
		\s_reg/NET0131 ,
		_w894_,
		_w928_
	);
	LUT2 #(
		.INIT('h8)
	) name804 (
		_w927_,
		_w928_,
		_w929_
	);
	LUT2 #(
		.INIT('h8)
	) name805 (
		_w885_,
		_w888_,
		_w930_
	);
	LUT2 #(
		.INIT('h2)
	) name806 (
		_w900_,
		_w901_,
		_w931_
	);
	LUT2 #(
		.INIT('h1)
	) name807 (
		_w930_,
		_w931_,
		_w932_
	);
	LUT2 #(
		.INIT('h2)
	) name808 (
		\counter_reg[2]/NET0131 ,
		_w932_,
		_w933_
	);
	LUT2 #(
		.INIT('h1)
	) name809 (
		\s_reg/NET0131 ,
		_w887_,
		_w934_
	);
	LUT2 #(
		.INIT('h4)
	) name810 (
		_w933_,
		_w934_,
		_w935_
	);
	LUT2 #(
		.INIT('h1)
	) name811 (
		_w929_,
		_w935_,
		_w936_
	);
	LUT2 #(
		.INIT('h1)
	) name812 (
		_w917_,
		_w920_,
		_w937_
	);
	LUT2 #(
		.INIT('h4)
	) name813 (
		_w923_,
		_w937_,
		_w938_
	);
	LUT2 #(
		.INIT('h4)
	) name814 (
		_w936_,
		_w938_,
		_w939_
	);
	LUT2 #(
		.INIT('h8)
	) name815 (
		\count_reg[0]/NET0131 ,
		_w225_,
		_w940_
	);
	LUT2 #(
		.INIT('h8)
	) name816 (
		_w174_,
		_w233_,
		_w941_
	);
	LUT2 #(
		.INIT('h8)
	) name817 (
		_w278_,
		_w625_,
		_w942_
	);
	LUT2 #(
		.INIT('h8)
	) name818 (
		_w941_,
		_w942_,
		_w943_
	);
	LUT2 #(
		.INIT('h8)
	) name819 (
		_w199_,
		_w243_,
		_w944_
	);
	LUT2 #(
		.INIT('h8)
	) name820 (
		_w943_,
		_w944_,
		_w945_
	);
	LUT2 #(
		.INIT('h8)
	) name821 (
		_w680_,
		_w945_,
		_w946_
	);
	LUT2 #(
		.INIT('h2)
	) name822 (
		\data_in_reg[0]/NET0131 ,
		_w946_,
		_w947_
	);
	LUT2 #(
		.INIT('h1)
	) name823 (
		_w940_,
		_w947_,
		_w948_
	);
	LUT2 #(
		.INIT('h8)
	) name824 (
		\count_reg[1]/NET0131 ,
		_w225_,
		_w949_
	);
	LUT2 #(
		.INIT('h2)
	) name825 (
		\data_in_reg[1]/NET0131 ,
		_w946_,
		_w950_
	);
	LUT2 #(
		.INIT('h1)
	) name826 (
		_w949_,
		_w950_,
		_w951_
	);
	LUT2 #(
		.INIT('h2)
	) name827 (
		\scan_reg[2]/NET0131 ,
		_w222_,
		_w952_
	);
	LUT2 #(
		.INIT('h2)
	) name828 (
		\max_reg[2]/NET0131 ,
		_w226_,
		_w953_
	);
	LUT2 #(
		.INIT('h2)
	) name829 (
		\address_reg[2]/NET0131 ,
		_w259_,
		_w954_
	);
	LUT2 #(
		.INIT('h1)
	) name830 (
		_w952_,
		_w953_,
		_w955_
	);
	LUT2 #(
		.INIT('h4)
	) name831 (
		_w954_,
		_w955_,
		_w956_
	);
	LUT2 #(
		.INIT('h2)
	) name832 (
		\scan_reg[3]/NET0131 ,
		_w222_,
		_w957_
	);
	LUT2 #(
		.INIT('h2)
	) name833 (
		\max_reg[3]/NET0131 ,
		_w226_,
		_w958_
	);
	LUT2 #(
		.INIT('h2)
	) name834 (
		\address_reg[3]/NET0131 ,
		_w259_,
		_w959_
	);
	LUT2 #(
		.INIT('h1)
	) name835 (
		_w957_,
		_w958_,
		_w960_
	);
	LUT2 #(
		.INIT('h4)
	) name836 (
		_w959_,
		_w960_,
		_w961_
	);
	LUT2 #(
		.INIT('h2)
	) name837 (
		\scan_reg[4]/NET0131 ,
		_w222_,
		_w962_
	);
	LUT2 #(
		.INIT('h2)
	) name838 (
		\max_reg[4]/NET0131 ,
		_w226_,
		_w963_
	);
	LUT2 #(
		.INIT('h2)
	) name839 (
		\address_reg[4]/NET0131 ,
		_w259_,
		_w964_
	);
	LUT2 #(
		.INIT('h1)
	) name840 (
		_w962_,
		_w963_,
		_w965_
	);
	LUT2 #(
		.INIT('h4)
	) name841 (
		_w964_,
		_w965_,
		_w966_
	);
	LUT2 #(
		.INIT('h2)
	) name842 (
		\scan_reg[1]/NET0131 ,
		_w222_,
		_w967_
	);
	LUT2 #(
		.INIT('h2)
	) name843 (
		\max_reg[1]/NET0131 ,
		_w226_,
		_w968_
	);
	LUT2 #(
		.INIT('h2)
	) name844 (
		\address_reg[1]/NET0131 ,
		_w259_,
		_w969_
	);
	LUT2 #(
		.INIT('h1)
	) name845 (
		_w967_,
		_w968_,
		_w970_
	);
	LUT2 #(
		.INIT('h4)
	) name846 (
		_w969_,
		_w970_,
		_w971_
	);
	LUT2 #(
		.INIT('h4)
	) name847 (
		\counter_reg[2]/NET0131 ,
		_w879_,
		_w972_
	);
	LUT2 #(
		.INIT('h1)
	) name848 (
		_w876_,
		_w972_,
		_w973_
	);
	LUT2 #(
		.INIT('h1)
	) name849 (
		_w871_,
		_w973_,
		_w974_
	);
	LUT2 #(
		.INIT('h2)
	) name850 (
		_w927_,
		_w974_,
		_w975_
	);
	LUT2 #(
		.INIT('h2)
	) name851 (
		\play_reg/NET0131 ,
		_w975_,
		_w976_
	);
	LUT2 #(
		.INIT('h1)
	) name852 (
		_w886_,
		_w889_,
		_w977_
	);
	LUT2 #(
		.INIT('h8)
	) name853 (
		_w976_,
		_w977_,
		_w978_
	);
	LUT2 #(
		.INIT('h1)
	) name854 (
		_w885_,
		_w901_,
		_w979_
	);
	LUT2 #(
		.INIT('h8)
	) name855 (
		_w976_,
		_w979_,
		_w980_
	);
	LUT2 #(
		.INIT('h4)
	) name856 (
		\counter_reg[0]/NET0131 ,
		_w976_,
		_w981_
	);
	LUT2 #(
		.INIT('h2)
	) name857 (
		\address_reg[2]/NET0131 ,
		\address_reg[3]/NET0131 ,
		_w982_
	);
	LUT2 #(
		.INIT('h4)
	) name858 (
		\address_reg[1]/NET0131 ,
		\address_reg[4]/NET0131 ,
		_w983_
	);
	LUT2 #(
		.INIT('h8)
	) name859 (
		_w982_,
		_w983_,
		_w984_
	);
	LUT2 #(
		.INIT('h8)
	) name860 (
		\memory_reg[20][0]/NET0131 ,
		_w984_,
		_w985_
	);
	LUT2 #(
		.INIT('h4)
	) name861 (
		\address_reg[2]/NET0131 ,
		\address_reg[3]/NET0131 ,
		_w986_
	);
	LUT2 #(
		.INIT('h1)
	) name862 (
		\address_reg[1]/NET0131 ,
		\address_reg[4]/NET0131 ,
		_w987_
	);
	LUT2 #(
		.INIT('h8)
	) name863 (
		_w986_,
		_w987_,
		_w988_
	);
	LUT2 #(
		.INIT('h8)
	) name864 (
		\memory_reg[8][0]/NET0131 ,
		_w988_,
		_w989_
	);
	LUT2 #(
		.INIT('h2)
	) name865 (
		\address_reg[1]/NET0131 ,
		\address_reg[4]/NET0131 ,
		_w990_
	);
	LUT2 #(
		.INIT('h8)
	) name866 (
		_w982_,
		_w990_,
		_w991_
	);
	LUT2 #(
		.INIT('h8)
	) name867 (
		\memory_reg[6][0]/NET0131 ,
		_w991_,
		_w992_
	);
	LUT2 #(
		.INIT('h1)
	) name868 (
		\address_reg[2]/NET0131 ,
		\address_reg[3]/NET0131 ,
		_w993_
	);
	LUT2 #(
		.INIT('h8)
	) name869 (
		_w990_,
		_w993_,
		_w994_
	);
	LUT2 #(
		.INIT('h8)
	) name870 (
		\memory_reg[2][0]/NET0131 ,
		_w994_,
		_w995_
	);
	LUT2 #(
		.INIT('h8)
	) name871 (
		_w983_,
		_w986_,
		_w996_
	);
	LUT2 #(
		.INIT('h8)
	) name872 (
		\memory_reg[24][0]/NET0131 ,
		_w996_,
		_w997_
	);
	LUT2 #(
		.INIT('h8)
	) name873 (
		_w982_,
		_w987_,
		_w998_
	);
	LUT2 #(
		.INIT('h8)
	) name874 (
		\memory_reg[4][0]/NET0131 ,
		_w998_,
		_w999_
	);
	LUT2 #(
		.INIT('h8)
	) name875 (
		_w983_,
		_w993_,
		_w1000_
	);
	LUT2 #(
		.INIT('h8)
	) name876 (
		\memory_reg[16][0]/NET0131 ,
		_w1000_,
		_w1001_
	);
	LUT2 #(
		.INIT('h8)
	) name877 (
		\address_reg[2]/NET0131 ,
		\address_reg[3]/NET0131 ,
		_w1002_
	);
	LUT2 #(
		.INIT('h8)
	) name878 (
		_w983_,
		_w1002_,
		_w1003_
	);
	LUT2 #(
		.INIT('h8)
	) name879 (
		\memory_reg[28][0]/NET0131 ,
		_w1003_,
		_w1004_
	);
	LUT2 #(
		.INIT('h8)
	) name880 (
		\address_reg[1]/NET0131 ,
		\address_reg[4]/NET0131 ,
		_w1005_
	);
	LUT2 #(
		.INIT('h8)
	) name881 (
		_w986_,
		_w1005_,
		_w1006_
	);
	LUT2 #(
		.INIT('h8)
	) name882 (
		\memory_reg[26][0]/NET0131 ,
		_w1006_,
		_w1007_
	);
	LUT2 #(
		.INIT('h8)
	) name883 (
		_w986_,
		_w990_,
		_w1008_
	);
	LUT2 #(
		.INIT('h8)
	) name884 (
		\memory_reg[10][0]/NET0131 ,
		_w1008_,
		_w1009_
	);
	LUT2 #(
		.INIT('h1)
	) name885 (
		\address_reg[0]/NET0131 ,
		_w985_,
		_w1010_
	);
	LUT2 #(
		.INIT('h1)
	) name886 (
		_w989_,
		_w992_,
		_w1011_
	);
	LUT2 #(
		.INIT('h1)
	) name887 (
		_w995_,
		_w997_,
		_w1012_
	);
	LUT2 #(
		.INIT('h1)
	) name888 (
		_w999_,
		_w1001_,
		_w1013_
	);
	LUT2 #(
		.INIT('h1)
	) name889 (
		_w1004_,
		_w1007_,
		_w1014_
	);
	LUT2 #(
		.INIT('h4)
	) name890 (
		_w1009_,
		_w1014_,
		_w1015_
	);
	LUT2 #(
		.INIT('h8)
	) name891 (
		_w1012_,
		_w1013_,
		_w1016_
	);
	LUT2 #(
		.INIT('h8)
	) name892 (
		_w1010_,
		_w1011_,
		_w1017_
	);
	LUT2 #(
		.INIT('h8)
	) name893 (
		_w1016_,
		_w1017_,
		_w1018_
	);
	LUT2 #(
		.INIT('h8)
	) name894 (
		_w1015_,
		_w1018_,
		_w1019_
	);
	LUT2 #(
		.INIT('h8)
	) name895 (
		_w990_,
		_w1002_,
		_w1020_
	);
	LUT2 #(
		.INIT('h8)
	) name896 (
		\memory_reg[15][0]/NET0131 ,
		_w1020_,
		_w1021_
	);
	LUT2 #(
		.INIT('h8)
	) name897 (
		\memory_reg[5][0]/NET0131 ,
		_w998_,
		_w1022_
	);
	LUT2 #(
		.INIT('h8)
	) name898 (
		\memory_reg[9][0]/NET0131 ,
		_w988_,
		_w1023_
	);
	LUT2 #(
		.INIT('h8)
	) name899 (
		\memory_reg[21][0]/NET0131 ,
		_w984_,
		_w1024_
	);
	LUT2 #(
		.INIT('h8)
	) name900 (
		\memory_reg[25][0]/NET0131 ,
		_w996_,
		_w1025_
	);
	LUT2 #(
		.INIT('h8)
	) name901 (
		_w993_,
		_w1005_,
		_w1026_
	);
	LUT2 #(
		.INIT('h8)
	) name902 (
		\memory_reg[19][0]/NET0131 ,
		_w1026_,
		_w1027_
	);
	LUT2 #(
		.INIT('h8)
	) name903 (
		\memory_reg[17][0]/NET0131 ,
		_w1000_,
		_w1028_
	);
	LUT2 #(
		.INIT('h8)
	) name904 (
		\memory_reg[27][0]/NET0131 ,
		_w1006_,
		_w1029_
	);
	LUT2 #(
		.INIT('h2)
	) name905 (
		\address_reg[0]/NET0131 ,
		_w1021_,
		_w1030_
	);
	LUT2 #(
		.INIT('h1)
	) name906 (
		_w1022_,
		_w1023_,
		_w1031_
	);
	LUT2 #(
		.INIT('h1)
	) name907 (
		_w1024_,
		_w1025_,
		_w1032_
	);
	LUT2 #(
		.INIT('h1)
	) name908 (
		_w1027_,
		_w1028_,
		_w1033_
	);
	LUT2 #(
		.INIT('h4)
	) name909 (
		_w1029_,
		_w1033_,
		_w1034_
	);
	LUT2 #(
		.INIT('h8)
	) name910 (
		_w1031_,
		_w1032_,
		_w1035_
	);
	LUT2 #(
		.INIT('h8)
	) name911 (
		_w1030_,
		_w1035_,
		_w1036_
	);
	LUT2 #(
		.INIT('h8)
	) name912 (
		_w1034_,
		_w1036_,
		_w1037_
	);
	LUT2 #(
		.INIT('h1)
	) name913 (
		_w1019_,
		_w1037_,
		_w1038_
	);
	LUT2 #(
		.INIT('h8)
	) name914 (
		\address_reg[0]/NET0131 ,
		_w1003_,
		_w1039_
	);
	LUT2 #(
		.INIT('h8)
	) name915 (
		\memory_reg[29][0]/NET0131 ,
		_w1039_,
		_w1040_
	);
	LUT2 #(
		.INIT('h8)
	) name916 (
		_w982_,
		_w1005_,
		_w1041_
	);
	LUT2 #(
		.INIT('h1)
	) name917 (
		\address_reg[0]/NET0131 ,
		\memory_reg[22][0]/NET0131 ,
		_w1042_
	);
	LUT2 #(
		.INIT('h2)
	) name918 (
		\address_reg[0]/NET0131 ,
		\memory_reg[23][0]/NET0131 ,
		_w1043_
	);
	LUT2 #(
		.INIT('h1)
	) name919 (
		_w1042_,
		_w1043_,
		_w1044_
	);
	LUT2 #(
		.INIT('h8)
	) name920 (
		_w1041_,
		_w1044_,
		_w1045_
	);
	LUT2 #(
		.INIT('h8)
	) name921 (
		_w1002_,
		_w1005_,
		_w1046_
	);
	LUT2 #(
		.INIT('h1)
	) name922 (
		\address_reg[0]/NET0131 ,
		\memory_reg[30][0]/NET0131 ,
		_w1047_
	);
	LUT2 #(
		.INIT('h2)
	) name923 (
		\address_reg[0]/NET0131 ,
		\memory_reg[31][0]/NET0131 ,
		_w1048_
	);
	LUT2 #(
		.INIT('h1)
	) name924 (
		_w1047_,
		_w1048_,
		_w1049_
	);
	LUT2 #(
		.INIT('h8)
	) name925 (
		_w1046_,
		_w1049_,
		_w1050_
	);
	LUT2 #(
		.INIT('h8)
	) name926 (
		_w987_,
		_w1002_,
		_w1051_
	);
	LUT2 #(
		.INIT('h1)
	) name927 (
		\address_reg[0]/NET0131 ,
		\memory_reg[12][0]/NET0131 ,
		_w1052_
	);
	LUT2 #(
		.INIT('h2)
	) name928 (
		\address_reg[0]/NET0131 ,
		\memory_reg[13][0]/NET0131 ,
		_w1053_
	);
	LUT2 #(
		.INIT('h1)
	) name929 (
		_w1052_,
		_w1053_,
		_w1054_
	);
	LUT2 #(
		.INIT('h8)
	) name930 (
		_w1051_,
		_w1054_,
		_w1055_
	);
	LUT2 #(
		.INIT('h8)
	) name931 (
		\memory_reg[18][0]/NET0131 ,
		_w1026_,
		_w1056_
	);
	LUT2 #(
		.INIT('h8)
	) name932 (
		\memory_reg[14][0]/NET0131 ,
		_w1020_,
		_w1057_
	);
	LUT2 #(
		.INIT('h1)
	) name933 (
		\address_reg[0]/NET0131 ,
		_w1056_,
		_w1058_
	);
	LUT2 #(
		.INIT('h4)
	) name934 (
		_w1057_,
		_w1058_,
		_w1059_
	);
	LUT2 #(
		.INIT('h8)
	) name935 (
		\memory_reg[3][0]/NET0131 ,
		_w994_,
		_w1060_
	);
	LUT2 #(
		.INIT('h8)
	) name936 (
		\memory_reg[11][0]/NET0131 ,
		_w1008_,
		_w1061_
	);
	LUT2 #(
		.INIT('h2)
	) name937 (
		\address_reg[0]/NET0131 ,
		_w1060_,
		_w1062_
	);
	LUT2 #(
		.INIT('h4)
	) name938 (
		_w1061_,
		_w1062_,
		_w1063_
	);
	LUT2 #(
		.INIT('h1)
	) name939 (
		_w1059_,
		_w1063_,
		_w1064_
	);
	LUT2 #(
		.INIT('h2)
	) name940 (
		\address_reg[0]/NET0131 ,
		\address_reg[3]/NET0131 ,
		_w1065_
	);
	LUT2 #(
		.INIT('h8)
	) name941 (
		\address_reg[2]/NET0131 ,
		_w1065_,
		_w1066_
	);
	LUT2 #(
		.INIT('h8)
	) name942 (
		\memory_reg[7][0]/NET0131 ,
		_w990_,
		_w1067_
	);
	LUT2 #(
		.INIT('h8)
	) name943 (
		_w1066_,
		_w1067_,
		_w1068_
	);
	LUT2 #(
		.INIT('h8)
	) name944 (
		_w987_,
		_w993_,
		_w1069_
	);
	LUT2 #(
		.INIT('h1)
	) name945 (
		\address_reg[0]/NET0131 ,
		\memory_reg[0][0]/NET0131 ,
		_w1070_
	);
	LUT2 #(
		.INIT('h2)
	) name946 (
		\address_reg[0]/NET0131 ,
		\memory_reg[1][0]/NET0131 ,
		_w1071_
	);
	LUT2 #(
		.INIT('h1)
	) name947 (
		_w1070_,
		_w1071_,
		_w1072_
	);
	LUT2 #(
		.INIT('h8)
	) name948 (
		_w1069_,
		_w1072_,
		_w1073_
	);
	LUT2 #(
		.INIT('h1)
	) name949 (
		_w1045_,
		_w1050_,
		_w1074_
	);
	LUT2 #(
		.INIT('h1)
	) name950 (
		_w1055_,
		_w1068_,
		_w1075_
	);
	LUT2 #(
		.INIT('h4)
	) name951 (
		_w1073_,
		_w1075_,
		_w1076_
	);
	LUT2 #(
		.INIT('h4)
	) name952 (
		_w1040_,
		_w1074_,
		_w1077_
	);
	LUT2 #(
		.INIT('h8)
	) name953 (
		_w1076_,
		_w1077_,
		_w1078_
	);
	LUT2 #(
		.INIT('h4)
	) name954 (
		_w1064_,
		_w1078_,
		_w1079_
	);
	LUT2 #(
		.INIT('h4)
	) name955 (
		_w1038_,
		_w1079_,
		_w1080_
	);
	LUT2 #(
		.INIT('h8)
	) name956 (
		\memory_reg[14][1]/NET0131 ,
		_w1020_,
		_w1081_
	);
	LUT2 #(
		.INIT('h8)
	) name957 (
		\memory_reg[2][1]/NET0131 ,
		_w994_,
		_w1082_
	);
	LUT2 #(
		.INIT('h8)
	) name958 (
		\memory_reg[6][1]/NET0131 ,
		_w991_,
		_w1083_
	);
	LUT2 #(
		.INIT('h8)
	) name959 (
		\memory_reg[8][1]/NET0131 ,
		_w988_,
		_w1084_
	);
	LUT2 #(
		.INIT('h8)
	) name960 (
		\memory_reg[16][1]/NET0131 ,
		_w1000_,
		_w1085_
	);
	LUT2 #(
		.INIT('h8)
	) name961 (
		\memory_reg[4][1]/NET0131 ,
		_w998_,
		_w1086_
	);
	LUT2 #(
		.INIT('h1)
	) name962 (
		\address_reg[0]/NET0131 ,
		_w1081_,
		_w1087_
	);
	LUT2 #(
		.INIT('h1)
	) name963 (
		_w1082_,
		_w1083_,
		_w1088_
	);
	LUT2 #(
		.INIT('h1)
	) name964 (
		_w1084_,
		_w1085_,
		_w1089_
	);
	LUT2 #(
		.INIT('h4)
	) name965 (
		_w1086_,
		_w1089_,
		_w1090_
	);
	LUT2 #(
		.INIT('h8)
	) name966 (
		_w1087_,
		_w1088_,
		_w1091_
	);
	LUT2 #(
		.INIT('h8)
	) name967 (
		_w1090_,
		_w1091_,
		_w1092_
	);
	LUT2 #(
		.INIT('h8)
	) name968 (
		\memory_reg[27][1]/NET0131 ,
		_w1006_,
		_w1093_
	);
	LUT2 #(
		.INIT('h8)
	) name969 (
		\memory_reg[19][1]/NET0131 ,
		_w1026_,
		_w1094_
	);
	LUT2 #(
		.INIT('h8)
	) name970 (
		\memory_reg[3][1]/NET0131 ,
		_w994_,
		_w1095_
	);
	LUT2 #(
		.INIT('h8)
	) name971 (
		\memory_reg[13][1]/NET0131 ,
		_w1051_,
		_w1096_
	);
	LUT2 #(
		.INIT('h8)
	) name972 (
		\memory_reg[25][1]/NET0131 ,
		_w996_,
		_w1097_
	);
	LUT2 #(
		.INIT('h8)
	) name973 (
		\memory_reg[9][1]/NET0131 ,
		_w988_,
		_w1098_
	);
	LUT2 #(
		.INIT('h2)
	) name974 (
		\address_reg[0]/NET0131 ,
		_w1093_,
		_w1099_
	);
	LUT2 #(
		.INIT('h1)
	) name975 (
		_w1094_,
		_w1095_,
		_w1100_
	);
	LUT2 #(
		.INIT('h1)
	) name976 (
		_w1096_,
		_w1097_,
		_w1101_
	);
	LUT2 #(
		.INIT('h4)
	) name977 (
		_w1098_,
		_w1101_,
		_w1102_
	);
	LUT2 #(
		.INIT('h8)
	) name978 (
		_w1099_,
		_w1100_,
		_w1103_
	);
	LUT2 #(
		.INIT('h8)
	) name979 (
		_w1102_,
		_w1103_,
		_w1104_
	);
	LUT2 #(
		.INIT('h1)
	) name980 (
		_w1092_,
		_w1104_,
		_w1105_
	);
	LUT2 #(
		.INIT('h8)
	) name981 (
		\memory_reg[29][1]/NET0131 ,
		_w1039_,
		_w1106_
	);
	LUT2 #(
		.INIT('h8)
	) name982 (
		\memory_reg[0][1]/NET0131 ,
		_w1069_,
		_w1107_
	);
	LUT2 #(
		.INIT('h8)
	) name983 (
		\memory_reg[18][1]/NET0131 ,
		_w1026_,
		_w1108_
	);
	LUT2 #(
		.INIT('h1)
	) name984 (
		\address_reg[0]/NET0131 ,
		_w1107_,
		_w1109_
	);
	LUT2 #(
		.INIT('h4)
	) name985 (
		_w1108_,
		_w1109_,
		_w1110_
	);
	LUT2 #(
		.INIT('h8)
	) name986 (
		\memory_reg[21][1]/NET0131 ,
		_w984_,
		_w1111_
	);
	LUT2 #(
		.INIT('h8)
	) name987 (
		\memory_reg[7][1]/NET0131 ,
		_w991_,
		_w1112_
	);
	LUT2 #(
		.INIT('h2)
	) name988 (
		\address_reg[0]/NET0131 ,
		_w1111_,
		_w1113_
	);
	LUT2 #(
		.INIT('h4)
	) name989 (
		_w1112_,
		_w1113_,
		_w1114_
	);
	LUT2 #(
		.INIT('h1)
	) name990 (
		_w1110_,
		_w1114_,
		_w1115_
	);
	LUT2 #(
		.INIT('h1)
	) name991 (
		\address_reg[0]/NET0131 ,
		\memory_reg[22][1]/NET0131 ,
		_w1116_
	);
	LUT2 #(
		.INIT('h2)
	) name992 (
		\address_reg[0]/NET0131 ,
		\memory_reg[23][1]/NET0131 ,
		_w1117_
	);
	LUT2 #(
		.INIT('h1)
	) name993 (
		_w1116_,
		_w1117_,
		_w1118_
	);
	LUT2 #(
		.INIT('h8)
	) name994 (
		_w1041_,
		_w1118_,
		_w1119_
	);
	LUT2 #(
		.INIT('h1)
	) name995 (
		\address_reg[0]/NET0131 ,
		\memory_reg[30][1]/NET0131 ,
		_w1120_
	);
	LUT2 #(
		.INIT('h2)
	) name996 (
		\address_reg[0]/NET0131 ,
		\memory_reg[31][1]/NET0131 ,
		_w1121_
	);
	LUT2 #(
		.INIT('h1)
	) name997 (
		_w1120_,
		_w1121_,
		_w1122_
	);
	LUT2 #(
		.INIT('h8)
	) name998 (
		_w1046_,
		_w1122_,
		_w1123_
	);
	LUT2 #(
		.INIT('h1)
	) name999 (
		\address_reg[0]/NET0131 ,
		\memory_reg[10][1]/NET0131 ,
		_w1124_
	);
	LUT2 #(
		.INIT('h2)
	) name1000 (
		\address_reg[0]/NET0131 ,
		\memory_reg[11][1]/NET0131 ,
		_w1125_
	);
	LUT2 #(
		.INIT('h1)
	) name1001 (
		_w1124_,
		_w1125_,
		_w1126_
	);
	LUT2 #(
		.INIT('h8)
	) name1002 (
		_w1008_,
		_w1126_,
		_w1127_
	);
	LUT2 #(
		.INIT('h8)
	) name1003 (
		\memory_reg[17][1]/NET0131 ,
		_w1000_,
		_w1128_
	);
	LUT2 #(
		.INIT('h8)
	) name1004 (
		\memory_reg[1][1]/NET0131 ,
		_w1069_,
		_w1129_
	);
	LUT2 #(
		.INIT('h8)
	) name1005 (
		\memory_reg[15][1]/NET0131 ,
		_w1020_,
		_w1130_
	);
	LUT2 #(
		.INIT('h8)
	) name1006 (
		\memory_reg[5][1]/NET0131 ,
		_w998_,
		_w1131_
	);
	LUT2 #(
		.INIT('h2)
	) name1007 (
		\address_reg[0]/NET0131 ,
		_w1128_,
		_w1132_
	);
	LUT2 #(
		.INIT('h1)
	) name1008 (
		_w1129_,
		_w1130_,
		_w1133_
	);
	LUT2 #(
		.INIT('h4)
	) name1009 (
		_w1131_,
		_w1133_,
		_w1134_
	);
	LUT2 #(
		.INIT('h8)
	) name1010 (
		_w1132_,
		_w1134_,
		_w1135_
	);
	LUT2 #(
		.INIT('h8)
	) name1011 (
		\memory_reg[12][1]/NET0131 ,
		_w1051_,
		_w1136_
	);
	LUT2 #(
		.INIT('h8)
	) name1012 (
		\memory_reg[28][1]/NET0131 ,
		_w1003_,
		_w1137_
	);
	LUT2 #(
		.INIT('h8)
	) name1013 (
		\memory_reg[20][1]/NET0131 ,
		_w984_,
		_w1138_
	);
	LUT2 #(
		.INIT('h8)
	) name1014 (
		\memory_reg[26][1]/NET0131 ,
		_w1006_,
		_w1139_
	);
	LUT2 #(
		.INIT('h8)
	) name1015 (
		\memory_reg[24][1]/NET0131 ,
		_w996_,
		_w1140_
	);
	LUT2 #(
		.INIT('h1)
	) name1016 (
		\address_reg[0]/NET0131 ,
		_w1136_,
		_w1141_
	);
	LUT2 #(
		.INIT('h1)
	) name1017 (
		_w1137_,
		_w1138_,
		_w1142_
	);
	LUT2 #(
		.INIT('h1)
	) name1018 (
		_w1139_,
		_w1140_,
		_w1143_
	);
	LUT2 #(
		.INIT('h8)
	) name1019 (
		_w1142_,
		_w1143_,
		_w1144_
	);
	LUT2 #(
		.INIT('h8)
	) name1020 (
		_w1141_,
		_w1144_,
		_w1145_
	);
	LUT2 #(
		.INIT('h1)
	) name1021 (
		_w1135_,
		_w1145_,
		_w1146_
	);
	LUT2 #(
		.INIT('h1)
	) name1022 (
		_w1119_,
		_w1123_,
		_w1147_
	);
	LUT2 #(
		.INIT('h4)
	) name1023 (
		_w1127_,
		_w1147_,
		_w1148_
	);
	LUT2 #(
		.INIT('h4)
	) name1024 (
		_w1106_,
		_w1148_,
		_w1149_
	);
	LUT2 #(
		.INIT('h4)
	) name1025 (
		_w1115_,
		_w1149_,
		_w1150_
	);
	LUT2 #(
		.INIT('h4)
	) name1026 (
		_w1105_,
		_w1150_,
		_w1151_
	);
	LUT2 #(
		.INIT('h4)
	) name1027 (
		_w1146_,
		_w1151_,
		_w1152_
	);
	LUT2 #(
		.INIT('h1)
	) name1028 (
		\address_reg[0]/NET0131 ,
		\address_reg[3]/NET0131 ,
		_w1153_
	);
	LUT2 #(
		.INIT('h4)
	) name1029 (
		\address_reg[2]/NET0131 ,
		_w1153_,
		_w1154_
	);
	LUT2 #(
		.INIT('h8)
	) name1030 (
		\wr_reg/NET0131 ,
		_w987_,
		_w1155_
	);
	LUT2 #(
		.INIT('h8)
	) name1031 (
		_w1154_,
		_w1155_,
		_w1156_
	);
	LUT2 #(
		.INIT('h4)
	) name1032 (
		\address_reg[0]/NET0131 ,
		\address_reg[3]/NET0131 ,
		_w1157_
	);
	LUT2 #(
		.INIT('h4)
	) name1033 (
		\address_reg[2]/NET0131 ,
		_w1157_,
		_w1158_
	);
	LUT2 #(
		.INIT('h8)
	) name1034 (
		\wr_reg/NET0131 ,
		_w990_,
		_w1159_
	);
	LUT2 #(
		.INIT('h8)
	) name1035 (
		_w1158_,
		_w1159_,
		_w1160_
	);
	LUT2 #(
		.INIT('h8)
	) name1036 (
		\address_reg[0]/NET0131 ,
		\address_reg[3]/NET0131 ,
		_w1161_
	);
	LUT2 #(
		.INIT('h4)
	) name1037 (
		\address_reg[2]/NET0131 ,
		_w1161_,
		_w1162_
	);
	LUT2 #(
		.INIT('h8)
	) name1038 (
		_w1159_,
		_w1162_,
		_w1163_
	);
	LUT2 #(
		.INIT('h8)
	) name1039 (
		\address_reg[2]/NET0131 ,
		_w1157_,
		_w1164_
	);
	LUT2 #(
		.INIT('h8)
	) name1040 (
		_w1155_,
		_w1164_,
		_w1165_
	);
	LUT2 #(
		.INIT('h8)
	) name1041 (
		\address_reg[2]/NET0131 ,
		_w1161_,
		_w1166_
	);
	LUT2 #(
		.INIT('h8)
	) name1042 (
		_w1155_,
		_w1166_,
		_w1167_
	);
	LUT2 #(
		.INIT('h8)
	) name1043 (
		_w1159_,
		_w1164_,
		_w1168_
	);
	LUT2 #(
		.INIT('h8)
	) name1044 (
		_w1159_,
		_w1166_,
		_w1169_
	);
	LUT2 #(
		.INIT('h8)
	) name1045 (
		\wr_reg/NET0131 ,
		_w983_,
		_w1170_
	);
	LUT2 #(
		.INIT('h8)
	) name1046 (
		_w1154_,
		_w1170_,
		_w1171_
	);
	LUT2 #(
		.INIT('h4)
	) name1047 (
		\address_reg[2]/NET0131 ,
		_w1065_,
		_w1172_
	);
	LUT2 #(
		.INIT('h8)
	) name1048 (
		_w1170_,
		_w1172_,
		_w1173_
	);
	LUT2 #(
		.INIT('h8)
	) name1049 (
		\wr_reg/NET0131 ,
		_w1005_,
		_w1174_
	);
	LUT2 #(
		.INIT('h8)
	) name1050 (
		_w1154_,
		_w1174_,
		_w1175_
	);
	LUT2 #(
		.INIT('h8)
	) name1051 (
		_w1172_,
		_w1174_,
		_w1176_
	);
	LUT2 #(
		.INIT('h8)
	) name1052 (
		_w1155_,
		_w1172_,
		_w1177_
	);
	LUT2 #(
		.INIT('h8)
	) name1053 (
		\address_reg[2]/NET0131 ,
		_w1153_,
		_w1178_
	);
	LUT2 #(
		.INIT('h8)
	) name1054 (
		_w1170_,
		_w1178_,
		_w1179_
	);
	LUT2 #(
		.INIT('h8)
	) name1055 (
		_w1066_,
		_w1170_,
		_w1180_
	);
	LUT2 #(
		.INIT('h8)
	) name1056 (
		_w1174_,
		_w1178_,
		_w1181_
	);
	LUT2 #(
		.INIT('h8)
	) name1057 (
		_w1066_,
		_w1174_,
		_w1182_
	);
	LUT2 #(
		.INIT('h8)
	) name1058 (
		_w1158_,
		_w1170_,
		_w1183_
	);
	LUT2 #(
		.INIT('h8)
	) name1059 (
		_w1162_,
		_w1170_,
		_w1184_
	);
	LUT2 #(
		.INIT('h8)
	) name1060 (
		_w1158_,
		_w1174_,
		_w1185_
	);
	LUT2 #(
		.INIT('h8)
	) name1061 (
		_w1162_,
		_w1174_,
		_w1186_
	);
	LUT2 #(
		.INIT('h8)
	) name1062 (
		_w1164_,
		_w1170_,
		_w1187_
	);
	LUT2 #(
		.INIT('h8)
	) name1063 (
		\wr_reg/NET0131 ,
		_w1039_,
		_w1188_
	);
	LUT2 #(
		.INIT('h8)
	) name1064 (
		_w1154_,
		_w1159_,
		_w1189_
	);
	LUT2 #(
		.INIT('h8)
	) name1065 (
		_w1164_,
		_w1174_,
		_w1190_
	);
	LUT2 #(
		.INIT('h8)
	) name1066 (
		_w1166_,
		_w1174_,
		_w1191_
	);
	LUT2 #(
		.INIT('h8)
	) name1067 (
		_w1159_,
		_w1172_,
		_w1192_
	);
	LUT2 #(
		.INIT('h8)
	) name1068 (
		_w1155_,
		_w1178_,
		_w1193_
	);
	LUT2 #(
		.INIT('h8)
	) name1069 (
		_w1066_,
		_w1155_,
		_w1194_
	);
	LUT2 #(
		.INIT('h8)
	) name1070 (
		_w1159_,
		_w1178_,
		_w1195_
	);
	LUT2 #(
		.INIT('h8)
	) name1071 (
		_w1066_,
		_w1159_,
		_w1196_
	);
	LUT2 #(
		.INIT('h8)
	) name1072 (
		_w1155_,
		_w1158_,
		_w1197_
	);
	LUT2 #(
		.INIT('h8)
	) name1073 (
		_w1155_,
		_w1162_,
		_w1198_
	);
	assign \_al_n0  = 1'b0;
	assign \_al_n1  = 1'b0;
	assign \count_reg[0]/P0001  = \count_reg[0]/NET0131 ;
	assign \g10376/_0_  = _w127_ ;
	assign \g11078/_0_  = _w219_ ;
	assign \g11102/_0_  = _w262_ ;
	assign \g11126/_0_  = _w315_ ;
	assign \g11156/_0_  = _w330_ ;
	assign \g11299/_0_  = _w372_ ;
	assign \g11308/_0_  = _w398_ ;
	assign \g11318/_0_  = _w414_ ;
	assign \g11346/_0_  = _w442_ ;
	assign \g11378/_0_  = _w451_ ;
	assign \g11516/_0_  = _w472_ ;
	assign \g63/_0_  = _w500_ ;
	assign \g8501/_0_  = _w525_ ;
	assign \g8516/_0_  = _w534_ ;
	assign \g8517/_0_  = _w551_ ;
	assign \g8519/_0_  = _w572_ ;
	assign \g8520/_0_  = _w585_ ;
	assign \g8522/_0_  = _w611_ ;
	assign \g8526/_0_  = _w634_ ;
	assign \g8529/_2_  = _w653_ ;
	assign \g8545/_0_  = _w667_ ;
	assign \g8546/_0_  = _w690_ ;
	assign \g8547/_0_  = _w702_ ;
	assign \g8555/_0_  = _w708_ ;
	assign \g8556/_0_  = _w720_ ;
	assign \g8557/_0_  = _w734_ ;
	assign \g8558/_0_  = _w747_ ;
	assign \g8559/_0_  = _w764_ ;
	assign \g8560/_0_  = _w771_ ;
	assign \g8562/_0_  = _w776_ ;
	assign \g8563/_0_  = _w781_ ;
	assign \g8581/_0_  = _w789_ ;
	assign \g8586/_0_  = _w802_ ;
	assign \g8591/_0_  = _w811_ ;
	assign \g8594/_0_  = _w824_ ;
	assign \g8606/_0_  = _w832_ ;
	assign \g8608/_0_  = _w845_ ;
	assign \g8647/_0_  = _w849_ ;
	assign \g8659/_0_  = _w859_ ;
	assign \g8695/_0_  = _w863_ ;
	assign \g8784/_0_  = _w912_ ;
	assign \g8797/_0_  = _w916_ ;
	assign \g8854/_2_  = _w939_ ;
	assign \g8869/_0_  = _w948_ ;
	assign \g8871/_0_  = _w951_ ;
	assign \g8889/_0_  = _w956_ ;
	assign \g8891/_0_  = _w961_ ;
	assign \g8892/_0_  = _w966_ ;
	assign \g8894/_0_  = _w971_ ;
	assign \g8970/_0_  = _w978_ ;
	assign \g8975/_0_  = _w980_ ;
	assign \g8992/_0_  = _w981_ ;
	assign \g9180/_0_  = _w1080_ ;
	assign \g9183/_0_  = _w1152_ ;
	assign \g9511/u3_syn_4  = _w1156_ ;
	assign \g9513/u3_syn_4  = _w1160_ ;
	assign \g9515/u3_syn_4  = _w1163_ ;
	assign \g9517/u3_syn_4  = _w1165_ ;
	assign \g9519/u3_syn_4  = _w1167_ ;
	assign \g9521/u3_syn_4  = _w1168_ ;
	assign \g9523/u3_syn_4  = _w1169_ ;
	assign \g9525/u3_syn_4  = _w1171_ ;
	assign \g9527/u3_syn_4  = _w1173_ ;
	assign \g9529/u3_syn_4  = _w1175_ ;
	assign \g9531/u3_syn_4  = _w1176_ ;
	assign \g9533/u3_syn_4  = _w1177_ ;
	assign \g9535/u3_syn_4  = _w1179_ ;
	assign \g9537/u3_syn_4  = _w1180_ ;
	assign \g9539/u3_syn_4  = _w1181_ ;
	assign \g9541/u3_syn_4  = _w1182_ ;
	assign \g9543/u3_syn_4  = _w1183_ ;
	assign \g9545/u3_syn_4  = _w1184_ ;
	assign \g9547/u3_syn_4  = _w1185_ ;
	assign \g9549/u3_syn_4  = _w1186_ ;
	assign \g9551/u3_syn_4  = _w1187_ ;
	assign \g9553/u3_syn_4  = _w1188_ ;
	assign \g9555/u3_syn_4  = _w1189_ ;
	assign \g9557/u3_syn_4  = _w1190_ ;
	assign \g9559/u3_syn_4  = _w1191_ ;
	assign \g9560/u3_syn_4  = _w1192_ ;
	assign \g9562/u3_syn_4  = _w1193_ ;
	assign \g9564/u3_syn_4  = _w1194_ ;
	assign \g9566/u3_syn_4  = _w1195_ ;
	assign \g9568/u3_syn_4  = _w1196_ ;
	assign \g9570/u3_syn_4  = _w1197_ ;
	assign \g9572/u3_syn_4  = _w1198_ ;
endmodule;