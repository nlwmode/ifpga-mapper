module top (\cont_reg[0]/NET0131 , \cont_reg[1]/NET0131 , \cont_reg[2]/NET0131 , \cont_reg[3]/NET0131 , \cont_reg[4]/NET0131 , \cont_reg[5]/NET0131 , \cont_reg[6]/NET0131 , \cont_reg[7]/NET0131 , \mar_reg[0]/NET0131 , \mar_reg[1]/NET0131 , \mar_reg[2]/NET0131 , \mar_reg[3]/NET0131 , \punti_retta[3]_pad , \punti_retta[4]_pad , \punti_retta[6]_pad , \punti_retta[7]_pad , \punti_retta_reg[0]/NET0131 , \punti_retta_reg[1]/NET0131 , \punti_retta_reg[2]/NET0131 , \punti_retta_reg[5]/NET0131 , start_pad, \stato_reg[0]/NET0131 , \stato_reg[1]/NET0131 , \stato_reg[2]/NET0131 , \t_reg[1]/NET0131 , \t_reg[2]/NET0131 , \t_reg[3]/NET0131 , \t_reg[4]/NET0131 , \t_reg[5]/NET0131 , \t_reg[6]/NET0131 , \x_reg[0]/NET0131 , \x_reg[1]/NET0131 , \x_reg[2]/NET0131 , \x_reg[3]/NET0131 , \x_reg[4]/NET0131 , \x_reg[5]/NET0131 , \x_reg[6]/NET0131 , \x_reg[7]/NET0131 , \y_reg[0]/NET0131 , \y_reg[1]/NET0131 , \y_reg[2]/NET0131 , \y_reg[3]/NET0131 , \_al_n0 , \_al_n1 , \g2119/_0_ , \g2123/_0_ , \g2129/_0_ , \g2133/_0_ , \g2136/_0_ , \g2140/_0_ , \g2141/_0_ , \g2151/_0_ , \g2152/_0_ , \g2166/_0_ , \g2167/_0_ , \g2180/_0_ , \g2181/_0_ , \g2199/_0_ , \g2225/_0_ , \g2227/_0_ , \g2242/_0_ , \g2243/_0_ , \g2272/_0_ , \g2273/_0_ , \g2274/_0_ , \g2275/_0_ , \g2284/_0_ , \g2289/_0_ , \g2303/_0_ , \g2304/_0_ , \g2308/_0_ , \g2309/_0_ , \g2310/_0_ , \g2311/_0_ , \g2312/_0_ , \g2346/_0_ , \g2973/_0_ , \g2984/_0_ , \g3052/_0_ , \g3176/_0_ , \g3277/_0_ , \g3306/_0_ , \g3366/_0_ , \g3371/_0_ , \g3398/_0_ );
	input \cont_reg[0]/NET0131  ;
	input \cont_reg[1]/NET0131  ;
	input \cont_reg[2]/NET0131  ;
	input \cont_reg[3]/NET0131  ;
	input \cont_reg[4]/NET0131  ;
	input \cont_reg[5]/NET0131  ;
	input \cont_reg[6]/NET0131  ;
	input \cont_reg[7]/NET0131  ;
	input \mar_reg[0]/NET0131  ;
	input \mar_reg[1]/NET0131  ;
	input \mar_reg[2]/NET0131  ;
	input \mar_reg[3]/NET0131  ;
	input \punti_retta[3]_pad  ;
	input \punti_retta[4]_pad  ;
	input \punti_retta[6]_pad  ;
	input \punti_retta[7]_pad  ;
	input \punti_retta_reg[0]/NET0131  ;
	input \punti_retta_reg[1]/NET0131  ;
	input \punti_retta_reg[2]/NET0131  ;
	input \punti_retta_reg[5]/NET0131  ;
	input start_pad ;
	input \stato_reg[0]/NET0131  ;
	input \stato_reg[1]/NET0131  ;
	input \stato_reg[2]/NET0131  ;
	input \t_reg[1]/NET0131  ;
	input \t_reg[2]/NET0131  ;
	input \t_reg[3]/NET0131  ;
	input \t_reg[4]/NET0131  ;
	input \t_reg[5]/NET0131  ;
	input \t_reg[6]/NET0131  ;
	input \x_reg[0]/NET0131  ;
	input \x_reg[1]/NET0131  ;
	input \x_reg[2]/NET0131  ;
	input \x_reg[3]/NET0131  ;
	input \x_reg[4]/NET0131  ;
	input \x_reg[5]/NET0131  ;
	input \x_reg[6]/NET0131  ;
	input \x_reg[7]/NET0131  ;
	input \y_reg[0]/NET0131  ;
	input \y_reg[1]/NET0131  ;
	input \y_reg[2]/NET0131  ;
	input \y_reg[3]/NET0131  ;
	output \_al_n0  ;
	output \_al_n1  ;
	output \g2119/_0_  ;
	output \g2123/_0_  ;
	output \g2129/_0_  ;
	output \g2133/_0_  ;
	output \g2136/_0_  ;
	output \g2140/_0_  ;
	output \g2141/_0_  ;
	output \g2151/_0_  ;
	output \g2152/_0_  ;
	output \g2166/_0_  ;
	output \g2167/_0_  ;
	output \g2180/_0_  ;
	output \g2181/_0_  ;
	output \g2199/_0_  ;
	output \g2225/_0_  ;
	output \g2227/_0_  ;
	output \g2242/_0_  ;
	output \g2243/_0_  ;
	output \g2272/_0_  ;
	output \g2273/_0_  ;
	output \g2274/_0_  ;
	output \g2275/_0_  ;
	output \g2284/_0_  ;
	output \g2289/_0_  ;
	output \g2303/_0_  ;
	output \g2304/_0_  ;
	output \g2308/_0_  ;
	output \g2309/_0_  ;
	output \g2310/_0_  ;
	output \g2311/_0_  ;
	output \g2312/_0_  ;
	output \g2346/_0_  ;
	output \g2973/_0_  ;
	output \g2984/_0_  ;
	output \g3052/_0_  ;
	output \g3176/_0_  ;
	output \g3277/_0_  ;
	output \g3306/_0_  ;
	output \g3366/_0_  ;
	output \g3371/_0_  ;
	output \g3398/_0_  ;
	wire _w274_ ;
	wire _w273_ ;
	wire _w272_ ;
	wire _w271_ ;
	wire _w270_ ;
	wire _w269_ ;
	wire _w268_ ;
	wire _w267_ ;
	wire _w266_ ;
	wire _w265_ ;
	wire _w264_ ;
	wire _w263_ ;
	wire _w262_ ;
	wire _w261_ ;
	wire _w260_ ;
	wire _w259_ ;
	wire _w258_ ;
	wire _w257_ ;
	wire _w256_ ;
	wire _w255_ ;
	wire _w254_ ;
	wire _w253_ ;
	wire _w252_ ;
	wire _w251_ ;
	wire _w250_ ;
	wire _w249_ ;
	wire _w248_ ;
	wire _w247_ ;
	wire _w246_ ;
	wire _w245_ ;
	wire _w244_ ;
	wire _w243_ ;
	wire _w242_ ;
	wire _w241_ ;
	wire _w240_ ;
	wire _w239_ ;
	wire _w238_ ;
	wire _w237_ ;
	wire _w236_ ;
	wire _w235_ ;
	wire _w234_ ;
	wire _w233_ ;
	wire _w232_ ;
	wire _w231_ ;
	wire _w230_ ;
	wire _w229_ ;
	wire _w228_ ;
	wire _w227_ ;
	wire _w226_ ;
	wire _w225_ ;
	wire _w224_ ;
	wire _w223_ ;
	wire _w222_ ;
	wire _w221_ ;
	wire _w220_ ;
	wire _w219_ ;
	wire _w218_ ;
	wire _w217_ ;
	wire _w216_ ;
	wire _w215_ ;
	wire _w214_ ;
	wire _w213_ ;
	wire _w212_ ;
	wire _w211_ ;
	wire _w210_ ;
	wire _w209_ ;
	wire _w208_ ;
	wire _w207_ ;
	wire _w206_ ;
	wire _w205_ ;
	wire _w204_ ;
	wire _w203_ ;
	wire _w202_ ;
	wire _w201_ ;
	wire _w200_ ;
	wire _w199_ ;
	wire _w198_ ;
	wire _w197_ ;
	wire _w196_ ;
	wire _w195_ ;
	wire _w194_ ;
	wire _w193_ ;
	wire _w192_ ;
	wire _w191_ ;
	wire _w190_ ;
	wire _w189_ ;
	wire _w188_ ;
	wire _w187_ ;
	wire _w186_ ;
	wire _w185_ ;
	wire _w184_ ;
	wire _w183_ ;
	wire _w182_ ;
	wire _w181_ ;
	wire _w180_ ;
	wire _w179_ ;
	wire _w178_ ;
	wire _w177_ ;
	wire _w176_ ;
	wire _w175_ ;
	wire _w174_ ;
	wire _w173_ ;
	wire _w172_ ;
	wire _w171_ ;
	wire _w102_ ;
	wire _w101_ ;
	wire _w100_ ;
	wire _w99_ ;
	wire _w98_ ;
	wire _w97_ ;
	wire _w96_ ;
	wire _w95_ ;
	wire _w94_ ;
	wire _w93_ ;
	wire _w92_ ;
	wire _w91_ ;
	wire _w90_ ;
	wire _w89_ ;
	wire _w88_ ;
	wire _w87_ ;
	wire _w86_ ;
	wire _w85_ ;
	wire _w84_ ;
	wire _w83_ ;
	wire _w82_ ;
	wire _w81_ ;
	wire _w80_ ;
	wire _w79_ ;
	wire _w78_ ;
	wire _w77_ ;
	wire _w76_ ;
	wire _w75_ ;
	wire _w74_ ;
	wire _w73_ ;
	wire _w56_ ;
	wire _w55_ ;
	wire _w54_ ;
	wire _w53_ ;
	wire _w52_ ;
	wire _w51_ ;
	wire _w50_ ;
	wire _w49_ ;
	wire _w48_ ;
	wire _w47_ ;
	wire _w46_ ;
	wire _w45_ ;
	wire _w44_ ;
	wire _w57_ ;
	wire _w58_ ;
	wire _w59_ ;
	wire _w60_ ;
	wire _w61_ ;
	wire _w62_ ;
	wire _w63_ ;
	wire _w64_ ;
	wire _w65_ ;
	wire _w66_ ;
	wire _w67_ ;
	wire _w68_ ;
	wire _w69_ ;
	wire _w70_ ;
	wire _w71_ ;
	wire _w72_ ;
	wire _w103_ ;
	wire _w104_ ;
	wire _w105_ ;
	wire _w106_ ;
	wire _w107_ ;
	wire _w108_ ;
	wire _w109_ ;
	wire _w110_ ;
	wire _w111_ ;
	wire _w112_ ;
	wire _w113_ ;
	wire _w114_ ;
	wire _w115_ ;
	wire _w116_ ;
	wire _w117_ ;
	wire _w118_ ;
	wire _w119_ ;
	wire _w120_ ;
	wire _w121_ ;
	wire _w122_ ;
	wire _w123_ ;
	wire _w124_ ;
	wire _w125_ ;
	wire _w126_ ;
	wire _w127_ ;
	wire _w128_ ;
	wire _w129_ ;
	wire _w130_ ;
	wire _w131_ ;
	wire _w132_ ;
	wire _w133_ ;
	wire _w134_ ;
	wire _w135_ ;
	wire _w136_ ;
	wire _w137_ ;
	wire _w138_ ;
	wire _w139_ ;
	wire _w140_ ;
	wire _w141_ ;
	wire _w142_ ;
	wire _w143_ ;
	wire _w144_ ;
	wire _w145_ ;
	wire _w146_ ;
	wire _w147_ ;
	wire _w148_ ;
	wire _w149_ ;
	wire _w150_ ;
	wire _w151_ ;
	wire _w152_ ;
	wire _w153_ ;
	wire _w154_ ;
	wire _w155_ ;
	wire _w156_ ;
	wire _w157_ ;
	wire _w158_ ;
	wire _w159_ ;
	wire _w160_ ;
	wire _w161_ ;
	wire _w162_ ;
	wire _w163_ ;
	wire _w164_ ;
	wire _w165_ ;
	wire _w166_ ;
	wire _w167_ ;
	wire _w168_ ;
	wire _w169_ ;
	wire _w170_ ;
	LUT3 #(
		.INIT('h40)
	) name0 (
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		\stato_reg[2]/NET0131 ,
		_w44_
	);
	LUT4 #(
		.INIT('h0001)
	) name1 (
		\x_reg[4]/NET0131 ,
		\x_reg[5]/NET0131 ,
		\x_reg[6]/NET0131 ,
		\x_reg[7]/NET0131 ,
		_w45_
	);
	LUT4 #(
		.INIT('h0004)
	) name2 (
		\x_reg[0]/NET0131 ,
		\x_reg[1]/NET0131 ,
		\x_reg[2]/NET0131 ,
		\x_reg[3]/NET0131 ,
		_w46_
	);
	LUT4 #(
		.INIT('h8000)
	) name3 (
		\cont_reg[0]/NET0131 ,
		\cont_reg[1]/NET0131 ,
		\cont_reg[2]/NET0131 ,
		\cont_reg[3]/NET0131 ,
		_w47_
	);
	LUT3 #(
		.INIT('h80)
	) name4 (
		_w45_,
		_w46_,
		_w47_,
		_w48_
	);
	LUT4 #(
		.INIT('h8000)
	) name5 (
		\cont_reg[4]/NET0131 ,
		_w45_,
		_w46_,
		_w47_,
		_w49_
	);
	LUT3 #(
		.INIT('h80)
	) name6 (
		\mar_reg[0]/NET0131 ,
		\mar_reg[1]/NET0131 ,
		\mar_reg[2]/NET0131 ,
		_w50_
	);
	LUT4 #(
		.INIT('h8000)
	) name7 (
		\mar_reg[0]/NET0131 ,
		\mar_reg[1]/NET0131 ,
		\mar_reg[2]/NET0131 ,
		\mar_reg[3]/NET0131 ,
		_w51_
	);
	LUT3 #(
		.INIT('h08)
	) name8 (
		\cont_reg[5]/NET0131 ,
		_w49_,
		_w51_,
		_w52_
	);
	LUT2 #(
		.INIT('h8)
	) name9 (
		\stato_reg[1]/NET0131 ,
		\stato_reg[2]/NET0131 ,
		_w53_
	);
	LUT4 #(
		.INIT('hf008)
	) name10 (
		start_pad,
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		\stato_reg[2]/NET0131 ,
		_w54_
	);
	LUT4 #(
		.INIT('h48ea)
	) name11 (
		\cont_reg[6]/NET0131 ,
		_w44_,
		_w52_,
		_w54_,
		_w55_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name12 (
		\cont_reg[4]/NET0131 ,
		_w45_,
		_w46_,
		_w47_,
		_w56_
	);
	LUT3 #(
		.INIT('h8c)
	) name13 (
		\cont_reg[4]/NET0131 ,
		_w44_,
		_w51_,
		_w57_
	);
	LUT2 #(
		.INIT('h2)
	) name14 (
		\cont_reg[4]/NET0131 ,
		_w54_,
		_w58_
	);
	LUT4 #(
		.INIT('hffe0)
	) name15 (
		_w51_,
		_w56_,
		_w57_,
		_w58_,
		_w59_
	);
	LUT2 #(
		.INIT('h2)
	) name16 (
		\cont_reg[7]/NET0131 ,
		_w54_,
		_w60_
	);
	LUT2 #(
		.INIT('h8)
	) name17 (
		\cont_reg[5]/NET0131 ,
		\cont_reg[6]/NET0131 ,
		_w61_
	);
	LUT4 #(
		.INIT('h0905)
	) name18 (
		\cont_reg[7]/NET0131 ,
		_w49_,
		_w51_,
		_w61_,
		_w62_
	);
	LUT3 #(
		.INIT('h8c)
	) name19 (
		\cont_reg[7]/NET0131 ,
		_w44_,
		_w51_,
		_w63_
	);
	LUT3 #(
		.INIT('hba)
	) name20 (
		_w60_,
		_w62_,
		_w63_,
		_w64_
	);
	LUT4 #(
		.INIT('hf004)
	) name21 (
		start_pad,
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		\stato_reg[2]/NET0131 ,
		_w65_
	);
	LUT2 #(
		.INIT('h4)
	) name22 (
		start_pad,
		_w51_,
		_w66_
	);
	LUT4 #(
		.INIT('h7300)
	) name23 (
		start_pad,
		_w44_,
		_w51_,
		_w65_,
		_w67_
	);
	LUT2 #(
		.INIT('h2)
	) name24 (
		\punti_retta[6]_pad ,
		_w67_,
		_w68_
	);
	LUT3 #(
		.INIT('h40)
	) name25 (
		start_pad,
		_w44_,
		_w51_,
		_w69_
	);
	LUT4 #(
		.INIT('h6c00)
	) name26 (
		\cont_reg[5]/NET0131 ,
		\cont_reg[6]/NET0131 ,
		_w49_,
		_w69_,
		_w70_
	);
	LUT2 #(
		.INIT('he)
	) name27 (
		_w68_,
		_w70_,
		_w71_
	);
	LUT2 #(
		.INIT('h2)
	) name28 (
		\cont_reg[3]/NET0131 ,
		_w54_,
		_w72_
	);
	LUT3 #(
		.INIT('h80)
	) name29 (
		\cont_reg[0]/NET0131 ,
		_w45_,
		_w46_,
		_w73_
	);
	LUT4 #(
		.INIT('h8000)
	) name30 (
		\cont_reg[0]/NET0131 ,
		\cont_reg[1]/NET0131 ,
		_w45_,
		_w46_,
		_w74_
	);
	LUT4 #(
		.INIT('h0e0c)
	) name31 (
		\cont_reg[2]/NET0131 ,
		\cont_reg[3]/NET0131 ,
		_w48_,
		_w74_,
		_w75_
	);
	LUT3 #(
		.INIT('h8c)
	) name32 (
		\cont_reg[3]/NET0131 ,
		_w44_,
		_w51_,
		_w76_
	);
	LUT4 #(
		.INIT('hfecc)
	) name33 (
		_w51_,
		_w72_,
		_w75_,
		_w76_,
		_w77_
	);
	LUT2 #(
		.INIT('h2)
	) name34 (
		\punti_retta_reg[2]/NET0131 ,
		_w65_,
		_w78_
	);
	LUT2 #(
		.INIT('h8)
	) name35 (
		\punti_retta_reg[2]/NET0131 ,
		start_pad,
		_w79_
	);
	LUT2 #(
		.INIT('h2)
	) name36 (
		_w51_,
		_w79_,
		_w80_
	);
	LUT4 #(
		.INIT('hed00)
	) name37 (
		\cont_reg[2]/NET0131 ,
		start_pad,
		_w74_,
		_w80_,
		_w81_
	);
	LUT3 #(
		.INIT('hc8)
	) name38 (
		\punti_retta_reg[2]/NET0131 ,
		_w44_,
		_w51_,
		_w82_
	);
	LUT3 #(
		.INIT('hba)
	) name39 (
		_w78_,
		_w81_,
		_w82_,
		_w83_
	);
	LUT2 #(
		.INIT('h8)
	) name40 (
		\punti_retta_reg[5]/NET0131 ,
		start_pad,
		_w84_
	);
	LUT2 #(
		.INIT('h2)
	) name41 (
		_w51_,
		_w84_,
		_w85_
	);
	LUT4 #(
		.INIT('hed00)
	) name42 (
		\cont_reg[5]/NET0131 ,
		start_pad,
		_w49_,
		_w85_,
		_w86_
	);
	LUT3 #(
		.INIT('hc8)
	) name43 (
		\punti_retta_reg[5]/NET0131 ,
		_w44_,
		_w51_,
		_w87_
	);
	LUT2 #(
		.INIT('h2)
	) name44 (
		\punti_retta_reg[5]/NET0131 ,
		_w65_,
		_w88_
	);
	LUT3 #(
		.INIT('hf4)
	) name45 (
		_w86_,
		_w87_,
		_w88_,
		_w89_
	);
	LUT3 #(
		.INIT('h6a)
	) name46 (
		\cont_reg[0]/NET0131 ,
		_w45_,
		_w46_,
		_w90_
	);
	LUT4 #(
		.INIT('h44c4)
	) name47 (
		_w44_,
		_w65_,
		_w66_,
		_w90_,
		_w91_
	);
	LUT3 #(
		.INIT('h80)
	) name48 (
		_w44_,
		_w66_,
		_w90_,
		_w92_
	);
	LUT3 #(
		.INIT('hf2)
	) name49 (
		\punti_retta_reg[0]/NET0131 ,
		_w91_,
		_w92_,
		_w93_
	);
	LUT2 #(
		.INIT('h2)
	) name50 (
		\punti_retta_reg[1]/NET0131 ,
		_w67_,
		_w94_
	);
	LUT3 #(
		.INIT('h48)
	) name51 (
		\cont_reg[1]/NET0131 ,
		_w69_,
		_w73_,
		_w95_
	);
	LUT2 #(
		.INIT('he)
	) name52 (
		_w94_,
		_w95_,
		_w96_
	);
	LUT3 #(
		.INIT('h8c)
	) name53 (
		\cont_reg[5]/NET0131 ,
		_w44_,
		_w51_,
		_w97_
	);
	LUT4 #(
		.INIT('hf600)
	) name54 (
		\cont_reg[5]/NET0131 ,
		_w49_,
		_w51_,
		_w97_,
		_w98_
	);
	LUT2 #(
		.INIT('h2)
	) name55 (
		\cont_reg[5]/NET0131 ,
		_w54_,
		_w99_
	);
	LUT2 #(
		.INIT('he)
	) name56 (
		_w98_,
		_w99_,
		_w100_
	);
	LUT3 #(
		.INIT('h8c)
	) name57 (
		\cont_reg[2]/NET0131 ,
		_w44_,
		_w51_,
		_w101_
	);
	LUT4 #(
		.INIT('hde00)
	) name58 (
		\cont_reg[2]/NET0131 ,
		_w51_,
		_w74_,
		_w101_,
		_w102_
	);
	LUT2 #(
		.INIT('h2)
	) name59 (
		\cont_reg[2]/NET0131 ,
		_w54_,
		_w103_
	);
	LUT2 #(
		.INIT('he)
	) name60 (
		_w102_,
		_w103_,
		_w104_
	);
	LUT4 #(
		.INIT('h0080)
	) name61 (
		\cont_reg[0]/NET0131 ,
		_w45_,
		_w46_,
		_w51_,
		_w105_
	);
	LUT4 #(
		.INIT('h4e8a)
	) name62 (
		\cont_reg[1]/NET0131 ,
		_w44_,
		_w54_,
		_w105_,
		_w106_
	);
	LUT4 #(
		.INIT('h0095)
	) name63 (
		\cont_reg[0]/NET0131 ,
		_w45_,
		_w46_,
		_w51_,
		_w107_
	);
	LUT3 #(
		.INIT('h8c)
	) name64 (
		\cont_reg[0]/NET0131 ,
		_w44_,
		_w51_,
		_w108_
	);
	LUT2 #(
		.INIT('h2)
	) name65 (
		\cont_reg[0]/NET0131 ,
		_w54_,
		_w109_
	);
	LUT3 #(
		.INIT('hf4)
	) name66 (
		_w107_,
		_w108_,
		_w109_,
		_w110_
	);
	LUT3 #(
		.INIT('h08)
	) name67 (
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		\stato_reg[2]/NET0131 ,
		_w111_
	);
	LUT4 #(
		.INIT('h0515)
	) name68 (
		\mar_reg[3]/NET0131 ,
		_w44_,
		_w50_,
		_w111_,
		_w112_
	);
	LUT4 #(
		.INIT('hf0c8)
	) name69 (
		start_pad,
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		\stato_reg[2]/NET0131 ,
		_w113_
	);
	LUT4 #(
		.INIT('h4500)
	) name70 (
		_w44_,
		_w51_,
		_w111_,
		_w113_,
		_w114_
	);
	LUT2 #(
		.INIT('h1)
	) name71 (
		_w112_,
		_w114_,
		_w115_
	);
	LUT2 #(
		.INIT('h2)
	) name72 (
		\mar_reg[0]/NET0131 ,
		_w113_,
		_w116_
	);
	LUT4 #(
		.INIT('h1040)
	) name73 (
		\mar_reg[0]/NET0131 ,
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		\stato_reg[2]/NET0131 ,
		_w117_
	);
	LUT3 #(
		.INIT('h07)
	) name74 (
		_w44_,
		_w51_,
		_w117_,
		_w118_
	);
	LUT2 #(
		.INIT('hb)
	) name75 (
		_w116_,
		_w118_,
		_w119_
	);
	LUT3 #(
		.INIT('h10)
	) name76 (
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		\stato_reg[2]/NET0131 ,
		_w120_
	);
	LUT2 #(
		.INIT('h6)
	) name77 (
		\t_reg[1]/NET0131 ,
		\x_reg[1]/NET0131 ,
		_w121_
	);
	LUT3 #(
		.INIT('h04)
	) name78 (
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		\stato_reg[2]/NET0131 ,
		_w122_
	);
	LUT4 #(
		.INIT('h59dd)
	) name79 (
		\mar_reg[0]/NET0131 ,
		\mar_reg[1]/NET0131 ,
		\mar_reg[2]/NET0131 ,
		\mar_reg[3]/NET0131 ,
		_w123_
	);
	LUT4 #(
		.INIT('h7707)
	) name80 (
		_w120_,
		_w121_,
		_w122_,
		_w123_,
		_w124_
	);
	LUT4 #(
		.INIT('h4b00)
	) name81 (
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		\stato_reg[2]/NET0131 ,
		\x_reg[1]/NET0131 ,
		_w125_
	);
	LUT2 #(
		.INIT('h8)
	) name82 (
		\x_reg[0]/NET0131 ,
		\y_reg[0]/NET0131 ,
		_w126_
	);
	LUT2 #(
		.INIT('h6)
	) name83 (
		\x_reg[1]/NET0131 ,
		\y_reg[1]/NET0131 ,
		_w127_
	);
	LUT3 #(
		.INIT('h20)
	) name84 (
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		\stato_reg[2]/NET0131 ,
		_w128_
	);
	LUT4 #(
		.INIT('h5115)
	) name85 (
		_w125_,
		_w128_,
		_w126_,
		_w127_,
		_w129_
	);
	LUT2 #(
		.INIT('h7)
	) name86 (
		_w124_,
		_w129_,
		_w130_
	);
	LUT2 #(
		.INIT('h2)
	) name87 (
		\mar_reg[1]/NET0131 ,
		_w113_,
		_w131_
	);
	LUT2 #(
		.INIT('h6)
	) name88 (
		\mar_reg[0]/NET0131 ,
		\mar_reg[1]/NET0131 ,
		_w132_
	);
	LUT4 #(
		.INIT('h0577)
	) name89 (
		_w44_,
		_w51_,
		_w111_,
		_w132_,
		_w133_
	);
	LUT2 #(
		.INIT('hb)
	) name90 (
		_w131_,
		_w133_,
		_w134_
	);
	LUT2 #(
		.INIT('h2)
	) name91 (
		\mar_reg[2]/NET0131 ,
		_w113_,
		_w135_
	);
	LUT3 #(
		.INIT('h78)
	) name92 (
		\mar_reg[0]/NET0131 ,
		\mar_reg[1]/NET0131 ,
		\mar_reg[2]/NET0131 ,
		_w136_
	);
	LUT4 #(
		.INIT('h0577)
	) name93 (
		_w44_,
		_w51_,
		_w111_,
		_w136_,
		_w137_
	);
	LUT2 #(
		.INIT('hb)
	) name94 (
		_w135_,
		_w137_,
		_w138_
	);
	LUT4 #(
		.INIT('h5b00)
	) name95 (
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		\stato_reg[2]/NET0131 ,
		\x_reg[0]/NET0131 ,
		_w139_
	);
	LUT3 #(
		.INIT('hde)
	) name96 (
		\mar_reg[1]/NET0131 ,
		\mar_reg[2]/NET0131 ,
		\mar_reg[3]/NET0131 ,
		_w140_
	);
	LUT2 #(
		.INIT('h6)
	) name97 (
		\x_reg[0]/NET0131 ,
		\y_reg[0]/NET0131 ,
		_w141_
	);
	LUT4 #(
		.INIT('h31f5)
	) name98 (
		_w122_,
		_w128_,
		_w140_,
		_w141_,
		_w142_
	);
	LUT2 #(
		.INIT('hb)
	) name99 (
		_w139_,
		_w142_,
		_w143_
	);
	LUT4 #(
		.INIT('h6f00)
	) name100 (
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		\stato_reg[2]/NET0131 ,
		\y_reg[1]/NET0131 ,
		_w144_
	);
	LUT3 #(
		.INIT('hf2)
	) name101 (
		_w120_,
		_w123_,
		_w144_,
		_w145_
	);
	LUT3 #(
		.INIT('h15)
	) name102 (
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		\stato_reg[2]/NET0131 ,
		_w146_
	);
	LUT4 #(
		.INIT('h4101)
	) name103 (
		start_pad,
		\stato_reg[1]/NET0131 ,
		\stato_reg[2]/NET0131 ,
		_w51_,
		_w147_
	);
	LUT2 #(
		.INIT('he)
	) name104 (
		_w146_,
		_w147_,
		_w148_
	);
	LUT4 #(
		.INIT('hf3c7)
	) name105 (
		start_pad,
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		\stato_reg[2]/NET0131 ,
		_w149_
	);
	LUT4 #(
		.INIT('hb0ff)
	) name106 (
		start_pad,
		_w51_,
		_w53_,
		_w149_,
		_w150_
	);
	LUT4 #(
		.INIT('h0800)
	) name107 (
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		\stato_reg[2]/NET0131 ,
		\x_reg[5]/NET0131 ,
		_w151_
	);
	LUT4 #(
		.INIT('h7700)
	) name108 (
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		\stato_reg[2]/NET0131 ,
		\t_reg[6]/NET0131 ,
		_w152_
	);
	LUT2 #(
		.INIT('he)
	) name109 (
		_w151_,
		_w152_,
		_w153_
	);
	LUT4 #(
		.INIT('h0800)
	) name110 (
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		\stato_reg[2]/NET0131 ,
		\x_reg[4]/NET0131 ,
		_w154_
	);
	LUT4 #(
		.INIT('h7700)
	) name111 (
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		\stato_reg[2]/NET0131 ,
		\t_reg[5]/NET0131 ,
		_w155_
	);
	LUT2 #(
		.INIT('he)
	) name112 (
		_w154_,
		_w155_,
		_w156_
	);
	LUT4 #(
		.INIT('hf3fd)
	) name113 (
		\mar_reg[0]/NET0131 ,
		\mar_reg[1]/NET0131 ,
		\mar_reg[2]/NET0131 ,
		\mar_reg[3]/NET0131 ,
		_w157_
	);
	LUT4 #(
		.INIT('h6f00)
	) name114 (
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		\stato_reg[2]/NET0131 ,
		\y_reg[2]/NET0131 ,
		_w158_
	);
	LUT3 #(
		.INIT('hf2)
	) name115 (
		_w120_,
		_w157_,
		_w158_,
		_w159_
	);
	LUT4 #(
		.INIT('hfbfd)
	) name116 (
		\mar_reg[0]/NET0131 ,
		\mar_reg[1]/NET0131 ,
		\mar_reg[2]/NET0131 ,
		\mar_reg[3]/NET0131 ,
		_w160_
	);
	LUT4 #(
		.INIT('h6f00)
	) name117 (
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		\stato_reg[2]/NET0131 ,
		\y_reg[3]/NET0131 ,
		_w161_
	);
	LUT3 #(
		.INIT('hf2)
	) name118 (
		_w120_,
		_w160_,
		_w161_,
		_w162_
	);
	LUT3 #(
		.INIT('hc7)
	) name119 (
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		\stato_reg[2]/NET0131 ,
		_w163_
	);
	LUT4 #(
		.INIT('h80ff)
	) name120 (
		start_pad,
		_w51_,
		_w53_,
		_w163_,
		_w164_
	);
	LUT4 #(
		.INIT('h0800)
	) name121 (
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		\stato_reg[2]/NET0131 ,
		\x_reg[0]/NET0131 ,
		_w165_
	);
	LUT4 #(
		.INIT('h7700)
	) name122 (
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		\stato_reg[2]/NET0131 ,
		\t_reg[1]/NET0131 ,
		_w166_
	);
	LUT2 #(
		.INIT('he)
	) name123 (
		_w165_,
		_w166_,
		_w167_
	);
	LUT4 #(
		.INIT('h0800)
	) name124 (
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		\stato_reg[2]/NET0131 ,
		\x_reg[1]/NET0131 ,
		_w168_
	);
	LUT4 #(
		.INIT('h7700)
	) name125 (
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		\stato_reg[2]/NET0131 ,
		\t_reg[2]/NET0131 ,
		_w169_
	);
	LUT2 #(
		.INIT('he)
	) name126 (
		_w168_,
		_w169_,
		_w170_
	);
	LUT4 #(
		.INIT('h0800)
	) name127 (
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		\stato_reg[2]/NET0131 ,
		\x_reg[2]/NET0131 ,
		_w171_
	);
	LUT4 #(
		.INIT('h7700)
	) name128 (
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		\stato_reg[2]/NET0131 ,
		\t_reg[3]/NET0131 ,
		_w172_
	);
	LUT2 #(
		.INIT('he)
	) name129 (
		_w171_,
		_w172_,
		_w173_
	);
	LUT4 #(
		.INIT('h0800)
	) name130 (
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		\stato_reg[2]/NET0131 ,
		\x_reg[3]/NET0131 ,
		_w174_
	);
	LUT4 #(
		.INIT('h7700)
	) name131 (
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		\stato_reg[2]/NET0131 ,
		\t_reg[4]/NET0131 ,
		_w175_
	);
	LUT2 #(
		.INIT('he)
	) name132 (
		_w174_,
		_w175_,
		_w176_
	);
	LUT4 #(
		.INIT('h6f00)
	) name133 (
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		\stato_reg[2]/NET0131 ,
		\y_reg[0]/NET0131 ,
		_w177_
	);
	LUT3 #(
		.INIT('hf2)
	) name134 (
		_w120_,
		_w140_,
		_w177_,
		_w178_
	);
	LUT2 #(
		.INIT('h2)
	) name135 (
		\punti_retta[4]_pad ,
		_w65_,
		_w179_
	);
	LUT2 #(
		.INIT('h8)
	) name136 (
		\punti_retta[4]_pad ,
		start_pad,
		_w180_
	);
	LUT2 #(
		.INIT('h2)
	) name137 (
		_w51_,
		_w180_,
		_w181_
	);
	LUT3 #(
		.INIT('hc8)
	) name138 (
		\punti_retta[4]_pad ,
		_w44_,
		_w51_,
		_w182_
	);
	LUT4 #(
		.INIT('h4f00)
	) name139 (
		start_pad,
		_w56_,
		_w181_,
		_w182_,
		_w183_
	);
	LUT2 #(
		.INIT('he)
	) name140 (
		_w179_,
		_w183_,
		_w184_
	);
	LUT2 #(
		.INIT('h1)
	) name141 (
		\x_reg[4]/NET0131 ,
		\y_reg[3]/NET0131 ,
		_w185_
	);
	LUT2 #(
		.INIT('h1)
	) name142 (
		\x_reg[2]/NET0131 ,
		\y_reg[2]/NET0131 ,
		_w186_
	);
	LUT4 #(
		.INIT('hec80)
	) name143 (
		\x_reg[0]/NET0131 ,
		\x_reg[1]/NET0131 ,
		\y_reg[0]/NET0131 ,
		\y_reg[1]/NET0131 ,
		_w187_
	);
	LUT2 #(
		.INIT('h1)
	) name144 (
		\x_reg[3]/NET0131 ,
		\y_reg[3]/NET0131 ,
		_w188_
	);
	LUT4 #(
		.INIT('h00e8)
	) name145 (
		\x_reg[2]/NET0131 ,
		\y_reg[2]/NET0131 ,
		_w187_,
		_w188_,
		_w189_
	);
	LUT3 #(
		.INIT('hf8)
	) name146 (
		\x_reg[5]/NET0131 ,
		\x_reg[6]/NET0131 ,
		\y_reg[3]/NET0131 ,
		_w190_
	);
	LUT2 #(
		.INIT('h8)
	) name147 (
		\x_reg[3]/NET0131 ,
		\y_reg[3]/NET0131 ,
		_w191_
	);
	LUT3 #(
		.INIT('h1f)
	) name148 (
		\x_reg[3]/NET0131 ,
		\x_reg[4]/NET0131 ,
		\y_reg[3]/NET0131 ,
		_w192_
	);
	LUT3 #(
		.INIT('h1f)
	) name149 (
		\x_reg[5]/NET0131 ,
		\x_reg[6]/NET0131 ,
		\y_reg[3]/NET0131 ,
		_w193_
	);
	LUT2 #(
		.INIT('h8)
	) name150 (
		_w192_,
		_w193_,
		_w194_
	);
	LUT4 #(
		.INIT('hbf00)
	) name151 (
		_w185_,
		_w189_,
		_w190_,
		_w194_,
		_w195_
	);
	LUT2 #(
		.INIT('h1)
	) name152 (
		\t_reg[5]/NET0131 ,
		\x_reg[5]/NET0131 ,
		_w196_
	);
	LUT2 #(
		.INIT('h1)
	) name153 (
		\t_reg[4]/NET0131 ,
		\x_reg[4]/NET0131 ,
		_w197_
	);
	LUT4 #(
		.INIT('ha080)
	) name154 (
		\t_reg[1]/NET0131 ,
		\t_reg[2]/NET0131 ,
		\x_reg[1]/NET0131 ,
		\x_reg[2]/NET0131 ,
		_w198_
	);
	LUT4 #(
		.INIT('h137f)
	) name155 (
		\t_reg[1]/NET0131 ,
		\t_reg[2]/NET0131 ,
		\x_reg[1]/NET0131 ,
		\x_reg[2]/NET0131 ,
		_w199_
	);
	LUT2 #(
		.INIT('h1)
	) name156 (
		\t_reg[3]/NET0131 ,
		\x_reg[3]/NET0131 ,
		_w200_
	);
	LUT2 #(
		.INIT('h8)
	) name157 (
		\t_reg[4]/NET0131 ,
		\x_reg[4]/NET0131 ,
		_w201_
	);
	LUT4 #(
		.INIT('h135f)
	) name158 (
		\t_reg[3]/NET0131 ,
		\t_reg[4]/NET0131 ,
		\x_reg[3]/NET0131 ,
		\x_reg[4]/NET0131 ,
		_w202_
	);
	LUT4 #(
		.INIT('h0155)
	) name159 (
		_w197_,
		_w199_,
		_w200_,
		_w202_,
		_w203_
	);
	LUT2 #(
		.INIT('h8)
	) name160 (
		\t_reg[5]/NET0131 ,
		\x_reg[5]/NET0131 ,
		_w204_
	);
	LUT4 #(
		.INIT('h135f)
	) name161 (
		\t_reg[5]/NET0131 ,
		\t_reg[6]/NET0131 ,
		\x_reg[5]/NET0131 ,
		\x_reg[6]/NET0131 ,
		_w205_
	);
	LUT2 #(
		.INIT('h1)
	) name162 (
		\t_reg[6]/NET0131 ,
		\x_reg[6]/NET0131 ,
		_w206_
	);
	LUT2 #(
		.INIT('h2)
	) name163 (
		_w120_,
		_w206_,
		_w207_
	);
	LUT4 #(
		.INIT('h4f00)
	) name164 (
		_w196_,
		_w203_,
		_w205_,
		_w207_,
		_w208_
	);
	LUT4 #(
		.INIT('h4b00)
	) name165 (
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		\stato_reg[2]/NET0131 ,
		\x_reg[7]/NET0131 ,
		_w209_
	);
	LUT3 #(
		.INIT('h0d)
	) name166 (
		_w122_,
		_w160_,
		_w209_,
		_w210_
	);
	LUT4 #(
		.INIT('hf2ff)
	) name167 (
		_w128_,
		_w195_,
		_w208_,
		_w210_,
		_w211_
	);
	LUT2 #(
		.INIT('h6)
	) name168 (
		\x_reg[2]/NET0131 ,
		\y_reg[2]/NET0131 ,
		_w212_
	);
	LUT3 #(
		.INIT('h28)
	) name169 (
		_w128_,
		_w187_,
		_w212_,
		_w213_
	);
	LUT4 #(
		.INIT('h2080)
	) name170 (
		\t_reg[1]/NET0131 ,
		\t_reg[2]/NET0131 ,
		\x_reg[1]/NET0131 ,
		\x_reg[2]/NET0131 ,
		_w214_
	);
	LUT4 #(
		.INIT('h4c13)
	) name171 (
		\t_reg[1]/NET0131 ,
		\t_reg[2]/NET0131 ,
		\x_reg[1]/NET0131 ,
		\x_reg[2]/NET0131 ,
		_w215_
	);
	LUT3 #(
		.INIT('h02)
	) name172 (
		_w120_,
		_w215_,
		_w214_,
		_w216_
	);
	LUT4 #(
		.INIT('h4b00)
	) name173 (
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		\stato_reg[2]/NET0131 ,
		\x_reg[2]/NET0131 ,
		_w217_
	);
	LUT3 #(
		.INIT('h0d)
	) name174 (
		_w122_,
		_w157_,
		_w217_,
		_w218_
	);
	LUT3 #(
		.INIT('hef)
	) name175 (
		_w216_,
		_w213_,
		_w218_,
		_w219_
	);
	LUT2 #(
		.INIT('h6)
	) name176 (
		\x_reg[3]/NET0131 ,
		\y_reg[3]/NET0131 ,
		_w220_
	);
	LUT4 #(
		.INIT('he800)
	) name177 (
		\x_reg[2]/NET0131 ,
		\y_reg[2]/NET0131 ,
		_w187_,
		_w220_,
		_w221_
	);
	LUT4 #(
		.INIT('h0017)
	) name178 (
		\x_reg[2]/NET0131 ,
		\y_reg[2]/NET0131 ,
		_w187_,
		_w220_,
		_w222_
	);
	LUT3 #(
		.INIT('h02)
	) name179 (
		_w128_,
		_w222_,
		_w221_,
		_w223_
	);
	LUT2 #(
		.INIT('h6)
	) name180 (
		\t_reg[3]/NET0131 ,
		\x_reg[3]/NET0131 ,
		_w224_
	);
	LUT3 #(
		.INIT('h82)
	) name181 (
		_w120_,
		_w199_,
		_w224_,
		_w225_
	);
	LUT4 #(
		.INIT('h4b00)
	) name182 (
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		\stato_reg[2]/NET0131 ,
		\x_reg[3]/NET0131 ,
		_w226_
	);
	LUT3 #(
		.INIT('h0d)
	) name183 (
		_w122_,
		_w160_,
		_w226_,
		_w227_
	);
	LUT2 #(
		.INIT('h4)
	) name184 (
		_w225_,
		_w227_,
		_w228_
	);
	LUT2 #(
		.INIT('hb)
	) name185 (
		_w223_,
		_w228_,
		_w229_
	);
	LUT2 #(
		.INIT('h6)
	) name186 (
		\x_reg[5]/NET0131 ,
		\y_reg[3]/NET0131 ,
		_w230_
	);
	LUT4 #(
		.INIT('h00b0)
	) name187 (
		_w185_,
		_w189_,
		_w192_,
		_w230_,
		_w231_
	);
	LUT4 #(
		.INIT('h4f00)
	) name188 (
		_w185_,
		_w189_,
		_w192_,
		_w230_,
		_w232_
	);
	LUT3 #(
		.INIT('h02)
	) name189 (
		_w128_,
		_w232_,
		_w231_,
		_w233_
	);
	LUT4 #(
		.INIT('h9060)
	) name190 (
		\t_reg[5]/NET0131 ,
		\x_reg[5]/NET0131 ,
		_w120_,
		_w203_,
		_w234_
	);
	LUT4 #(
		.INIT('h4b00)
	) name191 (
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		\stato_reg[2]/NET0131 ,
		\x_reg[5]/NET0131 ,
		_w235_
	);
	LUT3 #(
		.INIT('h0d)
	) name192 (
		_w122_,
		_w160_,
		_w235_,
		_w236_
	);
	LUT2 #(
		.INIT('h4)
	) name193 (
		_w234_,
		_w236_,
		_w237_
	);
	LUT2 #(
		.INIT('hb)
	) name194 (
		_w233_,
		_w237_,
		_w238_
	);
	LUT4 #(
		.INIT('h1222)
	) name195 (
		\cont_reg[7]/NET0131 ,
		start_pad,
		_w49_,
		_w61_,
		_w239_
	);
	LUT2 #(
		.INIT('h8)
	) name196 (
		\punti_retta[7]_pad ,
		start_pad,
		_w240_
	);
	LUT2 #(
		.INIT('h2)
	) name197 (
		_w51_,
		_w240_,
		_w241_
	);
	LUT3 #(
		.INIT('hc8)
	) name198 (
		\punti_retta[7]_pad ,
		_w44_,
		_w51_,
		_w242_
	);
	LUT2 #(
		.INIT('h2)
	) name199 (
		\punti_retta[7]_pad ,
		_w65_,
		_w243_
	);
	LUT4 #(
		.INIT('hffb0)
	) name200 (
		_w239_,
		_w241_,
		_w242_,
		_w243_,
		_w244_
	);
	LUT3 #(
		.INIT('hf8)
	) name201 (
		\x_reg[3]/NET0131 ,
		\x_reg[4]/NET0131 ,
		\y_reg[3]/NET0131 ,
		_w245_
	);
	LUT3 #(
		.INIT('h40)
	) name202 (
		_w186_,
		_w187_,
		_w245_,
		_w246_
	);
	LUT4 #(
		.INIT('ha080)
	) name203 (
		\x_reg[2]/NET0131 ,
		\x_reg[3]/NET0131 ,
		\y_reg[2]/NET0131 ,
		\y_reg[3]/NET0131 ,
		_w247_
	);
	LUT3 #(
		.INIT('h51)
	) name204 (
		_w185_,
		_w192_,
		_w247_,
		_w248_
	);
	LUT4 #(
		.INIT('h1117)
	) name205 (
		\x_reg[5]/NET0131 ,
		\y_reg[3]/NET0131 ,
		_w246_,
		_w248_,
		_w249_
	);
	LUT2 #(
		.INIT('h6)
	) name206 (
		\x_reg[6]/NET0131 ,
		\y_reg[3]/NET0131 ,
		_w250_
	);
	LUT3 #(
		.INIT('h82)
	) name207 (
		_w128_,
		_w249_,
		_w250_,
		_w251_
	);
	LUT2 #(
		.INIT('h6)
	) name208 (
		\t_reg[6]/NET0131 ,
		\x_reg[6]/NET0131 ,
		_w252_
	);
	LUT4 #(
		.INIT('h135f)
	) name209 (
		\t_reg[2]/NET0131 ,
		\t_reg[3]/NET0131 ,
		\x_reg[2]/NET0131 ,
		\x_reg[3]/NET0131 ,
		_w253_
	);
	LUT3 #(
		.INIT('h23)
	) name210 (
		_w198_,
		_w200_,
		_w253_,
		_w254_
	);
	LUT4 #(
		.INIT('h0d0c)
	) name211 (
		_w198_,
		_w200_,
		_w201_,
		_w253_,
		_w255_
	);
	LUT4 #(
		.INIT('hfac8)
	) name212 (
		\t_reg[4]/NET0131 ,
		\t_reg[5]/NET0131 ,
		\x_reg[4]/NET0131 ,
		\x_reg[5]/NET0131 ,
		_w256_
	);
	LUT3 #(
		.INIT('h45)
	) name213 (
		_w204_,
		_w255_,
		_w256_,
		_w257_
	);
	LUT4 #(
		.INIT('h4b00)
	) name214 (
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		\stato_reg[2]/NET0131 ,
		\x_reg[6]/NET0131 ,
		_w258_
	);
	LUT3 #(
		.INIT('h0d)
	) name215 (
		_w122_,
		_w160_,
		_w258_,
		_w259_
	);
	LUT4 #(
		.INIT('h7d00)
	) name216 (
		_w120_,
		_w252_,
		_w257_,
		_w259_,
		_w260_
	);
	LUT2 #(
		.INIT('hb)
	) name217 (
		_w251_,
		_w260_,
		_w261_
	);
	LUT2 #(
		.INIT('h2)
	) name218 (
		\punti_retta[3]_pad ,
		_w65_,
		_w262_
	);
	LUT2 #(
		.INIT('h8)
	) name219 (
		\punti_retta[3]_pad ,
		start_pad,
		_w263_
	);
	LUT2 #(
		.INIT('h2)
	) name220 (
		_w51_,
		_w263_,
		_w264_
	);
	LUT3 #(
		.INIT('hc8)
	) name221 (
		\punti_retta[3]_pad ,
		_w44_,
		_w51_,
		_w265_
	);
	LUT4 #(
		.INIT('h4f00)
	) name222 (
		start_pad,
		_w75_,
		_w264_,
		_w265_,
		_w266_
	);
	LUT2 #(
		.INIT('he)
	) name223 (
		_w262_,
		_w266_,
		_w267_
	);
	LUT2 #(
		.INIT('h6)
	) name224 (
		\x_reg[4]/NET0131 ,
		\y_reg[3]/NET0131 ,
		_w268_
	);
	LUT4 #(
		.INIT('h02a8)
	) name225 (
		_w128_,
		_w189_,
		_w191_,
		_w268_,
		_w269_
	);
	LUT2 #(
		.INIT('h6)
	) name226 (
		\t_reg[4]/NET0131 ,
		\x_reg[4]/NET0131 ,
		_w270_
	);
	LUT4 #(
		.INIT('h4b00)
	) name227 (
		\stato_reg[0]/NET0131 ,
		\stato_reg[1]/NET0131 ,
		\stato_reg[2]/NET0131 ,
		\x_reg[4]/NET0131 ,
		_w271_
	);
	LUT3 #(
		.INIT('h0d)
	) name228 (
		_w122_,
		_w160_,
		_w271_,
		_w272_
	);
	LUT4 #(
		.INIT('hd700)
	) name229 (
		_w120_,
		_w254_,
		_w270_,
		_w272_,
		_w273_
	);
	LUT2 #(
		.INIT('hb)
	) name230 (
		_w269_,
		_w273_,
		_w274_
	);
	assign \_al_n0  = 1'b0;
	assign \_al_n1  = 1'b1;
	assign \g2119/_0_  = _w55_ ;
	assign \g2123/_0_  = _w59_ ;
	assign \g2129/_0_  = _w64_ ;
	assign \g2133/_0_  = _w71_ ;
	assign \g2136/_0_  = _w77_ ;
	assign \g2140/_0_  = _w83_ ;
	assign \g2141/_0_  = _w89_ ;
	assign \g2151/_0_  = _w93_ ;
	assign \g2152/_0_  = _w96_ ;
	assign \g2166/_0_  = _w100_ ;
	assign \g2167/_0_  = _w104_ ;
	assign \g2180/_0_  = _w106_ ;
	assign \g2181/_0_  = _w110_ ;
	assign \g2199/_0_  = _w115_ ;
	assign \g2225/_0_  = _w119_ ;
	assign \g2227/_0_  = _w130_ ;
	assign \g2242/_0_  = _w134_ ;
	assign \g2243/_0_  = _w138_ ;
	assign \g2272/_0_  = _w143_ ;
	assign \g2273/_0_  = _w145_ ;
	assign \g2274/_0_  = _w148_ ;
	assign \g2275/_0_  = _w150_ ;
	assign \g2284/_0_  = _w153_ ;
	assign \g2289/_0_  = _w156_ ;
	assign \g2303/_0_  = _w159_ ;
	assign \g2304/_0_  = _w162_ ;
	assign \g2308/_0_  = _w164_ ;
	assign \g2309/_0_  = _w167_ ;
	assign \g2310/_0_  = _w170_ ;
	assign \g2311/_0_  = _w173_ ;
	assign \g2312/_0_  = _w176_ ;
	assign \g2346/_0_  = _w178_ ;
	assign \g2973/_0_  = _w184_ ;
	assign \g2984/_0_  = _w211_ ;
	assign \g3052/_0_  = _w219_ ;
	assign \g3176/_0_  = _w229_ ;
	assign \g3277/_0_  = _w238_ ;
	assign \g3306/_0_  = _w244_ ;
	assign \g3366/_0_  = _w261_ ;
	assign \g3371/_0_  = _w267_ ;
	assign \g3398/_0_  = _w274_ ;
endmodule;