module top( \G0_pad  , \G10_pad  , \G11_pad  , \G12_pad  , \G13_pad  , \G14_pad  , \G15_pad  , \G16_pad  , \G1_pad  , \G22_reg/NET0131  , \G23_reg/NET0131  , \G24_reg/NET0131  , \G25_reg/NET0131  , \G26_reg/NET0131  , \G27_reg/NET0131  , \G28_reg/NET0131  , \G29_reg/NET0131  , \G2_pad  , \G30_reg/NET0131  , \G31_reg/NET0131  , \G32_reg/NET0131  , \G33_reg/NET0131  , \G34_reg/NET0131  , \G35_reg/NET0131  , \G36_reg/NET0131  , \G37_reg/NET0131  , \G38_reg/NET0131  , \G39_reg/NET0131  , \G3_pad  , \G40_reg/NET0131  , \G41_reg/NET0131  , \G42_reg/NET0131  , \G43_reg/NET0131  , \G44_reg/NET0131  , \G45_reg/NET0131  , \G46_reg/NET0131  , \G47_reg/NET0131  , \G48_reg/NET0131  , \G49_reg/NET0131  , \G4_pad  , \G50_reg/NET0131  , \G51_reg/NET0131  , \G52_reg/NET0131  , \G53_reg/NET0131  , \G55_reg/NET0131  , \G56_reg/NET0131  , \G57_reg/NET0131  , \G58_reg/NET0131  , \G59_reg/NET0131  , \G5_pad  , \G60_reg/NET0131  , \G61_reg/NET0131  , \G62_reg/NET0131  , \G63_reg/NET0131  , \G64_reg/NET0131  , \G65_reg/NET0131  , \G66_reg/NET0131  , \G67_reg/NET0131  , \G68_reg/NET0131  , \G69_reg/NET0131  , \G6_pad  , \G70_reg/NET0131  , \G71_reg/NET0131  , \G72_reg/NET0131  , \G73_reg/NET0131  , \G74_reg/NET0131  , \G75_reg/NET0131  , \G76_reg/NET0131  , \G77_reg/NET0131  , \G78_reg/NET0131  , \G79_reg/NET0131  , \G7_pad  , \G80_reg/NET0131  , \G81_reg/NET0131  , \G82_reg/NET0131  , \G83_reg/NET0131  , \G84_reg/NET0131  , \G85_reg/NET0131  , \G86_reg/NET0131  , \G87_reg/NET0131  , \G88_reg/NET0131  , \G89_reg/NET0131  , \G8_pad  , \G90_reg/NET0131  , \G91_reg/NET0131  , \G92_reg/NET0131  , \G94_reg/NET0131  , \G9_pad  , \G701BF_pad  , \G702_pad  , \G727_pad  , \_al_n0  , \_al_n1  , \g2503/_0_  , \g2514/_0_  , \g2516/_0_  , \g2542/_0_  , \g2549/_0_  , \g2553/_0_  , \g2554/_0_  , \g2570/_0_  , \g2574/_0_  , \g2576/_0_  , \g2583/_0_  , \g2588/_0_  , \g2602/_0_  , \g2603/_0_  , \g2604/_0_  , \g2605/_0_  , \g2611/_0_  , \g2614/_0_  , \g2615/_0_  , \g2644/_0_  , \g2657/_0_  , \g2663/_0_  , \g2664/_0_  , \g2666/_0_  , \g2672/_0_  , \g2678/_0_  , \g2681/_0_  , \g2696/_00_  , \g2698/_0_  , \g2699/_0_  , \g2700/_00_  , \g2717/_0_  , \g2719/_0_  , \g2723/_0_  , \g2726/_3_  , \g2735/_0_  , \g2737/_0_  , \g2740/_0_  , \g2785/_0_  , \g2786/_0_  , \g2787/_1__syn_2  , \g2790/_1__syn_2  , \g2798/_2_  , \g2801/_0_  , \g2841/_0_  , \g2844/_0_  , \g2845/_0_  , \g2846/_0_  , \g2860/_0_  , \g2861/_0_  , \g2862/_0_  , \g2864/_0_  , \g2882/_3_  , \g2883/_3_  , \g2887/_3_  , \g2906/_0_  , \g2911/_0_  , \g3282/_0_  , \g3406/_0_  , \g3409/_0_  , \g3506/_0_  , \g3685/_3_  , \g3694/_0_  , \g3743/_0_  , \g3753/_0_  , \g3785/_0_  , \g3835/_0_  , \g3946/_2_  , \g3976/_0_  );
  input \G0_pad  ;
  input \G10_pad  ;
  input \G11_pad  ;
  input \G12_pad  ;
  input \G13_pad  ;
  input \G14_pad  ;
  input \G15_pad  ;
  input \G16_pad  ;
  input \G1_pad  ;
  input \G22_reg/NET0131  ;
  input \G23_reg/NET0131  ;
  input \G24_reg/NET0131  ;
  input \G25_reg/NET0131  ;
  input \G26_reg/NET0131  ;
  input \G27_reg/NET0131  ;
  input \G28_reg/NET0131  ;
  input \G29_reg/NET0131  ;
  input \G2_pad  ;
  input \G30_reg/NET0131  ;
  input \G31_reg/NET0131  ;
  input \G32_reg/NET0131  ;
  input \G33_reg/NET0131  ;
  input \G34_reg/NET0131  ;
  input \G35_reg/NET0131  ;
  input \G36_reg/NET0131  ;
  input \G37_reg/NET0131  ;
  input \G38_reg/NET0131  ;
  input \G39_reg/NET0131  ;
  input \G3_pad  ;
  input \G40_reg/NET0131  ;
  input \G41_reg/NET0131  ;
  input \G42_reg/NET0131  ;
  input \G43_reg/NET0131  ;
  input \G44_reg/NET0131  ;
  input \G45_reg/NET0131  ;
  input \G46_reg/NET0131  ;
  input \G47_reg/NET0131  ;
  input \G48_reg/NET0131  ;
  input \G49_reg/NET0131  ;
  input \G4_pad  ;
  input \G50_reg/NET0131  ;
  input \G51_reg/NET0131  ;
  input \G52_reg/NET0131  ;
  input \G53_reg/NET0131  ;
  input \G55_reg/NET0131  ;
  input \G56_reg/NET0131  ;
  input \G57_reg/NET0131  ;
  input \G58_reg/NET0131  ;
  input \G59_reg/NET0131  ;
  input \G5_pad  ;
  input \G60_reg/NET0131  ;
  input \G61_reg/NET0131  ;
  input \G62_reg/NET0131  ;
  input \G63_reg/NET0131  ;
  input \G64_reg/NET0131  ;
  input \G65_reg/NET0131  ;
  input \G66_reg/NET0131  ;
  input \G67_reg/NET0131  ;
  input \G68_reg/NET0131  ;
  input \G69_reg/NET0131  ;
  input \G6_pad  ;
  input \G70_reg/NET0131  ;
  input \G71_reg/NET0131  ;
  input \G72_reg/NET0131  ;
  input \G73_reg/NET0131  ;
  input \G74_reg/NET0131  ;
  input \G75_reg/NET0131  ;
  input \G76_reg/NET0131  ;
  input \G77_reg/NET0131  ;
  input \G78_reg/NET0131  ;
  input \G79_reg/NET0131  ;
  input \G7_pad  ;
  input \G80_reg/NET0131  ;
  input \G81_reg/NET0131  ;
  input \G82_reg/NET0131  ;
  input \G83_reg/NET0131  ;
  input \G84_reg/NET0131  ;
  input \G85_reg/NET0131  ;
  input \G86_reg/NET0131  ;
  input \G87_reg/NET0131  ;
  input \G88_reg/NET0131  ;
  input \G89_reg/NET0131  ;
  input \G8_pad  ;
  input \G90_reg/NET0131  ;
  input \G91_reg/NET0131  ;
  input \G92_reg/NET0131  ;
  input \G94_reg/NET0131  ;
  input \G9_pad  ;
  output \G701BF_pad  ;
  output \G702_pad  ;
  output \G727_pad  ;
  output \_al_n0  ;
  output \_al_n1  ;
  output \g2503/_0_  ;
  output \g2514/_0_  ;
  output \g2516/_0_  ;
  output \g2542/_0_  ;
  output \g2549/_0_  ;
  output \g2553/_0_  ;
  output \g2554/_0_  ;
  output \g2570/_0_  ;
  output \g2574/_0_  ;
  output \g2576/_0_  ;
  output \g2583/_0_  ;
  output \g2588/_0_  ;
  output \g2602/_0_  ;
  output \g2603/_0_  ;
  output \g2604/_0_  ;
  output \g2605/_0_  ;
  output \g2611/_0_  ;
  output \g2614/_0_  ;
  output \g2615/_0_  ;
  output \g2644/_0_  ;
  output \g2657/_0_  ;
  output \g2663/_0_  ;
  output \g2664/_0_  ;
  output \g2666/_0_  ;
  output \g2672/_0_  ;
  output \g2678/_0_  ;
  output \g2681/_0_  ;
  output \g2696/_00_  ;
  output \g2698/_0_  ;
  output \g2699/_0_  ;
  output \g2700/_00_  ;
  output \g2717/_0_  ;
  output \g2719/_0_  ;
  output \g2723/_0_  ;
  output \g2726/_3_  ;
  output \g2735/_0_  ;
  output \g2737/_0_  ;
  output \g2740/_0_  ;
  output \g2785/_0_  ;
  output \g2786/_0_  ;
  output \g2787/_1__syn_2  ;
  output \g2790/_1__syn_2  ;
  output \g2798/_2_  ;
  output \g2801/_0_  ;
  output \g2841/_0_  ;
  output \g2844/_0_  ;
  output \g2845/_0_  ;
  output \g2846/_0_  ;
  output \g2860/_0_  ;
  output \g2861/_0_  ;
  output \g2862/_0_  ;
  output \g2864/_0_  ;
  output \g2882/_3_  ;
  output \g2883/_3_  ;
  output \g2887/_3_  ;
  output \g2906/_0_  ;
  output \g2911/_0_  ;
  output \g3282/_0_  ;
  output \g3406/_0_  ;
  output \g3409/_0_  ;
  output \g3506/_0_  ;
  output \g3685/_3_  ;
  output \g3694/_0_  ;
  output \g3743/_0_  ;
  output \g3753/_0_  ;
  output \g3785/_0_  ;
  output \g3835/_0_  ;
  output \g3946/_2_  ;
  output \g3976/_0_  ;
  wire n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 ;
  assign n89 = ~\G4_pad  & ~\G90_reg/NET0131  ;
  assign n90 = ~\G64_reg/NET0131  & \G90_reg/NET0131  ;
  assign n91 = \G8_pad  & ~\G90_reg/NET0131  ;
  assign n92 = ~n90 & ~n91 ;
  assign n93 = ~\G84_reg/NET0131  & ~n92 ;
  assign n94 = ~\G85_reg/NET0131  & n92 ;
  assign n95 = ~n93 & ~n94 ;
  assign n96 = \G78_reg/NET0131  & \G90_reg/NET0131  ;
  assign n97 = n95 & n96 ;
  assign n98 = ~n89 & ~n97 ;
  assign n99 = ~\G46_reg/NET0131  & ~n98 ;
  assign n100 = ~\G3_pad  & ~\G90_reg/NET0131  ;
  assign n101 = \G77_reg/NET0131  & \G90_reg/NET0131  ;
  assign n102 = n95 & n101 ;
  assign n103 = ~n100 & ~n102 ;
  assign n104 = ~\G45_reg/NET0131  & ~n103 ;
  assign n105 = ~\G2_pad  & ~\G90_reg/NET0131  ;
  assign n106 = \G76_reg/NET0131  & \G90_reg/NET0131  ;
  assign n107 = n95 & n106 ;
  assign n108 = ~n105 & ~n107 ;
  assign n109 = \G44_reg/NET0131  & n108 ;
  assign n110 = \G45_reg/NET0131  & n103 ;
  assign n111 = ~n109 & ~n110 ;
  assign n112 = ~\G0_pad  & ~\G90_reg/NET0131  ;
  assign n113 = \G74_reg/NET0131  & \G90_reg/NET0131  ;
  assign n114 = n95 & n113 ;
  assign n115 = ~n112 & ~n114 ;
  assign n116 = \G42_reg/NET0131  & n115 ;
  assign n117 = ~\G1_pad  & ~\G90_reg/NET0131  ;
  assign n118 = \G75_reg/NET0131  & \G90_reg/NET0131  ;
  assign n119 = n95 & n118 ;
  assign n120 = ~n117 & ~n119 ;
  assign n121 = \G43_reg/NET0131  & n120 ;
  assign n122 = ~n116 & ~n121 ;
  assign n123 = ~\G44_reg/NET0131  & ~n108 ;
  assign n124 = ~\G43_reg/NET0131  & ~n120 ;
  assign n125 = ~n123 & ~n124 ;
  assign n126 = ~n122 & n125 ;
  assign n127 = n111 & ~n126 ;
  assign n128 = ~n104 & ~n127 ;
  assign n129 = \G46_reg/NET0131  & n98 ;
  assign n130 = ~n128 & ~n129 ;
  assign n131 = ~n99 & ~n130 ;
  assign n132 = ~\G24_reg/NET0131  & \G25_reg/NET0131  ;
  assign n133 = \G26_reg/NET0131  & ~\G27_reg/NET0131  ;
  assign n134 = n132 & n133 ;
  assign n135 = \G28_reg/NET0131  & n134 ;
  assign n136 = ~n131 & n135 ;
  assign n139 = ~\G29_reg/NET0131  & \G30_reg/NET0131  ;
  assign n138 = \G32_reg/NET0131  & \G33_reg/NET0131  ;
  assign n140 = \G31_reg/NET0131  & ~\G34_reg/NET0131  ;
  assign n141 = n138 & n140 ;
  assign n142 = n139 & n141 ;
  assign n143 = n136 & n142 ;
  assign n144 = \G92_reg/NET0131  & ~n143 ;
  assign n148 = ~\G79_reg/NET0131  & ~\G80_reg/NET0131  ;
  assign n149 = ~\G81_reg/NET0131  & ~\G82_reg/NET0131  ;
  assign n150 = n148 & n149 ;
  assign n151 = ~\G78_reg/NET0131  & ~n150 ;
  assign n152 = \G78_reg/NET0131  & n150 ;
  assign n153 = ~n151 & ~n152 ;
  assign n154 = \G77_reg/NET0131  & ~\G82_reg/NET0131  ;
  assign n155 = ~\G77_reg/NET0131  & \G82_reg/NET0131  ;
  assign n161 = ~n154 & ~n155 ;
  assign n156 = \G74_reg/NET0131  & ~\G79_reg/NET0131  ;
  assign n157 = ~\G74_reg/NET0131  & \G79_reg/NET0131  ;
  assign n162 = ~n156 & ~n157 ;
  assign n163 = n161 & n162 ;
  assign n145 = ~\G75_reg/NET0131  & ~\G80_reg/NET0131  ;
  assign n146 = \G75_reg/NET0131  & \G80_reg/NET0131  ;
  assign n147 = ~n145 & ~n146 ;
  assign n158 = ~\G76_reg/NET0131  & ~\G81_reg/NET0131  ;
  assign n159 = \G76_reg/NET0131  & \G81_reg/NET0131  ;
  assign n160 = ~n158 & ~n159 ;
  assign n164 = ~n147 & ~n160 ;
  assign n165 = n163 & n164 ;
  assign n166 = ~n153 & n165 ;
  assign n167 = \G16_pad  & ~\G66_reg/NET0131  ;
  assign n168 = ~\G83_reg/NET0131  & n167 ;
  assign n169 = n166 & n168 ;
  assign n170 = \G90_reg/NET0131  & ~n169 ;
  assign n171 = ~n144 & ~n170 ;
  assign n172 = \G58_reg/NET0131  & n171 ;
  assign n173 = \G91_reg/NET0131  & n144 ;
  assign n174 = ~\G36_reg/NET0131  & \G37_reg/NET0131  ;
  assign n175 = \G38_reg/NET0131  & n170 ;
  assign n176 = n174 & n175 ;
  assign n177 = ~\G39_reg/NET0131  & ~\G40_reg/NET0131  ;
  assign n178 = \G41_reg/NET0131  & n177 ;
  assign n179 = \G91_reg/NET0131  & ~n178 ;
  assign n180 = \G58_reg/NET0131  & ~n179 ;
  assign n181 = n176 & n180 ;
  assign n182 = ~n173 & n181 ;
  assign n183 = ~n172 & ~n182 ;
  assign n184 = \G59_reg/NET0131  & ~n183 ;
  assign n185 = \G91_reg/NET0131  & ~n184 ;
  assign n186 = \G53_reg/NET0131  & \G61_reg/NET0131  ;
  assign n187 = \G62_reg/NET0131  & n186 ;
  assign n188 = ~n185 & n187 ;
  assign n189 = \G89_reg/NET0131  & n188 ;
  assign n190 = ~n144 & n178 ;
  assign n191 = \G88_reg/NET0131  & n190 ;
  assign n192 = \G92_reg/NET0131  & ~n136 ;
  assign n193 = n142 & ~n192 ;
  assign n194 = \G87_reg/NET0131  & n193 ;
  assign n137 = ~\G94_reg/NET0131  & n136 ;
  assign n195 = ~\G90_reg/NET0131  & ~n137 ;
  assign n196 = ~n194 & n195 ;
  assign n197 = ~n191 & n196 ;
  assign n198 = ~n189 & n197 ;
  assign n199 = ~\G68_reg/NET0131  & \G72_reg/NET0131  ;
  assign n204 = \G67_reg/NET0131  & ~\G71_reg/NET0131  ;
  assign n209 = ~n199 & ~n204 ;
  assign n205 = \G69_reg/NET0131  & ~\G73_reg/NET0131  ;
  assign n206 = ~\G69_reg/NET0131  & \G73_reg/NET0131  ;
  assign n210 = ~n205 & ~n206 ;
  assign n207 = ~\G67_reg/NET0131  & \G71_reg/NET0131  ;
  assign n208 = \G68_reg/NET0131  & ~\G72_reg/NET0131  ;
  assign n211 = ~n207 & ~n208 ;
  assign n212 = n210 & n211 ;
  assign n213 = n209 & n212 ;
  assign n200 = ~\G71_reg/NET0131  & ~\G72_reg/NET0131  ;
  assign n201 = ~\G73_reg/NET0131  & n200 ;
  assign n202 = ~\G70_reg/NET0131  & n201 ;
  assign n203 = \G70_reg/NET0131  & ~n201 ;
  assign n214 = ~n202 & ~n203 ;
  assign n215 = n213 & n214 ;
  assign n216 = \G14_pad  & ~n215 ;
  assign n217 = ~\G90_reg/NET0131  & ~n216 ;
  assign n218 = ~n185 & n186 ;
  assign n219 = ~\G62_reg/NET0131  & ~n218 ;
  assign n220 = \G14_pad  & ~n188 ;
  assign n221 = ~n219 & n220 ;
  assign n223 = \G53_reg/NET0131  & ~n185 ;
  assign n224 = \G14_pad  & ~n223 ;
  assign n222 = \G51_reg/NET0131  & ~n185 ;
  assign n225 = ~\G51_reg/NET0131  & n185 ;
  assign n226 = ~n222 & ~n225 ;
  assign n227 = n224 & n226 ;
  assign n228 = ~\G52_reg/NET0131  & ~n222 ;
  assign n229 = \G52_reg/NET0131  & n222 ;
  assign n230 = n224 & ~n229 ;
  assign n231 = ~n228 & n230 ;
  assign n235 = \G91_reg/NET0131  & ~n190 ;
  assign n236 = n174 & ~n235 ;
  assign n237 = ~\G38_reg/NET0131  & n236 ;
  assign n238 = n170 & ~n237 ;
  assign n239 = n139 & ~n192 ;
  assign n240 = \G31_reg/NET0131  & n239 ;
  assign n241 = \G34_reg/NET0131  & n138 ;
  assign n242 = n240 & n241 ;
  assign n243 = \G92_reg/NET0131  & ~n170 ;
  assign n244 = ~n242 & n243 ;
  assign n245 = ~n166 & ~n244 ;
  assign n246 = ~n238 & n245 ;
  assign n248 = ~\G74_reg/NET0131  & ~n246 ;
  assign n232 = ~\G90_reg/NET0131  & \G9_pad  ;
  assign n233 = \G90_reg/NET0131  & ~n216 ;
  assign n234 = ~n232 & ~n233 ;
  assign n247 = \G74_reg/NET0131  & n246 ;
  assign n249 = n234 & ~n247 ;
  assign n250 = ~n248 & n249 ;
  assign n252 = n176 & ~n235 ;
  assign n253 = ~n171 & ~n252 ;
  assign n254 = \G57_reg/NET0131  & ~n253 ;
  assign n256 = ~\G58_reg/NET0131  & ~n254 ;
  assign n251 = \G14_pad  & n183 ;
  assign n255 = \G58_reg/NET0131  & n254 ;
  assign n257 = n251 & ~n255 ;
  assign n258 = ~n256 & n257 ;
  assign n259 = ~\G57_reg/NET0131  & n253 ;
  assign n260 = n251 & ~n254 ;
  assign n261 = ~n259 & n260 ;
  assign n262 = ~\G59_reg/NET0131  & n183 ;
  assign n263 = \G14_pad  & ~n184 ;
  assign n264 = ~n262 & n263 ;
  assign n265 = \G38_reg/NET0131  & ~n236 ;
  assign n266 = ~n237 & ~n265 ;
  assign n267 = \G14_pad  & ~n266 ;
  assign n268 = ~\G36_reg/NET0131  & ~n235 ;
  assign n269 = ~\G37_reg/NET0131  & ~n268 ;
  assign n270 = \G14_pad  & ~n236 ;
  assign n271 = ~n269 & n270 ;
  assign n272 = \G36_reg/NET0131  & n235 ;
  assign n273 = ~n268 & ~n272 ;
  assign n274 = \G14_pad  & ~n273 ;
  assign n275 = ~\G39_reg/NET0131  & ~n144 ;
  assign n276 = ~\G40_reg/NET0131  & n275 ;
  assign n277 = ~\G41_reg/NET0131  & ~n276 ;
  assign n278 = \G14_pad  & ~n190 ;
  assign n279 = ~n277 & n278 ;
  assign n280 = \G40_reg/NET0131  & ~n275 ;
  assign n281 = ~n276 & ~n280 ;
  assign n282 = \G14_pad  & ~n281 ;
  assign n283 = \G39_reg/NET0131  & ~n144 ;
  assign n284 = \G56_reg/NET0131  & n283 ;
  assign n285 = \G91_reg/NET0131  & ~n284 ;
  assign n287 = ~\G47_reg/NET0131  & n285 ;
  assign n286 = ~\G12_pad  & ~n285 ;
  assign n288 = \G14_pad  & ~n286 ;
  assign n289 = ~n287 & n288 ;
  assign n291 = ~\G49_reg/NET0131  & n285 ;
  assign n290 = ~\G48_reg/NET0131  & ~n285 ;
  assign n292 = \G14_pad  & ~n290 ;
  assign n293 = ~n291 & n292 ;
  assign n295 = ~\G48_reg/NET0131  & n285 ;
  assign n294 = ~\G47_reg/NET0131  & ~n285 ;
  assign n296 = \G14_pad  & ~n294 ;
  assign n297 = ~n295 & n296 ;
  assign n299 = ~\G50_reg/NET0131  & n285 ;
  assign n298 = ~\G49_reg/NET0131  & ~n285 ;
  assign n300 = \G14_pad  & ~n298 ;
  assign n301 = ~n299 & n300 ;
  assign n302 = \G55_reg/NET0131  & n283 ;
  assign n303 = ~\G56_reg/NET0131  & ~n302 ;
  assign n304 = \G14_pad  & ~n284 ;
  assign n305 = ~n303 & n304 ;
  assign n306 = ~\G55_reg/NET0131  & ~n283 ;
  assign n307 = ~n302 & ~n306 ;
  assign n308 = n304 & n307 ;
  assign n309 = ~\G39_reg/NET0131  & n144 ;
  assign n310 = \G14_pad  & ~n283 ;
  assign n311 = ~n309 & n310 ;
  assign n312 = \G32_reg/NET0131  & n240 ;
  assign n313 = \G33_reg/NET0131  & n312 ;
  assign n314 = \G34_reg/NET0131  & ~n313 ;
  assign n315 = ~n193 & ~n314 ;
  assign n316 = \G14_pad  & ~n315 ;
  assign n317 = ~\G33_reg/NET0131  & ~n312 ;
  assign n318 = \G14_pad  & ~n313 ;
  assign n319 = ~n317 & n318 ;
  assign n320 = ~\G29_reg/NET0131  & ~n192 ;
  assign n321 = ~\G30_reg/NET0131  & ~n320 ;
  assign n322 = \G14_pad  & ~n239 ;
  assign n323 = ~n321 & n322 ;
  assign n324 = ~\G32_reg/NET0131  & ~n240 ;
  assign n325 = \G14_pad  & ~n312 ;
  assign n326 = ~n324 & n325 ;
  assign n327 = \G29_reg/NET0131  & n192 ;
  assign n328 = ~n320 & ~n327 ;
  assign n329 = \G14_pad  & ~n328 ;
  assign n330 = ~\G31_reg/NET0131  & ~n239 ;
  assign n331 = \G14_pad  & ~n240 ;
  assign n332 = ~n330 & n331 ;
  assign n333 = ~n131 & n134 ;
  assign n334 = ~\G28_reg/NET0131  & ~n333 ;
  assign n335 = \G14_pad  & ~n136 ;
  assign n336 = ~n334 & n335 ;
  assign n337 = ~\G24_reg/NET0131  & ~n131 ;
  assign n338 = \G25_reg/NET0131  & n337 ;
  assign n339 = \G26_reg/NET0131  & n338 ;
  assign n340 = \G27_reg/NET0131  & ~n339 ;
  assign n341 = ~n333 & ~n340 ;
  assign n342 = \G14_pad  & ~n341 ;
  assign n343 = ~\G25_reg/NET0131  & ~n337 ;
  assign n344 = \G14_pad  & ~n338 ;
  assign n345 = ~n343 & n344 ;
  assign n346 = ~\G26_reg/NET0131  & ~n338 ;
  assign n347 = \G14_pad  & ~n339 ;
  assign n348 = ~n346 & n347 ;
  assign n349 = \G24_reg/NET0131  & n131 ;
  assign n350 = ~n337 & ~n349 ;
  assign n351 = \G14_pad  & ~n350 ;
  assign n352 = ~\G6_pad  & ~\G90_reg/NET0131  ;
  assign n353 = ~n170 & ~n352 ;
  assign n361 = ~\G5_pad  & ~\G90_reg/NET0131  ;
  assign n362 = ~\G83_reg/NET0131  & \G90_reg/NET0131  ;
  assign n363 = n166 & n362 ;
  assign n364 = ~n361 & ~n363 ;
  assign n366 = ~n99 & ~n104 ;
  assign n365 = ~\G42_reg/NET0131  & ~n115 ;
  assign n367 = ~n129 & ~n365 ;
  assign n368 = n366 & n367 ;
  assign n369 = n111 & n122 ;
  assign n370 = n125 & n369 ;
  assign n371 = n368 & n370 ;
  assign n372 = ~n364 & ~n371 ;
  assign n373 = ~\G35_reg/NET0131  & ~\G92_reg/NET0131  ;
  assign n374 = \G34_reg/NET0131  & \G92_reg/NET0131  ;
  assign n375 = ~n373 & ~n374 ;
  assign n376 = ~n170 & n375 ;
  assign n377 = ~n175 & ~n376 ;
  assign n378 = ~n372 & ~n377 ;
  assign n379 = ~n131 & ~n378 ;
  assign n380 = ~n353 & ~n379 ;
  assign n354 = \G59_reg/NET0131  & ~\G91_reg/NET0131  ;
  assign n355 = \G62_reg/NET0131  & \G91_reg/NET0131  ;
  assign n356 = ~n354 & ~n355 ;
  assign n357 = \G90_reg/NET0131  & ~n356 ;
  assign n358 = \G35_reg/NET0131  & ~\G90_reg/NET0131  ;
  assign n359 = ~n357 & ~n358 ;
  assign n360 = n353 & n359 ;
  assign n381 = \G14_pad  & ~n360 ;
  assign n382 = ~n380 & n381 ;
  assign n385 = ~\G15_pad  & ~\G23_reg/NET0131  ;
  assign n386 = \G15_pad  & ~\G22_reg/NET0131  ;
  assign n387 = ~n385 & ~n386 ;
  assign n388 = \G47_reg/NET0131  & \G48_reg/NET0131  ;
  assign n389 = \G49_reg/NET0131  & \G50_reg/NET0131  ;
  assign n390 = n388 & n389 ;
  assign n391 = ~n387 & n390 ;
  assign n392 = \G42_reg/NET0131  & n391 ;
  assign n393 = \G43_reg/NET0131  & n392 ;
  assign n394 = \G44_reg/NET0131  & n393 ;
  assign n395 = \G45_reg/NET0131  & n394 ;
  assign n397 = \G46_reg/NET0131  & n395 ;
  assign n383 = \G7_pad  & ~\G90_reg/NET0131  ;
  assign n384 = ~n233 & ~n383 ;
  assign n396 = ~\G46_reg/NET0131  & ~n395 ;
  assign n398 = n384 & ~n396 ;
  assign n399 = ~n397 & n398 ;
  assign n400 = ~\G63_reg/NET0131  & n377 ;
  assign n401 = \G14_pad  & ~n400 ;
  assign n402 = ~\G45_reg/NET0131  & ~n394 ;
  assign n403 = ~n395 & ~n402 ;
  assign n404 = n384 & n403 ;
  assign n405 = \G14_pad  & \G83_reg/NET0131  ;
  assign n406 = n95 & n405 ;
  assign n407 = ~n377 & n406 ;
  assign n408 = ~\G44_reg/NET0131  & ~n393 ;
  assign n409 = ~n394 & ~n408 ;
  assign n410 = n384 & n409 ;
  assign n411 = ~\G42_reg/NET0131  & ~n391 ;
  assign n412 = ~n392 & ~n411 ;
  assign n413 = n384 & n412 ;
  assign n414 = ~\G43_reg/NET0131  & ~n392 ;
  assign n415 = ~n393 & ~n414 ;
  assign n416 = n384 & n415 ;
  assign n418 = ~\G63_reg/NET0131  & n215 ;
  assign n417 = ~\G64_reg/NET0131  & ~n215 ;
  assign n419 = \G14_pad  & ~n417 ;
  assign n420 = ~n418 & n419 ;
  assign n422 = ~\G65_reg/NET0131  & n215 ;
  assign n421 = ~\G66_reg/NET0131  & ~n215 ;
  assign n423 = \G14_pad  & ~n421 ;
  assign n424 = ~n422 & n423 ;
  assign n425 = \G14_pad  & ~n233 ;
  assign n426 = \G91_reg/NET0131  & n215 ;
  assign n427 = \G14_pad  & ~n426 ;
  assign n428 = ~\G65_reg/NET0131  & ~n215 ;
  assign n429 = \G14_pad  & ~n428 ;
  assign n430 = \G13_pad  & \G14_pad  ;
  assign n431 = ~\G10_pad  & ~\G90_reg/NET0131  ;
  assign n432 = \G86_reg/NET0131  & ~n431 ;
  assign n433 = n430 & ~n432 ;
  assign n434 = ~n386 & n390 ;
  assign n435 = ~\G15_pad  & ~\G47_reg/NET0131  ;
  assign n436 = ~\G48_reg/NET0131  & ~\G49_reg/NET0131  ;
  assign n437 = ~\G50_reg/NET0131  & n436 ;
  assign n438 = n435 & n437 ;
  assign n439 = \G22_reg/NET0131  & ~n438 ;
  assign n440 = ~n434 & ~n439 ;
  assign n443 = ~\G10_pad  & ~\G92_reg/NET0131  ;
  assign n441 = \G10_pad  & ~\G91_reg/NET0131  ;
  assign n442 = \G13_pad  & ~\G86_reg/NET0131  ;
  assign n444 = ~n441 & ~n442 ;
  assign n445 = ~n443 & n444 ;
  assign n446 = n430 & ~n445 ;
  assign n448 = \G10_pad  & ~\G90_reg/NET0131  ;
  assign n447 = ~\G10_pad  & ~\G91_reg/NET0131  ;
  assign n449 = ~n442 & ~n447 ;
  assign n450 = ~n448 & n449 ;
  assign n451 = n430 & ~n450 ;
  assign n453 = \G11_pad  & \G94_reg/NET0131  ;
  assign n452 = ~\G11_pad  & ~\G87_reg/NET0131  ;
  assign n454 = \G14_pad  & ~n452 ;
  assign n455 = ~n453 & n454 ;
  assign n457 = \G11_pad  & ~\G87_reg/NET0131  ;
  assign n456 = ~\G11_pad  & ~\G88_reg/NET0131  ;
  assign n458 = \G14_pad  & ~n456 ;
  assign n459 = ~n457 & n458 ;
  assign n461 = \G11_pad  & ~\G88_reg/NET0131  ;
  assign n460 = ~\G11_pad  & ~\G89_reg/NET0131  ;
  assign n462 = \G14_pad  & ~n460 ;
  assign n463 = ~n461 & n462 ;
  assign n465 = \G11_pad  & \G89_reg/NET0131  ;
  assign n464 = ~\G11_pad  & ~\G94_reg/NET0131  ;
  assign n466 = \G14_pad  & ~n464 ;
  assign n467 = ~n465 & n466 ;
  assign n468 = \G4_pad  & \G63_reg/NET0131  ;
  assign n469 = \G1_pad  & ~\G63_reg/NET0131  ;
  assign n470 = ~n468 & ~n469 ;
  assign n471 = \G3_pad  & \G63_reg/NET0131  ;
  assign n472 = \G0_pad  & ~\G63_reg/NET0131  ;
  assign n473 = ~n471 & ~n472 ;
  assign n474 = \G5_pad  & \G63_reg/NET0131  ;
  assign n475 = \G2_pad  & ~\G63_reg/NET0131  ;
  assign n476 = ~n474 & ~n475 ;
  assign n477 = \G14_pad  & ~\G35_reg/NET0131  ;
  assign n478 = \G74_reg/NET0131  & \G75_reg/NET0131  ;
  assign n479 = n245 & n478 ;
  assign n480 = ~n238 & n479 ;
  assign n481 = \G76_reg/NET0131  & n480 ;
  assign n482 = \G77_reg/NET0131  & n481 ;
  assign n484 = \G78_reg/NET0131  & n482 ;
  assign n483 = ~\G78_reg/NET0131  & ~n482 ;
  assign n485 = n234 & ~n483 ;
  assign n486 = ~n484 & n485 ;
  assign n487 = ~\G75_reg/NET0131  & ~n247 ;
  assign n488 = n234 & ~n480 ;
  assign n489 = ~n487 & n488 ;
  assign n490 = n166 & n377 ;
  assign n491 = \G83_reg/NET0131  & ~n490 ;
  assign n492 = ~n246 & ~n491 ;
  assign n493 = n234 & ~n492 ;
  assign n494 = ~\G77_reg/NET0131  & ~n481 ;
  assign n495 = n234 & ~n482 ;
  assign n496 = ~n494 & n495 ;
  assign n497 = \G91_reg/NET0131  & ~n187 ;
  assign n498 = n184 & ~n497 ;
  assign n499 = \G90_reg/NET0131  & ~n498 ;
  assign n502 = \G67_reg/NET0131  & ~n499 ;
  assign n503 = ~\G68_reg/NET0131  & ~n502 ;
  assign n500 = \G67_reg/NET0131  & \G68_reg/NET0131  ;
  assign n501 = ~n499 & n500 ;
  assign n504 = n216 & ~n501 ;
  assign n505 = ~n503 & n504 ;
  assign n508 = ~\G60_reg/NET0131  & ~n223 ;
  assign n506 = \G60_reg/NET0131  & n223 ;
  assign n507 = \G14_pad  & ~n218 ;
  assign n509 = ~n506 & n507 ;
  assign n510 = ~n508 & n509 ;
  assign n511 = \G53_reg/NET0131  & n230 ;
  assign n512 = \G14_pad  & ~\G53_reg/NET0131  ;
  assign n513 = n229 & n512 ;
  assign n514 = ~n511 & ~n513 ;
  assign n515 = ~\G61_reg/NET0131  & ~n506 ;
  assign n516 = n507 & ~n515 ;
  assign n517 = ~\G76_reg/NET0131  & ~n480 ;
  assign n518 = n234 & ~n481 ;
  assign n519 = ~n517 & n518 ;
  assign n520 = ~\G67_reg/NET0131  & n499 ;
  assign n521 = n216 & ~n502 ;
  assign n522 = ~n520 & n521 ;
  assign n524 = \G69_reg/NET0131  & n501 ;
  assign n523 = ~\G69_reg/NET0131  & ~n501 ;
  assign n525 = n216 & ~n523 ;
  assign n526 = ~n524 & n525 ;
  assign n528 = \G70_reg/NET0131  & n524 ;
  assign n527 = ~\G70_reg/NET0131  & ~n524 ;
  assign n529 = n216 & ~n527 ;
  assign n530 = ~n528 & n529 ;
  assign \G701BF_pad  = ~\G15_pad  ;
  assign \G702_pad  = n198 ;
  assign \G727_pad  = n217 ;
  assign \_al_n0  = 1'b0 ;
  assign \_al_n1  = ~1'b0 ;
  assign \g2503/_0_  = n221 ;
  assign \g2514/_0_  = n227 ;
  assign \g2516/_0_  = n231 ;
  assign \g2542/_0_  = n250 ;
  assign \g2549/_0_  = n258 ;
  assign \g2553/_0_  = n261 ;
  assign \g2554/_0_  = n264 ;
  assign \g2570/_0_  = n267 ;
  assign \g2574/_0_  = n271 ;
  assign \g2576/_0_  = n274 ;
  assign \g2583/_0_  = n279 ;
  assign \g2588/_0_  = n282 ;
  assign \g2602/_0_  = n289 ;
  assign \g2603/_0_  = n293 ;
  assign \g2604/_0_  = n297 ;
  assign \g2605/_0_  = n301 ;
  assign \g2611/_0_  = n305 ;
  assign \g2614/_0_  = n308 ;
  assign \g2615/_0_  = n311 ;
  assign \g2644/_0_  = n316 ;
  assign \g2657/_0_  = n319 ;
  assign \g2663/_0_  = n323 ;
  assign \g2664/_0_  = n326 ;
  assign \g2666/_0_  = n329 ;
  assign \g2672/_0_  = n332 ;
  assign \g2678/_0_  = n336 ;
  assign \g2681/_0_  = n342 ;
  assign \g2696/_00_  = n345 ;
  assign \g2698/_0_  = n348 ;
  assign \g2699/_0_  = n351 ;
  assign \g2700/_00_  = n382 ;
  assign \g2717/_0_  = n399 ;
  assign \g2719/_0_  = n401 ;
  assign \g2723/_0_  = n404 ;
  assign \g2726/_3_  = n407 ;
  assign \g2735/_0_  = n410 ;
  assign \g2737/_0_  = n413 ;
  assign \g2740/_0_  = n416 ;
  assign \g2785/_0_  = n420 ;
  assign \g2786/_0_  = n424 ;
  assign \g2787/_1__syn_2  = ~n425 ;
  assign \g2790/_1__syn_2  = ~n427 ;
  assign \g2798/_2_  = n387 ;
  assign \g2801/_0_  = n429 ;
  assign \g2841/_0_  = ~n433 ;
  assign \g2844/_0_  = ~n440 ;
  assign \g2845/_0_  = ~n446 ;
  assign \g2846/_0_  = ~n451 ;
  assign \g2860/_0_  = n455 ;
  assign \g2861/_0_  = n459 ;
  assign \g2862/_0_  = n463 ;
  assign \g2864/_0_  = n467 ;
  assign \g2882/_3_  = ~n470 ;
  assign \g2883/_3_  = ~n473 ;
  assign \g2887/_3_  = ~n476 ;
  assign \g2906/_0_  = n477 ;
  assign \g2911/_0_  = n430 ;
  assign \g3282/_0_  = n486 ;
  assign \g3406/_0_  = n489 ;
  assign \g3409/_0_  = n493 ;
  assign \g3506/_0_  = n496 ;
  assign \g3685/_3_  = n505 ;
  assign \g3694/_0_  = n510 ;
  assign \g3743/_0_  = ~n514 ;
  assign \g3753/_0_  = n516 ;
  assign \g3785/_0_  = n519 ;
  assign \g3835/_0_  = n522 ;
  assign \g3946/_2_  = n526 ;
  assign \g3976/_0_  = n530 ;
endmodule
